`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502626c4f5072ee7e00c96883309c67
zc675df88ef861a52dd2f129df810467e044033b0d729925c27eaf52c821a8b7a56163f578aa4de
zb8fd5d6b9e7f667e4ab10f60feed11e9fc5ad8fa4c9c9a79248d557e12cc304f9792bb15616805
z2b129ef059be833f397c82efb8957eb2dce90ce95b4c5c997fec3ff5ee0374d38567ce60c3ad3d
zf600383ff0166c746b53ca01c91a992bb886b6ad33e641541f37dbff3d8808315c0473c6f8b91d
zba969f231eb2990a3bde7a36419db1dd158e1b287d9120f91450f17f5a796df59f0e7c9a28bda2
z0d8bd7aa2aa0a571c5e72f1c9957733aa2a0dbd0f38be779004d7c27301b7aed9f8829217783aa
zdc89f186b56d00a3a907a5c0a493eab85f332ebd9c17272010f70bdddd6b944550bd4b9285eef4
zf812537d3caf1f720e9efed5ef2e9f533525adca6ff2b4f4003d671c79ed5e76d2867cf3f97e52
z3e4f7d0a9df55808b817fe82ccc9b3f38c007e077689fdda0aee5439a783628704b88eab123667
zfe8b190721aa98ca1b48ab856a80fcf58c0cac3d441c6cbca4a8cf1442a9b4e9644cab465cab8f
zfc86274f370a2a07622ff8a4233800071596f86c9ba7276571f32a2ac93e77295a168e0825399d
z24d1969e237cbf4ad9f8ed2aef5323cef5f45751f330e57ddeac378c92c0c4df30746fe7aa0db0
zdfd29459d435c251ead37e4cd45918d0f744cf91f1886c530ec872fe3bff166b54319aa4b8b728
zc87f4b20d5e2fdc9c0ba29398b5c95c41566731e447edf32e178bb69e27c177615eb1ae9c31383
zb0b6e92c85ca9237d6ca2b1e5016faef574212f2b2092a832064dfefe265421dcd7cd2cba21821
ze2c1ec67a3dfc96ae83bd435fcf0dc93c05c5e563fe7e7c05ed3613c03ff7c3484468831642a44
zba42c7294a23245a678bd03fa382f845c22cbbdc816d0deb37e0aaacb94ec121a0a5951264cd98
z02055063f879ea50ca21d55d7e3848d1f8a55b87151aa2e44542c7d89f383192178dd967313844
z706e489f6520aae68d2ea5cf064e7c2052038ec9ef3e93c0a01033577ffdac1295305431e96c41
zd0d76371a688c1191af12ff2ec5c795747893a65207ac2b6d05a0ab4af503373a70c0844ad3331
z19d2a165cb001f15a30d5a4f3e39b8e3ef544acc378231dc0c440efa7f28626746f1632150d18a
zcf8bf53a9fba83f4ed0601d01ea5b143e1e618c01a404a77e4792f9ebb845fb5d5695c9f2c957e
zf7d6a0fa163586772d39f5fe2df0f1cbc9f7a375477bd7c4b28ad9ea08c4751caea390b3297590
z68ab4a8cbd8a802cae8d6ed038e163cfec649c19789d83ac8fa9ff111188ef013749f47fdb2335
zeb6678dc9ce858b803e6bb4a18edc8910c514ffa539cb82f22b54e0ba4c962b0a8687fe66daa39
z854e5ebc518f6e6364837510384dcb719dfc9501c618c9899c0f049f5185a8fc49700b1a041faa
z3fde7150178df0b874a8597963893d5c85efaa9167148aa508da68ec9cbc75288a5cffedaf6201
z8a02522c54eac4f9db697ca82612566299a00a763157d15a0ce7770265eecb90e296d131dad2ec
zea1a04ddb8cf022d917e992b11ac0154d37e0d7eb0af0da23457894b2771e8754acf8cbb662c89
z1d49a7073b0a1188b682c16bca620df55e76cdb4473883eeb322ba3d38432553948f1074413a24
z22a2fd1500a9be663f5ca286dea03bf91f87f55acd9d11342ee012e25519aec561750297056095
z40300cc7d05bf668194632e968e7af7e71987bd5d827aeacffffc5c343e929a36f956b17560c50
zd7119cbcb214f087aaae936fe3bed652dd0376e23be1d38ebb3e844466627c75746f0a8c5e56d1
za770e67e4835de09a7a9cab30f6f6281c6846322457d6ae17efaf2946c430fe5bd045c50854919
z0c999dbdf9661ab670a3a5fabb205c816fcca50724b7a991d636ffdc25387b52820e357ffd038d
z59804d81835a78bd5a38e55b160d83eee08aaad5293479cdaecdb5b4a3d0d4242761f9469395c5
z230f425b3d82f6b66c85555369844fd0804cc7df6ee7518dddddbade0a209d2ce931b836ffd3b1
ze944fb1edd7da3eb24a19f5cb525b083cbd29699b7aa4a75ec9def3dd91cc135076c99377478bd
zcf3a04940758add31b1a7daebff4bc9afc17bf43518b0419b83e617a8af9c8fd0a0b40351462ae
za1392465e83aca21100a5b6ba39e7c12320e89d5c0e9b4a16b886382d175421942ee245e7ce2c2
z92d7a407a33a2666a57809d02d3bb38cfffe254db835411f04ada3f5ac3ee3f2a39465517ffc2f
zc6907bf28feefd01d7418aa58e371e6f1ab6e421a029fef0bffa5363f28a644c70cde8ff36bca1
zeb770800b04c012d54921c70b4d141fe472f2368da9573f67f7ed333db245c4753f1ab41c2ff94
z1f1026a36203c14f3fe92532b787fc1d65b60dc27841e389634edbe1904475454c34a4ba284cb0
ze1f74443ab30b559d3a66bd0c46c74f6820eef76c9c288cca0b5339c798a0043d3b985a9a1eadd
z44ec2704976722435a8e9b5a27731874cd65c85ce6c769e5a8738c0063a6fae16a6f3567db538d
zbf7df8371406ae52a6e5be7619533a62b80f8d4acbb8bf7fffddf7eb8f66bad6dedb642afe85f4
z36bb8f9ea23238fb53fcfecc1499ff6f65d31a5e12269132093f41a597f22841024d71ce7ba1ba
zfc8f9fc6b1a41a3ad56dd8a2ce0a3127867bf6a6f2196313a2b5e1a6188628aa704522ac8d4fad
z93bc75807f4251c0b182cffb453139248bf12202e9f7a09a324b0a08b72594be569800e00ba1be
z0f5568ad52007f892e4d87b4102a6fc60629eb261479f9c6d4646fb6cfba204e349c6e0119c973
ze06212e808d32178b38fc3836d6fecdb8d8c40b96e6d7103344ade8fc223ddeae22f12a43729f9
z9fa466a21c3f61c7600114e9d69a29e67e6ec8af0acd4d1dc1329a1188700ab9010a6b66cf847c
z3dbd822e81eb7a37f289f5cbee3438dbcb9d04284647f7729005ef546b44c586be7dd8bb547fcd
z3d4ef20bef2e047c527d28aac129273473c3b58a0cb36c77f2b27653770150dd32ed07e5a91a9d
z90148c609c3078dc4808592814e2ab88c23b7dfe6e999b369fd0098125dfb0c1f7a1bf3de5a413
z54eec41507f7d5c8d7e0be02c2e983436243f0c1a58041e01e834c97d390b8153dcc8481969f6d
zcaabc67a3ef3adc1fd0a4cb026ce30def304467735403f9ccedc38552e5b7014a9fc5c552fe861
zcf144533596ecc70468777ea7f3ddeaca76df07e0f2a725dec8e271f1b239fc06cbec2bc98567f
z269d9b9bb797c6fa0bb90306f7e792c8f341bbab55a718d0e657376c17ef8816bde726ed9c822b
z98b8ae9e4beaf6fe406d1e0bf76a149c60283e48727e7a7e82e3642a08a8b29f0bb2ff4cd884f9
zd602ff2f155578124a72cfdeba6a48497c516ddfe456b0174058bd9796279b630aeb3939958821
z3bcfe092cec700a1c9bd9b617cc31e7509918cf1fd3c0cae011e6e94ab53a972932dd0ca2162d4
zbf296acf62ccf7b7e2720a20eed433b30a902917520ec90de7ea27aeed134c1db6f202fa225805
z2ca1fcb9651c38c6e8854adb21339577f8786b9b80132ac34d737c152157b815910f313cc4e419
z66c6eafba1ffb1234a7935f16cb8f260e7251fba248066d65ca3952e2de1886e58071beb9e2d8b
z047c540318831bba71be6c6188c4835cc52ba358b85fb79aef13d9ae2a85292756510d827bfb82
zfd7529556a0e55c26872d7b95e887ad4208c1e826ec3bfc103deab1d37748e7efc68c4122e8754
za9759b2c605e9f6783097649f7076e9555a6943070124881cf09330c4149445b2c8b9ccc972a1c
z1e9c944abf7076e531d4cb4dfbd46819bdb2d45ebfb661deab7c31adc97c70d202cf08572d97f8
z9f450c47d6fef2b2586c070e30b9ca85debbfed3748a17d0ad7c6f6346452ec46f7e143f40b8f5
zf8785ada7864c36138fe14fb11caab2742497bf097aed5d4deb2524bc3fa2ce16c532a17027080
z0b6cca22ae9d0dabecd6813eda9e898e5b8ba479203aa8faba0a7e5738284273f54cc9c4e95034
z16ed24984f06a32701611e87c136d8958bf6e2e5b68aaf97969ca19014c38538d7d8ff5830f357
z2f95f181ade34fdaeac8d2fadf9b576954a4c9d66f5d6f3c000364adc1ecaf56721140a87af4c1
zdd390c3b7d4d8edeec9a4cba08aae5285552f18ced9b7e8c3f31fd50d222067ac94e3a77c59e9e
z224a866b4e6bd542412df6e399959487dd30fa15530ade0faa3cb117be9f4fd84a42f84799ad36
zbf863e0cc1176c4e47dcacdf88b6be3f36ae9c7d7fd1496996c1779b2bd0fe736be6039c270b13
zb6e6ac9a9ca25cd1f3a3add3bcdca052cd6c399025717256c2c4cf063f7d37d768ee656340d8dc
z8cea03b03f54ea94e538dc44afee13e0611e50f0c1af869997f80a5d554f687f674a2f33c93d92
z3d9ea099b1ae0132373b812ec099149db88da9363b41a74114565f9ba33c1764a008e1cf3252fb
ze04275fba7e0a370ec7d4c7c2281ce8748783a99e99670e0ab3bd3daa7f680b70851a6e057f6fb
zab395e109fbfe561ada9c071d4b13e07c53a296af6df94ffa5513c9a932f57a1508058b2418dcf
z04edc337bf94ac05e972025630cf71f6089dd11d2315dae1a29d670ff9d5ad5fac0a23d013df60
z02a8199d7ae1283825b031da40c14451150e8e5166195c7f5d798f8dc97ede52c3cd9c615e20f3
z9c97a04ef431d9eba235dcfc67f80411e7a290ddf8dadae436be4313b49c7726b28b5dcd4f2be4
z79b0310c1caaa09d63fd9af6997c9276c3f9db338d56ce4c4321a771324abc523987525008d33f
z0abc62cd9942967d7c467eb3c10827786c0ff9c082952cc6ca93e0430e2fa4870a6003f505428b
zcf63250239d2f668ff30dd7199f6eae53be98ce5dd7ebb904a007782c38642e6992cc32a7aee4f
z19209b9972189f746bf221d34eb752a01f0a034fcc085d88765e46051d07742d1737df83b83c76
z73de9fd4228750c7b8ee2a4942b2131578ee86b864921f8fb03de252b822662592b9ab03602345
za1f0a85ed173ad0d2b5e97503dd8aa7a26f48ca8bca0410d40d79083e59c98604a1612a083d42e
z68d3f88e904816df88533b6f6394ff5b018f613a6490533f3c7fef30710ce0437b33cf72021495
z3de9282f5218e2c7ddd49f7e10612c047be4a6d502383fdc08fb00878ee6bbf3c0f526a4a8c33a
z8c23796165e6790a2ef3aaba1bdbf6646fa762b14892150d97f63959530421dc463567e16ec5fd
za9c683261ed883f4636f15e2abfabd734d7635dfa201c283fa8197eddff621d17e2c5c1a777a96
z32a84c6ed58de165befd54bf73b0097536eabafe8b3fbb7520fea6e89782af35fa51dbe83e33bd
z853f83e0df8b8daf6a3b63be406189471ea536bf503d23d6cdc00939f0bef09e25dce862ada093
za490288d11d408df8fb89d02e55061ad555f9d5eb46da26f397dc0dec1463c9f4ad1e95f4ee416
z4c808dcdce0e823685cce1cf1058053613e3138f8788834733b4fa65a67d929e4d5742821c155b
z1b081eaf8cfb70d39c37f5f71993f625182b58ec7283ea98a28227f724d2739d195dbd723263e7
z31b5a18439f9fdf04864bd92ad021cd0b43ec471f4786f5e9aa56fcc72a4a4c511f1a82c35bd8a
z52bde387dff717455a519950cc7e10592550c75744a81a05e549e839033c071f60a6bea8da1183
z711c422e7fb6da038a44d6454e184e6377ba76d0c4e5115d6e28524f903edac97126f1ce592df2
z3fca90c195cd29ad66a5c1b4e0aa32fea062965a1dc97065da012e95f4e62d9bcaf6501cee7934
zaa60124abcfde0f92590947156b5dd99804a229c5a8368262f5fe1f0027f253a4e438225e67385
zf0da53579997e37afaa24babe6d9371a6696a3aab6729262c5da08b5c7aedff5a4bc32d8d5e6f7
z08b1126067dce106abc6ab0264bd39803feb6bbe13ee8a32169ef7ab18c864d0990a8d011650d5
zac392fa48a17afb5e0d46a750292b0f90c052f4be3fd3be84af21c94a4556a829b341626ff320a
zacb11ad7d4293fc5e969796c448b5ce6f3e9323ed31e7698cf62248ca53da3d6624c434a583afd
z62f943a37a788ae5ad542e4ebce36adfa43bca22b8972ef41a4b60c6a6c3788930f7b5bb28ebe2
z2ce1ea43951b5666a71d95b748cca31d31152d3d297d25c1daef4752a51b2303d6d453489f2f4d
z2d8ed67ce4f1a82d5279dd16822906f6e371d28625afeca4935f988bb79091bbb4a41318392491
z84c8b766c436fab5e58862dc388c3e650f6a049756478d944b77431a6fc5ec4fc9c40bd1b8f33d
z3a120ba821f7e35d3277017f3c4b34fd7d9061cf5654c84c14f9ab3aaaa2c234df7d9b09e9273f
zdf7f07648d7e6206f4c3fcb1d0d5bb2837260bf438fa5a8a256636bbd22d4e02bd0f89d26ffd91
z7e4f4e635012f196c3877e67eb2d78366df1c1c0bfde97d97e3ef5f28b6f5e789121f29e5489ff
z8c07779d6bcc2a75c7a0a2e239dd3808528987749a7c9b396f2508137ef6c5d8e0aa4ded719c39
z9be933865ffac5953d02beda2b2a26d7442fd4e742bbc7e900fc759ae4435a32f7894321b75faa
zd75ac6d40807c01a7059cbae4d22bbccd73b303c06210a6a9c17de300ce1739556f3e17267611b
zafd6b10c4729e0745f6af47b4e2f31fed4e6b4eae298632b3385a8ce1c9f3e48b64955a17475ed
zfb0e1f670bace602c4ad1931710991ada16b4be5d99ac3d4be97167e51abc31c672f2017e3e630
za51532e288f12e78d7907800b4f02d3e80e3ea136f502390fb0da0c640b4d5e24856fa71963c3d
z9ac92e3fc69a18f65ec82126a831d8acac6ebf522b3f13f63f8201aced7fba4cae9926410c63d4
z821cd47bc61f6683c8ed6c579ce46512a994c59a2b08ce5f202640ddbedaf0817a7e1bcaae2f43
z1c83b1ff8786c442be9e53d5fdbc13d60bb5e19676da4897c7f92d97166ae09184f868c49ec0b7
z003b72253a7ecf63b50eb7b7b00deee93f4f64d692be18318f8d26564fa617f04f9875a9a10271
z21649ebb7974843f9fc769936ab7a15764d0b95839d76ff51af6fca9a646a2345d4de69192067a
z78c3b28f3827022c69bfecf9771f3702c11d099552138dcc258f97dfd14ca3a9fa8d9a7d958ac3
z0ef0ff84327e32cee520bc162d3425ed8054ff0a030a658355537159f9c427a18ee5de95892e50
z69f8513460711663e1d99b988c783368b075c5af95de9a0bb571c038d193c919a2cf8db984ff5f
z0b4ab7761946c5283684f178f249a582a42c28a43b3a664c048a784f553c394a1c1ebfdcbd56f4
z6109a88e69677511604f793110e3e5d50dcc0ecbff7a8ebad3f6f911955302fec5449f92c20c18
z6ff80ebb0b774d87149626c6ac39221632be67b90cab33cea565e7d9da6915e4b356a8ef23bb49
z2db4c8a5ab7f54d0d09688cfcc0be17b4924742afa9681c7dc0ed75b9e23f1e1cbde2323d2e581
zdf88a4fe95d9d3985111055fd042689390ec21e8f33797fbd9f8af7bfd27035f21d0b0b3f3903b
zf4b308dc00eee0fc7fcbc5626243d7c1c738a17a2230f328914fe412a04c550de45c7b4fb9ac95
zde7b793d5dea6da5c5e6ca4b4560bca26d8c5f3397b00be995e941a9118b8bb8823cfb51d4374d
zd53f70cf8a8eb02a863b4d7e99508f817a0a7ae75b2528a1fcad133e9cf02eac8eaa74db1fb513
z18e7a4b0b2ced0640d4d91f109a20808a5b728404a776cb73e2d603ae376284bb3555d08ef4be7
z4f37ebb1d5a6f138abe76ad40569e7128ae84e0fc7f8385bc7fc269b1c1127046ad4c673f34f9e
za3625c882da7dc324c8a566e43961a91041938bf140a805387791514695c0b6dcac7bfdbdea297
z696a0b078f47540647b43b828802d29fbb1335d896cd5b425baeb686e87383164c8d1ac5e25d74
za190fdc569435c32204270eece623095cf46b9233ef022adac975842b9d3c835d10de71c364199
z2431bf6f58e34ac03a129d11925359aa8aa2a60a2f4035c911eecaf3c6373df724a9096b16db49
zcdf8ff6632a9fff013b4a18a88bc65c6be124698dc2fec9a11c9b94c9ed485dada02be54727a32
z050b42e2f97bd596bf0c06da0a80a1a1581aee5b2f601a54bf9590b11c8e2f9bba068cabfb6a96
z7d3e40af2cd70f7a5a863b1c786fb3a8110ba36165ed0c3fd73a5d7ac5a9f9089b27d5c45e3ef4
z6cfe4a1e40e2204f770d15597bae0fc41d4866235441788130c0073821baab765891d70f6f9e74
zb00b02ef495e06f2eee31d7a4948dcd2ef22181d31aa96343fdb78fee2b6b158ad6253c72f1cec
z881dabb54ea30e60a2f23c631c2aea8d9a0aebcdd4ea131ac91c64c84b84a337d34faf0a966627
zb6743d5f42622791b00ef4a5daffa5fa2490a88249bb7c752524e04ea975356e9044bc9ea3e1e8
zb6c70d8e38e156d5ec6edc0da2d18c7e610369eb57aebd65acc7aec3bd59d3f3e07dcf9ae293dd
zc00092c9e0a646c60a5063ac4dc57bdf7bccd946d794a43098b4c263798bdaf65e348ddde432bd
z17626a2e31d93a8ded68b3ee0c4f5b8cf03c484ae167535907729606144ad4f2b3226e3ef25052
z903b87d1725071f718092f48bbad5737e1556ed73c6f0b2349c597b40f6650ad6659bf05419534
z83933190fc22f74c66e2e530ab296f1a4be111429b6d27401cda4e18ebc687288c3438a51ae9a7
z68c44f00164ec566b101afa417d655de3a87284f3ca149cbcf55a0fe95f7376c5a449cceab8ba7
zd747e52c2e6f1e02d2ff401f802c084e20029cfa78e81c9e784bdedfdecd3804953e89f7e1d70c
z569bc33f494ef403a1c4af21efcadd95dd9f1ae2cc86edf92306f6b0b79ea3add31d9adb02a802
z452136e22cb8b44ce1cf261830739b19d6063494ae475f5e5405690cc35ac0e3f1e3f6f621fca8
z48f0e4f4b02cd40f1a9ee8f04b6905bceaec727f170d0fb61d5ab703afa977182db75de669f7e1
z5c912e75670bce3d3e82ef56a8af114738c881321a0d36ac5cf2afcbe54e734ed77ef1b8b698fd
z0f2df7c641c1d635d07dad95391314350e3cba63a2c7ea1b5204331060dca50326a07e0e72f637
z92fd73ba5fa593d88717b3eae79c49a8a4a6f20e017de0563f5fc20ac2af2aac5ded95c0dab9ff
z8ac4a275d73c672b06969bd222033453dadc63dcc4d3a4c42ef7e77e2ceff51191cdb3ef59225e
z51c1d9df85bde63f1a890f41ec18b78b7d11c16a8da4cdc57e6715d7801cc6fcfa842fa40c9b9a
z345f5960d13d543fb785b2e57d6444184f50e857ddd6160e2b7774b49805382ead3f21889a1692
z4fd67a2f6d47031f2c17c1ee7bcacde6e8108566c5d0242c4cc1a0c9984f7ac8cb5c98c6281100
z57e37d249ec0a9d3d4ba3c9ed4178c66f033b0ade2df101379ff7eee6f6caff98a5a10b4c3f93f
zc6ce1721fe0cc0435e707007aa688e6c29700b7755d5d4ad426fa585056ea82b3eafb1c3d1b963
z6903cf562dcec9b666d363213b7f67a7e0c526b8afe196570e252edddfc5f652fd2cea668e6cb7
ze4cc69152bcabdb8d52a1e4d9a090c8ba37b5b7f63ca65a1e272623282788528ffae2aa3fca7ff
zc00615b6f172e6fe69efd41b9c412a25cba289e1035c5f4caa2a759c244e673830769cfd0ff1b7
zde4014c52b349b3a89ce478a1a4738a8daad23928d14ad2d3ba4aa2e45b865c5e4054e94d0e501
z5b1bb3eb16f97b28b334c2de423ab4353dbb7db055465aa599edcc59a582777f0677065231b5bb
zfaef0fa4c615c85ba4555e17c3bb75175da745e7ef9b8d0df508d2833cd731e1d5dc067096aa8f
z81f48c2e5752457c28f173aa7e895c9ae359b74116345cb9cffd08c2806899b9cf575ff8ad251d
za7ceb0d4cdefb6ff7a911a9df3167cc7f05d601169cb0c7c4882b10354d9bef01e82a411cf2967
z310ca8dccad861ca5d6c863ab79f42d18179e5b5bae2d0c08286ca6706eff39d6564fafd97a92d
zd8df4b25c00cd6a3ca04781802b67db1ecd65c5db962ccf60aabf068e95daf2cdcc75f5ceeaada
z879b440799295f02e85a8424b0ac7cc1c3650d4bab0850945314f66cd58359f2087ca3647ffde6
zae82b3dc4d3d402fc91d0471fdc273dc39b286f04f3bf04d70a54553d49a465e65f953a1981515
zc382f5a10ee2f19c5466d8ae69ce3fa67fa8ee4c1c4443df08d23eb66e5742fbb4a74831155497
zb283b9ed50c6e13f8b385e9a35752b99c2da1b33909d108d0be03dc2687e67e4c9c0b61866e7bb
zff7f6a6bd065fda49b247a18ea70614fd6c3249c6d4f8ea6aa04cdfad22a9bea7941a5413610aa
zc4713b39d5da71d642e7c6496aea6dc4d397a0d1da48896ec13cc7a50381c2975695a28011a145
z352d2d7b3024ca6e7b1a6657acf3becb60759ae332f4b0f689b8b2f36a41b19354fe2a3d65c195
z950602aa986db74b711c70836684e9f41e99743c9e5fee421d9ecdb19fc457fc6e64c1666cf18c
z3eb4b18f905c75e34ee9b41d927175bbb33ee98e4245236e10f86040269fb97e1c4176d1b714e1
zd27d993beff485d68e24985d40d18984a8ec8534bd2b7636a30285b561d518ed284231ad94eebd
za6964b8cb36f18b3f21d8be19575122467a3243a73d01f125257292f5b7655f42044f21188aee4
z547c1f3e8bef48588212a8e4f42fc66cbb1ae3bf0f54ee7a6352bf6c2f89801cdeff6e55ff4c80
zdc657ad948fea5a49dfbabe2525c741581fa1ce23350698cb7ec1d91daecc213d702a970b89b02
z88350763310d66832523cc6602ebcd3bcf2ef39d10195dcdb40fb65966b0d12dd3e7dca055c13a
z4f1f53bccfbfa9a52446f62d5f6f5a03238e68ec68abc5008db05d928d0a3524903e6ad77ffb7e
z6a606320e5f8939bae8a539670e0c2b7ab69bc373479973975bbaf6595ab7882bfe80ff091f920
z00e17f4ea4042123ce6cfc669c6da3809540d0628f9bc0fb55d4cf818ad240ceb6ba82da0ee5e9
zc68342e12d77b5531f436848b609d457fc8eb3efb0b0773f42232b60011988cbbc095531b1530f
zbd4bb2fb66210596ad33f73db94e80b53b8589f60b052d5197aae9747e68a66c927bd9f2d12ea7
z3e972529efce09dda3fab259580a86b414a37b01f9fb105f11ff87e47a98b3af3b0d9bec45c6cb
z5e9c91cac138215a316255debebcbdb910733c6800440b6cede3868c76d82e516b9f43e2c266f8
z94397a5b3f2b0f0f5d8713cb223eee6f7e994bc8da4351a2e9fe1c9ff2dd70e4d76ad9d38b7e39
zdbdd7129759635c24badb682693178a6357dc87ca06e131c4adc9bb29e7ae0d35a154c08f5fec9
zb6689735d520612051eae9ccc7531a7ff82ff5c7ed0edde2368ef26e5b6a2a66bab116a14936e6
z2d48ee7db6339b74c0ba3c59451fc936f7c026e951d4d8902793037ad004ce67f61aa252436655
zb12183ddc3681885f3f7713d90d109e8e974be5a1b6c20486e7e619111bffa25bcf9a0badd48d0
zf2c551c420a819ed293680f602478fd6e082883761d35f793b8457b9748ec3ee864752216a82c0
zede347e8cf0221181bd1dcfb39d08a82a442658ea85a326ceb1e66f11d7a2fc86612fba598211b
z822cae04e413a8412e845e527a304952781e338e9b852a44e4ec4f910f813850ab6e4d500e15a2
ze77b718de10aaecf85f853e84a9c2d04a0c75f6acbc0aea7d18ae1e956d4fa6425ad742be870ee
z9cac510281ad7444da3b4e428b473c5d696b3f0b5ba8e4b9dc361b93894e8a672605642b305d8f
zd05305dd63f8019893a6709eebcb669ed11c32840de623995228c7a033cbe50713bf125848228b
zb3a6337f7a723c0143d0d6dab8a17c400a11ed2bf43910ed27d97f529dfa1282b19c9e31165daa
z9e2b69472f29bbb08e9a07e3f923385a5175ec88b4d10dcd03e4c8fd258b0c0956887c0023f70c
za64af655ed63202ffbdebce8016da7fc7052f7931179f099c1ca7be9174bd067a0c6a23e12e179
z27c3e02cc2db159c57a91381cfbfdffb7dc1a8d99533ae5fe86782a2a2e6cf4749596b3b157d6d
za39b82fd1f87614414de1b6e91d77d4e216840046c728b3aa71d8166fc721cbe5cf79905940eb1
z3d1cb4b462c1f1e480ada9634d2d48afd7561727e19d0efc5ba518fe77299c5a413d9298be4d0f
z74977164f7c5ca2fe2238bf33946b699f2f1caec31476dd0aa1e7a6a3c51086836dcd25dd1589b
z22ac186eb474cc43ec624b1e69782da49d181fdd70248829f991dd2ac23b6a757ab80a80f3d832
z3fcfa0ac83d5715f47e2f7ffa23ed620e951c79bb5facef3cdfb594b3f0a172617831f5547ec2f
z386b2543cb361d3cfd15657f3881e39dda1d1f77d678e30f205c3b3f4862d1256f13bccf848596
z9017269e7cf5af60fa10f5aed6a43f3ce9ec09bf94ce0ccb3ac483185fc0418c2bd57233f12cb7
z313a63885e745d668291b55531041c6a233f88781abc7c2de03e359e85f2e4c39f70f417db441d
z14ffe280e227f29f4baefd4bfbc303b3e873b87faca75e9ab767faf75158a067674dabe3cdf090
zf21c023df238278d63414dc9736bd9dbe17eaa1127667b58ad5911eae30d437696862d74539d71
z382dc2555dc172a3d853c05d164fd451689d28c43f98ed92805fa29ae6c4dd97b1f7de0e19ac76
zf06c0d7a1c218dfad56400a24d7f0e5e1be9f6181004fc2cb8be9b6d0ca352abbccda5c1b66775
z538c85c7e5c0221c69dffcbfea17a127f28383ba58c5b02ac27979dfa721e9132465337a604269
z5c627c0ffa6c80394d4e9bf5c396ab7d131b014189ca6e0e0b4bd4cc0b2a2f051181e7953016fd
zf6a58f8d0bdc17442b16d61c43c0c9d101acb213b97f8df5c969713c909a7d9ab7badd407b5c1b
zff8e9e286c617613fa2d203e298ab10d84d6666a13e1d4aa1a221953e6b30e2d849e4abba34bee
z670fd6ea1dfa082108b0332df6700d16ae4824d873a63c3943eaac151d6c562976200107a4067b
z27c72766ccde3827fc2eaafe7b7f936a0c0073b2fe695b86c405fd6cf58612950e5c42391002ad
zd42ef440fddd93d9697ac23184eea48dd8ccd472d76aacbcc6d3a7b92b9e63dbc406fcdafbd035
zb9290a08273259332b1e84ee14275ddecc77e74439b2e37b55c381ede9a62b19f29f4ff3b80f4b
z6aee5e40cf2677d66355b31f55c0f7ca8141bdb144367ef0474b1e0d3932b65bf3b077ef683182
z115cd3049b2f16df5885c1b62ebbaba474996c5e8a6a12e49ea84038d6509deb7a8b1aea07c4c2
zdd54b03e4195538d5703e731aaa9bb951e39a55c1350a969f09e7ebce13aa1fb7913b41edcca00
zb8367535d4b2049c5f3c8549b5fb50c52bea2867c7079010dcede72830aa53a968289ff520d1fd
z68ca6b64254e56e6642b902a3058abcb960b9a3e9e345c2c2b6a27e224ab3bfcef6f9a1647e9ff
zb2dbd707e6915e7a74a7382b1874d3b7c06c53d778dabb1f9292ee3c815970e7ab0fff94d040d1
zb9d7f819b0b0a20a60238486bc4612a7e4bb3aa9805954a4a4f6a43351cc9ff7fc8513cf720026
z00bddb2d21991dab881cf938c03651bbbecdbe5f9b7b7f8eb5982f1fea82bc9888378e675e317b
zdad46757db97ca5f3bea4a8b9caecfac62445e9dd409f2e596c8a7ca14a133f195eb22f6d9140f
z1fe7d3602aa3afe54c8a7a5ac32affaa7d60c970b275487e2be5552664947fa61c1aea2fd5bc77
zbbb74eee8b4c5e6e61751e05a9ff309d9fbb8a4a3a5e19c858b8a181674c2a51e51ba83c35b2b2
zd3e60c46ea72652e14b04298619e9b835d256ee9927f3d8ada62223ade337c23eb394c5634243c
zef726863f1ffc7fc34fe23fd5be6010a65b83f9444390d91fa63dca897541de7eb14eac312ac5c
z1ac1f017abcd63b473a0d40064
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_apb_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
