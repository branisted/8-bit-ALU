`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab30857016fc53a
za25afc8341302f0c829d94450c399b8ff9b0386c187cb854ee330605b7b59da379b1f26f488e1d
z36e675f0b1336408b3a1ad87d0723054f952fbefc8d5a33eaca6ef5be8f42bc59870a29a5cc9dd
z4fec09ce6e44cac279651402e7e1f590df88ce49ec26ab39f12b4a02855703c6f03b1e85c797d7
za357087d98e5b1f45502e45892e5823d6fa4b762932009620038c05d74efcea7c3fdb38901d620
z36515d0824367e48d1bc182335f158c262d396cada6b0ad58add4f945eee634c2dceadbfb5118e
z14969c29a743830a07124bfa78707f3952b96b0db7af7c9ff36f77137d8c490c4f79328328069e
zd7d5280e4f95742c9841340368b9764f0f80413adb175ecfbdf3c40716abca7b8cef6f7fe92ab9
z6bd2453f1aef7f7899c5365c5c83793cacc7795c269413f6cf0dabad14d40e9285afde8c01a47e
zb61893788ec5060288cabde8fb553f21b02eac61ab0b48ad3d54f4d1d76508b22f0c600861b5ce
zcb30ba708be817b1f50f59c0f6fce449203e7355c1be55b662fef3f92ba58243d81537761af8d6
ze27d7864d2dae99372b2b75bacdc0437a4f7e011d68c3487a89759e3625548fcc920ad06471ee7
z2d701aabf726859343208b0a543c73eeff8406febf277e3babff437ec820fb49d6b78e73bc2353
z884917487d35a6cd06d7d73ccff5f05355122888b886d178a03d8eac5505df521c14d1e332b234
z86bc1de9891c0fe4654d9d65be6ba17e0f35eaa0e5fb8d4ffce747c7530d86192c5a60f63648d8
zec2b11ca4783a37281db3c8b2556885556aafa013f24449e0a06d5242cb51399b3e756b814a7f7
z7d2f3363d024adf895ee1f4c57fb3048cf14f737f4f7878d0d0c6b48a3aeecf0d16f61ec999e70
z8673047544b470019ece6d4e6f8a1469b42dc3022d4e7bf3ec62c2af4cfb08f5a5de608628cf8d
zd4665dcc3f4867d0a07a836531edfba94cdad9d90730ba8b6b2364b0eba1514c0246e78124c617
zf6a26bec02cd6601f40650424a431a340361b2120bfaaaee24cdba68de41a962bafca77ee84e80
za2da1ab25b494bec121443cfa771b7300360491417b42658f3967a20c16d3ac0978600bf5db91e
ze42f8327318524a1e54cc36e7ad8520c8c816f80b84c9f11b4be3894c99f3417e8266c7b37bd81
z2a58aa43a5270339ede7ac0dae624098412b66014ede9389544c6ee494d95ca24a6eddd5fafeb4
z4642068486f3401b6f5c6ac8709c356a046f328195de85c670a0e8d001bdc1491121cd886b733e
z28526543476e337e144daa4a1dbf26401f3e63488cee9ef8aa6872cbab5f394266eb372e1142a4
za17efde8f6d1ae853c8f6da33e3fe266c449d71dfa287e5541c7cbb3e701429e2170f3527acc83
z3eb481eb74a0f813899db8f2298c73ce5a01bee7f76a3b683ee69ea44786e2d53be7e4b73f4ccc
z658d4b2098ad050da2060ada973781798fdfb86e1f1fae5fade012756426deb407e6f910ada1f0
z2b9aeb6648c21f52cee2c85b5a73d793e6d737b55e6850695c76068f4fea945523d25f8969fd77
z809d98bb904a313f4feb676f6a7e870e3051fa5e3c6c008ec9a4ec9564ae9607e7ab863f0e2605
z29c3c861f21224b22bb4f337632d4ea4edb29bcab88a96d6fd1523841194350bde2ab7f0503656
z5ffea9b9d88bba0e7b2b014695015230503bc0e3c2a34c4419cb4878e0c1fae075efeecd58f9f6
zb3a9ac3d61201cbe60892fed26dc82a3749e147a537d0d68fe23f6d27a7423273a54d4635a1c9b
z3c56eb66cd1b79f217aab9419354ead9587bfa10e242a4154302731784b76fa9ea4de69c8cf525
z2f9fda6198c0a3111157327b9d8e4d4d87fc17bf63df440d208e017619807910318bc35f1937c0
z0e328efd7770799d84693edf5847e2eea20b0fabbbb9339016692bad574dc3f8c8f44d4597470e
z2cbaad500cdc82c2d67d871e04e28bfc30a08e6b1756c6b8900d80ec134e402bcab9514d5ef9f2
z350a4ea16ee76b194e26f138699bc6ff4a444ac4df1dda6f5b3c2c9f0e24f780cc796731a0e955
zed760e90c2cc5de57c6648262ab7cebcb8183c40978dd1ed55cfa4b3980c61ff9c0f90a4d77f69
z24633acdeabc6fcd71f8c22dc2f0702e531046d3e3bae66b70c4a35919528c1655a221fb21a67c
zdefb8b8a0cbfaae98da730219cb0e9ab675a7829cd7f844c48bcb4520637a575f52a1890f68c02
z03c017eb40b749b3c3828a3d67d77e6b2085ce1b6a11095923480b080590a7ad27ad03fbaa86a3
z77844aa29bcced92a7ab9d7743d8cb86f1fbb595de9b641546717eefee680334bab38df3e5e6f8
zf24e8f592a3668d6284455e6bdb0bebcd2e169a3ea397c4945cb94c0dcd894a6a1644f164fd19d
zcd0d2030b79262eb78e241a95de02841de08ac3939d49f93fbc73f56545a16393fe1fe4d8eec05
z4464a254deca398bc9c1092de9902a835e50841677c758609691156544faf344493ff1dfc8249a
z619864134bf934acf4fd85e0f70abffbeb8f1d57e534bed96cafe2cc819adedbdd70231bc89015
zca7167c0899ccbf376e40de5875dcadc41a308244841f048c0ab9f50c100c99b9bc1d7163c4ca3
ze8ef991ee786038f73eca3981fefc238299e2f93f68891c6295c173e41b2e20f7d823750d48e92
zdb3f19b8b6f0a4f7e9d97ec8b0b2ac19ae7671a5a82267d2bfe546db9ab26e2bb43feb1a030170
z4b125985f5b29c1e0eeafc543627685519d404998198f88cd271521960b10b672410bbc5909834
z84e09ae1a8d720a4703210d633b5f1fe87deda93d4e85a0a8001014ec80fe62df1ea9ff7921185
z16ab1d22b3a131c313763953de433361290b4a3ba4dc472930ed3aa94c2a3fedd2d92931caa472
z4c138c522553baba50ced771767f1d25c9739f28293ecb612be5a31179ae7f7b9aae060e3b1f45
z5f2c1821328c373b92dd5b9e7a5e4042ea433d509d1d0ac4ac400e46fca021b4cc9e54029c1fff
zed9718341c220c1b5adfb9943780521ec517ec8c8c24b87c4fdd4c4e87b04da6e0562664770ee5
zbfa56836825ecc532280b9ac736002aa0ce62697f16dcc023184b29b4c95dfe97bceb79d3d5fce
z8432a208282922194eec55866118c937c63293cbbeae0a01530123ecf36a1dae3c5cb4d7c306c8
z61fcdddb763d6ca97f9db42936da55c2c730dc286136538c752b41b84f47ba92908c1350b86524
z4855d45e6fcb37e8799d093a35eae7d377e41e244f600c95645ce5c3e4f45cfc0e05cdf216a7d4
zb78011cddd86fc49a17d7917e8279c64aa86a4f0fd42c35065cd185e21586eeb73b4209d4aa613
ze585b65c1834e895beca4fbee6142676685e61f099e0a40ce243a945bf972d50e060358e18aa47
z2e394dec7176eb130413fa36448fd186696ada2b02d164c206479c816ab581567269176f12e40b
z739b9bb926aa1d6c93b0ee5c541627b2bb4859e1a9c356539c481ecad7c3f44d76d27caff143fd
z9ae09ad7342137aad851f8d186de59e7030abc373865f1c2d67304b85c1b4fe8c10eba1420ce00
zf660a226dc17c7d51041b072c2c45b5b18b4d68c5873d405bf5a0cbf0886eb7076d7997ea61c8e
ze023aeb281afd62e77341d18d865afaa1ac06b933ba5f12e4ed63cbfb079c38282a768ac8a3ba8
z0dec848adfb567dab9a7857abb6bce2339f8d6efa5acbc924fb9bafc0dc87340dd8df60633b93e
z61798f022c08ad125f2b0c12e36fff400159b0cff3de0c702893a13526402ccac99916d099ec61
z4590f5ea89f2b7e443119f0f863ad821d75cd870dc26e9795cbdb3e7ce2f563a6af2ff2b075b3b
za4663858ea6963a274ba62296b8af54e91e85844d898e70ae71c27525a89b58e388aac72bc9280
zf17286546c1c88b41c9cd04951c19065bb352b1f64c50678a63c3cccdad4dc425b70fa22846939
z1aef64f74eb7746555368ff56b30a5c74dc82466be332140f72400aa1bd605c2850380ca6c268e
z0b13ebdff755e5b127ffac793b7a3e46ef987e9441d4a838bcaee01070a5b787f74a8ec54fc86e
z5015828576ee86e59af8f519b90e537f9b102adf99f78fa590ba806e62dcf68106126bc6e7158b
z03862529e1b1dc8d74255bbcf8b01d52991611b13fd0e01d53621a6020313b80c59154f7fcc577
z0fd892975b71aa416c05855a49db95f82e598a1511a4cbce5e6201ad834055c6abe1b3f4f8d98c
ze6fba4115150c375c7a9e1274a9af12e8e4711df8d349087be598ee6ba93c2ece9a39ffb4df45e
z12b992a707b16f9b53485d07afe31996eecffd990463a1ba61abf02d322fdb6f621b95694e0563
zed0e9194e682ae5848b9a15e6f720561e2561c80eb27551b7d72ebc12b3a06500d7058b61eb879
z9ccb7d5f36ce42f16bc99b008e59424142af92a7ccd47e13b71db6c8f7e6a3474c6d88bc6d5a1f
z3cb0a6a8c5d6f5c159e50f920c3daa13e64ec34edfb512aa6a39f70bb763e854fd82671307b81e
z173d209c70644949420b6c58b3597b2147bd2f5ad31d0d21af5b86915577f37209261132625217
zb0f2e68392241c7a90e8156a9f28d06a6a26a67979f36272b2995bd8965de91494a3048633fbf7
z7b364a6d8af61f396d7960926252ed2dd05532fd22e6f93a35854032981060304762cdb3af0778
zc2878435e0f5b364560784316af3f338689d942c0d51c81b3d7e89bdd9541e5650a9a551eb188a
z36209029c1208fb0c864d9f20b6835b041a2d334306d75c02bed60d1082bc624d5d899a8609437
z5841e56c8825dfcf41c57789dcb717273ce45ddac850f6a69af6e0f23076a14ef0f38de9ba5b21
zfaa176b2397e543b6b01561cefeafa952fd7497e958a166b1ec7cd537e49a268fdfc643782bbbb
zcf357961cde7fbb119252a1074cdc5f47fc356edc584750659fb0d28ab69008c26c460e9ec346f
z221d84ac55eabebada47ac19db23b7fbe7d03fe60444865f1c151fcf1787227216e54419fbd4f7
z64d41fd6704b0d72c89575d98ff10b08c3f08d11b7a7b3198a862a9648ab4f5e5d333622fd6911
z293d080148216f75edc94328209804fd96a7f41189b9538b7a011e2d498c0780f4a5d204b1f060
z978d03be38cc269e8cc3f811683d722b5e02d58cc9412f76729cf65306728a3799ec60f65807cb
z3dd39c79ce8cc769e721cdb7384f748dbe78e29e99b33d031cb5b627689e732a7c3bd31f069c7b
z8ca05c9eaa94eb95572e63d1d913e4eb6d6c1221c3c154c6b713a2191ef5029a3f87b2e625a92b
zf24ca495f7cb6d715cc167134451f3f300f89202953011fed35da1f93b7f6052e98b7d47735352
za7e3f34cf0fb17b1832afe8ebe607bc2cc35644fafd55cb35a0a6c0d312a6e4242007f0a2454fe
zd48df40fb3cc6e8f7385bd6d2b2c0fb2b51e20dd675913134580381e1b86c4225dd5eec1e02b82
z6e280190b99192230c91c424249ea2f6432fe515659eb2e7fc928fc2052dc3d77c8b2b3ffa9d44
zdb4af33a3424e90ffce36e1473a60b681835b37f80dd4df25d25aa8dba3adea76ae2fa443b9a10
zd85495970931df0d68535008fcd450f25efe7c632682e0fd868fc8ac3deec9cc07f464144e6e9f
z55a16cfcdfed3f7f45bf928291103d56d2c35c63f8f943d6b2d2b9ff1b500ada44e4820d163c19
ze2a2391176f0a5ccb973c323d68e7d82d2e3db5ce67bc7a7b6f53c7e32a6e6a00fe86db6845e5d
z251b27e76580d6b6741014829b75f814f9214c4c6e5118d33e584c319aa68764725cbe4da87cda
z73ecdba8cd0718ce37f13453e721119c70ad9972885b3ae32fbe5055d0b51fa8cb71268dae28bc
z68253fa801567ccab0174ebb4c193652ff8d093cc485bc1dad33d6388ea9cd81f3d2a5a00c764c
zad84feb1dafd47e6f14487a26229b18fed3f99ad37e8d4e96d6e0d8dba41fb375a0ebf07a5d1fe
zafedfbf96b357abe51a5551586d37ddd687ae52d06f10c593523c1b81604547b3b046267287234
zcdd821cd602cf52b0a6028d734aaf1eaf4b94761756ad91eefb69d8067953a9879b956df64f737
z3d99fce4fdbe05cbf2c3e0b5c1d0491fba92e5ca48cfa7af4464790873e05d9478cd30af1bacd9
zddbbd5f90b901ef93f3444929d698dd0d235fe5f56e4362e85bb02aa6eb2f3fbc867ccc6eb1b25
ze794081576d5e2376478adc9a1ed6015dcfd203c8b449ff2523941ce4cf9c2af588e5463dab919
zb1f6a46d11ac3c76d307674b7a22dc36248e67a8a92ee835a6a85d284dcd0ef3b3792d50d7ccde
z0d1ae1e195f9851ab2a50d6ea5bd7c43ae9780f378d89adffe6963195478e8b3009c9ee956cc5c
z204cbf98b805ed08b192760ba82bdd1ea7bb9ede7265ba992b884cf9ff55cd59f48eb21bdf4c76
z3114747efaac3cbb5e59526b026e28d597f07f4ec801e98f6758d224d451df935e8c7d0e07fa3b
z05bb16565528817d27d7ae9a00d4875b6d1f3bcd69828f9f0487e2d09e26e7426b1a470d92c1e4
zab2d405073c9a65fb0f3bb9980cf3a9c7132798970a5e8b1f809577716cac6de798de39c02e974
ze0e1d62eb972a014857099b6244a676488dff5e87120e1b2834161db18c979a600e19ecf342030
za93dc71bdbfbf168fbf4112c6bb8a2d77cdd2873bfd07167a5f4cb2622b3d3741ac736b1bfed5a
zcb542ad938f0797cbcebdbaa04387b8d1b45ce7a6a3c6ef889ddaed161992145191f2da7765522
z6301f31a08b6cfffe1f9b184687925abe23ef6080075f4e5c22c3f21e9d097a52071db75618ada
z76891d38b8cd4e3a0c3a3255999b1656f352e86a49abc150942168bfb6f876286c78e8b53b5d14
z83e052b64ab5529b35bd203e9d34a13fc3fc96859a64ee6a3247b1ee1cb3ec9826d9d0f1de31fd
zb20a562cfbc666a4b043b48bcca2e4023ac789870cb585c790e8d5d3b6fca14ebb267f9b9e2477
z805a7f05ca1902100eee098f27fd82f2f37276ed401bf6870a1190a8768afea7e3c45776db2016
zccef976880a22f2864311772f6145dd47c792dfd84ea5b41b818b24a70e3f6680f02e01e9fd2ae
z6cf25d233f43c1556e8569bee53f7c41b3c0a1b23ac1714e2168ed0e822403526c103e49db21b5
z495a48369cd23c95c3dd76eca73d05c06c2e5a5366824b01ed189356f23f792b25993d217a85b6
zfd45660ddaf1fcc0e4a6a0d2c9c9fbbea944bb7522f11481d68628a5260ca4ae16bafdb720e718
z5a01586fd69e648fd9ef36c71d0b84cc84fdee4976cad8369544aa9fc30defcd875b7ac4571da8
z818f966d81c2680624b6b3dfa4d680d2e1e0373d6a4a3b54d7a3d9cde5f8dd1c1e160e05385176
z8f6fcbc4007f9ee01aefe0df84c1cdfc90381e8c231134afa774d570f64fe3047575a3835fed53
zb1da08f5b9ef29e41d01339cc8f079c81275cffc3eb4cabaa88860d7692a7b8643294898178534
z5cebf496cf3c4a66978409483662f20cce6d966601954bc29fe31b04691333595e7e84ec3dba0c
zc956635955ee5df403c2e9fe8f31ee183db7d5efbcdbb8b0fc4437501d7e5aa6f057a35384d86e
zc7ddf624aa03b8bbc4d2e2ed8e50afa7fb6b9f8e86f51752b3637948be4f3dee4fff04991a71f6
z37e0a4307f2032566ac589e0f48aa5f81f18a3f249961d7a179eb77520e29dda170c7e29070b60
zff8155510b7389a4364284b90ee4af5ac71fcd7571638056d7c2ce9469d4098b404155db71bd88
zec4c9cf9623efd25f8d12209a9eef54c9de03efc03daee7470e25b9718844d9de6546f3fa9dd38
zfcc9e47fd68a2a1f22a99818313287e539ac6322f601f8ecb28086ba3e73b6be2e6c918b312b19
zc5de025bbadb2ef80ae38bf24b12a1e4d3787d8e1e39ed36df8a68b9c5d36988da612e3b7339a6
zd9a71f78babed59c8ed71e7561eba5886bd31ab1dc460c61773de1e585fc1aaaaeac4ee23f65a2
z08b744809042b98c599c5efee9a92614acafe17ad91c4cd456e812670b15cbffec5337c32d54fd
z0ec5f786e4323b328aa53a47a80a6cbd870dc5b13d57efff93e8d7121c8ca705092e272739d318
z631ee9b9b5f1ae606eb6863504aada8fc466cb3e5a99a373fc172f9588ac0d33295e97c73175cc
zf8637cda342c014250454d0b30993039643922910ad6e585f65c0ea25d18118124978777cf9207
zc0b4f5cc1c458680543c36d10bf1f63a1be820adbb00322a812068957fe1e0652d126631cbdcc3
zf274d2e56c36be30b085cb6ea7e680eb2a98e9448dde3a08a2a05d905ffb3439b000390903bcfb
z9490b822c769b77d1c410d7370fbbe68aaa0b61bee6ab3277933d2a0fc101f706502fb2b6118ff
zd395d5b0210aa5db1f25e20097beaf58fd96f0117719d9e360357af21e55c8e4f04f82942dacd0
z6f864d651596865e3f36fa7043189d86f446b51f213e53b7c7ae93f7d28a8ff717de44134be971
zf19d665458e502e4b1fa8789d9881625bc3d7f9d78fb1b0dcc41741083b4396928bb29d7a85e68
z76914d81c902e30cd0790d6812780774d08b1c2d8a6166246a211368d8132fc6e382728f612464
zf8128f4d0127f82740464861cee33f21212b62e28be983bd417b1801adde3ef2f57198a5507d9e
ze6c48bbce6ae82bcead6fc3bd5bd24fd5fdeb5bd3a39dede46a882d9bd1d7c628358a0169b8761
z7545af23ab88383dc0dfcda7d3fc9eacd2f6a338880a13bc28f09b2db5b909c7847cef9c5d0edc
z5f575141c0efb5d9c433008d1730108c5a4f09e8eccda18ac0a8da9f754882788e9fe3f5430cc5
z01b2fe62ae90846b881c2dbd7eee10dcb56e1a2f40f53b353cb99cc96ec1ba336b9b5e1f163acf
zd174f6e2de8032c92bb6bcc248fb2df5bcf529ef6925bac81669962f7342ddd80096fded12b850
zd3fcb794dba49f2cfd37b45582e6ee803f0a1266867e62fe2455c2a3e28355fd214e5bb1f5950f
zbdc4c2d6f71ff2acc364fd24f74b3c52a26f4dc724f9ed0a22d06296f6fca4dbe3dc4071471b94
z7e0d7420d3c97ffd90096b4143a238c5e7094c8a6f5b264d9769fc701f7bd8a8860664bef34471
z667023063f0e05e941e5048fae2b3f436c714e254c9187b6473c7df7be7700e3a5e6ad27a2ad62
z2ce0193d47f40c2f777f57b907cee5477318b38eed5d917a153f3a6b2e717e4e5ee56ef807cf4d
ze4f44a293fb19f8c514b78836a3c7517565f807bbf3654fe9c95879d86473aceb024f0c0ba8bec
z02b7e00a7d8c1213247668433a875c47d86717e5ebfae9384cac3a7a1c9a2365ff55b79c5a9b63
zad5f1adc1e27733ae0047d9ef0a8feca7f1b8831f06586ee804f0543c54b696b292ef2121b15d0
zc2212038ba8d12654b2d5a526bea22d04381b1908757d99cfae451a691509187a638005ffb4ae8
z34aeee9bd147c0d9d144ed7623c03d1b9f8af58319563fe6c909e79c27d8bf352e36d1886e02b4
z4857f090d12bcb5cdb0fb0164c24da656f43db43b021dcf1909762eee96af6cf2a75887b841945
zc0ac7fcce1d466b325d1e510e3322cd62c2bd9d81e1defac3036f9833b00ac21f719bb0fe46d79
zcaace94ba0013944f3c9d1a16e1fb999d6330ca9694c97fd4306465c3970a799815733fbaaafad
z0d05faf476d6e2f11670baa9706a54f0ab27b67d2fde55209116b9717bb0feeb14a0549d2909a1
z4f3ede56c0c5be8ecf56a1d5a88f0fd4272864ed729c62dcb5f0b05c845c64812085aae6e52975
z5f0fa7bbb1267588d2503a19de88d9c50052182d0f1f8587a6aab54b5b119daa1d9f4ce8d2f571
za4daf8d5fca12961982863db3bc53d186224c60d9d465f7e66df9181bb0edc3c04c4287a7de8a7
z483de07c83c6d1ea484152f95e717088a06149f75f4010511aa9291e7390b0a7268ec214a68362
z5a5c734f26500cce508ff579f17bfcc641a1fca39042c67b7b585ebd83d9e9b07f6aab38592f75
z10b334bbb873c62f82cf8ddc5a89f42d9962c154ba0f5fb41cb66a1d55628b4bcf56d9ccdc6157
z134f7f2abe4170677469ccaa534006425757fb659f8eac273ae89d8cd47818305cbdb6108fc9f9
z136002462692bd2c710f2bd76b5af8f48a90c3e594ee82085845a6af10abffb04c11ce15b6c623
z5f11b1169c010882ca3b2638cf52525170275844804a4b2b36ef326cc8c3495f622a247af50c3b
ze9c45978254d398204dbc7412c2164cbfc4e0620f4e53c5c7fc2634ed27cae2dc32073874332a7
z41e6b4a6744d2d8fd562fd83cf86adb99d0dba7ee3cf6af8e4ce5407baa30b06319fda1c2c90c9
z8d34f9e1e92b8e5736ae177ae3c5859eb1ef7a3e179484d6b98cd527751e3d60184ad52404b718
z205f7fcbad59994101d378aefb830f36a17a723cfec30da7b00a82e37d69091988157fbd432ace
z848675c6940fba7c3acb9d4d25c946e430d2f4a87b98c95b21ac623de53052f584ec67a0b80e0f
z24185e87919db764cf33b46bc2b1ac97a21f17c220a31301bb5b2b2d773e592d7a133dafdaf14d
zbf115048c32578e857c212c426bd3927cc0f1f57bace58b133c701bbc54c0bdc1f82e48b95fdf7
zb661b4175efcf99112d0589c9be824213efe2e15367181e4e7f6a779781d70dd1c902145ab6770
z9639bec06090b205e40cc17f56b0e2ab1896df3d3d1cf686de61ac727bf54d26978a842f66090b
z421e683d5120aa0a1bea3653078282d087da7d0844b0b9eb62d48a684f84bec2966b7f3b43b819
z7bf35a226a4d78728752731b42011e67bd19107a2b7f2dd8cd01f884b48477993e5ad943299332
zb2e0b955ca71fc2bc7f1148692ed9642a780b91d08992735eb92c6c9049d51b164da9350717325
zf0eb7c753132981c427ee6fc1853afb2d09236802908ebd558162a165322d2032209adf8b6c39b
z32bfdcb0bbadbc808e8329bad891895eefb2eb51b7f7e1b2cf40011f824e896d0d8955686138ff
zd4ee625766a534707476f968af78ea752eee0b0d8d960daae0354dd0d46a89b7f51d5b1fa9a3bb
z06fe63db1cfcab2a5bdc7e920e9985f06e8d19f28ff0c3046e7545ebf8345e2dfba91536b9e04b
z4ace9eb48e8bb38a076769f03d1d7e438a317d80d18488f98fd057decb03a2a07c9d0064217ddd
z64cebd8392abcd994740d73500569d2538e04b3df6aacd099ec65e2477a0d0f2219e0c6fc2d0b4
z2372c9adf4ef77cf8ec65edd1c94ba8b7379342a5056d73979842097fcc5def9fea776f3f79d5f
z9ebb61596eadd1c91174b319cf3fb509d16fa298b7c68bdb40872ed03f18bacdda97092d0e52ef
z39dd52be4b4374747ac177469682286b62a598deddcc61e3d6c47665ee8385eec8bab193666d95
zfd7222784ff95fffbbb0469f26c5cca8c288d37ccb1243ed6ec004825df920e407d2060cef66d2
z4bbe0fb461898bc03b99b9d8c0cb2ab848b174d7051bbbbaf54fcb26961d55565f096b0823f0b0
zedd921ac0ea03cb2aa49372bd7d90d550a4e28e8934c94d74a03ea5480b8d6a5b6c33077ea3811
z140a077c553ea893598716f09a58efc6028d601dbaeac13b0bbe9cf03756eb81467217f196ec59
zcf4d8a9c3de68ff6956849901bf1c09e6e5dd6965913b876b0816281ddca59eb3784d19c7f44c7
z31eff9aa29742872009bf8aa3d02bd44640737031f0bb506cbaf16ce8ab9f0cc27856987b7f3e4
zc58def4e2686a0f29ee3d790b06980130023d70b9c09a5cdcf6b57c6460021b99226d6c8c2a664
z9f285663f4252f661f16ec3e02624d7d76cb822f8a06b7ce745fc28b20e87a4c559a0e407f87ae
ze155902778c794b264089016336bab69d3df1d7575493ff9013bf01077d3c5356ef0540dfed5cf
z004f76a26cf349fd020cf3c82ebd037a7920622aae1f394677baca4583a3ba6a3d330599a9d689
za6d20f2ec016fba1230ffb6af8b7a3382e4b2448104606708f429d099b93de407a0ee6c465a95c
z6c0a71fd424327161fa8ef6d7016bc727d3d6426171172dcc798a2fe5a20c398d65045eed6760b
z29b9f47574bd586e88c0528247fd716cbae5bc3de03d39f6d6c078a233010be3e6fde0154505e3
za72475be14303b4d129e7a308d5e8058d03e5964730b97efaeeafbc394bee7f0dfbbe809a87f79
z594adc17c00b68dc7bc63acbead53653d6f4666a94bc8c516a4a01861d56b68c22f7e2b8ea88c7
zdaf79729280da487b8f0fdf1fb92773efef7eed397a4d3c97d581c5999d407177f18cde2d05f64
zaf87e086dde321bf13a3a277dc0f527634c182cc15e91ef76b10626e323bbe4b08010a61918baf
z4c9eaac910f4f989416cc7f0b5acdf0d000a07ba16ea73399af4a16d1d81c2e026c351d0746c57
z1de1723283c4681dee0116c6f34beae4a322bfb060e8df68c6a20a236ebbc45af352a724934de4
z8580d8028eac81ca089b8f3b7b4d039b1df284f977b49a9c624d201036c7e18132c3fd368cc710
z5246bc3d047cfc79c0751769c8580485d05d0b98796734ed7b10f8619c010714b875e1300210d8
z27088838ff97c9a1a50fc11c8c631bf657e43e85fb94af74bff55a808799f7b25f3b2872f2e8af
z58c4c34fbd72fbb426a69bd87b2de55f95f4ccaf308b245cab5c015b2d34cdb447080489fc9ea4
z93dac570d299f66b8201f8c1aa654fef8daee37e08d898db21825e55a17c84ef95bb0400031d94
zd37cc1ee920b4545f6eec0ebbdeea71e993030598d737cbdcabd9668155e53969bf8b3ac4e415c
z13b17f5e7882015ee51ec93d7d1dfc813d0df6a60a48adeaa1ad89b5b2c54cc9f58827fddb0b69
zfb5fe0ddb9c1896e073c400b8acfabcdb5fa80e158f035f56a156b8352c96a05996ad1b5bec2fb
z8150c029fbf04b8694fc9334d0c50bfdce655aafeb1927860a7cbab7e4e3411d9e2c925b0bd319
zae38804ee033775c40930e86759e64770c50806b1d4ecca2f64c8c3e98e6f8050734faf77d05d1
z70e93348678a88f734e0200364e38cce139dba55a6a15c1dd17919bd7eea6f4f6c9c3698429636
z55696a43f19016ba3e66b576fac77b58c41d4709b33c2e83a6dd7121eef711be290b1346157d3a
z5b69cbbd7ecf23eaa98ab4ce5e8a7616bdc18a11416785d9fffe3b77a31d4db0156ccdee56a253
zfbe7f263f4a235a816a007f0203ba79884274c62d15ee8eb2d1b5d432b5c99a174ca1eb00777de
z3b3df56f77c1333c2a36bb3fec15495812b485d63c54366c1388ad6e3b4b2377cf2d74b0196f27
z73c5c4dbf10ee417d690ee79509155743e1a8a80eaf2fe643a2b9fedb55a5bfb3744077151c92e
zcb01a21a183a562068a07a449c61411c8ce466d68689022a1a3d7999c854cba57af4e03425f46b
zee7b116c88785b6b5cb57232d1706815eaf9ddf12c8151d0ba5d0f2e418c3939de6667c946375e
z8ceae62328ac55966d67c3807791153848c15227814ece723d45c13589c4e1e5c40667c4acf56d
z2f8b548bc6d9369cc9d7505f699a16545fafbd611a86ac11d477a1f831688868cd75a563f45608
zdb4f2836afbded1c74fe1780320845f54962bccf0acc29fd368efc30a012def0be3774f5d38091
zbef6f1828b6a8e57dba46c5aa3443b43340fba48a741f13ab85c05865474b7e4ef3bf9665d0356
z62559bcda2b77d2d2f5adfad59fb9e075bbd9502f3adf90e1281bd783b77edcae9283d884a21db
z3f4892e6aab4cbeb5c22627fe39e51b609cb9c42721abc1c001dcc2dcf70f8a947fc3f2c1cdb64
ze0a83a191bc7ec498aaf2fef4c9622dba7a965332eedb01e1cc40177e2bdb838e85df356e59cba
zf8b5bd76d9ffaeb1f2ee63b11d3bca4035b9f79e999091b5f56a87ed84bc8c6143e21c2718adb7
z338d58d87a62fe3b59525c0688bf70253af353d22c203dcc90276aa6f08345b4485fd985de888a
z8e4ad96430e9bd66224fddf494b5ba41d0b1d1b3af52cdb01cb705cda71539f619bff2a1a7cdab
z711f487100afb62aa9af97f80d9b9996c0408abc0b76fafe0b02786a3fedb279f5c1c05d1cbc54
zb75e9b9112bfe8a4063cbfa07e5340dd910faf130cc33f13c06d0314b8982d24884621da1314fc
z39f6bd3d6d7e2ab1a6b19b56c69de9b008a52b4560cfcaedeee89fc95681c78df0350a76243c3e
z549a7e886d1d63c5f2f90559bae28f8c846b56f55b6b4d7a8e892acd5d8e4674090d3a9d536f16
z36d309886a2c18da3345a458d651d0c0e9c470eec7908e3c1e3a86a672fe96d361dd77cadc5e81
z794368d675dc3f50a33af38d1e8c0af8d7563e2489d7cef5fd8beffef5c632bb26835a75d4aba0
z1357c7225c54b466a4695bba1f74229237461533a37bf5c96b584a1a88633e931b69870ccbd6f4
z46be44dea4199a34e603c6465740d3b1f1e6ff4d3038baf8963236f5bed3b9ca706bbe47fd846e
z93ab1a4cc08c718753639e0189e28d66aea969535b749650521d9881fc9bd54434ad087049799c
zd1e595f2482cf315a8dc4338d62c0451db338a5688494533b2c65fc132bd7d5f1e4f7919482066
z60c00f2a4f365dc1f0b1738e2a33966ddd5390c2c5560e42dd8ea4521ad5f11f990613f57ab4d0
z808408c49340c1c091a63397f25bfa1ffa2b65418380e21d5033d89d5a9ed2f69c5337fc143063
z13f2c2aec2dd44376532054cf7084ed97f13dd02cfd4d901f7540da3ae76e79fc1a855c047fd9f
z1d291a65eee8c87557ce24c67855af7ef066ad0b21bc6fc88232eb9535188aeffb785ff800432e
zb7593017de9ba4fbab28dbcd0dfa32683e1de2acb4daa21aaf2a188dfdcde084bec08a76eab04e
z31f58b8d2b60fca72bceddda86d9f38cd2dbd83a5c96bf397b42774a6a1fdf3c0b004599c04a6d
z126f2016fce1667fcb7ce6e1d7f938d11fdcbbec7f79a33c025286ad7a21743f691c2ddcd1ded6
zea7061c13b93c3a8bb017fde4d9c9bb9dbd7eb7c56171f1b4aefd62dcfbaefa8a8ed6c68482b86
z3cb915d5dfc340b436bd40893d6e61b88eff82dc0e2364865db3059d27d65b5f08988b3310972b
z7c7cd5f974db7dcc0ec194a54c68b001eadfb8a43397be31263ab5465d737fac231c04b2664a9f
z907fbe6d8e7fd247de42a7c4bba6c57073234812ea75aee5d557c7ac87dd3c7c9a072dbfb7745b
z4b1ee7f85eb7fd1bd674f9ee7c80fd80b9801b7e34c9eab823de4535c45265bb2e07392c248646
z9a04a3faa312aea9751cd951cf169017433fe1c4fdc1fd4413c90802d2ac47b2da4a2b1c39b462
z89ee6a75a0bf153ea48fdab11d840fe26aff11f641a6c27e6a88a6057600342a7f42446cb1b237
z4ed6c35301aab053e06226907c2c496d1dae5732aaa2805ed677bbf4858483273ea0df40b26ee4
z9f8eb2429f8a3dc1589b6a67f053044b9b04e56f56576b04437753dd7f030b2749dc109d16e3e5
z8eadae0e9ac7ec21b66e892fc27cabb3816bbdc4499f61942076992680fc70b9d1d7d5d30f8882
z0cd3f59ed27999307618ac928f0a135667b2c5d5d396b0222cb618087c76471a4967967378331c
z49668090ee7ad246d3e30696374f6464cfd6f5d1bb8a27c384913eede5301646b31830663463e4
zd4702017923464636de8287fb9698d538d14d1cd6526ee89b2041f7e5998d0ca4e0867877ee351
z210ae75ad885787f0c42a7c5a2c5b61746ad36306fed5dae640f7ccdf062d6fd654ccf237c97bc
z6297779a6994d4cf599eb37b2a52ff94bc167e740c8aadf04adae645e4df984a915bb36a416bd5
zbd8696f0aaa63c411fb0e7e685e5c308877b5235c50b23aa99148962fb88b7cb493127decf76f8
z87ba2010c5f07cb42ce7cd2f9f2eff7368570dd40d9177360838b41f76eed4fc4b2c371a5694b1
ze5b631d86a602dec8dc9f2764814ce2a28c0ab4632481c5e904edf7bcafa7fabf7bbdd1c2be91c
z78325fdeb7cb5a89d197a82110e47423cd79ff704adc8463c55d042a0a3097f28c6072daefec08
zaeb7990a2f98ca67fa74aee94bd9fa1272fb5703866421b5ddc8c9b7bac819d48fb0d7b8e1772b
z9df9fe83714efb8a1b6ec557e1ad798a99f3d9eaf1f6497081d115e41911d12cdf8d8fade841ba
z97613e77b9648bdbc35355b3d228ca0a30a239fda4db4e331f8a943b6d1d7d108c70d586fae05c
zbdcdec8841d1f0b5000ead1479a99d1e2761adc6c264bf9b03a30bcf4a0536c87b892d9f3d9ad3
zdf9a4b63af34128938b9202231d3ee25a2c838a77aa68c99cc8df6023986ec080c8021503931cd
za6deb47f31e33b4d7cdfd4046e99134f3fe5a38f2958963d9d1fdd5fcc5576efbe4f4052271aac
z95c458bff54397c417b8d2363180ee0f62257080164a3aed43dbf4df2efc4b3598d85e0cf1bda4
z080fe54795f786fcbd4740ab1e43f8caa24a794521c054b2a5c7d2fc05b131ec1626cd1023f56b
zebb0134a452c7a2f79c3047e9f6c495dba5b4b9e57aa9c43361faf64b28da8225104a322f5938a
zf9da98a25823129ae3a88fc6a3dda2c30bb0b6cae0b62b7c78f8289d5861f3fb35eee37aced918
zabe3567ad3b1b97f30c6569a91ca2acdb5bc57bcdf28fa9232f5ba2e4f763dd0ca07179ea5d6d4
z289104f395c60ba800158a196abb168710124d8d7be297a66783535941dd156bea3cc2c52a0af2
z559a173b55b20f1465664c615c19af220b47ab6ecf1e71ebfe978a950c002a59e5c75ab72cda10
z5bb761af7c6a4390eeb74320442293f291058dfe2294e9de6454bd7379cb118bbd73101eebe5ed
z490e65f35ddd857c168f191d7a327203712d83a124a6b9706564fe76870d671e794d223a9fd91d
zc918a039925498fb6f7283247231f220df56e85bd73e05a277c7554917b7f685edf3c8123932b3
z84d694020aafe4c13427a37282dde3a0e4d9603c7e0e3380b93466aa98507166909e5135ee4786
z0756689495bb752cdfafc789baadbb8d1fbe68afb7eeb1f2b9b79821ad1f69ea07b25dcbc6ac87
z725457cde9b0856fc08bc33181005b79a00319e571937d112a4a2e30bbdf1eea8ef94944fe287d
z264de731ad5df417c4f1db37ac7b24b02cde082e44d7a2b6d10c4856cbe4715a7eda2d2e1d2c07
zee47b9719c26cca2c262910c0ac3c8ffecdd86594a3fc28896a6a60f0477ae4b9ce053124f1edb
zf2ecda19fcbb1b770c65aade5e43e41a2252fc12737a74f8a9366200cc6711207c08e03a3c2e7b
zac27084a29c54ade4bf6395c6bf6370c0a74e7f28684532a8717d081c30a0fd4132f5586ae9a32
zb87b619315903e85bdb722da5470bb5c7e06cf8357865d85ff22352ec2b625eee2b19768bea113
zf99133a8bb95bf9d23d9a2c7306d07e1a215bfa93ef8cb02dfebd090668a475dbc5f46bc23c89a
z734a975a0fd8b0ebe78ea615cea4e02f616ce9308d495b0e45d4bb1d070273a660bda10487547b
z7106d6648434a1eff33f8ca240a46569ec0a024ef0fc688541fdcd5c58f231e842d58c316e07e4
zafc52252015a79a06788751aeca0d49e1c837f6c325f0881289ec074d345c2af38facc398b81d4
z69b54f4613f5b386a39a125a577a4c6fe55923dd7d32ff8c1f926d69359ee670a53168cebc7224
z41dd6692c7f6997b58cff744b0eff66ad7056c548c0ec7b83dab3a8aea059440f8b678b37d009b
z948854a622489df01f076c399387ddfd4c8eef815891ce1e56c8eae798f37fd34b02b5b3ec9a1f
za5576f488c75744c7f05d3d46e04a46194d7a2ddfc10776a7132ec67cfbb04566a18e3b14ba429
z3adf5f787d40e2771b09de09fb3f1f1e2771a7ef3e9061ebb58f806cf18d0306d5e8c574c86d07
z0d265c073f31d3b46c72ffaf7502442687fd2f0c13259b1a31f9d6e20f1330d878c99145879897
z9d9c5ebb7682a159fe0042bea98d878bc979703e73b5a1d25f45bbbb9c9ecf2cbdd2bad3e49e38
zd7edfd28ffbde3aea6bde2848864bce9a1bdbd0364a0cc7000bfda50ec091716ea38412a5940f3
z944884e8e39b716c81ca8a31a34818fb77aca7d286b6ae4a0d0e35bbdd20b9efb39c7063f236d2
zb7cfb60a9c8ec3c49f7be204efd0ce1b49d8f2f46d074b37af5ea74ecc5bf3b44898d17c76b028
z6813eb4a26ede98076564d0063fb38f3f2df4dde29c41f11d98000ca2826e64d6e317c1258084d
z627f7a750b3fd149f390bfda6f9155ef3865b3393053fa7dc63f35f0bf9625472dd5770ac8f3f8
z9cb99827fd2c2c4063da1146f113d3d86eb61f9ff66ee6ab7c967c4a71293ab53a65dcfeb44c04
z6f50961d92687e6176be4a9002094c1c82ece0db364713de7907ad2e1f8bea69de0acb538aea83
ze5da60e3269f4dd0ecd2d1e1d90b1e93684d4f21821ea16e912ebd27c34ba6a07c9f9d2c073a05
z8788a31e90aef218b4930d225aab7a43e69fc55410ed435395e841150fdd9b5375aaf9f479a47e
zc1390fbbfef4c7e069c2cc34c13c26f0a165bafef4524e1be3c7e07df194bf7111ffd45f6e846e
z150d65606a1eba7de39eed5c2ecbd3d32b62245b4a2c9777e13ef5c76fc0c3c5422e6482e619d4
z2681cefdf523b65503b15b5b1c3748ac2bcd7042d71956b4b1314e0eb3aeb60926f3a03e430ad8
z07a70d2137d4013145df780097ba1ecd0f46f762d94c0ae587f732d3d049858469bda42437bc84
z8af603a630eb5d069cfb9f2f4d2eab5aed9fe0ff86f44034efaa001ce2112650eb86
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gigabit_ethernet_xsbi_block_sync.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
