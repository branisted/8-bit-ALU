`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc10ae40c1
z6b8a7053545f28cfde3a7a8170f836f6da5e0e5b2a569c0ffb6d279597cd02e015dcf0fe98e22d
z43d06265a264476e14500b9fdd10db3a0f09f891197432b6d7e8ea631250518c3d33258825a4b6
z61b77a3c7fb42f5e13da8f9543602a335f17883ea618d1d543729e2b72f28d76fe3358e9e796d1
z6da1176c22f501ed750baef288bf78876fcb706bd5adb9d51c6c460021f48b2459087350bdd701
z43bc692c17ce8ef19ee1b74ab860bc864d07dcf10939e8de50c042a72974d66c845560141b6d4a
zec940ea2302c45c073b008c2480572cccabf19d48b1d061d9c82ff0fd9c120edeb768f1fdcad13
z42fbcb275893459a47aa4def2f5ffc547b110edc7297d0bb14aa889b975cec2e97f16db658c1d7
zd50645f36d81b237c0bc2f5947f33fbfccbb8ebc6e3b79158d66d7b9d4353cd6a5c44d3569b168
z66c74935450356f1da3b3ae0c626601daf5253507547e258f004aeb9f37a6b7ff86e9067c292d0
z45822d42ab1c394df8f1c9994b27f3bb41f5ea4c772350a8f1ea55dc9e219d43b4b03625645b84
zed8be8dd294f51a821493f0fb90136cc5c9199bb36f14e95c4f7c4f838e467cef25a35f2297bab
z3e76e6cc820b76bf8d643b89c4a4f88ec075ebb8cf69cb7ea14715cf07b1df776df32505b508a5
zc86c7c42875dfcf7f97694aecc56fe1ee0542623df5012b13f9e40909127b4322dc0a5252a6f28
z90c0f6ddf40cb4e00bc80dbba2e48a6385baff907c393cd3c5d204abfdbe5f0da49d3eeafe791f
za2221ddbf5ac58dd8772037357654ac39ca15261708e78ade54c13879c4f8731747db65ee15cea
z32a020283ded1938653964496321e5d7c2daf6ff2c89858f500ec1181236c944f240980297a5ff
zb1ef4238f079ba8c531bf1100328a938e7734467fb61aa6cb1e31bb18faed66bb0f175bde403f4
zd65846ce7d7fe51a36a5ff8133ebb0312110c765d575dd76a8b6e8f7ebaff25e9a3ee34656ae6c
z52254c438bedfe4ebc8436eea779026e1c2e5ee71f1b7fa324118b386372ef48510cd152f8c4b8
zacaa246eae07fbf61e71abeac60e5a9eb848689d06838d5444ecf3f4d6160ef54f590072957c3c
zbe924fce033ce90890e0c34009696d9c68b05d88469f7b79708dcc2afa786f6abae4c03c7b1a7c
zdd8101d817a1ebcb602c50a82ea57a0af39065cf10d30015365831b5e6ed326d9f76e5ab055cbf
z5c4bd03209a89a7f767c0834fcb7a0cc395c3544704eb2a3ef7f4f874104362fbd95381511294e
z1a0faa5b2b44bc0083b271301a8011b4b6e08c5e6b4a9492ed12f54b8459d9629f60ded515b2fe
z63de2d6509513dbb88531fb7cbb8e2ef7b4d7cfefe2246dd290a9697cbc0dda87b538008de2cf5
zf7f5ee87d89e5287f89db46cd47250a0113e73e227fa08263f13540ecaa02b0d1fc4251eadcfb5
zbe364bdada07b013c284645f8d0c2d3cdb3e530dbb5b477455f65b53c1ec4c4a903c371afc5043
z983f42b498d3475b98fa70865d9ef3b5eb08221633eb871913e020467301063bb93ff12c600bfa
zad885e8a6b50a9b92f642dfd7df46ed1b553713c801266c67013217b1fc64565af4d54926d70e9
z84fe03aaceeb40946ec74fd682d4899fff9b6210b64294c3ec7a2001fe1fcad4b31f9be31aeb9f
z7008fb0f6ef2aa532c120c64b1fa7a9593a0c1e8d700f1d7cb715dd827d37eefb2e130b451231f
z0b777336f8c3b369461dd26e10bb2ed4559c71fbed675ad111460aad2807fd6ff86c247db84be5
z909c07d875c59eac9208c605d686339d9bb8c379b0126a648c166cfd542a7c7e41d8b9d99da5f4
z251d6146fae65115cf48bc1877e8bc8e3f7cf9db247e0e25222d2734c12bb3ed69f3013ce6e6f7
ze205907dc21d5feb7abc3a2d22a428061838cba2dfe9d623273ab4443eba89244f0918186a5c53
z19c73e32a6eb73e7a6623eb77cd9043815f4a0041ea680a1ade1850dbb1b6cd9e76c42a4457c1b
z6c4249ac441a7bf07556f0e6ed6bae08245eea686f0c636a076291b17d573123eea3cd1a3ceead
z529ed4c51cbf4be4c76e8e5c1db7ff619271f7c8ea0bca56e7b349abe84948e1a6df3cf9c451e4
z375a9b82426c8b2b0898bde7d8b3850913ac45baddbab6b78fa83dc1c7ec05d3fcc74ee7e4a071
ze8ba44ccb46a514362ceab2071f42279f7399854e8caa425d9b0e20721e9e73e7d61a6669ac95d
zff9df2ba8f7f02627cb923a6bdb9a4f4ba5cba10206f028c03139e0d24a92f9864f98c74d92df2
ze01cc68316d295521a1c86193cefa17726a541a25827425265c532fe34256d64cd3faa6428689c
za078e9b9abd252a79793c7f3b927aa342344a9c8c22b06ab6ebadcf37ce87bc0459d783e31e8af
z0cc6fbb30b2618c590442e7285fadbfa4dfd86cf05395ee8c2ec4b76611364bbc1b1d587c39248
z5902a82fe99a2191a0dd4dfe3aabd759e89d60ddf72e0093d06f5b0a50ed126da580de46c1305a
ze3264d21fa22c6b945a38d354b5ba64ee96d45eba96f1570e96de6db7f236169a3a38ababafd03
zfad83b7e03b899d4bd2435ae9f223ce526b805d67849ff68d80b4dddb3fe37aef9e19e1565299e
z056ff7ffb2561b5627d6a4ee507cb3e9681c52d3f6df09cf49ff916e199bc56c4ea533c556434b
z8c904c796a4da7caf65b19991901c4466785bef7b8e578fb291411b9612d18cb26bc58881a800a
z814982e6839defa511a43b63082f3d2aff531d38e4ba4886e7eb0b48481b72dbb942639a079d95
zf773b7e2ba914474e4b9db40ac735f6b70acf4d6dfe57eb1c334e6d1fc95597cc6c9a456ce95fe
z437bd5320ed56d15906fb08d5a3b88c60f1258475a3f45d75b62c04c88305312e73b430d498f47
zf1df22cbd5c2816196e9d0989dfe21dc72f380b65d941804a31acf56ce5fe7e3cf4b2bd8335b3e
z6251466a96f8aa2ee181c017b592fa0640e66535e7591da04265e7c720299a10a5998eda1648a7
za1debcf0d071190a855de014423691dee866c4639d980a44788f2f791e60b4c1077893c48c8c47
z6e227a7c5414e1e843c7167ae33bfbea4a2319cd90db732732dfd408c43e6ac83d6d90827d3b84
z0a1de7081b828b12bde0b4bac49c6f6e8586d34ea62edefd00dc48a78b6ff27a14ce345019763b
z60b00462e5f89edcfa44331b45528d5e21192e8d1676aa72c715b33be080ba24908a82fc723c54
z74d1d76c493ecead18c66a726c13069eb5e593f753a973950d405c9cb21ace88dc8fb016ff00b7
zce117a491dc4c77d3381ae5677bf471b4a3e3679c3f8a16c16972688412c374cfe0455ae04787c
zad7b3ef7d1b14cca835ff2d8059717f927b8be8ff196e4cf131c270a51c7eb64da2afd07612292
zbf813322e9916f0941674adc3019a8bfaaae6acb2d9b3411eb4b9cee95be924b91347e8f497d4e
z829ddc87d7e7edff2f241db9d6fb8690c5a87c092ab32025d6c7c234d28af7d8295fc36d6a0907
z708ee45f86236cc4b881e9ed128d82930a68380e834412105d79eda36e777797e58aa096d31325
za091c30ef1d850790bb6b4155bad0f3c52dff214b7ba44784b47e72491f124eb3c31d5bef0a779
za3228497e8c2ad4783218db9e69c4ce769b537f5379d59c95106901d586498b1c06d2936f68073
z92696c9d9f50abf4dfd425f6b3043cf31af44d22e71bb349cd0108a2b6fb8a01cc451c81f2ae6e
zb5d19f774ea21e2c55df3d9aab564deb3578bceaa9f4b6f9d4fd8ff69b6f92d415a7c52625bf5e
z3508b3499bf364e167adb08b3bce907e0edef46f8a5aa00c842f0983314019d4da24685987ef8e
zf4d7fca421ba2bc05d1275c16f59202177bab6ffe8f5af507eae0b2371f33c97f45dd692023e42
zb348bef5a7135345c2423f1fbf0c503c567ff65d69b8e4e5fc27ce67de8bf317250f2dd0ae62f9
z636a0f9d37870d4cda9b3349695e0facad2a8f24c9b36cf19646824a9814de992e06f8ec0ba374
zee692c35674dcfeb0b4000b6f7732bf75c8c38555fc6455e5062d762203380ab181b672dc4b81b
z83c562da2e7b4987052ba1b0a3982761a2481fcf1e54599e031cde009cf6d709d537d52a01152e
zea2e6402f8f70afe49600538911f36aa25fe9fdfdbc07a6377253be3d3367189d0b068dbc05afb
z9b4dae8f3b6c293769c42c503deeea5783c1ce27ed0371a4e7abfa9be02c94fd0bfc80857dcdf7
z74e3d8cff301265669d66e047df7f99f19ff0722dc3a429d88ed53c39ee899d3e332f8b48accaf
z4ce3c82eb3e9932eb03e3aeecedb09e56435e200a88d9a9e923dad24c6125f3a6f30cd326e61bf
z4ce4744af97484fe50f5d3619556572422c59143abfa2a82ff8e4d118df229f936bda3fd992721
zdbb19084bd2c54f7b9e427a76fd7b49088a9af53289a61d6a9b5946ef2a100f6ae989131a6882d
zcc9b55f81156a59e46f71ae9c66eb2081b1a24b19635b822a5bbbdb99738ba7a2dc940ca377511
z113d6196385436fa52fcc68d45323ac7ac5683b566c6f91cd20614953e94314b4ba5c343aa2aba
z2f793aee06059a0ec756fa6a5c387b6023f11479a563691be1a44241d83ad18766a8da15207279
zc9e784391e57212b9baa884e7a83fd825c518aaf5963eb8218a668539159acf68e5a8c20b5fd5b
zc547e56b25bdae03462219d86e3f7a09a27f6019de75c5829b088cf7bcc7be62856c7fbfd6d4be
z536949244af0a36ca9df75b3f795bfae8ff1ae1630a7cd0af893eb6f63f25baa3d61f04f0273d3
zc5153326611b32b14ff2e0b526cd55c10d0676f9384fd8ebb0b02c8350ccee1c462b3735b75e73
z7cf7cfc7d4b26deae880b4741248620149f5e86adfda613eb5b2d4aeba280969768c5c287e8a2a
z5ce975dd438165afa17aca4f826382b2fa4d8630c2367176bbb665c425c0ab09e898c6ef8714f7
z909871199d24b24431201e93a8307298ae7493a6a7adb338047c681052535b5fb1d684561d31c5
z03a6ae0ed9420b6305334a9311bf02efde1f9d33663f77affc2c93c7f1b0537758cff84c47a58e
zbaba2de90be34e4cd8fa76a53af245ca770ff7a04961dc00d05a0b84de2c3d3707b8c9745c07b5
z79f689ae570a18dcc2bb8552cc2b0086591c878d853ae1bfe6c2c0085115ef431f117ac4f53ce9
z935e3a5a6a201605257de03d20b7d930ba7988f5b46c2b1c1ce32b90c067f08ea031b869ca5e26
zb1c720ac10f5a03408fe9bafc41add3d9056c6e524124f6185cb9d80d09b5fe394c4d4884c0e55
z38ecccd2dd2bc63f33ba2f014a5b30cdfe06ea9e22a5bcabbd5710b738bdf2fa84137f02e121ea
z2ea5c4ae56d422f0f0ff0bacc6d9596f41fa0e849c9bd7194570e2c40cae4062ff2676b0b56932
zc91ffecba7cb1c621be64eaad3e7b65d11be041e6a44952277dbd71c79e9edd8aedf329dd4a901
z040e89b1405f1876db9bef8543b608d02386b4d92e36d0e634e38d8f5687701acc520d16f956ce
z94d0417d75ac4b6d9db0fa00f416be46a23f50abdabb57afd8f5cdfa8c1bc27f86aee8bc5d6ccc
zc23a840e85daf433be547d0632d6d769aa0171180477102eb389db2e8ce2fbc8f7e6c0c38c4262
z55548cbb43724e651229eb20c2f0648eda1cea1e5ade93b7107a2b442ddb3daa319ba38f635749
z7dbed148cd26f634d787b732027815cba8dc516565124b78e453e904b4c28207103eb8e9c1ed1d
zad9146e0f009d297fe224d37db6f7c70315d1223b9538dde0c7b5e522f3190af43335adf697228
z2e046476d965cc07042eded5abc6cdb80009cd174f1c7822ebb90eed79aa307c12403ef0747dd1
z86858d8156a26a0c9147aa2d7da52df37ca675765c0bd0d76130de4eb3ee618ae5fe1f675b7c48
zd9fdab0b400b616e605c4bddaac22d3180acca0e7af4ad3bb957d83c85066b3cc595f8407d09a0
zd63f27dbc63a149f5f1f751509f63ec0bdc0d1295aa106f208ff4c1ecb5a1944167bf7b96610c1
z05597baf16710085091d7458dd4d39b9ccc0d48ca5c3a1a86aeed0808b1779bd4b4726bdc988a6
za46e7d749fc09df2182936530d2772e6e98b30ffa3372c34b8a699c234a24aa8dbdc66624c5ddb
z16ee585a5cee5df6745dc41d45a9f6e8ce4bdc37d65f3c2dc224aa4c0cf95f0366eb5a4548f9fa
z3bb5e6248539c4582763edb8d57a7d11ad8f537ad64a377aa63a9dd0f62ea080e85e8cb2b4001d
z3deac4ae8a303bfcb7a65efda106bd608c33838f0f36291ca28c6b0325234caf075b257cc6aba1
z828b1767d213dd5a41031126987d0f18e2d864b0885c5ff7c2c17431d231a75cce00533247977a
ze9ab51320f0769fd93de271ce5a7b02f219165c7c0e97012adc7019eff33bd5820ef306a71bab6
za22c1c8f5ab08a34830b949e6e414fedd780d6065a2734ea3bbdccd495b492be1841b2e969607f
z5af227d9074bbc0d3eeee98ffc7114d450cc60f3affd4d85f54458eb059aa070b153cd947c5372
ze38555b44ac62c48390fea31566301b2eb98c47864492181b94b38998de05f66784df81fcd6888
z686b611eb525f627541d6b175c8e1144862e8263ce8c7362f87fa9be40b83a6ac8b76994375f08
zcdb7af3800072826937f4f08778523d12870accbe882992e3a96aed62bdc25007fbc3c16f514fc
z82bb520d7ee3fd984435346616cb92b25b790c8d8ab1b505dec7942b67c9206b9f17b970ba8ebf
z314d56f7c4b6e189453765a725efdc2e18b49b8de5d14d85e6227afbd11ea39e97e8f0c9f515d7
z20af36fa32f4c272b62609f894fcd148d583fc50a30704dc226b270c1f690bc64907404acce80c
z8c38b6792c62162967e1197157b6849ff785425d03f000899914b82495426103d5258c597b73c8
zee5504c93c50c04827db405284dbe4437ab9f88e15c748b5f57f1259faf31b5afb87a566a5db11
z1ca329f1b92b6dbac58644e6f83b91b8cb9959dbeb0f25277d2f22f2e3c66be86bf08fdc87b247
z3742eee75aa3e697c231bd84410ef44427d7f76882c849ed290cee30c86cf76fbd2f889416a386
zc3b9ac9e2ea5d4f36271be35a26dd5af53b523a689eede99fda8d8e4eabcadba85aa60ba4811ac
zc14c1c78e688f614e4d3315018d671423194496fe49707661634caf6d90bb0d68a255b9056c2cc
ze58320df3f6f98b1df43bdbe82b8dc66cba0e5eb2784f0f20730fdef2312467fb022a3af9ce737
zc3656721d3bd8705fdc0318c64a6c956c5d1d232a36bd1b934a95984e5b257c87571f35221704c
z0ab5b0a37e19ec39b4126ab58d3a179b90e6245ae6b92981284d5b0cf8d5048aa5f11866709664
z24b48fec04a3f9ff833ff6b24f5563a2e5813da97d83e088f622beac2bdc35e149a0e8699a11eb
zec30b7037f9ad374d675f81eee610f9a481559eeca6f21f7b8fd8f7ac1ce40a02f6f31f47a93de
z48af5f02de122b77c85c760fc98f0f8cb5e74eb1b2294e1223166425e75e24e6bc383c281f06ee
z6c9a947cb599f4f2ccb82251c840c93f5079db0635be64e1791d96320f368ade9e8352e30f94e8
z136375b2483e04efc1d0e9144b766cc50adbe46530af1f328a1deeb38d1f99e66277b7583e9e54
zc4ee6f3f82038348d494416b0ae0cf964c5bc4cf9dfa370b1ec93cbe1c0d81b9cb12fecb75c254
z1682598701c29252e82be6c8156012c93891e923c3074d754ea37b4bd013f46df6fe4a7429ce0b
z882cc6322a33a7ccbd158d9abc3d5b3678fd4ee7bf8fc821e5dc0ee1bec4dd6b92ee2a9c51ac4f
zf83cfae23a0b3472a8623806591ac2174b870504bac74a81b1ccee4b4cfd990b9c8f2798072963
zf426f4702972f1499e6847cccc48e75f4fe6468f4717b4852a691af4ddd1bdcce275199414fabf
zb4d1111de0635e9af86f0dc4c063fe8955610554ef3871d1ba0f4b3ebdeaa652f1e4b3f7264504
z913ed1fc69c61ae02f86a4d11917b41a27fc5942c5c887c965cc71577bc95155e86ad02ac1f1f3
z73980199355ff154416e8156bf2af2ac91e17b04b76ae3d8e97f1defc0cd44546aa1a73db9eaca
zfb2c3ddcedf440a83b81fd2edee3bf1ca1c417221969d6bc66be012d520ad270ab8c69514447cc
z7675e2a249fd3d1d4c71c5fec3683be617b30f1faaecaabfbd8470463184b42c1fe6575b19ce9d
zd856459c4fd218d91e82131da233b2c038d678f1e0d983177ff41bf596a25afc926b73e819fd9d
zc1dceba94a8c8587e171c847c3ee6311f29966f7e6f6b41a4b6d38f5f7b5b2bbd6f21b7a2e454e
z7d61448ce2a81efc234df8d033f72c2c016987bffb4d2b63c1dfd56fffb90aa26188da59fcc2bc
zaeac99aebc672e72cbd147eaa90b6f3dc3b6bd816522a228092151140bbac4ad2d7bd0d2a4d175
z0c3616d35f3f544e3898be049da9a28108ef137b260fcc5efe872a214f522dc37aa08a84171d88
z1e761972c797c44d68b205109b1bda8789f2d4c6e3a791a5943334ddd0cfd96bfb4815af5a7a2a
z64b4db112437432b514427cd55bd7e52d65db3ad913615ffea73813e6883124f9d0feb7da4c9df
z736821ae730d1caaa4ed013f7c7c52dc56434a7ed49d9248724005000546c5be753ddb3428eeef
zbb30445888310ef170dadf1daaf2bbb17cacf15d415af5ecd2de83a952966fc666bd1b1e43f7c6
z59d3c54a68a6bf815e7b9c1e017b86a54cf507f8da34b1ec17666703a38eea91bb21cb92656d65
z7f4e12b895f6294248129c783a722861fd635a7c4b1d8e5b9775a477208a791232514829a39bf7
z795c880fdc07be84e76927ce19263b5d9aebd57ca11e8b8dd8404cda8bc1476fb9401ffad94e81
zd74f5c88f2d6ae34c3ce95538faccf0646283f8f07dc88e9c494a0f6ff9934afeefdf62693acbc
z792b9f0a4bd7a5811c4f6b70a1c78b3daa00067fd90ae29b1f34e0fa70032d1eddad84c927bd7f
z69d28c5cee4536561ac1da0d14889303ec0bb14d0eafebc7b6b6e9e4885238575f532248f19226
zd9fd34ac0f1733f654a6fcd4744a341366e023291d7b5905955d939ab5528996bb717a98c9f040
z4aa162191bda2addf02d10061e0874b66a77ede38da9d65907caed465c6fc172a53990bcb76445
z1270eecc1f202dbe6805d615624c87961aad21395aa7818e9fa48bdfa8eb2f4c95def13a2e79f8
z2f53e99f4bd20a4e7d9b34a9474a1f86a9120d34b65d226c6e9b98275090e81c92d7dbf8ac81d0
z0ff0451094765fafd25e2df01f52a673214f71212cad23aa80120c39aa336d81716860adf1e24c
zc7f4624a329ea76978049b28c6b0daace4d5c5ef31f4c02f08b3876ba59b5fd66901e23a63595f
z078432bb4f843fdd13f56820dbbc6609bd6ff377fa4b367a5788213430a8f7ec6e9d3338da62a2
za1c3634a667e0b142979447f45d973f3d368dc1a18cddf04201b7191d84054e93462a629c81f60
zf3903d5863eefb82f3c1ab1dfb595e0d6f8bc045edbae090e135a0cd5bf6fe0b5eeb1233a85627
z26cdbaeeec984a64a7c27867e714c21bf83fe8595c95283979c894a95bacda6e09476692920a35
z6d869da560763bfe747aa89328f7ee24082fc79888be3d229a5491ecf38c1623fefa9282a4f99c
z4ddaaedb30dfd77a53296476ac8079ac5582e73356a045cd743f36a9963e8a5890b3e02ebb6c92
ze86b6a998bf2817ee57bcbb461831eaa6646f14c76c5d503a649620808bb872ee1666b18a6ca9a
ze56c38637ef1e3c9f544537b393267b91842b5adf9437ec2c95474cfa987916b9a7065f41588d6
z100f30d837609aaf298c2a113129508e16c5d9e08d608ba9992a5ff0a29b405a3255ad3b199611
z6335af8cf9833a77adb1399596b2a0e6e9fee45cb81d8651b31af805f4eeaf63e85663b24b4db6
z4df268fa5bfd438ed17d3fae6724519f495b29f4667ce2cea4e3c29ab047c17509a40ad003f94a
zb008fab2b8e96879e90b8ec74a1d276a89b5e0caaa35310f318705d52f3b9ae29a9d1b36f530ee
z3b4c8f4b6b3dce940b0826ace1774d4a859404bda6f5f3ada74e0b481a1061a5c5ef5ae1b50a3b
z5c16bd0d56637ebe43329c92275e09029f26bd0a65dd0848c0ce5795cb99e920358dae3a570ed9
zf23d5a8955c71453db331d322188266f0ad98896721fe9c894efd90977d31a5943276d1effb2d1
z02be3317a11db1acd8054e1ffe1ccf92e2d73e4de83c425ee890720d172d79c07a0d1c7c814a61
zbcf6d6287b5c839156948908b825bfa66b92f0dd9d556a3d5a8b74865c55d1a79ffd0cb6eacf12
z046e10bb548ecd7f618e4d9986fac0bd2f93c93ee51435d099c1d416227f8fe791033b87a30a28
z51afa23eb2ce67a901fda35546bfb9bfb0f17533affacc770fa385e7a1fd3b4e3ab5838bff4513
z269237d0eb82fd2257bb71a8393edbb0446dd4dfb2c1e624ed36b017fb665cc67f900c992d7456
z8100f6263767eac27afae316cf484b62c6692078b3cb864c8975f637f85bacb5d2a6a94761261b
zf77094a19aabac82b97e24e7957a768248b5ef758133265c7410a1b9f999db63c172439f1c8149
z07a4fda5e53d3d73223f3563f65232caa6e7124bb4a72903b247a52bf933eeb02d31f99d70e67f
z04499a2378305a71f28c92c1d30f42888ade851677fac1ec72c537f289b6f0c523008b0227879a
zfe4cbd2fb2ef1cc4b16d58c08a14b6fcc8b99c9af9416d6a945a13c38e59ca01b26ecc621d9828
z4b805e511eddd80c29a583951a368464c814adf3d788256ef4e8e67d5ab24e6c8878af5b2696cd
zbd7ffebd1f8a552da89a28b886e25a60e143cfcb4f56ea13ee1138ee45e2f81e6d8540873e1c95
z4acd0ceda7f7948fcc510c3ebd239b1ff5af192d576f180fdddf9c6faef1aa89e4032f21f1c583
zce74e3c9d5f63be163f1783a594caa22d6e943d8d9bed08c27eff268a2dbb4fb25d9140675209f
z8ad366331fb4280747b7fa93c3fd3a036d771943520452c05c94acfa0f217eb7bd4a2c84220042
z400c27e536793181481771201f6afea1045bcebc3e7a6403797dcd43f6150843be282ec34bfb8c
z30ae8a74b5af64d184e43457bbbd3202d943d8cd48dd5907c2a451291560c0c53498ba49f09bd6
z6dec2dd8012f1ada04088390921d2e47dd5b838ac5156c2fcf03082261f61a9de555a0da4068d0
ze72be8cb6b4b274bc3dbd5d40f95f19cfe1c287372cb7fe27033640a03510bbb0da132b7290eb3
z9108706021ea8fe778ff54324596376b96e093f6fa5f3edf248e116d153ab993da4cddc3790d27
z782bd2cf03a9994a9d952a306d14200ae6e2bd5db75a1e40c0b805c80cae801063be8568779c10
z850f4d0664826721cbc61ad248bc6a4a61c8805b57f9f6b15858eaf4ebb7891862fa70a455d518
za19a30f3a84e0df8710dec09c51337b4238d47e0a9916b4559abc89a7033aad2539ddfd641c6d3
zc2b398094dc94afe573aac1d5da314b18f037815ef3b0be7c6c6a228956686a450faf0564ddd2b
z5cf26b6608f1b62592bd83e431b12e89a39156d8d115f8a11ddcee079d1cb83bc2e30a8b20dbfb
za91286876eeae462d9402870339b2904fba26b6ad38a2172519a9f31364d15b04d2e1dfe792293
zc4137852020bb32ce87089fee9a7be69849a677494414c051faeee6b39ed03d74221a7db5b2346
z320de0db9b7ddc4f8e26d5f78bd556006217d8552cf0a73b22436aba66c5255b9e559af1a8cffc
z1d302b1d1adce7b4db98d690d6c6f915f71ad6e7e1b1fa8bd64b1d04a0ecdbd42c9c2d9cee38c1
z92aaa6de203dfaf960f54c6a4c35c52202a3cdcf0265bc43f94a7704c3535a7176d05958337930
z2b623f8225dbf0cdb2a02da47f4461c33dfa26607ad0765ce37ffdb207898a32fcfae27e288be0
zb5d69edc87d83e95ad5981305a49a0d8faaa309129397f2596686861436145c32dc129d3d9734f
zc61a34b83c688864c73b9ddcac032d9567865e4b7cb3dd0d9e83840c81d31ff8f7ee0599212f1e
z853e2e8278495e10cc8dcca80782b32769a011f585e8c6b0ba4917a4aba32a01fd7d6cb61ca06e
z4d5facc2e45152234085330dbafdc07c1088477fabc0df544ddd52f66acbce16df5e42f95de50e
z06308da94a89b0f9398a795a6bb85c3fb21c84e37234ff2bad1c0403f2777408470f15be245c7c
zd25512f06b9110504ecabf265284460f47297ba84f072b51d4ccdf9d31704bcd0c3c989e2e8f88
z47adb6446e1aa869d8562e232909492b07db29e78bd49eb37904fa93130d6cd19dd95b9a91b43e
zc3d1e4b30c95ca61ed89b945d2d468ff19cc9c73fb00348745ec8731973ea4c540f251b098da73
z64a62c03d49be86ca396decfc8cdd7335aa483ff094b63e874d448c2198f07d89dad03a6093d46
z36caa36992f86e7aeb193194b386e23221bf19b66a628235492f616629e406d06aab744030ce5f
zb3219cd05d033370c98e2c83e945088274739ccbe7a0ed3fbddacae2ff93378fb2b219dd011b64
ze5edf14263dfbdeb21c652a38e9ede285fc1a835f2ffdad9b41e8a83c4cbc4d9b07ad9d5ba819a
z41225d5a06be4be159f51122abf906203b06aa0c1fd767d8bc7d20a68a05adc70fc1fffd7ce397
za2a1021f3186d0229e918a069654e0b9480a6625189d3bb6c6964d161b122a05ac6746a755ae6f
z1c2cc67c65a3f38533a957d7d13070ecb35720c2f9f8e9730f5b47535c0cf5e785a4f5605deb08
z5330524f534f1b1c31bad52b129a9c41379128c0f82e0dba1e906bfb79dec0d21096dfe3f215c8
ze972677466bc624ae607608a075872899047430cfeb5dfdd48ef704d1e2d87827fd6ebbd129a55
zb25bafd25bcc04e4b31a4a931c56e5ff6fbecdadd05945f8e35375bfb74ef58605dffacf525891
zf934820851e8ff72744b15c1775a0e5d805e7379f818c30b02a54aac64b8d8bea96eec07ed6608
z11717bb2e15907ab4ad08921e0ec516ab6a80187f3e82de31e100df8cccdf96a3881a597587897
z1001acfdc93341de9c49d8b42ef8eaa25999c3ae19e7938095b5527c0414e793a042a469d85d24
z02e062979f0d05cb7628b30ffd39bb504ed81e891b9f432f32bd4fe7529554845979bef95c8335
z244122a56b5a042a94cf5d9ac8afb837f9b5f18bde0f37b5d91bfc64d7ffac1772719fc91510df
z35ee6ee37d08c26d046c5e76a37d91b06c2ce5e5d046275673948c832d4f61467751166ebe8bab
zb05a58df156364ff59ea3dc6dadef6c5b75bf13fc4c164db9f9c6da99db940baf3cc952b08721c
za7cb44e9e58ef32cceb18462e38135968f6ced971b296bea5d6318f9c7c29bc3491f81901ac210
zda26c4b8abf94fbe25bd43ec2397977c44093ed4780e46851f0b534792a11e15a09bc47c58a52d
z8e76f98d54802df06b1b751781d5be50f9017881375d190d57718bc0ea8af9b2b27a93e3cfc0d2
z0de73539427fa8a11215dd341af786d3071a2c9a2b418a0df6f9c424ae4dabf2b7f57478f3a016
z5f56904a6eec9ec4b460bd0d78e86a53ad77e76287ab8aa28dbbe46ec881215b813f317d60cfc1
z68a032cbc9bcdc8a58e9f6fe4811727a128cd0e244e48a08c6051a12bc363761a8145a31f01bdb
zc76e7d0510146d763ad44d19a4d6edd7726035cb7bbe9161785fbed85137d25903bdc3f4c1741c
z451f5a18c43a70430f45365e6641ee3461db7d702641a80c594ba166c1f10fddcfd56d6a6aacb8
z02ae378d1b379500e82d09c3417b2e046626f2bdc4aecb7fa936a5e469d864547d943cef3c7f31
z12b9d891af8de9e622c246da77b83c3049a0bc6066acfebed349d542e581ef89c6d8b3a998848a
z6ec8b9f306def8b4dc682a13e968bfd8a08d7a7344c8a71bb0bfe25db267a5e1ba0ca71222a8ce
z902d550101ac457c287cf4bd96726290550dbe3c961a4e4c336808c42b9c38a5cb48b93c269d18
z36e6bbf591ed553b02d61a1139704c3ac2a1e1a0c094a14ee4fa34907ec9fcc332f76a0f78badd
z64b2e6f3f3a421b1418effe243c0bad38125991cbc19338524ad243d2f4d4e0f6862b096bcafe6
z312d40146f33ca60903effe9f2fcaf34cac1490eaaf8ab1f53a2fc2eb753fc8fd86afcfedb4584
z5aa7b0b740301db262f44f2956f248d9568dcf9069ca78efc7d8c93d1d98ba731a6c13eb0f94eb
zf7d1041c400f1a5ab410aca83a3429c561e2d190d11ec0f0f3995af8631a0069dbf438acc096ba
zc91e42b5aaeb62dc80501037f4d3d1f2bffd4946f67b029452fd9e5408361d01b30b0b141309ce
zed24493d8d6460f47d79808a8c55b83f08e869531a4067f0d2292031240782ac76029964c2e44d
ze4a99917f9ae40cb28a82b652e22ce7df895de216949ca91b4c38b9766dbb4a91a058f264196b1
z89ef5cb285710b2f695d2c24184ff89aea60fa8cd38b80e5951fab8853ea2e77adaaaf6691d7a6
z032339afb79646ede658d6d97b32f2bddac8937c75c529a128bcbd03bfbdc4df78f64f713c41fb
z8da392b826e11a9ebf903552eeb54326a5f1c68da824ee797d288c32dfc607a4a059241a2ccd02
zb62f9f424b2ac08849c0aa90b51747eb1abb7973df5020c6b24d7117e46943698b597853e4d19f
ze8c0e8f58490430e46dd994f186abdf46d94864d14483e4b490c72b203960a0b720c195b1636b2
z1037d97b33c709503c9304711762fe42d7073afa774df925c31dbf2cc86759b3069568e3938a2b
zb49780ca0f9e056804b846102a665f023e65586e48b09af50fad2ae10accd7d92d4ce9d780b060
z305933c4fa7d6801e96c7b05a2f0742ff6a1be451afe607d96140b7e35688cda8d21a02ec4ded6
z013226342a662166e6cfcf38de30f1c1d37366ab6ebf9c3d01d5de65f34e1f2d1e6754071cd7f2
zae5fe30980f32eb131e6952eb68c0770a27c6f7add8008595dc066700e1179ce9192bdc32dc7d9
zb6908a764dc4b7d0bfefa671dc0c6ad6b419067f8b456dc87744ad68eec43e1c5313b6ec03c6ce
zaf2db64400f66c7b970d30a6312a568463a84dc36491cccc550347ff03b0e53b6b823c19dcc280
zbe97c47d0bd2ce8136d5cb9ca0c1f2f93c6004d16a88bc07d10bf9a2bf39484a0976cdfe87543e
zd8d750c847770c7ba3c8e9069956b59d8de4d3f953deae0d4a018c7c8f4d575a775d8fc198eca9
z78a913ad07d736a3c07c09d80705e701e63036719331949607c77f20c4922fb6f8eff59f39001b
zfab63da6e7498f36388963bc3c1b824d1c589f2be4f5889de7c31cbe87fed03102468761336cc5
zf87b94155b373034ad62747b5dbd29cb470eab60467eba0d46fc19502e20bc31b93451520cebfc
zb9b87a7841349bee64a2b3f83f6f2490d0f68109704a3b6f6ae9f7e61cba0fe4c936612bad01e2
zc822e3d43d3c127d229fcbf987b0c82f1a28bb67982bd4015c1fafe6afeb3fcb2904085a0ab0a4
z6399091fab1b6a20a57aa1f76ea2437d83d1384d6794187e81de296a648290063fb7266b0d09bd
za006dae9a2084bde9ae7f5ce1b3d359fb9541c6f79f33d859925cfd4e6dc542686fcf38807d11f
z243231f3f804181c4e1358340c5bbd46003334e4044e4f044021dba79c57788227c5a5ebec6e71
zca3389fbb2dc49190c440f22be5a90bd2acffb450a3043a9b34f035ec37fee73eb374d366c5d27
zd3e73899cb8679dbad9f2d0c9b499962edde80f8184ef9d3d3d980e9e514931c09bc685ac60ef5
zddeaec88df6e8e5f4165fc6ccc3b742d3f8ad95f298fad32a183c4f3b7c5c8d4b8b69bbc0a848f
zc84082efa20ee669908ab0b9495bf5026fd26557ec1d9e72232b125fee68f38a45bf0489d97f49
z7a9bcf0b7317294a2a0922002829e5b65cc3edfc530e71b881d9f7393a20f2a5d8d1c6bc82e241
zda591cafdf4e894506fbcda8129409f13e51fa64a1a9fea122d7dd0bd6f8ba8a30bf6bf72cdf29
z23521f6fb9be63fdfbaef7fcf4e8bcd3dcc949d77c3eb54cb809b7d393dea46caab2939e0e3d75
zb8857850324e9841b2e1f2b84dfcb39a6970ed08d5aa6283c9f4e81d795fc6380669901775d73a
z70e87f1f18fbbc28109b288e4f398c1d200bf40982f6f9679a3ff5b48af5b82b5995d4a96f304e
zaea436724e7a4678f7fcbd2ce7bc282e5380a8fce44d39e878f1cfe492d4287f01fd8b5e91f202
z5b445cb129e656d20b37a8691fc62ed11e5ced90f9b7486870f52841d99f397f4e689acaa8d557
z87a0bfffc6ea0f9c74a95c8c73cc7de7db8d4e36e56734b5896eef84bf6dbeb6e8c1e1243c0771
z608a2f3a9766f5f55d2c1f09737294d7a79adcd2c23b35fe17b7863628b21ef3e44063918f6797
ze09100e6cd765ba4c6d62ad3f099b050f7697d13adf5a104c59a93ba3f7161121532c511714e07
z9a27173f178fc260820cdc1dc76a90524e37c136a219add063678fdcefc430941177bc1b9ddb24
z5256c624f7a943ebfa75a5b74b66c782793960c3d9db155cdf4a2d31f7e2afae069b1282cbb31c
zd988795aae4fa62a23259749f12b55fa7e540174dcfa0b242bee95b60354286263dc0359bcaf37
z66226b6853cae50299489e067dfd0562465393892f84e409a196384912dbbcc7da171e816efa49
zd23728f1ec8e43cca693a5fd699366e631f8cc47e263cd3e7edf59447b39de79908446c4263da9
z6ba1e04d34b1777a962dcd51ec6c6477d8d2ccc41220c6c8c77b769e06a76e0d8d9535d11cc6fb
z559d3b815fa043de00df037693ad9e7907a3fdf6c91db39bf77e5769c3b03d2f370ee065d2b7d4
z2c8095e41674aab12f561d7b5d29a5876f4c9702cbc7480c01cb426352f917d38a745b664854e1
z90d077d1876a40092c18007a547083050641b9ea4810024d50c925c4b995272b601d93825e1e91
z1417da11671be379b7c2d1607fb26b645232d97bc6d581cd7fbeffe41098e74764c5e2b21b32ff
zaf037abdf26fa015dfaaa6ec3af43048b4290e511746bd4f6eebde8e27329834785f4224ea5af4
z7e4b5b9211b84a81698c82d86191e660bbd0dbaaaa8bb0acbedfb5b4a21ffe0950cc1fbf7fb4a2
z27a76e13ebf749d0ab333079b5a19e38967af0b2b0836512ba50d00a292c27cc35d9178dda6cd8
zb1823e56e2c3070218432406f70ee7e5636cc0a8421d3a34eabcfe88a2ab0039b3c06114b9d73d
zc508b8b03958eda0a72f6cdfe6825cbb92d7f64f065623cae824ed1d32b6a575f25d856626a8c2
zfc0bfa65fcc061c8e7c8c1dc9ddc30000bfb584bcc670e228784e65ccdf7e0bc7c4da282913168
za1dd5803306b8b00fcdc447bfebfe7f72b5b6df044b89a3f4d266817625cb031090e594c3b501b
zad02294bee183bb1df65824d05f15e023332dbe461d4aed936a97df11c59a49d7a7a0eb6af9d8b
z141ae0711a83b3a862be73de461b2979b6e9f1c701df843e4c6ec11b6b00828710ccbb0ec36d27
zb047de7e0ac87ceab0e8c686751c935500350fc9c97ed7d3e3e1a2356f09aea7f1a9f27cf0c57f
z7f82132172b2ee52483269e503e90a2b3450d5c832683a11d5c85e708d775707f0d0c129a53c9f
z497219e928edc94e057a0fcb3b7cadd467fb2e3ae996d883df04beeab141303f699ddb3f436ba6
z7641d5ec4afb1f61db516922a84472b9daf903030d24b41011883562218c1cf637098d60be14ea
za3a7cdf8fe52509dd8b4b9484778e5e1768c4c27eaacc9ec60f454df427e05390ba6106b798ebb
zf2b1cc39f63cee0658e1cd2cd2c2db4a528451d2e204b1fe69fd4ded257fca8be9147f8bc77dd8
z2688dd83d0014c0680be999950688e6d593c4bd5aeb6ca5009ddb435216122cb16554abde6251a
z577177af4ef5d2c83d0f9edaa7e20b3b7019977c4b50021f5f2ee35e14406992314be7f2340ede
z7f24446ff63900b5013b7587087c2cba070e279b15d0910c7c5501ade2ead9530b323a2268068a
z87be8d31f6cdef51623ae719dee76b9b0bb6264df477f7f826e5d0e8521fd7faf95234a9cbb2c4
z7c4234fbf8055c289f670a78da8ac3106b493dc2aebc635658a4884326c6c10ec67ba47e2ef1f4
z5d139bd02d285eaf480cc346d1600bcf8274ecb177e166b0202a67645c53cbc373072e8374ace6
z7da26f3e3ee3891ab0e806fb17089588aa39ed7b314aefcb1317487047bf4257fc54cfdacc45a0
z1e23058878b130cdfc2389d6326ea60d1de2a19e2c8eff1422c60586278a7208ab3520855c4e78
z5103dfcf29ed0b2be741cb847fcd6ddab471bde9fc021de45cf8e83076b10f15a8aa80a8aad9d9
zfe173e37483a670cec120bdaefd2b859090babd47580f593fc83f9f09355c06807815c4d11718d
ze130f28262e44c8855601cb7ff9d1e3a7ee584d755972c10566b5d81c834169213621b08221c5f
z76994187c4eb2c3f797c6e95b568d9ac97f068e78a0663edac1ac9894bb0a47d0898a6429dd03f
zcbd510a3c56359bdd1ba02cabb4aa7bc5bba692b9e1c98acfb0c618db43badd1c987ed4d9aba31
z57a9209049586d254a3b2dae12ca04fce67698908a4a37a9d2da4cffbcb81df9ba91a2e72594c1
zb31c257b6b54715f7e795e4a3352872a7d990ce0bae650e3bf63f9810dca1419dc026c98cbf8b0
z560b2396ff04dea6874b4f71f6ac125358e548148486d6b848283dc096864df09c49ce530a2c44
zfcc1bf2e50a9f30a1f283fe5fc0bf9a1b94033a012c1816138a9c984262faad069a31610b1ba26
z3d8acfda31a58b65e6c4ab33dc33aea1f0c022a9c12e5d938d367a4ecdbe7bcc96756cd174823c
z3f55ef08a6952f17a56408f2fd2c6492f85b0c44f166400ea8ac2cc2e16bf0883b7795c765c9ee
z6e4cfc2dff15ddadbee6be6247d47064955c5d04fe6760ba0c387a29b5cda4c07e539c18f034af
zd9da164e9b079edc5315db2f66e5eb30c72de164bd85dd91e7a123d15d0a5d4b803408e20e3223
z1c67d6a1bbe3d545e031b9647fbd1f3d726179134c45b796fe6c8693e03b8b56ee116de9a3b442
z61a1c270a61c097070dd231d185a542f3a90aa477a968aeae58b9916ae62149e2e8bb3eaf34928
za174636157f858f0200bf2c19ebbc19f1960c9b3371105a13dbd6a10c5f021cacb8ca3e26996f7
zcffdbbbe7db7253afc8bc77bab96882cb03e16be0b6c3c1ebb2e8220748808a0f3185413208459
z7aff73bc27e582aaf895afb8bc0dc3ed727a195011f247c506e3f7b0dbcf1d31ee9a5c01d682f4
zc3531f5744a9b6a9a559e379897a4f11931684d4baef49cee382eb11ae5184272939fad5938739
z2dbea54d7dae84f3ae6dc24de71fe58414b5b73fa93ea057149e15ffb8311331fa3b62fdcfc74e
z052b4eb42c70ac1832acb330291f00b90d9d3722a25cf1a4896663b77f8ae5dbaf53e37acf9f74
z8bdcc5d47673a8e04801f2da81b9462ef537ba9070ca998d53d0c108d460ce1ab8b142db4ddda2
z2645399f7dea96c45737b7f401578868aaf122181f20e2b47d0aeb8881d2d637ee44739f12c480
z26d4e966987e0adca0679171a45e5ee7781499d084dc48bd6b64c13183a09c9a6ca3a986e018bc
z11e9e208ab91c65787621e83775dfdd6ea004286a30f62dbfb611a4242a98652709e4cfb42ab24
z959fc7a298fa2d66bb4395f9b8b37d49f6ec39689eecf32c056d68c9c5efd39f4971ab6bd692ee
z95993f2e6119b536d4917e036f7a54d35d153ad6962ad5caaa1c38ccf0d97cac557e2870e1cca1
z57444a84ae293650cfbfbab37b9acdd4b009525bda68e94b522c208b69f767a5bf9a6d5e4c9ccf
z7a3eaf9fa914663c8277bc921351a9e4e6161b497d3407bab884dc25d00add0da7490fccc4a3ad
zf9cab70e2203a6154d2ac1ba145c759eb386ceda8d5776293ec5e087517eaf31ced34d31a58e67
ze879eaaf20457f99ab000f45f6c4ba73dd5aa2a44eaa4b3e51bb9314e468e2e56551202308d055
z954dc97e4669d69e8420d13da9c565eb0dbe03e7df87396c32a3e3d5c7c9254acfd7e4f21f0551
zaf8cb3b31a20f290cbde9fd714ff16a95c8726f634a285914dd2aaf1e923f935bfa5ef9ba0e8b7
zcea9d175b85bb8a5d8442ea23e84015cadf6f82a27702d05844e241a7f7fa846f8baf7cb70fdb0
za66ac15608c343c5b3e4a87396bbecee2f2bcf39886ccedeb0330f79cb560478dbc58e83ccab6a
ze66029b15423171e40630f7ab9e0856b489e1c9d942ba71d063d91116d481d54f92f3623c01f90
z2b4022c737fb47c7f87d015e7f27d907e3c4526a564323337f801a2c30de59d29023152b65d502
z822972868d1c5586d23464b11bd56a37fd3759eb815dd0c6c6e55b2b450b14d5381f2e7d7e04ef
ze23aa198743e2f518f6c512c96bb6902e29e1b1fe05c8b18753020a54671243c7d843011a1ce27
zcd331fad0725a8a3d8a9efe5d83bce51dfd2bd6072921d097cf2c7d2ff00d5096378cdcdeb59a6
zb65bf2938cca5f1ec95693a445a07b7a18b2d04f01beccca7d483c3aa4ea8be4b358f064f146c7
z0262a2c1c095a44f705aeab2f24dcd9d3a023efe37f122dfc74f892d910772dcd749d024d1bb2c
z4cfa36347670cd96585522a9cb879af0896556a2491b7526e374cc172086434a85bbb1d25be740
zbe7e06b3bcf4ddb0d3e36eee8343e3d76d72981d06c572317e9652978b8403541c4423d00f4bb1
z6e70f60c585db92e00d21cef4f88b7e55ad90f0c5e1e269e6659dd429a23107c656e523e0db2f9
zbb3f409482afd1f6aea1861d93cde2f1914ec905998d90aae6728d847b76fafd08981fd518955f
z67d2b429eb915451798a5da724c9c91cb4ade585d670723e0219bee234138551f939d03840ee2f
z21d88fe8dc4540871395f0868f9007a28fa4446578b46158560df0f0cc2f50e41741b3ad8bf18d
za2e9bf901c6556735b48996ae00d593255cd0bab9bcb562c14eed2d2ea38a78458e04f92693f66
z62f6b0ce5fd83f9cdb7971181f0ea77752186ec9ef0267928eaa91ef2230ad50ae24804e5b3690
z1f1063d313bcc70bdf2a068b3d6a7c1de0b4cc8a512b81770e86d33573ed37b18db4d6a3e518f2
zf2a9abdc2370e85d37fe7df5b007ccd96fa53491e434b169bb4694581e90ca6a1306157ca72463
z3458ddf68810856c405854122f2507a52c5fd5a99d51bf1c779c9ac9f96a830de71645a07f68cd
za9895c04d7a641d6400cc5a7c7ea4f619270ba8166db6e1ed835a177b2f7e14c9ab601edb9ff63
z612aa7c23e4653df5d60e7d9d05db676a95456a6072641b2f628e6f73864b6de8e8f2aac18fe64
z838f94663643f989826e6cd8128e259d928989319ec48f85999974d9b037acbbe5a216368ca924
zd6ec1c92d97664cb3080c1a3eba4d45151e16728c63026d968dd391b4465bdf2225e429ee242ab
z67a9513fe42e1f52799e2c6b7e673495a7b251e07b9c613f6e540f3ef46c60cb8ec73db6b09a1c
z9dbbdb279b8bb3c6325e07ca00a0a472298cd9d89ffa899432486911df660f2ef2baa7aaf41e65
za21ff30e355d9e3330e52bee70c89bcfb329bbf90c1e1a32c7f89aebdd79ef914c24de721367e5
z67d4aa334bf0a9434ff1a36e8074a40e933e4841305588e5b0b26b4c0388c21e4ff9365e87fe7d
z46970818972fe03ed27a46eb4601de72798897871f9963fab563db053387d3b748edcc307019bc
zb35f898550b22e157a0a5d2799df1c97af4950c35803eb6de3fb4c916c0409d9c1243edb0693ca
zec71eb9b6fdc51da21396989d7e9d0dc2552473da1a5ade2e1b39ade2a6ff87144a43e76a4cd77
zcf8b8756bd641e73a13afe73816466d0ffa9d1a22a742818600d2961b6771f900fddc6fb84e884
zdabff0009ac030068350b774f4a531a030a7a320533abfaec029efe3294ff2ecffda4edc8a00f6
z7ab8dbc40cccb58c6e3229d5d427486e30a722a5005b8d960c66091db11bbd0e7cbc89c3507189
z111a6408ef8d5a4cbac7b64c4ace25b1136045a016eddff7ed51ce6c7daf4466f4e4cdabbefe8d
z216ff6b332424b6bdc2237c85b0a5706db01acf5d1b74fca8c192f7ed61068789212f11ea79bd3
ze3fb4b7e9589500d3fe82f9160f22f3da3a42ad6b24b0a20ca7b92c81afc7460f0a7cdb8f0a135
z5b1b4c5d3553f0c00d5fcfb750495a25c07a3d519e102b9b4f6fdd1ca792be077a4aefda145bfa
z6cfe9c388ca08b059cd8253ff4576084570274a51fae8beb478f9d828f6193affaf6c105706e76
zf3d00da28b24a91e7a68c7275c7073fa0cfe3baab922fc3a93d2468bcd0de6c99b18f8d67b5388
z501fa6a92c798728d061d6084b37e9e46128f53b0e101ee1385b23246f1da120e04c0821ea8979
z18931ee5d282cc4a539caa7bc46d8842f2f760fb12526660a68496e6e6496643d4f9e3914f43f7
zaf1cfcfb6175278ad3f00fcb204f3afcef5658d95a9e39a7bbd0994af46fbe27b0d00b7eb3156f
z3129e22865bc26dc0f9a55ae19169b8a4d2ec24b0e061bbaa0b1fe72b4e56e0febccbd02305ba6
z2302d3531fd9c716b74412b2b9cd73f78baa12952b652c7b8a9e71d34824e600b828be097044d1
z5e710d6e424a59944132656d946e44112e9870333d1b159fc1116107f615b335e124b2d730fb66
z17dee02c149329e0235a4034fdd8ffb652eb0f61a16dcc911cc25b797a9652df423f8be33d6cc2
z51a0c9e30b570801bb07b5e9bd3457dec2658a9bb5e85dbd9873d83829e5e7cba199e51244e12e
zb7b6c25324f8aa6621ea967247b578fb89643175dcae9d27ac19f8899861f72e46a647b0a6721b
z65af593d790215d223e56b7ccd63481de3893fe5ab15a9818dc60f58a0d8b76fec1a601a13327f
z60367a5f382e7832d12360fb38b3e2dddae4ea8053d944385cd7e476f98ea5df83a20d2664e1ff
z1874a13262472cb1537af7969ea4706ea7d994311ed771ec6a06b69ea97a8ff521ad4bec288905
zae192cadd0a3efed7b0c5cf68ade7c85ce3fd7a3888cbd5bb4f7f0374e9ac237f1b1ef665c7a18
z188c3c67912a48e47b58841678f0517777c460b225aab3b8151c06e7c3c5d34aecf1a8428b4f28
zc1e9f50ddecee6cdfb0be4cb7e220158def0dd98d9262d99034dcb3a0a4253a34189c1be893656
z6d29b8bdaff358057874e5a922e9c1fcdba363b595092e6b147062ca44df13f2f18ff9690080d9
zafd8cc20bd7c32b6e8b21978681f68d3e6c165d8f0d756b7d1d7fe535156b06d84d06fc9697d5d
zd5b5c14878fe552814b5867cbdda22b1f43cb89db78f723e90e422ea7b4e86ecb8840e27a3b072
za7d4629cdabdacb571abc6f8b2138d48fba2fb274379a9c50377b8618b7ab98ccfee4fb12801a6
ze670b0edab2d827b22cd9a2607103db8896c81ec842c305691cb4239e707ae0c8dbdd5c1f6a487
ze7d16500d8d127d17b31ef2c120c0674ce3b32b00e6e862a397ef585f154e7df4e8e231f7884b9
z3305fa1eab6c4faeba3b55e77d09226a3adeb401cadbf4407f196217116b3c4ca5b09c05ec8554
z2cf2cf45c38879063df925c665087400151b408ca019714439e0e7738dda57bf217d9221d706ec
zef85c558f5c56b84b3a0d88728facffd08bfad64e3a80bd7a92c9de6107b2499bf83ef25035031
z5e916091c2f156bb7919c5f0208ddb57250c7c45c9fc6633be0173e4d99f1f3a0b32ac1136c39a
z96c7aa7b9bd18fc727f1810d0ddc1f4232450d8b0160ce99c0684454d549a2e67c540c4ca777a2
zb5959679bc6a7f08e7bdf938be920832994fc25d2121ae2cadde062f793cbf27a1c81c9f89ff1c
z837f604c0646b8b334fd7d352adc711ec7ccd4bb7066498fe711686b1755624842bbecd93d16ed
z9d1056a236a86a130d278782c934cf2386f8b1a81d3258555a897f8ddf4b126492438281c0ce8a
z02917f32fe68afb94a4e6ba8b0d2a1953f95a7b7a37d25f77d09c937697f6a9086946b5c94c8ff
z4c007746c891f0098e3ba35e8f00409eaad99b6f8df1786195105f4764bcaa08855fe3b30bd85a
zab6ed8c818b66bead2292f89d7356757ad62cc036a18c3575616e402bd900c5afd002a33b06b30
z5813c02a0b8a7803de8af988cb96cbd62a7704de814a3f72a539fe841729bd6d99c169da716999
za14389a42c73e66700f2ecb595920e4d218b2252c22b1e7720bc7c1ca22b3816b3ee8c83f8003c
z7c541a6a23081e41207a533fd9dc71ffcadb2ea1a4ae2e88edac942fc1c2ff40128e0fe8bf76d0
zf373dc72e35f5b79f15377d21932816dc1c958e2777b3d31cdf8b2c8dce97545d00ea94445dc51
z039f0896bbdfd1ec8473d2f9107a3522199a03238c6a1817adb1caf9a4b26692ed0142420fb25c
zdec0f35c56dc65d828502b0182712c9c008a4ff941c84868524565d90423798e5a15d8e23ea071
z0053f9fa9564af0619e18636963fc89d64dcfecfb626cb2cf671afb83c7c672f1005ce4e6b3253
z96d13b0baab663c61b9315be6d882ef71265581713ea0c36c775afbb2a8961550514a68b51603d
zcbe2341f64061ba6787e5e99240ad62eab22fd2ba3c709e68a601329edf0e4c7ba1301bf61f523
zf06378fd558b8cbf153e07925e97eb20ef6848ca21094b88bd5afc1ab019797e46cecf709d9413
z3741f0e603305287c502aeb73bf54eddaca2d07e7aed6dc62b5e6eb1e7fae10aed37d05ca06750
za519f593d6412d7918501391e08fe4b62026efc29105f91f49e6e2e91adefd12ab7d7b23dab99f
z556355eff8719eeccdfd0750a92f12d69991a38c534978b07d3d714609ea82468e2cf9f9b77d5d
z17bc1bba5ec8fcf73085caa42b50cc9bd06d584470f2fa92b03bc7228f44e05d71fc390d6fe9ac
z987bb733d9a7645f07fd96b89d0ac6df7020743a19e03682c72b55e1a6ba7c25ad74e0d625979b
z4bd04da153f3e7ea74b28c2b5c500c7c265fb03e3139474b2cfa044fadf301fca46d1944c389e3
zf76ccda35aea0a60cdfb780d36b4504715a3dc9bd13b3c85006ec2bada23e3e2058a1a78dd98c1
z01982fde3db557c1274893a0d5288d2e892e0b5915b21b6288978d4b4455e350919111f83310a9
z49d4e09f1afd8007c759a8fad5b747f9e3c195c0cac10f01e8f31f04294a28d93e8fb38dd43806
ze77068670d25c70c513d7f2afcbea2408c8d4ce9ba556fe26cb8f5618dfb4f8516d081ef1170fe
z0972f89e13249e2f7b2f26f37e389f8b83fadb3b8b88e987f3bdf90333927020c26911795931f9
z72f93df9f88830a55dcda21a952ff2d60e91303fa12a4272c17dc1bebd87b6fe92ae9babd33e05
zcfcbcb62dc2c4d4138fa8cfc42c76b1742d8df0de0584edebf5608be48c9c4340f38f017697f28
z9776af91f627e28fa4bcaf3c68cbff7c1c9f7a7fa6ae9a953479a21d33016080703247b94ce23d
z0a553aaac79414636219603018d7874e64b44f6112426451e710471505f6af587c16df2462bd16
z76b38bab81f07b03c56cbb1d63723afea09c24438f58544665845c7b10dd7ddfd5393e3b6c2052
z3ae51ad89c0a1083d524699f05fd28a42511c458be33df040e32d4e6c4a7946345ff27054e64cf
z5f3f73da58114526fab34b31aafe78e3ebe4031209c79dbd0caf952bf3e891914bd5d0d5188796
zde49eb322a42a4888b3e86ab6065c57382ecc4b3af51a20c0b868801162ad5b8c16f20e2376aef
zb8ca2e64708e252ff65b173060782f85a655514a7cbadef2ed40051a121d1503d256c0c40a50d3
z4618b2cd05711c8c985c34acd7ee5a1735808d8c2c6cfda4c8c596626fa4fc9a51c3917e7ace9a
z6ee5292793534626206b25db8062be22db52514a9d7c322f570ae4221d997b477fd17b405b9aee
z96d30664af91f1387d1b8b5f44d084b7e6a640ec474ed82842074405c155d3272f8ac546f73088
ze88abe03367441a89f1906e813007cc5fcd41f4bb6fc3fae652d398d6efde1b457bc39ceec205e
z304a1eb2b9cb3cf3bc9df2bfb92928c3d1180ee382f3c0cc9b36d9e7a303f7e9bcceaffb704710
z0a4d7f2e91b1e5b04d4c7782fbf8a932fc071748f683fd7920d331a836d33a18f180220f28c4c5
ze66a0b8307e08ccebd3a01e4aa954a3bb945ded549a762a0e9f9f6740c94baae29678236a01fc2
z3fc1bdc3cadf8ca52e5d9bb33b396a18a6efe074b3f92c43ded2dd6a1ef525b76c4b5c8717573a
z70bb3a80fc40369f493b46355d4b2d8d8e8f54818534f9f4f88d9774ec598733bed4d254ca9ef4
zced8d875b9afa92ddc5205802f2c7a7f7f64590b9d06f746f3c9a3d377e38f9e302eb86590894e
z8c7eb57d79fdb0fdbc2c5aaa454c7e4a00b2eed8177d053be7913c94409dddfb92b42b530d30c2
z7ac422885f6448b9bcc3ab155be7
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_bus_id_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
