
`include "deprecated/analysis_port.svh"
`include "deprecated/avm_global_analysis_ports.svh"
`include "deprecated/avm_stimulus.svh"
`include "deprecated/avm_verification_component.svh"
`include "deprecated/tlm_imps.svh"
