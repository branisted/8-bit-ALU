`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab30857016fc53a
za25afc8341302f0c829d94450c399b8ff9b0386c187cb854ee330605b7b59da379b1f26f488e1d
z36e675f0b1336408b3a1ad87d0723054f952fbefc8d5a33eaca6ef5be8f42bc59870a29a5cc9dd
z4fec09ce6e44cac279651402e7e1f590df88ce49ec26ab39f12b4a02855703c6f03b1e85c797d7
za357087d98e5b1f45502e45892e5823d6fa4b762932009620038c05d74efcea7c3fdb38901d620
z36515d0824367e48d1bc182335f158c262d396cada6b0ad58add4f945eee634c2dceadbfb5118e
z14969c29a743830a07124bfa78707f3952b96b0db7af7c9ff36f77137d8c490c4f79328328069e
zd7d5280e4f95742c9841340368b9764f0f80413adb175ecfbdf3c40716abca7b8cef6f7fe92ab9
z6bd2453f1aef7f7899c5365c5c83793cacc7795c269413f6cf0dabad14d40e9285afde8c01a47e
zb61893788ec5060288cabde8fb553f21b02eac61ab0b48ad3d54f4d1d76508b22f0c600861b5ce
zcb30ba708be817b1f50f59c0f6fce449203e7355c1be55b662fef3f92ba58243d81537761af8d6
ze27d7864d2dae99372b2b75bacdc0437a4f7e011d68c3487a89759e3625548fcc920ad06471ee7
z2d701aabf726859343208b0a543c73eeff8406febf277e3babff437ec820fb49d6b78e73bc2353
z884917487d35a6cd06d7d73ccff5f0292fb3df6f439aded7c8bc5dd0187f22a0fe1ead93318eb8
z8c6e90111edd2a748769a8d92e19030b0323140a1ef01d3a257fd16256b12b03810bb4a4e82398
z2704088d587398546935b6339280ed10cfe93a3a5b7a4f04e0a6f073f8fa718c2f9190d76f588f
ze9fdbb73c2c6c983be7680e758043939fdd6803162983f37193ecbd51d83a9df901bce5c960f7a
z91451ccc98f8cc68bcf6283cc3f9b8b51e819fc5551032ae29e1442013c19407df90f462e3e41b
z7c1aef3f9d51b70c68d822f0a422fa0d0e5ee892118ff089818bf687c336de5bd99d5e67e111a9
z0e2f62ed4ad8dae27eada5c5adafa4af6c21b4b091c6956691b57cd90801c3611d8f6c5efae18d
z0ca89bcbcec2ab7d43c1df3b639808f2cd136e5b0e449a403f6ca74fa9ce29d080fc4b6d260b41
z0bea847b489fc0e0988c2dd46437bcf4a79b2002d8c917fe4f67a6635bb4caa8fd752669f11436
z97f630fafe293d60a75d91cbb564256460b29007a8355b20b723f94098afa5ccfb198245ef0a34
ze2d50c0c0d30192c2d703aac3649c51f129c8a7ec465ed495d05c83e5fc7f2f432b0aa04a170e5
ze0ebe0a684a840087019b424a8c5698a4769a9d055b35782844f95ba152c91864daadde086267d
z28bb4ee6a4829f763dbf8d226ee067c490dbba97aaf738352a28c2cd120ed53e23b6846c1d43bc
z0de485a439515f3f53df85e009d272495b76219831ab3efeea240fa622b08698453ee00c9717dd
zea1b733fb28a66bf9fa2b0bbd1ac1b7f6b795d06d3af1afc682d40b6772aa903dc45589ae97018
z351d0f8c543f0f9cd6f9a7283a72f34d4b39673779bfd14e12b2447e8dc8a6531affc41757878b
ze2be06c3585e6f48703ac0acdb4360c70f8b1841b8ff983a90af20fb2f7aa84ccd27299ac9e397
z46f67a64f36c7149f94f07c521737536d56c03eefd8d678aa9f5c39752369c1c09876dec201748
zb430803c4c424fe74d904b77ff4f076d5f2d23635c7ad25abc2a77c23db6030c819848038efb15
zd2ffcb5988f590bee66dcb2211b478898acc83121cb18468b7340a1aad347cf34b464f956b446d
za9c6c554d3e8a22ba14041b6c233488cac03fc6cd60615b13f621e2a7bd3414a93449762d38b19
zad8a8c08ac4180b575e1c906df7cb1e8cf0c584b8e519a074336b1801f16e60fde5b716598968b
zb06171bc4dd5425e999af325482f5a83b4623874dc5d936a7533e8babeafe717f6b3d67b28654c
zff057f8e9fc8ce4a345bad5ce4a309107283828681129f4cc499a86928e235e99ff60be250bbdf
z595e35af95fd898babd1a013734c3bda778a3b0226109f9e2b80707b85190ae48a9e53ffd8afe9
z1102603dc7e391dc1d7b58c928b5e4acdea925efc23ace1d2b1d8ec32362c5084c6eae3859cfde
zcb34edaec7eac0753a5e8c38ce7342dc740a796b6ea6ff3d255da750cd15ce9482e40859423701
zd80baff85c3be48686f6b2136a793197b5739f7d86de8baae5f719d4bb83c017fb6e773019eb21
zea02396c91be63ecc9678b644737f45b95d74a65e9a82c6d69c06bb31f379a5868e820e9ac1c60
zdfdf65cd7d1eee75ae32288ed7dc0bb097a97779bd54b8164a5b7f528208a82f5dcb39b3f4d4e4
zb36e52783b2c8a67fc9a86bd07b1f7b68d32db8ab1ebb5b444b3495b7910d39bbafbcbce080c64
z3f06b7e067aac7a09ee230edab5549a23431b69f8ceb55fc0e43cc4d05b0ac812e86014db7cdae
z2eb9e2f09cae25701ebd0b3c498f910dff2b23f4c7b39cb545aabe0680e83d397b8887841bd161
zdc2ad208a7c7fe16a01d3bbcc66fa6687024bd6754da3c7e9ac358418e147803e44b426568e43b
z1f62d218b3b157d98b42e3c0280c4097e9d52d16ade9239025cc904b7ff795efdebdc0b43bdcf1
z4b55a093112f00589fa99de7ead3acba15ee3dcfcd661288cd9cc7cda04e7b9725cd12b3a29f8f
z8d3b09b440e67539a59bc9aa4d4a1081dd4cbdaebeb832f97ea2f476917ba1ef29ad7a7776540f
z5614e60a41ca2ce9682dceb8ddddd5f86b79edd3464bf17c030267dd87d7da0082a0847a5e35c0
z965704ffe903fb1a7ae20c6ac8f0b5a35772b702f9263ca1627aa618d561540648f3b846cb4f93
z9ad2f91a61a9326970bee42c1a36d6d32abc86f6231066b82afbb51da9f936d6beef86ed56ec2e
z8f871a7b41a7aa7545ec279f05ddec4d1b69a7595607708382ee0ed27e649b6df193bf95e73268
zeb2b2614609b5417df6f1ad8b340b005ccf74835ba9c743bf3a24eb73ad442b81b08cf19dae1c7
z767cc59a8fd79800dc9841033c400568f62d9a6569b6d477c1f47ceb594d1edac43fce2df56c7d
z2d3c0780a01d19b441f8334ec0804014745a7118c1857315b57ea95537c80c2500a77a616ed8d0
zb1d7f756f48a121c02f8d23cb4b3ebe7370dce591366b9324025645b0f7e715132b49efbe9a378
zf902903ce9a065ec8651317978b46cf3963dd96abfd64e4f1f9435deafe2a05da1afc48e026056
z37af1112997d2f0d55165368b8caa443f5129ac73e16cd764b1877f04558ddecab5534ff2a9b2a
zf7bf3f550628073ca35bc34c6e4908ce5f0fcca26bcb390a728f971b744fea065cb970bd9c6e6a
ze1e9e15a99f174d4e7b9c707e6a69a4653c5fd0e873ef7dd6d512137780c515c202321753acac3
z21837c2d3bd13e307a269a0466382380620cc15150a3680d49ea1ae72fb1863cc1fdf732b18498
z5cb70276a6b8a3f5d77b0e36af8061c87bcb547dcae37d23dc520363a26e1581264dcccfc77628
z7bd88e9c0bceec4b05b5df41a8f5b949a9434ad72d557194d96a93feeae69deb36cd36fabaeff4
z2dcccf2f27a5d59f2208dbd21898c78df7ab295ab834ba713100e7d7399f9fa75a4152b83b929c
ze41cb3746c963c080d5ee48ecbf53328b8a76562820c91bc62dd56b663f0887e0d58accfaadd9f
z73dd6e030a7b8af32f7150b52a7294b35721de8de633cae72ed708b820442b2de6ed999f1495f6
za4d2a0cb6c7056df0759e32c6e02199e548a1fa52783bdf25512939f5be288d0b8e6855cfbe932
ze1319cc312833869b1d40d7291356c36534f4b8da171bc5ab2b336c39aec0fb1e6e65b2504dcdb
zd1d5954654a0139a4759071a613005a897ccd5b1834b436d4ecb2501ae1fff26e36c65da54b210
z998a6d98e3ef94725cc4f76eb678b7a4cea6b375cf8fb50de9de0e88521655d0b462c971777751
z586c2ae40205e688711bd14d5fdb5de68633968be8345a6bdcc25bebf1aa261393af053847e083
z637edb0082345c287fe7782050ddea6c2be012e3a52197deea8800200d2991785d1d4bdf5685b8
ze7aa5758f48fe7624faf0fc47ad83fcdeeb5b02897cd92eb57ddbf3dde9266f6c617c5daea060e
zd925d7644f38fc9b99c06e8e3ed31f8d83b0268c76c4a8aed465da7920f2618b940f5a73cf9a39
z77fc86e380ede4dc4bc7cc5024548527a2f2c666ab28779654c32834f3bc0fe360d780c4b16c26
z6ce976eca6c38422fcc68ee1545c785f62e5cd23e5644977c1a0d7122362b647b3d0a086561bcf
z52218938c0001d128470bf26e429c47b76330025b9e433bdf06f488ab879d1d57420efeff7acc0
ze3c1f0e49448236dd69e40d225e7a9022a20a224e52c512ed2efe8d9ba2a118868b5dbe8546be9
zd7dcd7955d0e194620d08818b8c179bda4316fbe695f4edb1f2769cedc7fe93c183801ceb20f7a
z4a39228aedfe0910606a31bbd8e1a6290fd74a2119d0220ca21ac7d80cf60152f5cdcedc3afe71
z7629e2d475ac2a3dfb0c0f469f1c57e57dea699d4d5ac224f410d0ecb7a174f14422ba67364a83
z3717452720b35800e2e9fea09c76578072660cbdc948a7baca646a5b52387a6064242dcacba91a
zdf063a3816ab0a2c256ffabf2b7e803fa1535d7b7abd2176fbd8f639c4b44030a5fc321d31c3ca
ze1e237ee7ff7dddbd2f8a982afd3156f201822392e1d4ea8b4ab412090833fa4fb1d21cf9e6d4d
zda8e1d9af9cd6abd153267f7c0e6d28efe406e5a729dd4712268c4c5d33b0499f1b96ff76bbb6d
z89a49d21c25a168fb48fc85a0fcfa71a3b8352f24b2e2c3033257799b42fbc0059b20a1aac4e1d
zcb24f2b3917d3c5fd54852c9a2b1d3b45b96e9139118157cd66a7552e23a6f205001dd6feab3d8
z27c76d239ec94b5c4eb98019b8838e000fca48c35edaf3a9b2456cda7aab85af6e6ced8f5529d0
z15ac4e5b83054ab002b2c82d9620f5ca9d018b775a29fce95a9f358189735c66a3f96966aecf90
ze64e91f446e2bd6ad88fb728c40e741c972f3882f887f4a2bbf938c744ac44a6bc6d732af429af
za94745ccd8fab86ccb4fa44863bdd64987a03eef21f0f0da8fd40a146aa90a5d9dcad57af91514
zb724dc648e6447bc4951203b502fe2f84b689ec4dda18aa50aee5c22952c48c293a01481b63775
z5a3a7bedfe745fb6cbcf5ea98fe3086e3f523b1b53788634cc0d74d17baea89e2667d8960afc21
z37a92611386d4f250dab16a1f685a8a132afada2274df84426e53d83b567f50151335a3c3a3bbc
z33814bb13d089e8480c3180274029abb036d87d424715c1f8376227fd85a7c000f68f65c54f079
zdb6e5340868d35c5640e97b28433d5a0a03df9d8b8668ab9bf6fc525189e988b2356c426b15075
z4f70a0060e4181d898ce7c66de21cee186d20a5d10371e0d86f677b7fe7e3c8e9d8f4d28c15669
z7eb3e21b0712953b7ad5a4fad478cb5b740cb47b7c3fc4a9742ab48ed795d3190228ed9a63a9b6
zc041d613408ad714a0c123e5cb282b2df205ea1b1e22f2ca8a45c40a7577bf8e227ae638b0b0f6
z22f3b8d3404bcfd3270c4bf9ea42d647e4ffcc1bfe3d1170eb91edb436b446305e1b2dd9c7cdda
z7906d7cd19e344519e2cf2d004d38944f45e7c53c973a90405bebd47bbbf305f705616ce0758c4
z8ab79ca7a7daebcbb4b178ea88b7095511f9e363a0ba24cbffd0b93f9a66477b1a918470ba19da
za714ab24f2839a61a03c003d7737d9c5a5324dbbf996225be6f0d01b26ba2adf50feb41496abfb
zefff55c767e4f9b4fb56e68bdacc1816147064ce67f0a6640a88023b52810607b81230563d2cbd
z3dbf42ac62be7e70c1e36264048c95f251f6bcb675a1e5cc87c7d1cf8d64c0812c70e173fd37ac
zf27907bcdb9948ec99b68710978041d0a3bc7fd274166a2cfa9d15afc04adacf6dd12c9537a4a5
z315c71c081edd29f85167ff83b4bccebc4824a68851e0317af707dc054776d8e2feca333376181
z1d11fb79ce08ea080aa9d2ed781cbfe300d814168d32257fa9145ca09d020923efbf751a2703a1
ze83b507c2864e1df8a467f9b128bbb19962065b4817c5a8e000a085cbb0d1c428e57851d8be4a3
z00c7d6fc47b0142a7077fcbb8ab6b2055394f83552b6ed7865424979061e632b9744555f050ed6
zb30c0e7edb3248a8d23520dfee0ef53a0118d0a95ae2a6c3355b86fc417803270825a13a07ed75
z389a142d81c2683427b7339dfd0d9f2ffa8e8c3e3b6c917f79cf7fffb4b7027aa9d8d00dd45e57
z5a353ef4af7a57259a3fe8bcb1f06adf6bff775d2f9480976edbe2e800f4b8d1bb16040180cbd4
z407bae2e5f08a74c99367232cf67e4d6d508281a5d42310c21fdc612c3187456f67d95eb9616a1
zc80e8e36e789cdea8396222131aaa96054609782240059aa63034cab1fe6cad87ee41d0ed240f5
z449db8ffb5914fe21214fa59721579ce31ffe2c6acb7a621f523e5fbaaacc1ff436abb883ea753
z4f238662860f338ccfc920e97c7e82717baf3f21fc269b09dd2b9e4fa1c509851abd94c63d6bfc
zc6d86be4ce3c1fa710fab364048fe738fd6101f354a6a50004235fa4694858a9db38d1d62a589b
zc13eabfaffb1a2df00ed82b2d4da28873e03b1e362a46ddbf0388217723520022cdfea55b6344d
z64b15f9454dd2b8f07bc51bc5e0c590fd83e1a18173741eae4da81199c9a2d2928ab56a309507e
za59217b426129590ff64938973ef9192db53e4e46ab7ff881248cea00ace5ab9334f76c2707484
z0ccd2c4e8aab414810673306804eeaa6a97fa0aee9159400a1979a8437be3c6f00001531040013
z577b178556f2d8e02c56d69fcea027acd3dc3c49ebebf3f39e146c2c9d7c1811ca76f9836f1da6
zbf611a7aa285d626f58a2fc91e09ff02cdf31127d013d3ba61224f89234ce3262436a6031b7275
z99b094efeaf4668f4630ca4c9f276cfd8432f5544dbd84f1e3bd50b412bf43afa5c2db955af0a7
zcd87778042972231d9287118971fb6b11d5f7332efbc97245063a61267b9834468c065425455f0
zcb5888aa73d47c764e13028351a0044645ad645b0956ddc669ae13db872aa0e972a1446abf75ab
z6f103582dd2874f39e17bb7b964adc03fd8d6d2954aba30e67e4e287a9200d82675fee5a219513
z3f19a05653bf4360792c7a4982506a3d2bdb953e7a29c53266e6df7f2ff19b11f2c7691c9b8554
z986b57984e0f74b4e1ec369a5626d6cd11e0f4bfc575e71b312c1c640c21af5cd60ed35cbef086
z8ada597106bb8ceec06fad982510001642c99355470f82af301a9c1f4d823358709e07c792a92e
z0cae59c1856ec25a8bf8a0d97c2022d7f9c8f7997647a6ab348fabf64c5ea625801d984ec20ba1
zbcdbe482cb703d9787aaff2e2ac41dddabb2652ec3d2abfff233133edc4fd8d6a4cdca19019276
zb3747fbb32d0847ee6155671d96b2e09347bb05c4fc0353b6f54ffc7eb5b615e6a3dd198c196a4
zb13c176708d80866c43cc6aa4dc3a8f1a4e87a452f8c80164d70236bba5cceaf05944a1ec164dc
zd24e8791e15727c2dcfc32cb9d279c80b2c5876e639317faa45bd0f7bfbc9c1fd28f7d282c23d2
zfbaf341dd171e93091ba427da47e5691d195363b6e71c61fc5b43291142aabfcfa473c89b86c17
zed2cecdff7dbe22842424bc2294f37a84f3c2c6b3295890ba089ea4681131c8b36d6ebb5e6d4d7
zeb6f37b0cb883bd854bde73e904e4766e7bbfe5ac0b8f4f91a4353dfe1ba4bfd01a3ac29c9b7e4
z94d4099b492b70a3609e3d36f5dff9038a99ba70d3125a16996e8cdfbc2d1d5fcbeb3d0b270952
zf832bac4f6fa48557138a48fce021b2ef82c0a8d2481c9047252b7d1bed3fdcc2f341c2bb72018
zc03a39887b1f7d390e938f76ecef1e8e162cecaccaf4fafe9cb1b7e5565275005b85573ffe4064
z7b9a829c5bd89c2ba13b7fb321d87ca743eedb45c49af31d116b9c42bba6ebc2971327f58eb8b4
z207e466e4fd5cab07ccc06c8d8a478c312e31fae2369be61bae60a1d0b3297f90ac734df13b8f5
ze0569f90b129e08798d5b6cd23dffb0a50da4e86d301cb36b81ed5a6175d72db68378e08564094
z164a384ed930b1591adb5995b831ec63779a52fcd55e3498ac816d90e8ae7dc1067a69b7c264c6
z4eed94e5588a3c7cfd763fd183a8d46eacddb1ce06fc862643853e137a3361a891ae9d638f163a
zee205da54cf0505bc238f1916cb99dd987db8f8ef243759c295a54705b922109a0c611da4917fe
z626291c1a64359d4e32c53eb7284ac6eb62ba3785024e329a9cd1342e278a234c8ca66745c7340
ze51594456b395a766636d5f05102e3e948f58ac56a5ffdafdb20042fccd479b0a1940e055fb682
z50993a070dd615dcf872be08c93f3c5bbdf95bdbc80da3c46cf73937d66e199770bc6cccc7c3b9
z1c49b5fbc20b30af39493e1ef14d3a21b1b42d9d794a2b8535c56cc08142bedd6b629f0b3caca2
z2ac2de5b1754bad04e4cd77348e67c587387f549ad4c3dea41559f585cf5278d448f4b52a9028e
z85145087dc7ee8769ecda02fa585cc03c5f5602ab04451ced7f4f827b51d90623bce99ead0e7ca
z62be7cf10da6ca5031dbbe615c86350ab92c4344fcf82d9632a7e27ae142d80c17f7e9dd73008a
z30ecd64813cee737061ec07acbfe8ab2ff45187fdcbd58aed4feff4f55e3e83a74b4e70c72a5b6
z56743c54bf52a2bee461b5c421a318ab67f745de1c1b7625e9253f1fa301b915ea0d846acde671
z320cfe73ceb2710cfe806d3a150c6f76944c1fb81e7db282a85a3603960794ecedc1aade0865a3
z79eed4c17d1c07674925d9af68d5435fcfd0eb834904b25d6a208cd2a0d76f872193b9d06dfe68
z610a7afc7ba5694a5a8606a82bed48ec11379b77769a2d244a000a54423b0dc17531677c05ac57
zbca1fe082f3677b67d15a599fd0c50433572d9ed9d40d9f9fff0b40afd61d82423f9e7e969c5c5
z6a27307affc7ba5cdc3d170fd079e66bf7f982e0b6af8d7c41abaaacaccfee2f4be8b51493d030
z1b1e29db945578841a735a14210fb25888306ecfeaa06f2b809e7e8b080a9b48b9256e5e57764c
z1c4b824e2ba9d6fd68138cbb707131a9934bc7aa82d3200a508b46b4bbaf655ff7d861ba8d0ae8
z67d80765d4de8536a2055a69dfebb5f899a87d15a6bf2916e424b24f4c15fbe55b4c58cb4dbd45
z838747398aac003e7ad9c24956e3047c2ec5bde3152510f0340ba665981084b0c3475e51138aa3
z790d4e2ab8fc6c63ef61b5e648a88e8de5143ef6601b74a816781ddf5fa5a396cef04967544ded
z357d51599e8ce0a4bdefdb8b221a2a98b0404698305a97c4e65d77947da563287a2510559e6934
zb8f2f8cc66ca01cc8ec560483e14e93fa4e8051f23a8f548a3d041709211d3634af45d757e9f79
z770c570ca4e7e8e7cef6212102ea018dfb3d46ec9af44bc805b202b2147868d591b277a414a3db
zf6bf486f7e0307105a6d0e48b6d08fb579ae7c0d27840077f3aadcde4dfc0dd2e5829173c34364
z2aa28d9d0e6536be697aec2e9519d5179cc94c09874390aa520df5f4c8a4f48f2643bdb493c8ff
zc8ab72caf327cb047e2cacca4f3b17cd4566800fa5a3be0f9a28ac9983772a788ea08c88f37740
z18f62999ef8d84eab10ed957894c105274627446621da45594e859783f8c5efaa1421ec1a0471e
zd45e5859e790647c61203d4606fe7f49914e532fc8238d10d3a9e4538f0a0332763bf1f8bfb6dc
zd59093f060e99250f9805c907dea30fe2c071c3fbaa51908d50fe3e094f8bfe2988a38705d33cc
z96343ff25e6a05758b76b8942a6cef26fed8b5574d5ad3db026cd337d0dba17831020783fa4570
z3f9b95f1fc483a2e3900b38308f3cfe4b53c980eed79bf87fa179e3ec4b8187ce8202cfa827e3e
z980284fa8ee101a9429e5382a81819f7acf4c86272bc31c2a52340c997e65b914426b358565779
z97081a3d24d37f57889541641a25dbd639ab372e5ca6137298d007799175a8ce1ab776a69172de
zb3df3d01240cd93d6490ad0de07a902cdd810b5d8b38900853fd3569436bc5af7debbad65e8f9c
z2b9d42f52528d7b3294624dfde5334a13e4c77a7fe164ba17d9c9b243c01a8a1d0c73fc8e8072d
z1472a6167a1e6d1c7a2b4e61c4a6e805d16740134424fca42bbe5df1cc395e0d2952280d8e9133
z741abe1499b3cc891244e3cbd7a3059e083263f9748e9d1c7d778e71661bfd53aa499e9386d0a6
zf786039b57f61fb03b5b068871459b7bc7897449ed4e69bf583cb559da2735047b950f3ef8f22f
z0bbcec532bd3b6e800e80c711afd09d51bd82f045cf2c5d79256ea3044713a105d09b178837d79
z65ade3a74167500fc71ce1fbb54acd5098657a95a63cb9a86c4c09ef2a1f98a372103787d92d67
ze18384ad7d4957d12765d9e9a5058ace8baa94acba13732e9ced62b2e12ecfed5d221acf2825c0
z3b330abd0ea523b9904cec3237ad37523754c06abfdba79d5d89220a042e4c952cbbf36ff4d5f6
z8e407b41da99cf6492ec30b9838cd15416f8fb29088c491eee3eb7c4946ef49cf961841332d94c
z5c70bb8750e2e02b4ae8f15e1647ed65161372180ee4619ab6f6223e06509b772600c31f69ed0c
za6b0de361b1e974de896757b0a18f635f183e1d6e03620334d169e89e0c673cf608fefbdeee86a
zd70ca9d66692fc47b0f6618afc6dd24e0d89eb5ca239baddc1fee03c159adc8e9f2958f7480a3c
zff2c785946fc7979be62f87bf200a0858bc91e4d0aaf2ad8557ac3f959420a41a68137affe1f93
z058ea377f24bef1ec4acd81610da487df61c04ff6cf14740dd9c6722d5a92661ac0ad5a5d6b5a1
z146e9b965beeee1832642dc44ef308368c8e324c67c22dc4b345faaf87c4d377489f9938c2a62f
z8460173b776942e60ae7a1d49519f7cca0d1acd44c40ca52f383cfb6114373e4740d383b6a4dcd
z77d767229ce485dc4e2c1c65613f18d4bbd815cf197a89bfa0fdb6610ba46b07320057358741d9
zc77ed8437e6414f2bf3ea3474302a20ea01c05f5f03c92985ba828a0bbf0d1fd848a8733a4371a
zf452d5bfc3f68c74758138f0634a9e15c5bb0cff4e92c94ca27d1e0de04dda4842a9d51a93220a
zab31e4b14f4749860faa8b37cf1bf6d66522a92686b78f9c83fc219d3312251a32140adf23f0b7
z29a8afb401bb26099575dce9c0638189c4322c254b4f451d16c16eca9824cee0256ea0702954e5
z73d208d419968512f9ae20de1af192bd89f3f612b4301849c191e2bdb8c109c277f67e30cce85a
z36a1fe0b09f7d96d6fd159e13752f535a0f680a6551c8598d1196d819bc5dc6042cfb6b0b15385
z7e84541f485e683829f9ac817116282bcba823927e977adc5a0990e12d706260b1b58f53175450
zc568b65da2bc6ef822d7c45139c9723829e2deeb9b91cd2b2bfbf1fa1503ac2a88a08da60b2ca0
zc4e91ead91b732194bcc04d1bde7b479cd31a9625f69102fc570feaad04c8b8333954cfd7c7ef7
z7e48413d00b3fe740dea336ee50efca1bdd9deb962cd77f8c3dff81ea45c56150bc64a107026d5
z35dfb0c8208e643efaf84d31355ec412ddf258a41218a4bbae27d2c02de020217c9e41f19d00fd
z2570f1c7b0bb7340301bdcf3e90f927ed8ef5a4b167f1db22e8be4fe58f8ae30e932a0060cae6a
zb55b463c0185ed55ab1e677421648bf88867eccb71c7117ef77ff2a523064c88cfa59e38832a1a
za8b3f19666933f57b2d88ddf7630c2187ff6344bdb1496ebcc1658336c1f8e9e6933ea0a73b476
z92aa84a0b89f0926197f0ce488261e97a1e053a63f94ad71d7495534260e57a3e5af1a705d54ff
z6db5002295c9857328245c399264c33b659ded4bbf8d46f5c77c1d8242edf547e8c84c353f77af
zca02746bcbbb12ada559c546c51d5304c81f7af3293353f340542610cd7714c0b69c6eb2d6ba27
zb2ebd8463bded63eebc7883ce3ed99e8c61629e964ccf995cab32bfd27435098fc463cfdee2d62
z951c1ed892bfb4ee8056d073ff54da75bbbbaa70f10dcda7ad82b1089f218608c02f3cd921f8e7
z9dc2433f43d7acdd43f5ddf556b1455a330089e5303fd5673ee289313ae8f8d0fd1ad56948bc9b
zda06822f1add24f89b2181528a8b36534dc1b712ce13af29968c4dfe9ad234613744d18662d263
zdbceae291c847aeeca71dd72fd03d87fc82cd90674150752c2bd21c6a9064151e196f98a445d8d
z53dec18c9cdbd8c803c44d0ad5be0d2075c835483cc4a934fabce630a5a3c30b5b016a024ece48
za43c6318183621434dbff254c84d53afe9e3d39115930925c4942dee1d4a1f0660a290e0843a89
z014c3247020ca96082529d43bca4c515655f5b8f1506efc6a294fd57b94d0bfb99008d0bee6e0c
z78ccc3f1235b033fc9611d2f5956a7de3031da227a4ce54ef94f986aec0b1ecdbe41eeed113b13
z93b8f726b7e4b1c801fc39798457347202ce706234c060e35e972d2441b83f3b08c4f86efc969e
z750739863ca7ed904c1b727a03998031f0ceb8f70ca7086d6260a01af69d5a0ec6ce8aff025319
z6526e407dca031637d8b8520709fb950703de5a57e5431a362e9bcdd3bb286e834fb307ef6476b
zff4b117eb65841c536b1baa63d26c15fe7bf36137e7a262f960810263205a8b5db2c0f310ec579
zc8a32fd362771194607155c9b9eb4f2839ed95ed6da89fcbbb2e429158fbd21e9776f0dc050dac
z5a3fc2f33329a63ca64afe99eb7d559b58f4e1abdea4ebbe2185da737a5839df83355dfc505bbc
zfe61e883788f45c411d38da985dd4256d5208e8c1bf8dcfb421f4fae07bd76d6b6fbabe89f146f
zcfcf271967db26a890d9c6cb12049531fa0276fa03249b13d763c0acdafe33366da3050695e42e
zfda49c7d712ee0197aca4b03cdfa6f5f20f269e7d04d470c73e3fcee6260b4180f6fed150c6b55
zec96007c107a2676b64e3563c4a30d34e4c327fb6b43fca18991d046f6cd92e98933039bcdf252
ze80d396fb1f74f654e12d8c33df5d11faf3c8e5bd67f87643a732ed91659d6bf830fa495d1083a
z30d9444234df6a8f42af45a7e13405ec3b8484b4546252f25d30d9ee7f393334e30b49aed383bc
z25c108418bcc0e5b0e110355b0b74ac10b7bfae4407c710bb49412cb89ae962ffa5367c7e4a176
za10760efdb0ac169dd3be3d9c58ebad40382d1a6ca4d70a4d6160c2034dc9638e6ea5a0b25928b
z449933846a6b5e9b508040c60d403eeffc7a8012cfc8c06d079ed1ea5ef4949cdb8a34255d36f7
zc67cb2bbf1d8476e306e75db198a2e4151c903ac6426b47816ce3604396e7bbbfecc51e9b76117
z98d4e3d41249539d1858a5a099a56876b5f42cd14c68334c2424cb25fe7ba6bfd274b897657275
ze5ea741da36bc58115acc8db5cbc3f84c5f40e1da34245c398d52ed87d06a180b38c7c22cf5cc8
zdb7d3dacc03badb71173bc55c1c5e3f8359ad913b772201b2f91cf749e167ead370c7f6191dc55
z094c336da37e23322ec12a8e953c6795a639b3755c75359601e0600835d8b06bf64f8a072d37fe
z9bf7c6a30a49355396968db8195a64bdbbbf386ceef082f27ba0cf4f5d26126befa32f354063a9
zcf18d8d31fb36305d9ac5ef8486c33ad7c08e5badc0466ce1c3b2b17973babeacc5309262efc15
z8add64ba67dbee4e7df045056301cbdc6b90a6770b0aec8f9bfae51c674131c2e84c7951b33bc3
z7d97b0bbf83aa42803177ab5bb0b213a5d7489882e230720bba9b004339590454d8aa460894308
z8bff00b8caf302cb313455489245b938a726654b055f8defd27c531f466149fb25a0eb9526501d
z468b675054fdb7f88f9f46aa2ea6916f22b01f0e3acff5cc0f69290e373950bb7cbcc06d226014
z2df8a7f295914b353bdc49c25f941ccd33bd5a26c27b156f0cc6757ffd01801cebaf9ee746a137
z3e522009a9e3ee07f6fbea6d4bbab9b156aba88ce7c1acb4b510e22c0c8e58b4d654c40612637c
z387d5f99d78be0d1757dc6d8fd43604df6c3f0803d51b5fbc019f86cb3bae51d452098b2e2a271
z002313f4e036a45956f29bd696e657420dcab5c9bf9df2c9465dd2a31888f2471e74fd21b01038
zeae909d34879347482815941149ee0352d64e2d371481bf9517ada4490497cb46f5adf9844ece8
ze92e1e807f18cf87192575c461a2ae8f1e76f73d6e62e56554a8a8114d756ba41912dbae4acbb4
z6681f054bd972882530d901a62eb55b250110e02b501ffe4b62ac5589f919571caba39aa58b859
z89bb953809ccdba788f21de52ec8477dbe00421c09fa87d6e481c704e1b490d08488415662aa05
z340e8188a2ed9c8a36b12ae665b0ef24cc791e4f6f36e254490a4eb9be88042f093c74a8a761c5
z082432692f931c7fceb5bda7042298f891cbd4ab8ed563d7ba044b96c7c3cd0f60acad994ff733
zd37499140648931a93a114d995b82717c9686f7bb2aa4aea7f66d3dfebff7979278ad66a012429
z0b6a3f50bbad37a59c3a2ed64d641007b52b64f821703d8fb05832950b1919dd5ad306764d4595
z755d877f8d530a854b7186c96acc19e1cb499c301ddc9a53541c6f6905fbed1f4be1e0339c14a8
z1ae18b7b0155c8cad964e1fc49cdacc80eebb88d14ceeaa1aa8cf390c7c6e883961659d21ae1f8
z75c1b6397d0085df76065adde080b26742ee2426e0abddbdfa12781ced2cefe69c261c93091560
z2d668784ef0b797c2cb4c155d8320608efa10ce2d6350f852595da3cf5f4bc0c06b7d011567c0d
zc76f0149096a252e84bfb3bccd8be7d68aa4d4426a2ad8a9ee2657f344975e1517b7b4ae2b519f
zdbb3424accbbbcb802ab33dd8703f5fefd4afbc555c970d6c5d582fa758646e39a1431a4bdb758
z90ce934e0cd343abb48e8d5b0e9451352676b0aabe2f52e58b65e9da8423df6f84663a333ee2d7
z1e63a95cced2e9ffec73deceb02f7efeacbf9d7764c135bc9b5fe706327d2b35e09543f42f2100
z67cfed5c7d1f0ec32dc5eb2e1792aaec575c1de3a45b7da42d0e187d37bff563e536750d88b31e
z0a1960a5922c90324f3d6d4286ae48374886e10d2e3f1ef1c084429b23d2979fbacea65f7d51f7
z119576e31acf7e4cbf51eae9230c46533e8fbf970bb3ca5e40373c279c2962f758390bc7cf376a
z32916351fdf369fa4426f7077ac2a2c598dca672501d928ccdd0363770d4d2178e497fd5308be5
z37afa55745a0ff2324ef6da10adb0b41caf353b0cb7fdf398cdf8fc3ab8e560951a9490ca08518
z2614ff4d53dfba1885006822fc6d497445cc67f13ef4501132174213af699617334f28078662fd
z7596515814fd9a8da0b5fc1542c4e88d3670d1e9619584279dc21c30807ddd15d70dfcdd73b2b0
z151724d6d574fc007f6653b45a6b89f97dc0e97c1f143206c293a9455f1f4e0e74be2add1c183d
z9df1304e673010d27b6516161dc10cb7efb23b68bbc1c69a9ba7c59600203690cbd79182f8ea03
z69c677b30c703f750e2d3b9b6b4e8f4be74016c1d70a30ba938fb32a6c5d163e283966b8766707
zcea3d2d8b2836817399ae2ad4805cfcad326dbdf30da019857265bf60cd086c6ce97f0574e7453
zc4214312f3bd3e7b6b5762e8fa0aab768bced732b0d81d0b84a23b4823a82e65c7a04ee1a72e2c
zac45e753d97e4bacc44dec26ef4907a5938fbf84cc4c5503cf5188eacd96b77c777bb64b54ef8f
zf4265abfa01d7b03d81bd70b5e5c809cad9a4e52eee90e3b35332d9928a21c0be574036bff2e55
zdce7db3b2a93598679c2dcc8fe3f5a761081def50db4bf3d3a501dbf8f9ec58b77d2e0c921a1af
z9a3b843a15f117dfce0f708cf0c8b4cd1517fa388e1a2ea357f1cebbb932a25c45dcf5e831a7d4
z429e52988df64bd9c4007d981722d297b0ba87c96dfb8d1e19af5e7879ecf40bc37be2341d9dd5
z7d619aa1f89253cefb4a99376f6fd367a926eef9b17046873282087df259957371a7c0bb9c3451
z51a9cab46ebf2d1d195da457401beb8b2f6a93dab86dc0377fe830217e462e51edd1b83ed2f80a
z5cf964b74a77d047ec0d81220c2db3df2c3420cef284c6114a0fae48632dc56a742c4d5b409d7d
z906f9f41ebaa34fe2f02a1cb7344ca94d27ee1570c5f8c7f0255492a5c6de5f90381f8f228df88
zb0a7e4200c342771c3cd7561bd02f4895a4255665fe7904ff0898e9913a24b6c68662c28e265bd
zd8826f38c82a98d7cb28aad56b8a85063a5c3d5fb435cbb16a62a6dd1d657b4425a49da5210c85
z724cf9b05f51e9ea039871dce60ce250179879d8fb3634b62e797d69a0418bb77e50bc13f0910e
ze2928dabc55fba5a4e9957fec789b4fb88230ce67f3046d704329246749077243da75e87c77dfe
zb876fb48f39f0a6e88719bfa054c72d17c71f1650a1c02cb887a1aadf8cab5f2d276cded891d13
z6db34081227d86855977babc99d07e8c1a0a15ca038775fe330782e4a7c496b6dde1afd363921e
z9c9ae59a3a2a6c0311c82ccff3442c6770e7ad7af05d47c01f5e04a08bfe50bd68aa5a77097cc3
z39b2c8ea4d17ef97c28551d9b1592b251dc6d2e2e26d3e70c74c42f0b93cffd0551b0681cfe96b
z8458303af42ed90565c72ee6f8a3ec6e8bcad0c780effd47d64ed37680c87a726d3b50b8d6e2ed
zf2ba6aa4b3b0fc609fc42728105515ee591f127270c157b00c9a2a28de36066a107bc83379ed17
z25eb1439311985d70f56a01bbe4b8ad24c212b18e4b8012680d4ce3a81215e550ad8ad4fca24ff
z2c30683ee9b4b43b584452515ff88019597d458ad0d980a451007906c796b5e1d7bf55a4ede856
ze44244f06a1a918182070e3bd10128a1a937dd28ead67a0285358dfe1c7866e1864ea655d55eca
z5bd71ce0327765c8ba63d39186cebb82b51c71ae705f524cdca18222043e7e404b2cc31992794c
z9b854ecffefa068ad87cb82af18f7acfe678455fdf062030bf761b30486ecbc48ab0029282cbe5
z84f5d1c066a579703041421b12c8efd4d7a35400be12b24e2786709ce2a60616cbb6d76fa679d4
ze82acda90a42da36a7b326d53f1bd850808e98b3a7991c90de61e63aba96210bfb4370a715dfda
z82c8487650584d83a488bc51641ba514274d7fb60fdf3b96efe92f7ba120797c5fcce95a33f37e
z7f179759b1b48c9873a4cf90a0cee93b69360b31ea72265ba1b30ef70ad976bba500b3d63d1d65
za65f0b252bf060c91177ca43eae091c2052008370fbd00d8d934aabc121f9269886b37f5f472ee
z8ed89b917953a0ed647862f560c65742cedf8f63bf713e804d36133c2df9a94ea3798ed22203d2
z94bd92a1db13e60a0c286a8f65041e0e7c96be7f40568fe9f3dac2b831b7bb07038f7fd29324b2
za661c593db7655684faca12022cd819be26f4c2838e3f6da78d3c5a5c1bf63092ffeaa8d0ae432
zd48b9691a7e73acea44cb426e730991d8f62f04ab93b13dbbde93aaf3a8ddb0b0f86a5f2895ae7
z0b5c82e7fd733c8401ef0bf13c8865c578fbbf2b589923a2180bd30c69f568637e31a3f32d8008
z643ad636bd1bea83dbd766b9c521c0686a0eef14d780fd9ac88111dd0f73199006ddeac9d80e66
z50d70d2b411cdfdfb5df9cbb4872715dcda73dea54caf1e5ae574f0137dba2669b58ebadce0f66
z7b5671d1ec59ffc74a07ca34fa856acb4cb51242c52774a1f946efc9ff5a1a8031797e494753c1
z52f2aba687e098fa3e0ec185e6ffd07c590dab6cba15c1a22b37a9cea4b4aa28ba6530e349739c
z5b9745bd7a964a062632791ce4b1218886d8b3252970e958574f196db42c08d60b367eee9d70b7
z566e956c85475f43ea6e88dcc07bc0e7069034aac19f1b913a51f83ca350cbb67f1d3ec2d592a3
zf4a7e79fee81fac4457bb7b075c16dad6c48e6ab5c5bdffe2c3684cf0f22a6c55bb600094faa11
z7f269e888f155ad8d915232c3e6529bfcd679a8d6fd2153d1e207cf2af67f4723325972d42de71
z5714e6db1c3518d290894fc8f4f153835904edf396207e17fe918ecd352fd09fac40d75329acea
z257c0061d15363136b977d1456cb9ae00696fc5dfbeecf9b89578e0ef15108a58064ad5dce9aa6
z01b57c05dc916df1613a627468d25e7f381035626cd3c920170d2a3e7fb3bd3e5147c0b9f7bebf
zb3510f93ab370a8b4c52e80506547def10d829f788ac11841152d6c195af7f11afd841973d36b7
z61935032634aea00acf6a47ee4acc5973940a4b572b2461ff8cd69959a6dc02419533f5e80b94b
ze5dd1a22d0c79433aa35b328136c6e7f904f518bd9c5cdddbcdcb2e451556a77c6e16d57048289
z6ef59965ab7c0cfdbe932cec7a2522284f291a31ea4de4f28fec3c6a432b73c114c32691362005
z9fdaf8651fcb598c79778db2ec154a6cdec2202f4ec142a8a4a6ed7d4ff9289504f423807aff62
z03d6b8e9fc1aeb1f46d3d0be84d4418209052206cb440c92f6d1551e174a2450103029de73d76b
z6971d38108eca6451cf9b7906025311f08f77f9f5277e3b1da525e6d0c3d61ff48258b8db09d7b
za07288a5f5079fb5ab89fe52a1ed77f6536f7991742eddc57875047316e2ea5147974168af0228
z10a10843e375fb86bebc98e82622ce975b567dbf8ca8c824c899a183809e2c090a3b805ee4c639
z4f65b4b839f769fa136df5b3068573769240097e3e50cb269e1a52db34e36ae3c4af8bc875e818
zc9ac95a998dcab5fd91a5196348feed79223dda431fb05a1d628e459976d9eebc6cabedc18a610
z331658bd398b2b5d3d9c1df9ebc5f119096e570814bfd5efb5036f0f51ee652e15d7cd66b2c2af
zc1562f06d38f4e8c4e56c245fbb6ca842eb5b2a9cf3c39801592e7bfd0bf01c645b5e339a5c0e0
ze03eda7f1f6bf46c4d57a6c1a76fecf06f65efc0a86916722ee3e140dbf4e8415dbac907226f6c
z0c82debc46c81ac44bf3002671f92e64c64ae0bb0459f449e9f42c6f082cc3982e1f393c205424
z2ce6cf920c9854fd28d0ab23c4125aab01ebd63fcf5c2de3659622083e435fc18d5bd70be66156
z6c5d057e89da76b351399bf80071e806f9c3389323d687847deeaf1623b675a8e8ea5c27f00f36
z99d0f7d471c5429ea3be83635eb0beabc65c8e84c5933dbee4662982edcce4740455737b674cb2
zc0887a8f1dfe892f2b027e367c940b94553e2ec77f514ef0eb0606b02cafcf6c409f4d28062960
z5e6ed4f23dbf8c0bba690541f28fdfbbeddbcb4644eb67a6915314ab637854326967be723c99aa
z729b780ba500b92e6185eb7d8131bb88ed00dc69e7092693f4bc52d9490397e9614157c9b51cfd
z490da557e51eda81915355e73904f03858289aeaba38bbc8deb8dbcae6f79bf71713fff0d778a1
z3f3cbf2978b8109ffcc701a52c7cdfa6c5e511983e152a32f26ac26bd1d8203be9232318f6c4ce
z741386cc85b4d13665d3cb41e89d6a5b4fd5218a1bb24aad82eb9d44f4137ee1b0677c000d3e9f
z8f8891e0e2e38f77f8b88ed40056b28094014be4c79d6f69e8181c93cfa81bcd6af44a94afa66c
zedb872c92f367b6c2aa45766c5c8ede6ac34b1b0e25f7bfadc267c3937b34d1cd9c0c2e11ea51b
zd663026a89f29b0a865584c8a021c6f8969ffe2905016d463d29e5d4bc5de111a382c67b20dbe9
z3f1ef8c22e640b2ab68d1784e7cba2608fc5641e17f4aafa24564565880cd1158d9baa5bcae814
z721d93d78986a33b511de4dc591283f5e9ffb2ec658f33440c5cc3ea18a46d4da340352a588a15
z8433dc04df918b7e64d2df1ecf11b72d95c4d36999e0b44e453ef2ccfe1103da39f3175ae1d81d
z506ba900584e430045ac2e33f17c1320b2f92625c55826f7667eb2dd8dd74e5a4968171cf125b8
z28d530441a1252d5020d31a5307eceea6846988d1c7cb3064564a90162097df8e8bf7820f16a7b
z6ca5fbced832db5a4b84fa3b0f9aebbf4c1e64366e31d6d13970fb822660ffdd78504e084236e6
zdc2bab6bd58cf6d0b218ea66fd46d046a2c53802f30fca90b3a02984d757f14594c5e0fd03822a
z2f196939ca2fe89ca8fd3f2c8ee6d64ab0347dda11b6f4be930332b429fb21eb3a0b26dbff8d2f
z98bee7ae2b8a5a27ee62cfb8dc4a561098e32291ac8d3386892ab5506305e26330fa126bf93948
z7426b934a6c4b78a45fb4dc8dd09f2ccda5c6f0487b29281c925ab84b6d97c183745c8f56a0b01
z395b8bd86f443999bde82b819e9447a502c4d947b9d8c3ab50aaaa7551fd043014089b85eec0b8
z4948bf523f807550ca5a5d06c8a1d8fda34c53db39c1be25dd21e5eb5a2ee52db4a5bd14b4e674
z2dddbcc76acf77dd917d46ff5a9a5d9ccf1cfb2d09a7d5a2d10f7aa422582a25b232727a9515d0
za0a2bca559530b8e8212749883f991950e83da57d40105792a7da5a08989eabe505349ca211365
z36e1f101d27cb4942f2d1e9cb3b725f88895810473507de8db0aeb5b9df6c2e34fbce944ce43c3
z63bc015572c23a865987e64fe7e4c432ada9382f1686dc62263b63c1cf626a2f3d74f7daec7ac4
z5c845b63b21bab6ad68300385fb6ee5868b90cc7a8a97480b828a5a7d9bdc8648509f1205d1970
zb164009b60a20c2f976ac5ff03a2e081f26a903994f8d9ad21ea7a349ef00407b8cc8bf9850e2f
z68c70ddfff5795caaaf515f026f83e4d5c0246bba884ca641231490e7156dac2b0066d606198c5
z44b28ad3b6e8fd907dd91ec6d71caeb1ce1c60449b627f5c49d02f505c32355bae704a8ed4ec38
z69e713375d944bc8f8914472b745fe90726ded1ce1a3b5293d8b42f8780673fbccf5c524f6c3c8
z3fb4a8938590cf0dc1d09f471a9d8e65cb38b72a7464dc2ef049763c4639e57affc0cb79033422
z44dd6f0239667c59180707ecc6eb8ae6cdba6b0cbbd57503bda999933bb15de5ea045deba8c543
z39d733e1872c3f4737440c999c317df9d1605f194d9e04a7b803304de17a0ce3d3ed8f4afc1edb
z77646cad4ff81dc8385daf11703fa1ec7ba6d28f0ad4d6713fc8391a26940f5be5bf103fd70a48
z73db6f3b9f759aed142470d64a7a71a46603bfa91f09f30b40660c8dd492dae8f91388e07c4d0c
z8facc778d3cebeefa453272918ec2d5ed8c7be29771b63181d08ea84618872b97af55ab42022ae
z21f51fb525f68c3ae7fcea0463b959a50482b9c945b2350bf2b87f7b46af2f9c0f0f99eac53048
za0fcd2730e7b3ed5fdb18d50f6706e8b278de0d320a715ca640be9a5433011cefbd529c7d4ffad
zad511661e9498184e3fd75ff3557afe969a2e4754e533be8a8756695599d80cb94767c9cf2c818
z93319a0fe05e6505f9e53b9b98da181ef88c64eb7d8eaab51964e477e8c239618acdafe548989c
zb8733417a1e523eab6ad3638542397ff7b8e99be921df8899ca6228de3c30a4bffa3ee4fe66617
zc866cf3afc68398906d0fd856d38e84829ad27778aaac7e2d085c6c7ee6bd45ae29c50018fc426
z1e736c4d1993215669472e21ab32bf157de8d0de229b3b3ee32b55104679611d81639959195fec
zc5ea1a724b4f5eb8233a70f5f99debe3d54f477dbdb76525c7bb21a95d4dac21d7b143a1d60bdb
z34ff08eb4a5885d9a485830dffee443226b5f53e7b08bac7de6e8820a53a55a5f9dfa02bf22b81
z77d0ae495f488921c190104f7d1a3b90f147f53b35b2016cf7ae9acc7d170682f67efe9b9cc829
zcbdee9cf3bd7775d23cd265d23c646de546a4822b214c5adfef07f542c5832d064d7aea76d2603
z9bed274fb6c398c657eae503f8e3991fc5ce7e4343c107203d7bc04d34b42845b57edcb94c653f
z25c1332b9211a618e3a16b3b8debbda6b5be738b8a97b44a8aa3a2a8cd503f27f356be17b2b653
z5062a55501219cddf54cefce35f241a61fea3e7c4c679cde458a4ce445b1bd2e0c36dd496e1746
z6db5001db411aa08cb4997179a944e0ae8be4441a6f2ef996055928b9389098b2059c956b40086
z134e062c202319fa1c48e17467e0e09b4c2d2d542967ffb63741dda8d3e25dcfdba39c7fdcabd2
zb8996bec9850e7f6770b712f484277155e64056e3bc3ded8703997c7c51011a8820a528f66baab
zb372b089f6ee640f68eb355050608b280ffbc1cc64a5a601be7a1713543e4c840d4478a84328ce
z9c60bd397378145f946a8b4a2f69b41f4ef8e183b6858f8b2f8193ad7daca2939aabd954f3d231
z78f24a466310503799d581fb3cb40e1916fa965e4b2442a10158b8091d740249e5678d572f796a
z603d75df0ae82e26f734fdf6317f41a699b990f3c0e24a8d4dd5571767eee71da622204cc48a21
z0aa7d23c7b913498873bfc184390522fc4deb1e2417c799164dedbdf8100ce1b1cc32f9f5b4a30
z4d6b71360a6585f0a83d79fd531547f51038c38e63cebb8e6041b37dd7d92736592cf4cb0c15f7
z03bd033b90dfcd3bcc55498464b2efbd8687050c6f2762e4293523f95ddcd6a2e4752aa456fa19
z213dcdfbd27960c37a31579ad42cfaba6a8c232bbb2a9c46c404b04bda5dbbc64a757d80dba736
z4425b9932dfd30f5c8ea7636603a199f9471da2ef0f10036d017d978aba236712a233740bbe3cd
z7b9da928da846a0e0aa3c10f731371a99fd6be5209449ca7c715ee5ea1341dc3ec3561cf4c4056
z7ad274d29071b697b5ddae13f3ca9109248b2e824cef6c5e81498b47845b832b3a0086dabb2dd3
z1d2f52f4fbfffecda05b5b9805e53d1eb4028ac233771dd144029e70bcbd80db7b7f9c130de361
z4649fd721ba4099d75469146ecbcd4509b2272438a7a983f868b6f3d251e78891542ec75b350db
z87eb8e7df084299956f341c422ae3dd013a83b69e1e3fb2703c4fb78a9d76400c7478ce309d213
zce1e70bd6ca838c43f6c7cb6b7bb7028ce654228ee3ff264905cce2ca7c85d89cf55bc52cc9f67
z888011655446de2898b15468d4c8e5b0a0f1e8a5110d44a157f913d545b779b80ca70b4b87b534
zf173f41834842a5936af67e3e9cdc896e034c58c174d1b989f7aa0cc9466756ac0596a8663b901
z5f921620d07fe6cd6db997e6c0f59855ab9ddac42e8ef6320a33288d5eaff154a345d140c0fa99
zf1fdfcc3037b2b5b3b5ec6df1c79ffebf1d5fdd4658de4ba1f317d0e201b6da6285ed1cf3365c7
za876dbada71e790df098cc29947308e69d90fd540e7c663322df644bd3b7bd3a9966e882577156
zc338b241b7c05456b2f5a8a2b9437a738b725730767887e1daab469202499064fcb471a58b2661
zbdefec9b4ad7238cfecfec07a4d4b2c00c66536783f4e4a0209ebab4c1740364aada2bc20f43fd
z767e7121bd8b3ac746715a0e0a154863cd6b666e6bf2454b645503aa4e5953133f9cc2c307311f
z6ed251477054676832e741ac96fe637538fd44e18c75a689e3a41492ebed66b750a2ebd99afa34
z1b269945cb8196503e76784b25c88041f8e4e6f693136434eb7dea2cd1e6cf6c894bcf8f598eea
z302195835f0a4c7ebef1212b0bfda45209b3657175d308fbc04d8446bca3417cfcd341ffd1b616
z7b1dc9492a1e628c6386c2b9d4f68c8c8370bc6acd928b019218ae8eb3751a251b9c83627a17b9
z46e6cd84efbb097b5d3bfd5ec9cb2c906fb9b403fe7572cc30b7931bfdd90e377bfbc0489eb1ad
zb794f1c5c97b14434adb0053703a38cd6b0d3cc04ca7ea09c2c815b055484acc0cd36bb6d59346
z7a26ff14af172493e2317f11b6cccd1adb4e1d8e71e310ebf25799940ff779b2fbc1a8ac986318
zedebc3cb232d518f1d8a8b36da7e84a49e46c0feae8c45f76ab3ae35743d8f6d810226aebb5ca4
za7418a5e11ed8099bee3b8556f91153027377f5bf936d05527f93a7ac37941a267c8c61162b592
z576e3b422ce27d5aadb9dc58fb51e34c9e53a565e8b7c360828ea55ac9a58eb4f1b269c218e18b
zd980cd8a329db477af7db541915910ff8f690a6ef0fa24b5d7de12c1e36591544718798bb64cb9
z78b68d317f7ec5da7cc08f60006718d5c2b1cf9ffca9ea826ec0035dbb448a55ad047bc865527b
za1571e9129f11add9baf9ff3109f3c26ed5509af95f91f4fde43e2725dbe4cc721e48ab6a2f28c
z5e41cb5487710a835451e1b66d30908ffb9a28acbea197babadafe0799f66fbad8de12ce8949ff
z8f719844e2a409a07ed2b4935cee0de9231de06c67711428088981dd1fecf13f66f84731e99ba2
zf0d2f5397c6a8b0e009b73cc4a7801afe6fc8d1579662b799cca8fafbf665a1b3fd079a4bf886b
z43772e919a2acc58dc5b782d099b89ebc61d4eedbe543087fbf05f89811fcd381e4c25d46a5572
zf6ddfffa355414964185ec14d9d642b5c5eaada04058f16044fd0063fc65ca9950da8b22e8eea1
z10de1b4dad279b16c17fce6e74c9ef5b612faf47d59f3cfcdeec438a7f8f8910b956ef642f3ea3
zad689c82313ae5062fd046667ce7cbd67ace79f517aa277a727b08e029f00819ae4d6c0ddaf7ee
z53e1fb7d8d309acd1492561b265c2ccdf108c3508d83a1c196aaa39c75e10bf7ab90483368ac92
z7b1f3d6a760f3d37b40ab8b8c679dd9c3fc29b3b0b3d4be6bd95a0646e0ef4f3353e8cefc6a19a
zbbb87623465b4ce8e6fbc58c2847ce
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gigabit_ethernet_mii_link_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
