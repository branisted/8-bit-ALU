`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026201628cee5aae21fb892db766c4
zb5b1406e11aebfd6dfacc9da5ec03b70c276807a3eb15e28ec7ab1dddec42388b9424ea285623a
z248195c9f894b36317ca6e59c86f11031163f5f52d70922c037057ec65cf19cac58583b899d7e9
z5b165e80500bb14e47281dc3000df4f603e04a7828f6f0c74040d85c3c8ad036ef3bc1d66e3047
zcc69669174088ed23fe12190fcd63a31f35be060169ddeeba175f1a5c995cda14b83af0343baba
z3832b130fb9637d9da3492922c2a4f84c29b9c7a7bef95fac170307e5a87742cbde29d7e63d44a
z1ea2c32c161ee16971df5a176e10341b9071ea4477f60571cc3cffa95a787c8a550e8d32123773
zaed307dc63446b99b9a5f2b8ef593d323ec52af399ccbf7c699195a21573fab1e72ece05f53f24
zc0520b074b04c8b288e35c02c47a9f656b81224cedd0f8f2d79ebb9426303327f83ad71a9e5103
zcac99705cff89a76886ae658df437b82d4741125592642ab86d3b0cddbb81d698d2333951f1849
za8290cdfbef3db1ef9af7aafc890ecb5b4c7d4db1d98742c40cb5db3c2fcdb96c8b065a184427b
zdf066098df5235aec4bc777ad4883836ccbe62f4323aee1deb221ccb29e4a73005beb54f670f7f
z7ae73d8567352a488d47847415023a4339d7fb4a6afdff6230f9cc276ce1220d66fa7ee7d86055
z81de5c48f000511d81dd8d57a390a03cc2cba1961a7a8406296c57caa743dc542a6fa94df843bd
z05beeae15b1affeaaa23c9e79db0d9ce00b04f8a41da6666c51f2691f3fcc006d01117f314b0f5
z27d57795aa56df23eb5ab405ddaaa177b055b4b42f372c6c8949236b54d3ac3db45f4a45fd3dde
zc6895df7c034bf6e2b4a246c10331e286249031031b368483386fd209c2cc1d88b342f9bb738ac
z99bb8837c7639f5000051943ec4fddcdb70c0e50e86e3e6912b5b0453542bb67191754ca81b5df
z04a227aaff2fa46dd21ca8f7b814075947f684efd04404da5fb0fa9661fde5d31a8c7aff2950d9
za6bcbf246ce5cc9aa8eaea8f31e7b08e1d8d2f4929ec41a63d01ca828199b993ad4e9b6a205eaa
z8e4a0fde6f5469b630751747476a3b4d14ac27960771d084ccb29d4426f49f5c1a4d98e255b89b
z69d8c58885e2457aee4faff724d219a3a13f1cb6c59fa44592926e9e624ef6a68a2bdc71a55648
z7b4b585e317ed39b120451bae53dc77dd583558fe0018b594f52d20815cda5742134adbb422c63
z074455135f9f87a0a44cb830c782e157ee09436ab719adf855ad962af3efa24b222c4dd53c593f
zc568d2fe4a439d07d6b5ded8266de49d4547da55f90a85bc2adb30dc35bc78c57b4075a899b43d
z936e68ba90be82441a84e7c2b0043146b79ddf366366b254115cf0f30f7299086746c3c8e02468
zc9b9c265eb8d4d065d9d577e7e2b1559f92d73df021fcb80c85e1d6436ecbcc2af04ace8ad91e1
zf1368aada7bcd4c589832bbdc0ecc110a5a77671c31494f06da4020a4218ccbe9018bea295cf56
z1800352905a8581bd711e97b3b44982072d2145c0fc87a8bacf009562d918f91c2739f9ee191d6
zeb82d4c7e7aaddff1d355b07522e9fd623125be4a0e5b1996a346ffd3fbc76902cecb011cc0807
zae314c28ff1f5127847bcc022bc6b99dbb03c0d5e477f2f9abec33c07cb8a8728dc3f49fb79689
z2a69c9fccde9e30998a23f9a565f366e2f5c151e8e273b9375e30be9885ccb82c47afd55f4f61e
za49f47072075299f29e05ca05dfa884276df68eda53e96fcc7094fb5e756bf57117616b47c88dc
z9be5c56d0ad615a3ea5fdf22a3d713c9c6a2cab4a71c3878a64835bddffb665dd8206d24725a62
zfce3ffa5670b4934e7fec0d6b6dbd17a445cc0823d5982b1d340e7b24af4528f636be8578d9f0e
z24747c3399bdec6bfef9e15d7918c3d28b8f08847c4da57030d05394dcd18cdc4497aab8ef257b
z296fcce08dd8ed47acf458a79bf19817fa9c17453c6b884eaf1cd43852c8a94f5c61e05fc93580
zbb1d8feedc18abcf34a46198c8af355c02a4b55e5ff1ea4e6802e36958aa832f2c42711a4d5226
z7fd5d5061b005260239f006efeb7e2f0d9f536567e8fdbf788c56062ea1684b95762d4f4ac59b7
z5cb4416344b6d6210cd8a422702cc64c38653cf0a6ca3511728b45969a7759714cc8685c96708a
z74774bcdf739fdb024dc79dc00f8be5d85f5c625851cddea06326a52fa278c60b0dcbbba36d5c7
zcfc673b0f81b0fdff9b07e44a58486f7ff3a27aa48badb38afab4eece605b65f796083082ef3dd
z4d5a95b37c866739b363ebb7728f055f8e59cbd518b2e75e18fdfe23775d5dc5ae586a33f71b39
zdaf58aa153589fec064ba7e4fac73b555ea4a4da1d89e0125ba7bd5982940404999290932b90fa
zac079d8f1dd6549d61cc4efd7c834c4dfe77ae6454f5e80bc40d31103d7a36be7536196af76b7a
z0012eb1c69c2fb6981c3e948eaa1bea89fc0c5b7e35998a23632ae82aaffba0c25c50d8bef9df1
z772dceffa0f81de2b934df2eb0d365c4a47fd31cfd3ec0f7fd1eb5eb82fc8c76481c33266a0025
zec5871d60de78a5d473d80d58d54be69a7900eb37865198e34a8ca15cf37bdf2e454c9a9977f27
z5f45b2758b215dd9ff17b57fcd8b929f06263cdd399c62c6e82cc6ac39aa23547300506d96b970
za2779865cd62581006c89a25810b056b91457f8e94b62a762ceead4ccece2c3fd403c5d46ab36c
za50cf7d6e1901dbf21bcd17782f94c9b286850964b9f13c73dced4ee194f2592e03b5c43569ed5
z322177a5b21526fa444bb2c704383934c3ea34e802adeda09d8ce70ad69f47701e7bcc3ec36172
zb2225ad230b2fc8e5e2dc5f355b4ef88e3926e36b45d842d1481928798471e9f7e93e1dda633ac
ze12a0a85b07fd9a5ba363497226993c4ceadfb6719ce02f4bc62d2cdf65065b88ceb7257295cf2
z037ffa800eb7332adee4e9add4da0db0ea8a970245011b7b5e8ad985f3976e21d08cdc06cc777d
z9ba213268f4f7eb6229545e93bd018ffb910405e21bd68ea70ae70a023f91a3ac7355f3578dc36
zc44c29d1b955c0cbf2e78e8a39b573c3d23e12976073832a963e82ca6c009d9c54059f4e0e2925
z2bddc178b8540c1799d96889f04a2bcc76108fef713e813c577b6b687cd762042c912c9912fe4c
zd9121c3114daf34b1d9c7e21f1e79b272a9f8ad7e4fcf02fe7c65ae82770104ef3064dfac9cbcc
z97f79f9e7285f25a63267252ef55f81a0722694f63c9eb6cfc6a20b594752bbc7fecc43ae3111e
z59bc959deae306c58d042f378957886d743749ae45f05b83ac53c3fef162bc28dcd4b3ef3976eb
z041cafbc8331008295d545cb82f5d01f5d71fa7ca3c9d134de298ce019d4f218fdd9f603b053f0
zec3f0eb309520142cec31cf1d293e0112b44f9d25ff243c7bea34bc388ac51d2b40a14a7900599
za2033d1b5941943d7f8319ab6df5d4930ade7b545f4369c8955835e353e52e4aafe8996d71a32d
zc56e4798eaf823cb783bc314442dfc10bf90d567770b929fa4c1385ba7b0bbe247491b7799d10e
zbd536aec529d71b9c54114680879b89cfeabe901c9acd9fda1d7d15997f21286b1eb6635a90d84
z1dcfafc6e8a3dcf53a2b4c23426f600e972f485c88ecf8f9bc3a7478f1d3604ac8e77710a8ccea
zb166f9d72396bb54724335bc0ec3addfe417ebbb7920b71ca5f20a82589a0bdfd86c4c81cb1c28
zd02fd734e5cf9add8ddcab2b1f85f2d83519aa3e60cc22a8d2ed3901f74ea245e200e58879cee6
z6d62d9033af0907d8b5220ffa175216e8a97f1beef5613deeda6b54c70391da772a0b8cd056990
z57323eaecf0d33b33acd404461559e89166408cb6816482571ea0240e8bba810adf20fefd5f6d6
za4a8b74e2ec88bf45f777bae2efa5653f196e75ca71d0b627be93090ce03e47cb72f2a49ad673a
zc06e398c1dd61286fc992aa91a241243d470d802a9f3305511e199708d3d30d1e13d659a164377
z3f76731a9f4bcd0f496aefe32daeb83cf91934725a884eb318dc1cfcf057175aae619b93eb0c48
zf1a774f5c404f9a31579caa368dacb48e01f216274fdce3f3d75fbc5de01a3a56b9574816825c0
z791a5b1b2e1e0cef05720a1efb28b96e4b680589dd4e1aa997d3dce7ccb36257c0a98204bf26fb
ze789bf071c5c9fd49873be1bb222fe9d15e9cb09293a4a2d34194a36520269399f720f57bc8dc3
z91bdc86def0575a9c50cb8a2be651d416371deb79f60d796e97f5695acf3aa4d4c026805a99705
zcc9730620e53a3bdb16c4543c68270aeebb2deac6f770103af16dfd4f791b09d3353f9e7805afd
z5393e212cd6073ff0ca71db3cb0e59e845b38728f9aa6db56dc6aaa31fb0988837bec800aa57ea
z4b5af65603a2985de0ef9f00c2d77d0f97807b1a6904bb37ef5e6af25e45c663fb22e8a49cb714
z41f99efc850faed91fa37169a9ff264f6d0a078f78a02e023c37cfc6277bcb016ce85749095f4c
ze41718c2e9b6106c640b71764de841d5757e2e2ee3888db4acbff24748f0470ecfeec912c3b348
zc27e21e59f41f55c6df8d2f339e36f7761112409fe5a5c6532a2b7ac5322a1757729808ac8cd24
z399b896d81b19ab16b5d7579b85ce133d0aabcadf5722f1724606a5ab03a166627e3bbf13a63e0
z98674c58bd5c49aa345c5b2482ca7f9257159e8d80182d3e78b1bd30ebff496e8a4aaa34692b72
zca835fd749dfdf1e599face502ffd8908c4219bf3c1ea336dbf871fdfd14e7ac9f11b838544d0a
zded48f42206ca3207b3869bb1ca01d6f09a363503f96b2d40c152db81fcc2b5c8f7ff6380b47c2
z08c4d20eac5e551382a46b3cef6baf901720805822628f4c40ba744adce29b1a9e76ea72d0bed5
za6bccaaebf6986360986071b01117f0a8181f5b0bd9ffc82d8b86149e0898503dd9a438a1c2900
zac12b8d574d866a9be4499c541e9c1f9abbda66e30465ed47ee3162813044f4dbb89c06de2f726
z3fe163368734b406192cd7498679eaf264e6c1cab334340c0c558817720a075bfba9e604ebeef5
zdef68893f013269f00d0d3738ce9fcae1629c886b268593adf27c79a2029931be99b92abff207a
za51e34e8f74b07941452b4b0e3dbd0b75e4d898d4af9a99e17e8f9b69bac8ac3e7c2f618fac487
z45857eb3860b3b79265bc15c8825d573cbc65aea746915738f773a76e17779cba537d77becbbda
z5aad93c2820b642ea9bbb5c1c3247cd528f2702d93275123a6e094a1dc5bd8a306e71f3bcf39a7
z2030f5f1abdbd596c10eafab58146ec468ecd48c197f27d35435a9773b242b1d8b68c870451b98
z4953803ce2d35082069927c45cb272e2e6c743c7d808bdc15fc02d65c80bf220f63998b377d2eb
z6a8a816031a9a6f22863ee340b5282ecc3e3aac55f8f432b5f85f7b453d17dfd9f52a57a1e0da4
z4fd808752e71c2c9dc0cfb33c2e16c3dabdc64f186bb7968628034edfe989fbd9776513569f7c3
z9cb055c81f5b9b9bc7a9a5404c1ef069ae0b5f931609ac8189b4e900d358a4ff771a9e929d2033
zc6be18129b8e434819886f449e12ffe70d6569c64752c7869187c9ee1b5db1494fcccb6b7c0766
z2889b579ab1c8a512ae955ec8b76387b5323c5f5bf4243c7b13207acc954a8b0aa418c22ad453e
z4b98f376f5b1dcbcc18344c2e4c51c20563f2112acc876c6dab5ce6270a8f3ce9b99a246e1fe78
z4d7a7a48d3c35fe8b83ad2a002a12d29300ecf1ea60f8ffd8fa7e011433f7276fa973cee91f90e
za4179ace6bd9476f7341d2e386e90ffa86449a61d85572b5635dd10b6c7328493857aca6666080
z09523c437fb319f56a98d3eea7d1fe2cc83e1afe61be0590ef77b0ed6640e85af8b9967195bd2d
z1f870124fcfb39c3d305bd6ebc8e5bcf3b4573e8e51e3de8ec1a7ddd512e6285032d83f61f2960
z30d0368b492cd22597f4be6a67201e79d1116bf84b36caf6befb527085406690afa3dff3bb1d59
z121fa0b0b2a617cd4f5774cfbdcae2d199d7e004792ff288853b75e64d2be6aac79fef2476a61f
z5cf2b2309cd3863eabb3ed3dd5ea5c81bd3e5fadab2e456633b8f845b39bcb49747d08ba23a480
z94ba7781c155d3d0f51127423dadd8dafe3903390d74e036ec137c4b7ec8e5280107ffbfe8247b
z263b9d3e3f1f5bdddcfbb055f5ce0d2388961c3dacca7bab337a37a0a1d9c94282b980788aeedd
z95637f27473c7508608b0132e1da2ff4d0b73c62e1f1ce363a50c914b16aa5a25c515cbe3d1673
z2f54db78018dfd2fa6c7d7fcc6eff7aa725e34579922b38966472e85cc2c87a45d3de50bbd1bcb
z2f9b442d4e566ed781719dc338224613f710ee12e64b6f406af05bf2378e83e6fb681f22bf919a
z8e777a045a40cd0444cec9628b93e2cc6eb937cbe66f4678df6ff160f7ea1faeb4419da1247b08
zc950f28eddf149c7bf6394d611d3fb5b7fb50fbb181234de0a5625be6e23c247094bf6b793ce29
zc8a9b8a6e1f897f01e0f5992baa7feca51b942d5596ce1f774c397b739628dd30827a6bb167db1
zf9d7995c1a85364acb25dfcf716fe1a8f37be896e23c66c938a4f3e664408920d5f9a3d5895d7d
zd0c6ca09f0ef25bd214ba2834eaecb522ebb6b5175a56d67eaa2d9c542496b66d937b8434192d2
ze21f42d21104b34f930fe166458591540808ddc8ed0a2bdf26cd868b7101948445fc5e37082e82
z896ae6e78ab0bdc3f30c6ced4a21ae113df7c8ec99317da8f9e4dd2f1b7f483b6daae17c0caeb2
z0f7bb23908894d71d440e18c6f0b39fe873ecc806a427c6cd2e33a949dbc2b53bf36205ddab045
z20942a9e3c3f75fccbcdd2faa12483307ef2128264612ef212c4eebf393b5eaed036e7c8ac8068
zde96700cd0886a7e5715ae4311075ba455ab64b3057c929575d80dad75cbed817bebd9437d39bb
z057fc26176d1105fdc45f1fbe69c650ee5422a2b9b623fad7d227146074cf4ca88ddef9ce2a05e
zf6ee33cc69d67ac57d7c15c1d3c57e3379444a77c69f655c3eb431f7518a0fca2de7b1b1c30dd4
z7abbdb6721fbf5301511fd890a40ab4f4d1492305d094ccc91a97facd8e8522a370aa3a3b24844
z406f1200d7aeb1212cdfb54c819d1bffa8a9ac1771a464a5e06a7f59b4bfc22f73db2c9a6a8981
zd05697e674d63875216d0b60193e5d61998fd1f51470db2f6ec3fb4881a315cac08442c7fb895e
z8d8faa7c0da4a1d3e9bb9c412d8f3d895aeb07eecb80bd35e840a78be01d33033cbc9d6e28ef98
z28d1a3f3de299086bf056f0663b87ac0d7e2ae549848202565d3ae82354cbe75a9fceb2643d21c
z43ab1570515c81db5f916fc728c7e4465ce04286440f2019ed9b26168d207d5d0ad6fc63f45cde
zc2233c604803dcec032931493166f5f3fcd90b0ad37f5d4cda210d65f4011ec3ab3f0b5546e9cb
z44014e166a7bc6fdf1cc9fff883e4f5ec3c41cf627441a5099bf012e1e95fdbc9935e320790b97
zedef76d2ee572d4773f7d60a46e47e188872acd200167e6bff2554b467071d83883fb936d2f99e
z878abf01cf9a5ec5e5535a347b7242580772dcc90bb08cd02bb5cd667069c35a0361a5af2775ed
z572455ee7afcff6f98362abf4fb54eda858872398a8f2f063f0701c93dc6433ac810a14f64e8e9
z06b33ec6e533cf202fbc6890a2660d3e5e50a00c34954db7afb246b71764b7576c75c9967a54a3
z40b1cd9fe3758339a2da1a2a50ca5d1580f7cdbcde530a22670b3f96848323977ef51c8c92302f
z9bd33d3b0534f7e9f1fd5da0822cdd7cd622329a837f300c18fe723c525e92b4e20126176a94d6
z7a9f1b2b895d48d071823cfb0ca39bb73481de82e638eb1399e1b17fe5a4634b8e3ce7eb82da10
z0311a898d8d1200b04769b844e0dfb3dbaaa270ab763d876c83708d25bfa4a9d8840aff4cef459
zdcc79e65b67695dd8b3bfa43f7500de55820bb79d32fdfc0d2cfea888ee4e0fe6f5b2eedd364ed
zd02119da00b83e31c4767324bbd2970507850c21296aeffdf5816bebad643819bd1d339621e86d
z9b55b927b1263c3fd7d0e3fd120fa3e830ca79559dd8fedca32086216d45b1a074a246b9a8065d
zfb203c4c07370fbd22b796444a386cf0b61d76ba2be56021001be714163d8e166b236eca5a8a02
z02c40087413cbedd1e66cec2380951f74bc98041a10f87b4183102afc3b8d927d496c894b68f50
za4cc84e4a222ed7dd628c015127facb4484c5675664110f9d9a3d8b4b097cd3822196d53ff9906
zaa073c88b032b7991f131c20b9ec06ff9570ebf91f2199dc41bd2c38c53731577b7d2645cde7f9
ze1e93da7f852cb374ed3e7ee8bc271fb02b820c79b725ba8bdb5ff710dcd45021431bf88288fa5
z953c76de05e1e59996a8be664439355a2220cc9148e8f9c854225fb99442241bc7dfa4874d897a
z95f98949db8751fef9c701a780f6625e4c735e21fa27e0f2d4e75817cfa65671f73448c74a891e
z2f5037c85559bb2ff55c8b0a561b80a649554032dc5fd1d3bf41c77708fd20f231fc0dead7c725
z99df1369e98bc6e56c4f8b4499df4f8aa319143e96829fab034a98600d7d9d3ba9ba186af4b2d0
z2a4bc7f142369a94d8eb607e339b005e1e595da37fa811627b42d4dd6a30b35baf65f4f4ad9d41
z2adb2b98dce8b0b02a05906e6385b07b18422c9f749e03c6868515c57edd6983044893af1b6705
zae3fc86641576ade7329769057ee1241c0a6f155687f8188ff914c7129bb1d7d4bb9ced9915b47
z7072664cdf4c644072c628787e6adb18d10d08ba6afcdcd18314e9324bb2d129865c8bb7d1aaa5
z3527e6d2a770b01c158270bd20543c984a3e60bc32b302fe00a4ac8aa0cef50931f26493761bc8
z1ca3b9b6962e441309ca3e31a17346c273eaad9fabd48af5f624a10c3803b716a99d8dadbcd24f
z4cfa95e02be45b3d7477f611fe1bdf592f2ebee09c7d812e7fcaf596434624445cb787f4244dd7
zef456f7c848004dfc512d32d3631cab27be95ed9c9b6e5345a21d6811f959ab97d9cb9823781d4
z336a1b068af0cc1ebac2108181cfb1ca87f1409613deecd41e15eab238d7c91afe626115d9f67e
zfba6c576f81bc011dd87977a7759510b89d5ad1aa1e3d65221b3bd0522526dd00667e7dd369a95
z5612c2462d41e732da3987a84b6ec4645ac76bc23d970eba65594482a62663a0014e799e9827cd
z9150f398be598dcd628ba10ae8fe7e38196d9f90f829b1ca1f072517a8ca9384ede0f54ff51503
z66fa3cb29f1626f2efd76b145dc4465e09bc1dcb1b92b87444c02c0901d8b7da474fefc8d1d884
z2ba07c8bc7770ef001d592adf5858c54a12dd0b4731b35e70b797eb201f576da1a8e82186ef504
ze65aad89c06910ebc4cb60c336f7e3976c6443b8f5b236c4c52b749705492e3af344590b237a11
z668387aced446ba5fff8ff65ec3f4a941a286c0790452b2014a1206c1a15ab0bb689ff6d7e3eaf
z16546cd01a6b2cddb35cc4b3e21bd901e58247832d18659f6a38fa204701413d9a371d039e37b0
z17c367e1c8d59b1eadd8c17dd1a482dee667e8985c5af1ecb0a290940207fe162b4b3a44cb1bb7
zf5479ec3b40f975d182f1292136668d165e709bcbdfed6065c02ec353008170ba822da2a771870
zed0f55a7606bd63a926be4ea950704d34eedfd94ab6c9a3ec3d2ab717293ae27dd097f404ca224
z442bb1bd0a820416180185a1f0d8eeccf4ac7ad5aeeae915867025bb529605ad08aeabd4b48389
ze47b1e8ac364ac114cdf3f0f792dcfd90b25694944dc085b6308fe0c292fdaa4712d754d8c9a3f
zaa2533f403bc4c76c3ebe836efd00d7658042b9303b8ab55f7ddc4c3577f5808df8fa03dbe6d1a
z9694cd245d8cd6cf6f48c19b177063af06cc3217e7f012ec9e8f36401efe8fb7487094f44919a3
ze546d55147049d113e0ec3518ee33e411c1754c8bca0b31fa8de0b2dae67eeeaa68ca90df90ab5
zb2c23e1310e8078ccc137a9bce890b08cc235c23ca3c0ef6f30843e6cacdaae9f4e54d58558563
z65a4849ce2b27af9b9a0875a42bf325533d073991e0bb53ab83976bba0142324337bad092358e3
z0160f0968d50b15d9855b6c9adcac293d05f7d5caa8cba4340e56ddb9a9b6a845a09453db687bf
z02474d74883a2beab78a48807be1459be9ec864c4ddb6c1c1ac1aad2d479d38209f9d4adf1ad06
zf25574156339f08ae6d1710430804ce1d6d71b95ca3a76adf3fd03e62ae8d35e1907b5d9cd021e
z8ca540f1862a14e7b0ab89a494aa4bba64e007bae092030aeebb00867dab269ff2d8659d5116bc
z897ec87ade8c54bb5e40990dee5115551a4f09d656f72a36443ebe971cb30d6f08b64d1ec70d2d
z83ac1009de950ecc95e0a26dc17da9ce345703d8fe670626ea1e7c71f454a341975ffa313b3fc5
z49adcf66e01a57293c56a110d96e620c56b6422a00e4da97b03d19248476d83fa84c6f80fce68c
zda4c19bcb8839dbf7b3325cb04bf17d95dd7742957afd73d648dabb482888c0d28c4854ed180d9
zc7e2e0067fbac76b9fff1136b54c70bba421e2056f7f2ae01830d5f3e6d65e32ebcd5c93cd0891
z0dd9bec139c3de4104a0d210dc06c85b68921ab5c0602c13df8d05a9d0eb0f8a56fe5efddcb148
ze58da9715488993fb595e15f7b9f211fa52044ba9b601ecfb3ebfb67d6b04c407e3ad0e8c633f1
z2f8eec2bfd9b27310f2d258b419e8ae4d39297349bdd88b07bd36c30388034734242c6ba15bde3
z8d68bd904820dd90d9a2c29e90c5667f50abbe16447b44169cc5e26818b1d10201c3a8c8f37308
z3e9b04488af02ea0acdf82811131a55b867e0bf0e8084cdff567f1c10de3989b652a3cdff37ec2
z647f5f07b704e3689a03cb65c147e3c2120960c621c649cc1b4952feaa0e260900cb4503fe6c4d
z205dc676396024c5f693d2769c07bbc58733d0bfd577fb303b9b4ef003511dfc77c3b4db90efff
zd077cfebf1fbea0df7f7a04761a7804cc60acfc0ddff7e2430c70cb8411b9a6b30f09c3133a6ea
z28de693e196e33b4a6fcf638c3c201263753366b1af9f546e7ff33154b7677ec74b8277faaa6aa
z72b87ba016fa5e587208f4f249963c537fa97ffb75520e2b9a47f33f2f7044d7c349867900d0a2
z2e922ec9019f87f7d2112009aa98bc71dbf83df84f35f63756ff8138ecb39d9cecfdc9840258c3
z82f28b8be15a9a929f6b4eabf09c15d008f45f38c84edaca72f37a5d832c7a382d339776e29325
z85bbe5f8de2cb41f3361f7004b69737e6e931a9b28138fa578011b8c2029a6a2d751c88f07308c
z7d34a56af8b2ced4c07697d6c1d45de1c8349407bc443e7c9f9d47f897a305659166c15a9b2f7b
z099428fd14a2ebcb1427f2068134c4bccd614ca76bbf2faac378242e5148569e479debb2c6aca3
za4512a2d2d97cd8450659e6d72d986bfe4550111fd4d5c7a0c4b0448da7db3c4556e1d0e42ab64
z08be5f404d70e20e6c922eec09a19ce6d80678ba3fa6c22a40d013e92586420d340c9534d4b84b
z0e1f16f22f9cc74fff48902d488419fb9822009026d099e96230339d2465e3ca4e7f1d6d6de0d5
z5f62c92f80ae946c1c4ef8088a5c985146e661ec20cf4f1752f97214950c0f0c12dffd4bf4d3fa
z8969e051a5ee2eb4724d99da957b3495ba48f37e71bbb7b8f3698ce692f5227ad60e35d8f4fcac
z9ccfb38505611cf7a3f6beb30b89370df9e4969b64f6c32b76d7a18bb2fa557121f26ffc2f0d6d
z5be8571ad5f9c07f788b3fd384aced2f8e4dd13d6f259a0748c012065b25bba999be0b83f34276
zb043e036aa67d11b9c25777bd72bd72cc42f4fd0c3be77e1e3f72fb636a76da80fe1e98a8c7d9b
zeec0eabfc1b27cf6afd275700895cb2c116de437471bc20d364252386e9635de7235ab215d4599
z10f6709a8f335b9e08546a4ce1d9719c2adc645782507253eadc67ad2dfaeb9e2c36456c5fe9f0
z7b17fa5b1da2ad1d444440fce490359562878baef9f6c92b37d06e75303bcb1df71a814ebe819e
z66faec538a035c7ac6af48184d033ae324045008102e4152f49b0a125449fc921dce9e198305ac
z9423e07a0038accd4d5ddb4c77e6a77e3825d3a8833c829f13b3d145a67a567973c597ef276e1a
ze736e480c8558dd410a6d1e97c67d8a1f83105b5e35dc3571bb73684c231bc8be060e8479de8c3
z0d657e88a8b80bb079bb94e38d6b32c12086621e82377832d6b2cc1e0402e671d1b10b59934fc5
z245c9c20b15de1c8bc9b7ad6986cf674836a1e7162a2d6c6c74f1d0eb828220fe4465085071d23
z1f4e52c1f8c7a3146713f28c0859e9262fd3eb53dd8d1201aaedc2c020415ade5c5e73d873c4e4
zc4d635e3908189a199eeb5995c6a99c6d3ee0b32892527cafa023e6932a7d4395e3f306fa04351
z1653086f1eabd40d7055dad30b09b1fc6c12df24f8273f217b177d1e92e88263acfd32fecca167
zb0a2c56ad22dba1c3f19a2333c6b5dda086a344b1b275751bf980ce66062c32f78983fdc54e7ed
zc26021d9b2706728512776be44482906ae2e43290a747eafd7a621de5d04aba3b39c156bcdf91b
zd194c60d53ccb6f5ba2a13a94edc72a5c38056710061bdaba9c5788a9a122b48a34e62a7ac6609
z4915fa9e168c9a37469d0038ada7b972d2d413095c4fe0d37b8d596189b97b3be0493674ca9e05
z7644dbc52822561c03e9fb7632388fdc8522ab6c4a549cf57356bece2d4349c3aa7f6dbd9308e5
z25b1ab8aa743b1ea9a4a7448c2d91be315f54c169f0205e7ff287cc474c258b9bcaedb0a4b7b14
z1e5aae4de508affb97d529fddb17f0b637f0fc30a0845c0b1c63df459fdea803d04e3e59e2d363
z4bf6bab556d48b8af6b96469a3fe0e53db17d12cb7d63e32406a158e981831203c3d65f45e9aed
z09a6fc8fadf763a53e4a35b418ce726c8d1bf20a24b99ae0fab691671a5a41285ceaa48368a6a6
z6cd3e96a201229f058188639bfb449260814559589bae6c66123c43335d1d3300d33dc1388c4e7
z13a51d44ffdf8d44a52a646227d6cae98fe1e85e52c4bbe81f59fcd50681dbb8b8ff476ba76370
z4b7583e4434a41f59f4a3d6864e8623fd7a9c2b605b4214de4f9e51563feb8e3569180077d6230
z9511d4e4630f0d9f63c0ba28d663f5a2b90750332d7d3639fa769ebcb6e2e8a89bb4dcaaee19f0
za0a1c5146ee2539c6ca1c0c927ab78396a1df979816b71bfd1171d9ea539a6a7a4fd7c2896a86c
z936d237798558ecf99cfcb04a3fc233b8422b5fe3f7d1879c56af057242fffeb8f657fcdbd3ca0
z295af1bdefde7afc8220793552f4ffd612571ea27db9cc3fa66db4e66bf2adffa980403a08ee4f
z7f4a1d1ac22779aa03571689d4f27773f341f9de7c24f710eda0f83b792c759fb20b1da55fd1c2
z52398e4c669ae26248a923f5f0405ea257f32442edb8d473282c8911c86771be0af61e6fe9250b
zba0613ef18fbe18ea7f0de5de867474e35780d44d2630a09f466ce64a2c6477a75f0dc03acdee2
z0e04293d4049f9978e19ee2e0986646f2f696ba81f1eda004335484d6879fbb9a51df59b39d080
z6150c32e1c8532550ead743079b46de9ed01968eaa92f08a2d45d09f4da191b1bb10e8f6c7b4ad
zea3176619640be976386f692c25b1cabdb629c0f6057ead99cae8da6e5a5e4bf01c215f4f8b3e2
z738d25ca47bbdfe1ced5a1cf4f5f74ca22d179b72c2539cc014fba76c3d9ff0cfa926f7fb38fa3
z434421273483c68d1c17bbc00d5a91dfafad3cd24aa37ba86064cf6e44c26490dcf931d3f9d73e
z3e38014afdde07dccc9e62b5c01de16bfe7745708eb10808a96246e58d9f0dba8cfe3b07f2cbf8
z8362e873e60e01f1da1d9cd96a17a6370d0e312b7f5af917de09bc8b5844b2bb450de0e96c8ce1
zaf2aafd28790312261249829f386a05cf970c3dd0cda2f48d24ab9dfdfe1f10b0adfd491fb55d0
zadba72bfbe8df714a7108c9e8c1473cf090c3433010511de9ef33928b0eb206b04f8d13bfe0ea9
z7d2149de1020f28f575d764f18e970160e273760f4baa0e77463321fae4c617a7ce54ca7b9dd4a
z0016f024c6f7b8bb0a3bfc227d3662489b23ae2f0ea57e14d15954ae304108c8b74b8e9172af6a
z3eacee663d91b752e2d3b55d73b4af97026e468344f0e281c3c983145bbae6546061c038b25340
z995d965459dd82ccb95d10d623e90e9aae992607f5c0e5a54f5005041ab8551eb69b02b0ad9cde
z423082dd757e53316f49365ce28766406c2cef886a3a2d8fe4bc01c4affc543304f27ded3cb18f
z7071286d1295f27d5adb7f2e6b840f62a706ac50b963b973247cfa4e290a130f15c28c637957a8
zea2a3762aee4c695f1ca3639e4d86db1ec1b2bf983f841640e6314fa6b4abaa00489aa58b85a93
z441a0a53c8c123b6d735d8b164e79a636e471c7dc84b4223296c8da2757c0680eb9651a949570b
z1b69f5599533f6226723b36b6f975f44bfd124bee26eb479ba15f8b9e9e95795c6f4f5f5f19e7e
zd1913962fd9da13fc085ca8f624d341f35615686fa70d0989b7bf244a9c9870837f7bc0331717e
zca51788881e8c445dbe68661a179041109e6f036cfe8deab6606452e2ce5b8155c71c75b8eaa48
z4105017f30f3c004b8a39a41eb4770e198b3dc8b7553ceb91f4f122685e8ae45ace2d26563ad88
z7eda93227ed579f6ec5d29e56a33cf0119c2516051148459e9550ec7e04c724174bba3c7853786
z4a4bacf6d1e1abe77b5cc204e07d619887f9c68294ffd98ec0bd84460d4915591407fd2e3fc05b
z4f7ac60cc7a0771d77bbd2157de05de8f0f7af744cf35aa2c88501294fa26b4869ddc5041edbff
z89603a14eb69ab89909b8ad85163f2b2b2bc3c2ca8055996cec71575e9e96c99b19b2e9b84e977
z7de8b65abfbd4c0ac4dbe32741e33d565208fe52eada5e6a89aeb6a6568a780c76530081192ce3
z95d3fd558edb8166944f1076651f0e10bef4b10ad91b2d1ed90d633e19bbff15e79b6d3393dd82
zdda0b20e32dac84376c387b81a61888782f90e998bfb178a3433f872fe872cdc50e6d49e6ea8a7
zf624ab26c841df6871d76aad502e30cbb0aec79f5571476ee9589a988566c5ede37de338eb5b2c
zc9b13d05ab566c2681af42b29f0a54cb8d5ddcabd483f687bee4d99977fcfc38ba8c525c607362
zf3f68a0c3878ae86034930feec91cd67bf99af462d02d3aecee6aabdda6344d70e2da72c9a7b36
z37a27f9935886b39a80826796c980e575c0b8863f69dd3d3d51ac85eecb006494b80df69effdf7
za49e0ace7eac5e031d16a7f176bef302c7c0909e5c607993c325b71da398bcfbed28cea69c373d
zec1ba8de049309dbd007557ad96f499ccb4806809c91b033fa65e0131e44007e8454296cfa90f9
z6e5c6fe66713de44057f7728b02f4316c03586d05bf88fe6be46be1cf644d88eddb5fcf63e96d0
zaa0d78de12ff81aaea3f440fe319333d57d1e8181217d6e100004b45e74dc94a5e0edd28304d47
z252487514032bac7f5d6cae005d72f94be377c5908f7c285081a829eec32c406666743690ae52a
z5825ecd26147d0c03f4bc545a50da7827e7678301c3d93dc870c01c34fa248cd3594aa5a2434d1
z8a4e5173865d26b8dccf58b0364d037e6c09758cbf1bbd411cd24b3b59fa00ee97ed5373e998da
z07859b7ac81b0821a949c5d54b184abc6ae6e633f27a0ecb44d87d782c15f82faa0249ffb94185
za3a83e1b28b3b5bee44c532b9809c106a2f6eb6badce57117b701aa9d680ebd443fdd3050939a5
z257418fe7128f869d50a9c059c5f387293d5b21a1362b407958144c47c4f4ff541418ef719f603
z4f809f18f6dd5e94cab04221a50877412bb084c419cd094d337c2b974d47edcf89af0d04479942
z2a028d6e117688215e37a85b2dba560813a111c0a484a841f7d1b47f22d2b7e9ad184a409dc1a2
zfcf295342be02537b1865c99b6c3979b69a1f2a22e5addfc3d8e6e69ef7a6aac1134a9de845755
zce56babf71b333bec26b7ac6d97dc5de8ea528fbb792842c5b0a3335b4c95ab2871827a9e008a2
zcdffacc37654dfb1d20b0cdbf86e755efe948303b12a5903e3103c571588bb4987ba5d59a2161c
z24976739ee405406eb9c7e27b82da8123d17cf62566b531aee36c151b1c908d339f5df0b9194ea
za8915f38719228a39cfdd4bc8b6ac5e01dd464d94049b894ec3459d86f3d05cfba016856b4da8d
z71950ae61823a7de12ec88e6c43dc698fc9a0e5ff9bf37c33afa2077a435f11d1b46416cd4dc34
z2547e756b509272dc4c7937ab6da0f234b84332967709733d2d330017ad5bccb6f402fcf634ed4
z34792f66bd455a05aaf8a64661a61a69045d0c43432f3098db8486f228291910ca721ddc1268e4
z9c9a7a934e93f89993b548c5a7868092e2124cfe35e1c7be6661d9c8b88fe0606d5a0e70610071
zb36e9e51a0405650bd444f2d7a1d0a24253ed24fb368318bbe791db2271c0c1a06fdd369369685
z111cbbd133c1e269e724ad8acb71e2340837213720515087a47a02cdca1e1864778b57df865b43
zc168669cf792609034d2840693647c8f412cf08a19000141abfa0e49f0a1e8fe69d6a3046acae1
zc281048a4d736895d4883033ce4e43877235215af4728139098fd008482335f4fa9122586cc0f7
za6832b4427fd334d4b7fc52d27a975943bad735af514bc022e9d2150459f52639bbedc7fb9c257
z022e01ec8b5d210ee7e66f7c73f6dc744c288b80e9b251795ed82cf0ce9bcb78fad133b8169e6c
z08c4c40b5499f90e6ea3e63e7a7b4a3e77765ff0d06c2cbe352f23a63e4ef53eaf7902a246caff
z2dae1c1b97637c4baa3ab51f204ba9474ed75feb05c0c9b5dab67ac94d2eec4229f7d0ab46751e
z855f81e092afcbd1dad29fb47f082867ad0e129620222cacdfed4581f56dc73fb68546703b4686
zfc3236b955501862b0ea246a47a2f6f90eae5a3f563d79531acc34b3d874c06823239ea7507011
zcc3b23516c2434bc4aa8b265dccb0af10bb7c77185b5c4bb1f49aeab2b6acb36fae97a82f39a68
z716ec274a988cd03fcee130f9a31c9dc7cff0b96898f25d1eedb5a6b6e88ab0521f6940050db86
z334cd2e9d3188e69a4a78468e0033dbc9000d2b448a1a56e189842f15684078207dee5e345ea01
z4ce09a06e107119b132d76ffedda89bdcb1693dee619b95219d338a7c633bc13afe2f1bf35b5a4
ze4dd7fb290fab31c30422d7622c044ca53774d94118763e95fe3f14c6884a64d7287cde9b9f470
ze47745565c674b85a60ea6d6d63c60156c8d6657f7e4bfc4a494e4df7ef476f88e097a18a05ef3
z7ebe1cf37db8677d14495bc497014225bed49932739f7105f2d7afa9c9cb835b6177742384a746
z3e7ddfa309ae885046f7b7c8882db88a074717cc1b803bba3df127bbb20309fcd70e96b557cca7
zf94da3a8310d32fe76a470e745882b2c893c90bb5177bd6040b0c34772654d87d9688b2da600ae
zba24892817485918a32803f509e7fa5140ed85114154f07a3ec225774b0f0f8088ba31f1a7a188
zc996995a31762ba97eafa26d32b5ff90474f652c264e77d5a3d8d1ed96755afe02ce744944098c
z169871895700dc39905a7f393920421f71fd8ccf0d0a8ca42fc2e070d9e15d4eba84acbf8220c6
z516069bb033d7d3f479545a12ba84f56740d7f5d3729e1905c696aa8e4bdfecd5586279aa44e62
za3321590ff2e1da61089126ca6ae50b850ce502889aaa146955ba4cb73712bb05351c9163246ba
z556df0742b95a7958a28835a98d962932e758a289fa7c51d3f3e587a9796c7faf3f53b745bf4f4
z21efd2013aec9211b616ad99cf28e9010eb3ee40b69299751e1ec87bd543e5d75d4e434abed92f
z51bb3425a3b6771abca55b9c7b14074cd47d12a0fd6f8bbafa6d24ecff08bbd476e17bd831fc7c
z3a14c5823ef20523d3ab283663ab5fa41985efa048dca5d993a48bafb12090338734b4e110184c
zf08c05e507d0c0e9cc16ed44325863506b39b710b3d409605813d7018aa7e1c07e637996242796
za8a18232203e77cc0739d98e7ea5777d58d52f49e1e4dd91c4ab927238f7b4c07631aa7e6bfea0
z4c073ee1f95351d19a8324cdb30c4454c7dce2b1ed3a2f066c1668788d1430d940ddbfab5b8944
z45e5c5f06e778efd8b23d92837910b285fbfc2c5ca2d1fe3d1e313aab170a7d8111cf115d0308b
z546eb70320cd4f17868d9c9e395406ef11659868169d616188734b33c2e3118b847e38b8238856
z3b4518321703656cac6859d1c1c9d4c884b4e6638b1e32d7a2fb02a6325448f9e3e4596fdc13c0
z6354e3fadafb60abbd7a8fa575367cef617a195952b0c7841af727a4c8641c1e2663b880d60f10
z70991ddae8a7ca40a44170d3fe360260e50fefd9d86ee2b48368c320dd681c555925bb8ac6e335
z16afde3cc7eddcfbc68b3ec07c27de94dd0298045c3241fce17f5b0dcec52a2188447b314073ad
z7d0a67934161e0845acf401543e737e51125200838ab8bd8637d212d351c94f100802f632b1e5b
z5d48dd6bc6fb9515b2bf3802125287d11aa668c7556e4ef4e3067f31d8f0f7ab8bb064d060b3a8
z275e375c650f85582255f5c644158422fa7a0b695f4d04d1ecad0453da73ffb221442ed81fa8b1
z169a845a6a26ccb10f4c78ee84668fac56ac154217128beb989da3c9f368bc7f397a1798ff9b11
z7234ecd9e936b3ac8023dc22eb96829fdca7e59a52ac1d0d3b9979793b3b45cb9e8f30c7108248
z4874c2135dc9f2f61ff8bb91cb4a522c3f44ac2110ce2d91c823751bb1561f5493d59acae0c9cd
ze86bd8d0643a651b16e89846f84df8566d9d362432c11c3ec1b8c03ab5e70b84b826fe837ec03b
zc50b063340659a2ef77889b0794a49c817d3f26ac054e69da72c4baaa577185662ac455cbf980e
zf2e7be9a1798282709127693e75f4ad350b375d57c67809de9b8b175956e7078afd0e2c9a368a0
z9477eaeea4dd94c6024e56f6b752df21bfb10b389185cf63841c7020a9ea8aff52dee15aaea67b
zf4d4c25522fee39350a6f3bb9af052b06b4418a06ab719187c74be9cff53adc23cb55ca876a773
z5ed9a5616695c8ce77de2cc7e373f17038a776908993689d2bbe8cc196087609928fb677101a85
z15e549027a85cfccfc6887519ce76f603b144d1744540e9707ef03c0c20ebd6d1d7ab4c907f1a7
z200af3cbdb80139a79b391266c3d6d2962b3a35f70c1bb084bd83715ad969ab5663b9af48b863a
z5d370cadb7d959046cbc6256fc833634a5c0717042c297a9ce0cf1b69af11e1d8610b40f77d155
z9de7047d09952fe459c61c9da4c70eb126d8330876c890285739fa67812f716caae4bee4703fea
z1a9cb6b63869c93ffa2b6832d50856bf9956b387d92828d0dd7891ca503fc6b377c1e986c1e2f0
zb3c7e3ec3992bf0bef1ec280d3dbb30d90657edd1033933d5d0e891495e230e8f21dfff1f1796c
z878bfc56b0b9d9171798f3e12ac7a9267311ff01bbb222d972b4f326a7b439f1a15ca62dea0314
zd8cd9801e69111064bc985bedb137f4887e6ccd1cd7dee2ec073e9990e967d22da120a196e753a
z9cb92fa164a5fb5c42627e4ba4696cc4a0e28ee947be0404277861cdede285615bc025d87df7a9
z00785444a71293c36a4a8079c26d78a84cf5bf4b187486baaa6d925bffd2ccb06f53843d569a3b
z0e0c783e872ed72005a972a2295be5b57a10600eda539b3e200d3b37b847f8a70b12847109d63f
zcfdf368f727142d5d6f419169a2c5c74762888395c9eb45ec9203239117cc4038fdff066ea70d7
z6c74caa933c35786c7086cd7f87588b85f397a27d4ea8015d6ae4a45532f02e585c2a843a06c0f
z0f24a9e845568f816308f89a63aeb8d663b1ed3b250784af3cefb891df7fbcb80ee3a48f29a53b
ze346e42f449ddf8a6267164f7c3fc68e2bf811f2ed13156643f534a87fb622fa3fc558d55a07d0
zbaa9204eb0054b7300c489dec32326dad7c654fbc08d50dfc54cfad2e10ad0a3fa7c385797d4cf
z33cf88038aed7b8c573336b2eaec4859f754f346673804b147630483893c5e93152f7d3cf1480d
zc2fae5cb87cc0438abf38472dc0752f671294caf7d919caf0d3eca358b75bf7e646de2c6d5d182
zec7e276aa8e6013d8c35890028647d77272f30b15f27cda85f4b746d890fc8f8cc9421c6e5f690
zc0859ab38f720edd6ac0bd8cb8f26a4dee0e1779113cc7ab4f725b86dd545ba0afeceffa4a762a
z46ea1db97657a759f07a6b60eee2c223aeede12a31745ac1c1700225b27803e4d5bea098a7cfc3
zcf6d65527915de1575518f16514ade27146b1f7cd22ec5ba7abeb8908701c06e10be114a3d5db2
z5ce208e0950f8886b6b6e8eb595ad63fa4cb5a054c2acafa69ba1d9f49b8047ed3215fe4c0282a
z3143ee01f4e62c99c3dd3d774f756de3da82840dbe7157e44871b6bd5464424ab8e41ea06cd453
z9977161c672f1e80756ab8e7586cd0dbf2cf66df6366927cae8b999948559fddf30861e64643f9
z7f67b2b6af414c9bfd06171117176d8e3b77d86116fe4be341020b500e90c196f1ea7f198a3a83
zbaecb1a61d98ca02ed50a33a8ebd15c669f68c59ddfc0ca9a704d163226db41f0aa7eda2c2f342
z4bdbe0376ae559dbf55ddf6fea761ad30f2c752d9f2ad1bc23cba027e5160e13a15b9fae8c93ed
zaaed471d088a3758e77b3332b5b64bbbf290040322281e3ffd2ae2f6c5ced57682e22ca0102f07
z29d8e1ebaef66cbe24f41229983af8c649eab2ed00ab18e3fecc53a0ab34b5c4af134d32aabbb5
z0620ba69f446d7e6c21b03ba79cf6368c306572aab7de58daed6851a5b3c71f7269f5cabef870e
z8009e6e1b303cd996b760f2573e3d59138e619e568dca81c6d7c0278a238447e63f5bf455377aa
zeac681ede4a4c6bf891bca924d9ada15184ee012289859c189ebde9b0e1cc7107513b75c548134
z8a4588d6374fa87e7219fe8abc59a1eda2dfd54a389c966a3d7acb4b3680d89b9fecadb69c3634
z4d8e7f33f312be6eeb11c91bddda9a79847e0c9a6fa737163fb6588aeb8837e759492c8d486c9a
z547cbb9075345683db537824cf5a3839bfd5f18484ed136806078437dade9969d04c5fb47d53de
z3535318951f68f1cee0bd09826016add86361e0d7aeee2732714f4f31f03fadfb96fb27722c036
za8afa35b46b4178af9d14371b94844ad4a30e46b8ad7e69baa744f86104bfcb474cb633a2cfce7
z98d9ff41ba80c7601a9c35f7611ce97d2b97cfe6384afe181227796da36de0f147191642dcedd5
z951b9210d4af66e7c7706ed149f88802d6e769b283a017154001b1d4f7d37b77675d4c9134793c
z3f3c739757a8e18c167fec0c620ceeb143539c5a044f9ccc0a6cd8d1201aec6daf79326e8b4fe7
zd11c9b6b1ecba190bc4e1140966c3a147b52f32740dc2dab3d0e87d7b389ffe3f607a31be49374
zed16bd406d2bbb9ba336f2502b06a9dea50339ccdd934a3de5d0551a9a05ea54689239b5a3c730
zc6482fa2635632485bfa24b9e7cca21d2c1426172561156fb467d9f8743c6dcad2041667cc324d
z4e52b9b458a07ab8a2b83704d2bde3f166b448a859342d8f4bab8f316213e44b8bed1ada74b6a4
z2fd51c3d988e577d5eb01fe229390a358a8bd3f9dc7384e0e795fc0dd63af31620857f8ad44f95
z084970ee53336a882e7c47fa1394931545623a560dd6ec83004a7033e4a0d347e3c37412736bb8
zf5a763bbae93e8a791bfbf9b9a0aee1258f7f540f701c868e24516b336f14f939f170f940c0888
z1fa34473f0992cb71e660ed2a4537a4826e8ef61917977bd3ffbae1f05ae49b9a29a778bbd1ce6
z48036beb680b805de91ce79eb57e4cb0cbf0590d4110776c259c47472a574979679abc3475688f
z002053661a46b8a46e10f1acc9ad5dddd2542bfc7007626a796fb252ec5ea4663bef6663119825
z4c7b207aeaecd03c418b0b848937d5267304a49672f0ed7e3513d9a08d9f10a1a6d0db0a0fe057
zb32a48cbf2ff984f17d0a1686f989fc312d72bb60ca98e90f9341b7ea04f8379edf69f095fd2cd
za5ee76c885c59c3e1d1525fa3ca28cacc89753a4955c0b09c522a8d7b96b6b27ba313bc3b1eb94
z427d37d4c2a276e5edf71caf0e7e2bcd9f3e4b4d6e77864157ab1eba96efa488f618f453030fe1
zda37b3d562087690331ad6dcfc80349f810e602ed9dbd2ffbf82377f1dabcaa67ed5b62d1f90da
z6fdf2dfd371549aa2c6c6e05ad93fa89b0ab1ef73b153972b6b11d9512c5324a84d46e1049d387
zf283de5eb1c8d10e3920b2c0385b76dfe409e44ecf22b7a4d7ad66c7a39e458bc7a3c873c85527
zdfccf1cb72cc5c5cc2d5cada350001627f7e86ed42bc8e508a9b2e26a4a326587680d49020cae8
zc33d173bce02801e43d2a6fb60802d7dc7b37873919471030735178904b08fe5e251530339d768
zeb97bd5230c9460e06aae3c874b0816c9f0da409b5d2f552666d8a32c65b22726d62ced4f40a1a
z2298f91209bb65240a287040b566bd0df35b3282191b0b790efcfd11051445466d0ff5e063c4eb
zb660e1663eb57859d7edd2b855dd06ad02e69971f6d271252142843096a7d816d00e1d8f724978
z3676b435621e9858d492b73156a638e15194d0adc0f0a0ef6cadefe4f6d2c1a573bcde524aa28c
zc59895660b03af245091d32f159eb0ce8e2750c351b84f284ec8ab1abb473346b75fb076b3af9b
zc20af8dc3560ee603fe2f0199fb42c9d433ee91e40fbf660e62bf6c10c3bd1126baa9df5e76882
z59e338c4408b4427a2a508b7a3c2f9731c61ab14f5e225a52ba87976a88a62acc871773d9c36b4
z050d11e788bd408b13c7edbc7100866787e96c7c56f680c68ddafc2976bbf7308246f6352ec768
zf50551c62ada345e92a5e2dd7fcbdfd5fabf6377ca907e705b6b4a706e0162b475dbb2d0a4eba2
za97b2e9352eff2908e8c06193b13c2efb8f0f8730b7e3b2a43361f4aa0eb51cd03c110fffb71ac
z4e49a465da5c71709d850882fa992081e1c7698ea29d72acf97a39e1d715709eba7a8566af025e
z7725a9d5214e6d55268323fc8f2c453d4a254c88c4d6eab927d5f71ffed359f6310b982a019bd6
z17f6037ad66fade513574c4dc1c1796c61db01671bb77f2a731c9efb74133c5d266f5a5fc36e97
zc9c556e96768f1e9c5d66e3abbf98a6a8f8a2b13d192d629ea86cbc0e08b4fa4bcb8142060bf32
za46e77adac863fef923a4a18dad800ad881672aa99b23781ad3f0f38227b4d30a042814c32dcdd
zb295d90a1c7094d3db8c993f973f4ba2cec18a989d3af349e711dba57f7d1b98c50da7f08bc87e
zda1faf7edf446bfa84a0080bc6c507e1f86b32ec54b0b911b98f2535e72897937cca0c79051b2f
za474c8b185535d0a2786f253107c257a84395cbfd85f5582097c05094f4da6ab877d4e62d03935
ze71fca0ccd50f02f0f7916bf49c03940b3bb0558d66d3a61878927d1165c6a275f9d1e35186493
z8cc280251f40c2490269a9af68798ffefc3e55c1babf5f1351be062346640945ad8a05346007fa
z2a4842859e1f2150f980ab777a36f2b2b37f5ef06c26d7f7ccfd58d3f6f055d7ca7ba62d100a5a
z28ef50f331d5984dee2140f3980c2d0cb217c70a9c7a32dcf9d025e776d8e648d8b8f2534f005e
z9fdfba777c66e499dba0c22f44f5fe916d9de9e8409afb37a327ed95bfa51218c4317426cf30fd
zc7fccdf7e90a5c7281d58e97b1f541bf61edf30020fc8772f3c875af4fc40ef1703f241de61aea
zde6418f8780e1657b5a61d39d9d085bf0f2fd255329b16e3d85a4483d5984a772fd41e8c20c130
zacd51c8b6365e3d115657dbd87d388a521f666a6638f4eb5b73262e5e8152cc52c59a05ac72186
z3ac75692a69ba3b91f3528e653e019b28960f72c4527d1eea8b51a252f9edd6bfd6fad07c521ad
z758860ed2f8c70ae7b446cf0379bc8cd6e5dae70268dd45584d022a58105a1b707593bc7b788b1
z8de4fd978a6302fc0032ef64e0539f4da497b8f7b59f64e09902de8263a21fd9c255b3089626af
z4b15cf189c48d96ebf1f36bd7f5cf915cf8aa64b77a4b0dd9777904692e83c95d85458811242c6
z126baf1cd4956c430f4dfd169211e773a7b66ab662773852ca2ba32554356d329b745841f88387
z160436e8742c4be345d1c8267dad9ac80e9cd35df603f07598edcc39e8e3a9ee7413ead4977c2e
zb671862e4e28de3cd3cdd53e6ff79117f6f157dbd39931e164dcff5178b20f7a6a9097d5a2a513
z31463e6880eede9dce2900c14dd56ae46a7902d3d2135334e700bfbfa8ad84cc0484d589a2be05
z97f5ac6e6ad3b7fc3dc718813cd9b2e66f8c1e5f14074095b07349064ce68a655a2c21229ce1b1
z051d97fc957e69ea0a53cec30e7482a1ebb1f353be20f75496b7b69d13a8624381b0ef803c05e4
zdef6c54b5ed495e1f21f13b564d741094cd459beb64385c9eed960aff5267350e7ae4d60e0cd60
ze34409393f053a53345feedee64fce1f95d218a7b4de401d941c79f9c4e903c81a899dd424eb95
z8119f1d5c564ab23af40c92307e7c4590c58250c3092643c015a8b5265d475b0c7497b22102bd5
ze8b85b24958903e6cec3c365f211c5017d96ddd32abd06d9c68196b94a9f03ceb25ddd90d586cd
z7a3c9c0b0fca01c0d447591f4bac899aa4672e3d96c62d8da36cdc6ce9a8db072ce020977dc2e5
ze288edf3cf310a0dea2ddeb2a683e591b074e2b5f25523f6ff03085d9a5c85b5fc25a90bc74db5
z21c939618f3441d69e277a8005293e038c764890b90eaf78e01f111426c0b0cb7ab83d177591be
zb8c594fa8558107d350ecf9a3a8bf2c86da891c36a6b5a5abcc1719d6e13b6393b3fa462bf7fb5
zbacdbfae63600b10b202f294593506da0e4edbcab54d6f72a4b5cabaa780e345973d73e80138ef
z53d65bfadc5a7813208c0f698238d63cd67441a48244d0371058f8e8f403ffe15fede8da432cf0
z48974ac9d64c5133121470df4efe9a1bc6f93f051f8a6994450c2541faa5c2af250485324c7b43
z99a2de38ba66bac6f5ecd326240fc6b38ca0687e5bbaadd70b546a790c9609bca6d2f9393758e7
z0b42b5d9c108a9fa0ee729f303951f7a32de072c0daaf32c8f2b68682b3a8397a8fd6f15beab7a
z39ad8ca7d8e6387cfa039cad7924f2d258db1b6e34644463d027ceed4e7b1c23c79cc77d50c16a
z6dd752578a54a3b3df6287b13d157c87ca989cc1b04851a3adc147fdf280a85dda48cf25bec652
za0ae98976f42b2e75b229d8276198f22f2791bf0a3467cc85de28fd92f0e15a409e0d064a93114
z0440c1f60d4655c590725e45173a64556c51ea8f103b7e6d4f9235c3a5b5c559da2aca02153c21
z00b89dced4f0c02da22f3039b1e9d730870c7e45469bbcc63e33271a84d6b008745ccbf5454e88
z7ae791abaa73445bc9f7ae9389a37e55d9dc1c69a415f79553793b3e43e58c29e91cff6ab2fdc1
z75ede72e26d76a1087d1a9c86f1f5a30e981b8e1d0b19f8c68d97c08f96be907ba2c39d57ef38e
zc9b8a880ca74e96d86adc2028ffaf173acd649a14c494f75bc908cf5ebd26d9ce80e59370c365a
z699e117025dd824614865caf302b59c937ce3871cf1acc3cef709188f19d90e403a0138ad815e7
z2eb3d8e5e7f6b34b6e43566294d49c50a22267ab5d1234583a3aecd6ac0601b682f655225393e1
z52209cbce2c15c1ab5860f9dae5d934c28855b8608968fc6a66d4beff49278a8ad6ab7af0c0430
ze280365c5932fe9fe847b622ec5c4eaa79098b7416c614f9c89d667f198debae88087d845726e9
za8d16b5d35d27553225248fbb2c8764b7b4b214c2a0935d346840c9768751a0bc87e571cea4a19
z6abe06006978c346222f5fc919d8fbe61b6be2e6b48451497a68d0d662638b42d0fcfc6c76aef4
zcd21db3e6ccda1f611a8760d80f738ddba8b7cee4e3d2276036b65612a20513e6fd39993d84a0f
z1de2239652c393ce47d31d9f863289c830cc13b58b5ec874f481743829ddb189be0116f3702e2d
za4aefd060a223545de341cd6411fa8385fd86d809bd46f899cd8dc5d4e7ce9e58256568654b970
z706fa81a43a32c6634dd9a507c2487576bf141498071cdf6c4511d73025c9bf4d21a65428f2ca1
z7ec4e9750e43d6a3fe57ab7d38931afa997ada3ba1e6ff5a16ec8096296b069e13faa275ecaaae
z8d9cf82c33c831cba5598baff1a6d7b6f1dda1e8e8363018005839c4ef79e43d9f6ddd4ff8f050
z6555033fd50b42384219c570f0ec20c0ce241ff3e5b38693e5810d32e6e8235d024679e8c9dc3d
zf0d17b8a7c93166d5d0a87be0e626ea840806eed3457235ab840ea5b123fed6e16f7b31c8549b1
z112640c9c4f0cc297735581050193abc92203d02696f927f61e558c1019312219274e859432d75
z1f53384dafe46c7f53151193a15b47cb9a84a5f2db6e5b180e568397ab60232523d4467e251b2f
z346dba9e52a720b415b775ed141cd7d2bfa5375248ef16112bf5df7644045a8565b18b04ba9df0
z633abef17bf25d96b78ada02cc66ca48548fe44ca328a01d78939c0a7c0ff0dd4c4054af387c60
z70c55ed4348e53863a8a02e24606f72cb9d2e5e968ee45035c49a9f662a4de596fdeef4e132978
z3cfab6294001443a1d0c1582b5796e5c2ecb1bb2dcb1b09f43b99491d779ac49d423acd523b6ea
z1d397325589ab8ae4b987b6f878bec3b1739f28b828e7eaaf976ab7678fdbf4eda74fd258de738
z0b2af8b7aeb09be39891eb415452a814cdd330b89bf8637a3ba1199b41ae0f30b7468a568d71e6
ze0d99ed00d17d3ebe5e6bf0066515b0e9b077c6a8747f0c971d810745a709c36bfae73310d872a
zd769a1b22435e16d15d6a27d89cf1578e0a97bbb6752e7de021c657ccc103a0887e951d38c882d
z3a10aa8c0158c895fb9705f272fa93abed02761dadc299a2f2ddd14c36aa27326c6d53481e56b7
z0c99fce4a19c2059ec91fbfdf3b9dab22f35b2090387d3fd7e1d48600b2195bedd61d7053912a1
z8e8bf6d53fc7c350b22a81e798f4fd446415eef059db18d672f8f460b381ca6d5a5d8e947a392d
z25507b867e465eac6f2f4ebda5b38e13d13641a1692bb1ca2b3caf7bd80b77395119867807f636
z03eb8582c7a511828fc95d3e24a48c4852805d65cd31d1befd267bc85fa20e4ee4687fea799be4
zbb07b2254f853563a6a0eb34eceb565cfb63d6f446857075610814c6056152ace7018e8ceca06d
zeb678dafbf92e69703206c214943952218c23210b3f85d2f896459c42ca58e749e7e708a81d19e
z7337ef3766821a8739ff350c59e6ac1d3d465ec7840b9026263d4cc0075c6a95951c79ece325d7
zfb1a971f2022ae708ab550135f60f716d3d52d32992efef64747bac086629c241a66e2d99d9106
z3555530719130f0e05d65bd170a74f059bacb39b20874bf3f415e98181dc22d4aedbff667a97a5
z86a87fbc6ac51955a40ef594f34b6ccbb6df45db7ef84f87503c3d85676ac25f69d633497ab228
zdacbe3d2dfdd5e05c6f0dd95be0c3a284518d2f869a111ba8481f1ccdf0157dbba72db5446161c
zee9a84850d0c0e63e18372ee79e5e1fe18b2bc26769f362d8c81ee05e2f4a34703e617fafa64ea
z185d4679e22669e2a324d5d78102ea2bbd70a50802f8060b7d598d1207fdb59ef247becc96baef
za2fc50a268de5e15d6763fc2a6500b81eb094bac74eb7f6da57881a9e7b5ca76326f481f1aaf8a
z0e80871dfda16e2bac5ac532b3a528a8d92e824334ad49b49f5d349cf77a4f607ffe9dd8ac7295
z112c304afebfd064d21f553988631612fb45519b06e1e56c1da42159d114e92880eb9bc1fc50a8
ze4709461fc4c0535360ca7bb45d24a3d41f0e7a97ce9de0c960355d4d6e5e1006937bfc1a60db8
za41bd067a811106562595d1d3dfc69baa93e3bd220c26e531f6e7f800834b66dac113078791f5b
z138834fac3336c0c3ad94581c0e6190da0e2213dcd007458ea64be75d0f7c9a3a4addd2021ae0a
z9d18acdbb93271b50a3df053447a8fe116462ecfa59cf5659f5c96c7e04c0a920b9a9578728811
z003bec5d90da11c8d11b8a57d1f1a109f536450f277f4508b0c2cbbd661b5e8faa626df87998ff
z0441f5a7e300ca8c9fd619196033738fb99518f14f749021ce1f3e736197e4ea2c041c2ade0517
z769293dcf17babc0bbc1abc03d87090c1877134fffb46e73cd8334bf3a108a0d4b0d1544a97448
z6b579ba3cd9d0c878117e195053069db4c5394a1a5cea3fd33c142158d8496922ff2ce4011e1fe
z4d81af6bc81e447bc66bf4155d79544eb6252ccc3dc97094f0c51d944e19bf70d55251dec4a10c
z16a2ef8db31a21979bf48d7356042eff3470513c3bf2d688d32a98c54535e51608b4a89c36de9f
z387e05d5362442237e35da0be5991564defe1ffe5659e7d0b8dcee06c05d5d86f7799be2c03abf
zc6095e16e12bb1dc702a3a99e64a05bb62b992d035a065f7ab8664c3bd98242a2ac4027616fb43
z8ae6e8b20d4bffda8dfc0588d5b1b0388c23f6ac1ab4d18402f4397a87e5ee17b9487e0c370ec9
z2aaac0400471184455e95b075d1cc4da82201b3dff7ad701c4c7fa4e2371ec11db763b788df978
z20fec9a6d65d66b204ae72fe766227e8224f724a044831c6d3a50685a62c94f3be3c740074b699
z5e60b1356b348bb0348779f443b722160f28db699edde38907a1e87f4042e1910448a6359b37fe
zf5dc4d64b7a85ed9d7d91f808ceb7747a414f6cbc3f3064da103311f7327e9f80ed75707566054
z84c66efc2d0a67f8cf803826a1165587867003c6c3e975afa0426f7b3c1f7fa4e1c171f7ea7ca8
zadb2119cc7afabdd13fc98be6a6bd37f4c662146efe5fbbafe394491703864eae1dbd40ac772a9
z18319b95b8c5cac1fc0de14e3d21274adc9c549e797fa35ad68a0bc2a0b56cc7b14878c8b8e825
z24f4c4cabcfcca02f6db3b93c66b3d2a6ad838010e6a377b21e6a56fe66ba7590dada3eb3ffa2a
z6f8237f91a7a7a5b561bca8a564a3e512aece7b93cd98c6e7a30bd1b18b3dd8c2f91756ad16552
z08fecfbf025d3bfd586e59cb778b602c973e19a825e7078e6af266f6af85f50bab377a8346e8f7
z3a6610b863a2a2c7ce150471cf4e3ff781a9aa3f567a62f4754287e83f97fbd8d017ec7116b5d1
z7acc08628a978843ce103b9c2778bc7cdf9714cff1c3d506070337d271141351622bb70203677d
z3b5aa3445ec28d84cf91bc6e7154d0fb8d03409b032ff4030e718b54ff784934bc66e50ea117e4
z65d5ee5a22ee01b4580c4b05b2feb37066bf5a7286fe81e300390edcb4fd171cdd9d9a5cb9337b
zae1900aaa364078be38ee3e28faa95f261945d22086ff3f570e5a0db5b319a079623e2ec59dac8
z2813213fa007cb3db5bdb164c5a2471fd9b9b64af167e14938231f495b043d46af540031d5c96b
za26ea933d2da951e5a8f6a3d670e85aaad77d1b0b71e3e289caf391323abf94d5ec6627add9d54
zaf73b04f0a4dbd769c8befa3c3d5c9d6710836e187673293167aaa5143623798a6e2e4f372126c
z2aaf479509a7d8ae66a3ad8f3155e4958d221e2cf60c4adbd5e6e64947d57ed27df84600adfa82
zf3a6618b09ae5c0b81f96c9c3fced6da85ca82e0a986cf680d75a45909682c8ac1344c17b54033
ze151b89aeb088005b16cb4afa69d4ccfd915119fa58322621288828b111e9426326f1ed1d098e2
z77c8ffef0f6f8f7aca77eab4635fbcacb0b1f06f12597ea891ae26503c6ae0dde5a57621ef6f6a
zff09895bc82391612d4473734b3aa7f41796c39d608916ab50e3ee6766c2ebeacfc1d06204f9d0
z94a3efeaeb1b1565c719e965f9329c7cfa973dc1c7e7049c6ea94f8b7b0d0b145e8b2437ed003e
z6f2b1e102c6ed7fa6e358d624b87bdf9ecdf12b35a06c6b76a462a09c84602202b0239f8c4c8e9
z6767982a32f74e7559d0d37401e2fd0e7f8ffb084cfc661bbac4844cb02c52bcaecbd0a297d893
z9b7e06f328cf8c2e3aeb4eede9f64da1a6679c9b0a34fec6b1eb706679ad43277d0630c35ca241
zed8d3d875e3c95632f868473de3caec4187890d2a56524fd57302c7f08ad31af06ab00cad8f3a2
z7a947efe584ec69b8e0ae58e940407b8aafc3394ede1a4b3a31f91dd028a6b6075508024493de2
zc483d81552bb613848fe430c69bd136eff33690e459f00c2efafbf50dbb948ee105da5a64fba70
z73bfdcaacdc09203d176f0e8f364ab83e183fcb563d1b1484575680360f54df8d268bbc97703d8
z23ede07ee967ad1b706943fb3db40404c9b1f0b5fe632ae4da82cc61f1c077e1e736ccf4f62187
zb01c4e7f53ff24e517cb2b75cbc1e3e4f5be8fc9bcff7394991c06a2b61d733216931b80a4e5e8
ze46acd5e8b3588b4e85f04646feabaf15230fcbab3b25a1d1dcef2965c230ea13113d3fbe771a8
z5b7a35f2b03a496ada6562539152cd13957a2e256e48bedad343cbb2c630b4fae9147bf6a11607
z76df15feb73a06ae5c8f27608f813db44e6595fda4c67188d36c98a6b47bdaa2b42bfbb26b9471
ze933faf3938cf35ad1d472d4284f5969e59123dbaff3e10d48f41ca958eea584076e9e68b41f60
z6dd2f4f53196cc16acd511c6039e2cf2d948af64a1854eb1cf78a282f7ab48a948dd10ac130049
z0de78902c0a31780ff37799d3c267a321040a3cfa37c6fd2df252d26cc5cd58b5421fd70398f4e
z25cdb37b0625df750f8d8f417078ac05ac6356bfcc5ee933d693698d805f611c3088484845efe6
z6057d4506876241109af91bf35c311e9625043b3cd33f7cc0f8a2ce5270741ecc0fdd0f27eb246
z0cff4c9986e13421ff7c6af59ca20a48ab5cd2b9813bd2870354b6a89d0ae5c718209ae1117f98
ze974fd87dfac6387246e6eae6edb56b103e5b52b405a685c08834e1f4b036a9e77c7b6deb0d964
ze00623e85ad71b19c9ad2cde56613bdc303b45cd6f38e0c58b4e77095fd9426597134f1d06a344
z761e0b2bc390621d0ad0c4a8ad39aa2d2efa46dcb6c52bc3f83bb68246734aafd2bc6fa89a6ea9
z3dd2999b221010252a2ef5aa418ceaa2c007fa8e700c5dd741f56dfa374e6a07bc6b64eebaa991
zc5e2c3d9151443e775da8d9f85d2f6517f865bdc0617f930b42df08b3221eb1715dbc96be65d40
z73827bbb4622bdf9c758049c4a82fe83bd8f29db0ab09a06d3c765271f4da2d648500482552f2f
z438ea64d4477cc3add9e8f4d4c2ba1fe25a92a5d70c2c2e0eacce7e47009c60bff24bf999d2b96
z78e94894f0e56b968d64ddb89218c2fe7faf19e6c6df65311fb1f8bd367fa348b3e5037ef408d1
zd47e03c8bc9cfe2b4d3d7251470d4c67c9064727abafe3fb7de529960ba862fb705535890bc38d
z493b7ef2c0618468f8d93a205b5d482369839ce0d8dbf1340c77ebe926e5de87bb62dc369d642e
z8ae264db91eab3ba7dacf754d64ec24fdb8a4aa6d753cb9e62c84d89f05df0047290fbe8350ebd
z7c31aa4167c9eed4e28d66dd48230e67161d3c328d2c4ff8fe9fadc86f2d6089a0f17549cdcf19
zea83c2aa411224e2e96be99b03a505b362fb4fd565185d63e997925fc5e49aaba1b3244352c5a5
z6fdd3deb26688ae878fdcf69da730ac02ae25485b739bd86428c124caa833f08e6d83cafceb658
zc2d6ce29e50dc5a3b80152b8f9df8f9693d1d4200210e52c1bc0425b54b415f9f768f8fd778a4b
zaa677b8329e8540ae0d558fa16cb7a863de28dead41b884d55cb508a9fb2001b243631630deac2
zf91f40e9c3782b8a8faf15c2ec0a4d74f693b9b0a326c1fbee4ca9c68e15315cb96228b9cd7be8
z0c43f01897730e48aa61095e6731aeb86250c25b354ebbd5e04c3ade79fe07a684852e599b1c71
z8d037fab14e17fa5eceb18c6621653c47df5589a4f0fe621d6af873b56758e12324668c912e1b8
zf42e1e7fdb88682cfb0095e29803166cb6deefb512934137e37f9d6deb0a4d416f6526fd2a295a
z65f66d775d7f899460e1d7b96cc3555bc868ef71a837f8e4364fbc56c55b38d0fc863aabbcbc6c
z81f94d1db9764665b042bab66f0f3e78eb8ff4c8bf805a58e9d48e68e14788ef4b3a898dca54a7
z1b5829674ea8da61040b49499f1b6f73e726e704cc9621fa2ac8d2a5bb466224807f5415787bf8
z59e90e72efb399ad90e647f58c5eabf503a0f46a9bbb8018f6c6a7f15b71d2e006652c3d270fbe
zdf9cebe8c444e1e620ef427651543656d5f0d928aabc541175bca936614510305ad7efc205fe64
z66c7a7db7707e6e8f13ec628e986d16f3c567c12b1ac3de3b16d7f04908c10bc9307c126fff858
z32943aa6ff9899fee984df74f6864a47642d9142298a96d6854e769b2d3dba9f980bc29028101f
zd1253128355c3a9ca9517e3ba88b9aa03baf51f0e0312ee4d53f5c4ae3a949decea7f32c8e91ac
z364cf0658b6850ee2a930ccc23ffd75366f89dc0c285cf205d823c33f7ca9f1a519c550e7771d8
z09d58f49683b30fface9b93c92b041f00c28e8fa522f4deadc60cfc37eef409cf72f12735295d3
zbfb2b6364c31f2d3399c1ddb50499d03c205063668d4b58d9beae37d2ac1d667e12eddce61ed05
zfeb8153285bf8c67e97d81563c9faa7a11af7fb73d26459978aacbcafd0636031de61e0c7c6242
z98e366e0ef31cf01973ba7c04cc4f4294fc2fe26341e3af7eee024d206f4bf80561a7f3f1e7a57
z1195424fecc55429227df9824777622f810aee64e553dd7e6b248363d9379e1ec853ab13ee6730
zd21df762fa410f2b4a5b93bdd590279f0bb866ffef0a694ad31ebc8a475f84d0efac7fa4523855
z4d0ea5dda2e4fd657e1244353fcf173db4e7d988d9cad6193787deca0e036ed7a047e93734ea94
za3fa37a2beccbb4a053675b37478b8ee58ab25ef2721d532b78ef1f4da205d990e72c57fe14105
zbc6d5f00a4d45a4936fffe0b9dc89c59fb6a881dc1cde95cc8643b675f0959492f1e0c5d22ead2
za32a3bd832e972c7cd846cca4c202d0fcbe429dcbbd7f5714277df2de620f5366e39e89daaaf10
z3ae77e8b7edd96b977a3964dc68b2e90d1b05a7319b19c98bf5154d4fce6c3d0d703013e793c2a
z2543b27a46da70b9e72832be1eabebf3f32fa71622b9c3935b5ec52f64197883ba707385e58fca
z67c7acbec5e8d40eb17dd5c10f0d200e01543ec24fdde24e697897fc8fc2e3c0b8966f2e240226
z53bf11d8cb61b8c0017c597f4655b7b84439bea4d87d555595276e5e8056e0bd71fbb9658d0a77
z57d94288ad22ea29817e350dc9f4c8b8697f00fa529524deff153f954829f7112e62c82f17e9ca
z2b9030ab821cb13b71b67902bb48abfa424862250b53429bf191ca28d989044b8a82c90d543c86
z142ab8623e9751cf3efd1411141a5cb755603515248484513e6454ed126ede8c15f39b83e121c4
z976e7cdd649e6d92a30b7626c5db38b6b6e1b3e2293058ef2f6883b55cc070c5cbe5fcb61681a3
z72e58cfc5935973b03cdcf1229d9a91d32d1e4f3299666868792acd54e2ac8901cd4411f5376ee
z6a860c594a0e868de397893c8ddc34f8438bc1b1781aa9c8f20d669c301e558153213240765081
z0f053290643ffbeefb80ff47793b8b74effbe8f0170cf870ef93ab9d0c7e22782904f936ddd466
ze5191bb8a2fac0bf88a20c28be9d7cae91331b80815d51104207c38a1853b3fd75c0c1f4e14fc8
z56cb501bbdd3779b697b2715c4d295ffd9c58ba61f6b8d384a97e57dd0344573a121f67fc8558f
z4318d13ccc441e94f47ad4db118ef359fb74f10c51605ba78ec295be44d8065ca403f842a5b050
z7ebeef53dc4470ae2da80668a0954c694de2fef292352a051e3b635be55972119e899e63d23165
z76c68fe9a47f446726cf095674426788e64bd315151f57ddbf1e51d5c226ec45f5053ece64b6b3
z1946b505d36b05d6f45281e1422645e3d425e6dad8e33b8a372a6ec7a0cd45a6e489078ea1a5a6
ze41f58cf3fb48aef2610718bc9533302122665c753587e18bf046638879e60def260a0e819f885
zf71f5d730b1c1b16db05c758db9857f4fc36d302ae3b445e8d500ce0db6376381c5477fac6fea1
z14e8c2a3478f2a2a554a17a695b31f7b7959af83ef6947be5fb1a929383aaf4a7219d042527fb6
zafe0fdcdcc4e12ba30b1ed208bff8cb726e3cd3014bccd383daf2a44568c0899770e556d08da70
z5be523cffbfe47d789228ab8f41fe2fec76e2856fa6860303c6b76057e811287818a8d0a1d6e02
zfaf194e9a6f1537aafebd07b38172fb42803aa27cf3b367583dff1f82491003bb561d018be5ce2
z58c34e531f7e4d98b25f9323f65e8559cb312c7a437d6098aad162c87a9f190e57d61b91cf6e00
z7f83dfcf6179a74b6742a202750ca7b570e44dae49a178238b5b7306e5510f7c42e6b3ad684c47
zf6d9a4de72aad517a2995dc9833402b55114c2c548620db36fac68a1e423cc19ce304ef46be4db
za7e1d75a491a0d7ae8b40a65a274c5d31b85da1d2ba14b5e09df20a4fa55208056456c05fbab17
z9b3f87561f7489e20307a6ae6141774c87b12aaa4d60ba420825b936d05a6c0d7ff4963337c95a
z01061db963336aa6ae0ecbfb490735200e0ee927dfc612374f3be3b9efdf67ec0f06626e6029e5
z7f004f68a9a1d0c32f2abdc06ff2b0733afb80e5abb037b2695773423980ba38db8200411261e4
z5cb861812e90fadf556958def26293e81252e8f71b0dc3bad9f2dd013b64f0815a939d31a08523
z3286436b6def2068b4239cc84fc700fc7ca0a0c60ec19596b2a4daea1a29e950eb1a0278a8d6e2
z124cdb23f0a7507fd27768d30c3238e231965fef5f015e594a34598b2b647861c34ca38b0e5220
zc7aad1ded61d416fae04204222defd5e5aea2a1e5f1a1c1d3ec676adf2521b7ec497f15cc95072
ze20019bff0982915823cbf29a6033e08ddbd1cedafa8821c5b54636c0095c530005adf87cb8144
ze3495c00aac3422cdbf64360ffb2bca9960be66abb95ecd40f8ff06ed55e5d4d464d42fa4f9a37
z59989d0a73822e399d52bb59bdbf44c41776e1ff0893b813b271726b65bb02589ba07a71e09e8c
zf436f1de033a925f2913963c2667a28f902effcfdaca12b442448a928a4553cd5d0b0a5afecad3
z66b31f15609af1837d0f2d946e297f8e6721743383f95c117e0c297b603c6d8f47b4d7b884d524
z1767e29f00dda4123fdd24ee526ce8605403d9910747898ebeb4476d72845a69c9fa4b640f9777
zce4be292dff51a66a7618b5027a5206a9f63da50c30b87f2a79f692e7fd4154284f66e47693373
ze6aff27309f20ff99846fefc6a9ecedec3ed88acd716aea895ef897e0ddd6bcb6773025fa6b7d5
z30e609bd42e1e89bd8f7a9de1a72ca45c534afc61de9bd7ffd2e71952164cf080ebe9b2106a646
z18e7717945f950bd3d81bddd0ea67bc4c225f1dddef481dcd8ae9c52346e7c34df57d1e077a4cd
z6522f9cfd8a50c2e9799ff14e492971489a52af93516749b772100636d3ec955d54fc1666c3f6e
z7d17da381b766c32705140ad04ddb3e5281afab65165a102e9addf3830e35893a2a5c6c797d689
ze402f6afabc51a6916235a0f31e71c683ce5994173ad64fbda7a3044f367c2dc70af863ecb5e3c
zf2eabf42a0079ed455bff95a42e8da042b84bed5cd6849d3d58fa3d16de1c9fb3354756f8e417d
zef285e0cdf8b76c61168736be1f4e6fae9a54a64051043c6e332ecd7e57e8caf6df519500ffbb1
z7ed33182d9f92765ddef1a198ab708617c6e21ee5b5a9faa548b4977427f0f0fc310e10c80ea2e
z97f30b6c443844dbfaff82902bbd217b1f7be54f7f873a595fee6ee090e42630d02bc6e782be3d
zab1c5d59a7704fc62f7c05a6
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_ddr_sdram_data_checker.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
