`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1bf3f153bd631387c118a296ca10cbf0349426
zcf2ea5eb241fa84c8ecbbf7180f10eb9ddd4966d421e6ca571b198ed195474578ea51160ffbd6b
z0f73216703aef2bba31d04f6d0877540c760cd2535de4136d5bd4771107747c34c07fab3aaf6bd
z67c5eab3938266c996e67839bfd448cabe88dac2c17438997a3ee0a0543dc656070eb3dfe7c0a1
z57e24e01799b1ae1652a0133882b63649084f8bfaa3118d2448218b5c4119ef2134dee0d7a292d
z80c07e69250e6cb0856a07c01efe3f869b070b26474ff619f1ee9676ce10b0179ed9855d8e02bd
z3e17bd42a654e974019a7ca7de85bfb3ac5c169726f832c6b918eae789fa38ca70f5115a2ee7c1
zfb52b503ce6ce35b7dc5989bd64a1623ecf327040db427ea1518177d8423992586c82ca8ef5783
z63913b3bff1336b6e3685dbd63eb482c1694cc8e7bb0121103cb3f779f1afdb33a5dc4caad3fca
z3ad61f9e6798c7fdebf82270990759ec1a4107e22a744a216da0132a2888c982add83dedd55b92
z473c98e970f0292cb4fd1c6ac764bf3440c9b1318f8d50bc16bd1ece42ab2031f5f07b6b7ed034
z152d8af907ce476029716b8636a467a9c888befa1aad211cc2ca016bdda818d13849dd75a5839f
z6756c38996bf1fd29a8013133e827e1284f810b72d3e06603ef5817cc0da304a0a5dd1d1846808
zb2002160747a6add56b167a6c1fa52b0042118737a50f78acd43c7bf6e31a7ab7426d6848fb30e
z2fbd144a6372a039014a96b7d0a0f6c06013328415921a08bdf6673195dcdb181bf134f1327496
z7b875fbd1547314d474eca97cf3f7487bba890200e4ad7091b33286d12a39b1f291270e835931a
ze459d5c281d596e2aa36b1715b202d3777577d9ae416d9fbb86c58f4a29645564bc1aade9ce21a
z571168b79968822a475a731b4f6e290c8940ed32aaa35a19260485728c546f58e04fecf938af25
z68efc58a4ad673fd64c96c187bdb5a8ee0b31e18f7e7c38cb934e903ede0137723e43c24561fce
zc1f3ff874a78a1a9b91c53967f7cb6fa8de59e460ec73d056bd2c6a2fbc432aac0cb03e7898967
z06c8e9acb92a5beed4781f6d6513723dc52f8bdf020dbd6b9e2b5df059a6f9af2c5e68ade86441
z6896215ddbc5940d2207a63fce5e9f6a2b6715514952d68b1b7c1d5a7db26e7c3635c78a6ea416
z5093aa178b8ae0b7caf82146225f00a5677b9eeb32d4e4c8c675698d895747bc985b6b0bcc88ad
z3dc42300c364a9c3672a10dbf6cc9aa70893423158eb1a8315b345de133135ace76a956ade7979
z7a741749c2e45ba721a0702d813bf1c42f01ec8b8d5a536e01113c346a0b5700348f073b22b986
z5b84d17e4d3be8cfeae1a9858f26fc33c2385cb69693a3e3b0ff3e925de212a29ebfc1bf680406
z630a47b254fd3c108909a227b0806bd4da506abd65fff8fe955bb6f6accee14ed10820771b1f3c
z12538f8408c500aa38225cbd308569a60c2806523476479a738ea3d51e0121b3d578d57fbe338d
zf53fb6f643a1780ab40e05e9d1eb86591ddde1d3b6fc17feff07d4557b6b38268dec4a24007507
zbdf0353b73bc95ebd0ba3a073684a2ffa529bdba0d085b52339e58255d1ee1db22e2d40a23a791
z6dfdadac512978bfc4aab5a8b50448a8d0cb69a60e8a6ad0ee0ee61767cacb0219acf0530fd73f
zb38f737d59cdd78fa665845f1ab0d0db1c2939f7664e6fc1def54bb0830aae77853165686bd8d0
z20d845b7db468716953901ef0e185eb1d9df67c35f800c49d3739d67c18d03d1b7d83ee992647a
z8e1d39941253c2325d39b6388dbfa7fbd4d222094d0ccde69c8ef2418cbdfbe3663a0e518ba882
zf470fbf1b74b82132e20b96c3185a1262a7d06fa7bf2592fc8e5b6f31be95300300caf854ac595
z83f9766082323d4dbdb1332a4b2ed1284ba15eb2c3acbe280589c2cb6ee2df96ef8dd2d0f0f19c
zffbb593d062b535ee24dbc88b8c1920c00e7a756b3f094f568c3f444a57ef171af4946c3b40d1f
z80e2f6506de17f997c3553d7c347105d6d4856152abad776cbff9a42b51eaed23c6e73d784f739
z837d7eff23d3a7bfa68034f1f413b1070f5223561730bab3ae87edef96b04d9272da47f6014f76
zd3d4a18c41dc475c2ddf090e36d5e245fa0443b49672a9ee551178ed8a6ff663743418bd1f14ee
ze30701925acef9c8bbd22b73bdfca93d671809fb59109f0487318f4e45edfae7b35af1a1db8a35
z5d09e710001c7b754293a8ef45e2a4f4586b45b9f6966c77448ad65b673feb0a4b6ae0a8a7c808
z5b36063bfd9b50a5ea3fcd9d1637d5024a88eb8d2d50521ee1494ca13210f2a6a3eee09c3401aa
z7a339a04a3723eff3b5f5bd018b4ce03529ec5b2095d971e042f6664b78048730de792684caf66
z34324ea83bc2224df814242df9ec8139fc0b5e0dd5bf566b63cf34b10df36bfc9e5c72d58f63e0
z7fda37ee04333c7505a7441fbca6ebd46db17d35658042908f29047ae44d95ecd13368e94af5fc
z85cc4076f7ebe0fa5c9b79bb3a3009e9916c50a4a17f0ded7f93917d39eca8eed001e9d3db47b6
z05df5905352855919a25d89a62dc164498d0b15b0a33c7e81f3159b17e7fc12e8188039d168e51
z8dbd41aaa260dd5232602c5c1c11b362d4e17dfba19e13d4928462a6f439e75cedf4e7f9d050b6
z2c8d9fd45c4fe0e365c283ac98c27661b85b068c03df4e67f50c02845aff6792cd986b644a87b9
z5c1814c44b4380d9dccf47dee55dbf763580769f92d2bcccd53d58b8b0ff7ddb2729275039938d
z14df9791e195e6c36b98e3695f4373d24807187e62c7a75361484bc6eff0c4533aa023c86ca84b
z5aa4e5029289c362a38b162d604f8b31ec18c7f45464f56b7f715435f4cf2ecd07ee44dc1a531a
z1a3c2c373d9f0f14060e481490c83474fc6c08d545fed17eea42f9281e846f92f10a461a7b6149
zd75acb65fa3c8d92d5d391f669073ca3d9bdd6a8a8421acd8062d702c4a46e20234d68bc8846fc
zd9e61f6e45e7c58ebc7cefaaf749e96f1996eea327408b6ab5bc3fec6ea5e7dea609c3d0fb331e
z354e594081eb73c8540ecf5dfc521801c807be2f31e0435cb73ac8d799e8be502ed4b9308c88da
z8136b63791f5f8a794bc9f4b56330e1415a68d1fbf53badf2ae1a5e381868cf43f6183bac79478
za2a796cb0409c3c1a784c2ab6bf576be3c4c3ff776a8830a097e7d87ec5d45fdfdb2f9a35d3262
z13f8483be956db4c2fcabbc34fa6819449d0fdd95e6d0c0b36d298a791f000e9d737fa9894c4dd
zd3e3ff7f67ff2f4917a5a169dc0b0ca5786c687c5479ea6c2c5e1d1122a0c5abbf26435d3368e6
z96b87095c0d54a09070d3e5e2157e3dcf431c419dadfbba63d4c9208da8f62fad346e28621ffe2
z98e1c97ca5bb2c43aa05ab41d4f1e8c8480fd3bb519df070a22058732c5b40e53e93765af4b8c7
ze5a180b01d9d2621f37e95995f14ead97dc775a60eceee307e3bfc168ca04d1db3657b3214784d
z134b00d6c8a9243faf50b1c8148a60332b045f3c98730a8fb562f001eafdbed9af3d06fee2f750
z6b48bf259c5df62e721d40cfd34ce3c05be07f8c5532ce4e3e9be8dbf0befa39abadfa791c16fb
zbae084d969dd690c741ea195c154ca3aa02294ac92edf20ee1e9cce1e4602673d264d1d60bb3ca
z15719e0d44338f43c003fcba83dc6fb94d7ec080541fec10bf3977b91d667c17a472e6dfda7546
z776d4ff191abbe009c8cdd84be03e770d3e9d70a90f14abac1a2b2b795aca3b8e522af38f6b6e5
z6debf4c92fb2e971112bb0ffafd6a195159d827c89d632e615ea60024fe8f782e7b93daa5213e9
za7fed547f9c43edcb312ecbbb71d95689d2493ed4e99543b6b4e9f807a968df3db42280494e4aa
z3c08bde926a0a91fb99e84dd7826372d0eec019ede86c2c3ddb2a7687fbfee71114b9621ed09ad
zb0acc565d62a3a43b137a30f1385115dedf682d3d455b21f0819ba70bee4ed906793f0700c223c
z4214f46af5bc98183db91dc9404522932cce1cdfd9ca4349f506e6cbf8fa32a6a0efd390ad6476
z2ed2db95b6aafe832db4c7c6eda470945ae68658703b0433c5cba06d27d36e910b77c77e3e850b
ze5c711e9bb72207131a66ef372ee207ae901567d9bbb328dcaa73c1ae537954a35663876350f87
zda294715523bd98fa612921c8d5cd71a2e6e4df7e1ba6096e0569ba8497bb730f3eb0e9910a531
z26de7e53cbb2c118cdd20dd4969d71294f64acaf590fd761decde056b0d59c3f6c8e1cd47de767
za18511d68ed0a4dcc7b979060db15a594e72934e81e9f95e3d6cff75384227d3e29f288a8fc58c
zb4aa5c2a0d966a9420f40b0c1eec7b3e71007ed60a387f4d46d5d546833206d812221fb06e35b4
z17730db1cf3a6fda35880584f886026ae2c465fc241faeb56943e927ab567e6bdd93237e5cc9e2
z32fed8c2b6d931625e56b1fe149534e8654c13a0135ed684064b3e0fb8fdf1817e7bdff1581caf
zbb72ba7bff2c134ac585dd209491c2ab546158145a73aaef227ed39f673d62d2e6fb9606964f1b
z193f3cc924e45273c83b440877ca4490af83d212c5d40adbf7cf799dca06e1ad6f5cba3c99ace0
z765c59f366ffcb711f88f05f84065486fbec030a3c2438f7cf631ebc81d4617068863bb8800ef1
z786ac9104db5e45116f3e1c1d4713590ce46d36d0e62a7b297a8e5930134b7fa54c9f73a722469
zb825299d3c29db9cf3dd21270e424a8b132bccee7851f00727ec32ea4774c726fe537d43f4a58b
z6d54ec3ab85b4e26063d61bdb10c29d552871fafd661a02ea33296c411718356b2d84b228e97df
z10db62076afd0c3a4cd45d687c1def5dfc810caf143a603a6fe9efca2dd3e76c376ed5d1a08698
zc90121a85fb6c1b9493f0062fa76f17392643d8f56cfc569921bf359188227779467701402fc7c
z7a938a54c383d191ac63b50f53c365c4a7fe0691cdfb14da71f9734966ec2e9dc91a6648d70c6f
z99b8c9ac52b9d9b96d3d0ea31b1e39e286f7f2c57ab6dfcc8ea5ad312cbd6cb63a25e5cdf18b97
zb10caa3c93e625af6d260e04226ebd34673452a9ff1b6be57c5b5cbd67451ccf868e1c1f837903
z53315ab4e1ca1327fa54221caee6e4f5d48d0f3ec1109baff58a2e6e2726c878445ca8636bc32c
z5899cda09cf53ba2336a4743b5eff11d427b52646ea833e82ab0d9e2a562b6c9a19b953663929b
zadb8acb6e44ada4572375b90dab50f0abb0614890155828660750d31715b6ffd8d6bdbd1a1961c
z575383c2b58fef013a96b8744fd4d33b85ba905c97ba6058096f6dc3047668ed66b3dc6f1767f9
z626440d49e3fd184976beec05e1de2b3dd9441189e6f41e2e6fecca71f2cb89d51a1c968781cd6
z4febb6cec42b998b3a97bdeb5c4b2a9500b564674ed71635c903dba9b19640c25327307be584c6
z5d7877574624c30fdbd15c8277b91289bb4576cb8e9395b465aee2542294f535d7f1e34fe489f7
zb8966182d480b3456c9b0499d11bf0d509e8fb0baa615f5bed18f3d6a008a61bdd4985588bc959
z4bd8779fbfd93c390cf6c492619bed20a0a476c5a0c2372d13ea85883a24798738dddcfa3f7a54
zad0477860f84dae2ca6b439864890279faecad94c72fa8e0032557688a376aa66a56ff952f7f98
z6949d59e4b6f68662fc628db1becc740f6fbb895ae48bf26d57e679168bcd000f82749de61705b
z32017c93252292c718ed939c9e1ac23a5feeea6daffa9515ad17584fac7475c0b5ef3750fb83c9
z576955fc6e21ac0dc918f2e7c0a7a2e65ad2eaf42f296edb90821807587f2b89b8c14b48ea3031
z3fbc418deee47a019c191647c7b06503d7b2e5b912607a40ba4e83f08cb2e070a8dc2010ff3857
z1019bf5e992afbe173ee4047910fb2b0ca03565327776d8f75f1cfb3b4c1d2710f20bd17e73f94
za3e65b488a2856608e61518bc947eb9451ae640af5d080941196a000991f1c7392b302bcb2867c
ze79507a63897d8cad5d9b748d6b645e8fd5a7ec7000eb0aecc06e50aba0fa7a22174e4706a51d0
z31b94323a43d5ddbaa94c3eb209544bb1fc0599bcd3d07c5d9d8f72a223d4ef27f020d3fac0602
zed1b5abdb1ddd2a27ead9df4d35d9159750d2710a4671a1713854ab947812f634dca5da9b588fc
z04283e1119f9e8ad74165781cbb306d6c70f2f3e15cd0e888930da914724c2634ea2f371c87794
zad0fa7c864dcc7bbcedeff285b702948c308246455d6a918bbee4a434891d0bbf9ff1e8bff5cd6
za7d3f3f36be36665f719c95eef7071ad597cfae86ca6fab033014f45236ef4745584bc44ae61d1
z656f89200d1dd1e91de9424e08b66472378974d33566e4bab7a9556e5885836e0ba6ef12311007
z6972ebe4303f7b8f0df4700de8cd3bfab180f3a5130f3362ef7ba701a7b607d7fcaf89d5aac240
zba4a1cf2c7bea9980d9fe1fe0dd16f1d84e047a87050f045c5232c2af01f1224a7701d563d14f1
z75e5e9c894bcc0037d8da181994950a7bf9c52252171930c2b9e6a8a1c77eb52c7911d7e30d0dc
z1f239da3a9b0f799338847feb56c15d567343b12fbb8f97f8b166d635732eda1f44070e25194f5
z5be2e9e048bbcdaf595fe1c2c7387b4176305215d0f9b38461eb41d572d2c7091f41156cdfd130
zc0bb842d654e82dfa66c07401d503e8d1a9525421f0145cb20d4107a0cb116cedd53fdb15e0bfb
zee7dc7a7873da0ed71a2c5dc61b64020e627c6c209ec0d478af19c14eed036e50e0f9644690c60
z7c6d4e3b361ea94b2f723c531f319af793bbda35c5d2188b3a8308f0fc73db134423a7a2d71c88
zdcc7cd224aa0cc193173df92222503ac7e3d4ced4e1807d31e524565df68d86690d99323f9a67d
z3ea0a46db69a84760e532949f5277e1b97d663788c7456610ac698f7c7beaef0ec5cde2c4b7a6e
z11de2468b899d4a47d27446bbe8f9fc2dce22f41482b71153df043ba1638c7eae30cb7a6db3da6
z9db1104c192392daa4fb5f710f639eca31a67f33fbe0dfedcd25807837ec31d1cd556a415d30b1
z037554b83e5104b311e7e94de0d8911b70067163d390ea857542795f804eeb68dd16d22605fc9b
z417071bd43fe17130e5c7d37122bac347b08af811775cd368e1cafcb0899bedcef719fabe60671
zb32c99fc10e08c7412f9c1558f086241bbbf12484bdf0dc7b03f49ff61fc32f4971fe5493755ae
z29d15c1e47aeb33004f86fef41f6def970b5cb8c9f8317258c4fbf1e373a0a7f65e26c047cc89f
z0f75ae1baead39cc3c53b550fd0aa185d03b6bf57b724477c043dc64b5464e595a049c59919041
z5aabcff77db35d02d1d6de6c06031512eb3e2aed327508b8f67c292a8868ba939c68e82c996816
zc6494be711888af03298725038039900df6446547df4082708731e2cf1a9fcc6c6e0986c3c007c
z807ee01e7dfae5f520e49cebcfe75cfff9b29e0f10dfba67608480e8868e2df5a769119768a9c0
zf11d0e36e4b8e99c0d95c0efb74cd9fe65badf1e96743f5b833920e0ac0a7f79d72e96bc64fac5
zaf9401b14abb5090286333af5e92b8db98ba3b4c9fcff2f20b49af5078974eb7b151e01cefcfcf
zd1a9e7e8c90f6365fddbd3fefffacf4313647fea973f64c80f79ce2335a8361f6dd1c2441bf53d
zca82075e2e2a136ce96a9c1eefe3f8e02f375d73648d4e8bd76234a72adeb2adad7565bd7a557f
z7338d87c6ee6f543ec64a46ca293eb594c72b7622a16c8cbd83bf55be65245a37154f0db6cbcb9
zfd078a2fa700c0ada4d8f5a6192a3edc703cd8cbe4616671aee44a1024cc08eae7b1e0d27b763a
z15193e568a82f711cb5bd43e3a61879a75b94bd82c437bf111243ae069444f783a1fd85436d12a
z1e3a6bea966903cbe49ea2d53b780ec6a05812d5005f4ad226462f134d90a76bbb372e4abc865d
z993427cf191a34a483230100b0780ab8e8acf25b2f735473c6ff667f0b32adac078cff0bb61360
z2c8365dac0941b7a11f837d8a4c9baa7bdc7452ac871ed7a73606a3be0c17b49f9e8d5b3284ded
zd8ea3915d582368b728010b09fc7ba8ce8c38f4767f2ff66c97503d7424d2cfb51de191f0b790a
z806c08e7c569ebd206e4c79068567a7fec144673cbaf48a5c30ed5950efc2cb9dd92233b33d4cc
z7dbbba527b1cb7575379ae8b759e55e972b156d340226932dadf53d2d7f14ae76673e9619e0aeb
zd12a86767d6129c6a5c23995e0aa315b83972ec0425e39ee0a92697c2aa0ec011ab471e6582ad0
z5685b2445752a28ecce96b2f82d19013fc8bf350450faa3e3097be94f11debd3af09094116d7f2
z60ab9b8a09f1c835b3d3bd4e89e1fdc73d119caf1c0f867fa942a3b71765f760f4ecd30770668a
z20496161ccbaa4f186ffa9fac8d287b6f42e26a39d96190f762e5c2e09728230a8f131cb872472
z4034a4a4befc4963b988dc36105186756344159b628fe26437ac6fc2102d37cfc20667aa0f03b4
z09423f940b5a310eb5ba3ddc57974123e752e3ab85d715d5bc00a69def34e4bc6a53a61f720c63
za5efcd2f8f73e397015badd8ec646ef869f12d5fb2075c251d2cc95efe5e76ad54a7f3e1d4119c
z6b8a64ec73358b1e27556199f2417a7a21158d37ab4fa8c07eaee43e3e00368876214817479049
zb1e51a551e4af1b0a665763279de16c9a4b9019fbb67ad33a7a9e0e72df495afa0349363991fb7
z5445e570598009bf79993ee5e884d614bf7b4a0fe51dc566e182980ebfdc8657e3c13680cb6a8a
zad0961b9c12a78480cf750a0dc53791fc74c55718c84d22b658edc61bd682af835de7c7a31561d
z4f98d7de9ad82b6093e50656f2fe58864f90ba1c29e095155673a99aaf90cc3f00fb0faa054d4c
zd655af6d2d12f9521fbc295e30b8f189223653d487cec96165a250096af157001ba45efc6cfe2e
z18e14617fb0f11a324ee0cf5bb59d5fb54b5fbacf0d1490e96162c4bbb02981ea529a698564a14
z5839c201ef0405403d962d0caaa5015b0e7bb5c6e85c0faccbc62f0b267a57a7af110e0d403b60
z0b5db8e9d90c41565ed6382a044862374e8af4441cb98ea3961882f55d0fb95dd56634283b9a4d
z2402f5422420b6930d07a5e5e4c5bb0742d0ac8fa35f475cd864e34cc5d0e2936a41ce64920a8b
z1842a42aafd90098f8afdc91f2c4708bbb8d4b400615bcbbb7c89aa47ceb77424cefd4a7f9cf0b
z400b5b4a9d0fd0c08c641b77fbf9032fb38afb68ccd6624abd74e77f6d621c9f7065e6a3f131e6
z892b5eac6022b2b4924b1f12c9edc6ba23ecf4785e0fe30a90502a7770803fc46769c2a43466d8
z5c97915aa79dee5cdf76e4c8c77669238466124d46ca5899b2cf2327bc06b6f95757baaf0e07d4
z3b521b5f0600c7503c04bd27852e2b0c6ffc83cfcbbc2f3068ed10da451cc0d19cac7077e7ef8e
zdf05ac8504db090463502fdad3254f2b28740be4941916971373cbae45016743cd62f097144a5d
z80057704fa79decffd712c6a4ce198cefd9b55713fa24f945051dce387470b8e8e2b0ad260c999
z90ad566bd7db4a8d4efa40c79bec132c81f880c06c1c7d400a80816a3d0aefe1b89844db526e7a
zc1bc6c1a9021a106f62b812447a2dc6a063f073be77084a5976946e2995e2205288d5dc23172aa
ze83000a79d5fb71417625a29072d80c864b787edf0f1a850f707b3a0e852abc6118cba2b639c67
z406e36e5d37d31186d5bb0f7a1d6f8a85e926b57cfb19b0a726209f1da53a352648209073a5dba
z1389ec66164f515c1b5c6b63c4194c0e0959320ed7de602cda1a18116baff45c042ad544382af1
z44693ea56fe6b60d90563084a98b87a1884f7ef04615a37a5b9460b5027d2ec656db3c5ebed789
z94d50b4ebb13c86a304bdd5a1a400fdf31f9ac1f94fd304cd20857c1430d52bfbb378cf96f8c41
z11cead8305568aa03e7efda5b7c23d4a6e1241a6b1e50bbd1f01bbe3d8be6c34e55ead8982d409
z7db6dec0d13a348aed3652999482eef762dee337f5a645e27299c560123fc52e3dbca294c08004
z64213913140d71888e4daddd6b2e99e53b9e060f3c0fb2fd9a2afa096c981730b521020d93f3e2
z21d6aa9c084553faee287792511d805a1618079e80b762e42a2d3a1feb3ad1eab2f00130fa8f3f
z0f3bf5f0ca2a522dc705373360b3bead8ee7213d61d93b08583c11dcc41052c8eb5ab8892d2d7b
z64936be7b58da9b44ec45c5bfd3fe9ed1333b2619725e318ffee08c2263b0281a7983ab9b3f82a
za5332e546d4ec17cf3efc1ff217b21c3ec1940cabecc9ad210be983788d80abf9ce891e16a407d
zea0bd8e6d3e58825d26f7ad8d6892c0a1040813676277dcbcf4dca0c9154ba36842e00238e25a3
zfebbc5d7d439893b227e889f96edf70e33e34fe57bc92b3453813f037ae7b1222e552759957e9e
z9e3e35ea664e6242c5d2ab90af7f4351c5e232dbb250aa15f66ee59b864826e4af644d4c1fd24d
z563cce3a476460e7501139dfda056e4ae9f9dddd0110a84145daf515638837653ba7e2c265ac1f
z9971799bfdd53933d556df4792964ab44df0d192cb299923b79ee221062f2d2a8a81f5dbd44dbc
zd701cccc97d42f83fce92561eda1e1c8092eab2497674270d3914bacc3bbed38c49e90843ea271
z56791518e769033da3d739e4d01205177bbc96d91dd603fb6118b0c5f4e63b569871236b5482fc
z65a48daeca3075103992e69d178c7ef4f6d83dbe82e7f2fc080202b7fefc7806d728de5ba49470
z0eb99ce72b766a3f65c622a54221409ee9646fca81a83393d8e99c98c8550e8d39747d72ad9a0d
z9cee1c545e957e16b15bd5233c5d93f997d40705d78d370227ae5a64a661bc4402e9256588fbdc
zd4c50b55d712b1a1939d156a2914162a323686b06fbeac79749198330ef08d0910f8c27c5b4332
z1ba2d802f7ac74b02e35f9ecbad4108e1459f7343bc874f2e5416fba83fc73bd57055604160e92
ze4718712a545953b23390f4a85b2d5922f3fd64b4974798ec8ed6e9a78b980972675f464ad670c
z6667bc35b3e7825ce5cbcb94b5a953f0246670b60cbb956969afa3c820ca5bfd85d9e38f9b68ce
z7219157abc704064ac41e4ee15f794df512f6d02d3fbb6957d210dfdfacbbac213eb36fed43644
zb575c7f244e38a4559f6c475f809e1bca99af21e6b1a98d53c7c39f1d2d9cc7888c32b82d3471c
za66f39589f0e10996d4fa8febd8e3fee3077a89aefc65d532ec62edb15e4caaaa9475cf52ddf16
zd6296b42e86f188768d6c40afa350bca3159d03135eeb5dfb8f297ed795478fdff0e1e75023bf9
zfe94ef9410643dbba23937dc6e41f10f07af116dd3f1cf9c0c23502ab1eb526bae77d11cd7fea7
z7c499d6b460b00e1152d7d4e4f2247e722b81255b834ea963b742dc0b9555a69b52a9f361bfdf7
z83756594dbb09ccd0a516962738ecaf0fe44798bec1d5328971c13ce4a36c94debfcc3286c3316
z60b5308c6f4a0f7a961e390c8565fc148ea96140993e6e2befebe3724df4bc04b803619d6d0949
z7b1cc44c77c7757a1555f475d99eb6a0a2de475c1e1bbd60acf134e1167762e696ffcb31a11c9c
z5f861c2ae281447d5be234d6573e1835c539e88cdcf8fcc3b9f3461c69f8b3304a5ac49f9cb541
za7c80e03fb6fdedaa7e8bdc1139f728ba9f2867702949da4ec58fb0fb4cefd223202820c9cd612
z81d67d6cdfac0af61d1bcc44dd7a52c1f3004598dbc3ff1d831a8767d52ed8a295341e329bb7a4
zc7218e15aaa3eb52db29e2e93f0d2487270543569f3081323bccdf0513d3bef43824ca8ac270db
zfadd9bc2164b72794953770d0af6ad14cfe66646c8073908ed244c7923bdd4783d659c2d3ec5d5
z358d58809a39534c421860d88edd9176a67c0072a912290e7dfb6324378ad6893e37664a2e2983
z92cbbd56f81844d7a0c54457d7446e462a8a77aa9c0f8254d676ee896c162205df6786dc42686b
z147146907589406ef49e0c7a74e9cab49a9e8829b82dbc6dd1650372df8bc92c81ccb8ad7a15bf
zc19da6dbc60b4da51499b8099a13b532bc168d3bc1755a43134f9f5c1a572b44361f21ac31f4fe
z4b6b782479656d3e3d6b6fb6cb13f06bb2751d1c50d5ab33b89a074c67b1e0c2b818471576feee
zf04a09b23797eb46425ca61d820bababac1b5537fdf6099bf753a16a5509245f9bfcccdfb01e7a
zfcb8202178dff0ac1117b3aace71f1a3a9e9604d8597d432caa0d63a972ca3a3cf72feea6cda08
z3ab136a28c8610da86a6720b59eb595fc0f2ab314c85889ff6ad1a093af7de0188a09155410a63
z1b121fdc7efe393609d582a1c0ca9931d6758ca8191be72360feb8127bd26dc77761e12412a660
z5760d725e9b5185c782ba325783d15a1989de26b1608e2a9a72642d40f1ff98ac7184c227ce67b
z874629e72f7ac323885a7541192a67382b3b0bed88136b45e4aa51a5856abbab558e3c1f7002e6
zf88695a63807374137858e85837e45757ac348b44e93009bfb7371e47a2b75fd8a18c7472a9084
z2de9651a5ea24ae608bf22e47060e230c3c4b5e95394516521820748e5899bdb36277c965542d2
z6f4a54c3c9084acf615d7dc5a63a883387fe0780be263b935ec86321af72a33de22af31729ee2c
z52273f4648db3987251c2434afc4d1d0efab65a44137d168cec39f201e15b43445d7672cda156c
z176a4afe7c549a3c33e2d2b41351ba10f73a0e0bd7a948c80f0c15ece6597431de9f84a3fce102
z0dea38ca1b5a5709b409eead23cd808fe98fbc2e2c21af7a050e4b3fbffa605708d72982eb3b6c
za179f9318e491850ae259cc2a1026083d51b1626177835baed74aa503d35fecf0bf88ee7cb35d2
z91578b3b1f9c08d51b28c5cf9c4030b40d657852387c531e523879d88f50fbf20d7aa73e587b8f
z45120e421c40c9f6512e46c53af1cbe99036008e34517ba02d35757b6cbab9d7beea9f4656c53d
zbacfc5bd0351eb7828c190e0c9bc1c6a661831267dd9f05b4bccbd676c28a765905c7a8a901b26
z02fd9ea76368c0d2a0f658b516703ef3a5910457ba018049e8d718106487cca75c2229fd3ad593
z74ec568b0642d176bfaaab68ee45f9e8df41ac192ae6d11e1410a889ebb255c7ff78f9cad06a54
z52e7a4972bb66ce4e2823e7d98188051f3f1e2a8362bf69594d8b8d074ef97fa21a3d0ede8191f
zebb8c83e5686bbcc0d5601af6cdf2ba4b508b4205b5116c029dd889aedb24e4000f10526d6952d
z680271cc762f68cb5a5367a46b555b2f87b11ec61f8e6c9c3db9ad623e946295c989499cc11601
zd31124aa4d42fe39af3cea6ca157e45375c1e1af1731c5bf0362eaf115d36d0851dccea3c31c0c
z28fa24821d8a1c2d49b720746c679877b22c4d4876c7f564fcb81de906fbbccb97b428241129c0
z8c939675dfb5e065ed7e7423e4179692b35b197818ebd670c134d39de3a4ced6028e5b824f1fc8
z0bd584541b83a201c5213a9f15a5bb96fd258e71c1ecad79a2a343d51ea20f476d6c7740fc59a1
z11b010c7f8a85d82f5849955382aac2d47af525f85809c428c5b75a404d7b68758f7b3ef8b48e6
z4eea55392c956716651841816eddb9810238305d9efc5580c04febd809842beca3d4ef71460a91
z2ffe401a7c5bf115b11a86c9a71576fb09174f225e6af7b68880e793f245589baa8142e17f2cd3
zdc5286de7e05d884377734d752cf05a05aac44c46f02d2a42d5b87ea4f44e3e99facca32e12fd9
z6d035150d31fd65f90cf198c2c4d47343d0dc0663a20cb98efd26ef80ae8edd0d876c914ae5e6d
z4c2745e25ed5f3cf6e26e2b048653a9bf07dfd68b110d5c3f39134fc140bb40e0030cc89a14d7f
z27759ffe4a13b4fd6f1430ab49f7e3ec42a634b41b733ae06755b4cf904f5b77cf32b5920cc2b1
z7a2e15e8a946a402e0a8282d50f036052586318a0a4d88502993d1afd01f0def6aa69d014af1b7
zafb3e79a6f5559868e26071fb85307e30db7fc35fdb2113081debded499124e30cf80962d763c0
z53c0c1715d3fae95a789c6c6478c4850e72923928eb9f2f853f17347ad01b93d9a3fba2a245883
z399b89b2cc9a215e4d7148699a4840d2de87cdb2f8cde27f1d29d1eb95db150ee02bb61098de4f
z0838c742b4569507eed433fc4606b54aa93ac16138ef9c851b9d330040b723e937b4b7e3692a7d
ze167710cab987d761b4eae19fb16e92b8672ecb738b7b22e584d896d67b3014f2b74e21c2f894c
z40fbad26832704d7dcecdeba9fd18e183e9e57e3f85950a66a3e8e920adb8a034ad59308d5e003
z5332f0ddaeeb81137350d9b11f2ed8f3b965eaee654b22faad605aa06e886c66774c84b487e4ca
z61d9b9715bf74ea8da3fd8a75851932ed5d83e0c5ca4a9850e7c9d96025a7a9d8342fed02586b9
z13b8db192ceb989e027b20dcd45fe82668cd8c68b407cf00f8d6f215f48ff2cd7dc8d254bbf75e
z7660907201eb716fe44ffb4d105522624ddfb3a2051f85acbcce1cf62a2e13a6f0ca665eb996e1
zfef2b613bd8c851ee08398d180656838382878bffdb738395e8def6a430a89788b5760866466ed
zfcaa347e67e8121667e7bfd50c96a8384955726e21bf2e73c62c63d2107c919c77f86573f20c8c
zb78a42b8495ee8105668f547999f2708e0dc245123bb15a2d2aed9b02731fffc503ae45c62bea2
z902fe007a98ebba331161e9075537a6bfbf7618e54bba6077a8dddd4ed489bd76cbcec6a9376b9
za23f33b4cb46548eec9b54da2e3011ab206999633512276067708cfd3fc4762803651a22993f8e
za70e1dab8197aceb9260f079a0dbaff2cc45202068abf24dd5f9a146d00936f85304249cbfb7c7
zf264399726bb7fc767a7db5dcdcfde9e4a3b471a9f17d4e08bc941bed3d8874afc4222c3c3ca0f
z09521d295d0c668716d13af1053b02dd33644c91259960f24863b52408b02949f47665eac7b428
z5db281db3f009695e669246d6770765821b17eaeea9a1a77eafd4d51e3123e1273900fb8d9a5e8
z2ffe8a62544b025a1fa60777067e345e526aabeffb87e79bf7373a1d3cf90d0e0269f3da10a98f
z668751dded017efa68e500cce7317ab8b7805e3d8741986e012d36f1316de3bf97aa9f7055cd58
zb8e8ae6469279333d2cda8a8022130818cec5a191a9ad62b0dbea050157dc9f518e4488b4d3b7e
zbe93783b35c196f7a9dd4f3bbddda790ec3e6dd2b9471e34878e764567480098140bb38dbfec42
zc3f94a8c78b441ed190fb179c8a2f915dfd9572aa064e1a905dce430018ff8ed956139e4cb1544
ze4fa8c994d716f958d5c486111af36e3c24bf764010919bf66e97756331fd4601290a9186532b0
zc0b8f4d605a836a5817d694cc470a4ddeeecae5c4a7b50999533c9c74206513048222eb0402d23
zddac2ac51dbccd584d462bcad76aa3f4b44721a9cf0e6f108eb26f64fc3f0690344af95064a81a
z426d8ad3dcc9b49916949bcd100c63e8ff280e826dfbbbb2988c814e2c1de62b95f86464c590ab
z298719a1cedb156dd9f8b85ddd3c9a8df27650bb1b91e97791ba71a6960fe14036c236c3b8f2f8
z874445fb6a07687b05a9009c6e7811d570782e83ceacddc710bcd1b566c1aba2562748d2efd6e6
zbdc195feb9e2d52f8319cd88de0189f01b73601feedab2e7e497a8c9d46f717b30f9ff2893b776
za9f4ef26881f0aea6d2c246bb052d7bc42d716c622a46593fd863dc75ed9b1246f93c71b7be49f
z9c944fb7b02db03cfc84c5b63ead851379d8fb9ded0b0eb163fb8c179f1a9a48173aeb38880003
z46b2f5f21315baba0ff145a584fc4a757862bca699e63d5b63128bca315a686cdc9db85b024267
ze145416f58cba9541e35072ccef3f6dd769d8a075f72f8e411f16824389b4cf909b1ccc3871d76
z2d7f0345146720cc13db66b3092d12c3be4cfd32aff0a075e3890f186b9589260abc3d4366727b
zbfa03e8fdeb0bd89c52a95dbb798679a3f3f0816b6a9a23d0664b58769c2a7676bf0facb90aeb2
z818533ecc035b678ba86439281bc25e07a134eaf5f55df1fa76b417c17e207dc816041fd1ffb10
z3ce262bf1bbdff9a5d6cfcba67c2d6d41b946720c78855cbf058565d5fa253bd08c9460ffc7b74
z7c919379101b1d5d567f62bb5ce69559d808000c22f5c855886bb3556c6fa1ad70b251840564ae
z608ee4b5cabf1655ffab3edf04676560ab84b82b0c44b3124b866afab99f6a901e1dc65dcf0394
z6b5d47d0c275456a7c501277f46ab99902c9aff485d9b0c3678c48f46a184b9ee38b62c81aa35d
z09a5edb7d781dceef8f8ac93e7f76a6c6dd54ec0c74dac6125db8c99288ca7d71e7c17ca9dee5b
z1a55e6b0b8440ca590fbb0a59e588a7168b188a1dbd253377ee4f21955466077ef0392187ede3a
zd9611753bff147b9796e1a285e2c45cf49bf931aaaf4286b7f39ca3253d895f5d6f2feb0d0c4a3
zc69bdfd631a8f538fa345cd34a6146d9cb28f5e147e18948debf6c0afee67ec193c3958b9fbd80
zd38e994b4cc4441f886261c74cbe2b41fc6d3211c6bda227a4981dffaee9c43367b94e3301fb60
z3edc5af0c526ed8e78ca2799a7d2f45baccc435efdff3e248126b34ae235556656b95052cc2bc5
z2d676324038fe0b69138c1bd371be71be1b5583fbd566c3e047ed4542d94a6521df0ecde99df45
z236a275a904547e4553848ed8252bc55ced1dc6dfab7a77fa8b4456b94fd0d15a1844033c1d458
z666961f4a85ba35ad9a643ec3df8243e6e108a519422900cedc0b5e83b320918709fa5da523754
z53e210086ac0aaba9d5439a6f82bb41eb271d95376c0ddff58747c5af88182162749029eb563e8
z96a23f86113cfe48532d7c6431edd04f45dc9afcdfb4650238612daece4ec73e7db6493b20cbdb
z26ccf07e4a4fdc861c34d7b4ecf1a8d9738e96ca0908eedd1a53bdf61adf049299b61d377f14c2
z4c38d1704d3c18f1c501e7db06f7afc9453ef05a475ee7e14157f01bdb721914314a40cd4ae77c
z9de891de5e072d90e3e44854a6c551c32f17ee247fee5d5a805c9adc57b00ece6abb2997239075
z9f0e44905f4ffdb244301dceac07a99dca1e6e2d7064aa78a862caf81e71739d69751cc931e87a
z6e8c58bb8298508300d4dbe2e043f458432f8dbc30caa4ae676e16120a02c40615f0b6b467e28a
z703bdb9530471fa05f32e6b008327ccb1aa54ffd1918dec8d7052701ffd4dfdf39f8a413663d56
z6482aa324ed7f8b459e37ec7ba8338ec1b42d1e8698b98da93158d4ca17018034d0a6af0d2ce4b
z3d6a13e5a0cdc6920ead54b57b34cb0d99d62ed4f4e0e8dfddc585a9a9c8d4e6a288a1ca15c558
z0c3135328d2a63087ac775575681d9cec3d2602a568db511183994032d6a328ad63cc73637900e
z65d35f90f0df08b94a3148ac605f5c369858f4cc874f4069d9b96f455ae8557964b553f9a228c2
z58767c3e4f2d2fd3caf2b2b9fe90737d080967cde77ad893f461553b1efbec6c9823df96f415ea
z3cad2c98067326a62515dde0151684d9650b23471edcc6da3a31681f9f42a774401adc5aa74ace
za8e93fc0f73e806d2e21d410332295fc5b7d0b2c643c2ae28e4e5cd70f7b4417fc6e32edf8b3c1
zaf94c5226478a6e52229cacf37e45ca89a037202aa5eced66009426d605752c77f843c70888216
z7b3dff7b54aa6c720f2867d44b471a980bd85cbe3dd7f1e8f0f7ef8f07d4d8511cf096b345ec0d
z6d9799377b23477bc48359bc5b00f05a5d2755b03d86d5a5b66afa9a58b5ed97dfff97fcd9548a
zedb5f4b5a2753accfaaf715b152146533b9edfbfe4267b455d6c39ba5304f59106f08bcac1819b
z598364a86865c6e3a0f6a1a68e74d8db926209f38b254cb6b9b9ba9d307dc323a73dfd7e742703
z8fabecce5d7813bb104e008cf87caa0409eafc0972abc17e0a488827f0f603898cc3ba3645b0b4
z7edc5ca2575cf5d864cb68831bee717a7b96290287f8a4a9d37c3b41aff5686e55ff9db8816217
z20566e83c072bb5ba1a5334522b429e97420ec67a870ecf08f065056054518e08003d622ec86ce
z0fff59c70f8b499b8a9a74ab973ebfd33dae3b27c521fdac4f2735b9832f3a43ffffdbb773aeaa
zf4d04d053a0bc4b8594636f13693ba27922c20072a972d24c465fbfdb2984c1ed04223e14853f9
z33664adb96cdc31a377176f1d05a1088239a5ff47345dfb6de08310a627fc2b35eaec3a4aa69da
z1c7d99139883a0f8ae9b42d78561c3547d9ecdc1b53f644750d2f2957c6e61a4c323806625c791
z8d1b3f8ac19a06b83d9fa1ed175406e0581c378020c96b250265196b2e564e8caca7dbc578dc2a
z3754b9e7079e586363606c99e942a8c8f67f2804485af22238c3c6059a68dc51836a854278c9bf
z00e697c7baecafea21564635d9a2e58191a34d4ac02de46dd84f000912df5d4b34087a3b25c1a6
zc9da5b838d9a3a2349ff4b69164f01b5c3c06843f240d4d298788ebb50cae30070076a014511e1
z2ea0aa40c5597541ab7c4dd01df7d99c13f40a5840b8e7e217e83a5a366458f8d4d9468fcc71cb
zc83a2dd02d52b5fee73dd985edebd81cf7b5e9e50d1ce092ca09b3cc21f1ee9b7e1b256675c88c
zf0f1c694097c565370eee8c130a947f5b4674fd91cb815e91ce6d2b040cc57dc121f55b4bd7ca9
zb2221d3490d15b4e16275cdc7482b0968683b3d4c156221973a9c3cfbff4df9894875ccda4db3f
z11e96de6e55154050dac398bb0c1348563c3b2c0d5d114dc38e8f6a9ae7bc6b3f8519417663010
z488c057626808cfc005704ee112ecdef4e63beffca877d61bb041f00039153cb181c7371a00be4
zc98ea31ab1a300b80941716d5bc8529c57c10cbbc8aa1fd196bfcb1266bd2cf102ab9648b9edd9
z88c703f0a13f86e253b353241a213f18d42cc2a647836d359839528c52fc821898a302a6e52c68
z26d827ac8ff73ab216f9575ee1e92ddcf4818d68296782f6c794bb145b1f944fd6160bd8634618
z3cbf17d39f628da315ab899bd09d347b5eeaf7f58ea4ab66806cc3649ccec1abe10f2179c5e50d
z9648f26e7e9473c21a5b4e5f2b8509a38c3fb2045122c6f9b2b754f11df3898729f0ccd91490ca
zf6c40efe61a6b3bed439197ad5991083c4c2b9ee5d025bb88d52d1d497f821ce31e35c0200e172
z5fa94401d4a4275d5c8847db5c840187f877b78920a2c5459435e4f96e15c00bc80b5dddcdfff6
z43baf0b3cc4e2f4a2730a3c27c87f04ef7a3ba1a531b92b5e2510a0aab28eed4c5a5959f47428a
z0aa9de493bf5b9c379ce2ed28e0e4f4ae91125e9230cb57f7cce6e774be9d4eb61df4c34c0222c
zd10624f7fff4e77eeee4f797ccecc41c23c06222273bcda8a5f9483594afa6e41d50c8a75e6a15
zf07ca42347039b9dbe098e23d0d845ae0ebbbe9dfab5a3496d8a2623a543737bd4702a6265be7c
zac69d05624584dade75bcb99470dc81593af89357647349e5c836968c902a21f4d41020b85a152
z8b16c449f59e67c44942fdb5b1c1df66d2c8d9a599404d59abba5b02d927d25360c359e635a638
z0bded8b421296049ca7509982c829ec80284c028e3d5161f4d538aff3a161ec6d66f89aa6c9a85
z0317edef461d598c6876a408a435a50940442170453d4912df77b7d6c131e97b215951020b0d80
zbc579af7cf41b075bd2fbe88a351c9b60fe357e20dd1954ea94e4e4acaac29bfe429903c3233cd
zd2f53805ef55525d89feb541026c89e923f566a67a7a1c15a43bed6fb3406794c7d6d735247b84
z91be5422fafacfddf4a6534ec74b1546939083009dcadbf500f34e17a62d90b1b1e7588335bf7f
z352ec61f4765bff982f2dbdfdf40d2b737abd220c2b7a35bde111c8c97284bd0c1d7dd66450995
zc0cff6f2c0625090075d4811d230cf0df03e61d45422988000bdcd7c18aaaacbb33efb44271b4d
zba229375a2bd864a6a998ca56323e414acdb7d10004f1549546c952d79b73e4ab7324983b5ca0b
z8a3f3dccccced0f3c06564e2942066b9946ad13eb95385cd1ee15b194b0f19f6e2c6ed3cecf21c
zc19af6c995a3b39cc2a30424020b24a119713bdedd54be5beb83f98c7331c7f25dc5106dc42a29
z6089f7ab77b13a76fd305753cb866a9c245c52c43fd0636f6b2504407f85d7e4cebc28faa5faee
zb0eeb76ed62fd742aa8f1f4a86472647a42d6f6a537f0c30688e0999f1543e29bfddb9b69f6cc1
zbc35420d5cd16257fb3233952e107e63f4a7cf36e5373b99466b01fa60ac7932b3bf0d24661135
zc0ca72082da679885a048f7c7b8c51fc27fcab428170fd83415599ff448420d42c26bf7ab474e5
z84d44a7559561c7eb86a822e567c14cebce97bf2089ac6fbd245033caf16360384401817af33ec
z5aa5ccb68c804d7b4821ec2b317bc29aa75d98f539410e59cf1af2b3a60a505927039a1138affe
z9885d5b18cae473b5fc4d91ac0e6ccc222aa93483e6460642f94f7446bdace00b5ed74ff3e8433
z631de02cdb11059c0b0e17f4b0063097486a57f89ff3d8ba468af1431dc21d245613f7d143b641
z05fb4d3410b6c5dfb78a248ee21f7b02b03c89afa4eb54ef09306596617a5f8b3b57a4eae60f78
z33a7ccd4e4b88028a67b6bbd9e341243d3130f10874369875f3e65710130842f96d6934d077c99
z9321f010d7df6d19b42d2d36d84111599fe1f309e53a24595809c488f71e41b3486bd362cb2b38
zd13724c33251dc0c387e5e62fca867170b8974a8ed383ae0689497d1b5d392ae4fa909a8710ca4
z7039202d70a5d507d600f0b8d900b4024e08250fc3dd2e020adec24e21290b58279cf70df915db
z2573c58a4ab253b62a0098c72b0cd57c2c5ea0c0ae986f631772beb2bd1989260d5709ce01fdb5
zc28fe715a1f318c9f36c7a683626639f4cccc2af9e38942b30892ca71346d88ce7c8fb49a7cad8
zaab9c08bd5e14a6ff8c372e5e95313cae8fc5542c4404d6c6705280275eba701fda87e8308d025
z700db16ce9f5ce1d273af38f480effb790645426a8f7f56d396a8ddd30495d01a174f881c76f4a
za099ed445bf4d9dea3f7d1a92c0154e80400ef2c86c0461c7030d12ac0f93f97457d27fd735a59
zc0450b0ee4777ca5f1ff6edb6e4c3ad67c730b8a08888bb12b2fdb84ba97c0b038da2027f44214
z2340577a6772e96779276bc62f2b76c4db87782a70cd05e1c20cd006beaf58b572b811344ce86d
z8e8ed8fb7e9fe9c2d6e364f667dbe8544255687716eceb94c5bc0ec245d26584fdb69a34d27108
z96bf56408c682efa769bd111615115e7060d4ec65bea57ad44049782eb4065dc6354968a08c7c0
zadd4ab5fbe42b4ab7f3f49720058232b8b75a92cf9497b6976172f39c3fe4c594866e84134cdb1
zd467f86fa6cb62eb59fc98a8ceef21da1bf32979e980d412ecc78a1a98bc99761ed9a0acf76ea1
zd5b35234040ee8a12edad8dfa30a8497a8c3ca8caa78b05aaf0e2f16f86db2736ce2269c3a6f0c
z4f744ca516fa647b042a866494f071f715ba1c607bf899bc21918a138afaca12eb2f5ad8143064
z37c4f06c52814761e47db12525d0313f7688e831a1df3b20298c0728b327f14123eb8a941ace26
z7cc3d93229c518656a8f789d00f6a8a096a26cc52772b940c29079bb5eb4bfa506b19dd0a107b9
z56c9e9a8fa114fbd8e75370b3f944e92ecd47e408bc8b8893aaedd0d39553519b63b46d9c3549a
z6c006a9fc4ecdbc5438b9d0905f1c11a148f0f1308a392d1a5527212b54821f387511c1b7fa9ad
zedc4d746e7726af47e2ff4f7ed6370350578958a1ea340a161f1e3aed37a04665d6a1ba477a4eb
z257a3d731d21a1d1e5bd1c1b81ed6043969a5dbc25d220de2ba8330b875a2719a804d8860f16e8
zad47979c017e47e4471a89107a964ae7048a4e654893cd0c26d4e2dd0499dc335bc88769322bd5
z2cf7e0de6d86513edcd91e931d76bc5a49edc3edf18bf3e3533a20d12cd732312cf9532089ad6f
z72d9e244e449827f30b951f3164b7cac66ea1fcb97e463a1649f8f7879cdb217618b79577c6f40
z03591bddf53822cb11d189a6cd3f8c1e2563ec9b2f7c2002b55605f40b825367857c0ac9702d28
zeae701b8e2d5d2929685587f4f1a5478a29dc9027010cb6e3fbc80b2fc2bd7f1edc0004ab49907
zd80801eaaf3e77fcac5d7f86b7159dc2826755a46b63de06115e0ca5cc702bf283b69f44bae071
z3180c34697a5e753f8b7f317111e640c138d434fb96989e80dc222a089be876c7dc249f4e12424
z2dca9860f46a84b11ed9fcb8abe3910dba14c72188f09b4815356fce634b89be03599afbb913df
zdcd9482d12ea5439d2cd0176262ef256535a350910cf8ef156906a8802682f81f86a37dcf17f9d
z40516ce61e6203135e137f8823186e18febc1b69a3006ea58bd16159046055ad875f51bcdac2f2
zdb9a9d180ef890a600badfce3d0ad1810d579939175c1d4d293c5ce43a884cdb9716fcdd57751c
ze54bf9f8a0104d7c7626d9949783037eb6296b3d1740b559b3a6272ad64333866ca788be58a209
zb752c78b43d5148c710535da67699c81b25b76e1e81c3b2f9db0096ef2de83a9de5018194dc349
z309b71cdc087e171bcc7a3ce6781e2f510869a0e8874494014c77cc69cb8d9c17a8ab3b7db2a4f
z479e933081d4a9252d10b4a50bb409a153cef1eb0ee8d79ad6bd58302845f0145143ee02fa99f8
zfb7407ed121c339f40c6786cd38b7467af0df158b26bbe6f2e0037b111c23e41f9949c307ee60a
z93e7928bb83e04577587effd8107f712b79df419c43c6a2e187a1d7c462d44621295b6ed9f236b
z55c93657644e2fa8b433c5203ecbd65ed96e6fb819edf6b0dafd740ab6b977f7387b9a93a58c95
z4629bb564d23240329e066fb48d0a7061a81f31224e0e5e0baa5b16a0de2ab2f420d6b4be03be2
za266ef7fe4cac3db8cfc7fe2335d8f397bdd8b83c847efdb51969b5ba39a0bcab3f635eb5530a4
z6e2a721c975ccb8eb51d159da5a5f1005dcc523036be7e836391fbd64ec051737fc9ade6084c30
z5c1aeb55c535c1dae76e28a4e213c476c9d830e49e76a0eeeee9f6d14ae2088dfb38a163b9d80e
z56ade343ec5912b7f6f1aa1841595012af5d4cfb866d24b46b91d468469a6a31b5028c69f7be88
z9465b06f133f770e4c07d4efb8ee77d8c24d239a389cb5f9898748d3c24ee502b61810fe670ce3
zb95ee0135d5c3adbdc9358b4179b246c79618b8f33c34f14ae13a7fd73d743826f777fa49b3af8
z8016d25d89185aae697d7b82aa8d66ce211e6e8d965bca7c03c44d4cb95b380f4fe3ffb42661c6
zccef39a77768a93bcfa2fa4de3e6a00a799a003ebe4781554c58a0c8f0803b726d9c87c86b01ce
z2b28e485d800462d7ae314fd71fcb6c61ec7672ee5637811ac603a2682a91ae9046c214291590e
z6bfc0333e11e88d18481d8c15721faaa4d4bcdff7fc006e4ba3fab622b6146c5df534667537a94
z87cc82e1c2a8c47708c8853194da44f325697aa0343d81304e3234457cbca801af34f9727ed972
zc7baa9a5503aac7102793499dbb0aeefb190e1307293996420b119776c9b8751c6dc0ec890ee2b
zd9785be309708a05719f070236d1a58f82d7e425d57526e4bba3ee7c15d68eebd0fccba3f0dbda
zf27ee427d4b7fa5362a30372ecbbedd32be482dcba047fcb4fbd5bb1acaadc789fb65bc5c35c31
zbd58e81f5f599cb8a706146029cfa769ecc0f5744f714183c25e319ae995c1d879636bf721d8cd
z9306ae55b8afc51ef4419b00468db7b3f631cac2c563a4e462b3fcb66de08df118f33c266d940c
z224f3af1d511a7300edb8af602e341f4d94f370b065ce484f0b36783b59e506f470b1400826d33
zf2c1362413533f43c917ba0264c5b31ed834b9bceca73b1c3f118b9f2924eb723ff1b1c3d64d9a
z8d97336b09954f3695510c42eae092bf89b1a8c7d2fc38edfedd11a37629dcde34e779cdf04ef1
z0cc441b8f93e6cea661ff33982453f88884f5529226fe1e659914f375fff39b03300872f415c1a
z854ab7ac013609e46c811118ec0011619adced18a128d36e9c7165ca821c4c4a0eca6d27364ed2
z4407a68b0a81087e47558f1948bb26f5909a7c54853cba190ddd43235fe5b8a88bd9a55e348f7b
z287e77b7a8b8e3f5aeac841508e316e7346e48bba26611931049596f93c3884d849e5ebe798cab
z05b23680e65d089b180cb3cf64af3834db6eedbcef0ca7d24926e857947e3dcf8e1d54719a2d6e
z0e3d4037724166cd72a3f120a0519dbe60d38883123508cacc061794e8802aa2628968320637f9
zb62431d7ce2c59c96f2c66e8e77eb15006827b341cc967d2b8455dcf6cc5882e815e16d0078468
zaa240b7871727b593368d4cfa17bdba0c2a8c1ac1cd127b6e74b15d009b63b877264dfdb1fd281
z3e90b50768ddc925a33650f962d340034db11f29d137138f35b1bff6e58e36e200c0dcb98f4622
zf2b2c6d407a4df155871b5f8504a88dcca1849bf833a5fd0f51d2c3866d978630c52ff76babe02
z31d7da36d5b03a3774f758ceff48f3b2937ccf4cacb81d2fe3e99e1a2ce6d15172c620c8840aec
zed331094ad0011fe4ac7548dbb722b73291a808cfc7c9c0ac7190007eedbe9731379355e837f32
z21c6ed97dc9b2818e700b7d49a1f260ba5dea23a0372f482a52c79197397dd7659bd1aaa51e692
z9d3508c527c385cfc6c08ae3f467eeb599b6b06c4743d6dc112d10f342012af5e372f95d404e67
z42fbccac58d94f0c105aab45677f20a84a1f3e1525cd7b4b1f41fdebb678b4d821052f71aeda14
z9610e008542864b31aed73e1ae1d8a112d458842aff272beb0d55cbd9f121813df4b97e82f69a8
z52e5054dec6ec9b0bfe0a9cbbddab4ada1c0ce29f2dd975f35cf3b18b011407834fc628fbafd59
z2e8068e5d5efd3ad69472cd32c51237ad8b977844b8b398ab41748e60167544423d7ac1761e7cb
zf56bc37236de8b6f98a07d3e76d341ea61c1fef94c76ca14acbe8ea763c2ddceed516cb28dd3ba
zfb2fc2caa562d60ee518663eab8e60b30327f05da01c184d5142aa9e26cf91f2d1dc939c4cffbc
z6478e82736ec0a3d15a9ce497ca1248d61bb33255310cfa6dce00bfe15de80df76e986d6443f98
zd2da3631ea639e8d413550fa4ecb0db43d4ce692b7d29eefeac70610ff8b6470782076ee722974
z6a7719069a9d0b3f0fab03051406b067c783efd106d234de5c6c930d12dba3ebee41ed94ba2d3f
z69fecc699fe8e6da6eb4e7bb9c28b8777c1c702afc1fdd73986483486395521493ae91cb67a85d
z058dda464360cf03a9703da3be18bd656e79e6e6a061a1bebfac3b9cc814892387d2dafec0aed6
zf707a9d7b564e3d82590d75c090906682dbbd7fefc4c82c3ce53e80aed65de1b66544b73a5fe3f
ze2780adeebae0e00315edddd6b02599963226f0e8a6f726961a8a85cbeffad26f2285c2d010300
zd76b215b0225f616572fafa32f8368e7d9d4a7d8abb2bc4a0ad8a998364e51d87553417fa12200
zcd0f720244bffb579802166170cd57d01215976b2f08cf0bf5d211c74403567f9559273691f736
z19bb88ed74e1ae6f2983578b20d3eb7fd59765da77465eb9f5e365e31b215550bb34cefd7b085c
z9d62a59d3876509ae3e216b5c80e03a8f994ca6d18db9f88536b678f466f6daa9c2b25ad1ac836
ze87d3c97b54818ab8e1406d57625933631dd2c3836bf2be9b1fe1f18006636a1e15c7aeca8c4c1
zfac7af39cd45593db7a9794eafda31498bef479144255da7c530c091105d1be06387dc4a2d3d66
zf425f88283bc05875e44537b8da1e4d15bc4b97b46d898628760ffb7e0d3076ee476fc0e95341e
z8827839442a0f9055ce62e2328d6637943d032518bae1bc04e200d7229111e2188cb64131fc6d1
zbf27fff94cbcffa212b27b8445ff6335dba99ae9e69a2fd486227d679924f6b9ed4f47b5959668
zfbc0106ff3c9a1d6a31e573eb5a8f77cd91c005922e7e7b2c46be7e7a1b0ce07b88f28df1261f9
z9c0fe5b9e16aaf2850ab0a96d9ab39436786f4a335e474d94eace01fdc3d6294f33c52796ec35d
z1f665f501a0c8ae9e8ed3af01329106f8e37967fd1a08eae12cc2917f959730852b8b6a01a75ee
z26a3f8db54d3dda29b7e6217c06a562a0ba4a20c9a528df5316c698e36fe8618d6cbefd92b44f4
zc7eb3d191745e207f0be267047fbdb40d9fc2461423143dfbf3a62e823a2badfd35b19d8835baa
z2826826536ed802b34b1c231eb0642c7bf6acf478e02161544efbbce135e5d4204690a216a671f
z9ffca6d8d815fd92647783908d50075958dcf3496ddc6dbf80155d3532cff08b3f0dd19ea99b80
z92acbb453fcef9426a27f261dc6bc5fbad9685088bd784998037ec21a09025da17943ba2f4ddf6
zb2a8e064b671733f2ac689c6520d510784a62d2b96732000873c8f0d532def7081ea4fa02cbfb1
ze54e37a50a315e6311d4b81a3b337f0396f533e14e0c758db5f5632d626083cae82cd446a678dd
z68e9b54e932418c7ba68f27d926987f759af3e213ac18e426bf320f8fe7c7b8aeb64e121823b85
z8d6df3deaae4c15ff20e76c51a46a833391a05bca390b3b74481ac72e6c2340005efcad8ec6759
z5096a8ecf2e21b2b601ff6ea7a690d7ad9bc09fe5f71ed7307968f0977e3f8560168259e6829b1
z3c0c863a03b2f857c47802a81a8eb859c854d3b567a0c82332a4bacd5ecb30facd49f27cf82715
zb9540f4633a4c470fa1fb40a6404f069dfd456938fe3aa31d38ae3df5ba2e516eed6e96a613327
z3d4a83b4ead277d6a2eae8b4b6f4e0296be764f4f0a83f94d0dc63f7b2a36abcee03c346788534
ze96ef270ae3b9d0f4cbc3b76eb7ab494437bf0cb39f0994f454ea7588bca807b8cfda95f0bb85c
zf55c7092c0a3ca9da230fbe5cc618f22651255480460d335b601b568998ccd95d9a43e420060c9
zd5a0db8bbcfd7c79490106689bcbac1b33ebcd3973f5b05cfab83093195b0fb858a64d187b4c7e
zd75e25351fb206952c48a85169d4151f171cd3b1ba17de59db73eb3fc48d260ba5b59ac5447572
zf693ae19d120de23cf8d3ec0531123336a06dcf52b98f67f60a3818bd269dd50ee382403f1178b
z76b85add6acd2d1d06171709ab543051c06aefd8d60e27ca8edb1b7aaf1fbe4967dd6d41b4c960
z3010a4adc9c401f5c58192901252ffc70cc2d8b8d14927cde6637e6af099500a4badc407feb04f
zb357da04c8f1a40862822a4c6db4ba49304700808e87c77fa1c0e4010e8345df3f3fd8aaa02e88
zcbcfef1e09cf469e8be2d9f8ede405ed6d13db8d5fa4207979e17b34b34c59254bdad1cfbc0bf4
za469b68cd35e65488398ffe1f84216de4d62adc1bac680f980ddc13cf08ff937d30a48f6119959
za079a8724847311d4b20c3d848b711b5c1fc305a0e2569648e6aacd3a89bc5cf7bacd7d0daf198
z2e1eab27d47dcfdca63f3e1d189361f647c6b7937de0a5aace1725a817a8f47b56fa4a157fe4e7
ze1dbc122e44e4d989703dba8dcd32c762a745820de2764a7068fba1d1a212102b54793456d7d9c
z353600faf41985c1dd6e0ea1725e0612b9292fd84926cfbb5bc4159a5c6d94ee6352afed1d3eed
zc30b61dc99746c562f4980cd4fafb19baa218fc962731dc83ea6d2f04665331997f8142d988b6d
z5e016dcde4d19e04f7f4cb3b8d84d4c0b6be7a34eeadc246019e42950e431b116677dae99e7f23
zea967079e49e8dc2277ed077cf1f9537dac2809dd68ba6ebd6f2f83b9089e2c6b348372c5ede6d
z74bc1e8ea3aa03c49fa9e40aa9907989b8af390ef7a2c44aab909960468f493f29f5a281924a89
zc53cd1168b7970832d4e3351145040900afe8ccd17741bada908d4dc2962716f85c85af3621474
zaa352c2524fb97ff552ca1db41c090285a0c07b4ea28a5b4e804f1bad52c1f5de18510d8a1da11
za47637933fa87a6170082294447975007fe80426c0d6031a626092048b8c7f7cf8ec753f4f79a1
zb8d72864efd79ff0cecf7befa17a7388b23d7dc40ebe063577ee62d8038e39ee2e8f4957f733fe
za43cef3c98aba7fb3e95333a6d76b7d90806b33a2570c374afa9345e50a7e5d444f9ff76ea5b09
z17e77e10aeeb3b2e5b555e0968511338e01cc3431c6819f9f15898bd6d2a7614e2ab98cdc2e6eb
z54297e6692e5bdcc616326e1f3c3f9c15a61e3db1402d007781ebabd7cb8792f6fa43e063b89af
za668c1649b9848b573a19a41e1e7344c56fff59e22d65af1cd18cee0a34de784c208d490ed292e
z1b8b32a8b3dc1b407452f71817f809e992ba55a1bc7285136b85ca35ce10f79db99d08daa28c22
zf718c9b43aecb8d1e2cee590195e723c33971ebe040a04d6d4783bfe93161f0f6fd610f8956022
z2d997609dfe9d97117e8e2e43c987093c8bc70c31a306d666fafa1dfddaeea7d8927df40342c63
z05a6889b3d531141108324fcacf87f991e1858aab8a55313eab7a9806b9d5653bdf991d70d6759
z7c70900fdca64e1748502d1b426314c9c8ca30915df98966dfba9cb2591464ee01b2978ecf1b64
zb9aa654e7f1b6efe8eae50e0ce49ecacf244b116483dec9a161df9389df5c662efaa9e6a01cf24
z80dd4e8c1471205574248cb01c39a75776cc1c8bec1e705354ed45e4b90fc2123883bb1a4eec90
za6ced62d46c37cfaf90f216b8d2c877d0dc8c0c10c6b2ee2fde6b8f1104b15e6a4723274c155c2
z00a44dae81b13ea7ec8dd51dfd00acc01837ff0b589ebd9978eaf9f5c675c41e5693796d82809a
z8c0b01ae0fbcf7d514b0dd230d7e9f275385b1cff054dd412b4b9cc1c6533e34c1cb77c3ada64c
z4a0d186c79646382947252150af850ed7494f8eee505f8022b64803abbc2e59457fbe7000f34e4
z2aba02380c3cfa726a37a4fc95006e427fc2aa016bf3df292392022f0e5f16842da66c97000116
zcb23a1903a03317e6f30a18b1c9efeec251b5a73fe5c5e645fff092320278ef48fef02936ff885
z4e6a52c8e614b21a5e5c0cff5fa610582833d3396a67712515575334e3ec90a4a495eef7be037f
zee156cba7030413e16e905960591b301478f58ad9813cb06c4362bf286ec5a9d70c51516ff0132
z5501f9d4a63eceac1c8b87be1741b9f081f3212ea81c4c017bad10fdaa523d48877bed1bcd61e6
zfc86c6cd0e7464087fa007ce95a795415f3702cd0327ce016e2468e77a9de4b2c39e909955b6e3
zc80d124b7f63c63180f4cf18da03561c1900978d3f17b91688c9dc85ef3d000b94b2d807b6a57c
z1e23d92b726c6d685ef8bf0e763dc65178a165a00b9ab20a38b15ce7f803c9da624d29e6f3cbb9
z7efda85cdd257bfd446fb0f6a4dc35a662e8af4604457347ab68268fe3730396878938414a4cf3
ze1a2dc150920b5901246a05a2c927a22358a47417e87b1a73489f94834860c6064fd8d3861df94
za1078a878a214fba784e088e81a21c36ce04eb296971ae33c037a7f9cbce2e2f1cbb7066482080
zb67a88e311f2967cc9329eda3bee548ee448948daff9cb43881332cecd271fbc68273840c573b7
z35f23facb9a46cf7be9db29abb233588ddea6e7329db988d6b62b0b73eb57b45f606bd563c9561
zd1e74c3680d667f580860dedb7177451f54264d819ad02924ccbb13714c8eca298ac95e46f078d
zdf661b6c0fcfbe6fa2edcd8f4751887ec6fa3256d3b19112469a3afa603e29dc3f0a7a71f2624e
zf789fc6095ee5dccab915582ad5feaee85806e0008926a7c81d556d2e34fef96c05a027b4bc2a1
z469ad4a09bc61e055ee70345ad6bc1a2a5be14f5e1a736304374a161471f8c57e4e3c32b7098dc
ze940729f94d7c4cca3d22492f0120a3f555725826b6e1262b6f0d218e259f1038da3b26dc29c71
zf516ff0cf6c5412e5bf1a3481757bbbbe53a85db603dbff8cec6414107ad3389fe2b3603b754fc
za49255c733ad45387eb68c91286a93acde8e4c47db888292dffe38ac1290ff2828bb71e37c66be
zcabf5a3aaa69426a6c9a0e8478b7b6901d05e8a956e27bc0b9452589c7ed8a2ad4bdcc5c30cae3
z6d6123198cb57d53cd6a4b971cf43a18762c7166260461fa25be89e706985f476ca8b2ccd43776
z08337f087729ca33232cc604640f74c8b1fd5df0745038cd206b1cdd7e71565dfbcff9d0ee1bc6
zbab280c5ed8e37642f6447e52995cc91ea422ddfa339822758991f7a5a6c3418f5eb415baa954e
zcc24fd50227dcc4e0d369732bdee962b8f3c140931e5ae791cc899a7331a13e0e1caba3a1dc5d1
zaf135d231bc0fae13ead233f77e086fa1b1875d395b1508947e3c92ba28147e406409d31d56f8c
z3c46cdbc6641ff34dff5f38134c903656aed7e60c324dbc7046b8b1749fe52733cfa735eb6ee47
zc8fab536edc0c3278c435d1a87a25b3c4dfec350e2403a831b17f0afadf7481448a97a995da0d8
ze653041a35925aa76ada3a56eb90e3fd373fbedbd5ede75db794f3bf50dbbeb9be13c783bac8d8
z4db459241af5380c0f2f81656eadffdaa4a6393fd3952b6507b9a12003a9899d423de7ff8dc6b1
z533696c8bbac4b25f8915f6a3b8f8511e5fa495bd3beb4aa56b6de6815f91e3d446818fd7bab94
z412aff342e2f953f3ebbafd60f27742326aff70778754ed6157a5a46b2c68fe489f9ae834e6c82
zea273840d70daf4557c8060bad494b72c8240ea95b62f7d3e15028c2b209cc4bf8ee8edb6ca89d
z7ebad82d765a6389350ed413de874018f5ecddadd2c087d106f3a30797dfa1a57fb739db5e7bb2
z6b57be0a7d2da67be65fc7b56be741e213d09623ab7e6ddfcbab7ed15e1ff5eb9a5e1d491d01ab
z17de6a674c6be44c4ff7eb5a3d70c75732ccb1127dbd3333fafdf5b9b373f1467c059b0b9dc332
zfc5a4996287d770234ba6d6a97b11adbcb6e7be107fd0a155f3c9acd4df2c289b451f5a21a1f42
z6866a2e30556aa29ae3db0ef1d43d714cee94c2cb4f76f6b7407abeaabe2c4f893c73ff870baed
z045cfdd56ccc406259765f518cf786856b836e12598c8f6453c4fcaddb34f38cd4bfd511ea642c
z4f61721c96e93d3ab8effba97f2ae675233436f4bd34dbdff0e7c3f72e0a33c5ab2e0ccb03db1c
z6d49a39ca032d4503936c4f41cd628a2478c1c5d3e6cd30bdac277fa746a94a89a6fb204ad80db
zfa53464988b5dd8d38bd5ef196770ade7cea904474cdbb1659975eb6068727dc7a0c3f5691d357
z6610cb0221927f0f8f929aa916d22f0a736b93b1ae9e137036a51d9648370d97fd9cbe0da420cf
zdcd95d27778a5f12a33361a84641c6f645aa737271d5604822dd1912b119364dec97ba6cd0e36e
z2aa2975bc57292f2add0fbe9a4455e8ebad6e98f40c2031b5ad632e74a8164db39a6ec12cdea8c
z6dd833effcdb73cee28af9cbc0fa029d179b1c558bfeab2155ed6199029ecc9ffcf61eccbd06a3
z2de343dcac6735bbeef7622c83829d45aa84a573ceed166813b3589f6703ddebc3e8d400cdb70a
z597d9102962feab102895820d11839586636c737b4542ea13e5973b4874e6ba032e4d17d29ce1c
zc411b4263527988197823a3acdca30b441a2f079bc0d81342d7f5429983f3bdd087a4b4dcc8f04
z138b2ee7e744b5b2bcba3ecb6dc9ff568017755191a8ca820bf9d3c0e109fbb5f08c47b7bf1347
zb15e19c64dde9b899ea1ce98fa25232e52e362414ba71a6412f7840abdb4b6a9e7aa4cddb387c9
z6efed1b1ba7087fe9fde054edb0affc79189fbd617c23b51b5e4a2f149446a115d01ccdbafb376
z8c8c4d642c7c33370f6ed8e64123e3eabc29bcaffe4b5e25096dd59324fa8c9f7c074f5c2c7c89
zfcff134dd464c2f49c4af4b8e1cd93ef6cc812496d5c2570b856939ba47e4ff82c77abe20d3285
z58b84d776dc5099e66d27091d8bd35972a3622a6b4cacf44530c8ffeb25b4d17254971128d5506
z86345e5480535296c6a0a233f8560b6cd509cb694001d08ab6de64d167ec81943001aec0f6fcba
ze91f2388bb4903f904e33ff8745c1042e6fcb34f802221209733700b1d3ad778ade47812b1b10c
z34d6f8a69c54966b5eb3eeb624fd24af9d259166395a687bf2462524a07b47c2ff5f9838f5ae0d
zb835fe5d7f0a73a367b516c7d8d7999c37b96b2bb1313ede3b457ebe6f6012094f8f806ec9377a
z8c3dfbd5f469acd79a82c4b8c3f715c1569d1412b481e86e4b1dace5bd0f5f2716db0cbfe1c467
zda57a7fd2e924b8f3d66989167782a633ea229c2d49d15a3fe86ea474415d4c7b8b1d6b5efbb4b
z471e1fb5aee7e1cd1931ecf92697c66e1e76e169f8e53e9b0c204a650a6f88ee84ac0d749c3e98
z901169a437d3552ba3c0004ee168ade706f2fd3ea8b4ec199d0692547f41c177b910b405e36651
z600f84b650b91491f6c3ec75b9f7600a2813003ed903559bd374a8804ded5041d7020791ae7925
zc1006d6e5183ccbbe4c53a3516cf286c62111a70aa765b16c0e189745d00352a42d89a55ffd4b9
zbf34a91addbd7b5358d1aa2bc807bb7ab5bb04d2a9c50ed3f2ac37e7acb7dee5edcbf4cf1ad005
z8d28257d4fac477bb47e03520733a5b68b1d10a675b7844573dbd42c16e05ed3789b91cb54ef78
z0ddc50195b505e86aeecff7d58e57472039b59f9b2bf7c1f38c1d4609b7b65b06648a0e4072556
zba2edf1231eefbf65f7dfa53f197f18fee6cd523b06dd12507cf86aeea77c38a7e4748c84b237f
z616230004de00346730230466c778eea57ec2ff57a757e8e4a12f0661990b97e5cbf73a6f3ddc6
z52d2eadfc7691046e77a601be6c610b513b133b6d1142bc5a6a07977b5727009e7bc17aaf3afb9
zc1f8a5bd59e9eaa54949cc6f8fe1a6e3ecbfe09ec3e5c6f4deb03504fcb53879a152f34b1db6f9
z0ac1c5f06edb3e10f55ccb506aa62a5ba377a8660e33fa14249b26686c5b4ece693460472710e9
zbc2d02f709cb33b70d3007d7a4a819d3ffb4311f25e3184a9f94e2050b0d35dadd61846aaa6357
za5ab900d49d2efe94a28729b60575655860d56c302a52321c6c5706514df7587dd85987d6a68cf
zc2734aa01f32727d8487f98ffef3b6adb94ceda6e92efb2ce781c58744a02a8ba92f50419f6311
z0d312827b6f8e495ad0624307bc41a122b7b58224cb51904d6d0b59f814270880c8970cc070020
zd3bdd628bc98efabfc7c54809f7953202d061cd579157bbfac45fe4ac7ec178f30b59d1410d074
z7b39a3828df81ac799ddb98f9e4fa4d3084ed9cc02d94a50b38c592c22a41f05044818072ca4c4
z989595f17f0b04a5d4b30674ec0726f341af19fcbc33d07c9133ac301ecba100e385b369e71711
z79768017e365b453a95de78d2124777e968f7af012c23627472df2cdd6231792ae8c4ce486e60a
zf2713084adc4aaf51e12f6090088916cc59cff6b46a34b0d599ee3cc44774773b441f0e3523dd9
zfb4d641723643a4efa7de269abe10ce63825b40c6aaaa7107ec98140218b64f80a362d5274214f
z9cf7424c01030f0b181d2b18731c7fe6c3bb46a4255827198ab57932f45df0c2184472200f3743
z687e9d54fb0cb865be921b64853e9f214f309e13ad7f83dc6854a94f8ab64c4c14dc26608d63db
zbbe5ba4a63695484ccb313c37a2f2eda5e3cc82dd959dfcdef033d90d00651a4cf829bdb7fdbeb
z39240dad63804f91f2666ce8fe60b823d680b6cb94498cd7a15f23e0eae5a04da13745b880c058
zad9227b040c8cf8a7656b50e788bd33007ac0143042ec3c0022cde89dbcde31c25bac4e98d65b1
ze43bf472b0706b59c19c7800e8a84b3b1d7ef8abca52081d308fe16f125e3514121b8263b626c8
zebbe0230057f745320bd8674d460d32c649ec98f200fe3631639abc265e05f0149e17a6160e95c
z572612006d1a9b553b14cb0dfa52d51ded5609cc4665e6721c81595a0d9a333c74c8fba5a55403
z760a702229f8911960f160cbdf216d0de146ab164d2d54212ef0a2a01d4311747ccdc14313f39c
z2799252e33cc1a66dd905448b3fb57c87d8653fc59243ec4109a981d47fb09bdab5f5295f15608
z5d07b87a9dd9c4f25d3f430ff92d371898bce53c30295d0209eeb4b5f6af37336b3f3fcdb7c81b
za63fac16faed4562785f2a24ca6158d92c97dbba63f1c955cbf5db1025b887b1cea75110e069d1
zbdc5621dbfc5df3a99ea9008381a1255a7d3560d9db9a4c228f1668994c3856287ff1e1d913435
zb882664d7a9171d8af469ff5898f96be3fb1561291d5f31946ff343aaa676c9ad58bda749f1a20
z80fcd30f1c6b505014517fcf3d8ccc888a5d691b99e899eaf9be9939609d8935c7dff1d247962c
zca923fd90c0d5aede71be963af0cfb518c6c8813c7860e5eca1d99b5acd621f5c66d7dfcbb9e1e
zdc71159da305cfc48a3c7babd36afa988f3ffa5cc60cb7ae613750380ecdd276e7bf35f627b91a
za5b790472bea68b8660cf9b6e4a3f9288271ec3fce2cf06382901ac9ef3be8677ea3e9d12a8ea2
z8bca8216e50fa110df56f38d9177edee972cb746460c5bae9cae2d72756794187d28b38e35b946
z63d9d60a63b3736842bc93ecc65b09eb16326e8a51365b84579b0f166dcff64e49da6595f4e573
zd3a31fcf2beb1b42989d32356032bcf9b73e1df6cedde72bcf7a605138860b78e01a82eb55ed1c
z06bddb0966f44e6ba7cd1b3ff8da02d9599d45aa07594c2e39d2a849fd67423c982e6dfe81b288
z861dd2a827e3384bbede84e21431a2efa5e998f92966d64fc1f96ad738a6fee6e04765c59c2702
z8276b5fe3089d448a82c5ce5628547b2e24fae8ac66e9059b59855bdf72e0b97f92eb1e19b8386
zc5e7d9b3cda4228be8f58e8005fd0c9168d249c70be3dbda2e7db439fe4c7b1d832d6960768421
zc674b158c7aab637a5d34c8a814be5302a0323586b7865e53fa31d066ae0b027912313040ea6f3
z120c5323c217553c9665b264ba184b18c2df2617e5c1366c2520340b819093f253c8277ce8f7f4
zf82dc6492716d4ed0847e9a652f3a7b5eef7578154fe70f48363003a7a581db0db2b45efcb2bff
zd863952544c122326b2d47a37ca4e9c45ddc91733fe597c5143b6280c9a2df2a1b73f66c336f1e
zdc6fe4e8afed99163677dfc7a184f203731f159bcec393d8c4603f663d2f30c387bb2995f464b5
zcd66935dd2c09aa420b5b3ee3cef860aae98bb3c44ee8e3d03ae38aa68b726d8aabdba6901c067
z517531d6b7c1e33f4fdca96a6b1e775399ba389f3ccf23ea9e9db73399c0e726d1a3179831eecb
z8f86c09cdcc1bcd8198d957ce04d6b4f624fe4befc269376b3cf4b76778eabc0215688ed627191
zaed0470a3a77b9074e3e5ab0d74d71b55f8f36ac90abbd1b0b95a623475c8ee71ca726c2d639ea
zf796f5dc8b213ea477718760e4b840a37b699c7787a42b10ed1af6326cccea242612420a420fa5
ze2e8e438ac6cf04020693e170a92d9e47ef5b3a7805bdb3cc7578d6831320e5e45c79e236e62ea
z8579f73b4a12553b4d1877073014adbead1e8290aa78e5e05a740cdfd5514a40213b20af493558
z07fac757bc2751796641ebdeec3647b4d9fca6285bf114df823aedf7326bc332fe74cab463e3fb
z685392a48d621b5a822764fece0e85564170506696f43c35fb22c698a94fa558aa392610540a9f
z185452713b06da034efe404746f3662edcd05250175e03c7b65b2611c7d3827a7eaa2f15b8f888
z82996bcea49794255b838d5eb174da454fd1a4024ec4ca57f34f57152c8578299950384b464076
zd25431bbb62295eab2532812fc2509e87c9605bf5cfccc58747a7af840dc4fcbdb12c1d019ab6a
z161b161d84062429a6a74ff703947c984948ab4faeaaafeb4cdc392f71b58d2d060e3e0a9b084b
zd07ab8ff84318a8fc261eebd73729006d0a14e2af99ea3ec9347b70f70476f163a9f41cce98ca0
z67d65ca604c444b79ebc77cda07a2b5bf5a02549994d4388e305b2123d449650fe88cc323d3be5
z37e57edd62366a79443cd1f56a67d1de98745546dbdd4608b71b913032b590bcaf9bb68ae62f80
z63a9a311e66b76f518297c79d048fe29be480d9f9833d609a16aac8537c09872564d1dc49c4ece
z3b1ac31aa04b937d3b34b62e472cc5f314e280b045f0dbe0d058ddadec78891f2252572ef47196
z88e5f0afff4765971013f00a8c312dd13bc1ca46fc84031d66c184e0f5c6bed2c7ec22cfc1e615
z90f9f37104ef71a0dc772885bb1e1d47429dab7d9d736c3fe262e42a517eb3f0937e865f5b6105
z16cd9d0574a1d953dfa9490b0d9ca721388a3ebc3f427ecf85572e06d99add542d1639363a12c2
za08c960999f3da2558349213ad63d7723fda17f42fa2ce05e4f9a956e90a4e964cb2c4c59272c4
za0cbdeb418bf62d13adf9e60d702facf9b350a1d648f6446b238d449aafa59ce9f9d9f302c7f68
z6143fe63e9cacc2d1d83044694e2eb65442eceac1d4ad038eab87ec00c05a03879a2f21bcac641
z00af581ac7d4bfc497b403b51933f9eae38e577f753ce01b0227e01e2ba44391e6bc853067bf24
z8ac923e02e0ff971e61f5b73ac43681e34f46126b1f53c2ce96e857c372f8712ca9fa7b6da58f5
z3eac23beb2bfecd38b259053b797645a52a7348f82daa400f5e8e4b309911e19343b67aee914bb
z466cda689b539b2b40a2c5e8022835ec5387a1fa9be63189e64e3b65e6467e04e036da60f46b95
z17d667ebd3564a030aa12d6ca3c276684de1495bb2b7bba50a2f733c7a02d766196801c0cac4bd
zb6288742ab65d2559b208d50856244e2a2100b9696fcf324f04106b04829699ce47be196f435eb
z2667eb12f4192f37add8f028d0707e8bb50722113828dca075d1b919b7648a2273d23410c9d8be
z7d6b236609c69c3283d907580aa7413ba1954fc19a49e37b07230b398b0b60787ec7c8d7482110
zaa1a4eceb54903a5c0b95002c22ab72e8ec4954f863afc0b53518514016a29577f9bdbb280c1e1
zf50ea116124cf125eb0d84e24f9f1c2a264358cf66625b43268f726598b26b8886ba89361fd0de
zb95e7c3f73422862e04e01ed390b34fc8d87a26b38fe80ab9cc4e6f0c383240d68ea406b056310
z8be090e01e63ca48fde7c1b97b9def527bc6aca9cf0691cbc850d580e9eb7d2c0a9a20a8fd4b97
zd35bbb5e75cb49d96f0f91a2f1960ba8c4bd0217be70ef183d6b9d1ce0b6b5b97f5986a56e1ee4
z7783eaee82b7df7b972b3552c612c051e23a075d701b371903205e4a0ea148409146e73328355c
zc8518f6ac6b397ab2240a448f6e7417ca873c2b22323cb11b8c29599b7da328f43447dd39e85bb
z45584eb9bbbe4de2ffc82842ee085e8433eef7bab8de4581c12f54960302be8412844fdefb9e4f
z6621e237a56a24fc16d3d2d4cfbe2a277abbcd66dbea3197b59f4278f32bcb4f6c218e0370e71d
ze2fb173f80e78887996d1bce888d07e7be91fc4bd9527d16f3f9ad17c02b63fc22291661f0b3fb
z79775a8380cefced95a225151093dd126759096346a6e8148a71734b809860f888e82f0549e2d8
zcc61bf6c3a969d74333183659c3646666d183359eb50b10225f5dde83f4ae8fe77d49695f75643
zad10619bc74285cfb6c0699f986ec1f01f527be232124e697c076c9e127b45cbb5899e87f55342
zc9f07d6f47f0b4c8ecb855e038e7b997a2c0f9fa5530f37a9776270f8b97fbc48bec24e8ed904a
ze4bf2ceb0cdca11b0c99d352911b2599785b4a09f670255aed25bf98bb759fc50d565da14649a3
z80da8963c9a61687df3c4e00fb461bc3d59b73ea395a79e524c633cab40a63643e3f9a9a9668a6
z24e1497372cbb1b4294934cb8319f2de356518af0879aa2403e5467d18942134ee52d17e6d0625
zd667e4465d2d7cd5b97e2e9803dc5029038832dac2fe05168f0f62e8b433368ec5ad6cbab5403b
z6ad10c9cced3596f30e9f7bc79f9ec3a4d9d5771bcaadb0adc4615fa6552e66f4f79ba8b86c359
zca86d4958b027e45d0369d41c50a115194f237ccd95f7ab8650f86b16f0b0d7ca9fb529e730d38
z0ef2d4946a62e457e25aad18c9f55a2fb7d2de762ebbb6476ba8f6b5453f254a3412be35a31804
zb25c2f320753561b513f9c02c47ca6abec540de89a958a9327db885c941a0339cba5498d93624c
z25efe60a605350e6fa4d07125067c4c7e5f55c1b5cf4412369e099b2c32fba07530d050b68a542
ze3bf32652ea9cd31872a3b6d74a3e851d854a73912fa0370b35dce4bc1b80d2a031542adb17c90
zb875d2c670fb884136c69fc6cba540f1b8bec3687d49d6ea6bc02f33189e19632f60191963d86c
z14ff54826255e0ea4d0ab892c711dc428f088c15e2ef59f8718f227bdb56ad1dde4c5700c1ab11
z2d749f438c44b74de72271541fb9b2a16c3b092e1eeb8a8ff928425bc7e67e253a5dafb3648c66
zaf165e7d537202514520b0ad145a5d83903174e2df58ef63357de5fe5018f6e168467e7c5c9bce
zebfa250f6560d49a0da31e549ac81b8b7f51e98159f0f95b1f8524e5fe0adfa1c946fa054112b9
z9b6bf5d65536f53a57f7e8bf7464696aadcafd5008802186778f2bdc9c934e738cf8c667d3ab0c
z8c97c5baccb2576b660b5ed0d44597cc3f3137cd97e4e9d19a657491db821017c98e28749f5d3d
zba5cb3e5149ef870e50a9c7e5f9000ff3e0f12b1473c2c74051728722334d92f1600a913e69c11
z07d422f1b79d8742483e934717162c5eaaf9a1e30e9c50494ff4203fc61f8e9a3b5b1ef286bb11
zdc4c990b71821308b41549de732647325117fc2c02448acac0a8cb7a3f70e942ce17f23ab79e5d
zb25f3114a15b0db7b3c1cb1a7647af091907ebcecd3649353f843b206e6f9df02b4548f48c2a78
zd402cda29a2d05376e21a132dc271f396e8d10366fdab144122c08421b32234e8b91fcb3b1c3d4
zfa5e1b5c9f6eda66672218daca409cf48e2d17a917bc19c1116f1beb4141d475733d1f014cc56f
z29de8374bb26b53fd769dc41616c7df2b824d856ca7193a58fe88428a287039780b37bf7ae3244
z2ef18a1e5a20be3be7b66657d77befb7c8023162bb2464f3920d1f597dde2d40bbb38d1003ccf2
za0c449ead96f9cb7ab9b9987588c885aabe6038aaf2b607aa056ef95263fde8916cceb49086640
zb2725e2e244ed47db9fef4587e1344fab87438398e9718057345d4efee57bea0cd2d17dc4c84c5
z83edb9c10b2cfc79f0cae91dc17398137b557b3e0dc5f0619581cef97bf3b65fba7060d2926d71
z150cbfaac5003257594a65116d7a3a3185f3b5a303c1621470953aa1b8e7ecc63feead496f32b4
z6dbd1419c1bdbc10e388cde14d20c0428ee0693176f7dc2a0707ad9bbd517612246ac978deff1a
z6637d4998082e6a5891f2c098704dca62ff391bd5a0681846331d62860633765305c086bc84b9c
zf6254745dd1354da058525b34481fbd3695138dbd327ee768dd7d8240d462a31ff127664af5a49
z29f68824a6cda78c34b1c4fb5d8dfd1847f5134938f91f7645a8d273dd80c485bb6bc8a6f6eccf
zae70fcb4bce57e3c8f8f830c549398aa45b31ac75c5b6dd2ec6374e7ab8fe29fc00c8cc6f3f3f0
ze1bd01c0140670184c6ff700b9fd66ddb9f4e0c73350e39f46a41e336e1e751cc29a4b334a4ea2
zbaa0e0bd9ebcb21300f56a319a2b7ac1efed40471b171f9c716e5446da48c6749f78cb4587993e
z17d956c827e41f705caf381e8ac4f98e3891c58788bb695375828e379f841a7d10dee21276688c
z6e59d6bd728e8bb8457b4c5ae83256cfc507ae352c0f07973291fb849880c05f5f2d1914dd9268
zf021370e358e2e810cd7aa10ac58f8df83336cc6b3bf9d99d620befeef3cc091af03a0df397289
zeef50c230d8d79e493bfe25d8db9d556ac4fbfc5254c2fa24c6634d653f9a24ba260a8237a762a
ze31a0437e8a75ff02db611faa1558e3e8372b1712159f13200a8a16032e1a045b99d14663310cc
ze3f5fd73de6c38e2d96ae246ab91da1cf3c061f019e98720d83af370de79807a22355c2d9931dc
zb405c28082d4fe5a164b51326e6eb45d59b2e1f77016267367760f67951aad47cc9739b4d69806
z07725f649a360e6dc0d3ce664dd68bbcc1fa2ce4b656fc0e109b1296edbe08ccba6c39f31163bc
z6251c633ce62b8cbb6f28c820c366889ce32065f73fee24df6771ed547ac2a73e8a11970441c73
zf67816ec2920e40ac241a23ffaff0f726a2153f24155f76737e25e8a5504f68edbb79d66a5f4cd
z6f90398bce550661e58a2aeddf73867b6969567ffc10de5d645f9cd01a916612ba8452584148c6
z0170dbeb0eb009ea89cadb8d32541653baf04cd3db8b1604642f26a97abb7d466087db5bc64f75
z2ef66af986c5df116b5c4e07bfa0ec33db64192cde002a7214d6f24a8975b1ec0e40c75041a285
zebbc77bf8257331a1735b76e98082d7c961e38df99e2a559e8b6fd800a8558de4da5e27dcf6dda
zb108f9281129a41ad8986439b23a9f04ab3519190c03d201adcb30e9ae3ea2d7e60dbb293b772f
z4fcbe9370a8e76f04f1590b47eb7502b4a535347820b74329b5ba4942e176694c088201e4f15bf
z82b6fc75b7566f1639f0f48d5a55a29d6170b1f618978f9d02f2f52bb1e89554275542fe813e0e
z8b605e8802504592ef76000a95d8e54ced11e4facc4dfbf5033b718457e857845567c1711bde02
zeb2c8da62c4c59f88dc13b8693cb96ac09e1b365adb7062be454a01314416a7ea165c7bfaf6fc2
z9804022f80c4643ee7ad668bafdd7d304fd3d5149119a29d4bd175eec43245ee10f1ea8ce6c6b9
zd3dfe6b3727c42ebe40d3e47efbd0a04ff9e6d0651d1b83f0877ee56b7fb84e77526933e3ebe91
z78ee9e0393103a1131ee29cc7d0c1ba281187dfd0335918e8adce92d7d259a31e39754980742f1
z6c9dae9671153a652124dfc6ce0dc417213b1ea5bf9a5d7f29c3b1b30bb9ffa0df1ed95011d703
z55320a0156350340230041f393b4f7df19fd4f4d74a6dcae26eedfb116b38cb427110ae18db8f9
zdaa826f2965cb6fb5c256bbde22b847b132df8da852b95c943c430d6fd783cb5737b5b528fdd9f
z8f10e4ab070c36bfda4af8552d3ea7311a77530e1cbd38e345b8e2a6d4a7eebed70ef54021c4a3
z3bae2d39c2727a69ff4098f3e094ce93fe5a3ffb905ea8e16039d42d10315095474bafe65ba915
z2f48e8dd1a85290944eeb59fad3505bb5f19b6152991f6a5cc44b944f4523523aefc6406a2380e
zba00e98aee6ad6118caf0ac14805f842c05ff2a3d42e7e224b6c314b9afe2b682b1a8c5a547a77
z735653d38eb063a9eced40e2bfc128b5191d60cf343eaa21194068037a66e4089d265ecc71eb20
z03bdca0dec93e6097b88506216385bbf565f34063f6ea715e83e396a8881f5051450be8207abff
z98c13f31462303d27304170f6439a048f0642d50cc628578cedfec81ff0701cfff3411af3fc09f
ze252d2c8a87e7fa62b44c60f55bdf0aa3466d5b384ada65364d650920115487720a4b137270459
zd4a5fdeb7d021ee0cf71673dab3023c7d480a3f57258c86f5a8fc400a8435a454e32439b074199
z872744a203730c79ae88f6a6667032691cb8b68b6643d25c8f8dcb86143e81e35f8eded6e2e4ee
z1d675ab08944e1a8750f6e129bfaca0757b671fea5ef8df80727faf78c7d4dab864e6eba13e3b3
z4ee6f9d691579e0cf6fd09108cca34d3402c40b59793bc276febc54db8ea4ace0219242994862f
zf780d7b968807ec5e1f1832ac2cc417b12017968bed5dd6c3fc3208d95790e33508d82af5d8561
z1c1473bb6b8ffbc6d3f56761c2afa4c331059af74cef382c640ab94e9cf3df6bffa593e2e85e85
zabf25860e4f13fe6cfd32c8b9c203e584d3d8a500f779f692e18d17ef3c254b93e24863b2ce195
z25e5f7c50c79b3edf9071c2f7fb75ae63fddf29f1d1077500fc2444a132860fbd0eea9c29a469a
z88fd06c5da0027b55d252692481f0e643d16bef0ab929571ecc0d077a92f6d6905551a28d31027
zf9573e7142ea9a201bbad853b6e2959ddba0ba8377dd0add39d6cda5a6acb7dcf54d31372ecd99
zcc7883562fde2c3f9bbe945b7c91058d55e557a20bf68642d4f11412675b579ce7de6b4b98c302
zc60c4b8b79cbae3dbb3abbc8465cffd71afe80b2550a56bc6aa2f8dbedaf8801b9e42a9a190c82
z67506ba77180d10ba92c675389f8aafbb04e41e1bae9ea7b90b9750f6a286a6d4a267ef1b5f576
zc03d620b73d68a76351dee997d0c396232712b72bc0090b91dc3b7603413ba75595f3942845a86
z6efa9a7855cfd855c319901c684d82cf9275536620c9f0473a0f40d851bbf9cbebef429b8bdb1e
z1f3140beb072ec093c0920ecb3bed82effb9c3576aa8258e016149990ac9ead08337e3fe564f40
z6cfb2fb0760e945fe5cd3ad0c958c675730931ffd0b125c9a5716d013203c9bb0db2bc3039248f
zdae369a89c031ac8db4e6d09204e993712f72f3e66db628625b2246bfdd68af80ab1173c710b4e
z989c887ee065cb36f0d3489e5f432a20455903a19f5a1c1ff4be99f7c6ccda4905c3ebbda2d523
ze2b146371f199876cf20344135a451a0ec15e5dd6b2ce010e3da3cd90c8086820d55fa6d892fb1
z5a822d68a69f00038d4da28bb450645d9aa0941034eb72fb44240c350eabff619893371c63d227
zcf379e8affa3175777d2cf59df663666bc01d6791d985b0a1e0a282da644f2aa2e52e000a3e32d
z956e8b7716090dac0f9d8cdbb7cb319683335dd161044a7be2e16e0be7542a3d985a580fcef440
z515f5393a0ddbbd2d45814098f0719f8691b961cc76971f3254da2b904a4dbcdc888e29193fde7
z646b5b8597a5effeb9024aa4dc4a21aa199ffc1dd36cbda12d5b0cea99c7be862025db769b5d7e
z4e286dfd2ebd4ce06ba2595e543b2383c3e4e3596d734030dba9a115f0d111e8e1094a54e58a6b
z84d65336d06d3706bc993aa067baa2f5d5490d3b00c4e3aece5eaa9fe9e9fe12c3f51477599f65
z483939445bd07d5ca711b741f270a52d583120e70c68848c8ce9f791aa482d841a45401886df20
z3e21b38df266c54969ba218265ddf6b95c9014aee11c9457d188a3f141e538b8a746b22d892335
zb80b6cb5f65c2b38556f6dab17d29ed29b49b5143b30fe39745156b165eea3d45aa5a36f670705
za22b80cb22a9347bb12c5bbdde7397c8fa17fb6e8910204478651778395f5170638ff5e3fab056
z5997f458cdfb0c9f0b279d3ba33a55a606fdfc4fa4ed374b6a247d2b0d7d23518f5e7db6547f53
z8b128e68da251d5bd4aa17f8e5710de0ea0ceaab8bc97279d0c4532ddc428c273a36c30c4d5ff8
zaa1a181ed578a9bab3eff204968efb0e37740e113b80eef8f0f9aa8640c6960aaa472838756843
z5a83c4d1adb2a0382c5ea78aac29bfb61c778c916561afa911fe78d49468f1efa5079ca565c9be
z85cfcd7aacdad965f2e97235e7b8875a9b1612955b185ca93c89738850224564888a8d8b61eeaa
z5da6622e7a32a02efb27805adf073afc45d4c0eb8817ccb7fdcb0d2e6e4cd24d5bb3329c465a44
z3c51a9f7b249fdd053a15b03f4f9363c280bee8aa19d6b2a43b909c7428bf952389ac47012ef4f
z084335711370963a8de45576f1bfb4d2535b27c21b15c697fe2ed92b8eebdb41c37145883ddd3c
z9cb7a8d5dc06d7ca989ef9685a70949efbc9dbbaa999f9df32ed573ba18d2812a16ea1796ad318
zee4116e303c0ba6198a8e5d89b855a2915021e8e93e6636a61b2c26d5885f83105e414e40d1372
z854a13ec226374c792d173ab848327a5f77e96e7001800488720718ae041f79afc4422db379c42
za32a0b0614e92a7d0ddf535ee5bbf3a34ef41afbe8c32a96d20a6ceecaca169b19684d166f7098
zd7e188ebfeeae86d5da379a63cc3549c73284c7a7ab88e87d48402eb3ec62b2fd2217041e89fd8
zf312ba482f9bd2dfa7bc71cc88e59b262d19be6dc1a78af8b965126d7c2ba58b86460c4938d20f
z290a91d193dc3bf7a28ff50d0abcc0d14e62fc8be12f3245aded4b9963154e467a3d3e528f77a5
zf88df2695344cfb31effe8fa9c1878f2fce8004808c008abdd356052a4b5e3e161d78d38ca1467
z599f60db8778a33178c2dc22622829556b3de8d4e258a96406fc06472bb99711a4a05cfae91285
zb89b87639f84e7c96d9a694e7159678ee51e55bbfd9ba147b7e8f2b5af1fd1e84d23dbf9c7e56b
z730581704c4ee57f5d029a85b501b80da78b045c8be531820dea12acdeeb724b3738af7f8365d6
zb70854f80baeb365b6e560c4ced421ea933da2d47ded5a228dfda2e73a161c83efcfd4fdcc3f07
z44557a24e5d6a19a64db1d97b23fbae7d18e9efced2c504a33341c790048944b25565631c501fc
zad6343ffb4588d66e2ac834440c771d40b3831e636f0d329ebeb00055baa9869538a11b7c60174
z2b619bb32003c41fbfa6f586f8a6ee328baa558159c98989c31a726c318f773131cb60c2b64cea
z6e3eb2186b5908c1f0cef4462ef471970b8f0bf1ff5f9d28c98ba0429e0a3e61181c54931e9643
z0296c305db03a22b5e9a98fdf850e6d9346ee4649b964945496f8818ce213ae81a43f6bf977646
ze01465249d4934c42051116a056d8813e00f7149ea4ec0f338142080e868f777bdcfa0b80dfe67
ze1e559e0a808203821355aaa3c45069cacb73b45a61a3c2a70e9044461ba0c63882fd9f85946b0
z2af3f0297848aad643bbf7b38e6e9afe7b66de5c83f1cce4c17ee3ee6b1cbd3644d877c078f803
zd21213f1c6d09d51ac593d50d107b45011df0dd745d8dcf3e1fce84884e6730bf84b2b0934ec79
z0097cfd26108cbf085aa50660a215725a6439103464c294b35debd6b260534976637e17c58afb8
z222532c2e4967d1591bda04b2a775253b75c917e95324d902ca94b1a80fdbb5afa7fa87b1477d3
z38ef37fd441b5e3bb8ae1716954ac73994d926fb74d1c75ade233a2c905c92f244c2e3ca150ff6
z5f669bb36f4048eafb44ccb1e448aaf0c0a5f562b7b9c940aaa1a5dac797d8668f73ddf3c9d604
z74064099852ac89f7c53abb20065da00a3a35ee0cc20db2dae510551f1010d84e9d098c229594f
zd6e60a5b784f29a01ff35ef75e43b1ab2e8c9eb865988f9feb9464a44ba81332444bf7c4eae12a
z1616b4b15cf0615cdc4aad999b50c820972ad32385dc41505371b402e797e8cb0da194bf03c9c0
z02e587fa272f5b648de52edd946858c2d45d5a9ccfca15c5dfa517630dcde022571f75af1cfe83
zaf96279fd6b557af46006b7d751e9780a96a3c3d0f7634dbaf1045f842748def39378299296829
z3d49c224e21953c03fdf96941328949a209af5de9fcb15bd5f332525e8de7006572ed52b8e3ccd
zf94305927150e7ce39902eb26548dba63bfbdd982f788c9d5bae863eb240beb7f12107d30b38ef
z8c1dd05ac9451240267db3e85f3b59ca5df647a9156acd257eec82767b8d794da9ca817517f6cc
z182157c32c037de3b209e9dd1f0e39f394b0d0c73bd389a24235b3f1dfe6f8c05d1a7a53e1b8bf
za295f76b0750c9dd7a8def217d9fb2b7459970b45202345152e9d716052dc85286921833cb5641
z784f87cfab66274d0976da3e3b7ccf3946bc489c4d4d4654ecd1bbebe2c36f207ec456e637a633
zf3ae737eb0011b935209a47ec857b291e4f5ef3e26183f488b44b38ac0ebeafba22ff715ab1e01
zd8426aaa31080db0d413400cf646520eb0778d92f670de355b756fb28dd2b19e99d783084bc2d3
z06cd2a8c944fc37d582cd6e484640dec79337d3148f658640bec2428f8e3c18beefddbbaf87d5f
z328c749bc580331cb8a3a6e0311bb5fa6f470523e61aa38ca52e964d5ab9cc0e636bbaa242cb5a
zff76b24a254201771e77e575d1bc0a797f5c6a10e03994c79e9b61296b03c377233ee1b6fa50ee
z4fbcc85c68d99c043c80497473b36f8ce3006f90bee7231d0132896ed7817843ceac590d426e57
zb2cb6f487fb8d50cc782bd5d04ffef53d793d65970da115d0b6022207badf5c521e35eaa79ac51
ze1f87efee4eb9275ce38ea38fbf1b17c15726b869a7347bb22b2a8bd2f33667a383717e0829e37
z4004fe1db702be6061575cb85c41f99efa35c2be2446f70c06e94c72baf45b8ac4a6fc9ed3ef09
z6dbddbfa536c8995709d76bc0ec6eef7c89a7c24d920e37c186d542a3d7aff27fce571e66ade11
zc42e102ab0c726cee215684fe0e6d3d5852d0e497c011b521803e70caaaf5268544f1d0e6a278f
z759ad275ae094cc1dbbac1f16ae5a6e61ed4f167ee9f7e94c23e197bf128f84aea8acef240d223
zd6197148f7478ee1f25c8f9f03b2213e01d6c5f4b06ce2c2dd84313db8c44f0860dc3d54e3b2e1
ze99266f05ca3ce91ceaab074a7cec4cded460c9bfa96e87468c24a10289b6ee86fd3f4afbdbbf7
z2ce618b73ab2e72e05f39dc43ed2b95e916a41d201e6b850398c1afa9db7782adb120067b1cb46
zb48541464941e9a6273484f15977794d0e7a10e53e1cd930761249fbab88fab87557bea70a3baa
zd24355a066e502e2bffcfada11e2b0018ac14e71dffba92e498366bce1b291320beb55f2242fdb
z870391b429b40000167403ee86971a616361fd4dcb9c099d0884170d9b733997f0d2252102e2f8
zbef801dc254c8a21003193bab6f59ae35827da9915525150e194a7ccfffbdef9e91d583686329e
z6d8ef325b1c7e7de0aef5ef09ef9c91a1793d427e62d4474a391bfe99cd0c0e6f7a3bc82926cb8
zc0250323870a764123ecd82ee9322e6f31a219954f1d7b276294669625ce11da2e512e13a539e3
zf492391452ec13c7a3e620101d2c9db8f5aba3a3668f56dbf95344ab9e21dcc60e269dcddfea10
z705705fd9ca74487fd56adf0ee3a241f932fbe1c11700efe7c949a515d4fa2108090fa2698d709
za548bd217c9a05c1ce3123cd1fedacb528d35f2cba3a81ad794ff9782bea5686425e94b8b6a09e
z9211ea98c148981d09780b4dd4ee0bf819d8ed606fb6d7cb0aa6851fd97a81ee0fd0e7b626a977
zd1ee583d5169acd23829c3d558b5a1936a106e70cdb0353864174b5008fb75b244d0201a4f54de
zabfcf9e8e9135180769b22a1406dd7340187d6f05d49e7f867cba342127c4b05636fb9b12123b6
z5160a665956a432526b34b151c39ebdc64d6cd0b4a832966cf43376ce28520351ce2b725efe4e2
zc7dfd12a948aab370b4eebbe0bd765c70b545af4dddb14d8483c28943f4411f60ac68f54bac478
z6065863c0743fa6faabff9e74a3768aeaf330830ed4d6ef126daff0e060583975e85d0612e3e85
zb48f2efde08f5c1916b3d8be8396a78b74e679f2ed3d103ac7d937e9232d6e412f54b20fd61d02
z85e87c6f557e0b544290d858918b0bbcc672b4073e2387c51c9833291b8e8695be1990675c6a33
z8dd6ee084d3e62a8098e84aff719baec8f78b52bd177308919eb016a188db3f5f01d2e8e12c562
z96e19bf0cfabb3c1759c9d2a0fc3bada2e455a13931b997b07cdf016fbeea2ade652cfb9569666
z333e60187c0e6efa2f60e5178079304cb916f4409dceb18cb3c2c06f7bac86f9565b2ed36da2f0
z3ee841767b6298cfa93780d8e0a796d54c3c4bf936973e84bf31c36f6acdd1fb1ff9498da9df24
zb00616f4bed02d92f2e87a61b682f37c8e050300f881cfebbaa4dadd86a6c65ebbd42990a7ebb1
zefa51a34b42edd58dfec5bc4ac3e6668ef16604a71cb9a140dfb0a21b04cce2e5e1e4cd64c2da1
zddead75886a9729d529b1e3ac96c16b3ae2b622e4e9df35ccedc17169d45dd151ba646f5fcaa49
z5ae0f5536b612b4e3a01f428fd45537c45389a4db10c5daa70b1aa02f3385b9dd0a5b88ad3a154
z644232a12a07498f30547e222c596eb8ff4ee07aae49d89824eddeab4209428fc79425fde19624
zfe78f6f246090ac2133bbe6a881b43fed8b34257ab5c3449dbd47e88b4d0d6c04acb1decb7b458
z0d559736ebfff38f460e3c7e52c19d50bcf742419956f6a9dd51524a96d4eda49eda986c78e3e4
zdbadebfab91e3ce9a9b5241d750a3b7a764712bdc82fb3be1e4b3cfa715d96e1affbabd02c00bf
z84637dc9ac14797a4414373d8e0e9b0df13e94abbb4464656aa5614e485f67472775fad06f0efc
z89f9de6126155ce69118f102d8b1d6dfeddde340211ac2d03f52a7e74196e246615685166f0229
z161911a473cc528b7f6cf74525f82d345164abf906142c7bdbc388cbad35f7f7fe5a544d4f4be7
z2f1a529d51348320f39273ad607fe28cdc22825c9b1357af033e9640ee828427fb73c7592bc4f9
z4ce04da135684b47ca1e038531de130202c4518a83f082be20827ba12930dcd8c8d46a180cf710
z5f00cfc0bd1b5ce629557d6f007c885a78b5276b83af2d09ba1e2bea607ae6494dbbf6d22a9b78
zfbbe9e2db6f4c895df7f3d6a2453ef2bb83dc1d7e85ee0217cfe0788b573d2ea690cee47f0fb98
z9044512485f21b96bd551596409fae5ec1eeb17b37d9838042e9882fe1a69d4175abcbb7c888b1
z767311e87bb365811c863e4a2026b9c734380488aea1ddfa1db39d1b8ab8add64a0b31c050db12
zac6f9466f357d4f0920802dcc0ad49043a2ed4efa29ae579899589a7d52dc4587f586d7890e67a
z1de423c53d62ac03e54d6669e11c5d97b7ffa1a5c63469d6389351a1583cf369190b04960df7e5
z8d353959dc7eb1b20da125de9f4ca442a18db49cc0da28023beb9587b9802532c4974ae405ccf2
z1446763952bc394443473a3efeb546e3e5716c88d86b5bfc372fa232d5976210158c2a754d2bdb
z7280a2ca5172c37034be3a1c54fbf2dbf0d693e48ac57e162d8c658c18ad0e7d609383c1f950b3
z791903f2f0425a9c46fa24f71282dab173e41272fb745a33b207b198549d87aba0abe98984ab11
zfe1c2c4377b2e1c8e29a2ecf49933c2eca652382f79434968e9780db1e3ae88417e93a818d15f7
zf7b2aa7a7ab347b6cc45c354e53ee8c2e59c40339bbca3ec40d4b895881f9f99a8d810ed60748d
zc87e8589fcea99b9a152c31fd94e01ad456026b98ef0841faa0d8f7aa759ccb77a983eefe98ce1
zdbf8abe0c26ecd99434440512a3228976a47a97cd56cdd47e0910bf6fc00e75dbbda5c75b70850
z09de354c7b084db7daa2863dd36bb9683328fdadbcd31bd78e976c53a3fad43eaec6c99d45fe7c
ze27fd6b0970052ba03f4b271926e09d7aeef1230d14af30c9e061690900e58e51ac306af80a6c6
za9245ebffb56c490467980479a18762bb4fe1b41c238a82ad4fecec73060060a3cf79a218fe35c
z39f1f9e220faaa23169e6e8048889c8d8351b28bae52194254ebd59506c064144e70102428f2af
zebd3ec98261e547d79c3a3426934b7716f6090c961261c6e950aba7fb6495c247f25c095bbb2fd
z2f2a0ba65558d984769ac199705ab576d271bce7fc85159234509e79fdffc73a9e9e83be78ca04
z17abc09cc4bff1293cb63cc2d7a1406d416f7bd5cfa6d8be16eb4ca82c1be889b7a25882ba5474
z831ee7fd65016be7d9b10733a8ef2024edc97e065af3cdeebf93bdff8ee58fd8b58b71d43d6407
z6d82c3739e1bbb2f053ac299ae7cfe60fff3aa90dd33fdf685781c892f36b91338120a418fa852
z93dd13eda67e43f51e2e9052dc64db94b871635d808a0aba960b8a047b22ee786b28e2f30d8d4f
za1682e5acc4b206b406dc66e7d445e6c9fb14521050fb38a4dfa0db577f20fb1966ebc97ff5977
zaf1652a16aa3604d0565bda5bcccc42e6738d4ce1f4d2c50827f5ae43a6a3da67d7d42b138623a
zd05ec128f54698fcf6fe1ca36bd31f2cb1fa46be0b94f23071fa95ad4926ba93763f218434907d
ze85a7cff680a86e281fb81c1f1ab200ea3c7035755e2389dedcaa169806e0517d920733760c408
z675a3ce01c9e0a349c87c74d92ae017754f6583db8c30df5139a94deb1fe1eda66ef3feb4b853c
z178ff7c4a4a4a7815bbe5a7bc7f7fa0a21fe2c830c190745a0725e2298bf9aa2b43de8685352a7
z1fbe0c2f227103e3c03c38f680fb707bafe5e6cc8fa7bcc60e2d3ff44caa692beb5906f57478e8
z848279d3a549ce1d538a592b3fe91f2c846725c963af8264da6f0b9101b300c049caa6a1f8b50f
zcdf063e885b990e0696b5e29e9ad09f012f7577ee338f73a6d741f5c833470915d76a665eb4e65
za28ee10e610f6218739672b0d5758af5742b82a08126f805bf830a48c60f12575a5b2f81f5eae1
z7c1018a451abdea07266a04db82e6baa4c6e10c93aab7edc633fe5e5ff8ea4afebba017e57e0cb
z618b44f7929db4228e84036f429644e32d38fd80dd2f8cd011686eba1caf9ba20527179f71a8c6
z08161d869d83e0139c3b19bc9b40770477ea09cf660a672a16fb0467c878c39ec27046ed8f0ad6
z672ec7c948753d95839e3b3d88a44d7ff9a4352919f5b3e4c8eaf050557c151ee3cb6aab81b267
z13a52186e252db98f05df75e3f62a1482233d38c7411872284a1a984f4dc6d20098dacbb63b814
zdc66d9b3cf8aebe43e200c8cb8763aaf2c491a7d51faebe901e75cc8eb3d257cab60359a9b39c3
z7d58ad15a5a1616f6d0955134addf2ba7774cec8a9f7d92e21bc012d6cc0c44116570232cac74c
z8394abedee65d72adab7880ce042b862d2e8390068e9aa7a55e29235b6346a00ebba1fb7199944
ze19a741b213a637965afa21de5fe283df6b87218656e50cf75c206aafd5bcbf154ea1a79d876b2
ze380d154625756302f4743d17291fb2d30a6d7b32d1a10bf54ca1bc79a2c3fd7fce0f89b8901c2
z7202ea06c73c03b4fecc389fe5e1a9db3b2679d436ff1aa1a5c630ba3f444da85cb866c3002e1b
z169743c8ca19f03f4e4f2b4473e30db680dea2c7f27f9ef0f9e164c490a79f77cb90d97f0b0498
z57781386304f8692064de293c0330bc8d202783c005ad6d8b2bda8f0ba7e22141351f5cfbf9b54
z1f0c5cf20ad158fe97ae951dba32f0f7a0ec95e0328aba7aaf665a9c104d42384ebcd5ce77faee
z7513614423721369c5885e1fabbc8de1ea89170ee3d3386acfd5f631a58163fa87d8b7394d3eca
za64a1ec2a2b1b351833c77a4013e5ce0f3e36e22f6cebcd70c29e8452609f22d6177332d5deb6c
z92aeb8701d52190a82dd7c5b33a1deeb20b382e287361d3386a0d2af34aeac2e2b33e008ec9d90
z8ea8173c219c1c6e9409c0d228a494655e0b1cfbf5b9ecddd677cf377bf2e0fa16644816c70cfc
z0ecbaa018191e262878c583a2f8654e2b8aaddd8796528e29aa389a3fddcc40b5f7f16f76a64bf
z1a39e11b29afad3974c20effad6ce863e4a6348678faf75050a467dfc5b36ecdb56de7b9bf9e0b
ze80afb39308a1a730c9188e0f11e83f166f2daeb76db2773e259952721fdc826fc3383d0db770c
zc4008715dbc98ddfc3b4be31e03960339d18c36d5bfb699bce5b222d288a0fc36b9a3afc5660d4
zad693f87bd76335229b72e5f7bc796954c1753136e8e2a99e8bef81f136e5c537633976d7c60cd
z651aa62664a06a00ba6c2907e74310c11ccdc3293f9b951e03a086305be86bd95500953165f1f3
ze19a9ea329a04a4c979fcd09e78b23b35d6e81fc8f46ae661ddc6bfe1fab56877ff5522978e18f
zf4a814f0347c9925c1f4bef5a49e05219411bdbd5b3239270ad269384ea085326ad0f7feb08a3c
z9c699bac89da81b3adffcec4fc11eb4b8a9263296c249988741ed092cfaf5f1ef2484f92e6fbae
zaf84f9840ff8d1c0d6195331a183fb00ca92038f84f4bb076bf241cc1be14f75d866b3ad4d75dd
z87149f14cd9f7b63d9608ee9c2f5b0d576b4966ad782eb97d47503180a04c4e2a504f549752012
zd07e23d76ee88dcca249a77206a10276869cac8f1e2fd9fbc9ff0642e78cb647fb08150d62837a
z2ed942d7bfca25c45250c1e1bf813ecd2dd6d9aeab4df07c725a683794de494034e61d979f3707
z40bcb600ee362f861e238a639dbfe7f2e872cc76a5b67829881acfdb03e5ecd1de2551642ac8d9
z881ae3b1b05d3bac5a98c217f524f3b2ff2a939d3f2783bd45c622e663d6a563accf46f418e03f
z9b4f423bdef8e0102169a4dc0558da8a4b9d93b034613b117316d56699c13b387d01894ae1e76b
z0f531d310e3dc934382bd14f5ff2c6b4ac5596366cebb0acd5fd5c1d9d77190f7e9bea4a595c40
zc6b4938f3daaebcd5263cc6e996e58ff7c97dc8f6fa839646c82cc6afecbfca71fa0530df9813c
z1d39b923802333d2924bd54a6d8850893c47c522beb268fe955421d6c2a0d17c94bdbd9c305dc9
z95d28b7cd2f984aac07ad5e04d0d6ab059170e17c88eb418313dcc559d29e5339c6293e4269c38
z552ecedea39c05b61f6ae2f1440ce708c55f120b315fa244e3dff7f62589355a98e751b8cca8c5
z9bdd9963f9c9cc9ac9ac6e8c7f8c324acd36cf29bae8f329632a0b10cd00e145d6d44de995efff
z0244f351c8955ae769597d05d31869016741dbf8bbbe210e410ad2ae70a4b9001f4a4b2a881f30
ze16a86636c39bc2373af49d617f8f775e37ff47336457b008b74a9422bc1ac5cc507f6ba095de1
zaf17b8b720c2f6e4927e69f62af62da43e7970684745fc50e664b26dc4bda01b45ae6a03c24fd0
zc74f5093eb12b2c0a0f3f8c1a3259b66f852b69d8b99311ab1f12a2564790158b8cb201ba22005
z5a816d4a31e77958dffd31a60fcdae8fa6cf647d2832c8d4117f9d4e2459bdbb27cc7b269fd9b0
z2c52376c150704908ceeba884e95712ed69883a3e04a901fd1d19d260be8a06ced66bbc70018dd
ze7bec5552fe7207b420f63ffe4ba2fd4f4a466533f2b1640a89dbf1239dfa59454e86121abc1de
z751eb381e72e6d2585616f3e043027f6225cc8500cee56e05bfde1b35d19c28d34faecb61e55b9
z419549b5a34c7001830354bc25cb8ee4efa38502019277c39be9fa92d1bb7e2d8917abc3b2f4cf
zebc71ae3bb4f32a8e71806bf0fdfe32f8b5af2fe8a1c5ffb5ea0971077837c644c19cab4f2b709
z4589a90b918652d1226462c27fd233869d7d01175d5f0bbffff2e2cff0bb829b26961ab0d01b44
zd2bcf3f67ca36a2320b0c8d4319dd4d806462ae72dc219b780855b1388809061c93b4694dfe0ed
z9f6aea50ba8d97e43b8b879df2494ba394d22cf004f69622d72533137d8b0bfc74220fc591dbcc
ze41f2c0242b3c9785570a636ea94f6942d11cb5025ebf7760122fab629f8234c24d2994848a4e5
ze274723d0c76539108ee6c7f26781e2078cf95a93cf0d66c8d4d7be38774a089680d91188cacf1
zc4d9a840c5f83a947df65c095cf7753abf9186e20306f4fd5192df941806f091370731d16581b0
z9439fc99d97e1d117e34b8c54aaa2837bb4f3af06586d8047a6e3df0d1295b2adbe38099c6b26e
z4b7287db4c0c200eb70a02682799f86f303172dd4d5f71e567ba07483c479aa1e266bee73c7220
ze2ad574908fc4bb8e5c7b5fe93cea4b68d133528d74bbf14174e0d8708c346516205a2603a4e6c
z4c411191eea6ac9f2d33966f4b330ea34eeb70550524ceacb502512239e52beb066fddde0b2777
z222de4b1f8fee0baaaed16ba7a70943ebc29abc1dd693eb562a9ba0145b2444319f539254dda0b
zc4d2d9092f5e11d37b907f4896f30991477a5ad25627289f732d17c6f6dd9233a8ec9d34d9b6fe
z93ff919438eda75c82bb5169f0d24cbd3a07965489ccc2a9f89ec56570af87d53129ab57f1d7bc
ze7e49d95b9a5a253932453a2ede009f08fe156d6a2992b497ed858eb4e199aec22c80e42aaff52
zd41b40461c64f430e1311d1aac0b2a05cb12584842e7f64d4810d99a4e730ab081c5a9e15a730d
z1bcebb94a8a8e034df4df1c7a4a2beb8a36695985b8d991b6035826dda126811717b2544976891
zb956e35f48a0f83b7eeb96ee0ab053d08354238978bb8228ad5c769557cf2dc35359e865ead76d
z4ba3b1aa4bfdb0362b974197544b0dadb8f3be89f2021d85af9dcd07d7ec481f21c9e6a095561b
z181e34778ef7f0dd8e760f9a822460672d0126ee7bd91443bd4972458edf2ebffd7dc7ae7b5e28
zd23d62ea7643789e241105f45276f3a7acdc67bb8c5915e81910f52e6b2287fcd5eab2b9276da2
zb2d451dad3fad2c4d6d54f513bc2d383244d83133d037d4783e5fa722c820c8ccea2241b418800
zf21319ea4dbb21f045dbe2dcc1ab5059073292a5a318a95825b32ca873b04f28f9ff352e95a17e
z63eb6f7aee6db30529a44248e2a07575c25c84ba41de2e72df4ea703af7699b4bfe1e12a91611f
zf0b9025cb8192cc96efd66758226943062fc800304f5a24c9b81f68315677f20c34b01c26be638
za70c0a2bd7550ac70994fdc00e61d722cc71181176c3ddf6c257271159f81cb644d4178c09a6cd
z40acb96a04547a1a7441e30184b242d133f4cdc8e41ad5e617db70e32fc35ed9627ed3342b1432
z02d736aa3129e30c7cd7b3b5e61bc157649cc5717d99b2d2b6cc8cbcc508fc24033b2a4216707d
z922107dbc36b610f696cbc447734dc8a762abb9c1ecea1426b71d628cfad900dd2ba1f90636739
z2703eacbfa266fcc6f0d1804988392dcc75a1a4fef636f3e7dd59e8bc2dfa26b19edc295b73510
z9928fdd08cefd9d5f1134d9d9b4b0f46b2120be42fb2d74fa4ab4a40d9b703092664074ff7b3f4
zd470ceb6934b8bdb6f3ff366ce9b1cdd0ed2dcbe4e7556b307d1f3c54da0e015097f3aabf47b59
zfe7ab41eb2e280cea4a5576cf3e7087c992259d13f2661cf36dc2d5520c1ec1139c1b4d7d12977
za5cd1c900f3dc08a1776fa6ef993e04272a9c71d9f4360ca5c5b5b728385093391f2c709530243
zfb15ef2e58f8064e43555af0b35fe28e9518a6e28402eb485e2e63490f1e25a392fd76c9faa6c0
z221a856c8af4f308cfa720c248780b226c2449c2422256e9c1d7986b97dcc103f147637465992b
zd2cd0d2b709b360a262cdec5837ebdb8a60a9cf43c8330cbf387c836c14f15247a323d5373e581
z30b2aeb7481239984c250e083568f001e42c6788d20ad3c5911c131ea1b01b9c6285af8a0e8f13
z4df418848f1fe1ce24813021089297d66d845cff7629e3d44e7d081b854c693c67dc9f53142056
z6302e0ca2ea248ad1bc12f7fcd90fb91cafff23753133c1e6fb6c8916822cb8e99b9dd0d796b3a
ze2cce4c7535886d504c3d8dff842c0989def3702a3895a6c5d42391e8b263479950fc43abf7d14
z93aa4880c82f8b6563db89105800ff6f0389e7a2bb75c7c6bd27ceca2b464e0219b65305857c4c
z98dbff3d9cc4ac1984ab17a5ea9b2260153d3d2c8c2f05b1684a23e9df193c5b05040f71040d36
zf52236860ad89cbcbfcc3e9041a6f6fce141f79e168bd47924f3f1accfe85bbc3bae5b53f0b6c1
zf16817c96e56a721ce52182b7b8482e7db924c10f520f086f42380f1091942167f94ef2151fe3b
z4902533d0e3c6d74f74c07eb5dfae3c72585719650fd843aaaccceb7fa3a30516a7016af1aed18
zfa62f158581950af62f979328f857f32dd9f372758b1924cc8285ed442fe06e26b777dbec5d3a1
z89d2e8528a53849e4a77be73d1f5df8a9ededa591180921e3311d10a21c2ba1270f160585e208a
zc3e10369ed2141d03e4571743894c9986cf0be09b0e0362dfe53e4564540dfeee3a3717ac58096
z82cdb1e17f99e1485274b4bd3ac14b79f3b396f964fb75a07d6154184b2667798ee7e51a6599ac
zca971026a36fa053c7c3cf34b2baad6215d3bb96760b379562d31402ac45f05be1ed7bb920a7d1
zf41a7284488d611a5f89b59bff884fd3e8221dc5fac6e797ea41defea91b7a16dc304961e74b5d
z32e513fd7dcc1fab9c8fdf6acaf8577935e015b89bf0daaa25d55f30eba23c4813ae571831a8d1
z9f5db7dba687da094612b24df95b080bc7608cf86e46f4a8ba48b48d83eb5f03593b7aa57810bd
z611845d59c3370f4d19ad8872dfe894adc5c318f1e1295302ed6cb754f4fa4db5fc5781f12ec71
z69e68bd40ab794e7e752d00c354b241f5e1824b23ff83cebfa53e38ee5cf7fd64aeb889bfa71bc
zcb6207a8896a8084247582162a2da4aa73e639ab9579dc595ce039123b8626793386d92366b42e
z5cb93d6ebac0e493ce8f830e3b89e49461904f86c872acfe78f1acf25f05be927ccca79e1ede61
z71977ae31f912aeff62fd931f49ba944aca3c783b7ff4f3df7a3e5f84db8f453cc464ca6e173b6
zbe782e57eb8ff0db2100d6606d5d2c794e0e4e3b9640bd9ef3ee7abc093c007fedfd5a518f0b9b
z43f7d42386ca3e8f5bf7bbb30838b594528837ce8697f0233b081aea9f305138e8bfd7b981bbd5
zd4825b72a31fd9371994fbb773d72e983be611425b0cf9c609feb67684e644e77a290ee1dc5926
z2f5057f6b8dbeeaf0dd20522ba46456ce73a82be78ec51c9bd7a452cb06a7b2b8298ecdfd7bf4b
z84b91a2e81ee8a4760ec17e7e9615d195f09cb7a9bbc79a57a05eaabf1a30bc88bc1f7af40e1e0
zf0e273e8e3f2c5b7a8da096c8da7472f74614eb88e3fa82a82275590efd58d58b88ea54cd31363
z0445b7ef466ec25d17c018db15a28bc9a9a04739cd9086ca4f965a99c72fb2b859934027e253cb
z07b38ba8f99d7d39efcfeaf756e5f82a51caf4d91821b31767593de54525a7bef2ee78586916e5
z34c67b5849ba4fe500739a6ee22973c710701eafc51f5c29e963383e175f83b115d235bbff6476
zde73820362a77f70e417c85013f09274a5db175ed25a2902937b51d0a6800e22e83b62aaca8b1c
zc424a6c0bc6a001aebae53b116bf5892584da32df374f868a749bce1e5649f9d27845982e71dc8
z10db951873aebb3b9ffb190b3399d0f03b01751f7133dba51ac30a0f71d1c49399a60a49a98e08
z02ea79c5f5ca84d4cd8dfe7b599ad17e296c9023125f0f21fd2caa704a2f9cf364cce51c365f51
z770cce787fd6a8326ed2c6b5253e2850e130da24e4cb7df08fc42eede837f0a8bce6df4cfdafb5
z47ef50034c8d3788cc3663a73383285bfa76b5de65a81110829e0f8537c76c6ad9865b3b3ec46f
zbc173ad159780ee74d693fa2692e0c71830c7082cff63025c8a9f8c0edd50d80e10fc6ecb83c9f
zd61a02b262fd97536499469e03ac016e94c1db8ddf0bd1017bdb799f56e578cf0cc5e9601dcf42
z576b07db5f7ef4372e40fc9b34bfb09f60dcb915b8f84aa9c4ae417b53d690d76b187361b66355
z4992eb7d5c94e16ff0d47b7d7f7a22abc0f525d30468b64386af7f0386927f0247337d24192d7b
z85c8b716de0de0eae88bff1dd4f785163e3e2cb4eb97838647cb4b81747bbfdb315ed9700e5ca3
z87cf415b6a93f5708e2d3e3554c11b260729313502005456a084a22520a5195f2dcec832a2f66f
z21219711eee055270fa0c1f8f700c4e4482dc7e70755c94c07e399b297f6ebcbe4e93c0a50fb27
z1b356321142ea725ef388500a7ecf1a261e5b82e7d82d956ca4b6b11029290a241165539583128
z1af562f73affe6b632b7c14afd6fca2c5f283b5108521b2e0158b806cacd4c46eb8912d6146ffa
z21527fc86b83b3d79c3bbf77bb220a5d6c44956c7b562cd2a508552d91d0d66becff889329ac55
z0ec358532fbf4cc847d7a8fb61302b00bf366a93dc5ac325f6c9f3f16402206429ddd0dc0e4995
z5412f7c41427e53ac50678b5b94b8491815166b9ea99961bdac6f56d8b4dc520fa593ee39cf3e2
zb8545e09b290943adbe6cd270f464817c37ca5d1aa53b45fde24ce6f6fcf7a65a7bb4aafeef6fa
z1e7cae440991567ab674ee3af4ab5847f64c279fdcf4c14e76bd930e755a0277f35100b0658aa8
zb9e85df0173559b3cd4a05cdd2cb62f48cfd7b11a06989a747998619e01d14582992395aaab4bf
z2005cd70108f455e56f2491057cb90f6435f7c04eb8aa28fb4975384d42c7f035af9a9ee84f8dc
zf278cc336c26f8a2ee21635cc0eba8a6e77fa2465d14f0d71e0c293eb1df25075732ebdde72fc8
z14326c3c8c4f51b12fec2b5bad3dc9d7a656412fe9c64cb46787effe5242176e899e251be8b761
za803c4af5a172015474e4c2360340524fedf29db64548d8b1314561630d57b58e780116eb00e7e
zf64635ed81037f539ce7d132cc6a2bd650dc44071363f01a7bdcad70e343e9b8c4a6a7342b9764
z1bcd57ca17cdbc43eea47fd2f12fee14ed30b3a6097e1a3b0f418d5f5b31dd6a3dedbe1e901393
z4a188c095475d7c141bcd480a2abf6c8c70d109ba5a3b7567781ab574511d4f42b4a1538fd76a4
ze0aadd57257928f44759d4c410c6c70384938bb153e5dc18c7484a63c4f658fd819c564dee8fb7
z6e3ff41da734007dfef3c3c116d144f03aad4488d88c8acfff7b39003c0e6b950e9943b526c137
zf4d224bd146bbb4f842eb0ae79b84a864a381308b6ff3b0cde33367fbe34fed674061a41441adb
z64e1491910df70e6599f3770c01d434791585edd6b90f5f7546925fb5afbb0e6d51278007c509c
zd9e747cc02ebe682bc66b6e0e2fbb9d9e3b29f78beef19a9fd6ae3efdad6051e0c8ea0f74eacf5
z0cb5d702f2192aec45737a891032dfd1a58857089c07b8ee5ccde5035edd1b9d816aa5012d151b
z36d32087198b66c77be16393779623dfd3ccf635cdfc0d6c53cf0efddada88f0c42f11f0083562
zf32cc2ead30a162f246d0705178dff3a2fb4599f9cb6f5cf9f6f184a7d9eaeb8b35e937020a817
z8a8b5bb34c42877cf2b9a7b0707773f483af1dba7538ea0220612bcf1cf807bf4cfddd43ee04b0
ze738d9bcc75f81290615caee50b230bb442bb78e9570427f26ead1700322f96745ef82d594915e
z8b3a3f247570bf614d76451db3553437a311d9d159d7f3bab90a189feb7cefaa23581d99608b8f
z9d82c83fe0bd369fa29c4d71406c5870f702c3b8e4bdc835b6efeaf55a6c9044c572512a743354
z816d20e507dc3bc444126198cccdcd01c7d462848139aef83ec88cc8cfa633908b344ddd3cb539
z3984ba59ba8ec496a562d44d569f09d29ebacb791c58f3fe11b2660d5f0337efd00ed327b2aa03
zf4146d2e8fc55f09a015a704de573a065ec95d9d714488741e9f3d19366858164ba75d741c0030
zbba448ef9dd0edfdac976707c5d1c16dc39ff67eb07c02bc913d840ee9ecd80a06a1d9af6743dc
z664bddd8a95262f3ac7191356563099cf66bac1735cdbf9202d31c3f4c758ce8dc1b6dc33aa373
z33c5c5e21dec7088ddf20ed5b1addd57c9e89f47ad57879d1b2ee010216ef2578efa7f2b99274a
z1452851463ebd4bfb8c19903e5d63bbc040ca34a14aded49c87b753e3607735c7e689dc9b6211d
z6dbc673e7640c882696a23d8f17005eeb8333be29b17956d4d6947c62be29a6b9dbabd80aef0c9
z18cb7f7dacf321bf0ee83f57fed4bc407d5e7e3b881f53c212fa1623dbb6c05a12324ee75e7031
z3b66bee391f98c84c1bd515cace552c5f819ed3c8c8b486d042b8e75bd308c808bf289081e0bec
z1a18d7c9b77008ab2ddf85ff20bc579e53e7fbb99cc57232b0337c305c6c0b19826310a6a8e566
za586ddece1487efb603ddaa6283c0088d15f8eb5c7caf1af9fe29b99dc2c0ce886a805909161d9
z9810ba6898de2d44e0cd1358d1688d66d935eb7a25142d0503e5fac663f56875b68c17887eb5fb
z5074b653b5a84203ecdcd22f90aabbe9ec558a6b532b49784b440cf4f3568be627252dce2c1e75
z4eb07f8de47481d5c81dfa6996b233c86f0098ae3220acc78f943c141f2a3534308d19e0865c2e
zcd21a64dd770853be0c3ffc7e268fb6b476510e7c9c7977d825221d54f020c84c2e18e3cbf35e5
z02de4e8967015716f5a96df508d8fadeb3629bf8015df8a58013c7c8f5c997e34b2ad73595671e
z49561dd659bcaaa6f709a59a1ee0fd3a9ff76c612a4e18c2cfa1126bd1e57aa32fe0f18b877779
z5e17b87f2e759b3d05e50ce00858827d9b1df08ad1dddafc2551238395887d993fa7edfb7a7bdd
z388269324dd5763ef6b199101d4490ff53f1f57d4a6409b7ba928896bc8b93dcea0d4f16a73aef
zf046395011d8678acaa49aa8e3ec4c7a8d1f7d1f55de07c62364369e7fd961265f9d8306cc31a5
z2a0d1593514f62560066f0f1f14dc338bc9443cec23e531307392b496c76412f7abc8c330e5026
zb40fa0d9c0162215be0dedff28ade86891830645924bc3074647bcee9ec8d780f4bff7822cd041
z42a38666ba9457eed1e1fd1f94a01fcae29f1c818f737f3c4911afabfae91e1dcf3befc9cf020d
zfe99bfff82ee9f15e92c614a68e5b8112a9e6995d5f40478dd72c2e5713aae69350fbbaae97d9d
z2226996a6e6dfde6f3bf7edbc55c760dfeeabf999eb878f0699bd1e35e7f44ce8efce58a27fc84
zb82331f94cf3c57fb94c72667ecf20b1f3d6b6109fb55e0e27c1dd5163e756229ef2738893c2d7
z4f62793f006bccbbb3cb09ea8e243e50147438dd4c8ac779abd9922d49b79b9e8057c8dcf6bc6a
ze173ca72b3677a0e0ffb033b8eb2ec6842b4ae88f19e134ea1dbdef12a52e373456866eb3cb509
ze12857dacb51571f20b232e99890264536eda0be8e00b036cf55beb58ebd48fe69deedfb5ec653
z85fae5521048549d53433ddff6f8410f4e7bcce0aeea9111c21916542550b78fb6d46bb3d5982a
z872d76581b4e056c7e92c562225679ed817ce3475b85918cf535265d40393773555f5d15543fc7
zcf9b61ac78204d2910cc81a868ee5af2a91c7f93c77b112c4ab8fe0fb39a1b95ae21e272fc88c6
z403e1be242d720990f1573f6cf7d79b84221905cc6217b6a3386615ffc9277cfc0c36dc30c6176
zbdba8a2fd3bc9c0a331a5ebc945a9b7eab61724cf8ecddff847cd0893a1d8753c23693c6e43810
z1e3ad8f4d293e2d78555c173bdec0770dfa7363ee2a87fdd2960fae3d7545b10330ef8827632d1
zf255c9b535b0411a13e6837d95c285929de1b17fbceb9b7d64e667add760f2f1ba12cf43d49193
zbba461872b5b5a25393885699499ceb5b9231339ff6a94c953347dafe0dcadd9a5c26110b4172d
z4bd16fd8b60a90c6cc1777413713af7ef0969a64b79d8a1ecce02f4a927dfad4d0835c38db7369
z05c446cf6e060931c1ed79f2471770e1e3bfdc6584c8cf7268d99f6bbcd529f6d93131c8822a59
zf2f6770a689b279892fbc400b9648d8023417f453a27faf9ccbd6046ca58ead90652eef28de2d8
zdaca228e9c1148340ddbfcef3cf73a8549d6c6c336bafe141d29271233de43c35f294115cc9f04
z2ed2c53e6af66b5320e92df2448937d0d1c53fa73152228ac81635e77551f3da5ec810b6218c1f
z5ad03a134e1a636435737ce8b919a41dae62c780c04c7f3522df536e374bf5dce3a26b2b9205ed
zf25f3fca17001dbbf7343cdeb5dbd1f78fb869b12618844fda86fdcf92c1101b5d680e2f18f1fd
zf86c5b0406fde7267a5f84f58cd6c603d9238e9f2cc5e4e7b81c71544312522aac1b456c2ab576
z42e8d39ffacd17003d430c0a09f833b7632c39af228e7e9951db82a2af96ac5a42973dbe567651
z185b893cfba1b84f282f8308e7ee07b3dcf07cbdbd4f2a1a3c6142c8250995e5c39b8912f19794
z2b5830661f8bf6a8241bc55d2158016cd423c8fa49e268049c571ea246f8740e9aba04d15dfe49
z408ffc85e99d96c0dfbf07939b5b8231eacb667dec8dab78dcac1cf8539be13f6c15f075d8f34e
zcead2ae09e10625151984776874a7dec38db9ffa0db9f8f27b33872ec4cf9e678820bd9898566b
z6cd2f91d1044f7de8a8c8c4f7c6111c719c3d361c43cdbec92a5702c7de83b75f5aa9a6913b2bf
zfccfd63eeab3263c3c8352a2b890e94662583f17085f469b24b2458daef5bd10ea9ae1e48f7395
ze02004ea3975ca376aaa9698c5421df1c4238b8a4d408bb88c96dd0f533a8b4cae0f4816533944
zed3a011aa4bcc6e4ed3ef7b201976a32041d6039583d132323697b12e30e7e0c6f9462e0bf2440
z93b5c021bf68418519f612ae46661d53017234b1bc0f51338c42539379cd0851ed2e97d7d0912e
za3a30aab40ed3231963983d7725ee23fd5395950ff9f529550176835a9ed8c68e7d33092be112b
z0aee231a63b152879bf49ba3fe508523811e98a6686e4f4b43c2ec8d0acb829038d617f736c890
zd3f9bde19e82d2638438c76c053f67193b5b2b3f603d761ac0f695a45d175d11034d44fe2a38f2
zb6bec789cbd11d8404c7b8c1e0e04031387f4ce49ed8cd965d312481e6e2a8827fe124d4a57ffa
z111128a5f712d8283c0b0d05b7367a13c789e1bd279eb26c59e431925084ed27e6d700c7518641
zfe6e016e3d85ca2ffd3238a15feb23fc262a37ac97949b3a0e52f1518946013f4fdd8eabddd403
z65be2995f43b6a15e720f787c135e571d93c61c66551c9123433df1b5e6d1781726154fe9100da
z03f3ec7a0e1f0bc5016bb74129c44395bc0f21dfd209aafa86b449b6e0084e02b9568b6967fdbe
zaf8c8101bde1e674d160a57cc1335bc2d8bfce685896b259574cdc3bd2c10f28cb60aa36ca0b33
zcfd433c83c65b06753c274857b5f28f455e0c30bc6c63f0772ce94f56e3476396a439c662b6bd5
zccdc43d169468f1b1ccc7bf4ef812fc3ef62f654501f60c42866b2455ac8aefdfc138df23babdf
zb974edfe920ade0004db342ac4f6cf18068c5d317d7ad757fbe3f32fab4e9391841edab5f03cc0
z6c477ba131fd820a23a6a3d541691124aadff6f9367002db91e250c2ac25ea2871d126d518f23d
zf7f4ed45fa2f9aadd13f3e32413c9e3231341d94ab1d30329e5de15f007210f45576ede7d98b1f
zeda9ad52677bce61a95ffe1c778ba13f05b0a67c56ddd6ec851a0ca05f7bfbe1df4b1120ac9134
z5133a1e3cc1fd444ad0babc4dbc2083ab7ef0519d5b0b462d5b321e2e4e311f83f5f084d044290
z8cc80fb6f67fc8c97a80d4a1b016c76729ccd845a2c3bc77f838d8e5d6609089d9c6d628c3026a
zb5836316a96c722d5003fa7b7a4b1660b9c2909bd367052eca4ea3eea0093d84767e4df8a27fbe
zfee28c55d0812fde4a848abfe2d02ea9ad8851a53c9be1862494828d915da729987a1b52b52907
zcb017f47f917b968dee3a5a1d3d2c9fc2b5aec7c05fb111b3a32a0cfa690d5132de94a85a949f6
z96897ee4340ca4fb18275823d588e332aaf48b859f5d7b41541cac1aaf37c9ec3575800f7a6d45
z095807878958293ab63232f6a688dfa7c67ce2d8bfb03f4dd4c6036fdc8d07afa3896a58b54dac
z9640c9f6d014877ef8666435b34e193c108c7c3640115d4f262aed0143a9835f88811a38023f65
zd63466a7ba26e487aba85b515045ee49273f07f187061c307ab433ffe2144fdcfad6c9ca033264
z6eb2f72e6954bc9e283861fed8b0abd530d08d01a95f710574af8030b0ca877cdbd34d0eee6a59
zf09b6ba78ce72a7e2c02ea7803ece3c110a6ec3ba37c191325508455f3efcf328bea4ef336cc11
z27416fbe480f0fa56569304c84c04074b2ac7fc3e3179883e5145aefb51da0ad7f55c71c0cf4c5
z75e2645a331605d3627b2b8a156d30b6068858723668a54f503a84897b5f1bc548906ab3321fe8
zed65785f93f17d53be86e8b375dc28f7ceadd3807ade2e2c5784fe42710a599f97982ad3dcde16
ze21e7bfe37243a439d5209fd691f5144a6b6cd766158d6c3013c90897c655fb653a696526d1ae3
za85a0101cf746f7f49cf8387402242f4fa11f5e6ecb44b19fd2f2dcc9cf8c9a9a50f7bf1d28c07
ze2fab4bed50a2f869bc785b395afea9933dcf0278bdafaac233704000cedaa050fb68321642217
z841a170914c434a3dc7e8a9f3f13f4706d8e60a4796173e0b363bf347c97188e278879bb0221dd
z5959952071056d77daa59907f7e7b568714e3741dd93ee85e7c608715bdfad1c41f71eb219834b
z8805c467eef5f657021dfce873dcc7158c9ad272cbdcf86b6212e9c421ccc73f30f430dff78ec7
z19548476b0c5d4bbe7c804793163f0d4c049a4b2e1c3b34c2a2e6a02fbfabb5c064bd7c17c1425
z89d31717e0cffdaa10253d3ec769e376b04926410d071da2db559b18ad708c9ccdb4dc4b7ba715
z83f2a3d9f6ecabe8e0b1fd6021a3c8b731b07f91341fa2258d4c0eb54f29f01cb17cc9b165d56a
zc86eaa46c0f1785b328a73eb2260ca57f2edbffea58b0b2c95097fe0b6adc176401d76522b6dc8
z247bdea525974eb7f0586925dd7e5f0c83af00717a046ddd642744a480c8a8beb0c4ecf5ceb09e
z37c306dcfd4bc89f956055697aabf234825aba87f98036aeea78430cdc7e4775cffcb99a744597
z9c71e9b173dfcd81261f5a7b538ca1269bf97c5e3062f2c21597eb5d1b4e6ba072185e7f1e44af
zbfca3b6399e03deda64fb5ff418424d955ab81c9d9c654ad826b99c8189c2bb6cbc92d45362c54
z4b2997e1ed340bd713f125de17cd26fdff9f28831d56040e1edaf0e248a6a46158c8f215a4989e
z822415cdc6a7683ea082d6c987c01bbad1ab52ebd969622302e16b3a13a5215a4e9701d5e98d9a
z7f2c9c9d6bb81df3d8310f664c32c94c9113ebd46f2204b3722a944d339cea1b680d3ce9d2b3e8
zba9ba5ed113e9a46ff6fc48605edb05e6ddcbc4dc99629ef531ba8d41670dc1177f7d9c6e87b16
z4bcbaac46cb9a6130f9d95a1844d493a5761221dce2384c29d5621a610db49fe230e5c71ac3cab
z13d8f3530794262830c957cc535b4a2253a16b18017949eef6bce65bdaba76299a42c355f297bd
z9dd2d8d725f3fdd10ace7b27b0a7f92d0b3d073c461e27f26a3cf8952186fb8ed23768d41effbe
z3497e1a8df2b16ecf3c54654e74f3487129c48cbe941b3d76af8a08676352b1a210f88616db47f
z2551aa95f36477040493e068cafe3e31c86e7ca785f5143b388e86347b80678d95d68cec239efd
zbecd5f2888b0d1559e2647115a8c537880b8d524a9c9d17150aa8fef93db79a5d3ea2f87bded0f
zfcf028933c6315354d17d6d7c660d2af0cc03d01212418e0998b0766f2ca96de7b80cf2fc81201
z28935417b109a0e80e3d49cc555ed4eaa60baf0c7d80724e2b98a99735d4970f0cf00712632a81
zde6b1a4478d5775214e9302c9c4551c0bb75650330ef39f5876daf0f085a67cdecb6c87777ca09
za1d655fdbb6a91ba01d3c3ff1406602b77e5f262b0dbc6218647df4023a9874b947240dca457d7
zdcf58fdac1064d1f7f704fcdac2f5dd6befeb058df7dc4bb5c37baacab147f02efd3f907853595
zf5747c4845cacc7b3d32d981c9f7f0b325a86d9f872a4fe28abd7498be62cc1ecd13ee579eb632
zebc50591815087074ae8e9c4e02c1abf7b5cf7e19eff015bb77506665660b1eb6188e56402ae5d
zcbcd7a936bca9419cc787ae38e4b70097448c43bd1eac8b718a1d1c6ba7592903b2ccb93899269
zee8b5098b2d4eedc2d22adac7606e2d2af6a215d378d0d720b3229d5e2caef3d9e8a4d22570150
zcd4c2cb6b114f4e5dac9708c7afebe3793b7e53dc97705bc76cab11efaaa8876261405e12d9396
z45fe8d3571bdb5e869a86d0addda300b0fd530d22787172b0c3bbb1ce4803a6e8461effc3ac945
z285b5e400b7a87787528da1e35df60017cdb54de4495079317aac2aaf5d884f87633a97d7f3b73
z272b45c90199b79939f864fe7296060a4a45e10eecd020cfe99aee412d94b1ae3b6ffc1d6e4070
z14884f0595f84575f81a4d95f2c625a243a32acc249e1412198ec1469c524eea9c886a0c56b4d8
z4710eb021bb9903de5117a159befb9ed4d5a11796378ac336cf60e0e31204851ed9825e0817ce5
zd4a0182a64098bd6bbd517a63b7e2cfb6893ccb851bd983c10c09e5ae7090f8439e4f816455c81
zc12095495d1cb496434373b002dd80cf7a47a1aee270f95c3f2bb42c9861666e271565894cd374
z1adca992db29cebddc06a94e149a70bbd14a8b68e3a324ac350244d15064f63999064f5a4b467c
z578d441bf82a4f59a9470b1c3a3ec797b9d8aa1c0bd8a0dcaffb5c136af75de49034b747ae00c1
z097605ea2207468dea5387de85dd4a0e344e6aca427f02e48ebc82fe7c0f3daf87b8461218db44
z3a1fa1b6fe021f40014b5b147412c18bfe54ef43e4e7dbad4b7aadec5d31492fb71d9cbe4d6c5f
z84098058d80368cbefa8683eaf4b4db8dcc6ae8bf8f08ad10aa8f4dadea221afd2ce93b9336096
z773ecdd7d292f829651dbad95a2f9f1e14f225dd74f128c2e56917b66f000249d5bcd3bf9b6475
z1ec701d372ec957c76fd75834421407e086437adfa920f4813e02bc757f151d390b90888498223
z8252585a862ec1fd726dcb3e11c91760e7eae814cef0746a748f70f9b0d167074dba3b74ffedce
zdf32b68b1fde3e8c7ffd94f840b025bf1a29805ceee349e6546f4770ad808b819b3992a99f76c4
z17d1995332c2d37bd734ab61660df86c60a75621967ed3757b8599359036b0a6fe2acf8d283311
z9ca1d611e4de58b88560c76fc6f3443efd720edafe65d7b979869058d46fb41e12579d92041100
z9e2f982b5c14b1c3790feda322ff74c90e998bba56ab96b5527e41201415aeb79e53de34d37f52
zafe5dcdaab147ac2ccac510976870728550a735ddf8ceb710e7da84dd7d4954a316f8dc0d51eb6
zb5e5af9d5973497ab76c791c1d5c2b301afc9f69b6a366f8085dba3d67a86e169a8c8a1de89b59
z7b520d2dd33a420da2f14228c60a412bebfc88fd10f2e2a2a8de1a5d6854e0c51542b3ed1eb1ab
z0f4348cd4c1e61752a3b93f31c80b7281b1d8e9f7bba201f4e83fe2bd05e10e7091042d60207f0
zcce8f0b7c9fed216c011c0ae0b8bb58c06ce5b233e20dcd65c472e0e6800b00408253e8e6b87f8
z0d459d94aa14e3740497d8285926ab849d15b05b9b69c5260accef911f3635567602004d9c89c1
z57442b4eddf791227d95409a62e6c94d630855f7c82bfbb915bf831dd89048630fc7f947695463
ze1044c9b16dabaf15ad66b112949f016eed014edee6a53fca647e72370aca812af66b3557fd44a
z23c3bb96295a79c1c688dbab5c7481e0a67bb1aca8af8da4e09686b17abf5dc6b9a5f9b0182cd4
zbf337bb1b66f0e9c96c840bb78a3d620b6f4ae7483300c737dc56ef402fc4c34957d235b01bb3d
zf9e6f96f1a597569990eec65c34395bb9833a5b0d1559e945251b3a2ce443aef7249096efcf753
zbc9725e7ee2bf754fa18e0f3ee3fe8441e876e4875cf94d08237f5955ef8e3d47e37de9e9a651b
z01cc5a209c469acb98c55cec72c6ef161aa49de6819f4cfd229f8102a9a763526c3162765f9316
zfae77bee8c839b5d1ebea3c4e744a967204ce5b95652b76cf718016a123a4949adb8a45354abab
zdc06cea6442ea46832efe60453c2c81276b988c94e0af840bf533a253bc6664c8ef4b30c0049a5
z1c54895319117c1ebdf74c5908cca90cf4d062d5c333a27f73dab90eac74d82bcca029610ef490
ze5af9a29c7d05cfe20601dea9d79c4f1f6524d403039b472fb2dc9d1e5acc2682e95691158f96b
z065be3678908f647346f2b52e8c59de633b0bcce2c4685dcbb9e7ab3ff0dad98ed30da05bee2c9
zfa6b06fe193ab5dd7d0e0e262cb50713df6d441100c679beea81da215eda82867210d23498a35a
z2c4dd921f51c3826bc9fbf6c31c19f1070ce922ea2a4c88e47e7dfe946b3f681822e80081f52f9
z6d3bc23474832b73499ccea2e5e566b199fe908f941d59cc7870d9f5eaba01bd655bce93d323f5
z0a8db0498d623f8e6db87557678d6fdcbd73131a2ce4f932fe2610643736aad4f941f70a50e0b7
zba127ce5155b766f06330bc0c7dc6cf89c5956793da5a8e01ffb86c3c12e7df9b1630cb40e113d
zbf064922148f55839cb2168fb58e6ec17e2ed32e904c70a24f582030c5c9202811a9ce21a7006f
z2d667a3c0aa22a2494e9077f8b96fc63a19391a9a5772b33e45c136ea6150545b57f14c0cb82c9
z488d285592d5b0d467ebb8beb2d5a34cf9d42e52b7c2f11e5d5fe8c6f024ed8b82831a26afc30a
z6242fc1b99c282961ef8f8c403baa5bffdb2e80d888a411b7a769de0d291dcdfc63d92eef0df7e
zc6b6fd186013153928fa409f0de3448afe139a7889c096568433ca995e8faa09f07fe90d0529a2
zfef2095b6933b0cb71ef2834d188fc232556dec815f8272fdd958ebaf138734ed339ba558b4631
zcffec6c3c2e3e24f3865b3122d145bafc77e0a8db1b0bc2a3dfbe400aedaa118408c854f4ab4ae
zefd924ec378a7e691de037063b36b383bf874f98d78d17739679eea82f325631c6d1986c6e3aeb
z6fda18325c43c41e2c73ff8e7ba3be5af988a803a210b5e03e51d350ce758ba3492d860d91c79c
z4da470f9bd698e69e44cc9735b386fed19a7013b4d4af36fd6feed33cba0eee1124e9a0bf0268c
zde81526c5b3347564c9e63d4e43c9f415636ca7e08812af2c5b3fe611add8ab1b8440e6c0b4e63
z249f758e1fa61e8d4294a684e0440a14861bda9a88a492b677f6730513530e10e9b5754b7241ec
zf5d6b253f24e9624633f9cd08b195eb5786009d718250659889a2c221c7145f48ca9173ac9434a
zc391ae2173b0f09ab8bfc290905dfcb99bb7519c21873618768bfa9469f58174cd6bb3f2010879
zee4f8f7727de0bc235025876f7f4ddaddff4712479a14e839fca72533f47a22c17cb4609df3530
zd6bfa94ece1bf7905c422e8162262365397c0f280c6d2ee5e2a3d4ab220ffa28edd25c64623985
zedbfb80f7c5e18a9f3adb3a08d7025efcc7da2a0d989075b709abe1dd3d1f6dea378917496be62
z65bee2eee8defd433704755c1d181f8360e0ddda67ba761824191d8e57ebec26a8da1a8d05e95b
zebe6810e86a099a7a07cab0305b4d6d95803197f9d86eaab035ccf1bc363678136a950e3ae7e7c
z375452577ba2bcf22e56e31fb1930c42eab00ca2201f5dee13482fa44f9d5b31207626885abc81
za7ef1a9f099ffb5e16b7591e977c1c6d01623bc59a92c2653642cffd9e0cad508376d779cfa6b5
za715b4482be681827e7bd8001de25b7fa5aacc9edb9ad83b405fde997e354fce00c6bdb9604883
zde6768a1d132447ffc745c253bee3a498f134bad4cde4eabfc95b4ce00ed93dc6b3e9b1e6e1b7e
ze4eb10228357a4d0729ca48c2fab1aa3837383581426e6d68de2be67ef710f0365d153b6987867
z4b23ce7bab46daa01f15bca94cff4458ed628f997fe4362985634be5f6e3c2d3bf000b078257ed
zd4dac9415832f4130e2eb0d410fee638777f4116faeecd84dab8f2af9af404b125a4bb240da5cb
z92a5ebcbe4511c921dcec638336b6a8c50d54e7dedbc6bf3924cdfcca67d224ebcf6a880153fbb
z1f0a3f2e3f0a2156a74dc108b12e47fc240a76a04c1120c5a7523cb8c319571a5a38d99bc11dfc
z489bc2b2b6a4bf3051b5e471939cd2c746cc7964a56352172e06fb65de24a03d81574a9f52289f
z3de09bdc4a835efba3486b2f4a814f655b5eeab06dc503858f4e89d48b415e35f337b18c7aa00a
z4790409f3dc0d1103a8c12d77daf846da433d706e83bc253787d20593a5de4ce914a870e53d1d7
z8dbece07fb2ee05c1e64308a1f3d540fe86e4c7c6bbe5d301b230a3805e719a849075e4ecc8742
z0abdceeab4a811838dac1f929f84fdaa446d4e1d5c7b0354cfad20e358970b24116feb8934ef73
z8c70e142173056316d78480fdd3361f78dcf1403b0c174bf1f673f0e3b55e2d3f062ef043c1a2a
z2fa06b4b858aac0aef409daa8f8cafd813836876c587b6f76a69260ea41dc7c72cd42bf44ac9e7
zd0142776d7bdc7dc5bc12952c421615724da756978c9e82c87a8fb88a7e9a0748255ec5af96b9e
z4635818e10cd98d6e49bb7a5f3fd24b7625c3db6572f8dec165f2b8ad8c0fd52aad1f99040f191
zea6d6c18fac45122703818bd96d9864fe1ff611693ccba7e1d32f56c0d9f362158643943d04974
zc495f46629b05fd3ffc5ab362ac04ca789deeef3017b8a07e5654ab19095154e7ea2a4e0da1d68
z4210ca3c41c4933f17241958d0ba335f41ede55ece6ab106da684266bab558d7f3896535543c78
z6a1cb51778ac20c3c004de44809b4f99388c15e1cf5351b30b0397c60a882b9033df72a427da05
ze94b379e6de737fa828e596c9e33ce8ab08412d857c29752c32f647c2986b9df793ab448683ab9
z3314e1918c39e152f5ac88ca333d840b850fd750cf860358a59f9bcfb432313bb9466e08d82388
zce3f835eaa98890933ae0f1eaef5fc610109e39b77cb105cc446236db300f11c998133bb5d796c
z352a1d6f413a0105561452f720d38050df966b23d76ccb9a23fc3560a802d1668eddcfd4b532f8
z279d54df479e88e4ec84e4575d49ee79e419a0b031628b83de5e55b69a854c9fc25a2073ffc47c
za50420527372252bed7ed5a0fcf66c2cd3315a915ec6e56703fe796df20e56b748bf237516c114
z1cf8da0bc23cd44c42ad2e741f7ed38a5254501fdb4c1c6d76a144afe6a2feffac0231cda45cbe
zed151442b57fe8124c7ed81ccb7d55215a20d060ab72baea3879b193e63a178f1e59015c2797e2
zd484fd3352787e405789607764f700d01c3ff2202b39f52d22b24165290da5779632f0d8cfbee5
z8e4e3cf2dcdf64252e786f179a51be8d1324eb58aa44fd702646969f00661bfd55f36ad14e6400
zb721b90a34e11c3726cb61479a91fc1b39235155c7c189bdade308d4b29afa94421691319a403a
z08e1cd682d4aeb2a9ee13c0b3c53a68a88bc8392a746e2003a74087630825dd75c2f108b503bbe
z011b297a0ac36f3420bbb0383510fdc30fb594372256990ab7b32f808fdefc47afd2b2e802a170
z3e43a2ef36a8442eeecf7c0e107fbc8e5ae53ae9b5b8f1b853163267da17439dea959d0487d26a
z5dcddaed675f965c02bceb2c56bc1272220d358a669ee36886fe5c16ec75154c99cae05bc10371
za2be31c45dfbc2f8a7c9886cf2ef2b31a8ee3511e8c4ce5f856dc9281c96dee88209011276f205
z824dcfafa455b3b08255b8f4db6b359ae476fe375d2eb99d23355f76a27c934595d72046011be6
z68971d40ae3a4ba15ad88357f0801385a8f801135b161a5d588496aff78d0c00824fa727d42858
z55f8d7e46832ac655006454dd6f703f345cd3d9cc3bf4b0cf761f00f1038a26ceb44acbd4abb04
z83b22bb89b6ce0c912bbccf2382bbdaf9c368574ff622f634cb968f200488c7a06c422018b00be
zffd02eaed2c09bb71a48211f253a153720823a984ec09718ddf6108b7473ebc533e37f0e628fce
zed3d06b69bce9965b1188e7e54f72883ffeea452863ef2e574401ea2664260a3a2053dc3ee0ce2
z746934ce2e295ed312bd7a827b9e920dbb3a41a5e9c9fce48f028ec51578ed56aaef106f3303f0
z0689e66eadde7bc3ba313ea187ef664b584224f12ee91548955164558baa8b887864015d6c4e46
z8bb45e7bdf4757b3ec428024c88c043432e8b1b9dfaf0aab87e940b768070a48751df085b5c879
za7e520cc474a8fde1783d5fc98784ce559b08ee0920b18c2d785d4ac1b2688ed3c9da5c651175e
z45f20a7613730fcf2eea518f49f31cb5340b4f8c074b415d35a1aa2634eb31133e0a0642d6c492
z119b58436d8d1b505bb97fcf4835fc2967bcb0b36cc88a67d3c1d9a2ecf53be6eb17ee7ba49ab4
z8cba3ac7327f3ca000181be48e03f197f29a814be112ebdf33295022634b5a41ef74f5cba71dbd
zce969321377c213880d869eafea47511b2c915b9b0d513f05380d71319bd191a97a500181a5c90
ze45e7c8801167fb7f1e19dc5c7151f74f4bd976ca88844bd9aeefed3eced94111034c18e8ab0ee
z0616f2d6c023dac36a9fdb7b55db932e34e750ec71c9a25954c7da5d01859e689e832694b3065d
zdd3e95989a58ae1cf29d550ad248e26441c9e15083b1a879d653e7a70dbf0de1d849085ed1d09b
z6c229a78b9ddcc1fcf387e3c427da826eeed308d7e8eb2f1efb0827bc4252f545636934a0ff7b5
zc10fa9246aca6c854fd4bef035ccf393e5bc17a19143e86289cc11330944c6ca95897c130bc915
zcae2d291f7d9469c13d5599db554f4135fc952d75c68f9c4ce5a5de8d694582f751a2b7254d228
z0a2cb271259840384570ac6579566e1344d49663762d8de0556f5d92710c4cca3352afd8f81746
za9ccd4d1d10fa1d447c8877333ea4cb629a7eaf50ef7a5fc8fec8f253e8e29208618b98efdfaf2
zee2698878a88319f2b10ba18e6be55b1b998d5ea7adef4cca1af1a16e3dc6a16d7ab860821b3f4
z39391f36a007b07449e241e92dac274ca82dd61a07be5345e74c8fa628b6f5c0f6b67d769e674d
zbfdd8565db81b1275e04eb59f57c7af9fa8236eaebe7eb0553a5dd344cb7f2607aa013e6847093
z2002ad2dfe3c760987f1286d38ff7a2ab489ab1e7547fdf56c7db2481ebd97b836c1ebcc6b2a4f
z6efefc1e109c67f479f43098363a96f2189c16e75642d4111085bb76f55de59c4201457be914fd
z4e873d31618fdb3009eb20feb87b8a4953e4c81e90b6162d6271408010d8b31ddf583be1d07e24
z8b9f1bfe385fdce90b157716497254df6187b67bb84dae2b64c43588442213ac957dac16f29468
zb928b380fdfa1b9388c3e185e24cdabeeb5c656f515d8088fbc34fde06eaa33ffb6704f69ff0bd
zfab416832e4c5bd4a8429d981caa56bd4aa6266201f55ff6abcf30a6167e141edd4a50d1aaef59
z7f8e9176556ceee7a4cb0dfcbb13273f21d9d57e88fb6ab9797fff66c9abc6995c42b02efdeba6
z82fb9814a460494c99434e3417c7f797712d219999886337f4a6ac7dd95dd9d9cab0df242417c9
z29a3b9666cdc67bee58bf4f4507ff38d9811250bc5dea5ae2e811a9b148be5505b2c4b00eb40f0
ze1f85c4e2c434b44b039c2ac50a6b9b702c4667bdec97f35afbd788d95ce3494366dfb9f0e3275
z581905ddad2e5b5513953a66350a1cc84cfd6761fa053925abc34f361def70c524b99345f55b3b
z55a92d0fb3c2c6f18aee56d7deef941af32bd91df079c694ab72dc5b3a614cd700a1d3952ca755
ze10999dcefbecccacadddec8827f018f35546dc0b917ab9769d071e14d632db77a3aa09a3c725a
z8de5352b87e3154a91f52027f8b348747bfc0f5e9975edebfa89c65f94ad5358fe54d7151fafd8
z0834c5ef19cdeb3b84bffe7130094ea6598f28bab05b4b49b5670ee023678c9ee5a76388d39c29
z3314a13deafbecffbfb23a2e03b681344fd3101d6cc2a16c734412cbfe22dfc69a24a7c4f5c080
z1ffea745a0fb511c944c383e3a3a15ea17b60910cfffcc64bda777531dcca222f3067f6444c6c2
zcffe4ff4d3340db1879cfc64f9ae229f91ffe0792a3bb6ac6235529024b48131fa2a663d6448d7
z40815fe8195cd9cbac888f00e0ad2b694474767b395a3f6f11dfd7587cb561cd134635f7c24734
z68270879be44ca33824858d9f5b0c9b1dbffa7d2a0adc5ea27f39d9186f127b8929f970c1c892e
z5306cc48e91f8d60991d8862f45f0828feaf8a11f05d9b0d04333cfec8d26f2a3a586a2b394e66
z0fa10a374b9d9e92f7e9bbdb29d351ae59626b2a92bbf17ca30e427b0e90f1fa4ef3b1154e8705
zf86aeed2a8e4019cd6af2012abfae7251bb35133783eb9dcc52d0b88f096a732c3c0e4827f08db
z0f5577f88f31b7fba324913b50113a816a063b23a01479353114dfb3458a3bde70170744265ce8
z867ea6fabf4b6028affdc6dcc17c9d22ed5b840aff0cc7c0c0541e840178317e42a133b7bf8a27
zc86d7dc8505f335781cc78d2c6f3da0328669f51a3f0ca4b46e042a3dbdc120ea6982f018db62b
z1ee031368418c934b16bf36d7582a629db30148bbe1aa2553507138dbd6f48fa48aaad9994921b
zaf681d45ae68f5e384a2f1e68e75cb2274b3039d068405988ebf830612b0ba1876ce4bef33bc63
za962daf3a8a9bb27b96933528b473d107903f694f525d1022471237715f4c668844f61966afa95
z6a3d49b70bd6bb66e39cb743a5531eadda16342507f12427912f89964b963a9f8de6c1cdeb81ac
z024d618d30b6367d59de0014af7eda4069cec219b5f89020db4d538fac2b7f0b4e603a2cc0ced2
zea68a19fc3abb040a9f16dd575e44f915f6d7aed1663a14d43422761c4b94683315885812062a2
z9b70c438ab20182424c621deabb7b0e48bd8c1e46b9ee5dd64f043ca22e039cb6c02a94d02ca97
z61ae26b3062d2b988e0485342e92f0d17399966be1f34a0fed63530aaa7d7135c48db1f2513e3f
z61947417f841099feeae748299e7680a6d76f04bd3a94f4c7abf789051e640d26a048e13276325
z33a54e51d2aaa0a71934d65f86de32dc6b1a86db095d88a2a4a2f3ad501b716e7eff0c1d552a74
ze803299abe41201d18a4d45f64dec8d8b214f398f7806db400a8825f7a3ebc76612c6b1b747339
z6a45ff16d6065e136f151f71348dac4cda173c81856958ee15aeda659a021f450bd80c809ad22d
z96151469852b67cca4500ae055d07194f429273613ae8a0a3807b028bf04310668884a1e21af0a
z40491c1083fd759d81e3c8ae58e062158ff7aae9a2d4cec7815d37f09b469e148f674fae76cf34
z0e72b205fc0f178986e5c9df22a41bf7558a5dfd23c334f7d48d4db49d8d4abfb43c25cfa122f2
zee2ee5a4e15d0547c9da9eff2b88cf041f6debd54730e443f1c41bc49dc550cb5762572a86cc45
zbad268be2a440b5bd1712a2e62557eb6cf2094366a60e382c40a941440597867a32e7658113d61
z3ef4c7c801d0b438e7151e16f7f715a9743742642524029e994b826c652ff328772031ece33c42
z7ccc19d45a1810cd31ab2839d0847648c63c7906722738a6202f0f3fb4ff5ca2ce9cd80c0adbdb
zbc051e643dc482e6e6b6ea6bc144e20ed98a89c2a2bda418f855ddd1901101da872c41e006bd32
zea259219f7d23fe8666dbf814a4df042ce749bad0a7de0c6a699b0268200416b8257632cde6a8b
z9060103155ca0f37449471d9be1b45ca36f183d215783f1ea59c1cff101925052a5e5112a54738
zb9e90d9bb048141669d6c4b62edcdf0aa2dedec2ac5ca9b88c084ca7bd14d7577c8b899ae94d2d
z3fb454d254cf7efc8216760f358c15129b28d594a4ce4226a872fa6b827e13d85c3fa64c7daf83
z98875de55f37654c4eb2344f9b9116406a4710e571f7fadb6ae6dbb677ae5533af84987ff4a843
zf998d1332b57c99183d4496bbd11e6c506f6ab2c670fd72e14210ec077f183e2e21fa0d91c7101
z5b287c3b573ca6db8a15b983a5fdda4c322329b580b3a75157b825c5662169e7ce130f9df83560
zfd44498c37f4fdcc54214589812efabf11cf8e23657d7c5517f2009e558597d2c4489aa0bbcf3b
z76c33c6d652c539f72f6bce84732b0fbc00b363bae9399df6f45be7c66b1bcd239e4b006461bb6
z3296a609738a8f43c207857465923fa1bf9a354163da530519165b33b8756e2270002ec1e1a034
zd80fba4868b5684dab1c11a8bd27a074139a7ed61b464ba4f936899a9d868fbea5c5e26f0d16b6
zdb0a6e10b2e0dadb820d9492d6f24cb21ab8dfcffce676431450e5e108b417a383d1eac6389449
z3a0fa588b537a46287123a57d50dca505c199ced38dac51ccfa3d8af0b33fcef4f5af5653a9c2d
z95f058f2445342191be2f92688ca6ce16429259cbca01965694869dfada5dc53ec03a9f8234d1e
ze7475e91d9a9a4e8216e5afb239513e1336d52fc42bcc4227989e38c4b09282ee213b169330473
zcc60855e818c0c1371eb792a3a4ff4e26f6062d15ea61885231e728b2496c64e0486fb999fda75
z9ca86570d17360fa72ef11f44db07345f2f1b680c1ece0c09a8fc1a14a65d8549ff8099735b21a
z179494280234fda51e1b8e43fd2742156118382ebf3fcd97973fffef4bd1e567f35a48bc4c9eed
z0df7e79ff3c420c7edf173d45b0c665ad0673740a9b2acf7aba5173ee701d4a61bb3e1d62ec6a9
z6cbbc14bce4e451e851171b9622a181d7cab5a25f57730fc532045e8d0c240120e811c143f9a09
z6af06160001d9d27004af317dd23debfdd09c527d8cedb633fb79b7accbd5b364687792cedb6c9
za71ed3f5aef6a8f58ec603dc8241e45846c44df215402f6239cadabc5b7d75eba11a0ea8f691a4
z8356748a98534a97e2ba7b35152db475c5f3691c143cd80b8b458ea0298dd0f4cc8e84ccfe6716
z00ce86fb26dee2569f20004f18fb6e6ad2f6027222e57f77d5f304284b6aa9dfabb8f088164110
z8136f13c967217ddfd1e333b71e74473578519603c27ee904520881b9d90d2b45ba4ff5a53a540
z170c46bcbb115a06234181931ad9a096156767af53f68928b02bfdb4815f10094387b6cf87aaff
z9554dd48a7769e2b552ea99d002924609d57c6b4412f1460b787ded9aee9557e9d1bcd9a1dca5c
zf8e919a03b2f02efa863924521a6d3c66f00dd306b28478cc78a1f7cb855e8f35f2ccb4af57483
z11e5b6c2e5d83477b04c0f860a6c468efedbbb39ae1a9456b76350faefa07dfb21150bfd764d01
z8cc6c22765107fd16ad1bab863a914e6af8821f97a56f7cf14421ed7369d8bbde7b4cddc11d515
z28e60b9de4cabc67a9b8df8641e0f84a87dd831525ea04153a0bb9ec759ec78f6d8e22a5b2976c
zee9d6d8ee0f6e3efb09233c5b7448c2553a93a341ecb3c2e0e467b9fb60e1b4ea188c806b5fe99
z11f07bc52db4e263397cdb788d1a0eb3a2927f919f5a19d9f51f9c0e94397931cf5a80c41aea55
z406277b315f4996d9c16a950134a72d05e3d472156ef6e6693fe6d21df808704e79dd7d60e81b3
zc47744430dde992c9a3ef8f6422dcf8102a54ec1ebcf15c4d236227d1432d58943dc167abd3428
z7460f3cc825b2fa62df7c3c5e8437a37baefbe36cccec6bc16cc015a8dcd902ff24fc39afda3e4
z2bb6011e7465651fdf503fd6caf3a681647f42b06471b841bddf626b1fec3dff1a24394e15615b
zb22a0dcfc3afab5a05f239b3854d6d4c627f9dead41f37aa7e2e0f416991a0961deeea38c2b3bc
zfb72ce5278f64019229e98aaa3f0183037e40ed1dbb5f74537521c57aaf2c0ffc663e3f630cb65
z8809d669062cd04613fff09eb3883b5e881503c5dd0cc98aa501720070710b276291ddc9f4b272
z18fd7934f4ae0b7764c51d2fa986b4a223d616721c3658884b757ac345f2fda9072332cc7c5b61
z86f497d6a9bbe99742ff9f288e909f321e85e92f61a4626424e903d8475d32cf68694dba7b9f47
z9b639db1a1ea640b3ed80dd1e0bc1fd1e0684433d997e58b5307fb68d8abec42bce06524da9ae1
zfe87b8222ee71d9569a7fbaebeeeef5911f9a011c40ad5bf5d5514e30ef7a07ba75641a1abd78f
zc4fdfd720f5c8b0f32cef5682ef5c9576b727cac7ddc4aa2e50114dd98efaa0a0ca0a3a6a5de10
ze20ced1b368393d0619c106b347f0b8c40b1dea45a52ae4e5e87745788343abe9e109347494099
z8063d552142f371c407075619fd9ca30d177d4d9177ed2189d9144c49fd61dfc7d9d60d3bfb6a4
zd02e62865716fd555205d0c786da68e58f9ec59f2d05a1ccd4aec9b50bb94f2d690d09edcb38ab
zea33c2a17667a00d6cd00ebdbce60606e89f2c3257aa49ab7baa7d529129cc04c6e67fc727fb06
z109d3aa94efbce9f46bcf62858208aac6103fd8fd836e664bc1e7323593759e32bbc56f7800fec
z62417b58c5cfc5441f3ae39aec3d1d2c099c868bcddee37135eaad0f9e4e3c637049fb1187b490
zbba3180f1bbae3a8fca5f504b4cc75329d2da96d5b22c203804b7ce52413cb60d897bcb5fb30fa
zbe15853ead83a166485f367dafbfcb88682b2ba68e5e56d1a0a932ae1e41eab946338d954e4a01
z095776cb7c649af43be001e1090be2eb4542de2e3ce324448e9c6f0ffcca42d2d879dc3356d020
z7d8430c9c42c98a96008b072d869d9233969740cb03b39ff4b4e8fc7d4ff0327b7640217c53e14
z2fcbb0a22c304106c063ce6e5de313e4987bbdd7384bb7252cd2525abf43226ee7c4d6a16ecbf3
z359fe30aa5c4d56590ddb01c4ff1f62b3cb0809a9617ba6a69015170c0b3b30aad3e019efc5b5f
z677a4f0d7b859505bd5db5bd6774c82a4ec616ed19f00b1ba9aba3beaf25e8747cca16936b0327
zd3734b62ee115cf1385f7e8a313fe72cf6018981690fff215e3e15ff4d8435c481d62642e31c60
z5c3d875537046a8a830d6a0f7a97a365983f45a8cde029648ae24ea89e12a59de163b86f636168
zf3e7622d25a25b3d5c126fbcf310ce44b0df6e1be30fa471eb457e1a58145d28d313b331a0193f
zc3d1ca9af1488275c781eb6abb709cb34d7219aed24caad5b06ef2959492b9aefb0509da6634cd
zb7bab852fcdf7a78dfaa8500bcc8f4b2a2b9a83028a3d40c330ee6cf8fe4ea96e690088e7e055a
zba5a0b3701755a8ae73deb67391e0d6e963a3ca49c60c107a9a7357336032ba69f19be1ffd4ffe
zc5560a79b78e783a7b9082d75034cc3362750b6751f1c12e52c8acf656685cff93645b2131aac3
z5ed48b539637601d4801462bac535b74ac21354d8bd2641e43dd646a76bd1674b2d62690ff87ed
zc3b1221fcf80366c631170757547f991b71c1ad0e9e5d1592b077bccd6dc904058fdfc771741df
zf70ad7931f87e2c47cac23ae7c70106aaba46d6c39d13385e96b71657618c05694d3b5f3b04df3
za832147731857fd2045f53db6e9cba0491ad897a4c0879ec2db2c41e346d6618e9da182f0e3c7b
z965f0fd47eb3660eea3ac9a757a6e1ef61b6198a3839b1883c27af0500c11d3ddad9b1b15960e9
z421b6b81fce77f5b48f9a91fd05660fb16de40cf4e91a824035b0848cddaf62eae7f395d150c81
ze2bfeb859090eeb1ddb61656c21e86a1b3738eaa0f44c4c89dd58dd75af58362791533bdb6d0e0
z6e5526760ab21857688305179af89bb1a9409355baddf979c74e7d22804da2925c2a8a96e06d18
z183eaa839fce1fb50c86c9b7fa5798cdfd0c94cdc45696ef4331a9c4abe86bb03db654dcaaab96
z2b88f7719ec38a646199437058fb31c60b5793e338ca670fdcbe4b5cb19e90c4540fd2a1ff8b53
zc6e92314de4d5c2bab68629f637170552616b7d3211f3bdcaf9f065358d4bb3162f31b09a43aab
z3afbad57f3394d264f53e95d73fd52616c0c1ec1cf57089e4a2d83f0af65ffaa2945c6c49898b0
zfde370a53e3695a2242ae572d932792d4f53897c41b4b53835831da00a66faa793ae8941bfabd7
zd3014d27d9e5211ba1420567ea73769d4ca688adf590531afa8f2cc885dc72a85ae8c02dcf594c
z8128b465968beb18ac6ffc8748cf8b6b5a29840f8553b72d5148b44db6a4d35aeca5ab00f25d38
ze5cfbd81b888e43a001b337d781d7c79b3145ee89cbca46ef7c9a10e1377e08e591b36d40e19fe
ze1aff7785cb868e27082ac77ae334055cd2ed3020dcd09d363cf4abd5375c96330428fd40af853
zb7c5dcf311ca20b84e694099bf951c72405175cf498537ed86dcab1e1409b0046335ef2f54742e
z0e9a9f20b6e7e0d57daec55c1824f8ffac0cf12bf2490fadaabe48f88d21fd53287cf530ace66e
z3278e246dba608ad42bcd183f088947dde7f1b43cf2cbba511ee8927589428dce548bfa2d12976
z52dd5a8693f83ed1abd07be3468e3bbf08966ce82046231b613cd94d372c551d82f60461826bf0
ze4ccb37bc64d3fa5563484a46ba7cc75023e3adf98e766eadd84b1c1c056fd1ed513206d82d502
zd6a2b97e441ddd1d860f1da6808b3805db8777a170077a8d4e35853e4ea46c1b5b3d97567e8e27
z935bf24ab6e3e3f87a46407943241378dbf0fe17ac14ec71f78c17cbfbfdd59101a9f085511192
z20fd36da5254ad39a85a939cef36b0c3265c09f63661bca71240d30f62e0d2fc5196b1a4f7147f
zb1fefd6b6140b391d34b9374c146fad34b8856e2463c3429b1ef6bcfe0f5d3f9a1a28125e890e5
zc883b529f45a6a28677059a868eb90f1874acdee519a5c393d4ed71c4c433c3a0cc49bca97b91e
zfa73c73dc996255acf7c096a944b5e1030e594524f3b7ccb062461c051de53db21674c1d7c5463
z25b9807bee1c1caf290fe26b266617b9162b80de3665efcc2eba82d42350f0a254e770075cf8a7
z1b97693798f78522e99360d8b4d527c84fe24e61a3e9fc252e4d593f0566385f25cb91e47dcad6
zb12f6b05d8b1647e2c62821ae8649e0ad8e2ab8023a70430b765bb10cb05dc6d772628b67bb383
z060d4bfdf2f8645391e3211b7e73af6e803e98761a56d35050a217beea13bee2f44f47d84e9cea
zf016c3b177b5b2b96ca0f9a3542b15c12851faf2d564450701baf19c7e02ca7e6b43935faff5a6
zd2719318b3331a8ccbfe0b49980006945944f97a9d655275bcffa3a2f3012c097642489661b6e7
z97319fa9a9a74676e33acaa3ed40ada9c852f7f55f6621ba87641285009e1c3833a474c2cbb963
zd4e44d64b9b77f56bb944d5b7609ab13ec02fb2efd6abf083c68260109cacf3c78c3974af70143
z173a4ebd1239503007d513146e96d3168280865b4f133af93a780eb09f18dfebcd05ed33865671
z426005993f0eff8ca810e79d26d1f2ff861d160d33cccf52ae2bf4f9e252a00b76faa06499837a
z766802cbcfa03998fc96dab6e2cc5cd3a6b69d890a3bc4fc3331fd8b2fbccd3dcefb5d49ba6785
zbb1ce23ab50a248a82cf57755f60345e16d24b3e5391b47efd2587687c60877676b74a79fd35c3
z8ae18b8cbd71008ca401d178412c2f885f540b7ff5e957fbadc7bccf586f4bee2b7f811dcdcfb8
zdf474373afb18e9a4a05ed8ea598d94593e4396a3afc930a7652e056b52e5f4e2e40276a7db10f
zc3c7384bf9646bdc27ce53f2f6c4fc6d2063d4d5aa78113366fbcd448ebe53afcc61453d0e53ed
ze4df9be05ba558fe6a22832cb3f9986dddc861c6c3233c6195463ac76fbb65b9af8b4be855a854
z3aad992b4cf5c96143517799fe9e03e10752b06320f340c9cdb0fdc62e070c9323db445f50a9cd
z25e34b632c270ff7fb960f7d14209df449e98f564586e2cebcdf4c7579e9ba3148fc1bc859bc56
z2fb64ed2d8e1de036c8279bd21ff396f5d34890bf0a909c652634a1cf9a72eea7e95f5c6b2a130
za0e6d5e2435da16c346b2fa7b5b814be06c776ce695ab3dcdf413ddacda8134b132749e9a388aa
z57d15e7eaa30a72f470be2def9fe2fe690635b0d4f457593aed54e483aef6666f410c1dcd54215
zb30d2c4041f72068205926e9a52a5081c7d8a8d5ad7269ff81192fc515b97964e250c66840e393
z6258787ea08391b61b4086c5274f0697669411a29329cf660dd3c1b3faeba7d3e2a828137c569d
z44088d327a6f1e8d7323997151781080c36b421b1943fc4d23b5c987287831d4b8ef0d7344f5de
z62ebc63636196b6dabd66f26918aa3ad1519b06e454b2772fd505d60fddae6b5a5a66d8140019a
zed6ea6d8de77bf90f25c726c32ab0b6197652ae1cbcb88f47d99f874f6ec5aec8a4a16c29e3b2b
zbbbe1dd2fd1c84f380f2947484b71df557d14f0e855a8034af527f7f275bb776a26cd74925d525
z34bd9e09659631d9e1d3532d5806204c7c21d6a3eba905122b9ecb652abaa0a7a5abf05aaccbee
z610731da7f059396a349bbbbb57a0da0e2fa0eed32196674da7c0d13245b4c6c76ba15e06df435
z33f776d5ec517b80ddbf5880c7c694d205142db6dfaf126d0811d7f5081469ca316f21f726ee47
z882dc9290b792017808e6587b0c79c950904ca4d43055ebaeb3f4787a04750a3d7c749c160ae06
z931651b5ac6f013f7cf9d98238ebcf603cb4816ba4270898338d8bee75f3586f3a4155df501e57
zd7aa6dac6497558dd64151502e5d84f8ee6f458d70ec1ba1119e6631fe065f10bec5b3613e16e5
z50dc9833a8935593639e27cb62954a2a2ec5ef141ffd541fe3fc6b24d35dd9a51c4ebd2942bed1
zce3f384cd12aa9525c84288d8435ceb6979a7dccab2f64afef3e5d6dc8c8152ab168fefbd8d9f4
z55029d3aeb02f2558120d9cbce768420ed41e878c5046c1c07b18bd95601f95d5568011bfdbee3
z657685b38c55b2618cad5fd6b9da5ea1311fe10dbdf0e141f4fedd41ce5b2ed969f701f80258ae
za7d33297ec2a40c5d7269450affa027636fc44dec88ccb93b0486cda1d727ea33e5c3b22387362
z13418722c099426b7127719c27c2e81523905b4ca386a2e15c3f395e7b991365aa878035d97b2a
z2c1607bb8111df188f9dd2d49d29fa2308018b310133e0bf04f1812c5a4a5fe4077068cbc331f3
zcde7af31a7713b03924e1c0b342d62eb0d9a2f4a11651daa2d1e01c954a6d96335d6cf8f03ba06
ze8558c54bab83bcb97040c5f5002b13482baf7b9007678c7fb6e4afdfc8d3dcb4471e54f67c4fe
z5c88273d37f69db028b36deb84d3f2a1f02b2918f183fe83ee4c27eb6249ccd6bbd5320f4d10ff
zdd376626961db7347e83e0ae621dd26f6ca8b347c2092aa4f50045ee98db5db7efc582f11d4571
za15308913154856edef516820ada4807201d58b110d1f85d91b1268447da54ac740973f7b5178c
z88f5b552715773a61445cc1bdc5c3d0b05bb38edac14180d76e8a8cb7382d2a20da42b2552f846
z4ba9691b85b23ae307aef3c0a5e31e5f49b27e556193e79af2be86fa684ba279c3794de0191033
z35325c804e74237750d5fdd1b03958e83cc4077800020bff65f720f336e326ccd6f5a27b585d63
z6cefeb6f4615e7014c386b89d3e58cb0bbdf6e17451862fe171df3e0c05d0c13823b735ab09408
zbea3e3e63b3c43374787ed6d444f4f2f7b7027581a1502dc3db1aeefc230d493344fb4742a9ecc
z29cbc84278dc846c3363afb7ed0691ea92a79a9931aac900a84a343db4202b724bb763f0530e09
z262c647ec1b1abf1619dc64a1110ec1664bc1a8c984ddc53f008635fc93b8d46e59fd2e177e7ed
z89fdbfbb02685008a8eb80630e82186c4a899ed6cda43da0144959a318e1fec04f20882af3f474
z04ff939f31768654aeeb6c094d644f5c9df28146233bb9d7e8ddb3d4471b2b3f2aa4698b4d599b
zb434f7a483ae4a20fcb80c0a9ac8f9ab9220ad189284f2ef6186c4a80c197868c41b38bcbd2289
z7aee708c1c33e021f18e8f2c35ac7acce4722ee1ea2857bd6de20dcd31a36984812c1f9797d5fe
z13539eb306fb321d4037b51e28a07b8e32b6be529fa440e1106262bdb382e46aca62c17eb6f952
zf02671664da8801d8df6f5778a34d71d2721d6ce9f712b703b0bc741420d7621d022c680df46d1
z1fd89da2ed2df32c3efed06e008583d0ff0f28a6c419604dc0a7bb40998839922b9b57ae3536ee
z66644c352d1027304367eb0acc824a9f67b6a0d0a6b8f732b91c58824039ba271cc04ed38d25ea
zaf5b2ea3d9c1479cbb291fbbfd478b3e14ffa0b4385cbf0df8fc380d1f8a97428efb25e567a81e
z03e91401511ebc2190c4a87c1f0a6cbfe55efdec406fb40ca2ec2abb3928f8400d52bcc38daa9d
zf5da7039612f06006a463da90cb9ed202f76a0595363056b1c814d130b1754d15a544a98bbf36f
zb76420ea1785d27d155bcfaf111ae6b048bb8864ceef9fe2fb01e5f953fa0fc362b6c4c3106c3d
z4a05a845c39c1a7614a61e35145c7e3fda442d078905210c81ec0c78ecf2281da8edbfdcf2a522
z1f5d9b6fd23b2ed618d7f875b17922e3c1f1f24fe90cd1ec67b40d4b2af8277e5936c5ed487aef
z38030c79baac038216e71b107632bb571797ca28a0118c14506bd1d2416f2f40832bf06edd7c65
zb779a0b00a9a5c01cd2bf9bd0847086ccb7e6444c1265f4752e2a9d1bede1958f8865078fe769a
z2dcb5219c158f91d572e22af14c1cf121998ef567fbdad528559d762dab40f7b646c8c9cecea5c
z6d218050db6bb2b410a52ffc391ccb04ad20e4b23f406dd4dbd41f7a1ca085e0d962d853255fd5
zee0d43bb50394f725ad75d1b9ab4caf4f7aaefe2c1a9c28c3cdc47e2ef9ca7d72f42ef2d85beef
z0baf290ea79e04ffef4af233b57f2f709cd782ea8e8b231f2feb9e899e9be0849c7b482a0f0e0f
zeac464881f54f04a054b2f340655bf47628b7fffa85c5da0788efc1c3a8c4987c8aa6b7077fda0
zc9375b512cd997e0f266017af54388c8e23cdef11b302fa93305e175410631aa743c166a3fc5cc
z5b6d6a313d20bc3417576d55ca8174816c726b1d73953e22afbb5f3ebe5c8258851a2f53d57408
z89924b3338546f309a43d2556e3476d0ff3e3153181a2483450cfabb84c6cc41bb0626a99f87e0
zef44c782c5a95bbf890f812081de7e0b34ef8b19de1c87650d41f481fbc5f7662de4d6efc6cb07
z64d1e591da4803d7b62ad95a586e04bbfa3d98be315ba253c9d154516ef5a172c0b9f087f80909
z962e1db3ca88ef00183aaed32435e13dd4f1b74b9737193ceb4da991f1c7fecdec4413fc6989b9
zf50418820122595fad5ef719b52b68a1b5fd142fccdef17cdd22400cf71acf52d4a5934af354f8
z9b7c5e4ac4b2fd33d62f080888a431bcb5c745123f28a99aeb82f1834fdb31f9801d864768a0ca
z321f724f277892e04a66b6c1e9bf848198e0ff269ba4d532bcbb086ae4224163101c562f17c732
z541cd2789c29f033f11773af964081f6b7d47fe7e599cffb6c83e2dbb337ec4a4ad71e2c5d3b40
z42fc9b56314d0cdbae9361ea62d3de675d95d38016d45b1dace16081aa1a4450d387d935c06b39
z31039e6773293934c4b1886e6574ee0bcfcaf2e8a11daa0b9bda147f93c3626cda90d979b6e0cf
z1fc1e0a23c1e55f268095e572da53da910a0769e647f95647551d5d1fdc6648bda8c70b55d53e3
z93bc049e2c0dc59b0b380f18e7d74c39a03550311166c2809cd15236e84ff3b9081364322eb55c
zb6e52eb6e2c136014ff79392586eccd187d5b09bd7f2c399578ea60308cbcdc9e598a678729c79
z6e57dd2b8e51c4d7c8c1be367a33bf7ebb356281825aa34f82061e60ed40011fba74636bc160e3
z6f540de6b6a0cc134e297b16d817c885b3f527442cf912abb2eb1bf4491e99d6f03de4d4aca176
z3e2237307770e4c3b545a9233f7b185da39b2f44f3eab48d0de96d8757d554ee31ed0086b9ba99
z2f219c45186a0eab92693ddd1bbd2e452d33962536bfad38c4f0af110c378c112857e0dc25b97a
zbc17f5b72379ba46e03ce879452a8e3d4b85e91f7d520a1ec74ea2212d26e2c7775e32d86ae65f
z723079abb3d4a82c22634758e62c4e823cc30f436e85f8d80651363f6c7bbc590e4a8c2f9452f4
zd0f3b49ad3519fabaf444cf58792d7df30eeb8810dc54d9723cdde2b4a08fcfee0002971f9a9ff
z68d461abcf1be4cabd593fb2fc426d7818046a999df83aca1ed896591fc5e82fdc88a2f5896bf0
z0799ad573e59843902e346fdee1c190e646e5b5d51cb57ed0d2883984db81f011d5690827f85f3
z2006d89232010869b5cacd2bdb7219b11769d8c376765ea1289b7802623de5ad80112a4e8808ab
zad4049b896f140666df89bd2cecf36b92e81a2d79855f3230af397ca989c63c0c4b112ac580951
z6ceaed508787cca216d3b0f7bde9dba13127c9105c8ec844c9ca901a522f672b4cb0a70c585278
z60d0b0cad8ace775e0c127e98f7b9f7e90e4af0993e4f168a9a3fe6c23dcd03ef3dcb7036b226b
zd27f258cb9d1745be4be12bf93ab0a7b923e2a687f9b97d3cbe4c02066a66554dc94fd09a6c470
zec042a90bce40308568e488a4f642ef4532c24221099249d51be8bb361f7dfc876b31a90f8de8b
z75638f3b8d030606e87c093b21eb17de7f3fc94ffa2636458c875d2740876617ea22078ce27686
z1a4e7e2a5c7a3827331ddeb1276d0105ce985ee932ff5a336e7de242404782ccbdf73e087e95c2
z01a09c9657771a9dbdc6a0a7333e3f11bcfd926f53e9fd60faade17752941175b790a9b4d82aa6
z394bc7a1eecca68cf9b8cbc580dfacedc556490458c8dbcff07e00684bb6232a9c075a6195e29e
z02370361528dd92a2958225d1f4e6aa3f68432eec1b19ae66e110a96949cf36ee8fcf973475681
z9cae42a5c9028093d243da2f70bf6821d4ba7c5052f1ab2b978c64f7ff01894c87704420aa48b5
zd4b7e674270f0bd20009788d13a525ff1fab2b659cf85541e49ddb89511161f31dff7465a35d0b
zaf004b43baf7b48ef59cace1ab5351ef2d0709ab3fc07bb45fe70e476368e7e5eb1184e35ba374
zd23d20ebf9ac8483b156a701b3f2905349aa5a56dd8a54038bcc62b48aff73a316164df7bf2c42
zef6705cfc4876785d7125374e04cb8b2e06c1c1007d26ab7be2a59ca25f036ef2eec26c6459b4b
zbcd93a51aa89ce1a6822223f17a251a6d56992cb15a2777e024f660279e843e4ab8ebd0db80094
zffbad279832d150a211f4855b0423497a6ba3d870d9f463135a03cbd7f47ee165f90301e3d788f
zb0a47c4a5516ce8d6f9347490a8f6d16912ef3ab39b0932e2264c5575ce8c1006d31ae92d09de7
z5dad844174cb308a42fe3d5a05bdeefadd9b5daddb4503e63ddccb2a650eb8bb7478384e4689af
z7750f6277322d5daba354cef87e9284dc16d5cdd68b2587dcd189654d7d671c36fabf409566651
zfc515a8cca9b881ab3ceee60c967a566f3fb2f1389fd31215074498058e34baded37fb78fe0aed
zda8bb84f5ba41ddd8191513a47554866ba119572a794d91bf0fc2adf86d5c143aadfc423332305
zdb9768270bace08efa3ec182940494a5d77c71a93660b83181c5818d859c3a10217d7bec63a50c
z4cdd0f43e2da22be98cc24121ba0d124d3116e6299be2894d2e269f42769679b977513592e8bba
z0e9fd61f25f5869ee83ad742833f666b9871485b2cd471cfd7371d92a6345ae16a5e5db0f495ec
z685a1884641d743a367fcf4452fc972355af79fd4cf24629fb060ab818b155df268500cd2a3b65
zb85ce125e99d25ba36f79c015377a93fc1bbaa2fe163fae8fe7dcdde7afa198d32659a5bef17e7
zb167f5e3219c132ce8cc1d1cbc451d6de6c66ff5622d015d5506bd5c6519c058bc2b6e3d173d01
z7f4507bc3a7db2928cb8342dd14f4e5f217853ccb6dfe58004afdd0fd5ffc38571bb18060094ec
z162c60f49c0cf3dcbb71a1c4bdd834feef709bd3624c32202cd0f15dc103f185609b735cdbab44
z6e83e606f2bd78e5baa3dcb40b6e248009818225f599f6e99afed9ad82e09e0f6ab77c2830cb14
z020047d469a88fad814447c7ccccc7413f5c7ec7974abfa7511b22b5f1280a2df68b060e4d97f2
z4a51f12a7c91daae76aaeac5567daa17aec3953920daaa8cd0fc359161ac550335f3ce7bb136f7
zb7208a7e9746223ea9b276772845ac55ba33eb3ad97de85d37715b6996712f74145d34f860e5a3
zad8ee6be391d6fc756f08a3cdaef90f28532d0bfdd037046f99762f8b1790c12292814dcea176c
z1cde8b7a76c643dc1b34654d3a23d6550181dc3a76e83b89b38947802e18aa91e9b0deceaf9034
zd1aa6571e3d6fae849e8303b158c2ec076e6f4546290c7a185f477c309b240868fe601090e339a
z27040e9586da83d0121d5a987bb082e10e3e2d153efc4fdd2351c2c64010cc1854bd8ccc423c25
z8662ed4b9d02934503ff8650621f0e323235311c6ed568546f69db69833d70f19aec128ba995e9
z710deac8b62cb3689cd5ec1a21c039caaba8018a0c29edd51f94ea4e3e080be08a792da5461e4a
z675dfb913f261c2ceea1242b17187f7dafd5101e3e88a254b9f68160d3112bce10e9e2525e7c8b
zc8eb4fcb3e5bf966ed7daa384346439dd1bf49cecc67d9f6112b7400139acd2f15e43eb0bbf09b
z69dee96d781bd1f5cde17ca8192ab7a3297ac200e43e825c4ec81e777040797e40ce3d69069c0d
z8e8556435d1fc23b2e85c7b83b57e85ebad29fbde7dbe624719d90e1dc3dc97d7226ec76af8651
z5d81f0eead433897e602e05b722361d6d6c17ce15c7aa13d7c54e7dd67b76d5bdca62718b21c1c
zf38b6f6e91573d74c0e7cc27d88be7c176051d94003aed769d054689f499d8941ce90a2609de8c
zea1294eb952bbbf8b5928587f8744767fb39f947bb8b8d6c6ec1974d4d38d0e994ae35a45f3165
z29179e106420f0d8306e96d665f59380a8b55f7b68bcdf8cb77fcab881b151d635d1188b1f12ec
z9aaeb2b92c800d3f88a2216f45cdb1e26996446e3fc501489dfa9f4bd124531c5e50c9fbb14fd0
z2a281b45b12ba6d0d23adcd93600af99ee7c3c704fc7664b28cd97b6047c3b9386e81ba86fd969
z99a37317ce400a0e78818d6ee85ab3cb73fff1a630b0286ab778a63d422f70baa7b7cfb22ca73c
z026a4a8486001c7a7292be28f51e92c0e60c6784890b1ca76d4ff9f8c20f9dd76917ee7ad78f62
z8c498c3da35179e24aa626423f4d198bea1b018cc0745c9b3dcab7717e28edd16d2f5b9be24e3b
z4a34554bae95693ee537a99d1e0b45ffe2518772a9a2a8bb020997991f862163f29b89d052190f
zd13534a00f9c842d29ee046d17f4aa91d85a4a66419c8961ee3d79886d79dfed53872bb38941a8
z7fdeaf0c6fc1bdee866021a250fa8df4839e6aa4ef9c9c5774baa501b4e5ba25ad32b50c200307
z0e02f7e771489d89612f660be6938aa836a09feebdd0bacc6158c2a563bbe5c44e595674811115
z2a2bd7bf8f98ec936844af887ba343b994b891a5eb3e108ccc1ec8ed39638f4a8341b255debcab
z04e94aa11705f988f982641b5490de723b59c85a92ab8a5c11617a65df37a1479fafd7f1b5637f
z9a1750ab7c6790ba7089eb0d037e874729e8179eb602cc63bc9aa3f169ea65d0265dd4f43f2f1f
z62a3a26c58366d9ff050182174fe2b4ec5e83c9084b4ecfd0f088f105794dc97190977d4cac912
zfa49503b4cf86dacfaba2331ce20bd4167f8d78e9592bbb3ce803eb8c00f117f464832881fc097
zb1fd87d62659efbc0046a58b36e35740b9e541ab75246c9729e4f06e5bbd1ab436754f3dcc692f
z442ad5afa6ce20b8ca3ff593347232c94bccf92c5bb8e40971ade612bfc83f52e457ef126ae610
ze86e9ce4de66deefeefd323c3790f7da994c3b9fc4c38390b2497acb73bbb7a7b9738e88f7213c
z05e7f7322ebcef177aaff4ecd47b7a7ee8f94c0e6b0ad0c5320ea49175122eb9e70e25861d79d5
zbed5862a32e24e03de3568b2ddf15bd0859c97db5286612750de5a8b6f814fdef935cd1d55b090
zc751bd956ca179acafd1929a8a7091b63e858d33588ab2c6b5521fb71d6a7afba96b006c40f669
z3a1de281b4b03fcb92452f88e0afd20ba88915bfb37a1edf3c8937bafd4750b8efc6824f693059
z288d4f7dfe33b8c4d679d5b6a5c7159eb1be44e858b0415d20a77a1a6baff10ce86eeac893fb5f
z66d3210eb17f646a3bd5e80612d22ed9cfb6bf2b3fba725eca39f4e9ec14336a88d1d8a512985a
zb51d2a87437f46cb15cd2be624bdd760e850ed80ac4ec09508d445e45837d2b12b0902c3e9e336
zc45474ca093d9e70d6cc330fe694a412abef4725f6f8b7fe1e7eaec382d068e740ab15e49dca40
zaca5688a0214fd27b3bb20bb5e4bcd6bee141ac91dd4474908b6a028fabddfc1fdbaf78f9fdb84
z060fa0b68f107095b838a53dbb910182fc42f9b156ccd509ac46d9a0f96dc51b814c499d490951
ze31e05f84584a0ec3b92bab3cd0121d2c7bf6615a299efb2443a931f7b489170937f87358174cd
zd996570bf1bbd0ef462d1f196df62183113b0e241bbe28f56700a731d44184554dc91349572b4f
z03bb54ea57ff290cfedcd9ca50fd9a0e41281866fa630747032fd61912ea2cf34c682c27844a75
z0519db842c26bc5e8d30d66a7b7fa92cdda2c20aa25f11bde04c367fd9a69be948ac4c385b2480
z02f0710013e8967a191833afeff17301f1393811a4a1c0a540cbe7755e5fb5f53408f543cff73a
z195883d8adaad3542f38061727848807428a2c85c47eeb5760190ac8ddadce5a3b7fb7b2e4b58a
z0a54c4f04d7b09d8e6e69b2460d72b72ab27311b2e14ac19e8532c74b8d3761c500521978b5dd2
zfce4da0e2054e9209c0d48aa6d789d431fe3fb8d27bf22731cf87ebbffb349031a95302b24bd8c
za152cad2c6e1197cf6a49c013bbf3a49e250965924e2d319aaaca7ee3e55b44b93d1f483ca8055
ze674113442879413bc56b1413a5cfe3a4d4e96efbf72347e3d3c410f821c57e68af91afabea4b0
z532945b1ce7668e11b364ba7ce97f5fbc863877467a33e8b03596ae3d62706d64e3d969563692d
z95e5cbf94a679cee47347274130f3d62edfe234b5817a378ce62e8b9dadfcfba5b641c48301666
z3bb9d45356744b09a62d569c0c8212d38019737d8b4409735dd4872391894a539155312ca6b7f4
zcb8279286bcd3515e705b85118aebe3cdd289e7ee0536b7b1283e1dd3f14406421c39d52c4d4d2
z92c610335a2e3f191898de0931c02d689c42583e18771f9d9f660a05933d077490162f9645c144
z65a9ee40f6ec277c2b7926e7580c6763b656b5a612f143f88b9e972b7e8a11d1b6ed3e2ba24021
z3653bab7e4a3297005a8141047c5a7c5cefe6c8bf466474223a7ba715128414d709b6d09d9c7cb
zf457ac8ded2678dd4508c49e5eb512c0cd7252ae9f44f9979e9cded864d6f116f9993158a07973
zec0a02c267bf0b8d56f05cb9254c0d67a1028afb121590ddb0491587f9ab0f9f063435129f8662
z7545c637ffe5166f53cfc22a637a1596d3f27de7041e3f52c826389c2f032b512a3ab97a6bb7c3
ze864963a9b05d304bdfe424d60726052c73b36addb174d42bb8b41b043e528d750b4872d343601
z0f44a7ed97ba7415cbd0e9e12c83c4983ba72b446a418207a91f9abacee52ab86d95562bcfe7e4
z37b8e6cf18dbf8f376c0ed3955fbbc6ea8a4294e95bb50dc8f2647d08afc4fb32087b80f0804f5
zce4de7860b6afb22d49b404aa9b0e87a7acda5e23fc5a06b467c882e261dcb79f6d967447a75f3
z6b9bd5d449bc40fdfe28301adccdb37d49ae145ceef6733e3727ad8ea4016855ddd75dce491e03
z80603f147874c9d26986951679450a885df44c8e092bb83b0db9a3e5302f02f0d031380f66358a
z4c95a93a40c97ae3528159dd8ef8486dce97dc6d841235ea2022583728be441dd6fb77d90481d3
z3a9ce3c1b102f84eb7ab82c6eaaaabcf76d9c1f87cbc04d5d837172cbc8245af407e328a24f27d
zc51efdacbee7c1e0dd0d50b354f0a19e2e2b416db41a00fa8e53db675c5ac269b86afcbb0eb659
z1fdbda6345fdd53c3637514f744057d4486a06c73e8e93f52fc5d9f8ff73b7efa072ed6c6951f3
z356b71071b4a7abd1a08bdc6763d034de8a2b06f3c12c8296082600dad58cb8294a2a3f5f02427
zfe9462374b2748f196f1d7c3438ff55a9c49a8c54742d786b29059a974f01be41ff958f6b1f6cb
z3807509100728a1966962ee73806c83488b923bb4754528974c8e754e6e67e952ae9c61976b973
zcea779471360054ddbc8df43ecb4d9f5d467fd76bbc24f09c0175e02e93ecb2fd7d9031f1295c2
z8e452ebd22dd633a63e3e78ed67d98073e2dbae3fcac8959a88db1c297441a0d6ba068eda3438b
z0c09e67627e47405e052ecf01018f371d56d21e0c1be07d6943781a589ad740e0fd9882da1c66c
z529ee7ea25032f38c9fa06c86e389d463b8dcf500924881d94047b22b71a97acbccbab4975c27f
zd2afffa7bebb2da05ec59274fb97ee4a1d75fc67208d5f2cfddfa7ae086ed4f23c6a4d3203361f
z3918acfe53d59e75bc392d0d32b78971d201fccbb8fb5b967af89e649e971caa6cc6477dd3dccb
zae4d8217108a33992db59ed82f3d1ff52b03dbdd5ae1758f220637e31c7794fad20e8d6d998a83
zecd74c54566fc2f5f5337a981c18713d014686a73a2d2322f3d3fca8096bff9e686e9106c8934c
z1fe38be0878fe3e96ddbb14287d4d745693f48f903827f598db38b537c4bb2f7851404d6e387f4
zc18c89890f5ed9c990b195fdefb8f8b26f689da4a1f6266522d0c23fefaa364196ef4990381db5
z1da641d92d9b3e64d88fc480129d4421255676b174160b9d231444d2fb67d6dbb0cdf15bd63af9
z66e532ec3375e4649ddbc0bb302c65e5421a8d9d98e058fd5a5b639897d42089baec16cd19323a
z3dab9caf8770ce28593fc681d519d850b9c3f08a6250a678ae3c1c62a3e694cacd9c51801e60f7
z35750b683d9b2cbfa63619d2a24295e93b28573d545023fceda4371eb174a7623bcb2f5b903154
z01f620fc4dbd4641cd5a75e6b139c5dc9dcbd0da9fa2e04bc0e9a8cb630310a00335fc1b125a8f
z0462701d10cb1c777b6c110774215da322d45ebe4ed8385fddf0a3c5b22eb133006d01155072db
z872c45f1c246b9969d86fa8a0a3bf2cfb8a2ebc2094e08edf92ff7c11f0652eb36b931def6fe5e
zbf9ad672726edf9a71ce98b289ff37039bd62e3aec7f9770ac547a4bd01cfbf6fac79243d9438d
zc11b953df3bf3035374819a81818657d76c894840e7b1f487f0572a581c89551819bd11925a03d
z8798fb95265b82161b9c148ab6c5b09c65a0892489f40de445dd7e8ecf34149ff9c0c1ee17cb43
z585a3033b82932b78aeb739a739709a3bcd48973022a58ae0b150c8b99c0101611c98f0d7b0811
z3b1c60ccec1d8de7f47ed48e7480383105fb79a5cd65afa4ee72b93d32783c037c81936bf333d1
z75144a34c1e64d304c23a197b616bffa7f1dffd751f3d7730104514226a8c98983284794888c2e
zc6f9676fb5d67f53c55ca1956b2da9a4c5e6b8edc992c698142229522fd0d41c00563543f95523
z612ee4ee0d6c33d23da780259f6dfd4ee999a2db62527abdd5aa2db3c8867b7e132a4254cf41b0
z539bcc177fb815b3519b54ace43476537e15abd68b61dcd16b91e26e18ed7a7a8d567e6d8d0fb2
z821f8077a8d885ef8872184eebb212275efcb40fc1771fb28744857e0613c87838ea805e0da35b
z090bc07d156dfc0ce702ad2454e7af1773ce026c4c82cca0abeeca7d1b475a0b1eb90aed0d32e1
z5fbe7c26a28a362d31b479916a0d147915223efabd4e86381f9f1eb8ecf26989128815f7601fe8
z2d0458f7fb35131feecf5eb5b02ab19b531ad2b47b4eb14d4dddfcbe8855a04c94a5712a91ab1c
z9faca3bb7589c253d22f42695267a77197a5b9fc38d9057fafa137881ba59501e51a9a1e891e4f
zb8aaef9d7463d1600a2f17609b7b74c0e79697a7ba080684e2e467cc402df1d08db1b07baa5787
z2a9ab1561b64305608e0efb65779daa96482e5572b6ce368b415d463aef0700c5e259cdafe298c
zc3edd1bdfebef808a1660e8766f61288e0241c1dbc9f017d8ef564624dfcbb92ea231193532a8f
zc3281f3590e1f50640ecc54b5be229e66f1b125b5c24564210a8f4feb49709a0ec473333fb88ea
z565715c516b7a8cb1ab13360abca9f3d7d4061466e0ca189f143c19cac585e08357c066cd73fd5
z9a618fd2c0477cd10b556d3ad6961a5df6c22430bbd38b31c915dc3aa8384bc36bc55eff5aae23
z03c66b082d07919fed17ca8d55256bb4f000e2e05b7fd3f27d9121981f9f926f3efe13287a1c0a
z1694e86588cee44c11f9189525d07d24d64eafe9d659ed605e068db7f668daa76ae69eebf7445d
z08382ea633816f754856eb3ba147cbcebda8eae25819d38a595a15902677dda4f91d09a4891884
z66511d30c498d8af4b9f4a352a412513e2ea9e6fe3af71fd061e3da19744e75c516bd540e8eb0a
zb71ca1ceb5bccd5d778b61014550f70e1b594bd1cbfde409a4ca81586d024f082a63a88412a07b
z3706f0282d9d4d2c6c130a9834e6641177635132bd550628db711b1f4b91b1efc26d21f0118f89
z7815a1c9b631da8f0ff4e17d16ae0d6bfff209ee485b7f0c915779cc7c7bf1d823e39dbc053080
z18baf000722ceb8c73d3e930013fd3bea0c05ef1d79d3199ced923da4f8d4de47c0da1c7bd090a
z63d4dff13b64162f61dc6c0ecc6f5abd42129ff66ccb0400f9174bfc5f397a5b7700981786dc7c
zfa722501c0c9b908ef56ebc9bf4216faafdb178ffb138f46523c21a1523ed82331b3bf0535fc92
z9583d46e05eb356750611686cad8e15c5a509399914ad22a82ff6f5994a07a7ee207d81f0f9bef
z9d23c00cc44594f199e532c488a2f7e35993afb46ea6b72164bb83533e13a8678dcb051cb0a2ec
z48cf8ba110b40357907a17fde143a2aa80d2bcff4a29e66026ade345a04a591b6ff1f9a5c2a911
z142420cb8954cc02bef3d56e2d576da7ca99a2ee346778a66d766d882e96f907cbc1207dd39750
z50085a00d83108a42008e250a0fd02ef1269347171968793445045c98ebee2e9b03d5e016479b0
z2d1241ffec4c1647e2f286be65474fd68154d2215dc11fcc72ec7abc3d1ce4422264931f7bc915
zb1c4c82da4043306f117cb9a986109ba35d0b9de3331707e1b46353875846fa46a98afefe92b40
zae3ff06f27cd7a91d6cf10989abe79f7472fa4f0ec9fd8a3bc1645ba7a7c856d454b05e33a5d02
zbb16d3937a1f34bec34ac01e76ad6eae921ae6225cc051b8d274718b3846f51b0f97041535041d
z6433d8bf3aa8a3153870a81e107380e0295770c6e19d8f18406a0944e2c910d6a2604b8d2c5a11
zddec385d43a0dd898fa4d80c79d9555065303f7015bc4bcb600e24718e6db4214d1d32da5fa6f5
z80bc3c08e32132f3b6fda10aefa25361f09659cc165416415e9babdb4c3d7400e22a9e6304f6a0
z1dd0e4b392349bc1f88f1715b32b2b5821cc848871004efa2cbdc85644c25e89870cbbf1aebe5a
zf22b142db5960225497f2946085cd4949577c987b3c2e498e840ed3cca590063b381a7425617ba
zec29e5222ffab0e498fda5c578b32db26ff856995aeb1a70267a7d3e921fa8b1f9f89acae4d34d
z117b89a438e2feb1fc0dcf4ffa1f4537a53c81a282b104896c4dde445ea44221cae8b75f622f90
z0c873dbad87d26b2d4583485a157b021f7b029d1c4c0936d62a3ea123732e41c9c70909c0f7ae0
z81a75d9d52d10bc35fabfcf8d98a87742805981811dbc36e793fd67bf53e18e318e7e5942e3a74
z0c532d72ed0cf6530b402252d92937dcd5dafdc61140ae04c877ae4462457c6ccbf739e46b6c24
z6eb3a29e66bac6a4fe0f257af622bfe882b1f4b84e4ea27f022f4283c43fcc094cb5eab4399a30
z252bbe13cf57766f01cec95a4851c7d23bd0a4c8076c61f4f3642fff900e16aba605f82c877423
zdf047a086850f5756edb3d6c8edc2b066f3a66a6c5a6f5867abef69241f2cc8002460ecf5ca72c
z9c390ae673fe9250ec7aaac996a21d125a92538094bc26caf51afe1f70f0c2cb8e4a92ba17a407
z3729f4fd974ea22947f1ad6f9ea3ea89d3a20b1fd53a4d7e4468bea8ead4b18f832b9e8453ddcb
z54e33a23398397e43a346f51a358d6809212886ef246af2c0be1235648908688e6a937d0d049b2
z547cfd72f1180efc90ba7121ec896cc24c96838c9ebddae2eb9d45b5884b51c356a4f495fda3a3
z2de5b7c2e40dbaa3a8daa28d6b430b41a161fb7aa50a57c5c56159fa52a654a00fd67e26e0568e
z2744d3c391a7c30361ec2fbd4cdfefd4d90f5f22341e6372e1bf912dd3035b61b56555288ff507
zd9c1b68db4aef8c203eb49e2cc7d91c5b571138301edaa8573be02c9decda503d5ee0a4657c796
zc0dbbcfc37d055a1c097476963e64a31daf32ea95e2aefc998a7af33b2f24413437c5415fe966a
z98889aedc03e254d150fd9a91dec412c32b194d753beec51cf8f796f2b821e281c540950e49e48
z0abd61ebd706a164ec7797bb6296f05cc465c0e15e7f4c472f3afbdad420483c00ed260123bcc0
z617b27c804a5757199c6aa4524fdf978eb710936c641e2c95d5ba5056f16f04cd5a1eeaa3c0fef
z3e7282016258329c53440b3e82bc231a48fcd6e5f9e00ce79f25e9139c5242466d573ecc77cd02
z464f1a29c8475f971fc36acbb84234042db49d9924f3acd779898464d635dbd8737fe8f90df1fb
zb9c59c94917e861ba4e940f2ccf13ea5ab580910dc6028130f669e4cba2c5c3bdc2ddb1f3f9d6c
zaf9ca09b79c801ad688f8145c46b20cda3c9f8c95abaaedaf7435287c442a944c0e2fb9da50b5c
zd04d518ec25bbce668ea5cf2fcb3f4541875b6284cbc4ff0a20697067be681ca4072d54e3c0bc8
z266d25388fcb7ac43ff88719d09c42d53340f62441bcd47d89aad3a9cc19fff5cbcd3fa9392acb
zffeeae9ea498e34828e419f4cd0bf5a5746a17f0467b3f00269fbaf196ee3606139e07e962701d
zc017a6978a67f69074bfbe4cd7df8529d6ac41ea667a37367dc3ca32e1c575d923a410f3a814fa
z111f107eb0bd6aee7b64d1d4e92fdeb36011a70b67278e509bdc510a5048b9c748317bed52cfc4
z7fb5a1f954b27985c0667b8ab8fe28fc2a0946a9113bd5b7da2567d55ba9e9eaff47d0e0520ef7
zc713af05a590956e8a525aebfe01fd696f7d5d9ff819fef0ce8949be299ede9e3706a2be49e28e
z5a1eb68638dcd97e5e20b46c3530ffcfb0f60ba723e77b8190d68573d5a16af844cc1715c2ac71
z18f32602ae335391bad3a803327061c9fb8f70aec091ff3f4e6c091ab827d50b6e21a46a7fc5de
z777375bbd51fffec3260463eaab0b10a29258d812ffad447e0d68988162ea0d99d69ba3de7728c
z07ffb01cc7b93e76ec94e50f7c77b077bfd9e082c33a9c9cf0e9e3eb63c06b9e56f7410ddac0ab
z181679b2f9cb46b7710fa0066ba1d2b5efba8e334843e40c41c2dd29c0a49a86051230dc691cec
z1690642bcf718e96356726fa9b429674e7cf2ded8f8a142cceff70f359cb13ed4b65693bb6cede
z4d9703f878979ffd45d12202cb8cdceeecbfa7dfd05667376844f4c5b6434b11da18343f751156
z2d1cb5c5709b33f9d9805396cc417bba468500537e51dcda9edac1d0dff5fd281fc9d62760eea1
zc29bc2596c3251137949181a4e33d22c6b7f93e19439f467465b34d9cd5cf1e45512dafb49b31b
z23b5e5231dff1ae015cd26d3aee476d24c991af30ac227fd63968d3b7523eebca63d53644fe607
zd2aabab0c7fd934e3bfde0644a62a4a18c622916dffc17b2dd8e4b8b177c5623072b62db729c1b
z33a7020749a254a5c43eea2999e99bac3724d651078fcfa745a4abadf03acdd26769d9d1944168
z29ec8247468f6dc3ca8fa822f93805396ab1be177e14a03750e71dc24a5e50b5bc9ac0c2745c15
zdd3cb7992013c75db72f71494c5b89f31eaa6c0d240d9b9b772607ff64cc6b4346ee6f3ffe8953
z36e77de7656046d607d34e672d4b4c413adefe46cd3e04fd1fb84755f606828ad465833c40e023
z07d91ee2fe9af52b3d7a135db7c84dce24504c417fe7ede033d5ea60463001f4dbbbff7b63fefb
ze5c81aa2350e932bed4a4b02a3ad20273189ebfdedb32ff98890b8205e976d35d9f26e029f2910
z32c9ba0a8eb5f1a6bf35f8ea818970c1ef43c8f035ddc09494033715db9a9d5596a17af1485c84
zd41e732dcf3c9d21ea7b89a01404098827bc25e75f76775fac6ae5b1fb66ba80299efc1a8b8a63
ze99550e6dd54f2d8a8730c135273c22b848700c339bdef178403e0bd84e36e057e1d8157e382a1
z40671d64b27996dcea041bf803add67b78b71018691299a68732baf6905201077f416db077a7d7
z7ca6fe130ee728ea8510819956804936cf801b638afbdb48ae50616a64391b917956296b127bb7
zfe4f6e5fbcc2d6df1757f8eb8136d6e3eda13655d2b0209a5f745c2c6d10965f04ea6397cb86fe
z3c18d70f0091c03df0c98509876c27f8992328d7caf55ef7be0ffa40b49775fa6ea2ec015eca2a
z7b6c030050ee1652767c63d8671d37cdafb3072a60f6ad00d2188c1e067b7862ffae44f1920422
z60b788d0af136627404979c01b7007bd67658acd37ecd6ecf2ba96b071d12a9237b7eb2769202c
z76421a4d15f93e17233fb8a6f1d475d39a676b172c11560beb441dfa62ec1e9c38cbc92578decb
zb0b58e67945005790895032cddc52c45f3b3af9a615333ca0ec80bf6ebfde895de783b3d386aeb
z9c9a2083bec04ddf3f250dd8810c7f30dc909ab48027100d2415fc34376ea2f2005f3cfcaa222c
z07bd874351a881dde68450cad0853a248114cfdf13b4940c2bbbd0692274ebaa6a6d9e82c4817a
z6a7fa561c6ca8d707773e89d844eb910d44a3dc14763de7e074034eae718eae9e1e52fe4d9705d
zcf4f14bb384fc9e9e696466481393b0b9457f082be1452eb81b88acb9a405bc4c6fab86e5c7325
za9a6553fbc57019bb3198c2cd6f002553279610383462fb7eb13787bf8118242662341cdd38a2d
z721830206dfeb4cea6ab0650eec6d74b983a0e5bc062260b0e7564fe77860a82cb514cbab4523e
ze83f85b967f33906bef53fc72351027894dcb00e79f2537423665dca5dab5bf2c2e292344525df
zc4871c3d9f0e3b622dfa4d680b54a4f8661445eebb6550a23cd5c6cb484257da771e534a00f0f9
zebaff0a12600087dca9057811861e6e24805b9f8874b174a1dca4a0ec1b951edc48a5d796c1eb8
zbaac7ac5d843b7b62b37e7bd16c6f37039e122ce600dfc655ff212ac4ec3a841bb45898c22ac8d
z3bd31c25fbbbd6798e2aa6cf6fbd8695f759c7baaaf9b7183778469745fa8a00f517c987151da3
z65266c91c51160b077bf5ea539d7cafbe26843a262bb0ee00d8d270f5e16f88a69a5dc52623e55
zec00d89ed2a00f781a5ff8ebe3a65f26d18e4a87b1130d9766ec1b699413901f2884b4bf36523f
z80533b57960ec4906735e04fcdfa93951f6aa0ff731b6f40fd4c6512164ce9268486054a3d957b
z0840540d54ba6286e183acead793f175ddff41b9e59ab1a8b1fbe3fa0c81c2a2e3254dda219cf4
zd30eaf1b3bff5e2190559aab3ef267cbc883e7391d255a3ac7d4b1b307a947e5805005f9d5c3b6
z6270601b1ce040ffa02a0fffbe0915d87eb7fdd9830e6dade3d0129aa1ae9da57f0603d1486612
z9be54347d0ce142b61e397226bf2f7a924c7eb67ad71cb23c5eabc5b8c210a866b711eca05aff6
z6343c50c9fd0f8fa195c67a0d6591bf249bb76f56c55bd0e0440491d9359cbcd404309e7019008
z46576daed8b7c808805dc0865cf3327ca4992739e50d31c05426e90a9d9afb16c85b64dfe5e350
zd5f53cfb199db065eac82b2f29710e0630a6ffffa4c7233769668adb7cd1a9ad8a4f56f7b1d3ea
z67b73e25922b5903765f988fe65d1b9cfa6d8cf60a026fbe3ed77e05d4ce55a9851e454c81b5e6
z96229b030f3147ae719bd23b425a455f80643bfb02a2e7315e697137263942977420d6b33987dc
zf6780db050111b8e1d2238f4ac91216204da4f5c48181b907d186de66c7a44d0ea98b948ec2620
za4d759b0a4e01614bdf5b31ba7dea41a650e433301ba36b0f82870b71dd5036f87f0e05fef1e50
z098073a4e55288b3e872380d3e2aabc44d9b83fc0342fe4487028953d1936b094dd2aeb93f7897
z71dea4f48f088be53a09c1b868b3e5331367062610d0a8b3e8c14b00f62a70912609db63374521
z75bcef1b02372d4f8182497f767b17b852aa42018755d27eeb7feb3faccdf8abec5bfbbd1f30c9
z1efcc5eca3ba43fa93539166a01118fc9bf8197a0ef5ec07fa9e6379bd9ea395e6e7f3ab07f8e4
z82b39ced70d67a958f0eea091a83bfaf5c5ff6d995532fbd1988b55c6a576724b7e0d7366d8b14
z9858d30857e4d39a0f66428068e8061d83b61b078aac0199142e7457323ef399db72f042d5dbda
z3928c374ddf00da71eff871215cde31fbf87ae2daa27a5e8efcddd6261f393c907f18a35fef866
zf13b23670a6c5581046ba82046b0808c195955056f209dc7c42bdfaf0003ca1d729da3650b374e
zf0605a7f88d6cfc314c7caf9a729fece86d3eee927036521fe3416f035d2cbe00f2fc0c937e4e3
z589e0c4cd916fd5ce95e2c0ec06733f1ead2656e9eba84b82e17d3b5b284b3a65e0d4a8c0f32e9
z155fc3fd459766198a3de8a9a514f619664ad30a4f55f0b6d32690ac2b411930b80194ab785ea9
z81ee39e979d624383f9b83ec26b6fed492c3412b57cd5bd0fd3f40646fcab529daecc463473ffb
z24a6aff9efa737a1eee282460894c2c4582c517a97b1c257545e979e6302d6023cd27eca8d1966
zc08b245b167a3ed03f2ed711e9f456bd3444ceb0d084a5a3bd19d2ba80acc446b9bf30fe07febc
zc31c609f883ede5ca13617a3e56dd0bcd454272bf12ae7c648b9baf8e04afb3e7f4f1fb78c9a56
z4012f27a9ac831794f9790c037c5b15991adcd5d6aaaa974ce6d9be3339b27ba55f9a3219930c9
z52c0a3b1afbf02d016e56aa0e91f24e0921271fe6854b11ba0501e6aa0b2af27057c070e2c74de
z47ec98f1ea77c9f4c214e4403247978fe71844e4df858499c0f3852d992f050ed2ed4704e58ab5
ze0291d575da0b92c3d403fefb871cb4320fda15684162b0af5c493182a3a176ac704aa13325687
ze7b6c421c59295a4e56d9c358e55f342357d69eb501d209080b7af5878be6de531c517c237138d
z482c395a98eba6cf387e5f28c20e0011145ad66fd7583352567c454479a927e79edd1dce0e58da
zb166e1bb9c2e3bdc65db7ea594856ee7e20df67e823bded4cfad3e12a923e0dbece13b87c69cab
z0cbc58584f14d0b4c61466ae8970f1b19912a490d0a0dd3a9e5abe3566a055277ffff4fdecc569
za56c18f3d40ed397b45c46d3061f19b5d91af00c231bc346a7aadb87fc6491d8a38ccce8f2ecc1
zddba6e556876a7310902f564aaba0a4080bd44bd4b47b2492a8806db3835e6b5bd73d7e3539bae
za4425fbf8f1dd06e3cbf3a2104791fd5b042fce0cc81c6296a901910f3169ad138b84f0f9fc1c0
z6a04ca2d518a9ba316666750249d4da899408f10bd70e0f2e24634806bf2c3e9c7dd3298bd1995
zae5c63b35280ec07f3e96d4641de683e63ab6b2fac51b60282f500db495b94cd0cc80eace58985
z5dbeb3f8ee1b1fcde6d37a277d21807e8c3ffcc510c18b7b893795523ef8d4d138efe2f13209d7
z219fe44ebdce15240499d15e85b2f8ca1bc1e0f49771e2477fb8f9ceade4c008ec2219a26ffc06
z40f5e087eee68652527045b011212b7515919150012f71233ed57960b46256c69590b8cc260fc1
z64e0b3efe26173e06ccc28361bc29f64a6e4e9370e738fe81c9e31d6f2fbacb33aca120038db66
zcdb5f5169b8056f47a519d7939c3dcc729ffa990b6904c03129a196b3e6befdb1c1aee5061e428
z78c96cee076020740c00536b5a14a542efe429a2f3e1059046a70fd48590829f97ddcd32b19618
z97675370f6ecabf280758214a7c031051a4f4158a183e860031e4cb66afeb53a9d2af4ee915b3d
z0d2f552e7f2bcb93a0ce7869c54bf287a503f1ec61f2bd2eb8b624c7518b83359feff4753e17f2
z3b6674ddb1ef130fc74f3cd4985d00071a5fc93f8e09218c0c9c31fc71239b98cd9c2693d68990
z85d0344980ac30dc724fe29cac8e59fe7ca3cf7566791e9c8ca2e25c0efdd60d4fcc823d649db9
z1e16138fcbb6a799c50a8f92acfb4235654a7c54997c59d2bf92fc23ea831ccc3aaa4d8ba4eba4
zd157d279ce73fd280910fa44b53d4612829ce924c732c43dc777cdad2efb723298af2c0413a573
z58eeb7d54d0c02b2d8ae40c8c8b242a62aeaf52461d6d14d27ee84b690f10b0e3c48503b91443f
zec6e1f0613711520bce7c3d95323bcae6942fb2180c7363c47723f92d06b3da330eab27a748718
z5015c5990f28a6a24b403b4ed018e61736951f44e7dfacb801eecc3d936bb61b0125ddad5faf4b
z86a9b516dd7c262830946f3601120a4419ac91cd8be8ba333fc4f086bdf2c9030b9b61a9a4bc2e
z7328f4633b09e9680f03b196492a9c7f15b58e60c329e6a0e149cd65e8c7b646fef973bd5d0e81
z500ec28580ef614d92ee1e6a7e772ef743931fad895f1f38cdcbdbd3b9becab26e63aa9d33a2bc
z202d4a13290b89c28283a89fa794ed8a79d947fb6b88091abb8adf148b11b2eee500ef6f73db4d
z5b44d57294def745f8412093f97c02c563c1117599b9980ba27d3ce265b475f0a7e5fa64edcf06
z74db5509c454fb506c418aa52b5fba01d23c3dcc4690d7a9e564a4a03ed0e9630c92b2df20007b
z15370bf8dca59727c60b93d4207646e2bf00f444bc4a200095715149ed901a3dec07e5bc723590
z897ab0256e63a3bd5f971b959a4345bcfd270b436f252b1296d179596a4c7656edd6caf89b2f45
z8659aa0a6158ab09a0aa7d82031aaa7e57b0cd639ba0fc978def20e456992d014caac4eb76be83
z52ee4083c5ad4aa265269117843a3cfb5f9b146880f3d97c381967a857288f5f18a8ef70fb1d13
z79f8e9869fb917d5259098e1c9b8d7cdf3bbd281c68dbb0f46cea4e8e4716afc8548397b953721
z8341a0daa042fbc83320a1ce4c6684ee218fe690bb3e89cd371b737dc91271d949b04538e54efe
zf076a7c7be59c4c98e1909f07c0f87dc40d7c7e2ae414d4d11ac3eee36dd5945ea508953064842
ze0c10c7f762eafa1500fe80d38652546ee4319782a0f2802a0e442376c4f41e0b5f7edf0cbc4ff
z5037269f0f58bf43fad093b9fb21cc9fc2d69de830d082e52d4ff52f2a7e5ec2f9fc3c9dd7c30a
z3c8ca5341931fddbfc1ee3ac5812867f9020667f7ea23e2379e45071e43699f3b2f519060b4ca7
z29c9e02a45bea8b0293a25ec5559bc134fd79bf3aa6a0c7bc9323fcfc7386b85a29e8b1f8bfd43
z67e3e1322df33d8bc8ecfb33782f20551d55bf0a7beb208038a0065ec53ef833f6d2a41fb662e1
z6a9e443d9a80ff72c525a5e3dc077e6b1c6b4045feb631975398a80b900a994769fa57b0fe82e6
z637dc42879a15a88d5792597f477b3107fc20590cd854d72dbc393b15667645bdecb3e1ba9b5e0
ze77a3c92a8d9e30777f97c57500c6eef6ad1364a55a0166d89d3274de006e6d0b17e859fb39830
z53602cfbea86ebe20e045e6e7781b834d301681b78e2e01c3d8b8b7b990c7e32153d21ab72733d
z48ca501c5f3ccc90fb6dcaa0e2d5337a80db8d7ec55ec2448f05f61570dfcd561937ea19c58649
z20869f3872dc13aae6bb847d9636ea5b6738e04495b3cda4be39426f91ad8959c800080ae24d51
z73aba03ef06f619d0d95c1e603e524aed8fc86763cadda140d2ee397d50db83f20a93ebecd2d88
z3a323c0916622ad6a87e3924209caeb5832c4416b2d3b5352411d73849f185a2e9802675640dc0
z1fee63010661c7e31bb5a35253cbaf723a321c9b173ac2114312655451f189b0d4b3ae31376f5c
zba1d7fb8c3bc776aec16c37c456c6cd6fba69e04427aa6ec384056f35c40c17642307e3f584caa
z747685e227de23785527b4ab51a631a37aecd9184aa936e44e0693b3b602bc66de2e79f61adf27
z7cc890377babc49f2b47956db58311daa58af2d0323512343a899efa271470bcbd76dcc30baad3
zc93bd02964773c5c2809b19fd938423cea11762f225da9c1e1a7b9f9ca82fcbcd9768b93a22a86
z7c51ac9227923f1dcb1d623e8e5b8a0bde548a37e52ad262a0399404719e37b4b5be61bdda76bd
z1b426e44cc9f1c59d7077038b55c0690d219d2db321b4a884590d80a34fe2ccf77625c2d037ba3
zc0c43c7a04b511ddf74139e683fd9090aade98b42c66755ad0abbe711b99a724c674f14479477a
z1411dfb633c7497e78a07a41626215ed6d2e9f383eecab1f3a8d770446aded913b052e6959e852
z7548c36ddd098b958cec4fd87327ea18374d367e31379e7040e3838ab2381c39ab9d3b4ef72275
z1361e1333aeb38a7821acc1bfbb24de2e7e9a87f39496cc32f898aa9cb9b95c23f7cca6ddef92b
z466dc2c9d969dbaf26a025866c1c08be45c53daff05a851c34e513ead1bdd850b897a3294bd4eb
z0f3b13aebd929b64d4f7a9c13bf1b9c4fcae2a5a9bac052cd4f2bd338d19a5d0c38a8ef727d24c
zabe5edeb359cceecc68618c7a1b0a363b29a10e2dcaef5d74234eb8533b2746988408ed0fd04ce
z2ca9852cdab03959cfe22f97cdc9504e184dfe4d21122ab66e8527ad3d04b1bfbef5363856150e
z8d1f7847e8e14df60800bcc645483235f53e18f0b912afbada4aa4ab70e205a6a7ffe757427a15
ze71aa34a40bacd6a189f6e3edfb6c6a2f881de9cccf252c5fd578e6f937f7643cc96991721aaf2
z80343fe0e2a2ee68048fd9accb4852444f333babe930fe517b751b896d10359b7a86ce42187e7c
zf11f399899c93417304ad1434c81fb3af708b8ea1cb4456cfdb136da858180eab0119e94e2091a
zdb9cfefc0e3da07a2920178bec223d8c53d34f2b63acd117f09820346d561f771ae20a65ebddc6
zd40a7c2de45a28dfbaf90ac9d07379fd3d152ea7022271ff73876a7db01a1e33eb44bb0cfcafc5
z7cbedf520b0bc1b5bc1bf9d634c69f414f1e6be5984856c0f72695e810cc1e77ca5d7459ae5141
z36a0cba5fef7b6f669ea5ed71afea8a1e7263aa2193fd99a1e37f6c96a8796483a59a9d007d971
zebc02e29052959083a6306a1647f86199b3825ba4a1f532af0c442d51935228799d6b5a84bfd7f
z13bf950538d61cb608ac76cf734fe4a4f465611097009609b9d8af463ec36864b1a4b1305b2b96
z9b3f8d6b1e0132bd2e26a016940fff4af4c3af1f87ff5e7a199a9bf24205723ac70796dbf94bfd
z0b39c8f50e4db0c16b62241ea7abec1a96c76658ea57ccf2559431cba11a939062695fbf3562ee
zb6df94d7120d27bc289612b10680222ca2ee0b8603109a175ea700c02a8400e158c70a3b1ecac9
z997d46799b1d51f9059b0e6c82cbb02309dec3910bcaebd556535bd40a555eb17dced4bff6dd28
zb88a9f90aeb958a155f9fe105ca484fcb1f35b3cbd36827f014a106cdf86d933984211ad9001d6
zc0942745fc532384705a668f5c1fd670879d6744eb9f11ce80151b34d19ca71d4a78ad25b73d3a
z00ae281a111566592261e281f0ccfa5e2e9f73465c62f95c7cd0c1c2e10cb752d9a25c97dedbdf
zfe0304bb6363c4b22915dafa7668353b2786907b4a27947034cf34517b0ef8e4832005340d6ade
zd8c2a53e08a65235446f8d271368e7ddd250b28e687e32f88e5d1089bca65f66d565ffedc8a1ed
zb03c8a78fe42daf9b2499e4915ba7e4a718f8204dfdb0bd96df64a96f238330e2bc597766614f9
zfa49a82a237245ff57f1be30e98e983ae5126cacbfa8ea00ad72f9f9aca198f00015def6dcd4cf
z666bfc2fb66b68ae86d11c6dcfa53eaa1dc8090bb8c08feada09da7fb687df02ab4ea9656e4707
z8e806861e1496c7f29784cbe621253f8dd8b21bd142ad63fe8b3012931187ef84ccad483c280eb
z3072e935c11ef29955764a44cbdfac55646eff5f43e00d0b8393bf411e26ce2a05ca85e938fb7d
zdd79500357b8844a705a85564e7082d380b5ee0e979994480655822e22285a456a3e400b8eb2ca
zf18d70ffe9013eaf393614c3383ce0332d0a58271ec89bbeb3aa855d1e8f43d676d3dbd97edf3f
zf683ad5fa928112a4abe6774894bc606027cb4c15ba03a196a0044f9e925546417cf3cd0513ffa
z56ce560b79b98537d2ab46fcab86850e70eb2f7f12093cfbdff88857032f1e1a0b369b09689e67
zed511b48b3dde41fe7578c2c29ba0d546b4f342640a5cdc18e0366c0ede4d41dd17c62a02965dd
z8cdf4f1172c958555181f9b2b8d9661256982982e45e0a7d8be4b8e24b94441b8b32a2eb4a4a76
zf4f7fda8456e8d44b235e8ac149d30dfa173af0d36d33b918a1a79a184855ed28b4eb404e9ca00
z15a687d40576e29c0a7b14983b5aaeec7e9221a3c8863dfc1961f695d090368fc3180ffde1d0d3
z2aca8e63bee3d22991392dcc65cefb7d2b6b7d818da64fbda5e200d87107c3151f7f9721316f23
zcef1c1753656b59d9107bc955c5bc0701433963f205106532ddf63a390fed3c3db09c7f9630a18
z7dbd230aa120ec793d88daa59e9c3c406f5acd33d489e00b46c5f1f71e0715425269ffffe04bfa
z170a11fa5016102897493a9b790c1de63fb27a4ad5a6c70cbe019a93759fadf34551ba4e9f50a7
zb1042052f09eff392a9cc00bd1d6722844600b101d88f1a5d275f54bb4eff63778160d01c0226c
z1cdcea43ee118ee9620eb65c052529fa04a095a3a1d5dd16cf6d8fe3ee5680d35e4ea71e248acd
z5218df568deed8695f9baeb3b6cc795e763885d9d1c36d8633c77ff098dc6d1d9d401f196a36b2
z916255901e623b27086399c66bc8468b2777a9377101336a26eb6e6709f3b575b01850fd40fe0b
z4b669d0732e6e96a08c1ab3b27af95fd7b8adc91110bd470d1da529578b66ee5c93f22e35e4062
zac9b9069a269b17718582c030ec919a232f8e7b8491d539b57d82e055815d9d6acc41795d1148e
z0e1d74902c403e94cc0095c8abbecfe5e183257af4797b309cd2c6c8f7103027162d9140f05b31
zfedf0c7bbf55805a2c90f79d12f5a628f3227db5c139d923fc7a50cf93a03de7413c35d4832d81
z7e82915cf2578c74cd62acf11c02c6a0e085065145c0f92e745ce13afe31c50b43eaa08dc6d820
zbd1ce094d2f581fc02a4dbffcc82ef157e0070e539c4ee761141b96e544be829310ce5e779e561
zc347078250b3f70c33313fbc0e85e8a04555d542b0ee0d661476b3bb672e4b342eaa217f99a507
z0e1e8cd870cc5102f60005a790d4943d17821c1364f8f3c21bc4bdfee325e856252783951cb906
ze61cb44affcf0eaf00c40ce62ba6254b64de07eeae05cc823f4d851e2f1d402baf11d601099ac0
z8930c13d1486354b6e79622c523bd4d6421e1aa9e2e6214d168fd633c6bf14b0dc0482c0899ed8
zb4750d3b0da23400cef542fd8b3351a567b71ac1a391b25bf6f6ad202d99d8d3d3ffa753885915
z8edb76583bf9fa361e643d50a0dd5b6b0b9164bcbdfbd8f01874375e7212956aae692c87280389
zef0068c1d1e12cc8a491d881f9c046bab749b393bf5c6997970dc8bdc713d2a8daa8994c33325e
z0ae45834926cfa5fbe2dd8ee44e72ddc072a5225d8cb2b67b838648da8fbe7e6a6d50ca6acd7cb
z6e6ee02a83151f02748e281de125d4a792298e8946b9f6ad28f3f92153b5794e2bd1dab591645c
z2d6f93462d07421595b847f951017c7e8aae4f98217316f808d9d5743e40eb3a8e186aac517815
z05735832bcbe94e6a5a505807a1a2b911660207d567d193664334dc081e770553dbf5df281f004
z5ef8d0625ed058f2b28847b931874115309552fd006575a10999e17a3dfa43e6a1f04f1387754e
z415d6048ac0e2e4126eb70c7bae716e7f11aa080d3af48f2ef38dc38851f7db4d20bf92fb153eb
z1792c5c11247b5623cf1918b9828ca1113d39814aa35c98218af6bd03338ccfb257084a57c0277
z734c0b9ad297928827906b20f9e0e6d682a63b8ffe6c68f4b67d9878bb546d847f178fc9ceb7d5
z040427149201412135c99245f4b7c777f6310cc12558d18d3771ce88987ba4b7fb6204b881d4cf
zad0a3a24d0c59333bf375a1a77f3b685180ca5bfff65c279932a24b7e83256f570d956ddad4ab6
z431bfdf8900de2c35069821b955dcc2e40864c7bbf42ab096670af3172a2a1f35a5172d1f5b441
z5df5b4e9a13bc497ad87fff9674aca629748f70025ec49c4c505d70e71fac62756a8787d3627a7
z3701fc65e39ecdd77bf331e9a0b46f967cfc8ef8a235cffbbe7c57437a45d9e6e8b37671bd3b21
z66ffa8f95b81c5ee4d3c59ff9adf444c6becc8010d6bd7720d89bdb260ba5cb923d4c7624ac819
za2eb00863d6691760e2c5abc255c6dc5935c77da5174abce2e43d64b5717804c4f084608d48909
z05f2aed49a0b9ba8d5f4c7d8bd818d981a02ace08df12252771a92067814fe3e55614a59acea24
zb3bf6f0fb67668a6fc5b1437292d157cc0e462046e15d8decbba82eb4267f18657dc6b92a4d8f2
z3e4e8583a507d42b73724626cbe27b7523607b5ea8684bb10cfd73c97ecc4abcf00b8c2d517b67
zfaf9e887a7be99a998979ccf2eb9bc53e6a35fe574c99ff04f61e34dddcfadcf8dcda939baf051
za67932548bedfe0ed0db7505b7e95e77d2e4847809a1db95341ddfe81c8de7626128b23ab39f7d
z26f3bc84abf3a2291e9885a559f88bbd847417b1bbdc6fdfab62fd02a6557694449842b0d412bd
z70f85b1e8bb63074b4c25a1acd48e213d62bf4742be9cc97e4becdb80859def1bf68239fd268d2
z3f1384759cfbe59801683c846a7eeb89da5cb537f63454c3843cbefe0c23642ca3c97e4d183f9d
z07077b54198b10c94c721e00ddd3a80d7c18e5cccad694001401580620ea62bdf2feaa50416275
ze237d6af8d63ac011297909e112dd6c440e6331265c6c87d03d3abcce8deafd74cf8097dbb0e0e
z92f7cdd3c5f8f3525959d0120d401b088d88d4a2b61971de3b878498ff730b927ca388a48eb567
z871b7758e90588806ae02d428f8f849822f078bad73b39363ea0730fe5a8201fd138f36dc748ff
z87052a06bcd7cabf87b2b5bb800b896c37a1149b010347c3523febc55053700e6f7cfa4b8b2034
zba0fb7b291c3dd01a19e994de3cf1107c11080606b529e59bb80f3b2a358ad76b2fcb2b408cf3e
z9d8266badd386115bd4d50be52755565e3388c82d8ad0e1282b3f110eae56093f67e2872ca98db
zf0a1807f08b4e28fd6fff1f7d08bd77dcf24d5fe4526187b522345f5c0a9a092f46ffeb291dd31
za3de30250b5da92bdea7bc30bfb27afffcb465285d820d3f05048df9ab9f73e773c143624f6258
z242dc949968efc7931c3433f76a06bd5f3fdcaf5c31d66984c2ce445d6fea255d3ab1167d96e7c
z81c0ef774f4a313a01973de59348db1c2ff130dd658d7568cc98da05d92011d8eaed339cd73d84
zadc91bffffc9a6837379c7c7912b9699598614de24a2f96c46b9f679c198651afb2a4babde9f74
z9f8804d34ed3796bb1df2cc77fb55a7b940757cae365be473d4e1c4adb894ad2041e3d93549e02
z9f3462edd72a861b57afb2e3122c2ccc188cfd0494227ec503b3f1ce3220d2dc50befed8f2e757
z58a5e0f03b535dba4ad105a232b212d50be47437c2115dbca98e5b8bc855aea8a1a1beb2aa6003
zdd7506c1b3988e2a50fff2c5fe8156db19b30269351445e6f4cc74d8e41270cecffedafc7b85bb
z9c8424387718e50dcd4dc1f20d2cf092acbfa8445ba3ad4b14b680ad78c3335179475aa6c5caf0
zdbc3bc440a49e9528cee8de7e3337bf63179a37499145be8e516b8ac579cb50fa4141ef9c17ebd
zaabc194ab70fa318d59c1b8890df0b15d924d0e5b9622cdf3f4c15cde9b5148cf693498f24c469
ze9f4c8b9cb2067210fd9446a03815d0162f89e62fe76391c8606c49e560ab32be764694bfa14c4
z0a5152ca4a648107fbb20de8e5d066421a152a89df7985ef3fef981fa11a8d9f30c917f9d987ba
z40012ab45fdd2280f9cd58b71f63a427766dac91aca7e12e0af7997f6b1182fcb9675e31457c7a
z17b9b0403edb9a26c2a4b72a1ab256723476606d8be9f0a5f3daff6765b8f0013bbe7b9279fff1
z951e64d647305d75ee124da8270cb5063a2155675f4820f64b4ab85cddeaafde17ef887f112974
zcfe00d45afdf480c8ee19af290aa1127f0a25f2a6f53fb7ce65c3f262ba32b0f9d3d8e6e6745fb
zd290a82d42ea760f8998d63633f04e62918da1de3b1a9d4b27299ca6fd97203518e0c297375a4a
z828b7be024bd603ca376974129333d9a48358683b1efa47bf1583ee520b4bc8fb1860173bd6f20
zdf40fa0256ca5a665775189987c2f263b048028785c0bbefec2b30acf63e005204261285786ea3
zc2f3c02546a02a25606e976319394f45831c29cd4d62702db34a784e08541685f6a3335495ac83
z0994b52106ea27fa78f6d966a99b5e1b0f4c78d375d0a4d253a4bddd6006a82240bb9c42738bfe
z56a28d54a7950a69eca4ec8c9b3d09474a786e059a9b08e25501382acfcb19115bbdf7dbe30fe3
z14b95771e2cb14c34121efc3bb8c892d40348bfbed047b12f69bca03ca803e9b328c56d30d9884
zfadb5945ab186d4fdeaa8889040c495edc6d4c35e5d3639a7d1b5c7556c9ac5782eb6335537c0c
z07a6d36256670c6da947060e547e82857b7c1f68ce9f6f49194b59fafc683f4857becfa0eeda99
z9770f9e4459267797cf29c7b57d31b81de15fdde09ec0a7895e6c7c284e35118edf6bdf70bad65
z0f4f08a721ac5ef860de6769c3f9878ed74d39d83717aab49b0b11324ffc9316978215bea5e811
z7357bfa5eae3f28b1089adf390c42b61f475598abd8ffa5f5aa30ce7a04443d690edab0389cf5a
zafd2a419545cf3307414bb5e82263c735a6a73b797e1a1c6c2d771c9feed7a498593bb314b58e2
z5d1f3dbec135fd755e8952bf18d6bfc66e8cb97f635b76aba29d3dc9edf5a09c80198343b3c3b4
z804425cd1e67e2e69f01ca6313af39a31712e5c661e735d76e5a1d3294eb2e93d7fe78eadb5b96
z88fa457f3961a1375e33548c2e74342c6a590ebbca088f9d8a6f8f256c6c7754ace2155ee9f67e
z8f5ee13663a32b34cde222f22b6e0a7eacfe66fe88fcbba674a19f4827176e1ec8312180dc9adc
z24182e73e73721330772adb3aa0c52e1aa5e218a8fa74ea9d00a37e36fffa92ef00374cf8d52ea
z87870efb41b9e658efecc474c48cefc1da9ed266449280eafc3043d3569b522415ff6b859c05d2
z2a97f6aa37f0f10c56e4a06818d2d0dad92b2e6395f626cc614c0c7da76888b21aaabcdca99c15
ze598fa348e2edcc43642413034ed067c43bd8f1ce21509e92cdc8ae3d2eb050d65b755b663cf90
zf97f56fe3536297541d8b94fd18107b58c8f8e73e4d468572e64ab660ade82d56846f0761767b9
zb65fdeca778fa56393d82d7596d7999ed12d71ea032d6e94b186a584661a82019cd0786541892d
z1e2cc2b9b24b2ace7b9846731cafe0a76978f3825e45fe562de763d79710c50bcd3abdb0cdd021
z4269b4c4d56218796a26c462f642c910a1f41016a56a46e0a6e7debf8181355ff1ade470be2c52
ze87f7bece192c49a7070d696b963a7544279f63fa79f30faa96996cd6fcb32912352508dc97717
z8b1a5e7e9f3e80d437407874e9351582f60518939a704ef0a4c9de2b6d3dcbc1778aa9e5c2271a
z43aaf022890131b21db37da16ec3c7dd83c36e5e3d31ef7c7a0105eea2726812578b17007dda91
z89c0ea0891e8db83dd65deb12f12754dbb16a9316733744a9824f0a14083977676dd7b97e7ab09
z04d472b6fe2442bd31cd03b6a12b6ba819d76a3d88aaf8cf4f80e210573692b585705368a576c3
zdab0a3aab6207d368e5bd7329829156e7674a23ae810db5fd81d955688cf8659238942a0dee8bb
z73909bcdda66756ce4fbaf3357f4d212b6a728c6f8093694655d97cbd516ce1ce69ecb7ca083ef
z3b135e1ea7d61edc5b5b44f584ed1177e6223a979f3eb56bcc85744d4c0b286b0fff86946d5781
z94a69ff000260101f5be89a81d43170804498e4b24ab3e5f49bff419dd2564f0e577562f6be151
z12db5e403b53d759e69d1b43a4bc674c39a3d2c794218d7151ede1108f7a2f447454dcd221c89b
z2002fe9c164d31166f9a364eac7277c9cd73c05232e841c3df84c630d2b450e2252a155b0c40ea
z9294ec91cc1ce518d2c4360102b74b7352c9631209268b7eba6786577219a5198538876bc664b9
z592d84fd59fc6ffb727a64d787dd0e9b2aa6ddc517262f3bfbf8ccd6db61427bf9159ace13df22
z08de114602530b279187a9faf7d426177ead39a9673154368a2c96f5391ae93ac0b05767e927a5
ze0203579632e2882ea9d6fbc45bf56a6c8ea614740d32f29e73ad7d6cffe08e7e1d183593608fd
zd3dbbb5a723f4a9e7e7685e7b2237685eda5075da85aad4c1db0d16564a2364c671f7bf92c6f32
zf14514f54f0640a809c9f8ae91efa67994789c950c6f1ac7b618fb05165da33db5651ef9c1130d
ze1c26d97fb5dfac91bcdf5b9859b981a40daa7f8eca10faf7081142111a4de1611aa6824d18b51
z08ed7ff2f289ec47ce07d07704af5ce6f3c742dc04689a8fcd5a8bbc8fee8dfa8b68a37dddbac2
zaff1155e42cc49cdab182a71d2dcfd30a851abcbd6993173de1a15e5363f169eaf7c3b8e951447
zc32373f948da0b9013a8108b95e69990439f093939e242fc7b2116ea91ed9aba50a4d381e4917f
z8b84cf18926730b57e885079213c9287bd5ae01f5e42d246ff99a3739864ed0fa0c27983695ccb
zecd7a80f2ca59bb60d1f3c76cec6331a309e35ff4c2a0bbd1495c0386a09cf32684f65284d01d2
z71ff20fe3aa4d79c4a95ba8d6d2f37c94d8a3f73fd3199fe67dcc5b767a56e8db25c5d412f67e7
ze061db1888e5a6cb4f07ad75c459d43cdf0fcd9790b4acbc7f92a32185e8efd231bdf4c280744b
z3f61c0aacb064f3b8c43ecfc700c07ff7e536f337acdb3750c7e4e1e1855266faf8c2e9fed3266
zffbe3bd1c5226db9311ac6b54a4d4c3a12116e9d4d35940ff174a2392dbd0c72cb816ccbd95721
z93945f7dbc92b971b7ea97028b7e65d1a5eb4313007bafca1a4bb688e1e5299757871c2066405b
zd21427654b31e2949d9fa8553929db0984332abb41514acd2fd950cccecae9f9f92f9a3845cbc2
zd12123894cd582873739dd3cfed93dd599c57978fa1d37b802dc2d4bec323eadf8a3ee0292f427
z29a0cae9fff79455528f4de6f8ffef2307cd0ac5b74ba04cadfd98f9345cfac66009db970ff106
z4c8330215cccc9c4b905acf564b0ee91f0c41991a463bcbf29dddb14926337e5ec123da53f6e6c
zc0458b79bfa55223a669c50bbffcbf9e5040efa1927f2f5c6836cf8c0bcff8355c5735799a4ec9
z7fb11391c593b8bc4c4a402d3e16fd1b26c999ce1c582560b9bd0bd2c40514a83d0b4ff48b1432
z282dbc9017523acb87604ee6c068fbecb11b906736ce41e1dcf4ac403719448ef9153e174cd4b4
zc9cd45788bfe0f69e915d757b1837fe8ef3d51dd3de493200f44b51c3d843255042ef127fe7286
z3f079c189c30bb2adf8c4bb8acd355e5ae693fc30d702b7cf019d1154b28ff64716aaa6c0c7b1a
z6dfa2e1e1c0aa4906908248c99f83f5fe34bb2b6e08da8aac479bd11b74c452be765ad09af0782
za764304f00774048e1496bd2440519495997bd3b9d570e9cb897a5d9d7e8504efe1d2b75037945
za1d57b7850adcfe077229b591ebb53d5cc900eab2c03c3c2afaad55ce1a082d8ed51a4b71941dc
z40621f90acb55094d7c3328b715002f6dfb58122ba0cd4a3f4fc8f1f1fc557e40a104354e03d5a
z2e2298b0a1b07931b39ff5e595ae522cb6ed2753af772f2942888b27d599521ac14807d88779ac
zef094aaf9e02d4c091eeae5b7bb992472b264bf88ebe0f696de03fdd3fa62865e37104ed960098
z7f3f6c780bf183dff886c588c5ecb324346c1be307eaf64b70e3a536ea4f4b309e0bad8bc8b214
z8b023d00eed32840104c49d632ea8271ce344529acf6793ccfe34c2d5da8afddda757700c7c89d
z94aa67dd18b9d41b4df2bcbf4c4601c383deb841be645a2912be95acd425eb297e0ab996cdebd7
z14a47470bc86a0453139ba591538476322f24d5ed56a499eb0559d30aa7ccba3394d7b0921e300
zdf0be20accd6c736af34b8bc5adb86fed7b1478bb4f459418e478eb92afb1985dd50d7a5e90686
z4793ee41fb873585bd6edb60bb2eeef42399c1cd78f1423a6e52d5d17e974bce62cbcd3a0a8e40
zd84480bfd3a82802c00e8f273a30a29ee806f6586d2bddda38b8168c442796dd9cea887a224d22
zf659c89e37b469e138051c0d4aa569478ef9aec77146ea1a11d5cf5e53c0a4f32059dc3e030b90
z800dfb5d669e9a002fe037a3f31087f158ac71e6d6f3e79aaed240f7c09000c74308a86e6a89e2
zb115f0a3ccc46701e9c8cd8e44f218e6465e4f13660bc36e1965487aed799a0ebffb0ad661d23a
z10e0d91942d13e9295d7bf74505fbd638f5ea076724458e96cf9841f91b214eabc7fe683447576
ze3eec21109a5becb90cd5b1986f150133ccf0a64341aa8ac570007bc302938250f086f7528a49c
z409fcc7f6d8791ea5f93e7bfb8989e86d720bf4af6673e845c9a8690657dbd417427128dea89a6
zf055c801b9f3fc374ee2b411ede404ce1b0055e30c5e1b8aa2fdd69fc2144952b3e47ed96d8027
z786f0c382b46a85cbf016baebe496ceb3d7790bbc1f0f10c6ddfe82e37272aba25687c8cc9b1cc
z32fffeefafee84d20b7578d9f2cf2690159c17867b7980462c1fbedea93690381ca728307fa78b
zfbf5cb154366bcb249bed0e930298acdf06cad4c8834b4d1cb62742b08f1260c26ea6328634119
z762b86f10045b025fd51a3f54075e752be73f3a937a28e13162b2d4096bb5276d32c429a1059c1
z65a7b00cbdc32a50e0bafce6b875821391b1ea0b7d0ec84c15b43cdd7c855720b0e9b0f81614e7
z20bf144d9ea149a1715f0b1e3657ee35c8552e3def0fa0568dea16e616c8a2099f741205d1e9b1
z7420bc512e5341a0babd10feb2b159fb989690f87276c19ce3e4b155eb29a32ab34b1fbbe84e88
zb91864fe9239d3ff8db210513c5791f9a0192405d53050d03e75c20763ed71852717fd3fa28715
z4af7d22a0da8ee61ade7ef7d39fe450ce34e219fc08d0eb550f9049b9a6560c8614594fe23f46d
z0af16b6d068da0d70a4eee24b1d5c08a517da21fd5c03a1436e1d82a0e43276d030201d30663d9
z82f7aaff5434774835019a6d8b262d7bdb040c0e4cbf4904ce08ec8da567035eeecc5bbeb86ca3
z920f675353f66bc91bb5f226ca55c2909fbf572b6a224ca5329498a6464bfb42f66c158dbaa5bb
z9552b110192218d484e9ebbf8edff09224d78af33ff488879e12ee6d9b9e6e8e837f216f6ca23c
z55e35fc193532cdbff7f620ebf5e677bb9588e1fe0c857e9734b97a81114a7c6d9192c6c657383
ze291d33c885abfee7f85513ca11072c47238cf725ee32269c8dc099d68e24d35260c1a32ea3f33
zef66f423dcca76091eed40d806115e5823b138629166d45a6ed5f84ca8224e1a0c2f148c825b35
z4f2543501d8aafe22da13783d00d5df338b4dcc790149f59845890b225678870a096cceb1a6f1f
z46ec19b1a22834ee6c2cb05a5f7fc176bb49a7786a627833aa0a6b31357a099c48388028c67728
za96217834dcdebec301dc6d12b31a8bf946b02bc9a91f8412bc80f1100c6cf82a7c575d6966730
z87c32394339f721084b9cd8c114eca17e74ebf66754758a29f11bfd68065f410a7592f08390b46
z97bfedb967b689ed04e939f6e435dba3a9359473bcda401c98d25a0501bad96800df78739331a1
z713ce37b6379134f1ebd57fe880035d107c24f733b3e8a156b1f5daa6a79dd04243e21fd8565a0
z34140a805cc258585fe918ef4d9252409cc0022c243e96c0a695ffb671f30ed2f94c42fdfdaddd
z485df9e9f444d0dc2f447525d87e6c91ac54c52b8b74fc981940b6005b32574b5993852f8d3233
z0121a2915602c2f21d42cc05da5eeda0cc01a92d20ec9f62a2d62fff297916ce9d04335cd87cd6
zc3e8c8367b13e611dfae4c3ff9caea9daf58b4cd0eb2712031d3eb9826299b33339e27f5919b02
zb11b49f3b03d90d3113d3a0abbcb746cdf6ff3634c6b916e721f61e3e5ed093691692be37f181b
z6d7b5c9710117605cf656a8c55d9a1f1d731c25efe0e78f3a7970e143baaacdb41ec25f5ad72cc
za644779c0cabf09b0d39667b619bd10ac5a13ae93b4f39eaf1cce90077f76f477936f97d5375d6
za224968d6aba75cf0ec05390218776cf8f1442347dd741cca3a15c82ba7b01984d709e6a04f711
z264bb75b22af465a51f617e7a6fb39110c03281ae0360f418878105f2cbccb819981b021f94310
z92667607fe21996f2bb94891b5ba3efd8f17dc83d910dd30bfffe9bb5eaa72283b1167ce991b40
z05824c69699fc4d1c8b76ccd16f7d0bc465c0adfc2418a056abc94e972764a3e9a93e15c4acab7
z96a2243dfe8866906c68bb267163f30ce1648a4cc52bde2c93f94e877f0075692b4ee7bdbb3002
z2292ccea305ba5ec6b053cf4ff48d64fdabdb34ca476ba9acff22eb6c3493a84a346235029c246
z2d79eb265710549169eeb398735bb4d006df62ea424bce64065d9c72686cab79869820c3f67625
z46509c100455c51f7e0b43b1a58e34c1abf3a58a7133bfa5a685c68772fc25dc1492c5b3f3e124
z35f06f70ddfda70da784fbf9e08920b7efe0d27d3667751913c2d1a045f08f592c3ba2e9dfb8f2
z4005f777c5f0e3c3c933a920a88b7a2ec66eec6179ea529ad57fb573479c6f471f62c8e1ee0964
z04ca836c8703dff01dcb5a7a728df5c2de7594ecfbada02b6602ee889792b43ada9476e59fcc07
z9d9648cf02552021208a918abfdd1d2ff4c44352e72c8e43b1fc80960d63b70b4cc1d2ca66102f
za617393b6753999bac2853915f189f6c65df145b556deb2f08b83a8bc8614f43b3f7280de94053
z236af14b33e24310202701f220b4b0981d977dbf65f236c2edc72fdeedcfeac4f11ae5857cf3c6
zc2ded9b9eb19990b07273322b36689a6a2e83f2773fd7a63b74e5b48035334ccc526794897c44a
zd7247eacf4eb0472c4d46f937ef987b85494d111426c26bf029f0317b3ede8e2ad5c07df0b5ce4
z4288e2765d1e86964313574d23d7c3c677d64be1abe29adb8f3b49044b8cbbce30bf5959303f4a
z90cdb2a22e32578582ae7e10ed68309b61b6b893c9bc4f5c5ed4d6405908078ff01821f04fb35e
z99a510b093d35678373bc2bbadaaaa28d73613fd64b2f4be237d0bbb5796f3c6706cbf95340050
z99aa8a9936605598330a6ece3f20e5410482fb7edc4c382d5bbd1692fc8b3f174a14647ba6ce7d
z49841c53774d8094d73bba1dbc7116241e50f315a7981613646f1d51d9faa0f02d8cefb4a52a47
ze445eb86bda090ecf42d69d921d00fd610076ff6ef2d1c65aeb444c95fbc882092884c743e3b29
z614e6d389b30e488e6ac0ad4b099346b7ebeee0c962a7910beda973bc375ab66742bca51f4d94e
ze348253abe60fb021195cbd84eb7273e3ed305941c8622e2d1db9df56d6d1e4ff166681345ec9c
z8761c543c8ed94ec4a76f5c94671cdcd815b39c0756e30627531beb05a2a70263a10559e873d31
z7f69e6947c1881d2fc5e0dbdf7a02a207db12fdf897ce4029bcf0d73834ac500f06075fdf4e050
z356eb88fefab05280fe96809ebfa376592d1e55475c6e97b499ff466ba8bbcdce3c63168368281
ze0ec89003f6380a7526f32a2fd9d4724d2e1fb4c6379c149bc993ce54a5554416a750dee93280e
z78076ff9546ee6ab5c8b05828f3779e74f9a418a9facbd5c2c1adf54c7b634f0fa8e58be17371f
z0b188a85478c55454cea294763dbd057695f79c01ace640f261093d1a43e38d83db4559c909c8d
z5044c64cb5554ee9eac9aaa6eb91f2e4e62cd7195efad6bfa663e29fab11fbf9965aa5c07348cb
zd5e771d7072e99f1e668389398a82a169012d499304bd8a5641f75901834f32bba5c4e0bb31f92
z68495bab679a651153d994e05a4cff3bc0e98a0cb33d2e7977e90c479b0feceb1cbc993abd274c
zd89cf80c9e9bebca33180a14e0a18a9a913fce74b0c618812443fa140eea7f4d036e96cfafd5c9
z00e89764c91cd2940edd921a451700d21560e7de94884f7b93b9ce78ebe3e8b8ca59f7b2c6859b
z921d0f5c3958b6a199356f492418b97c56536317699d9808fe02e50452011257ca33972600d434
z633b214a4d37b7d518b9228734b1e246f7068d666aaae35db44719be00228ef98cb3defa0d44ef
zb211adb512870bd0e3e90faa3d6abd12b5db752de0c1dd22ea3fc5a845e10c0a69a30931116266
zdb7fccb63bd306d7fa45c215ce94170aa01ec3344add538ffae37388ba1738fd03931e0d20e95f
z4a4a98feac79cdf8e113555d2ee0addb459a69af4bf2e415606fdbc01077d79207eb6748479225
z252b558dafcd98b11f7ad99bab8dbac609243091174995c9376006ede56255bdca451954c88de8
zf4bdbb9bb47dd19dfc2d1fe396a11691de34465bbe9b9bbb5abb3e55b8d66453e50ee9ad3aac09
z2ea837cb7c8ad81007b0bb25345dde6ff0e91470ba747c77f0739483774d8a8941c6a44c564e92
z5b2a6c678e3b2b9f2d5bca0976e0b6194bf07e426856108c590f6e110a1a6df9ce67fca344f965
z1be8b935047615a902b57929d94c1b5bdcdcb95e09fbf3b85ecb01d836c56329fe86edd85de359
z25a924030a3e95d1d65ec1df24b83b42cd428706e5c240de79b509c6ae130a78a7909e34422821
zad8cca6a74852e28673195ad382f04945d8f8eb89c7185e4581485076698e9e76bdf5707e592cc
z646ec18320de3e10014e17462558523e4f633b4c7b9ca1611a56da940213531efd764a49f9d915
z25ea240d900db30c99d5c38fa8d61b3064042ff29d9e8fc429dd08c2f2aa2ebba1d0d549e948e7
z23a3b11f441a19c1fd6f4bad9288c8659142b9b62836b4020137cd0ed0b0cb4a5ddd6bcc782a4e
z2b4d4a65243050e4d529d64a8ece1aa361a57479364683a2869692fcab0c197307ae494fd8d77b
z049d4256f00dff8bafdffbaf94f00424b78f221e69a6493020eafa4830df3e5d1a614e1c5bdd93
za689f9ffa96c6a187eb616eaea1931fa37cad4566ffb7d9205050d997c9fb806a076bbe7a66f6c
z04b8c840a03fde0d96fcaee9f0e3faa9526ec17f91d894879485e4e13ee6f3c29b8e64f09e7534
zd01fae71c65e283254fa906fedb3ef4f22cdea48d883372e1da0a5b4b411b8498ee16bd5c79961
z5f610d8093334d541b151eac94b8f04a2bd6c8d3475e0d85c83e0150f6cc861823ab002c2893c0
z0b7c0e58685e859bc7b305bc9da781b5d6239e9cbfa268201e5a1cf69d73923e8639ec67ae14f7
z0a3070b685c1d8599c488e6dccb2349ffcf0baa13df42e5f116330850f53c5348fe6127209bfbc
z7a1a23298e2586ccb8905101a3b92e64da77656f0b0fae5114e133b787ba7d87e6cae67f746624
z45beafe89a3dd32fb1241885f7144aa911a4379f1748b59daee75ff5f48e0e6ac4a8476f6e3185
zab31d4e6c749fb208ecd4bf8292a1d5c7ae334cb72dc49c3e4ff96c456c66878ff1879bf389837
z04961c483f122f2470ab084493bd2d6e00082dc0ccbe58cff88aa5cba580425472c0a7b24fe6d6
z34661f92d5a6dc1ed2d3271d12177c4f99956aaf93f90b319ac004478253254dac83aaa5ab65e1
z30bae1c50d026b5f0b5c457819b4495ab70fd1707e5a0c4e4f42850baeb630096cc3d1b2e67a64
z9eb89b1255c6cdff6435e3fd6fb9ea83f28b69a74eaa12f3ebf9f0590d98fd2896a91ae0127804
z7b77dfe479d9a0ec8e34f5b77253f140c2d1f7142fdaf186ca4b9e04cc4ca990e3ba4ce44311a6
z83fa9f59b6d47f241d2cc33588210a8017612968b3edca2fa48afc782099d016daef74bc873d01
z667335bc7c25a59a1ea0e7c6a76b09bab2b3fd28ce0f1ac5bf571dbe1091d2796785bf1503a490
z71bcbd1adaf3bbb747d9c1cbd0c2fdd0eed304514df28edf7560aa1643153be2a85dc44984efb5
zf7b02f58af199ed413527a2702d94e9b3a479bfe99713b4f86d2c3ad98accac536949c3695e3d7
z16ed3b7d189ea0a4e731073e108d9cc9e804fd58f17c2f3628cd311703c916272198655a5e3317
z6b0c76c9df16448249b656bd32c04b7bea19385da0b31d83d4d2ffe12b96bf93601e00297df985
z07848bbc95acac8e5c13b1c033c01b97630c62bc44d43dd3db1823aaffffad385b883de0608be0
z14b4ebc366a7f2b3749f62e6b951bbf4e0816acff66267fdebd8d4c87db5f75a2d6281532a7996
zbfa89e7d180c37436b28408b2ac823b09c6d60e9394c3cdb4d3780180637dc9f42ad8c69bcdb33
zd6984cfbcc6b92d663effbdd77b45693aa90ffe808e050e46c8a1298b328b20c05ef55591d6d8b
z3c6aa997604fe5d98bcf50ed16c27733d1414351fd2310f57d31e34917a9631703261acec0f656
za26e7838108f35b02ba408bf90001bf10c56871f7a3719a2e024a6f9afd3c9478ca2eeb7b609de
zecc6c95a385a7330c4e183cf6045df7eaed2e94b40e1e55493345aef4fce6fd91b007e6cbed999
zbb0c7324b9d33823245748d2abcff953c1e6c01f4fa6236fd8fdec209875ed071130af8d998803
z3ddf4204f9acac8b7fd94d5677a17e541f5353776aa05c25bf7b3df59d1e16a99633a3df1fd133
z7a0370eae8b8ea886a707ea9a19c00f7582dbdb4d89a713fa7d311aa9fa6304d74376e8e9cecd1
z8a5697ccd75923f5efe6f0e63005dfa922c4c4202d651e4afc37d4022f935a7691609bb52e6247
z69cc3a76535c8a1dd3d8c292a807017463c0bd9f4c5efaa669f595e7896d8ff1af1cab64e2bf2c
z9e04643b221e27896d53ad29b0fdd37d109c95a1367e4dadd47b22b8d172a6a34007716228a6a2
zc198425ed679125e9c949f3021bd0894caf58df8144eac1ac22b8dd81c7d6bf8819af23ef761d6
z9a96740dd64a5c55de2e9cc2c5a423b0023d9e9db492bcf4be58e8ec7432ac23146dae53768ac3
z97f151a3660b265efcfb98c38c14e6f1f689dca1f4e1cbeb6cb8ce3d68368fcaad83de94321ee4
z9554567ab390edd53f79413095d94f161997f743fc3bae94197d534f64ec8279639226d1a3e716
z2539e9ea73b89f4add90d10ffcdc4074a23368bbacbb95a4a6b9507b093b795780c8c294a5aa87
z345912a6542d514d84be7556037921cf2f2411965ac57a60e8cff13af23056a8fb3a3cf0630804
z95529ed1aec6d9cee034aa263beddb12897b4ea19ae90174b2e80c79e54e1c31c2c64cbd28b6c5
z558afcb4209f83b360a67718f02264496ec8d0e51c1797ddf8f3bed500b9c5cef82119744825a0
z39d22efdc57d839a8cbd70cf60ae928c6820c1d92e38fd0d24136767d652b9af732379d6493892
zc2ee8f440bec442f3534f0adf94fb65b26a19461046431026b1e0533e1cc179319a573cbc590dc
zdd66ed394b3d787960202678af7e049b32ad965c8d6cc8cee7e27931fdb31123e4f67dd7d0eba9
zf7de1c16b95a72e0d36a1172b4f90a9177459146292db7846fe8465825ea7f0faf2b162aa852a7
za08415d5ec25a668a06d309d2447ad724bd5d3c711a3386a078da3a66026de20c59150263da05e
z41a1e3e7f5d7278b52f81ab9c6441c6a5a16990e4b87864a13629363d0bf4cb206057c4c988f5d
z0356d81a049f307665da3312804849f1abddc2642892a7888dc2daefe8927523c09454172c2154
za6784ca83caf0eb94cb8c89a586bdebd87894595b3bb6aee8be9950a17d2151007740fd5742afb
z4262e15da50d0547ef822047ad656c6f3e65e0505f1a943b46d4686946d33f3c1d5ee19b1de1c0
z402ec8206f81a01df47f95be218a7e158efd9b184e35354963c3a09b58effe8613592964081d0b
z4e48c0aa831d4d40c50bccc6ef8b25d0d5f21f0741b8141b7e172c013f8e6a1c9d70fe4790840f
z155e184277703761e8b0c03d0bfde8460f1b8bd84344d7a4e147a4361fe5700294b52c2c4c5df8
zaa0da928405fde17d6a2a8d81857cf870fa2a58cd2b8036578ba005e752d211098fb1dc096cbe2
z7fe009cc20ec6daa28cdf1729ea4566fbc5ace4ece7c246d624e759706dee8edb362bb543262b3
zc9fd550800763cff925c8cfc0c70577b16048b0420a859c7c364fe02972e8bd9a07099b5eb0d5d
zd86318168c19f55632b8e524b9b6e198c39afc87221a51bb3665d9423fdc3df174b36075aed702
z27c1b6896638452d4a446628eb6756118313bf0a912f222f258ea7fa2f0da3ee6d92738bfd41a2
zd079e09f6596f8542b3518f9ee337fe27749d03caa9a67b225cea074a6749852f9ffc5ecd611f8
zfbb530fc86384abfbf82f6af5289b872380120d0fc44c2d5ef5ceb83300535fab83c99d76f917e
z3fe3a84541e85b86e2b67b637787d1871f5223005123d0d50eed1292332e2fd004627cfe62d602
zcd387f7ba5836a8fba3f639f2f0e8f87bc2a01f03e6e39a97f5ad88b91c8051909cf995485c11b
zcb09ba88690b09de9e4cb6adf3dec295d87da2bacc11f0ed97897651fe101ce551eacb28838208
z39f5d836b0bd2ee5b4874a32f56c5699806c1b5036eaae36d9cea20983f4fc5d6771f1d45de13d
z63c44d2c02574b20184e4e4bd44fbb336a0604b1c71376e7e0e826605ee7002f721b4f411b0744
z0b1ee4b3c0418ab7644d82b71e53ebe3ffc287e733b4efdf7f4c9d5fb5ceaaf83d6848c55a7293
z058d7530f49e37f9d74e6bb021567cc0bcfdcd7d82b8385d2db6719cc7c32c5baaa506fbc2db4e
zada6b9bdcc75b4e1cfc1579310756e3b3003a5801dccd663edd8dcd9903b6aea99ce3525c91a08
z7fbc2ed93d97e490f6b7d0a48911b018fac1e1a304640314b20e564202cade318a7413eb4bcd85
z8e64d7cb8f7021db4cf3423d71c74120749592e9b2b4dd60614b3d7b7be92d071ddbb023eeb737
z35ce3e55e615747f712f33f8b2de4a8378febcd03e32f9ec05571729193933ce8dad4c15bae096
z6520779b234f7efd3d9640d3ed163612835b4ff2dfebbe934717ff1bb59e6d52228378f8511f9a
z6b06fe4ad8f0a4d68f22e6cb6e79fec2a340d48eaf7920ac4a96a2208b6f3a460896f38e8d54fb
ze35c20f22a8d933d9f81dd11ec0bfc377e600e9707ded0cb96d853e93c0f07049fc5de8e6004ce
z38c35970f7b8ee083ad843929a22db762419950d51aa5d3b926e2b06587d7084de3b1e8804a734
z32455da42a465c32724c64e041618650ca183124cfeb7a9651365b6b4ae2e4f2d040c670483242
z30bd95c277af948e5cc52e4647f7db105e6160ccff73eaaf1d7ef2f5b3e4fa849665c1aece308d
zf12eda7810b71c11e992d4b689f00f9273a24d04db296579107d6047dc39fb44d9b7053070a7b0
z7759fab07a5c16b35bf867af0b7b72f54533968e019a3f5856fe4985b8772bca86030d4627a015
zd0159681fdb1f4ee2c0781392a06fe104bc99602852008ef71bfcf6babb44f38ba6b83356db1cf
z5f1a5f210daf5b909b7053af17aea1908fe83cb71907abf3611cb556683eb05d305dd6cb512b2f
zb044d5c92b2f421b3f07dc447915e5e63b70f733361c52f3acc2e1f8b11cdc725c314e71162f2b
z6efb6da35603162e2e2a9f4e31a728e62e3205122418b7a833b11791ee57c83f4faffa51d53fe9
z35dc83ec69ab81f4421819f36fdd077f5ddb344c2c75cfe179d8027e48b278a1c60161ec28aa31
z8caad31a37ca967feedaa6cc3dcedf88402a0f08db95c2ccb00cf72bbc777f3782e96a13880965
zafba861b5205ef5c837f001c8cbd1bbd915224ba7a8d214855b1dbc8d770fd2360e781692437b9
z9e146a9e7ed510136c796e49bde5c7b952a903741c3f1c64e45d05828aa59695e061afb660a918
z705b90f9cd2758de48fe0e7f620a98b625aa50b301f1f2d0cfc9a7e6d5e0be8af2681e6f5348a4
z0b9164e6934cfdc5eaa50c85e700523d0b43fccefa67c607b60027a3fd90a2bde093f663d9e2d2
z7fa06fc80657d566fceaaccad8a13f1bb34cfb96a6edd2aec6a02c26606a0d8a5fea5e195808b9
z8a727f98b9104249cc8c5855a7e9dd0cf918c10d4b69f0d54d65e717e65c855e409ad5436d1480
zb81b40f58577982db09404158680defae6e65a065a2917523eabb4938e0940771e8aeb5426d582
z8a8cc33c5e7936a9be4c4fd8af5f16c158110a34e1cd04638a372cad321bfc13749bf245925d0a
zc55da5cc932c530468e99b7de0f1fbbe4e2436537caa4c7c81f64748d737c6612c61a85d34f9f7
z680b98982382127b90d1f906faa7a91fc98ebf7d72df327b1fdecdf5b0f668bd66135a33404959
z5ed0ef9a2f782a38e170f2eac84b0ee74f39979f48a7ff8d87a12f0b03c85fef0213f3621666a1
zfc32b31e1c1d5d286231c662760d19596b12c3595cd622f4b2a422c51ee91d859019d2253d6844
zf652bd994d37b5faab8ac5046b89c399588eceeefefbcb161d36a3105f7795c97fa69a0b952a3d
z77d94f503339436fb31449a70bbee4e5e82d6c56e6ca9c304deda6bb06c34942f868d99da35c29
z1064e0b0f28d2ec725e62bfe269e5d7bd4403bf06e929fb0e6a5c0d6c822f35c401f7b602d1df5
zf220720d4612b0785594ebbf4a4df2d795b279c5a9225fcb656e4c865468aad0282918a06e9caa
z0f07ec5ed7685c58cf5edfebcc63fc03d617831b612a69ba15f7bdb1ebadc93e84ae5e402aec96
zea52fdc4af04886e6dc088785f324f5065630ed185fef01f59c903c4f885e2b3589e3f72f91aeb
z629f78aed5b038e03d60959facb806967039cf911366713bbb5147895a7b78bf3715919aca5223
zafc012b7ccab9f09d8ea3a420ef6aa395a2d6651d2979a7928ced59fb3153a83e04dcf22a0dc4a
za31f2051e39d6c02cbc9f76f5fd470663c90af3550cc5a601ac0200dd4f45ef0626b30aa3b75d6
zc3b4ed3085841d95fd2241088be37771712fd1db68bcac7af1f7778dbc4aef0d360569891cbf90
z067a5cde1bca2c085741ff83880cb614c57f7c129cbcfac2c794a7f9464153047ed356641ccc8a
z4174bfc96d13fb5d7c460008d6d27387b781fe57b6b323560c42bcb53e4c386f7982c81f79e640
z7f4fc246d36aa46570f8f309ecf208a98c21ed41fc3bcff0efa76104073c80112b3b40eaf55ea3
z923fba58650950c5c7f65567c2bbdda29c71de435f2382d32994e7b561beb545ae638f282cf129
z438a0b57d3cddd7a891c7d16e461991bff037e4b7e599e424275a9f015997db43c4123d9f0c06f
z130351ef37eca3f2d346bce1f1b5541419ebd8a4884b29dc5d39b5a87c25fd46a7984e888e4cd1
z4fc2bdf10d332dab224aa6b4ed093e4f84184759d6e70bc22ca8072100b60bb9027abf3003423e
z5e85bfb17c774f7470e54824653123ddf3a47f1d481d3e2e8bf98a758466d1ad1a8e0785844160
zd607113e3bcbf78f386649752abfc94e8bd5dc9a0eba798268d2fbfa9bdd9db5dfadfb59242c13
za95dff1aac08ad78b310f5e043561fa63bf1b4380b4c4073d812363664d1bcc039fbb925be3049
zc4f22db225bdef50c7100270d690cd0573bfcd6345ab3a1bd57c507f6db48e232f3320edb61de5
z78bfc27e841569da6adc921a3553b5f7c46aea2efa95887fa6c24932227828495a95e56ae6852a
z3211a4b815edb32b2756c24f670590711a78d1a3530d1ffb2ee258584c1cc95755cac7085fa72f
zce0c4e50d9f7942d97b1bb71b36a5589900e24491ce97a08bd4569c01ef088258531329dd19ea5
za9745a70b8e890be34c9c360f393ea6af3717afa823ce9861dc99cdaa6a740d7d6026e48188a03
z779be728c2db4c5ebbc8fc7f97c5904863eaaf9cea373dedf0f1d245b9d43e23b64ba8f240498b
za1a86bb1b3a71078b5f754e58abd3a78693f8cf3a91210bf8bb100bf8862bce8e8e8015899f2db
z6bd35e78d7f9e7010c47a3227c45bda5f22c4640917d6712f650e590e449fd9b2547b8bee8fc71
z84f2d6af613f6483a0d7242631e25f3cc7486beb263e5268b2f1b2fa970c0e1694854c7fe8c8e0
zce66f27bb87f20345f289c552ec127b79e133764ce676cfe67539c42af26d7cb5c3cdbf3466e2a
z27f6fbedb09606602982d85226449c74dc0601d4e17ad9d1f6ddc232ee08b2eb643ac6d69283ea
z7439a678aa494303b61c30b043f0438de01daba9f1dff52a16184a667b9e7ec0c7585d6a2faa80
z960fdca62e9572bdc23db3aa922da0ca959d2b3724fbab840984221a18c58ff786cf137e2eb143
z02784927959c10d423e2bd99e0ef0bd55b0e5f12ab28418ef733a939c83e920fa65513aeb415af
z5736aff30b41e645e905b8ce221b4bda10e4bc4a38bdb1da9328cee9b3dbac67ae9aafd4e7e800
z683c172199aefcc8eaf1e0fc4f2f51053608bdb6856b7023c637b0870267a75b54f018b40ed2f1
z44b95b2d1deff01bb26bc623e4561801217603c11fafbbc133b0614a1d99fc252dbf6af66fb070
zed6f95739873a6cde7c4380ca3879b4e2822b99698bd3a9e7d01aaf993bd9b8fc59f34b07b49c3
z2e904497cfcc637b8a500d34d929746052b07119fd1e26807d60c87d6e43ec7ba0abae750d974b
zde73e97154803f4d51319b2e9fc97592f9fbfaeb27529fdee06beb3e1b829806e11f3fbb832d1f
ze20ebadd3938f0cc7275ae9ec46e91370861da6cdfa7b697f9b9d04ba737fd0fb6776d44a79dce
za42f7b7a7d6c1329f7d1f640c82bb4923b72936abe0d1a891cb2cef668b1d0d1d7e3f7978155a4
z024caa69678b4b107ff7ab2a5bd00a050747b559a2ba32a4de0731a8d2d9da62fe45f1c360bf38
zb671251b1d3cd826ac0b0e7a9584a42ea008481b38ead2bda9f263a960dfedb3e382df52243b5b
z70f1da0dda657bb9d578288b7002f9aea13f873a9b2c15651a02bef21c19e24c4b0bfab3b75b14
zc7daf08072757b77bb3245fc1051d7b4c08330b309e3390bcd0c07dd07d9854dcb5fb3e73f52e0
z2737ffa9cab04b37c3e7fa9ca8f6612b187941156a5f51331067c245f5fcd2d68d3c20d79af2e3
z887a08675c972ea7392060d830aa953906708677b816775a80d8f4e755cbd18a5733be041d4ecb
z2410a847f7e241722091fe52ef0060563c2276516288cccea6904dc48492d3700fd032d3cf9949
z093898d7bb044e543bce748f72a080bcee6936422e1272f56791bb019aa28749f68694d525d2c4
z37f62d745676415682047dcf7cdd79d61747f55fdb5e995a101f254011d00f020f684fb8e6505b
z7b6784a1e070022ac658018f457f7ef0edd5f4c5fe707215288e26342b3873fdb706dc2c294deb
z0b47b8cdc829cdce46461c92f29e99852d80d7f35df4737f0a8fb3980e21108245cdbaa9f82035
z8ac4d9323321a5dc2c4a0583b034d1e2fe720e671584164e2565df822f4c4914df3eea1abf28c6
zfe2c2a482f4c08af780a7b13e9f018e5da5149e56d587ba5bafff076b20e21186f0872bf8bbd42
z0989c2024834ef2b2bf785f8583e4e05ae4b7099829f8ed14d189989330d1cb243be21fbf9aa20
zdd12bc351693477b56e96152108a36095d87dd22bd1dbf352d7a9af0b009e916962f9d965aa6f3
z1f3e67948dad494f6572182d6bdcb25d9897fd120b7579764d6ec9a68762deeccc094f361424d6
z52611e3fad56edc266fe9a4ede83a70c43eacc8ae1aca50a20c2c6dea3b83c96f25415df5b13d6
z3890cc8c34be2c9d7dabfbf38d916e77a7a3d904bbd430077969a45dd3d849fa9a985eab1cc7bf
z57bbbea30ef5e922df6bcba8f05daae9f5d7aca54757501757c3969694d0a3a724ce637a6f0ef2
z19a1d1ab88361910059a002fdcf2f09a3be9e8f55879eda33d506b9ec2892489e3ad10cfeda0b1
z59808f9685d3c8ea8caa63ec4584fb07075d391a5979e3306198209b8cec29b5790a6264685a2b
zcebd48e10dcb1c1c09a1a1291971f778161c1687116c54f07d9eaeaffefaa54e37a2803d095360
z46b448d769ddd47a99b56ce23b5aa8847a8202e31b70b2b060c3ca3fce501a6acc1af9bf1ad788
zb9bf768f34da5ab01e64aa9a3cf50680d81e76a7816bb842094a1083a088b6e370cc9f0852fe88
za12a977917bea90da608891f0e6da1c28bb09c76f178037ea16e822964922f3a12d5ff6306f105
z3b86237efd65be5508675d256434aa01f4b7fe7b4f7b2cafb7cbb37d8f93f654ed226abb2a5fa9
zb143135a5f4cc7a11786dcb14f1e2f884fd36d88b68d37ca6376f5d5b651212bcb14da34a98974
z2bbccca0286acd80157836f8b161f2d47b40ffc2aec19dca16de3afcae9c6491bc0af6c5b01dea
z9142dd3e9fd49f24ce958ce306bb0c0c283147797842051c492d7f084be04b61eaa01bbb954f63
zbbc0f976d4771eef5a679de19831e44cab2549905a8593c83a8d9b3ef18cb739b83c2b0d7403cd
z4274c82d075c161bc50614bbe134ff9c39795791f8b9ecddd0a276dbac14491a66e5e5e53d6b04
z86ba979fd78e4b7374232e29acf71bc74398008cd8f6ee50f345ca08388997e36de9e39fa14f30
z557a5b2895c4047a112de55644d37a9934c8f06bb9ed22a91f768c89177b759d19a1e682bf7481
z38feb74beec32b63b6e2d357b2c9776c83383014290af9509a8556b5a922f5e70c05e219d1764b
z3cf535cab315696e79df7c37cb54c4795a164fb67fdf07815cd3982dd629476a26c3f083915ef4
z2f37dafa977b41c6dc8f49824f7b8faf0f2c4190786ad0e035bc3bec6b67958acacdb2ca430b4b
z9deaae52ed41253a2cb5eaa1abcf1e945a67929e4ffa5ab6e17993cd70d7e203d9fca997f5c3c8
z88a51b3bf400d5bd36f03133530fa38fad4f9be7352719e5c7a6460defe017606b8453db4e4a1b
zfe84f79fbd41bc22708b79b3de00e534c4765da79c095d1d36302377657cd2eb163f94e998d193
ze829a0a9444f68e82c42b383126f646ca7ecd02dcc2eb4be54d68e2db4388b8b94dc7a11956473
zfca52cc7355078c4b2e8ca410d5060226462ab8dbeae2a2e19514248bd360582a9c323e710e94f
z326e23cdd24eafb8d57a17a6a41e2ee2a795fc022fbac019d5a4b970b82350865755152ac45aa7
z835fd3a44cd98e1150af7ca366a64ef985da8ce782f605877580b4a25ba5a10ebf775983dd496c
zfdd8e81717c9574c4efbe4af6ac5f573c700955e70cd504bdb4ab2c36f8a6baf1fa6041c212c4d
zb07bb0f60a85c79fe7652a64d8eabad119e921f08a851a8b1f9dbbf4e4edae2eb7c0652d34489e
z51bcadfd2637800400af2e76999dd83f33d5bbe56e12db82c739740bbdfd01050205078dab459e
zc14bf04e202e4fd7acaad753ea7cde844a9851407913384140e748c39668d8f7de742538769330
zf67e4ac0909cdbb4ac3967a5d67d7b9ade5000c8294a0fd48df6cd8cc69bf9a3048af97fe69bf6
z11bb33cbb09c9c321d1882ab1614d60a17b00f92b56eb019157bc4d292f42477f6f0bfc2d5a859
z0b767be416fb36819972b1d9c7b935a8fc6179d0228d7c7ff62ea3717e49206df7695bfb589350
z53682e1c0caec4953045887d51b483abf40c0776cc6f03bba7f4d31763eebc109c0c2bfb73347d
z5a4a6a8b492ed385998ad2d9ff03d47164d4ee74ec55b4aeec087c42f7c62bf3f7cb4ebbfff271
z3bafdd13dba21c42e3da6a20295fe0c0d44dbf065db996dcf27895c5838b09d00685ccc5efa891
zdd718814f9269fe12c4795702b9873025a33ca1da3cf8cd22ddf6b85be57259cf9249242da8d06
z2bf80fe55054d802d19b5c77472c3b5e408e20279223eef56e9a7d282390a07bdd1f73f580e10b
zade1a1f7a21f433e95740f6dbf12a6ca29f320b52d0d9435d32646cf58bd32878299043938cffe
zd689e18890766d4bdd5c482132770f9927cd7bf36a999c3bc727b680dbd107babbf5d63cfe17dd
z7a267d14a5d75db684097fe139777020727b20eccccf7b498dc82564e3bd7c084810e4774bb21b
zc019ff58f9110c18fd82474cce53b74242d8d8cc6e3e73fdfcebfb9db16d6df5b3a2ceb668930b
z71068fc1b36fae560d40299f7abc9eec474a33084998b036fbe0775c3707a7c52692dcc6838fdf
z360e95de144c7f98b922fca04ca617ef98dfe0fffcf97883e6c1b7f9cd400a07c83d1bf61cb567
z53a57494890507de48d1af2769cb2852864638979e280dd66e39f0eff4aa3622f635aa1c46183f
z10140778dfb1262c5fa8ed59caf6de259d5db3394d9b884c661c23bea67e243b447bc634ef54c9
z9d730dd179750f443ada54df30b236ea60a6da9275fa55aa64567a20b899750e49eec18a062635
z04f8e7ce9d8c8e04cf04956de4c01fd863dc9e99494831851f82aaf81ede4e0fc191575c7691f2
z2639b454dced128ffbd2aa8c7ede6cfd8c334a2ebfb67fcc45121be94d245aee96a2718d2a02d4
z6e2b45778d8ebace6ff9085e6c0cfb5e759284b86058f5430c3ddfaa3f3c0e7c6500c995b2e790
ze07520624ece75f2456f9d32949987ddf4180faf868e3ed6aebf7cf26a65711f8eb0fcbf36e37a
zef72331bd6491d6ad55e2dd2d81a3d9952d0ad2fc92bc0884563a9d8c6298480bf84c7c9ecd754
zebfb21e6064678cc538078dcd84a24ba83de8741291132fa9e532dcaec7a532707489bf51688b8
z7c5a83432d8a170689b33e6e476b1507e3863a0972c08eab29f967584c30e31485d6f875e6c664
z3f28f5a9e866dc6af76804d3c9a7fd032cf69cb0a87001d93094396d5615cafca87c5214a16c3a
zcf58bf48df06a1ca69dff0751b2c6c2fa4f867d7c5ed9b901bf98bcded4e87332ff3d6873ab255
z73bf03fbbba3a9b23350fbf9b05907294872af2678c4268504c3bf9dbfc892fdc845468a197b39
z21f9c8116cb4240784ede9320b533843c5921a6f6b1a34837d6a58e0d4ba9e3f6d72174cca3e26
z925d0a69d607662ecf7b7f11aa834174e1612dd92149711bb7a6f93b957cbff2a1eb873b6dc476
zb26357dd44628e9621db83043b9312ebe1f313b9cd815c532b88ce3a163118f29ae703d2e02023
z8f349b5cdf89eb3a381de1a873c44149a8c47934c418ca99c326ce127f5711422ac1909bc1c7b5
zf06af230f54ae120fa0a4ed79d370b53f09d60042b1d4a53b7d8c6bd0701fd61eb051450e01d54
z9499bb7119e3ffbf7dc5c86dfdf0e30520bb7730b8380095fb3eb4008d7a6bf10df7a66e0375d2
z6a73805a6090b62c4f7ddf766661ede0025e7fe739360b9e726724e95c2c9975cd363fcb09c0b4
zb310356ab6da8781aa459f21536dc330c44c33a2431a230fe360f43aee081a7c65074bfb8afcf9
zf6b74f81898af5a46a4541d874662611863c92ff7ced26990dc59ed73016dff2e837d84b6dee19
z2588437f81a9b2359509e3d338f5d87415bbf9b99bb5f9f27b9bd749714138e5e4e104e2777af8
z7641d9160eb160b83048bd609671cb2d609df1a045f5b06b238768a207945bf0fda6b6e8453327
z401165654472f2ab0e67b30b147a6130e6292e4119fb208fe014afbda4e258faae3f444484936a
z757e38a100332e01727b9554e8225d305c3195d201ba070c8535d8b6e21ffdac1edf74273c8001
z527dd28aebb06e95b3af92430e29a502ad1a90c71957ed2c89b85c0e6c2ddab7c5654455c46190
zf2ae73de1cf14b2d121b6ecdebdfd34a0e88182b7c2b0e7818a64c9620bf4abbcff3279aa3a4ce
z4374d2210c6abf9865d69f5592ee70be60c5b6efa3344a3a58e7da37cc4d1147f8266f9f97d62a
z03b961eafaa01771fad7353e4095bc94c9857a43bf3ef5f9298bdee4bda62e400390c549f3b52b
z3bdee350dcb627fece24c51be3ac2bbdd296d1201ad06c8368730db599d1d414e5fbde3373d12d
z5047e40b17484db5645d59c8fc0d9be4e1dbdf849ae0f4e90632d2a8a218d71a2a400fb241939a
z18d583bce46500adf2725e4ddeb6fd60f54e06f54afbb70d6ead75d004ff9234442b7b2f083b9b
z2cbb0d5c4abecf8cb3c813670ab48d3fbfb711a7c58fc74dd4c1d5a65b3b25ac21b8410bec0122
z2c9fb78de8e8fa4874162ecf71cd6da6fe0e7fc2edb0c62894bfb5f2ae353361d51ac73596d20c
z6e60214c62c777f6dedbdc02d1cb6d3983f6523a3269f5ad5a5a3539ff8dc726e2694f2a3249e6
zfb3f2cbfb24dbf0b6532669a538afbb181c06e80699717ecac8c33657ce9b9b52f3e8ee5822f05
zfb52270b27b1fca1203f5e8f6d96098e438b5a27bcff8554ef2652a339249d07e845c6e58d4524
za85a96ce3006da6d9d513b2187a737f42e97d9cb8b08f52ae880937bfc1821690705510cc50f8b
zf73ca6f996ce798f76dacbe129782c5cef53e488847847aaaef62528be5d05a70d98a3490d5995
zaf06300775625325662958d0a4e882a652694c58c26b2a40a7fff5fd1961887ff8e11b42db91a8
z7d5e46da1c846467c8b90f590d0b6147bb4226a8e36e6377164e134eddecc2fffa276a213b8306
zd948ce17c2c25f68465fb395d9df8dd590e3083914de8a795e0af543b9d3d4a3d1130aa468b950
z9cc6a94f0c4e3abd6b0ba26fa68182fcc68b64b73da3949b21e6a62c9303745a432c8f59251000
zf05931a9ef97f3d41ec1c2c847095784eb2db6b341e16846a3580eb1e1d2bd0a1734ce054d23a3
zb68784e8744adaf297807eada750bd970d434cdb0cad32cf62bf1a05ee80adb4412a738243c9ea
zdac7b9e27bc675a2ba1abcd53b06df1e783413193368320c0ffa4c36b1f21d442c2b5d15e55c05
zb5637f1d4c12022c4c189d5dbf58fbdebd00ab6c5754704f88f6d9b78edd2c6624cc13db02d87d
z031f942cf4aa23cc90e6853d0db99417c37359cbdf562a01b75b9dbc91fa0012362ccb840e867b
z4318e9ad9cb6339a4bf7890e78f2feaa20aa4e921ea8c641fc65e7eb85f2d82b1fa3bf983c0299
ze9bdeb9e9fb8bf65594054d5cc38c45da4eed878b1ca8e6094e9001893ebecb35c00a640b4cf5b
zc9db0d4701b0231b5b2e3bf25625159f4c3bd35e934bb17d178f27b29cf0d636c5cc2b20421079
zef64710cb794423c04f0026942e086e0e77e22302f3a69f77f42ff8af89e98c1cf393442229b85
z613acc1278d55397f53f110896c25cb6c270482869fb615981d9c6cc2411722a90febc9585b089
z7062064184df7ac07357686689a0d71a040f82a8bf2c30e39fa205501e82cc2ec66e072bf828f8
z4c71b1b328fa1c5cf86275d5dc40a942d51ab1eb6f57aaa68517ace524628f374f70cd890e3d3a
za5edab03768f3033519248602b64a21debbbf0daf657d66249e0fea49a2e75bcefe738c64693b8
z056040349a9023b488297bf6512a9bacb9c5542280da29bd65db0a7d7b2fe18f88604d170f2797
z6446ea3aa3f652da5b143ad648f0d9968de11009d591f640fa3afe4a238b928eb0365415657946
z18ddc72078e792450c628f8056a7dd61c2f13b03fea06b99e739995fb5898101cd20cb5d07d2b1
z7f854dc996b7848294dc6367af6a462c730b68858491a2aab778ada4a693ce385b01546d6bf559
z8872bf1196e5d858caa0183aa104f6fb309abb1107909d5f973e721fa6a546b7d7198e877acd0d
z4152a8e99d6b617f3d454cfee5ca54514c2348d034bdab5bd65520b3384f855196bedb2bb5e178
zf08dac47cdd2226251f330687850b906b7ea475234649eaeb088448cd9069b19c1dbb53be90ef8
z0d9ec44b5614355d3db82475fd4a25f7fd301907e360fb5241149b8060435d7a6d0ad5088bf521
zb70eea2738edf85af07a3aabd73743ec0bc2f45c7be5dd2c35a4a54b743291fee6559de7fbb49b
z67e9a2459d852e0f27925c5c50a3a36d63f104490140b9315b03f8eafaa833d971ea86367bd23b
zb7d6513fce63f8791c8ba9119970f15c16dc70196a431d3a33ba478ef801c164737acf95177da3
z13f199041e2113f61b7542fff452ed98beed420bc1230a80bafcbcb55e139aa89f73dbc2c6d3dc
z8306a4de2e0193992e6de434d673a762fe72fd8ad695f3dc3a2098f39a3a7e8b8db6a2b9460cc2
zd4c831e28e5adf6d3ef2f0ef6d2b3fa4a29487edd56de665f4439b8be7854c9e71b7b13aba9567
z8c797a7397aebb66be4e534296c5d7bfdefc7062d18fb255512b16706d67dde11dcccea8c7f884
zc3206e914909db7482a525568a3429f8928b66e232b1dfa53ce14422b7b3914e876b057b911a15
zcf2e6037fb6ff8c3dae3fc3d9970634961f638a7dfc4d71b8bdcb5b86b81d9aa4dca6785119d0f
z1315801c86e3e3884166e5c998abf03f897d18bdcacc51363a8beba5d5bcc4d0cd165922a2fb5d
zb174c6642712f5321037cc440a8584e407d347118d3c861386cab893f3e41f05d405c4466ff71f
z23967c965611f83cdbcc0142a7e270f3d418555132e690f8cfe79d7fbb951fb2ba61cd5f20bfe0
zdb3ec80fa1e361db472b518881e7089fc7670a97f4ec3a45f6d014482425fa5be586357b661424
z201e0d5c9dd6c720fa49319fd9f35b401ddb8de7886d7cd400f3dcc70817a5eae9aba5cb1f1b80
z952f906c0c53c9702b94f4cb98c1dc03146d62338ab8767b43db5af41e16b8d0641acceaacbeca
z6be9e026d157d313472b53a5651be655de29ca546addbdc1e5b46b6c6f811c2e41a8875c20ed8a
zda98f46ab439dd0d898b4d0246ff3ecb2d8a667d56ae0a2a0f37b9b08a8927de1d84ca564fb643
za6addebb03715d639ca24756eabf4517d604459201bcc46c00cb6b7cbc3690725236d940f382f2
z2f6afbd2c3ed0ee39eb2e59398ba1eff814b2b9f9d96eb4c5e58c1f64dfbdb3c07f068996cee8b
zd99958d7a58ab99a638e99fecaf2771868ebc3bfd55a76e53fcd75cc6c2212357dda8a919653b2
zebc63110fc9f25726e2d5a1f9e6927dc9f6ef3206e2e55711f874c27a71b1efb2150e2fb0bff38
zdebea37c5f7b3a664a93309b88b146713ab066af5661c6e9d9fda4fad0a9894b01a31531924584
z45f2ddd3a23b360983b3fe1d4f822a2d4a003e85c32a32f44fe7a3de770d4648573c4d4dd24dbb
zde72f74f92319535d9c06b8ca33f671d66a2f231a909de833f0fc2cac9cfcd5a1aa2018f64e4a3
za560bf1e3733b2d23644819ca4a167a3bffe03ab9e2d2d87aea6cd450615a99220f6d51e1548a9
zfcec02adb3ac5817741f9f9384b82fa2344e9c72bd17893b7464cad653ee9e91173764f7442578
ze82a05e4a70971f87d1ce5a523d9d7d4532711e92740e73d19ce07ff7873ff6da1e63dde95b477
z19dff64721cc6bbda7ea1284a916e9bdc7c6a551772331e61db3e90c6e2471c1256a07fa8a927d
zd0f4c5241caf16c6c3e833228a41a2e1b23101b5daa9512225df484c66917437142b12344161f1
zf12093b8cbaa22d848192e50409ebaec2953f6702896a80b48085c5530699c32f6ff8be4d916c6
ze0933cad78b56e8ec497f8a2ad053adf6c095510d216d5f63c6f72001ff0e45b43ae47733f9604
z0a83360bb94cd700c67e66e9a53b04244e03cb4e0a59ddc0427764040b0eb4de019d50dedb39d9
zddc8a451fc1083b402919c333f7f99f6ca89edcbf55a76dcee64e11e354199c8fd4098fb0afa54
za379bc2ea96c09c76e948828ad969d6ec7105d9b52e65f8d782591184898c0c78c89ec2da6c599
zacd3b488fc9068d99671a41805b732030c6b8541f882c8c63a2af48fcc8349e60e0f947c10e7b5
z508b2d15ed589fb1b207d9fa198c2a434c090742ec186fe20a0357ae06bb4349ca4f57ac1528e1
z36044a5a0652bdb6aace13ae06d9e50978e991032936ac3632ebab7c2e73075dc21305876b8bbb
ze35aea4bdcc11f40189add4bc7910b62fb2a95d64c1a5dec43fc2ef6f8eed9b16e1e6858cffe88
z6bddb61ffbf6a66ac80ff834e709c6464fefd871ca3bec3fe90ce8098c03a86b07b2b17aad72ae
zd11df9c8275bfa5b290d91e77165f465cfca8047c2f088e490cca89461ce27906f18dbb09afacc
zca9285c41750b7872fe57cd371bffc20f239cf040d455b7065f6b1f43ee98377231deab895f4ed
z79f5f6ecb1aff923645f5b1af7c060a8217433da6a9f63e897118aa0d46fc02db115ea4d5e6d54
ze5600aa7f5ce118795c6531b27d082b746d27a36d056602a61d4c587feaf43e0f956311a49cb4e
zefd02822b9082e2fe16ef24e38557061bfd8730c5c495ede6aa909391a8ba1765e38df369ac17d
zaf6134b0b84b5736f4e668390f4a4d46844b9e620b9a1c5313d10d872112a1de96ada7adc52f0e
zd4163127d90f3836295218022421b6f5139ffb77bb7f5074ebb62d2d13982044f6ae06685dd516
z24b2f969ab72bcd9e033a25c4178df0ae71306ab7b02f4f95b14a494512c214459c32bef072952
z54e02971048819bb5ca10378d11ffcf0825faef9ee54426f5e657b6e9edac3c32434471be3e594
z4f7ce9b9938b36962da00f6304dca109f036dd7689c5f07ba89487bccf54ece2c49e12d3626988
z0ce181e043abffffbc162ebeb10159c989806b5f70561d5d84a8ad5a5453f5585a633fb76fcf75
z9c876181e1cb929dac2d06457070f034a34b8c8f0556448516cd3364d92b781d2cdb088168886c
z68b3663a89c5bee09110361a8952e475f5a43eb2d6ff920131645aabe425be45193cd8f731a246
zeaed834a3ededcecc705ab77028f0436244f4f1e80f589ac4f97fad7e3628b3ec66d5a69c33245
z96211a56349ba51129cee7dd780ceb171088ca4cb10940212cd1d2156591cbaa7b276526ffeddd
z4d6ed53f7f9d4f3f680100aa6fe93a9a973c2b90a3e87b173bad121a206dd66fb8b7bcb0f80a4f
z437a5ab770afd9f1eee5983354e1aeb9757151a0a202780bd710687aa24da4db4fcb838436932f
z684258cddb29e00628885de01d3da066faa9b5d5c009ac9119eaf505411776b4887424485086cd
ze3fefab854fa0691178069e0a7276954651306473600d6783a624939bdc4595c89136b251b19b2
zb6ab62efdbc147fc2edc158774be4586fc2457bc816b1ac9cd202e9a4aa1b46844cb942b66627c
z565b2a9b0afe3dacf8d483b0582c26f568573ce77c492fc35b5d39df5bff9edc83e9aca88890bc
z9dd79b43d8b9cbf48e90c4950ccc697f22d8249735252d2cfe9d3934a1bca686031c36caca7227
z8f699ae3929c63220b6ab6ecfb40b26f64266982e63359893ad1ff25dc80c82c58a3f5a9ad3332
zb0a9a7d955279a640236fad7ebd426a071c34901124bf3cd483a1b7aed60d28eb4faa35aaff564
zc90b85847ca846b2a643ed941254b2581f45e04e35b6d04f72db9c0b1375a02b79884e2b2e055e
z9351fc2b5c97df7319d65d30653fa5cbddf789ec4f83974406965f7204e561971f113f69908f9b
z1e864ea9e107d1c7decda2904eaa2b3cfe27225f323c48354365789e4c698cf55080d4124edeef
z30a1275a81255dc82ae1f88ebf78ecd13343432cd03cce3d770487b3c4312cfa60676b56525013
z637e4d2e4e4dda5ce64fc244e2be853ce00c35c62160ad094584bafe8b5de3a3b8e46af0f77caa
z6c98c7fe46bb5ac0f689dcc92c59a17effff14ff49cc778e56545d3976200b4eae77383e35dc8a
zd642f7570af24c4b56bd21d7f5aeb22eceb5cfd7e321e62223e8ca724aa4d48672bf89cd62d8c1
z63794a1a7356d687a97d75e0a1668755e693a1e5e806a69bc13e967fc87c8e750dc42dab4f5b1c
z54183f29209a6a814bb3705dce9e33738271b7417bccc3dcc5c7fa8ef32dd92b589ed10ff79d12
z714f8f0f54dfd8058142141db57716110aa4230aeb79313af2be1a967c8a7c137a2379e3ca3d72
z60858a7546103eac48f19b0fce017bcf0c04e2210d3e2123003b00ba61b15b5fd32f4b77f6b101
z3d02e20eb0db44d387fefadcb50437cefef7be8a8bff24fe18d6621127451445851ba33f38a41e
zf9aad6d2d0ceaacfa712ff1d07bf28d3470180e93e0a8f5e26d928e6c1d164a705404d1d860873
z59aad02a1bde0896230506cb050065b40849164813fedd08e46d3fac5c790c13bfc1cd38d32a77
z417b677f3bdb3981f97968d2b4ff0efaf91b3caa29cd697b678fc8c5369a87a61f8eccfc42dd65
za40a798fb2cd051993f0f53ac1646a276c034ea36b1d5da857c307275302dfa61a7ca82722a0b0
z77d8221ce5194b19b7bb6a3353fdbadd6687d5590ddb7e6bcae8312cc714d4e33423da2837f240
z5d6093c53de2763fbe47491c8e8adb841dbaac5f05d70ff7670f0e4024e5293549c00f88b1ff65
z06a1c35d20a2d6466341dbfde727be80b0e0d0ed76fbd2b08d3d5c508f0245d8274ec8969c0755
z8f10e9822e5511a70dee9d0ba07d7d395f50f309a294c47cafe27c81e3191b611f60d90d18e45f
zb5b46ab6089142a15de005261aaeb66b7c2bd201d97d3a20bb1887bb20e9a7aaea69dc49a608f5
z571aff19e9fecd0320295fe6a660e69946d5879904559c5298a63446b2dac1209b0c50931a8527
z9e3b231c0e1eca4de8311e5b902b376d553f793399906d6f23a5aae2d6dd776835a8fe8a0fdc59
za93f04b4d36c2638b194da917871c7e36b6c4956261edd8b0675539cdf3c29c85efa7676e3bb58
z0d31bd71aa6d70ba9425ae2df62a8c62c705dd0305803acf727fe56a66b5d592c34f24cfef360d
z1fdfe0f25d1ab9f6c48872f6702de463b5d810a38285da4eb5ad87bb92f413fbbcf36fda51e2b8
z5892e2de6cec9c5601df8e3819ee3e7e4d885b45b32111c5f5b3cb2e2cc2bca6e32e1a6ef0fcb7
z3b3727b72f84422dfbce6ada2c066904f897d54985b73c434149092d2b4b12ca61d7ef7c8dc964
ze288727c1561240390e029a8843c788e81780045461317925ba13ebc676c222f47d292a7927d43
zf92f2ec6de9f87928cbba06c4dc5a736ff3b115ce1de0931833b21661550d2a826519ca1de3948
z9116b77f11ed459a69989c4a5da805817fe3d6c1ac6889dd8e14904c6ccd2fc448be48848967ab
zf9c405d754e8462867bd4ae91265b4e4148168607571be063d725eb41831fbf30ee9d0a3850e3f
zf5e89de21f79be3e9ca41139d7cbcb0783cfd0be127ec80c3c8fb08af77c7925fdda61f2098df5
z637b53094c840cd7043a5e2945c325c8dad6041cf954fff501b67478fbbbac3dd2e9a239132704
z2f5fb7d8f556fa5fd6262fc631478c37d2c5c7b4f98f5a0c0684c37a09bdc8a357886e1cbf0f2b
zbec8fa6ed4fa8f243282a5f0fe79effdd546537855040b923f3dff8256300934b39adbb53f0556
ze249d7a072693ca4b05581921622844e3cb01346acbc1e6f0b4c59afa7bbb202c4892b657bdd10
z37ab7db59d01c61e6f6bf74cc02f75fdf1c72b61fe7e2503d427d723cba280b9d933c88938e505
za9981991072a945224bd38b8f0e8476e95f6beaf54eceb0456ec693e35aacbae16a70513e613b2
z803030c684a70168abfdc53622fef05895937c5e7fc40e260b39737535cb28e575ab3c9537e62d
z84730db6f344b2b24d96b3e013699a62f6073e7d64de1bc92aed6e64002a4c8d9b66d716de9fd7
z554163979a0b36958515dbb8e5ca08ce1d31359efd12410c35aea9430945943bc929f882c5afc5
z8b5866101b5e660c33d031d5942b26ebe7148ade7bc791e22a586d17db61c43a379e06573cea25
zb9e0ca624097bcbee9a8a9427a8efb0a89abe99e98c9dca4d5721e3045af7255000234e63f3cb6
z4431a8334375369408dd931e2948f367304c90dc128a668971603742cd60dc8e3fd22670e8be9b
z68015e14285d899a0f5c717e0418eb80cd51ef268a3ef1bd11b522494898591718a98717ffc041
z10d6b6908cb1dde082b6acbd481d126f5537b4f09f4c25b268360b064d00596a16151ba266f7e6
za0a405856c5ad251fd1787070134c22eac2c07d45918a4e5239be7017f35145f8bb09b043f6d78
z86810683fd92a5bf9f09eb109f392259faefd19067af9c672ae19d5c47239fe8f49151edb28705
z44ad0d1ac003cf0ab94ec34e99690adaa6b650ef54e8883d1cd867558bce602cd8416da4682a7c
zbff9aea22221be5e0c6cbcd13ac275f26caeca5dd3fc36da45a0c245cf7d2fc14f7a3e5513aa51
zfa8b0c0ffd1639cf9160a4b33b51c483a232f4268e9b41919b72d0069a1efc0caae7e01a0f5078
z0e70c427b5c88cabad22770317d41e46058738ad21d0e7ab05b44310751b1cd06773f0dd6fe232
z325382b0f68995a40e0a041ac48fcc17f2e87b2b8a78be9ce082880c4fca074471592079ac9a21
z8d0fbf9a2bcaa017e2da8f190fd4f7e7b9d678fd796e533a3a5ad8350e2289443db11838919168
zbe1191c697168cec09193953c787b8cda5ef67ba2b2dcc5966cf4078d302e5a37e4731940cdde3
za5fcec54e0d0ea5723f4089ebbcad3561d8a55da8a77cd39e7dec86fbf9dc2cd1c8b385edb4400
zb975e096cfee035de94ba9eb305b72aa2736f45e43264abf66967b9702d65119e29146051001e2
z1025ca960d646275ab11ce586a7b2fdfaa725d41cd409593e41eb661c0c0be0b093e02f2b96cc3
zd19eeccb4b7a57537c3fd4a3790678cf54158f29286e9673e1f8164c5c8e85c8bbe966af560d9c
z7427c2c7111bb3f534aa5ad161de722976b6a50fa9da398f08c26d639fb1844422121cac118bfa
z15fc675d205feefc1ef0c7c8b6ef5d88506c6aca64b1d12d965ae4eef33892e8662e85a25b04ab
z90adf127781a00d07b26b7987b0aa7c33f23fc354df2da38cc9105969f1f83b3d9f098b6ba4552
z45f92f6768848a167909d90e3f153264e85228f4e9580aaffecc4b339d2ce4888d0d28d343fa16
z7f5d586011753f6afc15ef103676d859339a414a1bd9a1657c8b10353260700101bb975404bd0c
z653f8dc9b9fe4637f6d4ec09581223d2c14bdb3412e1b1c28b26eb9c86fa23648d6d5475e898dd
z0a7234018d221fe5a6f9b670b41cc4d2654502ef37ff9e7290c914e37f382391173527a2b0928a
zfd959192d37193a39ab5898326de3db101542b4b3e9455f19a43c660e237f5063c51461038434f
za091d36404068eb3effd96930baf17b68b4d2e2aa3d046e4994ce764bc113c4c13f483d285d6bf
ze7f6de39280480d722a801a63b0e1c3a5cf3a27e9804e4becfd29e6b6e9acbe10bbabe32471897
z73a1b597e1621b4e49a70f185bbe787bcdc28b85d69a0ae7ed9f932fd53fcb7f41745de78a124d
z90e861375860c70fa94748508e097beb84641d776c25815894118addfbc3d38220e62ceffcf449
z43ac7780baeb40d8a9b13aea311f9bc5b0011da1cae1af6057d6d6294b3fc67acd3008e2d916e2
z9a459e31336be146dee90c0d564fbcfabffcca76e16555831d034940532edd6204680672a2b743
z153bc83618d28068d1edcdb5562a1cc3b9d996fee70f406ab2b42399d222b87327593fe4c49d1b
z6f3658dc08869a1bdc2accf3e720095b5dd298060320fab6ba5fd0eb1c120f8283d65efd92d5f7
z3649ad866f8385cb859a4a6dd148116d2343b9c7124ef2bb5620963a5b26eec20c4978a8bbf9a5
zabba4dc394d54cb6a93d09ae914d8033b549ec5c0623fc457daab24c0257d540ad80460a3f9d04
z9d70cf28330ab9c2ac082feb7b47df006eea92b2eea28491470c72f163fe5b930224e8c6d78e58
z8c19675d4bb2cb434aa3a5e067e9bd7d576f24bc1a786a78fa1b0d5de87e28b040187e3280dfbf
za1e1d6ac912d02be9da5e107cd2d40e2e8cb9ccd7dd45e894407d04f1e8e3997a5fe210f8621fd
zdcb0f895126ec45b50dc398a2c7df62f29e9b48a7eadf078ed9ed084b1d43dcad467cfac3b3d9b
zca0d6523101233741c4ac1009e134db48bfdb84df464f58bca62ec25d04e6cd18b91723d94b243
z755298d8ea84cd1c2f3ba1b103d3c7ba28c8b96372c365e168594526f0f2cdc401ea1c1e85f931
z550fd24750bbdfd24519c625bc69eb0b3bfdfe09b65323ac114283e5782dbf10d99362c7e40b10
z346a6c57cb9ea02236ae16f0a36bd2196ab1e43f7722192461af41a15a31dfafcae2bb05d7d2ab
z33bb90e083bd83cbd83a39f1837a02aa78f2bb1016c8189307d0ca7993a0ff15b3b8dfd7895443
zf827e6ff4fe9c894dceb3da3a6a1ff60f63544d267a4385e30feebe3b72e3bbf2d6cf248a07df6
ze347d90cda01f7d04e7fe81d7d6071159f2962ca6ef6ed12bc2f0638e87e57c8ec55f7d64fe38d
z83ff1cf0b08e61984b59cbe0afa5e06b73e89f187424f550a85ebf1ba9b574d1363b37db98cce6
z499d6540e0759a14521cb969e9af81b182f976ca3816cec8c3aeeff976fe7753c4064f67f7df0b
z6b4d9413aaf34733283842e79d04ae939475044c4aa999f18251c3763925e5b57c7ce4cf3fca35
z6a651425616af2db51574ffadffdd1d0b3f340d9a34a73d5b83192772e5116b9bcf991e22b5719
ze5df153caf3a3ca4f5bbf396dd7b5dbbc655fa44bfe35f40807c4a6620d9348123f7173cd0b0b5
z1a41df687dc6e8b1d0e1ce9f78f78b7251165892ec0ae2a4291c7c8ae1bc2d9f5b3a69ce820471
zefaae3fb73d4a7a9a42759a3749b9dff92ea9c7996336960d3b6f1329e282f2a52ef5d05c12a38
zb5a9e205c66d4ba5d217e65007d75f4fbee5e20875f0cd92ee26b919dbb9ffde562ed59255363a
z7e7ca025bab05577346c2495dab64ad98d095a2a7f8b19e51c3f7ad721fb5b2edf2b1685953a04
z3be6b18b645e99d3df9f2440ff69cedfc526fc29ab0d384c6a06ef643136593200b170a72be071
zda6bb3d5f449fa78d4433c15978842719fe8e85cc73d10ec8b01919674b3c94e1e5458d907043a
zd5ef7206f4a1d56d6f35f8b1f486bc24f9f1f8fd445d9b3154d4038c41c297d61742f23922b5bb
zd64a2f02949c82c10dc4ccc60b56df8fb93b6d741fa90bbd4be16bbc5d34959db203fbbc4910ee
z9b7a88c8cf031896ff9e35221d4d2ad896ca978023c208c50bff27adddd183bf5231bf393235cc
z97f06932f1d3d59b3de1af3a01921a1e5e007e7bba876d8a63764a738a08968ea30d12648af0da
z02c6255e4820ea506d7a97e3448ad8ad0510d78e8a7179959fe5eea8c1a94f1dc3ec0f1f0ba30b
z1e4435c2e17ec30cfff82d78bf6cb4575eeb73db7acf3f5c8087c5599b89e578022bc5314835a7
zf7168ba35c786d8613041138679e0563a1e089ce759f89a86e87c0cd619ec6d9a3ce3109e24466
zfb3e5b553c2dadd6a6b3f3cf08b58e9151a5114b8a3e87a3d1011951016ee56dfb885b22a8ddba
zc715bec9c946e14aa0445db2325525fa5d6ccb906713379d63f7a374c496de3cfc6be02c0b6433
ze76cf32d14b0afcc3ce89c8169e6685cc657d9e13191cc3d9c3535a196ec68e7915c117f985153
z35071fba87bf8dcf313b295a89969f392f573a7a52ce3375dce5f6abda102f0992d4ba26109a01
z25e866b15ecadbeea22a18d4d794c1dd12f27e5e5de46b87bcadf47a46334b44c84cd6c0ce6b59
z83b55351d49092426f0ad6ee47caecd12a809dd8436eafb537e97c5b03ae034781c392661ec245
z1c8f4a52f85e7784ad62a01b2ea78f2170d2cce4b9332af438d9cad70257a5c34bb4e57b85fa4b
z291a33d30b228dfcaff6245b3cdc6ee86e668f805fdf66d34354cac570a75c60fdc30fde6b88f9
zba25b2f5ceaba47bf35c6514c8c0eb97e78495d84d1c75ea723f117a6bb3652c3a1f2e60e02191
z10584c0cbd6027e45e350caf1837c54863966972fb77fa436f57de4da6ba4f3770ca628f0f252a
z03be9f6b144054299986c7a5083f5bc4cc1f7eab7035d285eb511e86c112354a6cbb999277fa81
zc389bde75f14d963bf0551e3f36ce666f7b8a8d9924197019d1072f390300260c9104734683dd2
zd77ea6a3593fffaa6b3897f6400e3e0e0f8916c632c0d369e467920193374f8edc2312a7c58e9d
z0ed8ac822ea500513e8e8cf9620a1079db1f84710a1e306ff866c285e7132e786f09568683e059
zd2f8ce77f1f153eb5f1f3585c276ae85baa713f5f734808987d1acb577b289497c6d9d9cb78262
zbd62228ba3cedc1b81093f6cdf9b3fe975db09fc43eecd10814f4afbc4634a6a88887f3a9cf629
zb989b3a4964c31b3ac179a80b507e5ea1d0e988a05146aa22db9f0694efaa23c6b109d761107c4
z1e75ae108816612e8c3ba180ed9583de1d82cb1cc5e1f673d687f837c747e58e1ba1f9ec80192e
zd54808fe22f0bef2a6ff7fc443341f7b9b7d59bd74a2b7a50e9653586bd00588ecd35f1cc03c99
z7c323a2df1dc92538e563e0dc3811a86f522b4bfd4ca8a83cab0d44438571278805cb341b6d4c4
z97928b291dcf3adc1f72589fa4245977b6dd58d80e3b67adb6227d06f15048ad60d61edd3208f5
z284449800ffe4e9d107559d686aa8cd5b9a522a3084da54863d4276e1475a1f8d204022339d7fe
ze7d1480cddf56fd8a2a9ef0701c930bf9024e388e904db3142d7b43c812e1b4d4236db0e573f31
zd6ecbe8538955d926f990496b10a6a3ea72925fb0baf5d3bee8adf2f54dd99f52d46cb754c5c9b
z7e0c635cae6ed0ce12714df290e73013c58628cc6f566fbfe51cfd3e04f937d56ab1a9df0683a9
z993d872da56de1bb775681fbf5fc3a486b58fa8701c8ab27a981fb413bd6974319726e25d31675
z7b289365b64dcd85a3bfd3657acfc812cb72e9ee22c45e53e7ced5d14a9503822b001dcd9a5eea
z7ef6702f5f800e65518e642467f116d8fea966fb6250b520f6a94b1880b48a04c35127ad633214
z3ffaf9483ca640577e96a914c4859b1f62038c0e34677b6d79aab0ab20e324e9641aaf474b5b06
zbc4979edb5dabad9e5d46cb98ba0e183499300ab35f94cff649dcab88ca6d641466cc6ed2a58f4
za6831376ffdac4cfd74d01ea28bacb33e25e5247527ba770969076478c3a870e77e37429a2d60f
z030c1505d55c8ff1b7cb4212a1540ee3360046e35ebfca498dd3973ddc63340ea2a0af34d89ad3
z91abf2ae5ba0b306a61e1c4e3941927eb3ffdb27e6b9b9ea7b2badfa81d21926f6091ef473852f
z3bd1004c1fc610531b188a07c858826f9daa1d4624390d6cfdef6b14ecf636ed45afa86a52952c
zfd776541c0712bc069ca42efd58e11b7b3a41e231c14879ab1732e81ab3697231a5127d3157843
z9d54ed444e772cfc132abe8bbb22a8cdb3e45fa184fca396ec7ef921937916db1b42c5c215a35f
zcb7052330f955ee008ec339d2499c4477f187de9713ae5772466da2b79e6bdfb31e5209f210141
zf28a1a689e9cb82745aa91ecf0e1fcd7517045c8864e87b74c2cbfe9606d8e6e21bf62a740992e
zf158d463068ea3654fea6f4cb0ad79b007e8a06cdf774ea40a74f6e6d0d90a5381dd634cd99523
z6dfd5794a138abd19f7d4b8862871180402c0502699d6ab4479d47e7ff8c3e121559944719ee03
z554e3b76faa111878f06dcde5db4275b7bea5c548b4da54ff272de521730afa0bf509c1763770d
z0adb48d1ef1afe6856724607a87e8fa3726fc0f8c2eda4480633bf2d757f2630b2d10710871c65
z55ae9ffaefbc0e62f455e294c99ae1f4b492ecd0be9498103dc29dba971dcb90f748d6deb20504
z9b64eb024314be1f2cf6d4443cdc45bdc2ae072a52c16769bb4d842d1ca362a6bc490e1be54a54
z8419313ac667ad91bfefb7f4a9f5daf10024f0abe4a0a60110ff4bb9b1af39eea046b03d8c7571
z1f24ef22cc5a6925443e7a8b510b1c5a5b0816b53e47a1616b9876c2dd375868b3bc53c67e4819
z8677d6fa121724947c7abbab97ec073e93f070937c9eb5d0bac5a7aae15733d34d5aa446c36d1f
zda6c622b2a152189ed2417a2ee5d1ca18ff069124835eca0b08bb8ef406c947e70305af764eb86
z03422a807f1c3fba3ca827480d68f92a9d8e97a361a6db4be7e419f0c74b8895daf482789ace86
z5353c42a66e934a17129f893350cbbdce52d828ef754d97795922ba2175e8d921a47b5850f0f51
z8ae580f4895bd2a60b8e5d60fab72034c0ed360730a4cc50589c25fe5d8935c964512b1a222b79
z6e1deaebc32a515489de32e47678df3540d77fadb76a7cd411ad98aab067c421b4d7104784f9f1
z94ed0d3bfdab6d7222d969cd20a5f9c8eb335ca5950fdee03fa5492be5c5204c671258d53ece1c
z0601b256b03c520870460da15156812f20e3e227736b84d63c7f015d08155e26c923f23f8c3498
zcdeb737ac3e5849cd0281eb65bbe39082ac1d5f026ff422c2b8081b9d4e41f916302a648720c9a
z15135215e1e7d583b48867213913bb8d57ee3e21493cd199b8583a158890b8df8b1071d8159deb
z3067968fb25ca13d52baf46fa5a9be980b0a08c34e2f2c6e12afdd26d8c646a3636fe3db7ab88b
zd764d9d4ade4b9a42d206af0b8937559fce590fe9904f15b0c274c4349139cf40c9fd5a41ba521
z24c1fb03ac3da97e0071cf7cdf10930c42b6ca269ff624ed187e631733bc255f36960c24f646d2
z105a21bf11f1cf932834071544ceb9aa62ba341da78fec03600b900d28e6c5c5ec9f91c41316e4
zd9acf941bffc2c665491d651597384e4a0195156676d294afb9bd670032ad871f1d259717e6da2
z382bab3a61260870f485bfa6aed927d1dbd53344a88372cc98a6033dfa02809d6a3e076a83b06e
z64c76312d6865dd49a965e45c9c36c8e01ff0542bebdeda7a5f10dcbd6c8615216834b6ad800a4
ze350633378e4eae44437dc67b90f465c801c7025b46ae0fed260484deb8506859948741000f50f
z5d5f6ebe5937c1d38f673d93c804c74ddab40e36717cf8c569cbe50ae1b28bc0ed2027f82f0697
z736a8413f7eaf274149a25b7e330c8800a289a087e53f8ee0f1d2ed2a8a8b9e6fc4e44f9a225f3
zb08150a06cfe1df6dded8c7c3fcb7570f1d3cc33fe44cfb717d7f6eaa6cdff68a9d7214ddce766
zbf976e7309cf01c8339b24568aac8443e4fd90ad3fa2732b8287973d6ce7ba9995b2fd16abcae9
z53720584c1261d2d0f6ce512a50e386323771d59aa467012d09e01dcbc608686061885cb3becf6
z69fc9408d0b25e8afdaa50cd9b4c55549d7320528e968caac19965553c3a9869003fc446832c24
zb436d075c9bbe4178ad26b497384bf91bab205606e22f93db621c32daa83d1d06066c34fe9efc9
zf33135759866b41bf3d45e1b8c01213002c71171c56b8d7a2d765be7d0a50b3bb5ba4766f0d038
z75ea4a755a9931e154a0c2862aaa3605da54467f9207e4630f79935b03b66af0fe387ca9ddc115
z470dd63728e63dd6c39220f3b0f4cb9cfad1ac62934f4dba5c369c1e1a861305df9d73214f966c
z910c3a72fb1154131ddf94ab80d301476d1c74b3984e1645d1e7db4a262abf4a6806cb483e18f8
z92b79671b5ce8b491043af284d56dd6d2f23ca28723280613ace457f0cbd26df5886f3512050ce
zd2dbae1d77f5023ad1651f6b10ef6b5b16041ebb5246c77990cc3781813c63862ae69470b33806
zcf1de10f2fa9fb389571444cbce1d0ce3bec0e29c0db42d1991d5008b54f41a5d6267301cb4c8b
zf7d04d17101b6b7d6a346b91892ba81bd3659d6d638c11f0024b5f1cd68b330dbb78ce8584cce9
z33b65618012b1a35db2079437da47f357b15b74134b850ad46e33356155e945fbc17d0b46d47eb
zfbb914ff760cc59fbf4c53764a2f004edeef67b1bea408d6232d5d5a47d93222aa906c6671c59e
zaa4693ada870027cbe1332fbd1cf4cf3e9099dfed7f24927a4a1af544c77bd1ac773600bb7ae65
z1c212f9a5d4ab433866517fd6e96fe0376a35e84da04cc562e0e8f9cda7206c81a75b4be20d40c
z67ce6d4113b6a14cf1ca69ef9c08143c23fc52fea11e1c4c223cd3ab93ea009cc3130fb8e862c6
z459786eb9134cb772e72e933898ed64800331344ed66c1c85d8a91589b7e2a1f5e059068d8ffe3
zfcb33e37024cb05456b636e9e4c50b32ef499f405ef0f4024ff0e2a35456aa630b9a169c748151
za8bcf790c9a4518e3fd0779dc3b86b90e3db95cef92ff7c09243f06f8f8713ac729196584e0a07
zcd6da1add563da9dc971c57c91eb5c35c10897b63d53bb192730e05d34893e542ea90a01cbba27
z58aa6863fff3dff126f9a78fdced56d24c4ff702757e14a6c67e99e369701b3a6aba732422a828
za58570e650e824807f0f4c9da363a4fe3dbf5ac1a66077dff885e089e9374459a9d7086deb3ecc
z40b2bd4ef3e7579c9db9a706cebeb754584a89b7a7b932dd8df9e1269614d8c37328d039073ba0
z0017342bb021ba6c085f934a3dd6a077ce9f0bc46f25640e54199f92d93f79cf134d4eefd4474b
z810bce61a4853e5d207ca5fe3b8f498e31dc50ee64cfa2acb6187d18745e3fe4756267dd651cf9
za21789836a10e8776bd3ff322ef100459d7c2b4b494e4818164a2f9fc9278b4f256211fe43e468
z1d6599b05f20b1a725d2e41b093ce72ea4b7f2df56813dbf323e02ccad8f02fc5284367c3e95ce
zbbb4ef3bc76e4bdb96b182345fc66161d1e7f6c0040452d378e1298794ddbb3a3adab2bf1be05c
zb836b81e1b734f0cc0e25fa43dd7838aec7b094664cb0a1c3f5a81e2bc091d69fe1b580ddae66f
z9c62b84fd911fa1ad2f64b9b7c12a528d7c5cd5ce9348ecd2eb02fda75c19ffe8a6743bf2db2e6
z14ab0ecaf28b286ea4c6d9830ad9107303d00f9ae0610c12c4bde227a10980270b4c5478cb7dfc
z333e0240ef83e423484b54662bb646ec181c969bd466f7602f98f4add01c771fb354a321b1f928
za41fd9c3b26472c5c055d42566d1249c9f38e6c9c4b3147df9657f9f4eb96b2e4969485c40bddf
zecb4feb30e02ce1e86067ef1c6b91d5c2357f65f6fb3df8d04d87e828bc2e8301acddbbf2390ae
z7ce5449c17248abf0fcbe0de6f37242133d559eaf18e18efdd13a8c3c1c25d70533dc38975b92a
z73aa90e786758893cedf6858bd895e863ea0f981d0206a52cc818ce7194e95e585e273c97f3dca
za0387f1fd7595bac19feb228d25acaea0f75a04280c80f201c7e784f7ced1a937cda29d852b19e
z2a2b90631cb0b44b8aed2f81d47e96af9a1d7db3fc114902e3a66debe66fc85cfca04e65fffb63
z460bf8e884da05bf3135bebfd891aa338b1a64cf475e6f13548cc56840efcf8c028d8fc5363ca7
z9093e9715c361d6787ac0075ddebd45c2bb2d6c026dbc9140f6975d6b6073b9ffc50b0cc2dca24
zfc5de2b41b2b759652da204d030eedea828f8723c84ba13ee72309b90f1aa194198ce3adcde63c
zfbc227c4645323fffaade76552f47c6124e01413cf19036e17742a1c6ca3754d48c5d6ad0afd83
zaf9722b4631e717702b26e73721b6562ac091091538c649dbe859a994f814dd6e9570ce49ad95b
z8586e5ba999714570f6d1939295d8a7fe0b4ef5bee1757000491455a5487cd700089eb9f0682ff
z8ae38f8df8eabe77aa9a03878d078eea697b3b7d08c31970734076341d07a4e8349d0390f895ed
z6273944931b67eb3fc4abed85bd771f88fb977afb5ae089bdb705e728993868262bb7dc617d5d7
z3db5433c200ef590f622920dc1daca4184a17721528c4a1395a6eae50ce1ec7064fde07fc6d120
z60c44f4189b58a31ad241539d2c7f91a4026a3a274e4113749f94c57267f8f5ab85b774451bab6
z2a9275c8329d93adca3c6e086d2696e0f857e9650b9a4874d7c18272d4ff8c6b8d8a7e636e3fee
zdc0739b8ae6416358444a298fa4b2466d6d6dfeaf8c9e20a94984ebf5891cfebc6b74e4b3cca20
za927f4b266f81c63120761b650ad64e1d809e1c2df82c79680f2ede341c4d7d30d0690080fa144
z36914299fbda13877f81ac95d2209dba3834cd31144b21883c8265bf672932caebdea3fef3a668
zb533443d9e26324b2e84befbf3a1e6643eb3be524ec3c738f4cae7e43cc364f7c391c60da91248
z807e1ed71d5ea480ddee1ea66d5262b034255c6f2972530e28bd42151b9eb6130165780739defd
z970f69d41a3fb5695795838aca99997220aff9e8e8771972e286ab6fd6760c616760305c110b94
z0b7baec330688d18106e8246fad631cb3c627c15b2b4cc127cec771c1c13b49a8bfc96dee0ff67
z873be22af9adc5f1a50732c6dca5e939d98d872ff4a4dce51cf28d9f898d3c5b3623fb760e0eb7
zc8b57665ef32befe99bd07ad9e5c9f7d8b0f6b14823324a56be3c0eb8a3e94d70dccb414f42030
za07f36717915ed1a7633fae5f1c00e926deddfca614b959c555f3b16691516afefc08fb06d1230
z844e60fd99d0d49963b429e3d9ee7320d13d218f896b466fa9cd17b08ba52bf2c5574786bb9f04
z3a4c725b9700b1b07ad665cf90df3feaacedb5a81ab5dc86eee9c2bb000df5db6cabe83f1e2e70
z5972d34ed495955f659d9433e170df7737b2314be6dbea38aa834c1728725c66c8a2ce96484031
z3be280db7ed7ea3742a56cc66a3e78ec47c8e537ac6331ef3cedeea003168d781ef227ed749d3d
z5e7b31d655479378f5ab08800014f0a7700ccd3ee9f7117d0bb74475453159251cdc7d0122736f
z59c529c2c2c4fcadbd6b187d94d229f0b104a31506d32a0cdfd540e47571d706d83b4feca9c9a1
zd192425f67b3c6a180e57a3021c993376baa3528e2ac7cb4bbb5a328d4f778c6c0fadb4f4c40f2
zeafeea699eb52ba9045324a89cb6084b47199d25a70029dbbf6e75e07ba373775142fd841d3811
z0af3e4e8310da54aa871ae4305a1c2950bed3d75ea19db7209171f5ba4a33095b69d237752b50f
ze618eb21b4498a30c31b13d65941890b549c853bf638088e91c6f28beeb449f46373112ad858d6
z70f34c12ef27962b3a235ad3b2aa3334420a5c37ed777b20ae94300f5039f24c794923f2c3cb44
ze002782ce031891a2a7e1d6e7a26086010099c7e4ff25ebf2753d9b53b692af626feda35af5669
zffaff4e8e56dab82277ebff89d9d2a6044c8bff31ecd988c27dbf312a6e54e0de929c8f1c91fba
z6d473729bca9c08a43f9357de8bd4bab7c0a599f51458b2c2026bff24e60f1982e0d3b15c88e9a
z00917eabd7b56537a9ce742c7404a4f324d9b44cc34c30a4e3b0ce7fb12dd074379c9b4bad66c3
z918d506a7035ba2ecd7fbd1ecd0cf679c2995201669a472daa38cbb229ff1be5f028b6097478cd
zf80a085c74433d24bf03adb3dba9579acc863ecd95b0ebba9e1c23e1c7a6c0c49066f10c45220d
z54da5257fd377b523e0962b3672c81474e8a8cc212cc1aed34b88c699552d8d591ad66605b66f0
z5036bd28dc1945d1b6883e4162d837bfc32901c561c206a0cd0ca34751f711b5ff8ba597fec173
za8141a66e5e445dad5f91bf1fe3b4cfa3fce39b8aac82b7cd10f5129465d855ebbe000e163d494
z2ff4bc32349745b46c9f0b80003b6b60a6ce1e63ee9f42fa58d429bd3066fdbc73063c8e2ff9c8
za34bb0765deb50d925ecd9feb65da41a07fd42fd81aa3ad47aae7109af94383837bf72d346138c
zb8088fad252e93b8f9200e02343ad34216d3cef79666c63d6ad7c26408cdd1e16cfe1a803d0f02
z88730989a1356f14db1689d9f2fac8f63f670dc8a9c33e2c8d5577cd0c621ffa31572f48776e17
zbdfc8b22c67041c89130128b8baa97acd7136f895b564131f3df2656aea09c766beddd1fd6f183
zd1152972fb82f35dda47d3510600f8dbfe940f59ac653db09cceac26bd1b4334cde337e3219149
zf553d947faaa16db5fa1187dde663fa51eb201617e0f7d2cd2e3de6468139beb8e7fd3fa62d723
z8d264e504cb0e6f4d93a41d4159ca7600289ca3daa0381bd65da8479dbe2b27774597f9e222e70
z5a5e682ea61830d05b3386feaae7cd75c41f324d5a2e8e04ea817f7bf1d85aa7bf3418d3b8cd4c
z44dec4f4c1c56ab5b9f3b188f02674ec7be1c3447d7d1a92151e9d3c81e351eee4209a671f20eb
z63b18ffd27be75cb253f03ee9dfd2fe26d40b51ca67f745650f631e27335657cb3960dfc600a3a
z2d2e7f549026b0d681085fd444870b49c53908e5269b74ac92b380fc2b7af1c69b0d29a31bf624
zd6420d18ea5733946937f49b4223891e9a0fedd92b5d45ab17fbe9fe9bd14c92e56cac68487a0a
za5807dcc1f873540d6dc1de268589b49cb15ff6b13f8f23a978fb3ae2447858d9436d8b9a3f832
z85959919c4d7d592d675c01243c360492cc361ab7eae5e79403fa373edffa674773f349e5b12aa
z4b5b8c1c3e55e8fba8e2adedeaf8f21bcb05d48427d8bd1c3cfc7bc31ce64e7314066961591116
z10582f06600007e12749f957c267108edcd4d4a8c07c6b456a551759a6f05aab1f5e5035b8e0a2
zef8e4c4cf03b5c16aea0a2cf9036160599cbd965b64bb4f867478287b0e67a933ef4305adbd203
zae41846f798cd3770861395d5c2c5c552855d19be8916a61e8777ee79bbe5911bbe822f3abd91b
z4ce24ef5d70c30d0a4715d83d0c5cf6202434669dd48483a6c79275cb58e3ce3a9a4dca3cde63b
z3d8dc44e42afd94330054e52b8d02c539741b0d7b1a50c3d7e99bfd9efa7a0c36df83d9df8eace
za1c9bbfda64c5f30a628021c5c7113cd159526f17ae22dd6aec289f3656eabb8414da3557ac25d
z6049b46359973acbd3872177981527d2f84d9a05e34edcbb60ab3bcd3f23543f61716182e509c9
z5c854eacac24564a500f9502328e263d61598ccbd368fda645c667a4d004961bfb733bd2457cb6
zcb93d12339e8634460b0842a0e87f46a335db21e93a764fbffe19374b3a9400b9140ec71cb0a47
zd10422e0a74f6623d0cd5ee91784e9b9386bd7255bdee98e9909321de0780be1ee9bdb54487a2c
z31c4a0fc13736c52ae2715cf3458d736bb24c1a5ef18fcfa610c814a99014e37fec2c6fb7e9306
z0482f32000769c2e3178291f41607e3ac9e672cae3cc410321abc36cd12814b8f9c8324d370a46
z1f034234f0095a83e12768fc21911f9014885b441c6d4c690236390c8c65de8719cc2f7226d9df
zbd881d3824b4b585de5ab4226fd60b0f505f9e2e4fc22959d078348db21a94d5c201268038b795
z07ff0533bd807d84b4a26a5928c06f17a4a46d084af7d6f8af71615dc8308b71f1b9cb05a48d98
z922ce3b73acd47f12e8082a2dbc6f1399d225654766ede568923081b2204355d17f93e4aca8e2c
z299b09b91ec124b77248fa7764fab269659d20ec779c2ee6be77271f98e64e5d641ca42e3785c5
z92256e75c4dd3ffd9642316b9a5b99b6615541f458fbef6b4200a82ec7ba591521794194847e50
z4ecccfa46bb34aa5950bdd1c2c5405e1e2564f253025ad47ec5e17a1db88acd6118982e512abf1
zb6b9ce9e70abb2400f6974216b20288389e7e74eb259df492e310c92caba972d53acb49d46d149
z5ca2d3c4742eadf3252442d15212eaac61f0c30ceeee981045b2bacca9cd232e8a69763ff3e465
z46612e544cc0acf83510d38d9796e0215719c6408d96822c3efb5e44e1d18879e15a05e0d8facb
zce9659118c510ffdda617045c627c5cf0827dc3b75507e91c2f6965794e673d7292bd49235ecdd
z705efd7c7b90437418c24e367338ac7c349ed45b1bf2386e42f099775fd3cc1917c0d5572a2aa5
z6c307996258f1158807a5f0bdeb61a53725636bfafe765aff0c9411b462cff9ede354d26908433
z33edd9da96906b6287c7dba0624ed8469e3ab1962ca1f1e792263e9396c0a3fddcc239c239124a
z81c138eca11ffb31c3cd0e0afe917401bd1f6b1a62769475fbc3785b9fce8ef48c254d0984f418
z3eb389d2d959a8336e2c02fb0a868b162f839c34b365e05b58118a783821f9acce2427a47e1773
z2b97369b91343cd37ea22456d8d76c37bb033840c948d9e020b57273ab6f779e6a8f3924ba82a4
z758fbbb4bab06e634247ba6d3f236af7f938f4d54ea768f151f98c17fd22901ad472ed0916385a
z5761f8c72208a92252374dfd0100d59e6fff7fd0e91d4718b3f45f0a2557ba99d8237742bacac3
z2aa7175d766d266fb99bfc67138f7c48320aa0521224790f787442ddd6ad564bb76087dc74525b
zd0dc873b1dd6bc7955da8321a98fc3fc5841c56464ddb2d535dc99ac8280f17c04cc4c1de9b030
z4668ae2188d9714d1d99c520a02b0eccf5d204ab5de15f63c30d80c2392cbb17e05bc6a938d98e
z8aef6b211d8ea006262f0d1d731be4292bcfaabf1faca4ff93092d62b4defe2475cbb0b7e4d8da
z728dd775d3e5df33610c955c11b4eba7dd2a9b846808e5bd03b666dfbef1c4282b7e433e188712
ze71c608097bfd70a9c9edbed6ed1034957f9fa5016f24ebb0c0377f22e7973d55c45d9ca0d6691
zd8fc88af147b254b216bd6bdab3d0ddda6511ed0462e14acd7bcd65171967129275554d3039a83
z79a7fc823349eaa50e5a184f0df801f366e0d1491a118648c49c52ae9158ecf7d20ffc73de71af
za1660f3be71d72dec76770fd526372b9e457398f9e1d19efadf815138c6a8cff176feebe56a16f
z27dea3526c855c6dedceaed50ed769cdd4ed7b4a369b51dd471a5f36c9cf8e68ce14325791bea0
z715c07c4e4e6745cae8c4ff46b4c283916c44b750ee74a6a15d2a1370f4e6cdecb343d7de23c5b
zcd9810a9b2ef1a50f090b81334234047ea6cf32b1284e1fe0b844603b282c32b5f69601063d665
za8a9961cb8c74070ff798adeaca9930a9ae33bd2ced9f133ff3ef77ea478089d1fe52ad65b79f4
zd7007191f90d253a7d6cb4ed9809e9fa5fe841b523d294dea9c0196c5c4f0dd6f6bcbcc67dcaf4
zcc91691c3f1e8ade8eaed4035534604d9609812902783b60f342387e4328bbe3bfe298d6470eba
z761e85c94fa8dc6883273f5d6401cdad3674a75eaa6087d0ac94e15d2479e22afb27697d2ad208
z2bd01a30db9819990745cb4451a725985eac80965a50ad7da585c2e80527d93bfdf7d85fd24c77
za1bc71898a8786a97f40e0b8424efa8143683da301b20bd3e80b08622e87fdbffb60162fa80826
z15cd9ddde2cbd656346d887b4e7d2b46765bb453209e4c1637efb203ec4542c5d72fa6d3140cc9
z0e7c45b36975ea60155ef66f43b30c398a0364f3b9e9739f4e1de1120cecfc90a1b288693bbd3e
zb549ca1f06a572d565622620f967d3a6d7ec5cc017149b882e2b02ba07b49d8ac8722722cd34be
z2cd87e12f1e1cebce0e8e483cf4f461fb7ec37dcbd9bec5f2c8b978d9461c48b6dc9bb8c5d7252
z1217ef06cfb81b94952ad466b373287fe0d55b94054466800c2acd8300a38cce57a9ede101d63b
z43d8f1984918705d67943d0e37cf678fea9487f1ac179dcf50a6a07efb51f0fb3caf5fb7d190a8
zf694ede44aff1854d4fd626f529b222c7210ac0ccacb7a0bc661416c36a3152286b61ed76b5133
zee72bd5ce39865e84ead585d397c2e22a62a72cd7b121a53c4016b5652703b170243bc36ec0bc3
za21b4b53c57b045248b0fc21c5886033ef876db08747d3b3a85e101a42dd5ae583101567cacaf2
z9254ce6fc991a32f1d67be6760881c2a02b860d3a7098f691c924a049bc6fd87b2fe61f0a21395
z9c1ae10f7931be30e01d79838eb5c99a2df944244bb9c93f0fea820e3cb876117dd7b998d08c04
z9f7ecb89776c6cc6092d0c0880de202bdf28b9afa0e6b02bd092b800fdcfc18749aa46e87f9882
zd04f2d5555bf8c333f2aa7cdd11a3cd85e39eef5ee3fee0bd8c930f259ea147ee02bedc6d7f529
z3bf68e477d461f224c176e50dba4b6275f28139cd6174bb68fda5dbd82154088dbb93cf59fd9a7
z6804aa1ea059162429f1b4c8ae66fd37d74db8eeef79b8549152e83fb7957516ac57cce44867b1
zd6495f1655dae20df4ae0b8108266c067d4c4e719e56026fa0f7fab98b48d2efaed9e83b17b863
zbdb34f33a7722d6d3bad18c8d6852288050081ef2db7770f0f2b79152dfea07f4b50e6aa98b2d4
ze94cfa9b73ceefe88bab6bdcfab0a367bdb35323019860ced5ae03d0b68b2fc32217e622f6a465
z57589dedfc438909d794fbecbdd55a099b50de31cdec7a05d1e547ae8f77f4ed21108654ae517d
zcb68a99e6dbce7f4aa9b9c16938c984e152e09b2b42f109e3eaadb3232d8f09421b1c31b95fe3f
z3f17b3aede6003a709880f64507587b146d660c09ca5610524dff2889d9514671bd05229986260
zfbb4a52afecde3790fe408341c3225ce257aaaf34734e8483a8d3c5a45f85f394756e680262e8b
z10e4188f2b9ba0e3e67953ffb7014b7d16a89936d2b6a996b15298cf50612ccd60550f83966c7a
z44a09a71f4d2b7ec0219f2ac883c5bba5b089c941dc5490ed42cb5ebb27a33e4ca945c91665dce
z8d15a50b5440a7797425f38e184f4b0288ea40b90ae008717fee2e02e3b8ee9fe1bda34ede4969
ze279369f498a47bc24d0f09167b53644d7d1e7c8fcb44e6e2eee51f2fbd2786ac9f5200175005d
z69a560dc84dbefa1b991cdd904f312027f9673414474fec6329ec8f90c92fd02142aa2046935b5
z4d6dee7c035abe124175937220e314bbe4bad1c45c9a2a17024e19441044460a84cb14f27ba927
zd979c329bcca444e799c1d81635655b3130118ea710fd01caee635b181f0c7770e332353e37f84
zd83a57e3899eeb32df64b0b658d5ba5de6670cbdb088119554db612dd4381d2b5a0932a8daf516
z7d5dbca4f0a171adbda5e5e9c206b5915f54eae72b35f95657ec0e2241998dce451f7e205da774
zef799179ea54986fe82c70b73b87fc8d74e34000bbc219c4d9856212b00a971aca75a377b5e0c4
zc2fa0d54c47927ca33bdc7bace1c2aabd2f0fbfe7528bbffdd7d9d4cc4dfe763027000cd3b1392
zcdd9509bd7eaf68098130f41e1eb1a25b54f5b043d468c51e79d61969dbfb283b406d7be7a169e
zaaf6557be6f085c8d6da281636d90b8b148160d57095294feb898c001a2d77689f5a8d6b27dc00
z33eeb45e73cfa605b4a4a11ab15bc7e762e114a0dadf7b713ceb698829936d7fe8cbe2dba1aeb0
zf69be4d8ae83d0b7022ca909bacd53b465d81248157bd0e3bd4c16f2a455d517e7b04a8efb72e0
zbfbb9769781ed5b1d66b06fe794f6d2a8ac7450af0d04e37bb1e5899b516bf15f3bda52cde71e6
zdf74209e3a2b2c8db88c1dcb44d56522461a7c979b44a52820d7b9614a7e97c710b72a2f244529
z6a127390754711c06c6f9fd8d46dcfc95792f6a20898dd267f42d61b81755025252eab673aadb1
z3b07c1e470b8e4b4370ee372dacd0f2de97f43f6c9035432c208336f41a5a8bb12a524dbe4e56d
z1a8d4046c5acf4ead1819a63c48164c8af075446f42002627a9d5012fdcd17c87e60d1174d316a
z7e1f7df792d77ebf31f544da54a3f88542a539c5bcd6194f8f948763b7e2af4ebf2c0d77eac27e
z81253af2cbd5cdce36dab1b9b2dff404f5bac767c665bb5d6322e3f8e1bba41ffb20626091d7e8
z51c039804807ac30fcf3988e86f7cb605d3d8083af25facbbabc01ec560ea2da161dfb96d625b5
z8abf796a9c41be3c801e88017cca85d3ca82af0765116eece328a0199f13fa1978fc75891db889
z282ee80c94eeab63086be121cdddda0fd33965f1376ca2379a8afed58c212e9cc479045779003e
zdf43b62e46c3c3171fa785e68d0f43cacaab07f2b4b149fa1408370adcfb03604d4f3ebf0e7629
zae5d5eb8e3381b10c283c2ff13844d1fb074e08f6bb166659060f7d08680de531df2581664a4cd
z6223a1054bcf7ab604ca53efa68d272f2a5e14947984b042fbc09a1a6d635a981f9447a4cf4db0
zd668b3c9e27ee63f3af3c9642e44fc7ba9a9ccf560009684841b2738e9e06e79b8945725256046
z9beb429c961d6ebd0955035b4018de8bdea6b3d1d2101b7ebdc3607a57ecc2d89138e2d8565117
ze80ea6ae3def7a74c1124daa4ae808a9a1c3afa1872bc8188a16370798f168e1fc1078862abd9d
ze846f60e77a180f57c7938837c2ca43d27168cc567b16b623cfa6708c156ef4814142c9e815cb3
z547ece6cd2f5f00863569e76b9a8ea87bf84e61a3175961bb461d46d496c90b70ed752607298ed
z20d87a0046b1a6c050089e9edf9799c60fcccd8f3f359e2b416de551139296ed46b1d26992aab0
z81339d7cb3abe8f51de00a3f677ab8b87bb51764b3bf67b0d59ccb2e7c342e65f1d09f0b6afdfe
z489a3778a8b7c4cbfda488d40dd81cabfba4f8e84199406d038ab3b869632d8af1415341ca33df
z0bf1b6bc8bbbea50d8b6c9ba966b02cb59611bf2acae5fc154291e6ff8520099047caaecea872a
zdf2cdf8ee4625c3ebb6c5bbf64fd0b736a5f9de2420b260b019a8d8400b3210de1f7b095cf7b52
zfd59fd0a63e2fbfcbf1e537d5f1f1f9581506eda5213242c8052b100f5320d02aa697579464f24
z3f882bf04d971ffa943ecd703884e45ac0bb245178880ee61ab8c588581aebea68541f008276d3
zbca102226d2666a679de6b0c4837b04bc92436fe6fddb0e62d37a500a647b2a80a188424ef6d33
zf52a30b8800ddceb63220c36f04dc71cafc08f5dee095fe93af05c5935d2ec93eb3594c7fd2a1e
zb21c923c05720cbd82e2fa730fd2a831746e5103f183da5d403502f8b3d8d061266b6f7953be8d
zc30a746461d3e3068cc519e927f8ca3f76f3103196d043c9f83e8d97f343ada85d3e38875103d5
z2d65e4374fe3b8e5d78f4766a8a4b36325d69a9c33047c6232ab2cfa8aada98fdf7c9f42a2ca81
z220a9e248e298a62d39ee5e19e4ddd38e6c081425f54d6352370318218221830857b3e2f7f1c4b
zf1f72ae05fa75bd46ef1a97ce010d86e60bc1f83db2a233172dce2ceef66e1881d61227c7a9e56
z6465f5906974e1faec07f5fc2c50a84d108ca7695a5a725323a8c588c5e303c2b9bdb86e092fa9
z741508e817234879ac5c8655a7442d2ac2a8cfe20ff578fdd87df15c1c68c890cc2e9547e71321
z3ae5622634019f8620ce33f7ef026c362564620cba2a34b2d0eeeea67109b3e5c7289ca8e16de6
z8233bf486a0051f22fc82d1ef07c69890ad6789ed0a2dca7ef3ed5b2f4f057c73717a4449464d4
z479f5ed2d141e9a2e28efddc6d03158ab11ff54f25ccbaa7c38dcdb014288cade67134d68a6bb4
z4bca01a3ec02238c706a6d9fb8514da4bf81cbf633745ac0c63c7e155b977607ea5c1add11ec29
z075530b1386b091315e080d1b0d6fcaabccb520207d46213995f6955b29f66fd4c4c2fdd20adac
zcdf8654e98faf2a932706b67dfe689cce96e3edc30a6f820c519b24c842b54b73f53334d3124f2
za14014fb53847d1aad01ca53dfbe551852278703054f6718cbf57031ec4a01d8c5dbdcd2bad455
z9f08e472cf52999f0e7b4f2a9a1eb5de36e35318cadddff2a3d60228db41415f85fe49543fed99
z20178357e1f092164721f3e4abc076b64eb3607a4ae8bd67c79b95b18d9376fc9d03dcf35385e1
z8050e1297c666b5de578c260aa7c7b4dc19e4285b18117bcd271a58c499dc69022faad387d299a
zb66ab279a5f6c027702205de100ac3c00118227ec51700d15748fe6018752981f5f282421c2ba0
z26f433e0d8560b03916a979f088617a41ce8219b9850c1bea1e00300e6e54fd91d5745d516f442
z252837d63723b7bac5094bdd8e3bd40f95ae801c5bceab86f8779e6e782204d4631d35b14c0f0d
z852460f13606664cadda1521b13d8ad9e61e294b28882c84722987fceac595151bd4c1cbcf2901
z57575dc06a1152526d8269591dc11f0061731a6bf8aa7a914c03232de796e89e7cdb100c7fcf52
z82f0d5601d319e33f875095bf33fef90956fd313fb4f180f3ea7f50a6ff722fb2fe03ac98b4105
z128e1fef809b6c8643a278e33f41901f209bedec3ac24d0721364183c83ec3d55d8375fc065e60
za4323168d65f6935f313dc4e81f103500b3dae248b03e151cfd5b83e54599a4d3de892603317a6
z55ff7509049a4a768c5b8c027d41febd521c8d6456c7dd0250882586f5058ee17981c40b0c3e27
z20ff6260f41dff4764928ef17f63826cb952853bdd9f60776a11f54f6f173cdf948ea025968b34
zea8ae8f1db9772b8eb7cac2f1478167bbc396ce74bee4f43e733e7bb97020057efbc3dcc722b36
z2db2149999658ad6a39ec35e92508fe96232410bfb03ac685c4a23fcbc72e9b15f36abe0facde2
z92c13c95dffe4b94c68cc2541388c6598a40047bf40f41764d2f58c0626b1c08669720c7c7f739
z696ca7f7ac3d254915ce72a93454fa93b78f535f4757e8f72d1f3937ef24348ce3010c28bb5211
z70171117195d7a656dfe18a2ad42a48daf19fa6cbe6798659c06d3fac4a5ede135b2ca2de834d5
z43abf10b031a9233537e85871d4dd2516cd40a9f8bbf0cfd9d0b2a22067ce9f51a0d0b64ecee58
z75aa6c877e2bd7cad77201718bb8be7b1fa86a24b590d2cd2409795c8926eeeca0377c8f436254
za004e15c6d0c553afe63ad3ae57a814aafcca99ee298ed89129dfd35b2fb1469cfec471f990d4b
z7c1b207dc47f67d2d1565a8afe96ce28b418077aa1ea8b2555aaa386fb5510d509a452f5919d6a
z801559dd00d1f09dead1d375a40a80ced7ebff70939ddfa53f3a2378274e52ba8d9d8bcf1487fa
z280292aac89417e07717e186942cebec0ea65cab59c6482b630e1c9144f7458469d06d0f5565b2
zf880ec385b8e2066430f952affeda67412ce3f2b3c3f9b8845808e40d482168b439bc5eaf489d0
z81a9aba9931bc73275087fc05497052863113e32429b1eb5e85e85241f5f0ebacd4b799651ff3e
z4609ab76847e4e06646db858f862a32c9a7cb035ba557dd9e7d8a6dd19b375bd67ed7fd1fc0955
z2fa3d348ccd933e9f88e138c1bb95be32bd21dafb03c96935ce755b905a9754fb7fb5e897d47f3
z4a1f3adbe84900921f6016dd808d8301c8b3cceb5c3e4ad7fef0058bdd48cc5713f62fc4d4e2e7
z763aa840719f447d753feb429980252245672fdc44d178b5a461caf54882b315ae5ae338daa960
z324929ff946ac0d945377685bcaf89eef0b135ed9bf7d94b818d15acb6c667d547682107b83716
z174b23639f80ea285cc52e166c3da9afa49b0dd99bad68aeb274a57ef81e4e513a54a680b25b14
z435cd8b9ba45a95bc24f60c0b975163a282c81acbedb8a2aa4f76bcef9da2feb137e443f17b3d7
z7badf094985fed01df586607acff149b7227b558d9f5b4273cffdd2ad9c4cf0584f51f956596c0
z6c1063d40318f041e367165bba0eac627c6dc28d83bbab7fc5a4645fc8cb6261173e6dc1dd47ff
zc96b855af4c7988103b3742c4bb87fea790454349e6a6596c16c2a035ce207a76418460c4a68fd
za49c68ee843e91725ef2a508b30bfa54a44ba18cf2b82bfdecceb078d6d4eb68938ed97c872c20
z5f59775b8e27cfe186ddb4cc0d74fa4b86c4b34b571a66159461a23c1ca70e9782cb4a2b2fb3b7
z9e55887547d53d2fe724978ff2a88c9ec5a0b82ef326e94ef7b4b710ab28ff1791a2c3a7bca9ac
z5877382e04bce760d8498f4c53a5a5794fd836cae353301c41f24bafe93697e13ac250adb6db57
z5d2fcb5fc82e1d3db801b9ff1727d03028452cc5924ae8d074d64e8967a847ddb0c28642727ded
zea8cf9719633be5f49e2bae197147f26b182e3abaf39b637a6af3f4e0d9f1961c01bdf18520eef
zb7cedce1387c1edec01708bfd244e128fe3702acb563401d9a255a15c075d01a764702978e47ee
zac4b386d5ead467adeee49a44dd4cd2603297e464e94449c8f045948f03e9ab058aaeb8fa9f291
z398395b8e5d80390e84cee3fb3d520abaa5d5b3ad5cc4e9f20b4c15c15188fb7b357837ec75df1
zf61f71baa69ccaf0f5f0d8d85b630178da0aa84732fdc80621b7afdc38a532136687ce6ac05925
zf87ff7a6af42a00430a3ac385131d2b349a2a6628df1f493a5d70fb64120cfb57df4271941f3f0
z919759abf54f779838ceaf48f6d1a8b5d1d321b4611126209f64a1483a9233727ea8ba3e8832f7
zf41023f24a1d740c28ca71e7d9d4d30334b5891e03fd67d88151bd35f57ba4f5695cd2685706d9
z260906db3fd46ca14ebc00ddf4b46f266e4627b525e2804d1c9b7c8880cbf707775ce958e7f106
z1243f175543805c2684e93e34f06e22ee2076ebbdf54f67ed0c00cd6015aaba786eb03ab3be7c5
zc250cad966d4364574ddf94332bea4d586622f9977ff9c06c614547d6426baff921128d81ea2f4
z6b864dd5ada718c686411b5592c5df9451bd8bcc44d73d7b6cf8a3e322733c789fbb995ccf5f4c
zf5f56072c982669f77258c0f3103e5a85e7f40eb3c1b3d238e96a1358cb05d2e2c89da703876c1
zf77ca218bc53898b5fa191b69610c775c16cfd82c64aabf284986d88dce93155495eac1825cf8b
z212b1c6002171fe1d395aea0d267b7ec3957fb8e3f9b93832fec4a2c587404d1b87d5d816cc583
z7aa08a9f1e2b5e8687de2757a584ad06277ddf6857e05e70f076d391d285f039f1bf6ba151439f
z5e32b62df18bcddd780c960ee892979b9cd160c6720d1c282499a26da9f5048f6b704203f6b145
z9b286c59ffb557816661b50ba73e1dcbee0361adf9d38d1fcb25eb81d117331a2793c51863d8b9
z8d5a92539c1cc0b26ffabc0397a2a59ad196eb777ee83eac4031b2f83ee8863a1e9c4f432f9f4d
zed93938c89c88577f9cc6f3817d12a62506c83684a16d0cce468606b4c5a55fabcfbf8f1d13412
zc843e338f1a4bda3ee154a78ba716a316bc61144805d202be0a78c5e56d4c2597854f8753323b0
z2a9cfa24d4848b3d35f49bb00b111bd50de253839c01cae8d21ebb945785dea5cdf4270481d126
zb30d70910f018e6de78adbfd8ce534d92078e9601d67edbacd1e28deeaca52f6c877c2eaab1e0d
z1f0f72d5bb12bf353118167272cb064c296fba94867660ae81f2cfea88e09ff55d447797e3015d
z52e1e964f2dff36aaeb27d32c071c14600c97bb076f6bbfedc26678fcd79a09e03249418b30bb4
zdb3b917ab190a0b0662615fc2b025f276eeb6817e1fdf86ae408be25d02f54f3c1b39fd93b5b2e
ze5f87203971c30753a022681837545ef9e4a5d26ccf801fb10503a0a28e1567ceba1634c1ca634
z70fea5c68e439fe28dc4460b6139aa4d13fc06d9675d5a059d9bbfcced2b8df306cbf27a99df6d
z8e356e5848da1c0cf6fd7748189948ec6dabab3b5d8dbfbe9642ba274b1c806033a184e768fa27
z02905fcb41f005e5ddd7e6c758d28f2acda5b77c0c429c98c149a96cd6c00c98bd773ff1ddf839
z57ed55cf827859bf0ce7d7a42bdc4d10cd69e8695060f725731b040b84f6323eefdd29f6fdbc9c
z50865997b3845e75c04b74b215f055d8857e7f800fd061206446b1f70b0a0ae2e0243b4b294ef1
z7593c1d8850eb2cc6515c3f7322c7351297045ea330c3af1733a29a3c16817e7f9100c178a9dab
z8ecb0c6456cd4a4017813a0ef1f6a17635ea8b65621c5c1441d9c007a6359e5ed5d8a99cd08fa6
z1a395e4c9c6ea303dc8f3669fae35fe124c531286c1ad46741ecd17a6d57819fbca7411ff1dbc0
zaf59f48af08e03b6ff07ec6384a21d6066221c553eda397d89acd2122b187e15908dc4e2b000ef
z8c9f2b13e033ddaaa641de09681e7e6efbf0556faaf65d5cbac615866248c48490e55238b3da3e
zecc3b0fba4fe5e5ce9f0a9665de93ad265814648723e064d026f106830a23dc28b1e8feb1a299b
z66c7f2a465c376168361d042833fe1f1cc1db4a1076c31b8d74a7d48362ca2bc31fb0a631d7565
z8ef75beb864b40cb00df9b08f61b2f4329ce1a32a0ba8f3614a8dd79439901006e45a730fc4a55
z39309347a28f293dd212d6bc6112ef48ad5b295b38acf4c42af8aff6fd2c39511e93305ac371f6
z3ae03303c049b6964b4800209930c136fe495e0572315d670988fc222904f346ffdfdef94cca6f
zc2b1b8ff889cf5f4d797861e4aa2cb5491f28f163df773c052ff1475aeb1358b30cbe9cc1598aa
zdd5e7f10f8f6ed791f6642f013c42bfde8ec7922ff6dcfc8a99e635fec24504e8cd00172ace194
zd5d9210641e944290451accfdf267393573c7f4bffc5256cb7ccb7d701cb8402a56b1c43c41b00
z7cf6f0a5a91d3e1255ebf254e3007bc7095aac96aa519d4881094e777962f6834124810b91330b
z1fb0ad4125806b0adf5bee04e24f2cc8f397f9eb2b2b28b676600e66e25e21f1e226b926e4499e
z76d753777c1e68ebacbbca80c98dd1ad82696d7385757ec3d98450e90856625b95e9add4f1d38b
z8804df8c57d332101f190a1c75a4610b97b9cf06f3f7aa7d1a7fef31a42d37488dbc1612642e8d
zf897a0eaba871c6c929ad73eab923bc8b11686779a9f599bd28599d39e49e08aa661cfb46753ad
zac32d6e4c9246d44fe1c5a8b084eaa8cd26a812d594361797d6d30c4e1a3e8dc39ba660de85111
z459c1daffc8e37c05ed495d3b5dcf05cb0e07ed8240bfb2e87d736e8a861b6167f8dccb2569d15
z7ca265a52e44e7f5b6c5a1867edeaf01552b69cd2f33bba37c14637f6ef78189056a55ee725cbf
zb6c5af78e62b34ce1d2e12670078250b823c885cfdbecdc794da6449ddc90472ac13f6412d7351
zd33d6d9bfb974aa2a344ad4bcb60a313b5bf687b27618cbe6757993d5085fc4484a9fedf1885ae
z617106cce347abf55e0f6e9a4b7683abd3ca7f683b6206b123faf3f1e6004b78ce2b65f673d488
z691648fe1e701a0367a1dc91a2f9740ef27edb71c386671bf6e387bb867ef8c04d6f3e2344b02f
z2d79edad4441eb4da0eb9f9934f65da0e0cbffbda0ef7566a1db78a0d731054c3a47722883adf8
z7b5a4d71146899872171a4ff1a33fccaecb64a03c495dee40cf53ab084bd51
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_express_lane_receiver.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
