module divider_non_restoring (...);
// TODO: Implement Non-Restoring Divider
endmodule