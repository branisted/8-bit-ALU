module tb_adder;
// TODO: Implement adder testbench
endmodule