`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bcbd1c7074
zed3c238338730fdeb978e5a05edb18654138d6fd72de6c4ab74d0ccb934b93c5751c4f139ef424
z3ce768762519ba13d8e379cc659fea22b625563d2adf866c5de8afd014ef918b19d2d6bcb18d35
z948f5452d4e20dc2ea05bb6e40f4e32834314559686f1fbe368d08f0a9551bf4bb639809d1b851
z338db16796b3bef2ac5caabdfe87a77eef6d358b1548ca3639f13833b5626ed1a21e9a16f5a1fd
z5c7a7701277779f801e0f7db33cc44c9f7f80e9db47e7cb2ba9e013fee56a8f94b35c7389a932d
z24b6c0d36de31c1f41c471424bee29273c160c357084842a10a3019c00659b30cb41614c553d16
z149608c4fd975663872cdc7cfbdf4f33eb2991e24ef2c7c15c0a850e4ade3db06b5f6d1f85f654
z01aa66786666c8cecdb89d336585a56892bd10ea46e156e4b73b4d8af46b0105ebf316d27c4cb1
z57c7361f7d6601c1a8a3dfcd544e2b8bd0179c39b50750a591a2b9bd23d8523bb479422c507e6b
z55a6abc75f1163acb8db4eed22d4815ea5d6be587aaacea14256de2cdec350bc11aa74f2ab476c
z718e10863152ce2c9de30369636eb4f89db1ebaa822ec9eafb619d4bf3d53ddb012f96b11745de
z95ad4b6c826369024888aebab6f8323a5e20670b3c3dcb8ef73fe0e76cd8121349bb1ac9c4139f
z65201a7b291fdc552a0cb4648d09b4482847ce7c4c4af82d98bedce518526ead6c590e20f03359
z0125ef235ea89952f36cbdebebdd3cd8ea01ffdaf254304f18a82d1f2f142eb5b24b9dc9494d32
z85f974a2f672c2635ca3caca623b343f1f91e47d3a0a40c676011db33e5a7002e8b1d437a0a13a
ze641ba29a4c65ca597f45436fd97e522a1333e15bb14c87a2d8aa1e94f450fa6b4ed163a08a7d2
zfaba8ec3116093944b84ef13118748a2913fe3297c67415d7349e1a27d99c1f3f32e148704f4fa
z46a3b458cff5b5b1996e651a6cb41314c44bc3cbf5dd777a1f7b6cdba544fd04ecf3ba5cf0bff0
z43f6739925aaa114e6bcbef0f56ed939ed0019d1a7418dad12fcbe2d3f4d4cef6f88ed93a73f9e
z2398947a73067b6c015eef4ce004ed4902c67ffb7d28a1e45ab50f67d3400b6f6575a45299534d
zc5b11f4966c78b6b50f0f7eb2bf281abbc44b085c3adba93f2a99917d1017c168e40527d29851d
z07b50647ba57835c8be31a9634ddb92d26dda9000798217e310c73fbc7923aec0468a4c704091f
z2662619d645130dd43937fcdd009a87974af826876a35f6292734740ab242133fe881873b248d9
z4fd61bff5b0ce68601b9d74ea7d3032a9495b8dcb6f310647653a8323d268fb0a485a5738a53be
zf8f7ab73000801085100d33e481987d68a942945441313629b281e815b4584678478f021ce832a
zd88e8f8171d6972e504ec3b963ffcc69808bc6653c37a8800aefe16791cfedffc76a21a311b4ac
z1bb24f688fe05cdd767ff7abe93d2944bb106849e9785dae28df6c4ff01bf4da7564c03c7313f2
zc6d9257c986b7c031236b36afd2bbd4d552aee78f7bf0e719388b3af84f7a9671bb9ad1cd38c1e
zdaa9f0a7ed0171287ca5416d628609915b6341ecbb0208976dddf19f1054054bebdf582f7bc62e
z1a6c482919a4de2ad9746418bebe6db87cb3e5d89b99369f5c23701a5e9a0ed56f4369e9658b23
za65790d14e92ab10ce074891a6eabf06a6a84fb99d4ffec19319c3eb73d31dcee0ca8235ee9d87
z6a46dc0ec72f1e3d08083060852e01db9d9769fa99040e401d1c7523c0344f9d7fd8786841e8f7
z40b1d68b0c885f7d3b5fb61f9efdef5da0d4dabae79dbb4143e431873687ed204451db423c71bd
z7c13eead616eca554f75da295c0b40e9012696c29d97fb4c65c90489cdbafbfe2b65915a383b06
z687d3a3a14514a72020146c7cb27bfe04c730ea1cf3f969c4af05bfdb93f7733fcfe302b2733ae
z341440bc5343d7e15a7b600e804376c2d18dcbf3d7234834cba3fd3b05cea1a53a776845bc7f30
zdfa8fd418a703ee910ae92ba497b6fd479da7792a75c99f29465cd536d45e8cffc50fb34b31468
z7e349dfb8fde0403f0b2b79b31c9340d4e4cd862dffcc1c8ea2576bc4cc82a7087c6f8d021d91c
ze53229af105cc9d5aa2d230f122202cf9a033402f6a9e6a424f91cceee5c8544796d194cd01171
zcfdfaf85b7ae50a43431bad41902f365cad0663fcd59dbf6086afde5d4d764bd3d0118f3127800
z0af21b87503c52ea2d6010f26ff8c64cb4c7cdc2641186897bdca5b1ee0f00bbab633dd9abdb7b
zef8add4783ca9971f1c66238a01f4d8d94d826d8279f7154efb02d1fbda58d8700842c4a80377a
zf1acf834a9fd7827f117b270ed52e3b29e99be3038c4bd3b05415c60796ff3366089f0a2d5a4a0
ze21bd7f8811011ab2c38b972ee0dee7274172c5cd7a6d4a25bf70a224805250c39a03483a160e9
z68f02da861f4c29ee0cfda5d289064b83605aa4037de50ceb330da723a72a92f0e6bdfaed62aa8
zb9f3248017b84003d345ba6b32af8cfa686e72bc656e691ca9170c919817d3d2ccbe15b2d99029
za239335d6d4aee98734406cb5b916ede2c0e6fc287bb09b0175af020731938ff660910df653165
z45eb8f6bb764178439eaf4ee2d242eedb5b05a3eab6c39b625702afc87e96ffb06cd58f8f111a9
zc8b97ee87e814952b2a427d014d2c6ce58c6c2b1cef4a7f984e7b14942945082f27c4882d28342
z968d53f5f1def09cdd5ee7fab14716332eb52410e0cf06f45af2af0027bccd2eef235c4e9151f1
z9b227905b7a7c5d718693189903327231a4f7bc97f77f5d851982fa34e60f0a4b834661ffb1125
z6ff5051923339df16763e2c88f6995b379fe779c69c5f04b7a19faa21b0b686a56cf45decc1728
zf60520a847b7e137bdb3b0ccebfdc3678278d29f8840136668b4e8e8ac5207841c8581111f910a
zf52b100345f6b476e4d781fc8fdce57aca93335d78bb70e47907efbf125aaaf4c167cf398098e3
zc27d9ac6e8d15908b02abf76af883f744c7477325775f4c020210237fab6c27e72b6fe6e777288
z8692091bf6e4e021d2c239e86c4072cd775cd0b441aa7f8db03af483d7d14f72a1cc4f1b21a9dc
zcceb1702c370e78d963ca26e55e916b786a5611ea6961d5b161ff290ff22ef751bb2d94918d1a4
z1a43270ff4e881ca3bac86a22b23eca87c9ced353ace333c3e357b96d67913d1aca47df981f10f
zf7d1619da8a09796c2b6ea6654c1153b1de6e2e5e082335603f9c118038b7c05e56e7133b8ebac
z9331508f30a58542af916e2201b2d31229cc6b7a18707e58f076ed610507bdcdf08a9d08eac8c3
z528ce7d8a1d4de5e80c24b7b9fd58c71f530008d0d056513c5a72dc471875ccabce1476d5cbb15
z20efb90d68019961a112faaf7b263a6f0db7385ff784a02cab57368f4ed8d0c45f643f8980861f
z0de314995823818342c10fe4940d525e69f0b4b16d5b7eca931663bd3c7e2bf3734a140491e97a
z85fff20125a2bfb0d7bb78c204a24b9c75051ae349daa05f7ef25d0cd4b13d587588921c4d9af7
zee880084e9d1971057f1b3b6c7edc3bb8f9ca9f8b40548101e8162e2e9ac1700083568f4333f93
zb65851780f0c9831b1cffd1fd4a9c6ab8426fc73dc27053c912aaf0f40cb55dafca09981d322f1
z37f7bc4b27f08fcc1d8866ead59013ec51e5cb05d64c05e200dd3e0c87c2f3bde0782ed8f92c15
z4d37b13ac597cc511303a88cdf1ca014fb54c17e6d73b9af43a4cd1ee7b2b4e438f7fbe0742b9c
z5ebbd26fea1e637c7919a1eab8d37ac2d7675a42ee0a37df097a5549aec07eba93e1e7fc0d9fb7
z204550434fbb6d12d33733b83200be3470d2a0e787540421b625d44e37a6f2e950e5e2303cfb77
z5d771a16de757f1b249e7fe0aedfc173cb0746c283bd7bce1501aa8c1d7d7f9a73f56ea0d1f366
zabd0185b76493080e05b62f8876159555c41d3718350b78b84ff0d659f723dbe24aaaffbb103fb
zd7c99413e8b0b2f2b75195b216f7334dcc91794cb1b17b56de8ef304d7ad71bde12aaf4099bdac
z4ff472366a42cf627ade42ddfb1c42f059d4223559bb03f05ab89438fd1b868aa060a6cc00dd1c
z312b2d646c5d09190666ec6fa2e8edca5d574e61a5dcec9329aeed386eafc6340934bd2a454717
z79d72382e1c419a419e353475305df4e171c05812ca75adfaf484dd9de81eb249fb6152d00911d
z36d1cac648f25024608dd3e408f3d6a9bd75c533a6fba3cbe789febd68ac52764820e55f142743
ze4ab0c344d16980ff09c53a5b4e4e0fcef6b804592b3646a9ae94dc6a34967798edf35a7804352
z1d1b7442fb1ed73c41181e5ee6c2e4c9db6fc5f32f70ad3d96b672aaa377d2bc0ce196a9b11c3d
z36a6f68fb033e467efedad1eeb4988a366f44b831c69763e3ff3204cbd5a264ec2aa3eeb61e235
zb4354fe1b81932c8d3951a0b5be9721b1777e38f072ae04700bd70e0a82cbeb88a0f5afa1d83b1
z0c35a569e12e1112eecf24c84690a00bce15d83bb68922e6694a07dadc5479d95767d217c69602
zf21c75425463234059eece241c08a8f0b46c5d75ecd0d78fab72f837bdc85f8ce15f77344f8c4f
z0197577c8bb930b29ab107bec60435f841fd62670ebe1a4f76e3b84f4ccc4bf4be713e4f942b9d
za170ce7e6686c9f21da4980479d59702fa5487741b2c490bc867ce129e01eeb22613582aa6f914
zdc1c2f48ab955fb38f65842d6e6b26286e04b32b8e180b22377c113f7d44fd40dfb2046d312331
z9c763f5c082c320b0dab5251a5ea95bc233343aeca7c966394e4fdecebdac40d70e9559f46a067
z98952ed6cff93d857bf75ce9d5d080273ff258a7ac02ed03655dfdaccded04d75dd82f131bdfde
z8464a984b3a7688c14347fc2ce2b5563155801926396a0515aba6bb9df25655face0d0485c506b
z17eff145b65fdf2692f4096550eb50cf67e978c6efc4dbc8b263afe4ad2c44de74f3c7c174b55e
zbf9ec21164f521179e19d5dd0385f5df792fedc1f6be387486d517caea03311ae468967e91a558
z6691aa82b3b7327d37f785aa64ed7118d88df544af881fe185636f7de323d2b7f07f5a63ac0b46
z6f93a5df644f7959d44b534158b09d92670baf1f2393ab4e141216e2c075bdfdcf778afc413c47
z8bfafd04008dc34dca5290e8ef96ba602f2aada1c76fb6ed5267b130711e6763a9bf83d2a60744
z1ed5c31de32e46501ec59d985012ea2a16e1f36193a8a589499376316425d596003e48cc1eaae9
z891df0a65743d5980cf48d61a4001b4c2ead20fc11210296bde8642f896079c0fc1b981abfcd41
z1b781de1efa274864878411b366708c396344cd3bb207c72383cf74ec2c1177d95c71f3098a617
z233620e04e34e4cf46e5646118111a748b79df5259983bd44332590ff610445740d041e4ebab1b
zabaada1d40c6447e3413d6cda92822aff563220c1d6d9efc7badede4f7891e1f6f4bf1a6d2919f
z6b3fb646a89836257ee733d9a6b79133dbaee14c6fcc22b99ebf172f98b06d98192d83789c6ea4
zae0e71464e1f042e33f7272b8dfa6ee7ce34d2569ea77964e116cc60ef6e4cb3d4a09044e9d106
z1308b0ed5a6c96ad3c3626a1e54520d6bbf1a5ef3196797b2602681a61fad37e181e093ee31e72
z290e1f16dad7484607f0ec4bac810449a7770e29db3b8a71bbffc66eb7e3084c29a2aa3d0a1f2c
z90b31544833dc5319b02b96c042d25b13b15803e77da998a32699cc252cee93b865c231cc2d5f3
zac6d893ec799f5c08775cde5d482c45923e5b0c78b87fcb7b105315be2f2b55eea5a91e1f4574c
z72e31c29309305d318713270f461ba58ee9075062aacf640e371aa2f6e7d7cfda041ce8937aea1
zd44a798f8168cb1bd58f4b016c7e90fe84553763dad98b2f1ddc87eb799c6633dffb67c13dc46a
zf78f0ccb80d19647c4bb4143e3934f1c37c9548b6df1b58c8f31393addf1010d7de38282acfea3
zc1b7c99c7e4f59a47387bbb6e5e7073cee34a494d5bd43a75c37bbc3b1c989d35d6927c832d8f9
zc3eb5b1525184ecb28a425336f186991419c3fe74e47fb05d7b4cfd558d118958d25a657101c9f
zc1313d1e8faae73adbabf55c28e0ef84776abe6a3fec2e90aa0635c21c30cf7ed71753dd4646a1
z88a19a56b1df6ae78479347f3de5da714498ed0314c07ce04b7341bfe9e621fa4b6be901f9301f
zbddf02a841b3a4880661e979238a2419e360a7f1f6bc0bfb98321693f7f61a6f300c31f55423c6
zd9a28652380f75fdae9c1dd08b109dc7cbc030e551f5f3538c88ee1715c2049787717182efd082
zb69191f74121638cb1264e44b755aa66986948437e62b07d39029a57f812d704dd488d7241360f
z66007cc3215e1d19c04c6536ca1129bfcddc2d0d53586a53baf0b38b06b168aa274b859c4f139a
zd9203bb0d20c347c2c487ca9482bbeca35b798c6203b60b4d99a23f5c018cca07292fbcb9af9c8
z76e2348e80ff1a056463b917006cf8c6260980a339fc863ef865fc14144443f0fd40add1c70e4f
z0020d773b060542e7ff464799f088175d8dc509892c6b84f778536f40854786de68039ae1abc9e
ze58523038a8c756fead0de1f678e6ff6bddc9d3521837836dfd3f1705da627aa5184089fd0c0e4
zd8155425cda5927a5d3903cad5702ccdf26185489c8bbb49e7ff497ae25443ec8fb6675978eec5
z6cfc5f354e1134fbe909ca86379a160c104a2b574bd0873a4ba3f2f9f3d651c11dd055e1afe817
z6a80dc991905fae17ebdf03a2d150efb84e1a28a980c8fffb96c62b860fb05b39bd1c500ef8fd8
z6137b8d0e50ce59e44ad5f832fc268844b6222799807b76428bcf0b3c6450e85bd1902ced7f14e
z727da167bcf54e535cfa247f63e41792b94852a5afd5e732829591bc6b7e484cb39d549ce560ee
z0a9436a72af13f19156168a408adb42f002ee7a19b2b0f763cf0fc5f0a98b1943d874d791b04d5
z69a0a462a5ea564d27a0304cc7194d24702cbfc5a7d900843dde080d5ab632aecdef14a2e7ea28
z9d495e6b59fdd9a8aa499b7ddbb0545ed609cde101b83a12ee89adc89fd56f004a86fae771919f
z5ed8e0637b3664d21918656016ba089c1df704f68d20e85894cfe229fd4b746c6d452fce989c76
z32c80de3340cf73553e313683428c8fe42a64fa6a004fc05a55bf3e3f550137f1b51cb26b1dd90
z979a61eee100da21ce9865bc8ba079a443ca1bb0525723db92539ce5125a8b0a4675710f453e87
z1307c01e1bb736a3c92e1f4e4a38b60aadfe6688d0e06b585df6e7b3a5998fd1b47d717caf8493
za1961d65e31029e1f29ac279cd2ac663372ba388b997a8c7a9a656c0eadf52c1ec9d5335255b65
z8e1880fa33de780b653992b4123770360062d472d9ca60bb664aed2910db56620abfbdd705b921
z8066eb6907dba22887b3cb85dac0af6fa3081cda9d99d45b3648990695d8643cd7a92807dce7f3
z75cd7e85947c9a06a495c6b56533383f683df0f9deaa7c871c49ad44649d5c0973c9153a93ee6b
zcb5372f75fa5fe05b5c5ad0a68640b691eb5d32d10c265df0e25ac43d69c2721ab7220482fcb2f
zf4fadc51b91bf1965d606604c79a2dcfe7fec81413c068e30e74de092c951f74e13dffb54a5454
z79bf63a5c896bc3c86a1b13d105bbb4b4435cac981613861dec0281eb788ec977d54c57ada573c
z3579577703581297aa519d6633ec93f1e8517b4617df6d3c0321bed4b38ee3c54e5a391c9a980b
zc45cb9c6df763c8fb7e2b97e44ba33ab2012d1d545fc23d0ec4e246d530f7306b1a9a2622d4030
z2890190b37f7ac393450cca4af94655a92db8e7f5779be27d88b11654ed9df68d2f87c24126d42
z5f95a6e39758617ed0932a0bd3d7fe427d894808fff5d85114881259a1a069c5eab99a41a5b951
za1f2abdea9b0d049df3145cfef8ed37484abb6d7c34fb2a593b555232c56693fe374f28bd34381
z82fa406668ac96ebb898b9f2f2e856cc36d2fef8f5eb7a48f01e984ddd750640cc613e174b8587
z6e85d9e11e16f15fd5472424477475c8be1fe0c7860a6b8cfa35726d6fbc5a4b1c5063e75a5e60
z1dfd86887ea53e5b32a540e5f6ba7aa5c79e8bbff72fbff88d26d7c7f4c903bc77adb4328b1b49
z8f0293232008dd0a58f9a9ff6a5a77efa21c67b39120ed4e4ca2db7e7798fc88708d224b6e6bb2
z343a63951bdddecbaf69d2c48c2830dbc803283d528130f21e0e55dd86cc9bdb964465510152d9
z04e1514445e0eed42f35680ee5b6852836b393466bd7878fc651184c307a3042b3ed5d6e9f1219
zb97dda87275cf0c0b6297f4fc21aace86592986adde4dc28a93a4adaa541439efdfd9ede80f891
z77735c861fa681b33d4689e747622cc38b76b9c0a0540d789d13525eada82b4bb8bee567690e8e
zb3ff20185edcb4f9d4df6e925700a18d047ef4797906bc0a981844cdec6000ceb34df4d333c4ce
zf1c191b6ca35381d6f41c26b6f153103d0f1237b54fb0043b1f7f0067876c6004ccf42fc9ce3af
z05871c9663f921be1cf28ca7bee64c1c40559a36ded0cef8613443100c075d69ee37a6ec74ff4b
z95c873b56231e671bcceb3b862ab77efeb1cc51b29e594009d9b44e8c2b2bafa229acd5809de29
z7f44b91afb604c9e29f42f4a04355e9b1409c2da473f0f7e4fa471b890acd4bd825064cef76ea3
z0855ee89c24e18c736f0f3dca919cbfc92c1b79fd5850c4603b5f28503b352c7910427d8ac056d
z0207b9ade19d5f81e6f17113c297108378495acb61bff1634f92a66fb54c68bdabd3cf6d37ebee
za6ec10d3bc7a84564d9077238739b657093017e8119a1da47287c17dcdf8799c19b635cca39f8c
zad53084664220735e29b615603381bf281f2927012c35db617d6e3c05f7e180e5468811e359540
z9ae0b013f27b7045e7c438daee1829d59414cadc28f7b4c7b69e00f2b5c092afe789f1484e0804
zad706a970bf21e55640ac6ef93d3233f4c9bf18e4336c914ef4a42885830888d54d7f32cc2a598
zfe23c05e8639600ccfe065675f7237afabfdab6586bb03d6ac32029d570e0cf69018fc3f347f49
z04af9ed8e71690193f75fedcc313acc07e3b2917d9a7c75a83efd825fbcebe44cbf7b09f0e121b
z5d9edee08e52ddeca4fa875b0f728c3ecf997660fb4e10c99a087b88e3e3bc22230aa0435f49ff
z678a11e4179e8cc8757ffa9b911068bbf3454b95d443d684facd6dc5251527c2611c4ac8915add
z3727812701e3ffe48bd5f825cfa6736c85f9d1bc16eaf3726ab52b83c63407d5a44abf5e98cf6c
z0f95458ff5fcc46adae8d7e088d508c4e70db7cea8db055a68e79630f66f95b1d48c8e8003141a
zc5946015748b8187da085e8a85374d01b36c7f4f3311529cd24ec92749dba84755e1a6ecfcf927
zba2f3a2c906c9105fdd6f3a60a7ae23d4a607b799536024042a2050e3f2326075a638f199412f4
ze4241c855dcf956802cd6defb63a44dca4aaf0573929a8647267f7dd214cddbd80e0a55a8b210e
z13010678506831d9215ef06be0ee3c05ef59f7b942e9216486e49fa7da3bb4bfc2f608be9eb372
z4fcc3dc21232764dea631e50c02dd1dadbf62c24205a28eeef434514ceecdf52249945b88db60b
z3e23fef42b0a741f3d4336ee293f435957e9a4f97afe4cdbd8e633dec1ceb6d787f875d89503d1
zad656f20fe45d22c87045a3968e2a3b71284bd8c63c8e645d960adff549681f38e84ac337d5ec0
zcbf8f3129a9d70f535d52e925904093c4e3a885c6b95864ac2ba4c47f5a959c4cc2c685c432fc7
zb845a72e0dfe8a97f9f96b2d0949aaf374b7a4f2fef49db2582672df6561e3e104bcc7722d4609
zb004e8eb06dd569f9ed49327c54f4ef294a6715ba2677ea25ad28340f090d4857188916a434c1c
z31128669d9848776bd59e9d97a816a41d5fb49cfa00550bf715b0de0bb984e903fdb4084240a28
z54f0b8e6a500a061db4c42a123b5629fb46dd74d822c92ebdbc80d275317e4de64e48bf9764dbb
za53cb7acb592a48fa32c09e10a4d9c8b03ee1cd9b3dfb42ae2fe146daedf2d6008fc62dbe1c00f
z24eb1e3f556bfec83134417f9ed17140e7913b5cfef1c853ddd2ec6980e8276a40dcba2243837e
z88c2c97183fdaf308fc14c02235f37ee9cca13d8078cc49d7f26088a5f975882f0d81a324f21a1
za1769575fb5eb75890a969b8d46fddb0edc4b421b861f941b82bca5ee408d3ae55c3a2e46ae74b
zd94cfe70011a6ce0f0e9c42b82b8429165aa30b2315597c33f1220509af41089b7e6d43630366c
zbeb1674a7c1159d9196493553059e115004cd1c30acdb8ae525a645994b3adb99354438932cbdc
z87386596b76153bc8e4296cd6c577616021455b9540d1363ed271aea5a8c0889a7fd0048753ff8
z7dee78a1b1cf3a60c47eb4ffb3f6cfdf3161f364c5d3dce12f60e3a5d785853ef39241c1cdc86e
z2b38f4ef1ca7168c4cd474579d35525cdcb086327307318da9ccd695e6e52c99ed994a52c36c6c
zf8569d5d156922dfc212251f1e0ffe0f976f014609ad3df87c27e477d40673db29808ec26a31c7
zea3fc5e87c8126d74a4b117437eb8f524e69d8665bbfa638e7ae0e04c3dd813d9408d7eac1d046
z0ac04b7c40d1027afca4bebca6ae44fc153c6fd783773dad7d86a597bf04ba186fe5aa79f01dfc
z4e3dd75fc4e98ac8ced77efde11fb729e3b1a8ca2a6ad74ce798df40fb569e79406c0f628a2d54
zb74a90647d30a00b3f775e0a5b2fd940fd3b7924682c6b948a4daa76bc27fea2fc72b78b9b9362
z7fb5149c8e235f5a8ef63fd8e755ebc3c1f8b9b8d3090138cb32f33e9c1cdd0cb774c4f50e5c53
z6c469921e307b1690411130747103efd1823244e55bcea0511e771d695875100e8e6fb802f0855
zc468018fbcf43aedc5476800a826f8767dfa72e778eee8cae8edb8df337cb2badfd5bdef6148e5
zbfceb04496e27e29f6157014450ad25c41be430d71dac9318a220136b2fd0ddcb6b4cb590faccf
z17279b4ca045f4874b1523eb0a41b4c7becf8a893761dc1ee5606a9fca00941e844bc446e20abc
z4c52596ab7ead14185164e70852e059cf2d365e5a011401ace4195d47ac5634c26f27c88aa7d3c
zc37be335a3463b4f2c2df0ab2c7a47c0297110bc4abb66c3e9b1d2af73da108b909cfcef5cae3c
za79de376e0f220e76e2bb3e547bcb48bf54aec7220e24ee0d5912d226d7fef42948d78ceabaadd
z0c9d212066a46748487e2b2753fcabf49fee7bd7e6db3bd6143b3ce6e80c4deed5086853a9d110
z2022aacc6b8bf7e54e93737dad9744c57378d9290e5fc1c85a865ea8c1dada81f849603291c026
zfe8d3f1ade76322979d51386946bb71a83025f41e1efb277897b32c4baa92c2f1f8f87f03cf679
z048eea092a1e5dc2d3989403fd06880289695cec8bda004a646428e3a2e24f6c28a69c02c702db
z66017fe6b1330b0aaeabf7ff4fc1586bcba78e1d2db01d846bbe393bc8eb98675c5c4dafce5389
z77c5dbf0f86ae53ddeec9854c8c04a2911a10d1efa9efdafd5f99b74e65ee5e71c7953cf6744c0
z456ae98d2143f6143d332b5699788dd0eed16ee8602112ee7ef62010821966fab627dc5fa19f74
zcf6764290c6c509ab12edbe4d56c25da4fba62f8ad8f27ca49dd9d26d978c762da6ad59bbf06d3
zf8b2cbe5c2f4b64ee032e467059e56ebe8e25102330274f5658719b6db03281aeba65b4632b3cd
zb6b466cf224ddb10be8c709fbdb1d8005ccda6a53e287a6310fe0d7314e5b3fb7c5b46eaa309a5
z2c54508afa54af0ebfc9312d8602e4d7e8d540ecc193938ab8a092f9e884ca05f7a8aedb58b1d5
z46137eeecf41c582cb33f386253e5288a54ae1710754d85ff4c452bf84006272c5635f4dbe1b72
z76f77176d90f484bb7e807d317b44d7b89474f913207fc9f665b79845de0017422c51437dc2e95
zd0db82f88dee2d5d8a2ac6521b4b5a816da2b9767e1bc903f1c05c4b0358a91c75ffc2171ff4dd
z6cfd347db83aca7ef74e08a3693ce7f038456e06b226c7b17887b67b93c9adf08db56664298c30
zf4ed4210f1b7165e352f85fff0d2fea66ed564c2f4da85099d3e316443f1e81d54a3b0b923871f
z08ddf96d350b61bc8085578237775134a5e9f2ee4d01bc6ace2a66798ec1e4aca4163ad8ef6356
z68bc9f63cf3a7d1681c5b025ed99d134c8d1a527a9ab72edc02e92e81a4685e7c7ac9f32adb89f
z8349ca18ed87c0debac6e6be173c1ce2351e574e6a6c190aa0f85dd8e15c6c77b3717a35120fb9
z7fea11781582c2518f992c0fd79a51586679810101f4a11b9021a2d125f35a72db43d07c1c59ec
zd1c47a7d729ef967c635b1c9dff4f7e05f40b443a57bef6a7a61339402091c4388b2a7ec871f53
z0d801bc45c3247b586c09a579670fe39d9c2b552bef6d9b1db6e8212946ed12d0d015d8c4793ba
za836064a9488e2e4006632755c3527d616a9d8cd8dd63cf1aeca78e7df336a385afcb4bb4fc21e
zeb4326b30ed6f4e7a8e21fd9430152d326251f9134e5ec1ac64076086017d0735b78bca1e5233e
z86839fde335204328d8a03ac75e7e593d45660c54f008e6c0541bf4551f6822b30e3af6e818286
zed29ec65cd33c850a37bed38289056547f9b4bacb3aee6d0285283c32837428eaa0035964cb6fd
z5baae75b60ccc6eb5a7167096eb6c8ba82a6bbadc4b6582127dae2037de4a5c83d682e4bba9b83
zfbebf567998b8eda179f9c4f0333d7d0ab0867740a08caf7f2c7fc717e001424c6489342fb569b
zfef2ffe8c09c49708f5e8dbbb955153b2128303ee2f88323a7676f8f0cd14933faca3f6384cd6c
z71a35171a04ac5c64830297a4cedbed0b9c52b7526ca5463046dd1560ed87928c5a3b874951aa1
za49aacc6e640bca4f4cfd69c54413c57224ea3f81c3f9a2f24523105d65a16eecab514981d0ba3
z91f476cd7e73d943936d2e868c363ca94dba829f166b4eb708872dc9eab4f34c4df84dedcb5e9a
zec23f3b8898a6cb9ca454b2897d3e055f81465aa862b5976f95e9ebcd274c4d44baa5c85aca260
z943fd31d47e52e86b295065df08042c9841a4530963118bb48bccc019b498ae5531b02174bf2ae
z1dd1ff6045dd8e100ddb1f700e166d3dbe25bdd136c46d5ed7cbdd1aeef1ca11fb7c494938bdcf
zdb766a5edc215d638d40ca59e43123cb472d83c8560c1ce9edf626512b3ccb90a621d2cc003374
z93768c9da5323557dc8ab1cac467a0e6260763ece82ea27b72cfff9f2bce38dee3abb7989b8542
z06530e74bff15578481acc45525b23fd52f4ead7bbe1df0da3cab8b25414131238b167b92c0cea
z23a10b016d14803a1318ee6a70ace6c1d8893b5f7f5107816366a66912760b2f586a69585f57ee
z7df99aa069e258b35361ba8ba1914fce1397b3843437aac08328b03b9414a24571530aab948c34
zf1b90c8fa70a5ae45078c7ad93dd21095fc92eeefc69c399adcb25704d538c4f8950496d7005c9
zba0cda9b9cc113591fba00edd06ac13b69632fa6b7832736d45ceca8e2d201dfec135bcf801d36
z0ff72b80b9c552eca415ac6a394b2b3c39de81d4510383546429cb618a28bf8000a8e555e53900
zb286081b78914e6ef40cd2c32f31317704c53f0069016f1c1242d526f65c5f82856b2cfccd2cc6
z6d248151d0ef018fcd7398969a5f358bf65defec6eca795496cf0a0fe40aa32db120ece79b2438
z2ab451a5cc57a82d55bd6d40c1573fa4b5eb5c1e9294c20b9912a7d29197e7ff168f51fdf71936
z20d5b77c02872876252452a8020ce166f04e4c972b54d0069228e6d60f477f4e2ef06527edef48
zf4c5aa2762a64ef084a6570eea6ec59ef7ca9c2f4f57282e04634a5fb22143a5fef61d7f9a273c
zb933ae249b4b14c1eb8f3c8ab442509b1d47bc0b1322e6a9ffddd6e7495bafdbd6901f0aa03ee4
zc56d83dccce0f2664a783c2907ba66b1281e5dd9181c960215ed558ebccd4c6ae72925967c5841
z2d6085f16b127ed10d2cb176da152cbc027fc4c9fcac4fcb172cb9faa47938cdf33c9f9cedaca7
z5bed68b8b40dbede256e72bc9fadfd50402d19ad5a16df4396a28d958fb1f2b1d61f9034c96469
z8eb401ed2c0967a74fdc8c9cc4e4fbfd030f5e533a67058ad1d111c727ad2409e718a037920a77
z4b077d35a275e15ef434df824b8788be8fb7d125ac76fd4bd64f5a873d767ddb1105fc82f347fd
zaf82f3b4ff318c75541b615df7fe322954e4ae8ef5379557b0fe4079a61a51c458c84cc4103c93
za8289c2ea16282e3962f12538fa09dbc944e967f25f1920217df198bf6a7fe1c3aecffdd7d0c42
zfd4e624761330b994b81a8907fff36107a0436e66a2416009298978e84a3352f0160a1a15d1000
z0f66e9931c1fbf8656c6be28eb3c7d06179aad722e2ec5998cf0a42974b47328edaa37d4bbbd81
z171b887c828fd23ccfe99883e343b7fa6e59a4dc81ad73a5417d604c50f7c3ea7903ac68e3ba16
zf67438518e0bb67518d3192944674bffb54543352c51f93561bcebd70c48b4200a093158b46073
zc8bbcfda61204b42e1ff77c16e046c20f01ee3e1ba16db8485fbbdffabf89fdac36782ca668f7b
zaee0a75ae3c26ca91903aa7fbb7bb93449e25efaabd2cffd2988abb1968565674169c8d246a07e
z4475b069549f63f827c3db6698de7f71d012b1669c8b2421739c0b35b8965435d407a8abfb5418
z9cfa77f3d854de09755678e0b0df9ae9209af643b34307bd8499b4957fc4475411eefedc18e60f
z46d8aeaef7b93c5f01cc163f68870429b331fd05666da8bfef56503a76269f17db4db76d7d48a2
z962c1ba7e09730531b371fc2ebe81247307fa2544768a5b68d73ed2a21b195bd90dd43ab1cd154
z255315305b6c55fe8405d8cac5fb2a5621297e016ba213baf5ebb5c70eb35745d3e58a381b511a
zd1a5e9431e41620b0c6aecedb80a2c9ba84146ca47ba06b23bcd8eae4d6bcf800e088f9a467fb2
zc9fdbbc6fbeed345cbc02ccfc065cd3a18724cdd79800241972a77d66228888705c2d732174c26
z3aa6757c1d44ce2e504dbe57f18b39c5834fd5e1c0535b0a9b67210d918f171e722a3f25588feb
z61481383d98ebc8a560b967c78e3e3aed8721822fbc5bafe608ed28a7b705944c02edfbba33286
zacd8ed59a7c1eccc894413a4ffca87795a1f39c74b40355dbed06af608fa35c69abdc68344d49d
z54161e884cd6e2fa3b19a1e3bb93e2c2412608599dc1c605c1428f5c75a23842b7c66bbb38544e
z1a90a8bf251713720a365e643b04c50d58ebb9f2c3ee1c073d1b9c9fefb181372485ba31217d33
zde12779974ae529e9b55cc53094a281bdbebe3f789aa418070bbde5b627041d65bb650485e6edc
zb846b18429b39c9699b4d5405ccb503b254490014c227ac3141855b24645614d1ef4ea971594c9
z9d153fa95c1d77e37f20e8a1892b2710c6fc8b921959e520d12c138082d72f778458e46c0a1c18
z0d407f37778c9d0f1a316f5004eb83f25ebfdface3c39a36c1d1cea7ed91522fa1b0479e8b8829
z1c64f57e649524520a3f92dbc7bf46ec8d0b31c586d0b1280ac80a3dc8839b36dce4eda4d42fb2
z9041f5072b57c8f071b6d901f6bdc5dfc6f20c167c63e7080dd23d2a4662ea00c05dc088cd48f9
z7668278ee9d5ec3e788c76751e25edbf9f4eb7cb521142286af79613789608da741ee48749be54
z1c9c5f1053c7221a28c0e5a3559fae5d069179b3fa2826e60965954245d64af6319a0f5d372d26
z30d52d3c2d2b1759e3f40e76c16d6bec3dda1c662331fba02cb6172b3dcc0fd3683e2b7d70e58b
z7da6ea26549d6de11f43e43724e30e70532e796d8404cb37c5572df01c5cbdbcf444c47f2b2021
z32ae0ef69905821e98aab50dcbf00ec75306e7a5f0019ba45c360654ef67386a59ca2a448fbe9a
z7c31d8255ec9d90908527ac3705915dbd2dc7782db292275fae820a8ed1f7f2ca4390d02f74c28
zd32fab12510cd33133046dabf73784e967561d569fdd63421e3d171b2f2f049336e8a352bd7dfd
z4794a4d4159860e5f751c1cccc7d79bdc8475bdd8883e997db01eac39d298a0431090f183f650c
z5988ed7d2fac129a85f4accfd7263a3227dce366c78db215da41311f7d2dc1762f5c50c848982a
z3d2bd0127563eaf18b971bb157154242d0c8969d4019cb0b50e9634be5957de794c283f96126ab
zdaca3a4d287de7412afe79ae69427185e5b27114aa52a8b2857dd203f363978a3acbe13cdeb75f
z6ff9aedbd03215b00acdd58e825eeb1a639effce08bb3c65984c0dce41f8dd1c304739bb7a6986
zd57cd472fe557c975a1ddc240f9c854c59c6b2cbf00b5eb451b68c5464872756d541a57ff0c30c
z1f392ef8d6a9b48d281d7cdf82e817e261011855e00665046513b11de765c647f432f8954c2b26
zf7b003409438e0073cdee9cdd732a5f09cbe9d65b817ec81b86679ae431b585fdac064ab177934
z56abefdfe86cda00367e8b2d66daa934680600897d7c978cfc686a3ebab52a0aa421d32282fa4d
zc5e59d69b4b9a34e1cb22199d01dbfa46f5b93427475c566b957c2a3fd0f6bdff611a3af51cf36
z88cdc4560df1293cc19e0e6d3c46470e2f90e7ebae16d5af3b039281b1fe8e768aac791232b813
z5f8ea1d8107c6e87b13845e366716ae39ab5c36e5ee3eba444e6ac28842562fdf5034410faf67d
z103f505e502cda52b70cc948cfc0b35807e712bb8b731597416bdaf8db0cfcc1dfb072ed537a12
z77e7ccb85450e30c994d5f47961e4c86bc0934cd41fb9ae8d88601f6bc0966d44e22ce6bd81f8c
za47282f521258e98091b0e0da84cbcb39ccbb4f9eab312ef77608f2bbd5f5fd2f3fd73e3a9527c
z3b537c6669f2690983d2c5b54558a74327f3013c635929b2cdce5e741ed62e0a008dcefac4fdbb
z036dbdf0a8129567aa130dcf7b7f6182b07462e28f5d944bd86a7b4443c7579809b5e8dee5aa48
z6af850330843f0435e6eb09b8bdff60fe38a1526e3420754d65e2ac4582fca512681bed0bfbaa0
zd2cd343761caa9f9d7cae240e544bd5e54a0697f8bdc8371e70fdbdb81140d80ff2bd6f38d6cdd
z93249bf48e1f31fc802f9d8c1db30dc5e5ca6bcd4cfb68b1e42bf4957db208a03233d6090a4e9a
zdb9d87934e05e61d5f42deba5c309880f28733de8bd1f1384c76b731ac4061e361700771460e72
zba8a459f25dbc061a7fa47357340b37bee2157485891c9d91e8e68f7616727e14601245b2944ee
zd3aa952ee46b1c3aae3638879d6ce1b96cbd153fab2c4f09a99494eadf00ea6216da121d161a11
z688c18e7484ce9cb527ec19aa79504d32f183defcc6b66706922147cbaff3bd07ae842d6a71adc
ze95c699f8b6c2e3135f0299336360d8a102c53370b12d7057e571022fd13f6499d7adb7816c977
zd320af9defb5ccafba69accd309cca098dec708ca9d538674560ee3a174628350db8efd486b86e
zafedd3455b26c8f4b00bc84193bb3d80e6bd06b3f21a947b77cfeaa0260da1a99d3ab54abbca5b
zebecb968835b200f346912a234de14c0fd759f758d8439c24df13dad5ce0aea0b8a06010b432fb
z987331cb34453b42c6a11c9555a634631517352e4bda281497daf2d9abd651fdee86304eab5876
z40ec34dd0e129506e649124332094197b49427adf9046bb9a390acb0e8c8abaa04a64c27887d31
z63a93ac2d726a00971027003a573634a5c1ce5a4a6c8d8718722d5c7d2078f4901288fb83fd73f
z34eecc428b99dda4fbca7c60b5025d7854b5654ba55b296c87c704ac7cb91a1e64077833ed63f8
z6c98d9afbfbe16b0dec8c743587765960423f20402ff8c6e5132d85ec52be7ae553a9327915528
z0d8c0536bc5256ceb69237b7d1e603c1ca39f3aa9fb35d3d6abf1dc7f08dffbb567b2a302be3d4
z052cedbb25155e99a893cf1524725500ca9306558c34fb78319b2e052db6a5024af8d40b2da976
z3ecc494bdf630dc4959bbb170da1350acd6ae0afc618c8cc58479a5a97098607f6d5dcfc5662b8
z9fa72bc842e7a32c18335a71d1af1c885c4bf7a556047146b48f7b45437f6e122f3a49db8498db
z684b564feed08e734edf97c3ab6319a33d678106e699c5031b8063cea158af234ef9903fd49d78
z58fa5b31e15d82cdea0d9e7a5af526d0ad05cd954706340301240a0596497e2f8f35ce8da39817
z8918aea3363f4dec1884dd62deaf4e8f53124badbeb259faf87d80ceddf57970fc1393af332f88
z62fce301496312fee7cb479d9e5f7e96bf8314f3b5e761d6f891d2fb33a086be44bf1cbe5ff921
z590f4b1d7206d8a4b6d1d745b2126bba9b1d99984819bf1f607f7b15ef53bbeecf70d470fcbad8
z31a4c100e39d01509ce724ac85b98246bf03c48b463da2bb4ccfc05b5237e79223f1b7e7878685
z78cc9d9e4f94b032dfbce3e863730f352b6d1253c44d547d1cbffc31ac65b33a1d6e1ccad9d6b0
z53a9e0e0bfdda89b539a29431ed384021164f5b6db8bbda521ae93a4adb8f64b4327960e512acd
z1ce86634344940d3e4e7f6306f8571a8b85872bbde8942d7f757fbe3fe27f73a24a772923edf68
zd0dc3cd0a6e7420691790405d1457ed8b48eb6d5d050e4ae26bdebf16037fdaa0b91b73cc8f38c
z8b5a0de6ff0642fe76bcbdc988d4a1dd896a11c74b6d5c4f1f0dde9cb84eb53f07a017c3cc96cf
z5d0e14a29065ba85bca87436dfb0fd48f762a70a58050c0fbe902cfb12c7e784d7b2b66b06a545
z6f7ae8fe9cf9c3f13e4185efc08d8e976660b63dff81ecccd6ff109f992b5d8180a12a1276a87e
zf5fea6434e2e4e11a04e21268330054702d1db92b0aa549981b7cbd426e729c95272d8b2db8e7d
z2aec876e77b5a0e9366dbf183f265589bb0c229a028212484e6c7a2908ce5e27cb7561cfdd62b8
z790c676a9385ee47cc415383545bee681f53b7fe31b2c817a0e1e25505712214d66fd09eeafd0d
zb6c1cc35c3b69bd81d78ffd3e98e313a103a9c8a797e51292956675fe31ba3ca8bb8f8b7df8066
zd992c212ef41ff9e65d4bc55ddd0bb0bed406fb55dd1cfa107f23592d6e76f80e38242e3218408
zb1e23ab21e4dca8a241d8010f123544f19179c9296109794539cc4b046bf64cc1b4c0a3442024c
z1f7ce3a5e24ec40bdd2b53eab48a9a1fd3e4dbbff8f01357eaf8041455604eebf8542919d9555d
z881abb320a7e54b04b221827afd968d76d38ef1b61e5eb94af3dc13be653c219b72a6dce0e42b9
zfb5445531b20146dd0dd4c37546584a0c841a19d93f167d08f5b06d9b2ed11e3986f5a42a9a1bf
z9c8ab69a2304f7a1e0f531f9e04a8e6b1bf049c15702307daf3810993d8959cfd10b57a91f99ac
z348155b4c2ba2b54fd575af1051a7d13ab7375ade889e07da65557fd09650704ff50956f6c0c55
z764919e6cfef8fe9b9983cc98a9d37cc92b0f129582f98156a3b2189c12eed12ca8a515f4f9000
ze168df16705ff7021e164c743db83c636c2509d5cbd20f7fa9cd86b338b63ab93164e37dbeb9c7
zbf88632a82564a1b2de860e11289cd43d80ebfbb2e504163f0aecee207f1b0d64b6f1f94babd5f
ze5a0ca590b00f406f0e431b9b52a85a35d34836bb565905a43101d409ddd90c064c0a33c0c6646
z80a6045ff19016475cd6a33a5744b86b3e694da9eaaa5e59ea17069292816b97fea40d21af199f
z45a414f4301f453214720bf1826b3cd28abd2c326ea24fc635da5f633b015f953cb407a7b5daad
z3532a93f73b82176bfdecaaaeee80cd1877ff52728baa9a1727dfab2eda4d3bbb501b5aa0c2a1b
zb269ea9d6007eeba5bdb2d7ea4320458cbb8db7ce4b2f9be32dac667a9022716db075017bf02fd
z32c28c438d705e86c58f2077a7e791ce8eb70c37c9669a0a07f1703063805a6d24b50980b50bb9
z369fb4383fc3cb420714a5adeac9cf40fa80092167c6de9cf2053e27853d3a16eca41b8fd5eefe
zc9f765b9703b4c77a2ff9b88492dfe08780a7b5acba4d005ef61d834f573f2098c64b805294615
z111bc17f4bf18380b640c1da1664c76658f809b209a0e1b061a80c4681dd196a32aeed4a1d7b72
z7a61408b458347104a8330e35c587087f119413b883b5a8e8e6ed38a6ef9beb6714c64b59d0b38
z1a0984832e8d54c715e12702d84ff4e2e62076184f4beb94217c5a9bfa94e9ecfd3ef3ae17d2e3
zb91eff4050f71a2d1bd04aac498bc8e10ef73f1064249dcfa8dd4dc482149a7f0bbc9ebbf1746f
z4c401b30363f87b8dfacdd38c76e7623bcf6b8a3f3f649f790b880c28f23d6347e11427615e866
z821c8b2d6120d752d24a6420a5eea79985deb4dda0ee70d91308abd4578af0b4ee58047d6b15fc
z7ba3f481c7400758fc19d62a4acf46f4e73a273e10dd47a94528cdb6155ecd2499860197e5a750
za82ad3039853bebb21b7c2927e066c55a95aca4e6c54a6af41e228cf4aadf34e0786bd2812f741
zbf76626a19645f0308a09f0cccf199905b43452d700a57fdb3f3d206f1bdf627d7f0217821482e
z065ab4e535776c6c034553550cb2583250c320d6cbb9b99ea35665eea535afdf4c89a2a68ad4e3
z45347ff7c0ab4ac728dde89e534012f556abaebd8ef3eb4aa4f42b2516f1929fd58488e949efff
zc5a9a6e97f44e867c2ab00b97503cd2a2feb77f9b6ecfd1dfbf0cf7f07007e318c0b91e561c649
zc77fcf167c7112a0899619b75298aca8e1785879924177edf88804b7fd0f444af87b6d4cabb1cb
zce34f1991980503590b0a8c57fe75d6897d5ac1e713199939ade6bcb6ad9339a8c4b1f64287410
z91276b78854f2006f3d188cb94706878ed7a1098ac427440c2307a6b5208b2673c85025b85b4e1
zafc9cdbd052425dc12821baba494f13dc458f8b8ca924f59e46f11f58bd21a5f5c2a046c1573aa
zbc555db5444ede2482e8091e75a0133595d6968ec1532b8d466b3e74669e2d37efbe21f767d7ea
zb602eec7f4bf2aaf5672bfc30c2d4a9bf0e9023bb711ec9c5b483a42ea64bf5b1470fee2b50937
za35fe1a3e6c9872feccf2ac45fb8862e8d94018f8c3d5b2d82d9888bded2520c434bbbd9847ac5
z93b9ea7d948bab9cdaa93a69d05649cb5b683227698b0408ca19995055546c97fb6863c28819ca
z16f429671b9878695461fa468c5c709dd14e09e4af6959397fe8efb20ae8a44ebc852b493d1d84
z633b83114ce8b8712faf36f053538e83d40f69dadfb04d2e9e2936abb43808185d981f511a6d62
zc287b3a9551f49a60f42aea413e6df8b52fa9490fdcecb6148518a09b017d7a0a37621aed4f4f0
z0aacc8bad40fe2ca0e31d3b5320b6b64fc17c775de6dee1caeaed33625f056720a722137563ced
z4c3608f854eb7b16d1cfbf63eaad160d2521090a54333bfa19c69f9243f3d3506df706b307107f
zb88b8cf1917670a559c5620e0e75e1e3dc6f019bdcf0ffc5b99a51bf0f818bc688828e70708a77
zf73b3453dbf21807659aa7cabca0d4f6da8ab4345690a7f07b94df53532ea5b88b985bcaed107f
z6af22b9d7c5cf67d30f0479e2b1c31c4ed490451704c9c0832114ab1755385d157a3d49f9f4d7c
z6e1e20a2592196866e209eb7bd2b65c0b381b234f666cfd7268e613892c6cb36b834f240a6c409
z138e869627b3f921301118264ec6ae7d40e26975ca3bec24d4593c5b1c2cf38963e839771311cd
z446260f2f3ffbb900abc83d8383b719de0161d125c958efdf8f5e32b4bff00dcab4c7df2cf6cb0
z667c9b94c3b3de0552847bf16769933e7377c49a597fc9b6c08e6ec665d1be2603fdb14fa12137
za237a316daef68188dd25fac1fdb680de4b298a19ce46e3fd202757ee25df3d5cf0a28b1acaf15
z52f2c7fcf66b0e098bc0ff283758428cd7f322950fcf427aa3c69a719b5f99e9f6e8881e69c82b
z648f3219b2ebbb82d0cf59290d1cffabc2af3275d2de4de682b4107f26741b4f573fdacd4f3e07
zc01b42551f9defc3e24eae120158b3029341d15ddb32124e5daf0cb75568ce4cc247ea56daab61
zaa5dff3e3d8df8edf273919a546fd1159906b85fb6ff2b79859a7d891d62e8315995d8b6e7411d
z4ed82ab2247bf764ad85c47669c97ed7a896503709a058b2c59735bdb8770b23325636132203dc
zaf962544988c80208cf98da3722fc398e6adec1a19164e575998d70d91de863d41bc389e4123e6
zfb824630ee7e720a689c1bcfa0d71144b431fb8a8d96f28d8a354ccb656845f870558dd21528da
z030b67e79b0c843430570ec67256084293617ff05418c47795dcb3d7e2f2043cf8299be7ed894a
z1453d96edbbd367c7594a924a5c9932a0ac14573798c571330ea84adfde4834b76642b9e68ab9d
ze7a21a5dee44723c2763ae3b1d40485ce0b2fbbf95fe064f4f28cdfd35b4316429d3b47860b124
z23321cedc105f7da597947a3df241693c01ccc9047311898f858d57639d225407ce0be4407844f
z6dd4b8a787a281dada51556e6931f7364ec95c6d66caf16cc07739228f5fb43e167a50683a9544
zfb79d5b4eb7e3ba58d6f363a397ae02fa89488d294c2473ced18f2a1a9ff0d66810481ddc70b80
zba0ace018436931233e857bb34660d8a891e33afda3e972beafcaa74a965183b87ba1e86e0af39
za661b8db53290c48a1ec3cb945937901da4f68393a266c160efa67ef373926f5c3bf29b9bd09a3
z8c08412950cdd94e661fb75e261da102f1553eb9efacc81f6457860cb85ad86a2834794ff3b469
z469336e7332f49cdff9ba7642b9d073034b9bb8124f2e5bd9ea84318d1341b7e4540347b974952
zda8ba94cf27e57b20f825b7d5d024c4f8910471f9938c8a31b26e3205495e3a0dc8dca343e9bad
z7b2636a790886eaabb144066fe32bc681f3cec6a023133ce01fb102f4f30fa66d5eaf00825832e
z3fab7d4006ff0b4b814198d1b15713af77efdd5888e6bd734a953ff0a3c493f102943b4c50cc25
ze3e7c1a1e28f27b368e1c7ce7207c6c0140f3acbf9db05b2b0c51c7720020004f65f47c572cea8
z79b51ab3a9898a50d2bd32666ac0862ee2cc8d809a78203c67130c41493bb17c20c4dfa155e02c
z17a3c2f9394e80e25af69eabce6373549f439bd3eec4235f928b566a10e7bb80d3774e1884406e
z31b249bfc67801a658e240a97946f3b0195a45562fe799bc4f548da62205d1e86dd9cf6a411f34
z746988cec1352773ccd5860a9e32365542143cdf7207997f7493598baf3e5b07610b39d5511a74
ze6a2b8a7367a7f6af56db2c0d0cb71887ec550181dd7ec28647c42ef7a2d66bffb089ef138164d
zb4244068cfcd2cb60a9c9871c6646c9d2c82bbf576a08a08dafbba4054e9a4df8b515f3c79b283
z8856a543db9778a3889e24fa023a39bafcd65a8412d04e7948b4872537dc6c0d8b451af2c68ed9
z49da5d7d592f4a1af9c53551d473a103cd9cdb92bd27e1dacd5137e1ce2ffbbc09e70ce8653da9
za1a59d7a0b8ed8941d35d68fd41e5088579430b5c707bd4a9d9abfc7ad727e2d00ec21c63256fe
ze3237d4d33ed6fc36c51741053a5d7bd34bc57fa7064fb332c2dc2dde2981ea6b3fe9009f08664
za4ccfa6aa4ca0a234c8c836ad6b607788b9f1ec95d38e4db4a67c491aa8d911019ed9c02c08a80
z1bcfff443636990a4ead018fb4644559777b7332ad6a81f344476a4ad61bc7b4b7f8f2911dbf4c
zfbee3e415a6d97d3ff26e3f3fea59fd8dcd507bd383acb0f6b6428c48c845a65e990ca985916e3
zc39a9e8053a421bb49bd0cb8dc089138b88b14d2ff23008b8a3a0f80b08eaef95dff445d700403
z550f420d7fb8576c77bcf6757c00e7aecb72e681244988a211ccf298cdc14f0d4099a3a1513dd8
ze2c3dc96a4df1174345e7a5e6007e62d744f28213614a90761afbfd8ed5cd0308ac1b518b0a847
z6d6d07124682716c68ab0e98531c34855d0c2ae8b11403aeadae0884f7019484dd5ed3c3b2a2ae
z0f90121578f3243575d61588fc6c02da735c356e0d836cfc9a26c575d0d461f84ac213b99ab198
z5d7ddb600165064588b50de0abf406b186a883c683531b0d86cd07908fcc1c257a516794ec067b
z484ff38961c7a2f28c0e03c4eccbd03c3ec1a2914596a3217af30d3f9495f170d5605e61b9bb92
z5a64919abac78ea2f0d4d2811f13c1c90cfc162fc2866da46d273721db2d41d1e3ab544f3148e8
ze0be96329f52b5c6e98c7e8813d3fb6c4a535e248e6c5dfd05e937ede0da858c00c43b4015b4f3
zc4c91b64768138fd187dc21b05c46f1e85f8d57452b609b82c15ca099334cf1caaadc9a58c3633
z86c43e804fc94b5524a40a4bb917202b4093279f6bfdf7085a56dc59efe7aa2bf8738fd45f388e
z876dc33955d13ce72019a9b84ef9072c13ceb8b57d4dfa997f87c87713be480f50dc3cfac16943
z06e4d376e7822fc8fa0b22d46fcc8fd373255edb278c4859d8150c244fd3d2fedeaba42a4c3258
zb450e2923d7b5ee21139778dfc682d5436a799214e17aecf35691f9b6f84ccf88c90bb4d7bb264
z50ee336d15e39cc7e418b187af44abe0b6cc0a794154daff7b031938ca7ed8ac223fad5540a83a
z4c2aef3166bfe1ce4e301a9e3b10004fe5e00fc9e683feb19ef577d43f67419f2df7657e66037b
ze153b228b8324384c18c23ece12c915597c7945b6d00485ba5f93ca667836774ee7e5e817f3bdb
zd5078562e4537c0adfe8217eefe771056eae76a0e569f069c3988631d624fcecedf5d70091d212
z758179653d9a5850a4eac17ccd964cc5a3ba1ab9187f045e79d71bdb55fb6318f4fa6a3c74b893
za8662e6d63d70783c1d6c7512e2aa572c608f9427e98c88927b981cdf16641f3d16dca55514034
zc5ad64a2228f1ee08897d3768d1b46b002ebd2ac5bdeb355bcc07ec71f65ba7b78087741339980
zc251639167b90da0a74e84a27cc76aaca6087169a5c19c052b6a6b7b29ddaa707ea25d42581615
z2f8f0492521ef9aab558db9eaeb29add42be8c1cf12ee150862da8c24ff9d1ae9a35c5ffb4ade9
z2f08df6d7f7391f68671a323e25e760265d78f355516bf287e407c20be9cf8d4f757193fbc5622
z879985db1e0135b6c447042a4bc62c18a9ab9e177041c14e3c75ea02e19be909c268e052554d61
zf32d22a923efae60004fc1394628609428417f0595bf74f16ef989ed29e29835357c1cde642d4b
za71b688a38eac896658799912c45fee28850d90bc47635c4df294ff0ae3305f83c4f38da1d7e28
z932ad503d226b065c2508f302e929f3111911831135161d79751ffdd4b9453dde345102fb46c20
za94f6af8e6b01dead884c8e0e3f40ca0e936c0018a27bc6319390dd67a96f74a5467778f1a8505
z2a68f8b5dc99ff6b2471e270b27561751ff0c3af3a4321d78636463460629d9577e22391a15222
z6950a005bd4d04db8f0e2fb615419d1ff8898b65b3d45f85b524f956191735cba4ca1f0990534b
z5a56fc36a9daf6575a4ac527d0dda6c9849dde31d53a715a865f1c44dc5056c589eaf2cb66eef3
z01d43be896e60a9dd0e4274922f5b0f5f02d091e2c3478bf35debf0c5bfbd30991eeb0577697bc
zf3948688ab44ffd2d3b58fc7052b51911862758ab0b5b7b76bf945409ce4ee2c3ed937e0099ab1
z65ab10c9399e9dac332ac5d77d7361045979fc67e41a36ec2df37644fa64cd3a063618c1f12333
z5a5529ca422db02bb29150a31f1b63fdd70cc2cb8ad85e9d425f2202bd5b135f5083ab0425fbb1
z6596bc2735fb94ef57ff5cf564508463b8cdebf1eb035e62247e85088417fd9a1c420375a5758c
z0c9e0a37a7c3aadd2f9a94d4bc3e4d3d8438d91b762f184e387ed4232b1e6009137b3a2411bb57
zd2c7a1ffa678c3e49230c12b45c8d38c7c86bd44185539e4607796eef537341d97b372cd42415a
z123f33224c4c5b4116d82e303e2eaf2671a95ef20eeda422d325c1f0f9a1c1eaad3e314064e18d
z780a80955bb885c218f46e18d64faa6dcc158d326ea7f0d6c6311150015f3d5c7bbad2b84ede57
z5a474dab755a4249faf67ce28c6ba83b0f1cc4c73c966c2fc3b98d2f6f1fd7f933fc089a72580f
zdb76ef8669e2c0d62a4ffb23ea09dc121738674d05fedbdf42830c107fb09d1085041c728aba20
za73de46ab17d6b00224fb8bbf4d67d6d359b65824e0d8ab77361432402e0ca0018bfd106a3e094
z4ee655523ff582d17dba3e1970d3f721033e1b90994a979882c8b79a001b5fae6900dee71c0b31
ze49d8a8f6b365a4082c8d39a1e6e5a2ab4cfbb4ebb46e7f35789de3d9f77bb226a6f919d258ffc
z11ee7bf7d568a82caaf2675fbbe8a1c69c25b546a8da16bbe9cbd44071e04d998b3d18f6e1bae6
z7e79a7d0191f3dd1dd05f2bf3088814f8355d324778f9d3f64d13b96434f0bed4a8c8be7cc8a5a
z5ee0b58f5130e42aa91b2aaa4804110a870b827e5915da13d742ed489e751431a4bc9666876fbe
z1996a4e78e380503ea27bf04e0c3fb9e024f8807652821659925eed6d1002ca804d40e3502b750
z29a3a1cc2fe0a2dfa97a07ab8dae049391d0e72d7ead13c9e9487c82520369212c0fac2567ddca
z85668fe445bc9774d9924c3882fac49721d5eb526c6f33a0f19f0a66ba9b518fa5ddc787a0af3b
zd5b1b5e91fc9fb33580bb92d6abb161d1ba494e8d4e77972f5b3fd5cc6675ef39f794aa94aa029
z71cee3de322888a3942901f8b326146759d014be65dadac60703236a9a6112028dc91ac0edf174
z662adb660f84a888065672e1c6e3d1f5475360d0d416a462077f5519dc54b0d3beee8e9567a5a9
z485e4a1ca6df30022d02a4e84f328436864f111838aa6398f4873b9e0c5e50e64880857f10cb3d
zaeb2cd2d7428a00755d67255d6dd795b3d54ee4eba9ad64d0795100bac99039e86b08d2e06c1b1
z0f33ca4d38bfb5da868665291f7cf2f55f232ea2b533ab99966060caf7069715a94559264250e7
z02b9e121ada5d406d5d2cc5c11e6a6b1d0076d52861668ab11ea5a69492420ed9b0d6baf505cd0
z77c0caa37eb056ec866fde29b61a1b941fa527618c6e8b1af6aabf068be82f170f65c3a01daa92
zf494bb7bcab252d861151d1c839da5cbd42c26ab26f81ecfa451652029249d6451bb365ebd6255
z61c657397dbcb2c8e39d1f5624b5ca642c84057ba0946b93732783e016f0d727ed009f495ea01d
z2f21e9274e5e54027ccd1a607e49ecb9308a6d68f5dcd9d8b2daa712cc0e500e1cf4c265ef8105
z1beb34dcaa098efbd6c51445c3d27ae2353413aebec2fd856389bdf338fb8c9d15cf370eeb1723
z18682ee4bcd3e8b7074c74f6353f3aa6b413b0c9d2af4c393ae0b4fa3b108cc1206aa6540d7b91
z9a881e3f3920036fce301a64111a3972d10557810efbfaa3cb907bae03e6ae1b58775d2d5056f4
zfa5e85ba9f31b9d31da7b8c4d513d3ef36eb66c36b64b56a20c3c8f31e38ad00346c398fcac50d
zb1353bd0a1f55480cf70497ff7fb9e25519980970bbef485f076d9756450a61706cab866502836
z522949d1ddac6ef668c9201162f842eb1a6ada4d619d73944d137b33d5e2d8f9e42bea9a94ca53
zf0ef26191a47979d5707ced86c29c335721f0bd97ad1fadb2179d6af0f1aab78409122b4f7b83b
z0793cc6aeceb93a81cbbd6fd67cf36ba88f0615e1d8c234bea33d8af6cb704dd9f368127497bf0
z9585f638910e6f45a49f6937c515e52540c405fb59b737ddbb24c10cdb509771400d5ab0884d76
zf00ae4aaeabf027b78d5bf476c6be90b4a6ed02c51f53cb6cde5332d75c1d906a459579c78fdd6
z96b83b78dcfdcafedcced4ec6e4785d63b1c4201c55db999c6dcdfa95105c38cb76905516306be
z468b88d6d5190fd6b98a0124afa7f70e17baba6135978692c3ce9fe6ebb1a747b8105fb022a136
z3928a5c577956503c969247fafe23f8bc1fae45b3bb83d438d4d76f2d21638aefaa6f160e0cd76
z6662b0b2a5c4b5b5c59f4df66d2a59b5a1bf6586d3391f4968858bacd95bd48cd24681b57c9f3c
z19197e6885fc50ba4bf1a9f8bdf932e9ca780857cc08aef778d702e7bb1634f54996c3890d1c2e
z935dc5f94f0a7475437296f76e6af93cf43753ff22aa69c4e75819a6f2ca2f8a08efb89327bd5d
z23e3dcdab4576b238dd658951d4b067fdd7ca7ef07fe4e3c2dba75f1b2c8110bd1a1f49413f0eb
z172abf854eb026f6eb44e9da5332a27f296386882dae966ce15d9d1b132fe3a47dde8c196a5e75
z66b8cf8bc7876e8ebf2e44a51d7d1f91c69c27627d1e1fad6a95cd7cac9190801b04e68d467e87
ze415da556db4106bb2bc5614d7bfa98720d2254d979454ef164bb71680143963067a5d17d5e780
ze455cd6c921375afa59c3364e42b0c0b7d2932d055d789b88eb63f428113d9f8986f5b03595fde
z7b476d89915cf9f70936733566ad956c36aaa2389d0cb1496643733dda5a455efa22aff79071d4
z098799de154673a3c7c6fd358981c277eb884409b84d51e67a57dfd5420fc44b9317c937b5d60c
zcdb27487c5b4389992a7dbd030d4ab29eb7cf8511f80730d5f403f87304bf00b02772ef0fe5226
z344f83b7934ef962ebb81f84a8313663e398c30f7c82a6cfe690e9baab9b226603a64a03714800
z43d42107ba587d6f0c037cab79c306f65f08eefd95a61dc74c6ea81543e19ad1414d38aaeec8c6
z370deded6c4b948d7d54d03c7a784e3ee0a400d645578969444526e9b5fe9d39235c51ce86136c
zf1747f7747cadab61762679fc259dec46aba49b200374c8b199f63f9787cde33e563e132521eda
zd9d74eb72f94a8a67fef0964ab4f7d2793ac7999f0270d37d4d88202f1ed8e9bc71b9205366dfb
z39c2c6b6bf5ae2a61b3b24bfabc5743d18aacb2cea82409d8b4a7956028735c0814b070cfc376b
zdfda74d0beb2cab2f80d10377c7fc904d2c2488c6770458aad94bf120b3e781e35c4e0356a4b8a
z497a51757bc7c2edf8ded9c034c742bbccb124f026060d08e6c84441305173e7e8dbcbfc369748
zc96d2f0ab0d937adcf9bb202a74c356864736e076d532a6cc9b0bee263ff9b9ce51c0fcd36d882
z8dfc832cc3ac3001fb914f6ca734d965709ffd578a1f9ccbeebea1c0d7ebc4d2c6752c053c353e
zf7306b318175994b8fdbdddf11beef67c5388c9553f84c2580308b6003d630c523c681c40e9730
zf08b39dee6bb208625158dca0f82e8333fa3f5a80d7e4657d149e9cf3199497a9f01165d82c0ce
z3eb934bb81a68561ba081d2cf57145436c03d8ab23dc4eda62cd0f7ae2f2592c842424c7badae4
z58c2cd892f48daba578e37ea547427c5fe2829266adb490834506436fe5c23e594cd515059b182
zb29f1e2231176c7e2d947937dcc36ff2eb90b33ce9c8725c3d24f2f39853e7c6985065c647b41a
z21ca32256d486314f5f1883b6957d5817ca68e4c25ba9027e181891e3d5695ab8a877c1814eb93
zefd239afef836a2390e2056b5a9c59b96556f4faec351b097d22b99f016b78c17da71d86b5c35c
za08bedbee5fc0d53369fbc56670c50c68ff38a3b5dd47e42c365039db7f52f530c0a0c6cd428d8
zad0d6c399ac06798fde0065eafcb2ae3cb621fd6f00810c33bdf6445fececc0a719b19894defd6
z255a1c5fd0493c1fb6ef731134f4bb269c891452c470c1a4e573de536874050fb41f83da74a2a4
z94dc7879dac60e5f48aa57398ee3acbfb6155e3be573c5f2889ed1d2e072a4818da61e93625614
zbebef442d166e734c2fc9569d45efb37d9d0d88cc7e16608a6eebbfd501499b9f765bf4d405155
z9027aecff188d741b565a4397e0125ec063326e9003f84ac4603c8c59525a2b86de00094bb9f32
z117c1d661a8d87cf6932963d6f684ea407833bbf545c996bc928d4ea39876288e77dd5b0114ce6
z569834bd0d2bb12bf93c6054c5ddd3b58e977b2f0d87768dc6640ae645ed2eb304ee82cd20ad81
z36a6253caaf48e0fa09606c487adb352fe3bb818db1fc834e44fe881d7ec158da1b95b77aa72a2
z934b7d4f9f73a8972c690721f4b01e5f6edc6942b1b6ed7dd09d36c21e7380ea65db5a91d78f22
z08c487931f57042e0c5bea9de360036bc65c1c25b6e69fd99165ef4e6c769e78c938fa64557acf
zf728415b8fb4ea51f93d4e887f4fc139f980435e22bf9f0fff6df9a58667cf84dd6e6332134382
z9c2fdd4a6baf2b87aca982bcbcb96a768a7424844604910516d2fc1313182059d18836f4e150c5
za6ca615903d027e1cbdb9161085b722fa3bdcf0f3aaec70b54c9cbd94daa4c90041e3423698ec2
z63fc800467306073fec0bc572bc42fbf446dd9c6c60c7870f1548f3613fe7dec2881808afff081
z16a0deebd53d084e61b449943250837a0e1ee591df8c351982bbce98393e98885e1fd8a2862edb
z1267e55be3f09c14afe643fa07cc23711e7f6e88c29380314f0af934687f76e202ecd9f4ab69ad
ze63d79b2c6bb607576484eff75d2968b730bbf0e3c8ad8c7b012f0c98147fdd0b29ba9af37c6df
zce485139c89cf5c2784647441d909bf50dddd7429bb5fe6fb35df3607118cb307a938666b7d071
z05f2ceaa2deb15264d0c7aebe7db54b8038a36a52d0dd36ec883ec27c5ee547c7b0adff80cee1d
zdd7aed46522a9c5e6f2d6ee8edf31729f9aea0b4f79b1d916b7f41b7c22eefe6b075d8120f273a
z48ab04066cd403cead20c904f711d44b60cc3203fc5aeee089b15f6629a960be0a212c54646be6
z34ce1c427ed1ad66b6ad4bc9434c787b258c77d61fc8cd4d25583f6dff97eab2f60c8dcd8fcbd4
zbefeea1351fef3d8e09be208c4ec7caaee8bd3078afe075d2bc428d0df0bcb934fcbfad877c8dc
ze8469cd8e3cd47b446166f17cf7864d81abc36ba0acabb4c38f32461e9bdffd1ced375190fc87f
z351cc10840525f8fc1a1dd5c97c4ee38038a9837f874e5b096a5f28bca1f9ccce443d9f675849e
ze5bbe1314768f05b5a615a49f21b82ae2914e2064da3c0268189c849aa80fc7044e0d25b260dfb
z2535e41b8e33fd5007f6252c3217e8b58dccec298c6758dd24c66ca1ca508359adfffede593ce4
z97ed74270fbdaac45f78f30dc319a66dd5d3646a6578370ccb961f66377154cc116015ca652eb4
z5625e8e46eb7a86ce1e70b751fbbe71f02a689733fccf0fffdcc8d63737c4af022a43528b22b34
z7250607d550d1cdf061cec49781d7fb91aea54e8b9532c388e5df651d97f1ef587f0047d82dc39
z0aaae31aa8830187c7a79d6d9e21178dbce69e7a964fbe102efaaf5211ddf597910f89ac966bd1
za1be47c4889e86f3b015b44d549816a87683180e2c91409dc468ba4b54fa92ba7e0d4fe94aa1bd
z6a840c86fe8a7da75982a0d7f9f18ca165ee96ba6837d75d24ce9d3c20c3184321777682ad088d
ze8234851f15825a3e9aa8274e9d71972c863c3d055c1f559ccb8ecf1eba4d79c9f8ca1cc0c45bd
z61fe4a9b434cd48d7a976f1d9a75d1df4ae44246e77437fbc19d63bfe1e86de70cdf1cca6ed4c8
zb55a353e8959c4fa8cd7ed1c0076ae4f7e8ecedec576907b7ce57efc690dbc11a5dcf888f8751c
z3874c9d44e51e88b5f51f22fec3867ad71e8b4ad30f96a81f39a6a2c2683a9dbcf1dd53b1f627f
z67a500c6e5723dc6e39c931b923676bb5cb9ab398a1bb60c236bd99430378c6800df6b8bf3fd9a
zc932016f15431b089a76ebf7110d00af6bd80411a5c927563389f8c4ff41e0b1b9650e9d3e1515
z45db0bea1b4ece84c0e88a858262f8ae2075f1ebf65bc5f2a01594d91c53f6d21a6bc00c3c4139
z8d292a8760c37106a0cf0ad593e059a1d71dcc8482687464da2919d860903dc7a4a51d8c3d4454
z226f12307292aff98129dbafb6cc488b74eb773f063ed507bbb1894e6adee6cd48ebc133df7fa4
z0e3db2360fed502dda332d485187414450b1073ef315883679ecf58a99689cbb28faa4a08e9770
z26b18870d9e2f28926989ea91df1a9d46bf8e59a3ef0f637e3073d44b1e6fc4030ebf19c64c912
zdae5eb4b5d9fd393f4a67cf69fd21851312227f8bba6c19568ffb8f2ffb48d9a3c4aed633b2b9b
zb7280e5b7fc25874dee6ae62f7cba9a4f784ef3e2dfb8eddd127cc269166f137737cc4fde807e3
zc8a8ca484ab72e15e076e597a1df374861aab9f6e7d05d23087b0c821535c0680eaa5b5310d625
zea7af2a1ddfce50ad4b8501ce7de2385b0c455c247dc67357324a22a863eb9d9fe943466952900
z8647666901b9774e9947a24f615027e7dfdc23b3696486d2245ff0d78aa8c87b6ea5e853e99878
zb28a1f03485321babc752bd5c3dfe52e2c2da6fd6de97f169f7819f16fa25821d2c53eaca1c732
z0d49ce2eb5f43087b1907769e4dd37275f20817ed349e3f0e1025a82bad6f9257806d8c8e636ef
z3222fcdf6fadb7fd2c641443fc12db0e9c8231e0bad8fdbb5d76d3d3965c28e40635940db4031f
z04d04aa09758492afb846353bb5db00315cd39c742f623a16898b839b7c42f8f88ef2f0295fa36
z98045c09529d577e5e26c15d8ec9f3d520401644563f5f48c5b141b5b7bcab87a1713d081941e4
z0823cda13ab836fe386fbf0c179fc2ad632e7fcdc287534caff9b93c2aebea51b2dd7f0e3516a4
z67f458f9de351e3544fb4d15d725edaff500342268c76fbfffbcf4e8cea87bbe8c6ce11ab8c380
z42cac18737d843eda09d7e491a78c6b9c90850f380cc21ede8253f172a990c2d463f83070f3980
z4fd0ef4652c0f5b7c8bc076a11f1da3603de53bc11f13255fb6ecfe35581921cec7c90dfad579c
z50fb9600d24f7ca797b6c51f0a360e7c65f64b4cfbe88fb69192b223c1a50d47a01a0768926068
z45b4860e44cf3c859c491cdcd86c243f17152852734f9116b9bf5e381bbd00249744a116785989
z71b2d8ec5d2147b011d3f633454c8dac2efeeba5247524768559c776b5c129be5e7bbf379582fa
z6603480bed52d554eb2a4320c9f8eb0c9069db14dcb2c89b6c5b215a6efc24e702bb153e973248
z1289ed04d3eab95c4ebcf21f85fc26ba21200e04abc1a5b7552cb2fc4741339c2da66cca04ab24
z967195f1de1d81030d09a2405a0cfd7b420f00f26b0acbe8d74664c8e59568e13c4b241069f18c
z5015e1806ddea4156aa1005c015b928ce93b743c4bd73461aab267634b04174f40bce268b89760
zb13c3b5b47158ad231dfd5cd80551fec05d5cd0e03b6f18ed15830d9c9c33035bc3d25539deab8
z91991f408d1d53766400b70b974d28bc12c3c6b8067dea984fd09cceb7f026a857c8152b5a3756
z9d4663875a4ce80e4d7a22381e83ad2446ea0945141ea70ead68ff257dab8b6dadd52208a4d7c2
z5733ba61c178efc8e667149f01baf613f13b769265ac26df5dd58dce32e6aa61b3fae0d06813fc
z219c0cdb459b500f7cbe10c6c25da3438cec68f66740a4e5f7ebacedf24bb177400b02851b5853
z0691d75c1c126360ba6d78b9ffc8c8104717d077f5ec376cb651c64c7188a7b6b96a8861d9a79e
z70b08912b0fac48056c0a727ba42d5b035cbaf8d26f04bf1da0b9939e0e8907041ef1a93b350b5
zb3fe546c54f93e9249ddb3fe12ab94aa4bd6f2bed1614d941322c81dd1b1e2958a8a93a7f500fa
z96851160fd0e26bd8c12d62d200543422374af2b10a4a906f9e9274c4c7c4fb0660a8abbc835f8
z4019908a87d3980da07b4d706489e9f645ab8cfe33eba582b51d8b1d42b7b25638b007c08385c4
zfdbe5698ca860710b43ef6935627098cc9391f4cc1e270f814e92a913b62d07a99d306f33adcc9
zd4762b65e372939f0d6aaa6bf2593d34e235b627bea53c7b7b1b1ff579a1b7fd85ca973814f0a1
zaefa91338ed3d190bed17719cee6c833dc1868e815550a5a6647e92ec2b0c646162da52f081368
zf4d84d2540fc16112fc8e49b133cb89c55182fe8795b4b3b1c75dba692f8c2042e42c6db7f4704
z9fa27fabca3565cbebd3e6247348cc79ed10d673ade445dfafea88e75866d7c8bdc57cd745980b
z27e42f5856f08bbd602130ff00c49662257fc94b3694a2f130de9a5c423c44f8d87ca80f0ef257
z2ee450314ef47fb166187dd2b68c6227e03d3ae4228ef62adec879a24a3e256a639e01c7f42dc5
zd9c0c8e210cda542d4b3e3d61a93415048d308367c1f22d8781e7edc187b2b0bf9a1effd384752
ze494dd46f7ca1e6ea1d7e59e275bfb119fc33f8a1c60023e305c27911a0ef53e881e8b7e4306e3
zd9a582f070902d0824fe1c3ba9b06e18a175d28c87337c5125d0e6808cbbbbf98b85ec5566871b
zb69602f971f0b3cd9ad36598d35afd51a18817df845bf4607c9c9bdbd12573766bf425555ebdbf
zb64ed93f68a325ede9be22a1cc5a5fdc49fcb950aff85e48de140101b7174928ba6a06729a1c0e
zb8c5b3581c96e7b4bca2ff03304fa370ce4218b54bd495877396bb1efb52fdfb86573f482f47b2
zc8886da68492c425af8b25be6309558b88a7f32b8cfa5c05e9f7d0c7e37fa83488c2d3e64afbb9
zf4964a27eeff67e0e301f5daa066370644cac17e9a4ce8ece77ca6c92d1fc24055337d8fb32426
zdd7876c4854e779c4e09d0e386838ae15b202f16f43af4fc214fa10cd621533a49de8f9ef54d74
z462b429a92ce7ad3763fcdc37ede3fde822d67b2de331d50f9aef84c07e384354d64b6db9f43fe
zdb7f154be24d83060fd367bcf7914b09fda0d393990c764527e77b80f9ec100e95d3bc00ab5754
z9bd60d1f08315eb52a4e080866ce5bb4dc6d7a19ca565a5fb6a7f7fa227cae87f4976b873752ae
zb8c6bea2829ba287b569dd58a0709745befcbe697fab7e7304cd5744721ec831ee029a6b63b789
z9686969434202a4f64fe43f5c96d477be876ada05b771e7717f8206212bddbc74fb5a49d750d17
z9b452aef394a9dbcea500adcbbdebfc10f4a5ffccd7e362726ed8a982ea7c7cd76dde799b40c36
z69fab6944dd0e14ba8120ce3ea9337e700ac5a6be8483bed073fd0f0dae855bd8ef04f12b8fd78
zd2263d208bf01bda6e5bbdecee9111f8ff29e2ac745e8083025a6eb11795aab2d4d1d5bdfb20be
za0d2afb57fe7931e79457c042230aa8f682bd4c0aef0de8c5e42da422f90ce1218157f053e0916
z1817e50ccb6ebe2dbf91bf9d0c7aa6eb732a51e137a89f57ef96fdb726d55c649fd85729213e3d
zeba1eb618866a38dda3a445d077bdb42fbc55b1eb2ce5cbe5b4d634b1a6e6895aa64cb6110b487
z609f6b0f583e5a5d5fee0f2e989342b2b7553bdbe1f2b02fc31c6d764a590fe48af61a8bb66a62
z8f21196b9b97da8a129b81cdc5a794213ada2c46093f39b19fae28f51e7b538bb102a968e9ce75
z2eb6e9cb7fdcdccbffe2d7a14c9a77c60b622ee219e77443b5046c257d379b075f19e9c16750cd
z447cf05e61de6c60f58aa427025657c466049607c34fdc0eaade72a9468c0b4ee0778a8ffa1cb8
za5e52562f8b755e3b039cca1e7c3f07408a4c1dc5a4361e8a087b1506d87ebdc0b9dff5875efb5
z7e7487de170afad1768be2d388e17f4d1d247c172328cf15798b22afc7b50f2cd102fc153d14fb
z543aaa59fe8a6a2ec342408c310901c6acfdab62cdc8bbb8f81b052fa8e6c2aeacadc1f3aa7f54
z408830962fbf87bd5774c6926301f85f82d6aca09e6d5d6a0be3fc92406ccd30c5762a035bcac6
z823fc2e761795af5ee8f390c446a4a1f7d13c35e013038f3d689548e9dd3481287f2a947dda304
z996c58e81743f29938dc13862f5f34f9adb16666aa918ade469460d162d05d3ce0301f059f064e
zcba71730cd4298d73ae5d98cbcb1b24aef5c15cafcff8d1ce87aeaba50350a235c900e4932609d
z4fc484a3ea0f4c32e0daa2bf850bd0750211dd1bb15093e63ac7dca36197a7bd6b175f9c4f8cda
zff6a51b61503fd382957ffb96b8d6e3ef6db402e8aa1871bddd1deff2052d921c4f4f22c1729a5
z38c2c2448ea355469de6e5808e07c39fbe8451ebf8fa3045b1f9edb555038969e416a360838735
z828c6225443e22a634bf6f784da768935c4c01ee461151760d483b08ddbe2b601d3d9541d8fd36
z2ee156290dfb2f0079d088d5ad8a312102e99ae002403bd5285787e12c091ba935d71960782100
ze946635faf2f29806dc5af778d5b21e4632dd1d3b798c9ae845e38691b72f40ada9d2bd420736f
z444e30a8d3f7f25d594e3b3e43793e7ae7ef55b11a8af313ce4ebeb00a21f60cae086ec05bc8a4
z97c5e08875073fbb047f7572f13e27835c6db8ba48bbde3c144734fbe07305f93f6f3fee7bc8c7
z4e66201ad970bfe4919af790174a44b5a8ad7ea440d12a231908f535e51d0551fa122de89d667e
z8fd51aa17c5feb4df744cb07584444c1ea11db398bcde69803344d714688841ac03e82eb084c3a
zd995daced62ad63bbf34ed8ead4ed350af52a255b1ea5b22c3b88998f98a1f38e4d6740d875045
zcc7752276a52b1740a228f71000f0ec34771cd3fad3a7cb80a48d450e984d9f5297711e84f8e2f
zb2c163caf30704bf923e09801b0cf9040a3e6e05ebc1aa2add63a9b7491a26de29e252f7e9dbf0
zc7682f0ea0ab1c84344c826c190e691eeed4c6d1d1883150d93e798760f365d826ae707cf84f44
z7267118bd15cce49cfce03785505b8b7a887b947c310ab7132b64b8a1c1cc16c3f2546c8e2e7af
z3fa643e91a37767a570a64229fcb99f3aa4a97fd5f94609033d0274f1a27a2dcc95d69745d11fd
zdf0c912a6f11636b56440a5e147f446ab81f244fa69cbf004c4186c900b64d8977210db24d11e7
z086c6e8584c1271d6f6c5b2d815dae2684371e465f01464d85efeb5e9dbcb98df6506423f95979
zb49d3947d2d819f958de24cf3bba82e5cdc5614320818713535fa2d374d1a28f4c8659dfef192d
ze35e8e3403664d7f4ef3ad09f3e5dbe6bc0a9de936fbda7fbdef868e179b04414014994dc21feb
z6bdf07e9e7952351237bb3752e355252085a50b53bc3c95a61e19016e113ae7a6f7c1c4f1bd208
z0ce6a67450e933c0459635a77782862546428b513fb8144f6ffeb9797cd8c876e2bf2310cd3062
zddda475825e17fa5fedfefe9dca96a1a6b719b483a8319d49205d4ef27d8904eef8694cc34b254
z625385ae712a74c15e02d2ab82f24b6cce0aa52a28f26512612583db4436241e90554b0ef948c3
z4a72f0ffc8247e9f097df5a9cfa028084dc9bcab16da653702de64d6c8ce381cb15130de7d3252
zd9507c6815e56a70c09c65b5cbc678c30c5b51656470707e1e2dfad4319f81c2fa25728f92efab
zeb7888a4cd07c15dacb05575eecdf27307755a221d30f271a7c11f6f2b457d4bcdf5c8208a7c85
zb3af4f74ff1de462dff3e018528f1e7cba1ad8b58c05d22d090ae561da64e9adb2e4ae1ece8c8b
zb3ae9733a1f812aa62df987253bf657ebb8c08b361315ca229d2d2c6e1f79db637b04d0342e709
z62a39d561b0e357ddb38fce52a6f18d365db065a2399f522935914a35fbe644135cf314f12e92f
z35a4e97c536f53144c5b3d11e33635023faeb67434819da08979362ad9f301674d6176343fe347
z198f1f3e521006e802766d157b9bdb2e9644f6ceabc7a362c4bc6591fee6f57012dcc64f9709e9
z0dc63047476835d75c2d30d63072e0ac76151d5c599e6dbb7207653270aed521328b05b36c02b2
z09b20f7cb3432da0fd0fb31e6815d1524336d592a47a93a17c4f76fc6b96acfa1308e0a9ee9d21
z33a3c4f13e22ed01fb27e0906c6920eedd7efac215dabe8279b0e4c6ecb5037647965c46052cba
z4a6a33442ffcf5d1f5e4c8c3c07fc4ca4706b86a98d1951aa9f54cf8160377234181fd2046128c
z66590ccf47adb9424dd592938646f064c614a2c06a63f31b4982fe8a5a6b4ead8901aa9fb2d95e
ze0be47c41cb174963696d9f91f56f90443df730ff67efdd62403087b2dbd836fe5e22bbe606ddc
z371a81887e7929134b27cff381f8b7db8577ddaa5509907347c238fc850a2e9d8f23a7933838f2
zf9fb48b4d6d7504c3a696b9a93f54a04f149fcfd39a35099076f6ec827080a4574b5d1d733d53a
z5172fee6c837ef87c4986aee6117e72a11d262517b32403dff48f6b0a4d9023e3d53e9c4c023db
zf007d13ff08550f5f592bbae460b335d46c73df7044f484ab0ca4187e8747b9f307d61679c6112
z3c68e613823dedff799de11f223ba28909f25113790d12052c44d16eda08d987bdee2f34d68bcc
z38aeff3eb67d5267da5207324b95677b55e9f42a2aaab79442d3f0e54908576a189aa0429868ad
z918a9c37a6cbf7211e1f17795f27f33bf32fddd07b144f3300c3495d9a5739c586af9235199895
z94ec8030875c3ff0c7f97739ab048cf58b9083563690b0540e516417a97cec9adeafe4dfd0ec5c
z0ceb1680cfc1baefd7e3dbfbf6a8885ebed5a1d4fdd16c8b7b540bc7507f0886d169438c27348e
z5bd1ef177f53f4a464846194ccecc025b1abfa9af02f4f6cff5e2d78fa4beed5558504ffd6a770
zfc8583ccd9a1fd66c19df53e805f5bb2eddae3644d990449670fc5029e0f9d4169e7256aff82dd
zc2a4c54ed658679fd2f73a843ef76301ace1fd9516f4cf5b1a3ce7fb1a666864c8f36e87c6801f
z1373bcf53e6b73e69b6a4149a1bbc0ddae6b41f560df1ea6b2ee62b9702e81d8e58ce041fe1262
z1c7df1e3245c0435717740cfa3d9bdbf16f47d0bfa640c0c23d9bc4db15e718ca253f8c8b5dbe4
zbf00e980913bcd104c90218a8d1609aef7722a8cf29aa0dd6dc80abdfd2743cc955ee84316d541
z8f88699c5d08700942193c49be25adefff20d9042dc1762680eee55cb615187075100cc9516b76
ze109d3a091913b798841cddb5c8e8597a8e0325a93e493f967f8436a52ec0b2970b1dcd9b3be27
z771a94bd93e1b82452e3e7a841edf0588d6728295f0cc46281d01dc63cd62777c06f4eda77bf94
zcb0ff029576dd59e15c3e09703870f5e6e772db271f28f3dc0b403bc7d2351fd08569d3dcccc87
za38486da949e6f4a46102af4e703a01c63a6577644185faff31cacdb72a2e9e821c3a8992735be
zd830922042c386589cf49069d11309df50bd75670af85a6ae6b84b1d87824251fe02c8a18ee8e9
z6145dc29849b410ed93faccae3f28aa17dbc9d117c3a1a0ebc25c99f968ae6041cd2881f07235e
z754f57c99d31bbf2cd499109b3bd294f49284cb98d50465664c4832f2a62d4a085896b9e71d0c8
z7db2062f59290323ddaa2ffdfd5bf5a070e549d7cce88eb2276f4d3e4fb76a8c91ee8c24aea48d
z286e83ead9e08101fd6690f5a9b0673cf6dc7a8020ca7f1c23de9b0e0acf7484ed9d04951c4bbd
zd352a28f35bbd90ee9cfc018b349ea18befaf14196f130715c981ad71e55977a6a41a5c413852c
z3ac937ec346cd0de7fdf352a4a0f9bc79ca9b80017283d1c8f02851d463341a1f5248692c252ce
zdf35d408a2031861a9b6962278c288ce8653c4b61ed387af3ca3f7a216e9f29a477949ca7af7a2
z75eef3ef5c5f364f7d35f77e2b9cccf7142d5d4c8402b838ad3966d0900d1abc5efe4663cb38cf
zfed457fc8c0302e3bf0e24b8d79eb165d704cf6af4427ec177d159755afb2f8559a506f1e71901
z5678703b6dda79bc7035ab5fa53f35bcc88abf0e9f293e46b12e2ab24c44db3778af1f3590a9e5
zbcbcbb6623ef3d93573b10587f167b57c6210d18a2cfcaa1d5fbb93070591d7f117c6aaff8c1f2
z8a8628c8f5fe2a9d7c7c50a29bd3c0cad71e2c61285d7c88d8dca622e2388293a47d08631ec34d
z8cb76e157e03bd3743ed6cb70382a2c1920884d492aef27f9a8c73c023357770879a809cd4e0a7
z750219498a881da9fda3d36bfa2bccbfdd9be7ff707a235abfd98ff260fc057443151ce0fd86f9
z0ac2174a2138cb0f5c7e83d00a7fff7fa559b358139896cf2d7c5140565514771491a4d7a1a98f
ze249a81ef4fd2f10be00a7277e392d48c7003c5ff408acd144e779d085b81e06d18136ead315a0
ze91b1af4d46fabbc0404ccc47822b52190676eb4c3236a2995af1a5fab8db12c14d5976d05ea89
zc6c2c58483c34a062696da7a42b655bd2d543a9dff9e468a2e0ac967c101d80ce98aff8d425f84
ze1780bdcf3af9b1bb2029c1434bdeb362811bc0dc37581dd5bff600248458c91f1f352da140522
z15e50915899a85d464b49746777252012f7c49bf2e2c6e1085f8af63e5971e036e214666546346
zdaad6aceb87cf481e140535153b2086f3db8aebde782fb1e109cd74b90df3b679beeb73aca272a
z6e8894840aba66f3ced0695140adee4b9766948a306f148c131082a1c1baf259b1aead2e0271d9
z0cb8d9ad9e63dd2a3be71b3586a651850a13732c7092b36634d044a09ce05da53fd3fa72b0b244
zb078287517470b6c96685614f4d23afe9e4132e3f67b33a36dada20d5b56533dce87b3ebaba042
zdbe48a50455e3ec66f047b1b4cbe949269c0542bc1fa2b49d364b19fed6983bc15a29549ace3ba
z32ef0c9d2fee4edaf996c0bd71e8a1e81139138e90a9f0865ed373385b133f4cfae0ae56620d1d
z3040140389a64b1a44ae04528e512e5a3531ccdfc31cf25f7b8effd3dd8edd117913f9bf884197
z3aea3ad9d6d7fd3478c91731722e104cbcc88755634ba47c6b32c850ea2e037b31e754d5be174e
z70222e687d21c09333ffa11d55b08015507770ddd759b0e2f9357d778e3ef4a28f9d424e5227a2
zfebb8a034ea68f31530814db21399d9ce7abed874c5c38a5354af310e789cb33185975a312e6bf
z1da3cbbd9f5b44d405fed2037d2215eb39f43a253ddc35b8d4cb5c884a9099d99f96647f5e070b
z4206077bd27c880bba36e02507e1b549298ed00715791db2420fdac396f91f1b8819ca7fd0550b
z6d280d5275e8884c91ed973cc6629553099813ea83bc38f48811a5c0d461d75e54c6c081bcdd28
z095fa65ad351506fd7b3bad799363b918c20d1b1ade6e6774de613aaf5382c7cafbdc80da9d62a
z4db67c3e07e0670bb6abba6f7f3b7469af19377a55ce8a7b140b79b6a634fc4f21f4ef4dcb5e03
z9630c0e2f807670ae2f5687e4f322906277948d6d4aa4a90c0c6b373aed7df4fccfdb431828c60
zde3ad6fcc58ebec149069bfe810a166e585d5d627cf6bfee166d10acadc40ada3e853d19744385
za88a341cc946ea4508a948d3c765df3a54b3fe58f2c706041a96b04987853d3b0dc80cc12dec2e
z1c22e89905579041fa3108bc6ba8f184249fb2bb4dc5a8e2bde6dc547faa6d80868b29ae2a07fd
za9c0644e941dbfdb4e01df91b8371ec8817172739de3955377daa372269d9e5c63230a05efa163
zac809421ea53b3814603fee1862ce28f3c2eb631f664db6626ae1397f8d326ab0b87d899df9c76
zfa548deee2333e6de48ab2665f783773a60f9b9a66cda022ff58af71b01b268607b25c7f75a7ac
z8082a87a9d5bd38deea5cf168656307abb53b513e08debbd3b12277aa2b79f662eb3f17874ba65
z3a603eb5501b512e3325683b9d9ebcc8b3732ce9786ce1cfbce91d09a0cc31c7e066677417b010
z7d9de5250435515096a74ed702cbac8bd85fbbb78e349b63d0510a466da65f827fad90cd66f86e
zc176657e44cc26df783030da137a77669a43ab702acc343b2faa513a35a2253af4483d20f5f985
z269105ed6857f3e1d9a82f866294dbefe9a1ef004a617e9bf4c686d62c6e7dafa548879d785c09
z717ae8b59a6752396078175aa911e5d283dd31a853960f667db52eb3531198efd9de985a5eb567
z4152f9042d7a18e22c945a1df46fec5d484e5a7a90acba3d10b8a73db1eb744b56a5df74371779
za5bd6881c76339d4cc6e8af1f5a32ef2b5c018c952697e547af7b2f46c42abd7e2e63c82d5d838
z987a41de6877fba29650554d910b193388722f5aa27a83f691dc8ba5529447e03620d66fb70be8
z154b88d50c10f28426c23c0ea3519205e1a87099cb2050c1066d88c2dc0398a928fa90b81b629e
zd65144fa45b46b8caa971d8178a8f587f2bef3e09fcf7b34e21bdc37289b42c9e9cf450aabb26b
z6acd4e760b137e41e901171145f73959b2152ae79211462d72de1a54803b170f792c238ba2af6c
za108b9ecff7100c80ce8faf5d1520a97de71bc2c51eae11ed1b0fa3a946acea7e47073733241c2
za21cbce6c1c2e3099b13b61030c7ac3a1ed19f7cc69a65cde99544510c9f8be000d93d629bbe8d
za72f59b149dadcbcb40130950e890f5fe2238cb658a1085a3cffdecf8f595f6ad7f43ff2b085dc
z31ad4e4ae34f40b4463afc8602ee39e309922bd2f74c8cbce0bd218f01a18ac8bd7d6fcb3bce96
zc0450553837b6e23a58933cd46ff78da1bcd4af044a8ae433232c62bb53780397b6d935a1dbdd2
zd6c9bb41109f2f32262159db349dbdc40e97c3e35a8e676b53c35141f0abad9ce31ea7b648167d
zb9b2866f7536dee2c9ecb897ecebee9a5745a7236c632aa64639288c19ac789937fbd9c84cfee3
z7e97b15d0879e07b3d5cf5697d0352b3c09fe7fe43d718a8367a4373eb4809d3fe6b6f65fdaa4c
z67c45d3f00afe3f56f4741f0f2871cc47275c72b3b9f2c1b0c7e95f0834fc0cd639e9ec43f3c24
zc1304fa3df94f6c0265888290c1a36eef92afea70817c7704fbb4b47b194edd85b2df03a34b143
z4086dca786e1fb406357fdc5066a6c0597e046702421a465f71b144b941ecf13cc5a03372f20d4
z55ec719e3c645f68a4e642476bcfd6d8dbabaae782ff1ad12bd129f444f4360cbe15766c08b31a
z7da448cd53710fc7bbf50048c288f6fd7a2dd0faa4390f42ce9cfe09fa86a1fb998307c8c00750
z3992f6db390d7dbfe8f25b48ae6fdad71fe87144a31833876f01f2928ceaae577f315d5fa9e757
zb320431ccf1a402e07cfef25002f470cf30fb4287f8dd9e411e85879c418ff8eaf77abf721012a
ze362bcfcf77d90fe293a33a7579a9fb3da1e4d43a22e1b8246dd2118f09c61fe0765605fe86b00
z9ea118475f5780fdc74ef11ebc02ff71ac7c9af65a038c99bd8a270e3639cca59468b870f8bb6c
z12779d9f21a1ba291e923b4f044c209168634e04df90bde4729536224c2467063f985999c78ba9
z1f1b541bff3e0a4d0f774611ebc18ee62ae4e50f8b23c7b12173c8be7765cd8ef1e3824699f0c5
z535647bcf9c33b21100cdae52ce5c5a2e4dcaef97038590292de665ebc5f3752ef0a045de2e63d
zff50ee60861263ffcce11b168ea584ef50613aa427212c7df4a733c35b26d3e2243deced852150
zb6b323680dee415089a7c990d00e80618aa8e00fe9a61f42cd8cf28259f47ddf969f858249c7a0
zc40ed08e8beef8059df44ba5955af477d381d8f2ed860c613477fa35f4765fc63ffff065aca623
z9d0142b637e3c37aaf2b935d152c2bd7558809e081355e029c1d409a69454ace10392950f68f5d
zd17c1d0a4710343284d31995dde48f049e9c505aa6d0c59bcf0c5d6e2443c95098402bb9ae31dd
z2984c42e599094203434c35c6c28cafd93d3ecd634d8ea5f6187546711a5eab06de9cad2b02e79
zf6c50662329e6910779afa21c7702abd6526f286789d6da25c061d39f0cc8ae1044ddeaf28a3ac
zface9b7105d13c05dad01bcbd16528b1538686886d0a211282cefaf6542e2d26516978e83d8905
z80cc537610b0a96be35c7a9f107e69ad8025e043e25503fa2a921afbbaa05e8f32963ac5016f76
z9b343d89e0364975e6c1eda413195dac6b23dce3011aa0cb435544ba9bc6bdc3f316dc0dd0d4f0
z97ef854cfd5e36daa940bde41dc62b0a1ec5467fd92d218d1d75bd17056272beb54c0d2136ed7e
zc3712d459ed49be62659d75f97e2ba378e5ef67270c2e232d5389b9e15701b3a4926a74cd18621
zd0305d103d364862d612c05041dcb99a3a5041da535faff24333e083189644dcc71572c8739d4e
z8554a3cf644e26d76d09c6594d7960852fd57a86806171854eb9f871de88a19b8edd90d78160c2
z1f282e94d037cba4e0ec254bd84e05f944b0c1defb9284997da2a79b66b84fb753f2c4932f460d
z87fc4200abc743b143d47cd71ce08d5b55cee5dc7d8ee42cbb661c6207f9006a415c6c79169d22
z37030c08e39a82414864f8c7a6d0fc6009d67af16a42f0887ddb02a408f114dc005c6ba23e9f17
z51ae9741e0b0c3b08b79b317356594168c26c5c2996898e4bbb028eb8b0699a6b3d135a63850f4
z81d82329331351b113c03346c3509200fc9c40483ae02e4a514d512db0fb2534998a27f31ee03c
zec68d753a9ac55a2650e6b028c861ec8661a0d0c9c3c5a390c7446cf669e3d4dddbdcf3c39fb45
z6e51fecb07113a04729661382b115c6d3f7a2d5ca802ab2f9ccb95a72866e099b2fe0b01cfba4a
zaec8f49dd3e15abf884e3b8f5369ba275978c66d8e7ad92b7063e35e331473fbd87a18d53af79d
z5e810131dbfa53ace0b81c5a56e42c6604e2056fb83a3c1cdcd1ce2579b2c0e1eba3f14f44f7d8
z5b75b70b26c88d672d51146a9391086296d32ac88ae980964d8daef1ac1d547f6ea47b5f035af4
z26d2bb7c05a96658a1d5f37b1d582c7349acededec45119dea2df38fe7b448c7cbf67312806354
z3ebfd81ebbee34d31d87fec0385245dfd953c98cb0a3baa03af25287731ef455c74cf1581c3a76
z2edaef7138093778d76e1d105380c695c5ff1e499913ff2e94e20b36d4d816af719e356ffd999f
za4f0d7f2e3a9880812a9837594fd7648191f29d69562d75832595ac15110643e04d2a0a347566d
z7368e787d46e1551d6170a0286a7e8be0b5db0cd7657e639c324c84f9d50976e089173537cb3cb
zf6f6931fcc64402b6f4c72a55e6901bd8307baacc5316a857d127ac2ca691bf135e0ce8d5e75ef
z97236412800fb68eb53b8e1273fff6dab108fdc7608b42b94a910e9825a592e9da5222087b0819
zb21a30f137473831a8e3b3422b59e7b7d7e676e2b763f525d00baab9fff4caba38ba76ff51e575
z75d1acc2570fe9d6fec720dc8fc2c2698ef5d857eff937e1faf989c6de8ba919cb12b606b01136
zbcf3f6f848af66197036af44f9941e237fc8e3dfc71059f6b2eb1826748ca1f2b20b5f9e0a3560
z0d946a122bf2998ebe5a65e2e16efefa6c2b658786c237bbf4db7510bae2e637c97358a3be5cd2
z91b672af54c0b45705d987755fb40c16e86a58ca766eeb866f0d246383100fc0620ebe3f4b60e5
za04641a6b616f834001d951db6738a2ec097abbc0de237d9be58f60073f4fdbf6c396afde8037e
zdf74ead2cdc1e60c92ff24b52dc03667ebb0bb6bc897798d0963f4edcf66ba130875327cc9c6fb
z5500822f324c464b06e9d03c4a10f0759dea91a92527dcb4f87b4e9086280207a5c16b92ee6f70
z3ed05c24e8ecabd3b9466a7f6afad3f7be0d9cefa20f0592aa74f053c40ca7fe91c4cd2a81e710
zf9f3459c0603760a09cf4e87e74a19610b2227a48e60b6ef60489e41cd0c0211a468c0d913deb0
ze1dc5526291717f233e8299437d63ff4616b7e58d58220f9d5c2f37f0d97ae22171b999cc7e7b6
z95055e938ce3143562701f11e1229178658a0ad0687ac92962b80fccb65d04cf931f250faed319
z2459beab97e1f8e6b5cbaf760750f179f6b78f51143eb800c5ca54d927ef5dab186c90995a808d
zf9116fb3bebf60530c230228e32f27a7012c15319e55850c1a97f2c3df2fb5b391ba693b5a1a6a
z7179d65cb8e1ccf3d03a9d19d4c23b5aba0d4ab71f9178b3a764275f030e2ca88cc86dc102be02
z91b46879e3e8ffdba1f642e644b08e10df3ce47b2b95ea016c0d564f60592dd549c6823b07b502
z6d9070a633b9bc686be505dbb3f8a2fe8896ed6cd90e775a1a973a96e127d07783cb497470a3ef
ze8c414688950cd76c9e842ef47d3edcd298d7d14252acfa68840fd05d7d73298c0486816e87c14
zf5959ebd1730b02fea800cd02edac13d180be801ab7d8bf0f4f9060b264d82a551ebb06afaea53
z53444467d1bcf508e95e43d3f088ed1d1e03e7143c483c2646904d239565b07bb700e2c76df48e
z370a2cc7b708eb400d0b5944466fbc20946542886dde4f584831fc377866e18a6e1390aaad0dbb
z2c4e28c8d2f6c531cfdc5c4346be4a08c00823564dc8a2c22dc1425ce64fd8bef23389e8d304da
z19ea2f764ccc1cd2dbdb06ab3e30c5eb5e6b2dab00d0ba64ff018e004885f9c218129a59d7c7b0
z3042ad35f0798e03d40d0fb8fe9d405f432e7867de7ed85dba9236d8b7689078f65069c74ac84f
zfd48325960cf3ef40de987e32ffc821fcac9231caae05bd9b07f1efb052157f6295b00ff91b69d
za91b4322690cd1e3d62d0fb3403bb76330da884e192e9c181cf828571de4a3d3ea6b42a3fe711b
zfb6b172d6399b7e7bac8a0719d29021bf55ed54a3a5fb0d9d67d0670531df4b1aa0814e93208a5
z97cf021c10ddfe5bc6864f10546ab0c7457aaf4e9011b8127e70b561609fdd97441170011728db
zb352c32185e7aa2e0dbd24b1fe3529ecaea422f9a7e31e2a7494e0f398d28d2d122e9d2630d3f4
z6508642ecca448b542e3f7a14b40036e84d7be0db899f0d91a06bc5ef569030093ce973d946dac
z2db4b3ed6167408fbad3aabab9a62a671b3cbd13bb47bd478256a058a6dbfd72dbf055b2cd4875
z919a0d4460e75556b9bf8a37b03aa41c6b5154c2d32c2d68f55d0a8333218893a475b0bdea107a
zc7b6cfa391431cdf943515364ee9bd7e75de3053b685a8ae15645675b9a7382c07c5de5bbf7e51
zde020323eede7d022c4a37f0ffaaa2ba078a94da3ad2a86fc5d1bdddbd5061bd82f572ddd248ac
z1c02e3d363cf8832ee97f277782c6dc8376f15a5bb1679babf15a05b66c314c8bd387d7ac90776
z550464c53b4418eba9761430533c3616ecf8209c3696c17bacb0a40c3017f5c8bf35edb344feed
z8027ead025c7f39abc2016826d67732e0bc08d0e6e2761fe043e50cceae5de024e5397d70f74bd
z2dcb277865944bb59cd08e0fe49f9f34d2a0eb495450fcab777e1c2d6ee8b20c0f8c250872e6f4
z12b7890a40157ee0cf86832f6acadd41ef0ff3452d06463c823cd95abf7ab69a9e4e8100df7f5b
z02c5194e8eb7e6a21209a04b2ff6f075d1f05236f3536c196c9e17d6ebfd5aef8953c6a40697ce
z93fbfd74f9d55dc71185c8d79cacb168d74795d50782a44a3da2d5f8a21e8687bb8bcd73c96314
z62e7510105ef763b517bf06cfabd0e7c680a61e9aa2af6eb10cb547a27a3b5ade8cff4e1fcbd45
z0b6cffdb2862b915a987cd1a7c8b5652b6cf42bcdd085ee950b032d64a78abd778de43aa6174eb
zc654040428d7442afcef51a42baffe9ef5b41b6d2e6de5c6fd7aed23d2a4ffcf24262d6324822c
zb66381bb6187a61053a02c2fc21ef96eabfa8ec914e2f6f657c0e97d8ae4a6e6176b39237e9425
z1736df686a3b517d73d80fbfa1527f5cfbb6d1749b5c92798d256548a9436a523773572fd42081
z2a0559d299e94a5cb99ddb080fd0e0917abef7e752e33ae8b556dbe8d4840e85bfaa2273628c0d
z6b039b6dc638a2468f3e2f5f5950064c9f10e2afc3d3ce082f44ec207144785c520253351715f3
ze728207cc97db1ef6835adaedcea4dfb1006523689834617f0b728e6c6b3ebe5d1a2ee8beb3326
zffd991ec9522660973d0ab736faf0db8db6db11d2d7a3f532115bb28cd91a5839c2bb94c929dc5
z33ba2d52ee21da99e26dc379c25bb1082897ff6a556de159f095d8597b0ffc76b08de3824da2ee
z0c062ee56058260b0662317d4b77abbe68196805e4602c5f5debd6cbaf8313c03e99468d05c897
ze38a3207c743d0cf465a67b0f687c0c063f711ccb5ec9ee52a1e21a7042f0657f524c6e4eb88ba
z70f5e164a1113c815e8266e3b1ffbd0d0bf94f1f2af7d4ac4149df1e51572f77ff47a9c1b22363
z342a52d3a81490f6fc86faf389a0e89331b542ea4d1d0dadb259c890c739a0aa912736f694b279
z252bc7b1d12401d970d17af197c9ef1f7ec45d4780481c524cde1a2ccb287b8b5b8ecf4cba7423
z333bdb5a5da9a795a93c76aff34571333161f207da9d584cc695886ad8562ade08dc5c4c3ddd47
z520ea041d843352690772df4f86bdc2a5ed59c4f2ac3e94d2ebb99f382d0ce789ce6afd300f97c
z3d0dc0172fb67481251271eebb5017a7ac510269da5acd68934d290b06a93cedbc114d37556b05
za7c358ac5eea398bbe3141a85bd505a8ef292b43ab5a8bf0aee3a4de7d47adb23bd0a020ef1924
z29a34bdb05e3f30ab21b6d6e8da1153590959b79f79ad8f666f739ec3f6ab8a5051438cd58ead7
z62f84a983fbc606b71342f21f05a697e480e2f4014dac57185fd2773286d87a05f7496567f25ff
zf2c0fca31b1a1e529948db4a0a348774267104695b787105e0f3c9fd2f7bdb7d5df77704042676
z43f0fcd8397e94e1fe722eaded6985ae84fe65e30e2b03696f2ffbf4991cbd3744819017de7963
z7867e381db45e1c384706e2778d5bfa85ae8910c1abced941ed7139618e6bb2dcff729c9ea228c
ze6477556e4fd41d7d89107a89832864c1b94ef6434972de800cba64a4b7c9c1222b8736b34791a
z87728f3005adf3d33cd7c8ecc13463bde49a50b2158c3397e01f7e0f5e72a719138c8db8767a8c
ze2fc689bc9f271da6bc0112049da799a237b22dddd25749846e7b1609adc5272bcf55c7dce0909
ze3219b82ef0cea06b9cd152ec4f6830f7be1fd918bc66e2312568075c6492de87871a10dc02e19
z64cd721f0bfa2b0e1fcbe81a94d27c03c1fea375134a7434f46b961d9baca94d5f17b885866729
zac940f34aaaf7f1dc48e8e0bc8a840a3858e31a559bd84d1e05e4ccee57fc8855e5b342d88c2ff
z22fad55d265c8e679d86440537ebe87f171fc075441b0834a318539da26b387b15af44c01a24b1
z692f19835afdacf9b5924479a96772b8ae08098089f00010caf60e0e05b40bb1dae568b55f9495
z28f2945586e2afb2f2bc9d4b7b72e102c14d85d06feb176585b1dd67433c0f9442bd18d936915a
z97820c1a4d8ffaa0a16471d31cf808f8568e0a5bd92529c9c2a3ca304cea2401fbae0236df9d03
z4177033eb231b48f239f61d8c0a44ea844c3dca9d6f1f455a4f8b8a4b1e6734d3f89828733d4e0
z44ff657ed478f3b09a284ab98668ba0845666f9abe0cc4de6e3b1c61d5573d908ee3441ec3d3ef
z32316fd92efc6e1fb7f1c3e22252a8e4b732b68c829e9483e66d700a9dd8dadd2453ee2170c948
z5f07fc4cb66ce1a1df282c0a5522fb68102e5b722e26e49f474904d6b558f8ec18bce2a94ae5e3
ze45d9ed30d104bfe793ab2041c53366ca47cfbd5e349c6bb164be6534ba8a630fac71f5ae22fc4
z96bfa1fee54233ce06e28ccee38995e61ebb632fa3998069907842aa2e24618e674d2b61f07cf4
zd4aced2c8d604e914ea7a8d3931133de6b7e4adaec81f59073b87f1c8d1f030141aa6083b40ec0
z630f475ef165c6bd336b0886c31bb2628aa8cbe48cef88484e854cda8240d04963706bf3ede96b
zdfedaf1fda11bfa72d74cc2da2dc37280210be3f42bbf721522fe6191fa2533716d89cbe89e451
z0cee2677009362e68402fe9de3e28988e1d2e3cd719ad42ccc6aeb4dcd78f358e26c8d2fa35628
zc51a12d5a5e5b1fd26e526d3f0ce63a288854d0e26aee68e918ef824fdee302f97fd0843728baf
z08b0fbaa77455f66cf5e3959b5ac350480c80052cd9a9c181ae1ceb14959f8fa23e67595a0bd7d
ze9b0400cfc7e21514091e3814f41187ebb5f3dcfba3283934a0df3af4d7f8ba0f92f2cde59f17b
z1d72972a0e425170916b3bf44a146245746bda007dcd8728e9174e6bc234ab47395bff5bbce409
z6456c3a694e05b968e2c9d85d3d4746e70c38abc7dd9f036c6320c5c9aeeb021699320a3113ff9
ze31884f08b138d52ff6edb0f096de80fbec46714c19f0810c100190862742f83d5cd4dd6adb904
zd0467624f90cdbd9022ddee9982c95aced444b525eea9f85c5731ead4bec90b4bb9aeb3b44f60f
z782b52df4d44af44c801db60e04f0d07701e71e785edde32b37c5d68b2221cc11de44ff490351f
z63adb94d988c4f19e7adf3d96047d849254d43adb5c58e442e0e11ad975097bb7065b0832e3760
z97c6c09ba0885ce90c6bd0d6b9669cefb3e718d39eeaa901463a3441d42079842ced087cd805e6
z36aedddef6052ec82ea7f23c62ab9db7637fdc08821ece821eafc30f63d6f27f87dc6527557e62
zb046bf0a3442c0f9aaa380c425c47064ab2e737cc447f67a544026b5d68d213fd20e7a40826cb6
zfbd8ba3b497c9c9fb1de7407f5bd63afbc4061070eeea9f0b9199233266510c679bad18d02d371
zae284bf3048056b5fc16b7df5caa5241c100db6bb3dfb2538bec4742814e8a504d6328302d994b
ze63e7f33fb60f1de772e1c93923364852c4f031fdaf8d9aa7ada4dbf0b2c9dc636e7e03c35b88f
z632df2805867092b005e1b5b40b202add42ad780231c1ba27851ec69daccda328d470d627bade2
z1a19c98c95d25a01421d8fb1cd43700bceee628717dec3fb612754dd1b0dbff133f0134d9ac601
zc64cf60c80299669b9eafe82dd3bd8a722f55c19101cfd4f6600d774a0c5fa84d4c6c683abc571
zb98799ff2d14eeba46babb09afa9444d95630a3148d079963df7a7874d4df2005cc117d38c6098
z0c4466ad541af0668f01a2525b3d955585bd48e11d01ac42a9ba86239f2915112d3aedf18d12b8
z89360417c441b66742b777ef7597f9776faaacf2c060fa6ee035469293126314667a9d77450ccc
z5becc118a5297da2cc7713a9f6a1a78a7e8e79726b17879c96d282e37252bff720930884674d84
zceee1c0a7755bdc97c0ddde63b15f013abef5143fd60c5ba878a3e3d0cf349446a4092c524b83b
z1e3f40510b7b0709d8519ca1b51c530c91944528fa6b0f07f13bb268b5c86365218bb365310b6a
zd4ea91f21fcb742b5274dbdca816e6e9d34c9c4192bc6c6435045391dc11f5907e4f57d9b0ddd6
z80a99527e279124d56e38b48cad498feee488b276021459f352aa0ef93d727ad2b7ffaaee67292
z8095074f14ef3759adcb40d963a51f86aa5a0b387a3c48479898e3cd7143b69ca142d4ec1d0cab
zc87861f59affda022275443c539ee0663202e8d7e78438bbf95216b51f9861efa740c97a966f14
z98faf1824377f3f8c98d176b3aa06a8a8411b6f9fa2cf62afb48ace0828f31e9f1d89359756eb7
z0f6907219e022c061bae9d6770e61c89c4b16b1bdd9afd798f38abeed22c3e50d4733b10c0acaf
zb653e6983a8af2c4897d28afd456a3db064c41fae8461c42739e763f58aec333c5bf30612faded
z2abb3907897c05c70f4e4de9b11300517883623b2acf3bfa0f6370e51283427c297ce92f04d39d
z6121f90a1c3f32863111ad3108a1ccd8c4e48a2f03338060a5fe9a5129acc12f633048bccd33c0
zf2228ef4fcc9e35702d799cf1e018953535971418f2e72a66fd9a1a7851edcb2bec6871f5bf134
z4c5c7a651962c90020f8fb0c3dd18d5e6ca8c66b053e21f9077080f4254240efe8a1db775b44b9
z0849e713a95439acb7e2c3782d982e9efa4378457e4d2efcecca80de860743e0876def1b5eb64a
zc1f7f3b6cb97cc6ade3926267b8107e68e4ffec8532294d44f1b5fb8b446d1e522af667860b861
zbdbf3a0480c346e211a99399081bfe9a0ca19f01e3183e2e3346636f2b3608f2089900e7df10fb
z7c7d358f2e195a4407754798e254e1f49d3b401d20d3c0f1039a0278849ac88690458682303f4e
z48e2a2c24c3cd51c85ca6b122ec44eeb67201b63f1de32c7ea903edf62a3de3db55f8d36972baf
zbc4c7cc5d2193bb8deea1bfccaaf3ca5131608d0d060eb7fdc690d65fd58c69ba6d86192dad1fc
zbf842f5654b250e04744e213b1ce1fa534e9f5762f478fee293cd3f09fa6a02aa316d329d2be63
zd4ecaa810bb60ee38485d68ffdd7cf70d1ade3230f2018bb8b62ff6cbe02e2ed0817ca62711615
zbba9d568d1167a3b4522979750d564561cab7b1e7dcb3636fcf4edeaf25b145a2bcfa3a0c1553d
z57f7551c66b49057d2ea2a726f6c9d5f361ec3d01479d95c27d83f754cb71b9bb3d03dc85893bc
za7442a3eba3aab772e72ae8ac01d89e58fc666fc5498892c3031ffde761ed83da6e7541f5ade4e
zff37116fed24fce06cc7ca7469c1df2cdf04f1a3e1c94ecab9170d6fbce26a4d5f9eb9debe5f85
zdb17f00fd6363fc9d133c0f8a6aea5281cc4b3b98185a3c7b303e735e792d676cb412f6781fdd3
zcfa694f0cdb76c59d3b8c34f983c8d823ef138383256a71881cb48b81781aacba1797080b41c1d
z7481a44b62580cc0999b842274a437377de07189745695c3b3e90afbb45c0f21d9e02b24028f19
z32be86e3a6b7006060e6f4f904403af4290bd715ad3137e2fb982819e81c4e058cc59fb85baaf5
z19f560711096004cb19e2147a3ba728ac0a385076342f8409896db042e4621c26e371e4f6d894a
zaec7eeca1be97e956b34c5919ae77d069b7362dcc760d5464f26c446778a45f79a27de311f3297
z221483d65cf62b1e85d1440957438adfef853ec44c8057730e88b061c0f14828914e11fe78914c
zb74bfe8f480536a5b580fbcb83445f2d0c68541f83069a5f486582887e6d7e988b487d97dcbea4
zba1170d5e1e46319ca83790ece8584367f7f93c82e383f76edd33c9f6945f5ba4015e9ed0e29c5
zcdc3b005ebe91ca420adc936d6b82ab40aa26b95446322a2b7aa8726c54b671b9b04fd642246f1
z2ac2089148f745a68360696455ae17d7de5399cf2773951945a778277f4a30632fa913cb6fc1fd
z96f89640083d2b688fe7464354d47eb3c3f1366735fd24da2523aff0c01c250d9fc97052873ce9
z09719bb1690072b7eaa5dca2cfa8d2ea17ef440af032b3afdf8f23df7200598acb5f5d9772dcde
z6039290aa1a7b536ffa794e1733f7a11801b3f45085cb821862be818616333bc1186297676a678
za3f719e496a7dd4b587e198d7ccda9f2d7dcad66af0bcb396caf3007f29632127cfdcb784a7c84
zc87276d8b3db2aefdbd6d460ee10ad1eb9eec2016995ef8c7814fc4e9971401250562b9ae3de98
z90ec6141226b4f8b4df5ad01e9ccf2346d90df844ce3e3918ae044bb3c1335c1e3b63f6cf09565
z6029b1cf505194fe5823af9d37dba0657764c3c704cd527d08efc20fb902fcf5f97c2c166a87f3
zf2a4360fe53d3c6bfeff83ffd4fb842d7ce126a5b340ba5fe62d8d7d828694c28c9693da30670d
zc015650d7a4fa7231f029790345ba92c575c8b9c215df8b0d99b97a9ee6267ecd78f2f219b56fa
zf091ada4b6da26ca50017122dc7f09b4a364007eb0b0594bd56be8e9dccad83da004003ca17e00
z38e488884067160563350922b3bbe3480cb307857310b99890deb027a0b2c19d75a8c67b9c992a
z8c9b60bca50ab01d46d17304228811ba4e540c5052a4b0f49ef2a01727880aa02edf0f1831bdbe
ze3b1d8031fd20ec3613a30fd8e4d6dcfa17556f97acb8c824dd6c99dcc86d6682be6b7fc157013
z9077b6de87b1d91c30ebe75253e488fee8a9de340dfca91fd91eb5f466d655145dd8f9d0e3712e
zdc396d5c42df2b5dbcc0352b89c6ca9e7d921b742b3d1a147f9e638b994ecfb6c2624b5858e099
z69d2f0d0fb74f550ea21dd6c1b68bb62d7be541c405e238b28686bccbce206999b78f91ba8ac7d
z2586a2e94cd7481889cc8feaab7c220621d0acc25f5dbedaf03b16c75a9ca46a3f93d52ce1f0dc
z742ad0a99ac49dada16c8fc8a8dec2e72fb0f4c7a912fe827e4682a20f8f89848d5433efaaf1f0
zc89d72004a3e60b31e0ed29197cfcb617de15431412b4f3238b18720530976cb95eaa46e58073b
zf5ad50a71e12d7e48e425f8953a5119cd2f95f68df5c9dae3bcc3b4332adf42acd4c033852026b
z3852a6cd3cc88ee862fa9dbf79d733574f91ffcccd121944868e853f0b6280e13a5021a918fb04
zce89cbf919a9fe469771aae3aaa35b8fe4e6e8ad02f5583b020913e8f14675ba18930e7ad41cef
z3c6cafc0175acb7a749ee053948a00b2e4be617aad5df2e89f86f470ce145493b661eba85b1936
z1254663f61b14b148bcd3fa1b01289d612e17a816cab1d5e134d2693e2eaf8aee0f5b4c17f456d
z99f88ad979ba215036811a6ec16a66956c62de05ecc97ef1e096401490ba2e2b3a73cbbeb60812
z4ae4dec72316bdf347353239f98e79f9d8cc7a041c643e80de879310ce14584a4d8994af8388c7
zcb8023a849cb1aeb86f49c0993fb4ecb3a0d5d775a147c9e725fbc309b5d279d3322b81432b527
zc5f51471d91a8801c2b1b4a1e99e5cdd14b140cc5a789816ee3c561427fc5c8a704b11fe409c6f
ze4313e4076b6ac991e8132ebc7de3c88d45ce7147bc936e45a2c67eb065d554d68498df8cb0e22
zff947e1b8a568e858650321d2f67c2f6d42496859250ddfc85d9102ad21db1d1fd422dfffc3e62
z01f008bea98bce77d749ceae4076ffe599fcd099276b7d5133ce36aaa7d669c6920cd916e893e5
z04c01184eccb3d68f67db787ea6560533d002a15049f55ddf16c43edea2a9236872f70cb4da997
ze47664e0594f09d4c1a136be7956531fd4e68eac9f17c71866f5aa5a2d73e5c76b848ec9d12e2b
z6de1f62c0aa4034efea1dcc66973b66da25c63541025b86d994e12a4f9b0b5cb2a34381820afe6
zde417d33aea39e6906aff037219ee55e4699d563cc97454f971f169c5365eb7ac95298863195eb
z366947029a5b2596e912e289562dae3a665132561c85c486ccefff122ed6f8549bb19866845f28
zb9fa7a44504ba579b99d35c60c2db0fe6d983b18caa84607084bd1c4988e30e06760d24268d81b
zae95d837bb32e845929e937faac174942a2d6c9fad3a93c7ac784cad7a82fe1c219c89e525663a
z0f4ab75ce02e43bd31c18368953f3cd9e80baa3de626623ce03b8beb6182e8a7c8e2285a0069e2
za70679fcb7d8be86342e983f352592376b8703867f13e80edcca8c5390f6d61d0fd7203c8c50a0
zf7d3e08877b7ab270767d6879a768a5f7740886c3f7460ef42ac085443ef388c9e01976f2b072e
z106f6457ca522ba615336dfeab11db0b643b8759cd3688828c685ea93d41674a57147302f84e0f
z99914e7cdfe4dc639dfccd3b6ed230df585685729950ee0e36acb86b5c4a2d626d433bf07ae4af
zefc711c0725af73a5ba41b485c5904ba2f0ad3a5e5b5092eb118b3f4ef5e88b675ac4236b4291c
z7637cb12b333f0c62cb2cc280c5d2631af4c818c103bdbdb26c94a7c111e3c4371a30aa9243bb7
z7877753e90feca8bdc3a91388d36bb96e7580f492443239b3cff4e692432fb248a68097f7de7c8
z0ccd0be530cfaaf5eaf2696d58e852db24285ef1d443dcc9d6ee4302ad0d680e3faea9d1591bb7
zf90290bc18f7e6ca0ad8bcb88fb31ba9b3a3b7c172bee121bec7aa8cdcb1cbacf8d1881882f6ab
zda02d46fb242288a397c8599db6b43e6baf553e94cb404198f0e58f89c37244e3478d7517ced3b
zcff96b0081f4ab652ce0ba01e0d8dad8cf3d00f7e0e1b7992be91cb43b7944ab804c8ac1ea2e0f
zce6704c7197944f399ab409a7441109553dde87ea179607f2986b10a66410da69f5fefa79359fa
zfd0b09fa3baf787af635e8d13790ddf6240a6f0bcf03d66787ec0bbeda52121b09d9a9c54395a1
zbea9b165d9f6cc4c87875d7f42ac21830da561b35d9aa6d1258559112fe3e775da7845c714a9fe
zb74d6d93d11f2dc0e79d92b5063c0975618c73fdded6ec90db8e6342d45acce5e03bc3dc8c4e2f
z357c2ea9ec355f300f127630ec76cb12d722b2e4a125cc92d3af56ca7d791640e966158a84a470
zfaf8feb79ca0ab4e7489c015a2a5afeaa2520d193242a0e4d55fe2439891781c994a7e3cf2ddd5
z8a14467477d140265dadf5f428fb38aa3774a2c7ee21c41d4c46eb6bc1a615c960f7cb8d8f1e14
z02c7822d1f23d2b937afd0926f5eb0b857705547569e36e1bacb519d8cb77e543b9537976ae742
z1b5e68397e1871545efbeeb4371aa5a94df14e2334bf1b8b7ee0e7c99a8766a1cf55840fa75fa1
z955ffbdc7cdbd40df62035199c6eee384f5a04d200611280e8f9fb7af5bdc9ace84a9aa9c0a191
z14501fd9ac243b6ab2ae25b93b1467dc1cdd69008fcffdffdc80cf61155a263b2af6db86b67fbc
z0ae965d59c44dbe12b9613f28d47503e9307eb0faa7677e1f9c2bfe2bd83aa7cc59bef7c3aa7f1
za0bbaf42cc66b5eb870b090d177c2a676d9960dcd657deb8105762642c6adf0b7a3ee79e8d011a
z30ab5232809d574f97742061b20967ac11660ddd3f3a0d34eed3db57c4ea3c51b9610b228e6479
z5d212e8cb580b08453bf90cbe92a9d580bda6ff7900b66fb24fbce98a4bd00a0da50b69bef0dba
z12aab97e6900b3893deeab1f926ab4a3544f2cfa376ea633797bd11078975cb7e97c218794b77d
zf71b239ffbd22bc71e20b9ba1751401e1b4acc00b9624909a8d3f1ef8c99b13b364a8f5746daee
z8f31fb7d739c3240cd12277c9cac339c6b6c084fbc7a493c161998fb3f0feee7cb0689f2d74fba
z9077760af43fb6b0a1441c8cc46894e93b0bc6e16a8fc266dd9dd3e64543796f25c752053a0e4e
z2d1d12075a23793f9b164bb092d1ed6db2d01b9c41c401b558fb47035fb636e22917381e26cc11
z0d9294e4c85797256c33ca7512b0302a298c5983cfaf03fae57be370797c49b26dcd051a069be9
zd3fe6f1bd2207643a28d35309d5ae4830dedebe1e3434db04d2e8d94b369b3324d27ec060f680e
zde7d5509a4f01af8a3cf6bae0bc202e71b46dbea74887986ed49cbd65723ded12021254e4ab6b5
zf2a410eec277deaacd08f1c5a86f44e066d98a4e828b709d95b2e58eb500173de1c13115726859
z82d371ac2ca63eef2b2e8774551aa2129a2c9e8484458ab5f7d66c302ffbebb3372165a7d06d25
zbe97c346bfa452c88292dfd24a8cc95873b5ea2fc5fac7242cc8ebdc526a6dcba16814433ca6e7
zc79a41cf739569a9d7c9aa60eedf3988a1aa84184577e80b73f456fbd7656d190b38f5967d8e0d
zf0c33227e5a9ec7429c5127ebd70bbb9d83ab4699b7b7388958a06c1a6867b4d3d948abad3cf7b
z75320ff11b27613ec9f3c9eaf1cb4d6e72440ccc778c31f48469bda3d98fd7c34e8e306ab998e2
zb8ff69d819c243fbff51afd0170f9ad1027f19a171215d42d1fe1956566e33dda85bcc1ba0164e
za549253fa54406a017efab7ba833f2ef4ac3e55029f087ac377c98133f5e03168e4abf34219ea9
z97355fd31348d78d5a3a9ed18419c1e7f86a3ac78c14771c5a6d6ed99735b87cfcbc9bb1670204
ze648719b57e26a8d5f0d19cb655f0b8086c76c70a980fe2c8483e26748a31c7869817fe65916c7
z7c4c59db429e79eb4579a9c6d8412398606e77bd1325dcca428daeb0358c5b0b23fa0a8fd0b3df
za37af1ca29b315e9eeaa408a3e3a8e75b72a358fd660ad1df929c5e7da94535b38109a276e0401
z370ded585f9c3265c501d7add42afb405e5c96cb4a1021c30dec6b9fbc5203b25b1b9a9102e463
zf18b9ee59b24dac5e5e7efb1e162ca903ad31a4be014b969d232eff8531bf1f03dad7b693c8aec
zb973b6a488f724531ca75642e56296c12dab81ea77559b96207ddbb5c5c12bfd630dc7d7b3f4c8
z6bf377e490c35c62a008e74bb1e77c38a04191a9a6525f1d45b68dcedf87a53f7e847c1afe5143
z729d0d44da211fdbec11f78e7f35802aaf4d3a03e8734797fc6b87ff95c09d3f0d25407467c858
za907edf25284848062f0df91b507b8ce9342725a755412d6eb5e2778550490c1fe04902c5bcde9
ze9c89335b8420af99a0a6dae6a1884701003b88b1a021794cbfd99a0aba4932763d7c8da6c0ea0
z7db1991b663736f21dc7fe0f0f2fdcb97e5bbad19f0f99bbd450f61801e7cd4da31e59d96f697b
z4a333edcebb1bdf0fbd382c56ecde0c82e0d6036b9479bee8b31059803202fed0992d6435d3fba
z0045aa3988dc947ba6b77bfa6e5ab5c72d5d282e66b0fdc781dfc8138f9c0f197732ca43db8683
z16c43956a5532977b6bca94f55a24829c1ce27cfc8170029fcaff1aa73de63f7d4be716db769a9
zbee72e64fac617e281cbc81c11ea82371becb38eff0d8c2e40df54867117a5737f20d77a198181
z0ffad1574a3e789197bce9a7cec933125c41bf395da9a99f9d9507989ef4529ef971e71cbb0175
z18f71e5d60c908914613a1490c932c51af47dbfff0b0f2ac0975c5d9770a1f41c0440062ab8e95
za5a7e968935e36b68e68e0d09ae227f594da0dea31b50011a35086482972b31eae0b67f2a5d8ea
z2930ccb63dad988ab9a06d99de34545b85558c2bf5f26e6562820999887d884c896e0fc32db334
zb6f1b8a14103b5444113923166e15fb70e6b073d1f667f1a175615f3d3d883d5edf5e9a4d2fa11
z24da44ac7dde15d797237adc94c08bce6d91a13fb85a70ca0088d6b89cb1577324c84651c31b84
z4f7430b3ebfac54233ab77fe3928a52cb6477605a2b1db395a02cfd744973e1e96e3dba40337b5
z642cf999494c48838cf4959fdc4e164f7ab5884c81999adb202f38ca8d5b95a2e00e3fa593505b
zc9aa9c11088a1f475203aa7de9e8ba908e4e59c2d0e8c0fa9b5e6e019d05ac40c39271eaf67402
z692b0379afe105ae49c04c008b8b9e4dd82a386ac0e8f8c6dd45c6c16c460e275b5de6f4e8d70e
z4e09d339fc19d84f123c22824eed0cac659f48729b99d95175a52177ea096c76830a237f65356c
z9d5fa0f3b9802741226dd59b4e7042c0479e66ab321f56ad4c8333065759fcae7524492f48cbec
z31bc2cb42226a6702c60a82c4671859dadb25234975a3bcc5d7bcc09d6dad65ff4a5e0716e7cee
z62cc79a7628391bdbf0e14ba750292e5bea7b39ec3910c46f736607c218130a671223e04f52082
z63799873b89943019ac33c62a956628153ef1b37b75a57827dd0aeb7bf95f741a60618b4817713
z54a3ff8cddbe23dbb4bee52174776c7e058459715896ec0194a851dbaeadd0c141f3f589c4da05
z1ced1fa8f85667b152f696997ee109e4300ce56b1f50851cf21f8b7fcedddfcc5efeb07da23229
ze8bda0f897f5433aabb7ed2e5512c6d7fa26c66982a6c0f133a489e07f546edf3f8d3999a82012
z9c4e2fd0d67a2cc72a18fce5ce33295326b6e387a78ddf01892c6eba0b259addce582e91a4ac17
z2974648489745778affb0a04dc010fe62d2435427e0aca9aa7f43cbe32eaa2bcd83f65768d0305
ze03d072e003239842f854e7201febf08e0f127b1a6cba8894f77d54dbe756634596e8fad1df0ab
z1752629381281e4b91e6312ae99a3859c120a113ff0a99548a5283e0ff96a027de6ca16892d13f
z1f2ecc0d81f4d52105325d2cfda92b4de009643304c55488c4c5f6f0c64e52e7b0d6c5419d7100
z1c9bcdb109a29d17d8bc97b84fe9b3ea95abc6589f9b83bf230f518e377954e50c7cc542177809
z716bcb401c49cb381b3db49c1d434530ca9033258630d7988b1c68da974c2c569ffa8391bd49e7
z4f445f909563eedfc51088152caf3d9086890eab2e65a8e7d2b4032994ac903e3cb3de99dbdc3a
zfc186262764f65e2449d71dc3c73cb9cdef9c0d80944b95f14adf770bd0f30e71afc80af5cc0db
z020918ba10d723bf6db3e23b7b5ab75b5cbb7a70adc1658204cf5bca1c34fd39cf7bf5ea9b2085
z831ee4cbbed9734c238403b1fa6d862e3b3447cbe091bc0885fbcd9d91114878480d9c303ab283
z15c88ec4fd7fa030d161071a60cce448257f50b7db4b11037ecbe4923fb02bdefe3366dec33a33
z51b3ec03e193925324992d8c67112eb75b78d45dbf681f53db2eef1bb0b15d37adcd2672976e5c
z954b0dca617e7c35f76e712bfce35e403efee9906f6f62b7e9b2b5d6015b5435e9973527c65fee
z7402daa6181298bcfda0a0c07cf0a0a5879dcccab74dc80fd2aa7a30d4037cf22e394eb43a97a4
za4aa970c0b6c4f56b811a7eca0a26b823cda2553dfa7674b291b176437099067f2a26c2695127e
z7f537b4bd819fef1c00d9b479211bc9dc9be00e719f05aa42089745b779994f0402df4d7b7b120
z163b23be0b41f72c6577cb00e286c65ee2afd23bcb4be51ba3461aad2fd3a029376488a904577e
zabfe366b0c5b12ec22dcf40e42aba609d079ede5c6d71f65cfa3790523d403a6d9611ddf19abc7
z59dea783e325d7e46d4e08436ec521967546e473e0a713247453da633f449184be8a1590d9a03c
z5986315a4b8902a32af751c6ddce7c95df126368463afc141d73e6e995858c9a752a704d8aa98e
z6d1d21d56a5ae669c77a32198784119802d4e5912794907eab597d6a6dd84923193d9bfed23857
zffa96036b3260be4e497749249227efef52efb5780b32b9cfaff084a85edd71d75062b7d7f6252
z32e3d55b8e110781a730539941443d3afe66ec234ad03435f6e0813d88e6ad1f1ddc39ff71a88b
z61ec0b81e71fbe369f019b2c5cc7f2682dd0813bac25671af28ffecd7e0a18970dd7b5702cb221
z7f27cc30a8fcfce01e836696ba8c9e823224ee57bf28cc98c04d473db09d9f2ade111d7f2bf54b
zfb62dc2b90763f76c1fc80ee3053f660704adb3eec2eafb8a7511185a6a5c50c30ec9bd6972da1
z6c6c9108763cdb89b6fb4e6965a4e18a0364cc9b04d1d74ecb9b104b535b390b209652e799bb8a
z9b172760d06d108cf87062124e957aaf1d1a060c12ab975989807dfa1b99654247fb093818738f
zd6f8aa7816ab6397ef51c55e8647c820ecd8d39a37abc2fa0de30ad7a60068abb3b2f0cba7245a
zf0c5c786fb2c4de5bd79043ce8de701a4cb79a2c84cf8c0a3e9e7397fce96fefb5de730e149740
z88c24a999e966d1993a99d0ed8a728bd8733f146d848f1f6eef0a8afb6a59aa4fc0b7f44d6df3a
z750ab1e220077046bd2199767408daf74a92ac958a2cafa5b3e5e0f848879dff0d948d5165ad12
zdd16010f6449a88997db811be585722fea80a01cbefae4027d4f7c683b9446838155bfed3b0eef
z73ad903f7b957229adb83f78dcbadc5550c15fc46d476621d249e1112acf7e6a4cf9777a36c4b3
zf10139c9dcda333ba128ce845669b489625c1d01c10ca2de89021b8bce47fcac7afcae14f2f1ba
z11b4aefb9d339d66fbe25a94c058480451a7147d72586a6d684ba3f7204751c99ce3cf63f3ba73
z1bfe884da4d9296a1c1f3fe226aedd24e81443fde70bd10a4846683ca5bcd01e73806d2c20f99e
z49ae3a1868741156148889ffd005f01648d0e4b3bcb6a737631a09660914cde341aba02200d048
z63f7784ba5727383073b6fa03628e3823262516135deb6bd4ba8b443c2a9711844b288a93d1c11
zd36a939bcc4be6cc935606e416df070cf7da39bbf9cd8676aaf8b22a9cbaae88b9f6b11162d85b
z480f85907805e4c8b31674cbc1ba746485f310d9fe81b0eb6c345015e037a62ba836fb02d45a7a
z4860e5846795d0c540ce837840185e1dc69a35779772c15e3a9a4ba1d163aa5a9e096acfff97aa
zff677ded98fbfff0ac815dc0645a6c8dc9254235b66859877361a28e2b332ba29d847f5770cd68
zf0803eeeb698f8acebf28372c21a60505da8eaa55753e249a1b364a7b863b4e4cef6c8f405f6e6
z7a99bea9be7034527716cddfab51a3cd2b4c2bd3c6f6adde0ad70793448bc7336f7320b2e5f5d3
z3cc21d18f9e3eff22e576c43ea83a8a3ae78dd95da48bf783690f32b0f7daf5aa0ebc4adfc2521
z913f5731e0a543eff1805c7a6e7e2f996decf914d9f81fa79c0b8d0a7478f82748f5008764449b
zef5e6b764d2fadc81263feacca28c7d57295ba83968ebfa60d8b98225b608c16bc07615ac2e7c0
zee5d23fddd7fc6d9c1d5af793d984ec9f4bc95b9d880cf8131fa07f8a89e367750de376fbdeee2
z97c722593d71e2e6391781b662161cd8d8b98da0d6c18987787c10cf5d5e6cf68608bc9d682dc1
z596adabe8b116aa450898bc41340c341870d9d618d948e0f7d6d568373f8345536efe1126fcd32
z7506fc559a6d23e5eb7033e2319574c47839a364352719453e5b91c107032ff107af320ea9fe59
z6b8a0fb563b3b84af113f440265ffd0d29cabdef94bfc02956d7919d6a36c49eaa6d1fd9c0e6e4
z13e3abdbe71bf06abdea3a80558974872b411a6be16e73ae30d44bee7d86b81f253761e7d48584
zd16323c37fb3bf287d79bed38bd092a0cb4f8fc388d918cbe7752776158679173fcd707973559c
zaaa29d68c69bcd220dcbfc98161bcfb668346387306c4cec65713f1284fdb98aaa303139fc7781
zc49aad2e7a09a48c7b35760b7521fc5f6eab1722b01f35122b738ef6fc6754b3f24f9171bb766a
z70df5d11b10e5ba3226febbd2545307dc25c3b9a80ef35993ada4235f474ef0aff6cd00ab1c0a9
z46d62b9bcde1ed9617f3ca4ccb8c85f2dae12e77cf5623373548ff67b020363449c2ffc6a2826c
ze92430bbd8a0b2fdcd9515bd1f1981d7099dcb7164e5043476d6f275b0d12bdef5037163bb3937
z7aa294cb60c0971216335e0215eefe6d6b1ca9312dec9cef6f64b220d48a95e57ebc27bd3932a1
zeefd7a8fe0b3835f3dc6f3b600b4a3c7d7f56e412c8b91b8a35c37bb80115369b02c39408bbba4
zb448d4ccbd5e1c5f7d51302fc719820cabd365e0bfc8566321f8d19b406b6a38404df635dd2086
z8f82e742598c7968947aad9da0b9a3afdf1fba1386731c2348c06ce4b336bd500020bf9375f10d
z11453f6a828fd7af219562eabd6fc56e5c2880d353a5bbd101ea2580c593434fb15b2d86558893
z38c84d708401ff480c24372b1ad71f3ac49b742247a376bbe58f998bfa42331e0573a1ed577ce2
z706ef74fc68fdc19a652f3ade8d852483ec080f39b9f934240307fe23b29b548785791b77c8b30
zc94ac840538bfdf471f650d072f4e81b7bebce1ab04e1d6d1daf6e8e59c5217670df644b85ecd0
zc88d12a169b333807e2f84f6433cc68eb570ddde422e4452ebe6065f469e2e4c28a474e511f06c
zd4dd4f02e1d3e09f17ea8c048a5f9e4ae0556ec0e9bb958b37875f78f5556150494c5d9c23d51b
z8400972a599088487d6024d85df00e733c84f013fd4b03bb5320455242e8c98be1b46582307940
z0afe1350c759f27da9e126bdbe9f9141180fb3b7b1604501cd70ff619ce495da12f59e2933080b
z634503cf0e96d5167b7daa3c627789651704d95012125c0a8d2ad2c7c42d14ca4a2481acf4a62d
z5330fe5c7951f428dda745b45bb567dccdc5cd3bd232321bb5fd7c6780e7350b5fef86665ee4d5
z91460a87809e7b7046ed07b4088d3ed1dbf9443ff81e0bd1e16d9f8a214c093ee108c92d09f9d4
z2e17f052a396a31246964b5e103c25fcc259d9d71613a32f61d05bb05990e95c744a16855065bf
ze0b1dfbdb94524d81049315632ac3b54c471243181aed34fd5c2aaf7f18ae0e013adac2d0a053f
zb3f6fd77adde70407a66ff9ac145c9481579425af9246c3185a0aa0389f45587eb27918cd218df
z47b899961a11a8d85c3147b32f220939d79c891c7688af20f50ca7c4e0d1288dc4b7349cd57e2d
z8fc8be42f380bd40d2d6f11da39b89f24d4d22ef6e1c4e8f9da231d07ec91ba090d4359f16bfa8
z541a78088f28f35d81ddad14792bebb8aba71d6e59ebfad22062ffe8aed0429b84827e2a17611d
z76c10b1c4b8217eb767e40d9422473d008a7b2f42920913d90d19803eef3e7c4d6bc0c7ffbb1b8
z160a0b713ffc9f6d86b5519dd1cb1b900703c41ca36292ee911474e76969ff2c143ad4e112002d
z7499104827d10842b90b1c5c1590767577f229e3e7562ca638816c351283dc200de0ffdc023fa9
z468c83421f75e73b12b929fa673797424f9736368b9959cdd10eeb073c6c48ea3297882ea7fbab
z2d18f0d3c000163ac29a7caf760ec4608c93802e5e533bd0fdea21454c2e553a3da3365254cbf1
z66f9f98f8e9eb6eb04d63d67d28c013afc133e4ce64a8f7429058db487ba4dfcaa3351a085ae31
zb66b9053f9b93ecf90d566b5f8cd708aabc1209bdbc3a82d1f694a3ce2bd70a6037f814377a23b
z6677deb1f004d421dc7c19f005e460d41e6530019ee968906ff101fef3195b3b26f5dd57d257eb
z40d849960ccf8217674c134ed497e1a09789756c27f338ebea949a35fa4b9e5757b2406b30b7fd
z502254bcf085a8de76f76caded5f2a56f8c68e0d69169c9020c6cab9f66553c12b15144d75e1d3
zcec67e147ece68f670d5746f9c514439ba7e0ccf8740b4f506efe1855796636f6c5e80249cc211
ze87cd3d5968a57e2a5b4e73abce342486d578fa6912726c836fa437a79a8701eac92a89e934127
z8875492a2c00cb12ae180c9c5b67fb804979f1db5b08d29ad00111c7754ffda7390668c543240d
zad3e217c4410b9f91be07af78472e80449750d449a17a11551c9e50a514edfbd0d8685bc409eae
z5e817be9a10bac16f4eb0474b8f6ec807c7bb09390cc97d5604a9f92904726c4a9dc4a452d5128
zc512561b3ff30ed3c6ba9d2b2526a5e0e347214973ff2a897840aca2d6232ff13ef703e53ac0b2
ze92eed065d3bf973b8c6268f52ad80d255c8f32d3308cca774413d79820420adcbad23bef31dd9
zfd14e5d3497c28c2d350244cc3bb1a1dc9fc74656527e338b6278f29a9893ba72d9bb1eb5268ec
z0556650703c94aa1cafd7b86eb38de9051b39758c01e446264159b580d6690a3f4a8ec52b6e0f5
ze38ad4f85cae6e5902e4e7eb1d7a0f91ffb7a293284503c013d4f064319834d866d320a97bb8e6
zdcdb9e0c7f5e16dc3048c342e4887e3ec53b07b592bd06a6867d4e86681a64b2fb41aa47ed1357
z3e442c4d4457da7907753a0fb7e380f80601b6a82f9ae5cd6f6f2cbaeb7a394c24b80aa70d0f9a
z2827db6159b7ef37b0fb3acf21f50a6d65adc69098411a524c5e0977d866209709614091fd15f5
z7946e93c12588bb4d625fc65c2748fbf369199dfa7cf315ea57f05324eb06e9dbb98e5168c7645
z3cb942d530b18492ad2f72a1f09276d7059f30286619888daabc323e58ea782a4ce67177b56e04
zf2078576b20be4c87f7787000f990bf9df83de78c51f3f38ae3f04e75616e332a0dea862f76fd8
z0fca58d01010b9c77983158e1b693f3895171d6f83bfc2b3365336dc18b78b6058b0fea759692e
zd61fb80f1a42a3bc985bb7407f68dd10d8f2755f0c3ffe9abdaf6d068cd0053ac6a0376d69fcbd
z8aded94ed66d805e2ce3b1899b964c2e2d7ec0f39af3d6324ba6f9774f6ddbc79c6cbabe7d02b0
zeac826ab21b86a83d7e429557ab59798ec178af2818f131922ef4896cf20a8bab15443ead4546b
za3f369eba7064b853949ace352b808d3c57e3ab1290e077ceeaf945b996dbcb55e30feb9e4720a
ze4986d220310d80162e4d7983024ed535eecaf2f3476af849aef56c6e4e2484cffd34989b5d75d
z83bb5777ad6eb872f9800512e9137af46830f364009823b68fdf93dfcb2747dc47d10c6969b116
z7553c7b75383e937bb1c08eace395a404d0cb75348264f27b3346b6891cd0853cac78a293df99e
z9e1f4709bb8fe4cf4b1580ae88add359ba498ed963d5b938b8db17e94a270d0088d501d8677543
z49262bf85ec4d57baeca759f138ec71037b3c89caf5d8332ed3ca97aa6f12a9845bb754d562974
zc7081ce01544fcb9338e6eefd3dfab585d2fafaae2fea3f4edb3561c4fed7b703f1874d52f0b32
z62db2b42fd34d412fe1ff00d2ec708968bd07afcdd02cb723173726b78272bf77be9449ff39be9
z27b3c3a1e0829f50a9875ed843d287ce926b575d016107e44b69fbc9d264102caebd90d116407f
z6e835187e8b14532483729b4c997ba9758436d2ed00be857ea7eb0ca943613879b2f4ad763c94c
z503977f5fcf773f7f9c0702a997bb17332307d1740a4ce8e042ab6d491abd4659bfb34132058fd
z8f3dd3d530fb6119603960d432f9e3bcf5ff687bd06d4c3c1b761cdca5ba466f8942d14e158eab
z61f1093d464fdc78adad9412629ea5230d9c3c73ac282fba970dfb2ffc84fb4c87854d21acb252
z7b56b1cd4b3719595c8aa793242b53777c4623fe1078032be430adf7d2139917d318326abc2135
zc1da3b5034a91fb1dd0a6b65ebf15e55cfc3ddb64604ecf64c87ba07c66fe6353665929ea3953b
zebfc2cec5386b5930e5c870dc3be1953937c964833e40a21985d6ebaaf98be041b6dd59fdc14bf
z7fd974e971b9332508db26bc3796d833aaa14c55ae965273233671329d1bdbc6e30341fe91765f
zb1cba0a96335bc33ec5d37f843f3599730ebd403093cfd12e1d6f54c83a069196cd4d7a58c3964
z3a36492243a7c7f367ed96d991111e564ee070af539c87642e491e5d0f500339837cb2fece5de2
z6f2045e2746330e551f001870ad29a887340211509bc6576962f82894d4eab210e88fdcb2eb34e
zdd0621fe35d377f1d43cbd7e5e1351fa0016841dbbdcf11347f0171d6a184f3e52bfa01b9b6386
z88787489574201a56b8e61cb753f5465893495952a9120bbb461039f4138c7b73f1b13f503c77f
zf6f1fcba50ee5068df83e39721f22b69fe2028efb6efba36352d6aabcdc943b048032b1b360815
zf347b12411f240b54692e49c3b0ec498ec50cd4092b008f4dffbb958083a3f17e774bc8239ee0c
zd9670e4ea5bf696eeadd6e21cff3102495662794a8dac5cd31f93e0a8b171fc5f3828280fb174a
z1fef7f5ac12e13afb377330157aec10f1fa5d6f1c1b9f926fca18e62c9636090edb57c5ddc732c
zf5db0120ab4f5349a3b22f7c8c5b8f5d690e0fe6e4386f60b479309437b3df795517db63e201bd
z8e620e324db7b670b88b9c7042158a86bf08ff1440c1d3ad6565501d9a016ff9a47090233a6498
z64d29729825ead9888f70a96d31b3a5f566472ab6af22528457bc407606552e3f452039ab3cd1c
z61ea1e75ea74e7e5fe0c7faae02ee45cd1f2b4b29d0e1d5b671c21b119c03e26f401d0b6046d4a
zfe6bed67d456c05159de0b9fb307182353f51d7404729238919e9c2d11e0dda3b3f6ea347d04d4
zb6642051f9c80c15e50ac779f402bb8c9e34991593bec99307bb44793e615ba54caee362c601e1
zd1ffd9e360f1fe279680fc1c416e1cba7b518b68af986ce8a68f7a558263169cacbfcfcf0185f0
zb43f50e8819c964906e92038b17e934c83ac9ef72c7741b25655dd73177621926069c78d77be70
z1b4cdb24cb6090acb9ce72e3738118fcfb68cfeeede11648e75567a6d6ffef31f3d2cbf67fb3e1
zd1c8c9e40c58043dfccda14cb53ede8ccd938c4c5c65e9fa7293cefd3efdbac18603de1b032641
z96c921b45a954ad231022e9e729cb4c72c9026a69836a954032220c86a96c61d833468c5bee0ff
z1a003045bf8fd17d4c1b3a3ceef2498d40272877efc436edb68d3c7f31f93b0d595061175fc33e
z65064291ea39e7eaa921d69a3c5ae3d170372e45c394e045f7b1a9dacbbbf8aaf3d408ded48bfb
za7bae467a350518df27a9f5b40a1ac99d5938fcf8c8af0ffb3d59a8e742d48bc41ad9a2f9cfb13
z0ef315854d249e24af22745856eb934039ea90168cacb80308464c997598e132d5c61df2e1b93b
zb0543b12cee1f3ed23e067899a4fc4a1d66e9ec3184ac541698dd43e0040424eab7af8e77ca719
z401a2ced3cb5ff6bb8d23f5d397c30214e900ce530243dacd7ae6a2264bd0ce43608a1306c6b7b
z82090c68a70f683611cd59a736c2cd6246054bf701ce9b46dae53d9043bba5d179327124c60653
zb953e8f282ca07eb6df6e8682b3284aca1163faf3e900815e45d8bd139e546930932f9bfa4dbb9
zaeec932a7f738271cbfbfb5fa993749210141573ac2d5650d8020168b6c784db0263d305103850
za86021df3428d2d77c7cbf3fc76a1b85ae874e0016c2d56746c40dcc8b0489cbf4a7d82a8e49de
zfeb0d7c337e6e30f2a3a4898c4d1967c661678ca2f964239a5df57f6dcce303cf5ebc2115ccbd3
z814f2f23411a2292352155773a2041b09d4b4695854543b72fee472fe49b38e13c49ab9616ff91
z803da31421065d12d77ad677d265dac104af6823f52b22591e59afa1e133f8c70dcbf325072dcf
z9cda00ac918ef6d1ed321e0fd53c3b915c027e8583d4b3433a65548ed592a117b5b81e546abc2c
z69a371a8fc690651ddabcdda3fc6d4b7a44231e74fa5baafe0f4ee9a58c379c057b871fc5d347f
z35316b2281de0e4eebedbe10b72fca35e0a8916f314f6b80b11dce54d690ad982eb81bf814f5fb
zc0e3bb8d7cf41bf973188146963a772f3dd6dbbc8d2a255d606630e0ce482d8c23662758b80a4c
zb791d25142cd89a1a82ae898cf3f4b2d0a372591f52f85787138e49abce48c4ea926da866963de
zc12a31ad8baef1dcd958f8a073ba5cc4af22f2b287d94eb1cc0cdc74de485c3b9777e58aa52a72
z15b1819dc22a26e68e6e47bd88cade50a538b9e8915a1dec08d5ccc86f31c6ad6509b277b70156
z6e8883a94e727b997055dda389513160c774e1211ad7dbdc43a856527f881115af21519c824b18
zecaceedc566aa034855af52f75e88e94e5a1ad10eef5de65c7c0172369ed949e6ee55c4abc3cb6
z2aa48c64ac0049f7545de1c9d35c916384e2ae805c3af087ac73e8f5a4f222558eb0155471ba45
z7a94a2dd90bf44a58afd1b7f74b86d0b0609e978751a76cba8a4f99c51b14fc5ec8d6c3493440a
z807cf262210f72694203c267bfcbfc5dd4b782808edbbc757f42ab09ca4b1e5f5df95f876c4948
z6d21684c3fdc1c0a8379696f37aa7d43d51c3ee3856e4d607a0c0388c1d2b6babee57090138409
z4f8bbd0232730a17885266e59ba65732348040de47ec7777c3247873ec6ee120454d06e461e1fd
z6b5fef9a10d1e350c64e19d8ed02b1905cb206008b01b232bc5e1686624ebe7da32250a6ba0e88
z4683bde5f195081989e15dfa9408074a96c1f621a8ef324ab37c7e614901529aaf7fc0e7762cd0
zae8ff2dc6411570ef46c44e583a953e30c9aebe619d5140b6a9f7b80ef6b9ce80b60967449eb4b
z3af511c05b1a4d7cda0da7addd91bf48367848ac27fffaae3f4ed42d3550972356bb0a912055f4
zc08296d549201c4e7765f3dc9125f4ec1463b735150cbee15973c365a7f147980a26c368b5ea2b
zafff413e9259eac4132d7f66561b31245210ceee1c3bf56c4784ca5b046faeb5385ea92a0ecd39
zc08f26e798a4524857888d56d9db1d9c6e0c2f993d3897f77e932ab0c20ba11e6fe0f6f8d1132c
z71da6b93c80671b5ea7706beff676745257c69aec03311bdf894e88f5904f174f7f429c5a66823
z34d15033f3764e9b7b9aceae68bae54cba97e77430510ddce89272ad39bb1f696f0132f6f7996a
z44dc5481816c06cee81fe6faa62e7e07010de16fc0c44763bb157a9f291c3c9bb8423a0a07a7cc
z943bc42b732907d01e8d7ca259d6d3d2fe9568d7e618922b2f956340bbfb2dd9f2c5f32bdf37de
z6322005558095c3644f426866e0306284ddd0f0316a822f8153ab9895bfc0b899d318675411e72
z6910fc31134b70abd2141ab55082da067dc01774d95239db5f6bf5ebb5b01b158839abfb24baec
zd24c96030737f0322fb78b86e9fd2a6bd971983ee419bad0b6ca6617250380fa47e7633075fadd
z4c50ee4cc27536a6e0487a9c5e8a8c0743a50a15ab38d51725bad485792a049c47188fa3e8d1d6
z032f926e865ef4bb5c47fb4549226f7b324ddf910386f72d745c6365a74a8deb203c31ca457581
z242bd002d3bfa7bab543de1aa9528cd77c0b3069238633e541c82e518468f2fa0160b582131b25
z71f2886f4c215aecb83a6d8d244597c89f32cee19fbf2e1fd94aeba2508f4165b29f702a5a5734
zbcd4f5ef2e7d2a0f158024096aa6ee034f4682a95bc3dc8f9b51fe9c235e3b33e70fec4f7ba8ac
z84324a4149b428f664ac72f47e96912b000c98a1600cc40b8990b255816855ce69363a13dd6842
z35c205c95173fbbfb3ef46352067e0993f261e94b872137b503ad703fc7861cea9fcc31ca7800c
zbe09a1018bd41b0358c18c7973633bef4a741e76d8d826b646ac3dcd4753d87fae472b5e062c08
z269289b797c8b084719eb918d5d5ea400ac0bd842334a53f2619b25d18b52e30d00f33f17941e2
z9b5e82c95bb40e685b3b67118d3ccb277743b64ad783818548542b48e84d511590b498d6134028
z47f1e3f6ff8427e13c792f8ac833e7affedd82c8f8920b4dd7a2f6efc99cfbb1fdd6653b710756
z8a2fec72ba2e20bf41ba4bf98152cd6426fae8355fe89b5113be1ea93a539d004647286f0e0b2d
z4511329ef9e137e241b37e73189f24f728103e90c9cd0c55c80c4c0bcb8cbd8f19e5a068bf162d
z35ed97476fad48ef1a4bfd41ada2ad1951321a697c39a8ddb81093d0250e42b6f964a0fa302f41
z06f1350dd5d889fd3e64a7f1ebd6a1fbc75cf7e32073822a2712d6b171917ce24984d52c50c6bb
z382c5abf94238c434f090427a3dd6d225d6c86addb6c1fab7e116b002ce58e5726510311f46a89
zfeec1546968081057eb0269d3c16eb3883dfd727352b267d94d9fae141059aa788fe0c381dbc7e
zb6e950f961018a16e916f0383908fdc002fd2302154e3f6cf1b163e13e316b08e1786e45ed9921
zf6ec1a12971de9439d4537a9d340f4bfb1a1302eeb238d4f161aa575e80545efe25bda38d66e04
z944e258c4f9782b9012467f4ce5dccca7534dd9b1d7b830b1a51f6cc38c0b085aa2d0470ab44a7
za142e76a5a414a2f2887b6f086d1757f5154e3ae43bc97bbc1bb7bfa3fdbada125f879a6a8c708
z6de8cc47973faab015306a000022c2fe940d55289c0db439c1e9a8762f27b51b31158b7afe3669
zbf24206dd2a18b70e5d5e9218cd5a04285089c9771330abfcca0739e344efffdb1b27490b67067
z11cd6a6349e9b523ed7e0d68239c1dd298134045ddab1a0fa0ebf7a9b695e4879a4ce05d8fd48c
zbe9dc830337e6d6ae5b7c2994a50ddd7d7a37f56e287b42af2af9b3f20acf72ed6fb60dddda025
z510f1a8d7d10ea9cd356d88f2b7c901ee9ba9a05c38e45f022e9cfe9f7c5fe3ff12ae13ab4941b
zecba85f7bd09e91d58b7ef960e8af6ed43b05fbfce8ef5ce7e3dbb4ca7a1c7d8e002e09b75c4f8
zbc539a982af225867794a5bc712dd33a99982e4140cb2d53ac58ebdc398d0b1ebc52620bc13521
zb9de5ca3e7e6b8e5a73b9d6720969cbecdbc3f4152f19747deb2435b279da9d78d05bb8e2c877d
z93ba8aa55f57d3eefdcb2a7b2417bbf210f37e1016c88c5a8951df96e057429a75ad8e5946e7c0
z22768342c48d181568aab12e172796f40af3a16dcf94e7b49c8631cd1869eacb829d450a22f20b
zb5395f524efdcc3e949b60e7ba9a0878d47d30e0dfb21bff372f232850f944c59f309c79a14517
z32d1fb54607059fc15c5e16b058790f6d0921c4e3cc37db2fbac4d4163fa54533672df49cdee3d
zd0a9c39aee0c6cd36979481e8c5356778aa8bed44b9ce669a9f443e13552af8250a31f7277e35b
z97e561b8a25d1eedc68ef89d0a25690e00e3675916b55d23cd2c31404e146a30ac2c812274a67c
z0dd5f0e83856b69cfa7e6e8b5a53c4c0cfa06d1bf2f487df1de1e0d28e8cba9ae38ab90f288b53
z3bdde2c0eec70702707ac6f2c78d6e8b3160e8a7793d3e96faf2d706e4352801ba03e53b6f19b5
za06efb08ddf983756f0b9a0fbad965aa97dc4a2887309ed9e44fa7b5504fae06440b6f5a0350de
za9ab2777290f4972a8ed14634622a93681b4a577a7ba00965942fa8edcc2b809cf0bde2969a754
z1b10bbf722196b934b46a928adac8694cfceed6e38c9ae1ddb653efe8c014692a051ab37a7669a
z336bb6b25d6fbebd54b0b28b985909dbfc90161de2aad02fa053d68668f048904efb108de69f4e
zff8997c5d596d3f7a73d41ddb0f0b56154deda2781d328f335f13cb4915c483d46288b89bd2e7a
z78f187e49b5fe64aa9d9d6f0408691bf1bffeecde81a91e3d95abb6799cbc9dd474c2b193ab27f
z1c0eaf82d8787233c1b872603181f5dedb6b9c05368310c1a16e70bb12392362a3e3a37464c8fe
z426cb76fde725e1f4576ab2639177a79045d43beb496f887c363b7e8a17734040e2732a72468af
z61657ef6230cb864d80481273f1719c3e91e23ea4056d6e096dae4391a52b7cc734158230401cd
z6848168dc12d664be496cb04fe07c6d41b2c48e4f6e4a9fde9d5cb6eea5909a1719b25b0647725
z1ea34f86b0e5cd12f84af8be35b9596961fa1443b2759a11d5216a570c828597c466cff2fe3149
z075bd71c70c0dceda3099c3343e7a91847bf342a99e5b50d7d8292bb980cd9b37ef070f581f2d6
z3d2c91a0518ebc9f013d8cc6cf3cf93336eb829b507173b1ae3fa4fc22338468b28c09f9acb5e5
zc79f6892cec3ca27da1b176983459e37d618bae2e489a2e729154e08b809b1106eaa206c6a28a7
z1fea83299440e6073b50e367294bbea2a764268f43b8f0b28fa8c20a36a8c6cce5b9d245e9fff7
za1afbdab47fbd1101ca43f785816e9fa4c20a71a1d91ee13be2911a4edaec80cf9edea1b722039
z80685c52c0226b57e8c4619d4ad24b5e5b729c9fa635f117fec0741bc819689088d662cf43d3d1
zb5056868c82073791eaa230393bba663462bc21adff5ac9495a76c4875d3513c3ce5414f53aaac
z7db6a4229d1a5014979260427b73cdc2980fbbead7869a7666a37b1fb7b735d7efe7983d5397fe
z3710e2b9173455ffa64c5e5004a51f9de73fa1a9c816727f1b6466545cdec12d0965b1335d3194
z428198d0d4899d2444c2583485ba42d3b5de4fd710d77f634a927ffe990f0c105ff0cede26caf2
zb3c28d6f04f29129bb09a26bee74444b4ceb3ce302f9de1c4b5c55bbb0a23540ec1a6e5029f5c5
zf814d562c571b4e0d3fa5c917eb13e94698ce5ad64375d69b6396985068218e4318f5ab9ca1269
z0449e4b10c464f318a944c921b2b0754f0b99a83dfad511d1c8e862f4573347ef9cff2b91b5804
z8a458aa17d8aec21e7002f439fec70a8208f7311daf7d25a7af7efa77f39fe6a68041685079643
z5ce03f1fada70ae6ff979c22d1d1abea2dda8810a299b2d2142039acd4e34c4c764c3b4abefbda
z5ad55d38cdbe984926b764bd1ac9d9235880a56615f096897f95e41db83ffdefc54f9145ff3bb6
zaf90dbea08f34b0f1bdcc4047d319e708cf7f439dacc3f1d3dbd50238e0f1a6a9f3e207861894e
z0e18cf0b6cdcd0a59d274bc8bfa368d4bb1235a16658158047cc2d43f965809827fc4fc9b6551a
z2e402ad2ee94769d6fe6331bcbf84f5fcda5caef1d99a1c1e20f23b54144bfa19450352294b876
zbfa38e4aaa11dc768a3f2246857d8a61a5d08af13baed9afed70a13fbf8cea65ed860ff91d1dd9
z61fef4d36b55ca1974e146b1419c9e082f12e6780a5d6594c8ac2e13ae4abe7c933caf921e6d83
z09b10c0ddb3a8f9d7499c0b8e3e99e6a927e59f6ebf1bb13b7b07bb671d625a36fdfe602465d6c
z9b592b1028fc120212d6c724b9b55d80cacb3460358d12e387ff6034760bb772353a98890d580a
zf659ef3b19a13148dc2be354519fbdeef54c4365f16336647e6e42886aed09c5d1cadcf3084a22
zb7adc7678f3063ecaa9e6302cb8d4fd52065b66e4f2926d483850f79714f029f4f7a225128a21b
z507a1c1c026a0d3ed2f3733a28fa0e3e7d96618429ccea087aaab0ce1a767f4fcb358179420e80
z024ec9ed372ec98434ec92048b385f61583335a2a7baba0dddc1ae90214e2be2b5f1c32afb4408
z39f30d6412a73ad4a3b0c8be4b61b74000f8646645cb5d85cf36b8f5360fd4a8066bc8720e57f6
zff25b09bf82511b20d10de5902b4f0db5e7c9d0411992ae1e4aacb08347336616c2245817080f0
z3c96474c6ea88f5b35a839f9b0082b9948fd44a82a0274bf23a99d02590c029323d25744ac5829
za067a0be15ded471fdfdf0985570f19e59a9e72a7400d3894313d761b6c9ee4d3d62d42b4eca22
zf3a09f2d8ef2e670a212472358782de3fc5d8cbca722a856f752c5f747a86f6fc01158edaf40bb
z939e70b249245b52c82ffa3ba0995ff47054959860180b106007eb0852e790b2ed7c50cd1cae5a
zaf1996159e56ac0b9432465e4feea22e92614d20e9b00d8dcc38a6b3444e08cfa76de04aefffbb
z01e36e0f84fc3fca8faa9e25e3a2183d626346dc21d336fd197ef1ea9e98d33bd890d0cd7e2d5f
z98fbb9eff4ce4ad17093df1b88b4476826c3351dec5564fe058525dceb083b7886643a77e97138
z24134cc7d7780bb5a5e5b6f0d11c3767ab14e73af5716e61a31c6044e0c1e0cb173a9be34657d8
z2db1226d5d92c7974df29675c03c80dd390bca16c83fa05dfc28a9743a6ce889606ac5a2bed2e8
z7b65b7ceb89d3db8a3bead11b0a024e8a2cdcaf5330d8b27db4d0c8533b7c96c2c6ba760843992
z72de348697b6df8ea2bcdb712d416a1bfbd2dca26dc085e53dc634317d2bfc7cd04d4ea4508a8e
z9ab7e3cb5f7a6e9fe32f107d2441f17e9e2279ef12ba9b9d54a2481c060071efe37e65e0f58f1b
za895cb3af5f784d97d37d2ec406d27f61817cd0261661752d8220bd53b3f54846f9c6186ef0612
zab41bf49892c2b89cf61a894ff33e73283a56bc498f9df4e1e902c3e8f411324a8cb1247d4e65e
ze4a5a98d8cec8ec8cac9e876125ba28baeb70d5e6f4cb99a69e2122e34609a4b6779e240d21525
z90aba81e5c5fa29d063164dcdeb7f4e8ab9a38b5af07ed65a4c507e88d53c5e3d6d3aaf8209565
z9bd6e6f57fe0fc39a73e9fa57b9dc6fa789b184a8cdab6988539544504c2b3a5195403fb174fec
z8368606359f1bd41fdacbbdcf7df127b25a7341c444e05e969d8eff054edc459f6c6af09124b80
z0e16cd18d1fc3b0133008ad179bf302036b39b2bcc4ca8a7e1df23bbf5b9e50c7dce5bedf8ca04
z803f0d038410db57ad4f01413d5016e8570219bc27f7448b873eadd77fbfd117f1a49be200b56c
z848b5d3fd84fb9a1b804298a66eeb2fa08bafb7d74ed05d3ed138bf77e011689c8452e751d4134
z2b64f447c4dabc96120d0e1391293b23ffd18747f77991bcfa03b68d43c9f9b9b442a1deb4d756
z9b5a2665e6c3c1e261e4f51012114defa19b9e88a4b82e323a03c3559cfa43cb0f7d5a9ed4f361
zce21dddf48234ea7c20a9814e92c22469ce31bb7c2ad6a9e827e2ceba9ca404389a3346532938d
zf561a1e383a6a59dba0489c2433a34fa59afa4f8498f129ef546a8ad937b936e1501d8cc89bad5
z94e20759340be872544a24bb7d7f6af6cb2632f4668f664d8957d1300ae325cf01b02295f4ada6
zddb59b734e7fe925f964fb304a77b18f1c4695b5ea479ab8834f5f29a188253082d85611081a49
z140cbd1990346218aa1b2d8cb803c26513fe0b911b2e4734d7587c9eb4b3a636c9662adfa10305
z205adfb742f86c0434823e7fc7e5425e6d56272143a67b411d917cffab4fdbe7780dd849f7f3d5
za98f168bebd275647181a820bfb3dee4395b5e6264184ee599dd9c2e25b71fd7c0004cbcde8d27
z71c35712c0031c0f91362e279157d37d8268af13b7fe493ff7c3203914aebb03496ddd5fd92931
zfa9163be4eab5f9e78cee8563baf4baf4d94037e7690d3ca0d5961b8f9b68ed75f28b3ed477f75
z1d875a68a93f5e2b51df183051c2fc0a232537e89de6fa8bd04c8bb05881545039fc07027386fa
z8bcb9331e510331f04397a289451af59020c3916dfbfbc5dc0f11cc8b8592827af7a347e0bbcc6
zfa824366b524ef52de44a6e570c4544980b0dea492363c72457aec315a2ddacb522a52ad2a2241
ze3d184562f8319e36a31015d9a9a8e1e0c0c2d15ac248529b418455ba6d35645506579f1d973f9
z3bdef9d3aa9f9ab553215de6668877ccb42d682aeddb5cf56af80930153bb8ed4e252da401d4ee
z0567f7bbeb29c27e8dcc2b8f4fbcc8a7aa5016cdbe7fbbca22ea0afa0a82aaccde6bf0069eef10
ze3e9f62dde2878159df193bcfd25162a5caa4b8084aa3b495c2a18babb55e11cf47577ad411ca1
zdffb7f1f09745646d68339232cd6a3cd36ecb4cc04afe69b934d14716b54bbf1037a07fe980c20
zf81cc48dd01e2f5d4eaac5dfbfa7038e23913a00812787ffbe4cc12df5e03c53d86b69d13e5c3f
za5dbeda39c5ca96aef5706a1ed14dc172cce5313ecba5bf57fa981956195c4c1a63c5da168f093
z014e680eb91a45e7b3d5ab4d6496240b1d9ed209261df71248f46cf8d9e57e9e4d3b6eecfb5c31
z0224e3c5669ab5379881f7705d315a31587f87d11957bb912575d2f831ef441632d5d36086ee38
z1774202ef44a5039e59dfcf869c853c158177915eb07f73704a87c1cb665ff04eb326c90b95afd
z5ad24e064284576a4e79d5fca34581257e826bcded3564ef124df49fe59e00ab56db569702ef52
zdb178d8b8f01d6c426a772aca1cd4bba19f68f73da7e23e7096ed901a7c69c0dc5fb61e674dbb9
za4973b036c62bf3e7d8a4f4edeb10e1fdd751a6ee80d55dd622d5155bbd7a8649cc825ece4f1ae
z9719e2652745ed4fb208483ae796c7678a37ef285796d9e668b973dbbc92e58c631a7081a154d9
za8dde91b4649036540bd270353e41f489617efedaa07db53cea24f39c188099c235195024ff5ed
z77d1730347b61ee93937d51c8a2448cf4f4722675373c2c96a74536f5d9e410bf9df20c1969b4c
zf85febe3b93877eab603216e246adc29ae69478cf3b8766dfe4c54f302c9114dc53f0e4f6bf5c5
z8202babb2aace29967aa5214ccf384b038a85ce6361aefd463c4805a6aab01c0c657e2a4fb2308
z5173463af947910f068370a8c8639074e08d7b0aa4bdc79fecf802dc68ce3c444bafb8d6d5c7c1
z0a44344ded9c425bc901cf21f53226a261ef23450ca6b10b1f4169c7438761db836f6a95f09444
z1b38adc0f5c858a2ef6e341217e305a9bb2f4810d17c931859a45c4f119080b3cc15684c4fb01c
ze920dae1650ab2580f9e9059b85b4c432234a9d0646407a12f5a0a3e5945b837a0b36e28ee6e16
z549b2b6e2e1fa0f45d61e38574b7dabf265112921afc1103ec26b7b2c162c046e321704f4a206a
z88fd5f20781cec65f3fe8fe3d5e41ee90b7464ac16e3a96f031a5a275c79f026367652ee24fd98
z928c30a7be4eade67ded10806077157192c1932372e4806fe197235aa5f3f501334ab9104f3f27
z989c77a3efdc33aa0f1bac58236e90e325e1dfb79ebde960bcf77cef630cd2a2903bd4beff42f4
zca9d7488123194274f9b5325e391fd932f069a98ecebdf61a97cf0ceff683316b6bd8ae423eb9c
z28157c6477debc319292cdb0a77ad1b41490546aadd3b0dabcfdb32e9ce18512d47a98c67edfcd
zf0985ba8e1a0d6ff721b310b3e0e1ab6f3dd8a0de42e80e52619b3cf83087a789567e7cbaaba95
z4ba274739a475ab8ecd2263982888f09ba749511a45399bb698a24edb0e8e5b0bef888a4318b13
zf529bde43d0e97f884befde6e0017b2bc1e0280553446782f4120ea060c6436c64d1a807101f5f
z3a0b195fa050d2b6ea23e766059d2a958a6417685ffedb92d616697e0b3979fbab7743d554a031
zb958d4131eefd74f719607cafbcfde94e1563df7cc8cb7f81601cd170a76daf00c80ae623e66ad
zb9928045da8bc52ca6c148940c7cc44c2f85d20269029259cdae378db0a6a9948e03751e27b810
z36ca9fa0a86b33ca55545693a3dfffaff49ba5dc32d5f285dc0173c39b9c58e61c1f9cc9ec6f19
ze053d47c141d91a9455bd6e9210fb33344441887b4feec8aea016b8b15ee4773f59689cff8ad12
zb2db8a1c4a7c09b31443e9b88a6a4d0870f18d7c4720385ef526618c14da76361fdf3633fb2bf8
za6c2e5eaf3ae1ff3b6ae58d7f63c5cf43b45f5a75038f9e8eea95c21bedb21608eece900b67ede
z2760701fe70b1c83f50d69f7830348fca061664527d70c352c247882a46d9c2d751f0dbd3a129a
z225f225cadd5b5c05a5252117a3b2dac259a7e1e59e29bd67156c886b2242460b0620c4bb13ebe
zf3fe5b2090d5df789e61098b873e39b147d4fd4242ae613f5638948b6f33f18845bc463b6aacc2
z7c89d41284c04f5a15e0c229345b23e377cde017cc0c2ae28d65df3c516320f4f9eb6031a715ec
z17b9c6f455a496a2257a6fc14228a18eda3814e399be6ccdefa2df0aaf42d5282254022e32ec11
zd79d170750a567af6d76126312ff16f857c27b1b29b3ab916afbbaf61632e0f9b6aaf9f4783797
z64ea737282d47da4012fc139d5a663401b06d81e2dfbc61671a1f39aac3435fba52e7e0cfe8625
z051f84afe59e6ebf22f30a02154b568ff1404b9d969006282e49b311d39cb6a7c1fed129a59451
z47ca985ba4640803299ae7c2dcc2f4caf40c38e68db5a8a9e4fd537cca8f11333c54b676fbc971
z053b46524a586ce4763ebcf9e1e1db68d0af4e2b291c83ad631fd017c085753ca7d57c38302a70
z77eeb84db72bffbfd858cff3774e9c7d993b7ece67d0ae892ddb772b00ef6d795b7b22afbd3710
zc771620fad131b2c4d3251c4c71be3985f6ff94bffcb7f5a16eb37f48036de541996fcde0f63de
z2705ff62c272e1c5b8aeb04819fe336ffb2192086d342c06ef8898074924cc1ec28f22e935f1a7
zdd46018d5bce4c5160cd295ee2a8674b824e946989954234ec41dbe869018ef333c1f5c1467a87
z6fb8d5ba0cad36a8865d15c0dc23fdc2eb56d38835d1fa3c2cda660693122253fbd4f1c05a569d
z92c00786b61f9eb2bd393c91125d657bdc991240716c852620d655a8bbda88996661e914502cd2
zf3da8b0370525ca5fb2e7a60328978852c62a5226dabc393b1421560171d79b95c19b2275d0f2d
z9059e935322671d7672cf0db5d620c1add1d52d475e47068d97d3effe3fd4781f8db045f6d948d
z7f1ea46845317a30afd65876ea1bec05e282174b8229f0be57983e17334e21dffdae293d531e4e
z0090ff9fa1e178ded2344eb780521abe3775087036192d390ac144059dbec359d7ab48f69642e8
zb894c243ab034400809d913101c6dde9c191d150cf367bd54534c5a266f05377d6138c6d442fe0
zd6a976e1ae60bc84d8e1e4b10c9b9d3878a63d4c4303ef8ca49e284811764f8d1a7bd91301e914
z0cf33b6edb68ceb167e5b13debc2f769b5f091394b06c5686b067c8a0d6652ca5632da5d8c9021
z583fe541d25aeca35f3781f11f797afa28f123e3af5fe5907fb7f8bec00672ef17d3f82208098c
zb9d9c936b0b3343579ebcf77452ae5840bd33b2fbd51af954c0166ab2f75bd2107631a1d90039a
z5e1e948d87a1bb8b5eb9772441d9bcc70c44f48939f18107e40a6fff49406a62bbfe65bcfba30f
z0ba108fa3ec56d05ea496387a2ab697757e07f61751c310695c7c5af98ad29ad5d86c7bbf2946d
zd0a73dbebed10a3b20cc4e522202c7174b9ca9c3a5c0bf6ad0845fefad772b88d3fd2191de895b
z4f5e0bfe18d135cc87083c7d0f48db8d906b80a6bf0cb2719485784865df6c75d95bf070e178b9
z9985d6d1f2e2d5b5cadc7467b3db9d2ff9ef8869af5281ff4637eb18f5c1b044a9d26a44b43500
z7b1bb1499ee7b0f76f2b122c70e1df421d0e26ac0222fe1a34dfa7f40cb73396f69b4cd81f6ad7
ze648b74a39dd9b7da0420edd28ec0eb3d19f96f3a880fc59c5953b6ddb81c9c022c6ced72ebb33
z86f32c5ec956be13887992fba30f48abc3ff51d3ae47d12d69e4068bae33b278dd661fc9df1938
z235d0c51d172d12aebf819d109c844230473ceb7a0d5a9f74338e9b5a0d2893ee75885e1367e62
z1ab20f1d318815149e8c184fe13c289e26235fab7a184ac8984b400d28849bf41f47dc173b3c0f
z30003edc2b8a90916a2abd61a5df845ae09ca41803ffbe19eb63f5f1e018e5c76b86858b72c42e
z0b109c931b30d3933843515622ad34b3f595c8d5c4e512b61496a396e7908fe35ee8262430b3c1
z26d62ccd1d29974dca3d39d7409fe99b7608d0fd67fa3cd8f477304688141bb35df0caa72b5e59
z86316d22d72dc5f4c8fc84025bc88791a0c79b30388cadb73a98ce78beb354c7f98980ac8fd472
z1aea7989b6fa88f6c30728e9e1712d60d2256430129b957eac39570805badedfbabfb93e791f76
zc1ff335ff9201856f6c32d66522937319787c27e4f478fa987987674a5057a2bde063247ee2ed8
z0b19eb054876a8683614ebb8c308388f57b3b12075aec9167c072849bed82f44b8f8c9b1d0816d
z0ab3eabdea02c57e23104edbd37e7cdd8cb826c22d533523bbb8e612d962054be3feba38095003
z4c88042265295aa98f0494b70c81d3163049c4aaa736ad90d3cb59ea8e5c3cfee79814e3357e88
z1dc7d429fce421d387fa7f0c366f8206e99ab4288fd92e76450552f0aeab4668d5b6376c3c1e4c
zfbdd3e5a30b1aa3d1ff0405d2fd3ebfbe0969dec5f2773699909ea8426c07da237c27876cc93b5
z5426c4756d34100aece4b770bb2f5ff828d284ed32fd8ad6a03e06999aae2dc6f385f39ee56e61
z536dbfb52e89e675c32858ac38a79718f7eebd26ce8e60be5c81b74368ef02da1a0acf44b770e7
ze6ccb03948ea0c4a5fa1e1bd76f47f69c5a93729227db986d482b5858d38cc7fa2ac012b5dda34
z73d363b8b78c95390044eccf92555d5dffd72f9545ca395146d55cf9a2a020b850d7ab31d668aa
zaf4c3f13385a302448cd382911a897655ffe2a9dc6599b1fde0e1a98277998e7bb4f2cac58ab2b
zc52d5b448b9bcff39aec7e1424627fa68000de6423fb9776af60b6241c3abc57feb242c2912ecc
zd8f6326dfb127861bafcdc81f26f0647fe17494b8a4251fe3a4d24eca5b5a1cd13de45fda5b6f2
z057757fd1f701642078d5dc242598748999b80059533482d1bc4879b33f0e7f489623b619e054d
ze1266da3cf903727cbe1589aa4190c53de9d2c550817745ee39ce5a7c983c3cb15c0db280e32f3
zee1a5b22f584bf09f72f08e9fcaa5bfdf9d11ef20c83afbaf087d5fb4ebc4748e6b725c3e3b85c
zd7c23689e11a72cbb0edd802024d6b9d14c8f842642e10fbd607dd0f723cab0ba052c6670ecb5c
zba9334e87792ef1464903d34bd261c17448f5074126f7c9af691644a389d48401107b91ef9d949
zd94e8e58bab52cbaf528d8dde522cf5b3a35d5adaf5356e5dfd276b077f3e59ebe437dfcef2474
z9b16dabf0a60354c0b57804d4e29b0f00b56690ab2d6081e1dd5796a7d605dcf5dba5310e6b636
z6819a0e0634369a74e3b291108238eecdfaa80f32ccd4c3bfffea866cafb0dd9d346fe47537cc4
z111027dab9a74abf3fa7ad32ca64a6dc00fc5f21869b14b0787d30dcdf2d01938ac538b67f989c
z6c5e9757f0616697ce1d348ba4a34103b1e9a3ef5b195b0f5744bf305ff05cb4fb0b3e66dd81e9
z608d83b7393a73e8c20761ac1eeab592eeb33e390fd524152a323c753a21743d782d74f23c9d70
zbcb024323177cace6e1df7bd97553a280b8762565631fdd437a249abeb2c2df4070d3ff62148c8
z70042ba18f852eeb12fb804a76357f3a73cb84dc24eaacfa15d2a1878f51eacf601d76ee28d167
z61ce41951a23054b352ea53624d81929f1f97622bf5976dab68b610317bf440b0744d99da57dda
ze348b9f53f7c4a23fcf2495b0f337faafac850a0a68500cba05e09b67d81655ac924474b4b5da1
z62fee82bd8119270e3d657086130bc7e7bf0f7253da7035d6ae4e04a8d50f2fef3621b4613b962
zc59e2eb52035a0af147b3f7dd886e0f80073141fe50ee360e425f1986b377124eb09c81968621c
z390277b3f56b86163c84f45a6ce72f77520326b2ceb614386fe53bbabbe98142d23ef107aecfc8
z661744f8919096ce70afa229919264f034b50b5520ae9d660c240f5c47bf7dfbb5a9c31f8c2a8f
zcf626400e91c1117227d3e293364d102bd74518f820c483b90d730c80a35c59531510628341739
zcb90914ae8675e2458820059f0cefccb33e65dfebbb51565f01652a55df201a5bfac3577dd1d83
z53c180b84ef1c114f081e5c79e109f1c50b2b88ecb6dc773fc4b10470d43e79b3fdc091de0e979
z4ae33ecb9b084e3e0b02bec22cdfd2c047198bfab7733d870a57049cf92b8631433901718f8d49
z9e4e83962726639c1e0e3b02ac48de06e759cff233751846ce667fb0f4a3083895fc80d0a7649a
zd4ccb4336ae34cd0089934f08b10ca1cc6bce273bff8d483808c7609d77b829d4cf21cd2a3092c
z688a68a1a563aa93ab46db1896278ee76c1348a594b89b7398296f2f2166b0f3ea9d4cb5cfe7b3
z8c1a8803a78df40426d43bd05516f7a4077260347d879a8534e79d995ed50e1505894908b7db6c
z1fe7b052a2a8e3d4041e6a192e7b840838670d1738bba6b6f18125b50e08ff432531fab04f5385
z788aeda227d6e541979c3ccc8ed48813539e4cae19ad891e50461118884d500cf649190ad8aa19
ze079362754dc6aad82fbafcb86a2b57534c74272817f2da82047dfd37313c920525be5b45402a0
zd4108e3f43e311b64ebc81cc0456dbac258eb60f727de3b9ef0112f80e6ef44caed95b1c865663
z1603bcfe56779ac4aade37c92fb629a2ce2cecf6a6b46f26fffd2f5594fa9c0e31e5ca6154a4b1
z264f942f255b43cd760b8bac81505b50eef223d58a7912d3567caf6d8da720df0b9c44e31b336b
z63946cb72d4db97e78c2f31ec064cbc7960d07cdb547c8285c4a3fc8aa9452117d6c55f5b67403
z9de699bf9e92b29bf4550b305e127b67c10b5d42723f0d961a113ac705078b3635092a5f3037ea
z9f09727e9d1c62b6b8826f6671c33c7eb84c3197634b8bf0d6762e2310cd83452e696b101b4553
zdd8db062ac20fa2f1afee3b2f638561f351474da6afe8fd0496c39a2571634386acfd59fff212b
z6a644d53d1b2055c863270b1c677a3d32fb132dc3b1c6ab2fda8442fecec0a71431fab28954369
zca377967b39732981e04b28e5337705694565349132eeedbfcf466f4790e65b20b6bc411fe724a
z9e2d1d5d771f5854c7672021a1bcfeb2e7ab23b5228f41d1b17994f1ed54178c77171fe75eccaa
zf636b9e9b83d81d2776691a569d31f49c4667420c9c6059ece1283deb753cc8e35b63bca969e60
z35f4362271934ec2ebfcbae9588010bbc2e799438cb161226159d217e19ea7a8101fc2a1f3ae29
z71aff45ba026134cd8ee9bfb3df00e23e3a568e68941a601d383967008160cca619f2a433a2b56
z358bddda5b51efcbb3ec306aff4f3cd943319c9bb099c361c283f24b45172ade54486050581bdf
z05007ce6ac6a77903118bda9a1d4b98b29c0a8c6fee6050dad1e92a07dc853469b2a7f80f1afef
zb516d7ba984e65cd272ec772de0287cfed8d6e2e8e920ad762e2e625e67e740462ec16a377baae
z27b5281e92a14e7a8fe5aa4ecaff160dda5323ec182c32360ee9789e0f65c15c89d6f487ef1a72
zdfce1f58edad49e61004286997c3981331148ea8231aa5da4f1b8bea15af1a8c9d67cf155b33b4
zdd5c90e906a47048d1265c228be2ecaaca5026100eb813bf642943a3b7cb14ab6b59a6fe52a73a
z80cd6765c42b26d608af470535c60357b41d6a2db98f267cf0106e6da1cdee00294aecf5b793e5
z5926e2b994917985458bc49fa73a46c1caf427807bb3410282758fe39c985f57723250496c9692
z9c62490cad138772d0a150971751b43df9adf619bf13293e6e4acb12f41cb1b3398c2b0c5d2104
z423d0d237cbc05b4805b4fbfd9952fef8ea10cbcbeefeeaa5fd5cc492527dfad68e54026181219
z8fe914938170296589875a2ecaff4f10b7c28398d3c0af900bdcd1e63d2adbcd1f4b9ba153a3f0
zd734b94c818224bef31131bebc90f23d40c993e8e6ffe2ab11296d9202188d959b57f2c33aa52f
z35c499cb8d114b674749ab46494925a5e3b258584ff736db55348c90b8e8da61bec802274cb0ba
ze7cbb94e8ec49e570c611c17f2b5361f4b9cb2e36ca954f0f7772c8f5779009db29fd83cbde3eb
z6210dadec3b22692de3048b09b4b9a832f7588ebd9bc4b14eecbe543113c0272ec35db6696ee91
z73cfc428b4f9ac53de301107f27e7356aa1466fd3bab5ad55b83d11741636461d520623ee14f95
z1bf007c78f0eea6dd53dff09befd22e636b33358faee5bc59ef7954483d0c8f0be6c3b3e3c4feb
zbd66be1eda2c2056cb9aa6d0f5712f7fe10eb86c62747ea7ae37773ce236be26edc93a1ef23d3a
z69bd7aad8142b5771e02cf447162a1551c634a2380d459a62509ed716a27e78316286eb13f6f46
z474d862ff093717d06b2467565e0d343e2ed2ced7c837867b71a8710d7c49325f2d350aef81aed
z4c7614a492a91bfdd2a6f8310e55a46ac8ccf04a4c7f68c38eedf3e4509bbc3e06bfda91fce004
z1968b27a7a4d8691d5e2978927d6cf3686923d1168f3497b515aafc4a64d69f056ee59966db591
z058fed5b1cb748f20bf94e9e606ec773aaa42569e5ff18c3dda3d7cbf4dcc2602a238b0ad32179
z16afe3bccc78ea8a8f2a58d949a3ab08917944115d580e0966126201046af862278f5c92f52d71
z9b4ece98b125be9de589979f962659f2e0acead9b63e6a0a3b74096c42b3c8ec10272c3f11b2c3
z262c9f762630f4bd8135bd317b17b9e7e0f14074886de2e133ae9595b1adacd23b17a4bd80d5b2
za0032027c04025bcbbc5759d406d0659bc8e99ae45d2739b4281f370d2b276b8056b1dc6aed588
z9c6d8efdd73cb819587f83e64c2284852fe185969c901d19ed6378e01a055842015e84ff2d6232
z72b42c74be06404ba86646549c2395fb22947dac7f23bc55082bad660195399381b45e847b8b47
zff88c0dfbcdfb5088dd162de1d1127ffa26590659c999129683ebf2bb642751a4ea49471b5e9cd
ze3dfd5e150da72baaa20f40122078a9fbefaf1dd8f27ec54a8a17511940fe2bfe5f885bd967afa
z4284c85b1673b2963945d20587811e56e97d288f8e287a7f5ca9e06e3340e6fcbe4601499c5aff
zfc6eaf6e0c0b1d874ee1b7bd194e132e5c005c45d4d0261f1fe78bfc8c7cf8eea3d17fc598af2e
z60a33214412d32386e5a043249a00a230be8a1138726bad14a979636783da9ff9ab9e4ba73fdef
z152ced966069a58be413eafcd4d51bc070f4bb22426b282bdb4aa1036f0fb318a945f23db36dfa
z3edd7607fb3d2fce5107b39c3fb8df90196b24fc50e13304118328f3d49f336da35d489b2879ac
zcee60cacdbe16ed14d0407ccc2dcfce5b46b5009ff77fcda48d3c2c2fe0b73cab31ba383998d45
z78cbeeed8788a00c5fd70713ae9177db28964dcee38a25f225a22514b0ea958d7eb0dfaeb29dee
z326528122247b82a833b1da158df5724c9fd217675eeeab9d2ca2e6017fc4f3fbe1c618ba830b3
z10dcda33746a82357701f682ca2e4e0d5e01a1e5e6903abd9663d12d288a64d6572f5bb609eb81
zc4cf41c95a758f218f019e241607d72cafd27ddf9edfb126d22ee49162553a77c7fddb6c3430d2
z076d58022e0582bf974fc36d7a6a295e2ea80a0b26674028ef48edceb898cfe7cdef70fc225e2c
z217bddf79ee950fc5a28a08971b07485f4d4d2d358644ae21f72fcb3bc078815bb7daba7774abf
z4e2ef22e0154e85e6a97090344442adefc54e36ae042d11d75b9184fdbed20b0d8c4e9a529a0f0
zb3d368eb44b51ccc2949518ed08a12ec13d277d64b975245e6a563c0bed05dcc4f6160e2959f4d
zbeab56a948c3f3551ef87985a04b38fdc50381b071651e943ac60b0bef0e453edb38abfd016ace
z2ad0ed0376062d488b33e05925ebc357210d3115be2459bcc10ad7cbb1421744978a01f027b28f
z9d0e2898802c9bbc39f1525c7fd802400668586e1546c900a88c81a6f4ce38a16ae894dd72aff0
z98555c2dd8bb0bf1669b83891f2a6dfc075c3b746f4540815acf5ad757a82be672b126e18a61d3
z07a9fb9e0dc96f150f1442a01611f79c879e7d8ede630dbaa6e801b761f32f69c640086d76bef2
z399b3c1c846a127397fcbf7adaf75e0f06b820b82e67cc4a65c9ceb6ad900d99016ca327c674db
z57de81828bd1929173d8de95249edc3b43b70e9b177120cccf07502d9cee214ec1b0ae11bf83b9
z6625fc01a5d1933ed55c6c5d51bc71d9102b454dfc50bb959f7d607ebf3ba1947215b4cdc74df2
z16bb26a68e77bb9eb00c90aa37c261d043971235f819930a5e473f6dec1bbad8774f931f82913d
zc23b1a9f07f5da6b70bb56b76788eea1282c6c4cd6782133bfb234e9a5e6630a078b81186d7c69
z9f145a9a9ffbbe2d1848506c3013cdc2ce157697fb935c02c12f01eee66dd2147d79306293d8f4
z031773133aa4fd332933b57338de9aa2d79afed32a29e655d039f90945b783e405c37604586af1
z3829a1de4036c7854a41f9c0ae608809f52e52d918e26d7552ca398f435269ca20f4254d78f08d
z40715aca72fc571197f6c3cb187eaa8a087c93d16d4c024ae9ccdccd3514cd5b26c2085f5f7b26
ze86227d4bf66e93ba26b6ce6ca8d38a6d8cb9070a8eaaf8dc726ce24286eaff9183a7d5c81b981
zb5532c2940fbb666614ddf6ae3ebfced262c0d0ee97918693b946939227eed9e18d6b073cc8688
zc7ec1c7a6a04c0ac554d83fc63ca544daefb8939853bd3c84508440a8686f5c02e55cd177c5a27
zd5536b342dd7de0e1a8930281b18544a32976be24eb871d6fc0e16558fd81273e8d1358fb798d4
zd3fd492a682a4fe105759c6ba4514e4cbf9e06e20294118daf2d82efad23df7f83f88f8abb86ae
z5382b4cd9e25a90eaeee9fd5b91318a5a84d8f72469f39abb540d60239bd977abb5c452c209235
z8ff9f7e65f1f7acd1c15f8fe24786a744ea9a596d71ffba7903489827087676ab87391f13de5b1
z212baac5436ca6fe11f4b83f6ecd83feadaeba300dc5e87a8441bbf0d3fac218191d48cc3771f2
z18e8845f5ac0942bf16a3cfc67f77829407f9932a8629de107fc1a1005cf4badb2564356ee70c2
z2d8f3a1f6e88ecf83e39788ad139a080159b7894d963743ed5c9b21f0114038e5c5c279edab89b
z61f10b1c89579d966aa5cd529b2f79f79f66bde50fae048f2b70901f1b6f82b53645aa372ca591
zdfb222bac291e5164e0faa56f60284b438c9ab7c4493073846feabe033330bfa9fbbcc1b3b68dd
zcc4b127b835e849f830e76961f9cbbbe5350f494b6af3bc84683063af0055488ea5f0d369734d8
z61440f20823358eff0c388054ac1271a9dfdd96483c7f2c4e838b696d19ba6dee87db4c404ccd1
zc08f5693807a716687c3182bb5321b19471995754393e327b1bed7633d5b47b346b229efabe44e
z954c96493592413e73fab6e552301aa5ad8d4885ab6bf5c6a0279365273c3d97684c9aa42d193f
z7cd618e0b72bffa432e66646138ce6b14fb966d19c02a0ff07652a03c35f4150744ee3f332920a
z2cb728b8c76bab4052b6e7fdc9af4009968e15fb6c6e18124dec3fd507555f6578eccac2c08357
z884996410ce8bb44e7de437af25958cd4d545643b56313e32938a12467ee916dd8f8f5047ba4d4
z57ee18680eddf5d78a9283a431bc35927a72c2ae6b5bc1ebf4b2308a72b34c8ac6ffcb3e9b8d0d
z87cbdc9dff11a58d389e6cc40b7147ab41bd40c310f243aa9ad587adcdf4d1a1afd9d04325925e
z7056a8c8bff1593829c9d0204edb059ec1c33bf310641f9d4057c569e381ef3d48fa03c4f4e9ef
zc363e9568f751a0e36cd726f057410767bdb47a357f9bb519e94557962de6cb92fa534c3faf544
z4007e96a2ee648fd367a8cbbf0f7545a00698ce5f2568436cc8a34622cc752832c286b8c9fe7f9
z0295ede2dfc3dc48976cae1fa0e6b4f1fdb2526a21b8f29025d7827ae401b5a41feae36008e582
z10f1444ac59e41b40f02236f594e983f46ac44aea8dcd469cd5b91eb44a360db1e8a9d93bba44b
z25f84ca9603e5238bdd1daa7c7778b24755a7a02ffab31e67a88b2d03ea1db743ae35517c94ddd
zd6400c0fd03ad6c84fe502e43c8d3e213fabfd8e28920e83f93adc6a0da3dc5752d1f8a94910bb
zc9bf02a09a68338a6542a0654034be5f1c88164ba0af636f9a684b2157172c3520985f86bdd246
z69b118e94eef746c93b921f83912bf7b39a39d65b5751811745b04fadaed9ffa80dc3b99214170
zc4099475697a41b4b8e947b19898f1342008f22eb3a66b816de82f5c121a4ebb05697e3c1dabe1
zbb90f10bf4069a91413d9226a076d91b98344774ef346f66f1d3c9b0a5ba9c0b1a7cb5702c60b4
zc3f9d7c76c306291a190dbcd20f8d1a5f0b505a355ec6178e8fe46d2f896bb5ded2e999639b996
zd4dc1545bea8722773ecbab3bcce7f7bae7a81e5dfe1e4ac9564040d4df7774038caa7d72c5c5c
z31cc29096117ca4645e03053c1ce0bd62ce9ab693de86ccd35b0dc1d2a673f1b5eb4263c73cdf3
z8c05b92ed43da6d3e993e4f876d7a8e97bd288cadb4395d6a18e616ae1e0125547d8a28cba09f0
z4f276142fdeef9ee76934db0f0be3bf83848bfabf3f9aac3857bdf64d9906af3bc8b81e3a39bc7
z79490537ff50075ecbfb037312e2f48888a4076ece78bae1ee148f675f6d9a8cbc510b1d8a3f84
zf7ada0f92ec59b9db8b5aba31ce5cdabb02b8bf1db803d56aaaca22db39dd775af99b01698dbb0
z547bb52e2b2b0e5968c97626949768d8d7854276544eae7906e449c1dbfcb82664f00ae432ad05
z6e1758b0733c77055806be556dc7b7d530a4b797c58579d9d98b119c66d56575f23f523c4c4b34
z0f3aa74bc1dcb9a3f5da4917579c157c82ac33f271fd418801ace4b0fc2c28e1d8eb7358ae28f7
z6b57f8acdcdf1e087e1c1a84c5fddd6e8c5a5d4354da0271710bc345a5486dde101c48131e4f1d
zadf86eaf951b0f2566dc786f4a854108a0ef582f069f1069c733b6ec4c4872f2b397a9d12d7c41
z8fad3f930e4353b99b753ad2487916fe5f0718b38ce46e11d92a22cf92f4d402955720fe77c3a9
zff9628f8a1b9b774d78be1d419a869b0442691516fb68e78ca5b4dc94d2716d4b21dd62f631d6e
z076c45ae725c65e535e9bd93b78c08d5b482a914452af0e1edb5fd24ed53c897f1d3ab12a35c4e
z84def95f8f12b8ffd6e1a8b982862a778ac75ecd91759c5f30b36f28f1c815e96888ca8f6760d2
z7fa1214f654b9849198e17ba3dbd0656a81a6a58e54d0aa7852d0018ef3014f48911a6e1941541
z5477084ccac74adeaba08e74bef268fdb963f45ad5438faf4c89368c85e247f221a5681efd9124
zf830beed61285a5850b778e8db1bfa682e8b41e1e7599c63424208f9cc0a5a4f03738d3b98afb1
zf0cc7359ef68be1fdb540ae58804903614307f258d6cc0361f162382f04e42bd5a1bf042e35aaf
z7c3d92aa63923d7f434f1d254796ec6dccfee98e3743ce6fd053034b616f7069ad4256964e67da
zbeaca0875b960f9a1170f54bd9651be9514c67eebe991863deac60a112bdaad92d8265f1a6caab
z2549153e51e33a7cd6675a4dbfffc49d4b68855c64331e49e74952d060e0aa4d1f11e579f116a8
z0bc5e679bed550237131417ef4d91c42b17868edf8f72d5206cba2305187648c13a294fd86bdff
z72ffdb9260924924ba948769b57cca13d7d20c16d25e869e61960b014fd3deb863b815caa8e0f5
z7055328dd3340b1efd31993ed71b3f01df3bfbb8f800570b8349e831b58472528541f6bc22568d
z7fe949182a7338b559bbcc0f870ee0537e87a476a7759ecab6b423a51f4c3be3e5d0d4a73603cc
za04f7eb89adced00e7b27edce8fcdb5bf60cbf9731f476cadce924737cdd8227a00bcaaf1ef273
z7d69cb8390ef267d4bc050dc1452e732b59f5f83124c136ac6190341b9b99460d6da4c8c1ccd0f
ze88c41bd8144053dcc2eb0605694fd9f788bfb01a711c7b8e2920a5325b4a84e4e889beac20578
z170804bf204f34a7642fc171e02ddfc6fc9be227924cd8a40e9cdf9e37dbaeed4a968ef7185bcf
zd8593a716635fca0f5817623ea8848ec0f7b3ab796706acebc0291f181155840325e625cd25bc4
za557ae729654d60980e809cf8bdd70e19fc5b8a512e69a9beeb02b7ede2b16716cb2b5d9bbe075
z4c05ace899ec63bc8769d7601c89fb2445a3408832102f335bffd3c1021ddc7b81f4510ccd4690
z9d9f23b9dfdbad3e38e068a11fdb96c7417687c6e9c558c2cb6d79f319fa790a69aa77ca4fccfb
zda9f7c6e6a450fad127af4c388e7cbbfe80fa0d06a0bd078eda622ce74008f9877ed3fbeaf963e
zf62a48bda0e40a3e610e8fe55e6cfbed06a4c335b5a00f6f2cc8a577056dec534b882af18259de
zf0edf102c8718e1aa4794fc7d02e74e62a223e4be34298d2160a5b7d22b23e9c20cf4b7c45ad9e
zcfdc251714501b2570cac3536702afa4614488fcc005ef94df28c1a1270032c1ebb633bcabfbf9
z8bfdfc9d623abeb0e506bd84a9e5ac543203b259d931ab9bbdfe33fcd81cc48c4af797c23b8196
z6c1dce6767972c637ed5166a53afc95c5c8187772fe5a2b680f5e7af5020e60bea28a754a5f17f
zb2e0e1b9d6322cc1bfe94443eac28ee11ebf8c2471307efd89deb5afdbc49c12e92f822ab4172f
z31ef08bb44fb7017f154ace40c7eb16f160d53f0e8125855b27030907bafc238b5f335c7b40521
z311405bb9bd5be1b8f8b4e83f84e04db6231626f1c7038dac68536656590c65422b338e218432b
zd9af394ec13da6cae989848adcc82583645e88dc6f32ba823a5f36b1a97eaab07034a9e63cc295
zb989d088666398b8b17ee2bb2577a663fa8a740dd52b436f7fc8635a12656e1d87633edb0117b5
z4d8a889fe438ea59c7a2a6b7308ccb4fefdd0c21fb928d9d4ffd7cf21d94275efb93820d1364c3
z88dba691b8c8d24287565fcc445f4e2cd8c24cdd5492ece1cea5a2932adcf206086cf90fb69f60
z073b84066e2a47f228bcfd62b0847602732faae09881c58f9c8f237fb2164ab3e4dbe31e4b0027
ze8b88a6bfacdcfe1329311142446fddd318fe93385770fad4e9cbc67fb4d39b489adcefb111f1a
z19a116b242b3b37590bce00a08fa5d1af2abf297e511c5e5b792a5413bba74aa556c9407b5c44d
zbdb20328f9834a4fd2d0697dbda914a5815a2ebe269ba60899edb23963db582a8d835167ead68d
z2053847c25e051420af6acd7fe756092c9239ca7210214cb90a316b24be39151d9681d4123a9e9
zfe7055ba29c563e66822f2af4534de60a20170c2ee5ee8c15a8cbbed66bd767ae06dc18c729af5
zc212e98db03e5c7f242ecb4180336c4889cfc2fae0d1fd6664e05dc8082e88d91e3a161ce20f11
zb3b9976ed5570edd81f9e5e180495cb664876a05e1623a873910fbdb2b876e4216787cce9a07e5
z38bdbbcc142146ef9caf3bf7d6865c8871d15fb431a407c63cb7af6437b8ef2281be382cb6f5ee
zca9a3e37cd6091ef090de2ca7a135dc053d30166f15e2d4157d4bb0128c2c8d2f703eceedb159e
z7c95fd26b475bbb76024c4e1c9e5cf775b18c66df2a37d5ed44a438c4c265cb7f4be2420a7380c
zd76999fc6faffa8dd82954572c7155dcb85ebb6d82a84602f2ac3d3295f653340c13658cfb222f
zb12f5b6bdc4855f8da4978ba7ff43d14cf20c473451124d4e9d170e75be439ef00e5fe6ed43e7c
z7ee77da55a54841a280feac480affd1b6cb3e9aa95e631bef13b3d54f222765b3a472e8c967d8d
z516c8f2e5cbf92d79d54185333012fba901477a2cecfacaeb06a92811922506a769cb1985fdab8
zf140e1706a46b97dce8ba19834a8c0775559f6d09e8d368a7097f11ea0fc167b1a9c34915f8f76
zcc4ce4a825408ee8a7692b25a808ff58d5c418792d3b890c155d10c7eedd4d9db2ad88325bfdda
z3f613af482a605c6ed59543c1e2c365acfa5e9740dc594163d598e3e24303493b22fb90eaa5f6a
z9e542145617224e9739e8aa5d9ef51f093a7a626d0bf7b846516a15804bb8281dfe4e4a474382e
z972ee8e43402c90e210f8e71a65bc1d0b14134c09bc2df144469015b217fec7bda209b0a3ea807
z87e8b55e0763c2d5ae7aca2972284a8e1367cd7da6bf8186beba7459318ac6296ab40e0fb4167d
zcf01e8df6cb5463d911cc83e99618a19c34064db804344a8a0ed0dd8be7515e534ac6baf32896d
z1f77b323884cfa1de21cec0e668f453f4c232591c3950d53716b25059cc15dde11205dd997eed4
zff60e8e0a7bc1a893d3156883e27e85997f613fbea5f6281d3c8be6f507345508f68752185c157
zfffa4c320f0ae2f4c0384201a2d07a48b23be529aa29a785aa94fddbcec87e0027f8574fe3a628
z3fac56dcacce8f61c78d32d132d8293d5a13adda0ff44382d10620670a7a5e85527d907122799b
z00c84847faef16715985cd74a6c96e5984a08515f4b7b010b8c1123bde1875db37209e00bc3ce0
z4803f76b6d1173e16cf0bd9fd215bd496f2a3dd91b1056e930d65ed62f746d51bd3b3e3a437d79
z767a4c8081c7bb79a4f99667d595d4fe1f4ec30cc191b6f7ff0e0f9cc9b8290709eea6b1167f3b
zfda65764a0d64b84dee32feb4c4d86f9c444b33d95f7dab8874d2bc70c6d784fe9b41fba0c403d
za8c80d93161a7db05635225a9ac209f66adb99118d8a46c62a7a6d12a0f6dd6e9e4e0ddda8a1e2
z9e906c8a10d8be3d7616fc899857341c25379994dd9752eec8392002eb619ce9153ce13670febf
z8a319c22a3c28e190f4e7b8f6278d0ac77c54ac496e49f3d35e1ca6c94939189e7dbbe8147749f
z7296284f75b914b2fbb685b021c39dc7af81cc9774198c4eaca1fc1620347e8e25c19bed5610f8
z271931d3859c584af31df2d550f99019037c436fef8d6355ff1d5be7027c02258f003742831140
z1bc7de20617f7d9b73c61b926b6b4886c3a752180c6a7785c3f24b8eb23fe903d9ee55660cec2d
z77703d524c3efbd9277d34a628d18bc4845db03466cda2770b1e745cd439a1b6b7328edff1f311
za48cb5f2abdbad7268971abdcb2dc24d9061799e7cab26668a9bdfdfa058ebb647d1c0194d2e35
z778785f27a4ce95d55d4752ff003a0da8e27603895c0bee6c2000240f9d8cc6840ebaa2283a419
z90425dc5dc06aaca8817164bd565ed06d3712e05808ba6423529c899762c4bc0116846d1dde320
z82271273742ca6aa8e2eaeeed4c069c2e05934450161360172cf6bf97b573a4e4b6d482519a553
z05c93f74fcc7838d5a203ef547f1d0d3df3acd2099cbd0ad7ec7a26ec40ef671a840bbc0755ac6
z638797278dabf46f2ed16142758fb0e1e2607bba3105d19f4f6da0ec142178fb1ea4f3bcce3f96
zb5cf08f5fc5530c62037c8bb65f9fbe008262bbe43250f3912fd5bf702e07aceb5cb7c214a6bc9
z2b5687fd411e129bd6d564ad683b6d292305f7d9d16e108c0ea535c692c6139686ec61cfd987bd
z4025175f743a04792b2c42bf66511c8183ce6a7940e9d2d0c011f318a3496251a472cac87aa3a3
z708e13f1e9c8484c0a5facfd70abd3df6b5861deb78d54721ca28de38397738b50739b8b4ec33d
z2ff16bfd15a92acea94bc1062e02788c088a27386abe715c5e072991c3c68906069a8518779609
z7f76b436de9cb24e7c267ac2af238efbb2cda930941abded9f805333b4e15c9e2cedf41104bde9
zb0877d75f1493efbdc10ea8678a1f48d786974744979dc3811d3acc1d2655aa55165a092147c8e
z3c47ce2f7886280c6433a63943c2f6db1609d4dfd8fa49997d81a2502859f0dd24b808931f3b90
z788faf07dc34048f9408346fd2e26c23913f1fc9ddcf15e92f490d3a37bc6a9c3131b57bb261e1
za5aee6cdab1295a00baef941de9a1df0ac75cd101425e9e90399027a08c78b5ad3ca6361cd902a
zc24ec850e3e9670a08b4aaf62db3a3bdbf18deebc1064a7686ac65e643df798134fe0059f37eb1
zc44d2093ea9f38fb0e0fa490ccf06074997cb544057ad728e477a80327be4a7776a702b4f800d0
zc3fdf5b986deb643a9a07971dcdefd931e6824429a1b74226442955408085280741be6dcfee2ff
za9ba67aa9eeedb8d90b2b770de013d4940fcede77d78b36e784d505f4fb5143dc00cd2f5c27916
z86004439274592f7458a60da1a70d449001c34628c0a0480ea64065d2bacd29ec49e2855050672
zaf45b13c4dbd5777d6bc6b3fa1adbbea1d4d4ba0ea369b5ec7ed1bbd21fb53f5243cd5a46cc0ce
z2772471c7d17d4ada5ee62fb0e2e0b562efb67274281b0b424c20c69cf1660302f20af0b447d82
z853269e08fce964faf2c8be9717c36db8a25fa569ad651c04634d6e4914d03ba2c52a1ff27136b
z3e5c315703f168cd80534d44161f66c51296f1e850066496abe06138d16d098187c90a3d2218ef
zbe4623a71a82995aae6d37465504c4571f8557d426187e3dbaaaa75f2abf2775f65c674c7b16e4
z3c0da5ad523debec9861191f38a2ba1d59d7108e388ad616b70cab1cf4e0ea197bb49a30135bae
zf9923f5248d89477346f97a2f73d5ec1408da0d4cc4e9643939c47b7a38d12fd8a691083b9fbac
z6e90575ae4ecd2b0da49ea6447442b9a9a85e9bfa5bd9053dbd35ea9e90f1989ead041dd571d4d
z34c95e17a25cea99ec9d3026c085af0c4945e88c1b41c8f4f3ba5050c18f29c2b6213c3cd080b5
zb0e0275364380e102fb9815f77de489bf135bd052657040034344f71e0444f2d8b9e2adf1637c9
ze2fc55fdf9015b97a258aa800ddefe19ff699f74ca7eb45378cae0615bcf99f8015b44fb3edf83
z5571cf68ad52f780fca3a5d9d242f2e62700235fe9ed169296e0e2d9c8f146e5422c6dedf9d1fb
zf15462794b7517e4a9dda01a56af775684466f4bfbd027dbc0e4887cf45e0fed5f9e684adbfeec
z4a5c9b179d753c57a9f51aff585dc2957dcbbeb1fa515c5e38470324e02c86fa6d62406913a08b
zef8439bc433382e561640707db6ea4a00922e1eafc588d19269db31dbf32ac090e77b008f63695
ze0d0657cf0e731f85564de8db0ae4cc2c42732214029f562d61eb69a939945a02a0dd8c1289f27
zfb0a515eb1683f4e22569e7a3227cdfb191951dd3c4535f3041dd23258ab8df057999cbfeead4e
zd5457ca93e678edea9bc3e575407961296e44ebef1fceb6aeaa9fce59b0d65a0b345db44796e60
z11dac10beedff237f73c4e5fc2af8bea613a5fe622f7dae62fb4657697aa100be6dffb72b0a0be
za11e73e1951072027f46fd543b0a07a4d892a1d6390e9270a753ef97beffa4aee9a5a3e8978973
z180465f0ed2b76b77ad040c9e41d3001bf3f85ea92a47063cc437393224811a844ef0674d98db3
zf6cd6c0b3a404d2b1bd4a820fb2ca71bb83a8137788175ad5de0354d92f534e8bb02a4b300f098
z393f9a6053cdee503c128cd6e1ee57a2949cbe63c5c5fc129d75f0db350836908caeb7058678fd
z41b596c55bf8f352d9cc0c7aa240344a85d7d150fc4bba56a5d8d82e53c2a65763e5877bd204f9
z3ef9890927e07467ff45cd89081bc22fd42fbebe641a29eebde4287ae46fc6bd91f9e31e172b4b
z4c09ca92b641e277524dc1d237b6e8df32cd06549e9e833f2d6a616b80aeccf282a5070014e1fd
zea74b52619c5441e88243dc956ca0acef388075bdec3e8de1a14aed3da64f2c6161f7af6f7b41e
z421a8fcdf83dd9d306c5d67b36ac7aa329e14f7b42366fb841bc376ff3bf78b7b8db19d750f1ed
z8bc8ee5132c2921df6c3d968eb3557c7ddb7bdf61d876e1bc52893335d8f5fac4bbb7c48fbb7af
z0774d7f2700d1a605d90333c9ea45e213547588983dc343eb667b87e1266397cf1364b4fd05a54
z22eaa674c0b0f6685826cc6780532ec678d0de5aa6923ab82faa0c9cc1d378f4d2d45f82e357fd
zbb7915d1512d549e9b7f9e66e250a3bf05c2cc599a7b05fcbad54952cacd1e9c8a4ebfb7bbc4ad
zd38ee0b22b2709b312b86297cfa06f0094da6305e059286024dbc7fbc8c12a8228f6d1249269f7
z7174be1c56dcd7a5dead48278f8b91852cce28853fd891f9df01794c5a4a81934510af4d4b5d68
z046d94483cbdcf5adce418a57ac61455e4bffe7a79a75b611878ec4eb73a0e7ee7f7b0dea218b1
zc7ff687fd92d8d1c5b1cc6f9294d4c6807a5debaffdea741c1534cd427c1eecb5085cdaa53156b
zaa4bc9965a18b7603868cd4adb34cde52e102e29275af15f25c373f36bc329a50c2ba6a74c95fb
zf18b8dece7cb622ccee0f21838d74c144c585110879657d12c016e62dc0261119775993c55ff04
zf22587e1eada5bed3ed9744f676aca2f9c4201dc8fd849bdc95f6bbff69a0ee93afb9e0770379a
z82b5b8902a2f8a4ca4f4b6843a4069287ec3c7ed3189b0b77bc2d939cf89a2562d452c17836c0b
zf4224cbb4a38e2f73f84be1a2a52bb7260f7d6bfccc1acc0cf8c88fa8b5dd6d5a71b51ab4d07cc
z4376cdea110945fa8564a7f9ca36d7acf031297ddbb6c280bc44f9e131b49e635c12f229e84647
z15a12798559d8f48af202514dc5f04c484b50d1d0f927321a33ccfa3dad38901664f003943cf4c
z744588658fc3d9b677f9f64809893e8fc4dbdf7d25156a27ea791e8e119c47ddb994f673d1adad
z04c421beec86e749f9e32cafdc19de0575c00165765fcc2eddcda4bf3d968d3f99d31ab5cadf78
zdfec67cb4336dcef22cfd8e1427f2e947cf4b64e6200af11978d832465906a500454cea86876ff
z1b4eb7bf6bec7702f949933f53a28e7b787907112cb83312a3e5d4dd6607f8c18d22a2d4b7cb2c
zd8b5a04be7fb3c947afee160960b33666840fb58fe28a93239c59b7cf21b6e74cddbd5508dabee
za2f6853aa7be9d4b94d8ad706907cfba1796485b9997e5526606e6d5817eed84a803dd5634b7dc
zeaa968d5a0df7b837796db07474d39f6e999c75c132d4b3bfb777bf024fae6295812cdf039775e
zdeceab1ae2c62b69a70bb89464cc364f6bde913fd95d8cbf7d64394c3a3a1f67502096b81dea59
z84f76aef34d77741600f1a1feaddf2680eace7bf23e54aa7d5a121c86d02fba879f1469c9545db
z96158fbcf9ba83c47fd3f50bf98dfaf44b4a64ce6eea9be9ebe0fd304c62b2a190caa2241a2360
z266025d3c48c4bd323997d91e310adadee639cde301da298e1fcf8cf745469bb68b3bf4f31802a
z53b9602337cc3fba3d8e8470635591dcb1763683389be769a1ecff8c6b8c5572701c51b4e9fef3
zf064704fd7099b21792a66003900e32b24217ef2beab08770a9b358d0f4926f9501dd4a659ebdd
z2e117978f905dd2f238ac0451d1233802af77dadb8656b2e45a7ae9f3cc4589a1983745c6490e1
zbf3f7c98ab30df2f6539aff48b3397d15dff00c31363541905c1d54cf1576ea7c3475c4b5e53a8
zf4bcac7c2c663ee8dbeffc51ff7ceda54e7b1a87be9a69c96d92dd27f884ddff6642ff38955bb3
ze7887764b66bc198773533d59de4a574a76b4415a04ee6cc8e48e9eef1320977c97939b4a4ecd1
za857978644a674a94870ae0ba359b86404e26832f5a1f774f2b6ae10e0eb8fe3baf0ce033339c5
z71523f92f58533b6eb07c172844bc79d1bb2aa6fb54c77623104e77c05b6de2477a79a5640afd4
zc53c57e8314fa9c629f2d4c937809f021c25e2280d12f902b13fe859bd4921193bf8105aab9c12
z721a9ea29e9bcb179773bc9424b6ca06bdb35586edfb7359ed875052105b6391a9654e709b6dbf
z9a741f7338d2f4059cf7fe92c93baaa935c971a2792a5a79f0f3fc5a533e22d21631a72b1cc45a
zf8885cf45d642ea2a2429fb6360c77e7a4c6c0dc1eeaa7934da6dc9156e441c60b6bd01f129201
z5f018a341bcf040bd3c907f6ac99b3f1c59fc3966c778ed94534f9113bc5b94dd56559f933efd8
z52eb17b264fec7dd8c5534f1dcc5c68f597a69acf46de0f8246bc40793b87484c2868c705bd1e1
z41cd0271417d4f3fc4891f090d38b88e234ab8ffa4b400557b447a417dc5c39fb028ed9b3b92cf
z01be67910567573fae3bca9554d0c04246249c87acc94c27a7872c31ae110008baf30cb0bc0c0f
z478a8bd8286cfd71aac5d4f7a1c7b70baa4a83d5ac1daf70eeb98db2e9810cecc0f22fb1314880
z4113a31e09bdce6d6438af97531d02db34c19b299d43d07e4e174926c66f1f882d1ee1f81ea7d4
z663917b98a8ec16a43cea52bf72ffec8731e064c1039fa92034273ab5df5b0e0e71412b0f7ca62
zff3ce483f116e2d0bdade46301274e31af1c61d2bf0d9847f2bb8cba9d55706a5f4338aac31101
zdadcfa338343137c9866053731c35d9b1824094432f7700b24e3763238501afa226a4fe668c499
z2513c706881036f5bf4ca1e26c7bb5fcf75c1b2fc33fc86d3f96dc7763a4fda4b6eec295673de8
z40b35580f2bb958fd59f1fcfb3c9582eaf1045bf6e18d19d34044fbe78c3731ff09d98e8e4962a
zbfc422b4034a6622f2d456386266c28b2dc8dfae9df5d19b86eeb0e5ecda384bd5555c659df529
z103b1080e966dc271409bbf4fc32a23c0036e7208130d1a4d09f330538098fbe58678431075fcb
zc2596dd66f5fdd8940442c741ee3b950d5c8caaaad39f8fb331ec16dc5f9181ff491f8cd31ce93
z5bff7352075be07f0f174a5c4d9a6eba6b8b1de5c333280a172d5f615b9dc31b3de44eafa114ff
ze28898cfb9b51426134a5a23451e1fd98dd4280be6f8f9b0960f927633920343ee696b12e9e3e3
zc4eaba8d6bd089dba015e2863786216b2dcb5b5ec8bbbe98fda555e674f608b091aceb76edc60c
z4a5b9da63911f1909a2e07416d6cb1643686950357f7afb6acf3bfcc003b775ae4ea9ec54a82c8
za5f5e295774c567d36f1e5c4177b43bff2d2a3137a5f835d6dfc33677282a4ecfd4bd1b833b949
z805abaea7485d4f1fc32eba6399f17a4561e1410b5a90864de65572c284a53e9d35d65c8eacdee
z22aef6658606ea10ad38074edb477f768f1f49c11f342649ea0a04938330054281af9688f60b8f
ze8c5a56ff8b94a09e170206dbd86db0f758944a78269b385bb9b6965852665d03bae910941cae0
z8b113f71872899c11d48feb44d86e6629e3b014f4045375dd3ec6286b3e6f1fba65b399b8e3fae
zbddb8251aaf20f5f26575d6d4c2db974f27b0af8768f522c46c194529e57a6d937e86373c52b82
zd0c98311784e7012cc32a1ddc6300ecc12d2c4d4464d39d786ae91e2061c865982cd6ee672d6f4
zaa44d14d3e93c8629602f64365c9c7593069bf556317258d8a50d13ea91189780bb013734a713f
zba2ab9191305efc6bc173d6a06246c7a23aa33e636082a8b846dc4e40d8dcb9a0dbe40c10f2429
z776ed8962063f96ad7ec077525ef87a94bb359057bf9d6e0a01d9ea14a79bd6b398b172ac9b53a
zc08dc928c3fe4815e58f4f2ff90b1120838bf469b5bcf56d4862ecd0db14d495662ee915291517
z5ad347a7136ed469000d788268c63fee30c1a32d2d6a66f3fcbc3cdcd4868599c1e1bb55cf1b46
z4eff50dbd16d07ed809f78188f8b6a795417155f3d3667dd63d35fd25f339fd22e33fadfc0208e
z92a1c65f89477ca58624f5bfd87d5d695737559cb21a540663c8e0e6c08248ef87f916f7fdb118
z89fdeea4ec6820019f815bacf776399538152b9855972b333e6e27a419c108f5185225c93ba2d3
z581cd884b484247f64f18bb03df18637c66221ecfc5dfb6999b59a86fa921247f31f3f8f8cfa7b
z223c6b8cfab503d976187905df075ba06a0cd5bdbd865cc6a57af49be14ec740f23103d1c422dd
z32d0e3f4a31da0c9bde350675183f7bf54b7df865e59af2c3c1c48288799a556b00f92a0484338
z29e71409cffb4eed42e3f7710fb78b7e6aca3fa0ae2a0fc0d1c5010256f70711bbddcae424b034
z19d306130aca6d9e88cd7443353641b7025b41b9a6d478a12c7dc44e3e1db1616fec4e1d881dd8
z91e06d2deaac9872214b277072bd1bfad8f760320c3f4caa9d58693b4db11fd8b77b47708a14d3
z1c55b4ab6ea6c05641b830b327d6cc87e26a023bfc5a76d9744d3f4dbfdd3420ca559aa446c649
z4a81526f8496dcc19f0dc92692f5258e7f86698690031b91ea8ed18041ef79043ee35ebb49a6fa
z7171c05a25187b9089170a68e66fa25db0fd1b5ccca27cc808f205b8dffd456841990608069a14
z8ea411769f072029161a198ccd815d9e4f07ece8fc7ad5d86487b674e62fae5c9d40b75798a782
zdb05c500571eb46b2a6a1b975ba39f15a7b9a1d808d5253d617f6b36f66903f89c13954c37a9bd
z877add3d3b352f0da59738f4872c24ab13a072262284f15d88b29e4ec264d5d3aa590df265a915
zb68324e833eae07477b13897f35fdc71c42d385d0db6bc9efdaeb7f5874234b163e348c9b3e013
z033114b06ed914fff436781ca36bd19c2bb376fc084221072925eb4d70d6468d3b4df85709b8d9
z0957e9498215844ed33bab88a045708154578fde599c01a85de634a9b2a7770195e7b1061cc51a
z3891b7d5849f07d05dbd8c58f27525846f8f1f0e1affa55cb2e24f9add466ad02215d286bf2ca0
zcd754ede3b770864d5b6548c37471885bac055b3b427c81abf5144dc8c83a1e9ce9b65b457ee07
z1b47a39e466407cadb7fb2f24e9f4d1752b4b5ce46ec0ccb8438c907e83664ff48a1109e800941
zfddf95ecd9fc2d6475a67e727da201327542fc974b08a5a24354291473ea2128ada173926066fd
zca24898e75d4ec8c9bfab042bf2547eeb45bbcb4808928f8828537aa6ee1e95f89f61a3f6f0bd7
z7f1c29cc19a64ac277cf43783019fdfe274006648b9442070389cbf5fc2e4cb4f696c62df2fa84
z303b397d29e70d96425617c47b3f8a7f4b110c41eb0d8cfbd6981789b761934a6907789921f040
zff9bd63e3cb2ad8e844f109884694642dfe9c404930c2101af9da12856cd32132fdf6efa468b89
ze065913f678d2a43cb68be80d393ed7f8a6f68422c93632f263e0dd9d73a6ad13257220246121c
zc4e4da2877f2b64fded8f9b3f7684fffde14bcbcf8550d4251dbf7966966caf48df09d1a590280
z47e7ba52ea600c2e78673ec5893bad7e623d8bee282f2c8403f576d6c684a659b1db97833d43dd
zea1979bc73206ccad0d04790b124ca99e394860122018c70215f089851b031bee9535b459be97b
z42df06239a8e56caec138f41e128092f596d2bbd3de66467df64d94a3fea0d4efbe28d56fafc64
zbc73e3b9f1faa2288a420ab9e137db43bcc8484d4d14ffc5cb7afe66462d60213fc573756b4d17
zd8dd7c7dd7e9d139e317cfe019db3bdc99aee77274bea96a43c7ed439c93806437901ec84ac2f8
z7c0642d68713cabdbfa8ab37c82f54b41d6a4f89b416450ff76bc50baa9b726963821026d936d4
zfd4559e9b42d109ba2a607f3fdd4a1bd3eee2cf28883dd77147903b238f422a2f86efc0e5118fe
z6e84815c30d40214308ff46137d76e9923dc9b10b9bbae155719d1da944c2f0e192589af5fd28b
z1ec71ac49cc93cf0fa6374db4bf0f32bc343427f7562a0542214023b10a1709d8dbdf8fa3242b3
z6982af4e4252d0f84360eee5653462ffbab8d2f20a30c5ab10ac38ed59a728040381301c2acbf9
z413053e6dc31bb7b32e13f1cdb24e0ef7d4cd57d5b0a8936df2296b980321b6f973029ada7c00d
zf432254443b9b838f225eb96daee3aad4248ab5124513db9414cdee48e62a43e0ed246607d1a80
zf24d4456c1be25f996b72655acbbf294ad78b73bfab102fa3f6cd3e927029f71d1611c037b7601
z3a91a90ff7c5f06136248586e24408e7691170e2d6b6ec04e2484c4afc43ef92e1487ed1f0286e
zbdb19aeb4866c32db3a1403d5e47358d6990dc55e6e222aa384158907c78ff671ded125ee9a14d
z7a38c42143dae568e1f91643c6490fba72ae61fe022ca92c17a1bf9c51a2d90594ab618a2e74e7
z182deae6d732aa799f6f7a81ed09337b915b1f63b0eafe3632dad22a943ef346bc9735d0d470ed
zbfd513e3d1db12fd06471bd5eb99b7281a06f3eb282e6b896426b32c8144b7d97f57a45c8cf24a
z51f3dd0dc99298408b3ea4167ea268071f14e40407f19dda83b2f2313e871ef812390986197cd4
z8122bba0b1ca421099d8dc42d8f4b30c5b0f228e9bbf3a3d1ceec200cfaf7ba9a36f2d176b7a1b
z087de87968609b53a8ef45b15daf3c05c4ce3b878904e29e4531d494fefcf11c80e891f7d3c322
z3f825774d1ca4248c99d9c17944a6d23c7fb88e35caf784c4168855c1d46530d03f544771b403f
za31bb97a99867f04dcb7aa421bd7d3a2d3ddea21a11405e85298067924027f1afa24ea2a2d5092
z7de0526be695376723d71e820dea86ae00b81c197d7273ce8960ef7e5701fa9e0998dba7f948b5
z6ebf8e4a213d77b3b402d33382c9d36e5c71de39342f9df556697959526cbd24b8e448e3a8ebc5
z7abeb8d543610a007bdfab123c2940a58143d602629a77e2508c9dce03d6e1db87b88ce3f36271
zce296b05f7b788cc6486d01b0bf99f4c2051d995b73d647066d9d42e3a0a5dfa4df62884ed5800
z55537e47f72502490b8d7fbd03da6b0fc53b4a346bc9fb38bdb577f9d7a77b5a93faef6828f618
z012020736467d253e8ffdb5284ec0182b4edd79d5bc9b8288acec2f2c4a5e8347c5541fcbd84dd
zc273a27f63fe4be557cff5be096e997760fc2038f7a1f603325e3f5cbfe9805e1f20fa7d8b450b
z3a3722e68612a7a53addbf3a36b2b34d427398b3440166239bbb9f6ff7dfd893cab8145321944e
zfa61faf9359c61b49dab68075bcb8a0a725523a1f0f4d7f2ba57b6c6305ff2f2ad013f8b92a8ad
z219519b01b43213b4581a81e6f7954d06017dd4555c9f802848a60970eb534a566e50b3db12d97
z874bf1131a74601069394f8bab156132c6b7a3c1d17ed8cf401647b095e9bf63a7b8d18aebd383
zbcfa66aa1179c6084171584dee3417e86a8ba280c360f6a8f04c7133ba78c60566086a1d82cf19
z2c2eaa5770e4e36a76e6bf60883fdc1ffd63399d331d1e753f801108ba77350a5ac316f37ca351
z26e2122a8a51ccaa25ccab9724670357b9a3c730e53c4dc352f207ae1d7d0c02fd323708214b48
z74509d0edb453d1c1dbb441b428e7f266aa0396bc59bc4063a54bb9fca79eda016674238744d93
za38dfdfd4b1dd68ab270d99067812f8015eb8d61be61d00bd58740f341ab341385b9fb44ba3a71
z966d5ea48de972833f835a1a4e588d20a0497e564889c1e534942b6a4b9a43fce3ac05f5e66d3f
z93f59434f1b27e3eb2630e88fa238015807fd6b564bc588fa24b3233880aab7d93ba9b341236e0
zb5adb0dd7a4c10e4c3244a98e6bf2073fb6f922f19ebd9d2d1bb467cb2c53a2017149058f2b5d4
zda6c7f80de438046ba69c023c76fdda4af4c14edef7a6003878185479e20910de72decbc7541cd
z40c2fdd7ec5829cda3b63ce1574041204d798cdbaec649d552ffbd8065a7bd975e399d97827c74
z63faddf8837044a811d8c545bfb21381c60918cf184d8785667e66d2bf2812319cdff83fed4e7e
z15fbb3a4afcd67fc98be627f691bfe529543221d6d2afb070d7a3f3e0a4c95cf58b736d167177a
zd37730e5e6b30ad5038a680817f3f0d396c21ca44d9a11b7b3b4f646f5d6c14ea27ba805c4d37c
z4503ea36e941e1eda90a69cf9e741fb90f2fc57a104edbb3a8eac97b3a8c80ab2c322ec96b3fa5
z53e29790b6c468b23ca3b7d7c0bd071b0bddb32815a7d0c2aea2207950dba980ad07b5caa12f4a
zf2ccb362088ad840afb5a1b5d689c827130701b753b343bb0190af397a9d7f65438e3404c3944e
zcc98e016d1de32806a87c41fa39427aaeaf2412778b8ffc8e0667ae83f26a7909056315b2a3944
z3e01cb80542c92168d8d3b7dc65f001a43df666851263729adcc028f1e5f1c2ad1eaf65476db75
z5a14ab783ec0d37931a22675d08265bd59a2cf34ad2c2e9a8d7ae3bb30b0f64d99d96a9d1b025e
zf6200112dfff101ad287d5b3c477640e14c885e57854f5af6f2da4d831f8bcd916f51147b99b27
z060c635d78fd1dcb95eb0faa65e2d113a06620600df8ba27ed8b2757d72d0a4c9dd8ae3bb0cca5
zeda2d2a21e71d9007307cf5c1f48c007521599e9787060c7a415186cdcbb79f4fa77c60f5e0b17
zab144e9719edee7eda93e1f1ccb2337bc04bb3c79d064f16c7131ef0d8804d04197cf7b5a75ff8
z5454bed95251ebd766cfe89f8e738e0a0f24e896a7691b306fb368b2ac3689f0fc4bc82637e606
zf2259ddb96f6905ee42d8f4d732280451982fc88324bbf2332d848809d9728b19b5d9b28cfdb25
z1d4d26e8c6f64fd0dd7ed1a09e7b318b6c8c02940d94da3253594fb1fcc250fe77f0e9c991af20
zcff0d91115664726f26302604e616150f6bf40a76ed3012598ab0951669509545075a976fe4d03
z48a753f5ab3942528eb29012f5b41d6fb282dc918c017dc07beb988962f38e31aa2c8b3eb416ec
zb2133007a53d454a0bc72364762e031fa820f5cdebe961021f67f8eeaeb7d2c4ae23217776e472
z0df32a885b5456c1b3d79c6fc4b5d7f4151c2262bb87c12ac847b2474e71a154e3fc48408cf0b5
ze4dbc8164d81bcc60ca1e626f748ecb116f119922d1a5e0c962c4d1efed332296f87d112555e79
z6f5fd69e2d18bc67f3c2a1750e83552a89a836e24469056cbdffb5dd867019b8381078831823d4
z52ab3986d42ea2053f5338e5a41b9d8d9037f75231a4a3e202f07ac7e5cdb3adc2e8ece707ee58
z70fed999bb4f1fd7c79821d445b48870347364a5f1e4694c694a8262d37a9e2d95e2afe5fe44c6
zf76f1b64a89bfa9af60783e5c77f6656c0a26ea32cbd5fdc0baf7819694379baade36c4eabdc74
z614a63c333b06849e5af704473c48ed8ef14fff5e1c75cd70b31bf680f0418128215a4cce282c0
z46751f4e6f51aae97a4e077afabd5027bb38383628bd725e50ac93952172f87fb963191a034310
z23a3c5742701dc5682db3bfd5cb2949a1e662c3ff4c6cb34a8c325a714de9fcbc6512af9256c93
zc47c4dd6723ea31b4866a7df66c29b6efe75d839aa1d77a5e2fe73b1960d0553d9d5d8eda1d0be
z4db593cfa4570a48693e64450f96406d9f0c72758684ed4f8ac0d1a615bdf2b38f8884e1901952
z71eb53fd0c1de72e769a89699c30baa9cd1157c860a95fd2e1956cc2db1418c28d99fba0086ee8
za9e237530ce046222ca46738f565d141d482991f4b678ea99c565ca832124434104d0e42624b57
ze8101ff6b445a8d67ec8cc744d32e70ad13d42df083ab315534d3a10e7fa28d03e7168e5d06205
zcb881374fd8c34a7a41b3c20f8a7df8fe120341d1c483fac437dec33fcdfc148056d6372afe7a4
z42a806d1e1e31aa842d62389a97a9b99a72edaa2156cbdb1746af2e3bac12355bcb6fd22741401
zdd1cae30345ac87a136663fa5777a1573fb36f4b06d39000081126aa1e908bfeb381f83f3e6b10
zf93cf9b2b913b2fa1824c497ba5c40043aaf558d58906a8aa7a7b3f1986a6a1c8a566c85a75566
z3a3d4d05af4c5c4ebc85aad2306bd71edb1036bfe29de8dd2846781221ad2685c79115db8f60db
zf3b25305f215eb3ffc543531abf7581c416ef41c571196d2b3c024324b2784cfc72414ed7c0a5f
z9899956521bdfb0c61e7fc8acfde0454712a4fc8adcb78a4d4201b75a4783bca6ecc2d10552708
zea8da6d2846bde6e9a3bfc9df5d64d1aa6c1054860693e16d6433b801051a93a001b9e61d8922c
z75f08710df57cd8e95c06b9c1d99df23436084d7c6ebfe0d4847735ab43274a5fb1c5a7f6da158
zd15a16b052b85074e94c3fdc99ec3c6139540837c529310bde64968e8ab3c5379d600fe5cdffd4
z764fb0361b33d02131cae186b1e7d8ab9d8853b7b77d5ba6022b7d1dd7fd846868ecc105a31532
z8c7356db2ddaa581e99d42558f111dbf888efe14392d6b91e34065a0d0ebd42c9528009f8ab30e
zb561ade7708867430326c9d2619e46913705d86e6a9606eef7a70c509dfa95df92cb001a2a8bc1
zb04ff0e9a6b1b75f237d89972a29f7017428c87b75abd05b0a27830d4203f41245fe825edc414a
zaeeae2f67b3125852ebc48d2c0d12e5a93b06013b9735e11f7e05f9b59f91094a6e522bf76d316
zb1e137a43b311f8c5d646bca458fddae82eae47a08633b5af46306b0c4af3b2e6a76e2b8f051c3
z61fe6204388bb3b716251564da6350c654f441a02f406e3621da93d3410b5a4d7461f7d0bc1c1a
z928575449e511305d11cf14960cad8deb7d737dd49f9c96ae93d63199ba696740627680af34664
zd05381e1199612b01e06c0944195806a211e8110dfaa9b53976b5d3b39a0e7756a001b167fa2ac
z15c190b9b3cb780fc6cb9f7e3611290dc3b2836093dd5366b7924105d26f563b46d22e507bfbfe
z9d34cf1748a386b268c1f1d685734983c77e0c01521ae23041f6dad49a2bc976bd5ca3283b03ed
zf626e3a27b6d4b5570b148fb14c98e93dce5215fba227685066569a50f6eb96eeccb665fb3df4e
z8614b22490e5551086a3068da18f3ce94b58f36230d1d596cc2e22dac6741e027befdf72193a5b
z2005234ca122b75bb8edef093f3a4d4daced06bc07d9e3f539f6f4c63d9752c76762f0285ea139
z2cae25b3036266ea5313389e7e22bff6da320aad03d755153aef7c1738ea21612b1e4407f0848f
z088ef8c14dbeea536d2dd481d9a3bc9e9ea19c0858ab6477acad7e71f4158db8d30226a903827b
zf8165039b73a2a53faef99fe2e9b21f0b9677c66b3993a02e22e18c2f3d55a5595a77276b45601
zbf8f20b439b0894623eda59779609cbe1cac54f1547e09cd6672402ae816191dadb27e5f2df853
zf3290f7a4166b07eee049aa18189dbddddad407d28200e594987c6d27eb198d520200e55e323a2
za368fa601b3eeaa087eca310c6fb8ce85d691554082eb9713cdd19d560547d33a2ef2d28489edf
z4c5049c3165154d0eb07c20e43ebc929de7e0634c813723e7a704bdd8393322f4bb5f06d24fcaf
z7ac21b8d07b73d878f0986d7d43e61ed35f043251264c4d71c2d305d220a9c3964fb9839b8689a
z9b5eb62315d560ae55702fe9b8c0cf8b7759286b6be3b23bbc1d41b839d959086509c544c98577
zdc6c7f9821e3425ffc3f58b95e775f960de52a8c4fbc74025c7a5097141a305449015caf4c39c9
z3dcac51934b6292c297b73a81b2517165f7b53c79577cd96fd797b9bc2b90b8f1daf86dda8ca74
z8d4f26eba5f35c4e4c45657a0c86d6d313b47021489626606be3196718f38e066715247ec74244
zc3dd161bded43bf00a32f928b87388b45c8e09d7ceab9bac8391f03129851bd03627e71bdfacb2
z161f9a13ad4c438bed2e7f8872dec5afca0e5b544c1f8ec22f8ae352c73b9e526bdbd7aea40390
ze88b90736d5c84b1b2f861b2f11a63d4b1f29aaf255e8a12dbcc6bc7616f8eb61eb94607762068
z43aec7aa133d2b9c61f980ed44a5e8002abdfe27d6236ed7ba6920a1d069e19e9ba98d4b54d8a0
z33009eeb665302f46bcf855838df31dbf78f66e318e733642ad5a5cec6e0968e5c4c69754d0f3a
zf97252b2f15ea11d29808f233a81cd3c5a3f42d11869bb19a57bc15148370b35e72844cc400a0c
z15b15a7cfe4c3d3a6ca0a777a85926f41efca892b46ebe4b8a451fa2c112ae04423c7a8a722af3
z0ec928e47e9615aed9f8733c060ce446fe45c4821f84c3a503ed56833daf5e30abe0bb7abc7e3d
z149f4e4fb1dd8d981e2bc67e0df93181aa8d5d33ebc2d3c54c439ffac7a2c30a875382d0a66c0d
z82b6571c79d1d3b2685127dd1100e3ee027764f22ba5cb2a8f3ae5ce8f68d337ba85c9060d95dd
z684adf0ff5db00a42c71752bd8e833b06d164be186a8e9798fb55b619a424495aced5b111f3811
zc2fd57f51c94012cfe85b5cc3d34884e05c213e12b0107c844be19bf9e7dea4f91534cf9419dc3
zb70314ad6e649d4e2f0fa984580700033f12c0b725ba8d4199fb706b6a422405d4190267e56a86
zfc661baacc8131505b118ed82364fe3950ef2aea3c870c7adde6360320101357c02f6b2bc931c4
z0df3f4f8e6af54973668540e5df8be6b1147ef2d5df60cea4129c86be6cf4568a2c4dbdf14380a
z8039ccb49af5138c00b3e25f0123514045850325bd7d304ef694a7d6bb1bf5eede83fca9f6a34c
zb1c20ab12e0ec8892ef3e9043a82acfa7b42e6dc2bb4b9e537b28cf68d7644d6d1d3b38b3ec62b
z0c632fdda961ce3e5813b1511ed77c64a071af7e3373f97a657a44367aad3717ba4df6b6e3e3ce
z6ff0e27e03cee1aa6060734f5b17a7a4f820f672af6662afbeec616f8826d4048da2d164bc5231
z1af65a46fa5b38f54627572ecdc60b790ebd697d04a22ba29acff5f79fbd92ed4e7e2c0fe6f9d4
zf3b20c8686d347dbc674c631bf64a1814133a11c7f37bde5853179908540f88a6f40d6e92aeae4
z8658d9495846745189aa6b007db83763bf5c0a8c85773ee859eac6919e09a9dbbb34b84f3929f1
z0e92617a76aadc5c88585cd5f3858f015f78ea0ce9f007ee3c1a2e04c7d18772af700db2cfa845
z0942c1ad598cf840c872c669e7b52ccad1bd84377e72a1df991bd319bcf2b23360e10ce3111f2d
z260fe3b9ce87b48e4fca28723c5d055afecaf7e58583b6c76222e5ed7d1f5856e8826a1b003623
za602c156ba4552c2a944afab3e9d31b9ee1b5f7925201268f97d1d1a6a0138dd5d85a591a1b0fc
z3e1e5f8a9c1c874cc5f0563cbc1b4694e601f623c02850605cd1f2643af600f58d557cd9c5d350
z3b545ba43386e6b0493b2593fe288f62d2ad01d4d47c9af20361e83b096575341b4a0f4bb401de
z005990387d7234a4100f16d91aa37ee5895d57edfabd909f370102dbcd2322959232a1366d23bf
zce57213a5576ea927362b1a110e67828b6171237010508f24fe0290471513c994302d7a73b14e8
ze70bef20fb89c84949ee9c9b90cbaef012be017144893536512e2d161e142649e74d8e6bdf4777
z48113e1da120aea3b1c5e3b1633a0f43c7ed220030644c617149ee8c73471cdbe34902103cd861
z2b3a0d9c686aea997a652998d6ce142aef9bc8678a20966458f920fadc8a8582e77ee2f78b8496
zd20b18d23956692a8bff90c74b685ae6e8db11d806d7005e633b3233ef5c2f8e911b315a7265ca
z74f0058b36b085fed2c5cd24b82813915aa3c38350e8e0e18f87b7dc98eff710c082e5f9e51120
zeff65c82b3a23a73035e529b622d98e12ea9ae201d88166808639fc1c3591a0f218858883c98bc
za5d0355ef760757ae7e8366a31d9182897b838b6660e1cc629316c983c48cd1dc33cc0be681e37
zba74134b732abf8556de5d80f8e50f55e40a0dc84c1a1cac209101cc771c1cf0f9d509de350a7e
zf8420e037fa0502ac5beaba85a42583e4a059732a275d20364ebc0562e4401b20cde0f27055882
z8568ccc42f9da8b96390dd92b14a735a71cb980995eafd6e9932728957a607df74896bbbfbcee7
z1403a6b75bc182687b38bd68911bae94aca7d452f259d0ad1dd023e0d001e395e786a476c4d359
zbbf72ac5da9046313e3194d9ac75942cbe303d9c23624047d3b0bc95b5612ae82ea82c34af2cfc
zf255fabad5f1bb435a7ee075f7b0888d1741a7b40131f810fd3fc859a1bb34ca399b8dbda041c4
zb7b70a6a479f8e74373b6ed82248eb514ac7811c0d3bf41b024f2abcf3e6e7e5e1dce27f796988
zeccf0d4ba92184388d6d4b23cad0d597dc282380d74ddd2781dff4c67ed6315b5c8b8bdc5f5885
z04f32022e81b94199cc071e2c1ef01444d139fb1231c58a4870c256c033ea504bfbe5e67241837
zf83f6db240ac0971bce279bf65d1ce6c335180eb6def1ddd2bc32accce17963a5317c53eacbe15
z43564c04491de7210413f93f462647ae5b2fe3139bc0d9df813e9a6d55e8f9804f1fa2023c994f
zea359b2273d2c101d70d6327a1d528b2257454e5f5d7c0336d3bb3016aeb29073322274a437695
z1c8f27ee6d1e4daa898a32d7161cb342f2f6794d5169ca6383ca9993fca44db370dda879c0a98d
z538411d278430116734c3affa08f44b77febe014cd04f96955510b221648a0262caf2934c22bad
z661cbc43bbee1ce7b438ceafeba0d27effbaefd6e74be82fcf192bc12d3ddd741036feb4575bb0
zd55ab7aa999cb8a1706116853142fcc3e16b9fe01f6575b10a22229107356e25e5a722c6568abc
z2f60d36f83ffee669d7ac35b99e4c7477a663fd00819bc1b71ffa704e7f76cf82f647396027679
z1a2cf817911a3b35972f02ec2d120bb2e40996e6b839468a62fe2a809bd7e382b80900cfc3f927
zc927645aada12641fa0aedfbfb4a465ecfaec99916cc57b381afd7b68c620604719d3b97652926
z12a99cce2b3159129456cdec6a0af2017979960234f2544527a1b1585b707ea96758d613ec3f36
zcf5f2ca0d9a839b24634af0e8d35de86610b00e8d4f04be6cf8d4171e1735faa5bc4e9b9df98e6
zac62244b72119dbc469f828b5df82bc9ca8fb46a25b3c7361efad904ab5f1041be480601e2c2c1
z03a5b1b1e372ad25d0365f21500d1623455aace5ee39e28a34ee41789572ac4b6c22c8038d55f5
zb7efe627cd4e2d14878bdac65df28669c922c0b4415f26c616be49545fea412160f2872c2fd03c
z10fe1b7fcead8835e27c4e41052936fc33ff1cc6def9eb3bac76159086c36029eea281041911aa
z5ebab5a1d066df4a9925a49f42dc8aaf73ebe4dd3f6e10ddfdd1f3b9fbf5a4482e1e7a00c0a97d
zbd2fc48a192f8164ffe3f81d3c9c4d58e5f6b5c2cb4ae160e036a1e23fb5b0ea7e850b9bbff8ca
z64b20352fc0323de3cf097a6971cc68d825931361c306f660ff3e7bf3a295408b3c99a19f8140d
zbeabe646f80443681373d7c8202bc29f21113540ef07644597d54227b503f9294270c68bc8a326
z056be262aa1e286ced85dcb5825cbd519f0b3a1b509f205767036681d6b6b5c5e9e455f2794a92
z2099f3e548d80c745c31bf0eedd2b14b2098f94818c9ac216816b9b5bb151b0dd29ef102c451b3
z4584f600db551bc391904bf0f333a97f26232d8f7615496790ff8c3b8ae6beefaf010d41853a6b
z07e11847238e993ccc8fcf4cccdc3c347693d613c34c40de12327843eb931f0f041198c4629904
z4f7ff24ae60aad62037fd963840796b6250f675bd5e3debc58bb66fd0a6c461158d9d806de5329
z598101c44810cd10a4ccac0a2560f70e0a98e281d4a307b913e22bbe002cc907d7352750a5bffa
z7a25e59060d34c843fb9c7ae27ad4f55a9f72a35a2219210b2bf7b2d10dbd850d549f7ff0783ec
z0ab8a45d1b9d56076e886554067af5791461d84fc9aa2e2ac0f963856feaff157103f3236a99fe
z5f99faa0ed9695a039ee0393603b5120838f899d498d3e166bcc39c434c64ff1bdbce0254eb74e
zd8cf0555a23f0610f3becef30f2b4dc8d1e95c3e064b380fa7d934dfbe43ead3aee92273ce349e
z85186399db4fdca864e10e720feede36a2c208eb85361f2ad80b9f6f9add6360574caa99b2d354
z9a5e166ccde71b7340da44788fae4fbe1eda4daa99120760227e5c1bf4aae9b412d72b8cacb2f0
z92a22e2c85c9b05f20f74c129eda408c7bcd88b625e2fda38fba0d1809ec10c939e25448a22395
zc908081c8d5bab2e943aee9fcef2c169810881f3eef21aa88a16f398f88ad1d9a6cb6c9e93b7e8
z3e8159797e7b951d36cd7f97af51cd14909e07b319063cf79dc1804495764928cb16d0b812bc00
z8d29b0385fc66c90d96e9615449587bd8011ec18c2cf6a6718fd1d899a5b8c8bb0cd45339534a6
z6fc78884035388653069c159831ece851dd3b48df6b25bdb2639f59599c204ac7ecc5cc2b9bd48
z8ebb33c18f89cb8018a4c3d3c838e946fae3afa2bb0e76fb496eda7ee52b87f7bf4a6b3c644542
z04c4f39e6fa38ad05c404cd11b0a2777f8319b5a88c1e0415e387c69dedba326c88385b9ad66f4
z61280aa939e417ebf4f6e704f2d15b26256be02cd3fb0ec6cccea82ebb53e99340dd7eba38fde2
z167e038b5eca3e11911b3d4a0fed04e4919250950cfc7319b8efb4e942dd330beaca3dc9d5b4e7
zed597e767141a94aa11359538a2147504d9d9e51e62f9f7b9af27318988a454c4fd4f4a0af2624
zd58e36a133374b3d61e446ff2eb7196b932da8084a80673fc006e62a79e4370f58a09d971e265d
zda9d150dbd1a79b1c19cba07cf1523a0974b2628f296b24523428a5724e04e80367123aaf3b99e
z38faaa67e179f130d0b4222e814567aa95627c5f89c1bdea785845137b607a8131127f246687eb
zcbd5e4cd53d463521150b1edfb0fa4380ed09cbfde1f7dda4c61ee54ee8675738abb72d8c055b1
z670e2a50fabf3b4df1b52130772595465b14639872b81fd4404c3a3dc7e16144142acc4515f341
z1b40300637c1aaab394ce2f5cf07d252768b9adf95a43551b39cf53b1fe75c133c3bcac9412863
z9a8c1c56d47e7cb53967a2a3f32efe5cfaa1a65f2cc74ed866e13afe7718517fe5d498b96cbecd
zd102c6589103463814b69d891fc93b148f1ac609f99c5b8ffb17fbe7825d8628200bee9cec23e9
zffafd5fe3102d42198680fc560c1fa84e5fe37cf87912691a9d680d7b7ea4a3889c8a218e26b64
z9accd1655514c58b73b4bbdf536afaf6472f58e0c58187069fd6377560315f9d23ad54b523c0c2
z6ea4a8339e0ad6b215fcdc098998ebc3fa3c603ece7773e08eae16817c77e77b89341602ac8c8e
ze1eb382f5effe04e7e5261c4c4c9c86b1f584b0232a4eeb3e09c9bf33176608a22e19bb8be31ed
z06e7d40d1d944a644970f66490d5f91fc4fb4c98d4fc6669b1ef9ceb1c125c185637853bcaf73b
zfb34ca10e1efaa66d51b47bfc2deac8306942bb0306ce7d7c5e1cc0f5eba66a3cd62038b42c4f2
za2b6d5d2e54c630c2d4d88afed53790f83ee63e3087e7ccf790fd641db5441b8f74a3343a6a1c1
zda3369280fa3e7e583b7552f8b600e80790229ff1a23c63045260b58b8a53fe9e1eda9cd2db618
ze7ef2c23997b531965ac61ec624bca4197be2737a84795e6fb18bf7446ddd97a136c756ade20c4
zaac038b619284a97a19805521052302bbac3ec92eaf5fd0057181e7001dae03d150e2e29c48212
z0825052e1bb487a39b6236ab7f6ad0b5f6b0ef6f4bf1746540734d1d9c4857679bf71ca0329b2c
z3a99efab3902b2648e3c00eff05b4462cc74b26b97251a94fa8d483ab41ac86c76ec5d67f26801
zc1a8877a45994a42dd6827d7b724a6109916c37a93920000935377d461997622e27fee0cb6d918
zb0a0226859415ee240d996a91bc906547d70c576bba340e9f675ba2d8e21fec0ffff49023c32fd
zdacfe7fb4f6697c799a1acba933e389bd25905e2bcee25434edb8d653b36f796c444124203beb1
z443910c0f68ef1c46d2b145423111355bc5d235bb3399fd1154c058334cd24bf8507059bd0b61e
z275865d067c18b3cea1b02d5258988045feb58e072acd28e7dfe2425b111f846913ae8e35bdf76
zc87ad86f2bd9464cac0e4bbff029077286b51e1a784413443d4451f5a5443007241e64c4a4cb9a
zad83f657ee79ab1b587b46d0092334ccef2259b670f0a319a2e1246fa8824ab23c0fe145e20cd6
z5405788e3dde600bbcc7c3ca2ad7cb499727e34a5409f428d7b1d72b087c7a27e74712a2782ad7
z689e28580f2995cc9311a33e4b51714d154aa45b7dede80230aa409e07b598f212385e9fbfa699
z924db0ab533c12dc60dfd88332e7658e40303982de481154a7175450fada3f22f96641b4911966
zf18022d1d57be05f39c2946b0c877e2f28efe3c68c8a0e0d95d660f07b8c83c61e8c3cf76f874d
ze33a54c2018a414d6d4658e9ff71883b235eea8ba59f2123fdd9393e5dc41073dcdae74a73f9f8
z8e222efe93e192367c007ce95bf1b5f1531e9f44194aaa1991006a700a9113f47fbb8c2dadf811
zf495c20e9ee45ec6ab2cf0adc9b0e8d05907f382ef7cd13a28d8c04cf5dd93a4d6a8d150e2100b
z595eaa1f42d13ce93d41aa00688f023feb0ed05177e8ce4004071cae8a506304df1fbca72c30dc
zf8f336274220034063cdb857556e9521b21c98c300fbcabb18ae56e7db268f45fde75775759768
z31b6f1eb1a24779ca80de72ea7caca66c45263760eeb06d510e9682eca7711b14de6ca77ba1104
z289f38947e7de3d3670140acc0eed155bce1d1945c0b6b62375bc77121caa976405ab3757db28c
z5cc9092ec370c52d314a21bd5e01996890355242dfc82610209d49600304c37585aa1347f4f8d0
zf8115705e5b261395e8159caf1dbfc607a21755aadabb6fc03658cca5593098282a610f812cf7e
z7dcdceed97ddce835dfbf08928d441f6b2fa369453022826613892fe794f84f4bb2228b34abfc7
z9c93eaa271885e50da68f861fe9cf5dbbdb02b36a21fdd4192805bf110af3fa554dec3e2e35eb1
zc422fd3d8dc755b153568b0fbcd96ec2938cb481fe2dd78a5d1d8e0f70fd7819904b0a2a680ab3
z3b0856ea5aeee9e0b4e5b175ce94365f740d5b7ded945d24640a702678bf55f44d3844667fff93
zc82a64361c8f6492feba2fd01b9e7f9e72a82d3f4c6538bbf0bb21015f6538d0ee099940961673
zd9a86c8a83e750a216fc8ebfad2ebcbf96872da8291715f349200cebeafd3dd7c1d54820cd4c08
z9d71f1306442e1975b7efe093ee2e67721975199be0555591cc6b3921038c92b4b8fab81707c93
zdb8c85f3c1d3f52c1f6d79fdd2e62b2938e1c9e996b65bb830c5b33a53bd277e5f94b79407bfa4
z887d3718525ad2c3b5e764f01519afc1c9677f64484550d61a8f35540a7835ae2a5cdfa3081639
zbf5f6d83991d514fba5a0ddb5f6f5148328c35b4e40531fdf02ee7c2a4f298265e959c446443ba
z9e01a9aeac519702bcebead2e20c3381e82009dd70c82dee4f408774c9794171f87b830d0833e7
z43e11fde2751fcecc5ee234e374e8b93a8d671edb4fb2e94d72c2bd236b4d72248f785496924c3
z550106ee7bcc859c0f59bf17ffdd6dbf2a130a8e2909a9e707f5cc59c3550603f69a8398c7534f
zd2853120e53aeb36757c3682ddfe0b8259797390ab411cfbd484973e728aad865bd582aafb6297
z41c7f981a46d680ce051474dc3f723c2ec1e07880ea0ad47b68460a85abf3809071af1082d8a57
z1dc73fa2269c200ff87aa38caee0956f8fdd378e14a922f8d3760b97364da26df99ccd17e8ef4a
z99fd34771a6005946c022891b4cf10fa0e2b96c72006a27761f4749240c4b590922c344b9d6fac
z561624b30480602e44c56cd090e69042f527eb7c00b395f60442c44a8372c465952652dc18877c
z6ecb98bdc4c7d1f39fe64b7dd2f51d6a76f1bf5a147ae9dfee01d3cfc7ba6ff30d6675baa7c0b9
z067a1a580186c4ba3bb923931e27a59dcccb8456b5afaea617918a03609fffede672d10d5870d9
z104b694c66e1da7c0b609c224b84abcfb998aa2abe88834e549b4fe21cd5961da54e589ee97b11
zf157d698d8de64b986fca78a986333b251d6a8f6fd7ef7db35252d3ec0e02a1999bf8a3b6afd09
zf319eaf55215f0ae132319bfb97b3b4cb7e258781e72adf2219a916aae1c6b1059cbb931fa6303
z6f63c165e534edde95008f3239dc94dbe366dd839864af9f64e4c0aea379dba89a5639f7d5bb03
z527b7f694d726b6af289cf39e45ca595fa3fb4d1b97249727bd1e12ccd092a84645904794e4e60
zaebffeeffc3297c4bf51907c55497cd0294b0aab46b3a9c840c03b6ee848bd9bb1581c8517fbd0
zf6372a2c14fbde7f3209b32171ef1e6be93e5db78e153c6a8feb118ff4fa9112173fa1cca12320
z8c2659f1f64fd206aecf60e85580b85af550170b1e31ac904de202d1b4558adf51880dfffa0e71
z9804505151af6d6a0b56112804ef937d65259f1d9042e8e6a0cabe161eaab32e0416f51041ec34
zeb89bf327060668e8ba56d4eb40dd8a154cc3def40b86c0fca083395595da7a3e8a8f9f87555a5
z76592748fe4f20a50c87633b862da5e92909b91c050dcb961790fac8a82489fe3919b6d161c337
z098c047e8517a3cc15b1103727f3747a569891c5e4c47045035d59858d85d2dc61ec74c5a05494
z58d731cac0cae1879d46a972a4ce82badc35695ae56cb4105446fe3bb05da9a947b6c945904a3e
z6bf98816c11f57cb4a18a7916e1e52ae1a34731aa7b920c2533044c51eb570f3bf21be37f6bddd
z910d59f767740806e0b1b9fab32c87b720b103773e4a8c8ec5f31abd3d03266c075ec343d6736f
z46aae962077abbb3b327a55dff754e2297b2f2b100ec502053ece43063168ba16058520142ed82
z4ebfcb7f526d42052c9eb56ffc992ef5e6f1f66d946161a7b21c58637d4fb4aa493107e5c39cf1
z0c7b5cbef1fa906ea188aa33e36f2d669f9776187a47fd32c18020babf06b4f79795c6612df974
z0eeae962dd4e74db1aafdeec271d8cc82c3a86049e566321e1c7f2ae4d7211ca5c37756ef191a7
zca5c6e027c1bd2c3acf930cea2783b526e65df844870d178438bc70badf16eba91ce72c27641e6
z28ea13c3c1ed1f226c08e954b1a115a4fdd102199319cf05dee2191f1e9e3801d83e22ea8c7bc7
za2b3d4cfdceee5f1088047b0b88914039a8dc3558e2f12af575822c7171a85502fdb148de22416
z92593bfd862f627989d2e6498718ac9d790d506698face9568671183ca697d034ad134c7e9984e
z6627c8d0cca676c13e094c44b40c1d89c2068b1188d4af92475a353ca0379c09e2a2433255fb85
zc234d483528e1ce3de122127b0a770b834028e3e86a40d46787e6504465f996f941e193af9b988
z1ed45103b8eb4e3e687fa97f30822b9fe2820c0f37401ff719a51043f2902a731cae30a30c34cd
z1cc99a67b84bb6bdc73d65f40e07ec219a15010d46e823c7c990933e7b0bc2df193181aaf7d366
zcbc36d125cfe7cea7ef37a10525f99022e5b58cdc1ace9e3393b36ca7a022c8f823f9e2a3d6f65
zcac0957d294274b96e64a89dedd986de5deea7c92176252a37155dd4d754e1388e6fe26e9823ea
z75513e29bdb780a918c8f93e6ef26fac0e6a65b94995736f0ae010493fac4112f6773c52dfb6d8
z6e5ad8fc46510db7cc1cafb59cb9dd6d8dfe94c938c8b5fda6e7a3d6c05c54c94a66c2b652b7e6
zd4bc07356f5c34d3653f04e71cbaa3ca75aaa70392eb936ddc58cd5c37da2450ee5f1c0ec7a692
z3bb6f938767e570763db01969d0e5ad2916e6e6a91eb32a572851c63a9ce5075ef0a936a39c0eb
z296055485bb3924474a7fa8d3f0d3bfd54c54465f467c44f284ae7257dbce20d5ec5f01e2daf3d
zd410027cd7f290d324e754a733be03b96e98dcdf708062e53ea0b652bf993623cef5ef593e4d0d
zf4f32206bd51b2dd1c5d7dfd899e50ec8df0a43a2839ecb68461485e6e4c73cbaf2e276f57bd6b
zb64817bc6ba293b27e918bced1bb50a5c907c75e98285a16e447bf6065e52a9af6291707666bc8
z938c56d259d30ae3843707e0f8debacac11599e0554885795c9b4fe720d636eed273d8acee71b7
z6224faccb3cf39f26fde68bc50e934520fa58c9f24cc054dbf5da16a07e53e98945d2616b4f666
z0db9eefaefe239f150a2700ff113908b3fa485e8ff6a2bfda058b405c90a9fc5006acc82d2558c
zcb405f3bdee7dc6151fa9167f4ee92c3d51791cc7f39f84da5ae0dbd31417eaf78519776d572bf
z4003574d0c11620bcdb1e66b2d0c11a7427ba023e2233ebbbeaacbc2d63629622dd82d8faed34f
z38c2e6a210a7e40b7ce9fe4ee1c48aff34948d99551f12ba7139f68decef67b95447f40d95011f
zacb3e1c21cbf677b6a7424e1046d3736374b3ae631f2ee5f040a595a85b0ce500db18dd12f6f1f
z99c45973c445225d06f1ab97beab998c12f0d3b1a51bb459514e7597c16f069e45479accd915a3
z2346c04c8798516a1abd1675e2c54d9bd601ac5a3b0c0e469be58feed9db0d2481eb91057266ab
z9cfcfb6a36aa03f6bd4814dff1c0608cb2e181bc0688174fe8a71038306c911661deca4ca27738
z93c015411946226c1c8564a0e9c22fd02c19f27d2c8fe004d0ba43f3228f90ad204cbd5a47a03f
ze386c932c811ae15861bd27221ac03a2ecaf13549df61eb002ee79bf7177e2107ff066bc24d5ed
z6c266581c9fba7648a5a1c7641c4e266750cd04b4964f47e83efdbc9036c398dfce11ffc500329
z9d8751470b69ab6440422f0283db316ecdf669437bba69d46437ea8e2719d0e59bac9e68b23a46
z1e41e911a06777431f3f14c222f63983f8bc59e1b10c7d9b532d222d271175d5d9cc6f226f9a70
zbe555c010969e8302fe4e8f2efd3ce12246b1019314a89704905ff043a762a40f76970c28eb011
z901ab347277da05cc19e05c2ee1d67493dc304a3aacdda81aba18651df6c96d318160525e048de
z967a9abe3c5b319ce3447b117ea8820c93fe52bf37800850f8c760e0c8a3591abb8aaf448756a8
z9305d41f5ca17eefb0af9dc6598b4e3388cc0733e16c47f34b9fbcc43fe5147dfd1fd903ceebd2
z6efc1fc860cbe01ea33398475177afb7d8ab6524a2ce3ba0753a535abd85598ded1bbc0018a108
z77e5b2ceca62555b59485ab50ffa2a6cb507468fb53f069f55041c52ae23f27c107c4ffdb9ce38
z7f6b21c2d20ae6b15538d2a0bd2bd84c6e0ced6a2976a93954935506f68ece2b46b7ce6b8b7126
z6317aa30988ed210ee10ae8ebbbaf8dd0ddab276c4a8884e8c6a46d31e21e6e472dbfd94d66b03
za26895c4de353595c661866334a3ce638444a1927e486b9ebb44c62cdf9e1a5745fc977a05a2a1
zdbf4fcc98364079e7afe7a9bd47bf88ba8c60785b5592f4323a82f9063e1bbe05188969adc8486
z4fc93b873172bb194981c0b880cd452c7c22ae47042d9051c70ce22c32f0c64ef932f6bcffefb9
z0100b12da191840afe386269f2ccb8e96d0b7b1d37d4a4a5b6f87df9f0814f0b12e5271d80e82d
z5485c03783083682685d910c6646a89a9b66231e0cdae418f6287238d947326f465bd8be3fa83f
z0816f3f3961df1b5fbc5f46d88228b6163e029103f65f005c82b0bf23abf72234becc388f7d7e9
zacc0b521f6bb06ed287f5d587aaf24af755e5854b308ed2235faded21aeb3c98b5e94a6d33f380
z0217e22d6263af0abc74157aed97203f00bf000e4744e353c39f744bf422d48caf22fbd36f60f3
z5d5cd714e259b37c21c2ab2f284278925a2d4026f9d39e35bcf62f80bfef2ba11b4ed9fc0ae49a
z046e9b13a90efa713bfaa4724707ac32604a8e36213a7d1d6c9d6c05e785b14b449ebb9c3fa916
z4293297aa623f84e3193942ddc1b286b5a49e61ac6d4f45eed850d9ae889c4dc7f48c500cf5eac
zfbc9f4a3b22384ca9e2a072a9415f079d908009493669ba75e7c783a3e60ab553a18c64346d62a
za7916103bad510870b80f4bec2bfac0f635d47431bd495a769133344cb4bbea6d3f339b1563e66
z0a8208e6cc8474015e50da7cae5871efa80636c852cf81cc2e6846a89563c2967746a15abac874
zd8474813bdadac6b7d6e11c2a0f1e7fcfc64032f7e0f3226c6f92811330e8be2f8bb3058171aca
z9f67182b036fa34ceaa3d7a043f7c6b64059be3c2743f3ca79c7f08b14f2692caf8695dff9eaf1
z9e572466776e018873a9912f675edb30800ad046cf62669464d2ccd586485f68e8a1ff9d14b3f2
zdcfa7edce21f61f9c541f1e27af251f2a834b42c884138abb208e123eb82d8ac7e3e6878f18a9f
z0ab7b3bbce2ac6a23502b99ff45246a03050932d9552cbf61a5fa18c6ad5bf4fe2f2684389cf10
z0ddbb43cc1beb808a08b8bf9c02636936357f0d74d3e9875214fa2c18a4d2e8fa423fb2ddc0e85
z3709177ef3c658754acb213f81c7c50f6218834deede2be4cf5eec2f4151f31bc427297f11ebf2
zc7e5ad8d154c27b5d1342e9d509b034fc09b123edce9cbd88b636d24a3707e5b63dcc1c5714e97
zb4d36b44ea05ea7eeb346cc009d70c5d7cfe227bf721029b5f353a3c0dba6db9ce7d7d2737d9b4
zcafcb76f2677e898072824e1bac351e3c781413c56f7549139209b81368076d3232f60fadfa166
z8d22a3a08d84edf4b0ea80eb84b81430b31311887b2b3567b98c1ee424b628e8eba5a2d81ee189
zf968aa7b9cc4e65cb4ec85ce922985ed30602698f83f099325782930622cfc09c4a18c6bfac622
z9c32cf5040f6e242055181b1c1c4bdba22cba338b63414f2fab9df2e01acb25d8be6f307054620
z7a5054a1104a5dce2d03993f6c8fd8eca692eea455d033ad4d7d28ccb3b6789935088d8cc19801
z963437aac3fcc6bb05df197844bc85eab24649ca376463df04d5b6eebf3bad61470e7ace485833
z96509e755d953c736afc97a8d18631fdcb7c9702927288025d6520b8af981aabb7f6c00fdb4b49
ze4619f1dae3a9a63d420a9492b6199a2a688ef7e154664c26204f8daa9d6fdfa5edcadeedd9e9c
z9825fdb9aca8e8472dbb019fddb835d8a88a9590c68b364e567f38e5ec818b0e93125d5e7c151a
z655d267a0bb8e1e727e1c5ef3c620618cbaddd2c787c76408332b4f3873ecc5bb12b2faf14bc29
z9744a6fdb6770db6f68e4876f849d9a1b423a0683b35e08ebb912e0d605188facfe1d347ca8b3b
z9194863650071bcda5f6ebd3fd2afdd0c03744a07b1f38f0433e3f5af8bb177d24cd08e531e766
zeb5b933ff948bf25d3833b50a4217b7b946c1bc69eeeef11ceb6271fef27f7735174984f887386
zcf5d723e8cde84ca5129948d2a2b95a0a8681528acd42073878fb745e6b28ebdb74ad8a50caa53
z5b1e6a19c3497dc5bc876787f0b84a7bce2d5b49d5ea6bde2776d4ee0fbd771b556ab2d2390431
z66c5c6c222545e3fa0b52ead756e5d082e1ac8220f4d29127ed3c0425999fdb0b2f0ec27ddde4b
z33b4d3d40587149d2fb2789dfa1d947241f271351c8eab0915e7971ee5299c05811819147d9221
zd0e21b33c3ada4a4a75b63942050805a12718839c9b3a7088d95ae264c2b39c785b06f095bce1e
z3968bb52c08b296dd6a032fbd4264ea8cd2f1faa00e485770c3e1c0ed53f3130510a131c3d12bb
z596140f37f0a01d945a051790f2fbd19b53b3c3e65bc167ac0428fa0a497f722f4bb23e1e549fb
z8b1fd21d5d8feff6f401edd8386334f79fda10fdee8bc9b69cbfe1c9a38a270d59e337d9e60044
z5826da7ffda8202d23f4634d556264faeb42099e521ad8c254275702d2422b6b138bd033ec1aa5
z97f4806a45707067238ccce292cd6e3af13b007fbbc5293843011976b4150570ebbba0ffd55265
z43297954d51d04830b2f36045091a2839a98534d0d5c7686e7aa27e620e8a1ad906982b20ba798
z900487e59697252715ef006e5fc61f9f2b70116b8d4d315370d2a63da0359875ff5a0d8b4be2b4
z15f4491a8f8f12818da7cb424fabab289a601bc2622401e051db06edb70ae853e9caf285718c97
z24ea8e4746bb6f8ce80f56d02fef7bf77c44b5108eaf1f768cf8efd6f67820cf3bcfefe4e1bcca
z9ddb07c7359054ed007b55e2dee1ffadbf1283eb91c72240c5a33da762080b34e5514cab519f3e
z9cf53e36b9e8ac2c906b1b920b163fc241e0b38b8e892604241fcd1dc625a9e9d9e9839fe7f7d6
ze732f199431fff6737da2e9730dc7b29cb40f0ba93ff11a5ae100594d0c11743e76a0d50bc7261
z54916587cb9508f64dc55a44b67ee7b07bc34863e54851b0ad3c4ea8331d7b8c96bb450633c9cf
zeed195da90de324c9fc9936ce4d71ffa0c041c254fa8f3e89c8ebb82a1eb11624ad6696df58032
z89e3110ef27935ba6f9595d33c7cbdc01efa984584ec34bfc0608af099dc6ad480d70d1acdd4b0
zca0798f4d25b153224ecd5d5eafabb2b054b1d13f3a973cde365376b25747abcd5f567167805fb
zc8db3802a4cea05fab98c84fc753b0ed33b4f6fda2956ba543401d8a97511af0c9e304abb0f7a0
z1a46a8e44703057ae3a506354bba3d740bd6f3e1f11e470f8a55138fed7339ecae4f9cc326875a
zd60a973e55cc85c88011b6491539455828732d344e748b378e7a1e3472512fd333b636eb236273
za7679e7931480ee2118b7b73d38565637a532afaf7cd5a7e2dfe6fc7e4da26f944aa92d9347818
z34418aecfb1e2218e192ebf241c8e3ec255115534c90c55d7dfd7493b364cc0b4ce488eb2fb0ab
zbf884c9c4aa6f11593fb88f4004df35200df0ed5373fc5b992d838e9a7c6533d5be81e2f9b4116
z4f8e7f2b84c91ec4212e9140ed4c14b25a62801aeffc8a412e47e5de5db405bc506778fa8c1f07
zb79ff15ea82994ce8c87cbbbd9dea1df4734a274c51b972aed77071505adcd2632a6a358301768
z06da8b5dfcd35b2a64b0f8e6f399f870d0c8f231e012543ecf9205fceac3c081dad7edb63df430
z81c994bab2d71b887832d53e158e38efcfa897679a059801e4abcabc403a8d4333f798090da2e5
z44577e2346d383ca8a1ddc9422f6c4436ee983dd422c231bea6e32ac3681becf01cc3b7d038f10
z6f6d22314e78b73c020b5e1c0e84b4f1265d27f28baf618094e1d54501713a057d0581000bd5dd
z255141d13af8db03587b2c5e55a813d232d86554532cabb0474f87d14eb53ce27a9d42c789774d
z9c5b6d8c4dc541f0691b075d61c2a445385606e19cbf26ba40386306e311b583e34e03c9eed1ef
z30657178df92d41bc6b646cd9e2e1f2e2867b4c725777f2684c617b667a3cb9334fd055fae1181
zc6f479a9d6c0218f829ea85a987e9cbd762d1413729fb5ed94f8e3f8d52f607c5480a1710d7152
ze7dbf2783ff1a80b5e8d3b02ffbcd77a464b7d33ceed59f4326e4449ae0e8d3ce62fb4c7eaac14
zcb545e0a0840d1513690ca6ad6ac36a52976cd0f5a33bbf079f31c771eb8c8183105f56218bd2c
zbad2deada965b45c66ca01b1dc146d482dfe876335a1589b3be6b14afd4afa125bf28faf611c08
zb4953323ce9a9720e2a806507534025952784b2ea468d09e1cfea9a852693a386f6209971c296b
z83f6a923a43ccfb0e6a0b43a0f020503d5dec8b7c90f3444ee9d24523cd1a9f137238a4f270b55
zea4f34128ddbbe6c4a22531d12614aa23d8431ff7b4b7ec3364d4f72b91c001c8d2fb617664c27
z916abb7e5ff216ae75c187c997e2e971305efcf88a933d0e40f270725511b78ef55ff7584b5497
z185601510a282002b31d889f2507afd3c9d4abb6a2c8cb7532e6d7b534da8e1f5d3c286f7b75db
z56978c7fe90ba30560445fc8c41267e4a285f70fed023e8d81053dfd1877fd65b79c2b48b720d9
zf9912f7a3985ebacb114839828e56e4f3360fd0f906f98e9473084a3495f220b244213a2c9c002
z39bd41a262aa54742644b47ea3db7184b46b0e33b85ac9601e39acdb48b30c6ba9f81ff99a1f18
z612988fd0eefce7d359820259005cc68ba2d076c2d6b0e9d59eda44560e31526faf89bb3e4eef9
zee16d30bde57c6b1cb9899c94e2cd64da1361a2497f1e8b41dcbae7f22669482a6940e2e03dbc8
z1f716c5965ec84235a61c19ccdb7414679c4344a9d0221524d2b0ec6bf129459f73f39ad48f2a9
z63f291e0c1da0fe17672499c4813cbd657335c5996ced42460ddc2398d4fb90dbdaeec1b284afa
za3ea2c4f88d486ce5fcb3364d21bd81d67c2b9b1fd3c59ecbed19398c287529ab2cf4cb4c0912a
za8c9e8c7316a82e4a8096aa206c72a97bbd946f9902cfd13b2772024d95c6a613ed1790f746747
z24c7835fdfd6407be6fc66839adadf0b9248897761c3f3f613b712dfc2290162470d7abe446fad
z99b901baafc0b0ae3c3c84452c041b54475215957957752b0aee4ed9867a12a3f2fb807f534259
zb416b7cc31e81940d986590f2f996c359e4db2cc5d67f6afa137a913d5087cf77f18b1f2fc7bcb
z4a74f446f41608dcc3fc022816374d1f566007006e0a4b85337066e550361abc284e49ba7c28f6
z9d6cf89b23046199b52d1ea9484da4561ac5903f2ea338c0be3b5d3b78aa848f593810ee58c327
z9510d4e2da4fbc05ee797a7a9e1e92b897b1192936b9a31a902af5b4d08c087bc5b866c4acb530
zaed5e1a4de2cdf075c0160fd772ec90fca3e0ba0c5593a84445638639c57c25b86ca5da730d54a
zc5b7f481d2cfe0d23c0fbcbbc551d4f1e3838fc6d7695bc0e1f0df927bb54e6534781f65e52833
z897c41df43c3668664b5ae5fcee20a59bc566b7428388baad6a17a72ac5ca45c2c5b6f83cbcfe2
zca8a93d337560b91ad04d39be26fc33a769cb402dbdabe7b314b4f21a4cb348afbf0b26593acd3
z0a01d12b0ab779266a8c5ae5625cef5db8d470a96b8a3e4c5e3b8abf67bf71194f6a658a42b373
zb8661a9830748747da78c99a6ad3b724e35141e8df42dd547aeb6718e3e27b96a56bdca6f9bdf8
z58f4cbed44f947ea4168f136eb379a085c9b05605a7d9237540181257d7dd28cae6810d33a9e3d
z897ad6e8df6f7d9196fd97632bfd9c44966158c756627b8de8933637ba6e781ef4f45e7a55c4b3
z1ebea00e7cf202bf41869cb8041d685b4d6bf34e98b8ca0b4e6599006a6d1ae65ce57b3955e7de
z550a1ee72f724d6743ff027913bd03b3f0b35da9fbbdb5ff21dbff1c4b4ca5d9e3a39133e180fd
z3b13e9395528917972f815cd50796e0f452c21a3375f86c5a567566a79ed11677a0a6f2751cd5d
z645acde27a2ec28d2f16181eebf129b32741534e9142e418c46d75e87718e1a39a95938ff66558
z64e3bfb90d7c8185e0a4ee5ddb57c88113e8e9fc70d495b4cf33418675efbf8e9014cbc2f88144
zf29a8cd005c4c45803577059147344d2cc44422307ff7ef3db56094f438bba88be464fb3d08c65
z40e2beb29a224e2b469b85e0e0a46ecfbadc49b7bd0ae40fc093233fd82563a53634bdace2056c
z3f2fa9fc66a3174be62b2e1a267c587173dcce2f1d84f94d8570298c71fc495f91c113b60a2090
z978d7ff9a19971689985444c6ef211a111f998b35d143f9744408cb1753944291871eb6b0d6e01
z1aa53a583cae86a11df980f8da978732e4be4764ed9db3d2073b086d53439e5054fb7f8be2e855
z4f0e8924ac6221730cae67361073d3214f9777a0bb458b8ebcf7662846e58a7e9209a66bd7e2c9
z3f172e21b778244d7bb6dff2a1603a8d9fd921e8bd42b056d9f12202b5ecd12456b59468bf1c2e
zbf967ed30bca29167e9bfeecd26f686f021c144870f77a2139a8363b4aadd1986bcc820d6b0e46
zce9995e5284934344b7529353aa2b4fe1bcdb55ed89573d286484b11d076f7aa9a7c8d82392337
z1e49bd64858f8be654fb705fe59f3cf3c527c95f1a1dde8ebfa8f78732a6ec74ba65b43d982891
z0471d722b589c6266f9352fbd2d12273d85d4468a3ae8894805fce7d5794ee21434f0d9ef72270
z3e1f60680edf8b3de6844505d452b76cc6bd65825fdc5e47c39f0b5a90bd5054d48f61eb6486b5
z204f3a47f5514eec6ad3f66e630c34448d7f3e4ac9a8503a772e41782aebfc46333afc49c969d3
zf282adf701e88b67ed03587e4f85959864b57e8b47b005b68bb1c79cee7d0991878e7886c7946a
z179a40dff5046bebab17f457833aa8fa615699a42e881bedb97d12a2a7fad714e93db81cb2d7f1
z627c66c85b4aa70e315610ca9e48288b7e475a3ce8056a13871de92394c672b8bcfd17753ecf67
zea4a2a4a18ae6d7920315c270dfbdc43f8fc265ac53da78c35a57bb24f829e9a248e35e21075c1
z5eecf8b38bee325f575794deda108f9677f581618c4f2a811a24fcf255df6dde5f35050072d41d
z308b2aec6a7e47c9bb87ea1490a7ba3505492d4bfcd98f956719aa4e989e56e46838547fbaa1f9
z3c9af3e60b3e8840362b06c85ec4934cb24025a064d3dd9c12215b8924c363517585fe87505748
z53cd5c79a473160bc98d10d11ba331a362a41a6c5b0629f475195cec4198ecce724e41be4ce3a5
z6ff13c401b82345637da3ed8150c076ec64d67814e6169044cf3e5c30dcf83428efa965cfd74aa
zfbc92344f2f02f4ab2153da7e53d9d6ce47e96937be280b57d093d03d6ca794126468faf6f17b2
z04d2acaa5896bc64ca213b664acad3d595afba9528808dd9da027b7f25dbfc22a95a677ad62981
z22db835c9f6852eda53392c652e4d87ca40764ab5c908063c5f9102857c31a9378d9237f931010
z309565f10f9a4e2545e9182d4b1812f65d7b98d0baf6e491e36440a948379f3766a3b1bd328e62
zce3bc594c719de2035dc42b825137f7bc629215a3dbf0ddc5aef34d95b35cf4d7dd449f8dd5fc9
z512ee29fa2ac94bbb577fff2008ec6f56e62b1b9bee53a148cc63dd34fa46754be13aeb229e672
zdd33f972b094c7b8e66d6db321b3794eff3bc13cc24fc9cef1596281c303a6e25f298ed5439c15
zb79142e26628863c9c4a4eeff673f52e9f55026b9ab1b560199091766e2c0439054f9b6d2b16d4
z8e9368b0e1a9732d236fba43bd188b6f7b5c396ebb67509e3a61ee3a724e81d63242bc935492c8
za208f65afad634d4893a7ea80bc9f6e746d4ff18d0100f3cb3c7682e5266f7443a1ffa5a68f188
z0955b3390e18beb990696fedfdd9999f00a9d7825797acf218f4a56dd2bac2c454202c7de8a1d3
zaad3940267193c3004ee08fc3305e9dacefdc6f933bdc76a4148818cb3f6e12f3089aeb6df8406
z9add9ce9cc119a3b3b456c4eb1e5cd6e1168acd2bc11b423177524b600ca2b65a1e884c3ad45bf
z6c969c403f3611360d74e304330fddd7d464b90e52d941dd48ba62b75efa643fbb3b41f3187df5
z569ea14235f0dc645a290a55fdbe4370a866f8eee572c590197203ab9d6e3da8cac20e4c600f6b
z01fe2c48be970e173d77259c9d0371c1197738ec72e0ad276578bef5b4620a8d4cf24cf976671e
zec7aec77864f8caff4121b26eca93a9e10e7973d13ec460b8dcd077ceeae5d506a3368bea5e7b1
z74b9509b1a3ebab4832a74fe5bddc36c87fc20ba5e86e3b1fc029ef4149154549257e203315407
z734a7490c9fc8995b6ba73de5e148f702afff122163ef2d1bfae7252b63bf9da44c53df878bfd9
z7e2f1d4751751388fccb5c3a3ab9be9a563213d06197c47200156ebfed6d38bb6954ab48670fbb
z950ce77577c07f6bee85551f6e35597047d9935b744f40d9225b5d6be32a81e1a50dbffaa24124
z63b651009ffd9db275727544f2a7f6cb837d31dcb3d8aee3002e6b4f21c4fd21333978243f699b
z5e75e978c3ab1d674a06b55ed22b37eb478193d56f21d40caaafe88b719cf2073c904bdf3f4fd3
z59a8a2413789f15cf60692799c5b9c9ed01aeb5c0cecd6e940bdc01da51e009ee72a83ffd60e60
z126ff7810d3d69f39cb917deae063c651a4565c1f18d108d1238fc3c8524323fb5854f5cfb10d9
z6b9016ffe15b992ad621c06b0feb53ffe0897c428dbb7c6238da6a7bd2ba182dcfaa10224f3edf
z70ffbb777f13a516a043d45438705e08755a375b94b41431c2bf01dbb65ae65205f84080bef093
z4b9dcee78c451f6ad10a62a078e5e0df6f3639a02e09a54f123dcf80da7a47e442e080364cbd4d
z96ba1c8616fb9b1895c0a49944813181c0a25e4d4bbab638057ad55d209467b231bd7ef25c3516
z0ff54110e675d11043c9a663e324d6f3ddbed390b98ae8f563f6acd0fb04ca4a1b26926e7d6285
z19f86ef7a07f588a95869195f61e0c4d39945d3252d9d4c654d4c2aa7ac3455ce31ea3b3ced81b
z7f8f7610cb5ca32befd9786cb808a65e9d64e2eabd6b19a886b4b5e74acad36e6f5729ddb7c62b
z072824a21fc0afe28ac8ce7982559fb97e69c7ab28f02fc0506681a74c78c365be0d295cb5bbab
z79e1878b2ec93be4916b5ed28ec2955a9a1425f745c9d2e1b603c06d6e6eada823c27c8a4631a8
zb670ca52bd23c0780e762b3de2a6b7c883bef6dec8f095da8aa53d5552f340b55a8a57c5514f6e
zf4b15a21139c0764b4776a522dc3990d0ea33e8a0c401caf8ea5b127f2efdff52f38466d2346b4
z3b502f8ae52e1ebec8484b916cca1ffe14382edee1c9bdb722e8772344f4afee7bc70f67b9fe21
z9e09a51f9a5248ed1c8a6374c0bc6ab5f687433f03f5f2e6a3ec5384f59b82c1c272f99ec16791
z093ea687bd4136f7d1cd26f333b6d8fb79348298befc73b01bba7ecee5e72bb746f718d399fdda
zc5282b05447d51b970508ddec441cf40d28986c834595d4fdb634dc3cc8f9baf308954c6a88246
za47306714882cde1ec1b50b4f44082dbc64035a00523e272425a440df611a8e55d5d9f61209b4f
za090f5b8266ff3a6d0dbc14cafcbf3dcab893859a6eb7a01bf9220966962598e16007339322110
z84ed67d9d51487a4337371969f780d08800f523415b7efbd2db8eb8509289c7d133f66ab16d2aa
z9f3c29e523c696d5348e4a1484ea1760b0d1466c441e51b000e184b2cea8f4679a69b8e7cb6a18
z1ee2315234f0058b5dedd1bd8bbe71b192a0346689bfba00b0a1fd4d495c21fdcdb75c8f3988a1
z1ffb81e8607660904cceb4ffb1413768759d6d39c1b59090f4e42010abf6bcace5c0dee6c3d230
z33a4c08299c4a103fb5352468518047228783c2d8c5caea90bff7d6e4624a1dc4f00fa3baf9c96
zc6b289816afd09663f4fd864b1d2347188046330df5ad0f5d649ff22e304d4986648db1a919f85
z86c9f0ea17a005f6357b6a099616bcf36505ba422d1f31cde3a510612579e4361476afd7886cd3
z0050515895641ecf47561bcc5a3dc186ca082d2ae42ce88b552f99c0b164af8a64c14baaa91029
z9a9e17f5eaeae8abfb0d8ef07cd9974a625201849b72f099225e17a3c7b5534994489aa6b23c6c
z908602a1ac66c473038eb317f0f78122f1abaff6f3bae54e2740794461f9cd91dfedfe059aa7a1
z3d83377368e5d97a8100f149ec2ce639c1df542485cce5d372934b7af51855a3fee67346fb1f24
z9c2e126ab3eb249a58af73e89d219e6d22c2fe1e17f81a7d914029e4e4bcceba876bb4a6de68cd
zd3213d470ccc39587ce9708418613ffac97c3af0d08a234b62f0ef192d4b08a0de7871fdf4e9ff
z28a3e5b02e07d8ac21c0eef5d7d38331bbe70580ad779ca82ff882b833e8cc7a27ca2c14250691
z553ad032e35938ca9aed3926670b195b41184b9580770ec88921c72f165f04b2358980185feea4
zb48b3cc5da73353584325cd521b6bfdd4dbd27345574e6e2d156c850a2d7189f702cbfa0829b0c
z263bcb2acd97402c237366dd2b98f822e8056b80e294d3b55b982430bba9ddd78b9b5a790faba2
z047d11b510bd43b3c337baa91a5c002c626b6689b613ec5c375317e83f71292f40b39437b6ca97
z81c4b52c72b364448faf9a9fb1c7f60acc90854e2c595b76a33b4cb4affbc07a3bbd6a14ec28ec
zde5d4cbf34f4715208093d5853b0b77834ea28cd64d2760f8cdedd435a156dc16a30200fbd6081
z53dab933e1a9360b2c8c5979a24a45bf3c5240a36dd1e5a46ddeca113a4e714cf6baed09fb5959
zd6435ee725b18771c43734a65e97dc1f27e4401bad3f7d47576ed0ccc7fd2b3c7deafa5d204668
z7c4cbd8abdea62608de2bcc21114777fe10228949560410dff9da579927e98bf81d5a75ee88538
zd0532c2b6921dab4003b1b532e9d6c47975651c64036182176a40974a505ffdff66839479ae931
z0041b7845eb88f5780bdc9ff887bc24d8e80c054a24d698c03ea5e0ee79daf50cabec6a8fe1bc4
zb17675e021cb72692949c368813cc7e616bbed08a4522476958012fa6d62aa6599ffb869d9aee5
z7f7745a6a6a1a46d23063a0ca8d1c753c0aeb764d3c98c2fb059595c905dc32f4c050d7cb04d15
z91a2d910fe327e2bc0261b784e7bd08bc899a62c78e67ab54701843ddb3b5bceba8398491e8556
zf05a56bd3b146ee08e4dd37b363a5366a91a2ba25ce00f36956153fcd37725c73cd7e90eabaf95
z53b6d4b67ba64e593bcc095ccf0028c0945418a687d99e07f052b4dad30a15a81c678888725236
z58d7a6e262fbef8714360af1b71e847ab1c5b27fc7f4d1589da3dfe03e462230d837e05d3dcacb
z5173283dc40a4a470cc04d791d51b57cd8125fdea686f65363dcbd4e917c7d9600c73c717d8ec9
zffa2e9ec4759ec5d805db94817d53f1a09bf1b3679c69728ed1bf8af39afc52d9b2fba955d9ba9
z92131c0cbcfee2c2459804db33296f852b96d6b82e2f5c5eab9339eaea97be205189a713ca8840
z2cf3aa59d2558c5f3eac277fa950edbf43cc5056dd6fb11177c8c456c0d58656e5241c04dcb854
z2d13245fdc14220217fc9d8185d4b89cea6b8887ca778eb145fe2604fbfb6a2e5d218622c1aaaa
zba6a282b353cff48ce5865f35aca23e0147ec4393bd1cd61f0e8da7ce134de5c0e2f12918a1f18
z51c4accb2dfd3e230ce08a700c9a14fef5997e220fbdf4ae4ec5f74fcf3195d78b2b94c91e8f3a
z5cf23c128bc46b8d3960e1ed54e5c5e8d49ed2750f99056fd3b08eee230efe4f8ba2287bd7fdb1
z3c779b6ef12ec33f8de47e42924669b7061029518b9fa01bd85896e99d5b5feed17e1863d3af1f
za2ff6ec155e7920b52816372c8316efb4d5a4c5b44c524aaaba1db8e3959754ef9ce6cedc6d7cb
z11c2f026d83bfe6a8bb913e4aacc3f72ecae810e8e3d6caeafbae32890ca33f5fe9583594a97ad
z9eb785697747fcbd749388e57408adf77ee639b6ec2abadbf4506da6a1ce309c17c6ef30cea70e
z28015a077e4bfcd3e92c336d2c85d51d22d89f965036fbb5d1f612f7f5f643603c84832f0fca1f
z0af8fcef6a5823044352e6a94bb0e53ebb1af7f8ee8f8ea620fbeeb35b34bf450cd3d1279381c2
z348e5063cad16a0d4d780654849cb451088d4c33aef93b6286634d9be73de8e014739236a15fa1
z8c14da9e15f899caefcbe102a9264bc082831a55a51b048c877225aa063e76f43b03de0639e0c5
ze8001cd8971979a99d56a177be93ddfa896060ccdae09de1cf2a804b4b85e4b2c6238cad087b94
z5a1d5c7dde2290b4c37759c202bbcea593039789fb19c0b439ae245ce2e96c624c29b856f9093d
zc8990e6360e13329b87c458708468527abb5aae8e37094957140ccddfc90a9aa6e648d35b1fd67
z827bb02a4be3fb70fb3b7685bde0caf2194a7ce1b35954d19a8b5faca78cb3a237042e44912a15
z263bc891927307897df8a2b4207ea2596fa44a47acac8404ff73047a50c30ba935f2844f12de27
zccebd3eadd0e00535b5943e4d9f7f079ad9ee808985b9d3bb6c7e588e146f792da41d3cc265c89
z96bc857e21fa62931ccbe407a68c04e89941d092a305fe28f8a7413a634e8a7103d973e3eba506
z20c7b225f432cccd19cfef9d5f05f4df9ff43c51a68cee78159297aad7562ae00d29204d32b342
z608b56179f8bdd546bd554c4da8c92e9207fbb7839478b7213dada3b3bd58875ac2113a2c9e3c8
z4b1d51f8ffc14f5d8b1883f374076e811702c139438fc64c9d6a54656072f7d0fc1efc8d8e249c
z64ad7cc0578747a0ef0ec84af37446b2e14add41c4824ecde76689e92c4b41f4a0bf0deeb66a0c
z1b5eac32118f7925a699fd7297433ec13a9c680af66fae75ee80c4b5c3d05a4961a82557c42b80
z8fd1713fc8f6a6cc65d476f0fed65a3cd272be2712e1dc5f8b21f36c183eb67ca3c0677a25ffcb
z197427cad5cbe75ca196f354f2d639a3ade9cd92b0785766f353bcd2ad5ee4be8217bcba6de054
zbb614e57b8d797809acef59a95d3947c67af04baa72028c14d43ceaea6fc0e4f2837cfe6a790d0
zf787ee9fd0c541a0318095734760c82d769a15459e12b9fc12a8b2b2ea026cb8d42d345a8b776f
z39d23584454123baed247d5c233a9a30a68c6aa5650b36cc75e464293ef0a3268ba6234d543bb8
zeda632d81e26828414707eeced04104aeb40b9f10b5a1cded701d4090edc5cb37714fe36f47fbe
z91d82c246aadd0d69e35001ba485a1e1fe7037a3a4937a6370b1a2842bdaedc531ae20d8bb2460
z893bfec07645610d1be3be9d454f735d0a8e080a2d6cc73b0b912681c17bf87b2584d2ef9be900
z0746f46e0130cc742f6a032ca08960ef811e3552a38ba05282b875c979d1a93d1ce69c189764ca
zc8e286a0d61fb4a395d50d51a9279b9766bdd1cc39f9e83ca3206323c4958ea6a4b37dffa12603
z2fb1ed5388a187556aecd8205952701b9f2c8d4f7e9a041881d7ef57428ed4a27ed15caa2c40c4
z9dc9594c5c052b7713731b6c69f2175f9d972806df12584608e4c190259c44bb87f27fae1c79ec
z89f4c20fbd3b8599239ab4ef7f937971f2317ed2173feef3424ad8bf60deb59c823689356ed2ce
z0accd04dcaf2ff7b58732d54c4974da28122051460534296f94f7a1b416f819b891c6359ef31b1
z131634c17b9532a199455c4ef61593ca5405d5389e8b523cc96fd9ab34acf1eed0bb613fd48005
zc6b7a22cfe0843e21b97d0947dfff18aab5951653c9217b2dc0fa52ac822afbf5bbb4ca8e4d5fe
zc55b2f61a1b9b8428749d2e32ccac194a9063bac963873e4ec0747495e3f3d3db57ef453f98c62
zbd2b62bea509122c1e624d776c1d482a95e65ecdd61ecd0d971e73b337364874ed954bef0bc47e
z20228bbde9e2fbd6fb4d8878611ad30a3edb0f2b53deadd43e8993d6659c1151314e685b70f282
zfff6bcd0a611f8ddefdfe737300a70d48e2f6cc3575e39c1abe4e07710981284b4b0577fa7a3a1
zc5239226c26d86b0e5cca243c037353a8f68c9302d0e33d2f4c966072a6957e410ebc7ccbb46d6
z6641c72e6051f0c110f564095adf54ae40b00901ab548800c5e03db7b5558505b3feebb7705601
z7be39e515e4f4db3a14484a0a7346591fed2387120ffc13f54b9313bec5bb90f43c94d00d9b02c
z84d7f0db6db7683dcc48c2b5a9b53b0d439f9a0d0228bbbcf21007cf0a90afc058cdbdd4377ea6
z675840c855ad6f60fc392f701db03ee16976975ac418d84e43631244c6ff2dfe727003cc1e00b3
zb8eacf5f53f64a271e499a90ea3fcdebac9b47d15ebc590175ed8b460cda802c309d74cf2eee56
zf04c27e4ecf13e7d43c484c10cba8e80a5f0284b8020c8724fcabcb02cdd59d8b8f949e1924116
z074b80ec6fdf65d87cd52d86b91b871e13cc797619de2c22aae2d88d1cf3e50b5e265c492dcf05
z060402e29b2c6c0f798c297f8141f65bbf4a8fe87d5bce52eb40868beb2f75c723cd570ff7bda7
z0e87b065cc6379a80a2925b8835325bf0ecc74501762644a0285dfbe2e1f6a7d6b6e0e3dd9fb74
z7f80f3a3923d1389bbd2d60158dc1f2759709d60bcf973045c699e530f9fb75cffb41e82be0d91
z0dd7dafc65c2ec1ca5416213f91b21a38cdf813c51abfa576a412e4aa83f41ccafef03fefbd60b
za5939eb1ca8d6876ab5d04e7b975287c229321830256ebd45014bb3086e480110e8f90d5d416f2
zef08b81484910bf5f38e54dd7f3b045387e05d140b18f1c3bd19f10575fb0d8d41bc24769fea85
z210d0453d656c4480d0050c954fa795b1ded479af868c01f5822e3a7a154aff482f1dfd8091f81
zcb22037da92565b74841503fcc6dd605f92d470ba8009d12473548a53ffc9dacb6cb6908fb0ad2
zee0dd502a2e0e8b049359bc287e9d1b7bdc8bab57114ee3157b9c6ddff9df9437dbd4b4f57d55c
zfac0552de405fe899c1ca895271c9e0c19e73f5400272395f8b01ea028ba38d7f5abbcbacbc33b
z698791153199735857fcc4a6fb873321415cadf41e574af6a89b0120a11cd9a91234a702c67145
z51262523da58cd5cd0d2a139ead35ec45161879ae9b57059b67df53a290c92258cd2def9a9df40
zf5239c984fe4983a97c1b1b59026e9f73bffc89f502f57d6c4a831799a1e3935e8b97af289e7c6
z3685d52941d54e6a3d8965e5b74556db0b0e503f702bf678db3f02482717c7abcd828367f0723b
z3d132fdbc04cc0f7efb82af157f7b15cf59f15d609c08fb1ada52db644a52a0332fbbc6dc4ec93
ze0150fa652262fe824e2870da91c578203467e0dd855279699e52ac0bfb4bca0aa7c29c656ccff
zc6394e2f36c05f017502355c4a3798dffa24c26f560703c91cf283affa6f92993af52fb324c0fb
z717ced26c1d6a58a1540898abd0fa7339c2948b30ee84742f7bdb6abcb637b2595aa8374c34e63
z8e8753dadc4b6be6bd9bc43d95fb548440e55b8336aabf19ad4d3c5a0515573fd8cbe73aad2119
z1d2425e6b078a1c9a1645bce3601e1733b5c75346dc0ff87137ca98e9851e7c2f124bc9d013b08
zc0c1239f54abacbbdbc9f3e5a1b3266783cf584db96fa19aa4b549e978e2cfbbf3b60082b70141
ze64fd94f9796a538263cbd03c3c4960b1ca9cbfe86642960f0997b7b7286e55384fdcef53e9593
z7691ae703476c705fd1f0ddf10b1a151ba629b84e045bab86a22c25f136b9fe369a034185e20e4
zfd122b32ef41ea668def3734359f684ad9da6fd5e635631b40a8493567f8baf5a2b17f9b925942
zcb9b22c5e7e0b965594dd4ce1843de2b54840dd0ad28bfe5f560f77754e54689072314103ef91c
ze2286337e9dd364ae31d24f7ff780147a79b0914252166fff5b0581afd3982214b1bf4a2ab0687
zef745fd06fd99a1aafbd8536aacc53dd4be1c283065d810b4d22cb316e7801582023cfefbfb7db
ze1867b55caa30eccc642e8c998c9707957912d0a03070c7c14f1c9f15bf1b49bbc8161d4865fa1
z87acb3a0645c342dc52ff248eb7268f94dffa37dd730bccd4934920104f98e0b5e7f040955d11c
z18f6aeb2b48b5647c823bb49fe66b089cfa6c88731cbb35e417376ee05ef29a6d6cc821a632bfd
z5413c92c5adfb1d52942c83965d583fcd5621a1db25da5ba2d0ceb16a1ebb174cec2d34eff39b6
z692f0ff242edeb122dc7a0bf66a790e20d81f061c5c3e468eeded99580a21c633874ac1d20ceee
zd33812f280e3bcf7a1dac1d102879baca979571c398d574dc09d2fac5064482c0bcdb6fcc8029b
z2df5266fa582d33c952bef1b4a66df4b06947fbaed1b0007359fc376f7b7e7104b63046426d230
ze8467e4c720b8b992f9df46caa795246cfcc955ff65a7c7d6087fe4799e39c4c145f1160bb4996
z7ea8cc6a8afd2e1743df730f6eca0dfa1c46e4575eb5c4ed15b37f5742ff386bf0408ca8a14a21
ze96ff7bc6b232d49fe9e2748e8e6e774ea9115fb593c8dd0918ae09c6f2e5b000139e763be8937
z3c2500400286d783f546456c04ed8de097bd08d2e9a5a187617f46c105ce8b9a22c3cbf7378971
zecaf7dd20973689e2191a585cede0357acf0a6198a39e9cbc1ad46324866a90e95118c569f88f0
z6ebaa78944bedb871810373f36622677ff7f919bbcc6b596d54a2b754dc2ce881c05b4f9a5f007
zc027d629ca4236388b0c47cf15e8db9f399bdfc797b69a3cc2ef5984816e4c36de9d5672d22755
z72975ded7ecd47c36fb1906f771bc79f53c6438cfefc16e74d99c7b18ee0223cad28e6bb1fd3b0
zb3cd2f1d3d4c4884f78f5a75a12c3a3931be0c46e180a1ede5df04d5ec0498cd5c91e364578090
z912177258a8a2b6d5becbd488860edf8c4c4685bd339f303948206de4c51293b363454afcd05b6
z5e5bf11c63a4387394d074daff109574418fe4648dfe15866c535008afd7a933f100fc5e8ef755
z3bcdb2348b46855a8397e7d674539ce33b8dad29356cf5c1622ba18b983f30655f18d47b9020a2
z0818fcc62555697fdb9ce114515da031647244f23ef18236af3369bc899a2cbf9ef048971ae6e6
z6fb673600641095dd231a6f8ca781d4671f69feeda94fba3031e85bda518875946681d355e1353
z384e8c874699f5a02a9891c422290bc191a226f54ef79ef067b184f00fe5c88daa4b55ed942101
z94db0692b8a98d88ca93fe1bc1c80391130a6b56b2d5a81dfa813f94c035a81fe4b6a3504de865
zece266a4d7ca10b1a7bb0881c12226d4299ed38e640cb8faf9621b21b2a4d2e8f652f6d26c0e7c
z820c57664b3494475d3f7bb051a21333a50f5704cd9f9adc2f7d517320181d40ba55bc0a730c6c
z0488d4726ecf9788cd4fbb936123b6c1db60e65b436c7a1add47f8fe00247e36383d5b0f622f0f
zeaf15a97f092ffd10f9bb29da6eb1294deeb0cfe135ebcf2fb005167ebc767f61761114e0b07ce
z384884f2f2c5a7c0837507130f866a4e4d8e55cab7eb64785fc9e3d3e9d74b20379e8ad90a2d6e
z349374721611a3cbf6e053958d81d0c8f18e8b25b343d07a5838e664f76093d41ba5030b435d53
za146458c3228784710cb2bc8348b09091a783e85856adb3a6ed7820c99ac82ace242d8e5f848fc
z8c1e4a629840e64d6d541812f64ea6166bbcdfbbcfc2d2d626c47080e2f22ab1c38840b8415fb4
z4404e17cefc5b810c6895223064af91999955ab8aa6a1889029fce150af19f496cc62a76eeae9d
z046a11026ad9be6b93269689cd672f457808f5c3567b7cfa89352a705b98167069a27e5c579116
zf5c8d7ad45b020f0829756676e77bb804952be45a10e17b1d56f9c2fe5377f559568aec8a93970
z6dbf1a23c6081b23a704b49718d94ac7c3656299d1d7b314d1aba3834327dcb8168b54e176d715
z4b2e7236790af5aea624829a09f96c5b92f8c1437ba25e92aeaaf578d23f6fdf006dd71f7f42c5
zf1f079c3d7e9201d823a48a89a1b043d9b9251e44aaf0698eaaf0d8513c9333a6bd6f6cf86256f
zd77007d31204f0f6f9b84989f95b98fde166df74dad8acd97c6eee3538def8f97d18f7ff51c9da
z10d17d6e8a1bfbae02b4446909a002f33480235700ca5258ddf4ca745008a0a9534be5307b059c
zb2795d1ce65526afdd61f6ce313b2168696a5c43a98971bac5a808d405dcd8d7672f10b3eb1d41
ze42634d892190857a00da307bfc86ca5ce1c40e514bd41992fbd0c76b6d193e2f087c17e84292e
z4ac1e9b3c2ad8677d44b37dc452d3414f7b495575b98e99965606bcc975300b0ecda307515d437
zb2e3fcd11bb94b2cf8f7eab8077c968d9ac163e3c98bac677493c78aa7b241affcb03522cd13b9
zec10845eeac016d046b4fc7c5239485e6fb11b5df38a1af8c738465add2024010baa6b17998d77
zcc463d1fdbdabe069a60ff95a6ed36ee917a08915bdc8e8875fac36c49bd07846d606991050062
za0423d122e88f0732536c310d38d86b30199d7db7306932e75b0f4136dddea5cc835e620084585
z4e3cd6d66620cc7640f7a8502cbf41726148780bb47173c957b532eb680ce9389b69c0c6bee5c8
za741f93a306b6f33ba94282ebdd3595884464974f9a52b0c82c2f73d1eb757bbf0a69848ce18c2
zfc7d24a59af339c7e5b616df210dbe579bf19d3c8fc7a9365fa6d8739985db140dc86d51d4cfd3
ze5b713cb0ff39defe3b781fd96545c1b558ee9045bf062bbbc48397897efb2955e9a33b925c646
zfd9445c1ea5768f4d67716a77904f5071fb6d2247620a8611cdf069cd5aa21bfb72584f74d10fd
za2c85be475411d275f560a64f7c098342772148fe05fb2d664ea6c414a1dad948c87b59c133a66
z744b9fea874ec438af3e9c084f7b6df50f15bfe9164f20bce9b7904c567359ed8bf0377c1af38f
z365bcf88f28d22028431c899cf1041f0cddc6f21bc44e20df1e8e30f67b3d6c2cb95df064ecb0b
z141dabfa09ca9a91b0ca2dae0388ad87672f718741d5030fd1cd901bd9adea5d6d93f4d2646f70
z0a9f183f773d115b9c9f45970ec44b8b6157f952dff473cf29593b13b7c6002fb175eb7ba5bf27
zae54069ce003f419bb079ae55fb0e16edf3f694b93dfffabc1ce8b214a9f60004720cfdc902eb4
z2b2c60b46f09af127999ae20d3dc761a5be439974110bc1e4bc5c819c51b096bf73c5342c75dd4
z129829877cb87a2e3b14538d8c6ec3b55c5afa6f35cb5a5ffc26c658bac8a887ec51228f7b54a1
z6bafccbc670f632ceaaa8619a66e195346bba03e8b8acea4af7bb2c04aaf93a23419dec4d54e3a
zb33537dbc3ebc6a1caac08e10928f557578d220bc3360eec82b0aeef4e525eeb1a08005882ed96
z5ff5e7c22d3a9db36e540490faf1ac271ad139f8ad777854ada55a7e1bce03aa03d588c334e492
z7c81dcaf5b46c3ee55010a835da4fc5b2b032e6efe46ca4c5875ebc467a0d67d8c83009ef35dbd
zdce6f15a9b4abd524bce8999a821260eb681df916ad992ed88a693fd592405cd14742292f44be9
z846bcc25f118d0fbd790ded849dcce4f8d04ba2c9884ca252ca4425472f93e444d18899cb86b97
z396dc79f575b6d9c78d4d6d88f275f1788bcf564961bb7cce7c29b13eafd6f5be7ede0590336d4
z3ca2c5d9b73feaae16c34e7a6c33095a8071f469fd174755098243ae6b71ef30b08456c4e880b2
z04e518f23a0bb6a0108d1a83ac13998705000b5c50bcec5113b4259d8b562d821364a22bbadf0f
z98260e7c69d5b7f4ca3331da7339216ac9c08daea9a39828b0bf1a5466065778b4ad1e59c00601
z642973d0a2aa5afb03b31f93a36b4b5c016e9d4f287d1e9f7afb3c764965b0110a9f681c7bbee0
z0ad4eba308a77529340d2669c9f722dfedb780e15d3d781ed42444b6bc3518557aad4a3d6dbd7b
z8bc09c0d278de51e0d8b630d519a924e83b75976bfd814bae52e5f88fa2c52bb42842bc82cbfe1
zf98b322a3b1ab7f3125b7eddc3422f450e0e39a13dfb46f6a19a76bea970c6e28263feb04f962e
zb82c05fb6785f2421d87b8ab8408bf75afac4d9c450c10954b2fa25a2083fdcbaa013d54d82cd3
z2649fe54abc9d0cc0e5d515e52188350e1dfdcfa97d83ef60231e0fcaade55d182cf8537bb374c
z4cee12d1efdaf09828e44a8acfb999fbde21dc6311cf7807183c707ae80c918cedc63c5845b999
zba2f178de4f11494fae854ab47fd388fff2a755aad4d367d0e6d3a31751a20c7b9ddde5e455ef5
z584248a1174f899b7ed988c04d4fed666987f47267b0c77261a33a80ce8a96f2570ac0d4065ddd
ze9228b9e254f44d5b7e3f1b10d267d6fb87f7f36f6f082def61e64c36d05db5b7da503a469acf9
z592a6f769ec3a5900020b4873a45f58c7dcc33f06bd780810c6b98bec0490bb392db531ed77d8f
zaf5bcb768d4b46a6c33c37f8cfbc4a7538f8d6d5a7c8f15ede7b75d5e62deced53045a3afdac7b
za5d5da02ec14ee887a5f248e6bf8750a7829994a59cf3e17d65cf8400545141375422d95ea9c68
zb17488aa5bff7136d032866d5552b15c33e4d3bbf42dee0348f97f369c6a7d68fe26915f31fc88
z381c65e6c331bdb35b7d1932716486e1d53e7c3f287eddf09d1bef8505e4cbe369a7a1ac4c4830
z50896a26fe8ff65a366636d1eba828e94347bd2b788a7b3b3ba65120bcb111c190df153fa53172
zdfb572fe2d93debeb457ad45e3a45ba528f42f8083935861a2e0a60a5d245356c0efbc61a78742
z6224e44234197218fa7c410831f9a6d3995871e30c3da98d21c6bb51c491c1ea4ce0a5fc02de13
z26069537096f323a7667a8263f2a3aa9ada8ac7de16f3e28fd001aa1fec5b41c60fad1fc440306
zf1abc62e6da7302e2004e8e96bd369ccf66d344b24296dda3238ba6c1963a264627eb7526060f0
z0e481d2d719dc7713a1a6ea4902ae354466c19dd795604eec54d1fdea88fb0da6f1fb8d643af0d
zd3f93c9d280b916c5cfba618db57f19d7d4ef12ee08930118e0ac6570f3a818322b11aea161d18
z02667732eb6d68c7be971a9b8078772bb7ea3f301ff28f942c9aefb6dd6bd9011974c16eb3af49
zb3b1727aecb4f57b026dad20e0bb0750b2eeee446849362e594b0d11261eddb12bff49f13ccf7f
z2e9cc67199b603d086e8ff89ea70ffcf0e4fdff4b88cd18fe68252126c70ae70e9c565bc3c1606
zba0f05fa5bb314d8c295271d893153596411f617cf4fc88c8ec867cd385f015d0427cf1060aae0
zcf1f2b816f45548b990119c6b11f8fd5cca18d74a5ab7f61eb9426d32658c66d1418f275ef7e11
z8f216dfe6f9c12cc2d5c83cab047df9e1571bd4bcf62c1750f3582c7edef05b87ac3a720495815
zb89435f70919a53c16fd0cbb4c3d54305c4dfe9c631b7affbef9b8d2121f6ba5acace80e3e9dee
z154b90af384f13c41fcffb4a7b1fdd7c43bbbb0d7d3a73129b9ff3b41a781741562e3aeb5a8dbc
z00234108dcbc3eb3e17468784ceb1a7c02803f44052a2bdb95ace72ced3a1cad63f89bf09993a8
z1cc66376849d2b274121ddb4737a46ab6d5b4e878f941fca37d8c4cf2b021dc4e15a0f81fc461c
z27d5e78a4ba894682de5c740da1a941b33d8c04a32b32e40ffd1d52ac2b4653e724376d37ba664
z64ebfab1806911f82b22f5eeeaa66ee4c11ff62f0af3adb5a470deaa2faaf51ceeeb1d6a5b2d6e
zfc54411b4e5bdbf91b9648afd18fb06b42260d26dda1ce327e8a71308e71af1e4d0dbe65147760
z56ae2ae06560fb86e8d1e01556d2bdb0491aafe0ab66b82dec6880f34210bd8e341953b1ce8fff
z4414aaa2ccb396895684da5d11072d8231d133aa4cb8f45fc89bfc3e74b2cc987715dbf9ffaf04
ze05514465545279b3ad45bedb2070bb491254752bb0e24574da4233d8ffafa80bf494f2c471eee
z5e1dacd5074a23a7a345cd17a4cc574881c2d66b5cb3fe4c69dfb5e2e43aeca68c3c17775fb843
z5d5313044f824ecc2ceed4207babadbdb76fdf50b7edb8a08b096eec9d691e0d06c15fa14c182a
z87e457ed2fc1701f214e82755f0d5b02fa8f166ccbf2d9a570f319802926b53246a501ae5fab92
za8b370b0371b32485f5e55f21023717c62d0f1164638f121e0dad8c5a95f63d207e3f79c2a044f
z7f7e54b9b32fe99cf5900e688f3ed18d71e2c5ec322352cfe96f14763f7858aeb6cf532e46f6e4
zba918d0296e6ac5d7d3bc4f8951cb9355434ef36ab7f26ae56268c049459f2a83b7aa9eae8afa1
zda35dd7f558f83865102249221e302c3735238d1d47370447207d784b5f8ab327dbe6ed068e5f9
zfc10ee40ac0eaf1bce660d5c652433e10c25ee0bef3ffe0dcc599d6e0c97deafc3ea72637bcceb
zc47d18af8d8daf0bfcdc53a4c5b40f9f87bffc3fd46c9cb50a252d84ac8f216944b3e4e5dbd6e4
zb55f3ec6fe29d545fad70ed251d7321be5781df8be9eae6908cb5e60594e26b3f5e4e8ab419821
z79255a8885c36cb0b94bb82f03f855376cfa264103afd4f633f82e7e4f510438472e080536c76a
z82501a9c3fd5f5abaeef033a47508439562abc771c44b06127a254c050b0c9e3c44c222182004b
z33624cffbc707a56823142012ec2703332365011a4f8277175b346c8d45c2181327070e9ff580b
ze26ad24ba38795227e20562b26e22d5550ae59616d81031315629de40a0c5f6cc9cf296ff52aad
z6e9ef6e58a5cd8ec04bba9a5e4eb21f4c2826f87cbf41d4a2a0aeafdf624f0d9bdbcf09f5ce96f
z8b6e8d42aca745466d20496749ed6a94a633a70ff261a8005c78dcd5ff56c55ab7c1ca0774e18e
ze74d2b98a60a77b6cf3b5f1c54c07050726b0fe4307df2f09d1610bc775f8c6421050cc314337f
zcdac43551820b6d1f454feef55370ffbe63220e74f5d0fc7111eb4272a2cf982ba12306d52d485
z0e4752fecd8903d0c412f01dca708a05b5ad447e08641beafdb68513c486885b2433ff50c533f1
z19f09ed132a94713b08d17663391022ed98cdbadf9fbc28556d2638e60fb8af81c24176cc7927b
z5444a3ee3461d898d5a26bc7ed39a5e593e4e80f97208c1608de9bf966d0772f17a2807ca0f4e6
zf9912b77bdccb2b003f5309205cec127c13459fe03721944088dd090e49213b3a7814cd1c0ea1c
zd9f7f88ea26ad794e2bdc6678975639a1b357d1713e29028c7127348d2f84bd5d0957f8c5384c3
z99b01b850995f6c03ed27dd775ff5767a917f88e8a0b0c3c8fc4355f1628771fe5ab2f0aa4c252
zb47fdc1e8ec853a259dae8db9118b74a3bc52f0a0d84f9271784e645daf82d8ad666a869fb3141
z1e114fba608e949c8007d24512360c737ff3e484410c67fa3f79433fd944dab153d744878a2249
za45ece62afab98c92547df53199e86328745d30cd02d3cf4ccb8c533c11bfa2c86c5e43e60f994
zc2c50d64804bb99d885a4af1d058ba3f404af051927fb9885a73cd3182a233c17e96859d970d33
z809bb0109407c61ff5ea212cd734352a8759602b1562f0c16ba22cec24b977b90569a2c8949d1c
z6f7cfdcf37cb4ea2fde1eeb567da606900bdbf2bfc15b192118f07d4fc2a41810e566f28ec25dd
ze1f9fe2c6035beb605df81d9f22cab0e3a654a93e1b8b1f0a8a2216c385f77cb63da557bdba08b
z5b936302a04834638043ebbbe8f1323ad4bb4789cfb2acf3ae84b7fe16c129580188ef943cdf33
z591d2f6fde8f1aebca43b9a307b5cf71d73b609c76964d4154b89a1177a9f603f28e668ab6d666
z79d7c73e60e5634bbc60265a853ee54304b42cdafab0a645173707dd32cac4a002430e401a7aa6
z3fe373a7cc9970cecfd16d9cedb0a0aba1b2e7091101237ed4c04271e8c75fb64e32efa28eafde
z5d8b433c98ef3e1eed200b4e164d83caf5e145c46d233bcd03218b59d4658e3548bdfe27faec48
z1a7b833c6f3dea7d0f9f2a99dbc0b034b54ddbfcb38a56cef7423d6e48fb7758897d2fccaeb4d5
ze0e94f0da03f8771bcbafa3c64a4785df31be8e6591aacd65528111d6c1e992856a9f5dcfed157
z491a254d8186142ac1c0d863da12e1d8528ba3265c57411ebe89be3a447d5e52111207f403dc2c
z7c240fa68590ab0674c7d328e703e0b8b3cb2acba5a7384c953b1e9ac662ebf9be088fd4f7c213
z1426dd19dc32813e4fe814b0fe7a65f6957e276cded1043b0621c0fec1de00786b1b1337edba79
ze60d3e1bc5ccea5dc479f94bc039a61b683d4d6a27d294f312b7f1f6703e71173d956fc7bdae30
z85a8eb53758308a45628e8367471d19ae618bde75365d6e4d73972bc0f2cf2f1407d11a1eceaa9
z4dc0136eb53eb43f735c01112a1801ffd018c90efdb9238ba50fcd0f56060e8f768e8766f6199c
z14b07f865193b849c71fe111ac02e727a404fcb92c90aa7cce3e3b459d4610fba10505425e02ae
zaaecbbe3a6b7841fed2e64ba6c335259c4a83357e35e0b12cc8ef455b984aed6015aac8db1ad29
ze690de3a29dda0
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_outstanding_id_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
