`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd318151217f11a0cddd946f7445050ecf57548e2aacae67432edc
z32627b1419acc732a30d902bc5f9bcfb47b2bb5b50a3a8f00cfba181ec0e0a57e1931059d0cb41
z6c3bf461d9862ce89aefcbebd983e9d61c301834fc52bfcad8d8671163e81057510f91f873bead
z999075def9c70301f71cf82ce8c57a46078af24b8b1bc7cb5b2e32e72968dbbf2b18bfff88ea60
zed5018a743e6da26ea4d593b105e7551f53c241f3e6fdc37471d9b7053cad8414a68630b379310
z3a0f725d61dfcaa35bd27b24d39163b4f66974056008423363e87ca6e89b4657953b18c51b97c7
z153bfb0faaea0cd5ebfaca7d287bfe6f60f298e363935d13e53f4efb7a3edbb6ea1b5f3bed79bf
z603a7c780c484183d4daa318d5d5b26d1ba95cbd5554e4889750ec2fc95c412902bfba464ddb4d
z573e5e78d62a8f78d8142e798fd2ace98e86d9ee0f1ad9f36931b49f0bf0704ca4e8db7e56a115
z5486877a7ea22549e9b92022fe5fc9fec146c94da84031f94a9c21ab94c0bcbd238ee12652a53c
z3764d7741318e0e9ca76b7f16b1318b5dfc6df1c0330c1da02fde41cbe320c015570eedc86b10c
z1bbed264ce5dbfbf5c8a20e7ab805245e60032019e3cef24769ce94646c6f06cb0465eb46cee4d
zd1fead29686a4094ae93a9864912d0ddf9a99b3c97fb189e07bc54804dc98519e5ec41b8af9298
za648c331cd2cd1deab3c6d915e3a77476a74c5909b0a2f46086abc032d95eaec4ecfe77bb13fd5
z023b98e39f74b0ef9fd159f1cfef74ad46c16fdf68c57a316a85c2ccaa57092540912d9185e345
z62473b1d4c74b02bdf1b5a88b5c0df9bbee913afcbdc05949a5f26dc8c48a707778e13d46fcb33
z92dac81eba9467da85236a846a36b0eb4944e2335e2206cbc78f7fd207479822947915a2316794
zba59f9f50e12cc4ad2e1ec50531a791396862eb367d56cdad7879850f6054735a24cd9c5b597f9
z6792acddefa14410df808134433ee1582430923a21d2264b2308c109749024ba3cddecf2cab189
z3cdc590a420e1fdc2b4b3b2159769acae9ffd25e0ac44dface5ea892b336a2d76c7bc7a22fb2df
z7e8b4a67638f565830cf61958d1a27de654bfdb6dd8a4758d08119f193d13192f28da11d1264fe
z687112786a4a5690e5921686018bd835f99d26515369451c7c05df092329160c89b3c8b9cbd226
z9088518a92d61e37ba6a7127129d639efab41dcb64e09df2a3789e1abf07282df9815214cfe214
za5f910af9012bfbf17acbb108f6ee56e11ac8d011361218d61fc22a5c7761d79deee1e99817b20
zd9f55487abdebdaf60b9e10ca70b75dbdf625204b8bede2602a0cc92cdabd899b06aab2585d39f
za7bd50ce8146b25d0031c32a77e1db3714827e3992f911aabf5e8f92e0581df86d84ae2ec96664
z42a1df5f26e845b35a8e73a0adf1b8e7e4bec154851b06fd0e13b2a2d35828247492bc88afd02b
z20dd32cd6abcab30f480ef095b65465fd3866ffef918723e2ec809f71f271e1e5608979b9004f0
z8587f1df2e0ca1a3355cef8920e978cd9b9bd1529be0adde1a6e287753ce9939f82f32d0b5cd93
z394b61a832ab7e6baf55b81e17566a64e5c3b151ac215bb108d515e649f2f95fae724fddb585e2
z3f4d95be73cde0a21585f42b635eedaf5f9f02dce3561e7ade624731f4e31f4eca6ab1129d131e
z72d02f73d56869189dda1884e784dff9c1dd54999712ab95c9753580e204541332d418ee16d30f
z924748df5304749beb15c1e6c7fbb23c4c548ef5bae4c8d9d213791d0afa8bfbdb8b6264e732f8
zc535e3358a80b1568634b5ae0d301878d81531b89150858e6186c700bc3a49054e3addc6fd0823
z827ef8c75da0fbb1b0a1518d03b096fa1080136f544b3c64c86b7075d8df60b423bad2c4e9615a
zb745bb23c772e075ca8494613ec14e188daedc7cd7e329ac229dd017523fe3c4d2c788e5337520
zce9aebab7001b9de43aa2d3b3783c00959235fe10b7ea182040317024940e139735de2d22516fb
z5cb6c47fbe11d37407a0c196cc4e52b3a5b648704e47856f95c5bdddd062dbf916b80d734005d5
zce01c6c6f578e61ed8eb6a8dd6c03306153306ba36df616ea8f46a41bc251372179d82a896b534
zaf88c1df49a04d944bb8d780b899c1d79a87ccb518bee6677c41459606e97d5c3ed56104438e3d
z584434a514fcae93aee0ea8bfdfded6715df2a98b16f726fd6f04748a126761694a6e2212c40ae
z45af644f74d519b74930a2b60f8c6337eeb78f95ee82bebf4c1c82ef0c218ee1823b10b118a9c1
zceec39b43520ea844f6ed59e5c774d4132adfaf309289da70d72521f493c89308f84525701cb13
z25a1613548393f04511e6f80c78834fd7a28289ea59551e5fabd0b2be14292219d0c712a1c5ac7
z1bb8005f989fc821a311f478e7b321d4b52c4532d29e439ae37e3c0620f372e958e33892323ed5
z63cf9e13b7555de5ec4a32fee8ccf64758315524bff31923ad94d406c1949fb1e50402cf2e9e55
zcdf02336b76a62975086cf4b41cd3f847b326968c968853ca4c7c3a6d3f9aa7acb43eaeb38f43d
z36174a5ea180012351fb7609bbf82d352152f935c7ea4fbe4524770386939cbf53081192381b4f
z2cc37c1f883e172666e735f225911c4b8f6c060656aa1990462f2cb16fc134ace028869c4199af
zfe5b34ba502bef74f59553719e5447985988f3dc11afb732367d359fcb8dc1d929520a210c1b74
z61b43536d8a63646f3402eb9941094282f2ef16d158604b1c9ecf835743b8f2f5cf017c1538219
ze15e4765b5cbfc910be3a50d77d4ba7e6a0b94a20c0ddd1196ff69b1a0e9cc9f85c9b395aedfca
z3050ff68585e1da092c79e3f76b9db5b7c82344e99802fcd003869fdf267c0909da00b7795c05c
zf08f43272bd1867ff20f591f770f0a9da5e13e3eec91247c97217c2a38badab187ad30aa00458a
z6556c714476f59029537933a2056002a2966830b8bb3997fde6e04a1685661d3f93b4dad395e15
z8affb81a8b96373592ba891ce294c5fd58fea35434a8301570e7249aaa0f7604007d430d714ab3
z32c10873e61f42b2dc2c746220aea8b5cc33a548774935782e2c87c304f3ff2d0728dd48dcfdba
z5f0fba628f2e2566c97b63ca3917d208bd41c13af4eed5742dad1797a1533bad0e2c827f0b4597
z4620f8ecc8f3557432b43db31320b9e57c18bd20b0f1e85f1c2099c439c38be6928abf810ef73b
z23f4d09a4b5933d398f4ca93a61d2669a883f55aa465a78573746b44dad495e461efbf9d3c2e50
z4f1179d98b866310826e0ce38748b8e4922f3b4739cd2dfee4ae765d97f293beaf821227f2748c
za92a4a413e96378ad5c7177b6d14f89d6c02dfa20cb257bda7dd08467d23d9fe2d007da3f2fabb
z04a04eaa5b6b0212d04a2cb3b121e468059b8f6fe061364a07a54a8df7ba45cf32aaa3dc7c16c7
zed48c84c0328f51d0389f9cff8b4ec074de437db89dd5f718ad9da06e874971226842964f1a28a
zd9df8dbc682636e5565cf3cd6579c235f62ec77622bf6565178e87c51885c783314e465772b174
z1132c78654e4b2c1a2606a0f4e61667ddc2bdf34eb12c903b708a2d9d38a840e140f7f2b08360b
zea8ea8715ac084215ac10a178b9f7db4b3a7f559e6624cf4b553594cc16c2068810119d61ee3bb
z8b403da89db75ab3bf2c1206cb69ed7b0a0432ada25b6ad5568d56a91239977dd353f00645bad3
z72ea436c78cce1b53b8c9aa176723a4edd78974d6cbc46eaaf46c8ed23fbab3cb8342e265bf0a2
zc8c322c9a4b5fcbff0bd5042fbe5ad0328bb723ed2b3044bfa17688cd91dc015c8e47f0a33fc95
z5be8e54a59cffab6bf1975d14722f975a1d64e0603a1cd0575562fce503e19cc100a206d479c46
z94e65f2cf59b80e9d8f7b58bcaa70fb6537252e7cbdc07195418500a26b900ec7e5b2cb6ced859
z908dc882bf0c381b9b534478cb5b66db35b649d1dede1ff94b54bda16e781b73f0ba1b5825e4a5
zaebb4b85ce004064eea100d6f004596b74a6e39cf02c0baf190b5395469d1215ef5a06cc35a500
z523b8ad150a49084806ef9546fdd5c8ad0df5cfc0d171677b33c9e9a0daaeefa2641b98ca995e7
z41da5548052d517c1f03157b688d096fc22b40cdaaf4837d143418aae0063bd67da8d5285886e1
z370492d29cf9a63fb600a7eeb5947ea6fe7a5ad30c70f25e6563b25857bb5b4ea5d3d3ad0cd868
z988f61afb5eea96fe714109efd55c2052b43d827f74d2e381e45b5b9a67430bc3a2d1483fdc95d
z9d5fa14c49694cf92c29a54074717573a03cd1d086dcadd0a544802a92b52985737826dfe0f2ba
zb90176e7150de13d7f36834dc605c657d23b84b79c8445d37b3e977ae3cfd91091cec66f409a0b
zc4e3046fce09d87e20e99c9f020daf77c7d6223b8f29a6874ef8b4de6876e98661f7f99c8be18f
zafbf8c349a07cbd63376c0ef6635393df0bac835c121843676ab8468f8900a66a0c5622159d0a9
z1446afdcc2e0432f6059ebcf5b2ca5005474a27ec4beb0d4098b767ea69de177eaf51f6ad12d68
z37e99397cd7f8a893f59a08b7f9237905d3914b6b5a3a9573a70ecf6e3d17df2c90da0253c25f6
z9f63a616126d08489bb5678f0fac6d980a5622a87955bc6db78354d80340ec1ea21940ba23ea0a
zec9938b104513b87219231f8bc08574c6669edcf7fe29dbc23c2e4685e8c68b6d6d75de9d7ae8e
zb209437fcca7673ee7fbdf30aa591d717cc7f99199e0a56f37062aac44478c92f9be14e63e89ef
za8e6f2dd2eb0cf3304a6ded6ce66649ec396fef6cda0e144149db5fd538c92e3b7d1b5e17c8a53
z28a333af8af248e7cdc23d24615ac047bb5ffbe8ffff3edaf84fac480c927f2da57d72bca6f1e8
z5e58a98dfbda768558798a0bfd97cd906485601382aac40e7b619fc72dc0deb5efe240b4d93199
z4ab8006704c90064b1983b07b78367fdc97cf073e536ba4b9ec557a79da1fac8375fa21fcacba5
zf8dd1ed06dcec6ccbe9f66069aae7026363114cd60bddd0093c8a7045afed7f504a24efcdcedf6
z589dfed4438a290edf03efe4f774ccfb73521ec902ea31add624c2ce6802a1258230900be7340a
zc89383f3b9bee13218c5673f32fd50e94a0611f5bf14e92508477c470c2c6f5d7656dc854570bb
zf4d4ab5fb5c15cad9cffac5189db061bc641a52c4d1e99007897671584f750cf22c49c0f93a264
z46085e0a3e09936f68b5506b3c10cc4a5fa1d3158426745927fab4a794e76c93c8aa297356a437
z2b60a39b986c443ce10a6747d9609975973e138a57577c95867600359e7d129043efa7d12498c6
z7ebd0dc3b12749a9cac620c030aaca64ca0c867de61c961f593785df322b53dc5846831058b2fb
z5ff18a4dcf205534a11100ca0ec72d983f375c07f8bb15930cc008b8ecbd456c4b1c94232b631a
zb7f53fbdb1ef940d9471d18c557b7504a382d3f6b86a04dbf49ec7f9216790fee29bfe7654f4de
z865cc4e764ca0e9f4d457aafa1550a0e6d6235cd99bb611fb38a796168507a9d2f6297f7f01b8f
z73eee95dc5eeb058a0fa4cd5d4143c1fe16b02d9b3fee94f360a3679b1518f8d371cb797e08989
zddcc7ae19ac34ffea134b0d9170ae17018bccfa11fbb864c1cd1333276519b2d5c30b6e1749ede
z7daaafafb1b7c24bdf6079f21ed7ddd8242935945db1016496dd86be29242befcb7fc7ef937607
z005b4afdcbc193b41dde97521d2c59b93f88cfc5d26765b208c809a0bd045e404d8430e1c4dd13
zcc8c22106db2b7b197f437dc7172c47736d8b73fb4e383e464faa03b1992127c4490b56d49e9f1
zd4076f02d8893f8402177fc860c36fa4b887260ae218b5be5cf54ff06a1ba2472e79b8ccb99986
z54cad57e35f391da1a4b1662d70278435b56bf046c37523dec1a0fa104b2ee84f708c04a399692
z928c0109d3464acae4f87b2d753bc545f70341f3c61b0b790064b80faca1f684e30373a81767ae
z33d5b21c3bdcaff1292e6bbe12c3a75f25a253bbc46eb25e23579c9da93dc1e978a37d4e8d853d
z1462499e9159a8449e0fb070b04fc7fd13b698a2f619b646f1e13e122312054630d354dac27e80
z06d589e86afc78531e48de0b4e9e9bdb1ac4bf92212a70a96bffffbec71911e97ec79481a688de
zd884b25075b55a80eba9bab7108a82ceed4ef05a503436983bcf919d85981ae6763a0db94a6bce
z2f23ac95bee9ff24598b2bfb8c22b21f48aaea148fe97788b2b7df0c7b173cde7b63b0a6fe36cc
zf634944a1483963bf94fe08414165f8b91c7695626e59ea1f76de4c8167e3415ea91bea644772c
z7d8b360fe489fee02a2924a5c100b2e08ad8fb9fed03df572919aa30f42cbdaf09da7d6d7f7950
z72389891c0f290add9f5900cf5ba5987903a76bfcf7e10afedcff2bced49c0ceb37c967cbac7f3
z19d655fd5bec21e92ab91362bd7d3a6f28788dcb9ed49f5b71d0ebd3cee26d2c5a1fa2e731c6c3
z924be0f1a5f032c890ca29b25dfa518222c966c6e69f3bc9ed5023a2276b7ce5a2a9bb41916071
z6369d7f7abd30383ca49f070cc2ceccb52f527109c71535d910ec696a58b33dde84fab00b0e9c3
z6415214ef81475c984fc2e2d18d30c7057d8cd73384a979ac573673e0e41f3093137928c46d642
z397946afce1036cc3814440f694e5c55c6e8599b4beb9fbd928889a526256c73edc716467892b7
ze85028a0ac7591a496811e20866f270371aae0c06367a4ed0d2d81dad1b3485fce6d36e59c944e
z55241113cf19951fcc6858e0ac8bcaf98ac6ea4b40ac6823263e2a4d2279ba1befeed05a62da34
zc1b4de3926c22c8a31a354fe6b8eb8af8e66f83a18f21f99664512ed18e5a2c842160c5762c961
z522abe7ee39174f084467eae23e952bd1f1104919a094149480dbdd10c12e2fc2ce557ddf16836
z48df6feac6c50da5bd193883e555aff3a1bbd7707ff2e5fcf3f03ea29c1111c729e42c91acffbf
z3081e9aca8c0b5c4a2bed272783a10c69fcf3ecff921b47d03986187ade55cefcafd3b9fee78a4
z69a746202b6f737933924e893b5886974f0e4fffa53d6dae9814013d92c408b4f20722aea0d5c4
zb92ca3606b4b886d6435e42f3f6ffb92417a79f0d961ab9947f8dbc1f6631420386c06ba0491f3
z4251c05dffe0035dfeb2304fa785119146c6829ccb12198a9409ebf27a3cb2f8b67fa1b1255923
z1719f09bf9126d3baa260dbdb59d8208d0baa53521ac3eb06afe2e4b32602a1c7345417de4c033
za484a7e7d0f0687335bc08f58249f60472d77e1d779ac8a49b00d47622d139cf46999998988391
z701df4957efee7bef5931d13d2044db083c2e7c7e1d879dee28823e50efeaff723c49515a901a9
z5c765d634e9136c4fa2c4fb84b92b6e44ebed46e282c9f4677e8c1f0c7772b5d50a3e0e095827b
zd90a94b05cdcddf8f7a44d748d5cc73fd1b77c759da59ff988fd16a844090dee6d8491bb6ce86e
z3c04a1fcf2da7eae4977b710b29fef6fdbec9844c6953915eca04ecffeb5c75348ff030f3c67f6
z24036d19cb944bddc9cff723395e8eead311b53738cb3757ea7f779b3ce555b5a8103b3dedd1b1
zec2d15b7ac9e4505b12011d71cb1da98dd872249a783f683d333a0ff5d0fb03c3145146d16bbc3
z8e3ff9f572e13ab9b6f199663bdeb08d5ae123adb0a2bdc37a4cb67a9f47612d53c173cd5d6377
z291737352ef2e3285841eeea1f87061c5adb2ab55b74d32ff61a58c34943a180d1570c45b04c25
zae75b48b0964932b052c38930a7d6226627677b115aabe9255bd91e03815474ad1b6916730f2b7
zd423164a37812f6a7e4aa8584b7d1186312b4140d77f9ad876ea4068bd6609fbd6bd8e869c7d66
z0cab2c8e5312e2e94e9fe6aadeebdbbbc9fcbb73c1507140d5a15db3a26fde6083469c805ef433
zdeafa45ed49c0effdfc48a743855bd2082ee6a69c02036b0fe4d741140bb0bcec16d3a3a82ef77
z7f651d0be29a205460b858776e62312c426fabb926e13859900681784ee6bdd69771659d8ba129
z0086da72369b343f5f5e4c17f47ed68ccf979f8edbef994c901474dc93e0cec17b119fadac7eba
z26ea81a604069972c3a7ea5fbcce4dbb8fce1d66d1cc845255101cdd2fde0fe303ddead753d896
z23cb112ad272cbac23ecf621f5b03bb1c6ff1be1c70b2f583d386c70ce32653b232c93cf0d6da9
z61c1b5fd811c257b22ac27591624cfcdb70ebe2c1d7622eed5a236c7137a453f862a8ffc11e04d
z1124e5bd4e083603a4f7e12386ba9d2b5aa60738543083143ff35135523b4ce786512647174b95
zfd8653738a297bc4722a399a931aa24c39b80ea1fcd3c8a70cd591558b8d984acdd7e1d8a02c01
zea7c89264a126c2ab72526386dd749b69f1f294fa71390916220de0318d8cd95c6080b793dcb65
zfba50ac59eee418c96cc9e96e1d190e0a0f9cd73d8ce750cf2c626a6f7dd5af6336c05f0f1572f
z7b931aab48effc75a6092dd0eea6d19c078d53bb3708fbfdbdb9400141d29f2c7326ab3529e21c
z08cf0135d31d81d847fdad9cb5068e98d00226ec4879cb30a1ac7290760f27a1ded9874a8c0b35
ze273d1bcb016619830fd9bcac61eae8f175f81ee0d09ba315c92e39053e550588a6b0339991b8b
zdbf87cc72243c951b77bd6b21785a1e013b76c61c5224553c39443f3b1dedb24e09fd59e8cee0c
z8fb6f2b630152536fe81d4f37401084db6bedc6d6e01bf6e4c1b3980b3b2cb3ce79d7d5f736ac2
z2d711d8068cd8ad417f975e6ceee351446c4f0c21177c69282ef73e1746af0f739dd28335fba5b
zb2c166be02e0a8432199bc61778a6fa4b628822056ffe11e21d576b41497717fd6c98b12290e6c
z34b9ad4f39b292f40518348a9363b1f898d27d378cac7dcf40e54e66a9e55e7a29101fd3ed6afb
z1ea8e613d582aa16e5df10588dbfad994e92db97e7b25b27f9528096c8403df5a61a563ab6b300
z76f5225b7f3331bfc1b9614e0affccb12f53fead4bab45939a3d8074f281396f676f9821c9af75
z529fe8bd8a150648f318db37d326f9fa9b9f8d13ef08b1827ee712a6dbde4e3d91df0aca7c547b
z502596d421234c592c8ebde91ccad6a55a31b6ff52c077202c113f6ed8c0e1dbbe93f81b55db5a
zd545dc619db631e97283ad39c9b278cf89e7ad2d7699e8de0441c6a864eac5b1bc5acc072801c5
zd0120052904bef0525fc38b28e7f14f6e1d2290078decd6c58f41bb47d6bd7da6879cd047a2574
za83934d33446b435ae94b57c539f9e967373d7266627f4138c45de6b34fc57d7c70ebbed0a08b1
zc687d35432591884244fc81db651f8884baa6946b32407abc021bdd92f2a2369579fe30f7fe825
z504e91e1c0834cf08066e78597ebb56823993299ad4d21dacc9bddc4dcdd595dc55b564bae24b1
zb90a553d95d40e59e575a536a9c330cbc2bad2d22574f1e20ea918156f1486b5438c11cf469f7e
z661aa59bfd6a4dff218b2027028a2ddddfb75abc577dd847ca15eadb42af5a073623a304bb30e1
z5f04a2f367a86f9310288fc468495b73dd5b5468d2dae509556649eeeefca8739ee2d3ff4e7d6e
z936e0a5b73c1beb32f03cf1f8714a20e6763522695e4f6f5175b6d76cbf35a775d3ea3e1db0ea2
z9ed9c3b697277d554b1aa49a3828698d2ee0739f227ce7534cb908b03eece24dd14ae221b37bb0
z7b98b6d2db44e3afcf83ada5b056f0b17afc4aa2a17112c181bdf8d2865ff40d66e4eb5dc66fc3
zbb8856610f23a207805c80c4f445779badd05e7859d9c6960d8b3effa3b171f0d037f68341391b
ze03bcad14fedc53fb719868b5d8304abbeebf065585ac2160c27de70de24d02dae807fe2771768
z095b930b7bcae066aaacecaed543d33052de20681f45824fad3a6b8d3c256cf9ceacf74454184b
z75d86d1245ba8a13e41196794bea9fbcd08f4d0a91e01ea3f705843a697f6e5ea26a8c665147a9
z49d8c1e9f87beb099843d67696d9c54194303ff0338bdd9b8167ddcae76a7ae3f812dec1ee7530
zbc9adc59f47a6b89b28f0559adedbf7491de5300f3dc1c346908eabfda08014923586d4eee21c1
za97c1e7095ec15cd4950de25e8edf55ffc2117839d7a95c630acdbbbdae5c96072c8e09d132aab
z9f6b8adea1812add0102869a06cca01de2c80004ce74695ec27646b7c47baa11048fce800ead7d
zd379f710e6e702cf3cdef324ae74c1c417535a037b11b27c4ff20c84a2a0f1f5163ed1377449de
z484e4f4ad9a46e506b419d010211d32bbc5d3f9621e16486af071e6091e46330b08f3e0eca97b2
z2be14076b969658ee7deb355b2ef170599e25e7315bc4d32324d6265f91fdc09a73f22408a67e9
z886408b9e7aaeaa81ab314289c21280b2941dafd1d29b0f6c5e83ceda6226ddcdc747b2f6332db
za2af23facbae584e934d5064a63bd57d9768db1ad255020bd6c2c3a7de16fa1abc3fcd97cfe0cd
ze7de524c6926e54f12928448eecaab205df9bd7fb55ce61f90ce3a6c91faf2d811611c06d4a37d
z2b5495834cf22bd2008505cb08abbd379d089e1caf13bca09e47a8baa59fb76d1673a34ecfc57c
ze0519640df9e05c8aab2ddd172dfbf53a192d6420e8e70c0b3a67aa74680e394fc3a4f0521db1a
z48921db1cc4604f6ee7ca37a3b780d067111ceafbabba9543f4ada01e0b1f124a7e59a63170cf7
zea4878caa88a1ea46914ef44014d6c40a9235c34f1f67c06b51bdc569b2d4d2a03e5d09446a210
z11beba816b0596bae8c1cb59efadeaa0a9aae5e4447b1f1bcb7587fe04d9cd0c52cf55c17a0b8c
z1672203caebaca1bf771deaac0da1496d48aaea2f4c78ca492d530ae3f6cf8e71058e84f222301
z1c1f49c4843528493af2d9667fdac1f988e486d89384367e44b205e80997a80277089ed28113d6
zdfdd4ef429cf33fc6f6953fd290115b386e0d697b74d1ee5c6c56e19f1d1529dbb213605fd464a
z33ea54ea0e070baa363c580666a00671b26b6f2768fa4009eba548a272a95a657b016552913337
z65c9ef221c4597268e1e9564d0524fadbf14eca3579733dcc74acab0546273cb6606e253bca1fa
zad32657ee3c28e1d3e03d4406bf50d2734188ab3e230db015d10a5eae06c14ddabbd4d6ad7bbfc
zb80b3e769ebfba4be91085ce153868e8ed623095ba5b7df9f3f7c4e538128809293571db720814
zfc14bf8fa8edc24e64122631159890739a62957ed9ea57e3d90ce69971e90427ef7b075c7a9660
z869445acfc9c72465b2860801d7648c116d997323e7608b03cdafffc8e9995fa4b9d49e9e66d8a
z6c3a8311ba0087c6f5547c84df235ee3792bf06ef62b4d48ee65ead5f650563a67ed25d445e6fb
z0c1368859dc4f84677c4db7b11aedf04eb0fe748fab450287a45da61ea1053395f1765e134676d
z4767847b2d06f5e1d319f3698f5ee13a49bf4839dece880dc8aae11acda0f6c0e918e2e2665e92
zc85e27de5d9ce9312fdee231722df87edd2c1b85eedd8325cebebf55766383b0891bde9db17ea8
z416b6fb2037505584614091576bffa203afc7ef93877c73fc0d2634fbe5dbaede1ca303d7c7cfc
za7cbc4fa3a1f319fd41d468238400bf1fb5a96f87f89aeb9a8b706edc3e1bf2c9b903a3d415e76
z46f67aaaad90b133cf375ed3d27a8e1637565b18c85dc608e4d7a7b74adf1543fb161482d356f3
zb16552b4d1bedae286a9f79c6465297d6f558e1a561a5ae92fc73cdc38f0dedfc0c899fe702d5f
z6039bb5b0e2c387971859ac444c7e8436a5e0a595c89c3c6ea8d723bc0d9cb09e97c1269eef157
z044278805c56f2371a71035a89e8b13fed44934bb47473037bf9dd5af8a2dcfe311925438c8380
zfe382c5ba770f24f641269a4df8c22ea4eb1b126bd4ad50a9250bd90311c8ce7ec14fe0cfdcb90
z151d8690b1aa9862ca466b99353c513747b1a00f613add991327bc871335075ac6c31bb38cca85
z0f708978317adb476e43014193ca4427a1ed2d42ad3aa50dc605993c1cb732be252604bca92f76
z5661f5b748d5ae9801f8378434bb9ce3a7f64839580a5f1fc6a64b09debddff33fa57c06a139b5
z0b63884ef5cb8e82ec54d3376d1e58f2d07a0276fbf2b7e7479b7a4163ef8a58f9225168c32833
za3c64b938bc1fb8ab9e93d23b44889b427c97ace3b9dec3f54f24be5b859a9c15f2e4d7be2ba2c
z560ae0fa4af03f45ea5146ac4d553b07063fbff553b868ae51ff2ff3e4fc635100997eb7994626
z874fbdb3c9d42fb2e52d299a1fb246b5737576f5ac0effd89efe504db0a6cfc9bcb24a8e885826
zde570be4b69269d5fee4cf1e7984a11e75f2daefa13779638ab13b8e67608ea43295b7f964736c
zf96c75aab25db4c2d65d30d28183f291d5a32764f4f8f01aef86e3c0435d18620bc6f49a92b80a
z3c0a0df288f6c4d2d4cb4471a3beb82e74aefe1ffe276c38dcd7af73322cd6475479c528f130f2
z1ea981a0146e8906f78940f85c332f7b37b6544d656ddcbf93663a1b231f9268d5d060d995b5ea
zd02f3b5efbfff1e199818028f4e4f3ab91a542eb96fd0e2728fabd55ff1403d9e33b066c289c8d
z0683289cbd6ed2982e67844be76bb7238db8780b27e2f2cfe6ad3b24395d7933e323613f86c4d9
z7c4b54e83005f0e787e294d7c77da5e261f5978deb78cba6390a171dcfb542edff9e0c000484e9
z48dd3f8010879f0e09a566c3bed7f5a1c429f9c2c92e6e7ef12929fef746cd819e32ac4d6f3732
zf5e83f1bffb895ac0090bfdf72793276b3dc7f7204379dd4342fe365d75412b5b75e8e05c8d347
zf42dfd6a8fa10995a6112ad05790f363e26734deb6f9b309ef1f4c5a67d47b8a1ca7947212428d
z0641bddd97550561b897f7507ad84bba93bfe78160fe8bebc142a7963dc2f56b89e6ac87e17c16
z3bb719925a450b51aa147b016d1343dad21d0b9bf22073f3ae7464288a8c689060e63509494e1c
z69f52c8cea4e7bb3d6e9cc3c3484b29f040d832bfa6facb51baa4763db57b172ef5cd2d822d5d1
zeb4a53e27c06929126930b0cbb5d5c0705eea012d9bf681f7ee73932717b16bba3790fc758ff50
z8f9373d2b2cfba899b6f7c9487b928b065b9fd51880b8caf831e3850e2939ca24f1f6ee325669c
za155019e63e7ad1d42dada2cf1860ca722661daf97f71aeb642871507e96d6e34ed9dd2cc9862d
zaa6c3a52579fb7f8691cbb5aaad49fb4ac8ea905352e81e377809c85e94d0212ae43109149e318
z6edc7571dc376a91334a3c67fc918caf7da5f21db9e0f3157f5f84ad270cb63dd832c88f2630b0
zed85e01b7534159b8605a7b276f812b668cefec94cc56f9324b60aee596c10e5d592ffa629443b
z9bf3f657825caabb584470c95e4866d58b1e81c85bd4bf343c2c75c0953dcb1d7581eb9a732f8c
z6269e909c3b0a4fc6f79ded950ad5cc0096ee8b4d12383b756584cd1cd80f0816db2029e038320
z460c560f15df72f7cbe0f9c33dbf44b48968cd5d5f9f8b3d4d2acacd1e7bcab4ec7452ea22394c
z5e5f77633dfea38371e27eed0166c59f87c8d331b4f694c696b3a84e7c04f812625f6cc1bd0e7b
z9dba2935e5df50632f14b3e1b9a2447c91561fc427f4f2048b72fd816261823b975e014c516460
zaef8345e14748987c5d4747b8572b498d90e07e65fe558cdf4c57bd2d2057a3ee3707207fcd718
z4808d3ac4b95e2a630b1faa70fb197278466f4d4c8d1bd597c6fea1fb19f83efa8afa16cbb30c7
zcbe6b98a07fc1ce56d33d268938efcb9a07c01e8d78ba77d80f06eabb698795a39f4fbd01bfa0f
z1360cf5df28d2e6ab35ce1e580caaaea54c26d317cacab9b2888e3aef37570cb6820dbe922e1d8
zf2d2b49c76b59425c196f895d78ed4df62cd8b4c60eda1b3885f3118fe7fa7b62aa14ed7042f46
z56135f963bdfc51954743635102d8072f08a6f136c838e5ee1029f6dddbc50f7b53eb3eeb6af8a
z4537d43f4aaee119256be402b74dc64c8b3d814962b20aba2029202089933f885e1b01e9db23d0
z6af4505a5950a8386b248557386be0d48649dee9ccad707d34ce7598a91e09bb739f185defb647
z6bee08dfcef35eae8cad5ffb4d0b6f24c7890a245d9690e5246d2adaee1c7f48a138ffb6307966
z8d058064a089b7081843362a281c34e043a40ffc8502ad8f12ff809e47cc2c24921cd4a7a5b5ba
z1158631081a5f80e9809e95713d48ea92fdb54aeae64a3583c15896e8c6b7653f76ba3ad501115
z28c5cd69c8ef16d3ae7251b97e9345557a3290658ce8b0d47f495a33a27ba49d08ea39a47abd5d
z9677edfd213bde53812a5343913434dc5e5549e1e9a2a3877cbe2d76731a771193f42970dba770
z6800d4e215f968fa2fdd457af15cf9507a5426ca145cc1f5eda62fcd47e1d308fd2f5eea5da519
z28d0d6745189857c0baee55f3cb3650c27270ad1ca64ec3c0f971b27f3e38ef4e37bda599feca6
z4f27b45bdfedabf4ff8a4d684fbba75a542fdc5cbb328c93c1aafc3984ec8b1440f2f87e224cd0
z58a65f1a3a6830b83fc830f6503656f0107435fe0ab8ab2917fa90ba2fbb4d1738725276f3d987
z3a97b7bf14ac7018ca66f8ed2a2ee088f86c5c381ea02c3a942f4a1a8361b62e87748980ab5303
zc1dc836d49a0cbf99c8348c7ac78d180297116dede0e49ed77256606c1b50aa6ce3a8e513994a6
z0bc5cf8ae8387e07e3395ce1d56d48b26439e0f416da7e2ec75d3e3e5d4b096744dbaf53575da8
zb511a06801048eeb9d0217080678a30d568212619b31c29fc7f94701570c2b7b61d33bb3e75c5e
z4d2266c6aaad1ce185c2b5ee8fc7badb1114448c825a18d0cf108cf52a8a89e858a1d1f2b16d6c
z60509e0256c49f08df2eb213b6b06fa3d6bfef8799d2d04b4f49faa7c40499955976de712b82f1
z99999ad0a80063cfca113acec43007194a0d5dfea0f46283ffd4ef971f2e53335912737319314f
zc98282cd629b0c61150745f855b1f7e4953079aec7a3230ba6760eebdb1793b47be9236cc90575
zac82afbe5188aee5e63ee89eb677b44b468cec5ff492c7557e01a11ee9887f91276001717f2250
z2d27f9159c377dcbee00d22d182bef2b05c40db0fb5c93beb4e1f7927a35ea84ed7f7817456099
z4f3a35814cc249a9ec0d9ad6ae48d1e2365a88dbdfc3eb1614590dda0190c7f80389c3adecb527
z0141cd5003108fa180e4439405ea5a22e1f8b958a3fe3a8cb23eaa47601c1605f163b70286d71d
z763794854e31965cbb0b6cbafc4f613304705adfceb6aabf74bcb58268c5702e702c981c76e1a9
zf792a58b8953cf0de6a64d08eadec2c5d0f19ddc10a82b27e8d169a1f9
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_minimum_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
