`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1b396e1048595951af798d8de75c23e123dcba
z74156e068eb331e95842c597f3ccd341bf87af84cccb15a44d811686c10b5caab6338f8bd390f9
z35e3850857fe16a4bd09a1f73b16fb4d985cb91a2a6e022108c6d66aed9c9b28b7bfcecdeb30c4
z21adcfcfd1d3a705ecb82a7cb228b602c508facae7d7277529f388f1ae749d3922daf9cba774a9
z7a2cdbe51bafb7233b5a04f9bb9c3d371ea04be74069b3a4dd10e4f6c35c82f6cb174014a35e2d
z402e001c822d16b1aa1074708a615899420d065a95dc28756fd5bbe26801945392ceec1550bc0e
z515f0fdcc539c420f798c16eb9b9a870afd7c2d087012d56c6f5d61f91202b9ec8e4e23c2f42e0
zcca954964eccf2c9a8fcbdb189ecbc1414ef7760444dd7b8da02d1eb9890fec73370650b4ebf34
z957ede5930c6977e92eedb14f0b7a339dc32f20f994d01dd3c5317c1c2082975bfc237a581d64d
zc8074e2c08f317cbe7f1667e3171ab757132d8b950b61bc2d35a431f66572bbd8eb14674623c29
zcb53df71e13cb1e1644ba85189af6e0b860a88e897e0a058efd779c076f821aa87c8804a441b2c
zc9a100d69e12be91b37bc1beca2ec7348e6cbd8c1e4bc31620d31f377592be45577bacebfdd441
z4e20fdf353524730f177690bccde50943390b2a7789fdf9526400d7411e69ea6a085eb65e4ad2f
z0d7d638e936b6a102c456673765021abd616e05824f91968d5d6ccc27b1f0c6f67e1e96ce455a5
z4dbef7fd70e2714ba0341c0577508c82e42e8c8030d3f0faf904e08b2c1f1f340799eceb62f7e2
ze74bb96e24be9fe8951ea1198fe141df3ba90d26679da18716e951fa32cf929f9810b631807ade
z4a38ba7766383654a2d658f532428391356709f028d564b6369be33b440953d31e459134bc7419
zda213e2f59a72cf99b59439794aa64fc9bce4cd215f18bf44e7221f22dbcd32da392b310a3ef8c
z428b82155c7d6871de64aa6dfb97f985334a4b641b59c9cb4e6a6d6c7c138ba2699377dac3753e
z9a5a830c3f12f887fe24ea7e27615af09dee1550fa1185e86d599a4e2d9cd123b76df3be401278
zab9e13dabfb01c3d04deb09383c967b0cbcc4500b23d7bfd93207a6c170779a27f5bf924d607cb
z9c8d07d33646e28302397b0af8f77115ba28ae577d69944747b4966a1bc9b1c507deca8358deb1
zf368d955a101bf59f781babe62be735d25011a568f08c43a41bc498c260bd887d46a1a0e452190
z8ae1e1780104d506f1532a8dde6198b43593fc95940b6b6a3d6803cfb764ef73eec1686cbe03f6
z266fcff63ec3bf7e3d6c8e479b787aa8d5573bfd9930dd2d05c314edae861b129a68e3dbc8ff91
z761b60466ff57d61d6c036522eb23399a529118249d02690c6358e6c3edbb438f332daed5abb6f
z16d414551810d913041e71390ae00c99dc030cb238fafc50b9a9baed68f31bf44b8f96c080be42
zea45e29bf16b3f717daa35685434becbf81a98349f2b7b1aa7937a1e690a28f762776f29fda63b
z673bd684dec5dc4ac412d31c731812adae23b7c568e0645c78120c878b18173ebdc6d0098cd010
zdb873803745baa288a86b0a36a6139cf4a1dad586e83b5e1f52d4a75641038a05a767d6ee1ae1e
z4342405310c6208ea7d736feb69ebfbbfb0176699b075b151addb5514ba20ae4e5e04b172962d9
z95980396a023ce07a6813ca070a1c3c6383db3d3be08c9036e65e978673ba3f009849994ccb301
ze5c6d73adc259804a3a41e82676e2681097081259400bfb28246cc184eed384d7b8f924abc5a81
zf5380353431369579688ef39e11040d9e3ad6ef768ee5d4a8edd8763997541e7510f603ba48fec
zeaeaf36169efb88c387bac091f4e7add8b58e2a5bc0e6a9a1d521a2170b6edd8a3db0d87bf338b
z56e795bba2bf4aba26e1f195b8530886bb21f5f84868735854a1f80cd033fcac93db6f2b0b8286
zbd2eed4f22cc122b099c0a145ee1c62b56d5a3709d97427298201b3608fe66ef8cd4f6e3e953aa
zb85e38909579815275c70d7e7f04a1e6a0bc58a68cbe66ba6ed5aa3e51c8622985d54984127195
z2b9d397d8d7c1591fb6643fbe5b64cfd303f21eaa85f18300d29fea43cb79b1feea817d1f72827
zbee83ab8e1a2d1ee6ab1deae01efd5839531595347ef09249c868ad36a686e19e09e5db6be61c8
zf7e7176baab959b29ce5dc930fbb98a09c66d052128b29a56b55a66f32d352fa3223044ff7a6dd
zb043710b276523ca208de2c1bb29b803b6f5f679f5a4b2799bad018b18855482f655b04194a706
z60710bafe36a63ffc2b0cac145a35805518ef57d3475bfcf107c0aa3ad208e5cbd304558e44f87
z90e9ee0c815938923794de29f17f2805ce2cd4ce3fe4e7b5d0f87c5ef42d723411ffb0dd5f874c
z20be030066ef7cbb6885e7d13bc6f5b4ff3d83a3be568321f13a3dd6945ed2054b2a2e30f95a66
z9044511d6bb4e6d1c7337c9eea53f939d154d793481bd6403da5b83e2dd8d64093293ca5e409f4
z31300deb07660944268d3e6218b15bc7fd58fd82d633fcdb266844f4dfb73e65c50353bc9cad37
zbc98bdc65dff38f7f292c8867af8f7620bd08c168dbd982c37e1553a54a978a4cae086364a59bf
zc8d8ba89b1bab014bf882bd34594fae2369f6d1bd8f8cd9739412ba8f68c58c1f3bc86afaa04eb
z74ca5f7d42ee325b3369f8cfb18a62fb802b238a047ed73683725ab67d277130d3fb8fff160347
z000ef579d814485cc98993a6041fbc57f37d83f61a44e46e4e6ef8e2ad752b225f68ef23a31760
ze14be1f26294d985062cc0dbe34c35e66d7446ce969b29b528fe9c443edce9ba0f453c7902e054
ze4200ad51f6de1b49c29dc703ff097b2986a0bf098b6f32ef3947cd6907efc691d8a16c60392e6
z4de33f6cfa4db39eeb44b9802af8d89a352485f266f852dc2bd2427f8b761982b17a3512cb8bb6
z3d6284f67abc9458a848dfe3bca45fa086a50c0c4b025bbb55eac82f6a1809e965596d09afbc32
zfab5c49575107efcf082212017cac9cea4b5e2c4d1314bb84be1297165da742ebcaa470ad5c7c4
z145117df618b38ccdf0a39f8b41edd0f3e7c92e485867ea4deff7172b23f89bbf0f3ee8bd57005
z74927c42cc502c77e882fe3c9cf568ed50312eda05b02ef44ab0c9a091ed51ee3831dfe73b8edd
z0e6f167e06c982cab03b80eb28d94c6fe6f0d0fd4f7d74597fbb55391ffdfdf2e98e30fe63d8da
z786d1f9983f50b8d7d6f5d20a1917508981c1c6fa79699b98b365e69c3e16bd7b1bf8e7cc86322
z3a41683147888c4bb29ce7572df43af52e3b512f67a1fe2e03a6a15583d0c562bc1015b0c2d5a5
z3fdc12060f49478bf92b44a0407cc1761981d7d431b8a33514c3d1f540e28dc770740b91a235b3
z81ea87d1383ad2f9a60f39b0ee7665c33e2a852d642ee026d71314796e4dff9be9bc55c1aa76e2
z939cd34761536fede715835375791d2cdab74c733f6d416557088b528fe89bda6782879287a10e
z7f52bdcc9206239df8a57eb6acdeed1e0143218413a1a485e312d2d666007e72bdca4a5c066743
z4230967186636b27a55ef414cafb8005f183bf535f986cd481b90141ce1932fa6e8521509e5104
ze8b9495a9a56ce370e8200bf23002362bc23bd22e5fb95fce2d8cddf78963b05033a1c0b14205b
zf763c1376bd318eb5317038715a09950ad2fcdaee95643df4d4e7fd08a35a22c6fe58ec9f10cbc
z35a3a18febcdd93ad2e60d7882a69c652cc20f46b70fb682fe4e7f5ce8aa3b3517c0cae06668ac
z77c5fa000fda9e1ea4dd2666f0fb81a0569e61c07cf158524b8bacf2aaafe1440a5dbdf64002cd
z28cff0db905e4aafa5f5b0c478a4edf608fc7c0f04fbab20899350686e4fd20505032d4159205e
zf7cee344fec3db3400896a39d96e8578b226df3215e5087dbcdb82d6a8b2f1c0bba551491588f0
z3d5d1fe612e848f827fc7608d1070a0e48176bfc230f74ca78094db31fd0f4fd1e70d637833858
z70e252ebab2200cff48725ad325732ea15521bf27ddfb2b171260c6944d35ab0874f778105f51c
z298d4546ddf9bf64613178384819ad2b34fbd738147ca1688f67fc7216318dada7ab5a27f121bc
za162941a8605aaca63f88ce5b6595efed543dd1f52857653bb37ae8ff5d843aa2ff6713b2dbae0
z89f98aa0ed693194367c0e2703370b2f8d3d313b307442081ed0d014392fab888f56110b8e5454
zd297f2e047fa5e5693102c5be0f1ee2210d31eef78bcc2b4e4ca9b1b448b9c32de8a5583424854
zf34e4d6398690ac8ee62247dc945164b21695428487c9f984bf1ee3c127e6a626253317a0db984
zb1a221d080455030b3a807df312c0ecaf26607189fb811db6a48dba262aa382f2694d1f7db1811
z421e3a0e0ca7357302fd9dd3e99dc105c1eec6660f9ade4e8c77fc60f36efb4d2b881d6414ab32
z2e6b1bc476e38f40239d1ec2a23d96a59a8502a6c10957494617e45ba2c08f5df81ae7e41b71f0
z5da93ec8deb5ec442f71c59561c621c632f7d37bd928d5fd4421f9a3f269770010e7335bcd65fd
z09ed73b5fd396046e604cb66a624c9857fc5e4abe345642bc5348446ebd285ab83212449960a3a
z63a68a83932bfa03b1d51bec5a8e90c3defa835e8d0bc8e56b99a645588ab063a4b1c0328c962c
zdc3ee420cfd24fffed40ba33ff84a9ec45c60fae5b50cc9cab7d4c21ec18d25a73e71244eb1ea0
z0502c69e489c20e8d145673815217122b4946bf064894e9bc582b146873e0f19b48edc65a02b06
z44cfe3bad508b31561dc644075d3d5fe09be26cf6b2f9b7d13a7b0ad3c24584b01b20b4e38e28d
z1c0a6d2d46e473987790eaa6f84ec02bc6783dfa22397112ceb69e8d43c1645ce30052813ad97f
z733a2934958ed1462548fa85a292e2b99a17ddc3f4b5a9d105004d515edd8d3351ea16dab7f339
zfae8aa9a282213212feae3ebf529fbb2c61aeb644e87aa10627d5ba6de9a407f1f47307b8dc13f
z350e336b4ecd5674a91083732c4ec32ac49c7dd88798e92277ea0c1725da39df1a20983f83e354
z510db528e1f6b1923a82add6e7d0878badbab6cea5f37bf88534ea7d6ebe5e743fbf90f5a66bb3
z7637b4aa437ab553ae4d00e41ecc5534c1ee70123a50986058c49f6af0e0093829bd5c429b6d10
zb4ebb919ba6f9c7b8fa51c88a810e024a437ad159bb6786d38f74e103c69cf7db0b648c3c6f6af
ze94709afaf367447479e5fee95768c4ba8fb72568c3cc402af1345cfdd5ca8932ca8bc7aa6a844
z2f504128128be69cc2eb7a3a08f80490c67607360d9700b97ee5ac76a09796c8559734cd1d2d86
z0d0bc1b2cf88a80da80e664f9c0faab5fe3f351106d46952fbacb813c8bfeb213b2b2e814f07c9
z8194e41d2c8efaeb8118071321f4ba234b965e89579ba635e03f0654c1980ba4f46ef775738cf8
z476e373a80324800ed9a54f7c780a89d34400fe947a0206db84bccbafe3a20510625baf9573706
z881dbcd5dcd4b55cb2b443b98f3910a4159b06c4a5c4de9d753d33c965879ee6223e1fa2611474
zfd53d11cac5d4ff1428bef15f745cc02e4703cf5449ede27ff066d35cb6e7381b0642f87ce3294
z87c933cb7db2a2c907237694ecdaf6ef7461e197d0a857805c04140031ad220fa1472ab2b3c274
z08ac01c848c72d7e81fc80608a556ca278103d4f00368e931513ab6791efa6e9bfe5aa3e2d57a4
ze3bce161c69e4e208133f76e1cb8f136c80985ab5db7dd0c2239ff7fedde238d8df7750eb294f6
z17f9d77e85841e8e84d2ee72d6498eaddec6f5562b2d45069a5ad4afd739db98096b46b2aae9be
za11be7ddb7788f81153566e2e6abfaff93bddae81467408248017876d5e330014053f6ca4bd438
zd64cb2dff407cac29d0fd714a78178e958977180e70db72d9da4430693a79a9966a2a3acf31dfe
z20b4d2312b7fc1666ba1e0ac9ce103d6dcef5d6a47c19a858879285973aebeffeab6455d74c339
ze6c5aad1d16d91889e000d31c11f723de74d3514e2c458ee3744e197463f9b3b4a6bae5b3e80ee
zb3db75b8f16abf5c24c0061b765fe50285b633e9348fd5c3927b38a2e3cec470c1db3e65f1ac22
zd653ab3311e39ad0813671f33f025968a0249b5e28bc1166580835146ffc72b0bc3ade6d8e906c
z2b594c2a6ee2852991c4edc58a584a6265db5046ab251ef8a77cc3547d61a783db25692d00a02c
z54110509b5d40f4d895e096bcdf87de296d139f8f3e8f0a45299671a1e5a76e66440195f5086d5
zac2ba6906952267637e5f6adb489f92284ff9c29a2ac3c346f8470589e1c5d1b206c0e3db5d08b
z5651a4693a6596ae156eea0442d4e7a94d274298c1af249ba96f527e1eece285646baaee658da2
z4bc732a82efe310f3243d1219520e89f5c33dc73d15d3ee87799ff594221699c9e22e36bb658b7
z6b35cf85324c6117d3d239c6a0c23f16bf6db7ed8949f7748e1ef47b1533685ee8ffa367b797f9
z02fc771c677509def16bee904c39ff8e8339714b8da243b040dfb6e87088d7f72781b81d402ddb
z48aff9785f30ae20ab5cf872cd43af1f035119db43bc8c40839abb181d614aa2a0c3428ff02b23
z4fbfadd8fb0f30aee118ecbe6bc857be49ba7715d55b37cb4d5027d4ba0bd7b0c84ad6f69731ee
z438a92f16934e038d269d0f49c63b4d933cff70c9e68818af4958a698bddabb85f40d993af158c
ze6b21ce379da6b9959ff721f5298ee5da0744c0a74b3ba2975a6a6490155000dee381fc3103ad8
zd3018f28572bbc57ce49d58afbfcc386a9db5cba38c9c787d4224bd8182a77ac0ec1233468a86f
z51d9a3829289d219c84839310781cdd60bf7ffd80909c8148b3a5cccb183cc775f88d6eeed0161
zea8af41f3cfefea7ec7db2db8f44abfdd8c438e8a9b1084654cba587614d3bdef78609503f89a7
z5e3e3586deb6b5362274737b534a3257e51ee52ce611587f5f97722d225d81b8b4858b133ffbac
z47cd6f0bebace318cf6c86bcdd0fd20d33ab4853247208571a46efa3b003a03008e36c003a7c2d
z503a35589b44791435d9b16c0182f0a55823909ef88302882f747f06a238a46cf297f09d5770cb
z656b7c94459d7fd9c5bead6086e64bd2dbdf6c5283729eadaefaeadb73c678824e2356fdd4aba3
zb5ae7d245cb53a836dba7088625ccd4a060b323b9c8cd1976845ccbb9b05575b68d1a4fb6829d1
z23a26cbe20d89265500129bb10f4528a235606766e90b69debdf211f40db0d9abe8b1de4bc0c7e
z3d0a94f886cba0c46de8752ea98cfe1cf8e7deed9af38f0939d529d48bc4a67eec5ec46bf3e5d4
z1197b8852ded5517a3046c179a600c81078ecf3ab5b57b484853ff947ffb850acc49821a773300
zdb4035196ccd1d2e5878221a35e955b36981f9bf930401df763ee04628e909a7ac79f789962ed0
zc0bb099d0c3171f9329e3b8ad5d90a4ddc68cc64896d7c53fec829a29792338b3d07464163d6e7
zc04973c63c6035f20198e1a4e3dabc05cd0e4fa823f80c1ac5e18cedb0911ee6d3b5ab2701ad22
zb63937667f2fbbf67ca1f853f7e4e088cb2217ddc4b350b81eed1ff4fc9fe473d0e31bb02859f1
z2a29fda54ffe70775583a3910eaee838399b95f910627560b87db3401980682dc83e8c0d46ea21
z9a0e18e9573e39917b9409fe2c959fdc60dd64bde240b9c18c293d920f733689be8f27322b3222
z458787fa4a3ee98e2cf489e76540a9f41e638f676172e8a5b99ada3660fad100cb12cb66de6e37
zf79cd883cb5d8972543764466295ba9ccecadbf92eca30c7d6ccc5361ecf2ea35c4e49efbd07d7
zce601f0391a64a0db2c1b626f0dedce7c7fb6a23495e9c5f1cc248e7bbe55db221072bb9c599c8
z8067fb2564006a1efd3ef81a7d722a03e7e57141e6845bf38080d9b7b7202766b17f18bfb51347
z967579fdd86fefc6116b6f4fe2c5182783141a7a5546d73bd5c6390e5df15949e8faffb7205439
zbae7b27e96c15ac7539f375d3728d4e3c92cda48d946ae1487566b552db73083ac1ff63970f35f
z0543d148a0733efedf56a3e49125d601777275c8279b3c6297e2a72af5e954d6717e6c4864e04a
z16d3bd7de14692b13605617224dd514bcb110ed01e9145e07e9b286c22b39bb6c225f3565d3baf
z12225c2b147756afa71a81b67a23921fc2d0dd1d509a381418f69f53055f26110b8dfd1933bf73
zde01c41c8705c2ff6e15e5a6c14daec2bedc675faba9bb06b874c641aeb452e3f429f394ba820a
z6113ba8637321f732117ee7e5f0d69943903f65a29392b7dd6670736e41b3bca1d0e775d705fe7
za7a97668b6b9064e8453109c30ee2d2710adce72cc0e98e54539f477f63fa84393f6e6b26b25e2
z8b4ce50529478db7462d4fe4eb5d9593325e03cb674218710e294d61f17ee2bf7d9e829d167e3f
zc5ac4320f40a61c39096d3724ccc7561263eebacf769fa01b1b42f7f38beb12dd079953e3c7b24
za235aad871c821504f1e136520b6ab119189e688c7054d515e60c18e9831088da85b65c4f275a2
z38ffad9d10e91c254a8bfbd39141dc9e9e590f727d6c1c63ae7727165446890c8271212cace0f5
zeab0f36fe5836a12105b6ae1ccdabc4a5be85c9c510e971ac0f863cf03de858aafdae1d11b6fa5
z21b8e80bbc88b72641b8ad825f25c6f12534dae1c726cf09cfb5d9f2eea5eea5099bbc2885c580
zb0ebd43eea8052f179773fdbccf5a68e5b28e49b0c8eda9d69945ea7b63c3166f9f68d98c3859a
zb9f6e815743eacf9cad7cc88ca3aa6c98db52f61d72a4c0a2376e28a95d51a72a71768987bd972
z6c9959e43cd09c190ef202f760a701f6d59d9591ba15459408932a0334e0252f73e7795e7390e9
zbd38b2eb16842fee778cd274ee3ab18a83e6f83ca51e249fb46e9439c892a9bdaab452758e7c38
z361f4ba0c8cd6e3829344086b8e59813ab81f55b82eaa096bce203bf5f55051ab56de4281bfa26
z85f5402f3fdfd7f14d679bfa29fedadb88291604e291e9ea00be82cbdb93cdfbf3149948b8e866
z074fdfc7511a47c4c5a7e55bd385f020b99641b20ad347b88a073a3e745d4052377cf1749cff1b
zbc624565f9dcb0edc40801615266dffc3a75b806682a4d82966e2a5434a1c7169ae495a0a426c8
z35a79a60541210ffdcf682562c6134261f3bcdeab8c6bf0ed8de6c482c667812b5d5615dafe3d6
ze207047a8f7f67640131c6f59bdd6356e855aae0bccb709da8e452c33569cc43c217f893433fa5
z9e606e36a4fe51141e11a4e802c4cb64c72f05b9a5489998c4ebdd0866ef2550334d7963019d58
z83605a87ca3d66315e325fc54c98a8059211d0cb3881090670f3b1d4a116784405b17ac099ba62
z357cab58c9d923f92c2921c85a32c01312c6c615d8d8b2bcc470da0f3da87139ed43c71341197b
z2214016e92f321ef84933654ff9b645c45fd881d813ce9adec67a7dd20f0e8d4993ede76356632
z544e9e3413a647c27eb4f3b9ffd494efbcb0a5c5a9fbacd3c4995daebeda0c746b1ea253217273
z44b7c60d2d1e6dc059a6f3b01c840a2e6ff041bb6b3054958d9cf996e6caf94bc88ad5002bd6f5
z5206a663dd7a04590b2cfb2a299bcc560dd2cf08df21826de2fc867a20bd7c2f333afa83bd8e6b
z9a7f59279b8bd4d17b834429c621e21a523735696c0737030ea86450b0916d9c04e46d07ca3433
zb1fe3faa3e2c19e30df676308e6b2de0dfcb2f694fc113319859448ce855e23b5232e93353fcb0
z6c2dfdee14900e94182c991148054289395c708a39d9d3c7c5c16d682efbcba06d9795613be956
z9be82ac7d7da0f861339061ab10a1c5ed428bc679a95ac5ae6f502ea50e829a6cf812524d3bd93
z59ff9aed0b9ab9bcd56372e26106dce478886068d48a735825fc0bb5b0de6e55a1122096417a09
z37850a05895a0a048f0072f1e8edb04d4f583c1f0f3d909d17d861c2f7b8756bc6cd76b66e31f0
z078d0e739710a5e2f4fc4b405f7eec68053ae5cdeaf6026ae4b75903e8a4635cd02503da4bcfc3
zfe009781372d49bd6f6341ba1df5e60e00f36d08a63c448826254c256cb6e115055abc7fc638e6
zcbc0a7c20f203e134aadac71340691183e06ae7a3c6e734a16959691d2dc5ab6706ed35a89bd7d
z820a76fc38e7cd51c2cc1723a843257094cf685663e53e574dc531ad6e21d0ad43ef04a07e0e12
z51c86696b696f3ddd0a025d91106338a84c15f3f360997f2881002fbe47b1cb897c2174a738ad4
zdaae7d86c405a37312d5790fe9d3fca0c1fce59036f1dad8dc5bd0a68ef34969eca2f0816d107e
zfdba2c5c9cb9c3fe2031c15875c7f47933283d95616915fc43849699f78a65ea4c4ab19fc60e11
zc8c7275c2046115ffd56e07da367dd8c3732d8722321e62c726aae62a9d6f85493f692269699cb
za7b8685cbbab8afe3929d6479ac0f79bfa64263d21d52089f9b97bd5f655425ef1017cd11fde47
z11a831c34ae181b3b858dc5ec0c6bee651c961dce1869e7c0f459da0f534138e0c2d9620b400a6
z50e19cdb1c68b4a596abf228c0cc3e037afa3c29820be051aaee94856735017e891a4fc13d4d66
zb058cbf0717dc972c253a453a57ca335fa0650ac1d0e3b60811376ded9b5f670c7906ac51d72c6
z9858ad09e36ef94781eccbf7253ce7c9b8f88c7204f626dbb6711586ba0b81921c1cbe77daae53
z5779d181f27510145375bf37f2710da6d0bb74d57489691d73f8a2cb17ad58030982760e02c716
z3e9283a8c1930ca119fb820ea60dd7cccce0b15ab715be487fef54f4bb80738135ee4e8b328505
zdbb9dcefe249b06add00aaa8637e27a0187cd20ff1e4e84b37cc0e45e946dd437619008fc1f425
z68dce0a06301e06aa26f31b38150a87af427a364557db89e02c26eed017111c7a9ae099f3d12c0
z804306302e0e7e6195f6eb30897f5f88668dac1d7f74bcc2a22d2a92cd975a7819502f9c78e138
z101a1b6521843c83731e2fa14e535c22bfd8a5a4de92d784551a853c15d7e752f41e1b1a9f46cb
zbe864ffb0b854314159a140094240d45f39eb758ebc7341d9a80bffa9c61ec4a18f2b9b5036097
zd5158df44814931a98e96c2b10fa150b0e7f65de5bd258e6d719dee7a2a580e78be338dcf8e0af
z1eada8d8dd7e57c21706b09bdca517ad6290178d2bd506addcc8318c18e1d39be4adb49d3f50f1
z5006afcb152043b24a9f982ddd51300554c1f2bb879f4e06cbb018beb36ea937352354aee8bab2
z05599df132396160304768e64ab72156765570facbc9db837651132444095444b0eac9d6c95c4c
z31794c4c05f1fc36d4b46dcbe5f511cbd996a2fda89454b13cd488f65d452d7cc6a0fcd444ae26
z128cc95efe4bbc07ece8bca753e0e84d03476d2a6bf5995edd2a4a8b3f9ed0fbc9e03d5a5b2b2a
z73a302163ffc0b2fd7152fe534023fa83ca076cd2910871992a1d0184b34ccb8bc76e4644c8527
zbda955f2d8c26d19554e6edf1f1d82fa4f10d30673990dad98efc329874360c744823e78e427b9
zef21497b1c0b7d6352d118246c77c29e5bfc0249e38bdc48a7a6e99ac42d3037a8b99e96570ee1
zb6b1198606d6afe6eeb02ce97d66b397156d794bb4ab77d304930fb857b2dc653922c28d3278f4
zfccf5a097d89e07f5132b02d93c5d10d2595b01cc49e1cfb0fcfd4d02a636588ee543a97d64e14
z4b6945ffc2abc625dff714eb5659341143fded1d8967e1e9cf7a7ca9fda5128d083c1043b9f8ff
z5701b3945569b5a9b8410688c4f3a792e7495657f2a9821fa5bc2fe2405b19a27a6cce82260b80
z4c2d358fa6d33aa8294fbe8f2dd0befb6cc72282249fb412c1fff211d39d600ba6f62f258ddc61
z82e250ce93395b2adb96206e040dd1f8444647e108b30d2597b1a49de39bd82bfab8248ad0eaba
zc57ec4b693b47aa608c76c329b71cb6e71b999c735c6601f706af83a10694b1ecbe9bd9350a2b1
zf9a1abf603092cf246494ceb62d0dc97a0497e90692afd27eb6ce12d9962641d8d89ab812d99ed
z6f0ce1a9155fc33b41e5013e7f63d06742f569ed9c4050224790597bfaa1e712450194127dd39b
za7096953e322c3b24cfc1f2fe8dffbc7a2ba52c25003431826b88660579fcd93422e34d5c44c8d
z756d96bb2e24cccb876778a3f674f3550d224014f2fe26ab5d4bd0e5f57d668ce1d2513e709863
zef28291ceb3816feb441e7311fa20197860dcbb4164b58b3a8879b58f0d8e62afef672044bb948
zb262f50e330a8540e59fc7ffd99758800b8eb9a7dd3f8d6b39e599be4a3c96e09b99fe227ae6d6
z53042818644a3e016de04f0bec8f6a0f2bf0ca4ff0b53a30d90e34e2c8ccbe52b3dc4dc72ce7ee
zced778a5c41575de47cdda2621cec65eadd772748a17e6d147f5dcb6b77b1b8e7979ced32cd672
za191c90891365398d5aaa28dee6680cfff8e356a804dd29d16cb25b84fd3eda6c685c6f9635f2f
z091b0449517d8e909e61c83f4f52798c941eb3d53c104e48f294e1a3c48ce0bb4bd37d5370714f
zc7cd9bd7038e149fe1aaacdb367c38441a3586afb8d83410712568eb4a30a55e4fe7357ada4e29
z482a814b4c45b72719296c32a45ba4d4f557f49e9da31392e9b0ee8b20bb974d09caf8fce55f03
zcf56f7232e645b6bea8c621260806db40f067bbc511e36b19aacec6e77bac7b71f3feada3e2357
z101124357a549acf26690a32b5eeba555e7de70dee8e7e4a806a87a1d77996e4fccca90929a712
z50f9816d98c05851e8910583918f813a98776cc9328e3f03b6fb997824aad60248c55ad408ed45
z7a877e4d062d1ed25fb290a5725853e8c2cf6c9366204a736b62a89bbb78b92a5d191d740c71d8
za3bda8f005b6abed50c9cf21d74d4b06c9977341e1282895792153ca23c1c56725c607b34ea041
z9d5f33b774898d983f4ebb6db9176d8b7b2352e28071fabee5be3302300ea3d54b9de5372592f6
z40bec29a5bbf628ed8d1c9a087246ee1adbe3bad1ad6620eac2a49cdfc68b11b4008474948650d
z3904fd314094627f81e23b56092a7e474557fb3c41e29923fbf185381eb517959151faf825af13
zc7582d2b4f11f1415348cf6e9c87d2b65f97244ff69d5f611401ee5241467efbf207ff471803c3
z814a8fb8f9d7925bc0fef1740ab329a184fc6d9b2c34d0031dff170c5bb70ac4afa7d43ae30326
z22cc24028769de3829b97b9e348481b13d10c85573f4d7dd4748a820e5791df549024199866481
z8da2a5bdb69811170feb524801428556b089e46d00d05ce2db0f0120d8b747a9b9eb2e16ec0412
zc0df102fa4f145deb1efd636d2c5cf3ed3173fd757085e9d0162eb041a457827b196d5996bb1b1
z1377d82709a95b1468f74c3562aa8e988633c11f42e5e50d6a63ca8538c87e1a0b6e20791d41dd
z3806a229e3cc8d16294301855b3f6b2fe6c91c84f1cf3743aa563655863d58ad8d2ff0c9a3649d
ze4c0e70020f0400ad65ae4fb761daad54a526af313016512837d7f4d397ad9cbfd829e938cf399
zd57900996d4c8ae787990179c782ed52dffd5d8c8959abd7e567b1f963a23ecbd3fc559a8b52e5
za15646aefa74805f983cc369aa0602cd4c1383583a645b82c0799ebfec2ee6605f21864f37f848
z774dee4ee00962f7b133de26319acee05f832a338b413b64b364cd19057b35a10de578a5306a3a
z0a5b1361eb0428bced4af30409a4c9289d13d303c75315f44c076e3537b9e30e97287f30aa8ab6
zf4afd35a120d688861751a5a64446b416d3c844aaf3bc13f364e1f3ec04f98559701da582e20ea
z452c46fcead45f3f7a615af747a207d9b4843828cb2cf6334ed45e6820256421125d06b9fa7106
za216722f7615037bd74f895d400c77d9bacade9da9b6fbaddae11804a5a784b5b5ab0b58cae819
zae196cc0af35bf6ce2fa8ba631a0044f7c361cd3f6fd9cb88a66bf297edb0a6095fe601f51ce11
z158da88c6d547083d35d21dff5fe5298fb9371524482bd0284047086147d7e215e595c56bc2dc8
z61e0232e835941f8020a4c4eb9d88dcd9ffd3437997537fbf49c87cf610e7abd4d0b58b4e2105f
zbe803d57ef7441f26640ac23daf4cb8e087924df7f30a0f6a5298912223e3410c48a9845570dca
z3c80ae30748223f6715b3b3283fc4fdf42e26df2ede5c5363add6d67417838d7b10af9359d820f
zd7ab232d425761b3b98e0f29d339ac5da5f2f77c0362a61a64101eec75e2d2002ce1316ca66b90
z415e211ad1c96923ea97e3b2b115be4816c7ddc5531edd6f0bd9e8f4d138a7edf8ae0d8c2dd61f
zcfc6990ad10335dcd2d880daf867b4ae4360d13be234351f75797d9a0c4542b6e961d90e354325
z01fffc3e5e6aa0783aa9759e65ca9cb19b202cbc4af650649889396de0b317a1ff91c404d3aebe
zd4a74672c83c60cfa6a30b52c4816fc7c380ae56116986a42d2b0b0eaf97ce70156773306afaf5
zaab4432ff1ae2572cec214a9a71f96bd9f9b1511e9faa865bb8daf04963cd431337ec319dadc39
z41d81d2b8ba179658b8b791165af0748106b4c3ffb5caf2a4ccd853ee7599ea03309a671085c8b
z05b8c474ad1b84b81ea2a6af10459c7c0871a55b19b9e2e075ab3d6abede70a92b01a719ed5441
z612d4c1269e4889b86e3f1f98bb79a7ea8aa70934ba2ca8d399ddddaf0b35315717e712bf20e32
z9a68f597c534513d1bed0076ea37a1b6909d9dff07235d0a90d80f636789baecfabe66593a263a
z8da7b8cad0a1c9629d527ee5f1a0c2cfadd9964d1af4e968b9263e59bc574fad148d02418d8f2c
zc265bc05508406ac26aeae7abde16968040513333480a7936c5594388de05d5f995293541e8119
zc4bd1f6b528c08f601d540617772b7e54e1835ff997cd3f131d984f034a36dabdb294f4b981009
z2f438f82a4369106da7065fea1310010a7fc73e08e9c7d2ffd70d9d2569abb7a66552375c2c8b9
z8c8d4e8170642934c94e225b877293455021194096b0fe050ec70c514b31b4157ff2833e6a88f1
zcf98702866b64c8e83d91103dfe00ce3d7c3d96f280b27bb1e0be097da5bc500aa82fca1a191bd
z5779e2b4de83bc088bc59b088afa21314322f76f89678f120f47ba2f2604eb3d72d9eb3d7b91ab
z2ea6f6d3fca2f7a3bd66c09fa3c247a7f871d97f800f361f80894b2cf2a6dbdf9cb1879d6c74ad
z2a1614f21ea2ba535fec5fa5525c61cb0dd1b665e919c5e558705eae9f981bf696df6c66d3bb45
za0419e2524066d6e346bf35d40697a705fd997caa1bbb1188bb058943afbe939450e18f95f18c8
zb3b6bdb47c2f503365d1ba0b127899f1a65b15c7a8b41837deb5b98e8eda76d3acd49f9ac79476
z59984bdd435e25d3ac43152337bbc463de23ee5b78159cf6305b50c77bcc6a3d666ab044a00bc2
za1a2234604e4db18b0ba4d30621bffeaa375408ac1d3735909a02bc664ac39d1f222e7f7f75c9b
z63e09d429148eae07ff8d5e3fe5aed7afa2de8b60bce89d085ae27bbaa697b836f36afa14415ff
zc5b2f21b31b2bb461cd736098a0778f22e9325a49c6492e3db12006320370ef557dab90e6dc37b
zc0f094f1f001025433b773e66fae5ea8be36be71a90eaa3c4342d6ce85c16730e4da674bc85510
z0cb5ad86a02f8bfeb83df35928b691258932b1ba0a3fdbf044f88c7529e20a7c20be11e923bb53
z311ddecf2a701f78c2f82b233059e4541177fa71744172d8a415365ff8b7fe7ce393a85d24efd6
z0103327d9c516b96f7653ca06c3547fade04394c27efe7c4fcbfcd23b724dcad70ce7118a2357e
z5dca88e1d3baf69225ea814a0e02c37b68963851ce7aa5a0caa7c09c12c2867b10925706cdbc99
z72d6adb5e47375f9006cf6da314dbfd484169e0a79c45f0a4f911e34c33faf7038fca528ee59e4
za29d854f4ce3b5ac41f248bd60e8a63b25d198f4c63bed8d4bebadd55018446adb2310403b5f4e
z3c142221f3aad1c8c241835cecb9882c59416e2c788a3a7d8a9f6761537b71da80ef695c09de9f
z14249ca032fb00d0c1446238cffe212491629bc2d77dacd54d7af5beb0efd5bf42e4dfc0fb57d7
z3bf912a8c48f678f7462bff55d0ec101cd69f9d1ff7a2a504de06b464ec3cedb89a433adfe8f02
z89027f7303df3cfa8d079d7b41154624d675ac7f670bb0ca53842f20831408cd727db2170fd309
z188d1a56629b3de5ee69fdac3588deb6d509f41fb051b677804d0bfd1c19ae3328be52be190edf
z1deb222d4aa4ed79cb83fd04c0ecc9fa052f13a4d50037236a10bd4d82c215b7bd8ad85237e3b4
zf9e3225f6f72aad1e48cb442fbcde5a04b4ce8961346f26b33893244cc5ae0e87c18a5446f5c35
z7c424307216daff610b7f26d190006821f053653892de645f49d1e85c8eeb1da064681ff1dc409
zd7a8346cf6913db1a1ba8f729d998147cba0fe4d59ae3ea18505cc27351131d2796e6e00f7ac67
z0d5827b7f6c231afa7533d61db25751ab9b1ce4eea5b7bba511d2e8259f64fcb6ba07475f9c37f
z54f913e82159561c1006e088153e05dc082b400b51f7e0c1f73d7d9011493d7e482cb6ce7acd9d
z58a44ebf2a962b1f96c5f8afdf3b9fdf2d8d5b692f92a46b9959966a0ba50539941acaa921937f
z85bd3753205a4cb1722c0e4ef7c9dc90022d7dc51342780dc65cdd2c5619deb937d19bd18a2e10
z98f82bc596f5003801d0fe0bf207e8d8b937c7778468ac776e24dc07789bd280f2f2eb45e0accd
zbbc068c5e9c3a626d06e4e1cef5c26b735c3e54a07fa6296cb55239f95956a930368de022dd1a9
zacc3dbc771d45e3e222e85e810eff6ceaacdb7617f399364687ec166ddc169d09e7057a0118534
z850545603cc772e6e9b5e9f139fffb86facdcdc058491d8c08eea4e20f1ce408f60fa20a00f5b6
z1ec71c260421d701dd93d46a2eff19aecfcbcfc65a860b2186f1701886da848d46677a07a02aa7
zdecf2af2139c7e667268e98ffdef7496d9dafc428213afbe1267c628de5aba6b4b4ca2d13db011
z3f52d4055d39ecd1d3381dd4b37a11c445ba904750b1c8d5cdb51a7ca70b8ab86e73c4f986f0f5
z9a0fabf0967e8510581c9a7b4d5afa0274ccfffd6e529bcb28d07b39c426b1beb7c361e561869a
zf70782c899b1584f7eaeb0fb944dffe7fe91ee50bfad99454f410781aa8b8a118b7d2e84725e43
z1c29cf71769d1814fb2be2c333cb428ba77840e75f9ab45acaa8260a70752cb07daa9afe729cae
z59b8e956f1dab7957100c3131843600aeeb0c2855f23a854a9746eb280773374d97396c4294bd7
z5d4f699d32e29bba0d68cc6a72cc65ad6a753916a530bd58827f6ba9b80b4cd023346ef3cb96c5
zf0fd24df4793ee592be2534c6a4778b246410137d89e7ae50a2165cf210e92d3579ab77187fec4
zb9e3756861ef05ef30dc601626f3c3db2698bef38e9985f480c614690d822af6e43a0e7429cb0c
zaa99e66c8d6bf4ca3a536cf6439dcda8c426932974453b0491a8620ec333b353c8ca9d6ba8794c
za1a14105ae3ec66e0d4db8228d1c6f3c5c7c722db2270736398ff8622157a744659dd2a38a59ff
zd9913a6ad4f8c1c83a0e8647c3cb3d8f0516dbe90386f75214d69952d231161934d821816bc288
z802efa1a8ca756e1dcb14097e9c048719823d891e3142d4eb2e199c5f70a519930da40e1a92443
z29cc74e0fcd142410289a99cf60abf605c81680ede9d22f707d4db3c19a51346eceee94bafa8d3
za879931c91b3c6917fac166b840e02b135f31431ea1e7db8259c964646194505ce5bdbb0aec8a2
zc318a2fdb50526d75e6db0fed96dca79ea80aa70448d5bb8ccd64dd6663c31efb692f284eed40b
z7d66a76c0c20ac5e7e6ec1ce1c0b0878d30f9b8f314a6fcf749c9bfc00d661b8c00d96e8816e4f
z387ecfe006ed1e505eaa5605a645a163b28d717229b312083be0f8ff86be1b3c31a1f6c247f67a
z4841ec7d9c95d06bb03ffcbb7496a8ea4ab2d6c061df019e21392483541f90e9beacbf6bb4e6c3
z5a4d3a6dcc630952ef4336f6c7dd9e6296feab1bc4d1bea5a20b9f5567e591e1568f667962f324
zb92aeac2ec11c833f84f0447478bfddb70ed2575e9eb70529a44096e68006d5a8c7040291c6e43
zcefe387f0124e656a4ee1f8062c6061c8b229ec0e2d586a64eeaa29f31ed20657b26f7ef0e717c
zecd564666b2a602252efa6ce08759255b1b6ca4641e8688f99d3037b69729ff6a172bc2d1787dc
zd5688b601f5fb2b5b60e6987c720c7aa5232d70ae08c41bfbed6ceddc241955bd5d289fc963608
z7558582975837fd0f5ddcda8e512dba004b7f50378f9106ca2478aeab3ba84a952f5db025fdbb4
z38ed1d0bb90778a409d28ad3400559b4829343aa8547efc83a95f51d7283652617f75610318396
z819f24c463a8fc74101f30d9c6ec250572ed33a35707c9d033f59227c8491dfe1beda4fba22bfa
z6460a4384c18d959742247f6c27180d76754d55e6d1bdf2adae47fb893e3664df9a07528397fd5
zaa99a51d29e1fad9e611c2f055222347b8a46f67fc0c43fac1b5d3adfb5c780842ae2f313306a8
zd7bcc6bee202d214f0dd7d0a8147eabd61ebf2ea7d1e533cc67148eabe50e28c6bcc8f112e2da9
z87fde6b68286cab135961dc5186483cabf5c1d53170483cbb2c16b355ab4010a4287a3e28c978c
zfd1c91818bc31063f4b3208e54cf0a39059ae502bc13f3d49889694b51fd94f50f7f3787c6ad1a
z6d0722a4e9e3ab499f2ab5055c7629319cf508df4340c64a61fb0a987e063befa2c0c742737726
zdd13960b815ac61b4902a8ac7046435d5daa3b631f64d9e7efb16eed7871a6ce99b04d9c530be7
z4755c4e583cd07f5e9839cbdfbb45f956ecb2e99d2d98249388dc352d56d6aa785c960be3df7fe
zcc469d506eb308f8168a4136814269c316f96b7fc22680cf6d4d2465016f5cf5248ed7ed243ee4
z3075107d97b34da45e569498aaeafb5bca0c9bb37bca0f288ba0cb5d767d04ffd4a88cbba573d4
zc49b75dc6fa4b9f88ac5014937112ecaa5cd17ad984f8477e8d5cbf4c14881df61f004aeb1903b
zbe2cc45a5eea896feaec9f0265c1c142a17fd32b705ca0b154d285493ef9eda8765beb745340b6
za3a84650d7eb9f78c46da614e07f85db423ab75b7a740211206c7a415f866155c1d74c8a0a3b7c
zf409005dfbdf399fc3f61dd09b1a760bd04567f9d14fd7c4d51c63e1e9b5f325f900ff396df29c
zaac35645091945a8af16354b5a99ebfde3cdc18d8523e99d12d93052b72fcfca9ade849496b135
z8118e036b277849d85a0cdbd218478941c52bea5744d75a308f0821fb537a2e65dff99e8f54942
z294a4a2a79a968cbddc3b04d0e33f04dcf8cab7f9c25d02f170e39ae27dd229a0837ef09446274
z93f08bc43ae6faf728c538b7c88e47d1fd8d2f38a0776c397fd1cf8d17ac660f5933a75f54038c
z3557392315da5b95abe318e80ca49af6f49855b52dbb34845e265588bd3656db45317bfce1d93f
z931a3b595371c010130f6883037eba49ee39309aa0e45ba5dba55198862b1e9e6eb028035d80f8
z70b58d22330dfa482f85925af59663cf5039387bf3a9ca454df72f05503c24c4160a8e9871cc70
z88dcec13da10832050c17baf74dce2d2075de719f30c1a3d55c97ed027246bfd7c6fe2c10c0b60
z54020062a2078107ef8ffcb8b5823d1d323aa4f6a7353b75b167c57efb4baeba1e2aec547df7ef
zb4c9a9f41ac87bc1acec18b8bfa22dbbc790db1f7bb93c5423cbb42b43116cf196c6871701a32f
z77ca00d05d3ffc8edb7903f41a64b09901afb649f53ce926c2ac5e19c6108f17e5a5efa535adfb
zdc75b0821c6db86e42390240532beccf37f7cdca35cd3ba3c4563d22812edd72e46b758efa2fdc
z23d07c241b49923b0c2cf9631ed1f5c22454b144e5997f8b85ddbb73ec54eadf73032bf40a3065
z671c3441b88a5b80094e53f2f8e93c27060e65faaf8c2c5943a168bb1eb9970d07f637190a98d6
za01045070dd00db079c5cd6c2e383dc9b6c28d12a0fa88441ddbaaaab3aaeecb76953636a24f09
z9e93c65774701f5f95121d840cbb8fac0b6830c059ef80410ca063a0d7d6c58a16a2b16d604836
ze1cee192fc8daa9ccc8eda33baf563e02c43e44c4b7a7706a3720b769c8bf25c32d0cf36afe3b2
z0259be95702d898ba34c0b54ec6ce1e39eae9ed15fcca6e395e9d184972c30c74aa7d111293b4d
zecbf7516507db1b946f0434125ea0a7aee67d4f3df04c6428aa16fe0024c538ec364a2e0e28874
z9c5450ff27b90fb5c47a4333d3f36399176901015424a543ffac6e18c73e882105ef11fea05824
z2ed704ecbdd9aa343bdaa88c6e14faf9ff884cdbf2a799c2f6d05354d1a1902b575acaaa14a49d
zef8399d06f850f268663a02f6ff452adfb9ec52529be4a3db071980908a50cdae6ac389395ef6b
zeec434dc6a0a9c0976938d66b3160af4d867ca3d0ee1df8852711d7dd46d6b4ed77cc1281f253c
zbe8e73df3782097f2f385e1a79351acf4b8bc8a139a0672876045d17705bf4f55ba5ec8afd2f12
z4cf7ed4a456ca749d60a7e1deebf9adf3bd58dae9430bdf87cb548263b81ad14e292feaa3ca01e
ze6d932808a34cdc984b04dfacc44bbf4cb221796f8940729f95d1ee19ed895ee0f44ba9855cdde
zf59b274ea20cae16eb81aa2c170c4a7a040cf695f4fee2b9a84b9fcfce373770518651778d7b86
z9ac51ed2e1d543b729949a2695d54d1830d7cdbd63d669f7c6a52aa8b3753b850f01a59e47a832
z1b896d5cc7cd88b5636f2d8e9dfac516d926e0ec5f3f2da4b47fe3eb6fd921456ca213e81edab7
zb9768cd09a0e9fe7e7107b6c81c0000c1798ef17969e5d907061e16091c827ee7bea8ce7c90a8b
zf1004918778068499cc9d109c70d1b007413f1ae54b0658c4a8594c9429c09efb46e2953453460
z420bd1b1a0f760b06d70d59fafa52b20398fce01cf5fa63224352c5b09bbb6990dec8184f55ad0
z9cd3ae7fa0ae7d44797de91adf51792c7818fbe9613ea780f08f73b24caf354b5287daa81c3f3c
zc9ab1876cc8b8fafce89d2edd4032c7222c866f26857d01f60d4b9e663d4606db1981e16862056
z9e9ff33ada3c97b6f3fe4a698a47b16eb02740c86c74b627c46fc8f848ebb0afe657b6bac79662
zd5d9a7df0ac3a9a9fc2f2d34e6f9f75c6fd2f5086b17de3f7b433ae7c7c06a92958d6f6840b99c
z7f84bac6b2fb9e74cc62c467236da3af6c9049a6fd48b2be465928d3631dfc4a538424af0720ee
za19e8d0772ab98ff79b32d84b6fdc65231733a6ca64834c26800c4a7defee79b10b2f7333db830
zefe5ffb4302926c3188cbdf812f50f36283b5a1aa688d73f4cd8cf37d84fdc89e49b750b31c3fb
za5b6fb4a11317a890c54ccbac5f3e962aa64e3c1f49c5a665199f6ad1b0e6f07c39904afad4658
z580fa3dcaf987e7cfc73249142d84ad211e0faf61609ddd54e14dc6bf2bf52094d8ccdf782571a
zee62e5ad5bfa725e5e6c346980d272e6bc747485d2103e707226f1341307dd0d93e53c75848552
z42b98502791a8a08b87e64ddb2d67a699d2f8d1a4f87568919243ff66f8023122458e49f53d385
z9aa29f010023d1f01211fad3cc115e2d3a49fcb6d3c25ca2e0114cf02e72768ce5013403bd5614
zbd83df25637e8ef0cfb2f6f0380f062fcf2e502f3789a293d31bf14a660b1eb75bdc6906ba58e5
zf199039ce06da3102eda3bf491a6c307a0c9e5906cd2b437b904271eaf39d827eae805783a9240
zb874fc9149046a1983cc46206a049b43e181fdb203693369474799ab80e7fddcb6aca53733e1a6
ze2cc8d8a389489dce560dc1599fe69e75ee2162b8279edf6554e109ff5cb81da00923dc05bcef9
z06a8e34b8771ad7dcf8285cf3aafca5b7942072cd96017cfb770daccc63b749bb52f88545b3ac1
z1d8f62e7f3efd92dd4fa18f879d88932eb2fa189d747b6939eec6c380c6725b729fb674d935aa3
z7984e2d64fb9320ac951e43f2a714236d9efe16f828f690c420d16f5a25e865b02eb3a42cffc6f
z02cd3cf0ccfe44ac94a244f8f283aa34c5a853bdd9427041898838f5e2bd72f515b1e443df7ec1
zc67d4684f0d9f0d233f2841148ed5cbb899a45b7814476940019cfc5f5c8117099a07240228589
zf13a21666a7b187dc6949a38eee01ab5531b44b2822a5b82f9322dba8fa52c74a532dd655cb669
zec1b9bbe3bcf9ae214b8487add25c038bf2add07b304ec35ded4daf5e8fe6abb612ea6e55b8dcb
z53961ba831a02c8a292bd42d3d6bdba5d16cf32e96389cf75b0eaf778d79870f38f1fb5f8e0a81
z92a0169190a7c515f5db5cb6252392baacfe395737455eacaa023d9ed133de7d9e9c2d8b2813ab
z624d5d0a0c1e3fbeb58c8e7b1b56956c1df1b2f75d53f520bbed07008545ecc9552822e4374f32
z9c89d9ce1922b0ee1670cb03353eac991987a418af053a1beb22ca00a919772a3b1521eba338bb
zb478f375a9db309961fc8372939ab2df36a6a0ca5c78bbe7dd1db415ff3e783a5a8506c581a6cb
z4878af1a4c2dbd531d6a6d5aadeb85502b133370701ccbc12f8f6ccfe31254ddeaa76145075eae
z60bd72de9b089e0a6efb87a622f0a8c6d45cbca2c053f06d728597de590faf1ce89bc74d4f6892
z6f6d95e692f7f4b6650b70f3d7b26cd5a3bfa572411a9fe22c7734421e553642ab1badb6d47b94
z734934757eb0c8b2d0f6999cbb5dc8c7b76d502399123fb445e325b7087692e21ddae8b5fe755d
z04383b379c4a4088f28b08ce011249fd61dd4df3fda4cb9fef7290524e8e44517ecbc226dccc73
z330d8ef68b5bf11ab4c4d8ed9c939358a5c7849bd457e78ef7f2764549ff135bf7eb04a8d67e9e
z1073867cd7294b4d196ad3dc76f9e7e27e6c983ffb505e482131f31d4ef49a2d6323835d964291
z49235034127621be02cdc7ec55093ce20d934dfd1f340527040c43378a96c2043985f0cd17e9bf
z101ce5332c445c5b3cc04996af88209f2e74c67d262b6d6844e4d0afdf51990d503eb858771d4f
z3f1fb9287d452d4cf73ccde115bd5304f42d8bf65d92483db05ecbde9c9d9cc8da16670a35c061
zeab67f30337f68b0e0c6b57f02aa39430c4a1e2ff23e845f11e38cb3f0c81f884679424b4f71f6
za5ed531dc5a75e0715b52497b9b5a13c33f8fbbbf1c05c18aa2c31df10dc44db60447de0971341
z3b58d9c2b031e78a4ae43b2dae622e85e1da32a7e3c552ce02c4fa8a56dee0b6d0e1ad69533567
ze669d5417b0ac6495fa1b56a3d1f8e443df6c3012864ed77d40819ee841c553f3d207a252449d9
z051ec790df4a7ceaaa18bff100c37e7e6f25fb07d2fc85f346f3518873a80637a10288df385868
z48e454a14c0bc950d70e5bee4808d2d41876ac3d2988b34d70a389fd14e7c85b55fb94168cfd6e
zcf211bc8f80e8bfc365038fa2f842dcc775143500682a076e7ef0cfbd547255eaef9d1c110b526
z978d108bda674904a69c5e4c1e903f259c46603e53500a43e97b948f1d6c6564b11645eebd5229
z21cf18e47106a58e73a59dbe29202bd5956c423ebccfc8a7b9e4805ada68999d3d09d22aaa4ea8
z0301609aeec0e3743a673affb8d59752301df00a188ea5716ae8e0e6c68a800a693bca023b0d43
z38f66b7d60eaf0433bb599a426503c79cf8696d156e28c6f787cf629de9b2083e8d9bb99e889e7
z69b17a562804b30cb9386673571235e556eab5abe1176221de6e71d1982ac05a51a364b8680cc9
ze359205b2250712d6438f5f87d4cc5d243c9d74149624ae1158a86ac76233d7e30cd13a7bc1507
z5976bc28747d93d1aa11579a40069578848c54fef7e70c8a66b6fbf088c3ca26332f57da96f51a
zb036a1199887d030fb69d5b1f7aa7e6171c1ce7ad1596c0bb5febf65d8fa7964fdf0423b23ca58
z5dffaf831a9c119d2d54b5d25f0c49d2bf084468a3dd8069fd9979002d359ceb1b4b4f86c19a55
z5371c2e1b92eff00c7b262104211399625a7cc93bc70a50081c8bb83ee4fcfaf295e89105956fe
z9801dfab9e4422768b829b0fc8585f616a679e53fbe4bed8e0042455a5921b72dcc0c9153d6c8f
z1fef203a224652164a1917dd5e0f01e2f3a40341ce338a5f23f6b39ce8f90322b7bca187b391e7
z9e9bf38054ef8aa017b33c710dca11342a2cd69742f858add466e23be8832d1ebbf78f7b12aba1
zbdf6dafbfbb102e67d471260a24ea230b951a58c898723d91a1630794feac258667c7b0d4aa1bb
z328fa1f6fd5df4972c1ef51e8f119b64090ccaeef5f3c56eed207414ae7724cb3e221430337c6a
zcfd95ecd60eb8b578b3f04036e41f09f068cb4596c1b2d46ae43e084cc581f2a24309018431d5c
zcf27fe9d0441b301c64e27936ae6883a1eb4c5139f3053ac73cd988f5e9b36ae06eff69bacb01b
za1014269aaf1a7a3c4392ad780cc0ec1de4297ebebe93d5c95d27ee1fe0407fa40dec9b3b509b0
zf5d9c5297b7d808e82068b960cd290441962489ec295890c1093cd2aa2aca0a64155b342014d50
ze01bffcf9d05984eca61ceb4f6cc73c1437f5b4db65706d2e8cc322788c409899a9e96746403b4
ze07c36603b9f982694a3cf58e7457935661ef1b4cee570d2e8047a3c61303abd50ece979a5e78c
z5028eaf7e83636af7fa915fc48ee93d089de51c6e4b5d8261bb607970a01af0764154d4a91cb47
z43dc39761172e6a67a3d1742053a42190572a53d0e9acbcf9f9de60f924d6ee71d235998b626f6
zbc52c48e0d48f4aa0765e7736a4a68b5a12caefa812fd7c589e37a7f3bd43e5f75deddec08541d
z277bf52016c51be0ccee7a247717acbe2e843f573bfb807e1be3f1d6ca2c586aaf687247a74965
z4e5f180b13ba4363919ba877130b1db5c210452cf99a08be820b6f311e741b679ab1a566bd0167
z7ad023885b24366ddf6f2134d2f7a9d89110b3d42396ccd24ce4c9eae9a5bd9169d5eb7a0e550b
zee72a36ed97094dbb13fbea33bfc75a844d992840f5b2a79a51d993faa02ee9819221feb136ce2
z53192ac4139592ea3533faf0bc78ec1c07c701babf0c305dc5cf98bf0a9168dc3aaf77391a6bdd
z909fb110ad64b37cc741a480ffedb406309f017f414a9956757e7a7b2f30f79fc4faa7ad832a4f
z16c58fbb3be6deb61e2e02c2a88dd913d580380973f5fbaa686126ee3c9190e35e5dd10500e1fd
z73d6b4138737fb538b69c8de439ee68d476090ccdabc6bb0384ba217d778a58a68a70d935b8e86
z312dd818b588991368c64df7b24a9a2e78cb27a6e795993b637be6e08b5a88a80f6de7cb58c2ab
z5fbe1f93a2b503bd786834493315b6d3e20908c96413fd16b728e61cc902508b56db39efd06141
zfff4146e989dd0a23754160625d3fe9d51f1e2a161e8dcddcf78daa848d2e40f1a13983e0af617
z98a2977a934fe567e01893562d73c0dc77f0db47590dd14817472063925a845263804cc9590cb3
z91d1cd7832bbcbf813b4c2d630bba817c23fdd398969236bd82dbedbf45dc3feafc9a74e7f0c84
z4b84c599ca6edeb840788258bc781ff76ac9141d5ecac350a838980c1dd2a5c6ab787b505563f1
z008e6f47741198178a30f4a3a59718e11bd84bcc5d1b866c41e9739190ad7ee1c000199728ecca
z7c795bf947d8962d12700eaddde3e53df5de7e279ec0afac74eb92b7424e59f06596e0a1ce89c3
z027e0e81d74f8f350022d78a9d4092fe2c25f2ce6c4e56382291d1abc0c2d1db71d7e465dc8cac
za3d3eed32ec46d350497fb500f680283ffa11582467b37987c9cc4084b2b94d1c100095a38019a
z3bee6194993c651c107a599d97d0b71264606109b356ab7509ce724cf3e372171a1aa3f7a5a443
zd8a9d247962846d41229dadbeea48358901ec0f99e37cc73f78f8c9a066c72decc12f21a28c68f
z5769bcac5d210094df02da868d0bbdb71a0b69c96a2ef546c656db2f77f11864bcb27a39c288a7
zf34759f304aa29fe012b12a42bd8c89dc0ce82a663b7392aa4f735f9dc22a754a9b6b83b10749c
z5b590a16639e1d7c7721791164e64f7e054e4ceecc42477f2cb35188f9c94782f8ddd5ac694b7d
zec97ef52d8beecbe0415b9def01f2ac9028148e7b926a7edabc42fd9b7b1e40871aa3385ee1fb5
z0a328deccb562c65ef0051381d84c3a40ee87f86e653833cc99aa3d02e47c7fd1d6bfe4acd1aa0
zdf947e6854b965ab6c5c6e1baf989f76d5307aa8b7903a173dd96523768d499f4c6080cbf61fd8
zee3cc091466268390555ad3d8df21dddbec83f3ad84301b9d4c91e9e656885f5eb9e8ca2e89717
zab951d04f619bf8bee770d9918ed98acbc1d71c2ad130a8ef85c19b598bfb87833a586186bcf9d
z4ddcc713545c122f01e5fe4e1210e94894022ced63393be6e0ebb6b9698d54825d4f66f2c2a3ed
zc3bf83edf85e4f910ba0f5abd4845ad8b29e4253ccc05737460d0e6a289bbd9beea995fb1185ba
z9b32069d79141e4f8f486522bed7d0724aceb13a32b69c43c5e16c61b4d870debf708f5c69237d
zb266cfeac7a0b063c5f8eb139bd8588e0340b16fb4097ef498b786624b467c98b40acfe45ee2de
z42f040254297f0a8b96abc9317cea25a7d1f0b418ddbc2b75d39ad318832d7a8a0b6d045e9a5f3
z76f56e89726c80e1877bb1f9636d47a6c080c1fd018a2b9da230995c6d84d819e55beb8bd63f02
z09aee058892346a40dbf4b983089f830b9d78fd9ef41801315f235fb235e6c7a3f5e0df48d3ac6
z61e07f111a64002d0f4e50da26a365b6f2c64aa473e7957ccbc0491044ef571dad7d7f86539b85
z5cc91d8d077eba38f819bc5e41e5cb46ac8f5feb857b7732efee9054da92e9aeda4fe7f4803840
z9c39ef1c9402fedd915782cd2a061b920ea94156184709e8da24262d3d89baffe03f2561046135
za90b1724e7946dab02dc49cc738533fc476845fbc8317793114d97c03ffa685732008bc5d6f3b0
z2c82543c6de4e1620de3acd4201fc964f47dc99fb94bb10cc6148c11a1d666f20b3cfe39a559ce
zbe27bfc78653e79502ba227fc55713e3ff4b5abe4ee045d1cda9db33cc623ee0472c6ba9a4ac18
z7faf06c22df4310ae54c5a4a6a3d3952318765d0bee22ba8a10b5a78937e929702c9b462cbb17e
z3370f72e37041dbd5b059893d1d6126b71cb8e5bbc55cc058d0813496d7734421a896f3d44fa0f
z3c2d999c97e34f42aa1ed8bfca06a8d8afaa63c0424af936dc95597e5c774f59e190fda10dc9f5
z5e8efab8a274b3eab8c9c938d39c0f4f32358658396a0a4aa0b93772e4de2a0cefbea631e504d6
z74fea4c6b64530adb2c5a0d2920c808d444ff9cc88e9932536d0972af59f27f63c7c5400c1c863
z2580dd3a33d7cb01c71ad1b251b0770a7295f37c343e22f39391d4104af65f24584baa423828aa
z2c396eec2e48a5fa127cdbfa4a118a9c9ee379ce89a9fcca3f336fd5ef6b2db1758e0a05437e69
z493767ee97338748aad39b664aec9158f62f761af30e22ca25f1f90c08e5ffb6612caf96cd5392
zf8c501dcb446b98d20c4198dcb349a14f6bef20795c38638306820ba2194f6aa12f002ddc0e2bc
z3155a5ba5b5f779076d9ace2e58a89f80829f5b00275a2a7f6e50ce75bc66a94d0e70e8648a27c
ze7f3c6934b73f165abb8414b5ae8376172dac8fb24d962a289586d47a8536e55d944fe683ab111
zf8dde2327b4058fb2348ffdf3023cc48eaf33e0b7152a15d6687cff6707a8c97561e3df0b7b999
z6a4a173e0505716742252d556bd933689efbc126a3b560f48bfac2d43bbeec918e58bb6b63cb25
z8bf013ba0ee6a27055a2c667c221dd73b24f6b7a453ffabde8c12c504d1af074c8c02514e5ccf6
zcd7f6f41b8aabe559df2899e58632bc0d99abeb8a8c8a7f41d4df4f9405e5640658719bdd3b6bb
z26875b26d8b2f737260c7067f6ed1f49d6d45c6fdf650b2fc0cb73f44236f3ac68b1ba26854d3b
ze58639c131f40e8987787a2e329825cb2b1deb2d87afe344656dd359e65a6dd66e2f2a976c9927
z8fc74afc0e05440b800269e260b6d2e4755fb6fd9171d0902a341e20bfe407a1b9bdee050d4cd5
zd251d2bd1d6cc6b2d999346e68c75bf01286616f86bfb2314605263c0f4e1ecc22d13ea07c6e57
z6ac0a10d9f66912ddf08d251852c11e29f8a5bd80d698f8cde769d21ec51561f3c170bcaa59a79
zcc3b821e761b9cf77fbaad778a76dcea6dbc3bd013bc4a728f81867a99fab3c131c4f07e8bf2e5
z91b7cb125c1ad2c456c0445674429c949c4b773a486219016daea8fbc17456406a30fee3443278
z1995f9b66a712e897f6da08a2cddfd624ccf2335534586ea248df5a3045c95ec215b0822b28a7e
z71a3363a05ac5d3faa0be299d3c5d7926b7dc5eb792b3b3e2074d8150dba945d0d7b5149deca72
z85dc669abf9f27afa8ee10e610911f7a7db051b353c8ed435aeb9ac7e1b2206d4a6bead7c47ec2
z38e8131f9e07b3a8b3ec5f55a02e5bc0976c4381a650fce46286f4d1c561bfa4c4db92d140d107
z64a20dd966cc3677f124388dc9fccc2decc90229ce93ba91dd396bc1066f4ae0b97e42fdb25b9c
z50a3caf119b56d41afac7dbc21e94ea19d535c8b697ad185aee2d965332ee1375d4378c4396f5a
z5882d97c6f5597ac269620fe874472f79951d088135e4fd40939f8a8978ba0dbd971d62121a710
zd1bd7b2998d090b7356d006b25211e436c6bacd60b9a11e4ffeee5a9fd4e65fcb736477a8740d6
z1c58ecc0dd8ea58a15a1feab81e0522a3cf97242a26758e0fe820bf0261d96453e0072aa834b70
zdfb8b96bb0cb54cefb160e19ce186add8bc73a78a849d0bed2f33e0a4b52461f7370fbf19f740a
zb96dc7f4cd4489de1dca39a906b280134f6539d70f7a7c536095d51cc0be722744f67af4c74efd
z010437579a966a3e122c2d3b45d8bccce8e130472f08c99782ccbe12fa6c26633e18066c0b1c95
z0e016a89a3a1f7589fb0cc2cbba88e90a42ed188214188ef9c6484866527a1a05d64069efc92e9
z0168d3fc2442629c98b8c36ed8f81ec854f260c599302127448bf391f5e290eacdc934b7aae977
za21ea2fc04b0d604e851b482ef533d54d4be54082e184c68ab62d2c9b929f8f7a65a39d065f9c7
z5fb5ca4dcf21a0aba5f6a51ac8dfc56fe209e726ba77c402bda4d779e064337bb07fb717fefdbb
z17138f2f2915dfaefba50e0d9e9d42554fa3205708a1d90b89de4cfc4acb4972212b06e0634f58
z6a3c2338bc57dd89ba53980a9044ac0e975235a700052e407d50ad9ae7a5394dcdf42c8a3acec4
za03b20c1e8735b54a648fadae04a407cd55913ce6170f249415859433b41d04cba519b8cafb50a
ze2cd59e82bb9ea13cabefcf1bcb18e1a1824f6ddb12ce3a1b32e6ec55f0d84f8ea89736e4fc173
zbf73a28d94b404d2f00a1aace9729933338ecc6c01935cede54457a633e2a6953e877f5ba4862d
zdaa95e83aceba1c81086804aed1b984d8452b5d593a46d52a952bcd822a93338fc155590ca73fc
zf0401d78ab55de071ea73e3e57012e2b59f75c8f0a884a5af39c6d664962ad23a291cded3143b4
z360bbf856fa3d5722a8ac988de6f39962c2492f9269ef7aa4e9e65a1f735e7dcd9c95f89fef4c7
ze99cbe8674774ccc5793b3e6311e1a556bfceb7e50ba490568bc3a051f1d8ebfe5c27b0457b5c3
za95db62a739023e74bbb93bb4416e42a3170a2a77ebed76fa488a9c6003cfaca388cbb12fba55b
z62caa89797f475f2c2a0e1cb0f3838eaee7915e1cfdb45724f2d50ee92b01ba73e71b4ad719ad8
z22759864e9d46f51df53623a0ba3dc148bdabc7df7fddd542bce0fc9f045673f52b890d331960d
z5779a8904c7619bfadeed383baef85c18e1067319f960898c4c8546eeab234c18163649be45dae
zb899163a9cab089a4263df570dfe18233d6e2c35d447736b2859fe2b84df75f037b8825870f0be
ze2a0e28960cadab3f04b0d625888d9571cf1f07908d50c236373fd892952f1b9b9fbd16f91abdc
z48bada32ba02e7ab0c5ac740f2b47f0c13a2553f9d2887f88ff0f83dbea7f51dfb3494f0089057
z432011229547f5f9d9c26ee85b768e612c0c826d6f7302206f883603f5c600449fb0560ba83dff
z4c9b401f15610c60af64a68679a0c499631056af1036c973d3ddd95a5e25ea4e8d226ad114881d
z521fbfe431fff97ff047f0ce56b2f64adc59c5df931d9638c6b2843ce4cc5c9e9b28a5c021c31c
z49c83c7b2c13babdbef8a0e812edb5df250879a2df1376d63a198d366dff7f181882c347e0c9ae
z42a4c0e2fb56f99ee3ecc2ed2b4607c3faa4dea054a6579c04a45f1d30f22d081ef47e5fbcdeec
z17d8cea84ad8a7fb0d3c7c878147718d6239f9f89d38c8d60ffd22ef31bcdc9eab1c167b292a8e
z81ed28a029f21a24ef30a8f7b77f611c70c1bcd5114e0abf4c43fcea621b3b59877d2c7caf4f88
z866d901edb187e41cd8a5e03571d31b90154fd722666a8538cdb344396ee337783cfdf6dc78ee9
z982dd479641b0ecb866297054251d392bf3d5400b82be7796bdc5f3e279519066523bbd983372a
z8ce61635013923bcd8ec07cc1150b6e48a76e4e567838bfdd017001a4b6a524615b3b6ed980c27
z26aba9d8b74f4e8589708f27d0a14662242d380a9514c77fdf61dab2e3e3b4c5ac0ad162629151
z5b804a1308476e6f75b10869a3ec83fea3935637841e7042de81112b8125059f19841322024723
zda3e5e0d2891d4e849c75b68ea143cd93729bbc78d1c5143462b986337b84ddfd5258022cd8dc9
z9db48e8b9c926a3166c2a8925405642e1a125503eec9a85cb756a8b2c848ec30b9c45ca53288b6
zfb5f41262f7a216df5bf2479bd1f93c94f9cc41e78d94d622824094d5e16ef20a156df9b9a8088
zf422e217ff648709f0749b35abeabea5526a450a121a7895806cd73b58b3ef54a7ae8e8f55474f
z907369e497c829da19b5559265a6592e4a7920b54f517bc61e45e0d6892998e40856ded0e193d8
z60e8c09c0ea06dfd9946087f2a7fd18a60281df84ddf67df0c78fb2299527920b3fd1602c61048
zc7774eddce8974814e5c3cf7d79d4b49615aa38c4cf23f4654b4cc990505eedd20833d3f9c063d
z3a6424c6c7966c00234458fa5d0132fc4ae35ba6d5a1dd6f5079ee3d38b9050eb4d955c8db320a
za6400f8de66ec293ae6dad860867459a2849f0c9d155a47c207b396f00276213b10698a5e264f5
z8de4c93f8470c447fd04242fdf1ea94c6f2beb7bfb85f2e11847431289db1f0fee97a366caf8ef
z78d5a757774d500fc8926ebd1dfda4e7d9bce397601e50c083f37a7707090756406aab70630944
za687eb13171d62dd6acb48ef27d9b6427ff3dc9de63efb81889e23cf2faf5ddfb275c03d13670d
zb3998091e29819fcdcb1d9d77fe4f4c90b9e77f9046d706b2743ad8bee3cfc8802febae1b630fe
zc0e46be7692fa891bbf3ab427a4b9e18b2fa67e0e8b475ea2dc0717c9faad1976f4bddb72bea5f
z7fecf865f89536b02f3fdd9a962e91a349c481e0060c11cff61c004a102b9f8b4c97a37f0bb118
z3c5a93db2f5f8eec774d9cd16207b12855ae6c49c51f105ee34e5942100bfd5b30e6a4a1bae26a
z2323858204acf658124a465f65520796c78f14b385dd28a964be798c7b1739991894773d469e23
z41cebec251fcf451cfd9dfd0217349973d263715f38555891f814fe4880ee49631d97118eda268
zbee62a338bfff0449ef8323b0aab5fcbc68e4dadb0e333dbbcb5edf20ea837c4c59f8d1d3a4759
za4b723ece7a47ef107a6b0f688475234bc616541dfbc282d586eed4bc7ec2f1fed17c9c0823eea
zd787757926be7175c54cdaae927a6bc67de9ac9990cb56d60fcaaa42e787957a86e74090465187
z53c13202cf9186c41e6a4d57b54ad9b0215d62950730f6507df9f4f2b0817d4f7944d354a7dd13
z5569114e9db7b85510ed0ee77480153fa9c060442f6c0f8cc5bb70cdecc5bedd1ed4ba46d87d17
zc32ec5f7beda33bec35a8c4c653dc639a9f9e17e9d1fffc674e47522ce89cf38def7c757337972
z59e148666f9bb4f2255daea33fb0e43c6d9531283107f2ac96bc6a34d178edcf3610073e3114ba
z189b36c35e9edfb9f10d7bc0c324d467fbe8491fd3b55890cd806b37cc9576295ab461ffa1f94c
z743526ee92db52516e8b403ff405c0782581eec5a73c680cc933594f540409911a26738aa1ebf2
z007fcc27e337d3c34f0643236dbdbbf3e4cd8db667b7bb956664b26416dc7e1c9faec2c52b8a8d
z892547e86040aa0355ad59a479b1095dd92eb2916b17056267e499693c231ae7c829c541a3ceec
zda067f55bc85d2f362ba4f75aea90483d1f0c60a1ac13df4ab05dcd8539b2c8629a28c08a5b4cf
z0ce6cb2f193f52602f0a6147507565974b0a4c7ffb6f0ce2f8b1b4c4ff8d308393ec94c5b0d0a1
z61ea7e85bc3ef6280b9087d13377d322b8e4c9ec5cad94aa252bd9ed8ec7a59608e8315a1d550d
zfbc72b33660fa7b7a23b7f85553a08239e29a93150920b094033fd88be65fca2632845668de2aa
z6a26dc66d74b0a37207d6faff45550fe60314ba2882fb77a83c51749168744d31236f97d378dd4
zaff2e75861d3c0b547e4107f586cef68922fc184437f6cdd12f4e9a203da3a11cc9295cc4aaa72
z1c42de28010f8fead113eeed1eed65d24caad43995342e1f843ff6ad461ca40f8ee0ef1d8f11ac
zbb52554f36a9eabac82469cd8e59ef21de3272cb48c483f6e23f01cd6ccc53d7fba97c7784d264
zcd057e772a03b26d45bf6084d152bb85984f4c591e3cb7b4999895d60d6f88dbdb496d662e7277
zd8c537d6732c7d8d95320596ccba230551b5d7ea9c0673ba7439ae4626cd88be06a64e49dcb294
zb504c6ac768b24d83b965925a5aa075d30706d374989c9c73e4be9fcd8fee7cacaef64922050f0
z3a3376a363c4304a5e7321c3b6c9190c3c29121bfc99b6dbc957d6ba88095cabef8d3a5c5836dc
zcf8a42196906add9cee90b27b03d9738aa8a8a147307b81cc1066fdbebefd3822f8d952c1d47af
z6fca79096d7610ee9e4c59e44500d4ef8c038e48a4651c984ed6591a4012d03d4de6f07aec8a39
z0fd0f15a9c559436b57053c303e5201c9d38e00ab139da88f4670c891d8503fc3aaf96e233f8e1
z87dd6cefb5ed3e3c5e9ec903a359b0c54b4410660188c7aac0167ebc9e43fac05a7b569f4a6cb2
zeb9965fdb9e302411a1274d5d1b884ae670e466f0cc138bebc34d12b24411b36551d9fe4a19e9e
z2ed34e3e8786fc8aecf4dad3fb5bbde6d38f865f39c8a0d6486afc282a8cf14073ab572c3216bb
z6fcca679d936685b72fcc2c41507ab58699b5fb2f756a7584fd7808a7a1cbad588ef4be7a08d93
zf244eca89e34d3bc36bcc3a7768327efb3648de0d71ea2c4826a4b3d7f27e5eddafc0e0bee9ac7
z1cca5d8cbfeda5553b63761d5bbf49766ae297e4eb93cf274d72d10c8f1852c868a2eb570e25cd
zb424fec54c13497ddb3f8dde823aa84f5d82b380efdb276aa24d5f29bce5e7623992cb4e0fb47c
z4201bc753e58eacafb6a6c11081cf55984608ef773343718fc28c485172bc3bddbeaff88d111f2
z2e220a267df1ef98892471c554f4560018ab5627c77df6b5f2232b3899d3f5f48d414f25ae6b12
z4164cb000fffb96a57023ab6ec9984c817cc38f0c55c158e2b2a7a70e7d455e262d2b56725045f
zf926ec03bb9768cdbf456be13eb7a420236f1565441f468fb98c6a2a16bc13a6a1f6fa551bcf18
zb0efe7dda1fac94b64d5f99ac164efb3f96909b6382dee1c9debc2b457568531f61d549d3f5316
z7f948f7636ab608c63a8fa8e50030ee1fb74a98a8dcc9ff03d6e5dd3532fda505b5b1ffeb89e28
zb693708b34cf0bf031981e366a12fe55f2effb3330c015a9d5b321a3209c6b3925f7cd66827b3a
zea16a033f50581e3287ab2ffbb90ee8902631c9c2781a2b62f8f560dabcc696a714ad85a2094ee
zfa1097b9bd2de84260e8d8cb4b10802cc94d54ea23e0927051f8c30c1c8863f03135d86c5d808e
zc1ead2d04099ed8c25eb739bca936ac28baa6cc801d6a1e07e38bdd0922d32c3a34606f8c6e855
z46c21e99b04c81ca028d9e2064c39d2cdef0f163476dd16129df31e268b8cb75b0ada8e3cbef15
zd6a593ff9237e27fca60a6452d632ef1558c7f138548d5b71163409420e3897448fb27fbdf0311
z43c7563303bb34c13ec77dca1179afadc49a79cdf572def2ba4a7dd5b0a380b6bf374114c699f2
z25f9cbaf7ac83af9869ba3bc78023a808b71e830e037d1bfb1b9fb279c3b64b64258300e48b632
z13f6e9c026205a14f6d80438e9fc270728ab7c51b4819ae36aee1b8fae7e82c84adee6edb0ed75
za2350fce34cc81110577615793bc1291702327d26552671ecc0658d2af573a52388bd23ece3dcb
z702a680b063034e3f398c39ec69bce9bdd0a2eaee4792b89a7a27fe393e8a48739c61d3834be57
zf76de3aea1348c99bf30acd34844cf8b51661f42ed3ab5703eb89679129c40ca731827d0d322e7
zeeea7cde3fe9fe463ccb94211bf26f615a234dfb4d2403adce301844976793d1c67c6ed8df4f05
zaefef0795e5e0f340cbdc86eab71257dfeff1bb7c8319f60c133d9f3e665eb522530af5a76b095
zd26ffbd0915e2c059e99e72dc2033cfe8b28a86a9b1f814d590052b325ff7024a31f1cf9084b80
zb35297a31fe576d76745bf2d439aefb66d27176c7864feff48735e0893ac3c5f369bd3346d7f2c
zbd92cfd3032a40264545b6e7c67209b08fec06bba389d4c0819fcf785b65d46262cafadc170c78
z24bbded782be0a6d3783c740c88f7eecf51b3f90c131bc0834653e7fecd9ea0f3418ecca3c3774
z23dd0c726c11ac9ebaf26b43bff9f131f7b4f104b1008d0b8b448f8ee277d47f29113e18a5dbf2
z6fc4a1376ffa4af32bc0902edc69343a40b495e0a640c3824a21d5a858df330898d741ef409420
z366642a947557fbcb8fbecf149b36c8be7cf607eb3e39bb933aff4098f493153b6a6292ecc4c08
z908bd3cf072dd7030bf3178458f15da0d15da3acd90e595122e0f75834cea017ba614a205d40a1
z66254534084b95f50d76f59db0191541b0c98c8258cedf758af8c55bcac4deccc1937d78cbcd9b
z4854cd3b5a33f7971a0d2439cefffc55555d74d5bb389eb85dcac9add9d07c8c8d6683ce5e24d2
z212a0ac36ad9993ff8880ecdf4f7f9e79658f2c8305526a69aa55eb4c3fd4e63e6b8e4f2a4fe11
za668a37c44ed22b49cc2c520ea540d1bb2d59c3c7fc12e2b458f9e9c86876d425c2556756cce1c
zb584bd6d96a1257481f500194ca77a78ffc44af446e455dd8fd2b24592b628630c8e845fd3707e
z035d6705a928a205f390c82270ebd6cbed83acbfe3fd162b748d081e4823c976dc51f1e6c8e6b7
z39056a40f9766b6bdd652761cf13e7ae15a0d4bc30d871906e4dd765e2a1b0ec23bfe0fc1c7690
ze79b714d5426403203b90d9d4c9ed9f4dca9cb302d4c7d82bba576c22399716c20e6fdd396ed9c
zf660c9f63e6e112950f3bb50896c95583c87ab81a31fcdf14168e6bc398554ad160ecb51309504
z11b2f370143af7d86f98a22d2a08fcf3056c1690d93abcbe9650ab689bf7b0930e01c13fedee5d
z735e43689e2401f43da105899d05456f7ea30807af7b35c480cad074b1d8269bbd0f27dbcdecb4
z201868ab66bae3230ef555a5018661cb166f748254a01ee477d9983438551455744319a7c8a039
z1beb37e3a184934d211808512a8948a05882883f090c26b1a30a04ec5208caae3345f00a76b8d0
z406f38e420a28a55ab7ee8f585228fa511dd8adc52bbb440268d18739e55725ab8d6dfc9329e39
z4d7089297691efc0e047456780eaec2878042e9ae61fd948722714fc035a28a50efbeb7d80dc81
za6c1bd14ba371a1af214b58f2103ebfac3b79c28a6efdbdc2f7d7234a363016c62268652282bbd
z32a72f90887735527a5c864c4b41e8ba31f87270a81cd87a3f36136970eed67d213940dabe4a4c
z9ec5509eedb50bfdbde49a844c237dbaeab76ee17ab189269ee711455e947bc892af13610587a7
ze03db43ed9cb46df64e4cde892ff457419ded5ce943574b44aaf504e482db378d51bf5d4a0c217
za846c659ccefbcc6354aafa74572f742f2df2ca69fb3c7f32c2d9d22b75ef6e4669d5d5319908d
zda581c995a917826413a548f02b26e79ec4aae5678cdd4d5cbb92bda39f493574a04422aeb3594
zd0ef26538a63dfe15297acfdb9db960c9dc89c1025c97ec6ac8b7c124fbec17a44796ab76ad4a2
z9cc8a2b0dc98aec8f3fa89dc31b88426a7d45976b7f225dad5d7117eb65b4e90a19936430277dc
ze6ee21c5e6398728c0cb1c00d6ee603ff113e7c8fcdd15e52cae27fda52522f766dd44efffed10
z4b656846049f417ae3728ff2aeca78917d8504809c3444547fe8ff48dc51a72d52399e3bf17685
z4a4987d382b27796b2a672d9f0506238e0783117034448c81a9cba0e568218db3bffb92178d245
z15f93613366e8b8d993663f96b1215cfcf9221b4df14cd074f35d0d1a610c0993067f119eba42d
zdfb3f0a3b7f07b77ec324bdc52c41aa8a1fc034878cfbecce9c1344004f900cc6dcb61103af1ca
za70c3c4013e47e12b020227952c0ebd5ff93e1bfee9555f5c0ae55bf0f9adc4878c4acf8b41c44
z3ee09b72f590dc80d50d60e5f2060ac51c9bedefcc7b882950e71b9e9beef37af53210aadbb605
z1cd669e43bba2040ced19cf72e6113029eb5d47bf489ebe60e38e926404bf8128e3b69ea48e452
z6d8f48b2a543687acbca7fdde2febc4971cc1fee042cd91f2ddf61c5167472c7f2add19b9d3461
zffa49d7bfd2cb8f03bc3f56796a8442fa28894293193374b4a6fe72bddaeb95e909dd3dc542ecc
zeddfd55fa510eb155f8894bd625bf281cea6b256a5ddb1c3fe525b1c6bddecb15d01fc5a7cd1f7
zb1b6ff1eb1b05adbecb427330110533399a0f750bb2072e0273aa1cd1f154f9b41be5e8d083617
z89fbf2d0c7391ada0b651228dc892912e589f29928c15eaa93555bdd37bee2b03800705e77e7d5
z8b543a264d6df0590b11f22f982a5ccaed1a5ae6b4d283595366c002e48a3c0bd4e73957d28baf
zc0fff799995060e041b6d1e34213918b25fa94393b7a1e1988cf7cfed3e50414d14096ffcfbea2
z92fabf1238c98acf5745937e03c0202b060a23e967f63220a67f2fd24dd53a0b9e514ee0cbc59a
z0fb018dfc4f94ddb002363243738f00836e51931f22e783edf27ff35d95139c00e6742384da220
z6186342fc334bec04f8829b39a24587fe0aa594189f10e4cf2649ee208b8a18ffef3c16b6bb1e6
z036c0a7d9e433abcf0180e2360edb5b953cd683c8282f1683d98e8322763f5d5dbb5df923806f1
z131cb86c6af2b16fbf48df72e273bb960cf49bbbcef3735ca39975ce12952a54d823962e75073c
zf2053388c1dfea2c66c69ae93c1c5246589183874bfce6477692b796d5d7fe86b34c1628577b57
z3664109b405e3909b1c39e6b33de657f7be6b021cbe93c31567906d9b0ee77294cdd7be81dd29d
z2df6af619545cd237c24a58c1fb20c73b02676932b5eade1ac4d7669face993b141daa7f34f005
z43542d9537b2197b78f9c37ade6c51551cdbe1e8a901d888cb1aadc39ebe7c9d6c25ae6d60b276
z1dee33394c55d42c46531ea184ee3c5da6fb528dd17a1eb1ac790696a34b1c6753b24c93d4cf66
zeaaad3aecd017ed2d8764f73659d54b05fe31edb3a13371cf85d59ec95586feaae527728751039
z5f0336b961b82e69be59a6caa23f5339588d7dadc51fb576bc7413cf2a755744aafce41d1a7f0a
zf05eff5c94240146e95525599108c493879bca5156e0223a764efb609d877c84e59b0214d08226
z18fd973b7edacbc4f4cb5403df7ae4307c2795883bbf084625f7bcdc95e599ce369acdd38ce4cb
z8c03df5b77c1cf3a13bd03bd368c2d656b2c2b75ead3ba7cb20da8b6c9d2ccb0aa5926a330fbf5
z1f293d36276e21c06281fa2905d941b49011060a19e2e5d8062b1cb7d9fa4c14df4ba8442b5ab9
z9f9d4ec2d09bb9e66cd92bc21cb7ea43d7ae65c5ea00c8fd2e9cc744fcaf28a9db59d8f749ac36
z148697351e17c648bb996d4317fae409790dfe2cf049a00d8b2acebdbd056f4f50a607f1b14832
zddf7b558731407e4001695e1a7c468671f2f1e3c3a95800e6e6fc735ee9c33732ecb7944b563d2
zd2c7ef2fa33356eb44c4de602063ee756d66254ecd3a35db10315c06a9c172a4d39a69fa6b9409
z1f7de559d8ca1a253237a2c81f62b472643dc998ea32c96ce916768cac0cdd84d91a77d6c456ec
z44903896ef36265c0700d396a858e5884725d79d7ac93f4f34d6fb3cb54b96c1badada898e111f
zd72e7ba41445bd3e4601c72814be8fc9d7e4965ab62ba70be6f99621a33bce56af25b52901f74d
ze377a5af6590d9d5b1858ba0a01a2d670fcfa9f307f09834557d1de18d6c96121f850b45fca2ba
z1ff63f5d5955266d8bd733356f742c344bad2427031d1bb797e8134c1b6abf65c9b31b98dd60b1
z43680fc6786264eceb101fe68d9e57fcca7a4c856dee570436056b0c4badaee8c9b52a112e4421
z5ce327698ede0c7afdb9b620c662288685d1061e968df1d4583402c62a0174765a9972461d938c
z0d826c048877aceae6788736c1dae0e1f87a9acfa41f20690749ad4cc4f44d6723e066d4303625
zf6eb1ca8685c4466dbe721a555b16a5bc29c892676139d9283c9d610427596fe7ebb76d4ff1ff3
z6dc19f84a3b86bfd50e2ab5a951dd6681a57044a83181e03907e9ef8dd5eacf18b4ee47c88468d
z09c85e29e2a29d80d5fb0d183f778fbca7f844a0cb84749547eda1e4e631e07dc65cc4be5ca5c6
z19c000dd2f31261026e3eb89496d75fb51c0943b55bcbd46d9b78edadb676b70e653f1d2b75aaf
z19b1d9b9eab4efd8db744cf089846bcd73466daf8b736ddcbddba786211cc98347ac6ffebdb479
z1a9ea59f7d2cc3c02d25b7594195844422c93b069e2d7dc2d4686a23c402ac280daea359daf5c8
z9fb6223b5627d6fab51aa6accda32f3ffb4ebbc49f33de26cb3d1883b1a1f2d03197890f001f50
z60fa4ebd74ac96ef1459ff42425ee093caedaefda43ca262b630b5e432fecfd5e3d9ff803e6dcd
zfcdf781a932122ad6aaffba1184b011976e37a7dc34bf6de68a23a4a5825babb9ac04cbcd875aa
z9f1f409f2755eb4912a729a83012e9e0d3ba433cbdf71e2d7d6d8b5e29d3dad33406067fe213c9
z8f04c837502ee649ed8469e6b6b3cf2d03dfdded1947d8d9b7715c1189e8d4a4ffb159b40a1465
z6fa46a51cad8ee0b5543165d02093177bc81d2b34d059dc84caec834243ff87c8560b6b9d4e0b9
zd85caa4faa0af0a82256266dc1e76e9c607cdaf9fccc276f993639512c8ee150155ed6caca09bf
z44e62a005eb331a6cd43e4c113bed3765301e64171b746154500dd28c80acb139b6d96a7cdd98e
z4ccedb6af9c1c70bd6b971986b89fa4afb407c934c35dd73f0a17b1d69ca6f602e06f63bf6b934
z61583dccfc576399631f23a203a44c880d7e9ac118967576e685feacef79f6a072ecd651a443eb
ze601297e01b1139c7dd3d4d7ba4bc119c182bb26cd95bc6f516159d5b5073437f6fce2d5425ea9
zc828a778cc34e75ddf42cf00af3d1ebaade76984d7e634aa8814b4b333615603c39f85fbb4bddb
zc3e8a7c48ae7a94a765f34819d7c0f2335f26f08132536f2c1ed5bf8d3f10391301fddcd8a5e38
zf63ac0e2588c2f6d784144ed225a0910d5ac25668b43999dbbf4a6d810f21deec2ce73ba1a6675
z4b3142f0daaa58f4a5f6a958b6196d1a308163bd6f40ae01578ce2e7c9dd6fec43564598ecd98c
ze451d3da148b330959d088c63b27902dc4d53a4260fa92ecbf81a39ebd9223f259059517656508
zc7008b8b89b6566664722fe03c820fb66ee60c65f1cb6d9534abcc526171af081d6005f3889b71
zd6a8aba66e4f37f8a87c1fa1a3dbfc75f752bf1b6d5ac0613b73f9c110cce6a3a7d8fe3757a572
zb3e3cb5f939b6087b863a19965aeb3484edfabd7254ccb82247d09f3bc56346db50431c8a80ea1
z6ffc2f70480da335e153cd0077ac8a8f0d7024aedf04f88102363da9e86ef529e0cffb21b005f7
z9aa0226c6b180b1f52fb0d0ccbbbaa6054c141d66fd9961d6cd5952a04fe1aef592bf778532974
z0d7446c2a649a1b97ca04b6a5cdab193fdd3fde02634b9fd6131f953b8738643c5a7056ace0b36
z095533ae44d9e6d24854d9b6e8aa8c5ab54adcfc0b29cb11df45a77e004fc89eb1450b5760ad92
z1ccaf9af272ab9c302fc5320ed5930b694015773a784d6c72a5b6566ee8fead8fbbd3238a1114c
z999da37a8d135d5814f8b433f5109d49058c10b56286f9e6410664e096026f4a06a087bb9a4536
zd0da66b7417cd70496dc0351ade9bb69d822c224a42819141c9f1ae663f7942bb0c5587b98c8de
zf0b6ff908bf9f31c7cb56007c74609ed0bd6ce46daee4ee4c1f9b30990e10c10023dc90b360ef9
zeae12db7a2a1cb3478b0ffd5220fe006460d4b8aa6917ac4d88af9832bebb0dbf1ece428847e76
z3ec871ec637d02f78edb73acd644fc27e4c22a0a7d3f1258bb7106fbb134a7203b40bad66776cd
z311205797c9722031aada827bd480b694b36e04a50d97abba233bb228ecb772c5f7b397ae29e93
zabdee9896b6dc1c3e35e0b2dbf7cb6f4d1abb1714a3b0b51516d549e3145252e30864df9e8b36b
zc24b1031678b51b44b4c1f3a178b5c22feeb82de12714d5723b34cfc0cf4f35e0149cd8d9fa109
z1630947a045f9abe43e0f7837293e6d1f6d89949f4e08faee3931b6e00e469a6cfbf053831549e
z40dbd648bae4d118bf9a8785311ed2109830b2ae5cd51fa3afa5c840d8acad561da348f37b6e8d
zf6e19712a76e97dc04dc9c8d2c977475933052fb71f24826141566c5ff73dd5160ab188c0cb90f
z926b8d09e45e351297ad80574890611cffb03f13e3b552648df2c67ced916b61073498312bca58
zb7d1ba3c9cb24f5173755bdcf652cd8db2a2a8c66b9732bc1599316a0cb41e235a30f8718fc60e
za1f0871bcdec970a27d22a492b1215a4db431f07b8e0e1308da28b605f7e52a764e950e6cc1491
z3ccba206536b16b74ac2f02c476d2b335a2db1d0e02fb6e24344123a39e36dc899753d175010b6
z22166a44b37646138405c9a018626b70c3975a8d03cb43e0decfffdc40299f5e69e7edae954859
z5f5886063def63dc6ebf1eb97de4c1aace3f7079509699c5844b955377274c78e48a73fbce6961
z8a1728308620dc7c654de6aa058e687bd1888cb83e271b9abb224548373238fff790aabbe3bc06
zcf05cf6c76532d3d51fbd3290aa82b261f3db8553a04b5b89079e2c60cf3085261020b794d23dd
z5891f5a1484c5272b9b312aa9fdd3c0f462d8d29f689bbfabfdc39ac831b935040d3979c3fb826
z6ad31daf1ca37de7d53080504f0aa0c444d2a3e1b663678aea872bc500980d5346f416cce69859
z555e4778d3281b1d0b36f2ed205c1e4564355cd031f5bf0e489f0b0636c2f7c57fe4073af2975f
z262aa400fef9b1e338587a7bb0615eb34ec48bc27765cdf0a99304d1ef953ab27ea1c575b41c44
zce3f6b1e2d7c17546b75621f644e2e584ed58d2da25dc953e7431d346e7ae4aa1ffb0cf9fb62cc
z1f3004f44ec5009ac48d061a0c3596ff8a31bc4145fff1effc62d5cc0887eef166d8331a2d8688
z7f882062896245a0d91425a6003be156b5cbb1e33056ffb8ea62e1850c12de50f9a5462d726d00
za68d7ace6e12d97ac5003c9d8089063fc13792f97f5a6c1e74de22fbe52cf1266de54b5055d342
z27c1eb4102d116428e43924c8f39fed7ba871b2e122010d45827bcef77ad0b73d05019a33ee3ac
z551356b985fa4b5458d300eaf5a3bd46b184b9238da3089934a218cd980ac1a9615935d5a007da
za06475bd1b56346986ed6ee3c4ebcd9631399347670d95c5a6fa1b42ffc29462d020facdcb5967
zf506e265d629185fd47d8596d4348aec0b357e0c34a08e8eeb7a5c2003d3a68fdaa02b6a3e06e1
z95797219ecd0cf7e6f251911253de5da0a8abe6f79ecb09468865787eaa812299c931442034c9b
zc314613a25df77bfb944cb49347a86d8173d32a52b161a61cf81cf7b96c1c6a820cafede38f464
z3cd466a185f895003a360fb21f269b93ae50ffb0c300b711a924108e88ad91168b13078ada9ceb
zf9e4b1e00ce3cc5905a49f0a651c65824f4a8861191f75cc57771563064f6dd56cf6f541309b85
z4ca66a88fa0bd4492623c9126d17f8bc995bea327457c69c56d514a8345635e0e910769f38cc93
z1f998496aa0e231efbcbf078d77cd48ce54b1f5a2c0bc3e89024e1539a8606ff25eef8efd59bb8
zf1e523a7e4e8e3ddd276fd807864acd33edb3e7d6891957c2a084f5e86052e2be5a48dcf1bd085
za67b37db3b431cc7ebf439a612612b1bfb99850e751e1f1259940119467d41b47c599cc7ea1a02
za4d35d1fba6dd8f691928f1d454fdc0e340f6631735cdc2e00ba57005241276cd86da5f226fb5e
z3f8be05b1259c3d039cdbb44b73d570e158d3f29157d21037711a4ad6e02c4f108bd2f9fd4aea3
za4daa30f9265ca1f65b34618cbc3816fa73b8a8ee27bf87c0248f76a8b17c8461f53a81ef98714
z292987eb7b34133c2e9ad5a328432700852298cf66820ed7cc16156802a5b457139e20521d5a83
zc444c0fdbd948f4a74534ab3444ce889edca1b77161ad2064730f390e55a96a3a0198489f949a5
z4f3d2ee3b8edb4537ee93ab8271c63572bb8ace4ac8d1ba60237018ba4624dfb547f4b55355768
zf8bc166907394ffe343c82c2b7726d2c21891b7711a4c117f13ee87c00d3e0ef8e01b26d3aa662
z249d0fb05321f40587ced96b5db51ad361225782b2b11a35b9b428174a5d89fb3a3f68fb7dae66
z8545ca8f2b4435a12a1a3c8dd0c391938308c5b8dcd909ee778834fe94f7cf3634882d6704d593
z4322769e6fdda4f6048c019a7174467d01815d287412ef77f97eb7d7c9ae499572d969bff59e75
z987a7843444c0a4621964b2e382f7fb7c481f2eb606d08c2800bcb2aeb07ccda82ec84f3d10836
zb931ddcb0666abd9285f70eefb963bd84658b7ebff023865ad23ec10b054db1b6ca6b9527b07ea
z7beb02e513d0888d74a0ea81264c0bed21beb1ffa77259d22921b0fc4a20d61429981985c584ac
zba56a9ee5424af27c35ed318d2d1d16e85c608cf0fbed1e95ffc93800fdc485be8fce4fd893363
zb5a0d8ba1887a0c489500c67ce02e20362fdb043abec6ce8c9ccfff41628dc687964b653e82c79
zbda9a29da2600439c7581bc669f282559e144f46a66bc968f7f96539edbb2e570352b3322faf41
za96b980084c0957ba04eb77a194cc3d87c1381a0f054d643881e41ebaf6ce77a99ad1b670b8912
z72d689564fb74c78f64f9ce0e90f2e7b33c582e2684dec7aa3e41e097923d027e6eaff1b401cca
z656f635c7d69355309aefadd48dd374db5f8cc0458fa54da58e411384a339b867e7b4c8c6a63ab
za54a09ba8b804733992838bd934fb9a9d2e068560476c2ad5dc77c11fc6ac881f9ccf4a177bffd
z6041253d94724a9f4c245ad3fcb8f6eb89d20ccb367b8d7b7f60205bd739af3b899eee964a625a
z412632a2e8a045cfb9ca27203da671977cc56274d7a7cfb22b7e6cf164d4f6613a316fa3383a3f
z479a7170ed2e76878d417f5b56bc84b4a76764f0dfd06bd0f5a3e470735d0f23c94b98556a5722
zc3df49941320e5bd0d4b73c0515dba46d58b1d8ce47b321f3e851f137740d10f4d8cd6f53800be
z7f042a7f539204b06b32d9ddb202204e6bd07850b807d2511288b2ed7f391e650b358e63753a16
ze5a8bc2ae256723abe198955ffca6dfd500ab96e347fbc058ae9025ea9efd1e1aef9c85fe0061e
z9e4365cc81a58a1ca44cd902477c570f327c9567d62ff8daff6930b1aa9ea777e42a755d0ae6b5
z12ed339bc54cd6b51f8dbc09b24c25249b3698fde42f8968ebdda2e343e9e3b4c3f3dbd57ccd3d
z01951ea039314ae8daeef034cf043564aa5d33503ec137960f7241a5dd3a691be55412003c7682
zc0015e49ee5a2bc9a145d58a1c25e8887f1ba51cbcfafed460068c25422543d976e35fd2a5fd76
z008a81b2f00ba24358b6a0081afa47c8035991bac1779a7039180f9fdfd3daf2a23bd587ae2f82
z9979ecdafa169456226286d0da071b13d9f7b95dac79e7aadf71708ccf0bf29e5aefbe65abeb42
z220f64928b4f9310337371ad6ebf36a0ec2aa7208896348bee0b2c6d51eddb6f4a2e76176faecf
z943bd548eb0e5e12498a37ee0c407f5655fa718b03f97c9418ea324f01facf7bb5ab0ade7672a5
z09d80ee70cd01658eb857da8f2fae29a93d54208dfed2dbbc1dbf09bb95e4eec4664d6d3882ecd
z726af2d71275145f1e53e232ddd56d393d7c9c5f8f36050b3ade2da234f165ec8d9924df8e421f
zd90db36b7c8d25dbaaede5bf603fb343d87ec05b85a7742e8ea83f3104431b984348655b0bd4d5
z2683fa44956a5309a471d9c5df1c20c574184f1b435f7e190bf7c5769b24af04ccfc45d6c29343
zec3391003eb6b4088476f865ea53264ffcf6456ec82fc8c2067dc31faeee1449edbc6746d647b0
z359c988a738ca3c5166f47c69c2db6424ab053554908bd5bc668ff8c293d4a4eccc74a4973e765
z048828b6f1289277a2bb8094091790d3da1144a16f533091da5b7112d346f82c5814d1b5c8e390
z85124e8888da147ccc3ef718e4e20f3665695f88736ae64cebef6a5cc5f832520ddcdea8eb7d86
z417a4a4d33fbb690bae4aed630037159527476fe6b0c4ac9022a516a74423c886765a0653f18d2
z3cf844452f441a2b5d65dc9a7ce65a0c922a3b585226da1fe40516ff8aa6851f329ebbec0d1788
z30113e1c01ca02631c1fac5bab048499de1991a5eb8aacb914dfa704194c8be923234b269f8c00
z84754c1f617042f1671b540fb592be5fc5503c6f2f993ecae365efcecb42bebf34b14e01bec124
zdc1a3fe05b74ccf6b31c530d3584a1269441ad2fcf22c65b5ee608fb4f6beef0e4993236f64e2b
z97b6317b6a3c9bceb8b9ca5e282ed5570e261d70f76eebe0bd04a6404f8be9a80806c7c3ed4719
zabb0cb94d60f0be4d36b103d7bb50a9de9652775d1bdfbc820d9b4a7b9ec65770022de9e0876a9
zd7feb7e4f36b343b031b6f1d5ea7b816b5b028edeb593f423e3c76896393cc2314a2462b18ed7e
zb9035d921d9e8ad4d7006003d54c99b2c520a7c685592a900995bf383a70b4d7cf32f7fe4a52ba
z052b639e6a5aca4d0f11468d521df93de9b13ed6689e5451e65a7704c018ad83a8bf7df53fde1c
z51094cb1636859921f2710b75c33245618ad327a9e13e1dd13b4906b7e44fe3f85a29bbf531025
z2554e569b1501d2a59e04377e0c3d57ffd47cef52edd4469892be9350e4c349ccd202e98c1f7a4
z866ee84b8ba65ef5453591d7987f2aae50c7f2c2178114d9f785b7449a99734da188e12914a842
zcbeac759ab8ac77e4326340f881a0976aac48a0459556eb1356b3d88ad9d6d7b3dedddd8ab4ce9
zac507df691b435da74242105ed03cb7545bd444519551d193c8fc691fd820e7684378b6a4a9e70
zf21740e168c5f959da7e6a7e74b21d34ebce16a4b2f58e03077f03bac4e110a5bd6c0289355731
zdcd00266e3ee9681e862466d00c6c0e6a17371deb55834708befb76e8aa7e286166f2920f2d5a5
zeff603cb112c6097c99c29259652dc020bae0d19eff0d4c05fda212cc9dd9bc2f215b5ebd4b52d
z77dd4632687c721219cd9195d4a002f369b3af4f3ff9dd23d0d71b0d65493da8ebf92a2a8938ee
zc4b949196806d027e73ec922af163e7a08982ec928bcb8b6d43945f79de0466f33669ad7b7becf
z9da99729f0d0f5f59c329d800d5d61bff75170d103ee702cff143bfbb43b2ea3ae822b741ef0e7
z5c6a49183e7b94decc95920cacf089c98e9fba6bc43e1312abe52934c10d1e3bc7622574ea578f
z48c7b4d55365d58bc2f84848acb7705ce6eb6df6b0c0f07fe120983e42d318777628f2aa45dd6c
z76879ca74c463c771ebe47ffab32d54172727bab16b377c6c8df6839b277098526fd9de48753cc
ze7f2dc1ec894cdc5b80aa35d2c5b41bf5f5012d5d9b8d5edae058d993bdfbbf9b7d99e2315df06
z7f563a04d5c0f5471e8e03a477cf06e1d580c87c392b3a9f0e32311937adea00be00baa0b83863
z40bb59f2f23effe38eae8c8a8457ea8f3e56004966aadb2a93332ce6f7da29279f462af95b74b5
z539ba77886351ceead108b61a7a2fe47da1c4068eeb9af556b9ef8b99a72cd6aa8091955b7021a
z729bcabf76e34468bc1a96d0124bb048f3930c0a6ea373ad98acf6d89c6bce3bffdda13dbafd5a
zb162c278759e036fb1bb3296a4fb67486671a8bd84ff7bf6213fcedcd43415588a8fb6e7b37cb3
zea4c0e67b1a2219b9127c78cbeb91d6b1a36ed46688f56052739a1fc40a2a4888baa2405aedd1b
z83c52c05c8b814fc2fbba84999e70892a68f034ca11502c2fc9d4e2c5b72982f49304c9e0ae9c6
z930f6f903ce27085a80c0e9049a2f1a60ccc913ead7c7cffd465d9454f66741c4d9575e1c93125
zeb8e22ee467f4d2e6d6333804a8ca99c08bc4d42eb7942b4f3e1631e0ff8b1dcf4937b41a55270
z0ba1a64ea39189dc60e6b089f966068e1b087762d68ac4fd47beb48c5170f4a56d3d67b6d82525
zb6d28b1e1aa3edb129da073e0746785b66ea9e5915f38e645d9f32862b4dde1e4e95cab8e24b5a
z7f10ffd2bd49f9e1bf377df2c8c66d388c48d465681e57d989457cfdff331ae10465f4ea40ee1b
zffd4362a92546b235a3db753ea010695a2c093be7feb0955e8c897418c8520430bdc2c29e8ed6f
zffdf2f59ab9e414b682e9e0f7b95c7be20fc0c7acc50c648873d5b842c41ff0c7fa4c9c00e7871
z0aa738a0a65b2fb36cd45d78b9b9e97f0593ff20c856560e9ff8b556a1e4815cef297b49599a48
zcb784a2a324ebf8cc41c10cd53bf49225204e7ce162827b4d8beb84ed5677ba2c990e141352df9
z6f589652c8c8be6bc299fb6369c3ddedcc9097a133fd98667b69e0aca5f2a0da800c6210a628b2
z554f2b659a5b860a6ca003ac8ff98504a2e57a42dda2467e5134d043ca00b332e8ee1ab834e30d
z90862596ddaa9a7a862c10ae03971b07bcd52d3ba3820df15c8452d818810cf09c6827c8652545
zf373384b46bc255981f6b96631123f0559594f23f70585c52a47dc58c5d09ea741b2eb7c44b7f8
z53a81c6d8c37dcabf95cba40fc73f1037684402919beda536bd3c4cd9e787ff2b67ae4ea57cfac
zb9eb0d66edb7626c1c0428b83a021b8375f762c47c4cc3376cbe7b28cfe355bce8cb97244e4bdd
z63249d09a45349c360d1c192c7a37de6a9114a44e57bf673cda78a9a165587ca6d260492ac30d3
z089859fc37f3ec4420c053b9206b914c533fd61c3264d274e0640b911670d701096c204078d1d9
z1bbb673eb83867de34171978dba31789c323e6ad190523ebd037e57fff501353a996db9a2abe3f
z680cb480710a43802895f8d58ffe9cde59f9954755d11940c46f893cdce401d723650f6b4396b2
zab8309c54b094595fddf9595f0ccdcb6f5665e6d6aecb2231555970da7be010152683e66485e40
zc4834ebce1979c9e8fc74e22d0cee4d0c386899ebc0da1a15854a050531a617d30bd88788d43a5
z75ab81f1c7a74011f20e089871fbf113bd4d25341dbe67d250c16302c63ff23378f8517546fe48
za3e5ee924a03ff44bebb0d13d8b2eac4a1cdb8d48eb8600aaa6e89d28c5c25e2991d87d2c361c9
z0ffbe44c1c614f5d19e7120fd49a5e0d8f0c74efecf399253998df7477fe3f3901fd4fe26e0720
z285d6d42ab0bd82fb5a0fb26afd8f111da06f26f2a2b185f1633cdd3c567f2e5a45ef285cddd26
z650e986b956215fba9d92b49a4964172a89baeb84f4a03b2a7d4c043716f513a7d8df74779d137
zb7bae438d2be0819335a35e5cbf8f6980f6799e2cc3f06baaef4c3d8d50db941ee8cab050135b4
z4df42a2c4ddeadda6e5bf07bed9bd8210e9dff413016c23a0a474a4ea8fd76f459a7df022e76a5
z0d49a5e4d0c15dda17d232cb8959cbb70312c17aa952cc8e768cf753988c763b0ecd3468f63dca
zddafc789cfbf42f100634a3faa6f2b4875e8459be6b80eb7354eabf657c567b10ed8e8c71c8492
zae3f86140c7f3965efa741771d8430b2211bfbffb80e7e1d55d99f7bb604bcdb0915a8ed304a38
z3570ce0796817fa0d4d32ee99bec2e160002ddc46d1bf20e42a5b8e3734a7b164c01e835f3a62b
z9bdd7c589676296b8e1e42aeecbcdcde7509a0728a6bb98689937292cab363c09f7858764ca407
z7c3472cd01ded96a56dc575f5234056c8f2158bc847323b4544e37f3bbc5348db3320ed37872c8
z13b84595acb4e626683d9171e7a2a280089a182e0de20044cd432d04f999e2c0a2b0cc82e49f93
ze01bb72e1134babf3dde05e9a75fd2e5887d22bd4f90ca37a3754187d546f81b9e56edb1a067d0
z063c06417da499887e2be57384a9bbb05c801dedaedf7c097ec729d2bf67e7d8ba84b7bf2971ec
za7eeb0b5151e59ecd3d8f8a030e13d9a4e2c5ee539733ce7bf2a17ae613c3563a97c375dd1482a
z8d999e8478c12926af5d00f3cc4899491c3aed3a7acd603385092d221667800a34b1e9cba98c69
ze8540f5720fbeb628c603a60cd36d05fe7c3409118c8244dee395ee7328032234c98ea5203e8d8
z46f351d1021efcb87e1b6a3c06045cba7610d7a0708cad52bffb4a04a9c9deac652a7f79bd664a
z759d55883da3b5c85d41b04bd5b10bcd736ed3a8615e4ff86fb381426e797c894a1fb7ac462fd0
z4798a0eea3acf4147f85ff404ffa3316ad9d9082954b1c0928ecca6581e133523750638cbcc72f
z2a5e344bb290412977948e069c28c18b043ecfedcb7df7682088cfd154be318d8f0ebbf8b702f5
zbf48573020ae2fb6ad4941818809dd935863b857d62254741bf1c1281d88f2b5b5b544fd4587ab
zd79676c4e3117cec684312c2b48a709bef83ecc600cf4cc0e6008e21eb4b4cd4e767010a95e514
z99f834c3d897651247afb57b314044d9999796cd230951301690bab757ad7cdd8da7ab5debd8f1
z512da2f38b495e2320d3188206ec3b03b3ce0af652c1a817bb8cff9e7379bdc5f0b63c348e1549
z0f5202baae3c77ee9dc9ce963f78c0684832c180525f569648eb27ae96f76accaaba7b9d627b17
z754de0b49677b1bd853161839ff9da085ccfb4592cb183c649fde7d88814e034687b60d16bd3c3
z975caac7f3171b1c05fcfc5f4d1062a06630694f503a7f6ebf285b60b9c733c1db22b3a02a27a5
z709c747bc248d18ba22197cb3b128d8fad41e8deb46fa06b056c941a643e64552059e80be5fbbf
za8f96f3c17737153851a127efaa1dc2bc5a3207f0070b4eaf713727b6189f63904796f2a1d8f1e
z869a40c91224c40638cefaebf2379b86a589dad2407fedbb2b6da2eee498ab38fe02d09146c575
z7fb36c3e5746d8defd633487a4a0579fad02e829a717a3a42e06009eacc66f1ef284d4f900909c
z3a89861876e03cb011991bf94ec2b89a9e3e7c9985646b009280b33aef1cde4430dc78c8281a7e
zc72b2a3754e4e1aa6cdac76cd564ac76c0c968d33a02f79e3fc635e2745564b333ec8f41500dee
z0d105f18e7a17b8cd5d0b206d3d9bd725bca372992a760047a3e90ef611779bb9b7ba230868870
z5aa2395c671006edc33be8177f459137d130e3080f290a9faff1d8bebba08c5a155f1f79e1f8fc
zf454a9cecb645488e479c37ec7898ecde6c6141c1aed20d8917c506c33fc8de11080385263e657
zbdf17805e9391f0cedfba05757fd530b6a0a704a32ceb60e9ff31dfbfad091a98afe8fb0186c18
z2f4887ec8356d953458f5742c2f899278c32c2af5dde0065fb58055a84648c711ecff56825e02a
zf17dde2e8f73036e26f91569328ad3dabd0eebdd0d4517eb176daeab48c9e13e578bc1275e2197
zc20dbd7e444dee2322ddd7009012a9a296c02773ca214380e910e26c48b9c2a3a5f8583de52d0f
zc21c49dde644344c8003a2c8273e9b5ff59bdc5979cd30c983cc6ddb059ab68de4713f108d7a14
z390365f3e24cb8e3b20930f3f551e4f3e40cc37415935f9b26cf3790603082e47f4e08df45beee
z2b48f81c014e7724ab8dafd5f35ced3f822652284f2d6e402aef1ea808f696fdc25d50244daf06
zffe3f294c768063621f1e3b889a582c7560783e85b46e13d195a4d2fb83044239427bf5489d91b
zded0cc658e0cb410ee99cebd3b180460654f9b019b5c6ea61d12765e05496bb0dc02a9810b035b
z49be60bfb3474a0b101f1e0625d12a165bb529c4e2e7f21e060ab8e15119c6c5e74893e7b488bf
z4b8932763ba4d4f25cb8cd8989006f13a9b919298a9e8792be83bb0f96526b87b1db3b37385845
z5bf0a8b4b909e90f208e78a8237040cb4cd38fea0142a0b7ae04bd631f5605973023cf9af1e746
z0a6709608abc512c8bd2b29087188febe5015fb2d6d5da4ddae7771d0fda2a4f1e67af9d50b489
z8e91d447694df50c7cf2bf600a20d8937878c36374690811a16f68ca0e1fafaa2bb5316c04534e
z55acbcda63000ce48a740ea98ed9f75c532b6b8b027727e0b5375c2e355674739090ba962266db
zcf6472f95f48c13bc6064aa903b073dc11df13aba276b7b5c1ba83a09bb144511a05c32887f98a
zbe575cfdcf7246b7e64439ad281818d0ad687f80641b480e99ca421e5c2f203bf9bcea108cd363
zd70929d51538c4ac941745ba512ac3d9c3578be09cf68adca791dd7c108fd344efac5911f84d0d
zc4b9dae98334f5101e0e9d24fffc605ee8b5dd86f25c34e099122430286b08a7dea5dc8490390e
zdf50bd9fb16c927445dd37b073d560ab49a441da91df70b8910298ce10abab307abe2aa29029ff
z5f486234a6fd51be345aa0d49ce26cdac2e1d85433c4bf089bd6e011b3a5aa3c0c3907d847833a
zcdcf36db260e4e5005d6580cbecad24304a03eeb17e269b87d75e42149dc9fc349c42809c69d00
z94edbca5cc1e88410d9b8f7d4e016db7939b11ebb67a3552ee9c0eea50e1d87df64edccb61b913
zaccf317cd0fbf69cce872f74f57281698aa88aa4422692f17c8fbbb5b1806efe00cf56952f80ee
zff42cae0423c96d579aad290b0fc0695c1726d1a0c27bb9ad80df6a222225fbc885d5da4905d20
z54088ed3d07555709df7f82a66eaaf550b723cd5d4644d9dae573a2156fa6ec09c855e9ec047e2
ze4283b8297e058f8f0ed67727a17c5dcd512cc81189ec5521c35aebce6502fa3922042a392e969
z143b364020bcf28a8bb656c4e0741eef752eeecd0f0908da4618627affef50a79ca0f7c79a1059
zdf37383a5ba1a852203e22b96cc773596baa3df2b422fd47a1445220525bd6dffac28593a13329
zb1e248a976fe8f206e98e0a193417a3e6750532af002caafbfe16fcdc4566c1633090b6b46144c
z2b4e3aec3b79ce279d19487f3f12cc490a42ae407d1792a89117edf41e871517f1a85c61e2ed5d
z738ec08c35e4424dd893c738846882af0e73f67ea04191d80e8c1702c89aae63b2102cf5a590bc
z27c35b207c3c41c750998dfe9f834be447a13d5e4c7f3e73e6075785d05bb091dee234858f8ac5
z996eb7dd95aab223f66b48df3dd5ebdb7d778e90712771be11de3819d0bf0d81595a8a10c2d1be
zcf6cfeee26db99b72f651a3d88011ec0fb54ae1b11fa35f586bd824596ea889a354f51b88e8a4d
za7470140fe64b0d13fd7725314da49ac2c5ef907e23cae152e654ec5e4b8be3012eeecc430ced1
zd34f752cc3cb3cb4eb6500c82099954912550b81d9fcef163182bc851687495ffb97cde2bac463
zad5d57ef449ddc1bfb371e7c5b2b12fbd406fe185b215682bb652d4f4327cb690ab11418f7f8fa
z8ee5877adfe9473d9a5eb9b75f0f6b3eba6794022c23fcb7b187d44b56e9f98c0e90b63641d48d
z3071099346de5163d1d1baeba3f119884a7abea5436d07dc7fea198d17db6122eabac4244ad3a0
zc1fee0dd3c470f93bfbc0125365f4a560488601aaff9f8d7f782e8113019e3679d4e2eef4c1106
z74df2e8c0deb75b7fac7336a12bb44085435ad4e5bf8645fea0cf14a3892a64e994bb2b705a2e3
z56c5edf72419dd290c678423774e7d162899cd9ff9d46062d983124b3a1602684cf3b7b68c1285
z7ebcf21a75e18a0389e72397f36e39d9ce2709fe369e1afcdf1ecc526708c69f62a84187541ca6
zbb291f9571eb1cc34037afb7eccbf58dd2cc8168ad31dfb17dc3a3daca26f4a5ad4aaf7e80ca60
z56d7d90d6d9af7ebacb9797da08bb323fc08d3535a15aa46b54cebf0c54a8a4768205f3b13c3a2
zf7d814b6483670f104909a98639166818d890fcde25e0e6cf7370b669bf577f4a00075be97a74c
zbe4e0c6b1a5134cd865b7b2db24b20a01657f15e3cac7225fd27d5eeba4661ecfc22312c0cc195
z6f91c50b3bc4167fbe9f12857df31b359993a3929af132f2efe46496667bf54388764e8df0d44c
zb6169cded9031dd7bf35acffcc0761785f24a9555a6e82ee085c934595e77fc6511fca963453b7
z4ba69930c579a5e2a22d6b4b6311edd116126b5b156d0d691e8809f626c80242273f2cfde91ad2
z1c6ab4b2639579a320e31fa50d640f3747ccb18843c7f52cf444d228da50ade40c952f846cd0d3
zd9e4a12571df544827673864f92e3d49d604257b1a4cdfdfd3b51be2c361aed863f150454c0d1a
z911de4c02dba8b9903a08057801567ae7cf94046973edc7e3a05a91aedd6bcaa640b6f13d90e2c
z12971b9c8485ca521fab05cf8b27481b6ceef8f7e4ef1e89ddb3d8f202b7fc45af3441cdd76de7
z5e1c80d480b71d63af0a638bd680ded3217178195e5947aa266692601a8f3a47b449a681b28769
zb8702886f2057987624ea2c526d1db4afcd4f454e3fbb6273e77f200a0eaa7e103abca1595fb8b
z845f0351ad5e3f95a647426291e26bfbc784d47fb45b4585823755b22b698de3745670f2803509
z985a7346081aa8bf16acb932f0de3abcc30d5272996c4789e448723134ebc804c1b4223c030729
z3c05dbadc6c005f88e475b242942896a53021a1efac0cacc17935c20499653dfb228fa7c66b943
z9fbed2331e91946ca7a6759d3fbf9112d42ae5d771078b34f8b87275e41f7e312d4fc68a50f73c
z7db8318abae27681e312ff2d824aaf882b2c1a48b1a915b8d3be96abfc585870ec35791db29330
zec222f2afb2e50bb35cadd8a0a53df086975f80b6d2a22c577eaa31cd07cd837d2728ba07d58f5
z9c861a6e6e79a140203d18fb9a044fea929e1937fdff3dcff07188d3ea2f9c81960c9924fde9c3
za992ef10153d08b2b1577d26d2dcd7d0040c74a6ebcbd2d0c5dbe4106bf788a4d25abea14145f7
z4de5f06269972731dece624258f3eea2a47fb5340b09abfca8a37efb68625d652bcbdf9c5a94f9
z738d8cd7c35d92f2dc631b29e4b12f89a1cae5fd2846bf794d1d617a99237b0bea402deb1537fc
z5b73f4e2f5ad2f8a097eb9a9e4a83d72a65fad4ead4b7df18402c831a18c7ea74e576e1955ab78
z71b6d9b640883a09bbfcef1ec17b742fb1a0234e64f3bb81ac3c126dd3dfabe45859aa6e5fafb7
zae3caa9bcab7cd558bcc30be7dd7980a1fb8bda53ad0587cfef773f48b492b66aee7876ba5ad44
zf1a20bb1d2888918f4b5237387bd00a9e8285b24a0d1e3c84dbe4a09417644806e1ab23c4b3fc9
z2eb67b98076b91e1dd75076f6ba60d9edfdbd7b10a5c127f3816c328f3a5ffcf3176413135b5bc
z9fe4e2d75b1720dba90783b30ac7c88586b7b1b1cf48b8d078b4a6991db629bfa271797f1c44bb
zb1378eefb869bc7f04d62453c2dcb9f17f0912379f61a7b24c1c277b4af71b3471a30733510b33
zcbba76a11d44cccc9317e1bfed74a5044c3407f42f302c04478b4433204dad2c3670a8790f8357
z7dd8d409b8be8583029d7f1d2f1ee5f64baa01e29451cb2842988a711366079a3ca5514ad611b6
z8d579f7a16507c6f21c1265ba89c0e8e925f8137b257dc7b24370d9561af04eec73adaa2371c7f
zfb8f044573a58bca21750521802e8b5987c798175053d2bd4c8767e915f7035ccc5eb55e00b0de
z76041d2ca32d8bb7d6c70fe7292cb23e8cc14b6872365fceeffd1459b12fb3f0f35b25e66fe8ed
za9b1f2524dc48ce9dd622ae33541de569cd34b1c0eabd449c9a2d966755a3d70af88474dcf03f0
zf356d7fed72c6bb05394aa660af401d41c11a2dfb917049df67fed9895dbe31fa5055b55f35e9e
z141601daf774be66474c44638e86b858cda2c8ca87f9a7aacb9f7acd2e7ceb2e3f571cd83c0cb8
z7350e8ef76f10278fa8acee146a2e1a44d77a09a7f970e6e4976fb59091b1bd79374c594586111
z7f24c2fd7ddea01ed41b5266ac40b81f71997ab909cad09e3de6c6b2b247be8e5a2aacbb9dcacd
z4cbe1222d9b8eaff6f6bd3b9e04730e464da80d8915807212278871162bdd3af2556355702626d
z1e32ed77b9b806ae495d28f7f294ab301f9f98b572a09c0464a8c1dfc2df848ebb5fc433b48918
zb85674e81216a54a59ccc7065758719a9b3bc058c7ad610679d89567651d7cc3c7a5bb8a013695
z5946f319ec0eea6e0b6693aa0cbf786678efd1cc862ccd8d13f311a0b04ec268a013821820fb95
z9411c0c47d19fda421a77fae27dbca687cb13435c34bc8c009bfcfe785f18036920cbe31a06bf3
zb13a9cc771624ce42e6a91f0a59c75386c77a75ec6b2e705c6c422a580464e042d68a4d8de0bcc
z3404d2aaa502d66d4c188c8803cfd9c6cc7a80b7ca08250174416afdbe29ac5ec5787991fe1e80
z22718d470dfb8b16e7a503add283427c036072787ff9e7612d6e846e4407e5ce720bf05bc95c64
zbe78ddee818eabdcb819bfde9613b4dc54cbacb0353cafa1ce05d9bf5c42e2004cfb92e02c71b6
z6fbdf590a3173be1320251aef2c3caacdb7428d68de7c178e03f1668655247cdf4062e6cfa80a1
zc6f91a4c38a0aff4fdac1e0c6c651fab18426533d40abc1fb12e3a931ce677399e2d3dc254c2f8
z8da7c6b94717c4ea24d56e09330a1ee56f33859dfaed5a44fd4b436f935626cdaa0f912758cd9d
z119ac97866d14f61a35ba1570d978028674ad1502715f4984040319c97bba4e72dee5ccc387a2f
z6bd171f0bf37a59ce2c1ee14c9f6afc6d3d35b24b0789d43eee95c9ba6a64bef6bd4a1ceb313eb
z5d92f9e8618603564ca3d3b4b7d3c5117a5c298366305a5054f184584833900943758a11f7d486
zdddd8ffcac3a2cfc41fadfe36a3a0815f522cec48004b1963b49070fae591cc062aa17de7aadd2
z09392e6b434cfe7f39461b8f61ce953eb0987cec55446348c1f24d94be6dd36545e823d660b29b
z25ef65de5e9829459980664e57c1dda01405a0729d2da2f684d0b4e82b399ee1957a27728306ef
z7c16bf208b75cf6d00c46c407aebe3e73364a5c93e4d970db68c12868e23e540b1eab1bb6ab88e
z858a3699255e1f61986cdba2d97b4f807a62dbf21726791bf603430326cb161c9d5172f971169e
z3c3b3d4d94e99f0cc7aae8302545d1dabec72aa9bd892a543e6a99e686eca6e0a987d13b5c6bf2
zee05847d929ac5859a187cb34cd5f980dab15f95fe50ef307caf12c52369c80be7cfe5a7c366ff
z23ae62f39fbc9253106caeb3f48442327f150badf9be90774a679b38955d7c4c9a0fc77d285887
z28a4ff4ffc31eb32b4db5969dde7312cf740fc7a9916062061645f89941108fa91ccfb366d3706
zb832dbaa9318c7e408848f58ed127ac5a35e987af0e62368ae76b21203fed6a95271651b8e22a1
z0ba675d5bc838e286edae48eda87319bae3c1791d1baaa8623ada3beeb7aa4903608da3070f7b8
zcea0e209022e606de805585bf29f6a2c3fc675ab52de40b2bf94041536befa08f185afbc632db5
z8979cd6124469fc13e42ba1374d030cbac7cf8120b9934d878a8ae44fd45d762ddb1e77ed5c0bd
zecfcb3655b660aef92f18279fc7b754f1bc7eb2122d4f1db0abbf5f9a478c6e4818e855a4438be
zafef7732a04b139efe09e6dadce715772ca575d42645c266d041e7d4bec066490344788f809d3d
zbcdad547c8fb3cb5a9d25844ce8f771eb7f3a594b0272647196a96282e72e52df670ffe69d283a
zb466695a774f22c7ecc4e262a02bbea6c02dda70568f32de0ad6a26b05a4deab476ae001ebb77a
z5d125cc98f0bf601407e8963daf090c67f09014907ce5e0ac5371dfeec6e374ab3832435c11268
zfe84ca1145744e2b96b78b6aad15d0c922865f7eaf5fda9ce8a4832563b435fcd1d6e9b1b005a0
zc1b2fbbf13ec90d18d90216ef79e37d504256a4f3bdb85e9780a564baf1ec80e6838856aa356f9
za73d51e4c2d008dfc19572bdd58d3848858eacc17015cdc7c42451875c0db5883cc1a1e2d2573c
z59d5ab817c1ee3048ddd4d885a1d3fc983df3d1a5548eac2ee46cb44fe516eb3a4dba15ab8bff6
zbc2f5ba2262eae1fdcad7375f872664d008a7791cb0b8df2d748f449a006f290640895c661395b
z640fd3d54df509d18902e142cc3976ef9dbb17b13cf77a44da6fa073a70c1307e66b94cce91e11
zf6893cfd181bd01e56955da3c68943aa1d1b229386a44fe5c11d75297093a324282165e5026b04
z8174b4ae3f4cd4e9fd6f3d3d964957009fe2ff4f199ce485248d521299364ae162410d55e46f74
zae0d71ed8a49c12d279b47b4fb32e1fb94b2eacd8db62654da8698ae8f600832a7721731b7154f
z01f5f2e77f699e7104599994dceed6a7d9b867328dd7440a580e33209cd4b913dbe71f1e8cea87
zbc1f867d8ce2ade9a5b16d7018127d8b3ce40131ae26f33e1b8748f4d68916484ba384273ae61b
zd2513db452321d309804b45df76c61b49664a56e33eb6bfad3f6b53353320a2948cb833f32b6cf
z79f4ed94463de5da5fe0c247911649011c98056390cd7d62bb347b28eb852d24c2ddc72e477276
z73b9c34e35a784026080ce4ab718309e1a9dd860d0292a7f5f8e9f86d621b294a6ffb7f1549264
zf603322d2d7e7f4e4aa522c858fe46589a34d76eb81773529b4ed969b93614827f2ed03f9a9f25
zd620367bf3df6a4f2a117f9cb1185efbfaf24e547965f74d4d6d14b66582de90140594a62cf4e6
z47f246a067ea38411ea93d04adbd0d7ef7c605b3ca4b51e47ee504c78972bda509d93e207392f1
ze2852f8346af420159a24681da1ac4f81750dd39834d2674064cd83186776211f731d58de44267
z93e4e828c2a74c1b04746e716b3620019346cf84a260372e4e5ed9956f728c3bbf18786add1a47
z6ff8d2745d779e3f1227e3a4ce83d5353f350efb18a65eb0289346bd2b4ef8206080f9b1a072b9
z9f5e1f4e0e309f2bce69932ecaaf501b7f6253dce9fc5187917a649027e8c98211e9d0c05d5f04
z0a0d8e259454600e956a34e4b1c7096156909f22a8734c5602393f8740101fdef8f0dedd44ae8e
z0c401922bbb75a2905b10e1c7fa915ef548c2b38272798a912688d45ce9a4747bb64062f0958db
zb299f7f6ca0f535c892b691e8da9a385fa39e48f33644fea7a116bf01ab6d51765727925fd5913
zf667f03c7feea0b7077bc0723848e96abd684d8d4ac0264aa268875f103c1638323bf07eaad839
zab47a73bed77ce6c14fc8d3c9099102151157fb83736045d96afeefad0be36e9c2df73d8cb499c
z9be208d4b5396da1dafd627d4440689d13f90e94849102e1a9f52c74145f59598709d7c58e20ed
zb513c7d7de90e7c8dc60f31aa6641f484bea65acb15a68b529fa3f713b37ea39a664958a4c4e25
zdb9f72214470e04a5091f88a1a31ef74d92da1396e65901971c9098a7a4d0454001c4472ad8613
zdff182a44f30f8271a40cfce9d41b4a83d86ad8c20735ef2b576fff4e9212601920c436d28a148
zef01050f24042459b128fcec61eb48deb6eee9c575cc1de10b6cd991919e3efbfbb9c3395d5e09
zbbacf5d07fed313a2c549a5964af27315a00cc7f6adaa58685b87a2854e7991cfc4d248c40c320
z95b2895691aece6aed31ef0f35c2a00212c6de6551fd17c92c25e344f5a06b40a2e8009e4ec2f8
zfec3fe9068a714b23ca5a91efabb6fcc18e564563da26039545012b8f98a388e0ab6c2b6c98bd4
zc71fc0aebfa91881ca7a5755e6f534b2c3cd249d8d72802141a7ef17446433b3e9fc837a414c70
z01ddcb93ab9eb15dba7570422718e691b77100f8c35242a90318000e792640c83d11f1ab079a64
z08b668c14f0e2cf962ea72025c8d94695be8296f5ce9f708505d812e84f4637ed6385ca6ea4d98
z94fbe87a5ad1cbc9d795a39c7475305a975aaf9a7462dd72f8efff8e0083ee8cd8e0dd2b9187d8
z3f4a028be1874416af6776421591325d97f17df1a56e7324f54eb374f1fffd31a818b599877b60
z22ab5e908d26fd006361943315f597595329f9690f67a7f0c68d90fc3aca71bd60852fd5b9caef
z6be010cdbedd6dbbb263c7a7f376db69271043f00fb0722f810e9e4c8fc9de74827c35abc3f6e8
z23c0eb8765cbbc4bd22cfeff922f0c4050b85a4a8e7d0a6a18f68f1bcbb76b3f69dc7e6a09e6d4
z41e38ee70ff132196b94fa85043c7ec50da06b82d49035f701e7ca5f94223117ccec533bcbc400
zb70040ce5787e10a87c443cdba083ec8b4dc067a70eef5bb7ee68a5d6939fb586a0784b1fd42b3
z32bbbec61a2059e55738a5fbf9f05a83d968ba514ec4c7b903757613b3bb6aaee0471c528607b0
za3e527517b51932998f71d1be697da0640487e1ea477c6dfe06f7805dcd8a0254a0e7b8fccb88c
z4be0dec960e563e11e6c57473be2072c1f85af1331eddac61f90d21c1de96f860ecdf556329eeb
z3f5f2495da483292fd5befe6837818a18fe0db8366baf23ce80743f708b0cdd6923f6f438016e8
z8f0f3034bdca002ffe4b77da659c1df131d58467d712201053f0db9533079bc7fdbece3010a44d
z083aff411d5c132ef1d4dfb3458301d59ad954c6eb92ed4004b6c9f445fc805069197c66e3ee71
z1f721917feb9cd2605f3fb128b449e42e34d1658b8361e823f1fc1acacb72cedd5c6c20564012f
z901147d6daa6ddfd68868ec194b15007fd02ba1eea27a648084d49b2eca220b5a9ae6f5a69859b
z36e4cb9fe6361d9b505b61dcfbbb246bb3687847b5b057d4f5338dc39325a085febb6c49e47190
z49d1fc93fa1ca570b605bbbb3844471133c535ba7b496a8dead8176a3d1622e1e2c35f02110b44
z1dd74bd590f16fcacd55b85bf5b995aaef43e5118fee523d21ab294ba2887d83463c08d3525c07
zbede450316053477dc2174a340b367d4cd4346a4a2ce5fcef3b77f487a074514687de49ac0ab77
zbc359e6f668fa83d2a73ee6a32de0b2b8c9d869cc55df89a0f82a1b5dce0f14c4b558102989389
z4ee4594bb837410f18c45fc8991b4c8a19b91c8f1822c06d7842a61961c05689cc540bed92ac58
zc5f225409073307377cbcb71c7f5c89dae7d012d5910abbc6220680075b317923977942a93e280
z6448fc59a7aa89fab57f8ea72050dbe666d8b14583ea8544070d11726bc762709c805fe13795ba
zae51a189854b5213499fca3a51606f307c72647de30b2ebf9b430d73b174e77d21de4896ae202d
z47acee5f1861be9b92a581c0ad221a759ee9d33c8890831dc7b8a933f8f4a751a6c6dacd7cb729
ze0436752450b43b920453ef40015a9d1619e87e3fc8324c3aa3e0896ef7eedd4402a35b659ba4c
zc9493284fd7fe2be76ceb51f91648c0538673e54e94e7180d9901328f02683002b1e900f2dbe75
z09d01a211ebf92ae738942e938e16787fde27e4c9437a3fbd85c15558c3869bafc56591a80b88d
z9143899a16446b0bb3c073f4c1e435d4495bfba9c311ff7f097cfda568a144dc2136b749cf2173
z23b1bb44651b91fccf2219c50a56708d2ec370842e3ea236f7ece12672ea584eeda62737c38faf
z7398c0f6c720ff27c3ad5dcf500f7d91f3c98bb85e014b31db15084e6e20f559f654ca239c03ba
z206874cc3692600864219651d7cd87543286a85f3a4918781f4e53fa21ab87804738ddc8586b4e
ze3fa8f807975a6263f30db76520ee0a007dc9dc5ba9eece2257ba8b07c87bdf6351d348a54f6e5
z9e03bd63d150911f7b511c67071d672ca17b639f6e291317f5b1c79c427d70667cb213bc9cc946
z1b94d9402dc61fc340bbd40d3e6579ee7181062ede20b1b25118c28d4abbf63453957ea5c27f43
zf00d91df1ea71c01284078d4a915699f2d7f0688d41e62122266a0e8f7f71604279e1a2e878eae
z32f20e160a00178a80b0a40b33538338ce30083a90be5dbd27b95d95e80ea432676de1fe314ede
zd77a84bbd9c070ddb0b0fa59d24b0281d016c1fdf95f6a3b9e553d4a7ae7fe6bb6ceda92cb2a9b
z9fee1f6b4ded3c20f70ae2ba41f82b522ecdee50e4c5af8369c2ea66143784bb09727a4a013a8f
z1be54727a6711ee9495e2ba3bb5d99cae3756b1b998f92b93f7f483a97c934df188255d293a034
z31500182edd42c3bc3f418a89b4b5048afa2418cb64920be935c125eea669cadac378d3295578b
z3c118f93d93a7c88ae05bae5f2f1338266087ed630b82e691d0ecf4c14a569442e30f98d162c8f
zd8a7f7e057b51b4ddaa2ad5c5a1269b42801765cfbce7bcbad88aa45563ab0ef28a8a447b04519
zedd3b219e35a5b2f6a1c66650ce6efba6b5bd542104ec0baefa497fef13afa9f82df73cd4b6d77
z24395d3aad902fa31c257d35c3965d330cff78e71c4c20338db97b482f1b30be83fe3d69d03724
z270cb744058172474a27350ae7341d991f14370d9e5ce43e7fbd061c543ffe563f81573cf2c763
z72d5f686b61754e5914856239aac18061050b0e8886daacbee6d1fafb13416228e2a9acabb0391
z5a9d7ac818fab7488ef3cb1c3779ec0d999e79ceed92052aa490a30e21ecc0ace9f7596a4790a7
zd82a12f85d8bcf48dcffc3ca40d4acfdd5357a019ecc74b8817d64be839f844ab205ce9c078680
z093ecc7290f7f09f203009411af7e1b26a1b9772b762fac8c85cbaef806697cd59d93d4514edee
zd40e1d6f441d6c0518a25ecc35b9b516a405c33eee17064b0d2fcc700640499ff399c55028eb4e
z776c47f83cbe1e722dbfb81773414c07789c3f6c305d1e8d5db039da34054e9fc31168cb1c1b10
zaada1bbecea0cf17dca6773224986c8c238d77d9c06565127be338442b8de193dbeb5872c0bacc
zc2400d2859e7540de2ed8ae49bfc3fa48e4f7ea50dfbfcacf1db13211943085335878899458d47
zb8636f706443b60f2717394048ee06e018d812b5ee62c6de6c07f3e31ded5819529b2ed68bc0b2
z324701070bfd924f4f351b732cc2e10795d60e96de94b52d6ea4a9b6172597a935a86d37817110
zef72f8773979ca894f73ccd96358659e4c0f9a5201069767358cbbeacb6ebde27881bad236cfa3
zbff11a8ad76c85a97f16e7188e9bad30a0fde2a8f0f906678cdfbd7dabc36ae4b9dc6974deee3e
zde7bd01ea7698f0887d294790fad667c858b12c8c3cbe497da236e1e23143272da2dcffb0b4dc1
zb97267604e6a2cf00cc464f27d01fdcbac3d2a93cc6fb1a5f183bdc69dfc9346dfdb46d8f6f0d0
z5809dfafbd9947f2d942baddd11468a43077f6094ea00435e1a8a863d176a6b742a8e25083b136
zde9b1f925e3f9f936da26d726e1c809c4293e1617d38f2fbaeacd9282a82e60ecee3825503dd0c
zb5fcdf2de7443f78a36f47c58829367d944d41a787534d22b04b674ecb321388eae3cbe32cf55b
zc10ef4bc12ebbdeb31396139ffa955719cc6f7c3d05f7194928caaacc6967ba3883a1f28c5b6c4
z17d3ce90007ef5510eb90c9b84831d0fd70adb7f01e0de18b2204b578f59956bceb14ce13168e3
z4f0426bb2d8f3319eb22b078050eaff233a1af7fdc652581259d3374fe4431a21f035885e7f863
z6b256df40f8ab55b92475794433c6736c7354199b7a9b39ced74494845418383f1a567392ac0ea
z32534115a75bf2f655652669a6bf022cd59e5858e871654480453e632b76c4868119c435945f18
zb5eb9ca32e0e9b3d0edf1a2a35a720bcbff569596d6e3169ffd9f41ee612cc1ba0d214bd4472b4
z8d240ed0c3ad4522d525c2ed9f3f7349724b0295258f002e4902300086d71bc4ec5125820030b2
zc3320c2fd87ac59ca6918ccf84fb98fcb4ded3e4a86e8731bc9540df794aefbe7bb49df2d0b57c
zd85ec1d69e5f68757a7d40653a08721d4c60e67714aacde1e07a663cc14da50bf57ddadf4b2f6d
z8950018e767a544cebb5fbd73d4d39b81c36f8bff203b0863b9eab6622da7f5e2ef24f766e77e5
ze66f21ee8da1d7bbf3af3a176b6272b4f442ef7d8eb4935a576bd6942cda256cbe5438a728a4c2
z67f9073d8f77dab23be4aa39035174228e4fa8fbc1dc363da93d08dea61464a9f4658b52159e06
z982e86a2574d5b6330526c2450444a0e158b261be7bf615d9941126853b17f85d722aa2fe5d183
z2f211df1a4af46148739a0b31f3889688ec37fcfe24dfe85620d958462e80f558bfdf4a2d0019e
z5934e3783e644b77f5d6dcc644d0b6e1e85117690af725bf1d9850379566176162eb8c428f1103
za06ec9ee594cb74ba6f28b3f086d3bae31451d8aad0c5e795f368c6786166b455bb5979f513bd9
z260642296e6c82b496ef0a0547ebb27ba903457d9b29516f883223ff08bf2774764cb263d42042
z751b48928767532e89eb06bf13d522c616c68ffc9a2315ceaf02918a9db42c16d2c0772d7788a7
z33a61d03db89aaa3625cbeaf171472707cc1d07849741b3573d11e6a38de3785b3f66b0ea6097e
z6a6c7314d92a865bb3ec705043504a67b8fa8e172aef98d66103f6143fa705e3fc07d08feeb3a3
zdf3b80bf64eef922d46340406a53ce757ef7e66ebb42dac8ae06c76b8fd13e2663e3aad9e5d336
zad1656d77728f7f27870c7169b214323cfe4bbe5a6ec377532c347c268a569035d0d8d5c97825e
z9ff60d2c8604a806242abe79be1d78c6c63be5aa7edba71678c9ba50143d7c9af721d096444d32
z5f4097a8ad0cd5ac400f7ee9e9fca35230ffd329c42d518a7be8b534f442848678088135219a30
z9c4cb3c7a1441e982ad392a6924f1b906ccb76ca2d6fecf884a4f8593ca866b441969f5cb95387
z479eb769488357416cacb11425ea4b9cca38435eb0e177415e475a9fa85ca47dd249be56891eb9
zb33145bbf47854e0014e1dcfc87306257a50e8ca9d52e948fef3bf010a8467f7ae4f3fe407ef76
zc4f06ec830c2688c3f855adba6307cd1c89378ed252ade3fc2382844045151297e857e4927af1b
z03b28d30150ecb6179a05bf0f749a871c8cd1c5de58351cbfe8852e1c52560f8bd99c87904030c
z1c4464555f3a749696e865f0f5d6ac87ed7c2016f08afe57eab3912d6339ac2d322d8210d73d47
z7759f0829d87ef79f44ae786f515e09b3bff676280f17300a9434f20c334aa545826c889ea6077
z5a6c98c17306ce1766cfc6a9e882af770370bac68af7dbfc9a8137096176b91f0bf0cf0658a7de
z39a68bbef97de141b70addf9a33de5bab19a4c064bbf21e642b4e08f8064b52ac28c643a68ade5
zfb6bb1d2b9836bde7c1547955a50e0cccd51eafbfddcce9c0bed1954adc9baabf9042d23f29095
z63df389d332a17ef70d98bf2157521ebc3c7b9343b5ad88d9c1be4e56454cf4d84896e1f135e6f
zfb5e7c07eb2b0e114f7f663f571928a6e6768f10f942f37d78e55c4b825dee0981aef0e253c94d
z3d15958d4e6030c83c9a94e88c2744d5c9e331464603f173bae5693da7c55bf156df72e54e561f
zb5854250ed79bed179f9222eaa5e94722a53613491b1efc774f16e09c967fe7d91c84bca99ad75
z4044ba6ed5ce457155845c8f74febcf5a7a8c249de89703343afdd489ca24d4e956d08555424d3
ze7e5ec3400ad71545b764791dcec99b121c2c7b72ee8f7d4d045d53994ba55dd54b6638efa91a0
zbc91874cc25e7e9d5396a7fe798f28e57f61446e57d754d219c460a19bb0e5043e4d11a7d8ca60
za2aefc7d21ed4cfdb05974cfa80daae136ec4945de1b94ed852441d7da3d164fe4db62da1c0af7
z5c91039c513527044e18cdd41dfba70a4c7f71edd53a8aab0c1c3f96771a2219f91cbf0d3bb5dc
zf456671320af44d1bf2e9c5a373e4a55ee7d0fa8fa173c487efbe4535ce2ce94ce7f5f05a448bf
z3804a3b905f7bd8c36fbdac466e896d40618625701d5f126d6ef6739ef7e265fa2beeee9c29eef
z8443560d2605c6cbe9e17fd254ecee7d3f0ed0d163ba454cb829ea838e1dc39c20446a7afdd4b8
z1caa708f2dea36c8f2e7a5435ca9c0730b7cf7ad9e3a26f03abeca9410308b4a9429011c24286e
z94787bee13e2c4a6d3c5c9ab5b7e909f5676dc395ae23274f873dd107aa9dcdfc57cb54a3f16ff
zac968de31e16e56e8c5cfd6e1a8c5dd1327d0c0975b63e1dfce6d6aaae8287dd10975c4687f6b6
z0bbfcd3acb14393f0b7e8028619d032021342e5e8cabbc8dadecc8c22c5eb3ccd3ac1f2a3177b3
z514e0b0e1ef8e5f82ce033a2372ca8e069d9c9692f513c837e1fd6e974897f09e998eef47f0964
z3349659d35c2dc088d598be62a5c38c6534ab25f92959d1c75dea534b3a65039ea344d870375dc
z59cc6d46f98f5aee04f8cfd2381f979d58ea297062ca6b90a9f33a725a8c4ce12f4be6c2076c2e
z133639bec47e94af31948c45c962ed96ef029236b530bd301e4f70d58f18171b0e6ca54b1fa4ea
zb016db90ae29cc3f3c63d6eb745a2af01f570331bb96bd166a2d3783e419a51d27e74c0472efab
z4ea335399d6dadf724b2797f33ceb4387ab915ea6e671ce7247502cbd0e0f3d2007d788ea18c61
z4ee3b135aeb6fea8efa74c0d3ef1a32c81f2b6208bb6e17d674afd48eb0867106978f96fea503b
z1f1c8dc2125246d505a00704dc573c6d119922bc26e6420da9ecee9d9ccc2719dfee0fbe66ba72
z3b1eac547cd96a8af08552b142eeeac762c635dc1cf9d5c32c2f5962049de6651f139c4c28b3f5
zf8a8760e6380c9cfbee0eec2755eecf53880fadb27595ec5c6f28dfe5f6534b9cfa87eb2461594
z15eef59a37cf067e5507fd0c774197b39d05376b1f9a9385276ccfc7ba2cc74fcedeb1e7c9f06f
ze30c26c54cd58e1d01f22606cb6db2eaa11640c9e666e83023bed3cbf255caaa563d0fa1f0ba53
zd6155a316e06da3c8abe8e6171a4dde1d76929829c149f2b96ca9fd8f9c9e7955cbac498f490ea
zfb0a388996d02b6eee6832f961c3b7f7b2e6567237f818e90b2ff003620d6db8007497261924c9
ze05c0b788da5052acbd195a8444b94dc5d88286c187bd55c09e3d787c8763e13bafffded6aed55
za602a9ba9752c09b0f91179ffd1deb2832a98b186cb043ddf52bf85d08f347f95239b06b499d18
zfafc223e7ab7c4cc19091dceed6197329401a6a8d3f11b25ad6b7b221ae59206f3125605edbb11
z57649d74c03a3f1c979cfbe4bd9d3ec9c227d48a3c8c44e85f0bac149b3e0916ef9d2ab4a5ff9a
z8b89e8f23d55d5bacda998b19462e3732a46c101c3e38e3f3ac14e755397e34464bb815d3a4e48
zdd50999906c7acdb53d6f60828892e0ef061b7cfb31cd6174bc05e44aba31f4abff81bbe46795f
z300ef6732e9f093f9eb7eacb7687b52910afe122335df2873bb1f43eecbc651764c0f07fe5abae
z765dce5166ae69555fe4bd48c7f30e57d014ff6298ea5eb2973a1967cc097dbfa8886f19d25bcc
zfd89fb1503835d1099bf7d4bb54b0b077faa7afa0642fa425486150b3ce704858fee5d89e6e64e
z4c70a7076603873ae3103b6919f5e6fc6062fde537f7ece2fb95a9d7e7a7e88ab5fafbf4f045a1
z87d6a416380cb52b7ac416ae302895e3ee73a7a03642497e965ce78afefe1113ce07bd5c554dff
z449467c4270322575a42d596b719dc5a693cc1dd8e58afd8526ba7778bff569eeb22723dc30a8d
zd984ef43a508d71c32995b78dae063d59f453d487c86bec2ae00c573a1f2f23b14c668077a8dc1
zb52a40ae215c20cdc9f1733f422f36a376b363256e7cce47daf8f96253e13d5a66e9ca39f8a007
z54dabce105300ded097d2796d28a122413c1de2e2d6bdb8967f9cb57ca245a8f140b5400dc551e
zefc24103a5f2415a5b42bb975b24049183532618f8daadcbe6d0406047b6b00b9b2e869bace183
zdb8a26c974abd1519855fd4a5817f10169c5ffca04c922cad12c29b97a9899779a2cffe8354b45
z6be72b84fc90f6924a0fdd48afbb1bb919c283ee32219574bf0c830eb63aeaaae7197bde6695a4
za4644de585dc34fa90a2882bb873f9317b8ef18b317f779a4edcbf843b1cc74586fe43209a1685
ze7cdf8ac919dc04fbba1c21f304a3557053e7ed675ced2b261b55792fe214ded43301276c10c33
zf7068c883fd2d7caa1bfcb7bc2ffb536db782dbc26bd947779aed052400d6c27d34e0407a5c643
z80e76ea73c3f5873f9b4bd155dbebdc77d46697c50e075ce7f34a41752035243220e89e1af0fa0
zc4104e575097a069942c97b7b2adbcbc03c55716c5f070b9f49bd5a5e9f49e36bffddd78c21cdd
z2c1909e9f63c38e057644c4812d76ee8ca9eccc833691bdd7849ad3981177550a8bde91f8561ea
z53f9bbe10ee9788115db440ee2291fa71c1cb63b743cca16756f1aa12b3799d9989d918de18ca8
z805e92a9a9130a80c30092118610ca20fea68a7986df1d663bff9ae9f37631573d2d0e530bfb9b
za95b8cf47b842a402777395f7aae6a6d0e92c58d113d509cf5abc05a71224c49a34bbba8e89f8f
z54aa75c195f4814a7d26ca40161eba68182ab5f21dfd901bd19a862028d4e1c02bddb2e18d7076
zdbe2e2b144e4448cf128faca84b38e84284b293f68458eb741b9dcfacb12958e9c8e63dd189b94
ze9722e73a28a015f7ead4916dff4dc8a8ae3803d7f4a45749f9bf0008f755f0d5315b0b87bc48b
zdcf0c0b8dcac6a047b964f33509f146731714213fc2e827b0a602213ce05dccf84f0f1bd872574
z01e11b90e9083997d079d5c776754ecce947ce91d416e20dd749c1e11ad31646b18ca91b1a4bfd
za6c0d866a1e47c3ac99c828947029899f48f5269e8f17461549d5531c04cb952b96271a989199a
z47502143729ea5dfdd22bb2129eb0a2aaff4a6597aee99bbf56509fa1d75ecd23cf75f3c91da6c
zc8e7d7ebcf73523291253745adf5a5613b75ef53b7d1731461b40e7d660e60fd95de7fe27e221b
z88e0c45dade7137dd53b9d7386fa6593a9e52582b622404854e2e13bf713d58df5d838d388ba28
zaf2d2be3534f5f09596b1969332240990edd4b078dfdee7d495deeb3933aa90b05cfa8f2fe9932
z5efcf449609f5c339ff7803279127687c488116515e462830b3e40f37ed9eae90b999538374c70
z81f64a72e1d9094faf14c45d7daba33675102e41a8913b0b07dd16430a9dcba83e0f1efe8fab48
z21d6973fc1ad1abb11998a9b7a0149fe5af7e38a2d17dc1159a99b9fd09aeeea8e5811b8c2599a
z5c3d5239b52cdbdd77a2351a1527f4b03d353300e4e3195adf6deb6f97dc63c46dfa8482f134bf
z93b11044324e5f7a3bcb27367cfa7e57ef6f84e39adcdf2caae571156f14d33e69a668bcdb87a8
z6da6f3e6fcca1fcd755db469386f15051c89ea0b57da8007ea7529e9a3e862aa39e32c239643d1
zeac30a8a5f8b0602022a6a197ed8945cd126f0fa6b51b284c72585cf3dfd944c1ca50e4d75a17a
z4b6b6caa10dd17b620cfaae1cd1a338508a7dcf7f3167e1b55fcde4d29411d8e4b091fe433d37a
zacf6776ebfe03a2f5a4048d5ee4a24cbd2102a0b910151268b16f085c29ceed356946c0bb52141
z0631c67208613ee4b4355d00110d635e7de233624af38cdc019aa67db5b3407d68d17a1f74714a
z7d5339997ca1a6f42bb430bdbc2e587b28688b0de519b9386d43d7ad49ad0ceaaaab52632dc5aa
z3f9631b6e8cb43027fcd7fb83c428fc43c6fd6db2ed2001c5c64e1a0b8934089045326e1787b20
zcbbe17a6f8cc64192ee71964b8da3010fc3db26064c9791fc0044b7fce22fae0484bd382d1e2f7
zdbab64e87361e9be81e75680d4bbf13ae3e4c861b8869ce8d74660e43820bb60bdd50a029d2800
zc1738bfc906162270e4a30a36cd6ad02f924aef75cff4e637e4501d3b82760d73594ce6f247b07
z6b32ef7a0b7a9184d33932621dee91964d801e0539bf424230641727a2a93ce12cc7aba8fc3d94
za9e253b0560384a6233bdc8e975621035ae689fae56cf2c5761b544737f0b33e5eeeab2acf62b4
z36a4299992bbcc29eae08e6b1ca8997e5c77d1601ea4de67f4d5cc815160671c727061362a9f9d
z1989b880acf615ee2d1e85bcd071f584f885529e46f05ad304cbeb0190f8b3bc3093528db6bdf7
ze2a794c8de0670d47b5fb3b1ff11b0e5b0d53b88fe820b41e8e1298e6f42858d94fe6dad53a4be
zf845a0dd15e0dc5303658fb7c1bbecbb52c104f49d539a8fa547c34b2ed44091ea6348e43123fb
z3a7eda596abc7c9f8a45f9891b0e5a9d9e4dd1d90967d1f7431cca7f6e59d3c9dbfff22afd66d3
zbeed15b66083d660f45d8e3d30318f6338418266975e0b3f320c976fc55d606f9e4494e7f09e60
zd6489dca98f77b3b1d8a57b75454dadcf84bd5b0c6ea40de960471aa8b5e8af1fc557b39e33f6f
zab98f9418e69937c890022892049e510d034df7275c938c7de10383db2ea5cfc09383b12a7390c
z616f6c93a12007af0ed76a83ac2287f400aefc4717fc699357e44bede45631ccae9092fd4c0148
z4a32a23f101190e8f54eb6908463876d05298888ec24e2bb43c138dfce1ff3dc774d9b5fc50bca
z8f7ce57374efb022e4dc48cbd47cd288ab89d218241fcd8b84f273212dfb42f6d922a339c8d40a
ze019ac8332d3bfd6685aecad6f19ee0a2e8cfd6f4526b8572d9880517104e0fab8d5ed57012271
zd4c818a7ed371279db7ce0c7a6de5d0b43b8cf9ac814e7acca009d544b2bd4ab65dc357bbb0352
zd87da1c8b35366b0bf4f2db3a4b9e5036818fec758950666b0c3b67ffe7c513500dd1c20fe680f
za91c316d8a8c35e97633c6cb0bd87b53e00ab6fee96226f0f2d07473db6b1aeaec0bb54b5f749b
z82512129f2b72866f17e598144793cd67dd9f1fa5f7d9ddff3624720cbf3a9cd2b01fee44bf0ea
zd34b9eed594caea2b15b33ff0862b21f20e093435510cdefc96a0de1e4892e13ad517350e0a616
zfff6cdc6d3a77d050ee565d87716cee3d9186bf225a7e614ad03f61d7fca8214f51cfb52bfab4e
z1502672db3a4044093e251ec920598be4cf2e61aafcd2c24487d4c971c57c32c5511820b3ca69e
zbcbb3743dba9a4c91d6f3b7bea9ea0570e9ba6013ecb5388b8960d76574505b4130d3ea9123b56
z671d8477b1db475e3fab8affc4b8f2e8cef3da9a94adf798aab774dc13547a372ff14d461fb498
zc0cf417e35bb5b94c3b9008d1ff158295864a502f8055443cfa5686f8beca598a7177ab1ee8992
z2efd0dea92bdc35d8181d64611719515c53a2c49683476e3f4001fd1917aaae12193950574f959
z9778b00a710f1d75c4e649409a0dea8b9d2ac9f2b291d82c6533b646dd7441c86a63b453669763
zb6a73c9cd0d2936c9f4432054f84046ccf1a1eda75cb8b4239a0e75ed61e1fa4574f600e954930
z5c9bb7b29c448b1d381667e2d8422eba804b34101e5177552cb1058b63948a70f7e0e14baf009d
z7eb562679f42072b5e8dae10d07bbf086db417ac83ccab03e26f6344216f4c36e229cf4a26469b
zd75de6422aa5d1f0d079e75478368bf7b9a33e828905c9e582f7a490bba709a34c675855900b4b
z620bea2c3fa284f34024b7da47772ed0127f3a0957b392c276a140aca10e476c19ef1a4772ae2d
zf40322d068369824ee74542aa938cd31252e95b1a39f53b74bf6e684a36902676f779685910478
z972efce0d5dba373a96089baaa534e5e854e8c037c2e58f33122089c228dbb07ddd2ceda984afc
z4185f69fe69a96175afba8b381d53c4b9d850901961a18c330791b06193c4077cb3d43c32d2171
z78795a29f5e88d664c18b9d2320caed1a8d7d638a20eb316e6590ec6f61ba500a76646e25f342c
z4fbf82d51a73ac27e0c494fdd978bca5c74134068930ecec1374f14a767e735bc9c426fb167a6c
z7a824e6dafc7810e91656d071ca141e565841a8308b8581bfb418745248ca47cef2ea8238d2709
ze36273bf86a668f4cfc2a11f4a3f243461f8f7254373300a09afe0e1703ca7fc13e030909ff760
za20a1601eff45b2de191d35e8b9163df329d0b2d92c73cbf15965e5d6978acc709152c6d498ee0
z75708ad191a5d65408a5fa33425cad532b1fd4af9e62c40e4cbb4a5a59dc7097b01f3dbbf22cc6
z43c17dae457918064067cdadf8823dd3d69b411b122aac4b29161f460911ba4c4cfa1c14b11c74
ze2bfc1751bcc2ccfc72e3b685cc31a3d09d2b66866baf5d377ba2e66ac609d3d5486c09a3dc302
z1d3857ce9c172f26d8b5a358e029d30f5332c02c4da3927afd162b9928f1587e3ae84516894023
z264a5019d61e68c04f596b2986e7892c8dcee53b4d6616966a1690c94918c49c1320ff805e7b1f
z49a8f0b027f8c79a4117893a0796ac38ab04a583be3d0e7c258726907b2707b3c1084917c92ed4
z5da04c29a87f350917a11b7c21aeb9248e1e51c82598c7e27db224b468e060d0e47a780852e66c
z1e6c54fd6f26da84106507c18f7bfec53e1d8fba8019f121299c75cc0e16b382298d7f3e8a8af1
z7b36992c90c60be61fc6879b63695df5b1fbe83c171e6deff38db1dde0c69f10b41282330abc70
z1f1141998ca6f032f46baac4936f5fecd6f7e263b8e7fbfb651b8343a14f96809966fa2d48a504
z2eb621da851a004d24a56488c750809d7dc6c59105eb510ebd8eddfe44dc13c7b858a3a636b6c7
z7dc5fb872ee86ba7642908ced398e22c9cf8446cb3de3d5c396cff8d5be9dead3f2dd3cf9fad6b
z039f44d71f0f5bb4f3b74626d0cd8f77b2986359eed3e15cc822a1278a895cf2ef5cf64279a27d
zfd02024fdbb60754916a59ca5f3abeca624908ffad67ba6cf4cbc2332d52ab69b9b642b2d7aa84
z5e94d5314bb40d20284b74dd15810240b77c61a4c3cc5b8913b90df88caa24ddc1f1911dcc0962
zdc3a17b766229c48eb3156dc9cc530f63fbda3fd91152f08b24fa340ca549ac941b7e5ba18d08e
za0a1b16d02e53c7e081db2591b98c47b5ea4417e106bec213d8ef06663fbfa925730cadbbb570d
za9cdad4b9d7494020eb3e1f73af8cb31290b1f3f6c832846c68894a3ceb1c9702ebed8e44bedcb
z220c81399fe92c5cd30498ec6f5590d1405ade316e4a09aa6d457e1c011a0e045879ca984fe8f4
z1cddb992db51204502bb42987641cf6923f134fa28ce405aa6087175f5c3ceeef23d5134000090
z307bc8295b2a2e4bdc74242e14d294e6e0a10105038d03c9c768fe8a7f8026155b9c5900198e78
zc99f9f1f11f46e18c669037d84d0708045278a2c8692a75735df6c145c055f11b9650e5e6d3cf6
z1aa65890e9f697c353fc24794947e4497e4a574f8ac54ad61fc0129628d5592ba85cc73fcce0bf
zfb685ca1919bc963589580a89e278a3371fa29e93b5e758269637b7b10cdc66000390144b53bb9
z4a9db0ea3347d49242ccd557e885eba0824cf27500573fa2a3839615bf12cd18f1803eb367fed9
z0999dc0efd74e9458a48317ddf96cb1c74374fa4d66a1fdee4b4e7059c37d29fe615982b1055f9
z0cb503d0c47d0b50f0c852c9b88867dd36cf8e9c646ee177a874f0f7f19b15472225bd0d88597e
zfa0f724328a83cd612498e5231d7f33b1be7948b4a854f9b1233cd8b1bbab6e6bbb3c9031d6669
z48ea91daa32d659a50ef2f71af44cb4b90f6ba8b619fb75779c7bca6bbc76e9f27577fd0b8f68e
z2cce5bc1276548ce4031a7302d6d2343f5cbf4ab1ee41a9de922d76a12d1d850c5f57ba720365e
z63149c6f0e9ffe313a34bbf1cddcb28e808f5ac1d2a863bff01602fe12262355b9c6342b907baf
z4d010b89c09a85fa4537ca015e4060f0ec46458d6def361d7d4c33c3c31fe60166b38f72443d5b
z7ff80e546b7663d2ed39ecac327b202dfe85226f28657b901746526148e4fdc58244d6b2df60e2
z07b4cb19e2c1a1171fa515ae22c5a9f8ba60c1b7e33b0771b3b7b258e390040cf8ff8f2e4d7b83
z600ab5dd02f432dc40500343a33f2a8c4f6f6d48c709c8feb24bfb8e3482713e01847282a1ae3d
z3e5bfd1540de0337f0a031095ca79b9b8cb353b5c2405577fe813eca303f9f2ebf3217f5665456
z04d2766da7d27d7a0fff86ae056be1ac6b5e869c24157d1b51205de6918dba2bedb0bf7d1266a1
z5ea9104595a8378531125a799bed003a44f33be755784ef7134d27f776a177f702624dd5503c78
z42bf6d427a48fbbd710fe6df39b0204939c4a1a6f32359f6778f9fb1f6202a44b2355f147cac76
z5ddc1383ed2bb657feb9c6ed42565208c5ab759fd60bd065882a29946262800f2d3b58afa3163d
zc8c4a14289080bba4b73793ad2ae0aae5d97339c9350c66ee498e88b22ef89e640bdd47ea8f330
z5e740c9222cd1a98055cd23e3fb30d2aaf016acd2e8a33dfe6c7c9b8ed17b397926516fb5b57b0
z00c063ed9ccf1a1e6fa9ffb7cc6b355bd3c8eb5b0aac2562822fb6ef29fdd971ef75e9c3d23112
zfc395fd09c71672f47d6855a8d8a0b2e76f865794e3a1e517b0c83031e5d15f2ac2d54c08bd01e
zb3baeb660956bb22a0bfad066d831f4100d97c70fb7b587ba8a4e0c5df611a5ec78d1e0034edca
ze70d8516a38ed6f9cac5b206e877daf6c040b9ea84cdad07e981b43bca3ac1e65e7b4aeb1628a3
z59df3c936848ee29ca4a9e1095c3584da1ab8389085a695d44c8ddd8ef0e2b8342f507b8585bab
zf3db98427ddd27e779b47d13a9a8d9dd04347cb2cfe4b4fd730c3c88eb9ca3e709b7f5e6d9b396
zcb64deb2e9a1500abb3cbd26f2380a0eeca52e147688d9e9d4e788a609c297a6ac83c0fa4d70ee
z4930d8121a617acbf34ba3aa05d2def00c5629442bf41b5b8aee5d630c90249f7490048b8911dd
z423a4f1a2ebb481918dab7ab4a801e398b70379cf7f99519b37c78b3f6fe2c3103c7cb5664698b
zf90bd374059b5155b0837625df28a0c9f73cca83a69e444859e1dbd09bbdd876cd978b69aa02a2
z100323b48c4abc46954ce15647e4747bc56d7c6a96b98d6f092f56e631f93c15fab1efaa7529f5
za2b3a879439445746db7de68f56e2d6c58312e56fca2fa1cb35daa05f780133a105ea3ef3125a9
z86e0f51a1472ef855aa6d50e4eff6b9dcc93deaf2df47f0337b450c40a7fa2d45a7b80cfd83a79
z5bf9a9d9ff4109cbbeb435259950b5a55983fcc6a843994fe1d0db4e38c9fbbabfad05b624ae59
zbdb64f504a2c20b9a4dc79e37dcea2ff804c2eca5879f40bc4d843f51dea8107c7188f80fd2ead
zc58ecddc9b3bb2e1366ce41cf323f25aa44f39c5d07372b0e6d22b88af9a01535a985c14b2c1f5
ze55e4a75a2cbb00ac74bd9a6089ee6c5b5817305d8532e97c77fefae9ce5d1299ec7b5c2f21306
zc338a77e97f33ba704f59c02a7fbb1358ae2d5dba00a060ce8c173660941aa26d095e7692c4e39
z9fcfcb7a4433d595574db1e4ac89529ebb7a9aa95e8371d0912dacc847badec9715a1cde9ae9f9
z4a4d25b1d5393096cdaea239d965e9ecf57abd2d14a8420a22d5b58110ee6de6b106115728fddb
zd2e3905b1d324ebcc60560c0fb2e521e1ffe6e7935f9c8ed51bb2d2f926fd68434f6a9804e07ed
z161761cd22b03c9b9d30a325734b9deb43965db7c072eb6e2ccf504bce24fbd97cc2261ca8970a
z51e542725ea619cca84647ad86529db4b9dd4721c5e23aea294cdbc7faa24b59f94d75835d5ce4
zfbf9cf7747b0d17adb9bef580ce966401adafe47d147d8afcdb78b67de79c7a3358fa409321cd6
zaae5e227935475eeca967895826ae120566b1e63d08639b0558ef44647f54ff2214b3c9e825230
z524e62f1dfb2b8e0f8c43c62f5867811894de7a837eaa990b382451601fcd19c5db18afffa1f31
z87d43e31225628c64d43fc5a51317e4b9c2f535b7a038ac8a78f3b6e198d0bcb5630695482cd2f
z9995ac6bb23cc2cb265cbb0e190e40d079799df80b2a600bb89637377d148cd17e8932a4308c74
zb6e2aed73a53bf111a986266fee80d3da8cda67a6db13e2c6c9ccfe368bb3df6d89bcab77cdc1f
zd56adbecb2648e190b7f633b17609a49c56d2aa0a21c988f663e797ec2afd96d29130d87b45fbe
zdb5e17fcac1b41eca3ebd30063bc794d2c736a4d2f0e995c970953a5482b9634824f591932b217
za4ade828fa52213756b0824656b3d26a5b454585116f990cbe02e6ad265254357066b9d3638312
zb170ef766c0b726fbd84c93618268340629a32f7fafaa64cfd18db81bbdb1bd802ce235ec536f4
z645eae7d380a234e38bde18590cde606bce7371f8e2432d09a92f13888faa8bf027efd03f269ce
z2d64f19d6e629a7ce4c641ecea33239270ef1174c2e98b93a94731a5e48016c7651e30e4972475
za40f4451f41124bf888acf9ed6b1cc0faa451c11f7569f6a4edb0c70377125634caa4b9743fe0d
zf7d96a464defa3988fef9986fa623b6002f775230a8ca611816fdc57f72771eeb7a304d4a7f858
zfa362fa1781d0559f7c583640c260d9b986a24daeb68505436ef5b36e1b33e546a80aa326fb5c0
z2c1b8ce396f501f7501365e2d15185559971347df843f5b760e8084f995a3e07dd067c37657684
z32c077e2d7545b3ebaa009dc79175d3302c4e31133b266e2f5c7f1e735fcb0cb1cd49fb62ac791
z2b05ec0e896c3ed379e996a7d6a21d17bb2c8763a93b518d63631d51a71a76a4ee96f004dcfe14
zd57a1b8376b6a104e07f1fe38db8789a72dd53553bb6da3a295cfc576fe8e60097aeee19be0932
z8a672de987f7f52b9bc55928ab40046921baeebdc4f965ff4b03eab5167711568b404cbadbbffd
z1e80afc6a17f81d5cb03325d9e829bc3475ecfd81b6d8f548855881a28dc0f60dea5f31863d60f
zac72d07c5efc73dab2ce2befa19589c6b4ccf8c2848061b96519faa5ebc2cc6a865d0291563ded
z1d71de6938e70f8bd51b18d79abc9cd179c2692d9f88bcd4e09ea852970fc8997434d053aaefa9
zcc4605a4c2c1199cc0b76bb20c5f337bceac00493e22121516a7d5f770f30219b4523fbf24e43f
zad55b1e5b4198e98a9bf5f21a24fcb2e2c6c75f713965579890483bdea3724fee5676005a5e1a5
z95d50bf673cb21b80b5fec4ac035a5b8aa2164074f25d1daec5aedecd879be1fa78eb17386cb6e
zb935583d5e9060626be58429f55b42b6a21bea4b25aed3609ca30d04e19e774d0a5d9a70823db8
z63826c0c5a91a77858d7b377a889d61a2f35986550aaf7b55a2f55d4c3e5e57f16d21009770436
zce14be72affb85fa095fa5adf9d2afeb21a0f813b6f74493515b664593a1590da8c4f3d7dc687b
zcc179b06a4924e4259e7b3fc046b3323614ece95293319ee61d68031db596307d61a7eef6f2244
zc5b359310453062b73d3f5cebce6febcf82dfd4e507269b476ede4d88bc292dd21a542ce6f85a4
z50bbb229a8622a0d104e6713f672b764a84577823dd9a8a201d16caf4f8a0904b536a0303550f8
z36be51a712627afbaa5f84a631125cf246e77ebc32cb21044003f5259ebff5c7a51a3714260417
z0680c23899887ff539ea96cf5cfd6c015f9fd724ade7dbc8d1b4d7c6ae69f63de5cd15866e9790
z1d268f37789edaba15655ca3669611167e6ef8e34d561581e508f491224e729e2ee1c4ed349150
z0ef24185e80d6046ce9b48e51bc7d723dba3946917db670b4d0fed45f52371586e93f7f555ed8d
zc852ffe3c0255aadf64900c9c3ab2b952fd734a06bc8dd3cdd45dcba83ba1d8c83f70b0c52667c
z8e9f018027aa004a23a2968ce457953cb9b81a6a58a4f2dd0f05deef03753ae0669c71dba87ccb
zb116894a543e22426d1fbf5b085369103b5760f40266a985e30c387ad6929776ee6f1cd13ff0f0
z7d0f79dcd5a3be7ac8ccb95e11e73d0bf9f3fa064e360ef290f0517b44cfff8b4ed36765770d02
z591babf8a5e5ebabd044bfe53ab88d108f4da87390133f2288aba0a375079b6ce7e1dd17ad8ee8
z4f705690762d274f2dbc514f19d638f079f2b35432c1906fdbd2a547aab52864d80e67d2dff813
z047af28a19518f1c70415ffbdf282dda5f3a839ba7a43b87afe69d0c0ba4dfa31a0eb6d557fa0a
z4223e2c11d5236f06cc3d876ce0de739e66230a2d2fe4d617905a7dc3c7aa12143157b8522bcbc
zeb5a07db47d44b91586fb9db4cc8d49b7d87a06b0b8546e1dfa65cf0cbe262e38b48d86b430944
zf51ad1f5a30eb99f9c27139d07d2ad90b4d45e25d95fc63219c0e01cbe0782f7beb7efb7b780ba
z692b2b4f94609ff2c5e2ca98da4a248102e133e01cacab96d99fd6c18ca72ccc705c5fe8b9b350
z7aa65ee2a7a35f2371056690413c80e7311ec5c9afdc2a97721a25f7bace7ea48d718bffea2f8b
z0978e205b3d7f4e75f59724cdf58a1c4a8825e3dbe43e65086235f08278bd367e55eef70254493
z4037fb8d3c527e0bf75e2ffa895f28e39274088c50b07fd1da71df9a4967f48be728d8cb91fce5
z078dbc86011d81136fdec93429fc0b852091f29dd71586913377f63047ca322c6f3371c48387ab
z3be90be3cf6ec47d07915af732629a248af97f71ea3d43583f13786601c89447e7d5da1099f7d0
z608329d76b4c63e9315e981384069692c03e8d726abe2a06c20062a605c7a4d29da440c17cfe2a
zdc308c09265bdf6cf4ea387b5324d697b09a2b4df89e473fe8601155c8260cf0f97bb2a497f91d
zdc059a6147eade2ec3affce0f2f4a1a2f8cc3173e9fe9f439bae075662b36f810dbc5b509fc500
zd3917a3dd9171f29929fe3bd7a5e51f1ce6f1f604d2a557e1fd08c96e59dbce1139ddeb4b9161f
z99404c187dbf454e59575b96b619543b53c4981cce775a713177d14ed114e62d3f8fa83f3c7618
z8325d2bf5a6fe1e817b913fd4592dc57029de5f853ae3dc41492f2cac45cd787e84849cce4dc61
z78c79894a05578cd176eec9e9ded27972f472bed3e580e96893545fcd30230616e4ec6f964cdbc
zd7a4bad55d8afd92a6ca81753c1273fec26f07ae3580898852b0687e6929731e5babab705f59ca
z0c78026d1eef3e38d6c035bb21ae5d3630c5112d114a4ec990073820afb3af6770af995fca2d23
zb11f2134d056f4f8ac7b81de9e0a48a7c632f8dcd615ba4232ae66f8644bc383e8062248cf21b8
z6b42d9a0da5e8e74582916326b926cb9d75d505d4b9034636663e29987c2f091224ddb79fea054
z306f6b9f7fd53a33a0ae2aecac5904bd71b7568fef2c1726545cbb792eb92573a8a46f0dadc695
z974366324e8ae3e09b9372b0a95ced370fa7cc091b0834fbebe6a0dcc43aa85c8518c7d5671bfa
zb47c6dc37077b15c6d0ea6cebeaf12eb826fb3ad6360ea5de685375840a0b3518aaa674a4d9469
z46387bf63ac76313e7e70136b4d27274e2cddde32028fff069047bfd91be984427a05b993eacfa
zdc259dc9db340e8cc8ce2e49205c33f7d0f9391106f3f87688f4bc66ed4f9259a40740d5b8b9ac
z899c9e415cd328bc665cbca7b386381902a4c07489e64a80244a61a4503764d686a8c002fa6671
zd02346c31460bab0bfd97f11b3ac7aad0f7edae4f5b8cf97f1f50203dff22a6bd3ca0b4a785867
ze86ab8879e27ea6bb8777e0d4b0c9b9841d7188f28b02b2481bf9241d23e2ee1aa5bc8af583c2b
z0555e2ec247c146bf12c0cbf0fc494d5764dc7ff27f3e4c95c6e4a18156b157a04f16318a25581
zdc99067019efaf5e5681fb98d2c7a395e9e0009283910f9cc2054a5e704d300e82617083c7d245
zb4be896d4267fe68b019924cccadc89ca80bc41839869ba89c49ef2451e56b918dafde708f960c
z3e6820219a638e4f2acc523a784f351d7fd8bd714fce0a5448a30297105c19122d2717faa64be5
zdfd04d058a22be8ecc175c69acbbe479fe1efda8aefa6dcfce79772d04ad428220bdfbf0a8f542
z3249333dd7c681216a88722fafd57cd05989ad7c1155fb0dfc3d548f9f7b8eaff23b41b526e0dd
z2361b3b39b3e5064c9922b5c929e313bbde92a53af1cd1dc4926112bf5a4b57bb592e5ac16b322
z74463f05bdf71985eaed047fa97700ccc387b761b600ae4fc74b104de1362106587f60e49bbecf
z2118e6e480f9b1c522f7f02d2096a128e31b48d8f740d902b1ccf62f6acebd428a0c187b9c57e4
z249f903ad719cb3bca0f8f582025e53501ab88563930147dafc92eef9144464b9146f7ce577a87
z7bfe6578650f361885cc1fac074487ec1d5d3f5ad854582bf963eb859b69a3318dc3bdc25cf5cb
zc0d2f025b6988463dafb6e5ab6d04e809da85630d200c4120cdd99e839855ed613540716957904
zc986efe1eea100afc4b4cdeb829c71c6f260f1260fb36d64b36542ba9a7877362420991ed95400
z51ee79ef5f802f26b1bb3a55880c82ee081d989503e3b3d63d1991aa0b180edbdd4526d84998d6
z283fb3e3a521dac10492f90d06206e8b2070fdd4708a2bc5e31f16782a7c651d3b3f54b1ab2351
z942a0d819cc58f7dd364c3adbbe370a648069c806150951bc415bb79eace64d758179f7322826e
z51732d0b3d4ad25ba62922d4e3a5f0ff11ba378b229547c814456199cd9e2cfd5ffdba80be8da2
ze8f5782d4d4c9b593e8156f07fb969a73d7cee383f9beaf5a17f223ccec89995f2a7f2f1d3c720
z36938a06125aa0db9283aad95ed6f0213ef66c25398b0ad8bb920e09b413d8d20e3315132f7df7
ze3af9cf0f13c993fd3fffb8421cb0afe8e3eaf110bfe181bb14ae245cb7e3e082f4caf6f23b5f1
z1d64e17cfa9939ac4a892a84752f3f295deef83df70c445fe769537040104025162e998eb12585
zfd733fced1afe1a0fb4949f322dd4d9b107b5171b586ffa760e358eac1b782be440a9c142b212c
z9e554a94ab1a844dfaf0fafb207b1ea96b699585d804b923a1e1380418f964c6b1dfd6c196237d
z62f6721db0201e366182db091d627cb96e80311f66ebdfe28d1cb0487753bbf4e0840fb58ae964
za1ec8709fbb6d5e8fb9b92d66f8063870c6b94bd42b00144f348cfff39eec89b8f1b25ec777474
z05aead5b1967bf0624059319e4eb1a7d1fab64e74c3ed835e23b02d55fa0a1509316456ac51595
z44a3a216d77d2eee8a32ec20b6cb782d0774ad8e78181e985adf049d7b2836aa8eeab63e0e71ce
z4fa895a38bfe838733494e48ce079f77fe9e38f60edef50ad808c081eed13ffb606a555ad577ad
z43f32dd48f779070c5e59e82131d5b4395009cedf55872f5c71771c19f17274d66c436b97bb5b4
z3dbc76cd6ffbe8813996bf21c290e9e317176d74a8f2adabf493556a5932442a09762d49758af7
zc614db411ea595e8231935dc80c7c53d8cb89cc15bbaf6125a7a806782077cf9c7858a5a0b2789
z758dac21e3dec75146be7c5fd06b73fd167d8596bc185b6d3aed48605390680109437eaabcea41
z58d4767eec63b851bb6408ec5181fc4b7017522b15de4b53f6e30390df203c734c4ea1791d730c
z422bcb5538013ef9a745f2d8cba08bcc8b35163b7620d33c3c038fde1fd4fefb0ebbca5f55b9df
z146acc7c7c06efa6c5b37fa61e56cef9d0726be9cb5b532711f253b734e71ed4c078036c4a8ab3
z50409285a13b1c58836b9a362f2eb5055714bfe70577fd2a827addd0bc35e789ba5e9e11c7e87a
z53a0c8b5c9009e31fe18204239f466c8f4aecf4c7d3aa4e9f51dff1c960c1a040c8f38e286443a
z91f90afa69eeb09b80915e1dbfcdb99847ef76fc591637f62ddd0d7edcfc01f1e55367223ae22a
z857e3990f66434c30e13591f63c419bd97ae80b2ca8aeaee8a31da4e4a5e5ecbcb69dc7c53d5eb
zbfc47630a8cd2666288282280730c20b49dd88055547aa2875bab89fa8a07fefc8d3a10ec7ec89
z333a31d7ac5f51fe0545f8a23742a140b9dc312744d30551a0416ab5b680a37b462fb779c46551
zeb45ba8f7f4b442828167fdbbabbcc679eb5b91166da57375cddd6510acf9467e204174bb6227c
zec285eda35be30c18a972ed6533cf2a2d93273809e404ba578d3ee3b0d4910ccb6b8f2c5640bc7
z13349f124ea9b780ab4bc62b0d12c8f5d5132c4ea3b3ff4e68bcda792936de7cb2f0e5c40e2430
z3e4ca09dd73457246da13d443f3776ce97110992f95af9aa9b5585cacc87423d8961f4ab73b5b3
zc76d17b233314b6e7dd56b573b6ccec1237b3a1fd83a1cd1a4dbd119fb0a07166d18f81e8b0045
zba7f9e8a71febba093cc1a15589a1cd1d0874b3a8ec718bfe290d884c478b1498d40b70b501a73
z3e67443a210b31c3b4221702b2678acbb48be16fdbc44957785b4e29832742222c387cffdf5397
z3b18ac91c9ddafc471a88c3975d996f59fac6687b1458807f535fc772aa465082cdd6384b04541
ze53be7f02aa99fb0a7059e460941f8d92139a36750a0f5d0e39e267dc84c58fc7090d8073cba45
z7e0dd7d184569400b44d755a4e5979ab8090cb4d07f67d03a8711d91dc47fa4ba12761ef750ba9
zf8fd189f17a4cba2d349de19b6cdccf413735b243c4e537986f1a589f227fc3bddc422a0c60711
zeb30a57e380178cf66d62d134de546ecf5f3977fa8cfad2d0e05b05a19a2df1f6b97862d6af13b
zcb404cc5671c9e5201eef2428599e02737515bc35f340f82bab11a8ea7d6ce19575e913a0a1a64
zbf484b386b789bf84873914254cb368b4d12aebe561041a37f20a292f74ad8528c02b2b03196a8
z3c1bc3dc8df0348f8814b64da55fc5e64d860325e3a26d6890a14dd78fd85c11102751e9bed63e
z87ef09054195eb0ed78cfe9814edfad558b2d569b2ce26b34b5af2b407c75ceb3b2eb5cfef2d30
za454846b85ad160858d3f40b6d405a52b290a5718db065c6a03cd47dbd39e6fd17261b90d8790b
z044ea83908b398392f3b6809686b498fdfc40ebd475d258423c00d3e84dbb2c065adfff35bc834
za2ee67f118feac6a5b636cfe0c75c25e91766f46423c01613a171ff3ba0f051a7eb3c9acf3dce9
z2dfeac88709c0ebf9ec3d2cda6cc14d325b52177edc7accc7aca25ab0728c49386adc53292f0fc
zda232a3c75978f7f921086e0ea3e6de21dc799da07e36e9dddde2e4094f362df7d79d0d88138bb
z060c2236598e3f3088949d1cd4f303c642028c27f73aed64d0990b82143e7e079540a5a99e90bd
z60158a28104aae727c3ef6e04024ce1b055ffafeb3bf9fdfb957ed60599064480f1e779982de46
z2d769681305522eaa69f21378dcae6df24d920a34b190f0564a01663640369ac94ae9f488fba41
zd0f372b3a5ba6e6d060a9efd5666cf87c3b3d8522fda776220f94b1f4304f33377bb29156132db
z44a7c227a5d6ced8f10966107ad48a33d5cbf044b284d665f70235bd517a9e2e0c903306075e7a
zb01b2c4252a87739e994700b4a4c9b6fc7911e2a6878b8af37e840b82d5296094d4dd680b43963
zcb12cf6984655b598cea1d31d36854e4e8da85ee7fe2f94f6e0531b9bde9e61f74b149e1c46978
zbef05ee8c7c40595cf639c29a2019063072747ab8adc1f277089465ac30885208115d0582c4384
zc71ade9257ca17956bb569272c7925688a9bb84d2d4aa5c4598845e5ed12b9d70e0f383e1c2c40
zfd80d654086046a501d8039c2f20962755b21a85e5017fe087a1566631b815622d21d8e4436fd7
z3d0a95828e1a729226027a054a412d8a740c16664909d68c4071bf7f9ff242870ada8a079ee9ec
za7415e8e872d24331d865bc1222c84844f7ffd7e4a2df29fa55e8d99fa305d587b4950facfd904
za7fc562315030e40b0c79d7bc7ddf2d98a4b16d27d1665aa0f29ae9b006cdf342c8fe6e39a8b18
zc115836081a6807954581a61fd15836e22be7bef501a45a814e8f868215c91c3b446f0144ecaf5
z9b0cc7bad586c3e227d9c2d2012eff033637885dc262205a1da4d69216482ea3ffb9261fd2cfaf
za6f54e4dc0aee26155bf487ba52e0a8d7cedeb73a670ab5196a89027180d1a71ef34fd241ab589
z5a3ad58759335d6ca2b9781cec7994d4c0bd77aa71fe489346f54f9863a8f40915a06955bc1229
zec1e2a18f31a43f125b8f36e9b812102eabfe0efaad11a2c47e07bd2106b93319384d9f01f04bd
zcc21f1d747c0ad5ec48f7f85776cfe6cd9b4aa6f611d752e4f2f85e8e7591d9f16c9e431c3c0b6
zbebb248cd778e78c5d5608269135b3fc753f0ddb3a6a3503f48a05c22b61824b31d1a5847d12d6
z1308d7fdb02b3e02e42b3bbea546a70075a076f96854e2c756fc4826d4abbd8ed0f7978e6193e5
zefb5ef4cb0993ea25785c8eda07a500e419ce61d0afa7863e98203b3f45d585b6042ecaaa26288
zd00541d6d18997cc20a5995251576695eed4c8df2ba54dca4c0c3a8feb4cc6ab44b220a5ad85af
zaf88043f67d70d46ca2415fb357a17b4bbd34b14193fda3e6dfdd38a0ad0aa60117f9b35ad108e
z41b5b2402808450d5bcd488e2a2b6a8353534ff0e42ba37f5371467e72ad28ac00db648229af91
z1cf741e97156dd6efb69de4ac8c44be3a3367217f5c89c7064abdb8ad16ddf3e73dde9d4d1f79c
za152fe496f92a2cef55a9b1e46502aebe79e8fedb99791ca2f8097425e4e1c4cf717af8278073c
z22909fecd796fac716b0257b049b64427b41abf6de4aee8faf21147b647e0b1224ee920040b5f9
z1194ff7331d7825604768922638f95cc935541b5f73e060b461b2d54a01a0be1325849693805e0
ze644cda997fb47be0b01b2b8e265317651c5b7c69d827537f0f4af52230e5a7ce44d6ac6084376
zf34922fe4f155b1c25772a53a4490d1ff5859da5b4768050d5599a045513185ba2350192474bbf
z68c6050d632251de3cd57877b1feae27c2141138404146b4256252d55c14148359873523317a18
z807ac4ca13d0e36b4c4b6d702159beab927661ce6b5877323b90089caa7152d3a39bee26c01320
za356de1b1803852ac952cb82f0e90a9daf6819a68b8d96fedbe3f7f286ec3a79fa7d04c5e171e9
z6e0956490ef73c597779fbbd2a2069f5b3c97ec1ee354496e97b2149ac2bb3b1d49b208d78bdfd
zed40bc25fcf5ae84822ca2ba6558825faaeb5cd34c13870c5601ce0f2a783c6bdc97054c039b85
z31e96913c4ee631d66ff82b4e6adca7e6584ccec97fd8735af3f85184d714bc80cbfc555095ca1
z63871a253bc65c7e0b960747d8eef4fd2ef4c89164912e83d65fefb3062d5032612987acd1f80d
z564b6275a834646990ca21a21d6b92031c400dfc5317d2cf8188a884c5030926ee1ca2844e9150
z6ed2f50b87c37a3b9aa7890f9f6b46d233e6b758b285582c0d27c7b48ce803be9724148f99913e
z5757e680813734678b91609d0048d0215f2ced9cf81caea6706fdcd086521fc521bf59cd8c90cf
zd1f7874fefb74e09b60d6965c7905dd2900699a08dee4b542dd88538c3bd45b0f95e69cd03f48a
z0b13ade6efb9787b014a22e8e9892ff4797037852577a9d795a77d8b6be7108d2b0d96241f13d6
ze74b1aadbed9530783b5325af1dd9678c4e7fc0a0bdcd77b645b58c7b7ee7c64262ae502363a68
ze074643972d9ed32fbf44e03d0dbd677721f4efebd921d107d161ea00e271ea26b087ca785041c
zf7a732489920385863389ceea83444de0f870f64bcd33ac664971e5280605a9216049102aa6c8f
z26e275b9487bf86e2b9fe63f6ab15c730a0b02307a48b5244b2da90456fa6a23f303f37ef43e0d
z771f3293f999fae5f9dd33875550868499a3c0fd5d43010e95a4e343895b758eaf467c4ef29542
z12b4a770331dcf29a78a5cc4208d44d96b1fdc72d4990a34ed8ed615f37ea97500547c9e75bdb8
z95b68d489712112e70de20fe7d1beae906d24505c3a0d638313c87be8a0579c95494800a54c4d5
z062644bf55329fcedaf4aa88471f237314daaeb6ad147be5386158431bbec21a5473cb588fb49c
zddb3e2b0daaee77ddaa83fffd96944778ce56fc7131c505b3962ae2d9dcf254ed60b62222fb073
z3be279da71be0082b5215d6040a706ab8b2cf25d5c2a632ce56dfe5edcf284ebb695e410713dc4
zf6b15af023b4a9450e0fda52cbb6e66c1a10774195e8ce7a575ed5c67e1356ace7dfeb80d35c4c
zba10c4be592a9cdc87b552b84f67866ea40782e13c1875167af4279d40c7dd9b6a699210c60834
z012e2244eb43e6229fef03fde18924a62a8d24e842a057bc30c7859a2ee9fb943664a9ec6a18ce
za70835bded61b291396c3a1b0d5b7bb51e2b34a3eddd8d9c87a30cab401863dff11f1c2c3ff269
z9077162d92284ab6e86fad564783ad810679355347d8cc617bf4db08fe50e9ae95722083228bfb
z58848ad720c3734d07a616d6ba6cb6cd4012f9cdfad6b5c133b9b61dafe926b482be6ff0a569c1
z1a42e7c09552bca809f3eeeffb8af91ed7c534ba1e714b22e06ffdcb7f5680ae9b1ef161caf8a3
z4c214741c265a6d5370147d28061b4ee640479a25cd3cbbb08d6efde0d9b53b4d5a7281e01088d
za1a0e0bbb4a376f54e94ddc697aca203eda41d64d9919f8d90601d4a28ea000cca324c789fa0c7
zd4ca6a03838e2e7036876e04a9979f0c225a9b6eb903c475b89440b4adeceb45923fe014fc28ba
z7ac81babeda063a0f9e2464ce5bc691be60534597a382d8e1af4a727a22d57973c961b26ed0f1e
z16092951ea62aa43bd08b75d7e37db463d23ab5dfeae7b15b18bf6609f896c57c29a4d493440b7
z63cca1e77d425b986282e2cd4160081fb5d08dfb60cab3a065a49ace9c860fe39353b7aa4e194c
z07507dd354efa31c676bd2057c89dcf46cc42955d607fb8dc32f76ba3c9e5c123561ac70798d95
zdbecce1deb07ee8656ff9e6db610ffc3dc13fa50c54f19a5b5be81e38ed4ad7ca40df81ae97dfa
z36d81113e6b7bae6f45207069002138e879ab2bccd0d1b2c72210430decb581934830256113289
z36c9753512735a4abb733f732b6e883db7a4861ebf19f64240585caef898f4cc2491c0f149002f
z1e6af83a546440ec86e97244baf449446d5fa46b716f3ef289dd07c5a7798616388cd4edcf5be4
z655d3344b52c6ffc0ae24dce78c0d048e5cf07bed46a52203a33d7f3123211bfba3cb6dee444d9
z8b0a6bcacd3205133179c011081ff4f9a7e451eae766aedb2de659327ef89b0f6c31ff12fd60e1
zb8c705c760ce701dce2a436008e6d1be3635f393e3edc94c6a490ae68bb0150b81d7e9f62c221b
zba77e97ea52cf65deffd71f81338bc5e155921b4fec2da63ca2c32711e332b7389d6e8a6aecc9e
zf3e812d89078ad97b4f5c8ecc1410e4b8906ae815061a7e832a5cbc4ea910d12a02bfb8c1dab33
z7209dfb532fad4ec589759861b14fdbff4105256ec3de2d98ec0dd3f3bb8ada938a5eb10a14a43
ze00f10f57a3e733949d987304fbede0f4be16c6b9698ab0d3d436befe0c39bdf2f06cae3e5a265
z875da561f831157ed8a52a64907a2269f247b481740afdd65bd416c124088ac117346eb8331f29
zcb675ed56213cabadca38d3a15cf260aab24b15afa9b6c37b03f6085f0020db9d722a869c623b9
zd51e4d1462ae5fee01662061f5b41d23972d2770783f041f26b757bec3db44686a961f30e8ae3b
z013b266b103ad2d12cac40d8166cba6823db08f34468e2aa162c469599f9c444b495dc0e276f25
zc85438e95cc169a6738f4423acea2d990af676dcedc6cb2d660967f45d08795498a1bc9f2a6043
z31ee8771031c179b2bf6d4641da49b78ea6007642d18ff77f8493800cd1a7e7990a94f944b13b5
zc4a8a0450e74193d93afc03e44a56fedcd0d3aa49cb4cf98018da8542511cdb92ce9af08c0e2e3
z6090b26c001a9d00a09eb55bc16b0ffc7dbb2accdd6eed4a7ca762a3aa83f45f5aea8e35fb73b2
z7be3cf53194d1b6a2e3889a6962044e2eab5cde89c16ed50cd342b86c83a52d8d06413b7ad6b63
zb025ab08c7aceb1861a49746f5300842f5e9b2690348f923a94604bb24dac9f3efb768a74e310a
z8dc5fbad67ef957aeb2f3464e0b20ff3f420828832817c4b17bcf8ffd8d1107fb92debb364f139
z54152af83d030289c295eb2cf59322d3270a7c54436267c5ca25b497f7d5087121c04bee5f164a
z6328fbab24eb2da85cb39b5d3cbf2a3f25ca6cd0179392e91ac3265e5394a96c33955c66ee0226
z4b3e376a156dbe1c5ba40329a2c38747f143278d7a8f757f7bf78e78e834e9041e5fb4ee951813
zd7beb49025ad8b6f4260460e41bd53a45eacc16280d13225f28557ea509e47193294acd423611a
z6d090e6e3b055d0ffd36f70c978200f154d9053d649b9f5f335a546ab2dace5c22e29ebef171f5
z8c51248edc54b9bb01975a788b4352ae0a6c1a6458a5ce2790e2a7ea7c06f070b7193a7f0556ed
z587425d6a8c2f12c8ad02288dc6ece12ab63c706aabcb2dfba7155a008e54a9250063859b803d1
z95dff6bcf8faac4a74cc128a931cc14cd560bea8a925577edaf3ac091689bd8d1633dc6d227273
z7979ce25920c0bead8d79498341da214a557e1693f3daca7fd620fdb4a43a8cfb3dabc31eb8ce5
zff2a6e8a4ab7869956f1f783053e948753fe3ab421405c719599f90e6a6007c56277405ec6b5b4
z8f654c24d6b2a874be9256e8174831477e3eb04eb03d24305869f910081488768baeb9c0e699bc
z72afc34b101a20b23ac2b131e68ec8b660dc6ef28aadd4932eddcff47651dae377f5edcc8e4bcf
z0af711eb4fa68a5bf0cb01709629b28ccb7382db344c6f59b05c9a1fec57dcc50fc3b22103e07f
z6a1262eb7891c2ee6cbacb8e065f89e77cdfafdc62354dd9e8cbfcdd6475df0d794b3bcaa6d69e
z7e5354eee3f04663404460b2c887961b592490d17322f71da83928f675d2dc6094e81ea0ad494e
zdc75a62a78e977f17e116d4128f8dd430d7760d484d5a9f3885a7355fe84cbb80cfe578bac5f03
z8303f1ff41bbea131e72608b4d7be332a8fbd112d6c6c63f2b620046966fa58ba4b6efe94d8b8f
zb6c762edf210c0ccad912dbef8f6ba223f42982e3477d8dfa2645e6fb3b87eba8669ae555a472c
z7dca15cc88e203cacbdd1480f5493c648ce3039093e7c99db6b77e0602537f8b01d81b503fba6a
zf12ee9124d9f8ba4c94901588944d37bb4002052b1a3aaed913f759b152c1d584f70c67e1c9745
zfc0c8bd4b1c43ea72af4157d02284bdcad53823bf12e38cdfbc360b3d6e3ae6b22c6673abc2eea
z6ff82cc4b751fbf916515f77c138d32672f9c11ad32258f407219a67c51b9c669c4f283d39e238
zd1d9b12c1e55518e5b25e131ce320c4eb4049a3e309d40c0a8d82260592e57c7434ffec0c6616e
z757fbc4cc672c73217ec577d88964555bc8f20d855a71af24ee30a1976f5c954eb6b4f7e9e90d3
zbe4b8781a8b609b309bff6a498084ee1afbd7008d7a9d917d5aaf3b1b3b950a4f6d8ac5d4062a2
zc9dda77f0f41e33fc8dabaecde27414bbd1c79e288a7f1c5bf4e75a066cac4f08f208ccb2bddbf
z143b1466866b2968a3413cfc9510ef79c11f8f45c3e4ee34b77cfa693e64eccd9ed21eaba3f57a
zc15679f42c475b4c9e0b764f55a60f9fc3bc4c616e40942ad9f372b09ff52d2a6bdfb1ad7d3936
zbe846173585220b595e3038f5a9eb571b5c7444833ee4c8430e74857775f021f409a4ed4eccd5c
z15b65f04075187d81cff2c98fd9f7048f06d5c5fe093a864a5543310d3112e264cc8137c2c80b1
z430bd7dff61c163139ec06e57c3085fc8774c29aa64d4ec8bbb971e773f49e01b1eb7fa0972ba0
z01ce6591415c137416a74fe1d32c1cc6d41b7afb44de7c211be49da5ac9ab431c3f628b1001542
z6d7466bc9b7134f46c4fb0b1b2714aef73c937dfc0cac1a9d90bd5eafc6ed65713c27fbe8f5c96
z4e17548a104946b147967406ef6bcf0c4f48f774b99e1885c4cc89447069189f51d96fbdeffb11
z681bade0e810ea5724f78d52c61d532fdef4271c24dc56c17f289403fc667b2d6247acb5f0fb2d
z18646302b6ebbeb2d26321cee89cc8acf35d59e3fffa912f074996b40ed402f8ee737fa5070cbd
zd0312b301480b95038b283f72248fa35f918635d7b2d22c45016696b1177d42ee0738576aa6adc
z2a00dfea8858bd3778c83d3c2d3e2cee85e43f376c206064dc8be213ea96e35e9e0fe81f1b470f
zc1c06605fbaa2fd1c3f9e4fabf8b4c2fcb03aa0c4be50bab28170d0994672fbde41e08412181dd
z91b20647164458de24390575a38dc501f6ca5bbd38bfd49f08d99b1ade51c2c4942ae3f6986460
z9f10676a52b3497009ff746b99197c553a1da31cbd0fe66fc9c5f35f29f6d05f08390782a065df
z7eee4055455acaaf507c6f90448f0d26892ba93b99cf0991fcfd139367c8514a70a3e29625552c
z7f145f587134d0e65bb67d220110678d250af03d0f0bd5fb3069d122cea03e64f1d8986fad6383
z7ecd6e4b46ec65f3587c74e7955c5f6cc1b0cc76dfc0819d389b0e71fe6e5a5706d4df57d43f9d
z28b998d0cc19f3465a2bad9b924347f09d303174b5592da521b85abc815e46a650ba1e4cdc18b2
z4ff163fe25c6aa4b812bdc4355cf7ac40e138d97089a82145b9753f09c92500f5c5160200deb38
z74e32d3ec548cda7a01b3e33280f49eba5b03ca06763915bd7bbb79c86882910861123a7f47a45
za294cc483e5ac5bfffc981874bc45749f102b4e6c78889fce16f39a69b64de2d11afd520957f2e
zc32049d06010198a0ce9f4cfa63f06c10ee7ff774140be44fa990fcef3e618edb0b973a696786a
zd3d92f28ccd3436bcaf8aacce2a8ad2b630484e6134b262e93f47038a69504365009ba2cf9a4bd
zaea6734914e9132bdb127e8e1b8defab28ef4b09164213b70e7dbb0f86311785a04375c5dd09d5
z6e56d2afaa07e6633930198d1f826fbb332e06ca945eaba18c51aaf24a594b0e764d255753e8f5
z963b765d9680cf57dc5ad4f88fc5ccd2068ada5e4f90084758be8c097591b8fc65a812f530f2fe
z362e7dc6185081fd3694eeee49b3522b0f66fdea2ac15ca36c1a2c52040b9f273267d42985f109
z2097da8af3492a2676740954ac304d0cf5ed2b065bfc02ee0634c14d027c6f03361d2bf71040ba
ze2709adf137ea364302760b74120a06fbbd38f1e047fc071bfd23e81eacbd962fcfd638c351fab
z7b72ec677be4b187d2ac34b9e306fab7461cdaa0a305b6bc913224e50f1b071bf5f21a7c4a9fdf
z08621519e00b94546761ec9a17a0d9dae9dcf260826c45bf9bc6baff9f8ec953851d159e4c3614
z769e4fe2e032012c829b00e25dff21ff68faf2a617f8ddc9d87ef1926395a3421686683f7176f5
z95ab66f6eb7438af23905a28fb0da39db2fcffe2b2ee548f73a3a9e83f1093343629e7e7e8c2cb
z6d1918414b1a20a0fc557517fd40880facd70135aac3e5218b1dbbd94580717f7274aa84f640e2
z40b3739e160b5d8e3af74e171cdcf2534a9d9798c067ffc2ffc26ee4d4ce2c961d68c454ac0062
z20aa861fef6c7fa5ab87789f478eb9db3ef316e07438005a5843e0353518dcd1dd8003ae42918b
z3094e963c5d11be333df33d6f474ef07179a39673fb64ed5f1fcdec26b6cec2e1c787566a8690c
z98eb739411d63d62df24e71bb72ae4bb45f97e936c985a4d839723688f42d8fa1e48c78ffbe13e
zf0966ec6852965af778bddee08c19f8349ad09f0d092c38f3faa065e6a4cd63a3cebd92489e9af
z2eae926efc1ed9d3b6917a3a8ef9ca1422246d918557780c74ec35452d08ff46301836d26a81b8
z0c4a15de52b5a3bc62cbd67d0cedf2303a4b5134d94cff3e507d674247ae7bb80e7e87486f9141
zdcd4bf4b24acaecb3995296628c0ddac4863151a967b7b75e052411d407517020db3b8ae6ca88c
zc2fb8ff9bf0adeea6f6cde6019f9c95c2b1f3aa499e3bb7813b451e71d372fd1f979359d25430d
z4ca715a62bef5e7b5a469bd3e97dc8e58b2aad67bd4cb7896086999d5975488666793f677325a0
z61177a768f90b3a1d0c318bc92a70f6a1612df516e06a4cbfb8c77eeffa100c6f66128f2e0b798
z94c5f8385971200a1c7391d3e723323033c77fa541085f431760c410f1732b6ada75fa99fbe31c
z066b7c45f3d05f58ab4a9d96b1ce6073214d09a1eba61b276652382096bcd99e41e4f388aa020d
zb865345f15336b7fc832c10b55066ea972df40e37734a70d2f4d92bca5df177330431b884a1a0b
z2cd31c59948634a82656c3cea48dd9070682fb47395252382068c51d6f8e6965e33e6248fdd764
z53e281cfb7cad7742e0a87939dc96550b397e9af4d04de39bffdf8a745c01dac87d2fef7abbeba
zb4709fce7d718cc1c115449aa25f0fb324745903432860564c8da677f4ec9bb29f749472d6606b
z2b0b393d54f73202658f170e5a87d86fa3a3a9540d7188c656d32fbc526b1d7ac800550c0d9590
z5312226c86c49925a5998cd729c9ef9abdab5b7a004aed2cf9ca7a8982f447b36fa09c54078cc1
za5f091925746010ff72d3c2b541e5a6fee08bbcb027798a146c6a49af6d4875533c205c50d75a4
zb13bc4c1f7adb2e3cbff8b079b1ba709cab3604ed3754744958b1ff37724fec67476ce1938bcb4
zd8a15eb68e598bb57a37f175478ddaaeafac706ecae44a84ee9f0056438a5823fddef51c63b7d8
za9eb84ca9cf7d256ba20719d894c0a8efae4bda7442db57a6d9d81ae6dfd6ad9cde62bbf671d0b
zf39f016728c9651be587a745f6eb980bad81b467b558acc7c4ecc0af2c78ee00eaf18ea04b8a2c
z12613065e86207f44e5a3031aa9aeb512070ccdcd5a06ee0aed0e8fac9aa60cbe2bd47a176807f
z2ab16b5ef7ddae28744b51d45ce91eb35e501a1c913760a577b04b49f21772e7d43378dec3dfda
z55af967d4b839d1e0060b78eb59b03f836b262567d1604c7903908c3b3ef585cc456564f5929bc
z648a61abd08eaf8067951587f9f97eaadaf4fb111cc2f9d21bac913a5488ea794d8dea21b92c09
z01604d184b57ad09b8e01d643a05d7b86a5442c908a5a0f1d0a4438dfc191ebffa9d32afa1e061
z9c2c267a327b44bf48a1104164f5a9a44467507d6f3e49321aae65fdcbe119c233eb40d000a520
z87b8099e905ffea64754e529e6ba5ee0287c12772f47336b28292e2001f6cb7d840123a4ad789a
zfb0c806d6784cba68250f6e437dc7c5a2f3bce049d273e7a7250d1467aa2e10c15c6274385a787
z91ca4897e8a890c626b5dc825f25ee765e25f0edf004d35668fb70e27ea5d7987b2d49cc5eb3f7
z66d85397f5875e66b8e24466ce3f26ebb5423f7f51bde8fe206c4400b0b6e52523aa06cadec342
z0dbf0057076d7913e3f5a3413e9e3aa438617784701bd5d6831abdf6b057b2bb363dcef7c7939d
z50b8562b71ee34314e118e55c89b2a923a1ac138464eb8e5ecdfeba6e4e782ee0e9a2297433b74
z151147313108da2b9015a93ea20624cb9b024e2b561ac853937074ac8071665c3c8cd846ddc944
z6e92f123623cdf0eab2cd34eaa5905ca2a6b8a01e6e90858a87d32a59f81b815daf48bffe2f485
z5bb262b36d7501494dbdc2abd9543954c81435c684c32c36c39c407a54717bc61b765e450c5436
zd767704d9d1b2bc205092e0382711e954d1f812f76e537995c769ca8e9697a876ba800e054d4c5
zf007d41c45d815c6d84cce78648c4b541067856cc5fe22c06b5f9a13b1722399440e7b9c073309
z3a9ffc02ab940e15d5e1981d13734720baa20a25e6aa820340ae5f32790c8b85019b18d99db31b
zdecfa7af520ec51f517e99e67329458c7fe0fb4376aaf384a968bf95d44069308ea3762522a272
z2a6a7fc640a394c2905f4a4c83ee49a17ab1534e35b122bec7d5442aefe3b211590a822af35067
z527cfea6b46274552e01cbf8f7bc00a9f0ee303c57ff867e2e1cea8054c60f03a5222d6750cbb7
zd19d938a1bb9c68f06b9cb2f2afb1323e0ee2b03a6f73c7b46dfc3d83acb76da11e525d77b52c6
z0ff08bdc5a236e9302904cf546372a4cb3128b7ac572407c3e07ae69107b99fb9bffa6f59a0728
z0c3d656549f1512322a7108f113716c1f3d358045298c84ef8a36957b21c3ef6c4b03d58e46062
z046d5b151830e4e6265eda09630ff75e56dbda2117b896d0cfe71e794a7ed7307121e87a562107
ze5cd395fcea81efb224eba57aa1a95b42978982525f6815390aad9151e8cb6d9b83c3cbdb4159a
z83d9b2897d8d2272543333f2e98f307a4dee0d8beeea86c484635a3960885f343ea51b6f171530
zd6e14d2ec7cb17c446afa831fd019221c13463fbf838b142070381e189cd86db3ba28821fa847b
z00cbd91c765f8eee684c1768c67425d78867d9a44b214fe0d0fe1158bbab191bfc441d5add1eca
z3859cbb309445364e1f7f009b6f001a23db26ab8dba0bec9076400012e0e36fc872df3325cc4fc
zf442de6bb0838d18c280074deae2a2049bf533c2bee23610df0ad8ff038cd1bfa354e23aeda87c
zcf534f8a38d4ea7e76d5a737695de2b1720c67c71f14c5504b64cf1e77dc7742531c72564e459f
za585ee80ffcea288862677fd4f040a5a6b8cf613b4657f878c7f572589fa0250f7c4c881a7ae09
z69bc111a99a8c30ac1eda8c4b31bd2d0518d83c4a984fc012970e42bd0c1a218662c6c4da811cb
z71f97621e83aec16dfb94d192c1c121e1c023d47812495d719a5d44759cac952c63d804529e044
z92704cf7d45c08439e73997cf25dc37eee7cf31fbdae64f0a938758e76865b99c179a0215da52f
z26f1e94e9225a4557230154408d3f00a13d86ce22fef8342a4f336fae0d5da698b0f9bc64300ee
z503be336b848031366ef7a82097f20e35f25012d2cbc23f635d2e2cd5f2702d1494aa38c2c58b6
z8da21298f31139b1931020d0c8c8ec38864fe2ed8ed54057c1034994b5bdad9856e46d6be28b37
z0baa32ff2e81ec0e8f42d335ab7edfb6f824e95aa4d21e7c6fc74017c799dd4d28b83c2a5bf97b
z78494704debf33c7214aefeaab01b8aa79bbc8d66ed54a368551f9d97613cbf3e9472b5ba5d752
z51b685c708b0741f1830e43e8ea945cd13863b543d576de8ea45e3d359005716b3afdc413c35ae
z7dd5bcef302231355e8a6511b1a879df128bd5aa9c9fddc8ee1f4d5c8b5f2510a93361722c7f9a
z22e7be9e63fae67f6fe676a32f939ae0043ce4b0422545b3a036d9a992116ea7483a58f44de2ea
zbe76ee6c2c7f931116756f8acb6a1c056f167bfe9426a9040232f5ac27c58411b103dda1b11b36
zfb79df7c62bcf15d3bad381ee1aa6f9ee2e2a148d0f3bcd28d0ed180c9c526cea1358dc89289fc
zfa0f5eb50e01aff59cea18b6083befe6413f8818e1d368f8da70067cb56b76618be823ae89a043
z50edf967849fead42ab4e44baa06a68fa4de6d714015dd85763b5f236cbda794acd4d07f299c90
za006ab0c67e6438833cae922332b36cfaff9be7516d593ff7a988b98eb3f90e7f23d884ee2efc9
z709335ac55dee6541a64e4ffa4f8fdd4acee351ea51f88e34d567a130ad783b3c83ad2b1e27be4
zc150738132346b16f288e89221b70227b7bfda54e48701df60596ebd27f21a1e6ee986f12fc10a
z769e39407cef16136172ed66a158cf5ecea4ab8aa0dad2d8a6b3ce772a8f3ac397cd0e57fc3516
z8b13b29f1b1c2a3c94b4f7464c5eb17af1e7e9063e6d5a189c97cf3a69562a637eb98ef58b2ee9
z6145b2322f8ebd5c19cd537b3005e3348f0f99737a80ee6c4a80f485fc90ced16c2a57e935f69f
zc845439d0b2766b5297412ad2a7e9179a2cbe7774da21287c5970fd43b6eac9eb03bf5d6550aea
zbd958887afe9502fc51c02ccead314d9582acba1c2dbe99fdc20a530d8c05b2942fe5e3c82fd25
z20684633810c49ff02a7d11d1570d963d5533cfe3a0e061f333c1e66a5ed2c865bdd98907bfb90
z9597290b2e74fc09449322e2178ff0e8f59a3967d92d847a6a1c49ff0ae626712989e74d7b975d
zd90515318ec0f3adf38b66b543b4433af9fe20a1744a2eda3034128933d2d81d17aeefd84229a8
zf34b03d12da30da88534a3f0212321a3ec6555b0a5dd718a55eac496b311bad242a556d6757989
z73ac71d0e9d7985086b7648baeb6173e53ed943a996170c224f90c17df2aa7cfd0d27fa08181f4
z6912e65ca52752f02227dce26a10777007fb99c2f56cf4146e59d0a79c442a3adca8c939947d72
z1e8350c67a589d6aed0b629437a054561fcb18ca5959adbf4e3141ac0c27881dfe23b63fcb6424
z487fad77e830a6d15c68bd99881b2619501908683b6de3ae57e14f2a3612f2adf33185733ee410
zc0d453511556482a9e9ffdc1c31d6642c2451207e574378988520fc9180061f1c75282835f5e1e
zad2a679e6d46dc993b9e6e1f86f01f51dd1eb2ef981553994606771b8b0398011bf42a47e37523
z0ff953fe009ce53306206b5b3c264a21c4c54278eda93a86a894851a1be3ff927104574e2b97d5
z7d06f3c4bb9b3bb2d63f463d8c71c0b831b3b75aa474bb1ab5cc8602cb60da0444e4eb6a811121
zf83581bdaf7e4471ac385a147957532cfd3c63b410f896cdf9d758124cbeff5fcba66b6218875d
zc6f728b9dcfa578ab0d6aa5db27f70c3b4e9431fa7b761d6bc4c4827a77ff8b111c40b77e58beb
zdf6dd6ffbcab6e954a529f2afc401da2d30b3f4cc2d1600c2e644048fe8a8b36dd7c587aeafac1
zf09e0b2550eaf7615cfda3f738b5dfa1ce2a39f47555bf5f366bf247e15e0b30e48fc46dcf4f24
zab8e56ac0f54621e9e93195fa67e288dbaeef22dd0c714b8451f9fe35cc956584a6d6082287d61
zaffb56db811f211c038e989ba57d2025dab09d2f00c25e21340a2a5cbf0a22a09be563244701b9
zda623ca46ba0bddc0cc765ade419990fbd67a8fd1893a55c9cd2de69b57d3bd782a3f546a6b9b8
zde39bfc74e6946c144101339f6262848aadf81738de3a0f59c44a1b2cb17f906e1de9864b4e7ac
z8868972c2b4662bc23c9716b57867305ad406a9e75b52d5dda7b47133bbd8fcacc14556bc4cf36
zbe5555a7381cfdffb426fe7b55e770b64ceb3e4cfa270a0e4425a6ea09cfea1747efcf41eedc55
zc7f8db9dcaad34c1fe21ea82ddbb30e0277f5ee8af0b2e1f11b76900644ed8f918ce84f5b09b11
zec52a4b494670bdf18802811140743257becc869fcf550ea929f4a86849d01513a15fd8d0b17c5
z05f689258d1405d27f5ff2a25cc9f174b2c7a2a603255d863013eee8ea69c3d1ad5b71209c34db
z32a9d06510f780f134fe53adc1c94a582cd88c7be43572e2b27cd5f8bf865425c1efe21dd9a23a
z080dab1354de0c1dd8507a14151edfa7df1a93562d4a74950c2b72f4e32cd372de2b88cd099ce4
z629b37ef94c93c4550ac4ccfd3c4e1f100096f4d5ff70605ef300245ee7652fe6436fb91f77a59
z3462550dd91ca88ca5ea69db3292b7458bb81caebd126d3709f4a26037eac2fa23f5f7872070e3
ze2e11dbe747ff0e86c79a335b271bbd91e24a3abcfe2d5a2ac37d0ad001df428f1b7560a9230e8
z16bd7c361234a6176f716df3f7981eeb519a2247c44481fa03e501eb530f2f38b463f6f675dcd5
z791a71d6bd3e7487b2ee414107ae80b18e91a7cc9b130ee2156273e121474d6d34c7d317f6265d
zf3332db8602b1e6c1f5ff6d0a6641b834be4b77357262482782bbe062f10c4f46d6e83c697edad
zdeadb496d01b285888aa39870df7e26237db23c765e281b0060adb87142f83ea59fa4a0887c72e
za6f767f62c4108f63fecc6ac409200efee66ecac16e6c4f88ab5e9d1f61c4205f3ae97c8e3396c
z9b49f11ab385688cef499ba813643dae63205a28187a37b5cd145f834cd384f7a00c541ceac8b9
z1a707b8b9fc62bbabf976db2b2dbb86a1a7b655d79a5712178d88c6d6fcffab7187b1da1654908
z204658a9fffa1d503261016506bab77855ddbb7ab288b67291bde870048ec363794c84fe9fdf1e
z4c32762bb4b491fa8a54054b01399e4e39171cc15bac5b6ce632a791d6eef2073b81cebcf78922
z3655012ed0dd118afbe7feeeccfbccf3e07a7c8beeb6851c516c38a11241b38389efefcce2595d
z237ef209d81dffbb8ee826c521a89abc9b9d6e26cf3c90a752e91def81411e8500396d46f5b660
z39f8ba6442c16e3592e725de0ebe10d2a3518d11c52c50d38dc22d1548f9253c3bc3f2296e1ade
z686fe971a3cbd0e300af8618f8defaf602e5f9426a4b0f744a2d516ecd3f491eaf207df077ca86
z1a6b2e3a5752c23dbc0a1ee481d13eb42ae0d8f0f9134893f694dd2aa7ce61d5986faf98eab635
za4b1b6aafd631560dd76c8d3d177cb2a5aa99081f33bc0a318b02e8237d2a6bb262f39a8946048
z52e779b2094c87a34f9ccf122908201a8f3cbb52af96288aa3ad2ec8e089baceddd8dedc2af5e7
z800d16223019fa14633e6770472ed8553f764bff8b6a101f9aaa59ed9b143e76a1ec6139dae73f
z8ed36c4fbfc0719dc4a9782cead91389f4e758e7e841597212ea482e6136df2dbfdd0c8c0a5e9c
zef8c9bbab736b97dd77d2d22517868cd9996e7b92fdcf8aaf5c45fe6cef731f0d2a57018afc855
zdc882c3a5cf098baeed23ac702323cfa5951f6602fac66c1b562451a5e5248b5c1fc1893280da6
z2c8bf391c80018aeed29330dcbfd9330b3093a9129125b9f58f6df26ec5194ad8fe67dc602b47b
ze779798305894c9dac0c6271f35a6d39bac956231c7819bac052240eb186e955d08f31d2537a62
z417ddcf60f31f3fc94235ef5390bf234a22fc645765aac287d092778831d7bc94e547e380e9916
z1f5cea1164174bf7d5d1c02bd686a436f24fbb1cd35422ceb1afeeea0a69a212cbb0abecabdd82
zbbf6e3697dfa0338f91bf50c08a1783fd838dfb268831595ff45869f26ff2204fc8c5697218f9b
ze8d5c2fd4a17d848054015d339e8b31dbba182e095b4e622902e661683408566861e56aa775c3a
z499798de41900f5e89e7bfdcba22423bec1fd3cf0852b21e90bdbebd9302fa276579b804f470c2
ze0eeaee956646ed61b9bcfc0127a95b061e07d05de66737f3be02f9cda34f92b54d8c044a54291
z4dde0603d110f93fdfa9e73227222ae8ef65bd66efc8d1c4f9de569e62c9795ab793ffd25647f8
z039e76c1276b0e3e560a595826b87abf4408fd00a477894752fdb6085a652e3c32a44d8053f04f
z206e902058d3b8781c8c0c37cddbe9164ddf6b4ea2594d85d5ed334634b5fe6422545596af092c
z42bba9501e2d5a401077375356041770cc906d553b5f0a1b8872d555810d89742029355adc5230
z793fdbe4067d2c92056dda6e1ee2e2ee4e8729e741ba34a5fe52df48c73147662813dfac95a512
z039e4e75e8b455705a6aab3be09ffba236e6291932c3aa7c28c7d21e439dc2f00aaf56bd1afbdf
z5af313815ee6bbf79b6b6c40958fceca7840e492421724cf8837e54f14868ece1bc082a7d29d12
z1e6056bfb20ced1b25cce5d9ae290468ef6c49495b06e50bac430ebb56fb23572dfdd9fe222f03
z9b2824caf5308c4568b0811f0a8dd5cee21a0caac69f935276dd191f939e187ab49a297a146a17
z6192936ccf00a11f9dbb7e8b865664cb6a3c73564ebefc74efc1a618dee90d9a49f20ce9f01b99
zea46b082e67f916d98ec322eb4c77594fe115ceb7ff23888db5c2e578ba23fee223eefb8ae39d1
z9bdfc8d8a6e59a412595f9a54ec16c4f634df240be0b3adfc330ed34ea155152de718e4f825276
z6aa021d8153cf18ed673c2a798784018f34d51612965f26451d2670b76a503f908d18b5b7ee15a
za876eb69f2765c8b06c1f67d4941104343ccd7e270a7a8386c5b948354eecbd2616c7b85cca426
z5b8ea3f6f41627c4896ff15942d83d134e9a555aeed676b7e108fa800005e67433d8ad2e2c8395
z5a331403e73c70abe37a46a2f2690fa61f80ee3d12ca9f5e52b8882c0cbe715bc01f0c0520c91b
z95fa48fd34917c18f09a336f57a64fecd47a08058a79cfdeb6bd7617b7f27fcfdff398399e9cc1
z870294e78b9af2e48e69ddf39a02c082fda19906569290a6f93bf5deef79a570ecc8bda592e34c
z92ccbc43d580a600945761eff71114fde878bc94c177fbc18de950ef8b33d57956349a01412f66
zc3df05b36da87d89d74bd360ae3f39ba0717dddff771928023aa2c0ace3544ee590897761fd272
zc00a9ffdb94d5fc4b324dcb7cef366763fb1aa662a4c5fee8f697b81a18a6bc171c798b6ad5aa5
zc0c088ec6f883274535ba75b77d298b17b77115dc96411841c5199d59b271e6eb9fe5279781387
z14bd5b61725a9da082d516b00663aafef799b3a3628f06c00be8963159189ff1837dd72589a55e
z2672551031797e46ce1ca6ca7643e477c94bfb8afd2518e29dc93194a0cf14ec48159c1ca45906
za6031ec3f2691c0712bbca5b0f627cfbce37bada261e04d4f60d865d8c1b05cca4d343a8be4c46
z6906f4f42426f83a6ca5bb1759474b83c8cd106925b11d4eb15439dce2889a86fa0c2a76ba7b83
z42474d6b8e83df3e3f546c46a4b2d9ee904e05bea342f8a246edb7ae89c608e4c1f4bc2a2abb90
z03fd94cf8851a871ef2642e15315028765d2227c5e9dfa7a2da9baf7b8372932effa594dc88454
za7e01f468209fc9e14827a4eb47992eda1176feba053ae847e8a95018df3c2b71b91eaf2c4b9df
za76c284a8e36336fe7b1dc05af683aab1988210e91f9e34ff3ec2c7587fa9b607325e946d3afa4
zb56b4dea4acd29fc18a4a073c62c2a94729570e4090c0ae7b268173998bbc64cb6037deb53a525
zc164bb6b3a4e5ad8eb3fb6b504936f6a782cbac42d7bb0e1a71bd5dc0186758d41b65719107366
zf3a934cd86db7493277d6ae38e33a6beb897483961cdc32e77f1869becd857572e9dcbab43bd98
z5b115ec96a64beb3a0f48bb5cee821286bef69c6f55f1303ca013a4203f72c9b060bd91de28edf
z2abcbb0f2bd5164465f763130e4b07c67669e71783d57d121e1b60bea0f1a9606d09b3f50b220b
z22aca75421fb02b039f5f68103f7966fd212bf4217799cd603d5d4596807a85ab9e699e6b0224b
z82de11dbc1040a39ea858dfea56e697f37673d8ee493ce1c18c51528d4931985eb64b359a3d20f
za254be45a728fbb9b7e9c3785c3c7c2dd95098b75165ad7ece3162088a566105f43dd5ed343c5d
zefe944509fd879544847d71f6845a26ba8ba0e1692925e7e1b0ee357fd3fd5c9e473ea7296c511
z63b74da83ba35803bd9d35967447c78e8f0d74deaf6a75bcc681c8ab82311cee125e18ef33eebd
z5db958b9df45e11a891dd279da756233558793ca30ecdb926b94d04f81f558355637cddd050108
zb957b24b8a7295f125bdc22bf13349bcc0c6a4db1d5abf668116673560750344bc7869318c4c66
z7f033643df20c18906d1e8f7d6e10f42e970c194c9ae45aaeafc80dbe10fbe6c000be9ead215a4
z0830ba2dc6529d1cd5dafb1da5a6178a6beb1636a3486b3b6db578a1010c7211eb454c3d713545
zfa1db1b056462c62a337876257278a808a81276b8e4ddfd9ad61647a195fa2b2a0bdedb73aff5e
z5298e0041efc0cc32828861a21a3c5bd9431b9f8275bb9d8f7c8020e62763b8273a8d69a18e821
z6a4efd80505c05c4ab95073c5231618f39827c239159a74825965f0f64b500892f5d9b33417f00
zf901597c9e9e2ada06a8173983c4f65e52be9ea07bab95e35878f0f566012b9f12a4dbb3d7597a
ze5a32d7c6b9d483df325f431da6c53c427bbe0c4dd2725ad40e6c83e8653dd26631a218e4ec234
zfb7e0da34f83dfc518166a388078ccb66da42b788029ef1a5d9b0a9960fd8710e41b1d682c12c5
zd2f5e683f4501baffed081ec4fd3a846f308921925c96fb1a0df7db366622e888c05fa87d262c6
z15afbb7e4a5f2c241da29a3ac47c16a7f9794b1ec259630dd33c2a1d927160d3ef9982c7537beb
z5deff35afb297e88d389de42067ab9cd8d378c18597f31363a64673a72fe8748a1a64ab472f4e6
z0a88abf717d3246d758538a6f1251c0b641cebf769dbfac564fdd420ba3552237f262229713f66
z0fb8e437f344b1f01390541dc57692eb15390e1ffcc159f8e03be8390be21c0f23a1c53b52f62b
zf7abbf8ced1b56e15b316be90483b6674dd61d49316ed70918a964b271c766ea598b044674648c
z3c319ee048074c241a22e4eaf4c2cbd47bee824b405962a15ad6aecc964fbaf9b457b55124f701
z7b79d4016ae53407d2bef046237b98447fd6052dac5e297e74330d43d5ab223dc8333d37df5756
z8c98edce51dfaf943010495c3f8d0ad4e2db0c956377b9b9f19e73b6079556e9cb867d22cb2df7
zfa69985ffe4c3932e9662fec1a68b10c73a04414843219d679e07a647f66477b5cda1cb23ec3b2
z48e930a3da5b53204424ed5b89fdac5c0ae90ce66858eeaeb7d2c821302f5bd71c50f6f39b0e21
z220d7e6f1adcc7fb4da23458aac21fd03e11c21b0511fbd63cca0ba39e782a7395526d200752b7
z71e47c26bd29e61e8c2e9102068956e202c3a872066dd962d0570f1214209e32404207e795bf57
z40730b02ab80af373979da3173b87be9558a974c321390f83274f4821fdd26a46742f0c6e3eabb
zd7d2b3571dce1f84fae9ef194c647785820708b6867a3158c961f7199ca07ce1112a14b718bffd
z8bfe09556227084fbbc4d2f8fbe7474f9935b4fb3a5a0189f31db0d2d36b69cd6ff5f0bc19a622
zc990f03ccb8d1b429f0c2d6429e5b582068784f96f8bcfdc00d46d5abf062ecdc503fdf3efd7d1
z10d73ac97e365013f3d2cb54f3571859b0a6a0bc9657f038e96db59892f40a6ae17df96e800655
z0ca176ec56d3dcc6dc88f944d7ae83b8d71869e87b4173796933b61ea2f1b23de1c5990e5a8c3c
z91786c4883ee62dde335fc5dc6feb9d26c2f49e1b6b36caaa07a1efc14b5db11205c7caac5caae
z6f081a25a4a0edb71213ead97ca1c618e6a88f4dd7bdccd5a3bfc12ad3b8cea2cf0d5b97df201a
za6283404470fa928d7c8ce6bcbbac6f805353903e15ccbb2e6e59d3865f1211afa895c774f3f17
z10854a0b2f088019935b6e521209554a425dfc3e39bdddca148f1f24a60dd900d8c53d1d7dd857
z71d15e938d2ee0131727a62a09d7e72879a8d5d5b72d275a007ac2fe3e63826fca93e1175b7615
z7d9ad0762b3d55234a9645fa94e31037c9d825b817a8987daea6a8ab8e77ec193e1f1999fc78f8
z4c9202133517adee9730e93fdb0745f1ad74b525d4624af4ef6c94dc77caa1c23f6f1080ef9641
zb1486fbc5847a9c5cc08bfcaac9979b609c9f780e78dc2fb9a40555b98456d9a9ddbee084bc3a6
z106d9eefe2593f3fc7508696dfa3ff8267417e0c2366379867b3a2d1f3963360b27de207014558
zced30301e8930c19d8c3f3b7ed22d9409ea7c9e18a8472a26b09387b536262a7067f74bdfb6fee
z1ac400a6d736781862e2f9812d87c5c94253679e3f9baaca0e2f2a29598b112858c79d39230334
z6132af2595c9bc282d2f0c882ac43406f2acb711baae051b0ab7b4c54cfe9779655875e681c724
z2dc2335adb036769c56f959d276db72fed030a1bb120af1401885c493de2c04a092a955cd50ee8
z7da0582ad82f07fb309a713090cbce4aa4cc5334f8456abf856331d398a5b4dd8f16590be6c92d
ze4519f42a14c5c235804039c40500a2630dc7f8280471669a5bb48bccfd45ad180555aa7873ef4
zdd9db97212ddab069b532aa00fb6a2c8d538edf0eb895b262e0390b7ad06c89169a420ebc5f461
zb9a9c58a3942edf54cc459961f2674c15fe2c0cfdeb3fd52dfb2f16f1ae3e48dc87012df74b5bc
zeaf7540ebf3bd36ece49fecb8c9039a3c7a0702d17098f1e66c51a3315b455f19c263a8a177f1a
zb033a6c1eab40a63544f6b1d212e191f308da51a695f5da9984528354b440603d6c766bcebb0c3
z873792797dd94ca2343dc93d236e7d3208f47157d1591c6e689611a1a23e7e870815683e8c5c25
z18cdec691aedc14b3b5e1a5ff4c889a5cabd613b19d7bf25ff93872950a843238054221b8eba91
z7ea4561ca70603c6bc4927aa6c589438d71efd794a4e53e86adc8d020d2cc472ea46d6057b38d1
zc53b9a2b829e64ee0edb6a77427fdf6bbad174daddc7b5e5895fe59c6cb2507eebf5d29f042457
z71cd3ae44ae0242e6ff8e30d11170c885dd89b5ccba3529c28a62b36c87740ff9e7496d0567657
z819d0745c7381679b152ac4312061560a80c29627f2c1f89a6d2a1e24eef9518d7a84decb64a92
z0afb64b343226ca4fb4deafec18ab6c9fd2e1e7a952be4986580ae5ebab3d15dc54264f4221870
z9c0d75c6f78a719e84a535b81bfd582cc157aab59d1609b0bbebcce8051dc83f95073118fa8ed4
z8e407e40a3dcffa46fc59e0cc5d32ec62ec2935c88893d90e6467fc2a0dafc40c0625ef3c45c7b
z357955de3dd7ce1cefb5a65a349a650af99cea56ba88e86f0fc1beb983c07c7abea2171551d446
zf8fbcc69df5de1dbba05ae5859bb7267dc042d00c415df8baa84f2f29911f6d8e426651a127464
z47e9e60498c82cada760d4b9c9599c095c316fd0f56513550f6f8b205b7a472e25da6c03402df5
zf72acc22fc5bba109825d08e103bf1526308b628b70fb565c3b6ce20bc761ba338eb25ba7a2203
zc327dd7033a52966f323a6c61f2345729c58367f7d00e9930d080f61472a9eff9d1adf137b2436
zd421e640f0236feda598f4f5c013855800e66ce4fde77e7f1bec46faed0b00a7c687f1d43fa7af
z8bbf0075d2bd0efe76517e75f22bc26c6f69fe67770fdc03d701873845e4d69e94cfeb0e187c9a
zba2d6e8a1488a9bbd08a7ae33f7d0aec3d26a236aeac4a3271f1ae4d74e3e8366561d26bff9462
zfe2c44d275b0a52d3e6be5bc464dce83609d8ae14ddd6c079f058e2b18a84e59b898154e9fb6ff
za2abb4c9e093f3f9f8e60a35417252a43ad725df0ef4c2459264ca65326a73d7a93225282aa0d6
zd2404a36e936aeb19253e28f87cf1fde31ea06eb79fa023c3a8c92d1d750eacd8cff3337cead9c
z1629ebf91ee8a5ffa772ce680034499f99c03adbae35f0799ae9c23252d7aac903bda59827b145
zaa5ea122cd6748232c4e1108834a8ee59884b4d10c52df90ce6748c99a7a78f0ecf68708ee7098
zaafdce9859df7766e9e32900d1cb683a04d2fdcc93d0b2233876dd14f50290c15d65e2e468875f
z4f3de6b83cb684878bf677af7bfe2f9eae970cf1fe85126d95f770f56e98fe4db65230755be48f
zcf04dd5e2e0da9679026bbc42355ce61f37ffc915344f6e34733bf1a7979b9da370aff6d25d285
z84a3f71ccbc70e44799807a7ef5a6ce4ee1250b48c91c7cc9ba9f6d32220ab0a040bac870ae187
z9cb4f183bf92a29b967ae83ba17aa6095625373d0c6fbe7af4437c147c562871f94266ec84d5c3
z8abdff101fecbfdb392c30990e91cfc4776ef661816a8defd246a9041cb1e002bd0ba64be9d0ff
zd82ee9b1d34b25936f2c6b5110a24c490a4884bacd01c6e811fd812d9851733ddd0b0b83b9ee1e
z426926d3310ea592dcc2bd218eb085c373290c28220249437e5738073e11eb542ab3af31a21349
zd179071de2cc62181f74de5f74790efa8b7366391122c73869cf123357ecba35a9d8f809e4b685
z8cf5f6ef861175ae3768d5fb1970597f0723d72bf6723169c1f091f16806931f008c62e6760c49
z25fabbb62e5cfa47c44a04c0ff927472baf4876ee1fe3a50523a53bc87f9e31e18eae9880a20b2
z2619d0e1561fc46d38a0c84b5d63c5d45537666c4068405b1eb971ef6be3bc1fd7af8b37d58617
z7206f015be832b65a92091bcb4e4fe0865e3639da14c84bdf1a29b2af4e99d665436d229355d94
ze4dbe96ff374e6a037b11de591cc0d81064c7d175a0fb8b82414f3ff35d5e357d5df323f1f9ac1
z2ec1356230a085ba603a0bdeb8b7044fb6992a4564bc1c074eb65876ad167e11caf502486db59e
z917e577c59c37da8df17e936d7cc9444af3aae717edc934ca07dba44ae31938acecc92aa3f07f2
z449d15cb75c98e9c3d4b92e57758e4b499ef84ea11d3700fead8d7475d0fc3f41ba845965edab5
zf7bd28b6d24172611d6b3588049f0f6c8ae263dd7e49a6e7d5d858ebef55d66027c2caacf60e85
za1d989a1690327a11b70ef898ee094ef6ab539fb2f145425f81072af174356cedc550d095c2029
z0db27a648f6a026bf7c8bad33918bd3b3652018fa29de3cb679baf2ba2bca2cf020e8c0c8e6e31
z7c59ed5e42e9827a3898ba43dc3511f1ffad659ba2d3f8a6785e6ebbee3f5ebc6c08a8402f2d3d
z3e1fb4ae3d94c1b99a1e42a5bc23a9f34fa23dda43e092f0ad09a9d8a13ca6aeb9d8346aee54ab
z39e4d4d3e4f25d9e3f7fa24787dd32ed5a1c99619cb27d026a569254796bc0cda186cdb1e45824
z3c679b99e0790595247395bdafa4e6f809b7bbe462272316cae70f37f4cce3ba7c2d33f31fbcb9
z9d1cd780c509628c2eb04b6577853cbf6b4dd84bc0f02b07fa02abd3cb07e68b69c286ee5dd5ad
ze226b5a05e82f051304d1038f49bfd1721d43bd921fd3c463cf991fbadde84803df46f249f1658
zb465bbaefde009f7b3df84ba020cedbbe358c30c346e4515919289dc3159bcd0613f9be34a7750
z09aad34e143d77af76328c652f810066dd0d47f24bdeded5e3066bcf6ac966d52443bad153571f
z75aaa87d73ed3890db0b801e8188036ea614807d4f58ddbcd7a2420b279b57e610dd7bc0568851
z966af382b25afe9a8e31bb5875b5144858670ab2084898d7c6ae81b7316e83d741dd5d8c354591
z713756a563843de2f65c1b4ff461d7119518beaefe69fe8401f3bac897bcea3e17ab80c172deae
z0cdd155a5019f0ef75c840a8684b799699fcfeac3a162c49d435e82ef32a2b1fa67b206110aa0b
z440a5fb6be3a7efe79500baa940fd5ec382ae9f7db106af1b506541406fa4dcc396f9cf428dc36
zf76db563eebbc269cd0561074ce2668a71c69020f2a629433583344531ae2b53934d4dd126cdb8
zcba1b743ddd52ae1edbef0ece7583dcae9f2270ea72dcc22275e4d225c511674d5ea5ebb81f0a5
z10de7071fefcce1fbb083eba390dc2728addde28ecb34ad896766322348c8f57f43e4d0412a687
zc244dae763ec94991d74afa57496ea2f7780f9ea730129f18ff875ff6023bcc1732858d25e737e
z942faba7ccded9e9ac08582b3b8eb3d4e426a9bb0b0ee2f7d97d27895152f231487704c7fb7371
za27039380069ac71d374d5795209dc2e28055ef20c540bc6a554a5827c93c5d20241b6530745b6
zd6e0b5cb03ec8e416e8610b5ae7ac7088e100cb77932d1e6239ebf0b3e6e28438ca1bc96a9611a
zc591f0cf6dd8e3dbadd9f7bf9351d07c6befe6444d30c27c2dfb8e052fae7ef5d7d4fa74a5d976
z09b76f6db5c049111f6e55419a33f9029886ceb87434ce9eb909e75ebdc16cc57c35140f31f36a
zff8eacd5e0c48ce9b678362f360b9be053a69f9d649a047245be661d12a9092a44d6caf362ee52
z1b0f8edb787c65cda4e2edb6ca5aba07cbf03354a608e740b52c0ceb8c6236cf5adcf9e7e1f86d
z4ffa74ee2abb469ebf92157c7f556dddaae733295c44fb0a180a11771a07000180c2a22a1f6434
z51644502b89fce14a9cb3c845e745a2363e35fe7f9a35e74c48260fa428714cb67a9f91e8922e5
z68c816a61620645849f7207dee511fd647b11f18c744aa2783f2f661fa59f62347715f6e3d4ca7
zf8a05f88c206cee8811b40c3cedfae3ba4f6fa365cefdc2e3218891115e2f60abd6f2dfb271f12
z2b7f3834161ae87f0f1586608e53870f92d60dc0a72fc8cd4e0b1a586ecd18fd61e3beb6440977
z726395f0c4546974b0a5916e12c68bbcd1396fb185f527b2bb5e0fe644854379ff1e3508c4e785
z0c8e961cfbb0deaf0ef782f531a1f4992e94b78bf0546cf728656fda66a0a18cca46bbac9f3ea1
zaf5a9ec98e93ae374f012e49e6d4fddbf067953445bc25adf561761378fbd0509d9819d3464103
zd70c86914852c1621bcd3975aa6b428cad042807e32c32e60e8d148b18341e92e2a4f940d4b77b
z497f9ac3aa07f2f70184a521cc7736a33994f76ae0e4a7443ea519b02be2e1bb520a6c767e557d
z670483231284f5278db0bbc1fa1648e1a37f20c72efbb9c66e61f031d2c08337b61cfcf474bca5
zea00abdbd47490bedcdbf73b068a2247f37965e26035ac6861609d677178854ec4c46520a36bf2
zc34f51856dfb4860fa46dd088fc4b3545733a9ac908e3e2f3969937c4f04c6cdeb98e12b877e01
z8c9992c2e99de84a36085023080c4e0306b22b6b71f88cb1ddad65d12b9786073a3ef249e0d3ef
za1bd08560e76894ac6a23e448822f2179d717850db7814b7156a5592e682786f8038e06ea823ca
zb299e453201ac4f0349cd0da13760c5ae341feb5df06bf9138bd205255f3224100be0669aade14
z476c7c1e838e6c32109f6d0b6073286f6d3baca6ec3b34ff5e5f31d81b03f116a7ed4fd62defaa
z81f1ae0f54f11702992fa0105d0e5068b909843835cb6c4941f31c08ec293fe30892472bb27a4d
zc3bd4546c90b1edf2e706223462aee8f9555e01bd5926d0bb83bcb996440be616c6d7eb4ed5851
z8615ca96b3a4e24789832c0eee34b8e233db69e5752c42ea59f69bb45c051cd0b770d4cb994154
z2a553f3f3edc39a2e4e59731328a5a2473cf7018f5450f3f95216b887d0a5cd94dd2f23e2757f4
z202609eb107bb4064be6bccb8f0b3dacab373bd09749a4e67ebda0bab9cb43bebaa7b318b354f5
z03de255134723b070d5c193836dc2dabefe954fd28cb0e4159eaa85177281dfcd7e25fc92f3bfe
zb54ea3751136195a8d7917b741bf663f3a5f65ed1f86794e495fc5ef0f7e999d3a512e66677761
z497198f508d5a2cae9300c70005448a1cad8ea0cbced3008eb441e64fa6e0748b31bfcce6ca2ee
zccfa02c5f41a976ad08e20fbdc3567163bad76e0254f4fa26e52ad6ae59dadbab0652fa842c8bc
z574e3d587000eee8bf40536d6f8aa825382b7a09c85c91d6f40ed43bcfcaed29644caf85a47eff
z9dc7c035924979b4d8cf28fdc8c5c77068c15a788cb43f5800761a61969f502afc57243abd534e
z1b97c9f94a700fcb9eaf66eb0ee7e68a5006be989916cb869a2c211e01da0cc96e9db3cd256bb1
zb2b7d3208473b4dafacd7c97f1320a481e5dfdc54469b658994620bb67e17bc5178f9d25018de0
zf14a2c5fa3f9acb0e43f7d5360d74a4d3fe45170c2b6b707252d866748d575e0b9b86b8be02971
z9b74cdd6edf61815767c88bb7a9cd3722d8810bb986953cca9e0c29246763c99e2710d1c2a8d5a
z66eabc4ffd8cc6d5b159dc18909c69bab59c6e99704873662938061383f979473a9e5553ab038a
z575ce5f952bf014eec7f20bcddbdc2e5bafd23428c62d6ac880487411c7ce2e74f02009149cc8c
z54c746d42d1327e140198b5cf023bd84abb8470df050dd19a66c88f2a58b071453510f7ca3d44a
z90711cc5fe3891eb4168615ecd79caf07a73954c2fdbb31f3a325c3fd644f62bbef7ec8fbff81e
ze7cfbe1e881df8ebc19dc538cb24cf43f884a5cadc6681b49fb48fe619f6d38415477b9042cfdd
z903f2eb616fa195976cade69d1c92f8e8e07f35bde63d70312a6b1800fbed21798bdf395ff2f03
z9bbf85ee3d9c5c253a57c6f54f761600d0f595d07b31b89a20fa865d4abe69a78c250400065dca
za7bf60848830d1ef3a422d7402ffa5e7a55327326e294def8887020bf0b8fd8e00fa0ff334357a
zc16350f2fa99e9b674597366b7a7453c523a9b3ca2ab0e918fa596c8ad7ba033dd3aa9906f0850
zc357f0c63ef7490b12ac76990c3bfd8ada6a0553d6ddf4b289c5c705f9325fd58472136a3d9583
z8130282a87616fdb461d11cfbfcebd41fb05a03882d81ce7a14cf6a940aee2960f14efcc2be2d1
z85764bb32c9b76d43b48c5157e2a97899fbb205d9993707e5a8e24cbc87b13bb5c4606970186a1
z9688760bc15237e772244b51d7b8941bd7eb295a76f95ced408ad7a6513621828d6d6627969d3e
z4cc9cca2b93a101046fcd6c5d894d713e38fe84ac9121802d621ddb6cc87cfa8bff9226bc0b4ec
z5778a4ac375a6434593d808f6076bac705fc8cc7ac61e6438e49a743ad8574c7f11205fc65f183
zb2bbf6043e31dd88d142707fec457f2ba173623c552db0e46cd5f70d0380198f179f850c7fcf2e
zc0b22a518b8fe4aea7227d29e06ecd9a14d4730da8f9b4f787aa3e20d4a88f1a5e5ea9d6753124
z5e196bec4ebb0ecd25cd1b486bdfabf31445749e9ef8f64aac725bfb803691c8a9defbb376170c
zcc3b8dba48a57cdb5fc977a0ad709a4667947c62a7071210a6132a28aed36fd458dde8cfbc3b11
z0e7b218c2b83671fb38cdd4465c5f492d515ddca19290200db50de98f712363172ddc99fc2f1b9
z90f52ff5abb4d4f8547034a8113323bf049c3e2c13ee562ed6e7e6bc4e4b91aac5b3bc1f479291
z2e3a3a0c6ce6f27405328f4855c63c8da13bef2317ea5a9a19a5f1aef345fc8925116ca45ece7d
z26a08c7f3124578d12b0c2c10f2ecea6bc0fc44b41952d017fc1e305e7eab0501299b4db6b8929
zf635924f192c6606ac6e5216c8c6fb040dac094216764ce6b2204537f48a4836119e37d0e8a8a5
zfe59a4270ccfa3c27a4f4a7e00336b4ea3e60182177db3a67e6d4189581ab1afa37b65cbb98266
za7355c3620970e0f2132106453c5c527b7ca1dc28be126a85bb83be4461215873634a9d74eca0a
z48b0e7cb889fb37fc8a4a0fe1406056b39daf6542d75c51ee9b41a6841c2abc1b29f435161a587
z3f95a1a877096d97e99e7fc4f505c2d8f192a9ad38f5fc04070f15ea52008028478c137eb03e53
z12893ae765cdfe538d87fdaa6347944451e1b83e4f5787ec637c3abd410036a642156ae1b31c69
z77a545057c4a3aa1893d6871e0aa0aea3fba41cc86424a7c4e5a59466c34f30afc3271b8df5a90
z35a6dc000f56f107cc06a9ef02edd0852fc858fb593378e55775dc8f97f9a4c5937bcbac447c45
zb6dda967fd6501a476d497303e4ecaeb83a973efcd45ed89a30a06bf886388d2e1055b24542241
zf0bb53922299025c4a4e50db65d2966a302d2906e9d6c0cbf3eb00f68065fd3e3d936dab5c2b4b
zf652f7b467f299b45f569e2bc7e1edcb19207bd9060618477e9674388fc07ba87dd04fcd4b48ce
z46c5b6bc1f9c984af8081e9c2da8e2832aa25d3d9413195a7e90f4f107636d1868cd2c65059c06
zc0295988c586d1ba903f3d623f06ef1919eb5a36f03b37e6336259de4f56230f40b5ed423be971
z5ca6b4b18de1b755785e89f4dee17b29b5aa22bce40bb56b33f6334ef19360203e5787386d5855
z111c886a6ccdb3cd516ccc29b082e31701ea6a7397d21ef1606ca4bb3a013f591161a57e61e562
z13794bb90bada8f33623d4f95392f2782f49ff1398a05baa505904e6469b8572f0fcc92afcc3a8
z7394a0f623711c7d3867ae52d73a1ca331af951eb4f376c9705af74411c37a442d2e394c19b34e
z3b76a88755e4b7ec84d5cf4f67120f345bef09ad3b579c8812f40a71d11e32d7511f2a1993363b
z9311b81e46fd883df24ad18001e2b9cd7baf59e874c0f3209e01e29703ce9dc89a57bbf643166f
zb3f61faa834a70d2c41d7082be4995eea436f86833ffba820da239a0bf2e2ce5ae4685584dd9e1
z17801af03036d79c9f7dd2747d10e3f9caddd4c760c7e28e97cd58879e4f9780914e0831a58522
z2e3a11d8a8fa73ee4247443b7ce4dd13471f9c137ea55fa2d894e0465a51c0274b7234d688b9d2
z275feaaf610015dfa01616a2545f73660f5aab2cc721e1c8fb016685ccfd78186f79229027e69e
zef6c21c1deb0fcacc2ead979e0f5c295e786b3813a5472f0db184b91f19578a5ed490b24ac65f0
z64b3571d7bf8f24262f80802c53a12af6bc87b303d987d57ad1581263666cd1a332deb5bb80f31
z45200e0693439e8f3d3eabed2e7b0c534eb0a19b290e77c97429e408bd2bad0a2693b8eddf62bb
z07a4a01d970a057274c6e263010fedd20416c567ba5a2614607c725e3fa4160eec3eeedaa34237
ze53524225194f1ead1345b9a9c0360328592a951453aab8c20b54cfbfacfce28bf2103a7ac0c10
zd989a7a52140569ff5d37d739e8c5db2854d806ffb403170e843edbfa11fdd96508941d84b5a62
za8d8da4fe4ba9d3b5ddb4b6bc3023cee589d18546671b30643eba2fa7e4bf1b51fd0f38fb8f05c
za2e3783d571d8960b43af4af324165faaab0356d402732cdfa5b561ea1dda87a0264c3d0e1cfd0
z629b42b1fe468c4e8c7cef3c7cb3d36d09419bf308ea944ee94179f7f4c0e94f9898fbdeade689
z7e860e118cb9673b695f19e28e623d32865c5f076fd0581388b32936ee5968f3918ce9b4d68ed2
z52ecd25698702e9d7ed8ece1e6c034594f7c6efcd887fc3e26195aac84b893ec81a4967c138f67
z21f37a535bb7c6c22ccaf9f68efda32368e4c0b08be900421616582dfadeffaedebdda57eac5f2
z636a00a6a0bfa61843650aeddc879320b87f28bf141c151db2a1c9e9c2fd72f929cd3948fd4a2d
zdd36903e00721ea5da46dfbcd074ada0f1d04626300d059ec25917a2898cc3a57dbbf4abc2d851
z0eb7917c3477506c558c1c255a73e1fc045e4b76a857052f66b043d0ea4fd6df4424526de54b63
z48f0bf86e388e12b7b3a57f505985d40eb616b75e31378b0931aaf0bbd1d4db84b28033aa32965
z594feb24c29fcf79ae844ed2def66885c5b63635d08bfb0293aa6bfd32f05e3353d5b3aad49c8a
zc8b706ff2f49b86d08141ee96086f0d6ae2da13270120eea6e0e48fec242a0ab2871a996641bbf
zc3f1e008674057c9ebad6b5a6f806d4c54fd3d582c649d7db84bbe070e2d9d58780cd5c6b6b6c5
z7ac39f54908874a6f9405ace20cc18f22632d283d97578a4807a8ec995881dea3ebba28d2d9d33
zbc98b3b4372aaf80f657df3a54a9b4aa7011a39fc65e4512e95e529c6d5c3029a3e1326da0fed8
z4c91ee69bc289783a6ca5dfff789d8ac784c969a03a19a10e278f5a37b654c534041e29f0f20f0
zbd52abc15f049ada6e8256013715a6c89df5d7d16d00202d0d0c1d0fc5f721244d27647db8b23d
zca80609574c228048a6bbf0162ad64445533f06e82263185a9179557c22567130833bd6ed319a4
z898065ad89e1124ee82cef3a8c3f71512e4b5da1972bf7ea12ecd999cd03e885bf13021ea7e300
zb4c16085b497ff4d3d2c192d3cae5d9f7327475a91a75f4f37c322b4353bcfbf755bb0b8674fcb
z0fba17cf971ab1ff7f3243424492a3fe519006bfbec2619af1f48023e19054baee47a363d158ba
ze23e749519632a0dd188b6ff114c8965efc242e70342e931afc396e9d4e01a01ff357fdd00795e
z6b2dc1dcf14f7c09b8462c76346cea18ffa00d1b2ac33b75e8f0679305058a2e10891bdc8e5aa9
z816c8c1f390ed91c893ba26ef7226aa105cfc77a97f3283cafff2ab72d79960afdf90decb18d7d
z880cd9907ba7f8da88e03416eae3e63149cfb04fdf09007d14efd9c50b0b10eb321a2293f1a61a
z3d5fe723e3b6cc4e7cf85eef18b85f301a1d115f7044adf02d1c3cbe717c9689100cab73e64fee
z3667ac6a82d129e7d9a8754117510614f4231a716385f726af81ef138bae8315f5be32b8d429b4
z42e5a8b28b7c9a4fd55834fab8e2e21fa67e3bd7e8808a7e61be01b19b560e3c8b3ce8a4f65a8f
z0df2196d50b05d63c640ecfd06e1aaf1d363d74518eaf674e361fd31cfa1ec57b208bb1e142860
z1243e7bdd27665fd4d80d2b81f6f336a7c9b95ad4a36cd3cf74ff7cc22e7edae2050dfc2f26487
zfc8908b32168ee3ad017a3b2c60df29991a6568277b3b272f55499f30a448e99a2dba87d75d0b3
ze2808dcdb34fb8897a133aed29bbb31dd30d78558588f44dab4859b4c1fe0211d9d664208b8a74
z5cbcd420e7f92812c872bd718a523048ff2b954181678794c1ad7a5e0823c1ec5d803986321014
ze2675cd4dd5a6a4717acbb90dc301cdafbf71f9e0a5bbf05dcf3e0e3e1adf508cde56e82bc2f05
z12386e49fd336e44f8544dafcbab4a3b6122f7d03836383513ad55c70ebe9cd982486ebbd324fc
z3f56d73ceccabe70af5c9c0b53f68f7d0e1767c3944a13b38f57c37ce1e1c5bb2c0e2360af741a
z3f94a7bdb06900660916e493ad15281e6604c69cb00ffed811adbb9c8f9bcb52e95541084d8f51
z6cc469dbb0f7cad5bd0a7d6f3e45baf9802026eb94d39123cc9a3f2501d1a8c2a4e22f33156771
z0897a8a6073fe48f91ab6968726265a418008527da13273376b65b2e979b465cbeb621ee2455ca
z247b3ff30e0e626851ea0075486b6bda194c2ee81d5bae90a6d5428576c044f6330b2d68e52477
zadbd033eb00204fda27192565b4cfdcc8270500be71567d9a3f1bc2db1db0aab2fd008c829ec58
z80b96e8ed045ab94029eb384c4c67c4a680dc2ff48356aae7499c8bdb5bf02025bd66f2bbaa3a0
zfdbce208597fb7b1b2c438c1b3f3248a96be725288ac33977cfa265a91e1726dacd5c10ff045c3
zea5e4a94608b127a5e934353002403deeb1385ce6ba94b6bb0b97587301e9fd113235f24f82483
zfa7b05612ec99876152d4dc0be75cc71de84172a68205ffcafb5945e6e67fafc3ccf160116d5a9
z3a41782febb20087e026c370b9aea48a5e49e2559ae4899ab3380a118ccad608e039d3413a1ec0
z3962eeac4d75b6c551f9ad13df16e21a4978a449c2baff1b6ec40f4cc37a8e43dc0b9d485338b2
ze2747681526cfe8e15d97e5c368e12f6576b341e44d029cace265e46f7b2b2907a5b6af1ebc1b4
zc02fed5baed011e22a741f98f2dbc63c4343a2f59e8299f961e60845270512820d9ec37573cbb3
z70962d37357301eee36e33a0b578239d59f7eba77274e7f04bc771fd5852f78d57ff8a16dd2ecf
z203fc73964fbf6899e40aa66f22bf635a6820b85e2c61927b63cff9234c441e34bd8dce77fb022
zc9b461d7093289a61834c67ac3cc1f6a82c67d05dcc6b6bdaf67989a9752095ad1e41be7a2f1f0
z5b84891bf8d91e5c857369622a2c6aebac89a9a62cd9170e1f3434eadfef202af03a7825570e5d
z8e6214c4bddd373e69f9245bb52986ea1901f0f318d6855ee699bfc96c3c4cd6db895e2dd65db5
z5055d695c7f8f5469b6d8cefe8e2a10bdbc2f6d0015683569846fd8d6420e768b6492adff40ff8
zbaf9aa809af326033081a20388c08d2e8dd2aec1e9c0f5c34370b90d29133758e157b01b2b95b3
z7bd774ca799e40c15e59a2dbcbe76a53111ab1788e374bf98f2f3d1cc5af9f337e0ca013106c38
z23e5526f23c645794aa9fb588b1dafdee2326205a97861a12c5daa48a9aa3fa9493d81dd7f7577
z9d122f5d640267b9a427e3a9e21befd74eade30746d09cb9fd4ad34f44ed54cbf2406aa8e140c9
z2f4ee4f0848dfb144f696a8d0af6e40edcab2ce5e4a82c9cc674ce2fcebce5af868f0eaf6a1746
z6793cee2b29602b8fb43ddf9b68d8c85f95c8de2fe05330de9e4a0ff470ef617c2d21f7119db45
z1b051efe365925575746321b469b7cadddebd4c18d7177bd6c0173288a74b21e0d3a653b594d91
z937d1cfc5cc23fcecdaf1977f97889f00dafe4526316a2e0a23836d9f948411bf15d63cbd7a24f
zebf8d7dbabcc5db66c7bfaf1ccab07440da2b9cd03e4d664e623863daf2580549225e8d1a77f17
z06acd665ff3450073d2ed04605ce4c210f0be16956bd5dfe3156ebc392146414fdcf0b52b12f1b
zc09574b399f1839ebb6edde875b9379e050d18d9bd1169be96282975edf93517bd4a2706c4fb8c
z485f1a4335b1efe24d324f6a3b61b3e1cf4bda32b526d5f4cf475e0ef1f50efc927f56c1433bc8
zead64b7d7e50d85597b9e45380cbc4209ea9b4b540bff298f7bffa68459c234b8ef31d6072e1d5
z308048407e8b5e3613c48a89b2a79c8298d4ee16c496d80a1692d6f0b6572be9203345cb0794b1
z7241bcd617a8a4aaa860e47d182fdf04831b563064a3a332d463042f60dd30a960c54f3939291e
zad40df49b58a13fe3fcf34380d34d8433806c58bd0772f5267d2b8ad86a17ecb09611046bc75a5
zcf68f1b7fb843bb12021335f5ab2d6c084e1aed15e4347f3578a5ff99869deaeba8706ccaade9f
z1364365f3c44827faf5191fcfe1a3245c080640b147238c5cdd75a056333d399253c2f7cfe0294
zd5f214562a93200167c66e51af14ca2eaecf8995e143c2908baebb0005864a923069f165fd59cc
zfa066fc2608886073180c22b21ddfdd504518ca6c80bdb044f073efb90ef4638fe8bbe22bbe9a9
z782324b774f993be14b09c74dc5b6055b4e59276bfeb909f035fc90d55d7caeccf9a4bc28ae944
z209f9d58a1c7e42edec6d61fb4f3e260ab0e9864d1d662e46056722cc2c075329098ac1b6219bf
z0403cfb7f61c1baba6839fb583d3625fad3030e62ae230613f5e69bdf733e17d03f7a7c261799e
z9bdaab096e4b396fc977b52e811e666ab887ca79dab2880ae7eb8da3168585bcbc078723500be1
zfcc3da1f2b7ddd31a436368c8820962619151ee7a337521db99f844af2fdc21fed9143bd5d09f5
z9c5115465d9d65ff4c421c6515ad354b3dd3e77d79209ca946404a162f8506442592cd4c24110f
z8609f03b456999729bb77a57001f296c1ab3d4ba0e3b259621917179a82726d756948f83ce11d4
z7e15c30b79e385246201938fedf9ab9369decafd20cada52f3f1035e72ec7103e9b7fcb49fdd8f
z0610053d6408aa0f1ce1f06e788d55bbbb5e8c6703ac6337b229cbeb3c74e76e8c47aab97ccb8d
z2d73ab777450a5c88954356cf0b4e6b997a88e76bd14f05090d017ecd322e86291e87698fe2388
z27dc62796a0b200db00d9df3e38cf9896a4aed079f15764a5ea333df6a2bda77457b41a25dd80c
z67aa62461c5e6fca22eaa1e8bc3133e103569a72df8ad5e86fc38f5db44598154b215eb841ba6e
zcb4678e4d86e5d6a400b5c4b1d31d446bef2ccc9bcb3f44414ff74608aa98666c4f6e62a625859
z31c49405ea7d62f3a4fcf83bd73f41ebaeb41c79ad02ef192fd99bff6791c0a6de68d9d40dbf97
z3bdfd823d60ba1fdfb2d842c025967673ece9896de7347bb9fc191f2fbb5d300ac84e30b2043bc
z3c84a7887a4129b84aad714fd1c6abf209e6faa0ed5f99df90deba9bb7286f9766fd3244472911
z4056413d355ab166439f1a75336bd5fb8c95020d6721fd30003b1c2e2736cb8299b3b69715368d
z3f76f6c3b08200ec9ca8691f805e6e65debe9d631597264b09ee55fb8c0eed1b29928c4b448c77
zd9fc19b31af8c4b26182bf5e6da8d8b687c42f5585ea1fbc6ec25f4fbd63af7aa18b85f3424b59
zfeda0aedd3057552c7c3eb72294ccc0c0fa8a55c45070b3e3f837ea90c4c6cb95ae55f7b0ef617
za1505dc93244bd548f59e59b9bef631b92d0ba011afa74cc2f33b87c74e86436715af4aa18b3ae
za8e5ed61037b49d2ece99206d292a14fce73d27f6209f60e25bdc2e54d2730a6df092ff376b8b8
z2a3c2dfa91983cbd7db5ab4baac252ed09fef7cd57cec456c6be9a5e96d46c46ba246e0a56ca52
z5ae8b3723cb313a2fa84650d4d00e52f0d9b97bff7eeee5cea8d6de69ca4506d06359bedede088
z43ef9c8ff329ecb6ada5e721a6f39ff6b6d60c0e435959eb0113225b75ba2061ba64165ca4521d
z4252ed08a4737c399bb3fd1dd4437b5a389a91ce31fa694907cda92ef8317406e18eb9d5f509d9
zca4a7539447ffece3efcbbd539001ea10e751b2bd3e4faff3cff094540830a0ab4da1a700d7602
z2f83a5070567305a91a1888539b41d59f217dc0b514b5198a65c169c904f9d37448afc83fe37f5
z77258d437d3390e54229a496488787005d85eeee4c21523e4cee6fbdb57ec54ab1346910991ac0
z66a3543a4387db8d1898dee67be01e26d8004cfb30d875f8816be5ee6bf2fd0416cf8e22074af6
z18ea0122b43b7c2787cb1b58648c0837ffee986af97cbfe4e84838122955cab2c0c4575198530f
zdfc86e197b5ba4c12344a8692d28449bea2de05332fea351b1de7a2235f841d1522f96c60b779c
zac600c4f94ad2bcc1346623770e6cc4e6ea064fb4c81eb1b12a77ac52ec44e72e54cb6cdab47d9
z0366cb85d468d2d75c7563e97951e85a0df9d3205c0240410353711689d487a62ce00b10efb763
z655e6218d0a377b6110f61d2732ade04f8638a102483b3ab81a51fa65b0a6a4f2bdae02305bc40
zfb9223ff605a08d2204f2f779f2c119f8368ea1be8fb111de64c719f0512aae3cf12a0bfb51097
zf92333ac8acd81de88c39bdc8ecf9150deecfaee9038f4d827bd652e9246c5d52b60f3c8d8ca68
zc1aa626497a97d2889701f0eb8141f7279ee0051be2bbf87c86ccc76de867ae210b3dd441a4edc
z4e04486d92f94da4ccb2631bc39cd0fea32e3f67ac961460e1abec85f8bfafd31dcad4e4f67e31
z181e2b5a2a9625e098d118484f0c3a54d9969f1d315cf3aacf6356fc54c90182c70291e632b149
z2776b220831e79c014dfb16d9017960e83643d921e2198935cb424f45cb521589e9392b2bdf6a5
z10dd0c1930b9c3668b65325a0f810737ebb343d5b7cb80f184f8847a71f1ca16567621e0e9ffcf
z699931945a1e1a16d052d3de4e018899931e078128561eb3e16138f055661d2d19866d3c5451a3
z1372d35537185b49bbcd615aa9134df150a1cd496c45c8296ef0c3e7000edb2841d28ca56c6870
zd6bc32a224483f0cc3fed195a2bc869a15e2a560f35bcf459667ad45b0502fbd28bd0047ce54c7
zbdf28c89ccdf1c4879af2ea78c38dea7963a6c0c34fac31ca3dc3c29f124729882715a64ae0871
ze7b6102027145115a9c7097da0c133c023519fedc6d7a6e5d01651b2ab09f3425ee55a3c3f88c8
zaa89fb1b81271d28b86a903d5f0391dd4ad742951e959de1947600f92bc4893e1e9fcdea1a8461
z867188aaad60ac5faf60aac3da43e6b68f7c11a3833d2346dd1c21361bc8db86f883524657ad8c
z4883479282da6a565a93f9675ead1376b22bf903cbc3e7a39391afe6801a722da83829e1b5466f
z79a210e84630adf57aeb96acd0fc0ac31289341c5c508702f302b1b328bb0b909992081a8d0554
z4ed5a8ad9bb24c5b50d69db8a06804a21938ba942539b9f5f134b9fe8f27aa5dc5a1f996b182c2
zfa82c4a4ccd13ea3a4095a7a95f7dc6a63f0b900bc0a0572d6a57ea6734bbd4a56453a4aa4b722
z0dcc835a8e14c24d24330500851a9d31aa1fc95e3f5802e9dc9b639a76e6c7de4d9e04aa96b7a8
z76a2e40680c0e2c9686e02f42e0fc05f3117f115692603f27402a57003aed6712fb74c8e76390c
z362b4d68db87e9c83ebf125315c5d3ccfee9b4eb4ff1f3d8de22a2af761d949e81dbe2e0cf53df
z0ed4a3a1af396f72fcdb1013d87528e536845d257e3d18adbf9b6869b3ddf4bcfa964c2c011eb9
zf27a1ad02168ce04874867d30fb4300fc372767bca62752c87b274a8f1fce8256a776d493e23d4
z1c7addb2431c968ea91f65051a443dda9496702439f18f38b448c1e8ae905fef05fa2014751d8b
zaf041c7fc5279e0ce44bd40e6b6793169fd926716efb882c757f2703a07e57ae95ff2768081f25
z72e2c0b05545cc3b541687128e457effc8601cb43f82e6e64b8ceb5b18c16cf534dd6252b430b0
zc2f39fc02948e6c6c14318e681093311583b9f0caf2ed95aa85f5665e1633a02faecfaf837daf5
z5dd04e23c896900aa3ededd6f311c538dbae88862a7861a862567a48b0ad04e4aa55864a9bb201
za91c5824c532fd2f2c1619bf80dee992b62de04505a843bb8134b9cb26d86ab09916a5cd93a2b8
z4a7f1513bddff5eef6d086b09d5b4e9a9b69c1886480ebda12fff60a05bb8c69ed2204a67218ee
z50f06c3ee4590de9dd041775d0bd743a0dd60be35f862107d3b19d2e73313cd4fdd042150ed896
z8df7db1ccdfe5a8d0d7c9e88cce49d0b87e809084aba49dab0619138c47d66ab8c7e0610e678d9
z4d2bb7fd5a5c3f3b4e4b7533c455fa4acf79adae823b14eaefd11220ecf819dfab09cfd93ceed9
z1e52ed735d75b7dc70bbf5a0ab42824eb56dd40c26ee91800b7ee685dd8dcd8a0fa7a5a43fd01f
z33a551a8fb46383723ebdc401bb3a3ad438daf9c52341d1d1bf5634b922c1441a91e312ff59849
z21027ee5389b803460664a56e99bcf5f2fe2cdd48ec6f0c40e36b2f0da950c92484f18b74cafbe
z8263aaca4c0bd17713a917a9c0624f0499db6418253e9b834705074c10e1fef37f0cd47d744a86
zb1f3b465806a9157f998a9611069461418644a9ac0848650d2f6385c0563418d4ee40a929fa06b
z82ea132ddac4835d554a6dc82f9bf46b11176f5ac5e695c0c3fe23ccf6d54a3af74c1cb331d5a8
z310f34daab389c9b8cd401e03539b6625c438dcb5d1e41c15b1b5d70e15b9635771b17c4e1d7b2
z2d041dafbc082aaa3e37db17c808dd35d165d68f691c621f7c185b52efe040c1fc6ae9e4617f2d
z329544cedb897217d2084781ccf1b15dc8783c12db3e1be9be6b235f0109b571a214a49e42cf8d
z10fabf40d7327a01b77dd2a878a21beb0d371989a8c564f56ecf81eb15ecef706a013f1161e083
z03194f681bdb5b264e72f5f5ae38515a5aea190e90caf4af8c23d4f6c94c2d520ddd16cce3b791
z4d2b5c8bdea8a271eda6470940b3bf00e97ad687b033a6f5f85a9ea5a5130967c4e866a680a113
zb9f60d1436752c93e069881445fc550e6147630545de03800cd695c349f7086de299beec1e36f7
z3cf87c30cf3bfa367fbd61f61e36233880b63474e43c1250708c11300d9a11408b7b47a8cf492e
ze3cfddc4860709ac18f053d093c6f5967887e623fb0b82a090ada7afd0a1b0d3ab36ac38dd6abf
z7564e241bbd96fd44b7b1c60c3553af8925109c1c316b4e5c8eb7e57c5097aea821e6af8e52879
z7b3300420da93dd37e1c7bb237fc4f26fc57057abdcda82080b07be0a97a19a32f9a0177e0f77e
z63be8e90a088410c6561c0dca5aadf2a1224894d09695822a8a5d1a2f92dc3afc1e51263dfa3d2
za216c38a707d06ef3d714a7912b84c1bde610e8ef4dbe33ff79dd2920db4ac0aa5131ba44a2021
zcd92972dcdb33f8a4f8cb6d945d357808d54e449f9863d208789080cd0e4f86c5a425cf21824de
z076a03d97a9736b4ded4c5cc6095ed0764327f22798b32ebfece7feb3f87028e69797217583c68
z86e04bffcb42d3e868c9213c8ef92160ab1104e01424aa9240679d2d2d863b10b83007dc9bf9bd
zd94c6f8668ac86a11384a6c9a494bc1d1aada1f7f470fe652856bd271bafe0fa28450c3fba4f5f
z9f2b2531b5a7f1bde9e8d2dd4d8c5ebccb6db3dba74aa93659a6c62bd214b6027e93b929f7d5ee
z5824b2560863350d49f19c6d0f539bba39cfe5fc43f674f340177abf7ced3b2e0934453a4561c3
zfbf8e0050e2b570d74a9d75b74d2ddb3953e2f52e4a69b7d60f668e880f8f1611a812716e85605
z3539f0ed07558f26b03144f4ed08231cc3775340e954fe06ad1b9030183d2011fad5469b119eec
z936583ff83ae1075410f3dd1b6c5b5d97bc5ab89d3a6dcc9fc0c9f86e0e3bfe414832fa19457eb
zc6aa3fea1bd47400cd30de37aaa290c7a2ec5e9c670652a8abc6a06248bb75c5bd33eeed25472b
ze224beb1a35e20907adadd4f3d00906ab326e9088a0ce2caca1e00b658d5aa34496b2c4a914335
z5d51e00c2c57d3ac1098ad1e00372e4f4aaa8bb5584a2556cec0e3fadf5cfac027b4d36d455c1a
z641d9ef193b96e4ef9d92f8a57184f687e1123ad60acfa7bf9195ba46e1308f9fceb8b8d79e378
zc23963d976d46a2d4ab3e133d4676f2e19f5e3382e0881fbdf865edff378791f6dc1b741bcc62c
z3c1f01301664e68accbfdfc306dedab2b48ef7f51790cb4dfce6e5eb31a2a206c6aed24a3289e6
z0141fea38e3a46b1435d25fb5e29f865c6cce271f9961ce4f5ee88d4d7b25ca53e7357af600d9d
z2d6dde300cf29e2de8aa2c66c5300b9d272307a44c5163ea0c8d20c2db466fc894c4f4be86670e
z4c9dcd06c1e54076c3b88ae8d70727800d06839b97b8afea012cb8e1e68e51fa62381714819427
z3694478418e95a07d17f4f37a4b527e8a850dc7e2dd18099bba4bc5fe8f0e31586ec3b93379aa0
z668a6109f7444a0a3202f90e9107248920686b77f37e4e067aa0c57c7cb9625b8c04bd97f8257b
z2bb67a57d7d3349b8b72154a1b44f68728a8a4e8d95b28346fecfa1be84d84c14e217dcb0666da
zfbe504f9574d2952010c120686f913bd2a888828900d14d1fd0044d976b988e09606db4442ae8e
z1068efdf0f4ab06280982d98c37b638edcaff1cb66852962caed3bb2a81d0cb97fc66e0854ebba
z1b3a03360afd75cd1464ccf89a76b63190ca0ce81d2cef0f9bdefadf28850ffd7ec3e5eb397f81
z3d12b662e8b5e8a0c056b7f431cb71a9e7811643aada3e634a9a3a8dd461135c6e8265b304b7a2
z337e1b85df6d604735b9f90b619f8e89a8241a206cd363b784434294e29594e2ce95c68a48d27d
z10471323634eb25bc0efe9fcf430d2d91fc7df6e61601af8cd34c50121ba3ceeaf2c85806ac8a3
z1645a8789a1a87d2cbaf38736d783184379f1bb919144a937ed247dea6027a2e5c99b503d23c55
zcf08088e59e9411cb5f01a4439a03cb656d6f39c27415ec8daa975dde8d40281580fa6f8382df8
zde19cc45a95acbf89953f0a475327a44dc545d83d1bc9559765e70b612abea5116ffe94204c575
zacefd0a6944fe702711d8a003a77e4d3bc6d65ecf6ace27d929ace8e157e7c6c87987fe1a1b9f4
z3bf299e10aa2c50fc5f27f711ae179a749680d40447ed9d1cdf8e0bf56f5dbb966ed514bd9e4ce
zc7b009559353bd664103e7ec81be7c5f76958998fd96dfb134c162c37e544ef4f11c6d0b8aaa59
zd87df6668a64119d794f9ae2996bba8cb9af2ba707ebdb9a2dbfa546a16280452d4030a54a17d3
z84aa16ee5541dad49eacdb332931db1e482fe8ab9f1d0e89bf937cbbadd615b5c063aca6546944
z4f499cb1c1f1626b75a186af2b9d0a2a75ceba95f98a79320c4c4d7fa3f4f8c8ab08829c635538
zcec1d0d1cfa72bafa78e2e24dcd3efdc3f524d62da7653c1704a3dcca775a1cde8940a09076502
z2055c71058102935b74d3768260ca1f40aae0bb6d1588e0322fba2f55762676e2821ed247bb920
z63f12712b06658e1fe0f2f83bd400804a4eb303922823f4d6fba4f0a322bb783da2e73bf6abb7d
ze7233edd762b591164800784873ba47bb42fbaf82e6735f4ef7241f08b3a126b853f0850f77f31
zddbb6331373e68fcb694073619a66211deaf22bcd500bad9d4dfd998d205ab946354c4a114221e
zda396aa386de74062057420736318ee3beebc44a8f81efb61e81120f813fbf5e5bdf95d83fefc4
z63b98d29b348998daa34bd8447158114568577504b82f8db6b322d3da9ba00826149f25b7a879b
zbc77ccfb0f53f8777d8ca0249620fd1077d91c18ccb660e74e62cee7e2bd7f0269e814e858c6bb
z6b16ac5c86204a618ccd554b919b26c8bdc14783483cf9969690d6f086a670058eb57a350c7953
z505f55dd4098574b81ce1fc8b94d10dbeb08b8450313aa9e32e5f858b99c313f1cf792b480a6cd
z0f21ce275b41eba5c6cc5e7fde5485f8d9ce01a717e0a60521a35873cafd96f180a8849a15ceba
za1cf1073e3c9192235f9a14b787921c40b23e9d83d8be91802cc56b2080fb66dc97eb799f5a814
z1b2b39e054caf158a69314e60bc1d18610c3930b6599ae532ca97e4b045b194875f7e70bfa29f5
z9ae47df6b873b0ce3d0dffe84ec64bbf6b501350b0cc78c6f9fd338f446ec58e4eff84ebee700e
z898ce9f4ed14b63904fa4f5b42527ce14e0c9fd98ed556f595378c16bdc615e4bcaabf2b82eafe
z6ddc9d6def183aae231a43b9ce247bc3f5714c6f8088bf23dc5bbb6a9e0f1ebaf887dfa98deb2c
zf31f1ef6af20a5d8f7f8191dcaf923caf0d6fc82c90bc6a0f93a7d06a960b71118611294c83219
zb43a04412a831123ef704effcd1bfa7b1a65643e1f4bbe6ef68b5cfc03a9cfafaed37ca67bf457
z8c14b8fb21c0af1a0b8343368af49dae3104e91a3339e8c9405b1c3c4a0efa04dc48ae5fedfe34
z0071750e6e2c4303bcb6a539ef70894b9cc9aba9e99b076405971c22f4c9f61d6cb778d3c07f75
z0d3c2296b2cb7b41dbd04ac62f4ef112fe816729fecb1749e5cdb18522685ca1420db50100909a
z1d72637056afb83ca46788e9317972e79f43a184ddfba6c2b0d634f9db772de3af80eb671f81df
z0ea07857f99ffa1b6c7ca09246318830c9a836739d83e93065385d60e949e7d37bd3f5ae1633e3
z4e457882ef9947859afb6f3e2ccd23f541b32083fdbb55a5959b8b8c656400c510449abb0e1914
z64c4fbea4900d16918344d0936ff65daf38574adcd47d1b6d6cef5fe4ff3f9e83ef4d9090c1be8
z01b645e711c60ebf6703fc9e53f06ab1b50c3669973db36caa460ec712166cffa90a304289ab48
z963d9db20181e24dc8ef90d8d786e11ec6b3935147c01cd161831a20c971574f5dd9d9196767d4
z2f0ce725e3e018555eaf9b98784f906ae02ad83f4adcac91243c7be9757c6c4ea70126266a32f1
z5b594c2f96bb901670386fd243c315e61d74adca3cbf3db445297ab08121697757aa5beaa288cc
z9d8ea8025ca32a54c8ea78cb9844153ae0750941b5d65db37300f2cdb5e6f115dff7e863d7a672
z40ae15dbf6826abdeaeb07fad7b778cd285968fd530942b30d3d49544669e536e3222465157be8
z84a0328bc1e32349038ee218fca7477699d35ed76c1849c7fafba04f9507c7338fc0cd884ac0b3
za57609acd131c5cf0e99f6094708fa236e196d0fc7af976dd85140018d8fdef3a3fa29db869d04
z4f429e2ffbdb10208c8fcdcfde25d60fc32153cf0589710d3a46562d23a9ae8cee8c827945961c
za5566eabf32ae68158752aabd19241c6a38dd92c5b48035274ad598ee3f973c355e40c3d9c1bc5
z0b3e8646fc37f2dd251b6ce19325fa29debf0b3aa362d6d4e3e17279f6921847f176bb1a6770e3
z37bbe77a1f8873fa085218d19ce53a3b6d52bce16eda67029d938f0731acd3975a434af13b94f0
ze87b5cdf438bc0ee4ebcc472e849123d82220263c3c9f179ad3c660872beffffd977ada8f5347c
z6afe00bb8fc55245f9391647973de72140e4b135c761ee23ecb1981a6f647843bf8acc2fb5653b
z7dbb54d66fd94fe600ec63310562657efbf4e3d7a310e8cf26323c309be4e702401339e509f17c
zfd7b09015919d09e7c465f7a2cee256c83b20b86d3273511d3544733869c903cc31edf80830574
z324fa1a115d42e18e66a0a11cdd1459540b9443998658f43da741cde984ad874b14a70fddbcff7
zf42ef6eb2e58eb78ca111199fa8fb6d0e2d9a4cec8d57523ee0d1a9404ce9b410d6ead27a74525
z380f859677d1349d5af12cbca38ec3d8402e98fdf69738f473fcdbccba18804a91f0b13bef4d6a
zae4e485de8df7e18eab49450cadaacfe2e44e740d5eb10296491d0f1189582582992f1d69d8cac
z4d61ba93df4126555b5fbd3acca671de40651a162bc6000a62134373ec1919753ff5f6b5464246
z60b269e5a7b65a0da50cb6258c0b689d49a38b999a8a8ce3b14aa8d2e0ab90e8803b06bf409c51
z5961894e36a5f62883886a12161a7f0beca5dcf1d79a855f0ad6bcadfd393049161f7a2ccf8dc0
zb0cbfdad522ed36bb8d2c1dddcc157c9d0a2cf04469c01cac9b637bff7e02eabd1e19904c555bc
z0a8f0832b73afdadd1eb8e5afd427e435475f3ac6949ade93aa0b9e5fc231a742c66e04bb9cd41
z4534e65e51507cc95d6adef55f315534200e90c1e50c0d25193e1fd646d524f6038b09fac9d49f
za18f307ff5fb79d849a24b2ebe73ab368ab09ce64deaaa3e80b107a33fbcd9664655b2fd9e47b0
z0c52ea5bfe861501dfa6c6c075ea4342a1fe3cb3354c70d5cfc08b7246d11f2c9b14b0cb1d1c02
z5a75d641f173e81e426ca9c0e2e697aac94422f5c0c8bed13673e470f048ee294ea936998f655f
zd68fdf8bac4e7cd9aefe35a5f7d91e4037358639062db3ea5057e42f74ab0c7505c144a1704515
zb4092e93061de4d02b48622315e55772ffdc1c444b1b8daa1fa789a900194685482c67da64390f
z20dbbe0c6cf711a19a552e3bb605c5ae8994eb4d236c55210fe85f86a98c1d85e213524ed2d4bf
z6d8b2ee9afd75b18b49709a5d4d3711ff2ca4944d3cdc46fa49831742ede41399d735f55897cbf
zcb94bedf16bf989e592803f35a6558974299d97bcb2a340c9b66d06f4d1f765a479e8e8b7187fe
zb346851f1825c7e7c8bd84838565d5cd4bdb7e8d4e84d975c1c2f0097ca3daf4dcf440c65e39f9
zb0fe6ef48afa72fa03eb66a97a95825a07ee25be7746bf7a924efcee6c7749d723ae91b3ec0e13
z686819b9368cd5cb5778f09d916ccff6e11786be35e4a4ad6d15b48014a53cddbda7b51ab25d36
z5f526a20a7bce066ef5757336987380420d47f7ddc3c0011406dc0563356bbc2635780dd1909fb
z141c48ec0b915e61469a054e6f339422025bd1f2f6740a26bd3c7aabc5041bff0401ed17144528
z0f417b139c3e22c3b3ea69ab973f9f5e2064765cd4451477e66e82b9b91af3e4c88290b432f742
z0f9677b9f994405f2a1d5f123f277e07b1042c65c0bbf0fc02846d8d2d61a7dc103914754f9f63
zb02e0f8bccca70e5fba9f0931e80ffec24addcbd16738acefad8e4dc289e9136bbfdb5e72ddd0f
z71178c08b95332cc4d89b70a74dec2d030092d4a4ad89f0ac6aeb7936d77c35364d4d48c3dedf7
z702899504d9adb20c257ad41e7236655c9dee1ea9019698617a3a2013df356c74eabf7bd21cda5
z3b10845101ca6f97ea5b23b044fff14818f4773baae67fc92d52e115df58d8a6904d5db946ac47
z00d495b2d7c0de5c92fd0da25347ff8c24659a4dd3fc6940477fc01a7713adf79161471339fbb0
z41d559ce49557132c0ece05c7ceb60e96e3e8c4056bdb5ed17cab5cd4134935088fbea933b6cd9
za92a48d67eecdd9792e18c2d0cfef748c75b24b3746a6adfaea55171273b726a1c2acf1a8f2e79
z9a715c45b54d39e6bd4b0ecb2fceebe8783e23cc558bd2d4be69e6cb5420ce85dadfcc255f3692
zb3c67102d0ffee043b76782401620ed2e3724de714224789ccdc982ace10e44e1f9d4a0eaa4fa1
z486251ea2ae6d0620f824005a1d23c8e846f71c2b5f4a376a0bcf8ac34b3249bff07b858cf83cd
z5b76e133c14cda95a098223e25e19bc2f288547b9e739aa297e32efec372dd16cebc8ecd724f5e
z9012d97deee54cbf43aab4fd88d95dea7db12c370f54b9a36abb53fc3b77822183d6adcccc623d
zf77d92b835391913af7798d758c9b35a3ed7494869fb871200d853d30401ac36f8fef4280155f3
z56adfa7f0effa796b75543f5bd6b3d60f6e4621b0886bba575447e74e4a315e709dc511de2a496
z12d801ff0f31b4eccc808a6730dde4d6ea57f07c6aeebaf2efcea8ed1a39fed65c07e069de8adc
za6b64f5847482464740e8fa0ae79b5a28551d72343aa44223ce62ae12f48af95ae6f4ea65827b7
z1e051ed15353b32afccae08e56b5a9a1fe1f3ace7ae0346e7da3ccdf3732d2b59805a98846c726
zffd6047852c550ddaea2191ebcd08aedeef9f5553de927de234fcf4e2fe562ef66252f2bd1e256
z005151fc90afd206cebb8edfff54d701383fb9a78af65db975eb930659c7c8930eb421e71baba1
z3f0c303c7c2993945a761b6b5be2de01508c330fe5ef7ee998de29b6ac915e041e7da83ec7b588
zb630850d4f4ffb2228ba1041aeaf5c84ba236178f10ec29d72178bf4f771f82e1eb0a96a98e197
zb1c1f97e5ad5707ef93f846206e837e383a10eeba726a0b96aba26300843627d522a1beca52ddc
zc92a187de5be4af95e99961ec1dcd8c88793478b38456e71dbe37eae6dfe60cda2d09b1669ad08
zb71289d9b3a80296b296cf346da2e524c35a18f1344dc6e708e34ab6794849f010e9b97be47ba2
zca866d19c2a7f203eb39c592bcf83fd3bf578affe057ddf6c1f8cf650900ab8b5184b1ec78cd00
z6ab155e6f718691d52230f7b6695c629b1728be327f6fa97c70379f8d30f3a194f01ef72b0a6e8
z0a756bf75482a5f4e9a6b9890381a7ccbeb4f4c6d2bcff5dd2b1c6f7875e5c7bb65df0612369ab
z8bd2a564ffeb34fae1c78c95e71816cc5dc0b0c21c3d28d001cadee9f53ac3f5d9702b22916516
z6254b4fe9863960a27c4fd21196836d9d4d7673df3ab919503d1b37f3c467b0e7ad409320f00c0
z765a1bfc30b750dd7646a58e123304e93ccd1fb69af1568e86ebc7288706300e445b0cb88a2939
z3b97b9397aaa4afd293f4d7cd1158f1cc501024f7ba5cc7d4613663065e36d4d055eb1666d2610
zcc5653f5219067d49aff860b14b3378ba10bb870e8e235fe6fe419de7fdc95d5f18c7555a537bb
zb96d957f6c8219533372d6b2c126969f61fd8eebdee0defdd7352529c904c9dc8ded64fc1dc6fb
z8a7036ec0a793b78b4ce3058d1fe972542c53bd25cb893b116434db716a55060c0c99bbc311531
zfbaed347340fd6c010ab02a65478655a1128dc36782267868624a164df612a9dee3b81fc50b18b
z0d7f0bd7a67669def1ed40a39e856359a32fddfdc619e63bf50e11160a13519885cfc60cf86bbf
z20426e87084ae0da37bca1b0e6b274d8514b881f3586ceff1c45d9b6e311829cfd3327ea1c9707
z828ca276ba281654c41a0d6bba5e961a3adee9460fd2ba3a040eed5b6f92eb979b5c6e176efd8e
z872c592a0e30bb568d1fe273626d4c3bbadc3b46586a287cac048728c8be035548bace3111cb23
z5404c37ec0a513ca36f6a78aae5d9b382d6ca59450b712795fb4e1af5ef64c492cbcbfb186b799
zc069a25aa9c788cdc81997fcb29f0e78ced77c06c9c5147fe071cebad2f71571cf77016f12bfd3
z4b80bbce3cbdd2c9a10834c9751331fce1e8a7fa61deb8a7dec8cd7ef6f59f02a581a90f034cc9
zbb8397ddf8e93bde9f2a043ca68285bb2832e6f6c46c93267ccd5eae188e21c733786a9e07a9bd
zbb0c035b8d510fdc76df263871cb4a94055007a0d0aff90e19eebbe86029eb9254bb1be6860879
z377c08323ed76e9f657c78faffd76fa85e05ff438c95b4c426a9a7a967ad490017ed196543a6bd
z7794168365b8dbd22238eaf46032fc4fbc4f9807c3e7be3d1294d1286821af1a5157212596d9cb
z3f517b8870e81e5fac01d8776cd7fa9c6b397f03187bf474ff52b4da46593bb76647d0775e2397
zbc906ec61f4f8561d7e47c9aace913c9984dfade741359216e65ee46bb2539d5de924d0527ad14
z1dfea181a2e63c0717b4781483115242e0d04eb396475ef74ffce14186eee3e7ebe9ec75d70e81
z392acefa32a8c6fb0fedfff8cae34408f138eae94752033a7dcd8134fd97bf0f9da8e3ebda4569
z549e6fc6853595c0c72497121eda6fbbdd839891a2736f78841bae439448d5499822d984855d18
z4510d2003c1d7efa67db3f47b534b6367a3bc471e0eb123bb9bb03884d86992f5c80978f5ccd35
z814aaa92045ef7de2ebf83d890d8b81296539a4919a4c3d82e90c6331410e9622d741172437c27
zcdedbfdcd857fb90b6a077ebd1cc98da241816b8feba4e2ba421ca0db95d94354a1866b6c6bee5
z48d72446395d9d3b7b0db53f32a504c0ea0a405bd860ffafacb2ddf5221711656472994e8dcf50
zba1cb7e8afb19b99025b68b6e93b3ff7128fc613e5f0692d19aa75a70f2c2cb98f4c636a28ffa8
z7c9a729ac21be2559c5730dbec34ce2d1a4a2453b036051ab934c76b9270bf50f76eaf2f0a8599
zc7cff6ec3bd0bd3974074e1c2dbaf816fba223eb06f2804cf9646223ed4041f7162a69f3953a9a
z3c0d0c93d8d620ec85c5697b71f7d057f74c630e2da07ffc6ec9bdcf2388a199697545576326cc
zc687950bee6986c6cce4af8e04498e4f437abced0bc7c6aba72d3c073b2bfdc0d141895280c6b1
zbaac8c6181c9403e5273187b22665acafa7eb150c5b4a1780f90a7b435654faafb1c24ad3630d7
z0275111a7dae90647222274ce91b98af8f5d7451953dd07d100cf8650fa38e4f52166067252765
ze84e274b21753a252e4cdc159982e10cf117828bc86742c35c78fb87e0185640eeb1d4f6f8f2f1
z54463211e7718be8e75f2ddfbdd05c136a8a67ac4fa47e9cb5888123e6432b73ea5a65ac2fefe9
z285bfe0511d1eb985e26c10d4d6cb235d3ab58838352a8eb20047fc647f75677145cfa7ff14873
z0a81704a49bcdcc6ef30253f924add295feae289714a7e51f548320f64ef84519efe69f3e14cee
z52caba871aa572c7f9651ee3257639aa2b0c37d7d73c22477972b63903b1ae8269075fa5fbd66a
z01be6414574b62267fc75c7eeb9b92d56af36991dbd94b57e666b4b2409fba6e81d230fde50fcf
zb3960b7ad412e6476aed63ccf35c7044b9ba385da3a91a4b7796c98c8161927d24eec0cdd2689a
z2f0120b51c0c99e36390e19eedf1d8a599617d9a30b6bde00d60a45eedecb02cfc6383b9f5e1f1
z3f1cc4814318e52bd71fb2b1178ece5d0b05ff9602180427c80b1effbdd2e936fe7c3faf81ad18
zf95a5e340a0ea8b7a93eeb6396226fa68458d1a3b954e68674acdaa57bdb406297fe7a589b99a5
z894e70a6d7ce76535c65c83c7fafae47ba6186ecfddaf7c303dc904f50b203fa942566fe38dc44
zf0afbc21cdb9dc8c47f81de2ffeafa8ed73621de6d4e3acc32b11c77afff62f99a3ee752755b92
ze8e0f7264c1b238542054bfdf4913cc7820c2099d99d29eff0938a494189e78cf1e89f76f6c8b2
z6ec5b39f3fb6a995917f43097bad1fc21880a03f49bc65b5d4021355c02cc7f2e1f1676baf6bf6
z50454867bdaa0298d5d65172bc84007889704b1e3995ba8ec5e4484cd5b8962c584d6e868d57af
z724b8b1f0a9252a080b4e6a68ad2f818ee33ae91b4d8cb219513e0b36c0dc5783799cdc2203bf1
z1f757bd506370ad60f9eac482989c4ae2f6221753b8da04a1ff84cd7aae00e62cc18b6a0db3859
zccce943b4374cf010797ce8cbc7782ae0fe681b2b120e301cf2d093476bdfad4a1d26a605ecac0
z46df549d7c537a0a0cbeff2875cbc3ee92050b5de62e97611d658e3f3692e7d2d61fba5204a185
z068c923097da23141649615b57ee575bf65034fc3a36dd3599137005f52ea13fd2b226a5a21a5e
z3aa113337db90be06521c2d2849bce22e66cde2ad4b9d15f57f6d5568cedc603e3449dba89f4c1
z394cae16ad6846469c34d37547f2d5e9a5f418e3f1303d4d260dab37f48544e5dad5086d7b25ab
z675dc3ce863def5a7ed02e9b60100e13498b494dab7467bae7698799bd9d023623902eea83115a
z8b7ee07fdaca7253124474e2c71ed77116ad2e7c3a1c66116d01dd4d4d9d48f7c7b9fa4d77deb6
zc5b3ef1a75fd58632c9276e62aaab5e65e5c0b5b42dac98d6e24e3f51440837cbdbf74488af06f
z51f7be5fd514aa58f9e1940598b076580cc4b732a25aeb70e8a9cf3e0f6042bd5417a3966dbc60
za0de17745dc7fee35caffc09e766bbca852eb49a8393264621fb4c469ba05188af5762e3afd095
zdb9028a15cd79878e5d779adfb43afd72deeec13b1a881dd64d1a9023820d8bf50cdb35e411ab0
z11a5c8b19b3b6cf6e1cb6f6055d453098381265f3aa1835e83bfc022675dad4858da46cc8dc6e7
z112925b2ea24b729f0f9cb2b7a5113a5cd2f64bd25e7527f35c2a4ed27afbc95593868100fdde8
z9256fdfe1a1d15e29415c6b34fd33736511163e1e191337bd2b31bfa5ffc14f25e4c4857ee99e6
z35e00e35e4027bc48fc78315c347ba6e3fec01270e91313bdaf4b2459580459eee186cca158bb2
z9ea9aa082f8de7a052967fd772ddcd0008fd4f9489cbc067d5ad36ea0c4616aaf9a17786e6eb91
zb3c7ab912052da45b931a7514a2cf0e411918b1efd2d3309eb91182fc82fa73af223a7adad6a64
z9b63bcf24765984802098f20cca2dad62e6f34a5bf66caba2dba6ef1bf6775b7199b35f056c409
zb7e0147bc79b7eeba5c5ba5d43c0f32e63f74887330444145407ff1c85bfe30e6d967ac49f7ca7
z782ab7f6f815990f100ab4286e3d0673eb7d509290924a2608129565d13f64fd78467c160fae2a
zce03383ddf97389a874213a112717996f6d078e18358e532e19be0e1e677c44d20db80b37256ec
z2847e062704eeba7c7b67bc95f298ed1cf92952eb5b877419023220dffb8ff75bc3dc9a49672e8
z772569a63d5f2f7a04d98027b7213f9a8c15a6d5fc9fa47ee438cbf9f468c51f52b02fc7550009
z23438d8f88e3e3d35f647401d488fc30e4d7dcf8a3291b9a902cc765ec6583974ee073551a3e11
zdc8403719905a5773132c95d01cefc9114a1f8545d361a80b186e429ac803c36d6f26a265abfb2
z1a43a282f1061e1ee727a5efcead8985ca65915365d114003f799e843d938fe8925a5fb2e9c502
z5f517ba1ce502b126d9e6d318dd65df828f58873da567477e5db42c42f9090df310f41eb5ae0b3
ze95d54e2c4b114e04290e9c4bed32353be7705fe6f08fefe73b2d335db0c3bf58d74865272225f
z5e1abf476764cf1420b63b921609d1c47f07065c4c3e85e34829f372324529162f6b2c40dcf492
zbc3fe9d1105b7c5edf722bc221586555c1e03ef208c2275668ac41a80d8d03597cbcff41a619fc
z23ee3bab102f35a073406dfb56c4e51f513f14e79b60c6ee0acc993ebd2d5b8cfdbb0f88cb5e46
z4f62ccf46ae5c5d1f60502946596baa67de0d27be30e03bf8847c61ef72ad46cb74fa26b780161
zde89e2048402ba58db9106c12d5ea4edb5f52b0980f0e0026856cd43d48a135afccdcfd50ef644
z6d390f8f8756bf91ef6be8b408ad65a0518272390f8cffa2cb1eaf622690bd5f8a0bd3625fe3a6
zb7f34117067fa2fd7a3059af2a26b0ef01f9f9c5958cc9461d8c678c54611d4a9355200624d27d
z998e031223677d8ca9e3f077d29492077127581eac51e5619b03e2a90f44936933007a2a63d7d7
zf0d5f261f825fcc95e97f2db9425e649f0b6177e91b18ae2f40290c3bc18303850c0220be69276
ze945f20e07195c9ee50f8ba112f1883e8900122d004106f48cb70052405d5f85fc6d465d56b2b1
z85345d31224476316d0d9a08e22ceeeb3d676372686e2ee0f8dc26e4391d5ce6a3ded6e902c671
z3509bc9a2e072e3fe5abc1c69c2a66128ca84771ccf869fd27280968ebb2cac30937a051d4e28e
z634a3ccd6c31f1e3d473984ee7aec3c782c4d2ab92167dc62124c80ae727872d1b01cd023fdb40
z174e993d31a289a88819c98356960302f1850a07238859152940069d003250df54066d9bc58c26
z9fd65eeb3595b10a1069807da3297f18b8e1ac7d9c08f1e1b1d30b447722121a1b785b963d2a5e
zc7fcba0f6815ff80e591bb55be967f74b8501ac45b8007692cce00f4539e4356cef4da0a7c035a
z0947589097a8f93bcc854bbff2733eb54a5f242f4ecc16f5c1ff7bb6ba56ea860e58b9215dc13e
zeeca7c09bb55d88360c1feb4ae8354dfc408a17ff3977e738876d8f35fe6fff6136bca8c5fa123
z1564a5ed48cff0ba04024fa3c90e1b3bceafa3c47ed08b4b063f0c04756c3a9f805b11bae93d55
zafce28be17a8a957fc30e2c3893ced4d521725c17ee753fc59661c6c34ebea7183d27f415c1afb
z848185b64825d6a4e55324d13a87dd3701b7a02406f0ed4db12b0fc3ec1cc7af2a434347f23522
z3a683a0519577b42bd3cc547036de86a01f20b7cda1538076538385d44668b369b8733bf238498
z7c132148952ebba618d61a89eada971c5e79946d0faf06cae29c8f9af1f75e32e74519312fb261
za19d203db13565dfe1ab6d43c7599e5c5f89179f3593d27ea9cb98967b5f75b16dc1e520110320
z6d5ce0db1844f2c75afe130618bc7cab867004c9e776a49cd5f4999c9a996416f244f0d0e04659
z9e3165f3550f2f8e4adca9b794dbaf8764a8cc3eef96056458895e9962a3fc8a15fb6c80239fc8
zd99b320aed03174e848f72f3d8d7b4d5a52a895e2dfce9e6bbd26733a048b0fa38efaa32576a45
z88da0e3638cc776970696f900864d195b42118eeb74ce1f7f53f95790517088f806a8e06bd82b0
zea1a0601b2f7aae8b9774fb7e9f6beab4495a43d066e27be311dccd41b827c06790cd92b2f7bb4
z816a42c8ceaf10bea6968ec0c565ee6d6e8fd9c5e0bb1c61492362c0f8198eaeada597740ab680
zb740b7949a742877dfc6630e81864b4400b3613833c609a04e7151a4c34dcbfc173c25966b5565
zeb7ae5ce980dc46a9c545ddd591868a23a45983e0cba558baa2029ea49e59e4d11ef1a584492a8
z968698bb4157953c0098bc760b6e7a19f9eb9835deca08f873e685ca42d188212a84a16373623e
z60be13e02eab856cf5647307f260c083347dd89c34ef20499f277cab0abee4094889322956c333
za28fea347b1bf4a0ab5bf6d57b1a41a7e9e8bf9b21320e07c35666f8a4629e1083fbae831ae15f
z91ee4e7aa3e61ca69a60dc0c7e7472267b540782cf8682b712c1e5eab99ac0174f18630f2d834c
ze8ddc38b8989c14610814c7b219c9eb4a39f60b5d8a6dfaa8a31321d9a9ee7a085df0a660474b8
zac3080a13074861bf00a43558282e367d2f6d3adc2e84d38dcf69c6c910f18c792fad853398c31
z0f95502338417449efd158a661432b9195bb2da68ffd8c6d1c749532f32aef9e72b610fb60547f
z1514b1f9074015050997c37f37398f905ce0e22263ac730d2108e16f2f72f2df27a2ca3d6a8e5e
z05b1d4dd4bb49225be8809c55b50bf25d372edaa425ab11a67bddd75d5752ddb3b3970e8f76fc3
zd8f6f0b5d71475b1cdfd222d1c2a2f3e0674ce783df51277b06848feb0dfd3daae9e9866cf7d1d
z793baac3938f0a134fd1fe1389c8340153ecea26cef705638595117915dffe2f136ebd9e0a6a7b
z4312aacc2eca8d50c89605a8e3f74e8da38d3f45ee61694a66fc1aa1eb8c9ef2468151b2352aed
z397a9c5c1042d4a2240524c03224b85b73977da9ed10fca8a4e23fdb9593e648cfa6a2693a5f44
z730e40441322deff3ec3777680e903c6ffce953eea85fdd433d7046dee58bbab09b4acc932f749
zbec404e7645932cab4cdc087734a47d610cb850e0959e9bcbff839c2b5e3ae167f1271ae36ef87
zab4125bb479b7cb4c3a383066801d9121ee25015ad3923d270b03092a5b0d73267c0ce555b9346
zd7354aa4bb3d9f82211c2fb277d26ef172c531cbb1d07671ae315e2ec902c3f73a14b5d7796f43
z1fd518baebda139044dd4448a6aded0c3ea8a89739121783fd06db7a0c607a3ceeab5092876813
zc1ef726979ccc2afa43451669b6f2a81bec22d927dc8a71aa906682195669b5795f31993d97e35
zd79d4994e13ba336060094a18c92126a0f9c43dc85e165285c063c63a00c0737d40c56173571cf
z22ab7f0cc39c257a3e32eaa2e4ac9265b8cf8b03f3fc89426d43364b2e743c1cb20128d5286be4
zb74731796e6d397ad95e70fc9e9307fba447703283fef0f20037927883e8d842a4b6364321a217
zd83661de1ed400f9622fc54144cf05aa0c369c2a749e1695e0e8c6e83715bfa1eeb14387dd4db3
zbe9fbd597c9ca70b407e3cdab97f3968507fdc518988dade9061ceb292d1de80b324da3b01cad3
za42c59364fef24f0408dc072539e127288856a10f7307487cc1d40cef2790d93f3c351a9deb97a
z337f3fd097cfbcc5f457e6e09c4a448b0a569aff332a85f882c95b217c8f6a49de3e74593fd6bd
ze7cb71c8a88d6642d424ac62ba414037371f74324ceefa7fc382924a336815d15aec6419d1f3ff
z456742773922c5318ab7cde7d196e40748ee35b1a7bc8d5ad2b4ba69668dbcb10317a82d770256
ze12b1c39af01f63f9f025947691b3d31008320e4ddbd342a14ef2d642a33578ed6748265596390
z358c3574e5b229707ab77a2ad6cec24bdfb3d10afa6b9b1adc5bac119110190b2b0cd4e4e7501f
z90e72bf611ad3f554f5107122339b09c87331e2f52376290029a713b635df04734b5213bf92a28
z308982629d23c162d3529e701f9092a19024d5e94ccc6fd8232b08e171f7378676450e857e0992
z090e20fa4acf9986ec259bca8e635254db78f0275cb841cb45fb6f210b1871eff437db3a7ab0fb
z4a9284a1ced80b4964ea02fb6c63788f73577b121e550d80b7514d5c97fe2e19b6c35a53fcbb99
zf9d2edb588f57f59db718140a0647b7d6e5ab61fde28b4c10b6788a97baa0a5ac7f4409e7f0887
z8cfe79620d97352e9836cd617733cd7e26b504658e82fba11ba0887a77ceeb66a810e1b546681c
z113790967475af7e65ffde7cadd98e674a9d7b393daa1684ea1e10df58e50678dbe89bc07c6de7
z692e59916bfdbe1dfb11c5c27d1ee31f5aee89303484cde6ef9906e8c04d636e8509386a286618
zbda6a93f7d8b4cbfc717064dbee51947936ae230f7097cd973f26ec35231fe782aa29e9752ae28
zd17e4b556a54fcced5692004d1b3de074bf0c823bc131011532c3915f85129a78923979a8c1260
zd11eda27f410e9b9c19f70921816a7a177da1d2c7a8e5b4ba5fcff44dae16b31542cbbb9096615
ze3a41100a9649552f8aadced9e436a31befcc7753b4d1cec1304d1592dadcb6bef1980c710cda1
za9a7ca6fb09690b460ba3c88797b2ecf77bfc3ad446f982f6ad243433357c7eea516fd07b629ef
zf7d63fc9d87261e3c2482acbc34f3dbdc132adb06ef0f2883900b9371855d3cc47356f6ff04d1a
z2f73eb22fd55a73c451b17907d8e003e27d8464f2b9df15d155d30f54610b7234bd88ef66e8e1e
zf9808d46fe109fe5c26c2caa5eb2d767a163d0c12cadbc5167d563ccaa35e6550579226b80ec91
ze91766903f6b3bfc005485e202e5c5783584b5b9662b6294396a22da8e613697d37946b3bf6b81
zbd7998e5cf2498fcdf51427f7c8b0d92cd9b9a53059cf66981d2a9271bbccd5d27a616285bff76
z698badca572ed68e5ebb4e9102fddd9b2f98194e0a375da1517a2b51f3adc55c03ecac2d8686cf
z493b89808bc1c09e6fc380d0d487eeab8c94803a66ceb1bea7538a4dccf6fed485941d543b21d9
z948981995d742065bd9a275c71f1d1933c73f6616cc7240723bd806a53f5bf740896ce1d269336
z9f25180e6b47392890d55855eae350a7c8e18aa2b968ec97e290468baf4e27590f07064036435b
z22592d9fc865e6322f7485a6defe084649b1be54bb18187313b6b6ec0bc7f1d54e3e5db7e77a2f
z6cc18c8d8eb242756d1294f0ac53b3b58afcf28bf4c3b6f2aec92da2036c68c3e0d4b142cc1683
z88ae9f19892f0ee7a226c60037b3d3fb34794c96cc8e21ed918f02ee34446c18bd4630afdb8825
z7945f5959dff23c43e72c44f14e9acf12e6994de9eaabb97281cd6e9d4df67b59c82941e4eb108
z0d18290d52bc46b0517059546bdd93d1bb2e4f11cf69861358e24b7d5e0ebe044b166c514ae95d
zf058501d77fa45712b8ab889547592e385d77cb885593532c7e2c286edb1df24383c111256dc26
z8e3e40a84ff2808f815b79f4fffce91dbaec82618b962308e65d832aea793946d5de3ce1de707e
z06ca772839f8492f94e1a53b14c6db9398a3b452ec5ba8a38992e99c72ed7dc8d9b44954336590
z32958610f89a9a5abd4902841fa96d13b53907305a67c8b4b61754418829e2319676d85ca20740
zd829e99c938333e5cd13a9f1accde89a99468d54810c1b608ee0b128238e15c442cbd7074c740e
z78bc1146332f39e2233c5815303006c8bdc1cf920747c22f34143c6f9cacb8135ca749407a3093
z22a1b23093e5974eb2d5516bf15384a9f5a99eb2f7161a0a3ea1d2390895b39e4e3799f342e10b
zc7d4c436726a5cfb71560c1962ae16863636121dd588fc291c30317055afa3a464dceb126746ec
z0d41f3d87925b077e4eae5ef809255c3296b93d0f109e36dbe707cd935d3fcc7fc87e15f6ef49b
zef01d9639f18f3959e6a36b808285684743fbce23e90ea9132281f57aaef610770bd1fd872cdbd
zd080f7b2263395ae585458b26b1f3bb9dfbda383addd9ec072e53586b8f817d94f8227676a01f8
z669e441c028fa9d5181b903cd6590a1b61ce6a18874a2834acff4c39513add93357c4bd0fada8f
z5ab420b697b32ed8a5a902fdb5ad1d0319699268f666162604ed78463e5b6b9346e881bd43daa4
za1e788a4571eddcd64e540704cfe948aa56948f82fa8b922965877b8489570af1eef954ad923fc
z16ddd6748065037f7c96f918b231e586394f5b362e51a08ee813b939902c1c7a896e0e739fe795
z160ab338265efc7ceb6e65483645961f3147dde1c71da74a8c6dbd0b41a724b29277dc20cc53a4
z6ca0bacecdad503c6f32efa475826d162d21542623a62aed8f3f422a84d1392383415481390c00
z0d7574d2bd1102796718499321c7de9479f9ea44c63e0ffd2b29ecc8b49f2f3ec0a9adee2dded1
z1cb3d2388f07e54e4f722fbddffba380805c034f5178e731fde194e41aafb6f03ee7358e62a0a1
z4513bc542ae4babb24259aadc3147fee350a2333414b2bfbb22b7f48ab4f418fd55237d39726e2
z3b746be18a26309ab38d7bb2736aaa682d9bdcb2d3673fc4b5b02960885ee429028c5292b13c67
z27164ff2c7c101e31151e3e5a400237d2fca508dee041aa4f7822fafc37904f44b743169f8de6f
z61f872ce6316e639760dc7888ce7f3f5ba2fdaf8333ca3b420e07be381221ad4e11c3bcfdcb410
z02ac2b0da44a285ee503405d66264f000fced65a8be1c226c4d50c6b57309b3a6b949ef5a897ae
z37cb2852662998f07ae711509556b2bcf8a9265e3a903194210cff0830c2f4aa6180d197e76708
z14fa47f668d2bb0154820b2e8737a43c7d602bb6e867c3f04fbb7fa9f5a779521ab41a876b5941
z8873fdb8c11c666eeaed55ffcd260bc2ed43e2af8f7c63ad518cf950f55828817a50009c6b0955
zeb6d3a87048ae33c547a983a21d07ad47653eeb6f0fed919e8514d4a191e172b3c74566bf61b2f
za34a3ccd3d90e15923fe73a9eeb5b2a52f4e3544162ba69b476b97164ea12f9ac37dfbcc265a26
zc72858febbade4539728ce19d11e0827adcf5ec7e8b78f0d53ad9c89d34504a0b50dc50cf383ee
z02bbe5ff7e00b5ef6fb946c6f97259df69767e736eb830fffe9adc43e4be4505fbf3dfb9491265
z7f34a485c524d4506dac4adefa89ee5f7024cf8e3920b576cd42ccc96ec3381a1e80427b846e9c
zac843f135db7684c79462504b2249d2c5838d860a19bd6f7a716dc58423761a0c112e0af73494d
z80f1a42083dc7f9a78c605c7c953115dee06b700133c93d84664d766d2320fba560ca2ce359eb7
z3ed5ef6b4ddd2194dadb29b86445dd036889740a3caecc321c474882648c4c2e7b69435b4e72a9
z944b334695c5433ea8b77b1ff6dcd87726cd48f333909b5b9a66815374992c25c2103063415719
z60d2be4139ae3c5dc8e878bbcfafd418b276960ea27db3f28b13800d1cba1b068b0d6cea72dbd6
ze07dfb9f7064f0def7030d87c68393ee62c069a046649b2e867589131f9106bfa0b1ba21467aa7
z74a0add709903bd2743fa0be2824bffe0a379ff35a05654aedef73b92406c98d46ea949270c285
z51fb92686870da370e0ad2bac8b5f5df358744fad1599ac536a7df07783dfa04d680f3302b82cb
z4a260064842c87c995ad2644328e165a9ef143856932117b73bc1fa2e4f402549562a9d07c47f7
z415197e01615af08805c727ef0e4a35eafafd924b1b0346f86171d6c9593eb5400f15e33dd7ae9
z9a7f920e2f005efe7327be81fadd6c472055eca54d19a52b4401b08f04d6f067eb9bb91acc28bb
z7c4c29a7aaf61a722ac5366841b4bf988938aa899ceefa19c8c6e01e6ff8763dfbd6f5af857c14
zd7496cf0ca137b8ddb482a556e3138aa6ff71bcf83560290931661d73b9cb0fd877573ffe89a21
zaac417d112744418724790d59d96309a4c53a2237304adb91c6313613c1ba524ae0fc4b0c448a8
z64bc3f4f1b686ed1c0db3577aa3cf7a2303699bf05a57539d82f7e7ea3f9ea4ac83b49d96a3b8f
zd1f1edb553ba2e07660a17a509881859228bdae419158c6939e14b3d89d3ba55715f087cae40af
zc397e1f1ff905f1bbacdf5b72cdce1f57081c79575878f955a47645a1007702909aba24bcaa89d
ze0a402265c1f164ee0e043c792510f7467743e2075a38aaaec1fec8357b011a8549d6994cfd851
zfd63299862807daf881747f0b7381382ecdcc5676fe766d9287a56676f2f8a2d0762fe287a7b3a
z8e3d88fcd525457f8c3b22cd2c64748f35206229ce2ff5612518e5314891cb2618c81e52eaf1fc
z4d8ab7ddf230cedb1fe1f43d8657ab1f8ee0071b43633f8425854fa3773639432c5c0a583a8744
zd2e15dc76aefd1ce8ff8d0b9524adafa599ad0ccc9776feb38ca6826b03a8f1b32fac28cd2d002
z5dd2c0a062eb48229f0268fb5d6d9e96f9f50ac95a4cab54eafde7385b4c4252cf947c093909a3
z70eb5c14e7043e1971763f29307b9f24109e1421c4ef8bbb7a7a5143abc9849b5aa5092b0a0929
z568304742e55640427c5403f41073a673e2f4c3e09e864cbbe798c931804ce7ce374715a2b7a25
z8baac31faf7de6228da185057910cf0bb9b9935be47280cb22d4ad51fcdb0984228ddb8541151b
zd025a6bfcd4388cad9aff27d34a859486cd91e59a98f3e2aa3e8b1c254c2c4256eaf8aca53cd8c
zb551ad73f986f793701364ba112f52f63df5b1489acd0b8497fcc21fcd0ceb10328d9c7b4850f8
z1cbef3a05e159321a106fb28692be99cb230ffa06b23fd7bfd2bb06b8fd5cc756f1a31ba21385a
za3b07dfa0064f5154f923bf3d36065b86254304ddf592532f4e6895b6ed6ba173ebb51b24f8a23
z25df14c2730d28f9c87775201b5a8cef77c11dd840b5216c59db7a09b7e4ed4267e121581aa86a
z4527dc19740902543f07a9482cfb19832826d803716ba09d00960011b595442b72a3cd42139be4
z6bd2acc72cb72ac44355557bd2f98567ab9799eb82753a9e2e4f7cecf4538ddc1a6b9764a9cec9
z20fa8b8950057f3e579a56a2ff90a1b66c673525e594710e6373b4b4f955a5c2b8e3b07a47751e
z81e7df2aa2f21e264032b757290d6f9d0ed1a3acfefa8443ef1c05397bbd73ff7565a0df506012
zf80c7d6286d050b46b6c5e33ecfaf36e5473e0d1182eb2f75ec643ed4b1d900a54c91ab77bf105
zda960d21fe7e0541bc3c57678df92440609f8a1907800b6cf15fa96a5b606a58e9bdfb99eedcc5
z45a2b3766b06254b51603f39aeb5520395f45558992a51d8e049596bd1c207824469d703f3f585
z91caecb4ccd994469d01904ac9d122178f4f751df54daf11ba844143f50e7fb7330da76c5a1d15
z72f1039447a704679ebb08cc450f9023784caf0b876bdb25dffae1414671b184e41376307837c8
z97cdef88beaac31db1deef43e6ee5320a2e2fbdaff14e86489270d3102c9816084d9a39604f6ae
z1e8b4f6d139785cc465ef0e3264659e7864c8f3b121737b16a9f03c53232fa5a8654f014607526
z9606efd5dafadd4b0762ff8a318c2bc3a9f94b3bb76fa2b3656f3b8e6dc6f0e428c9026c9334fc
z92bf8443452978fcbc3b5bf664fd27ee6dcc46df97bf0aaeb675867558589f9c75d04b2da509fb
z2702bfe98990b23ea623cff5641e574bed455eff3f72bd2a905eba943c4bbca991926d6a213023
z8c89f00077bca348c1cc89aa1a7de192e62a61960590a4ee835b11bc14cfe5d410274b33f2c005
za96f34cb9ce5c004fd6cdfe9550aa6cd05cffd81d562a2be12837f81e2e40c960d6823b8d70bad
z70b2a4f0f7c33c5e5247d3e8fca30a802bbef9aaa8c1f28dc26dfffbd056218afc4a3d1119448b
zede69f3c895ab1db5254ba8864629e2c5dabe5fa0a0372a5b0a1d4e7a51b2901192970ef0c653d
z95661ef9477836be143b10a4047f86906d4470b84454b1854e0281570cbaf2c744718008d68c58
z90c62fe5975a62da81c98d61c109b92a0924a6ce493232c4515d65e8cb5ad913f8f049d4b56338
z05809445c220ab4ca16c31dfbd7696c2459185281c98cadb9873b1a37b70350394fd2a7e5bf120
z2edcb5ac004640f93efe93adf8066c08019548d5f3aaa8fd1dedbaf84a3e7cb9e42db3e190e107
zd4efb689b8face67dff60ce1299f3d1205a1315857df4076c3bfcc5f878961a325bcbf2487d7ac
z82f8c227aa3a71187828d868996cab109ce54bde1c8e29b2a4ba08cac4a10538b3f44af4465038
z14e90f70d7769c82cf5c39287792c93bbff8118fc3d8d8208fc0ab24585bfb266deb7608d1c157
z87397e0bf653aba1188d981adfb95f830a09b735064746943271b7ff578c9a3169ef816cfe961a
z98338b0d1a582ad53af8b71e75212bc8b57fc50b64d1d603cc31cd6e06707d60b4d9a513f4983a
z15415e518a4cedb1676c713b677508e4b82f4bba9442f87e05a795f0de22ec99d59cea37a138a8
zfca755333c35c699bf5fb2f1a888264068ec3d6c16e7ba001795bada3506f809f1cb18c0d74881
zbebefe048c99f75359cafb27b049e857d95d3ca4faa65a0813058f766bab0d3502aa88b3773f16
z245aaa0e7bdb03b0c29680af4c4bca41e781cf9af302918870ad16b232b7b29b6bf34a84acd915
zc2569fcd627842c525d7e32f1a46af14c026e88e96a240b32ab774242b46a492e97ebbd65af544
ze1a4829a522765bc2f647dc9d8ba3e6ebbac6fe812408bd75eb5025a76f05883b834de03595e7a
z187b2036de1871bf3e25ef8d24f270bc62de4e8077028b24a5c5cc03376021dd05b10a1b2f8fb1
zbd8782815ad97a6cf33a05af66a78f4b3fe1cca10e99f323c7181ecd5b1003c1f0ee7a3ab3bd05
z997e7f7078c919c59a8c3269b3dde525816550042cf256fdddc7876a97462fed979edf4f72e48b
z6ab22f86dff428c9277ef3e5176f4f84fe312a47358956f60c53db35d031ae4bf74b6b4565ae5f
z0e6f2ce48466be61696da0c0d4ddcd28dd809ac4c98fb7f91a394606e1edd09f3b93f69799945f
za976efc9136fe3b347f91078a404d72aef85f928420bc0a374e35dbf6ac44cc36910ba7ad3128e
z150c3c0898aebb2039ae39dce198e2aa004db380be4939927644c800ab0c883c8cfcb0136781f9
z61d1485adca277da40b88d33b5b7630c939536d80127f54a174cbe169c82c452b36430d37b6d10
zfcbec152b0ddd98899b9b798e5c64bd981c223cd0a3156cb63cbec16cdbb13b1d4c5c7855f7c62
ze595a4327ef26b65f061fa6101dda30b8786fb6849084ea0ba21a6a8ead4d53a08b7d415cc5d1f
z744d986c2dc45724b89c713d9ee6f9c0cab6fc6e848c1a9fd53320f71fbdee8e2467a33a450f3c
z68b550fb27d50f5e04af77e4258cd667a1ef31707859ed259b8d5a39cdd7d6af13fcecce5003de
zca62feb56cb986ebd29e104f2d3b0a44c7c874fc6f3237fd09156061e60dbf05ff2efc65d630d9
z785cbce268605a0d7cff5c32227435ae0523e26bb25de31b13c0976e22b2754e0e0e819da81bcc
z162f2c4deb0f0fc0145fd987598a4f730535033c70816c39512a1ba8461035a2b9ee227fa288eb
z26d84f27a8821f469247c90c19aeea78b9b9da0927a081781592fb258306e338c14205c57de93c
z713bf631e01ecf1dad43864bafea94b7f3b7e01f832ecffcb74e3abe9cec4fd608146ba7f8062d
z1c06145b1e771cd46ac391a39accd236bc928f26fab5bfeec5089b972e4f1b80c7b090c6c68ad4
z09d47f49662bb1e824c0baa92ae4a0a1efb008ff4de8e3c0373528f7353228603f67249175d45e
zaacd65f4ab8c36486997c54404c71cac726bac244b6df197c727eff99bc436f57dc3e599cff555
z4909a1e89352ab05a50c05cde59fbdbd82ab0e34cb16e2256578c6df785c702ad823c29d747f76
zb7932e37fa7bcdfa5e6c8f724d486763da3dbfd16a0680ea5b48ecfc5d5390e5c682364e45d561
zeabd71fe330c1401374aa3c8cedb5327157c47fe3a9afc052c57a48bb35d4d1da005c56feafab6
z312822d84e1450497ae953874f4f8adf0667d33b804538f8ef929d717028da4513c0819e6c68fa
zb92567e88fee4e7a63af404ff8700f576f4a1b25fabad8c6ce9df78d300a61fcd3e1f8f0bf7b70
z9fa2a001abf42237670eaba94a82afb7a67827ea99d3f66e9ecb9a1f0597357c90e240e84a762d
z9fa4ba33004b8e74d06c8cf0957afbf969ea69c3d7a1fe331d7b715551ec966efca967ebbea3dd
z06c14b12f32accdde51bc9201018e3f703738209a2372c9bd42d0f1c2d9fb4a82ec65211a90d8a
za87e6b34e359153df2baad09977a5903df2a2917e3c52791bf8ad27c5888b8762cc5ebe32ce49b
za321e62d7d1adba8169c7aaa79c40f4e071d118c747d82aac06b16eaf8faf9db00e08dbb8aa4a2
z6fc9a24a4155761241d2fe9ce99bdae21d7114f5de782cc0381100f90632d681e40f95e6859d89
z4a5eb0ca8b428630488c1db83f5eee97564db34660b301b36b5b0b7e0b35f28827dd92f13552d3
zb1f27b9ef5c6e96dcfb9c7c1e3e74ebbc3c69c06c180b0db208903ed96f1f195576f55b4841d48
z837db6daea9b11e3755e5af56085fe1e4b4c812af9769cf4d118b0a5898d9ff75c731b7258b9d5
z1c231d45641141f7952b10beb08ee7131ede61e7eddf53f8091f01afcef04a4d8c47d64aa5cbfd
z1e3278032db88791ba9ba4d45813597c494bbdd8788d04e9c7a09acdfb1076645954343089f0a6
zbc730e3ee213a8171c1d91047e9418d3c6ab64dde425432828043ef1a10e595193145a19d35b02
zcfcc05175c23c83faac4220e77d60c347b6ee32ce2af17a297a930e8957fce3d04ffe12e5eee28
z16119625951665d3dbd7f36f7e6b809d3c975715eebe7b65356eddaa1eaff243a68b2ea452c2e2
z6ae8f24fbd6e7a3b2af3d957994cc21bfd1339701215a238d939949ee483e34037f36f403217ae
zb8a36872baa3ee92fc340cf8a1717314901163022f8d7db524496fe9c5e43859f88f81fc646636
z08df09f49253afcca038a3a4cf1d35173186f8e7fb0b4a10251c5dbf158d8438eb605f4e9666ca
z48959ef5cd67086b41ff46a17072806ef3ca38091a03102120ba56093ea01bc73300e21e5f2e9a
zddd18bce31c5ff2eeeb036a9261420a44d11463a9ece2a5655c015c65f61d164a6ae2e38cf071f
z91fdf47880762141bd9b34c38b8c020640d37102a1a3830fdbd165f021dc4d26e59361f2b47a1f
z43bc651ef68a1a8cc8908e0b0a2ce9921bb1ec4912d49491f4bba506f5d3be91f3c3c26efd5cb2
z6adb9d26b4c95bfb0d60d1c7a8ead44777a88e8cd9d4e3c6840276b5a55222d2950bd4fbe96bb5
zed877baa87233bcaaab5cbdff13c4f9a407648b2a652ba3add33a0d12e5295d14d02b56ef06d62
z36b11f13aef2fdcc63560ff8f99f3f5845dd28e49373d4ffeb867ff131d656e86d189aa0ea4d2a
z12beb2485652ac787b5e03ca88169fe3b10a37cc769aa25e9bdd78b3d357fc2d832d1b1928ca06
zca729874fce2ad5cbfd5ba20036d32f730f32b9a669958e6c2c40b1f167dcb8c05efb3013aa017
z82e8da346f5711482761cde1b8a672e8548435e7129f36c6e800f5564deefb8eae88d768ee036b
zf20e7f9c2e0fe334168513c0ce4b3cb00bde47f163206bae4d5b3126eed3db9e08d1169f9663c4
zf928e05023e2ca0731decb155d93dec33f582f5f55863568524d0e920e06d408d17949bf547147
z5fb58790d4008b0a0408e42e632af2930d2d5dedf830ba0836c96629d7ecc42685a004dcd1389b
zc82389026fda3688e69d7c25ef4a2f83fbb688ae1c37de0a74107f2b5e8bd5776abf7ab7577b96
z620e9719bf4c318ddf5b81b926da3df75867a7f695c7b9192e126d6bf75e26aea3e6aefca2fa5e
z5a4e3c18536b9d2a9e1068663da3d8f2162cfe98341ebb1f34775a086ead03dfd5dd256d46df1d
ze9852aaef651579d11976443b925aaccb3993df054827f01c2ec7ea6024bdc2f3b43b667033998
zb670049008bf03ba75e525672dc617930991bdd6101accb73398d37f37959f3cfd8e72949b5213
ze29aae9874e3731cf1563c481c7ebdb3cf7195cda589a47309cb7dc174900b59382e07fb45986f
z448e85233e55bd1acc310d8a07b0038cc7120874c12528d3e54640dd37eb838a62cef4a924c4c4
z6000249561ba3237ee709829f6b2d45c301ae26db7ec238a1bacb27a481a3d5641d45a352851c0
z7c2c459333dafb83510b7f0bf04b5c54b8e7de2bf963792a457cb6358d5befc04269009d184238
z1ac24a8840354516cda3ddd706acafa391f5c8720c748678a3f63b7d1b6cf8d71338bb682dac71
za6461fcc251b55a1b775cbe55f3d189ef8b3ea13ab61c398af439e9320ec0e92a704590b03d0f9
z927bd11dd8fcb85464939ebe56830ebe804d6d8fe4527824f8481723867e72ef7499495d59b9d3
z2795528957faec7574d190c7b7884b79466d8a346079a0480555e6be07b4014b12daf3208c14a4
z0417e9d55272d26bb1679e90005647ce4fb7d10028e667c9e6a27c39f06e0f68acf92ad73511c8
zbb9559c01f11c0ec518b5deb96e962b231d21c0901a8bcb24c9366c0bd1bdac48a519fe609b525
z63b5f1e614cc6d2f3316a6634db5934daf2f39928653defee396a63cacb6cc671bb6783181ac04
z8d45965221f1a70f2a7f1afdb62e0758482f8d03663748714283706ffe0ba10a6a48966cc2fd82
zb2c13ea24d28240a40d4c482ef4c7fc7540be5d4ecc962351efc8d0cc6028b81d604eb8889eb06
z7ac28fbfd21817957d743722ecaf48562860a0110be55e45db827e58b387d19fe680b2fc80b203
zf88c69910754d079a92005c846eeacbe82c71060c2ba796b15504d9198f11ce86959f621808614
z36505d0d54468622fea43ae2a4a8a080916b9033bdebf07fa8b5199f9db7b77d217528c9448c97
z97366dc1a13a19a67c77e404bb4e0694c62ac02bbf3013b89bb571aeea0be1ee014d2b3213b970
zde1a89c92a46f7542c045a0ed8743476d377d17f2250e8c06a1ca3ca8fa219ad3c6f2d9c0e6795
z0face06c431bafa822e0b632e6380ca05b14ca75141356d2b520234b2f1ee9340ca7412479c1ea
z7bc31aa9d81f873e9c6768693ccdbc77547eb792a548351c2fada9f96c0a8278af9ea5808643c1
z28dc3e64b3a9638f533edf41add887012c20ac52897b1497791ba36b89ee0331c9b4f9ae03eddf
z387cacd6b8164a2500d4c29081d2774b63d5e327ce0303874dc66f03eb76d76b61a2fedd0b0703
z6e54f46428dbdf79d615bb89d8dc47c813b7f6ffeb2c5659130170aa0c5647a82571eccf02f420
z02ab9c86747903b547c50ee193b3797fc74ad8971ec130dbc4fe5d3f8d21d0079281f5241f66a4
z989c64ab48c05b93b5ddbbad6af9cf80927ffc081c17a7cc9984cc9af95d45fe3d19d600182600
z4d029c7246b78d73deb8731da95ee552a8ddaee8b2f8ea24865d290fc02670119f51aa0558fc56
zd47b0122a5e91c1fe6baddc18a0100991e6007fade90d5541419b3d3356d355380b0177b6cedef
z60e3aaa0381e3d4bff6ef387548c07da06f882301e8fee0b38a0931a301f73b928e3315944a52b
z7561e798e65590f3548947b52e368e7ee06426dfac0529673a83316b7243c85d700d10532727e1
z9d6f6173dc6b9b32030c2da03929a93b93424cd6cc672927a61cbcd1263f5efa24e5052b5a2687
zef89a0e731295939ebde3dc1e28d873b1b338e2d65fa817d74f7abf911a09e1ac10c4247dc14be
z7b646403d3004dc8490f7128a4ca908519cfb1090b225e26b4f8aee223e35b6d138b79fe0a56c0
z3090a876fcf48d9432df8f8966226421ce65b2b13eee8c272717c149552907dc656eda032cb2b3
zeaa1c328bf8c30b59684982149cd0714a7622b83531c7dabc353f036027e87e8e326036439d825
za1fcce6fb9d25f5e4244382d3c8094e18e183941072dbd206ff5e28406ded502e787bda9451fa8
zc783b06ab3f14039c695a0852ab6d718033904c52ce7ca14cffc6a310c9fba0dd6b24d45572f6b
z0a177ea7c5a96c7b891e1cf8b1ba2ec5ef72da12d3c0e26fa835b884f747b31fbea0a23fb0bc8f
z9e0da6d45118dca904c6baf429427aebe7bab272b224efc2fe7ec542fa3f517e293d0dfe5458c4
z4e458ec0348b84f29d99d29b9ce82717b47883770cd9ca56ca1c08314c688b3f97a228565fb2b7
z899dd6770ff709a5a6675536edfdecb3235b376988e463cb89414838206df3073730258613f8ce
zae2875fb31b2937c0fcfd606f3c2238dba4a9e048debbfa2768d8716098ed34b9b5fbeac9aed40
z17ad9a64eca7955af782a56f52f958c9713c6b32b8bbb490ab02606cbbf74c445ba2e99ccd9183
zabb7f890998193014a4e7f2febcd854606baacd5f0290a7faf352a481cf7cdc261bfed362cd949
z210f9435eda90ce421b7e5ccc2238a747e7fb5a6416f3226b572675c2cc2150d222aab21b44bf8
z7d4085fa17335800a5b6710b17c6c3371b13550ac0d07582736626cf1af12f1d7838e252983cb9
zd3e05cdbd82addd16a6bf6601d4e8ade21e1b84e202b1cd33f8560ac9220a739644c023893a895
z7327b7373f524f780f0203a18fa17da8797fccbf1ebbacdc40b7aec15e33b1cd6ae0db475a476f
z2465686b05b34db62c30c6d54a535dc12ff84d84361a5a9eed6b5b46ed3bcbdb235126312b9de1
z4aa36fec91b03ed157107929a39d8b3a51913d1b4b7ba26261cfe7f5eed95c06d8dd3ba8ad4901
z3f3bf47845ece83cd7374fc8a6f1955795b0c10ff74a373062166cf1a203bd5137ae0461859ba4
zf586eb6312d4a62bc8fa53436bca0f1c6f930b96b589eb9ad4a87d93b65aaa7b2ba7476e040ac2
zb08e76c7220dfda264ae2f7b0c2d91722da2338df6f0ff6ae80a374c3d1ab285408deca8bbd806
z1918a3514439d9ee5eb477c8a310991a2964791c0b7aeea49d799b5322a5d063903eecc231db44
zc20f55e9d41049c6fcbaf0ea46cd0e5ad83ea256dddf433f3b8258f2d31b1ef34b8d84f7c22b40
zb75c0bfbf14434a6528aa93c8ee62d4d5e3b549ae16ff56e1682bbc1967c7e5df96761d5513086
z2b664e44c2c8e1f08f4103f764bcd5fe13da135b31ff1f308a062c2bf3a96da866c57ce813fef1
zdb4469adc50690f9f5365f834e53b353341307745b0c706d8ad45b7cd62143b8cf630827f28638
z7e48304ea78671b897cff86c9c23877cdc59228c6f18ad505ca66c1ab2b2130892412934316e1e
z8940a19389966186a08c89699d6bf83a80f9bee18220c2085b6e218b9df364f7e90432dc7a40eb
z67f7ed1ac1c6483c61e8405b830503b9ea3210240d7c31ea2e5237c3467226c90e40f19fc6dacc
z6b57ea68ff84ff24845241aedec84ed9415098979e0d1f756d81bec65a6fa6d1045d61eb7688c9
za98005d192db1d1cae58b342573c9380059856731d388ab9a5e2fb4e0fab54d13aeb45d7ac247a
z117ca1a8be83472d92f7403d72781f7e4c26372586fac60eb326b75a940cb54521f75c0ccea6d0
z8d582fe7fe4b2f85a3bfff7f65034117b829c1fc3642b2e26070a0e874f66c16fdd99bb7c31628
z13989faecaaa3bb1987e81fde392f5c4573d892ca2f5529ac1012f0fe45e777d9734e34a6cc30e
ze1dab53f2adfff446fe711006a90ba9adb6b71482e7c1764e9b68a1fc925829f48f4105e885e54
zccc65a1b26cd237107d4007abbe299959c24459a56cae132985af78d07a8613f4cb8b6561a576d
z0e3e4d6e6dc11f45e81425b8e000935d239fb16f4ec4ff73d9be4d2597988d982e9c238b7ce5c3
z7b44928facc3e6be4713f3a330afaa32fac95a0103685d390f85c042dfff0d7a31c8f917f0df6a
zbe02551d8c31f72ef55f83e1739bd07450c29fed2d7b6450f5d8da85f722e3d55f00f0d9fb50d8
zd5585705e3e2bf5759f9d0a15dfc4813b41fd7bb9ea40279e41873326a98afb9c9f40c5af87308
z847325ab05a5afa9096b46c4aae410330a7ac53fe7b8649b53fc775ea1f01e43a7fa8b3640fc5b
zf5d8beb3b31492dd0ac00856d9deb0d5c41c9affd104e59b193ecb72b9f896f75b977fea8c6f29
zff8c8efb4d4fcfe322d5be326151bf5fc6d2973d441f0d8d2472150f36d6728dbaceb64998d38f
zc056f7e8da11e49a072f1a17a077a9792bfa145c622d8ffaa0b469ca0131707c1cad708dfddfcf
z3a66876820f276d9d11cde0acf4b0cc616426483d6f472851726d7247726d2af2162eb7ca12191
z8c67ffc0da1bc3cb2296f4b094136aed47b4bd47fe002dbd383220820bf6ec5f35a8d82e8a0c26
ze5d3017e1c742431b5307f605f5018919b37b5f2ebb5c04cd431f4ba79e3724461c58bc3e0ef3e
zaa3628073dab19c3418398bc76e4fd9b9b537ff855cb7e3372f27f1040e9e73d5ad4d795779480
z615887e5813b3fc83833da47d6799b01805b294778bf2096dc535a815d2d6c8b95bab562483ed0
z407eacdfbfddcf963be1eb7525a1c75699f300ba0f74deba72a3b970eb801714af11861dbda6fa
zac873295ca45a92faa72e1f5e4b81e252d9af5a69f73fd5f36edf3e18ce25e80ec3da796ae364c
zb8834c256720802d1c7ed6d356b735447282faf466e12468b196fd4c6ad2691b65e028b3f3da7b
z1fdbbcdccb88c86a0e78b587ba5b83bddc336a72fafedf6bc2859ca9dd7b22db461e63cae2a6a9
zd55d6f8992a198f0a629f3f154b8ea24e0bf1d2e72ff85b9cc172f8bb82ae312b1ea792f0f18e5
zeac288a58e1525bfeb1868cc514619b1a1efaf0615bba7d65a8b7ae3e650e310497616fd9d6874
z2c1fbd1e8c2a0f531ff5e115c37319049f3dcdaf65a7136fbe3c106a07f91bda3cb9086e749b4c
ze8ec69e2be84bc7f204d6fcedeb74b225a89ba319a3f6621a544b9fb4819abd350549c0d131add
z986dfabb3e785d649abb627ede2481b9c7ef08fdd4d2c8c6cc0ad225f585ab3df86a86b1676d3f
zfb4d9cb7cf648bcb21d6b30ba9ba1c957dfa01cadb47a414a955f4d63784c23a8333ed2670d766
zaf5d94c4655d16bd17f54b088de1c84885cf42a02ecb9f5b0a0faa974c4246d7163d55683bb565
z1259b60f2b3b810f0152353f43fd994ee0ebd4084f4902185b4962b8f9a41e2b61a2fae96b3c0f
z8af7a8731b0411672b6ceb307754eca099b8044661cc3b65c9e9a1791252118dc06aa0220c9035
z6ca41dd05e60c4c3e8fdcc423d168e3cfdd08daf507a2399cb62e84683b3b6eb0c82eafed88f66
ze36bf63ece57edb8cec32944e03d4c0ac9823567be664e2f2c8320c43713f8ea08267e99701951
zc8ecfefd2f96971ce52820abf46c3a73569536b2b540b72b184de462f3b07f0f9a94d01e819bf8
z0285ee059ff371aafc0b9d469575c1a7050dc160074695aa107ffcc3cc465ccc2aae973a71724a
zd45bb54a844c2d1a35f1701a7d8a451ca4867a4ccc5d661c165a4c8a328e8fbca10f1170be7410
z64303267077570e1c292ac71c322c9f9a100e1587823e80de7f0bc99b85b35126b659defb93e49
ze2635aabe4f947f6eb64d66aecc0b13f66e5c777fb638fdeb3cffc4042f1769e6c76296733f913
z9da9c980f33ce15fcbc98671fb6f2724223dc67b4fc30271ccc41e28b314779f2d2922dd13a345
z9e0769b19df157ed40a93b30f5a4d576d05e383c6aa83193b1748e76e600f1da8d89d162a7edf7
z1f6fe57b5eb5115e638b574f3b0f11ab507dc3315da012f62980af2517be223db58c6016b4b44d
z57018e51470976774950e11a32f234497b4d07fe2423afaca499620fdb59c19b644b0ef0eb82b4
z3903a90e92764da3121809f1c3460db03baf31128a8b4eaa877892c4845b32eb90c041eeac9c2d
z4cfbf532aaf8dcf0d3686c5cd6390401c6187c3c0c63c45e2775c3cddb7ae14a05727dfeb8ddec
zaf83887db3866aeab5f1c75ee30b30545e0e0cf555390ee333c488662191dcbab6e5506cfc5bc6
ze699df55f1a8b96dc49b729202a4328c23a38b8ded66a41fb596c031b0ed47d18e76051037319c
z9d44c04590f15c26a7bc620dcc33b6e76def61c830e35fe761caf05b88d8bffac351d1a0eaec7a
z90c99c6815c2659a240f4c7ea8af25e17eb81e4e39e828dac8ca368ad947e99130ca3ca1ee26e4
z98619477eac347427e9134021491dc23d86962ab5935bf7cab49cc1200301854c3bcc34e6f6058
zf7f2899557db005d881deb7acdb9343b3ab7807b79ddcd22e22b5bc6f8709577a8436b1bb3573a
z501b1b22b1b2effdb95982fa173d51915879b2a1cf2fe23a67acb3307022dbc489ef8416d64316
z144bf677338721596eecd2ffa9f78a1d3247f591edfa8c438116ca28cef0e33b3432bb11fa9aaa
z0c3428e2b8eb4c953a0ea5ac437f4666f0f29b60f21466fac40aaeb4af16f84d138dde9f4b3bbf
zf84a1ea0771eb502c33e1f1e5f5fca15a31b47ce8957b35fbed51bba6261b907172072a6527c57
zb2dc382bc7328b8db0cb608d4e1b08672fb15e139bbeab5e3d8657e3ca6ea5870a97a0cf46f21b
z59605aaeed93ef37679ddc59bc054b1e3d0cc298aa49b95e4517a2c804d1d7f717e21f2bb39a50
z8f6029ea9cd8fb0a80591d8dadac3b2b1ea6a2d1f13147f46f0e1f30dc3b0f624a9aa09ddb2993
zf10b47cd6f9625f28dee96599b4c64c7b832727bc74199f5887c7b4f73c7ceaf6bd0a0b873e6b0
zffc09e94a7b6f28396030924959e3deedc7623b4f71c11fc3330a7323dc7e1ae996c02d3ec7ff8
z79eb2425e769939504a8a1d42f3ba9e57bac7fd22bdcc74a610e95d497d048ed34f25a0c6560e6
z5b0268bcace3f0f09bb35560de454ced000991cb28d48cec7affbfc8cd38ab4428e108880ef9e5
z1b57fc9f15ad2cc131e6b06e6fafa7fd7d68ea5fb2ca0ab899272f44cf0f7dc15916a207d99fec
z55696dd7d61c33e503ce82c3387523329fe5c0fb5b30f712def8b78d4b9ddbd32fbac2caf6796b
z0442366855279aa77aae6640d95ff47d3ce48300106e5b4b6871f02411b0136d8e354946493e6c
z3b509c32700d28962c3f144d498b062b3f133aab1b2e1f68b27676ecc5d9a2231c3512d7cd68b6
z6c94495f2656f0a35a4aa541982106a17e7a1c1bedb3e3a465048d05fa62b95bcbde385f27ba38
z66c706ce538a2e2d4f3b188d5f0fd511489e4495acfaa9ebd53d5b62ce46a21bf4c8f2d9c53a96
zdc7c12cd7bf4b3eb9676ae93333f3851af272c4768246c4d77bbc2feec30935e1d2aabcce55ccb
z8a180dca749625982b59f0244f54eab3b09c4ab4e17a0ac1ac09188ab87c3bd2b3df0ce83694b8
z6234821f223721b4c0df1f95c21e582ae1f47c3f88f6daca610ae29a1cb91a80d5b6fb356cb04c
z745d06aecfc11d080b82ce64fd6f72796688f8e3bf3eaf99b917fa2944d3d0417ed1ec6fc11335
zb90dd7a4c3e4dea34b011c1f15c0271cc6898d34d3f8b0eac1481cc027d5a7911c295376027362
z057ca73b0cbc8b6cf4804c1f285b44e8bbe47b744b1333d1aa491af2bd608ab27796007df68cf1
z83955fc90d12c4412f2bf1e4196bd4ac334c8ceccc92359984ce568db283039cce713626479308
z3b0ae46e9470c2b272267060467eea2be043e90fa78e25bf9ee6066a4139dc7b3d05bfcf48ad22
z9d08b5b949bf2e27028f9092b3870682cfed0edca6a58a9369e24d99ad51ff05ecae2caaad9bff
zc43a928f72e82b2e9404ccd0004b335a64797f53057f81550236b6631177c7680d8e61ca6fed16
z64fe4364ade067e70787946218ad079b0df435cc9011facc46af5f7112154873a4b8111b5c15f1
ze24f82da707ea18f3404848242d35fa37039fbe8574f85a1a8a47c34a598e3bc18f08fa9c6b219
z5ac6b4c81ad48db00bab9f2b2f5410ee46a0bac44e937f76b7b497f3ba277b3db0d88370543001
z88f3bdb0fcab776ba8e0bcbed29f6ac1ed2b6a5d610f3b08b0b0bf400e7e842099bedc4da6bd31
z0f68f538f9ca9c2043e09f4dd9bc6a93e7d9246727eea72746a321ad26c62234e852c58785d0f4
z52b3d44c8808cdc2b9a31f813255210fff6265dae0b7bf0c6b465d3a43a53dba08d94e66cc49fa
z2f9d2e88201c72eadbdb825de96b589e4f800a0b71664520098853b44ed776b3160b0613317621
zc7cfb63df1f37f48d64587c2895af3fd585b69bfff3f078678600eaa37f429e0c1ec1acf5a40d9
zcb8831f1640eb7d4434d6d73594006d8600841012af612786b3181d101592f596da80ceb6133ce
zcb2e67bb879ad73b5e29fc5775cf92b8968bac1ea56924e07ec5a00b76f02a11062d606257e05e
zf127a7503b3ec0d6c1da35efd9266fd3899c8b8fc2ac774c577b348ff9190efda6c54da43bc644
zff3689912767b58a13bbe8fad8e5e445646e07a80d66deaaa261cd1ed9b4105a954d76bf299d2d
zfcc39bc22fe1eb3f85336364e0f323cbd86df8443cf982fad63c5c30472055bcd7a279497bd334
zedad7da8d244338dad9eaa228800557d4622f8b1f1494ed696b8916998807b35cad7efb1a2bec7
zf64393062fab184e1f249d4f5acee4b0c54bd467778f583e6fd13d2332cd6086026eedb64dd73a
zaf1d525ed8615a3ec4dae2682f9c2a376d47e3a321aab63adb6530ec65b26c6397927d0b629463
z57fc3916555f963a5dadaaa73f394b0f1e3baea07d0502f6d4b3ff42c2dae0925b3bfd421148b1
z46eed1dfa1b1e13e74e4000dc9dbb01822daa84e8f586cf75c97b62116e0e3762fb434e9c55b23
z1f8e1e498686e1446b859eb3a80e7bb05887f116dac45cb87caa001c9eac2ef495b1eb69162e78
ze5dc6809c37f538c9ac66335cc2b869b4d56d7cc0cf62de6b5916e63be8806cec2aabe6154c868
z8a6f5b98046be72a4c68f37efc19d27155c06752342edfe197467ab237cc305eacc78f9e95f7c9
z3b9e4e1796ecc43c69c59f29c6147983f497759fe4281b0ba00886f6a52be6e5307e7a943780dd
z92b638a7caf60d7dfb37061eb0eb396cdf27a2f127077326c0d719b88f5ed0a7c6c056aa298d46
zef7ad9cbef39dd04a53b0dc4a63c0a1e79354a55b19c78b515c7f62349057fd367b1c5bbc06b78
z8abd5d0d1ce7b49aa9f2a977baa26189110a9fb02f7f26c1b38f1f6aa61341cbd1014428bc0e6b
zbe1d92ba44f4cc8c70596ade90654abf2bdbd340d0e9241ab2fd49e928f09161efa3d3596126b3
zf27c2b29ab92f629d843cef29bd9ee1214aaf743fdb106e18ce2507baf0b762ad1ab4ba6372e60
z204da354d78d1c62b206b9ce18258f6738a14d14627b77ad167fd5736d6a3bc11822af1ca0b8ef
z727a1af47545b154db1a0c972ec7a865b497ad3abe71120943162cf75f7743456824521d0b38bb
za61ff2ba9387415d181fabc234b85348cd9daf072dda435ae90db8e1d1fd5d1c586b005e43b3ed
zd7a43509bf4312241a865eccae4d0f09829347f116f01c808c5e899ad297cb3d0fa5051395796d
z199a265aef78baf5e942555da17454aa83fb4c04f59d629eb52469e711e890b81dc157a7a01f99
zcfc9f037198ecf9029afcac9b97d2c14292dfa2182d382e700c8cd158c4a7073497c8c72287b3f
z4d6d23b898856af484876f955a45e2f0848d781bc8b30ffa976aa26899a02826266019a4b4b046
z87987534eeef36840aed2a71110bd71a7936c040de5bdf16364dad22e5a52f775bc14ea2b4429c
zc4290a4e6acfda124f505eba1bc91f036edbe03e5af32fbc1fe1646e73d9b8903938d4826a077f
z912e62256375186f4adef4cf1d8e683ac6a8a6218abd57d338b8e8ec32f8628ddb30e3fd81d828
z77edf9b5ce36a11befc188b7c86343fa55bd4dd411ef2a5376a29b8d63b0e97f50ccfdcd7e2016
zaf324f462563671fcefad8c1646d15423813918cbc70d14f1d2816084b32b7773aec27b9d414a4
ze005c40307296059f8ae607c4165aec56c240e54904069193881cd86c8796e1348896579277373
z11cd16c02845a7ecd4324dd20452a7040cefe33b0da471212f1f6095250426cba8172ab329d6c6
zda1e44005ced5778c1f55e0ff3b1f5d321aa05829f619427ac494eea580445a22a226da60ccc95
zc7ccaa02b1f635b2f1186258547c2499f4051fe72908ea1da0f9eda411ea8616e66383df61b5c2
z12e665493473de96cdf7959c1bec2f1d48346fb034f9e5ab8867622f19a160f763ae30fec08871
z785673be325a07e1813ba1c61cb0754ece0e970095d35c82f94a50edf96e74c0ba631ee220b8a9
z44e1fd05ab825ed7930678d10f8b38e4cdc9f63499f0b063baf9342f8955b1d36cea5103d5ab35
z20e5eb7bda605ea64505d0837505711f05ca3fb93c2ab8af4c3c2902d2ebafba32858d98083f98
z4377a637af73c4be71546ca19c97ceee2fd6f6a371519bdd4f1d4162f081f774556aea99a38d72
z6c7b96ceb68865c7dec2a66fadc95975c16b93a3c58b3aa286b4aef626b0b09e0cc01686bfb427
z0d61602ed859ec2812981ce8cc418cec1db5aa314534b8d051bedcd8825214f2d4c3331c11ff08
z04c796ee3ff322a446c94326e0da122c92416f8731019ad9b7842f203590e2e9c2190719177487
z0744215d5232168507eb5f831de3c209482ed5b2d46ce3956dcff64b130221f7dad597f307fd17
zf1a63b85f984de5dc6268f72887491dbf515f1ebd7c366f07f2aaddad42f782819e4da63797a6c
z7402377bcccb7a5b124ba8463d33c97c6160e69809a94752a0506aa321020537adcdbcd5c40c02
z50881b0d8ae09347c50215a81f153514da969578e612e83127a1dbf3cd5e3f22f67777a1a94f12
z3fc802ffedfcad9e2a0d223857d0a9fcba1feae52c5300299bd8db3a7ee6a8d0f28f29a94307ba
z187082f73c470463254c0c9a2228017c3b304ba99dbbcfea09b88162536d7708ab314816e4ae18
z27435192a15adac437d4a3b304c721b074572042fc4daa6e21e48ae87c54bd965211e3dd3488f0
z075f1ef84369b807a52a548479b12c0cc102c6836ac74d33ddb2bd85a56242906b28000a4110e5
z0531f7cad88648bf19d5afbca1e70623821f8ba7acda8e4482b25a762d6c71042749301b0a0611
z0475cb1eb851e9c83bd1a7853b6343d9e1152f28e637d4538dd8d254b059e7f00c14fc05a558bd
zbdc72451023396633811dba8d9443b8aab6ba7d6f1c7a9b0c35b276fb1ff8659f5f0d91d5c682d
z22b70a8cafc83efa801a072b41625d3b017ddeac39def08d916de615b3fb93d6e7c882373217fd
z615d7f2e834785ebb5d511ed49120f815db5da8e7bf9944a04979ecbf5d5c5549c1c3012cac53c
z2f65b81bec360c2b733e8d1d5cbb8ad7265969c89f6b60e4859afbb7497a153a3089dac039ae8c
z77805198e8798899545a05200986615b0cf6d790466f88fa846f9487d13a0471f74ad48acaec6e
z0b3e5143823dc692badb84b3462793f3be29e703ca7243581393c9d04a0d4c44a36ffa6695294a
z26e7c25bfc7e2f33ea43ffe8bda5d054a71b1e6267349baa5ae0808a86620eba264ba277f13b64
z85f00ac9437cce90d9622605459f8159eb47369d5599c315bd485607eb433a4a50124167a3bcae
z8cc2778ce404c2ceb07e8b88769a568e3772919130b2d1e8d87072cd06f5d63b7afb6b284b4edf
z4101a3638e7187f3c2c9d4e1782d70b22236b2052d3ce7f02b856ccf22c082b2a4fa3c73968497
z68a80578f36a573551fc9af815fa1974407ce2ae577bcdb097eda86ee2e4f10d90888afd06a6be
z6244f26902978091e6ec4effba8dd974413867315d3cd41faa7abec4041ffc0ac63a7c24290cdc
za21af966869df3a0918fff29fc2aebd56fac725d544658983ad0ddfd8e5312c1fa0ba2166f6167
z8b44c952b68191d4133e0f15473cc8d3af07ff35542425adbcf7ad61233d0514c6cdbd3abf9993
z750193fb86721e63f6a3f5b373130085709c6492e9da9437357b3c37ad1d88a2604c6a29e3bfd2
z41f084b968cf7afb896d550913357c11dea3d4ca9d6b24003f5c1a694b94877bd5c7f74c3f741c
z47b8e8312e977fe730369e90e0fe4e3a349508c0960dccb3484c92a67999570be31c5f2df316d0
zd3ec2115e6f41692e8531d730dc739dcd73cfa9c11a9a41401baf019cc5b24de7d5eb2bf58c061
zdb83c6de353bc01a194634cbdb0a67c4430589648c809eedd3edd11e87e94fea8057d8570c53e9
zd87bd89ea8aabbb95acd00aa4a32bcb0ad0b4c1da324f6fcd6678262acfadd3ff895b38a78e9a3
zad956a51028a9d1191628e05278e185a91ffedd3955871f0b1c1d5cf4d2636bfcd04776f916b8e
zd0edd78e7ab4370e1e74812d72e2e4c8375bf8e22894d69a7576bbcb677630eb014e1471d32ee0
zb1c7545e9ba9434d55ca980d0f171b8ba34929f7270d8711e0416be648e837d538b07307dbbd0a
za916b6a193c26512b3b37277b44e0ee3f3a87f41a8244cb9c82f82d6557889dd46458b1796325b
z65562df0b3f94e80a65b1c2f66c858e9c3406476238a2c128cb3d02fddeb39be7b5e508bcd150b
zd7eee31de6596bbffc316c1ce0f6c49a95724c6c43088f0b60fd3ad620fca3b050079c4796a278
z7a5eb881860cd8c04a27caf9872db9e4d60e3f2ef9ceeacba1723083b1afb888d127309036baf7
ze7e6944901b7c47f53d4795889c6637838d4bbf76d0b38359557bff0b602ad5922049f3dd86be3
z72af9f5f7d4fd218cc66ff21639eb57b47f319547b8b6eab7e5c4a5a6896a6ba94f36270c7afeb
z0b41b289c3389dc8b5fa17f98cd1b9a688a13b4d934cf982cf5b574d8ac300123c4670f6e042fd
za73142c8c08d24c2e7854d88c362a81c4cc255b9b6ae826422b08c4b716b0f9264069ce17b2633
z32bf131bb7849976ee103c9cb1cedc7bb517886b17505956d455b268a950259e293ae499f3b0ba
z459b5596f2ed60aa53cfd9b547bfd049441b00ca4377468873ec772729a6497904a2f8eb982037
z3477df1e51bffecdac202bec31b0f1e05969253487289aedf8a4e6054e6b02e920840006077416
z15bb29243e1071e53bc765d3f1b74ee2ab6651c944a8570c9942f80b1ac984411d21d2ba62e521
z2fd1c0201985f70912dbd58c4fddf1f075dde29b87e209f10514d9f31c76c0bf9d7135677bff15
z77aaaefa386b7eb563542dad25c77df4574b2b505fad65512c92f9e9e2c54bcb7ff8bb2f2a487e
z9ac1350c0d6882bd8a37253d69f246f023b102633478324e9a19c5c85cf812c6769a39db4136cb
zd1803305fef2639f19cbcebad3616378f91a97df0894d68c38ebbc55c10c00c19827d32dffbbbb
z5213db0dc66d7c383d9ef4df2bcb161bf1d2aacc25698bcb01a4cef2c7f8617f911162dec66ad6
z4f544ec329dde902e4ccb52111d06a410b403ccad233d159df53fee2c9c39107d4ca1691106a8c
zcbeab1a277385bfb343c238cf5e9c1a6d74d5e5413f2075cf58c366c7241ade267545db6edaf17
z303e5e7649e7d4e985cb3e72e8f94daf32248a1e0fd6272e7a42057632e38b2560ba89539a170f
zf41f38b20c5a877178e42a99909c3411e08dd76d852329f6cacadef4085b8238780932bb48dd6d
z4ef0c5f0a5c84a727627e6d915accd00be7eac9861b77fc8ea6648aef6516b3df8461bb9093794
zbb095c52b56f46c792725e3d826e6023213752deabb7a055bfdd58bb3d7f72828cdbde35d8306a
z9c17b00c8ae63ec76c33df0355b6bbd8d0673dda3587d70608be4b6eb2b024e0f912e7e6280614
zbfa882c999d816f6459235002c9ac296409d7e3c184b2e15ea68c58846b6e44434b536ac5fa8ef
zfa817ee9b470985fc1aa1300f1fa871e8d84eaaf2db55a49c1f9d39fcd6a8eaaca79ddea633e8d
z4b0036cf617b7f3fd88a781ccd99cfc0cbe3475e4ffbe5eac0d4ac6fda0c676fbcc82181bb099e
z284cfb7de362744480784acc50eaf4cd62b88c29f5557cf9cb7ddd85a8f1beb21e0863534e8d80
z2d8df7421724a563f28bec3a7e0068ea346c22334ccf2e1755bcc874d72777fb4189d4019c2bd3
zdcb5b94cec2290b58128d38d50192648b42eed32099b9e0f3e346442e22c90b15887d0490430c9
ze1541dab42376941b913078ebc662b105d2663287c7e672f406ee8cedb0688626d1845a274970f
z674d3a0d765e0c6e5cf40a2a07250319be0571b5deb9bd5ad224878ad755fb4bb2a46e554e0693
z3909682076967bec06cbc5e3e29bbb4ba6e471ef3815c043445155ae62946771d9115d7aab5443
z578f1080357c2ae67ebd67ea414d2e5125fcfa9301b5ac7b84fd45651540f1bc37cb1e78bf3ad1
zde96cd0ff9f18bd700e959b1a377352ec3471e5ed3c1c4bc5b56e810580782ae41cb11e978544f
z0c9a73b344ad1da573fcee7daf478966b554a2447da863c6e3c740bb89c68855d0e1fc3c91d4bc
z1c9949c23dc3a1e82a4218d44823a4cc3981574e5f8b9c0bb6d1350085adfcca646c65109980c9
zeaa7187c0bf3afca6a9c5f8ca400a367f6e944a6526b57caaa6cb617625b67300747a69a241e4f
z2ac53ec197f969bfb0df0776d08f0ad46ef628946bd66f2819448f454bc683b2a33c0d018315b1
z02a2d11378d8b7ddba86027b8c55b86678e05e69fd2907408e4c8c54469c42018fd73534f80cc5
z9709621b207251f9d372dcd9a1e8b513efd9f60c814578a5fe2b796f81cefffc8f158d7bd952a0
zf449567c0f2dea71417761c6e09428a42c11a9969b46f0e85b9a2647754e8ec23c0c252f046735
za0ddfbc8278a7c0e0f82b23d0f817456242befa6773c5a48c28f7b60e1985736c5ed444e26e8d1
zc407e84fba8d50babfcf2971db5fbd52fe4fcba93b9a6a3614244fe7386e356b4cb02fc29f989d
z7c20fa08d36724a8e152ab53f076356f0725bbbeccf80ccc0a46a36785204ce85db664cd0300e3
z0367a9da08cfeadcef95e177612f303baba04750e78f484e17fecf64e23452ad30ff370e97f7a3
zc9fae761f4deeef9a54399b2e2ba4a039bdbf4b0e4cdff0005519ce86131f8e23267635e557825
z8cadf8d95ecf2ceec26f61d0b7a209fb36f5281d94c9b778b92ab55f0e42605a5008f9ae7d570b
z05741ad00cb656c501234de87dfaf86a8be74d598f9a6cbc9a5340d63d130067b4b94096079d41
z128dcb69aeff8aecaca7b5dcaf472fe3fe4e7a7703f093b8cfbc8aa5d5bb68bdcf98b5ca6966ba
z6493830adb75b62ed94e87d6c8c6cd6ccdc011cc776e03942e9869cc29ba28991147b0b226ca7e
zb143b57a7cbb86149e38c358e6066ee5b34532b2438a69a0253888d541de8e1955bce022ea792e
z734be98ce1053739ef7b8ee65d30f542eaadbe3831b8a06dbaac5c3c2252615369de6078656034
z3e7423d04a479f3d61d7214d18659625bee3850f8e3068f64e0115c08017da67f0cf6c5db018a2
z93d7d1c292f55007f9874c6420c94c473509d48aefda2d1ab5b1e4735b537a3be61f269f9fb9bf
z80ae43709d38427821616df00eb0eb405287818946f08a8dc3436876064222bb1544fa9b91daf8
z6d713b42c67d4d06e82984d5ea29aafa738221c0f6cc2ba27ae0d2959b5abd81af0adb5cc486d7
z0843c62d2c8ee5b41c5f050cecc17fa64fa4245387ddb1d1d070b12a996659d57b5cf3bca423df
z7ca08a279754ae6fbd27adaed2be52be2bce8a5a3e69300ce285e004f247ba041f9fe42306a091
za803ad8622fc002aba6ecb03eee565b6f03d4cfd9ea57d88be0728127ec10fbd4303c6e83652f6
z889c4e29f917975f99dddc8d5973ad03dfa95a88acf3f9b6af6e03b7659a85aae03f91f34a6390
z7054e62676e1d82e530ed8815406171b092a53f1a374bf768e1f907de080ea3d76a210edc60e9f
zeb7e5e93a39aa74435494f159c7ff2852bf8ec52c5271982bfbd733ac1b1d896b5dc477c91326c
z840cb3aa12b00293428acce98ad8171131068e5a8e6f13b0aadded186167556b678428d0fa9efa
ze9fa0c3ff7dbeb7f490d17335190d9854b8b94ec3139b33f4f1e5899bad70e7b60ae3a9e4954b7
z70bd395f987d3a3692cdcf577c3b26c46015808aba9c2f4ead114cf56ae0ef47753ff7561fbf73
z72e4d2603ce892df6b26ee222074743b5724c5169e38730d98d8cf27f9272ed6255440c44dab90
zf5c0d92c48913722b41034e798a16bd48f1aefaea52633f92e81504a5df0d50f1c5fef25b24765
z6e1816ac3a96f8d2dad6fe8d2849f96a023f2fee83e23054e8036ada2f8845d318932d3ff700eb
z9180911a72aa84cd308ca86f81489125e9cd42433de72dd28864521f057257f3072fe1c0f955a2
zb126b2f461891ee27062383933924c45d7d16c107e4f3f5b7cff3a810f2ed3cc7c0d4c18c12b0a
z0290788d2edef08c3fef90ed398070799ac948d116a22c307f25f25023498bc31df6ff05571614
z09e78661488dbedb59c960926a2451bec0a2f5ad97d7e413bdfd395f725d452d0082c24996e884
zb25a5fd608f97b3f8234b3da1f1dc1ad774d54cd77480be6eecc6a8fdc194bc479b034d07e2965
z0778fe0e6f29016c28997e240e7399d1943eba0e3d51541acf70b98da2fc29dced8e45161a122a
zfd643bbf0949b2677cb6b3b05699f4d63c2792b69b8de9739f474c67b259b79deb70b5baa0366a
zb00190dec73b965f5fe44ccfc90dc3616485e1e6e7e703108a681764127bcfd40f7be52d868c84
zb075532d42f36f510d73408d7d470f4e41d68bd2b429b67a21c5f4683e9d5cd238e1edee7d93cd
z83861b614fe8bfa5f2c11b5c0150d79e233557d09ffacd16b23f45846267e14b6459f2f9e9ecf1
z53ff729e3dcb2cabfba0615aa5d6a797ce8ded6b3e82fd4de30125d0fc767bb72a8e3ebb9769eb
z9fe30dbbc3190382097ddba6f355acbde2fe5473b3283b312ec39364be2eac6c8edd283fd96e85
z3d39ebc1ed78e88a08f147ab713004dabfce8675faf84d6a807274737bf7fe2e8cf05ece9bb94a
z5bceb9722bb1c3f34fcf9c5f4e4207de89ec6a22c0cd5400b52da7fc4b050560c387846df44381
z5a5f040b3df0eb5cab8b3b7e5a80a26424b9a0b25aeb75096f0e3362e347bd19600d5bbb02fa07
z001db2141ff6fd1d14ef76641c2770d8c0cd15c4ed551d0930e4f524601573a8d5f3dd156398c5
zca4f832806950ae4fe56e6d62338dacc3fd22f3c4408f9f8b46b5fc82a9a165e18f47480d90181
zd75f6903789f622b7fb5a48b84fde965ccd5f68ae224d6a7793fd9c0b5c173e5b710cca44e6428
zc92f56e3479c91639f262e0043e5de326c270091b74db15a4110df6ba4d2d0dd9730cfe49d4f0b
z5deeba6278899a8a8e53f8b59ee9e0ce88f0292d84fdb8583d64f24282a3692bfafd6e3b0b0154
z25af34c9665da8f85700d89022e427ca4368d83fb613d3e9dbfec4b86706b789eff61fd33bdfae
zb6b065940ec8608e58892527f1e2f207f216a25185ea238414f5da396b0f237c70aebeeb27ced7
z4d88fd077b39b4e2e016dea72ab616e4789dc583bf523c803daa631cdfb4e7ef77fd3db776716a
zace6a4bc2191ff46009e775d39fcb07683e59af5f022e8046eba330281abc92f0a449e79d508ee
z31db5f1ac8f49945e6132a86d2c9a77b9d6a38dece44e8f679a3745ea2aa3917005e5f676ccdca
zf619fa7a7dec60f982c164e1fe4f9ed6e9e31e8e3e0e71f50ca86a851d220d0a55392910cdb806
z475e6f5f7ebdee4ea93e0598ab4798e1b178f091dca45758ec308dacd3e16bf1cc91e9c9e003c6
zfaea69af45965c4c3e45253ad8f893f19f247cf37cc3f1055404c656219ee92634892e8541ad1c
z2b5e72e008d776eaff3208ba24da59ce601c892e68dd66551f062209fff126dad049543f7ed363
ze9a09c332690b66977b0381538c663886dc06c217d81529ed6242e200b8412dfb4779d0bf555b0
za4489a6852dc49cfe48e82cd7aa1aab9d6ed0a46f318c32c1b4d3337cb74ccf85815f409cc83ff
z5ebb93b0fd2cb816b046ff2c3dfe06a995a35db49ff0d25eca368c74ca41ecfd75a1a1873f182d
z9c01e7b85b06c6d87da077abaadfcf453f221871aeaa402dcd2897e8ce67901935f4a3d011094c
z02997b43edfb0c091fdb1048b90a6d2e27935b616dcf8037baac55c05002955554b9f41d766152
z4996d8c6ba4a1f8284a50a6d77c627a3bf1406b6af21f4fc7e8fb92b059a6470c84988dfa224c1
zec6e013f5bc655acc10aa0948dc6e191ebb0e784b8861b5a78e92e4582c60c4d68ea12e910138d
z8621bba8c0ae600ebaca89f16e059f617d5ec98729514c1a6ac298a52bc73ac0563fff53486a6f
z024e290fd17d2aa7554db310aa96d4b8842996ea84f8c519d00ba71cca068ffb0f2a140c64eeb7
z766890300d1b8f099fa99feaa4dba2d64e3706c73fb55449e7962fa03634ab2e7c6f1e2bdd90a8
z67cac12905a75521f8ba2027fa97e6188777acc519b5a631aa2569a5b9e71d722cf09688c29098
z9d337f6e65696a9890cda57c7a788db82e39a38b5ac1f61338645c21329008e258beb3ccf9c8f0
zf551f660187b305a2fce2e6d6582d1a4c12a12c37b5f57781aa9303062eab6dd23c91adcffccb3
z35a3e316a7a68e9306ab12f30537c14fa06457a6c481a15c775d6e9dfa3b884e233a2aa54c0dba
za34e777e9d2412451b70e8f3d09cf1ba6ad34722b79a82c873e0885d8fa612652c3db3bb10c6ec
z08a0a56a789c78485a53908b65bd99982477f813b3b9c0c5b2074d79f960ce06a8baac086580a1
zfce2c1e4eed285ca14b2bf525c6f4018e51ff111b0f5e9a361361d1f48bd83b438c32847236600
zae6f5ee5dd8dcea496a9c81825bc58c203844db198153893fb0700e6b7a3ac1cd71f0c9eee0bcb
z64cbf09a732b17a50f7263251c8b13806ef9b16cb143d60a81a9f20a8d6741968b0bb99ccbda9e
z2bedea3be7535f016417f18d646c7a41173c35884841f0b31f8c9ad2aa91d91a966cac39167ec1
z4efbddffbca5ec26b84828f2cfe3012517bd903b385331a6fd942bad6fa5e067f139e8dceec73d
z93b48d28f99f65e40e93c4341e6965fdbf5d7be0a151b5f12335506b273bdbf33e85b5a88e793f
za341eacd556c445821d9b28ba014fdabfd64ba653e83ba01bd5492475849f156a616690cb50603
za63c49749358f87445bb9581433b1c006e6a4a277badd7fde639ffdbe1dd4df1a4aff683872c42
z7819341910fe6a1ead9f8c1984398642986b087ba122ddcc5cf2fef43c7ac03a57cccbcfbda124
zfb0e10ed45fcdfe4ae2c267b22c2a0ec78c424321efefa9acb973a5fea43410acc9d37bf491226
z71218545187b45650237788f08b6f33d89974d3b6e746b74097163d2951a4fa4e51bd519146226
ze8c7a3467da215924dd3f877fdf2af90a48e821daa874ac79522fb94fda6ffa8707d6208002ce3
z6cefdf41da0a89a3a6b87467b9235690a3bd3f781be94da354f105ac0b0bf7cd8bbbe48aeebb25
zb7ea83bfe92db7ca14c005c5b40d0ff7fd6cf09ed2c8b4d18ad6151c6286430e1e43ed9ae21533
z1bb164f60a4a9e7724d36102f117ce3dd6b835a60846d64752bb799ef17d5ce898db1586c0d7a2
z3ca3df76a9fe88a62f4a532ec78326b6f475c19d2f3f38896eaa776b609b5d0efd9f5722ea67e0
zb56e4846e94d3feda4a16bcb08933e6d72b6f2131768cd14e5f011e8daeae3faaab5af2f2ffc8e
z89287304206380fc011bab69095a2080d0dde177f53b33b7f849487aeed1e18cf6ba404ccdbe57
zaa54611d22789d2785dc8407e23e65a0139e5874cefe4d2071ad1002c32e9eb607782f58683740
zb9410b42cf9837b7165d06acbdb8958a9be083c8e190e5b8e228b04e441c03455fb0507a3b0ad1
z29789b46cde8717d3d940a64f37cc49a0ea781c8b46e0f53ef5853f073e6ecd347a6231657ddb2
z05645d07b4a7237e430d157450547b87f5143f01cc5cee987dfb60a24a1d5937ccb4447f0077c0
z9ed2dea4350ae49717456d284b3b7c37b1e7c3cda35885bf0e2c99c63627337ebf2212da1ce3f2
z1b364511344920c4c6893e179d9b3f1aaf0a81ae45ce1b60b566900be415b682d236ef90fda8ed
z78e3775875f50c14b1f3bc98508fb1779e97944ff26d17fd670f7098a14d04e563c62923527a20
z18429033f9b5e54e517f00db9c90f2ba9e565ecd3b4d022cda0571f4fff7f8a5dd5046e1709454
z74c9c7760954dde05644a4665eb760c5cbe0c620219873ba095e4b354ada31c6d41507c55f94f5
z1faa989256517a78bb1017f476be2b09c0b06e45bf3711255a77b9f0f6e41b34dc76a39cdcc1b2
ze1cd39404faf2c711275a9fb5bccce26b56175ccd6097673eef69edac6be0ca693df3aa3254be0
z52c80ac1027e886d946a78218230754b3ffeb2bbdad44fb224c85eed8cfd2c734232fe0919c7ac
z3c73deaf55c602a687c20b3d714014339296146383bafeb10cc99be56e8943da02bc352639c27f
z19b6f29753354e9e4c995fdc7e23a13c2e628ca6eacdbae291f15e3545b9101ee71b1c22fe4c96
z5e703ce08ed0bcbac7af4598d8c2cf0b1a4d4b9348ca99eeef4cdc2335a563197cc876ca861ff3
z9481997f23c5d08b09c310ef610499ec55528d5521db68719d45b9ef41e38163acbc93fe112d38
zc52a35595b4b1d94b8d5563876bab489898eb38278c9a8ae97ea436010f6e9360c46a8f6949270
z4c04907c4f1229c666d462515ba98dae4774f181eb6a9eeaa65a4dfab5c8dae34f8566c63c0448
zf14909a6db90a656bb8e6324aa443def556c659ba1b7c669b43d9e7192bea97251338dfffdf8e2
ze7623e674851d77607e7c3324798a3f8974e4273773a6c5b275c077d8cf6c8fd102ffe994ad2fa
z640769cf7ba8d834f63f0a98236ac9405e0bfab0eb25081c01000e86300ac64b211756be572276
z66f57fcc0269231dd673c90b1a342a5103eab1d4e14897d43deff47af4da5b7d08249abfaae9ff
z56ad2d950b74e18b69e8150aa940b96d9067ddd8cda7b229b6f1dd848db1a33b8f8e11d09c2378
z1676ea588d6ebf26f388a510e5ab3b559c4480d0aae48caaa7f95b021e7d5d97968c7c311bf555
z50adde9160c3a243af4f8309bc7efa530d4e5002153311a613c9d997275a93f96d7a98329b0a4e
z2d3facbd4e392f8c116eea6abf65995a20a1357cb8094bd8e8136f69e128fca2beee6ec7c37454
zeb6019c4da6a87065fd3447414ec7b300cd84cee070da5072569ac600feae9f52451db40a6766b
z6496205df86a1cd409e0b5ed387c9f71be22415e547f276e452594ae7ceb83094cebd106771333
z83ac2a600fd507b10fc205cd64ec86d73d08e968424a96ea0b40d9f26b7b80e06048d4d3a0c03e
z2f258f67b8be67ff69c2d1077dfbf7e1fba9130aaf9c778e29c6d99f9e43ba5bbd30d3af1b62f3
z2d5e06749c67f16dfcb6d2719cafb0ddcee81962037fe1b0a2fc1d41d66415683b3d2bca845530
z7b34962b8a766b625ea7f7e420d8a4e07062842022f9a02b81c00e091784278f8a8785728aa0cc
zaffe66eae994a993a2f569514f5e2ba4be7a6abb93f2c1082f1cec35992415822c8fa9a2fa1654
z2a96bc5e68f749f193a56bf7f6e35a5d2320b28bf4af37b6ed06c81fa2788a4b549020717c1ade
zfde894239088f64901e18482f840a08c28f635fd1c633cb937ba97379688484dc05ae8146808a9
z7d5b150a7b7df327bea7656c98a111eeea8fabd63eae5e626a648dc96948c6c1216a80795edc41
ze8595b9ffdf7c1ca2d09de24346aeea59a36057cef2b0958b57ae6cf1211cf9e77b4b7dde3348d
z352c89c7d081ff95afb893875aa246795d286a289fc7420a0d7869d72a739c70915b8849c63215
z045064baf1f3fa67453423181b4298f71038338df6d5e5be6c315e2c262a5cfbcfeeef977e0068
z956eef5ee31568b6aebddb47ca9c7f23270828aae45436d9a8f10ee237178527734e9990bcfda9
z04ebb6f8fdb49968ec6c64b78057c612cb8f925e7febc3c76bc4ccbf75ea6a30273c70c977bc93
zd2c6526853adefd20d765f6b3c9d2288824c96be212800889bcda2a701fdee1096132a90e49153
ze485de3f29ca8419566b02b35ed7d72c4e536ff374b102e3a6d82e264bcaf37686e0d8b45207a6
z16e206852c5eee7c03ea6d085d9c803e1f8e0afb0e5ef5ec03b7279045dae10978774c634bdfc5
zfbbf8404a9b34b0695e0865647f368fdd87b40a166c29ac16458919a3b4119abd5882681965653
za8919a51d531b2ca6dae445e0bb95c52182e71a6b77ff72ebd59aff95f5f5c435f6c77b52deb15
z2c8705279f71853036f1454133d89b89e14d322cfa794dd136b65ed2cc0c6e596aca0107855087
z4e8b2f533dceac4a7b3d699a8c073f6dee19dda7910561b508e54855ea015d9bae03fffc37d14a
z301051064b32d28532b8fe3297c094f8dbece8ed5649037f0f445273cce0ddb5bdf0e2fb155f7d
zaa94257a2fa593a9498692565548b996cf14a3eef3a30187cf16cebae5159f7dfd0f8b878ddbf4
zfcef9708251397d986abadcd6d943f8f4a68e5ad7568822d6e070e38308da57a485d6af81cff1c
z22bb8d5322917e08f5fbbf9636ef5b5b1aa85f95699a716a629bc17d37dc167671a58d9ea662e7
z71ee34fa5ef06cfa6f33c63b02a91107cc8451164e34aa82658aa25b8f6b1d5f03ea2d1f788813
z439d0abf91707fb4d6369a473adb953a51f0809d190ccc6fa4dfe533c4a2341bcb12422acfff60
z95126c1d69c08a772c79b50dd4fe07b3438b4a4a51acbddab0f162fa5f0d84a3c17c1cb0a1cb30
z1c42e2cd51ef86c6d0dfe1b67ff9a15b1603711b0853718487621be8216fe28ff5e2a2b4309a6f
z63748ca36e6f2f0e6f070228d1cc9a3dbf7095deaee39497562cbb942627d7d06e169acc5fef1e
z87a769dbdf814ab6336fe13e692349094c395467f8be609feb8dde1353512d2cfa0737d544ff9f
z27ed5718ec659f6b54512eb7c9e23fc13cb10d29a4461793b5c74cb9a5d86bd630f1b645f217ac
z243413cd5de115c9205b84ed482e58da3e0c86d69a329c4ec22fa4eea79d8320481900dc21ab1a
zd0377384cd086881bc518cb01807ba3906b4607e6c686def8966a5ce1d98e86cc156acb57978ee
z73a80130286b85b415c4eb40255a62093c56c8746c56cb19a24e3229f57ea6fd705983dd107817
z46d2fd8f20118a7ee2d0693d1aa7d941cb17c125755529df888146c8090f3c67a85a98088be39e
z5df78302183746726eed4832b9288116390fce5b40397f462124a6293272087170473cf1e9e02d
z22fa644090478e50103addc0652250071b4ee6c3b7c5e23b4cb02aff45cc7a9e5b616422978f05
z7540e3ff7f1320f61908eed9e887213461e2455847cffce5796cfe1d0d66cd530dc35d5312d10a
z766df70c21701b2e24921a216a7ea6eb67d335b0e2a9c034ba91349b81a23d366a9d0220ddc3bd
z0d441f3b27bed4a692e751358746bda4fce52e942663cf80261d155a6eecbc9a19a090d7d94253
z6800082c2caa69e5b1faf7d54fb16b5adf4bc0087e8c365be3ccd16f54f9a9939f3cb42c5b9467
zd35167c0a1221947300359a58c9bde2700b322d1c1f0031e5ec8d621fa3066112be761165904dc
z6df7cb81884d3d1d29691e9c9f88524751609382133ddd1106b74437b24f0eaf7673924914907e
z5edac5711f19c7cc6b258bdbc60ae9730c8f6ccc2e2638cfa8be0f49257ae74c70cdf3717bd78d
z9231a3384d5f5060e7332bf39c265d178a9d34ec7ce46466499974a834f6bfc0bc156090597757
z7a4229d12674d5247379de0628ad73157f963728064d2b566873a733aa6872ceab3170d2a4aa3a
z2ab502a2096f916119b776ca886a1c470a2faab727eb1b2a7cd82e8fbc23868825e3a48315da3e
zd43341d70597fe75bfd2aaae37bf03f62c3e52f5bdde7a4934bc8d509a8bcea3baef362e63d4bf
z7383d2d14089f6a3f137c0c59f03ec7d68b1e3bc086d5b234f0f5e5d37f9728d8fb50f246875b2
z0b92f952863f566d637edf79bf5a962e91cc076c7030269a7ac8be8fe9563cd1061229eb017784
zbc925b6f0b3e1905f5c02c4cc4f6b09de610abe3e2ec865553f5abd8b4b5c112fad09917b6bae1
zd5d9771b1f5b692ac48d4567e5908ec4de36361849f08bdf9d14280bcfb83dc3a3255942ec2b96
za19ad12a3ff83a63e22ad7863797d9787f676768e4450f62de2ce695dd60869ef090df977c2790
zb230f70d685304cb9386b6a3daf26d63b0fc266e04c175acbe68d77d52f05daa69a4271cf943b0
z1d1b3acacfac7c10e34215cce58eab89ec6012934f44f40a339586dbe7b0c7ec50e26c01117c8e
zaa56a9bbada7018558b35fc98f74623384879ddee21266edd1dea06b302c68a9c1cb3652087fe7
zfa971eb6031743f19cd2321b7333bc9a2294c83ce361b673fa6321c6c4eec6b3fef5e328f8922c
zb6e27ca6c350db682dad58e085d2d7c78a6a1dd83abb6d732ee9c4af38ebece32c407db9cd5e2b
z2cc3f627673bc228d33f347cc63b21a88e42bcb22bb7df08855ab597cd25bf08b03ed8732d574b
zcb0dce160eb2e98b903bfb78f446c88bed755371325fc45832ad74f90e0a439dd4ef8b3873e4a0
z4af379c8eb566a6834633e09566eb429a169ca6af6a30a11d5328b05ace91d3e1438d1321c46d2
z3bd4b103e3f4f93905a6901e5a0ca57f58f04c32c57c85f01be7099492c2ca391aa239c16fc2f3
z8d5be3002069e112839b9d389cd2648c2fa32e7b8b51d6152ec9c08a6a5d157e6b58ada8b35eb1
z04f70290430e57f16c8c30f5466e2859f063a79e8944fced96ddbd6de7b1bf8ea6111098916aa7
z54c0c584e660a5e7dddf7afd380a9be59655f9698adcf08dda0284b13f2af0213a0fd1377aa517
z01570ebfdd9bad9078405f38b7388181f46c6cd2d6a72896affaf1ddadf43b3eb1855c03b317f6
z0fa29eee1396cf6609d3c738cd01b198798c41e19bb26dc75b1c26c25e35ad4161ad6824308fdf
z84381d6e73fd71a95cd7e57eb78eb9ad53b2149180b4ae1ca06a133ab4e61bdeca1831c078a2f7
z24e61c02a1684a2a4c549eb7f81458f044a020e3c37e1a7d97f3012432f4fbbd3c74dfff61d205
z9cf877f484ce74a006567f7a90502f5dc77adad40389255f5f4be1aebf7a7139fef88aac783d30
z469cc8454c8cc79ec27213e1b16cb9ec34d1c56cec71f090a67d33c0ee68c8d4bd80f0ba5ac0d4
zbbe71bfba3775763b4c6ed2a29bdd38a633fc293d149e0dcf693618fa87a26b040217e5156da9f
z059e8d70ac5730ee44ed70a7d4f058d50b75bc8f8852ebfe8932dbb78ef5706aeb8ff6553bab71
z9f8d6728e99bdd0071b70da9410fe6bfb5dda557bda61cccac68a5c1d26104a501dca8418a4c53
zafef69373826b13ede22dc430368666e7b2750bdb0f4f3b146267f9d5c751271270aaf1be5d74a
z5066fbf4a99cdd860b01022c492defc825f4cf268471116e1b22d5f01a614137c799be1d33c9bf
z94d435c328e0ba2c909816c7d81dab3f1dc6109a9a11c42f277eabdd9b5d33eb9eebb360afd755
z2236eb84763165a89b2171b6b4edb8e40c3110e46f077963d0f7752bf1e025066049ea56291c47
z51e232b8f98e40a9c769c571937726c3ab4222217ed074a15732168d7ab786dc1d5a4966fe8237
zafa8ebf1c6a0ebfabeff96a2b8851d03e5e006bd5ae62f03fc89eb41abd45953d3daa521087074
z19de7665fd2b3ac9dc379829c51c6f796ca27049dfd80cb8a8d6b6a3a44a128e12fe05bf685646
zaf601321eb06a142320280d95c060a25a66e909ec26b76916209caf4b03de06415d4a4bbf6e047
z61b5195784c398af2f433ba525314bfb3f4bee9901df814211fcf59324ae7090672c489bac98f1
z13ce82ae23fedef0f72ba0299d65fd3a435bc0cfcb48aba2d84084ac9f2096102db64aad0f3d30
z5c88b46776f0d24e7fe9ed8dd37f3ffda1547ed3b0e391750c4d56d6e0a50dcd3ec815a5768c28
z1b3b3922c88cb05e3b01fb5b6f0fac9955db4d4fb2dfb8d4ac098a8562351ae81daf0f6d688d5f
zc83647a4a21c4f8c124a1e06ebcd103d1784ce1e785dc6ad219974c3f781f5f2beb4f205a0ab20
z6664b4643b8d12d5a8ddc37cee0cc11899180f81761d846c9977324870995cea76f55916182f6e
z2170f778545ab895ba3e5dde5b383eddb9dffa7858caa6e7b35ab5cc5699d4bc1d8f0f7e6c4540
z609df83659f001629a238cb51f90a373e0a7eb2bab3bcb2baad4ac13cc6dcdcb8638754771eaea
z37e5205a17e9535dc195e0ff02233c3d734a3006bc450c20d396b153b1a748411644753b9694ec
zf2a40e9bda0de04b68594321e88ec21b1ef79e69bc3857e9e2b111b4b381bbaf0cf2fc78324d4c
z20e7a6a53927fe8ea43c141990753838f90384850ec4cdc681e03c0c2fee9eaa7f875bcdec7bb9
zd3e6c18669d531c57236cd6a3c2efb1a1b53c1dd8c8ba2369f2f94a201ff4a391f6e5a36a7f07f
z1ae9b520b0ceea2f463d99dc1112803af0e879eade57dc5530b2002b5fdf3c0c0ef58d4048a706
z031eb9cd4401e9ffacd7d2881c3c78f3f14d73837a19392122bc1e2a3470c8a04621fa14f22575
zaad4eff686d0d190c7330a8865fc918ae1cc04c9b4144c1f6b35cf4d849f054a59cb6f3c0c76d5
za6555bc87be251f3689a9704dd9c1712e4211c13ce356c11cb4b21f92e89fbce04a1d1aa425aff
zaab0551fbc76b808cbaceba4fd8fab88b17ca0e28720682150c4ef93dcd6ba33d1ff0a5f12fbfa
zb1cd9ede2d06bcc57f0f738f1d6b77f106a3bd78c9240820fee134bf3f1d1053ca515350d1c7a7
zb077563efcd82e5617fb5157e06d0379445626f309cdc40ded61dbb1f178daca77369d8f97b071
z601f94d4226b97c364fcf3ad488c4248d445a0354d48e23f6425b691bd260c7ec85d73b8dcdc64
z48be59712127eb66881b2fafe97873f898ed532a89d29e87ea10d1d7dec0dcb5e904f622e1f91b
zdfe8ae9f4fe3d2ee5386e7907a3eb2cf99d12a019fab90c44a5af47f8ed0f6a9360a7292997761
za0ed600c307236ce2f020c503f42e0b8074dec01346b60ec45e76425eb6c4b6f7a951ad738c37c
za6ab2543945d7eacfdbf2a68311a992a37ba9559532d7d281bcad593123d28b944fcd0200da149
z523e7daff7dea3a606dfcfd9e872da1edf6fba1b94f0af6294b7f8d32ecb00dc6f18b38104951f
z93655eada586610aa0c764a9c2a4d6369f2ed95c6a926b30873b08772035f7c09efda20b2a98ba
z613c75c1d911bfe999ded471a11228bb91341cc56995222d4bd34f1f6abca9dc603f850f363e5c
z533236830528a7561c2ef4c11af5593000a8ba05f34d33d35fdd4d1a0ea74fbecbf0acb89e1f06
z9915edcc08016ff0898f95b2a670593481c68f4dfcc687fb32288805ebf71e17f61f3633193a93
z4eb78630501aceec10564cee4caad4ab331b0a1841af80d1040ee9842b20f5aba2e17645a57a32
ze3a6af2782edf97f5ab75db5b2ada17effb94aa28e3b943cea115493cc22aeaf6a8966f37d65d2
zedaf305d5bddc5fd0d9108b396530e5374a0353176bfe939012b11e929a4c6a5fb49f12b0db3f8
zb91286c2087cb6601dcd9d0bff7efb4ca3830c6283b6c9515be9311a8e3ab0c7a7acb6c53ce393
zd1b71eced1b2c92ab48aceb82652872b232dc4541aad24957923afef8aae370f83bd1dbb7fa903
z575889dadef1247ba96bc614e954730c7f5c9048cb68c513d74ebd858cd02d8988423897ab759b
z0be8b7d94d84e124f3bdf28810cac0490618263d1a7f60515bfd47cfa7fcb581f0ac9214b39e67
z2e1c55f04ebab4d6adcb9932eb725894b106965cb2543310a8fa256a910c1cabc3a04ae0cff863
zca77bc483c57bd545ca26cfdb6e5f0bea941972f25a7e51d49d2ef39520ce64e151066c2b591e2
z8cbf9495068de5593888286a3a03a7e5497330f3991311c72d63321796f9c0b5664a61dca750bf
z7cc7278c30ce617e35401b55681f519391aff027d3f53b908be55d8f11b5b1852ae5d0b6292952
zb020c8b0f605a0d4566adca2b1047bf06035ad3181fc24c1000e3f8b37693d5cbf456d15208ca0
z760d25dfc4a1cadc3428cb36f0cc36adc8290a1e599d4a57db7d303a84438b8a644385516eca7f
z5da2927fadaee61801dee9652a2e442da44abc989dd85c9585142965e6822303227b74234c75ee
z3923531726e23b9a4bbb8c254059924c0549ebed5b4c893d7f5559d8c944320ae35fc2de1bb352
z139c1604cb37c3885640302b103a9280ada0ee3d5b74cbbe8c0a0e9ace278c3604053b61c1714b
z3a4b8dd291c7744ac65725bedbba16bfa0b43b791890a9d8602c795e9b6a4277bc2d239bd271f9
zc2b99cbdca60afcf20220c282df87f3b1d7d9a94bc89aa5fe5bd984ea42bdba5619a59c5d04944
z75d76ea98f70de887fbcfaf8834e0d9efa8bef556d4177435c6d3f45323ed37122f235104070c4
z3104136ede405105ebc5d55aa70885d4fce91a5c993fca97ece4ca52fee474323a7d543be4b6df
z23bfa1d611f144076b997eca50edef8645ab25e5ab771b05054f462a96590d976518811d486db1
z01cf958aa4895f3948df72e667042badf4e56975a87faa6f1cd51383df488898777de60ccb1e77
z1877202b91a84dccc68ceb07cc594ff7d85b7f677571016fff0232db9429c5d9c0e5df71fc37e9
z7125806c0dc4d29661688f3ecb53df76e13aca905b033001a135221f2208e3c3422be94915999d
z6ca897ce514490582afbdf59ad2014b32d8ae1d6db73dca3181b6103ae18804ceb8c2a9a2f7bee
z58109482c4462d1c58e40f1d86cbb5da360ac50160b610386cbb44805b01d11bea643d44892586
z64a3a97baeda8daa1604abe7e0e568add4366cebcebd9f9b30069f69c33d15d175acce5dd420e8
z6e76fae5172905c3d2a8dd522119e103e20f8a12fcc3fbb3cd0164e7a6bcd7c96c1b4ac21a0cd3
ze5038e066e53bebd1096de6aa3477486be6f3850231979c4e4dd81f61ff0960e926ac5205c8625
ze3871693ccfa1668073754591dfc4f59209680a7fecd22a7c382959f945fc5ca50286829be79d1
zd57244b1e18ca3aa22e2fdd9382209786a1a9b56fb642f5c4142bffa2d2f7c23e9cbf19178155c
z4ef1dc6ff0f8b5165e0bf02e7720cce8d6f8ab8707a2e4f9be3cfdba81d3271c54392a2c8fa1d2
z49a1eae8691073625238e89073e4a3395fed7c00d9e6f6851d59f610d049312161bf13f059feb1
z53d65de6fce0737a861c12c04fff6aa0a4df76b20320982faefa07dc0bca5141719b4686ad8ff4
zd3399eff1ade9cb35c6ff87f9c02413d5280001670c1cc59e8d7cafeaa2262d047c06fe91beca6
z700b716e0fc940f5e3f09366dd21cee72e96ad15efce997e4cf50e01df785fd9bcf9326a8ea2c5
z437c9fdbbacd5be9d8ae96558ee1445535d3c632d5fb5538f1aa4f18f3258d83aa7e803015430b
za985a35bd0e825ca4e70b44688e3bc03b6ff1844a38f73ab7313f88a3516d7c258a9f3a53da9ad
z5efe8292b0b8b717a36baea45b5b726efcc13d511e8f8ab57423094c5bf4e950a07009a673181b
z0b670c7b0e1057d88d3dd5f156990a987a870cc7394e4d0142382eb505f3096489f5118a79e684
z658a69b949a27dd62c445ac7b8f62655f4b04993f59d4ea902e03ae022216031fb4829776bbc7f
zb96779bd840ebe17a34f02726f7c43dc03f4c88ddadf9604446eb40b886e366b3c31ab12ce4b2d
z77d6bbdf75c97365cdc475330da5a2ef0497f24cf7f3921bb406bdfd23927f7c363fc2f0d5af29
zcd528061c7f5f6662a52d8b94879d06c6ad4e545669cbe9d6ff6a211c34146f5756b5425476c11
zc1be42393dbd62df779274ac087d00f936d7c21615496b5e106c6d6d9a652fefdb31dab7940986
zec46ba8dcc1d84e16fe388ed65888bf9056575a8cf15003116c323a3c39c02fa74a9d339646bf9
z644e1bf246214544fbf89037be3b2c6b3350e17548bb02eb41ecdcad3202558509b48386a7635f
z3350b024fcfe8cad432ce8b225312cdc3771703657ab577652124036a917a1e6c86d91fddf36f9
z4650bc8f6ffb8d819d1bbe8114031964755e737435541624625c93e2e36fcefd425ed245d79311
z65e85f50c67710edf460f2124ccf09a74f05fee4deb177eb2ffd4fd10bc351fc80d8b4480675dc
z1405c69dd927ec9a85507b4098dd920621b1d689970db89c55642026a34afc548f0a766ce7d1f3
zd20dee7506770c12ac284fdbc6af44f5a6fd93c7623ff4af70e019227931ae804dd96aceac359a
z6f6ea197790e98e032d30a59d66c7f5ed99225519d57e4e6311f29270a3bb409b75f0cd9475e0b
z4e53b5046a5b20542662b38496f4f408bd273e012c300fef28bd678f4542d6d1cd32672d36009a
z5d41b212e145a3362e9e9d573d540c05cba593de7c669d4775a0dd66d50ec31e39cafce81a9ac7
z38fa812fd48564c32463ce170be09370c317e842547001f8c8fe186a72b8f95eb62ed0f21eb8ee
z46c1b43cb58853b95dcce59a1a2f73b04e15eddc423676ecdae28a8b72ab72f6e3468e745d5eee
zf25a839f963d9cb069b662f5da4b051703f8df4f40549f7e028734a52f9174d4bf000868871853
zc9ef45401e61ba39282f33b9dbc39f99ace4868cb8c3941d3419495331843459f9c1f3960359a7
z76e36d54e79406104c5974b1f76a794c44d9d3c0c1d09476c6e297fc3fae6b614eb48f587e3631
z477bbc7df263f8337a68166421ac5b66a08fc8cf965cb0235488e4b6d9b4f867ad318ea634e79b
zc091033ad8dd27f4d458c5c8a71b0024448d2d26b4cc5d5bd8677b101bd3aa9b9d8538c4edd3f1
zf9e684cbf3d1a19c78801f21d665c057c9901cc30ae42d9b6ad94b10f9b21f948a6e03f54df1c6
z7788967797c2a209604d99911e90b18cfa042a8bf5dbb5a8b32c30ad78295b877124c125d78722
zeddedc12f72ecf3b008105d27ca0c1039aebcc0e2fc763d7a45a7fd542e6a2f3b73e65a6d8c673
zfe807d8266e42cbf6a9186e9cb0daf04cab8b3774df2501bf7961dc9f798df9ab24d99f542c4b3
z42b34df4929295e47c02317c75b8d0d278a9d295dc7a6220d5a1b5f31f39d7d2eb7481465236e7
z775654302c179eae3373c44c3c7138f2b93e55549acd98d9056404cca575537b94474ed42c7485
z903d9812f6fdac2f8d30ab366e4d015d38ee6c6d3872695348d38f66f12a866fd5173c4b814424
z0830240d1de5f2fda909f8bf8c22d9098605d0678d7ad00133fa902f586489eb9b64026e21f180
z00663fe3969bb184146ba5d217d9b512a10d43ca9e242fa687b2c04987e4b372d887c9c86adabd
z443a32cc8122505b5aee387c645dca5d172f357d8873067379fcffea0d6a125c8d6ac4f146c86b
z05da608f4a256cbcb9c9299b1a2efbdc03fb542645f3f9187d319fa1175a477b21c22cf1b308ae
z02ba3e0ddf626f303aaf17729c0d3e4b5d6c3ef1d22a7e2465e7f2985efb5923519ddcbff45a06
z914a629a01bc7909a5ddf137badd8f9fc3ca23832f37bf4b2281e43b2e2f868c9dc83b598d2ac4
z98f1300d221477181fa8669c45b8a6697dab935edadf778de91e1338e1be65faffc56f4df7a7c7
z758c5fb983701e43dea407b9bcc531c442cdabf9a264631316ea841a3358389911df047a7115fb
zf6658af34a2ef1fa520e72a5ed5372a513617ef8bb930773c238c9437342e0c43b75d0c4b6fa5c
z392f9107cd626949fdf179a7121976064f6ef182875fda40d8ab123f4701ab245649be69b33b31
z603eeb202ca8b90a764850b5848ab4af69ac85c9b9c2dc0647c07b7f6a80bb1096172c322b13cd
z222e9b5798e7834a394f448cfc84426b714b475a4d27f280ba63551809a7fa7bbf64f652558422
zea25562cb2b9c4e37bede7ae6b2d90a5cfa991a859bfd7361a6b0fd4db9798ed56003627718071
z8fa1a0bd7950d85d095655883bbfce68b59ee3e412f4d8dd156ce70638d68a1322b1fbca0d49eb
zd65b1e993804a9041df1dc2e52b9fcf8c6cee42b9d0fbfa56e91f96d06e7905792c56d79a34c11
z04c97fa38aac3c526b280b843c1039efbebc0d2e317ea747500f7b231ebb3636dae24ca9c2a749
zd37ffe584763daec99a57003cace2f2bf748380d7122a2456779be7b78610da1955711afae5d19
z3498a677f8682d907413dc5d6b60e3be6f916f10bdd3a404fc62b7049dc34e7539f859ce01f1ac
z15f087a217a1b0bb5f7609abfb774278527821229f32cea80ab1881014a99cd6a2861e5cc5a44e
zf9017e0a3cc0514888a885f7d8141e95c8c69b072ab019a9abc9ed5ec93dbe96dee77dcfd140c1
z67605d5c72a1e408b2ee86ff201cee32e7c20c24872e1373a46b541aa835d8e034e3baffac6a82
z927e890c39d0c6b65d957962649e23f9134779bd67cfeba8832921d80dd44b14237b337d9abe3c
z8f3adc0fa46e5192a9bf5a63ac687f8ddb8f409f4b65786a4b475b2662ec8f954f9dca104d7eb2
z9462c0890732b47e6ed51eec24effb618ad8444af5c8ca2880313a4476b4e2f05d8a17d73fd12e
z5b9c9ddfa9be1fc097747f32c3b818b196271a5509e79d532baea65e5c2abc0dd55a7b77f20c99
z5fc95f8197b9f862152e3da0374a8b635ac3d6a961ae9e934186ee072c67cc74050df418cac9fe
zcdbbfb219388c56c1853e4c80768492e1a55c6b863cd64ee6720bef9b29a1aa4c3ce1667c45837
z0344645082d2c560aa9840bb030e6b19a8edc396daf38f89a9c1225a95e812b6850a2a36c738b7
z2f72d19cf06dd5203cd20a995091bfa5f5f16169f918c2b6c65dc8a27d1c24119f136aa98d9a47
zd4743d53a4d948d0e657dca07c64a8e6b23b9cc10fc4f1991856a9a7171209bffee64f329b09c9
zb28442e46f5c4b4d91625d20ddd859ad44c5375a4d0bb2bcc6824af655bfffd41a75fa4e7862d9
z759522fac46f719718cb6bd284e1783db88e528627a6a7a3aab43c191a21e0655a0dba3307ed46
z70220d2aba6db200fd16b9c5b9811d25158fe29f7f0ac28bd4961fcafa9dd7180265a1eb65b6e3
zbf3aacce0f0c3fa9375ed79deb97f912cc5800e44a6cdcf4098c6417c09692497d6574ca3f766d
z2f3d474e0e26ad71d8287f40236826feaccfb43a8021504367def04cc0539291141ebe4ffa39bd
zc014b81ee041df180a0abe201384c29e4985f819e3433370f6c63849a237a4967b7042ed718b6b
zcbf2c6484f589ada0cba6ff02ad0c1c08ac0b7d6f62e106b96863c4534416955ad6b7bc6ec103d
z4cb6ffeeff883b655dff071764ff8ab8d0415a128636e97915eec5462718729c95f6e73a66cfa0
z31c53ef6d805cf2efd6c6fccf8ab4d7849b68dac2235f061c7399ac0885c1cd4cf5343235ece6c
z056cc0e4c3c5e36aec127efa386dbb136f5dab6699e2da824a3c95988bb9fc3f8db73f46cac782
zb4ba6b276281b8b9d6613c391c40d6774512cca6a4788794ad32383b46d3ba5b4f64fc1547d691
z22de6125e7a7e36f4d61a0dfc926632939de21c37b976ffcc03c31b18031bbef8c5d75b51ae1db
z9cc67fa48e7938520df59ba2cd210c7a7619b7ddded21e39734bab842533cc4443ee91d633b5d8
zd0bf7487126acaab20f7045806358bdc7c7acc77764c94fdcea678bc9f37cad6ca2d29342a4a24
z041a427ef1219a916e8806d9acc92ed36d2b6a43c6f2a6d06318c50e87e13b98ccb8258deb05ea
z2fe61280ea964a9a5a326132b1cb0406d6e4f0d7e82ce8ae221195d379564d50164fba83ad3a8a
z5b67c7415092325d98a3be80a429dcd4634635c4205816ac717907854121831c5412c207a8122a
zc087c38f0c2e4a3bf4fb2d4f51ed9e075f13a04195104bf496b24bb9899f15da5b377f95f41ebb
zbb782868aa1c16dc2bfc9243dc3354ff87194ff2db4ad158c238d12d95826ea0aaa52456d38bb6
z964c8c6d658fa25f265dfe00c8c2d9d3ace69816f72cae24f3e4abe65e7528d6f6ee20ce8803a8
zbf9a3c637046941845201cd76bb2e92bbf901daeb83597197ca3395becae1dbf41e8083c457afb
z287ee998661f686832f3aa852e832ba4cad15b0b41b860094167ced8ab15cb2af075db3e63d8de
z2c5568a63c02fa08313b92fe1a6ef4c73909a9d48de0861f20ee62d95d7770536c8e739460c0fa
zdb4314c7c70441a282e9947fcbe18d629be38fa9512c795a073356681ed2f012f0fe769ab70e2b
z750a74d58aace3431a78f8c3228d37199190365cd2e3bf3005b0e30bcbb1a9340fe679ac189f58
zae111022ffb5ed17534aef44f6e45c2835a70d61cc3465589797905822ca9f2c0c19604de7cfa7
z3027bdb3bbf87691cb7ba8845d8729571a68204cafda0e65f8f127d7082bf1c82c3747ba024d69
z8c86b336ca6aba82383c0245f39de7f65ad75704a2130e36c3eab4835304d32a2b960d735a4661
z2ac084f31f1ea45ad2bc84d7e1731c576e9098154357a7b9e5cbcf249337fb718b7cc61d14e5af
z0ee4c87aba1bffa03e897d7a3022d2903422a3097a66adb73929478ac4d7af590ef1ada91c857d
z020f1337ae49e0eca36f20aba5592a34efb7581a22c4f9b082333e1a6676a3838b324d6459d86f
z1c603556dfc2964ef611b53adb472149b22509f53acbc8df5497d7c477b06fb9b2fead7734683a
ze0e516be08ce34674dcbe655166641b75c94e033b08aef3b1037bb40d7fdfd82ea01efa25afe6b
z4f224f636dfee3d1aa1b81a6e4bef762e3ea046e64ca626514e174570c4bb73784572f79f40c3a
zc08294b6bc47822dd7f677f21c27a90aa1d4b278bc1316609552a06dd6138730e1ff39f1ecba8f
z4b8d2b275cfbcd17e49dc9031f9b2a39ff1ce763e5f11b1d9e4f9df7d3a5720a94833e3af940e4
zade184e6a9e6f38d2b08c61f2dc6b9933c68b3846607a6b90efc5eda9020bda86b6a19a7c470a5
z9b662f9eee9718e8a378b63d59ff8ba5626f6e7e41d3c821c9c9f5e565efa8d8fd4d71d4f2a7c5
z6d5076aaf85560d788f6b94be623c36689c1373654c604261ac916d9e83ea50edba8f72974a3e7
z04a4e981e3965321c35428e23d88fbd79b58ad99303a8f4677706470822ca64323513b2e9eae5c
z9621e990c3870d8bac0ec82a8ed22f97c1eae36fd22d74a037ad7ca9493330230704414f5917a5
z7f884af2b07bc8ebe8f2006078a8ab006ab9e6f83addfcebe5bd2c46a836f5bd9ce83e214fa547
ze95fd660b553f549216d842e2ff9433c87d36ef62c9f72c822cb2e860540bea1286048e9030f95
z424bbd30dde8541103bb7ae58b308f5433d7830b1e8b9a943703eb5bac3159c1e11d7999bbea3d
zb290d0e36c29054a1e45bc7bea44dd4e4d44535dbf56ebe3330d7e25030259cdd9cf10aba06169
zf7dfeea07ca989e02e63741be4474c639fc552daebd2fd190f224f988eeb06cabe10a95ac5868c
z80e4b7add6e1a9af4cd121e389a25d49d6c5e6eae3dcafe806ac9f3445ce1331c1404d42bdd852
ze0e4c02dadd0d74ae94bb7eb212d5b6f66886e11ff68e8dd6e401a537c35ad4d60e1f6bf7880fa
z38f280da61b050465d7e2c4690c6896d0d45305a0619c3b68910549dc6825a1a4f895229fa7ff3
z2ad3d9bd970d631f6f1cd20130ec799b9d3e3dea2e717c83a4e5ae15f592911fd64267e5943766
zb83b52700db37d4801661494f6ecdddc58dd9baf92c3c33de8c90796e05015eaa61852a5fa9c6d
za46d354da3dbd48580cfd6f509e9028811c588fc3ecf585d28a68f12dd19d3d62ee59a29ea0a3a
z75f658f8caaafcced80d73b31cd5e09811e5dafecab2ffa9a7cc6e885aea53641076d6685cb9c5
z2f629610c7b6202107a7f0c5318dbde41d7ed7617b2dcb9e5de7c315aff47a370a3b6f0c0ab5a5
z543231774525f3cea08dcf488af36c84d84b2a7cbdf44fe121e5afdaccc1d89cc376638d104018
z5359be5e4de34b9ff249bafcd6c387da30fb7a7e6c5da91b03234a10ea685ac92130f0df816fb3
z264021eeecb2a0a3ac28afb3ff250444dab73171fcd30663e62f830f960bf160ed1ed8ba5e6c64
z2629b5af541a5561582e4542ba0dc8d8fef0e7b156499b5a854e7f0b231c4c1583dd8759d02981
zcb8bf265906c20cdad7045e1360b22b9c24058c296d9e40a049d2ed02c8d8faa22a16a16c9c370
zee32ef4bfcdc9a5cf81b821a1032b379957a3b0a4aefbb74ba908c6b528c6e9d431c2a8116e5d6
za56a8cb2df502cbc0a663204f71c1436108bbc8cc52bf96f3bc612a43ad0bb0ba97cd38fb0d091
za8c54b318dc2e25998beec9c2d6805840f7a643da8343f4b1714d4f1d643ff3e3cd281d3301087
ze3662a8dcf49d3f2ba2536d1e9d580fc15b03bbd949a14c38d94a661fef4b30d368c6a24016cbd
z1113e0c98f9461218d943a6ac2d5a7b7768e813cc50a830adf70c8ec2a6dd782369e7e8ef259ed
z9083399a132c11876226092b53a39f4853b72783ae4e4109d8a6eb4658cdd5e43f90432a9d4c72
zc875cf6d4ce0d74c581705753e4a0b8c808b3e7e6df7bf29c0aa7079b98122d67678dac69033fd
zf29404a1f86f7df975a3fe7f591d0f6abf2c41a75e64965ba946fa3da9966a1ddc30dd6a5f1fb6
z1347c85a3e7eb5f920531a1f0034a38ae7e2d708c6b7fadc143bc13f0e703b9593c66dbab92eee
zc024802a3323579d693a66954a6504b1c1ebab9a8e7183374a40506d7fae7a84be754de1b60773
z02cad4b67aa52138b4c99d1e47688262dad42bf4c75052441ffc792901f6219a7390d3f71819e9
z367571314d1cb01c310b485777f0f0bda530954c8710bb79c01be50a11c6becd7b64c5e7ea794a
z134ea44546948da4d78baca08b74c88e6eceb05b2bf20aadd5c6fdb2afa246f5ab77321c401f5d
z22f7ce8384eda2807068a326a4c2f16214c71fb6189d8f035a6b77511873a73c93dc13fb53d250
z38b8abfcc40189c81838a3458479702fa0e683d9f833ad70ae9dbc859de2b9107c10a7c873ed22
z1a1c89970df190e2a260a7f27ee617c7a65c441e4b220181f2fc26cce10c90342fd17cc478fb68
z0439496665869bfa9a562d676d9a8aeb6bfa43aefa8c6db36ed03d54a25dd58f445aed0ddd088c
z8cf5e8a280411f3751162605e002085ab4c09dcb0db923fdd5b9c826c82894de47dc83f4a69879
za978ba75559eb7eebe1b9a1a5ef3a7a32d8a9ed0656d0084f836091ee2cc88cca1fe109ca1cb48
z4a62176ebf2d1afa4c5a867b624410bcd36720e3611e95431174765f7eb72ab3e5118375510e89
zba9ba66502fa507b8bbf884e9da7742ae02c0a1d22c4ec8c23d8c83130d289024bc4db1534b7df
z5ee29c667ea2468d86a3d67c0d019fe7d8b90c29331d726c56427bd35e23872784795c7cfa3211
z4313f5dfd93f9267d6fb88d780725cc35654014c096fb602e13ee73aa58205a11f99ccfdc3a1dd
zd1c2565deeef67852abbd1861607fcb7e87c2fc3b8068602fb71881eb3fdd7bddd870757bd89a8
zba2fdf68104cab55a46b2a100792f28791a338fb9c301e359c908083a91fc482134e883b1b930d
za4d902a8fe39ad7c2427573b47199589f2f318af6e1f7715c01d680953e6fbeb8c3a815a9efeee
z778e9273827be90668d662cc242cffbc9b2618ef22de0539ee6c71f9d3ed0aea9e5ff4bfa12c05
z1b6301f5d18e8709a19fc1d829b9c340211bef52a8ff26458b4ad2f5e49e7f63abaa524faef5fa
zfeff620933730c25b500dac33b5381a06cbac11518b6393980e9751ce7a9fc8006ffb5ea668f40
z26d82dd1f6b75edf2d87fe2056e9b97a4f87ddd40c592ed201a663fded93acc1e90bed634219f7
zf03525e42db8c11e7538bde649bdfb2be93b944741ed1fce96f8cedea3d2c8c9a299b24ee669d4
zd21bbee7b5e60b24ed776c8ea45ccf2e30c76607d610eb1bbe19a1de658614dde678c4ba8289ec
z199b34c86ebe98fcde4ca739598785f11fe19d310deb3f9f8ecea650ff9f479bc7ca67cd8945f2
z6400345dcf92120de53843fc36a84c0c8ed221f0495bd29c9882879926e03375eabaa68d7a051e
zb49872f33a6b7aaf09ffc9b877e47ad3856bdc8d0decafe90d6a746322e06dfe959d6083f13f90
zbf563f9fb0cd0ba234df6170f0d24eec78df096d4469df371b5f277c8deab546ac937e9b05d763
z3dcb1176367219d70806e8fb9f153dd55bbdca25a718a409275912719ee48a7cd0fb88fa6fbeb7
z492b2518de2a4fdff95932ce82f5478a2ed17bf6e1a9e4a09e9ebdd83155a3ff8a3d57421703b8
zd7c3ebe74ad35437fc836fe85a1ebee893a2243e779ea013f87d60c30a3bb5304463d5c84bf687
zaba06fc48a995298c677250f095202d22c4facc1a07e39931f144fa800a63fbb104c1d5caefc62
z601c2dd0e9c6e9f9f08d0191a36539f20202238d64ba084ae4c3d4470de7b5c9e192d4e3b69f79
z47eb504f23e0e52ae8df2e37d2f312b3d3136489c4a6bfddafc22aeb1e95143e7ad6368a44f374
z16f937e8e38a366f612140b72a94e54a77b131750ba49a9c6fa58b8af96b0cf43a06338ff8b063
za462fdaa3531e08a51c957f387f12d0789947239d421a5b375c6ea04a78f0205a7a41c215ceff7
z0abe3d682b56c82fcf08cffb65172b748c517fe70c00fa6d0031a9cac2dccddca23e069502497a
zb36764bc8fcdca3aa7fdbde57adc76b2972b58e5e568cdcc14d5fcf91c497a65b344d9c57dc70d
z32cca19bb338e97e330a3648e3e2d5b390fc27476e1804a4b828743ec603f41c8290c106c7d52b
zb48d5c00b5c043a520f7fd8f14ac541f47d2466c8d52922938c71377799489004b2bc9a085a27c
zbdbb77b74652d998523c4de81b848f8888a8df6b51315cbeee3a621c10d4267ca27bdaa156bf43
z60091ba5cb454bba631a57b033fcd98f01e64a8c69722aa3dc854a1a3b45c8d650626045228da9
zf50b135664ea442ada027215762b07d96ede467fd1e605ceffe1ad42d8be625257cf69792756a8
za36ca07ff3fdd7fdfd49b275f8ddb4b0d4a32a56b86e2d84ee1da131db9ab6db1f0c939cd9e470
z453a59152c6198ade866e8c5b753d28f37a52c49a3bcb9915d0500c49719ea6d01713fe065848e
zc9864ab3c6a28780bb16033f3ab2a360e7fd09d2f7377387011133ee04d994c0d3e68894e81f3a
z084184dd11542a114953a6870246d731dcdf71b4f511063eb5e61206a295fa5520cbce2fc5fd12
zf2604349a6331c6b36dbd011bb5aa21fd2be868c0beb5f63b6be7c99387bedcbc510c828ba850c
z63631ee04cfed652b1928fb4b939ee49bc965d945e6421164e795904e82ec64708a9f2d317ae6d
z9ddacff8a90b263f0aa10732a26853828d756bf1c6b581ee366ca8e64df988ab12420d9c1c7066
z9e2708486c0707de485b3a77ee483a70dc510f4cd69a4c531d23a37c2795cb9b5f1a27b9cd0265
z77f7a2921e1c72f97cdb6004b5885774b9a11d6ad1355238d65ef266853820728a62e18daa5e4b
z20db95ac89a62191cdc24ba50af2cd450f564330be3596ffb66174726d0902adb3cb04741f588b
zf3c99ce44cdfb6c44d3671924dd51931778efd9cd3cf3690369ef6bf00a9a923638140e5372a30
z13942d304004666d619a03b9ac4667f41cbe21976d0439c15e65506e7062923bc2d9c1dc4d3e9d
zfa9772fe282e9ed997cdd8b7350ae188cd69c48b1ca56df87300eedadcaede809d6698d469d0b0
za2f5c800d2fb69444ffbefebc8589eb4f40d0acdc1dd0523d8394f8b6dab302e5b0cb0959177b4
zc85eaf6d90fc999ecc7151728ad7137e14e0e4180754a1b6fc6dbf3e670a2698ee734d8af6de23
z40423d6b7bab938de13dbcec4f832f84c3d01cb2424b19b0369ba5615a504abbda92284f3c1996
z1a05001ead32577d2ba646594c3e7e33fc1332a7838e12c112cb2d0a5359d439c1e49b4995bd22
zb828d48291e3380eb752371fcaf0cabe5e337df7cec7717c18f9fbcf5145d62a903c7d41c04c93
z472bcfda05155fe5605b32bdaab3b24cfb768877295c0d98b1393ef7d1aadb8695e66a6bdb181b
zbb9065b1c1a4717548a231fccbd88a089351f74ec8e2a8f11a0f9433153a7058a6bc5f59bcb036
z1006232e7b3b612eaab3da29fd400078c5cbddfcb0dd4b309a43441be6dad97ce2d0f6bb6cdf44
z6d9d0cffc922bc29b1b61a0d643d434d600b5b57e910c4c5d5d282ca70148d9586258123733a10
z24e44b52e436321230d2af3cf779e2345293e58cd1a3fb8872aea1cb4022e6bed979a1e9b086cb
z58976d126ba1e1da42be7f7607ff27ea83a1fa69de5a97c30c9a8d1b53d71c520a3c531593d051
z3a22f46397b0bb4bebd196790571a26c6c56651a24c6f4ea23fec3cb87ab539a4dd7ba1eb34ac3
za47adc277031cb6cd7c564bf9f93aae23dd19a1fd940d04bf3963a34006acd6ba48003a7e38195
z7d0dec523e51ed3688006e40c2afa1a6bc5b5bbffa0721262bbcafba5df85d3303eb2dbcd44607
zb7ece7c00ca54add587214d3cfee50bd9f01752078d715f4bf44de9d895dc65df79b08478113c3
z5255ab231ec34a2570f9f384d3cad299b7ae27ad4026bd60f3ae140e4650d72783ce21b5899341
z142961ec4087d90689909aa9468d45fed31a84f10d9396402b3cddf680b92e15e1f5ab44351304
z657b3188a7ec52c28d0e210de27e3726dd6b3fb5b181a9fec34fd3b9f1e62a27469b58103059af
z2c6a8d5136a10957f90849294d0177eb1a0d78eb57e89fec048f8e70aff78fbfadfeaa687d16fc
z6f12ba7586901aa5867dad05ab41a5a80a8ca92f836bade57f1bee67288b20127214827ea0cce2
z729b9a86a594fd0ed51bf029f72c857781f9535386b53e647fee252a35e5f4dc988444a13a275b
z8f5b20e5cb1395e47910e5bb3c9313d1cad885fa42a437ee93dd16d83ba89dfb6bd14933479e4c
z2316a83c277a2e4ad180c1383987ea872c4d767e5eebe553c2afe8d77259520951d990c7c47d0d
z9d83c52b208fe142e7ecd8bf8a3ad1dde79f015b62505f6a5a22be618aa90cd729c2ab0cac293e
z103182ac3990e9d5a00b3b362ba7c6de70ce06a6f11757370d448e72109d8bca11c23b498b1308
z9c9217f626c9a9d328b8c154531f1327241ff7e51eaa0d44aeba31a757a07ecb9719490789f214
z7a758ac72de1bbeec04e95205fe0a4961f536d68c8fed6784eec4495112e7c487132acd3b4f7e7
z29a3ff314d4e8d570687039b035908949ec4d78521cc3f1cee46484ca6a429768b77fab7fc3f9f
z8cf30e4a38a5b14d8a8feadd1ccc9b68d3f1b634e6ca44fd4a954dc0c6dee3f05ecd3ee3b94e49
zde9a0d2a1e428303d8d82b7284f074f4e3605d426247dc577fc4fd62c20baaedf9ca2c2e94887a
z17e52bce65e8c8fd7ceb5fc1c9f0021c4be411a18ab611192248f731314f5ed60a07726ae215f6
z2a15838d01d7c95f854887bdcca7c56909651b3fe6047df280202c3fcd49c22853c38544280bad
zbb0b8aa04905b3b168544ae7e21549d4c59aada287cea87b7a894a1cd1dfbb5ab939197591d5fb
zda1c464479bd0037cac41cbc6a093a029385e305e0d39af28e31597e0600be7cefa40480dd921d
z5a8ecdd6fda68acd024a3c7136195bbb97e663895989c8f299ca94388980674855d470af24c438
z9e671db890a3df442bbc29ad08db49e875a7938f6d1816001a2ecaa1c9e7f50046dc46cb3dc110
zf156949363fba950ed96516f607cac86fe73b6b78eb00ec0813d975a1400cf647733bdaa59d77b
z0e6a1cd4bbd3e77f0f0a248d13952d3b1154309d548cab412ae7845bd5e4a9d2f69c844873b6d1
z85cc797c73c06f909e16f20ad18d5e76ca28b32918a32f9c451e0ea838b63cf1ae970c69e085aa
zbb80092af2de818f0683cd9389bacf5143619913a183788a5367744cd04744fadfec23307ff353
zfc787be2095d49102af61c6583cc8fea46ba408d55f135a0e35815209943ed25a3d8797d3c6df8
ze2556a534d398150b1cda62643f90ecdd9cbd4f4593ec3669513afd1494f9a06c9a2236462e7c8
z4a2b6399f71d907a6a24e08feffd9b2b078b11c6bc162fbb8f50f0903bea1abdb223f7e28f4542
z3399642a683bbf53e7cac2fc587fd197b85234144f89f94472e408b6675253c7efb9bf06f2cdf6
zedf9ed508a60bfef9f605fbc9d2a2c546ef0cb5382f82cf0a9c20d31d9bdc6cf4e95aa211512ef
z1fb5c35929062a3afcb217525592059e9a3f3fd0917a525568e37e05e16cf92bb741c3e57d710d
z48844466000ef856168bb99b6e2a7e8f9b58fbb5fa993d7b17c2675479c130de94850110e2f7fb
zbdb9dcfff763b7c89525c85cde830e9f212784e80d3ff6996d2b377de6798aa695630f55bf9917
z6b71d8ad23d98a3a433c6efb019688e2c82e79cf849d6a6ed4e7fb6aab5c7e45aa8b5eeae7c6ba
zd45e21acd32ad2d5088f114991ac279690a3693f75a006571bbc257fa6255685f64c9803b87caa
zc5ac9b7dee20305e42a5c97cd4919270fbb24e375647749ab7d0532e1322a7a456a5250a1a2292
z881327864ac8edfad134af7533b3a02254fd47e4c1c5049814f8915dce24ca0b6fe7f5f26e2997
z7dc05192b873fc0a16458dd88dcaa0b510582d81b79965dae1d94fe317dbc15fa6de69b4fab4a0
z0ee9166ead9ea41be7410ced18e67b0aca6bb402868d55648bfc4f9ddf24df54a8bbb9dba9ab84
za54b39c988e920c9916b5a46ad768f28b8170fc64d889fe9f20898ed6ae4202d3bd53c5ce8416a
z07264424b937f6249d80ebaf4b8195323f5adf7fed7e3f6f4fac9a20b57d6ad71a02c87134b6ec
z7312fe99410e9dbe1b7cc0d1ef6001786f2e0c2f99a5e4d8cadccb9a88c9931d0a30856b0413e4
zb02be4c481c597e4d5e390d7d3e2862d529c4d93d9704ad65d790fcb5f93e36ed41d2f100b97d7
z47a0f5a235ba7e36a98273582263f9af2b8b56d2f3efabaf1520a01a55259b09881208aa64584b
z182d48f32da08d63f9f38ffa2ae875f176c02789109bc5ebaefc49ba224d888ee2268fa7159911
z021389bcac32ba6c82c8b5144865ffc48e2c4e2237b4038a14f36673259489f8451eb509b5cf0e
z7d63f9037f0340d6603323c5c689559dbb9af52e1550d5914ca00d9ca714c7610d116bf852e906
z40c4c7e8bbcbd3781f27e9708445ce4537f19633cde89898bec42491873a93f7057526098d5b5f
zdd249ffb96e2eb29245d4f58338a97012e4efc1b30d9fc4c4f35742c08e32ab0d0d79518f2b35b
z2577a3717681f97016a4a07fd6884e33c7165a23352c3f232d5236672de92caad19df9b62aca4b
z1a0fbb762705e85a7ca964f15db393d8f703159e41ea03b19bfbca84efa12dd5eb2efce16397c9
z18aa2a1202078cc67579c20f617a9a66dca9e0b59f354d2eb28fdf6bf4efe11d217f739854370b
za2ce3fcfe95b0f9eec906a679c58ed92bec81f4c3a02c7df22cefc2b1d52d5143406893613eb90
z01cbe830a61ee447e20a6924711fdb7df49b0aa983e5342037e7083acdf50fe16bc57e97d048ec
zaffe63604c744b237019e7eeecd51d11da536d59f3cb1ea726c104c6b7474142401a95b58218a0
zbc6fa79b72ff0461f7e6901820513bf1191b06d39ba5d2dd3d9dca7ba565cb0c5d793dec6fd94d
zb6b87b8ff0abc627e6cc9bded9024b236a329f4bc0a77fffc39cfa51b4e05349d0de6d0678d88a
z4a99f8c7414de0687b75b73b7bb3300d1344b5d668dc8ea815999022a49d645c9dd87a2329964d
z91de0534307d6c5132ee545d86ab43eeeab7d8e9e84f56a539f9589141aa3cccd30570616b5b63
zf7b63e76b5bb5f0d0611b9d86cae564501a44cb70972ba1bdb2d6d16910c22dbb8b8b0b7516fc5
z3cd8f9d161d3975b5546e8701c02ee8e42a95f03dd9991c74d265efe1efd1dd3fa5481cb93d6bc
z214f70de47874fa2b5eecd39d547c34871e1beb173e6bfcdd2666dd371507291f81718c2781b94
zfaacb184b1c99a537d0cae7863526249f66fdd89e97f4f490d7c0703999b410258a3912656fb23
z0d50b53d64d71c7b6ece827a56d2b7c943d63c0be63cf776a634e8d731f8d58968b63f6e0a7266
ze402d493abbafd493ae0a89bbf0d6ffee2e85cc04781220747b6c92d28995e475389a97abf3ec2
zb43a4ed45ff67f7c53fd53c1630e2c6e48486cd8e60c9dc3f1208e4ac1dd1b48f16cb6387e3b89
z7eb9a908ca8a4155e29d76f7cf04100a4d94051c7faf947b512570802c1882ca9a1946945c0eb8
z4f896a22ba9fb930aea6402749f2d2bf43bf6b68f5892ca6e54744702f68024a5c17b3e1975384
z6da9dfbd5f55998157aec02e7933603dd4891307c16a909b17d349dc918cea65177d5e7edad5a0
z5afbb32218da6259fd21312741d43bfebd1335c2dc82110ecde192aae9830f9db0e0370ffb7f21
za1aa31374cb42c4bab555647a27df175d4f65b96d28350d030591790f0a051325b96bf18b8effe
zd493a7ce6d3dcd0f764fb9da53a8514dc63c01157573dbc845ca9e13ffe73d8ba6a27bb04adfa7
ze187807d18ebb99072a1b1c14d0d43b3140dd5558a6e045022001a14677891d9722beaac81aa07
z27fef808189f61043187cd2642991e9c22c4c1210666ba15092ed397c93852472239cabf766435
z1bd26c98e897577ca2009b897af5ce5afc91837f5fe9da3c979e37060fa5a437ab33467037ce94
z617fb9085c533340e07e36a9d959b3c746359f4759cdbf6fdb4651541059c73aa435ad77c0b916
z7b9308405d5b495c9549338938c39977e55505675634b209e57cd187b72eb77e6a4524c2f577ba
zb0e001c8363891a6aa0115402205fab1b17549871ea2d23d535ef8fbd65f0d3d3f08cc969ebbf7
zcbd1f21a4bf8eba373a4a03414ea86723762b5ee3f461ed8a5ce8d73f22c7ca6c467fe7bbbfa08
zfa96b438c11cad8e8b65164bdfb4f359c64b6c98625e43eb11d82e3a4d74a50cb3b79f277522c1
z9f047ed6fd55855cb73a2c88e1d452d1f4a9e2299dd3815b27eba2e4f41ba193daf5b59d940fbd
zdea2ab1d646bf421f280746d0ccba64e474a1d692a8cdde1c4e3c52a57ad2315f99cb1b3a92bcc
z0e61617cddf5fb137afc1d88e892352b34e71bc91400364fff733fa9e2b2889ff78c3a3d8597ef
zfc2f53bc91af71736652e11d8faa46ec7b89ab78df00a1c286a069086d7b4fd68ad568f2f1c4af
z178c9e7c49f513cc9932584176d663e0247a02fee63ad253397812f3f5166774213d3d8acd2191
z681c6096210d12e2996f35b4078949d3441ad4bd02dc9a61834c8c49e4a446934cfd2aa91b55f6
zdb5f67892ed729d5a1e85f0760ea280f0f4a175ffe0c1ab1a2529a9bf2d322a615f4dba28e775f
z37bc32b478c517a5e82e1b6477918a461daaf3f905d036b69d3408e0664a52f6afd2c81393bb9a
zd383b3716c1aec9bebbe5bfc24484bc323d1182bfc91faf36206302e3222356526e8716df37dd5
z9eaf2b295c1f874acb370b917d4b3e442b82896335a6434c21c4573884c75943227c1028b43f24
z128d742adb424442e0e0bfb5b4da0ae114ab4b053d11076419329a97a1a778f1c1bf849f1e071f
z505999cec537f6409c00ba5d0c195ceff9f245a090955246611db5f6f52f3599e20bbb2355ad86
zc0a701e52e682833fc27f7932f46334e821defcea2173ef6b004f46c67af79396ec95dd16a5126
z44cd5d183f40a8ef85de5fac7299b6526a7003c1c18867767bca208a927c89cc3f324217558c32
zaeeb18d724156aff555b756405d45b54bf291d8cadcdd152536839e2fba06137a8f7667fe9e94f
z753a491dae2e82b1824c69f1a98015cd3522348aebea0d8e3b62b7f23e471b95dc9554b3e0b682
z23ce131e583f6a9806ddb5afb4f7c1d54531714027d9ea673177f0f7c849ae341892f7c6082c43
zdb955dbedf3833e5d03d8592669ebda5f49b5b4ea60a56fb7611c8e750e4feb6bd0f2f0b3c033f
zd8a659b28d0d2d0cd51f7a9a5995e52354b5851f04554ec59e4cf421d67bd6b79111121ada498a
z8acc3fdb713ea94ac54702ab99e5c0a914ec4f0f1c3cf6db91610928c869321a98a084100d0f50
zaed615752314a4f88d2686db09c1668227399eebd8a5bd5d40d4b03771093a1afcb13ea46b910e
z1ce97a9b3b912c8ddd3d42e3f552853d1834c71b534f3b6617e1c63ed421c4f740253d3ecbf2d2
zcd6c7977a234983aaebcf9807c82205a785b17cfc7bfebfe99dbd3cf34a9e579d13023b9c54c1e
z8f67b1aa8ffe6fdd8d5fa97a50a1113490e782a9e1e60fb29a265c6a3b21e42f29ce090af16476
z64800f4bb62ef12d52911b9dd3c777d587da27649d42f6f76147d77c21d78e032120946db79a4e
zfa25a3add8e83d9c1bb3808c52347b9941fe6acbc78638b2b985c5ee83aabf8e4743743cabb264
za7f8bc0578c8a68321fde60c5e1d8105c52caaec0ba4bfbd3c3c0c0e21138926b5e417ff6dd3c1
zbac4890840c61fa50a0069fd9271bfc91e1f68aab6422fef5a57ec8184d7ecb740a0df61fbe617
z9f09273190576aff579fee43ad3918f26a58d1e35a5c11023af64a6d6c1c5cf6f2902e22cd341a
zbe4fcb478817b8b6ef0530374fa913a53d7ac03e23cb2f4498819f225a8fbb652f347a827e89d1
zcb14de74fe382586c05b624dd2db0edb13f9d272a5660c9f9acc06d531db1cb3622165a8eb9f6e
z90ed15ed3ad678995799b7eca2c408dfc5b05fb4b4d0591902d86b1c7e7e9c84ce0ff60b14b775
zfc4ba86d5516dcddaa1b377faaeaf144040ba78c7c637af2be6f76da542f0c1b23bc0c58f10c8e
z5024e8778725b6037d2135d6a1be5b8e8a5627e54b1787dcd359ff6339417065677174ba80669b
z0ddad57d4d62a0b4e4dbac40c4f4bd5c22ffb76654dae95c85daf1bfc1972532a42f5123fb984b
z8cccc893b1f5fc169e93839a4e78ef1cd86d4077dd036cb9fa141d2e920f5e72760d8df3e33183
z5f93219fa996c237e25293ffe09683fbefe95a296d2243559c60df8247cbf2b06a2aad97849fea
z6aa0299d8f7933fdd8e0613b3382a4636a57425e32e4cc2b54fcf75c126e5461b4e6b631c0b610
z94acf61667a58a3089847f3824db94cd9b45a799509bd53b456125ffc9128cf3574d513a8f405b
z8171c54aa1860670f09a7f8ad66df99f4e74d16e45bd38c8f586de5154ec9fdff265340ba44b94
z3f65f7f6f834f986022552e9002ddce74769e99ac0d61cdf720f12b276ee85d06f7c4000671cce
z15b4aff402a1d5fe3f02f4684e1431b08c4b9cad563dd8cbddb7994abaa92e9709be5fb30815c9
ze36c64ef08170f8f53ca0675552ab01845b9b2d1518ed4cffabfc1ead5931524c4053a8b016b5b
zbe074ce3107fb51a76b715a69a878f39e3d6ab6e1e9ceb69059655c87a599aeb2ca600ced02828
za90905273c209aa1b055c31f63cf8e6dd6a4a748ee24f5d78d0c655d64b4c37dab2d82344840da
z36cd67b34f5faec8ff5c51efc88b636899dd4da91d162e906a1a87185106d6eeb920f4f9d15a7a
zd5bdf01e2e0512701b2585c630f022840864fe9b0c1fbd6451b9206a234738f6fb7abda8704d66
zce1a78af44edf3a25920ccd68fe159366435f4085f70cfedcfccb013b468640ec207b1b8dd1cae
z800639290db98f6f60b39b3afb3c7ca9865fcbc5534090e70e89952c8b1cfc48a4e9703467993c
zfd1a2659dc3fe360ebad3a021ceb7b41e12912624a6abbdd31a79ee0c163cef8df37d825ff7d96
z8beadf9615f553d6393f905c57f68a743e047ce020cf74476842200cc0e91dffc3d5dd9bb421ce
z1078975a11c3f22b41e6d125f75dfeed67101898acd675c2d03c251a54410888bb1a65969595a1
z448d47944c5eefd9a9a7bf7b7cb12497c36160368f2a1cd69ff4894c72c435d539fd8dfc65b6ec
z66a715e5ee6682a591a6820cc42dd84050e7161acd4fc243c4f3e603805a496aaab5a55988715e
z614115f3a1c298bd330b84e3edf76fcc39ba8312bccc29355cb1fff9184edbfc02dc4e18f495a7
z0d7d17d145e7f9c1920ec686a0dadab1950791d9a9228a4867d5a9e60402ab541a95523688e27a
z09b3834c033e067c2932ee923cde56fbd45ae92dd75acf5a955cf97dc961d90c1c66ee84fa2f25
z8d60d9a3b2c0c427982f2a4dc0c9f44b30fade30e5449b99343726ddf80ddd6cfbd17c9b00f67c
zb36927b686a3d5c104de84fdb007731b40c4573dcc21f56f3d4a40b60ede1e840a006e5f2f5b1f
zd6ae3ab88677b4cc70ead9ac06e90372ebf0e31cd2f95ef99e9ec45e1cb459c4a309d26b01c9e7
z953cb1a3bd842320c2dafd860758bfd54f74a076362933cdaa056f38257a5dc498c8bc1f382c0d
ze2c97236a3487c3dbae76ca6fde2ebffef93ff98a836987779e47c5d39cf310b0ab90bb94ab273
z9790b3c004eaccadea8a0b0c58b7ef16dbb5b890e1643fafb15db1dc4fa77ee277af5157d3670a
z5cf2df90e5f5dfda86bcff27e8307d4797833f4e796cab365307e698dbdd7805247195df777a03
za24dbf408ddb08fc6d3d389f56fae34fa36a32b2dc5a16d99e8ff1e4f8bea6a66461925c27af88
zdecbed3bc7ffc687ea49700cced022051a96f6976013a7f88c125e2b28444e5ca2579644aaf469
z361627feaaf66e1b22f6d94d56d029e39d37812c1768687f2154615dc1326c2a8f4f875c83ee06
z107939e96b926c0e8cba95a6b53cb8ecaa1de76dd072fa2d8beae396b06a8e971b1623f49621cb
z0f62a359852d8593759dc4abeb9427cfff8bbc3beae5df2adc77a55663a56a9186655c4536ff55
z3a3ead40efe0098b587b977fd5bba320ec18f944d1e96290ae0631973b554d4ed3a785787fd017
zae8f48126245903cad9a7730a60427c1c7a5e79d2bd395468fbfdbe8c7fa35766f8dc7d34fc509
za387038a3d1f655c23973a45b7df503289d62412334e336ddc6a62a1564b680dcc221510a693cc
ze5060d18cb7b91c7230ff843aa59c43c2db4f29ee9f78eac71c65ce33de2c72cf4372f6c5d390f
z358ad2da9e311fc960ac204fac693b79509be471fef091b3aa591296781adb08e8791ed5f9a1d3
z8adfb3e8f70b986e5506070682e5f6e56d3437849e9c5f2eaf9142a1366855a93e07cf0cc3ea63
zbe9532776a45ec3c0bf89f52c0595fab979a8d6946467b918be7385e82ea22112661cd01f04b89
ze4a328a589170d96d4f3649d6ae60ad297ba6dcf6eae62181232ce7c1449589b2510cba971c0a1
z19167f6f2538ff7c831aa32ac6ba375ace0aa32389153f739ae303ddf77118dd4deb5efe3c84e9
zdb5d08a9b47b3ff4c6667bacac1a0bcab385a17e33ea905cd32a3efb0f77af81c3432001269642
zf7b844b10dabb26fab0e93553f55c937e4f425fbdc3a88a74b07c78907a7eb8c9d699afcc03513
zad3e249f64bc10154a19f7c4673b93d276f289788257edac64702a96c83f2d32f23d60e79939c3
ze8b7c7d7524646f0f5ca071afefc14db4b087c0a1b094e80b9337f76ff7a045dadc7cf9654ff37
zc546dc445ad967d0d90b3d2c2f4d9418d9cb400f2ce13c98371d4bc4cd0bba83a22ee12d4b0d25
ze750f8c832f2ed780ef9fdb28c5b7befaf05739be8555f00b5d91c26dbc06e5d355fe614195a84
z068c913bd24344c83b9a4393199d08d8c37deb87dbdba4dfbbbefcf2992704aae5247fb695ed10
z71289aabbd252952a7bbcf2d5da5ee5853b3dd96e7b550f7261b163611e4ddeb3a6b040e364435
z11fde5283ed38c12e5eba5e29adb8b93d6c2d2f7460f5bcf5dddb952544dc08a252d847948f1dd
zc794d0e82f925fc7a68d444b8f3cbd1789dc43b91af156d48e329e5a8a844896d602a064b8899d
z59c10f2407ce64280bb8f1a7b9f17a7855b331562881bd06b1397bc1324efb134a8798740dc1a9
z71d79c17c4dfc4e7e8909737eada8b26c48006ef75e41780909edb2c0ddd143fdda5bc045393be
z1d57553791eebd5f23149dc60345ab7f41f8415139723430402c0c6e2d016f8a2ddf8125fe6c6d
zcc3fefcdf0b4e2a2be055b1a210b827181ff4ebe6fa1d24b72d89bf5d755d182a6206977311169
zcf645198ed68dc629ad448ee7b3b2acdd7a56f0b167681825fc1aa64d3467078624034280d358f
ze42fd09739076f33e4560f8f6a09d8ecbc48fa2d3ca103844ee4f4362c92e6d2057846514484c3
z3d0b5b5c06239891219935c49776220e69ac72f942ac0713938f1593c60aaf79e7bcf9b57a4810
z64171650d9edf7b027c0a2c3215dd29f2b7936601b96343b554e75da237d79576391b0b6b82970
z8d7ba196befd9f1c75675748fe74daef9956e773eacadcbfaace7630ead0ef665ef48537f322af
za04ff6a87e221ffbf5cefef7e46d2e7e2ff47ef2cd6bd0e68cf48b01aac203d7049cee99bb6157
z6d66b55f7d66418dc566276ea0ef95639918b9b5d757cd30a1b876d223c24c58a5ab6eed091949
z6d2d5b7e1ea8faeeebdd0b1efd7226f3df2090c0f67f9703b86dcba38c92a510a71ebd49abebac
z7538efa7cf67a3a9286cf46f75e29039d05b249945eb88b380cd1ead9fa1bdef0c66cfc0aae893
zc0038be922a5928e28dede97eef744213b7b865c7f583a9c07b37ea9858263f24eb2e6a6dc54cf
z833ce44bc952d57949c5a14a66cb5766c9cce74dd35ddc5be140b6d324e49680d4c01f27b27d10
z0edbdc0fa809606babcd3107373184e7cf53001f35f8f6f3db6c3d28cf11c52d15c4f257882b8e
z37133cd692e5df53eb8151ce269edcf2d7d5ea69207a61c0d94ccaacb6379e60ad4ad67c4e2290
zdd9b40d6980b1014cd827bfb06ffaa1f5148233f9fa77e995ef6352a8f6693d7bc74d841b2d9fc
zb21ccffdfe68b9c6c16dcb31fec24235a0667ddd2ea28a35a8db9d856040a1a5dd661d6e4a5913
z63b9f4fa10d42c208c6587bb49c47df8e384c859919176e84606d05be983b0ab663edc87ae1837
z69a75c73bea811e437d28d6043b7f6da0fea40b7f25decbc21fffeee171071db39b58c34bb0797
z0f0d82140ae35fbc401810f37819d410ab152da8493b819bb6c06189d35b8edfbb79902955cfeb
za781ba5c0a0043a9c136e16bff50f6d69f832fb8d83b81e54dd792801d689523d18bc6d25b64b3
z5b8ea144da8c10b3fb1d58cdda28dde15ecf2406cf7d11e81faeb06e5c51d4bbf0d5ad5ebebe17
ze92dcd9a5b92db2904b530120385977cf6d949281567deb1eecf301be82e5dd3198f4909ae9208
zd64ef6f6e61eceacace94099582cdcd5c17fae53e966ceea92933c61e2f7a3bd892410170a4774
zdde5b5c8aaf15e8b3b24c0fe600e79e7f72aba486b6c4a0eaf49e1f781f97a3925bb98343a4483
z99c78dde589dcbac38809158b7d53e7a69b3b2e3ae0130e04510716f181070267fadc677f9bfb4
z2fce6b0ed3941acd5e01fc6ccbe2483286252bcb42fdb0ba018677bfaecb4fa268e1ed9ec02682
zb16930ba1b6a528315ccd55ffe4219cf5c78af690fbfa5eca77f1a735d3280191b68a3e73abf20
zec4ed496c159b7739623b2c15fea01edff74992ec1aa2dddf7c41c0e495e6d2614b991c5d9ec6e
zc97bd9addc14454226c04f684d16d21beb1d3483dacf96082da48a7e0ce913456c389b59cd1437
zcb8aa2ac9b27cd4491718f8db97af6e91b760e9d2c08f885185d02573410e85763a8c498165d2a
zbceeeb2cee95be51a9526280b4102085b1f1c07aaa3fe1ae1c4dde8913aebd492d0e89ce3c660e
z98534dccb5a01109edff30f133f2b21e7744fa758930e38726071b9b647c96370688a683ad115d
z4d6fb246d03fc48e2bc1711239bf35179d1992d18d255452413e686a283fcce58b7e57c5c512f4
z60a9c40a8b7ae93bd583a2d65c5cbc143d88c80af6d5cf35d2b53d1491eb26c4cacd61c9a1e417
z4c2c26d93e55923629afc389580c4d2392bdab68702d50015630ed05f7c040280a7843cf28f8d1
zf542948c2ec41beedf1ab6adcb8da29073031690ff6fb5f85285a7641571d47d08200dc74981db
z2003dd598ba0f7ff8771a28b2baa524d5042803fe4589c0dc4a2957e1a4ae0cdb1c9b7850a9fa0
z1acb78e78facab8309cfd31b422a6bb553e9dd163730ef1a2c60fa8910ff4f493dbba357f80e19
zbc4ef86c92b33826a6e600654a031cdcc0f5bd295ab5b60192d21544cec5ca2dfe7bebbf4b9a3c
z9adc2db883ca9565e23d9edc03d1c70b1ec59d18b2307ce64fd5fc70ff50a6dc46c2efbc9343d3
z9f3875b0bf9cc39cdfdfda10bba5dd4810e0f7906fdd8a9bf8c9b4a29ca6873c8ccac0ca7ac26c
z9615393fefed10dc5abc828dca50e6a7276652c903dc09966adee5af4de7704ad593e4dd2de14d
z7e1a8a639cf1a81e290c667d4f4e25e194b4f324fd2def1f31029fd5776d711f1ef2c7d0b56442
z22e6db48bea809bb7cb3748a629d7dd86f0c11882f32c72ebb8ecb70647b710de3b96aed295e2b
zc47c6be6733c76685e3aacbfd55c26e4ef51fceebd88ae5bb81340b0b443fefda59e92e653c053
z608e76a38ee767c714cc3c6f51607ebbf6ccb72072ba0fb423895d6328bf816159227aad6d1b86
z371cae96e06ae40ec7c9a7fb60559f1824e982e9671354393980049b3ac3242c9731be7a31b2af
zaeae8b547416b8f20a6fa2d9f7bbbd773ca6adb4044f147e46dd69fb3fc4d0ba457522e4601f50
z46fa06620879e7f8a7eddce1d8b3b593da8227d10b637f9e198a0f3abf9192683194166cdcb5d2
z42a04caead7beb02c7aef8d82005cdcacab0050701c2830da56991444fa8bb3a8486a7daad2caa
zfcba6abdbb8a44208468db470d04304a5f7bc811589f0fb40bde71fc5edbbed82486135065dedd
z82cd65535ef089e24b832811a2980b1f866986017ced643351d550e761bd825becc929881ea4f0
z6a10c6e7eac9a3efe0c21f56923f40c0a87e959283dd9bcaf95808fa68ea05be4b30e50a683a4b
z64cf75a452ecb7650141064ba7dbf298a9e6c346a19a9e39807e16b40eedc122900d6146ba2e06
z9af67c29dfffa512d93af721b63375c81e2529df56c4d2a5a37ca3896333bbf9b15604d716e5d3
z11d5c54eb999bc708a2ca48d40fc81696c17270485a9ec9a9616a6d2fe159cdef3c8f8b23539f9
z6f31572371e14dcece2c3c1b8a674acc21ac4d92d8d63fcb2939b84a1d61614d48a6150b668252
ze9df85a9edd8634d39748d3cf0b3c97ac5f5c3c7459d309628d51746a4c21f5dcb084b013fe299
z6ac44db8e7d1a0ea9b09999ffca0c65a7b5a6b23f01b3defea693e2b328547080ac92cb00a2577
zf97dd5e768cd365a57a6eb595a9818306d5a9957e8f4137cb0b2eef7c56fc86de4b7af97ab68b4
zead4fb061e2996bd629c4c6705e935cfb6bec9382b632aa688a7e0a51f3dcfbc62a704e59f49a9
za115f9b21c9299d91107ccb738ecaac6a9ca3e77084a5ba6f821d9ec513b5f5a6cf2df6d71a09f
z1092eda30f0030bd5cc09aa37a99ea2674cd6d79a5e7301c654b20e5285f3979e2e21d35d6e669
zfc989ea24023e5f949468bd607cd0d4ab0091416ecb1e996b7e9e218e462681b56d0f9cefd3bf7
z6f4a09a5ab31769e8deab8b81e1466312b554032f45ba5e276f0557ef21173d98335bf47a6e69e
z588c422731ff864d2e6fb489bbb6435cba317834d8d262439aa767409cfee7b22f69b80c4fbf9e
z70447b35e88dc1d4c2abf548a2841f63bda1c27afe04554292ee67ee9cb70994d88fb7adb81318
zb98430cc73e07fd2e45518244447c806fb07e46816bbd0c5e177f1112e573fb8622fc0d9574d54
za0fe7edb72e461ed1ba3017deb5e02053bafa6bfe0379a6d1bc15e617a73333f64ff0468ea4cb3
zeb6754aaa6d4c3e07f20a9d12a119cb66756818bfeca001bd8012acd969c058a3cccde729b81db
z9ea853b2235d180687b9d89eb4a06a4f5a47540cb86c6419d304d670496a5a3429017639b5b2ec
z1dd2e0538f6605f6566470ce415309c22d0f1b315c5f5d59fb0b1a6ca053023c3b3336f79e78bc
z6cb1008928d4c24c1e6c251c03d339b255fd25a716bc09e8f23e5b6a659c07e9a03c3a92395996
zc808dd13aa2f0e6e6bdac7439397057651fbdb31fbaf120cc24fab6a01cd43088fae5d65b64867
zeebb04ef198f202cf48026aa8d56824997a596da51cff2e963f51ea218114ed52be699cba7fc3e
z7ad997e2aa11186da1fb3203c7fcb70629b5eeac72a9309b688c2eb9a213341116e41328fcbc1f
z2c85c0e1d15a35350800922511437790518d826d2d6e7cb7f20ee91c79ae15ebbbb9b2d92da2c1
zb75300b2e87213f22f1074366ccd69446f9911315916bf60cf3bc88817c863548201fbbfe02b47
zf478f4207325309159153169b7b420e7b145581cbd62b0306f0076a08a2e8aa1ed980460de3002
zddf42f440925c1ad8eadea5ceaae54495045830c0c39e83ad8c87c41c3f48c64a2f6da56fbe228
zf3dd6287605b32545e528c95e304605630e966c3378766d79e40070825f5a776f6d342ceeec2f8
zc724bc53e77761b67e402367126f35ac88732d25d16d2825d337c3546c25c0216660c2e2894c0b
za2546399c0cbe53fd96d0adda2cf11177f41b3a68906d7759110635bb1b7b42630a7982adf0521
z54a8ec368413af68d05fb1b5d200b33e9cd881cf02b4b1ec942d076cf1cf59338e597dbee74c30
z9ed7dc13a70331e8be7c1f935b251b98f38775318cc0aeab892f05211a572dad255594c48bc4c4
z93bd9f6b83cec1b75c8e5712b3b00d8ef346ab9ed3ad663a871dc330e5c93feb7a3d513fd740fb
z2af2387d73998c6086ee2b193ded9004d2a8596aa2156d7dfe2da469c6c9debf999ba25b23ace9
z1092cb5dd5c7546c6a3af00d5ca93a76da9a5c6998ad995084118ee6402d7b8a1e87eb641d083f
z41db8cefe0d0a9e1a3322b1bbbe615045dce7b9f57c2b90fb44808c27dd59244b34903166817fd
zbdb8645b09cb362d77982adb6e6140622ca1b4bbba06bab58deb32dd67db8498e1467c7407de3f
z5c89cfbdb8713ba59572c853a3828cdf6c21d72ece52cd6997a445182be1bc410099e0f95466e9
z665ed29edd16abf2b9b1d91d2514d5277945439039e7d07291a1eaa3cfd280abef6d54b27b3ccc
z9f0cc5861bcc36bae566d7f09ba49040d7510c85013fb4d6b9a83d711b8d3cde15f3515f849ec0
z5280674fe8386135a0005fd6b61eb23ddf03f0e8d920a5396e01a956b0ae2ddc9088f6da3ca3dd
z1306645a75700073bcdbda3f35c3102418efa4c246b2ec976803f492d9907c33e2452aac284738
zf6c250b899b8522ee744889aba7883fe39dba746a8c2bebbaefff53969b808f0608d7a7fb3555d
z9ac9fa53da1d905152a1fa97aa2680fa277620b8751f47dfab6b284c85bba3c15c9834d202e883
za64d54c572f5045fab1424ead281adcdc73e45499e172f7def6b1f073e4edd0dc609f695583a39
z7874d9aaa20d1926a06a166e3db9d7d7709906e4e78c41731895d4275c09010fa0b500dc62e103
z240ac83ac1bcb261afda5c8cd4fc9f6dc9b97eb089d7ad4ce1b084b5efa6ca3781edf9b06162a7
z2278b1ad48998bd1346e67f3af896917c7cb5dc3da7249f52c529c62454d5c22f6fc9578587eb1
z6abb010589b24103ea1348bda7756e642f2b7fc66182d4346cd3c4c28b14ee080d2e15e2ab8540
z831850e11988f3cf98f87e7485a4842422bee17346f4d28c8deaaa3da2326835821483a62c3655
z6c58ea63e7ac795985319b01a9ab51056a6aa2f3fa94d77eff204fe216993232bcae5550d13787
zcb41b929421a138537b4bfe68ed5c51e71ef35d8a9693ff940319d5e9d0de662b2e3475a4d506b
z8c9681e6db0fe76c159348eeb485582726eaf89d8834782b601dfbd3b1e759484002d22ac0795d
z39ed3c6c33cbd1baa4fe792045fb09fc11ee29358630da6bbbafb7971551b8c876a59c4c6c30fd
ze33b49e7fd8dd5c62783516f34a8e99d3f1247ff8ff12faee13a5aed63ffc7b402947e2cd4b9b8
zcedf7ce7320c4e1ad263a1c15718ccbaaded2704b30b3c5c4d15f1ef2bf7d1630fe308c0779783
z19a68a10c54d11cd883c8c0b8d05849f09b99d7ce271759a9b9f498f747e112c663ce41f0dd10f
za37e3d23dbf2d62cf4851929bcc227cfe90482a5062655bf74e2d5700f29ffebedca538ea12a45
z93c10f5b9dfecbb5950e755365381f53664a1e4d6ae7f808f34cdc42381b75cf8d374c41cc9a7d
z8ff5c0bf0354e6147c09845492f7213f756ce56dd73df5090d8db3e302d15a4b5e4ea19a28aaea
z5981424035ec01fba7570d4342bc6eb45e66a187b06379abb5b822c2f382002e53538c93
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_express_transaction_layer_pkt_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
