`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bcb1767abf
z37912b984147c77602346f6d603de593bd477dc820be44e98597d42ac91ff344a7c650ca9c35d7
z2dec3a4f295b97023b5602d92e73b63093515db470e10a4f3769defa41ef4fd47de24f99af10eb
z78f3ef7556c4fda5c71d69e1ad83f774da504357fdca409a1c619be026593bb02e8b3b03f9f49e
z9bba8ba53ea44a39924348812e26745252cf500b272354e895b1dcda769518cb4bc749836dee04
zb6ad97bd27485684b617a2d0dbe522a6d6b081272b0ef8f7c2ffd9abe41b89a8b8a564bca73bfe
z649dcafb25f868e84e18e45d5f8b7bcb43245c5e94642324fee7f443b286f1c6b44abc0f2352fc
z8c05a4d18815434145c8dfb51f9aaab5b672069bbe930ac14fb8932ea5b215aedffbaa5ffffe5b
z211d36c55a87441c5405a9c8f513d830f09e8da53d241ad3c74aa222555fc855a89ded2685816a
z4d68306efb7c2d9d0ba8b931a37bdc4fcd68662b113fff9ff23fe809abd7e7bd1e5735f9529eb7
z2bf252c1dc3395b2f81548349cadc32c481b07a5e87b8f6269380c5520cde6e205042bd3e52f04
z7567d5f686902a4e74b660622ce3d2ffd45777a5e1b504768d98b263979f89be1b13d595f2f82b
z36560edd610e4d4c8348bf7446c4d204c964a5e28a85222d1ed0ae3619ccca85ac6e7452a93232
z149c49a57b55c774ebfdc63e21c4353ff479eb6051e40ddd047b19c637821cd3a0069583732b27
z7853ba83477bf0895b8014a6f73e81e2861e5554d86c503b055559f7b038702ee6bb2146ccb062
z03726cadb116f96b933d423b324365884d6e1585c4efeb0f2f3ee241de918c857daf753619f963
z81ab8bc103f4933c05196a08cdbd561f0a0e0161b7f68dee14f4df64180b37c508cd2d33496f65
z62651b327fc8982ac1dacd131ff2ebb5e3b284071b9e4854eb78acb672f7c6e079d565259fb240
z840f4362ca135c2125aa1bbd903c14d0007073c774a8c659bcde1276541fb0ab56197810498b94
z932d266b6472a76ca5f474c7d3e656dbc697b9f574fb33bfba679fdcc2ee774625fd60296e5695
zefae799b86efa5ddf1586cce8b7bb26c303dc8053799dcf9620fed3f5a3d59588093dda9e000ed
z113818848ac8449d5fa420338dfa5842bd5cd8c65f864da14a8cd82406e84e161b54eb851240b9
zb9e6597ae273753470fc833236b58efb08f9054123f1bcf3284a2d51afe8f643762e491ffccdac
zd1ab9cd20f8a5553fb4b244bc9bdf0c922633ffca218854e64a2a9600e438cdf7a8d43a5506579
zddaae296548584ce5ae31120de73e179bd7a0d02fefb7056a681c69619ed96619612eb5bb3c006
z41a92cf9b67affd17ad0a0d143d64b884a46443dda3c9009fceb22170a58bf3bfaa199c0b078de
zd0e39e458b92f4342ff01251a9e7247b19d8a923b9dc74e61984bec6a83cabcc6f8fd7a0387c40
z9eb9ccc074989553de4ea8996ee38d49c63d67a93a64daaafe9ae5b6d8c9149dfac126f2e0c822
z93281650d7bf17decafa3fcaa129769e78e907005dc22f9d5f8c4f5c53be3cbbdef04bfccffcfe
zf5c31b0fe775c35f79dfd33081be5f24b5af1648cc353190b0f1e06875081ec6ebdc65cd52dfee
z6863ecf050b35f58d4a54d4e758bf842c2776a8e3a1d14928d426043b52c28546436a493163b5b
z654d37144bd7f0b1cfad224f52f65f02046798e43754aa50e8e5604ba43a1b7e74f51a54a66b13
zb8191947a354a55d4db66745c9a3826adbb73530a2f8355f80ec0f6548564b95ef4118fe43679d
zf485d9729d1b66bf898ad2721e208d924809db4c5156a16d41e4694e287f69f68e29fcdbbc8f51
z84fa0991d795465fbc2ed8da92f624ff87a33af99f027cfb66c7b1995a399a9326df95f6e11962
z2f48a45fad82d42247a8cf98cc89eca9a3b4e463e1493dcb27ac67e79a723cd5db9b3e3f74e181
z010614045ca2f64d3403311183e15233bcdeb02f1cbb347858f9bc5827d0d177cf53af9c380923
z6287c51b3054447fb1a7469174ad22292ae60f3577233e28beb9958a79c8a59c6240a9615937dd
zd8a1bb86d9be23417dd58f466d938343c332a29fae0922ac402f61b38ca3a348942087972dc26f
z7949192f807928406307cc82307b5edbb5752d34b4791cc3125f84ac250d6adef0ca3c4485324c
z5fdeb656c9402b3bae2e6bd3dbaaffdcd2ed632bd7dbd49ec49094f26dc185755476dea119ff45
za1a2b4fd6f911849c01827e640c2eed1ea1b0e14b599768ed07746ae4fbf2d299f16b3610bef86
z974292b69ac2e52ff7f069a12ea48432ee8b47838753da0efd97e134ee1df225c5dd191422e695
z45754578a52ccfd3efdd69111635f7362f501e5d5bda28205159ce973dbd32c4a93f377a1181f4
z560631a9745315ef99d30a87bc74e99fd087e7be9ba21d6e262f25ab4ff10e995becaa4372a357
z77539776d13a49812fb281c77de668b4ad6ab3de91f30fa70f956843ed710b5848d77c2a4a3922
z9159fb361f89e42a648f30d2e29892031ac79b645d65fa4d68bce85ac9d396ea7603732f49be3f
zb3b7bbd6e365ceeb9904c749753be0583fc9c40437570b5e86a7f5e006ab1e93212288701c255d
z342eb3e7379c3cfa1d2a8991a045608fe594fef5f6a214b43b2170179a441fdff9481979a386ec
z3844d7fe4ecdc35adf389514a52b93ccee559c3aef1cf16f89b35e036d036fdffac67cce985798
z77f8901d035a837a063ee62cb2257d6385d8f30bb7398c5b6d658177b933ae31029a4e23c87b4e
z61d63664ec124343df0ddc51cdb099055f4f21379d80d84a21f7330d0776959cd62dbaa5419f8d
z35672df1d1812dadf0b2a773a8087254819388619bad9c68633905298b336483ade4744cab84da
z1873a2c05d9da1531b9518da2652f428de688d821c0ee7dea5c1841f48414cff85b0cd3131b8be
z27da8d178a5c19a55b348951e3ba4a2f39edad234bc0211623d52d93896ae4bc825e4fc4bf8373
z3ffaa9640ae812619df215a67aa86a02aacd9d7cadccc89c1ceb87cd2b86774a11a43260881fda
zb0871eb1d2b8888803448914fe1b0e2a1627b195aa310ecfeea57de2436ed2fbc4bc3b584e1d3f
z4f34ed61bedbf4ee974f941d0d68775b5461fb8b509b8cb20b97e04898eb3a3ba7bea4ea32843c
zf99e4c5a11734fa5fa1b0131c59d7eac8e18b435b0233481b61eff62a211ff8064029ee5e59212
zff98db913738f5d1ac1c2dd87f9a69ba9bff51dfee33f9f57202c24ca35085678a40e2923cabd5
zddae871174391461c47f93d6c5c1e2f935a9b1c7f74b5c40058e65cd2a6bea76cf40e01903b077
zc014afe0e954215e3eceb38306aa8da546c639040cc8bdcbb3ef84fcba8432751123be8eaac750
z7e3fb4a5690c9d00d881de94d112c0655d62d47b68dfd4ed64d30455d33422de04080895253ffb
z52deef5862d9b9f5867903e6002d80f4ea33b4c64bf9a26a4ccec777f17b498936b8b2909e2d24
zcf3068a50a01097aaea49d6cfbb92cd39a666478270a45bdbdf2760fda132faedf7deabc19498f
zb62e12aab57b53dd01bc82cc119c34a54f3b2041f9ddc5c0f6644d333e016295b487c2ec72c929
z0f016158f949c8e8c2de82304f3ffb51b26d76f0d0d48cd45b4d47eeef57bebc5dd5bfd5c753ce
ze24a0adb70b0156015ec16fe1fa8b9d59961049ba2dcd79a9ebbab20757faf151a045ff4ae7b9a
z6f553aebc8e4fb94fa90391f784300aa1983bf9aae0eaae81526be1c5ce4a91456e4b0140f3f4f
ze0ead715b0cf13419c09d9999c624394ef2cee78a72c91713c5f804fd497b49795c20e215404b5
z038ff0f7029e35d0610de084b0e97d7658338af4bd1d1cb0ef197cd0e8f51476abe0755806dcda
z35edc56348eef3d65c739c46bc8f4bd39e55ffd10c570229e306dd5716a237c89b6d14f10a8aad
z713c0a295293ca664276b0a190f9f03c58dd4ae0681e11ae987d5288c00e1664c8288f7324ba96
zd137c9c0f317cc1de1c779bbba7547a21090741e73e79249f5e8820d912f080d218ddf14004591
z7c2f564413d335aa5afe6b7cd3350c38c2a476082f377318c8e4322256f5aad4386ab2892f2594
zf6b106d0118f3275fd327fd4dfc043ea3a7171109c233a4260f26a9dfbd16d149ccac5c8c7b9dd
zf73ded882f00cd3d4890506d77565778e81c6b9e94c2b96d8c69e19b02d052f8467d9442d32b08
zdd8c7af470ba1a3483b531d79c261370bdf346c5c3b3919e6732bf6d254c3b3b301798dc78d104
z175fd7da2060a15ff1c825b86887b20c5e7e3d667aaa2c19f4f1d3bd083cd6165b6c0a66d3bb20
zac574f770d50004530c464ac1c67c62e7bd67901422379ca92e40ef54219165c1c4530376e0394
z8d73cd029f75238f25d73de0126979e159c2a641b100fc9bf109e3724e1c92d5e6ee5663486448
zd8e96ee666852aa3e8e907b7cb43dde14314d21228135632cad7982426a4630aa6817076bd4c6a
zf6ab23df883b42c9d0f52e3e4d51612db2a3742555c982e29a7b6e447fd4da31759bbd1b9f031b
zbb4d3c6515f58638a04aee13637c2840a0e478033c428e67039abae744732f13e5594d256da102
z576bd9ee2db843ee538d96c326491b05ef25e00459fed33fe0f81be2bd91ceaa9cbf9e96d47ff0
ze2f11221e52a51b5022a99c45c8a9acd4881858ec57b68148a831d8051406a81084e972ed16b85
z60a42778da5dd29792bbda6db912356b4a9c6216c36f9a4641b2cc698400cd707848a6911a7b26
zdcd218c150e493f73d1359335ed3f217b4f5f87cf1f8214cd4aa431f3e6f656a9adeba67b9ce5c
z58cbca34e31595369285b4b2cd79f3b2021ac8f88d68fcfb6e471a58f7f5a6c3b9f7432604f61a
z9adaf7c1966248b9b905581e4353947ab875ff38c257c07f8d5d4107919851fad9dfd0ac0bfc2a
z9ce0289ad8c862375b128b8a949c8c8b71c15c97b025d3fe00ef0b4b4e51a79b57e80a02582b5c
zb52698d8291f41663d8641d6cb0475094b3626f4167c54665fe1c98278dea9db1d8998885093f8
zfe54fbb5d1c2b9c56545b5a9b7608ae1c3eeff88d611128267a6f73937cd68675c4f3984c090b2
z8d4b7c04270921110b8c5ae2d42ae84ffe4dc574b57b58b8fffb7c7882afeb55573454c5f949f4
z52f4e1146cbf2a6f659fc7001e8f97deb4a37025a99e29414d2533d6912427901a0088fd7e538b
z68ff2a6de1c007dddb0d4a34d70fa8a309b62c6e89c028dd5e85b38ee8409359ee79c013da8990
z9351ca8aaad129facf1c069e91ff0a40cff909ffea115e11ca403708b79e3f388bac03676644e8
z164fae805ca8ebbc08e77fb33cfada5e01ec9df88718842bbacce3c58d1d046929a28d9320edbf
z3c5b65556c7cb6a83a2bf79aeaa3aeb43e004a8d67673deaa34d32a5bd67b1aedca36bdcd6d45d
z2af0bcc571a1898e011cfab106a1f73df63fd86a76cfae1175e3cf78552640a6d2c47589ab228e
za07e98543e633c6c5ddd4efadb50de87a686079462734c20c86cbcefd9122c2feffc3f90130aaa
z5be8819f2d5a46d422c8825ec55ec335f6724d83bb4f48a81040b220360c2dbf35886fd999ccd9
zb7016dffd0c9e168f42793a62482a4fcc3240f72d783dec3c2e29cf15ada314293ee45f498ae0d
za280bae78cada097fcaf682ef2dfaada3a48bed5f297b8fdcd8294b6edaaf6844f331653b2e553
z7513772d40762aa980f9fcd6b94461185a3bd4f633a983e2f86a74470f64e85b44111cf9a8dfe8
z43916aa52f4d8e111226377a964f81f2ac1025da15815613861944d110cdf1791f073292a0a3c8
z7a6d4de0a05c73761887b31c4cf9222809c2d75348ebfdcd74501b501754ef4d5201b1ab025f81
z001a0961ff30b3ae1c87cd135686fe97f968a89a19b80f3b76a04cbbea896f971926af54bf4d37
zfd143a080232e4704528361507478c12ba0fe1b68ae83b5aa1b4d88d70baf95b7c6999c648bca5
zeabc826a6708f11fcaec2905d92bec409840c8b2ec9e96933a08cd9e0c17aea3f128b2f18c5f7e
z885484f939b458c293c100f4acab5766fb64137796af28d017b604c052d8d252ab44b090e5671d
z3df4ec86ccc9b98d18c990e29e6760ae2e549e7f52c3db0e79a630670c29c2cf84f1878cf5ca20
za8dededdd2a449bf59c1d3f8b8408dd0111d3787521c412595284f2f55c94d97269c14e703f59d
z611c599a836c414ff523543ee6b2db6780ddeaac3de9d95d9a28a83f73685684106f07ee22ae3a
z8f1d9493864c91a5cd192487afd673676115545762721b46d7cf033ddaa86ce9181dcaa3deed1e
z7fd0444781a611dcfc4af32d9e0e85a78cd818fd3956067e5205fe52eef6adae8ca1fbf60b5cfc
zee0c51a269cafcce97fba4787dd7cc3ea92ed3415b56a8eaa01de0dfc123a1cc925893d804419d
z6a7ef2694ab59c7e69bd2956079d973e1bd63ead46cb043b29a80a33cab563322e9b37603e401b
z4fbde572b1bd9d6fec005ceb3e1741b817d8d00630e2e2f2e3d7c2942d6210cb4f33df59b8dc49
z2391408c5f489ac8f38ecab46a6436e16cfd1498b5b3ace28bbd7e2b4be2c5363ecbd5bc8c1789
z2b0a76310de216dc741cdf696f8e21c05e024b239a76f595cda68b06cbe78ed488a51aa368817e
z8e1e18480db117d2c0be3c95cd998081ddda1dac7bb46add3776a1d8836830f151e85e9dee4855
z48c60b4690da8968a1e05f5caa599bc05445b4b3433c511e90466a976bfb8f813fce576288555b
z6e0096e5667286a05613a61b0df00ce6c2da49bc7b1ad834f86778a6dc94d2ff371a8f857593ab
z876ebdb312cb70ee20ce00e6aeb6f86f4f2223987c55a1dbd78c59c3258f342fada55868f4089c
zc4fa3a7ee1fa401b0884a2d673ad6e0839baab33c5a4e86f0cbf49f8e2d1a011ee9a0e921d59d8
z008e464e571bc5809c07453f40d81bf25316f4485ea871069b68ebc2baed2f61054c8a25bfff78
zdd8f6752c2cf9fcde6f580e8600a27902c1cb7bb8ac3f695417d5944b0027f5c5b331247007e38
za4191e2cf5cd4ea1b0138b9775b1be04b1ef22487984f8030fe7cb25aedf1626bf880044b76ac5
z3f64ae354f8ded4025bd3af6825b5cfb49f107d11290c4e7b73b8554f344c40d2097d05053f71d
z714463060f1828507f082a2f4738a40856b826471515ba481f215ab547b47f1995021dc1a22538
z50481b57b945140d92aff448208f02e124a02085ccb81d7ce89cecb73b1fd10fd8e18276012781
z7cf6fc95191a7943d563d2510eaf0b7a7598fd9832b9cea6d3b61c061c02c23c740225b1ccf47c
z92dabb66543fc357dd8a605ece4b677e8dfb746f205a014a3af65cae415c185b976aa342d335b5
zb5cde93733e400ea9e8ee3c6673a648de139ecd362f7422d2352533478b7dfb090913d715b7025
zc60ba492bdd10c85389edcc6ddcff5a388eefc323fd5a492fa20a01395b437706ba8d1ec91c79f
z9622879f509d993008f87b915d170e38c0d433b4442706c16e9f3dc7af846cc18ed62635ff843e
z08bdd5a2179daafdd4101990c8e3edd5ba49a0dd2daa9138b723793f1a274b2d154ad2bba30eed
z63b24617963d99c9804d915337d5505a06685473d15babfd4e36c6522deec61c1c81cc98966984
z9ac431d9608a2f53cc5b1c43d0af260c03abeeaae5f8b96d449b8d65693543c4ce57306d84ff84
zc08fc1ee41dd54b5d99b725686674e92f27572be611e3042f476d7cbccdb88cedea4477793f198
z79bffd1672bb8f6534a6b287ced16ef320e3bf84d745d109c6ff0592025968ff3f07daccd1b75e
z1bc0ec39f7b040c763904ad3d409c3c92c03e2c4ae1aab23d22087d27873b634391c03bb70f09d
zc5e45756f0e09f45e711091afc81a8d10197daa4c2c59a2ae9bd68246b99ece6734807ef85ffa3
z644eb38f15d5c289214bf59bc1e25a90ef2c6975b916256268048c2841caa9ef53f59c3239da23
z903157007d335782cefe0f62b771367f59413db545702bbc0def7dad0c4b3a8ac030c2616e1bb4
z1123bdd6f04520d0c3c522e0901ace87622345f1882bff88deb2f071bb86a00ca7e7c457d17659
z13048404bab3db5416ea9024e3b49ec5b5b9418f99ec90b87c7837dbc81c87bfd12a14ccb93dba
z1ff2be1b4393170b0a29684d191e7fbe327eafcf1707e460bf815d167d82a00eeb7e81a57b637f
z4dc39aa6c3f487e667896e1314190f6dfd85a48ba51f6abada8958e44543d18fa1b5324e104966
zc94a5910eaa8fff55757c6e8c01df8ffb78183de6ef8f023823709732f289122dd2785cfe04ebe
z758a7762443a145c09abf3723daefa2f60c8a735bf194dffdbe3b91a4b598de968165496822436
z89f48176a3a85079110ebe8a0e596ef07530999983799b480865b10d1dc829ca3b7f602499645c
z5a2b1f8a38c73ebebbbf7414e60017ce0da12ffcfa08cb4793c50a4de9390c5e230f2801a5aeb6
z9416172a9ea010a73a341385d85c085f12a8b53eab126da250d2dc221607fbe3d407b6e1505f05
zd4d9bd5e55e73f25c2ca2847b1595b3a59341097e2885c6082301ea2ff00c756784c113360888e
z2a764c6df6f859d6b10282eb5fd1560dac922f5ca3ba539ade25addafc4a23f71eae9d59251816
z8208a42eff8ed22b29e55a238f04c09273e4d579d380dd648adc33a9ba2b58aa6bc18715a9209e
z32ad4952aafcbc575e1ce04b1814b601baf9236ef6e06673db162f7d768f170688cb64fbff0cff
zbf9241fe6755e2ad7a24211d886c68c18e94e29a54cd571685c0018917781e1dd0231ce1be8b1c
zfa2b0f37d43d0c7efc18465c73d1c19874624329f87aad524035cab0597508206ff3db9fe9f8f4
zde0d49540e0b9e3d10be979071d278ea520d358feba326219437b2265a618f854b3bc4a8f35c47
zff042925b30ced1f5c40de888ef121d4002260c5d172a08921b76f36e1aaa9ce02276acbe63f56
zec2bf7ff5860cb4ca3c94c8f0310ed67c34cce448d249181a4b36da024cf79b1761de8649b77c9
z03c01721a68fb8d9372dcfeef47ec3b8a4e70b90fedab1f137fa96b5228907176edda00678e163
z868674bec1bc135df426020d8b57352fd269d830bc5962da50bf59195ec9ca7c5f1542a025187b
zf062f83b29d512d2c9b08574af2d0a3b9eceee321bf8a04c364fd868e73524a53fd56cb59057a4
za81439d5302173e322fbb13c5425201317996e846c3d388beed2d997a86f5c6c6659ef97ed8dc9
z29dc9f080a1eef770326ff64af2400a8170f2e25eb814a9f934d3567eb3b534f4dffd0e0f9ea1b
z99522e16959bc1f61fa1dc4a15fb93af60ed86b5a7819d9b5cf68ed2319afc2a4b60800999d601
z3f816b28c961ef36fc45c5b579222924922f5e3cafc0026e44b9f84be7e514c8c22dd49de2d782
z63ee04ced273cebea18a942fba38c41af24fbe19ff04ac11d0f52101bafae8914d5db2f6aacc8b
z2fbd1d3933e083cf8b92003e23e5c9f602665160d6bcdbbfba92ee70da3df65816561bd01ab6a1
zeb6cd5d28538f610a0839c1d6a4c550211961da16fc1a5da7880e0fea4dc6a00f884a18b8b10d0
z5618317d6ed5c6b5bb1acd1f3b08b337ce524c9da5a645a43211af6d92e64f4d7425fec3bd0e3c
zc27f775c3baffc4f2a1f7e0e2ad31242eee3f55f6d998caab49f4275c06dabf381ec3eca632093
z235867748cafb34be32bc5aceec744a8cc8d0d10a382cf6118673914547c126a623e563315bc68
z0c4c3bdb7ac5c69cff4f11c3db1736e2c9815b1f91f474ae6b13603491e5e1e490e286c8b1536d
z110c4f4ec3918391bea8a79ed8200164fc1218284e91b71366b9d08d259e4d2db607811bbae6c1
za3752a48482c6bd35a8d63a7e4a3f8561c7f6fbc4185521ddc3a02cc4f63791558c68a6e42872a
ze887cb4c8c0ca1691103fa64bb4b6ce2d81893e0355c9f30e0abe057148fbfc4a5953f31c7097f
z3cd5a006a12695340c96f2f317da86b0e22ae33c729e7600c73aa5df8a02e72335c97d513acac6
zf99edb380193b1f3d92ac7dfda1ac808802deca878ec712957289745a327cfa86d1aaae2e32c39
z668084d2d2e023a22bbba6923a6d9926ec5e721be1527a8fee58fdd095b99a78f1eab577ae66fc
zc4744983dd75c75cf50bf0353ca415ed1378ebff17508415525aa22939056a3185d7af346dc86c
z0bc53d405b37f4de89d0e24d02255f0f7a2dcc5cc02375c2c8afc811c57ea4788f93c25101b5f0
z7be513b7dfd5f41fec6a5e8554311ae1249811cceafc9671048c8e2698b4e41f81d0c965a46fb0
zb975197d19e1cb36fc4975cba5955d514d70b86a2e991b1619df3de9abe67dd4848e1dff82ec95
z8063ebea535c72207ee3f56ffbc5258d0ac1226643cd860dc043215aee122b5f9a65944e1c7931
ze75982780b08aa27c8effbcbafe00aac5aeca3a398100a9dd6958bc0ec31523397aa2dd769e421
z9be19b50ae7b4fffe56444624f8c92b59f664817cf42b12e0f838acb7306fdaa89ec677920e96c
z7aa89607fe582dc1f14060e7817d1ff7c546dfaa8f0204d8801a431ab3f0302d9759bf03137605
z79470be6c85ed74397005cd91cc7ffc37da6ec7441b1c139a4e484013cad966d94a143bc206286
z43b5ca92302d8b032cafe182ebff7e90a3947f3f65f20ea317bdf82f76166d862654c05a3bcc9a
z4b86b384a577a72e4fc36006babc4ef488b1592b07f90189fffc1d2307941c0ccdc62b9c058f3b
z63ee6da36daf40e610049711cfd30edb3c0d209b2f93c5472cda01ad5baa926b2fa83af8f93f43
z6384215c0f4c90d2d23bf9d6d6cd6c779974e9168a586036a53ce3c3cfb458b40374da419cbe74
zc9701a8721ba3c7def34cd10be9786c2f655ebd58f81a10f92ba5247f2fed0fc5b454504bcc08e
ze6650538bfe65e356f4ca96cd5adb8d7da729d45d9287c1336fa5ce789c4338aa1ad6e143591c0
z5f5ee083779220cab466eb9b524a026b1ec67a0d86c6e73499de81fdbf28e62283e2b60081753e
z8f69d01aed6feadd74efbc4abddc8b3f4e0b316bf24c8b2fec858027843215a50de9962b4bb92b
za6a7df5d7efe06a9e695893a0c6d3c943cc473ccf313157482e6f3570181c6f688b36c1a72e92e
zf224c890196bf4b5b77cc39d9c7fdcd21131ef18b95890f5bf223156feb008050b96088d32a63e
za0f70cc8c774763bee880c8af8176302493431b70b9a83fc4c48b888dc96e27ccff60a6b3317da
z6ce34d6f50b7debf8bea655586b17328b46484911c913fe2f70ff400bd6032540f4b8e63b9ca76
zc9dd5606d19b69eab74d2e88b703c4b084bae8a43aa3f562a26a6d5cf9dad234743eccc84c63b3
z0baa0915a299a2346538173f99663705ee6fddc20dacc0e066b839be787c088cf35e0d7fec9752
z122775b853c06aeab1f2252306700ef1e862b96fc41b3bd68ee201ce527fc75069b2495cf41526
z9cd3dc8ca9ac5b4f8b0948de5c52e8435e5cfed1df0b8f5831b3aacc1b9fac83eb399613d44bce
z7d5d74813ee280535a63f0f6b961cdfc4b58260d5c430bdc9ed26a6cd457054390f6b92fc073ad
z4f7dd50f983d0ab1a4a670f291be69e643bbb15c292bb5ac74672854bc4eecbdb3968394a2f255
z3b3147b258a08dc0cc76c7f6fbe9588529ced122e3bd7043f761d7eaec78007720ed946dd3faff
zb222a38e3917244cd0f1cb67f7df3ace621436ce5f427958df1a8017a2cc53e887efcccd0a6c59
z372756fffef5910ee329f9ba651df84aae231435769ed260beec4300c7ae2d1fd8b19443f9cb8e
z8e46b51ddd6249016fc4ae1a2e68fad3010a75057da2aa6046930d0072ffc28320dd2d888da973
z2e5db86d5bc17120f2ad26821be49375edda2ad69d9f94d95502f2f696b48e33a1f754a2a3b2bd
z8241c9f9fb9de20cfe569e00b6210c2c1ea702377af71cd4cd00f2cf145a528cf5f734a0cc2f28
z7376af4550f5f46418b471117b5e15dd982e1aa906cf4a7575a54fa9353d98c3d6c680e32cfaf9
ze9bcc9b2ed4828197070ef2010518d4f6763c56332193464f507f5443c881f3c6fbad26a2391d0
zbf4594582ec8e3987f50dbd9e59b0afebcd11fd54843c3cd92db46eb4809aacbbdd9782a357f7d
zecb3a42898bd0847414f1517350612ecfb96cc24384c51f38543b596eb6652c7e8a4ca6fa5139c
z24371141b97c7469aa1754f65dbc2535e9f6062199191a295230e85d78dd610119ad1265ea19ed
z53d0f1e92b82ad9e2274e7dcf142b495f30e8db52e7ccf894370da45684c1a109e18f63c96eff2
z165f1d960cda1b94cea23f181d0c6ed34b1cc04b9b18a6e8713b22eed799f25fc2e8d3a99a8d0b
zbc8d712f8d49322edc12bf4145e68625aaa2884361af30b81cab3c42eb776dc4f0b5ce525f006a
z99a92658fbdd84d36e302a78c7180c663080d069bbf2c5009a228dd9de8c3b26946aab334da5cf
zdee272b796740d2b68cd469f9ee704d779fda4daed33f03b97bd199739b086e02e3088b597499d
z3b178255837336a27b6f9eacee45c7c7db1843afe4c34669bc2b91d964bcf7db128e3a8088798d
z2bd0e86ecc75c3bee76c31c02553eaed033fb7f7acc6a0684185ee92991636a256a6298e389a6f
zfc9b70822f208a5e89a6cd384f8cf89329e3bda464a71c6aeb0e72c26fb4065432a5fcc9c6bfd3
z0c47128dd3b4570e5d135d12061b52db538c821cc4c7fb9ea2dd2674b8a8318f8a079dbe692dab
zc71f7a556683c52cabc5c2fc3d1bc5f926ae8064966b53469aae99721c29695ac568cec5f542f2
zf3bb136a80c4fdd8aa747292f7cd8aae33640557f23e1de8fce69ddaefa1d3636efb751b949a8c
z17271899606535610544368c033170f56188aa50464c0188acd83c21f0cac017e99d164fa859ea
z2848ad6ffdad97f4cda459d6439f109ec36f5af9cfa4100bcf9d8a6c1a4b0592c42cf31f094829
z552f31aa72e8e5a5cc10b33fe315a588f0dee3f128edb4001903a4794034486c068fdea0599d3f
z2e54fc75b35b31f34a9e164e178db67c8d2979bc7259ea27a81b6b5fc3bbe3b961f8b12214e4d4
zaee90b437d57c3c024195823a131626ea1c97c708f6e8ffe4702d5ff3f60f19ff6c5028018c626
z9566d3520eae7e00728a3d4cc45228a8b43cff124d5f6578bd48c7878fc8fad1b3de950fdc73b4
z404317ade33160a0186400cffaa19aa29a3fc2ad887680e2e658bf318700c440929536d79669ac
z42731f78014f33e4e36957a2f84dd3ac420158d21656d0a94754467b06d54d6e219f29cc6495a7
z00fb6c634ba8e1647af71e45176a6b0afd73b6b0123581b673929b054a7a1be7ebfe09fce1e045
z71cf01f8f3eb1400c6c94aa2575d0111f5bdf188d4bbfe8316e2f5d86f182accfd77034e618c5d
z87892350ce83b6038d4968a08f41bfc0f5d1dc3b86a09604d26f6cc882febc51aa16c0179464d9
z79db72c746068003cdf004a7e407cbd6824d4e72315a06e93db958b936dbebf754f7ca7fa82dcd
z7f9217950454e62b94f13ee11cd5d79d1bcbf6d5bafa795fe0fa89d163ecdc90df523c2c2db4f6
zcfa92f68bccc3e62fe39c1a57f5d3540d30bc8538a07c6396984c24fcc3f7dfaadbeee0afb331b
za8cbc0b386f8e7dcba2d487a6f6fee6507bfc90dbd137855bd5632ab0ec27207f967ba7e7170ba
z5b530d63fb819ff006eae82e46bd5df8e4034a34fdf261234a2f62b292ffa1778ef7e17fc39cbb
z11047a7a161a25a9078f9be26ea16a9c5fbb920fe00fd146d65f8aa155bfe29628b5a7cd506984
z5eedede2dae37a08d6c87288caf434233312d0d694c30ac65642a2643175bc29812704d959ba93
z17dcb16eb15ac76155e3a17bbbc45f34bb41a1d38114a78901bc7b325ab85a9dd5fbda64ddf7f4
z37225225a844bacbe64ac52c021987beeee1650d2eb209373dfc9e7c5cfa0d8b653d689ef0cb1a
z5f0da80680863b014df163733bcbd81fd74144f53907b47a7e00ed1c090606c40c5b22e2c056e9
zb399cbbb3756a7dbce2743629db95361ff8517afc72a81452c6faea562964ed009648620d94f96
z84a6b2e114c41fe7841a033230be0519b811d689a6b9a025d1c83ebddb7619dac61a6f8132e3ff
ze55edd8f530a027b5aa12604768846261d51b5d72d22ec2690433ce67d4efa8809048644790129
z880ffed242668ed9d6d437ac6595fd5d329297957a234dca8b158dd88f58dc07da543ea69d180f
zb42d46668d8097fb6b8b800d44ca9506f0224f6a278bda8e803282da9ab9325b8809c52dc88bc3
ze3f3fcb92ec8adaea6243f69824202e13db072592917f4a81502bce2b890502a627f708b200973
zb0405a3cbfd18b38d6acf0cd71de43068d52e36725121f93f7fe9b45a7db9c0baa26e3de8aee56
zc1d54ac2d0860182828326bb382d1e426ad782116d4d9a3de9b877067c71dc0a8ca299d3c09a80
za978dfc52bcf0ec47afb83a9e3ff1544f8caade348c6268b9ed8156cf568a1958c80b70a4215e7
z9e386cbb1bfe4155d46cc7fa9857431fa22cb1cc856a2ab4061f4b3901b29f1ad4d254d9c95392
z67af72c3d5831aeb33d196fd7ed6f708b2da07a116f53b6b8cf4856e7d52e3cbfc52ba7a396c94
z7d3133843d704cc6a2e27b17bfe0b7e8dd368763706706b571919adf5659f1ace782824dee9064
z9436a1738724acd63bd4b1835d91fe6e578ddaaeb7412fcd5f48fc81bf1022f1ea455f47e88890
zf1523b17c7f1013bee7f107218b157bdcb3ec76ae2ed1091600f43e0d774a31cdb3e5752559c3e
zae437262c736d89524d380099f66bd793b48dbce24302c96fafbbce87650b966df8211a7d42a75
zefb5554d831d8834c4aa94c6698bc96aa0425df825f31b2abc94a891ab93633e878e46ab83055c
zaec17c2450e734b3ca495218327129f9c3fcc56ad303e73dd73c1c22bb54565e2f5b46cacf939a
z160ca1f99b485a91fb21bed2e6aa750994f1f2688013676021b6a08b3a22e985a1cb4305e2b986
z1cdd13c4689f6cf8054b75184cd38cea91517cdd917cac3f3bcf0801622a2c305973c07986aaf2
zf2056ca015a77ece094f0d741253a5d812851139c1ef607b9ca16fca2cd673d42d591405a96cda
zede1715fcbc7c08dcc239cd4bd1d99d31ce8f3fd1bab41dae462e7f1dbcb8441ba61dc74b47813
zb054cd49794e182b31edc3c56e45c1d64f2b49ae33046e354e88b406f32141cffd25ea1b15638f
z6c74ff0ff75bf56d555b8f72688197e4425122c7f809a51fd0b9798f24055ca04c762722d6bbea
z9c19a32c56bae6f8a9bd34de62b0173d5cf3d38bd6d45b23bb76200fc94dae5ec711ce37d031c4
ze385c1157e3e86b3c985f120ce9a44500314d9d9a8990faed5ad2afbb1f463f721334f74f9d1c6
z1923cc3a61f621b9b365ac0439507d5093cf3784c1d9bc62254447ccb4906690d171ad310367a9
z5871a0c55f2ba3a44b65a934ae7d556143d670eb0973ddaf2abbb3192cec80cf1c44912f55c65f
z5e032ad4a1cefa0512f26ffcf5eec5cd2c7946e48ae31d437e903efecaa8809cfa0678d677ae4b
z2af11ade45547ee5651e68a6f1bcb3bac28c334885b37596dfe35803e1a124247d89535d2911d7
zc5d77abf12df924bde7b3bfcafc2e58dbc14028c87578700417798ce79a7f9b17595e3bd74f35d
z0d5a77a47350f7a62b2d8ae502048a82f45d3b5650db21b33b19d80b0956e22aca561cea9970a0
z1d4f8de0463a6b68d12e43d7cc32ba8e5e1cc058d96dcbcad6ecaf1c2a4b164aaac31141182874
z0db8c8fa01a842a887d6b76f24dbcc895772f347aefddd8eee24fd47cf833626650f436ac87d1a
zf8f11f79812ed44a78ccc1349bb0e74a8cdc6e5936c562bd3bb6bd201e0b701f41455cbd53be9e
zde56d4af4d5fcdaadc1c4e20850ae8abcf8e289c4b6db0235584463d23ddd6f1017c82824580bb
zfe17e243fc8d98b3c637ff62ef657e5e9f28e76a334210e6e6f2b2b17b53a6000d665eeaf4ffc4
z2b50f487d423cc3f0cdee223981b4bf6c6ed865e92edefaf04f884f063286435153865c695b97e
ze41a8a0f46377874372fb2ac36043ddbf8a89fe13fba5970d71d9baeec49b512b69d5b5a120c2b
z273a61d3d1c972e93bf8efbbac919f3b0e5d28c173bceff2e113196fd8ebf593428cc653d82c24
z0d046f26d882221b2ce0de3367b149c1379c9bffe92e289551300053deb1f664185dd165ad88fd
z85547c913db782ca958cf0c9e251afd6fce56ca8d65b159984299bb3485d6a11277dfe6685d3ee
z7b020e89d0687460d046cc86eab4298220c21f34180a2f7212a209f73e69cccb4b473ad8fe1abf
z30b1cf8c0dc9b286ec61aa0c34bdb70d9816c1ee36600c99eb34d1e95fb4cbe0a8abb676f76d7a
zaef5a92a42fc677b3e0e20b3bd069a55c297b61257a5c919cf1cc696fb657b2fd1819f9eb4ea12
zb36336dcb101f38b5609a5a001793275eeeec0eda009c253c50cc240621159c67571a55c636212
z5414c62c5c7c3b567e815af40b48791580414cb0cdfda9feceaf12544b80e98f02a6a6cfc8500e
zd537d147c20dae6b2ecf4c7034ac7aeea125d35bd161591db5ce425459fa2776c75d8a6e209db9
z1b76d4245f6ed3a0a7e15dfe488502153935e1c7ae87070ebfa9f07873b35652209cdca6f30175
z9e6266f69d77feb3f862ce05cbd01cde99187a3b11a574c5adba353aa825a23e2f0a70d29b5d4f
za40fc30079b283e94ccab7d4d594d3a79fbed6d65b2e2f2d157873927488252c49317a8e1935b7
z3cdb566b9d1d13b6c9d6b3333a55e0f2c8189da8be41ddf372f319b0f3576089c2418616f5e101
z9a6e0da816c1a7d67bdff3618a99c61a7adb0c661df6da072be9ff85a21b9b830ff0f52be94295
z51ae019837caac174f22a92f45ab6b5b99a21cca6671c22e61e63bf108a1e9460b40725d368e1a
z021c20408d919d91a68e0f75c3aa6ef0b6e73853e004d2ef52461ee6534143000390c5b63625a5
zcda9b3176b9011c0764d6756ceb7ecdd442aee282d9d005cb43b31eded7c30b7531ddf2fd21a15
zcbee953ba40ccad7daa0597189d4a2f84c271edd18c3410e474429a3b751d32b861641e30e91ec
zb1c2c556f4f04b2e9c984f3a4a3ca9a1708d0248f8610ea86c08ec49bf73603c97cf9296580a45
zabd9ffbfaa9bcaa148d08e8bd2b69efc1a9257e6e1a0ce13ba2b23e52cf61dffcecd9dbdae87d4
z73cd5a3964bdeef720ea47e971ac69646761e06451f35a7f388e167344ce6f3e5cebd0426c0367
z57098800a8cd7ae18fab29a5928bacb48a8b74b4f45c28ca91a0ea894b9f8adb6cb8e99de0f341
z58ca3e9d62a84f09390c4c9ed824895d6d5c12a875870df87ec8fc1db6a423dfda685f5983a53b
z7e298a09aa3c1e2a03cebfe7a8b0c8a161be429399b6a9ad5eae05ad2903bfea14d6f08feccc2b
z67bfa83bee6816133d4fd0a5bc9a8eb9e3f6e8b4be7f882f6a5b168a92569f6340bb3f48798d72
z177c608e8022c72fa5037469aa6ac9d0f9a9782717deae62bfbe1e9ade7a1ef6dca4be43bd31fa
z38ed75569e7df7f4915b463eb3e6815b007aeb63492bb382186b4bc3f9cfb9264355bdf6048de5
z241d42188559498c1b87c33afc4c5c033ee624e32539740fbbc8dafa9c5741ef1824125633fa7c
zb2afe42e1c5b6c033eed961af4bca5b5dbb837eb2bfa8d93c90ecdb1c2488eb8932cfe10b0de45
z61a29e2ae559b21333c257ff4e03efce61f90be8be9bbb6099c2518f646d3c1a0e877022564133
z89e55215b61878f21e0929883a78c4e7716b8f6cd9a54eab066cc901189fcfd06bf5b8cb42a4d9
z5a1ecf0b09a6ded1f9867bf3241a53a4ecf9c9fb17ef1804eb1c1a413d827fb29931f10c11f68b
zb5efa2c2b7f257bb53cbab67437414ec62c566a27ca0c78b27f2e58610b27ee279066461682822
z7c987a35450824bdc134116ac8a1ee48e01698d726ea95bcf88154e46f3ad7aa2ccba9666ccabe
z10bcb3c4a935ad25700190be6cc27670725d60b5c48a0a1a6b040648dbc23f5863a33c79dd7360
z05b92bfb550727e6766f15a12df5c571dbf2839adc4b311f60b9e0858aaeea7ebcbc80e4e4e23a
zb128726ab9c6190179ff5e302702da6b8fe9476cffa7854e7811358681375279fbb84a7dfddd6a
z539021f4422f765c784148ec5e8d0baa8c4ae656f270998397172c704463fc3c9632a7921e032c
z62cfa8d27a92e95a3a4f9473ef66816855c6988b817c9834d03e8eaf5829e64fcb44fada5970b8
z00a483459db66d9f6213307db9466c7b664cecdff48b514710c2631a5eb58ecc251c8237aa643f
z9cde03fa71d14036e579d12df6dd20ce81e12b46af643768b02af9aa545fe6faf5eb6326c04871
z99affbd0900ff0ee38b106a9dab81cdcd72472851e4b42b0623a377c6e70c0ba5b0d7ff2552c0e
z302f7e7097a487be1723ec78f4cc382e84d14329ff53c3fe224ab92ce120b6eeea0673573952f6
z6a2d3bfb8002b5ad004adba0f10472487dae7bb422d1f2cbbf81aa73990e7b6061908e7787e97b
zae3c282504d1aeb7863f2a5a019d659375791b66a57bbdb0b38f4598b6afdefcc51b20a2929ee8
z74df665d8ba79b8b6995dfe46a26b59350222a727212cfe1d4021d8fba1f88145116fab6938183
zccc7cb7a8a68e3b5baa89c541abb6c98d352cb1a26ac5b3e9a09320085cae7d290f618900b92bb
ze96846c51cb128d3e0b14147d324108c312a3eace836ac4091d451ced53f617bb1fb326fa09726
zd7ffe65746ad65a957b1525f4d3abdd54344295cbfea83b8be6bbaf26fd9af2bb27160ae00bce4
za6646578fb26e0eed69de486227c7f294bd3acb15029beab9a04cf92182fe048af733d642d0e81
z491f25cef6e9644ccd058755333458f0ba0aaa43083a0ffa558db4977f5087ff38a21d400bfed1
z3ae8aeefd27c3f93b461c309cee9e7f20636e690326cfa211273e9d661f04b344f1ee314d39615
zc23a22c0d9251c1cfa088965f7014bd0eb94898a07e47e8d69370bd7e5ff163f56c3cc9862236b
z49e375496751d896b2c66e565907b7e6bfa2934283710e5254b31d9776f3ded4cd99705002673c
z226be3409ab8307125efbfd859300351de9be3aa6f0de4e7336b3b8af416bff935240a18c96041
zaa80afc8439e06b2629a497bb561aca282c0392b49151bd9824c1299858fda99acdc08d77701ad
z7fbdaed8fbd7ad8d34130b9d8f94d7f6b50ecb763041d2dfce8039b83db58b489fac0f95721e02
z00b689a20439a2de69b588c1917e55fd6a44660f2d940fb7259300be0823a247800a3aae5ab61c
z8685c86a8e4c0c549348963468012c6a5e04b8b43b757ace56462e44cfb8b7e6ce504b1cbe833c
z9e6b9c2c84b98ef4e3f3af92abf609a6d7c7e1e45c32d93c7a36f9f1bf7d18cd346094adc4c992
z2424d96dfa63603b9316234438a4e604c4f076e735f102e38b386678ad26c727115d501281bc7c
z9b3af2d6e14fb58de7ff4642be05f35eb123adfcb7197f14589c994c0f2248853f488043de4ca6
z409d54cd5dfc6c02526391ce55d09643f48a708f3870e5cce6f3e9561462960c0618d1474ff6ef
z80775631c8acefdca6b5df289721547774bd5b113184bad49ede97ca5bb97a6d55a17e79542b18
zab73de4eda5de9a9a3e89d7f865fb703311dc15f88222c3c834299626f8a4f367f84b9573d939c
zdf4e5faf23614c42f02a22281fc3d3581a98a3a0119525ae81b17cf13e371deee395e901e55531
z0fac2582f13687b9892c9989179236cf240510a2e73ea8efa1dc0319b950c68c7beb888da8d5c5
z66a5435a5c40b2fa6964d79a416c0e7c2a4df288719cbc8e91e950272c3d52037b511055c91ffa
zec550c822bced604ca7993f377ab9b485083e90ecdbd3e3e19d12cf704b5914c3aa9d0d168cd34
z8f145fddb95c9c1f38316b921a05403397c68f2b9527d9e8b8255e27a25aead683a8b843a13748
z89fbebf2acf8467c09ca6899614f704618128a081614b5fac743b524e18f48a561342f40228d23
zcb96b3356bdc565f9d80239736bfaf22794325be0a419fbb927498433655c7c4d55c6c1a5ca0e4
zf9054c622c66dbc8bbe2fd9cf8c3c2476655d8a1f46601c10e8df4b558960b0e1d60221a988946
zecc72d8f313a54b968f730ab08e3bb5cf58ed4f7fc209e76161f336cfaaf3c17d896ebc433e642
z4ce8a8400578055fb4e54a804309665f10d8a5797d5e640dcd8438431715a4da3a7aaa55983ed6
z501d5be06d19482c7898616886c0244153c8b17dd6514c37bf8624f11df198fc00ba40604ff08f
z5017d4395b7379bee5e966105e6a42faa080db6728fdb1cb05ae1083d53dae83c326990026cf37
zd7209f6dfe7b957035b612cc0ac317d06cabc174cfb846e3059d6ad37b83b54976cd86468a8556
ze83c21d7273c5c503bbbb6fbe71f4a0b6e811decc2aec0ec81396fe96ec41cdd54c8d052849b9a
z50c0b195012715ad40ea29cb91e914a620c4c00295dcd2cdddfa2ca3077bb47a75b32d71d8b1c7
z235e00ef7db78de58290dd088abe6e989cda6711bb3376715f2e94849c280144d7a07862f49f9c
z06a59ffb4754583fe1a274d60a5d7c62999d2ad36f5a2aa987a51c0ca42fc2b938292903a616ae
z89f066462f6a8a3da7dde7270dc2738025752379e456610e90c80262f27241d80f9dbe14981afe
z13a9feb28bf3de39f94039c7fb56e15a0a7732a69761b0dddde785b983ac99068cfc9205237370
za3837d03529aa3203f0349e66108ebb937e40dfe26ccc167d8d3eda216d51121c7c93c0277a475
z349b32de957c10be6ffac31baf37bfa56138d9ea32f24fc75ef86fda3a9f707ac785e1fec8d95c
z620cff48b03ae34a17b0d3a4d7c48981d41c7883d1d9f1ba031227823cf80844c1cd3e1785005c
zd749a5c37d6a86903068afff0b7685c2061eb31bf54136988adf23e77979cf6f4515018564ef8f
z4ec632e9550ef5bdb26fb29c5ffe50f48d5b3dace3a97ee91ed99c99c2e78de838c2d6d95196b9
z0f15e9c7cdb0b3f2a65385f8ebe2ac2c132e3c92edc466a07d1f7138166d81c031d1b8fae7b44a
z89d5d0420499864a574519961765c78feb6780ebbae6d0c408f0f312e4f3b2736acf01868e1163
zaafd5a188a727ac5e5f495ae8946715d7e30b605c817df06b8282c600fd810abf6453d213c706c
z7f0a4d2f185cb0fd6b1992deb45c3b23636d27bae2dbecf1096f9ced9e0269836d27264fe8f12c
z044783e42be09b6f6dea094b9d3be97452ee02a8d662a8e4de893f57b369ffa56b72897678547f
z3437ca42c5d5c857950e2ee4a60fac463e53016fcb691f9417b28f35a35cb77b993ef33d57adb1
z0e69bd527a53dfc764de4d1a22eaf77e776fab856c1f76a5d4665785f292fce1bf387ff3314802
z7cddef583260dd0973a5e60bd41ed1354eee945b7274496bb32131b83d7c6662518513508da8fa
z025d69bd5ca5292fe25052f1e1f5e6ae13ea481ab25845400bb6aaf116832477d5f39b0b18876e
z5678b14bc67219f35d6f5947f16faa5f8cb9d5f930a311dce20a2b87bb4b62b145dc5f3d827e02
zca1dc9eddf10ecee226e7e28d97f818f0645a47399148646954f15e05bca4cfc361a18715a6b7d
zd9fe1162a7efaab5dd0d8149ebb0268ff4a23a05c5cbda8caf1314dd53edd03188c60fef0cd6bd
z2306499ba72aaf406b2d541680a150648803d3e69c272d0aa520f42342f1284fba08a5c9be54e5
z40e2aeca39ea3307a5088853b38c1f103f38aa343ff9c3655486a131b18ddb847c3388ac879b2c
zc91b0ac18a4e0582e617aad28fc5db150e3d0741747f11f478cd88c934fae573da47b6a62f9052
z5c68cb12e30698c58fb38a3e15e57db08122763a8000dec744e30d3b1a2c105d3382a1c86f9a08
z4d795b26c700791d6792b409f20b14ffa940a2b887e85924a433678da7d0dea4ec9f077ba602dc
z44ae2ae0e98593365af2a04562c4b75219612c057e359b3c3fc4037e91f8b4b7fab439ac808886
z5b9bc0c7ad7861791e2a25fce324423cb108c009ff007d682d6208c5461a08223db597097af244
z26f186d7f3661cb4f0369ea890aaf27186238b48e95655d8890f92e08746c9035e732ef85ea8dd
zb0e4bee31b21c6c21b29c9cd8046cba7bc50f088d5d9e9e8fe54fabad4a4093900232ad9aba41e
z2da8dba7a7971fe36ba5bf4784e15cc3f4a91364ae53be740e59b7172ea9e5bfcdb88339c4629a
z4d6df13109cc72a7a4b17a5989c1b85b6662ed9df7a02571097c61172961ad16e01415f5896112
zc497ea214ca7584517ae3f2f6d6a2c1c66aeed5d2a790497903a47b35dde77831303cffdbc0a6d
z73d1166ef7699fb31fdc9bf1b1d587c3aa6ffee2a1044b797d613255d5358f631ddb9725bdba18
z3995c7a11c664c5bfcea8897f3e47c267f94050c1d2e20bad2201e55b377aea65d98c294469df5
zc56564544e26992b1482951780ac50a7bdf7012dc60649802b1e6b815c55985f6780ff3385d22c
za2643e78939f8c19b9bcfae113abdf372a3a0d2d67428e6f7b7c1b9c931edaefefe1762b5cd9de
zdd30123098d877633883870fd7751ca4d35d8347006b5e5d9eae0da592c5d9c988d69979a4af55
zdaa0c499bb2f33827fd9265f88a1198facab3abbebe01169dee836b1c47ed36e3c920ebdc31b26
zf9898c89494456a7a00c6aa729897f8c59178fe087745e804d06d328115dbf0e952022d826fd38
z8346c64ff23199bea39ab939fdc2bc4a09b1db4ebbef5df4abb18a286a4eae30fe0600574f3f51
z3c9e00772f7fa8898252b38c48a14bcbc17cdbf32e3544e46a0dc68d4d37b798552abb62c63bef
zfa3fb793c362a6dc96db003baa2a90450f3cfa593eb23c1c2b1da79578fc741e52d28fa6153da9
z2f2eb494ac4fd89b95e6e355c2705ab498cde9ff3e0f801cce240dc605820ccfd1e2dab142e805
zf48ef76dd092c3961bba67cf0aa32433f9827b2bc0c9367dfeff600f2e4f5acd0de1506e73a07a
z61aa244d0d0097c9df746d8ad7e13ea4e32b9ce0e32840be7daac7f0ed8be6b2f0815a4b1ed7c3
zd1ea380e19ad46281ec317d4295579afdcc37ad4ac2c48261e3908626cd8e8b1e20a4c9c5f69d8
zb40ea68ba6276eb8c26e33a8db771992a78fdb8877091d450d619ffe5bea289b8ffd4e8900347c
z7ab1a373b9c72b6bcf59d388503984b06ca488d7f304903e019537e93058e978b5a3c6ca63f699
z4ead49a9f6613dc2f87b23e65fb705734766b72dfa7ae39927ddd29051d903a3cb8d33192b8e96
z854be8cdddc07015cd2fe983965ddfea27b4e0886b0bb8880f07bc136d6d49cbc70dbd9c6d87f9
z4dac2e296fdbb97cd9db132e84970c5cb7688fac087c570bfffca4acd46f9c9a780ae6c7ee3962
z96ac79117eb8dbe65fea77106bded7b0f4a050d9e93919cd1c6543a812e06404ca77b1de98bc11
zc23d9403986606db1275f40976a7261cca2eb7c31810b61249914f1f55a267a40c39b94a6dffff
zca9fbb58a229ca6443749d9796ab4ddb16de2db8c59489a1343726d46567ff1b95cf41974d8fe1
ze5e56c5f48294c03f9387c00a0a654c633aa7e6a9e96a4620d7f9caeab1a417c648b77900ac7b0
z3898740f722dbe387c16ad487eb7653643c3db5aaa0f0aecbf5cb217166e5760b6407b861c57bb
z5d8708af9852882342f68be988ff12a75eefa6f2a3784ca4dd2785b463aebbdc6d0361123e3ae4
z84e316c3e8c1918affc2dbe245f3416b624db45f1c44c8efa3b77d4f1b88111528eecfb373c383
zbdb23674feaa3eeb51a72c9d1002cb0e4fde66bc582029b1076a89b9c0cb7919c309e686f4e238
z69c4fed5b99e1371a85e62653e1618e2e763c1d941fbc3c990243bf40c69a3ca4f221a006bca3a
z12c5e9b382b4f1e3551f3888429a039b49b222cfcd109806d54449e4ac20a1db2207da9319ee03
zb9a37b0ff32a6097ceec6e83e7ae3f8704bd1c9597c47ba2f623a7d25db3065b740de19b2ad7c4
zc4637687007871341d6c29f100112f677b3f99d65881e49250e4a9347fbedbd858fdddf8aa91d6
za63f8280057b32904319bae709b05ed0058a686c06c60160b4b6d06ae7f6c88f35925be0d85cb5
z008dedf122437311ecb22c372d21a42a9e9b6efca3a6c75011a96da7e4ea615bd3b8736530d293
z67567b9c2ad5b19f1ea316f25a9a512acd845af0a0ea74f5198f7e2b4187ad48bbcac67d5f600e
z2f61106fba9bf04911c8d1ddba7467a4cc0e3bcee3e1f2e69c6bb6aee79f7ac6a2658189abc99a
z3a47a2431bc62a934b74784f2a1594e7dfeb7437f1e0b4922c414963dd5971142f98aecd5fbaab
zed9c2b134f7ce2c4a5fa0628070f67fdef4e01c9c52edec8652ab9a340ad4b3d1c587014f69912
z638652fb387cdb16576e328ac8e79566c58f844fa7cd520c360cea51a336c5c381c339ef26fa7d
za73e1a55bd1538d54b468251de23983a7c0a1af8e2e79e4e0580fa1bd746ca6fc067e69416c9c0
z14d30eda3ecfe62e6c7badc4401d9a821c6dad9c76c30d33c238962a5b2b11f656e2fbd613af66
z77e0b7d5490f202e7a87bc6090b1e4fc2b4892982171230e6ad342563bbb0646e19ef5a9230e6c
z0836630a9d65b0bf860a05bcba128a9ca7b4aafe936c7c8a735904e7867f704e29944c90cc378b
z018f805880247cbd5dfae44a413d9a8a4398c0a98c48662b6ce06a6e01c11609429d6e90c54b3a
zdb37d0f88405a5022c479becaa14eda4a6b01055598578f2522308dfa179972c3085d00086db86
z4fffc0f36e88f7f5274ff5917c399c0c609f02c58980e53b0d1101348609d86024a46e6e36a79f
z5dd7ddc5bebeae7874bbca9cb8e4e4140575f0b9d9e2010fe35593ddac462a6919fb97f6ed34b9
ze909dcda099b26fb16c0b4609a1477a1b1d4dab0d5b30cc0548f53cf2c5c5ef4dd955cff5b7d86
zba1722c6782de4e7c2cc914613eaf7fcb829914c657439e91ac201bd54a7de3f4b365eab9cf0f9
zba88431adebb952c34ac52bcf3ae8b3882092a671bfae2bdb74a57239ba366450ca6fb39fcfa2f
z15006054eb534a9812a8a57bfe4b0fbc20c2e5cca33fd21c4a5316382a15658ca1f3aa7f946eca
z9d6f70e7d9b929a96d0eb913087f08601b466929cdd22b89cc9c2e30772cae814ec0a44fd0111f
z1f9a1a4d7c85c5e9be718009386f0ae8c6394387752b0e5ce09c3762679d4c56c7940cf6958bb1
z2e3a5a90a1956515c76b8884098953558d2f9e068540f1c215f180d7548a64e577713149c7ac3d
zf24cfc7930aad6bca890e6b88bab2dcb3d7e3a1b67d6ff98889e05a91c9bc3366c64070515b446
z13b4980c080478599d75cd0cb283a95767d4f6016e834d0b14fd4cf77c72aeaec826cfdaf7f8cd
z8d4a4e7fec5e97df4638603cc3648650bb36ce7574ff2a09ad1f5b7d795315ad98dc5e0b9f4f4d
z982a2edcb38d678797ff30b9bd7d3d8d9829f36bbdd432ddb0a19202605fe6a320e4c0745d7c00
z8dbffa88ca9072443ddebfdc171654cf42818ea30ec99562cbd1a5d97bf3d8b95f452a1235befd
z7f0cf7699dd61ea7a36d33661d969c541c99dd7da77b8f9ab0312c6ea7d22e23000e083e1423f0
zd5ed6f37a7657f5c0aecc34347a4aadb22a299a43c029f719b371b5bc90ebd88e6d6e172475e84
zbc745188b915ef5ee82cdcd074c0348bb982c6f2725f2a4f12d646e08db4f524a5d8fbe067f0ef
z05a673ec0f2ba82614a8dfe122135a5914df5bd4aa99735b8435e3053ba1f5cba9620c860f705a
z5df5dde1ae6648d5ed633b5687c67e6aed8e022235ccdca14aca2d15256c45c05e8fa4d2573930
zf0cee513992b2b61e968fa83bec549fefa057fd26d3292d59029f8e0bf725bd610f0612c14721b
zd552b5b25837749d4745806901082a516e3399bd2174149b6931e5f90184e5159cfe05145fc763
zc31bf3b55ff4852efe31ce3b051395df77207d4298723c2bbe19d6e530e60ff639a0659b23a5c2
zd62a070806db055403613d9a0a687b879d431c252d7e54cd03d76cfed9c36bd5b64edf1faed8b8
z2d3eaf8ac02bce6fe7d0aa9530016252ae0db712a96bf10f1621b47d32ddf1c1d88f9444350b6d
zf26eaad0163bc10a3a82506eea3efe55594b17bf2e755309661527812feeb44b8b4e302be2d7c9
z3d52fd8724b69554699074250f15b8d95280509cf05527b3185259a0b0e43a0a2ac840a8cde982
zb041ab8b7aa1d1af207f3a163df1c437c996db96518ae83c1374e0936339ee823c495ddeee4f97
zc833e4096baaeb93a807ca74abfc71790ae038777c5b20714db3ebb1be3018d905bf0ffaebbfb3
zc8fdba8b3cbe52a6d4a4984499dbd0eb345bfd7e36a023dae759f6eeb833e3385757d310587c4d
zbb6678383763b073252a4b7fd0441aa787a60481958d2d6738e743c21f834a5f324837ce6b2ccb
z9486f283552156ec67a8d7e1faa77707dac0d18650ee2591bfe1e09204226aeb6a2a40000fa608
za21f6e8117ea160fc38906b2a73a4bec48e663ad3b76bdc8c8a45d64bf7d54b12964295efd6f4d
z689b89a5b9d322cf21e87519dbb98b04a12174dfe5ca4273584f90340497580d7303a87511c0f4
z91b3e412010a02ff550f5d1d8cd0901dc8df1bdd216e3e4afe3e736ad295dbb592457cfcc6c8f9
z16583d503499121758fb47bde0527308d26971fe9231a8752cd6b3c35d4b37f2ccfb92e1b9dd8c
z76a676fe53aef9b2c066fc768c8a0dbf19b8a61c52f953a49c88ad15fe945111fa42bbcabbf938
z2503d88321ce838ac6b677fd27e9cdc117ae8c31a850b047f6fc7dd39ab8d6eddc8a19a9d1c5d6
z5d07eaafe561bbf1ebe08edc3d2253348f571e22e0b2287b187b43d5e87a8c5f1a3548a282f795
z5711ea391f436bb32934a3c8e51617ad9cbc7ecc1daaa0e51cfcb57a4410161bf3e516b0a2831d
z80339c5981d8b12bf42efa28c849dd235d0d02068d5a9d4dcaa5d8365c513e9cd5c4c955d7d9cd
ze3cea8acc5208a975e0a202e0a5d3c1a580fcdb93f105577a3c0eaf51c40509d91161b9cf7699e
ze124d0ce1ffaa6a23fe8c97c437e729708c1f1d8bb62b54130d788337d2be42227d4f10c52a208
zcdf3198b40efd788a9068ae84d1e4bf45594576d03829c1b54953aa227a784462a698dd4415c1b
z2de39d3a761344ac8b00412c113b24a5f0911113a72763f69ed1b5ab4748bf46f986dd4b246f0a
zf9f0444b6cd68a1406d9df046ec29e684017a57e383bafa4d74993d1d23807249bf4a766612eb3
zea78578a12fcbcf7b4f138bd40faaac8ac886fb8e7b92f35406438356a232a14c263f143855699
z6f134574831ddb518f89cad2c78c448ee84fe987046d916ed019aa1d5e51ee18090c2d7e3be29e
z0cfc2e32a3d4464aa28d2cba3f0ff4b88b36393d359ae18810f304deff287915aec3f84f818c24
zce7387e991b6ed1b2e8d7bc368cf9046caf3ddb91ccbee731c5345faa75acc23afa6ac18fb2881
z5babc2281e892b17dc1f640ca99739f659d6d45540dfc05ff00654aaf45a01d3ceaae777b783cb
z90b14d0fe0b65e624e6ba187d9f9204c7179d3a2a18121b8206d176f376b6fed5597cdab918ad9
z5c069ad080c62cca7ecde33c5a6850ab6f6281383ab3e6d084a2976ca22415fd1a206e5ac04367
z9dca7bb50f8255a5623df69da96a0b8267e6cd706a16010dfb73449e7a4e342124dff8f7f29041
zda2142bf0b3f70bea9795387c3b41e8ea6a61e144f8353956d06e2dd8057f06d37e75f9d12b5a0
z5336326f04ddc9bf6406916f771e3e5718e7bab08555a2f0a4f98993254d44eae7a14acb72fa97
zee5baf9035fe5d5d40d8910ff1cd4453301285a58e4e3cd848f794a8b5d060a1379c1eddce612f
z18a6fbe8f413c497f1f1ca0694d362880b1a746a96ca6fb88162b4db8b2ec23892db3994c538b0
zcd4bbedef569edb79e28568fb96cd9d500dabc2ff30893ed88072d734f0550a770543c10d81f60
zcbf6fcf2960606f2c86104f24533fdded736dfd02f3e5781add498604f98333bab791fdecf8765
zab9c9c4f248de313109117acf6fabcc4b803b99ff782f8a7fc7919f5e494d854bf00056f57cc40
z2543ad9adf3b5f6ef5caf0a16e3d64bef5cce8d5acb26b9a54023e2eabfa08c8a229b972bcbd02
z81d02e7c04fa53596531a66f4bfcf0919f5951f38047d336d5900de7792d5c0ab9399d180e993c
ze89f5ed6e3a36f39b223f6c740ceba3fdba4311aa47484687a9cd40907c342d86dab40c12dfbe4
zf33db4b84c13818dad01022f45d8b12de28ff40242e105c709be37885c8ec3cfc9f5d8ac352068
z97cac914515fe1ad935ae1bd92c19df1d2a3bf1ebbd099ba3bfa62d6659d249a872e0d30b08b22
zcd3723af3a80078c2521549b6590fd974f6dee9e125eef17330804b2cdfa79e5c9a20eceee4bc4
z9c0c35bb8a42b15758b3c373790a23e7fabd039a32940f880841eafccab328df0707bfc0596467
z9ca42dd7dde87e74142288c357b66a3c6060e68ace2f293c0edbd5f4d15a686fd24d4d6a9f931f
z446e7d03490a41c5f7c43f5e83251e05238511161f070a947885d4647e8a20ed9227343bce3c4e
zdfbc5ca84da589743abe84607c918db1f2dcf8865411eebc51fc3a59a943005ccdce12f6b684d9
z7e3f67b1e4eebd8729d24ddc095fb7119a20a6271efc819a7b75e3c21238cc4090917f12edb5cb
z7249bc68785aaa103b4fc66fee0e8467607b8a646fdf35cdfb27ab164a399714636bc521470f65
z25746226aba2334d84ef0710f0df562033ba2a660079ad73e153b5c751cfac7d589e44b7c96bc9
z2911418bb50666f54655b385424ddb9c804683de9bf8c3e5c006a141ef211f437b154e07f3e674
z21c10c5b7dbc20c4c910c66a2f37c9ebce077b7f91fe887ec8eef8b9c6b623e74523c5c3bdb686
z5bb5f0a464af33eb58cafae928835d9c967b3c622ac723cb61a2a4623899decf84a278271e7db2
zf0b45593a1c32b7933e87ab5e7030415bcb0bc3520958176a9fe9ffe68a3016f9d27babc392c63
z8e325f85147471c7dd0279986419f1a7aa1f23794ed6fc750247e9d16411df18a3f5ed30978045
z8c8e5549857bdb148c53617b6bc76aefd49e3d17be008e23523bf14132ca622bd0f856625f2aa8
z4b5526879d1bffb2c2df25644eb48c90aaabd978394b256f43096ab21075e38d68de913f168448
zf4b069513bbda6aa8acff59a257d80b922cbcdf9b41cb993ff31cb3c8ef80b9f252781da7fc4bf
z677b2852e46583f8f3c37fd10fe42137db0aa7606c250af8dd8ecb7246a6ea14211e5a5244d51f
z27b67defa151e7b86f64e2cb7137e2e88d04ba5ba414940987e8e705bc9cbbdfbb2664ddcf44bd
z61ecaa62a29f9b757a1dd7c823e3ce607306d8f6793890e591aec31888636aabe78db8a64179b1
zaa9ee2843fd0f534dc48e8fe5ff7c0a8ab9a072ff7b060bc844f2e8c968a7b1448b70a55a214b3
zf5cd358d290799d615ad5d21d9bf218004afd4ca294a6cc0146cd7cdefb333d1a5960d7dad3d5d
zc0a86ae4212b6deebf6bbad681f8c1956a91b87bba9a3d88ea348592303d8013ae1b5e54eb2a14
z1bc8ea65e7a41d008e02cdd0702857e9da7f22a5fec5ba6ca41a7879be4518bd947ce02cc222f7
zc269437ba5d22e3989ef1272650aa228cb50e005417b91e24f09cd0b3036326379181a08e98b78
z11e122d41f4afbc137d3f48538cc43c75f1d03f27470d63c5ea758c219298e2826b9864fb757be
z6a20c0fd63ea8f32b165c10daffed8e85fbfa38147a9606c93c6c4e8fb2d18e738b237ac5dec31
z9d8b1730ef9bf68d8f1802efab98674e8691ff20d458d0460e48d5400591afea4c8150106d7041
z885a22406c8d5c5784c027fcea20352b8fbf38ed0dc0bd994fd5a62dce0afd74f8e6f8ee35b465
z85a59d587811285b668fd2dca0c7ac738de81f276eb7b8bd0f62468a036e6cdcf3b22300746328
z02097ce2a24d190981b39ef77db476684c537fd77eda5683d34bb174d270862e22d46ef358f49d
zdf2b1233ac4f4b41016f2aab01dfe8ae1ca841333f377d784b14213916e5523ed1eb7b7eab6f78
z3cecd20eaa0680597c2d02c914b007abae240309e84c30b7a720acffd7b548139e9a125ae6713e
zb21f8d4435d5a3d923cf4ef2126ad2fd7c7315ee818501a0f6fac47e105132ff3fc6e27c5746f3
zaed03378b18434242250ae68218ed87a561328ac440ca18bcbcae6e9985308bce7564b0d377003
z7f033369b4fb8fb044a653f6ebe318f42da6918aee7af79ae84e6c01a7850de1846eda65529d34
z5063873516975dc1cb352e316769ee6632698a3efb7e578aae360f258cba7fea8e2b0531a15634
zad94a64afe894c33157f072874e62cd4a2b1e78b7aa0293d4a0a2441264cb9ad13875295c40d92
z8d552d97bd733949a69395ca5fb09e475b6cee79461eb646037cbad2db46a53daf2d32fa684c75
z072d0adcc3ba053916dfdfeaa1586e5af06fb8759628e7738cf598507b8d278785ee281909ed83
z851a819d2adef4729aa48af1eac48a25b90bff5c198b4284f997bad51f4620273004f038479712
z6ed59e907c6a5c41692b24938b784f30e378e4616ea5e1c445d152ac61868c06f2381e420b26b1
z92bf4220102f851084611f440c1d2861714d0934fcff7157ce85834c51dfeaa8c0f63261b23bf8
z58b07e8b5ba3e41f3819d5600929aa943cf41cdeef0a20fc313f6a01fb5da5d1bfe9b56ca26e03
z6c46da30a586caefca6e99d7cdd59bcc945255d0ba33567e6d138da8fd8f0d5e0d10d66cf64688
zf868b45b91f0c6e279a2630cc44afaadfb39f533063dc4ca02458a1a9addd5ea4e22be206d775b
z179dd74e2e807df46807bdc96f7c0045fd56649c2c7490395d0b5a7892b0d89b9b1f3b666d8062
ze891456e73f22561ded59ee744943167ef97b7d7c87e0c8335fe093c6ac5d94ec5361a1377a5d7
zc086ccc740456aefcc2b6dd97aee3ace5bffbbda89f36d895a0c17e613c28c1033e0bf1b37d9b2
z8924407d9f803d8a5a40788ba2fd9e3a6a9a71bb48cc52143187cd779aec18967a03c5cc35302b
zdd22c6d136375d7a9cdd50e8861d0ba9f9e00360b7cd6dec3be3e9cf67852b55478503d03111ce
zc349170d27921c4afffbfb0c3e0bee3e49819a36a9cc3fd3c574facc202ffbaeeb91bfe9ebea49
z821168cd6eba384b210afb3a36a90f1f60ed051ca910f9c3c7ba4bc8aa2ed06551708952cbde54
zf56763a2902ca25962980d9c71f7c56eb7f01188cbe48979615cd4f3250448f7d9bd7a1a8d51a7
ze5a951d322fbecaf827fcc146b6a8a12c556dcb85653ba0ffd263f037e2dac495dcb9151f4c961
z65c1cf9cdaa0d9acc0393d697ba24a96c0131605a91f9a73964c6b4045f77c6c00a661a3076303
zb2cdc30d434ac83662bd4e1066ccac7672f6f8028be70432cc344a0cc92a51ef9aa07ebead12f4
za86a7d21ebc13ae551e782af6302809a2f7abaf8de740eb2c111063e836a2b8971da22d7b3df5e
zf87fe648f198b138e81b90220734fc4dafded30bada3f0ef37c55c486c64f28fe87e654a6e343d
z2eb481c692d74c948c6378378b4a4a0fcf174254b98e6727f1a2224f1cca7e71c2debaf5b2f1ee
z74e5acf12560e39ad3a76d1b7d79b6f2dbb733f0d8c962ebf33525c73bbdf5323259c0b43a85c4
z026d64d4033b10b20ddcdf4cfac89dbc5f708f5868c2e8dee42eabb24b934c2de534a02f9e7907
ze5f7f50fd0e890098970b3ff93a5cec23fc8a5b1e90e4d6584bfb2df1f9e9bf334ce53eca8cf90
zf4c014a5544935519016fcc9ffa3951cd3aad9961850f2c52fb59a61cf56bf599a1467968eeee4
zce92624cc0523d34b6cda6ced1aa78d2a1ff605c508b29db052b9240e87ab68814d21154932d99
z15b15de7a4419f6a04a30d5b2e4390e560e916e76cd50658cac1c094ec9cac18668465998c0721
ze1172213fce539021c503b41ce4ba1999d25bfa9243fd4bb7877f0fa1a89f0fd0289ac696c15b6
z307cb37ce23c1bbeb9d4fe8c7360f6808ca4a1fca84efdcb441b2dd70f6afaae14de62a29a6a2d
z481f61dee46d7c86ab1f175985795c337144f36604ef92c6f40075497807fe524377191d0efe22
zd9d91c3a6e943759a7b3f4501b6f72e5c972cab417e3d95d161ad65dc9bb548617797f6f180db4
z185942fc66f568c94a00eb7e3c760b44bc24924e7e9e2394ff6a3b886b400916af4eafaff6f972
z33b34d8b00ae2936720a31033c5fb879321e43a35b2c9128d233d2e9af1cba3363738112a81938
zc2e12d23eb100a271f8af4dbcca6f53b32b041a143ee665b8d61fedf1f477bcaf727c1635585a3
z1a5291d5e4ab48c519a832136e7f401eec6ee940425dbd00f9ec013ad3bef5e555cd6fb0456bd8
zef59692e726bbdf94d006e5102fcb541d3db533297ae9caad24ad69cd3d52e03e5c37eb1157cbf
zc441f435c4bd60de0b115c96feae0059bd076f089ed83c857d35efc651f9919d76966b16cb1517
z72fce4f4d4909b27168171d130de21edea18496ae7b19c91e4d78c902024c9e208308650742652
zfeda8dfc8b9dbfcc12ceded9fd1a87ca1c5a7de63e15fc0f9eb9dbb7f21ff9db60d3a1a9b30fbc
zeaa38f526c09eeb73a4aed509cc64a30de1da1b88a5a400d45bf5cd7799710b84cfa1782a1e7f8
z576a0e49082f56242184930512bdd4cb852a776df786c80e72d224b17423bdb26a58fac5fb3dad
z4b1d036826ad485108466ffd61df92ee711117229b9cd3a9f22d9cd579107739793a5ffd7c25f1
z00326d5328c615064b932b134f8b82dbdbb0a5ed665f85a852b7ba4fb360a226ca0d3d22cb7186
zd31541dd61385f2cd171648a7f2ea2a0ad69452328679acf98117df7af3051932f69eb33d654b0
z549687a2e77fedb9a7b6cdb6e731fd589779796731b09206c385e6744d3a59fbdd3383045faa6b
zf8aee624a3963812b34de061ac66619ad31321916c5b9d4d24bb5b6a24a60b46c62f8ff09f1dcc
zd205a9e7fd9073e0308b3483a8d28b432924438ea7c9385f2d70bfc3df6c286ff18af97900caf2
z193f9fb1252fdadb46dbe5a43da091d17650764251308cf8b2789413c01c704482f0d7301bcab4
z3b220cdcbc2e0670a262e7d5058a2f32d47f5b3d7c26f6380030af54b77dec6523d150ad516c03
z25713a383c6cacf444c458cdcfa506470cf899b514293cd44a8f0e28c7b8f4582a88bdbfce6cb5
z81790fb576b5f22d63a6f68be00636a605a1d4fc140b89e3b84a1da74c050f717764b283fe2fd4
z2852c26e42be67291815e2ed77bf733019955efc7543756a200abb59730c58b4828894e6155324
z65c4493a35c7766547652b4f0f54e971b927682fed470254249272a6b7c24efb4fe820115df1bc
z798101d580b5db684f7288d47c9a461577919e3773e786b96cc4ae0db9d4d815dd34ed4255f555
zb80dff81d763b390fc70c1fe1880237a397699c2d508a9d086bfb354421beb2e1755b1707d84a9
z00cc1139af7c94717511696ed581c01f717d60e70debbc74c329434ee21d27210a447580deb9ec
za438f91b98ac2ae910a755d3c7e58a57bbe6055e256510f93ac9a37f1c199d86e95d058b0a8fe2
z85baf9e45c972cb1709540b7f7bd407b2dc201f05529a5ded52bb5713bf49ee8c4273be200a4c3
zfe59e54911ebb3738c4c0b8f8d571e7e27c530a60f10b3c2bccaed37220e61a861f0ce1201e802
z6935621472ba56ab1d3aeb8fb83a7bf1cdf6aab2c8ce88a18e83bfbc8f0d105b2aac62760ef92d
z42e9d8906dc2fe806aed3147ff4a02bb799aae79c8388732cd56b7e1fd23073707ddd019d03120
zdd6a50d54f20154f4125ee40d328ce43ff0f6bf35a1001c0251f846f996c19f4a9f7b384522de0
zc9b958cb6d25fd31ca0ffabb7e2e6f84fdb9b6bfafb6b792593879bdbb58147115195daa73c738
zfddbbd8117cc2dd72548af93911ba352c3801c01515de710e1c3476663f3c25eff45b691072b39
zc35d610397096163181135c275726c5fb15d3c84ea39966778c616d24af9592bfe3b35287aee14
z2d1c9cc435569bbb5bb81cdf321bee878a83a836c4b911853c937be05d1828d06cda92829b6021
z702c3fa8c215193af760e7f25153c4e4c61994b58a808976823e8cdfb7f3a51e3daee3000f22a4
zfd410800221ff870dd987049a6b1cc4e7c791e9b4c02cfe74b448f466ba9086216fb17e9a0f2f9
z844b5d2f8d1e782e180dd5fd912ace8945766fc0188caafa2011db2f0a791fda0c84cb99aeaf07
z2dd940b4fb7cc962c98f92aa6a31dc24cd6a8df42be2c5a3cb84c8f658022960eb644b3c369d4c
z314ed66a85c46f17f412c67b92e2c6b745577957f5f7deb933cdafbe897779d4a688c8c805d4bd
zc8f6518fe27c66bd98c6f4177386f3c00edec671096ec7dc8825f69bb7710478db323628d629c6
zdb16cbb4ec42c1f60fac84dbfa52fb287ad6156953cb580b3773cb323e9c355262e23f86d1fe24
zd41a72406fc427832007ecfaada8c2b8c97ee8f8b925c2de4cbf62ea2fc0801d49c841c63a0e72
ze93550337abd50546ec741773d8a2e8ce832bb66def92ddc8a24b9dcbcbaeb65a047a43a682f78
z00f2a287b112eb09279a675e9be421b7db5dff8dc84690abb4a74601f7edb50b9453478f8c2e45
z9b457389d1564974ee849c32c7d77d970a75843c64736c6ef5cfd7f6577cba0172217c35cd976b
z128b9eb83aef645c695846ca63794a773a3de197f2973287902db04c9f2e884a8606c7d95aad23
z104366ff1f1632cef139847db969ce24d155701993f47721b6e2d7dfb31f23d52ec517f76a6814
z1fd47de81021735bcf2a2ba92b0ceabc99fa99151e1e197e1764628c73ff99426e2a53460a009a
z6bd5fdd1841825c5038f4323c14566d3ddb0e01cc2db25e41aa5d32006d2cd09e387648225566a
zab26d4835c2f29e3f01e779fd1cd4c5c4f6ab396e2b15a9608043630a6ffea46439439b07cab36
z66b5adc4650f39801566debf13fc66628b76bcd35757b6752fff6ec8b2f9e0698f50808597e395
z32b53cc50625afa734415ffa47d6c3c1fa8cfdad76c8b1f025322086c71bf5ded9cbf7040fe345
z98296b254412515827aa3231e2a4cb308870db39555b030db8c203e3b231749c33d0672225f9bc
z610df1f0b8ff484dcf08f8667924d0bb65b954f521607a2e39991e6dc9676aa4897f837351a652
z2a9f0cb113294a1bfd558a9a61755dd73f8edb021cf06bf26418fb368e10361f4c67f2706fb526
z6979f6770f5f74ca802a3b94c6aaf926844ef853a0adb4752c9a8a8bbe2817dd09a5d96a6d7546
z7e6205e421c0575139de14d41397d530f8bfb4f5440423a2334cea072a048f4bb900047789caa4
z1e2535ac5d343a4a1721cb1fcf67de09e20a5b77076bb05d597127380dc6dd2e0d92fb0cf9e035
zafe6af007a69b8e7e3232740dcccee1f63af2c3fb6f6103682225fc6c0405d7173aa8debe5e597
zc11eda7354bf7b28b0b929d43dc86205e8bf79dd907a0e1538f37cb4f983815f02454a89e5a071
z7515031d0e0896e8532957e4568135e1f3c54aca91d91e17b95007dba1439c0cbeefd4e8b08e53
z9659fbc2f132275e11906c7c579ae3b5f70727c51b2270f0be0cad8e7ba477295a6c4be8ca41bc
za94e96a989dc2145009e8b9a50e3809550165ba12f22c5a20bb24ea5d6c81b2999bb1bd9eb57cb
z86fbeca85d678ab30f22dca0274e4aee713ea42fc2ccc30a233495cde6512efbbfbf3a99d63fa7
z410c953b67e12aa8e143b02e3889b0a03ed85d956e069613ee21743d3d6e898f16f4b52ad0955c
zf9402025a35751e3979962832054ae0ba491d6c538da4c7430eecfb87d6964c0cb844b044ea58a
z89bd927ba8104dea61a61b15b7396a93d6b84fa90b8056bfc0e5f65b2d30d53dbc83f6eb284d42
za9e62676410a1588599c738863b3f85aaca5241add4e8040f00aea5488db7d3f86fb1ea496da60
zbdc52a9f85fb79cc91eee411a6acf3c9f7d2ad910f06fdd32afeeac6770d93a9ae7cd39bf04ea1
z16b11f2c03af64a8c80f9b75dfa9cb58c58abc20793f6d6fdb74f6f0c277ccbb8375d1f24ba46b
z05f1a5b6c703d46ba8510a8e2e0221d7075f98dbd0138367e809964f40f8ff8475dceae0bf89e4
z91980c187e20ac336b05fea639d36f044ad25346f2812776c760d71970501c34890383276ffdcc
za2c7c4cb294aa01a941f082910580cb520d9c9ecb4c0aae9f71e430054f41cddc9a63abe51ec39
zb859b9f9da2768297de89e138d193b5a426d0ef64de4971ffbae5d5b7f33cc179e1cfac45c74b2
zda3926d0b4bdff97d7ad16bda9001b112bb1ac966b80823c69415b605170e287f56ba9760ab635
z540e8600802f8e7e77f74fa8ae143a060b020060e10381bc135b93950abb880f96bea51951c685
z3471bf5a35a3ace590751a79acfc71b0d53f32cdf9efda49494adc7302e0eb083e77f96781d492
zcd094813bd1f5580ad2af1dab3705fb36cc8569e22ea9ac6a98cd0f931ad72d4c2b1383145e6e2
zac131693ab0f60794c8e82360bbe5ea57bece2b25d677fadba2d7764b2c5c15f2d9e715f349a9f
zd12deae359aa72dd94ee27034d5e35ba16a850cedfe99e084e11e418c4fe80a5a6f6bc07af2317
z3e805bd16f14c0669bf3c4448b35e23d800c33a4c87d8433cde0c01f8b281ec35a0016484b5404
z39535f38070983b6075a5d247bf0420a2ee85e1e01b181d047ff7e8c7d51008e855319eb2b23d5
zb074aeb10fb30641455da290e7642d86e6e6fd159d3d4e2e9f74809ae1a76d664f65c583cbadb4
z988665937d33530bcd5c0d2eb10aa265d852ed42ee196e6983c6bdbcd8a3d13b34a75fd10bb566
z7badf3cce705f8fd7bc6b1631d2bf0db2945b4ea36bbd1f765b2809427443177887c45b195cf5e
z274e10149793fa587fa1809ae23361c92feb791b07834738fbebbd65ed3f5a83bca2e6b3a1841a
zc70428cbb2be6518bcd42c7b2ba16285d228df9929a8f740864e3a7913659599519397c4be7003
z3223b85ee02eefb30180ffed1036345b1ad159bea7a38f591e29c4b567635b935bf7bb36642517
z04caa0f4a3a6bc7c65d3c2937a3a7a4e990a5bd15da89f5405c6ed86d7dfe2b3a32db462189c5e
zd514130ad33e9aaf372789e842bc9704b5af6d8622ac3575bed51e2af6c7e0e939327586bbf91c
z894290784c700da3ba969588a94c6a4e3f0ccc25376f22c439aca57d13942e191d9fd7c933421a
z7e30ed530157e6c0fb3755201ece35eea7d7364bdbd2672181c9b753b178902a63d3ac399efa6e
z4098d8d2e72f3acef05f373a4518c80c634e11b3ad8a9940ccc13d695b89a7717e52c8c0917948
z8b7bb9a05e001ef8c7a0cc7840a40fc52c5bbed2cac79666b592bf14366c2c97cc251b5f63ee98
z104958c7d4c9e3777d5b6e90d444bb3202dce9bee87af7ce13be28a87b86ea76f7fae05dfb28d7
z7a3366e9bd465de7f09594f06845ba6274daa669d121dbc4e7e68b6913bc24a624d5974ccb23f5
z31adecce34cedbde5189bb0e9c10559093e60703daa504451155581de4da105bcc55dbc2cb0875
z85dbfa7d41b110b00d553dc71cd4f355b7dcb222fb57eb0a4fb49aec1cd0ff1b71ca72ce3fff06
zeb53ff4441757ffb41fed2662de4e81e0d5597c1bca2c12a23fcde8a9a75e7b1af822ff0ea0d8b
zbefc4ef5626ad3390e2f0396afe2a095e2aea0a3b4c5d6db6414d207afc2976ad926fca1de4f6a
zca5339d3c76ca58e6c174fcb56a3860fb40e0d30513c10a82ea20dc2521fa6ad130a4d05da1c06
z3417c945ae68134c8cf3040116610bcff4eedeeb439a5d8aaebc5056a7709828823511ac693e18
z9530b43ab14bda4622e005cee2d94dba5f2bd261b1b49621f4954c1f43d04e413ac2eb1cc619da
z9db5ae25ce34adcc723a68367909e35d5c90b74e0d0b82ab71d1264db32fc8f1a06b7e1c1a976d
z2573f9f729e42b616e2ced94fd5f100d920f47246d0476d49852134598492125f224b248c8eee6
zf775908439ec64ae7af2560089078b46b2399846dc94952612ef396d5cf5a8864b6718bff1c565
z167726d4c6ca98161b6842cdf27f389a1dc2713754221fee6dc5d4a0c87566db8767a0b674ed34
z6fc6dfe846fff4fce2cdc1387cf17285442c1b5f5fd8265387d961910588ee2c6e1f8e62bb606e
z1ed2df15b0bda2017d5efdecc5295366239ae3a4096b7f29ed6a15c1d14ec5750aaf7055312e49
zc1392903f558536347dea727ff435eba515e1446039dad414812da2317280105a2143dc083e40c
zd6db1a286e1fe8b938d8f4e0d6fd596da6e36ccb09b905bc9c492e0ba7c2eaa789b72b6ec68578
zc1610cad88f322c06df4f0536cf62d8071004e6af8ce106135dcbcbe54050ff3bee65320858704
z6e864aab274aa6175f800351fff2a617acde329f266fba5ed57f4875f9f9a50b9262264a191783
z376185768623e00c86c36dd73af780cbd526dd091734cc5e6e0dca9384a6c3b0882fea106235bc
z6c53391dac206081ebe914f817604bb2c6bd43f2aa207452bd5ec7e95c9019c81cb1e884b57364
zb6e1227aa5e5f6113d7efb1bb02c0a8ff6e4dd680d25c22307035393b842bba01280ef4d43b2cd
zcbe3a398e3ab44d0d68482f1089713ce163afc82c75fbe37e3e23d2f6f47bed2bdb87c6b142541
z2bd7acc1f27bfeb3cbdaac64787800708da4f5d63e12f9b7d8c96c1d1b8ad78f833c05114fc587
z5eda560800cc4cd180c2e66108b96919a8bd7136f7d7d6d6f90d9f7320bd1af4d747b4810f2897
z091e97f4f7f75a7b48036583112afc0a561d9cf138c9af5cbebef1c5405cdce573af8137f9b193
za3943e2f0fe7c877cbe91955b1dec318f0942b4d72774b0dbe4ab45ee20804026167490973357e
zcf081420eb1d608139143d157da0906017665a7b8148453f25740163acc56ac66eb0a5a8dda7ae
z908066e7602c8b3a7a76589645dd66521c6b2b6736b47fe72509c4ab5df0ea3c8a024cbb87b4ea
zd84a376e0ef044b02c034c278c9fb2e9fa3b5f8785bb9a442985ac004c01b99c586c9ad27bc63e
zbd690d6ec2ce5f194e495e8fea19a4967d0875220a2f707332111812c13de826b11f2e678750ad
zb58bc8b5d80ec8d82a99b88972ac70ce7d3402aefdb57c033dfdc3f622fc0bf38d7156814b06c9
zb3dcc3a8afca8063541b30dfc95c4692d8eb93515bc6b063ca07a8136b7a99d29cc286ecb05f50
zd5ffbb15ac7b9e6ed951efb99610f2110b8a008d48c1317b18f0cbbdfa70f4fd552f5ccdd75126
z9e423bc40735bb2d06868f0326aa3d0a780a6e901d9aa8ea84f1b9999e3274063575656eab21a0
zf378cb18047611a4dff710845e4eceaaf9ab3c1629b88663a859f9031385a6038148502e7f6542
z6f12cd1f6e4abfa4769f8c001370a86e43747dfb88d195d1fd62ea0472978a4984abb8ebc718b2
z6e14833d166a1abb1cdb42e84d1d51858f275eceaa1a1591fe4118c8a4ce37613b2cc7a80aec52
z7f7fc81930a003ad3299535c3229067511738270a9f33f49586b7fa5ccadef715746f43d369eb5
ze37f878eecc95fe5139f5de304ce1feb822bbed7478d50d8d9ab58b10736eda83fbc2d08adba1d
z997c4329d7c759ecd594efa7f3471ebd2c6cd8f8881e30bad4876af72a3daf518706c4d15f2a60
z92a120b4276e9711f76e3562ad965ede10b7e03ae7495e8fe7529a30f788855bba292e63920a2a
zd7ec9ae0b447882bd033eac3c6f3229e22217fff590a7c053c51afbcda9c43ee5758c56cc208d8
z26918c5c52a7a02afa0a249e23a5d4d5bc2a09fc873cf711028993a4c2864be6486b1db60db427
zc97a415982a403fdc4642fff9c6a8fd7914cf85e7aee213ccd0f603b33b5a52ef053947971867e
z641203c2334966f7b0dd51efbbb8ac8cce4c4a9e3c91afad6786e5a0c2e6678d0b86954d9fe35e
z78d312ad7a21b0311018c03940912ff6d33ed9a5b4ea8102698dc89476cf8e0e43faab19f3eaf0
ze513bed773cead993e824ed5e5decaedf4d617e31b01e8a21e28b533c2c0ea49fd30aa6bc89856
z7fd59fd643ae6ffc4e2caad4d172f4038ca68b3f921b5f2af4b1adb2499faf589286bbca95c556
zdb5bffc5e00000c96c607b9af4a090db43adcac77289b4c6385caf6afc6480345748fa7758dc88
z73bbef99a4b37cbd91d1fe92d9794ec8fed7193b03f1dcf1e1eedef66c24c43ef137b9e759afe9
z321a7e582e5033779c9a9df6a8505965afe9e587ccf36a99eb845aa1270f62b076cc0b1c4621ee
z7bca76fdf3223e1d74cfe48155f0489823b1b2b7af9ce9119297ed329f526fdf7cd217d54186c7
z882d20a7d4ae0cda76ffc88e25150c29442370c0a11e50640fb9b513eaf23c3e851e03f6bc8825
z6ba0990bcea3d2cb3f2c84b6da356f5b142a77418840f8bdb378d653fe3a38e03783bb03fc49b9
zea7252d6e73e157a834f7317f94606a2233d90d8afa51217b082bfd9c9019ded20ab550abe28b3
z41c2a52e5fa9cdca3b4615f5be645b44c5bfd4f88e603718e62d99898106ceb1b7d634071def57
zc493bf4b6dd62a26a0ac62ca6c8879c4442ada730c3f82e9940c659b9e3e060bd73705b9e7f628
z1141b76839c91f1b70444b456e83af13e563e166793b6d89ad289507a54df9c1f9396c86e26106
zc571ce7f342d7d61ed046b7768f717c60d452463a2029a6947e86a58701798c16c060b91b04a0a
zb8ec9fd51f6a3def678703c87b38ed9bdd357974415f0625be8f771a9e10465dd8a217c5abfe4a
zf112065fc0f23ba067604ef2d9c3fb9dcc87d2d5ff938c29d27a748b711fe23eb8940631b8a17f
z6888d3014994a8a4c1d8ec589810f99412bc28418eaeb4ee36f62b6ab8f9c7d55c8a9951964172
zbbb92550a935a830e1c544321dede1b05e8b0cd17b8b4b820fdf7c903bf051c2a89c25a8dbfcf6
zb652beb5d98ecf3fceae09665e410718d4b5d421d359f7f7e2749b9230d7de45d7c67f487d9867
zee80b41c6933c6c8638da0feb28610c7d890287c54ea8ab0376bf94075341e1e76272620b26b91
z2cdf27c92dc5e5f9f62cbe7b05f156f3824b87eeae5f271fbfb8af02378d60c3182c044a92df03
zfd4523ba2a4508a37026a2041b76234f3b0efd97d0f5575632706e0ac5e7f8d9ffe6b7e0196499
zba246ae92f527e811ebd540575b55996ffb137af5bcc08dff5f9eee6be74945bc905b3c561abe8
z86971be257d06f9c2e10c371dac337a141d110b3b1a571c14b70df84c31ef28685febb39c2aae4
z6a645f3f0e23e916153014bc3d81ed259c0b0e6d8c3c94859cc555ae5b1466f1f52185979ad44a
zb097eed089af017ba398a1de34837d5e52786c59c669df7c0cdeb3e67f5d40e8f42df0b376fcf6
z3f4b6bab8cc0a5a826acc2401904ea9814e33c94aed5664979de390d09917c3492903229541512
za6e065bdc7dcd68b2cdb9b4aa684c7daa6a45407b4a54c76400066963f2fd678f1e6e431c8eaa2
z06dc5a41ef898fb317084e61e7847e0bee7ba1eafb3e738006ed206282e658673337630f1be938
z2c7ce049154a2d0136466fa6e2eaebdf7b866813295127613206daae0fac30a3ec197f4983120d
z7461f99142582da4dca9b1599e13982e439f810fc9f8d05fb03e8bc4ee18c070048ee28dbb7731
z48575ec1634b1d670647a63882ab956c0f0d0f75282914c4fc8923d4ba36e7dfc27161ac2eb805
zd788fee3868574678fa0200f79b51250c2e358b6f3fa0d96791f8e312ad074a9420cc63860b531
z24f64ebd87e3f39b541debe9f1aadc940b7f4f5ce1e4ef8ba7775d62f1b331e4508553fed62ac8
zb28b2f93ea99ee44a2809f5311dd2b16028bbc06ff5666601995abe6562dfa10a97ced50a19e11
za766123d6150ce2cc70600ef38c62422a3ab64a8ce33cb61d75fe61a0c2f29dc4f00c4f1ac4a3e
z04749a57af7c7355e27173243b60f77d2d31448809b99c007fe7ce0c4a57c5246df5692f5176a0
z681269cd83c43c55a8b29d3f646de364a0c73073cc8c533115ec550cad57a0f668a9a9660e145f
zd3359458d1e7c876306bc2e1de248c5938562e6c4f1afea38c9db740d2e3151a3eb4f65521d689
z58d6c3a2f7a383e6a5d97efe1a05b5de7014c1485084f4dc5610a9cbf68099adeb08fbf2e82c70
zcf1c122f1480f3eaf200eb50f2302e11f8534dfc999562fe4587b64d15fedf7f8ccf204df7e2f0
z846d35b61295b0b25531ccfd2c9efd127b670b2c0374c19c4473165f44cb5b673b12dc0d6042b1
z628d569235349f37495fcb5418544e7fa0eab26a652de1a93880bbd290f48b64d7ed560ccdde45
zfd6374d7bac3fb890bb1287ce7b6cb05a8d0b295016206beb3c8f6da32665c06669046e48ef47a
z354dda97589fc4a0af9fe1a6d1301579647f37b64d2cf0c5800822c95a561e2f4afce4cba5ceed
zff5305ada83a636f72b9372e92d4793f2a447205027e6ae0943159184866e74f9f84d5d8b0d6e3
z6923b3b5f7a8576d6c354ec8a84a15677484f580804b6a8930426f2b6fdeb128e95b64a7790da7
z90548eb4a2216c414e4c9e29501851a7e44228faba731ddfc11fddd4a4bf836e0f3bffe1f16d4f
zd1d10cb7291b1106086942207b1bd4208e9024a7263bf237c13cd13298f03122b4a28d39dcc1b4
zbb639085fd04eb2b3fef12c1a80a93691ed841e8b4449a2f9503b433a3499a6f4ee3b2ff3012d9
zddf3ed2ec25f5017627eb48c7a7bdee859fe460a7b8878a6157152283b5ce8aeebcb6cae70d930
zbe29cd7308574d4fca639c900f20d86a30246ebbd86cf89ce5a927015c53b229f7182df5037041
zf6af98e8058f4074665f39f1efe03f210986b823e812ea46e9ac358642b02afd3ba5ea823ea09b
zde761a2e387e4bcdf77dfa1f7c9308dafcb83003677e47776ae50a962c52f01056b964e6c61df7
z2fe8a9a64348d992b8ed6c3fbaa36e0a8169e2a277030a05e928a21e995352bb4c5e920e6a5715
z9ed8f25f7e26d955cb28445b3d3112d8f59d71483970b9f1ae48341cfd80c820d727f72717df92
zbc790f0b1e82c87e0fc97b355f402470a7ef7ae2c456feab318f6d1c04c823ff8321ae0c567dff
z9798c5d59add153e1cdfb73f1e8239cf670b2060c6354e9daa47a1f9a0383011814d42f4507692
z5676cace232d25fd67f70c328639a076a1ed5658a9811158ca2fe1dfb62f62d940b41fd5ded3fe
z132d79138171919d36ed2a9a1bd91de9c07902dd33b88ce5c6d0c23358c694a7935143a38d97b4
z405dd9a1325aedacc877e4548586bd77f5d343b1ee398a5f0b15eccaf447097821383d2d6b4ac5
z0adc60b3b8082fb39d2c3368ff9c8c8ac3d9d35aea6c557ab70f1dd6292b993ddf75d9767a9093
z029dc8f14213e65c52fbdebd9a767a951d3bbd4329958d0e23b54f509b2f6c7abc0475e1834893
z26e5b88a9646a7af157060c465343a4fa75b27a68f1465bed250c5ac7bf400249c0379a796cf6f
z9a6c304e5d487213f02e649f5be656cd140d298177b10076d61034bc9dc089208bdaf3fe74c95d
ze1d75ea675ac587c4a8d8e424ba28084c566ee7559b4d6e327d1665d7659eaad679cde878cbe5e
z1adc20b4602a5f76407f6fde0be9ab5661ded7dc77324b158158e291e162f623bc895f51401026
z09e8585815400e384337b560c0cf5df5697bfd0eae6b32467402b3c7bb89e7fee4b1c1552e0692
z6b60980e42f96c3c0ad493e91110a30f8829135bc40a90b9219f1adc0ccd7e178e828c37ff7dad
z75300330f2830f9f499b48e578585558798104077e45d2120ce3dbf12b53fcbfccb42abf0375fe
z030cb779719bb93eabb3387fbfdf4d3e95fbea77cc75599515e2d27dc69be2965ae60dd207e34c
zcee3d0208ea01bf08a14b88d6138c26e9a5151ad57a098c79af8f81556ac8af56f5db67fb14223
zc3f05d4575298589e943847a1e874f3925467c0414ac1e455f5864969d9b1fdb7053b6f63218b7
z9b2c53284257253982c81a79cbfdddc83d0f590c72d74ccf31a11c194ed37584359056673ce1a1
z4f21aed58bb0d52ffdd35dafbfcd946f0ba45231732a05c76129869aa3ef9c2e581679e08dec57
z92a6116649ac615247cd9fb1b2277cfaf8cc48227074f4356c21f8cbd5fd752f9576280c4d4cba
z5df052560e8b2f9ac0216a2fd91b48fbc7f2f20f714b3866d7f58fcdd906b8e4352ac8460a8af3
zb2206b042527a8f0e8162610bc1254c05d2e0cf02a54cfe9589026406d75c3870539deacc4aa98
z739e4dc1da5c2420f28b9b29620f3b6f474bbd5b747f3143857eb64dd0e9f5ff4ea32ac738acbb
z8e151d878c47ea718cba32c5091c9e8a5020d1e2257022ff943ca58eca0ffb6f02b8a576003cce
zbf7d09e99a99c8ec9f91461d59f976f1a2c3fc691527cd3fe7bacc8fdc9ac10814b2dd4a11de43
za47e6589b797bd39ec7de33b82ab45a843790412b5fbdf07c5af984f4db787b47229faf2d12c2f
z88ea40326e78a5457897849705272b93a8ea834b87302f5f363f5279f00137e4ad23a2c88c3598
z8ba46ae23441c335e2cb58c9b89c98b79035a4680bee929c52c081df915d79859166ea0e6548cd
z09df559330dc08e41b0f3a9a215ffd5338ee29de2425c31c856a0e96db8a2a81bf2a6887d6d9a8
z183ba908589708e64d1621a789e62fd9b3c970620fa1fe6e78c143b5949bd1555fd7ce4e8dad3d
ze067f15c673a0821ee7ff17fcd209c49f14a7a16a3acac9c7f14990b2034bbaebc4655d60536cd
zd2679fe6ed630d35c12207411a33d2d723d8392225fa15b638cd66c8a2537b0edf13a17dca3316
zd4451ff2136d77339a81ab6b9a3e2e490cd6fca403c32a1bc2f5ebcd4ecdf324e6c265663ce575
z3fc7d2bf05f43f953e889446894c31f3d3b7014fec4d4a73eb6cd5bd2162f04b42dde6370f7d94
z069ff1b3753d6fb8b11010a9f911d0a8bf7e1efc1e4cbfded00004e51f89064fd9bd93bb5e70c5
z632a5b36f911511015ec4423d9bdac2ac46978af980ec1cb7578ec18d301c18fffff5114043a60
ze281a9801566e3d4bc0b6a38f979e2fb8c8c3dce5a842da766af7822d9d90942ab40109cb259ac
z5ee93b663d1b288c51c391f85e253cf56f1896f5e6cc7b8eee030eccd22447696cd7ad404e4ebc
zf03ec9666bd51fc81f1d1504edf5697ff800891e49ca03e27df78a3bc6977f5fc67343ae0c8f69
z9152fd4933f7e342ad99802a6e4d9423b819abbf27adf81f537f4becf118fd342f969651d1afc3
zc9df0330b37ba2747aeb91136d96504125c1c307b0745849ae3a24f9047662b1daecd67c86a9c1
z1aaf537fa3198657c9e8e51e1b5bd4f8269948b94ea0ac3d6a5f296a14d25372bdac8fd712523f
z388abbf92652a98c0bd1046e5147b35a756e70a135f1de61e385db2d30e3362a34bc8d2c479a6f
z00b0045113984c4f121edb4e60e1ef4dee528ff9ae5330395d43d78da88352c09734243c0cb5aa
zd7a33cc1826bfda18935d2163d1c7517fb5f2683f35db73da80f2938d6c269c262dcf32bb9a7b7
z2987f9d93df84551dd486e60aaa5fd0d53e2d4fa4c4d978054a41683c380d0d61c3e2ab79938fe
z44809a53f85ec0231a057f5e2920d381a89d72488116c93e01e3df69efe2dd8523ee703c95cf8c
z6d3a7426c7daee16d6df0bf9ef749eff4896a7db6c7f4693e1969c5924cfd5c8533899f47f4852
z791966cbfecc4aea7501522199f7d606acb55a69264834d953f731b0989dae554ea221a26dfd89
zfc1a47007111cd66e1c3fc1c5ce97ddea491c88687903605434ac20dc0eccace80a36a5b740bae
z58bfa89a1a839ef0969306ca4d5791a5ae7c9af8129237582ac85e8b0c8e889247a97b331bc158
z9cdc4ca1b52ef93ba908246ee93524f89359a886fe716b75d5d577175ddd87d3971d51c42c0d3b
zbf3ea46015a815b7f76ca17ec7fc157a762af5eced301a8fa9c80645973d4c1a4d53e6c0b6e703
zf0faa8e83fc51c5ce950b1baed13f5f98f0d3f7f5d86c0debb50b066ec9f63b82f65f526f8d921
zd8930b24d7850ecc55a00ab4bb7f2b1172c35b64e8d540f94809d3d2e287c5deafee4cd6e4e346
za7176786207112c25cfbdfd2d224b1dd298de6d29cbdd451d23f0c0cba9cf5b0a6842308cddae3
zf02c22cea48518d2e275b50dc0f93601120a61117818f262710416732d2d030bc9858537cf7cf6
zeed1cd3efcf1a7af3318e610b81c225341bb7c61c2a1531ce02254399af72e927dea8624f85bb9
za2d485572397f0f35c979f008a654a02fbf0c8cf2d73e2406836344994efd85d0a9d4aaec39666
z1057ef248c19d1d590a4fdbbafb79790234bf1f476564f10d199b8c3609aa4821ad1e5b34acb37
zad7492e2c90e6a483a6f43383ffb68c35c82c7c9c48b6f495f84b5637916d7510a7c1f2be608bd
z39c2cf925ba1d54e52d16ab50c3fb1819cb60917067139f2b1b9cfdef7610260917f2512a45f53
zf75c443e3a15f746317e30d6277480a75f446100544e42dd0dae3e754cfb5d3c98d1adf5587aea
z1e8aa8a8cbab37b551e73a4c544baca629a26f35c4d85bbd4f72c42c36423f13847f401ee0124a
zf7eb512aea117b08cee5f54c796a480b51359ad7bc2d49187b3316a540c9494c254eb96cdba32f
ze874461213c2d66e0641dba9dc2b1489a293638d52ec2cc2a8b7ad68d9fc797fe7acdf3b57c5d8
ze0871a086fe32c63c192b44d5cdc22106ccefc0943a408cdae0624cd4065760049e1d7e6331f48
z8771cc5e5da5f7b4d94dac74010d59977b84b75d4e17759524f81224248bebdfd972f80d8dd243
zca5802fec2e58b9761342942f73c3827ef26fb7bbf0fef67e3bb422a8b96cafc59e54b12bceae6
z964f29229345caa921690f7745be500275b42c45c71c249e59f07fdaeea3bc00dfb8f3d658ba35
z3169d3c0611e733b050295c3fb77522e26e70dbefab1a4ae51a8a9fbcfa44169909a903a1a0325
z729b4ff425d5772ff758614993cca7a9a807133c612a9b11b7d85990d4793c13a004d598ed2fc0
z7893f5c9ab2dc25a7941f89143cf019861763cfb554b6bf060e71fb4743888ad7e04d189634f12
z4db6401e965867e12dc8414b3841f966640921dd8316fad6b986b39c5a530290b402ad23e4d285
zf6fe43eb323e6db21595ccc3db79710fb9bceee6539b673213b494eb3c8dc378e3fe905a941853
z34d3dc81dcc8107bf5bbd90355e475449c010d598649dc5ccefbf65895bc133ae72fe6aa8d1158
z4c924a6194f74d8ea05e8a9246241d6082c007d44a9fbd64b43248c3c11c57a985332d17ad92a8
zd079da0295a0b66c354fefb61dd9767646c34daa92b89274098205618df53d619f8ee416de7074
z647c2031cfdfdea757829c53fe34e3e55ee87816d2b720cc33af752a3d7e9db1716d5ff13b9ce5
z97354d3505d9adf2ce1f461030c35d41564ea483f1e0e19f16e7e318b367532dc63535f98044fa
z48db31b88f74df01315be801e7c97f123070118b499dba27427113130213ba362cd0036716a5cc
zb656f824839aec4eeaa16ea35a77d56bec62f499f2616eb00a9bea383179516382654deaf6f112
zafc37848c697067d3663d25828384217ba21c195cb7b232cba369319c30f4e1d62c5de67c90ea8
zaa73c9a5849499d79980379392164ab00483062b71da40a1cfceef0b56cddb6b7f28b25a69c83a
z9aebe5fad250ab41c6da680674521e29985131704886839e956900b769bb6a3b38a546fc3b4307
zf94ea2bdf8de89147c922c6559dc55748f5ff25c683f4730255f402b41296361f9dc31d1245206
z1cc2e58d9fe90236e14ea4259d9cd24cf0ad636b36bedd90800618fba7efe50ecc23dc8cc657d6
zd597ee4dbecf6b5d7d552155fd20470df75c20773e56ef1fe4ebaa8d4a6ad509a5c4b3702a70bd
z2f38d832add347a9f1c5568bb2d4c6ca948cbb60d5e97d6466b6ef7ee356cd22dde500d9d53ba1
z3925e70caa3229dc035ed67ab61903fb8ba9441cd9e5c64e713fb44b668a15226b7a5dec5d4b77
zebc34e46f521bb853d8613501045f36d0a9e78409f85b15cffe295f575f853b9c35ba9e252fe29
z4e630d7d38ed697dbdc8eaecbb97f332a07f2e5267c89d39a4ff6bfd4e46827e2f144ea67abaed
zad3d7d707679fc8255062438d39aa52f70c48280811aa1e4cd90f58e2e9f325d42582c0d17c7ba
zd46fdf306a2811146cf933a025c6d6cb277a567a9eb4200973e014954c0da17da5b00da62a34a4
z7d338cec67c598256d6da08eefbbff3772f287ccc0e08be26493e2ee96d10cc4a7667ffec9bc76
z2f3b7fa5149a44c940338c57840e14868c45c393c8cc13909009334795a848d74b64642fc9f129
z63b2230f5905aebc276160cc5b7946431636ac7987e4bba11d1dae9edd935ae21651df9cef025c
z8fd8f389bb66ab7d71aefacad190d0777a8c5ee4f1965f153d679a30c9d28b1dd3e968c2fadc77
z3ab9b52c6969b6639288226f687d49a7a6be11e9118909592a8365befa2c96b2406999959290c8
z40439e755635290f55ae8a9e02c6af751dad2dc8bb5a1a5df6cdc909f9770456818620671fd39f
zf6d9d8c13b97b86b604027d4be01f67a2a15a9893bf76a56bdad5883f73a372869c131aa8d36cd
z07981da6da657616c239e896707f79a5e7cc08eaba219ae7df63e82f0a9c1a95c7dcf2d916d57f
z568ce2b019136ac20443c12e3bb9940279a70fb28cd4182c628239d53bef878bbc1adc88995964
z52d40a500a1f87cf3c7df6cd5c522c733a75da74bff924302f819e59ae27e6f5814ae648bf13c1
z3647918b2bc25707ca312a7c10eb717d9fed8d3282ed77cd24dee54e1de104b9c7f445d9b063c9
zc862b4dcd58636748fd5ce2104a48724c4fb6c620fce5ec3d5744c14c4ede70af8171796cb285c
ze4eddb97f597fcbd2f1ac53511f558311a3f519fab360396862cba0888bcf1767bdaac3ed70664
z9695387f9f300cde4038764daf4bb394791cc9d58069e0c47a0ba207fb70126e5f4543d0354fa3
zd4b6b268e6767221b5f10cad632ba3655d43d38e86f796e21a3f2dc35618b607c20063bfff1a4a
zb8749b7f91597697fb09349cd3eea54756410eaffd3ff0e376a43956505984c03a584e2ab10694
zbfd4d6f8b303b82bc7cc26ef8599fdd86444893689be1bf313722e5e647d9dc1fdff4e9373d7ce
z12ba9ebdd2de41b1319bb91299b4c1f9dd8e98f2d75f49339ba1022e4ea33ef9b7e6001e547597
z941eb2eff58300cf133b993e0e328dfd08725ec96fea0284a55c3b4aa41ed4e3bf799fb7c795b3
zd45261fa65f7d86bac3fd71e2bd7c8a6548ed5e04d32bb513d27948b7fea0d673839475b42b279
z4ccaca04d8e254fe9a445c6559f574c64836fadd98a2fd9c39556495fc38a0c1d3e9f91e10a081
ze7e2e247defa11ab08520f39a24b537ddef059e9f4dd93d22458d783282a194782beafe116ab3f
z54a43d39f6c9683ac3b5955799d7ffde0f916d3e11d5bfb713de581956b7cf834bd522a3a1e6b7
z015baff0bcd61e21b48ee5e305907247611b44cf66c7fc0218d051a6af11dbdcf1a8a1b8bea0b9
z19f5a30e0b741eba13db688235f23be5f05542beb606c1334fe89c0bba5bb2829592e42e7e8aa2
zfae32f9f46b04aa717a15568c2357b82ef2e16d40c9efc884d16a8edbaf5f3a3265682d72ad90b
z37892d4491f379ee992f1fb0ec52de93e8fca033b24294099928161c6d1c95155948ead9ea2cb7
z264298b1e6b7f1d3968e9f683b7f81f620b51c95564433965e409f2fd5d1474427b57d76b4f63d
zc39721e7ef52057f6a31cdb01991511fc302a758b2fe1dd5fc81c2760f026b5bdf7f565e805cd6
z99adc84d321ddca99917bfcf942e7e1f97b8cdda960844b74651d460df9e291d9da2ab0982ed8d
zc7c3ca536e023c8b8b6cd4a8749547d4883bc1ea03ccca55dccf2510fd8b17ac4abd04a813464f
za63fc9846f8336e56e1732f106d1e263c5a143a5576d3b0f244e89c523bb7baf9fdfb63e565704
zf832708dcf7885a7bafc95d20f0695efc7616c9ea64426ad34be0cf246a06962186be9e4bb1531
za3080b8c796c4e7154a1b830b41cd431dec5c29b3f3b322ceda315486fc866b2bde075a2c559e5
z7d0cb6d4da91a572d236dd1d6358e49d6e3dc4eae30e8032705ff71b46909e76d287b2ac7dd11b
z58c658a0cb10910848e96fb166f4c62f8a60c8a95a3cf2174d43c83db6ba5b0d2e49bb394a9fad
z8ecf658b9b7ad0e0744fe8d0e51d5400416d9ab854edac1ac98f57c5c8fe36247f90b023a97699
z6d7baf7c6b3ef62a3dc8d8a3bf3d6b33841dccd1e2218676b367f41bbb516c294d18579dfff9c2
zdcaeed99ec79c949327c94f320eb72132d3f9ec58877a8ec42f7fa57e6d6837e6aac78baa08da0
z049592c51fc9d3a5c5e0da3c178047e7db97ce9b0eee61182d6e6c057a1566b4ec1f7388c41822
z9aebc65d775473d892ed4dcde3c92fe8895cc8ee2d7e6c4e1db7bd3b3eff2a4d1d2029d39536e6
z6466aebdeb56b76f7513381360aab7c88e67487299400aef6c9b254d8d4827f730728a7aa1b7fb
zbb6461127828af01413d895c91b2f3b46825fb68be1b06afabf91d09c2847aee58beb35dacc9a4
z987f0693f51e7115bf18ccddb73a5a417c15bad77f0d5f680f02f3fa64d7e6f473dba4bf9a7967
z437391fd4009cf8326b71b69a5bad0a9ca21ef6f0297704b14c14e4b87dfae06cf1d2daa1bf6a7
z80ab8ee7b53de8134097c83f3f904d18185c877fff6383971c36b6bd9f3a107b2bc5ad7bd8f19d
za4e2b55bbade29b15a7891ecd465be7793f90d75352b0d1a3db92a9ce09fc40c9aeb0f4e8448d2
zcd170a43466325caf553d437fcf68ee5cd91e736d16b85457a7e26f5a67b3d9f7d0ce70df47802
z0d1feb403925e3edd80189e75bea5b0512a5b8bbb19e4b34ab356d70217dddd54226dcfeb12b84
z0cd2b99e8b2b715eb1a03a253c982a445bb081964b3c1dd16a28c3edd1bc2c9299589279cea68c
zdb66bbb9acdbc7e43d48b5374725ee374b2a57328fd48e934d1103f531256ec13984bf728e66e0
z150defbc2e4af386b84af7f1a78515e0a4d5833c811727e3484fcafbcec91e202a100a950c826c
z8e2761861d2eeac4599b295e3be549cbe8fa0eb3f8417cca002a76d9d81f5c517c508c30c1fe1c
zd91baca7c1fecfd0ae25a0c5d2792216be8105bb4df02782a57f0bef3317917a585150372f79cd
z53272d67363de57ef43eb345d6f13bca7bef6b52a280a10656e8be9846ff37de66a46d0700c650
zc74e2f766fc467baddc30b8afd2a1175507ac18983cf55f05b26c3e1d8615c1f4c045befe81f30
z905778cf57e6e70ec5417610b72ff5ace4bc0c5677eec0b95f3b0cdeb8b23178640e1bb3203ea7
z445477f596c4e0f3cae1e9b40bc94ccbed15b24b60849c44a427bb05c2e2ecc977030c278353e6
zefab6c5c6c2f27f01f78702ce3653a1fd0be4a9318118ce73bab9ea80a4a583e8daaff6e17b301
zb0053103d68666c5282f0d1cd477b032969dc651272ab301aaee8b2077ddffb8e863fb6d60ef1b
z856b5984703bce64db5f5ae2dafbf03b67b6c6f300bb8fa1077dbe7a24501fd257bc4b8042a75b
zf54f6b5db201d5e0fd4678fc138c4aaea5d84f43d97bff212aa4e9469321883afcc1b194ada547
z9fcc69fc87b8a9f21c6a9774ff182a3f0487d3701c4c7a1038703cf5d4c6d3dbcbcabf39b4016b
z1244e347b22bb1c645ef55f9607ae2c81c4591947f1f53b3c5051977482a389d8dcabffa801d01
z22c3122df2f649423c5c4f23eefb1be23d13e0e54d35c97adf13bac0138a2ce1f9502481c4ce46
z8fee80c3733f87365aa6ebcf8822dd87338ce1d77abb3adcf6bd74d078a8d5a3c9771b2ade9605
z09e40f5106754e1dfab851b059c9706fff3679d541e1496599f4c48d7071089541b2dabc275f4e
zb799fd6f3f9dbf5faefc4718bcf47eda49a76e2aa7c1c52befc4179aff6a9898e8593feee362da
z39aeea6e38e86805a8cd636bb25e534961acb248b9c4662bc7b60674e13d2bec0f9dd5d8dde052
z809b87d7bd94f32b00f4334588c70165484c66bacfdc1245506073694c690c78bb55fea88b9cc5
za9b29820f3982d3c295e9b7e1a0c0301441003ef2ded7083f6bfc66a6915e5bea575c109ba49e4
z239fdfd1aabcd5b39e5a258aa39a7770df3b246e9a4c87738ecc112166010c7d42bc760b3c1f39
zdca6c2a5cb423d47167911b123f6c74bd45789d5d73f4bbb64fa1d1e973aa4e275316606bde03e
z328ee345b9d42488e993c4e8354d5aa1fa66e309304e56432c3340de9d5f2ca2e7282eca7a2f70
z996c5f5673a3a21cf5ab04389a7ed0040be0e230e12f04db8d5020962c098c68810140b2c57284
z4b36111d52fd04f72343bec24b0ecf79a3f0808fd7af60191e4758bc8296ce77cef33a47ec4e2a
zdab40e3d542f604b0d94cf61a48c19495c4f183a9730d2756c6dde1d928d74dab32d8dc9d9de02
z9e0bc0145ff2e528b65aa9957fc6930e99a11a6f2b397cf4379cb24a563e7df94a4957b1c3a2e0
za87a59a7fc04f541ae418ba445bec3ef55d464dd75c1319a8fb7fa76ef24093e4c187001a34b6a
zc908c544c7f22ef6c03dbe0a1e4742e76dd64458efb81ff5cb8a81e24ee6cf728b6df62f48c908
zb9aff93a3938e938c6b07466bcfff482f6bd30fb65fe9b9b9ada87760e87cd0f71c19b9232ea29
za9312dfaa367e08407e877201f5f2ba00c2f434557201e6e3c10b76b84c86edee0eaa64933b389
z166f36a9eee258146c03ec74cf962db27d1cc7a78d0b472c4cb47f6c5d965c1c2225c883ed5d64
z418c401e9b332b53dfa052a9be812eb6de863c1eabf3198bc2801cb12154c435a22f84b91ffb05
zf7e4888de4bbdcc0cdd49a10b01dbf8e391f49b3f3ec09d555fbff4841722aa13d965afa83a818
z240712909068427e23cbdfd8071cb926da9f3545dd3e138313c9088b13d1f61a480a147dd5158c
zaa95436869163e428830244e675f74fed8cb54a75ad21c39efff841b16e5b99a3939d5f1262694
z0849ef1b4bec1c799d137247b2c1b893f2a5b5768de48cc05bdfd41d7d5810f48a91d6e7eee395
z94fbbcc0c3d7abc62f7605045e5176c7c99dc9b1ff09b9dc9a3ff7dc55f2a8fdfcfeaac56caa6c
z1b5933c7bc0a3772786c89172e715bdacef00ffc35fdabf883507f228f96bb516f82b5cb474ac8
zc93f3b14fb6ea9f71513ce1d7c3a83ed9e40f6bd5ed3442460ce9780913c0b4a18914aab64b07f
z29692f225e8f205e85dd552cec5fd33db349465f37d6288e7446d1a3f62c7d277941511f765828
z3c4e11b10f9f181c75a23b851379ad4600d01a1d6eb1f34432cbb1bdea89a39b8fdac570647e42
z1e0949deeba88b2c8ae83b3bf9df8ba40f0f20636a27a5cdbbd3b09ccc67c822467b711fdaab16
z2cfc10ba646a67520e2ff19761916e70305d85a09045307f4514aa1f67f4829b67f7c5a73be92f
zc90deadc4d29d2c0af08a505c73b610ed8b1087ac5dfb0e65c401b5bc017bb0a7c97dd47c4ee54
z5efeffa4aca8d7536fb78ef111d8404a72437b8d4aa65c8a10da26e03fd026cc5e6c2b528b2aaf
z87a80da70377f09480c85f7c01bef1b9809bc65edd3aea92b8b5f9f8eada06d8cb8bbc649b4810
z5f67ad14ba38b706ad1e7df4e12857d5b5b8ca56f7aaa234928aeabe7a1950605c043631568fff
z6d5d89622109a41814091005690f731a4740bf2cbad845d185b0232e2dbf31246070f6e9283a34
z5186962fb2df7584181ba9501dcd366d44a3b26f9b87fc18a2b5fdc67dcd3e20697ff461cae2d3
z5884db6401162602baf32188f822f91fc1422ac322bcc4293c816671783fd6a024e548c7876145
zcb4893a0feb9a72c4dfb2ecba24d2ed18f1245ac7392177e3c9297cc8a24377b6a9d62f3858190
z50afca59b9a76c3eaa46dcbb0fa579bf6226ebc9c31d8d9076da59c250c36eccb017451499c72f
z5edbc66dc747b0613170088f4c1784d2e9ac13fa6d44b53c8d97821dabbb9a0cf80d16e233c03d
z536b6ff0d3c1eea00fcdbd341b1c8462c3aea26e9bb5581fd5da4577be20694bcaf552cbe63a72
z2029c68af1d700b29faa7e1b99956da9698138afdeaad84dc3dff4cdc0578be82903a34310a397
zd385288dafccd584042a388423e2edcc4740bf8d55df195ee818fb9f0ea7c0ecb8d3a98e25f44a
zc3749daf7fc6cb238137b7d3d003d4467f9e9fb33b21e934e707c500f23bec6e4d6bced3da5b2c
zfd90f3f67e70548da33bb36ea8a2784cb174486c07f45f2064f1d512826cb75f7cc3d70431344b
z95f1d57e6737d5af0589b779edbb333ea658914968678f91f6f94a7b6e868d00277172fdcac86c
z7666f3be68e0c80328920f3868bf82477aad32a04f64f1528bf846f3f0248d3de2119027410eec
z688d8b61d531caba52d7c86d7127a7c3611ca3f2c98690108effda48305b242246ee1d33a44654
zcd9f7a26bf2859c72bda4d735b0d6dffaf3ab1adb696b1cbc173561dbf75f83f8e6e9ae4218be6
z7df17bdd8a0b39b48b3530b205df922142a461f4443d9b47752b81341aad139a3da852dd982c65
z354d496518fd1ca6f9aa10349a3a33dd9dc90e1a713c912cb0cd24ab36a1f7dc3fce13523fdc2a
ze31c0470e448ccf9435f2b69081482d5a703b7da02fa3195d7c0e307a4460a992b048b3dcf3803
zdc275589beab7c864a9355fbc74732adf22dd5a2d6e7bcc3fb974be130c7308f1c2edcfb2dd9c3
zd0c5d559600e362a39a38e7d396c196722545c568d7ae98f119a3954a67498ce46fc4655653df0
z894ec905d82ae60c925e8777f575bffe1591e4fa5e1d51d52cbd990658377386d244f279c5bd6e
z6bf55bbf878a923c257614377a273e813c5f09fb60a5932d5d84839c9f9e9b9d0e82d8e4ef7c93
zaceb03d30fe5c453167a97607c0cda0caf41bb175ba3d98cd708464003736e1ecfa68e32073edb
z18c6fe61d27d26922ec9b5c8d2454e11554a8a2782f0bb90d000cde8767268c5d172a0dab6e31d
zcd32d5ba2acef696f1c3fac152109c94189a8bfdc14da4dde24a5ab632d0d656cf401ce109d1e6
z467cd25efbdb6aeb7aabe584dce3054f754b44fd24f8bd73c4b4f840604bc7368e53caa2eb8c09
zef93df2c7fe5f575e70c21d7a4fe682df79b4ab2b821ff6085fbaad110314957e9e35ad02a2ff7
zdfc465ddec7f88cee56e01cf6e2dc6c17de725b88c7451152e762ce8923173738d0abd183d1138
z45febed00eab7dfcd681d5386f043f940baa078ba07eae833ce62f9b03172a9e00d3401cc42ae7
zd18e9cd0b0569b36b2b7ccdce1925f9f5ca34c8197cb7fb91531418f6d01ad1995fe5589ad69f1
z82dc389ae79f41c8464f871195ad3e9ffa41b7af510971652e305474ec3b7cabf536fb79f0b2ab
z270e164eed0019bc5c396278ac92f58cf719794bd5a00263f3cc2bdef75f52d6d8e61adf57894b
zfe7d1df83daf79224356867ca2b02d8228de327b72822f3d5035c751e4da5a6183cd5351e8bd49
ze1433cd5dd014bb78921d808e964e55aae6bccaf086c572f9fb969e41eb3e9781f9bdbb71556c8
z9352bd551d511db5df138854584344ef0d9c0e2ee7eebae23b39a072c219fff5fc6e490321fe0e
z54d3d6db76e6e72e10637a96d4e6bf63bc3744524606dde43c3dc6ada244b2e21b1f907aa00089
z46cbbcd6c173cd4c6656d6da20a6c805d9ed6b379623a6570d6d6b0c77a700a547b261ce9e523e
zef045816c309bfbde178eee5e813076cd48eca28523f3f113985e8067acba257fe9dd67576b392
zd5b0df7bb93b56e0d64b94ef4eff740db81e9227c0e65da985763f87b84cc399a25a423d874fc0
z896e686afb921bd462be97e1b40bab1c24837f4f6a662f5eb025a3ab2c9304c3a88d4b1f9fecc3
zeb494e5290885a1520f2aad57482416c19ffafbc29d2aa2db3167b468f0cc1e69542f7b86c6b0a
zfb3491c8668e7c960c9462a74c46229405cbd022382024c2182ae806ff04f0107189bd8ffa9cef
z8e9d69c3fecba095cdb51664b6554fab4c1cad2b546dd182f8f68eecadc65d414a630b592d8b1e
z68ba447b1df3048763857e1fa515f6e2eacda246d9c5c022203405c8d6bd7fe96a7dce0586f602
z85fa3c6f66d19e18094a776fb78632cf717b66cd4a813dc4f9ba3710078508ab622c4ea38bf1c8
z12de356575c144ac6e7e46a4b87de0c43126842bf48b4562cd70190633997049220b42fcc20f3b
z66f899d0a21be90b66a9191fcb47a35598f6ea11bc8a44f9ec7b2d4c6e2b4d9082b1adfd2d7353
zf51fda1aa01531de09acbfa5b04852a7b595927b32e3e9afdddcedc15df9729a4045a38e9ac2c4
z13250c08398ed2e9434199efda0b4b15b6f5c27ef6768b1b30a12aad2b644f0d8c1c9453b1c1f7
z139ca9793a973ed7ca3b632d1fc3d6254409d783ba858947a6e9ecd15f06740489caf6bbed1586
z35337dbe8c7e88904c55d7395de6522135a8bfbe7b107a5f276df6104924f699f425f0c095d7e7
z5acb08be315c6f323711863bc404a5f8e581e4cfc63c00b602a1a9b105a96f0f4be9085fcd268d
zf285e473db6e4b4066d780ffb4b68623518ea201f1075e0cda14d49ae1acd83d2aafe8b4b72bf6
z90e162a2c7369e2d10285510425cb2eec1cab62b231244eee96ff592cdba89a1d36757c1c2063b
z35db79edff242b3f3dbba572dfe04e7ab1ad1b9248f3c1db8932d5a9bbb8194999a894b6ff71d2
z62ec06ec01a760da5b8d1af3556fef7b8f9e94b42dd4b99775b66409f560766e296109cc4db94a
z59afcaee0579a6e67a13ff51ba29c5ce532ee16438f4a61c86e7bc2761df9d13ac7aabf032a771
zba789145c5a05953615ddd23cb41d6f45f895bbf4672a98ba6a69a81f21040d1edccde98ce4c93
z4e4916d58167031691d0b0e9de4ccf007cc7dcee0fe5feb76be82a9d79ed06bedf500313d78a1a
zbdee3faf3874c142dc5634a882e67b7028d12eaa15aafb564aebdf88b5ab56f34deb45511cb200
zdfb3384d2febc6032fe22d136fbc9c714d986701ab66906c90f9e04765c4aaf030eedb9eb28cd5
zb229149b90d04055d6e377e275ba4ec81530b9418604cb6fba11e615fdf81b6a02c4affd526ca1
zddd262ee8f215a129b5bed879d90952087f8bb51c76395630b591611452717242117dbbf263a80
z3020bcd2d5f843e0ba0a07903915b7bc9aad8181431b2519e79a33c5606af4e163df9e39fe2816
z191fbb0609fbb1dc0d82b75a3bc1ef341e5f1764c08337cf1998a2980de0365616204fc52a1178
z4c110e0d00e389f981cefb8654895897303a24867703a0cab555f9071aa6ad702f217382de8674
z081a8755b051374041d0b132443c362531de7676d7969b150d2c5082ce2575be4e0a515d62dd0b
zeb65091fce088ff3ce2a314a17bd9b47d8fbb9a6296576f7059a9d216a351dcfb514c1746a1a19
zffa2329e6835ba0aa770debb33ec1a80bcf0b0d7ad31e440d6520457bfce447cf2cdac8064346c
z82b174530005024060da8dc88726fdc4aec0cab466c5a7667c69073fa152e73ee20b58892b9081
zf08c34599009f2a270ab5066bdc8077ec36c6df11fb5776ef88e52e0e31a0ea69023e30db5f81d
z8d555988309cdf75f8251696b156fdf6c1667abf072d6f0a6146a9cf260e66fbb57ca647eeb9aa
z261b56855e06a222121d4f598bfabcd4c52f5bc002e1494731b4106e31062e494e66d0131fc219
z397f099d640eb14c0e877b6df0c1c49af56ba248425710f5c73a2a09a9ca3f86a0802b7d769e21
z1a80e302193c39007be5ce0e4a8314d1e34774d4bd82e27c1f7e66ada522256c0078cb51077fcd
zbb2b9cd4375cb1d697d2e4dc569c02aa994ed368f4828a0b4da952358323ebb542b0c832c24e75
z1b3e816c2fd57cfbdcd2d83b4735ecb0a5800217564b53a277048c35a4dcd60d0468f81eb9da07
z1c61eab9eb341bc8cc2f5cc91cea7d8d08b5a43da5be1f357b5400943089a914e955dd825843a5
zfcce4d3e4bd862ace0a3e43d4ce89f6b2bf1d52e6fc7c2ded3c6c38b8df3bd8a69506b74db02d3
z3815812af19b0ac3e465848a3573d2802483a4e5b3fcca406dc513d0d915c97c95ac235bd42972
z112bd82e5f3eb9bc87700cb6bf6b73a1b3fc37c3cd418085a7cad9a6c3e55126ed7d9e98fb6907
z045811adea966ad9da32f1410cf09ed9087212282dfede62a6b67b6fcc39c1cb6ec3ac8c121d64
z504f95a4afc5a341d28cacefbdf9fb822f719c6d1d60fb7ffa299bf88de88de83d340127bd594f
z50fa58e47aeb1e0e1ed263a04188aaf64fec90a1d1dd82cfdf3e69b7a1314c24138a15997af8ea
za21f59b17c0a1799248790afb37fad1e4050608fdfa847647963302dfd42bf43cd40f90f3b6279
zf3508fed4c2650b1ebd255a1b561980bd0b0b58cec7746c1989545cd0f566f946a26863bb2dd55
zd41c91eb56b35dfde136d2d5a92abf7c263ec834baa21e087c8ae43c054024a39c78f24e3edc8d
zf1f3039e42bddfd37dce506dc8f98ffb205e49f4a0268e9f67e4f3702865fbc4b9984070b4f451
z22b07a230c263a7e4e7490024d735031cb67cbc449243ecc9b327b63cb0bafd356a46df266aa42
zafb010d0e6adde45081c24a6fe7a2053376252483ce6baf699c2fb6c719383e71a5f353b13c30b
z85b57f9903501647165aa565509f212121cc3be4aa1ce821b03541210bb552bf43683f48ea64c0
zbbdcf037b639e3f2a357ab44f02a43d6f74bebcdf3f58203b102ccadc81e4b255705b4708a16c1
z48adba577470e496cb35779132bacd4c7b03bb6e1bdc418e6e2a5ee869066fe678e9068871347c
zc2235430264c26bd973067c6b97bf3f7f7dfa7adb1d053d23d150135704b1baa6b8738e2d5e146
zab6c1bb151fd762e9f9561a1b916fb119d1ab35ad8f32769534492f1e11cc965b2d405cf0b83b5
z3565c464760fbb58ea48270eb0adaf75129e8bc766c013ed1acfff3374704b87805754cedca681
z3acabd696fe33ae94ae06db0b20b86fa9c9a6dcc7d0410044b134c19a25b3d94c709f259b8f5da
z9a62ac859076a687ab721784a153895a03643a33988f2cd6862f703be9a5bd010afbcade1b8a93
ze735b1fef170dfdc9eae5371c50e7ca88bf7250ab422a0de2bf18deb6f8132dbb27bc78f368599
za8a7b46b324bd512b33053ee8e874ceae24b6786d3a9e1493af31d1700f082d2d35c94261f8f37
z3ed69a85510631167660fe3c5330f75428326ba93da0fedcb624439f1d8c4680bb083870ac5d55
zb17441b038552690c27abcd5ade86bb1bd83257356f17c8f8546e7b4e1d527808cf1f1aba35d79
z86f546eff09e924cb87e6519a435269ea93f057ef726d6920b70d639918a57b610a5276b57b607
z469b793ff944a727a4048db2498edcf992b1f05d87c69293424951bfc0f90ec4efa60bfbb8ee9b
z818df6a19b3a0a9044a3eab405013d778ccb7987ea0cb1f50cb331d087a5275ed1b87a0f31b32d
z5ab9ac5c22f814d2a6393924865ef383de1e63386ed0a7316927a3fb4308bd9a94d57fcd130ab8
z40a31417da0533c438c07c1b51d6aff48d17715169504ad57244c15d9bdfbcf3e44bec1233fbc6
z32f9a1a2ed17c9a28b410de77d39a262fc00e548b3ceb29263d937343f57165eca301606662844
za4f03a1867771b503ab4ffc1841ca4e82f5c2757d813b39f6e05d317e336680b0111488971fedc
z80935cc550b25f2809e9480c99a96086290a8cee6107d05ca4f91fc73df1aba9f27a88521bdbef
zabf5a300b716ae8a9a3f97dd5d8e8469096658bbba42b065dd1d09b266646b5f1c878ef863165e
z3a2499467307fef75d5c4d149870b8011a3e5aa1a5ad7a44dec3a384a04b099af1c01610207a9c
z019ee62a9c3b7fc09b4483b27e4b8c96092dc58e36048c806db7818c8b3ff470cf0506970ab923
zcd0a7d885379648b05bc08aebf84683978e6e718fab8240b792edccca50ad51eca154361883cac
z61fa538080da3b5a409542d7ef4beacf82d3c42ab8cd9667a5c4d01d6c6063f8cecc84ba2ba53e
z715a5e5489c2509856293943b9def3916bc53491127616e3aa47bf4703d2176b4925c7076ff801
z7c0eb867fcdaeab82febe65684769218f039877e237465c8a20ae3ec33f371bb155a49beba4ce9
zeb04d7ec8eae5152fb5d9bb3486ce654ab17d8dc479cc8b34769ff0062b66aa5421c9c71ac0283
ze574b43fe5f70f96c9c18eb4841a3f1a30a22b079fa1b148cddbea1bf44f14d6bd871ce84b2ccb
z10adee3ff0a3e30493b19784d2a852f9e6acb3814545a914d02983261d57022b0739a26e20f00a
z70cb68546b9ae8fa5e0a79d10e4e487dfe2187db202b2fcfcd153f5e2397285cc3e8a8432ff89e
z7f3c2f6fd39b149d7ee46dc49576c8065c11de90bc87b043955fe2751f86235af6400dbff91f6b
zd08550a2aec75da290a772e55db84f3cdde2c54296e4e534702c413dfbde5135617cbde962281a
z99abeac986815657383ce4f751baaaba7a521a09cf9e036cbf6fa056fc947b6990d55529812fe8
z42766c3829a0e5c1434aaf735af2b7e2203a8294d72ece17cc44d0b7a521e9ac21cedea1533bb9
z9ba874b7a21eef2da5e0b3bcbabcfb10a39d8d97b61f0fe2480c4aa84926a420ea4a1160855596
z2cb8c595b4a2bb85e8389c3c47f1b5304968d9f0d81ea5ec746975db1d4cb1dea0539e33bcc15e
z0645eda166d24a8bf264fecd8b40d7e42a4b710eb467b681e4a897e276b58d2c0f2120f47f2640
z278b86b7f5b2db030063f9b45d2e1586bf48c364a6f3c396516097c16b7090d664b4d396d84dbf
zaa06da3aab86bff020720ca15382444e3aba85e844ed3951672320ec0fa37905170fe429c7579d
z306a3d04e02dafcdd2c3ebf61169b941bbf9d02f9a5767459c0f4c35e08c36262db84176ba7531
zc3b593d700082329093257b817fe149dbc3ee9b4e6c1a523c69e143e978b6e4526916f35796091
z1081b3dce6c28ae491441dcf3ee4dd622e27c67c82421890ea56cf8b22263fc1e6d3e2fe0436f8
z03f825c2259f2e67b0ba61c6daac5abb2737a6d2ef229fe69c0ba3c9281d21a353ce93f4e04288
zdc8f677c3b476ac808ffc20fb6b241cb7a93e430de00d85d26d6926cdac6f77c90148db6832f97
zc25e5cf566069a527381356e99e7a6cea8a3d3393265b0326d94a8e56c090e8bdecfd7a4227b71
z86175f0d9fd2627e42734afc665687b6eaf87b8a954ca110e41452ca2d13b3eff5fe46f36e3fdc
z8e8df02b6a3f20cd49b8716d11254dcaa32dbf2c9be3b526fd2cda5c159b03fb2bb82e553e87ff
za43e48b05df38b5e894132e16f444543b209ecd1761e80db4556b87750db3e92aac0371359c126
z145fff9d8262bfcdf6a09ec7c3e4efbbccff78d99936820f3032ed70fd96817dd47a4e9355ca6b
zfa6687fa7ce3a35a34c0db9bd832cc07010cb5df09f38a79172840536b99474eff615892ea3d1a
zb889fdea4184bfa9dbe1a8cc47deed27e7dcd5a8c466c6cd583c2f4fa96640d9b024b80428717e
za81ed72fa6445574e89a67e5b563e41ec346ff9a58fe0cd372ffd27c4bf8561858fc7c2908b925
z97c625656d6cc10fec5fd5449d8591550fdffce74840a30e11083bdd93424b491185eefc49a325
z30bf002f0d4470e61fd97f2ed71b9c3df14dd56b3de8124112f6c64f8b65a6693607673919ffd3
zd7ed86102d970ef0378be207e378c2a3b32d794b2664556a8851875b2d4f12e8ab3a1cb1b30192
za9bfa1ff9ad64aa5d1129d4c97964f29cc4476e82190400ecedf2e875b58e11a171406e78bb75e
z97dddeca85b238587278c44d55197728f7a78f5437d8702455a39eb1d020d587405d17612ac2d9
z39d3aaf0d554316bcff16c6a55ec524f77ae9e30a7dc4bdabe3362bb7875cabd57ecdddf5b6edd
z44b39789a2e87d5ea73be9fe0d52794a3f9f28fc6a724d10bb5723087123fac2d58a8bd1d27788
z2b721c7fccd5cad94de9d2b90555159af4fa481edb03381dd87c875310f72fc7c285d95568d25b
z67d447c6d53edb7f4f9c136280d24845963e34ee9a43b7c7c740be05d2bb86e4711ac944970b5a
zf4b2820cd77f96d599a9714490537441b33c535bac784fe186b3d4af5961011d374fc6aafcb3e3
z56998bac9565993047394930016470ee94b4b76d7ac4d112c97403996bd75788b239b1b2bdabb5
z9c11a13697106c3c567ca12e6617f242bc4be99df80e844ae25f14bbb5e0a4135c113468fe696f
z3754324acff2c496889a9f41e2715d21a3afd86c9560eeb32a0cc54e730bfb2d3c464644c2e835
zfff3ddf4cfa1b8093ae0a68f214f4a7ea0dc0be7e707a50407d633727ab4c286ca4bef44d3c50d
zd8c789346da3d77913cad9e546da227573e7de298d533d6d4682a13b105c63b48175b132147519
z39ffb41100d0b71edd228910aabd43f839e4612548f17e9272bb57cc30a25a2c2c96bb8b264129
zae0f4e992ca14289c00341d7b4ef01bfcad81a19425960e4bcc766a595b92d84c198d45471bfb5
z39b475ee0c6dd8bc837dea8ce759f16ef672d1e65c38698f8b1aacdbda0da78a8a46f150a93f2e
z05b9fb06deb399d577a695dc0895d119d15065784f3287f9f1d6290ef9e5ed05526b831466889c
z1e132d9d8cce1667c18732f9b445314d9815ea5a3968c1139b420d1d5fde59f1fd89148f2ae8b6
zd7ad1e629960d66401e8cc6a50c86bed2b13172e435999305198700bdbc7de1919b2b1210877a6
z5abe85d945fbe0793fc81c7a2e0bd94d8d0ece613de3bfe3f376ec945f8ec041e3d4a1cbccf976
zc9ef0f77618d5308118d384058b4ec059d2f5105bdcdb0573b6c014f5240617cb2b020b097516b
z2e098a8316d3c6232e58c147f6400aeeb39bccf7f8717874a3e65568ef30d183d4d1a12a9a7177
z246dc3e953e8f64790a6e3cb71af08e1e441401db4bf0b42c4d9d31a87af452f229c6055212bcb
z63864cd13645ae076b20dee660adc82b7d19eeee996577253cc3a8bf4a4f3a389c43b9029456f1
z38c54bd627e750e50152490ff4dd06707922809ba2f0d2016e07a02daee9bf11e02f397be50266
z7b2a1a6af6d1e9bbd0b5dff63d707f4e0338a3d11895831c846a8fa715dd9e9b1b33bcb6944119
zb11c4f5f4bde97122b2fc1aab3457b2faeb8012ad09ed5432e6bb886b6c059551460b3aee9a060
zfcf7b9e8514fed06a3c4c449b851e6a60f9ec1ff198b3b28163783e614855e279e40a8c1422d30
z1fd2cab3070ae6a385aae0307cfa430e382df7cc692f1b0e4f28274d3c0c6323178ed9de601170
z94851be48bfc04409fda6bf8caa509544e18e88b0d2b5adc72a4089487f48b9ae35bffc5739e01
zd8703d35be1b9cf42eed245535769653928ea7b338e52925e61f7e8f7324561855050cb08068e7
z85cae598abc06ff4fe07f1d66465832925da92c5010a17d1a4ddca616900d449b3c661fae5c2ab
z96fc1a14cc7abea74d154a79c53fefc7a8040f64bcbb71e80e5d1767fd13972f7adfe07bf5897f
zda83dd6c50029aebf1766de513134a626dce0a93563c2f81a8ca7fe2855b635eae93cba6c28bf1
z5e895ebbc159d0bbdbbb1a996a35b50a4701caabeaa61d877231c0d89da42681184be70f505a5d
z1e5e522cbf70e5954ef9b64121f05a24e862d3ada9bc6a997c3b18eb8651924158e9949308fc7b
z8a9fda98a6dd5edbe4c2aff811495881246f148b9e1fdac65c739efeb69381365368841779b716
z9a4b2c0622548ae19945789f66518d1950508de59e305f4dded63a2d91b8716706428094b519e3
z149b00859653f11bbe86e256531d6a197d2797230a03216457144a5bf3a483c88e2e4b6a8d63de
zb9b7c6513128c5fe417b74a9a4c9d3cde43699e2a68bb62eaf6f0415d764f007f8ab109525b828
z4947f0ad396588ea00efccc9a47eae1fe313558aa6020d32b92e9f79fbc6d794f25c138ad0dd85
zb40ff7666ecad436239f03bacfa7e1f84c9e5a78eb8f712c23178a22da2a1eb1c4e235ee1f83bb
z988d9ee854d23befbf80f0e36a4d036c4b522d65cd7c526c9ee7c6a6d2beab8984b0546dcb01ea
zcffadf0d6f1de9a415053a69a8e5df451f9c9c72ed9598f9ab1b80a3063510801a976b6d26958b
z4938beeb6fb7d943939fd11eacfa8d81db7db36dd44e6204c8de8f3845ee70b3b613aff62649ed
z633548979d4ba18100b1fff892af967f0fa2d9a0e6e6bf54d54bfc8a88fa31c33bee5cf7f7996b
zb640dac605810472b0528f97dcda25b6c04f54938e6f97fe29963d76c5a56d167b969aff949aee
zbceea225ceb8d224f62b2ca67908c7a67524016756b60760fc6aa8221f2f0496a6236b5368a548
z8d9209dfbdcffb922a29c9a84dedbb587a32678388a0713e9969122ca2ac3af956f4059e050df8
z20fa676f6d44b0fc11e93206b829735a206c55566a4ca54418984c8768ddf454beba70a297ccfa
z68cb0313dd801fee566586b69059dcbf54fa1a8d26177f8f847ba02af89e236db74fc1f87040b9
zadb5fcafaaf73db4890d2a13a53c8ed7e00b0a10a8d81d49b9760b86abc8f54e42131505820fb9
z616c045ad6c2718b031d51b2ca4527998544a75e023242765c089ae2b29a5f6ba64d33fee7b31a
z4c88d9241ff0bbe12ee902686d926b6453a0568ae6f14bccd4fe162c3fbce56aea09a8cfe56929
z08f2be29824516c92ee13db73595b65e870b0e279d01b20dc8f6c65567a8a39356b5cded87df8f
z52f7b2b52c94ac59336b29cb1b10a21adb42fb5ef737ab84f62ea8f0a86d1e0ed6489bfaf81e1d
zc22734995030efa31d3a7af30d0ed4306f492de7313a4795d5e00e8ccf9b8fe0a753c427fb8cfa
zab9c47a2b9aa0620af320c6733ffffe0f0c89700e0d374ab59553847d12236a53b23303892c2ed
zbb310868aaa49ab5b8e9f298f0860b822782e29b978400ba440747a0d535327d8865e46e3b08d2
zdb2ef13a8ee1da5614745dee55e92565f425c04d014adf32733388e13ffdca61544db8b9ee2c94
z6a395265e5b87520c69daa5019400d745c5906f5f2f1000424c5d9c0f85adce27c68f86a0d974d
zfc1ef28511e7a44a0603e04f0374d8177710f8e048d5ff06932a5851447e867f5a8589bc302f96
zc2b728cfc612bdd50206f4a1b7f520123b3650b4c003cc9050865ad2c5e94e1c7b0fa9a3563ce3
z813934d97928bc04d483849eefa6459a0fd4e94b11b1ac807b42d674d921111c42d63934bf1a16
z01447200c1c682d9a478a41e832f9f3db529099ab19b561ebf04357ee3b6fe803bd1d5b8d91aa3
z53e868dca8f1b215ae351373a465ed9b24e56103361eebfe5d3674478a287a99647784a80a27a4
z6db84b79a8809526e4101894bea97d7a54033e9ba048e01273577ea4fa6091c882919b93542e27
z50b13c903f20762a4892d182897ec299118b76a5c8147d5ea4df075ae65a192c1193cc8e169da6
zf00984e186bdb89f852ebabb26d2c62585f54c272736bce3c42e6fac0578c038a62a1132a783eb
z7ce738addcc8932bebac05b46299e202a3d9f5dc24ad8472ca3eac5d7743ef7205d588fa4dcd1f
z10115e4618269ba5080ccc2746f9870111590ec7be6f24358fc6452b4c9c4b614e5cd116a55da5
z423cd38bdafcab5b2f0a532b67a8ef209b42768d182b294a0085aff2ce94e1736aa19ddfd26c00
za6e43b184fb5ee42b1c29b60e022f6f6b1cf7afbada987219ead8579c21a97fea37c163c13129a
z4f479a5190136e7e0a00e488c31a195024887c3c67903c718bb441b84ca5ed4aad140d25205680
z5e256da87ae1835108dbc91a6d8c02e3c35e298cd0e5eb7bf11c5eb901336697f99d108cd0fe40
z7effdc5dad9fe5cf2185dd81584b7f4b9c78152094cd923c746f1b1c7944893f24e0719d7e27d6
z11748c06175c9a47b3700c75b42abc18b6a7870f5e69d11864a4acc1ecc17140db560802c775da
zfb9c78e08681aea11afbf055e7741b464188b81a92b0e6e245c0f96fe5deca7bf1aca7200025e7
zc21ff0da58a60c6fc56400278ce647d82b9b378d3ef6b90d75d0f4be43d4102cf34ea84057448f
zb90179b270890e3ae82ef4ad3fe887d4fa9b03e136822d72dd971b2ba1ec47773f7f964f9b40c0
zff5a210fa585e5e1da201741d38d418d6b04a37c4772db768e1b176d81d350d099d61a0a1d02ce
z3adac5088e8a24f85b3c9ad3d91337295a786db27974425a23b6ed3216d73daf917944356bf443
zc039193255cf27edc295e892270923a76c5895f9019b13ee40c7e9a46ed3e3fd8b4d7d8881578d
zf515d97846fe163af0275dfe1689b8ce7a6077c1872906718307c132e2f00272c085e2e81072d2
z8a746cacd6b35e164717a414b39ca58a1190110caa67b10fb5a17546c13a9ac2c2155d3421f4aa
zeb96f9b470bc172286f57c9f7e77f6ab99c08462716458a420e2f9400da0f14c5a64a2e15e0f36
z5205d1472ba2ff81a5bfd0c934665590fcbf5701c0def2d6da537f7d82f658c3f32dfb1c44ea02
z08cd1086e100db2e7d1816f7ab50a7f5baeb79cbf49dea69cb4bf4ddd66cd7c4b4576f3823a57a
z5a9605fdfa18b7985dc79abc3131671f41e3638aabca8d31d4943939f5dce9b7f2a2ddc4f314d8
z318b52216a4851211f986d3906afcb5749d972163c5479f24b443aef3f9d6ed099dd13df70f0c2
z51705944286e5b4bc5fad58c5633a75add62182514ef4e019ecc191f3448a8979ffbf8bc6a5a62
z6ee894172d6ca06af317e20dba6172907b64c759085b43f870f6942d13e9408343f8c2ff18186c
z7fe9f1bd109b1ee5d0f885f67a4d019c854eb4acbb5db131748b3cf8501582ace1d2031ba50f25
z540eae197321672e99c690a89ed2b52b2018a021507b31ba0521d353f04ac0fc32cddbb3c1a543
zc8c78d16160be83e5385ec87968c04391eda1a04324e58e150a16ebe26e1d7bd106266c36d83b2
z1c536d4794b3edf8481a52c1c252e24fbd30cfd796687ecb37764c2be3b93eddecdc3b2792550e
zfe29369c33e71e5d7f606e9e3c2164b37f6266b25f837e52e0efdba1f4b917c140468ce14a95ab
z830049004b1cae1697ca78cf7ec1949ecfc2c4c50e81cc2c18d51ec8ac77af9034a177f1304c92
z16d65afd1b842cc7e9aee7db29674e69c0b88a3c347ce6b544c02a3c4c8aa6253b6ddfceeea084
z91adb5bf2602da6031c3441ab581d543b45150a2d48799e31909bd3eab1f99e1d280de095fb701
z1d3db924d9ec0a530caf5315965794e3b9f207a330c92b16d4545bdb9777354a27c0191da7ae3d
zbd3c205d6ead887fc523d8f2f1fa9e6b38d214ec3eba62d864364798d621aa8585384d266b41d8
z7ff4a87faa05b3d23dd0298d89373b19ad2dbc799a21016e9a865805747d9b142adb1588472f94
z3932aa3f663427eec205a9b61bd9277a59b9ef15d4301eeb9096773bdd67482bb82da6f3690634
z635c9ee658f449c4b009a456fd532f083fc7f71da6257be7ac913af18dc2f2d7df942f0a95d4b5
zbf03143ef0e5da605bb3c1229360ffeac267ebf3b60d5d1b443bd6e5e12353f0cdefa848c10f7c
z2336f39343cde1ed0257d54f2aee824e8d6f9941751c563767d0f20c7eacdfc49da646acd753dc
ze5d936e50f35d75856254a49c981a98602d524ece50a73625efbc5c94959b94a4584a2e6e65852
z3e98e07764940abe654f024a6eb2911d855cd47ffe8d80414592df2118040ea097dfe906e4aef2
zdcd623dfaa68688b38f344c3efb9f5b8473ba15ceb5de480a9ac94bf5a2150633b216e49f99584
zad123c8be9aeada34dfbf39ddf17f52d82ed44f1d1085b7215444a23640e6581a3f1feb24efde7
z9bb0c0bcc7ed6e8efe8ba259998365cafaaf52474194f1718e6f619af72d206fd989c928ce738a
z2690af2e0d212c9516063b238a9d4fa83f187a8a4c92584a620644646e8d309d18ea45cf2a75b0
z6cdfc8a94958637149b62814ccc98e5e126eda10db03f3074842af027d3523892b88cda69bb53d
zbb7517cef02142783bf97eeda0cf1277d076949e1f1177aef53110f33816e474ad02e66ec8e892
zf05a0cc6fdedac16b352d431c06ab205bfde1e00912f421c4d40c48d6f0099bf997dd0a8cebf73
zb9312f52d65a2f49fc3b4ef4268dc0f0aeb44238f3d6447e1baf8be06a4dc6973a9e642c84c23a
zd904a44cd48e06909ba6de2b0cc3d4176a4e4650743f1c64f9cd954226927a6e445c0fca7d9bd7
zecfe356408fb3f75c33e2002a8174e4b040d83daabcb983b5d3fa32356a29eed04bef28d649e0d
z04a1db8dc424bcd238830ff6356d35a8ee035e97f61e2c4ab0528a8d300f61badac30a327cad0e
z0cdc005eb3771ec2800162b29d8414a7cd328c2e1b8ade6646b515ad30381e278de604fc71be69
z5234ee069f05a9a827b2fdf396ec6a7473831b2143ffa9a6a66d223e4fee4a4a77d1fc1ca6ca2d
z0b0bdd33a9ecfac1bade0d76f794c72c61daf615c468c7cf01a395f7c6b58736dcb2c3777450c7
z09826fb9083980e544b8832fa584af7b116c567fec57347161cdb3ea0155afd827070df30cde24
z6b0811c57961e0806ea4afb1f9d51de333cf5bbc1abdb521ac4a0a45c1e4d0955ec89beeded39c
zadbb5c79239eec906a068938fd86b908737c383ea004bf63485d02928c95b23e941c3063dacaf1
z1ba74e524059fd80383ff7ea589ba12e7aa88430c94ee00b238562c7645cd4b49e3223cf274f2a
z49beb8a8bfec9787de7f355605366e3d617e7802fca14fe35a8e903c965754eaa0238587d155bc
z29ab1e2379125f740972e22094affcab024e54a4904100f00d9a2d75b2c0c04d85f58cd62f4775
z6908d38661ef753572eeb9a3d17511c5f3c0754e9726341e826b50993888a96266905dfbcd4d31
zbd4711ab356f18bbf6a7f416f02b4faa101aad129759b42c8e7c1479112c71c03f07da0f92449d
z0b33db2c36868b534f18b28b21606be81de0320fd7c329541eaa3d8a0a5b00cdfa4c677742ef36
z9510b763e9540734cd531644f79de67623dfcf84e6b7508496b3016deb1b11ea9b6319740e4458
z40c32b730a870f15d29dfbf6b1cce346641cd8fe2257f9f9edb8100c1b90a35d33bb93b8be8147
z4410e31c1d14da3b9b0a3e019cc9f9d89ee1fdee0448b59ac3dd2520a6c24ae7f0126cf3f85dc2
ze2b3be6069db8e02657e82c6da634a1dc328de5f9eb393a6ece2385adcb05b34815aba90a18093
z8c9d9a132f6995671791cb0be6463d03276870f740f3acf7647595a203cd9cebed3cc18c407414
z3ffab5a08fc447e05eeccd070decbefdffda066e298d99beecee605c3efbff2834fbfa2c9bddc0
z4efe9a45f00777d47d5ed05cded6e07bbb45c526e2c7ad0b05f42044c710f4c8a9442d893767bb
z354247dddb9c8c4ca20a1a56a0713fef5e2ba60a1b487c341e6eb34c7f06ce0c8baa3230a93ced
z67860a914e25842fac11683c7642a2fb2a852b3623f42b98f92e1cd0ba417c3d24fdab2e20d7b3
z59ac865ece253d4131b17b56cc7a9ab0a3f2e425664afdab9bd6a9bec05fdc1e5175a923c6f8ff
z287a0ff8d3dc79b949b5b095c24619a7b3ff4d374312280027c22a7fec2e406e7fe0ae5cb9dc86
zf035afe50f4c9ce9203b4b234415525564c228a542dda4aede6ec9c0b64de2b1f3c2626cf82d25
z1729f210c9665ce4ea77374f7e32dad2722b8215d6c37489c39f2fcaeb66dbc6e570132b4eb7d7
za323a88cd37597a907fa77fcf0a1427d844308d7567f89a9fe140e61486a7f3557e36a2f485c1c
z458901187f7709fd5b492ec4f65b18bc3c16d9518c21321de188329b280c954f232ec6ba7ea84b
zf0c67cbcfdc3cdb81bcde4a2b4702c96bea7f5224087cb8a50f01aa729df56d0e5b8916880fabc
za6948c4b43e25577a61b83dd10498cd4b472883959eca2da4913f26ae063f7f04861c0812c742f
z8bdf532e777abfb33802ff3b9fb8d7cc7724d5ae64b515ced341ac2561daca145232e92d127a3e
z8256fd3771b490a95b97f2cb4b0e2382ac2846f706dbd371235a033f5b4205f22ea937f5acc8a5
zb784cee25b669d7c08a9d81daa072e1ce75739b1981975b4750d9e09a7058d2c28e30440a3f83c
z606a8cb815e99bbddd45644d486eae5c737a21396fe9d711b42f15ddc9bc85fc06d304adbbc5fb
z8a57c19d4e908077e9420f4ad3b4f992afcd14928a2a9272f7ff9148725483a753fed5f2a761e0
z181a46063726576395bf37d957a02dd23e768071da4eab9e4e3c566a61b776723cdeebef1cd41d
zfca4cf59b700cab22316f8f7067b6a1d22540a839a98caf151d7538c47c8c0a8ab29a1416de3a2
z736704f8bfe5e04ade7ef6a3e9e8a0ee22f48ba64d7aab8951e0142263419b79e636a055467c59
z44d6d3b807557f90297113216a15140f791a10c9df72060330f14ec4498dc828504e61424436b2
zdfcc07e96ffc6af0ed3db4e8d395cf67e7e688c643a1969d208b262d39684862a8c0e6c1be8dfa
za9ce7963200efa7abcf8555b77dfa2b3f5394d1071544a4d404744b048ff15e88e8e56b9d4a15c
z0611c3df79e13f28d0d4b3cedbd6b644574f022f56336db73bd721de27a2ffece50aa17f1e1d34
z203217104c872e0bcfc0944989a6b9b00f46b14f596d7c2f53d386b993fe2ee4cd7a7a8d545d59
z6f4c28edac659490c35537d207b9082923b91811e745049f4b3b6d55af93c9b2d9581bde217a4b
z6cf8511bc3736e6017a40f8f9b62d4059ffebabaa9dbe72510bce3cd97cf4586f0be69ad3442d2
z0efc00a6f102fa0fdac458327fded2480d44214664a8d673b2a87611da8767be2bd134e6fe4dfa
z47ea189d0ffd513d0033cc8ed4ddec41869037f72e1a852cb0d1558ad80521e3dabacf44149655
z6b78c709cee326e1d4283edc175efe7ff90bf66ebedb47a12e8c7f7bbce392c29126ea28260f3c
ze81c74006dd7af6e95938bf33e0ba23f34243ad3b72095f4d91746d8f1c7f63708c3b82140f667
zcdbf00ea923e4d4fe8be758b759bb0e2e2d44e884d6f59d8787e935d5bdbaadb032a582547ef4f
z8c86d579092d30d07d9ad41817d8a4443a537e5b5c8e2720a6cfaf268e7cae6ce469a7069445c8
z8af42248629b32ec4c6f43ce948cf6296b80390070e8062c7a0e5c80b4d2027e80bea93af3a45c
z7f7c91873a5b4fab80594257fa953989078ee32b85e4354c4c781a12223a7ea84e9fa4f428cc3c
zad07bfb64329a359c7907536b72b2f4828864d43563db12986af69cd9232566310418ccae13d53
z2e301ba3a673289e5ed574726564dfdece34a03e3619348f5c899bad054dccfc91307f007b507e
z8d346b36f3165a88abdc1f9cee8447288d41d1b1e1347794e0e96af8f65d9d5aa57ada78df1a79
zb3df1761f1520a9a964dc678664d335fc3807259c6dca4e6445c67cdb2b71d8cdf039fde7c0081
ze04e3c07afb246e8e39a49e69dc8e0c0bb1b76ea02429c07cd5988d5ee972aa295414c50dd7642
z047742c3d2d1113580ac6270d8a14a695cb221ff1d7fc600d8dc4a41b51a6ba29fc4d5a3a53824
z806d72be9b6c773ee7190cdd50884d986ec0eba52cc2db05025497475f360ca46920714f23c932
zddeba4974e30517e182b1178f111116ca65ae0411f5e6332df9341283008fc28bcf32cdd6b266a
zcc0e454c2e76438b404355e3c5ee8fbb4c858a3810a3adbe7c31eabf141cfbdfc083b0bedfb692
zcfd5415a02a6cefeaee9683b14afd4bf6e3f6b190fd37ab18c8d15658e82be1b452bfd1196928f
z3961f76a53933c2373a2fe78289087d1b1ba2e677b81899c902d672fa8297c8ce42ad3ad81eb78
ze71128a808546f25ef0645074ff36368fcb987b46698f2da73f9b10b92a1b2ad08344fdaa6021e
z414f374421c1271015a106b94962caaca3777c640c35fbba4be8e3ed43bd18c7c1f7ad56315e8e
z0359128605db74722e85cd8a725498b7447c335da83f8d63050fc6c6455acc34a2060108303911
zf0267841dd5fc2a907faf1dabac9874889678dc4b746d80b6128065ed9cdaafa0c413c4ae61832
z2a582d183f3220b55ac119d751c30d4f631d9f20650217b48e1db9a4cf05335cc2ee883b343c39
zd28ac0047318a60436f6a1023a913ed1610f24e0a4fd431f5345af2b3a02a32efa191886d675f9
z5a5fc05c301d91e9c36ff6f3ce09186fac72821ee4b1030b2a8a3daae20ef7251228df6e0f61da
zf5fb6fdd5afaae93895e7061ff27f917926c6625e60d444621af83d718eb014100a93afcfe7c47
z0418ddbab4a781c26e68a6b22c7d6457bfecddffa95d4c995f8f1d3333f31e53cb8193eb9e294d
z3a27931eca1893f736f749ee100d0557dab47d08ddb6a54fc47c1d1a60bbd2ea14f33b8b49d957
z1c1cf52a58318edc42086dba05bc06ad4dde6ae0789a3077637df64a137a34637d6e4e3da71827
zd16b36d512ca577dcfa8994f2519e6c8b2395e2e272b07b1e9837bd3d2a736e859ed00d90133db
z23f25e141ce47c8b3f5337b6db35d0ddddd9466d9d574be2f47cf0a4b0bcf3e9667e02abe4b897
z76f62cc5b25c160fb5a9e17de851589b58b56eb88203fa5e337d016bc42a386d6e0809d2947548
zc7ff952185bd22011f7a982ebd6039f759195d016067e9683788b7bbcefda94dd78665ee41106f
zb9d87ea08acb70fceb0e2a3776f23ad1d8f10327609770db3638ade8b7beb8c9db1ea52a65a06a
z5cca40d77ec9ca57b7c7d262a79c720df477ac20b294b2d2b194d29387b67eb741b2865c900c5a
z64b8c2dfb5a8b393dcdbe1d9811a4389b02a564e48182b5aaf0900660cf7bfdb2eda3a3eb6cd46
z4ac106a43df551428dd3621eb69cf851718e2601b4c9d7140f574a07f54f7d1ef5f30fd7c45799
z7d4b4c92bbd493323140bf2370fc36aaf1bd57cf92680a80ded9a85f556c90818b81c398fa5cce
z93de1dd38670619dbfb7a81fb255b7cfcfdb4dee2c02cc7c4861bdaccc5340c3653b0bc0d33263
zea93f302e34d47e6e33ffe5e743c0530fcf4c497b2fa7ab2121c06516733d1b0282921295106f9
zb6bbf00d6ec3be9eac254b6fe28bbf51c52f2994637a11fb1003334a00e01797ffaf0111b70b38
z8a49e375d0d9292c6cd5c7300f326539c5f68dbd66bab6d3e0a7efee507811feab27f8fd646a8e
z51ebfcb05afc5f867ac8cd192ef931151493855502d347bd8d836b7cf0a18905b90c4240372827
zd3d6a9cde9b6ada7ae597d897ed34488ebcc6e06e841392c917640d04bd94c297e4ac6f6849538
z45af458602c005f4a8b51ec9537433221baea20ca7b2bda9d0d874db203959229654da56b65638
ze1799a1321d5e9d134a9d35d97adcd56595b2b65ccb910c128e445dbd81c9b0e5c4248a95d2155
z087f1b10afac54e10324ced4a4d59a3339cf8a3706784c8532443d547acbd87bbcd0375779603d
zb4ab0bee51b75a1bc50d5d4e88d406b686df54bd25f16448e86ffa6c058e97ec4edab174e704e7
z06ec628f6c2eaa6f9c3024646bd68d21c0d06081957440fb622a4ce839a5df07fbe3bf42f3f35c
zb76a00ec7982e029a0014ca281bf5caaacf638fbd82fa6d5d63ffd6b6749a01ced8bc4d67ab7a4
z745484a16c35bc244021a9598fedac3f1c2a071cc5a61c9cc706f74e3bddeb9af6ead2f56695a2
z254b6acefbce3ad9dcfca9dc36cf9e53f2b994d1e018eef2e11c3a116193169863811415151c96
ze323b7b60c543d62defc98e70176c23238f299304bb2988149aaff1887521efc36290b2a5457da
z11b29bd378406292c051c95e9ad2bc6b10da2941a8ae855e1bf8dd736d5345c0c2d5277513491d
z18e324022064cf1bcdf56320d2aa7367fbf5764bbf3235914fc81ef61526a8da60f2ea3d8e5125
zb1a715a707ae635c971d014df9f748c0a596ea00860adfd0318f90ab5714414d58c14d2d7aee7b
z25de07dd9074a65ec0ec12f8333ce19928f82fa21174f2c9107e55909818148ea16c95cadae679
zc2b0700d55a57855a0d8a19e5b44ff2ca469f7afc786f59cc16c895d610acb3ec510bef79f6f95
zb943c4f71518d84bc6c87c801dc7e8739a0ec602bb364e888d3e1e6d589928495a80af368b188b
zab29da5880323d026afb82373bcd4cdd00093f27982e7ca15b2cfd873f8f93f44fc604fc379b41
z6ce209b0b73f2b720835be1b7d99a7d50b295c58a6d930f21478cd2c4fdfc8aee027188f644856
za89e8c5f80c963ceeef972961670b1a32bbaed51f7cd273b2ac2371000e47c2fe326121d9940f1
z497f648dac890fe3dae4086318434bc10115053f9c5b19f738c3826766655584ade526f221d8ef
zd3721b65e9a221ec4b8adc255031a7ec3a4360f750946293bc5b83b659c281758065815f08c410
z04a25825f01dc27a5d028cc9c4f0fdb30578fb1549820caf77b038d5e85409d599217a00dd62e6
z24bbd8626baaecb769e77dcb12d1bd6864cf833dc03bdb7a6143551394e1d29954b48a492544be
z292aa6e54daf813d88350df50886ee5d1172fdf35d5e678d6e7e6b983197cccc48f75a49080305
zdede87bf7022e8b5390d84198c5356af25e4a340e8195a744b666485e5ff00b72957f0a418e201
zdf2ee3c5075186c8d286f21503de5e970796bc1396778a1153b25272d0f60ff88df8f097f6b2c0
z4b57de409dcadaeaeabfce22773e2b5bf46fef95543c672c7cef897f834337fb5a8821ca69b7d5
zc60889415ff332506d7e76e4bb64271d6b613c49a3d24e045d2140709e81fb45f82ddeb9334289
z3a07ad68905dcf0a0f42ca717f035e52d89e407e3136aed5cb0bfe781b08d17696108de088a488
z5053f6e32f9f15f9ef60a216716b1fe5def807abebe7c3e961738116e1b2a368ba8ee84250c402
za875b27fa1f9826c064980f63f0e6a6ea1e1e6a8510623cef830d55f91f3c1b0e0ceef0add9bde
zf515c6a93dd849600414fb8f753fe1de9818fcaf8c02d0b4c772e1cec0d710c34658b13e729d2d
ze8de8535e2dcbfa29e75d177282033bfe5ef76f4d031e7dc50713ea136a9dd5a400a654f8cea91
z2c104030e682c17785358f3e65a23ebb9b85a4d351a83ef74d6db94b6d85ad849e47397c12ce64
z7320ec7ac354ce646f811ac58e9357efbdb797ee5fad729652d87325c7b236e9bc5fda3882d827
ze030c61054bf5d4ea9d291d532fe84b30977b65f398484d358afc40f5fd39fb36af4ee720bc174
zb37ef4d96a0ba7648b84fff8a6c281b7b9a07f06757934dd0b41286e95951a70a7505b965ac85a
z896331e1eebca2f344f12ab6efc2989372ee658cc05bc7864c5bf032964fe019f9d105e44fec6f
z6666a9498315557b8464e3865cb83389806c7e66604ca2410eb0f6135bf64a9db02c80956fa482
z03e934d70e670d67b9794aad44296b11cf14cb21cc9a0b1314a6eb0cd59ada24d26a3dd762e68a
z21fa69b4a6ff350b5e777782a4e703f3a7a5c1acbd9054e477121cbce52862b00eb6c3ec8287d0
za4fd99256312d8d3de7366f07c27149236b3a49420d978503222289d4b7a5630302b4d259376f1
z50f1ac9d9ea9239e51b4559e32111a7687f8d6cfe12f0315b16ea8696cee2ee9da9a559247e05a
z603e316b3080ab7757bbaab7e34cb81a936e0719621e547a0ea528c8549db5c5a52c13bdcbfb0a
z7843ef688b025d48bbe35731cd0e9880959e4e1a587643f2fc95ae7fbc480e8e674de6f67684af
zfe5ff960f0ef10d76025243baf07ce9a8b4d1f1463e06548feb27d30147764ffa0f3fd38321b1c
z86775769c901b8a8ddfc32acb35af74569c1e6ebf0f2fd271b20853abd4f234fea05848e3abb59
z0350ec79129e85a33d709e7b3391b0d979b31ec3831f9c93c407b06a30d6b39005b2fda5122ee6
z9e78e13a1aad48aebb221b652f810e5081ad6e5c0375eb791b7ca33689f998ccb922042cb3b271
z44b75218b030d0a8fb20eb6218ee44acb83c6410d8307612a43253b852775996f6b45055538392
zf70fb881ca3172ddfc51f03f2ee5af893679243efeb93dfce8886cf03666d774ce13aae26d7693
z30239a106f05ea195f7eda62dd94d644db698b07d36e1070a85be457d3e09091fe54f9e0541cb8
zf561c582d866e379535b03721f2cba67e06184b79be02baf3447db7e4ca0901cc7a99eb02b1d8d
zc65c9723283770a2c61bed2c6c4fb2682e4bf2084aa91bddd28deb8e22cbc6f1136ff4a32b65e1
zd148fcd3dd356b5f28b1e10aa24cdece155c77eb9e3029168902e371c9b2b439fe51df5839c53e
zbe61d4143391b363858c659b012de6e4b3144ea3117de0d73d8a3a84521927867af262f2216e1a
z07065cc5a97b1bc098c31b99734f56eb1995e825a3fe3b3e55d8a5287596a6479ef8e36128efee
zd96e254624517781b54d3bacbac44bbfc715cb09b7730444b3b5820e91154ca18ea79e48ec6622
za6ef9175c88007154ba00354faf7750d533ad4bab1038c319b3add1d7f4afaf1a5d3f462ca897d
zeb91663ae4bd51d527dc0755180a3596e401d11c16d567d22e4092861a738e98290aef2e4f2c37
z378e71eb072e9bd9ead55af3943e40813fc6bb0d823bc0db78c4a19d45661faf8885bdf6b50c95
z2da1f964a5434c2e6f541fd75ad03ec0c9409826c240bb8728745a2256857c7f8c22952ae95c24
z63c846a4f1425edbd9203e9b13a9d4565b82c5dc07e9bfca748c9979493186e5d44c9a177b13e8
z8a244860832690401b0cef96fe1575a15610746e7d13c2ce94f340d880919611c774301017d794
z6d50374d699a06a6be3420c4f610dfbe0e0d008d9793c044e083c0d683c468dab663d1b45fe92c
z5ec234fc2bcda421467f9a0d10971d0cbfc9080cb6d5485143bb7e4327f5b5ae3d6c62857b0225
zb8a9f574174b264241967f07307b310934f3ae7e940bfc82c9483d2209b2fd3774c1a16ab8a88b
z16a5ad6f42e8ddf81448fa53db5e4e08d1646191eeec14cf5fbeb24312a5de7677c05bbe478903
z3a6168cd89fcecfd46393e3c1236cdbcde126c2f1893fc137fdd3c2db7e05a6e8293ca01ac8a95
zf9cf1890ce71683013721afd93482075fbe72599570b0ee0f55023447bd2d72c1e8bfdbe4bd7f4
zb27e5f2f99aadb786ba36f839f252072532a8e264a06bb57c043320f9cab53b440391da948874d
z6fd94131a73a1902f9f72be78090898492cd967d46ac6ec408d06fe5b8fb35dca6878f7a415e3b
z77bca259278c212a62febfe2f538e04060bb06076f37ca5b37de03c887f7d81f8718b693bbc2d7
z56bdbdfb71e99fc7c8c8114875967721194aca280fc7bd3e1bbf25fc199c247118cf4ddf0d73bd
z4bb8eaf9d1ce3d1ce31ba937c0837b1c80f83093aa687bcaeab4a936979a6261945066ba3cd1be
zeca9e5a0422db3f26de2681c7a6d01194b9871ba55d14cb0ac7b6bf761d534aa5b7e4bf032c3f4
zd104faec3520a9cb1c9c8816ab530f13247902ce526cceb738ee36509b1a6bc6b08a5a400fd4a3
zc49c2461d010f7e066e6a2d398c2da015099d5dcba67b65bc238e69ce76b21609ba33d644702bd
z711264de619b3dfc7fb7ac2dc679df24d82ff2c5725d15bda782a9c78b4d834630a864c6a9939a
zbbffc316f820ca33c225120fc8eb3c9d925bbe9b819293aff0a117e8a0c2137ee460e65360da4e
z0bda4e5a5f531ae05e0728138536700f413e9a36961524b7e6b57550b0c66107e5bfb98a31b411
za31dc5261a7cef8ece79eed1d4fc59dc6f29886543f2b85e5c8469a510cddb64a42afe1b2b9087
z625aaf95ded4ffbe0cb04ca5ca8fcfa3d26c1784640df8a878a1e879738fd4eedce99eca62afd6
z95c5a23a8b69c4d9afeb1a21e774f015842af34c162c4a8f1364f398e0ecb532338d417dff8b3c
z06dfeb0ead98d08235a41635d66ea0a597baaf456fd7eb750c05225a0a25a8188114f84d165325
z18fe02b10eb92acb8cd3206f1f01f55298118270e733e9b554f4188249e105553526d80b2e59f4
z78a27976aea632a427c0af0ceadae6b5f6981c926702401c67dacddba981956ca592ab1789ce1e
zcc902dcebbc02645982e8b5f16ae33c126cda1280f25c4a919786c30c4b0b15efe2cd9a69898d0
zf2f30cae9b18a59663d0624305367fb1b3f31973acbfa0c31f740aa36d9d153c080cba56308d23
z207b9322566ca80a05c012928ac083fa44b50a11fe34d421e168d065c415d8a04f493ea13baf8d
zc7d9d48c02ae6820ae04d00df215e2b5e1f17fbaa4663ea10473569d81c97731abdf0f045dde51
z91d1962d74b49b6a134ad2197885e91178ac32da3c974a380c83e26b35b97a745415f6ea6e7c36
zfaa0d78b02
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_memory_access_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
