`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bcdf89e5c5
z7abb926401d524244d2de5706f8053a718c0490e35498fdbb323e8418acdb983005bbfd4168c4c
z065114e49e569cb0b4c3be537315e2985fb5b676f19120754c6b52c2fb9bd4801fc7940f663314
zd22f70055102b16f02c09a64ebf4cbfe24309ad9e4450ecf55111c65231140a0ac900cf4b30c8c
z492ede28c89a0a28f888dd159e201be4a2ead1e1cc38300bd778e3d728623de2d88c9f2d02c85c
za17a17fe68b809286b42bafbbee1a53f68575c711a5076fd1d87c4a93e1fd6fffabcaff4cce54e
zafe0dc802b14743001c2d52ce21d046aaaf7d98aa78588f974b487c3e435df3df58736b9f1acdb
z9e729f8960fde6b334fc17000b0cab325e30efa8f9ba6833cf904b29d85ad56dce2b898c99bca9
z52350cef57f8100833215ad679d917ee4bf36ac63409be771b74f55147108edd16bff2eb4ecee3
z34e72b9016c44ee8bbac0e6203d7a3cc04a0aa4577283106d7a08a6558ec0ada312b7bda9f8da4
zebfa4d7cae98eae827a23b41db48051f54c5cd4d44b8073eb4682dbc3625f06c971afbb35f3721
zb2647c1a6f8d04b1034850d7c58138ec0254ca64030190e968fdaa45fa7258c6463bd3c63b9974
z46fe31cdc1999a94e7efe8fa66ea16ab706caad110abfc9418275071a9279c08fed7fab87c6f8a
z324d61fc005a8a503554c3e2089bb1e520025c85fba0e5b811090239cb7ba28e5270058f41db71
z975855baafd0546c3f34fd5f6c3d0f6958588c453ffc87df37358506143014afcc66eabe4b1ce3
z5b793505dd2725c05564def38a9f79ddc235cad25fd459f4ad3830ae5d25c247e71b900681a664
za48b1851525a9db1fd13ca91353edc5266f1ab4287646b0bb87d91d198d1ddb8df040add6986d0
z23ab28be9163539525eda47041b677acaa914481660d3dee525a88ccc96e82767a565267ff21c8
z019da2f68cecfc40ae8aa3eea21cace43cdb0afae80bd5553cf86eae767f43aadfb86d6a0da398
z2132d04efe4a70b5acefaf3f0d5a9fbf740cf38e3f28a6409a9b11ddedfbe9d22867fc1c6e3868
za9f68d60f01c726f24de13fbb26625627547ec6afd46fd72d498a87d99174e261a9f7be4013c5b
zb1128556c02ddfb2969845ac565efe268cac51c45d3c3a5ace024b875f240947f3d3b87c19154b
z64cc408a750a1809238f8baa1222607a3704f66e2603a93d2e19d8e4abcc79f79fd1f57ce9e901
z2a34227ee7f1ec4f68c334898388d1da688d7a2fd1d2a48dec8b3f1535b67eecdf3125c54a0bff
z92827e26ad2b26674cbce7997f4131f66f43f7765841ad5350287f83fe458bc484327b1922152c
z33cb459c9812959ad16cea3187ffa72269cf9686c1653abb5767d5c18f1ce5b5e6b9fc0c91a47e
zba5e96d7aa15ece2bb660cb22eeb8409383fdb8dffa532afe57bb8feca48637d45647222cdd92c
z88ceb156b8480d789cdd5d947b9a2addb1faeaedda5ecf1fe3c55eca6357bf7d9a93895c20c669
z45e6c3a2631a4f37d6a18f9457af6ee51049d3db81e4e81985ba5b1f974d726e4cce825e4afdc5
z8adf01d97d3c2b95963ce1589887e8f600005dbdfbc6a8db39e29d6ee7d37f55bce47604ad7def
z6e13f8ee2e0c1e08966951f4b937ec36f505e7ebac33c47b215fee11f42e54b584e8832ecf8a16
zb8d9379a53abc96f2f19e967d103f2a068398a636f827b3499c423269750de5230cffeef98711a
z4c80b892a2e3478dbbc6d0b85ba2693bd857f22ce373992dc4ccf17e2cce9768b64581172e30ed
z076f22036209a21da30810a90f592156d4d3e3c0b1fc0bd1d0a8889c35f8c77067b5c5cc49cc1a
z51213ee6b4d2386e0e85e8407e4286f95acf3c2236d6f40e4c01e60cf43c720e6aeb390bd51fca
z03ccda58fed7b8604065c43292cb8a7e1472af1060a24a2ed118926ff3519cbf9294bb7efbfad4
z7bd5ae25e5b7e5cb5b0385300cbba27194aca4aa56fc87f7cdc0e0628300dd281a6b15d4c7237a
zaeab2a433a5c3c82d847fb4d0fa64c69a79778ca37f3cffbd5e6b20efd4580a419c9c754241edb
zad547a5e8fbe8175d2bd1abd9c49bd32e7883ae6f430328bbb50a135c307879210e3555631c4e9
zf5025d1e8f25586b50eec1d490af5843d26e65f8bfcc747d67924bf4e794fba6c8d09e1936a2bd
z32c4be648c04ba6e3ffc4f51a6d583f60c9a0b314e50927c6981664c573e03a66c171d8b5ef589
zccb08f3ae375e87dc93d11dfe064264832f0858f2dd86ca8888ad7328c8e905d4ab5f377c01610
z0c482969a0fdb7c3dc034999bf9535295302c4b599e46f9df8c6e3b5ed73f06dcb4a1460cdd46f
zb591d3eafbf78fbb098c24fc7a696fbf6d9fead178baf4a744b5ac36015dca3b84a3f3a85a750d
za95a0594d7c13eee7768c5009fbfd71c3e751135076f4b6f2ad575baa25f80dd999b19653d23bf
z93e64309be22e5742c7d90fc63b1baabff292f7ffcd117a25f0eda14f144e58c7c3822faee70c0
z6bd48f8566edded5b2d06f4a27063b4b63c497dce6f9026b56fed4acb2084bfe6b54d752836fe8
zbbcd0beb6a5eaafede9acb06aefba23afa99f4231b1a5572c85e64ca522e41c0e6fbddaebbb4ca
z8fb4a3149e738587bde151e71399994ade518f23ea830a11d46be0c52da30a102d93a9654ea7cd
zd0be5e5f4a30d53ce2f833d189b5f5da299d70ca3304dca3ccbe1e3383f3010476cf32faeadc5f
zbd990608ea19ceb2162082675bccfe3f3766d76a022ea86531b6f66604eaaa03ddd696ae663927
zc6c0596f233fbfa2db5a327850d7eba15a643860f368e08b4221f327861ec5512fed23d6889ccc
za9dc9a5a82dc4d0fa1241710f2d1310c466a4c131a5467d3729abe931031144540d89f34b048c6
z2ca11d9c5bcddb5e89bd334de7395078db63c700335be67a14584ee90752ede4c622b28d384bb2
zb851ee22bb475dd690dcdb5017fcd38c7a347b851d3ded9ea21a69ff0a185a60d841047e0d356b
z70a5bf65a1f737e0e767f60828bd893e20109fdfb3d33a6a86a9b2c8999155244818f8b54c3293
zd505a8ac3b58f695325decd9cc9a336a2c57cbdb9f42666f9321674b8b4bc51dfe0c6a23bbfddc
z7ffa0b09190989526902de10f4b7a6fffa0d2059cb3aff5e59896a0cb422d899f6d8351c8dfc9c
zbd6f07b070c3d5ae2cd7921c8474f253dce23f83adcd634865f859c28b9f8a88f82e4086012124
z2ab095d9325e24154a8d0de78f1b8c6ea19a66f13dbfb588c668b9df164c52a20f095dfb152ef9
za0fff1481cd708710ee989c2ac3b534d7bc21aec73904ab448d88d2e9ca1f32aca8ad9c00f8706
zfdf007835a24f381d5193ef59ad73d587a8caaaf1f0af799cb40796940c27522e0a5f5ba9903e6
zf2ba320005e365f5de2a6b7b07e220ae6bfec175127e1e3743869fc291699ee91622783e6b7a24
zcdc0b993e5c0b7bfff1a5160c32e4e05358a088331b7204acb55f2988adea15245e37a0f9ab8dc
zf13fabfa947f94a4d3a8b2c02a2c0bb4e314eb882cd001f038e695af038a29d1e76885db570eb0
zae4056077786703f13664589863140fbe3956ba6d4f7e1e8e2b71e620cfe26232a18f7c1aee603
z5bb015b874d9d441428c007f786b7a7f080f09a355683d7c4750a27854d5517bbe68d8416949de
zc67ccaf080db23408c1a24467b44210312faae3c407a913d2667ba50c6ccb4c9ad4b115fdf4a3a
z31fc138b4b9124107d6661bc7890d26fcb2244ebcb56a80b74e720cc27776f4ffa03466cce0971
zd11a7f4a49330906c273b5822e29203e6d01121c2b9da913e02c73b6e0341ddf7f25c408901ce6
z2d47a4aadc772a555f18d71758f291e5b485e971f2dd927837464ce13edd865bcd9794a4cde48f
zb94cb54cbe40ff506d7788c3aec03bba9f2cd5b9f1049ef7331bfd89391ccebc5dba99c0241df2
z1d7bee1f82eed4a97d0bb8f3129b25b9ed45c44f6fd160ec41d5431b720d61e6333d0a990dbe73
zd1bca91b802780c458c03f0907d85a63393439455fd9f4a66b11094be8e9caa90f6107a1a46247
zdb365d1733cabca3577df685d58777bf9647699ab66f837fee74a2e96032359c3b7635d464f682
zb4e9767f9b91e2ed5ce3c982d4eb06d223442a7260a8cf9af91a521581d262a3a965a8e71ffc23
z9aec650b30d13a6449dcc9877798ede3a7b298aa8183b7a2c8f3bad23c706e2ef44a43825d80d8
z8631b73ae6537ad7b0181e545860d32c405eb71f3017381f4dee13aae4addd786b7f509e3f4b2d
zf56471bde78119ca9b033410dd07ba8f1f39079367565418d6ecca30cd10001fe0d7c48960fcca
z78820e33a21ed344a001345859edc40594f2884068fb4f82d184ccd8e0266dca5136904c89cb37
zd4dacfefdc62fd9ad090247b7705de46154dfef4fd39a9a1d50a8c3db575538508a89d3cc061f0
z40960b647142a8dfb353a83fc4bc979efd730709e3e4b11dccafae705c78561e5c072a8d22b06a
z04505cc31fb889ce8ed0ce75cfca915f148aad9d6962348e065ad31d31b60397b2c0beecfd5b7a
z0d139a44504f5126b6ec075b9f25a8182abf8ca478d5c48291ee9ed3e7a756cd1c94a3e08cbe58
zcaad96f682614add638e95b04d928bcf905d9a7f3afe1bb3dca6dd2970db7b6dedded849661966
zda061e09a5b34410a7db1de65673c1bb8aeddd3db08f9e418331a6501e8fe70d66f14faf42a71d
z8c1b6c40930f775b80587e185d98b46f3b502a39345cf8078f74a380c246ac5428bfe3039322ff
z960ac2caefd1847249f1b00ec2e9959b2f152c1e8e7ce820b03f86ae09131fc65959109bbf7750
zb29ebf5368d0a2e7cf8ce91d4ceec5e0673871d2088fa8afa6b5e3c10a1c31d7b3037a386dbcf8
zcdb6274e5be6bcc93b29813e42ed57e1fb75a4cdbca09b229be03d0bf4859d4915058845718a1c
zbbd3fccd4768abb232e9744de4e1091b529c6efcfa5cd48ce2a8fd78833ba3ef853add6db30ee3
z21bda60b7e6b6d69a82fc8d911d4caf03b7dfd3eb1ef2b7bc09834cc993697c0c14274d149d284
zb4d113110ee8177d1147efee993391e332a7b4e7657ea9f1a314e8d30ac5dc056155c2dc01686c
z9bc5ca72ae54093703ade3b19d1e33693c1f2516afed3adc9f75175e031c24079da8caff8d81a7
zf3278cab8ce67ecf138174dc39b80901c6f82ea6112f7185f08cc1e8661ca518853d1714fd9977
z5afc485cc6ee3858f1789c03d6b4268e0f378590cbbd50f1c124078097530b1e35414049292a5a
z045580b5c6694e45279ea64a008a88bd50f7d98b465b5577e8821a41554c1090ed59afcce3cecc
zbc83c66ce1e9bdea887586fe9dead21c04d40b034268e5aecce5b7979a62952a65834555ac7a26
z5c4f42422028295eceae139783fb8f94c06e5d5db53a788c638035350a31a8e81356c9704f9a71
z0d35db4fb7a670aabc37354d0d35fd0a06bd97f39fedaf2760e55c6f5c52bc1608d44c0dbdab04
za336e8ba06bb56a84b55a0633b7d1db9d9ca31054c7c0c0ed9505afa6f751e80c0f32982b0dbda
z819425c2271759407d94200cd91e107305c84182087d3536227a0e48f3904087090d54dad9aae4
z4e818990de904b5e5506bda5d06344981f75ff6550c4c2a5c41b95eb9a7a64254d0d9ae75702dd
z58076130abf2ce4aa8d3c54fc3f84d74c5968dd4dfe5ab3fb59adde54b327bc4ae591fd498afe4
z89634285bb11c088e76ca5b885421ecf4a0a3ea4b3a18d4636a3a45fb082999117a485285ba515
za237b3b02e28f86b0aef39072df79de44dcb7cac882a0e618268253279a32f5a108de60ac6a5e8
z613b415c32ef19a18c9ec8d967d2e98d33b44ca8d5250fbc9802b646736db49a20416dfd752695
z21d2527adb3de92d0a57b94c1b9f039c47996ce6f1f98a95ff18f1636f35089a729aa5bc502ff2
z3c88340086d19a53ec160421f45dfb20643a18c9ed332a6c9c97bbca2b57c5da6b599b75bece73
zf53773803454e7feb68e8d20a1cf4f722c6053ca9711ec88c2c7947d2b5c1cee17b993a4500fb1
zd3f878a5fc80cd33b03daf766104d1c3d5b1fd0082c14a4ecf61862380bbbc5d07a1530e4382c0
z90d627492ce31636b215c95a2cb07f941ce2df9cad5afe47946d6f342770e1a5b484aa50c17a8a
z230bab546c0219729d656755f3dba27d71083d68661fc8e41ad1e68ad9385c6dead11a7ad4a7fc
z4377e7b04a2991681f9e8623f3c2a3feb41766a92f5bc03edc74a937ce1558ca4c7b6b71881159
z4b1310076b32129098e3f79c81c319a9b0671d4e6633f8bc690a69473e1bb4157409e88a13b980
z1a5ed5e6c09b7692725759025d03df8e9a0a547beafaf03d96ab17a82006e3edb500f559d60eaa
zb0d436be31ac06c28726bf150dfc60332ebbffc50ae047e2c1fb9499b70c8edf3df1a27181c9e6
zf24b33cb56b00c89b74820585a7e6a5c510afa1a59b6ade25a7112a4bc971797c1923eb429260a
zf3becb3ae800dddc77d1205eae5cc6c2944e706fd664878b6117e69eefc3088768bd48c886be7f
z979c5bb48171232122641f7e808676c5a56fabc1820fab3bcc82391972afda6859751ae3c06c75
zfdf9ac7e9aa3d49010c5ab7b0571854ea96eeb9bfc4d6a18fc1ff48b91318e45b59ba60b27b9db
z48aeb87bb120bd4356f15fcc4c941c46c9fe222a63f35da5a30a56d7a06bc9680247f73b1ec5ac
ze56da788666e30d64f8b958d80d370096a534f936b4132d851697cde95398a5b4ad0f99422d7f3
zecd7ba78857d739b77e5704ac00b0d975eb01afbd2ccdf649dd68d15563aa054b8ca79159af5fe
z7b1e8e1b70660c4827b860479c1b9534d9441677f7ebb89d823b934ced6fa7056b490806d81e60
zee20a91ad53bd7574956d70bba9444d57da4b3842fd251cd5895f53750b2c9fa7b8cc9c38cb0b3
ze3383d89286c29f93d70fea23081bb3375401a1d377ffa8c47796f02e425597059c8d29bc71fd4
z2a64d30f03c281bea659947c0ccc345ba6f2eef037ce422db0d723e44446df068ec200a1d4ea6b
zcb0462c26c3f133c49ebe08382ddb47536e18265fe92ba8805e48fe4913e01cb1ee4f24bc79488
zdf0b3833c8e5d1b27b933f37d89d0fd274847955aeed9cd8b8a31b7f08f2c93d85198e90bb4a44
z0c9e5eb49b60c6f059e6ca8eea66dc3de2033183521d4c78caf61d5458576803a68ab4dbcab4a8
z78b1d244d2dd988e6bf87dc72b02a8c4810ab4bc9e0903910e00a30dcbd3f4030d9028d899aaa8
za9ec7c1e79e29c5de559d96f897122ae76b51c3b4a77017adf2047c5f74cd4e723122ca8222cd3
zf5cd6c51cdf1a4620e3d728273260877c3c26fdd4a68161f0243569a2d53c104c4493106908a17
z0a45bf3b2b671fb8570ef81f373600dd681f8cd95b5c82e398c71b28145d152413b83b93fa2c70
z507508659a79bb097be31fbcce5c7aaa856a54b5e18fe43755195c6a614a3c6f83feb476068577
z468165d3f1e9c25849a491a3808a2ed2249f55e6d688a504d5b352eb3ef920dd65fd3fe412f9dc
z242757993d29079ce14a6a8f70d83111735b45c624c86ad3bce874a570f9f1e263798d9db51d27
zb09cece99bc9cbce044deff0544f2733053cb8645ad71c989eac7be2548dec8b969fb6228b168f
z8fac9e53e75aad5301317e4787e061c0ff715bbddc70d08906042dcc4dc85ebe5a97e13797c86b
z625fd669bfe3ec0cb0dbbcf46d015657b9894549e06ba6805a1dc328db6e71d7b2832b8d52ff30
z7e7d5c2a4afd119a9286160d8aba183cd9b0cb55692f82b12a6cd6e1ef1aa9c5542bc05bc2df65
z90268842cf7eb872ee43ea19be6b1524ce8237934de49356fb0797eb72e420d6ede58a3904afcd
z88db804cbf6e83abad5f0d59d998d919b0671724d551e0bd289b69beede00a2517732e7416c7ed
z37b0120fd00b17f11a179a5af83f3a774c1f0fc96835a7f4baa868cef5245512cedf7417ddf2ff
z3bfe294ef555ff2a79d12ee411af7d0c623395a21ac93cc0ee6bd5ce1096d3a838304578f64e46
zc253969bc7531c6aea01617b81f5291e1d44f7469ade8f22a78a0582196267e4dc9d20777c03b8
zc8aa12b0888c35bdfe23b50b66f7c6ed3332a92094f28debabb67066b0a7833ed0a76c08665348
z718c910767d97ac0145cb4d10db48de0dcf53acbc93dc77fa2ace07178e8b980625bbd2af47396
zaa66315a7aaba7c9d052140101cf5c90fe44939e7aca54c56e6d8d12e412516611bef31e3bf4a1
z522247dd59827979657e16a6e0746fcbd91ed21b286e8b2e58b0878b12ff2b6f174fca9368eab6
z99a83df7a6504ee02e49834821871d3d6fdcf4bc1996eb522399d2d6e5b3bcb9c5dcdeaaae5f7f
zed2f22d19d45a5080869a8cc19ce98092d830bbe534683880a0232c805bcf8b7628f8e1e41094b
z5be4a6b85848836dbbf44828e1a7abcdcc957da0aeabb660f293101792f005e2c6b253f370f49c
z03c4bccf7f0ac46d8ed616a8d57d1ef4f481137266c4e6294040fc8b18ec0c84175f75b0a9a367
za3aff589ea281e38691b672fd621b2a0967953d3cf7d0ee8cb1efb227fca9324407548518ebb1f
z5bf536f91a43db829ed65f9334eb85810ef635d5a66099237ce36026e55917705dee1533acd30e
zaa63b8dbc36cf2587e90e7f93c86f50240178d64d3d18a191061fb340d6c38d133db9bf77728a0
z9fccda2ceb93c383948fe4ba746ce748060bcb28f6a4e19d84db81442b3286182281f9917ff494
za37ce411b803cd3e8987334a99efb3a17e047d081f88ed8380310d0487464bb4b23b6ddc427d69
zedae0adc56d808007f2ac42ccf2be259e6f3bcb5b8cba5ccbc28c6b5aa9f3bca10bbd7275e7dac
zdb1e72bcd3cd116809014f8483e3cb1e8e8f8c60d218e31dce78af7f2bead5f70a8f6bad40841c
z766fbd1916a6ca2d45b3c62668a0341a60b6c7075b90709c6360392a4cfb812a0f4e217d6b25e3
z67512e1d2e6f934a8c34e19fab7b5e2bc3172fb049fd5640ffe0932cde16d609968681cc5c427a
z2bbe80f699d95a96b972d5d2fef5cb8f7c8f675cb7c1e0fcfa13b9e39d9572fd5aa7a9077de9e3
z257f1618cc195f53c18544b82a49ee41504eda4fc942f2f91cd1cc12a188a5a01b402a2c78711c
za46248bdcf016e82e16a71765cf5166905b52371c3283219dd7af8576242facb5d1ed45e1f89d0
z2525191cbdd79584a166966db890d4b5890257f30f448dc6c1958722ea3977e1d2df9a7e0d99c8
z37b4f28800ca31916854a4748993930ed0451e8f69689a4cc2187a661a567a2fa742cd92036ae3
z182d9fc8aca6a8e6087d2444c536534d6dd2980e9a77bb57409b9e3fbe73e9a492de97e4bc4cc2
z96e9dfddccf751cd5d24dfbf7ab694b959d0481ce95e034a10e25eefbda0b328385919008cefae
z9da5eb8e7ec358bc9eb909a340d4631c8e62015ea7c4af8f4f911bec9425e4c5c5eee9b4f9d724
zae1176652492f27177971b488db5e811c885f14a044ed59e253be943187761b71221ea51aec65f
zc5c5a36ccdee144add0003dfdbe237d27dc3abc692d6a8bba1902111cecee8bae824691c1f6f9b
zc84a961afdcb252d2786bff1ba9bbf7574a29afc171044d91e925bb83baf45bcc2b805191beb44
zf55eb2aa6fbd279392f38ef98455dd9f5d9e8d8afee4aeffdb2783945f221ec3418a78cba08073
z2b2431785382f46f1023f68c03c61368a62a51dd3d39439ad7837a183fc170cf6ab40538f98f67
z000bdfb8efcad6e38784bc5f1a9fbf6e0242bdae2a9a0f13e3166b9569196c8c3714acab2fab36
z950e868085cdd1329be215c3325c16c62a4182aa95f23b528bcc185cab22563a1377b80eb2e30d
z429fab6d131159857529eb49b7d88cc777216ff6529a717e4d0ec06ebce2ba7eef6af8edd240d9
za8fb77bfcb1784ca4a97e8f2f0185f32be6436747f5980131e5c97c8107e0dfff3159411c82927
z6f68581f1c9f48f84ec16aa94aed199957f93d8a1eb8ac7a83da1b35e7bdf8dc7d9c7e39822167
zc713ffc137abb03610163f1465ea22e19d122d0c1b2046e5c6cf84ce2637bda4234a93e58e013d
z47e1d47fb17af8c73c9279fe19e4745072d5704ffdc49bb2cb180843e1f3b4077b6ca95fff9cc3
ze9822e4194efbfd164e67c16e1eeddc0f49a5ed96b09a76e1bc87f0e05478bf381b649496959c5
z64ebe4e9d3ae19f4f1e52707d2288e26458c583c5eae5adcf539f27f281b8802c13619084cde56
z2e9da7ca06bcb28bc011e6fe5848c1a4eceedb53be5443910ad2dc14a8a02d6d3ce0c3627e2cf3
z2d661ef9584737485aedcef9b74343532f949275ab422dcb9867308a36940968ea0bf58dccc9eb
z748224e3edb8e6697814150b7dba10d13304cb8c203aeb7797624b054258b0bf1e2231b3db2f70
z812fd19d017ca835f354243997abf2af0b4752ad1270cfacd6cb01c838e00471a77249b0c3b82b
zeacf36f8aba843c1f49ca6c4240114a166f3d23e28bace18c8e0c569ae92aa57cb078f13fec982
z2628bd2bb6f55caed58bec0dfde7645c2d7eb7dd6734880b10aa830e82a752008306ab38ccf881
z358bcbba1e181de5f73c2cb2b2303abd2d0ccefbaea7ab52afaa5dfa9f82261b65e4e2221da599
ze192181ca245ce7705a8d4ff0fba6fdbce1a46f79ba28e440a850a48a3131ce43a51edf3a38575
zfae196c9595a9717bc46b3716435ef479d3a9ef8559ab2f4eeee23b86c517ddf6e84e89d2e1f5d
z1e6066ddd387f6c40e711b1e3af4a9f9a1ed346bb3f970ad850a2baf5e2646ac5ee64fd8019155
z0128a6173e2f17814e0bc8d4902c1e49c2a66e10a00945c76e37719d3deec32690830ee89eae43
zc50eb479d9c1286a09e976a59b5bbeba6873624074eaf409e3093ccba1af8fb85985245810b575
zc3c879a5c2296836a48736730d3013257e0b9f931405c0d9376e1cb9ff1215d4a71f5767e59eac
zcf105966c4f90d438ffafe17f75ce3587857de6022131e491167b74df36bb9851a8a7ae2431dd9
z01a5d1c58e8e2457a3c55a35111c770eec0a0ca54731c3bed03e8286c24e5f77b52e2d955b5ba9
z44de4874b57ecaa206ee6d75009d539fd2a4e8aa24b441a947c4d696f0da4ade873b08cf50b07c
z0cb1c40803edb8e213864eb09422c96af618bb444945e8789616c7e8aad47317c626a6f2f285ca
z2f4cb3b38730c9eb1047b54cc77d2c1e705a41d38a74bac77a66b22ee5c5201787075323631ebf
z64d34ba6be9495ea0674deebd481121140d6c72a94c6f89f05ec0c5355c338af1c82d97f54925a
za3bc180752ef381d4e4f668a2965b8c56ef77073f12def6e906168012b691693c164777bfcc1f9
z613a33c77925a6595f2971f982c00a69e25575e8309dc6b64e790cd257394c7c82508b0ed22e5f
z37ba15cd51f356ea7d28155676f440a1085a751fb9747c712d20e9c55c6cecb40e910a7778c93c
zfc6af6dd96574d1dd9db0effd42cffe6fba5b16ba77d003e74e7d2890e307c5fcc763418685d8a
z7950bd6e74b5136426fa99a2bf42799669cf1998bf2b46c8493ea70bf6a33f3ee18e7242afea8a
z0bfe906268dbeb9db46863899e4f2af1fefdb1258fad34ee814bb4206effcf2f19c9a8f1d6ccc2
z504362955c774526d0c20f6a0c930c7e1ae7b8ac6b0121555ae5e63ff2c2e6e2346dd6bab2da53
z31732fca769063a73c9b4c7cb0399acebb919940dbd19f8cac9785d80c06c188862191b3b6f6c9
zdb8fb84a94973909fe2df78c505cb127fb1a40e509585453dd5d372086bdd1425e3c78b263a2f0
z444d9e48e3f257a44deda1b69142272a3f41102d23fbc0f7df8a89e35d1aea638a54b70b7f7a33
z9ccdbfe3a6bfbf9c3bf5711ce8c31608ba22e89de13b586774534a163d0275360947dfd0f110bb
zf0a1caccfb6a01ad669f07a2e95cab33f550972a63acd52ec2b036ff081be972f13b5b2cfc003a
z7ee0ff4f926970ecdc0044d55ce4387937714013ebd7e7cb681091c6574a8e5fa02ef555e555ae
zf5b833cec0b15253902356b38ca7b965af24fe6f82c08e74b23bccfdf0f13d7100b0f75bf3147f
z336333e92d216e8a8cce2b50276d6db190677867ea6e9fcae7540629ffa9a96dec4a1906b5de3b
z6306e577fba40674d9d5b69879c5c0b979269654863bc236843c6de0237ee57063bb20884ef9a3
zf3bf813e828a29722798055dcb06f797b8458016753320a919cced32f5b0f40bf72bb1376009e4
z2a9a1c3a7113b4413f92aa286b77d0e82223b63347509b812c8f40d05941c69062244008694697
z09cc6511cd3a07888940a71b51f7865f695d2abf9e796a4761b825bc0c072c45700e96b444b35a
z1305158a5082223f409965415888618162e96777cfe914de229f7370aa595026a70b577635b409
zcdd32cba3aefe124d6493a31c2db81bbc48a7b802319a3c7fa5cd8810c8514b37f61d53fc47991
z9d407b815184271cd8297a133a9ad20638313494f5b0680782b13bc2321117d9191cc6aee1a9cd
zf46c5d002fa7fe2824b096f2d64174bd51c15826b6f3102dc739399162f39fc5b592fef8e3d734
zf1ddc7ca4cc9830fbbb2b7c70e17b70ecf7091ea972991c64d7f6ca92f1d6a81afc43021a9cf55
zcf793b89866db19f2999d22644bdd3270680477440ae11891b459249b2871fe83f2bbf4130214a
zb14cebcd27d6fbc700e866cdd37ea22d33e22c828ea17f4315f6cd9bf6f60cb794d7a8ac4859b8
z985995962a5442c38bf6f005efd8065210e13fa0e56f5bc049fcd490db2aead0fa10ba144cad84
z27ba0946eeb929267fa3a1c34353127131d890420f217956548a40bb9f957e6211c920938379cf
z9112eb9143733705e936dc08263d965fcdff8310511319367775940106cb4dac651f42e3c454c2
z88d11a36c70fa5742bad9883ebc37857e04d54151f7fb282c3fa4bdeafd374f07ede14e83cefc0
z0c571c664a22555c7eeefad7b5d5244b4028f9b2f41e538c7fd28591d007e5eb3caca6983a416e
zf561ab38a96a015605b85f80e0026ec836b6ea9da73a4c444d6625d444d330ffebefb330225836
za63c44fe9049228ba889509c2fd542200e1027fe5023db700fa820e5af870912b22131a1518e3e
z16118ea580eea59d3695a4ac3e8326c7ed3293aef72466fc6ee9a3d8f98d3dac932eeb0ec52200
zfbd135980db95fdbe0263d9bd037804f22ffd805ee4e15a326537ddd4b4c289335827ce71c4f70
zbc5b371bfdb897b0a5ced2a345452690e8abb89b166346aaab5dff2a01a051101f29d9ef79f649
z87d7ef4d52e2005e4ffa38460f5131645b61c627016834b9cef57949df077ac1731f45d94fd9d3
z27784477ef62fcb3f7dc93b782eb41d33aeed6a39f4114a4bf6d14ff9043403b01c10389f7cf26
zd52c404acdfcb1f1d1b56376715ed4bcb0d2a78f099671fbb0fe31611e28a0cc4be3db70ff21f1
z72e17a191b93c42386772f5a1c25102c341f5197fd7d34233452c1233e2867b8e94228b39dd378
z0ac48769a08a8b406cbac82f0edc61a19cca35fb35b274a34e8a3d026a583648d4dc444b39ee52
z123f521e4918964fa1a76905b75543d162b8b16232fd0a55147310f63702b98ca23e1ea8b4b443
za898e8fd300fa60ee4f06a8c5a5335424497eef4c30580fb28213ec73cb23f19887922591f8537
z238c3b58fe0a6ca761280ba03beb9515b20794f3e1caf54378dc10d84975efd0612f1019fa1fcb
z581dc815eca9fe706e83ab609e5a3ea361700d80a35cd0418a07e8f75b4f6bcfc12f212d7d86c0
z7247afdda859c55d61040bcafdf9bd0dd86db50731b5bf5debe2a7eca2f959e48846a06634caf8
zd5cfffdd4c3b8a0b6b1dce28bd784f7f2dd87eb497e060660e6afc3adc5cafb46aa47086a70a20
zf909dc8c156d04c8eb73592a0a385c8889f5073522cfb40228649d7d1325fb506737ed8b045e94
z3bafd5b929356924e9efa9a87a6f5050a775f1188a3a947f110e17afbd855ac2067d3feb7d48cd
z6dceb6d5d01cc9bc746027fec8b6e7335a6b8f9b019e631583c9e76d74830e276ae636019aef5b
z8ecae320b85aa504e962cb94eab7a9d0e84e8a8960aa97051cd972327839cb72d39e56769e4403
z1dd116936c4e138706e6591f8f3a33a3937501304df914b709776ffef73405a5439da92c0d161c
z7eb26bf9e7a69d424fb53b36b49b72ab7d001f1564d51d04fe0fdcc021e00f7cb0d51e623a7ff9
z8d300255a298bbebc67a31053c9a1cd144cd669d361687e49f85400d8c567cc05bb5381d89ca50
z2d770efe4c7cfc70448af92ee9fdc3b85cfeb20a5076df829dfe683b2e8dbd5b52b661c5cb4279
z75c6d5d57f3817f3fc562da237fb0d1c710ecb1539a98e5f84127eeff8e814a9d0232126c5d4a2
z5b8fa60d9c167867868a82975a2f8268b05b9e7f6d00811d8cba173d39f10a2053f21e27fa827b
z94c4aebaa45a3f0f39ba22f84ea6d7e6fc3719f75d2c0fc99b7aa828ea5ce46ad7661b40166c5d
z4f1f2694fa2180daa35976e2fb7522ae354ecf9823fc43e207df36192bb6b7ac3b9191714f2632
z4db1bfef5d087afc0963b50d5b10361e83eb6f2c740b8939022b76fa51fac3ea591edf871b5501
zea8fa583203433790524131df5a21224e6ea4f31167c9b4c1c78aafce9280501d9e0dbd866ab84
z690ee3475f7a5951bfcae75a33d9b88aa1b9b9908ffee2d0e96c4ff8bb9a531c8a6658bfcc3798
z16986e5a666496691e564eb25477e09b79452cb8627902e473f7e4a5a028b591908a835d5b5547
ze5dd168be14ffba7624654dcfc9ea16697103e64ac45eb7ef9b72af2be02ead54bb91696646fd8
z0f25ef7b1a2fe25bdfd2b3c72e97789539c70b5914b6b9ee0829763c6794cbccd1ea96e425d5fa
z90c10281647eb2075b9a2d8426305cb918f277a58a860b2bae2f5e24ab2714d5e832928af77f97
z47a6a874209509223432bf7d31cd1ef7bbc7233e8a0eae011565e596a72d67b0d74291c80a5dd2
zfa8b56025f658f1616ae3fcbc28e2e2aef3b5e234ffa4fe67ba05d26e99cd598064e7091518345
zdc7c19a2c184cbe74893faef412eb6cb89db2efb2b8a1cd8524df2a2c08f612f4c7d89981a7447
zce556000b01b36eca09f64cfea3c2681a91f27d3c4221e338d1d2baa1e0898862deea2e96242c6
z4fc7e9fb7ea5561111a856e984ec00bafe6402a24f9fc80507c656522fffbb8a8a7aa270fa4aef
zef0840de69e66b625400674248a4d09f98e72728caa390efb7ffb03f292c5471e996c47a78c70e
zcc140e5d7f9cff2c1d9c2b0d7e2816333091e2a65f13aa94ad00eb573a8180f775c047c332dbf8
za042a57fa60350fef314488a635d1b11e85fb7b6bdcff9661d2e396e6394ddcd9d220f513e6726
z4562413f3389d432f2f2f025f4117a57b71f1b65694bae655532abef83f9cc0ad021f646be8396
z42ff0860158a99313450080cac28465f6b71f4059efef9ea1d9046789b10134344761a9f3d72dd
z2c4d141c6041aad201aa9a210f0e799c16d05422fc0ade998bd6d65115703060c46d297b5f69ed
zbe636df741b7a184f80dd419b24c0adc6b7eee60e2af41685b9c8db6a5187d8580b9097c9e10a9
z2652c67e0836c97f3499ac980cea17e63f3ca6df8449bafc48c4dfac812380efe1d0d7e2166ece
z789e810bc4f53f23619c9619e6576ef2314fc647e402342c379e92b70273eef70781bf8c7d04b9
z046bccb0171118da5bf0669a46500bfcdbdacf39edff65880776865331ca1b56785bd0f943c6a7
z957e7cc695714e82098a9debea73a1445b95f935b8714c480122eebdbc9f826340bbc94065d485
z3d7ed76db722cfdd0b97fa1f6d01541391f0a135731687d81f9f7a6ebf199c44eaafc2d23eabd9
z42b8402c5c3d8c2fee71f0d783fac8782b81952cdedba4c23e5b25769a1d39185612459a86b42f
z70c4ca16a3d0caa4728a7c4ff06e4cd3ef8dd4f160baf1f532e21222fd299394ad4ea4bc281300
zcc5f2754b094f2ab4e3e5c311abde66c54893855398a267e19ec475cca94102d8047095c7ea0cf
zf6bbf8df2163a289daf404d56a35c1bbc2d3b6fd1e3981d441ffeb6073a5f1ef8777963f9facb8
zdeef7984f8ed4410e558567452d397371abf3dcf3e9c70f8c3f4a4d130051a3d6a9b2be02be040
z8c93d68fcc818fc55af30933f5cc6a91ea6ea7405ab31a6a7d3799e8374601b664f9bfdba270d8
ze3452ab7383298476923ba32a3a5b59b79fbf79668f3967596becce379477d4e9a971738397bf2
z4703c47e8466bd4b06e224f1a41e065d3f791229eafc960ddd1f8e1004672a256b2970ec99b2eb
z4053a50409eafc1ce977d111863a96fa5a5f1b82cae891faa09fa0cdd64b7dc4cf95a1e9fd9860
zc158b786ea96f04253b3802b26c5d28bb2c78fa205572167d69341cca183aa358bafb51d53bd05
zd79178561c5028549253c7a34551b21131065e5e2eff5267773fb06db5fc693c1359ec28cd53cb
z071ce4cec6f4935581420e7d6711d7d9253d4dbc14acf396f9556e470d6d07161f3fddead99f8f
z1accabc0cebbf9f67e8a33b47e4adcb49608ca974a05f82437300a7b242adf0eece4d31ab56090
za05084ebe9582ef94eb76009ae7c4b56308f6e1559562cbf2afc1e374276008e426cd0714f26bb
z802e8c7ee0442da879ebfa4be9ecfe00950784c2ced4ff5d98539a1cd35a45eee0ee10ab92fdf9
z13a6d6611670f821188d9a39b9478272f818b7e66e66db83b358e976ede0aff0f34797683e65ff
z07f3f4be1d1e8b350b71cede0cfff308da24766cab24c692d86f0c08c41f2efcb133ec6a3481fe
z993eacc9814a7d42646ac3fbfcdb4c677495cdbedb1f57a714fcdf0f7ba0f8ccb12a8b14a73729
z4b1b0840003f3193cf24ae6dd4d823d77ba1f54ddd0876ecd449e20c874ece17e8b6d3bc4f8c95
zb26f9f6455046e05493bb7efde7a3491ae26f373f1d92c51143dd1a947ed46926168fc263b0cd5
zfcde912a27393765c3ddbdd2eb36b832bd175aaa1f8d3986fcb6443a966f1a315be165b94381c2
zaec347afb32db90436be6bb074a2b356a9d93560f736f651f2b6cf1be8bcd07034ba79c52f3d5b
z43676df34e9d81773c0fba32ab037467d68576c4370c86e98ea4fc3813b1cb2fed0562fe51881b
z5317774a9d2659b310bf959fc36488547d8651624c67e9ffed0a94d261b71032ae915ea6cacece
zbe361a6f4ca0a192445f2d3557071828fed91b20c6f47e08d1e6b3ee96b1ffca6671223d62cee7
z242fe87c76c5678ae4de455394736cf22089d9414b48e5b4999e96d12044905698b0d0c0c502e9
zc62e7acfaccfa0e9e506228423b6b054066933db312ce181665d8ac8da5f9d57ceb5ffbdf1253a
z2dc09a61df41f8d45a2d7e94bbe990908d922743e87014c3bfb3b4ce0766c3d6938badf48a2421
zbd6b61c18aff5093549981face31592e834992280f36c0a08d04c9a7c4df26a638187871ff139a
zbe7ee26b739df73311ef9df7719d17f72f8f43db0832c09b478fe87e21d9d8408aa073a0ab483c
z7d1a84206fc668770d53f39275330243d12f33061050cac6afcea773b98b9b18b6959c00019b9b
zd798e6c16767747f218a36172b93f2608fe9018fcd0e1f9a6aab87bdff9f38034dcb2acda72fb8
z49de1a7906bda1bbf6cdf40bfad7fb39bdeb94889beff9dd2cca4f60ffdaecd0c617411a0f7306
z591bd2e83f5e2d706aad46ed1368101a0ddb974b2b764f6551f2bdb30c374b94ebc56d3659c4c7
z52c91418fba98fca835d674fb1f555c0f4dcbe0c98c94ce7e00ba866a3ecde381aa050fa3cff6d
z33dfa2db17295601c269815cbb2a25e3a045a3fac27cd70092232ac207849796e1a482c23f4297
zf8a8d77251874f7b2a009ed0f62cf419b92ece7323210b96e82d7cda8c9ba33d327e4cf07c12dd
zeb8330cdc3b81f3c78e9a9a262108e22c976229e06258146a090160b6e830308546601a54a6dd4
z044a19281e7b62a901113e1f7bf18a7abea64cbf607a6ccfdaed83e8f42b953f3ba3371c1d54df
z87ca9d3a90b5542d2ad24d050c19b3cab6ada3e7a25fd4b08c6d35603f91f87f6b527c4ec5f5b4
z72b854454d231c0fa24b7bc9dac5cfbef7a9b8af32ee2cb4701e6abcbd088e016c3714fcfbdd7b
z6bd701f7dc2aec89f8abfafd1875f537ec2ea005fb396551b41e2328f4f6c20f63ace1e313a960
z4a00cbd09f1bf02e130c2d5a1f070656cf035df049b8562b91d32263d5c289322e7ac6ceb9b46b
zff70b94717c7e9db732f07c78833d6304ba35aa91784a33ce0edd00aaadae2eee4003845df27a9
zbc922a3ceb56f184cf52750691a442acf22d3e976a0d2f33b363f6cbc78a9a71379c028d1a28a5
z757e1079ca7ea3b9d3d47ae0166446be632f1d94d825af3714152421c5418777a92c1fc87f69f9
zf0aad1444ee460b2b8a7189347ebab0a0b244f0e435c4f15ac51e4aa770ffcaf23a80de3d44ed2
z204a4191981d32da4f116db0a6532acf4e6c93339540db36e2fc1834cba52cdace08aa71873d0e
z424e969aa0a2c771628e0b0867a4b8f70b037f17047d2c0f3400261b03f0a367d7c08268277714
zd2789255276630c792f6f1ce2d3b74f1928aba2acb0ff5eb3833691195cc84e129ef458de74330
z285e5a95489a0205ccd9c48362b0549460ce793e1b0585f2078c05ac3f2fc5e97bbaea2231922e
z9b54c48de3a72019339d5064f5e5f5676e901369ee6c1b5d132167cd75ad4159b4fcb0ad62a73a
z750d781ceda2ef79ba0343be4f3b2be4c8d14c1ca7b9d8c0829cedeb3a26a86eff6925e1aa4c8a
z402d3e16d7152aaeb39e4a9a1e818f0e70aa84404e7b8f6daa6b2a7a4e7d1f01e2bd0c1db16b79
z38f42fdb5e420297985de1678e6e4aa0f24dcd102cfba7ee768ef9087abf51a9a9484dee6aee6b
z1f8bdc6ae05c17824a908d5543b5666841ae8b0c6ab01f0fdd158e67b2196f89ac1c96b8ad4bc5
z870afdf1dde77f1e9015659d8f054ecebf0adbdfd5dc09778f6cc9d04de219eb557b7e7fa6f84c
z8db4c68115041011605c9dfe91eaa96cad95e4094de44a56d396ea63f6de9e5f0d77811a412646
zc3bf12c9296ab2b7eaef3a7fc9bc9371fa33000e396c561a8ae955e58fa73ee27127fe18ada3a0
za31aff14f3e1b11e289e130d9fd6a97b762c9658e9fdff6a04832727916dcbb8beadbe73ae2b2f
za2d98b9d7d7fb22f6c38bd076ff376ca07852878b32e96f9891156852743add4db493a2e995f54
z9c94ceba9879d83906fdbb40db618ce86544c4f2dd4d957cce5edd990b423dce13dd8cbad1b9e3
z9e0bb2d7a11303064eef5a59943c867b4f4d7fcee4647dc3fa6c94eb3ad8c1c3228e253887596a
z9d95216e4bc1442d564e2d733634df288ad35a4210110dcfe5ef2200984b68718eed21f78c3189
z520a7706c864fd152e79af9004788a0fe39260c2f6ce099bdac3fd16fd5b9b4883e474e0df2845
z314de58d77a528bf2b2f4444791f549f8e0c3623088aba328e612fd57a2a16f5474b1c85bf5718
zd47a965a5e35c9d3f2d53bb137dc627873e3a81f0c8958e534134fb88e12fd55415440a1f18511
z1b87210a61b5eb481fcf843cd84fbda4fd89ee3093009817c5bae180ceee7c2e15cc9ea7c53296
zb3ad28962404c5bf72ff9e9bebd95dccdde92bfb319cac2b49ddc2e3860de4aa1d567bca42e140
z51c31a045877e7a510655ede70b68be98bc7ceace334547988d250ce00f77c17365798c3bd5270
z0c5bd7f3a0cff2ab575311adc5971e8ee8d09f57253067b6c1b92b5dcc287c397c40c1f01783ae
z656e276bd517276a6553aba8196ef7e19eb3e52703d1028f306d8cdc3ca15016ecc811a2795bfa
zdcdf9f5b4ebfbc76a7e97651c1a67a6057644df14f60af66ac0145f630cd33bb2779438851cdff
z40ca4334c1a6619781326f6fa324fe03bc3c485ce9420df9b258d583d9443d5b6b866b74946f12
zaaba6934f3b36e9384dbd65082d292f0168ee4a74e6e20cbbfe7385f7acc878e15b203dfdce4b8
zfbf3913da4e8fe4ab11969c382ebc7f4f50bb4e6a3239db9385a9efe2de212d6fdee4deadf2fab
zbb81a89b3a8f8a7900965792bfb272db7c5a46c73941c7ef5c14d2093c65cbcdfea6e9a0040caf
z91b2f9a0c9257baa10e74e81288ff23f87ab8c671d8804b26ff7ded7596dc5802b6defd9fb838a
z276048312a95ef660c3dc5c390da3c1487c08050dee2bc507f52427ba59bd92dc5949e2a040c9e
z9a6f792bb1f922af1d77eb23e63b627d4aa0123f1ad2b95b733d5e5a3f4f3df1e8cde34a5cf29f
ze86334963dfe70a3281ef5c50cba14ffc0cbb97a0a4685f50443c7fecd8daf97a44d55bdfec6c9
zbb71086becffce9e98a84a0b8c8952e6d7f3afeb0bce15cdb092fdb3354eca283983150ff3450e
z93ce33c52163fb55f64288245bf59a5646ac3960b3042141dd4a65e162cb39f5f11e7b7dcb62f7
zd593d1555f7b951539be1314e1fa2149d7b6f98d805412d330a7e98893a24e7a689ab2a4289323
ze4cdf209c9c85fd8e97ac63d726f78177d7b61957c8452c6e92d8cf47a307abb3209b388bfb683
z89ad3e1987839ef1761c8caebae22785fa55f2ac269705d4fa66ddaf90e7ccce745e39b8a483e2
zb40af42dbde7482e1c86700e7d185165d88122bca29655ded5e4b057a2bf5927557180113f9bdb
ze4436e7b9e4887e52d01a67812b2c951581089414afd5f37ff476c7c93c690ccc3914a8c38b05a
z6c3ee145e289dd39b399122b020f4ac1adfad9159d1edee2cae4d7da186cccfbb5b07b54057bd8
z30b2c4ea26c2d874284d30b97fe9d85d2a8ef9912fc6e1130ab4931f9c37630749f89b09bc6dad
z833141f17700795c5e788b079f34d1a1ae51c29c9ccdcdbaf57a5b4e42c63d1382880d040468a6
z8eb35fd21011225f22971a1a17934fd5b08d1bb779e0ab781c7a591be5351390d9bc78bad6fc4f
z0554674ba0e08c18f3a07a1198530143b9742a72d97aa65ecb40dd62f71008a0baf685169d0644
z304f555973d4497f7e0a48995b2f8d80beda65e4ff55d3bdbad32ac19faae108e7f7b0f3a8574f
z1f94711b69e21c6e130eb47ccb18154f0f88cf939c561d2da7572713229d7d6dc356e0c4c1bdee
z3152a84fbcf5a781d1ac4058238a64335ecbc2b5e874f0eb96d77b797ac75df9ce3b09f6099de0
zf38860bf867b9e2f7dc63d5107e7e7f8b815e1aa1bc1d576512dface23ea3efc595800e1e9ee2f
z93e3283f12b2a91b5842c9cf196f00b1b368fa06b5f7a3b66433ed46d4cdc51671ff86fbd87b62
zfce5867a8f9c74df48c96face73ded76491c7d9e407320bfa7b00d8359d45986aea2f33ca3c6d3
z535501a6f6ca48d08e693bb71e78f4f409c482236a7b2617ef04b12f4093ffad68e9d5be8c0c52
zc4ae81b46c286113dd85b63646a2a7b36772a570e46df193ecb92e73a265fd30b67e9275b0d7a8
ze9d0ed8201d9ab2ccd4266c574a2e6a38549cc9f77a4e8909ec9e73565f14edc2d078dd320f780
z9d878f18d89d99fbb7199014d4a92f87e7157a5e578167410f4172312ba497f5224e1ed1d500d5
ze18a53d78fdfe3a9adf1835534178524d9813d489286830f9f854ff5f0643d034f4143a8f9fa76
z1000c44ef5d2d7959e0e88e8637af42c8273cc385d51f2f0fb3940f6a9c1a2ff7b076d7863a64c
zfd114ff78e51c35a88db57315ed2c040fd76cd8a08a409a85a0224b13cedc5b76375d9a9cc8324
z1499dc89a1424962c954c8f9b196aedb35fd1cf4433c088a6a2cd4147831623a67a0bb38e9c62c
z01dd79c99549544efa34a6702d62d553c1693240de6db0c63ff5ff68e88e3f6f52f48fe31d44c2
z6b1f443757178fd5b49dca36dbbb8c2627df9cec875ba6a3098b57e04cdea7c9cdbf28dcec320a
z4e66314a8f2c9a4818d4a708309fd4a11ac3d5d30c06f55444bc638ed6ed0c12806feb93a843cc
zd000f454da0821de4f795d5aef35319d3e020a60c447a3cde10b7e30c04fd73e8be2bf18b4ad54
zfd51dd05f49c9d79ef8fbc4e63778a7f6756d923b919040bb657235764758c077914c834f519a2
zf978033f646e6ac1e4955268ee1074eedbdb0cbf5e593ee7d12b43016579f2c7e2be3e386ec1a4
z57ea406540a164890eec33abf8b68b3069bbb951068944bff255a9f5616ac62374c9b41353c994
z881d655945f616e84e3fdb797162689084361c817bc008e96db0caf24b9a0ab81327153e2cf545
z0c26e3bad4afb53c6f0b10034ef96ba547a1842412a0d8a6096788968822f63765c088869bd49f
za619f4bf1b32802372517168e9209c536e0d00ecda0a32fb5a05d70cdfe8bf9f16300cc4324565
z8b814d41c09f5149bf7881766851b73437719dc596d8a99a1c05faa3e3d588f46ff39eb80ca385
z86b17769bb986fb7d2ba606396a5d3a2208ed996288b4b019b3248e991fd6de9d621b95a9a3106
za788b80aae5241377b563d7a6a212294af743ef8d1606ed52d72a6cfc52a5d5db1c728bf6500a3
z389f0790da72acdc0d834de6fdaf18aaa3cef0f08aa92b1acf687a61e1bfe43f1604a2fcb555a7
z556bcb9d83abe5b9c4d1cc3be0d0a1779841684cf6ee0cdb54c6f1cf3866878a9f9a78ee3fe98e
zc2117fd57a785723684297ae08faab22addfc5009e0991f27966358beb4a65c982d898304fe5df
z67d3a647e51b0242d3ba49683da4b06b1dbd3fc40be796ff9a819c8815cfc29ebb2b6247a0a746
z22e699f9e85c821dffc55e4d4488b96249c90261ff5db4de017571c345c940a2c99c309b7a3c1f
z1127012d0b5d5bbaa8a2b589ffc83702dd1bc8a4f8ba3a36cdda497a2fd68dcbe060fa748fa4f7
z6b94dfe0a3ae4d13cd961645a82b5ca26620de83aa15fcbe21711195563285d42366ed10708f31
z98a3ef28cec5c840e62d8ebe457ae5227c48328f5b111d75c1b6aec8fb9c89f3b2861da0a0b81d
zeb72864421165968123a83ee36c6f024bebc4fe71b996c42069475f31835d7a02d9966221f45f4
zb6578a4033c89059bcd769a3884c64d767570a9e850f22f8f3ab64c7fea189c3528307148b978f
zc5f1e3262e9d9ec60c16e179bc8653ccbbe9b8a06d27713c4c2b0dcfc03be77b0b67f14c83228f
ze55dbd4aaafdf136a448c8d872d9b4583cb7ae4881a51e38b8f84bb24d473fe09a6d7b1f1cea09
z5e4830b55c03b43e75c5ab75f5c79cdc3aa9dd81841505b9a26c394cd8502c4dd1d3d3d69fb762
z008ca13f8ffe92f31f985ead7745204f09fb844bb984ee828a69a21a641caf6e48be4d55f4858e
zb6af0fcc304ed781643f4e2a46d76e65c39c4c6dee9010c44b1730e923610a77ba69d00dd80ae4
z6075cba480a1940c126b83dfd536bd71b1657064392d3f0111aeedb240e2596110da4d9cff3003
z606970604ac0b16a77be0be8da3f9239db31a3d20ece27a494fd6319007254053d7d520ee5be8a
z831e7e1201d9a501e5bcb5569d8172d6afd4fda1cba010b1fc85d15b29c7a740580246e22edf61
z0ea536c5725308b0fa3d56db9ead3c735b6f06b2861cce2a40c0a79121b7e79d4f1714c10fb10b
z36ab1e0febe5e873be7d306bea7e64be05ef7f6c53e151e208c92682bda363bf3c99afd67881aa
z5b90cb5bc13631f93ea34cb0f3aa3a99c79c76a2e35a625d499dd37160f927082077c5b67f92cd
z756f423bf972299eb6210d26f0c16f15bd4fbf3d1d38956e24fb098312c617c91c410ac518a035
zc91af7a05b4362612ae20b1acda69fb4bf64e836dafd1a7cdae67757453b192b4e9f216f892cd2
z798fd3d9bddb248b751f560a4fe32484cce62319ed92023288bc70956c28e9d3be175d989c67c9
zb0dc342a5fbc2d5644224a73b7f1d26f9eb1bccd65a2d748b1f04956295e0a4ea11a675e403014
z3aa8a75d009ecfad1c821ec600ae576b20dc1782e3e5ca37fab197f064838f7b788d15e84bf29f
zbed3dd3c72c931fd87f52052f0a812dbb974240216b8727f13f3608e603a2b1df1ab087d38773b
ze3132df5e676068b399387f4005dbe235d457f349abf7a8c840e84b8d429f793cad88b87806494
za4cb224361dbefa46ed9b4dc52672dcf6e7da7a144dae5a846f7adf816f987728ac51825c4e7e6
zaafcc4c9a768ac21199c6f15abf1ee65291fb21611fc751fc93041b95b1c622681ee6fca137820
z70a38b67fe4e657c62b5459c6b715737954839795f7fd68b9cd1825b312aedc280b3cc8c55a6f0
zc08e9001658f12a60fff4669937bc897cb1b2e7da26bab29255be88b240ae9a2c83967a4f5c154
z81fb62e7fa70dc5d69319b3f46440d6bb50c67be2889539b8323b50fc42705a04b69e3a6f59848
z84c205b5552309b0679888b7a3b5b7d897bb5e61b211d51f0bce7c6abf04792818fc68afd040a3
z125cf4e5979b6fc1727210ffc2d57bfc935893b7ca238c79bd148d5571a3845df6cf3862e60f53
zb91d3fd87adf6b7541b0f26cfe4cafd00bc75adf1bf6bd660f994b1f391a067ce7e89b5bd2f52d
zed999dc980ca8d727c5aae6264daddad1d94e11ac747202b4431207a280fc12d34510768a03fee
z2f641b105c0ef8a80b1cd594bf3d8af341fefc248d78f650adaf36f2003ef3734f1739d898e4f6
z2978d90d659733556eb6fe3939942122768e561d19d620c8a4efe5eb80e749ebce388c794c92ac
zbe7f12ef6cf6cc487993cb068cac4ca7c99c8a7934995fcc30904300379f174cb00e2d1b2b9106
zffd676ad359ab75d2b8384f0a4c00601a0093d498709a073e43d7c79a8434e7b62b0f23264cb7a
zca7ca92327ee36abbb592d26196b437b995b7b9005dc0a92126ceb743a373dda02ffb28d6851f2
z243735059eaeb2f4c919344a7425a23a62c20f7968257c14bfe79ccc729c7d3916b403624da1d2
z7f05ae87ba0ef91e3b33be756dac8b39f0148390fce526bc956fcb48b2f0b2545f589336f42ff6
ze1074a92ccda9bd176e10a11ee68f41bc235a2f608fdddf0ecaebdb3038d17f508d11b904fcdca
zd1d1acca2e7c34cef3cf05fd62c01eaaf13196e2fe6a688e129e1067db9be614a41ee9487e0ede
z6beaa6376daa57b07409f16dad625d7aa52767b77bdb09e91994e9922ae631e7321d788a9d2c5f
zaa792235bebce126db805306a26bf76b7b2d036220f0fddd39f4fa053efbcb8b1057779672d6b0
z1ac1f5a42c0ea0118ca52f169d335830fc00120d075ba51c3f5a38774a7e1990dcebb2e2bf469f
z5b681ea158168fd3057a08a6a0c236d8b7573790f33d25c7c797b7857cea13f65f4456cc571803
zf71b73cf0234dfa52081c50e8c267b91a24d23c949963c061d8e202868cb49aa9277b5c6effe97
z3145598a0499afdb40fb627bbb94e2370ea0dc69bcb9972809f90cbffad0778daee57c5dd6a245
z43f1c60ca2931b0b4700761e2607650961f1d9322465d44678dc79e7a236736294486e8256ab5d
z9ecf850c60c315c4
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_multiplexor_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
