`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bcfc372064
ze5f6eeec6b0ab5dfbe69335ab6a8a923f7dd5c547592dcd951c059c73294a78e116af77bc6504a
z04fa390e3436886ecf752ab5bfeef2027639a08581a2775d95d1dbc69823be774fa35e22514e73
z499809e221173b877ac31614b0101373697dc3695088bab8f2f6d0f33565322ad9505cb05fd61f
z34e7702d26dc096be0fc4f224d2dd38bc726ae2986c657c0737c3d296e21547a69efa382a7937f
ze767b9ebb455776be9ecaac4ff5574c22b737d797b57485b038c7992f697ae1efbaa1dc907795a
z023d4dfe17ec8b3980b8e5574beb503b16af4292f28411b30bb40cdfdb5802a088e4f57fe8b648
z94403bfc0b6f66cbcb80ecf1e3eca463e0a7be00ce3c5934845ac82c103f26b0ba150152e3d18f
za11c9b1fa6807024481fdd3cc73c186bf2d889491bb79bcc4ec3ebfa907d90812e9ec15dc35d74
z2116936175b8b5ed1c3639d5a35522c3afd99b75613f7540ee4d2b3b873bee8ff2a0b927af8e58
z04673d20cb6993d92b18720ff30935967013f0863562b3aafc56e05f6aa3a73600cbed11b1b695
ze5f5e3491d22ab0c1727f175ce43e40bff39f9f3f445321019f2e78ffe9d7af6527c4cad75b6de
zbbed264057ce0bb59b47bca8e57c09dcda72168aa80f70852ce0d279980e0c2607a0cfe80f9a4e
zbb3d19ff5f2ca0378d2174f0dae2da4a1395a2db605b44ff3698a094a7d3a68d9a875272b7fa34
z4b79e90aacd62d07fb9ea5d382e3797a4cef80bd9942ffdb500a3b7b9856536cb92ba4925c02c5
zfeac846ba7b8490248452d4bcb622c408f1910f96df6ad6d7a39185ad1c9b7003df7d61518624d
zc4121f4c656d5172905a0bfa9313b7ae7c15038def6fc403c0c43b7db01179f1dc8e011e5b9182
zbbe9b0449d291c0a2d6e3236bc70ccaefbbabd454d59709de506aa75178d0fcd03bba3127a542c
z65242bd1bfc2a28f8a0ec181fdb199cffecf46f8b3d0b0179155fe8a856df0231bc16c2b494ec9
z11f7506714d35c9c729931c79660f468e7fcf13b9ee8ccdd10dc94ffed3882daf1f152989cf9d4
zab23c29b7f32a985d50db5091e61a89e7c411a5cba1d1337b6eab0977f7c218d25e86271a146c0
z8117e70d408fb76aebaf42baa0d3f8fe36a92ffe925a2a75ac3b17cd2dea03a544ae6ed825b00d
zfca273f8cdaa809226be9b89f0996ce7c858c0c99a3c0d314a4fa689b3f2babe8cabbb4a213d73
z3bd2d063c098c74e762b7476e494836560bc4abea7b60e42ca0914095dcc3fb46c7a2122b7b135
zbe4879b64830507caf02ba15219aa2cb9b5bd4e8f8e39dd5ca9909caabb9f8162594c9fe457877
ze1361be230b4303129380de8d4b91cc9f4d6cd03204a512f7d78a9713edae518d328b00075c518
zbf38207ca83f0a21a5f200ef25ff6ec1c3feb37c7da3fa19371f4e595b818a2ad0cf3a18673319
z890ef455a93f8003455141b95d21b6c1f1ee40f19c76b69b6a07363ac24a4cb240d41038f1ab28
z34cb775af8e293089be0fda1a3e706a5aaa65d4f265ada6163a45cc42a582b9de49d4ab2f058da
z074d73f61375cd42d41a206fe948e397ac0d5cd107ef1d8bbf174a11626679f2fd3c8bc46a1748
z13da2b32dfc3620d1f620b36ebd6e331c0457f3db0e9934f5e42788fddcafab9da2fc336626282
z3884b294d09b1949d13f56ae421744ca13ba9dc36df9cbbb468e3eef940998fa8dfdb4eb6b97bb
z80d4f229edbee8cf4a77cef84da6930c0b9bd5ad4a55f0167165a7824fd4f00fffb7ee5320077b
z9fe6601e3e3397cbf20cbc7eee7eafb92b08e5cb8eff556a1d4b7c91b3fd0e1c4391c18fcd28ba
z16c2ebc9c84e3f79fb8a6ead32d77e6fb793e945cea0314c5b1dbb8e29652626a30059d3d30f76
zfacf7c4d6b21f2b0c4e9ec62a2b4170d7df8286ad4b1c7648b137bad9e6667423174454852792c
z7e02b4226ecf6dcc0948573fa5a3d475cfe8a6c394ca9880736539086a20987a56c6e331ed0f49
z07d9adc226916b071c87817324183268574d44f941d01f2143681f405518dd3640095e1923da6c
ze38e03a981d29f3f146d7c62184ee4a41788da22e10a04a1d82a98940ee5fcf554ed3e11b968d8
z9b1ed0881ce97e5dd52c58cea4e46ac93601d22d1a122c86e0737e288a71e5642c86e02f73b86a
z4226aeb52fbf028a78b81820bf07ae7b030b97a897c734dd3fe07351b2e4263f03ba8e78982a20
za68b4a0c7f6164f8258fbdf6aec7c82fd5a4f6b7ee984ece8b0e1aca351a7c66a9474afec645e5
zc1fbee7df5e1d10a5a9609a597b174e09c481b5b7f3ba31897670b4dbb57de9473a195da26697e
z4bbfd0c78ca8eca1795135057ce6be3eea77f9049557a09d28e4256fca8a92c85200cedd0f9dd3
za8cd79c80af177a4090c32a99fc2857774bdf325666e3557a443d15c50c172cef2a146e3feb1e6
z51236c049e4de8f6085fea3eff762f863044cf756d6b7281e1712112d3dc420991aec93657bfde
z857360bb2b511d111ba8fe7536d1cd5d8ff0820aea6d431608f7206391134df000c0b171c0e625
z20a2dd6cc87f65fe11a1388c852959efb3852e6a7740f0e9c1878f507bb30ac9f913153434e2b1
z07489ad574cfdc8e28a01b42f8b6e6e3b0ca939f39f85434acb46af59c702fe4c2b30b657f6907
zd53a46a30e730f768a5eafc48a3051b463044306c0b979750aec1c6f1c8f773cd2eefef971ff67
z640602c08e1fc7c13e3f88bede2a638b6c52a704eb93d4f0cb632400fc386cc8ee83174686abe9
z8d029c5fbbe3b2d72c79592b66fecc89ea377b5880d8704e60c66d0308cf18e0aedc5740b4577c
zaa12e74a017284fa4addfbb3ef7b45838e552bbe705e65e47aa2bca26f17ee590a1f5ef1cfd4e6
z298e7de60b1633049a78d8b2238e84fb3d7ae7c3da95952e94013492cfe026218a2baacd8553f4
zbb29cb6535fd97204ea23ec9bc4598c2d70851b42e22fa329bdee5fa136319b65dbd38e381ded8
z6cad1b2646e261982493c71fd85654cb930b77e4a894ef193c2fea85775de3aa1f3f37af837237
z344e0d10252ff55673ebae4ad5c2eb74a1c0b7ca3bf75fc2af761078e3a885c03af575acd09662
z10474caa9e1633ccbe03b8c1c1f7d59958824849fe27e0b988f7756444c95bef2f9266bd000acb
z9d382af088aa1ed80737e012306ec4943157a88a6a71907d217afdeef53e43ade3d0b093f58eec
zcc6fbd4926601cb7a486711167a2e8b340195896bd73ae8bb1b2ff082caee14ebd8cac6e8045ac
zdaef0e7e01d9f5f17d021027a1aa0a86d48eaaece2831ea8168fb2fe94de4ecb501e3c44c5d0fd
z4874bf1a7d8e78663297c4fab72066138938aa3b949848b80372885ce3529ba8b8fedfb5218ee6
z11b8fd466591fec8d648ecefb49d94965541e286d2c17a30dd8609fd5239f57c4b4958b1c2cb86
zcb6a74f2c7091411bfe4c242ead7671fecc8d33226e0c4cdb44d9535607cf822b58765c9c39981
z4d421a4922fd725a1e882232d1b4fdcb75bf7dd026ec631b13453a176760f15fa96c31154ff139
zbdbc44732516fc1c964ada0a8a3472651a7975f867e6b13ca96978e8721da18d2486667e035660
z2cde253fafb42a4b1847cc51dfb2daefc708d8a173c7b62578263fc6223407d789547d6e52b21f
zf72d90353498723f5f6c7b637a13493fed892cf815711500dd54c717df9265880276208d5e8c1f
z59fc0aff093544b8224dd288e294cf47fe3b9a062275dba6c2e9413e19b574ff682b62f7cac899
z8401ddf43ae8d36bfe8cabfab1b056a84571a673a79420b6c7c2bac038dd82d4f9b00b3ae8283e
z6524ee37656b428dace4b3d2f5d78f3db18f757f6fb422f9d6529ade60a805e6973f8423868184
z9faf6feefc5e5f9c2ca3507306088f776d41a3dfeb594e7b1123046021a3932d35c87526d20cd1
z52bf16d70c665285bb6a50c034bc48070e78c66706b509790563704b3d06797347fbef3b201db9
z7751c885c37969dd0dccb6427f963d3a3023987a3d558e48e131d2e23c85e63463a19a055a95a2
z37202d596d8a29d6946bc0c0945e6ec5d256f4165e45b5830038c18f5997b637c712baff5cab00
z6e9630c9cf6990a1d6ae32deb9074a80039c446ca6943852221ec7f10b041bfc5fe8657cab9f60
zb89260f4aa9b78c578008e41140194c3686d86b6c31bdc5d0f2586ae702f71062c57f7d50ce320
z71df8d9fb6cad0773b6b4359cfd33220084d065c39038ec026c82a32ecb5bbf7aad3090f7222e8
z8fbbafc09b3624ce2f9b382fa5c5ab5ed97fdfa9fec6a25e8fa4957f0653efb38a812d3dbb1fc7
zce3208de2e947b3bf6630d757ca10ad8b0474b86844d97c180cbba385d30e71f25c867a1787f01
z3284965df675187c6ba8ca8acb0fbcd549e39b309bb53f10409ab4ecd92511107b7c85e881f597
zcc177a4eecc7eca53169518b2bb469231741702ebaa1ba0f3122dfd53cb62f2df50a81cd98d2be
z1f8807f237c61df51cd2fa30fe027b1d2549415dfc474a8b6f66dc14c86a6845055976c73af7ee
zc01ccb1bacf7592789c2a6b9b975513933e32f4e28d6f0920fff9a1410d5cf3afb928a9aee18a3
zdf7a3daaab99f550ae49a0b5bcbd77a89701927d94c2bfc6cc5a307e90f238fcbc9dd87a18eedc
z5ca1aa777442f035ccf620a767d8fc8ee3a51d34bdb6074b9c8cc65e08e400b66e2571dc51e989
zc52934b05aa662add43b73af3d80e1625cd808646db17ba6190c5a0af6019924a0ad96a3bb17ec
zf7740225db87f9a6c2b133f7c452fd960a5e4e76fc893edc68d902cfa833d6cd2a449ef379368a
z6e0a1cba675c74d63b1e0f92d0c01174e8102c121c9ec78e4ca277446a87730c776a1b2725933f
z3009847e32ae65f77b21e189b07b9292a9ac9d1b905828a627e8edde7fbac891a59bab37dbf66d
zce1c5095e426d8b7ee81cfdab4c621fbc4498fc16cfdc75012e5f934a3056b234a2f7fadb0b7c6
z620b2a6e38616a2987100818d8daeaa18c4747f537991576b668cf46a794bfc7fe3b3dcc123ce8
z32f3ad08987b99a3efe3858df4993f893af490f5ddd9ca9a24ae1ed876a36451ae84f44a80ae62
z2b18aa9909591d0043af506d648f2fcc0b6bb0e76aec5ab3c7f8e8b1db3b4f58cdcd843b0661f4
zdad3ab46c5e8c28fa9684e58845942e2fb1597602fa4937f3550ec3d9af06a82c2551b735742c5
z72244ebfa5e392ec23726e3d476b42407b957eed20cfd439d0ca59759988fc611576a673c91c72
z15a546b1eb4982fa7947f415d9f09c9e2728e142ded2130e42ec94f33110b6d16a6b87b86be842
z9ca7091e6b63422847fe7197b47321024e8cbe8583f63df2ab3033791c9a1b3e08ad07dc2cb8ae
z8acba199d1b98c78aae6d96d01e54cfaefd4c32717858e8d49b5904e5a1cdcbac972e5bb3b3536
z874b2d53d6ef291823eee1e7264c4d1ccbae9b231c6c92892e2993616bb92944feeb412b05126a
z1e552217bb1e4d2e503cad59adc7209e9691d64a791850a4d6ba275a0bda9556d6c6e9d561bb6b
z3abf27580494ab9349baed5cc7c60ee8fec941d08e58dccf6f066d90d69f04c956658a395c6eb2
z07903a556574259a2a79fd1016e8c7db7ecb1436de8dca6d2bb8adc14bcbed35d8b72fd1dc1b23
z8022b432ee37110f375410e1d7f515b1d7ad38c0482ebc92bb5e77d3690352ba8ded8f777b06dd
zc9a087aa428e27e545d82fd6a30dc2e967a103bf49d02022558484782ac9ccc875812baf27dff2
za1a0c40475a50b890b7b8101b8f0c0c6175df9669ca4b9992d2576546abd830841ec7649d276b7
z83dc78cae6e2df44d7b908d039df9ea05527d9481efb32726859aa90128ba62fac640990e28d71
zeab67a9ba6449f2919af391f13d88b4f51e4ba88cb8ab41b97943ddf3fdf218afe2d26c0877307
zbe6bc9859911736ab1570d9eaae322d59298bd91a7ea91a6370bbddd27d0e7a17b1bf5bbc7a499
z13faf5bd4f1ff974cedf31a4b6aaed53098638e279bda54dcad533b18d86af4c9d64583b825f5c
ze2a675f3dc3dcb40ea9a0bbb8bd8893ae2a78b79223e252b1a506679542227c645bbf27d44ff21
z0f9158ebadf7206a81dc6ba9f3a77228c11b3e13848668ff9740d1daaef89946ad0d928818744d
zaa0f1245caead4846b647e37407c571b0f94291b9be64ab7ab90d4ef2bf4ebe1b5c4deb0199eb5
zcd7d800c5dba8215e7f40acf6cc22ab33d322e10842fd62ec94932d7b24547199c457f1431da11
z1998a150d8e847d2391e8028ce9ddf474a453d5632fd2afc8323b4c0f23fd8b3fb5f56e96dc721
z4b586af5c6d22801a74d9cf3e23441b15c1d5dd7ee34eb3689c29c9e48201bfd306125b6e015dd
z767c61149652caeebc06d302b4ba30d152ccb9b368bd5697bfe1db52f970de223ee4065b14c615
z8ad9a1282efe31cb6f0f39925ded9bfa4ea023762ddde39dc5ec8ce76be843b3d4ede88e75425c
z84d4f59bcdb4801f504f51025016a8aeb84b4471c80b6d7319bedf4c4e997d3be81b82fecb1d7d
z2e7ee46ee50ae53eb41437a0cccea5ee9d4c5116d4b5f8cec45b02f346fdb9901212e142201663
z77372eac3d7fc2a4c190862828a91e2793de8f07e9da4a7623eed86fd60943f65fb931afe6a17f
z8e50c09323153b4131c535c4d62d1eff60b2c97672ee730292225a1d3797934e0397b0f33d23a9
z4644fb2ee69c2fe322f6615e293ec16ef9107384c6e8aaf53144f98d1b5df6ca8b58178f20ca64
zb16c4dfae1d1d84c37b5cf7c8288575bdd9c70175a41e98fa1d06b50a4bb36d96ad08aac3d207f
z05ecf81005e4f5e86b85181b7d7313b234300f402e2a97cd7e1d2389c69a2e3e42f4e6e2d0d93d
zadb476612e05d90590d8cc6fff9248f5de0846e8f39fb3ff92223b9c3eaeec3c85e2a921c2b853
zc6cf25f724ce789301fd4c99a0ff41d93d33c3c476128c78500eaa5c3c6e07e8212ead9aff505f
z53ad952f6fffa8566a71ea9a024c79c86b0058e1cf908783a58abfda0f746cedd6624a23281163
z6a3a33663a17299387159b59dd7b28d0a6eaece7be3a3105be03e68abdc275ea35d41b222a8151
z40aceef49d63f2feae3a162ec5e9212c5b49f02ccde6be609487ac8e69221699f573e12361c243
z933f4b16587fa3dcd1fb726e20def1ee58dd9cc9c4c321413b414a783a7ef745157034bd426835
z10ce0866981e742daed7f74d36c492fa58d462abd6319bb88bd8bc198cfb3476389c61856eb44b
z990d20d1b35c92335ae621cef5057081603e13a209a7aa186f98b024c34dd35bfb56f7147ae390
z95dae78faf382fa50a6ae2a54273deb9f5cadae2b062c562eb0fe72298f5112df6b35beb30beaf
z3475132742839a7a00b3d2430646c03faa7805a6c5041c3a290dc84f1d845c8fd3e6fe600e414c
z43de598bfc31cdac4e96c40e4c71fd66672f1ee9428f942eb7c6b52e666b6022c42dbbaac56c60
z11162bd47136a3609e64f767e4eb0d44ebf89b626ed38453cd57ba5e2ada0349db75e125ca2b15
zfed89f9fd7495544338abc961244919ddf20f4a980fffb9a512828c08b24ef64db9bfe4e7c46cb
z4a7470543cac187f6c67470a4da8e30c3544753d1ea6361939d03b7346ad33960f67b8d857e74d
zb1b47611ed6c698b72b7db89c7c2da8c8838b734724701139895c1dda7612251fed4c9100381c6
z4c110a9e135c83679fb232969de6e80fda79cd1c0968bfa91964c0625a7906fc5808f0a230118c
z37f6caaafd17697a58db0a70daaa0eff51ae15ef1d9020cfcd790960db9fb1d1d20099494fb34f
z3891d040c1f563302b282f75f09ae5991bd0188fe3dab41db5ef3b7cc33927b6112aee27a4cfe0
zdbcb429d33c79b703e140912ecbd470047e3ed5399fbabb867087229c9a1eef757acc66644a5ed
zb94fdd85b58386f98067aefef6503557a23a8577ef43682842a18e8326e95e8c6a37cf08ed2139
z2f625ad414b2898e1fdd0fc45d28816af577b5d7413062cb7d9ba6b3167b5d3fdc22cd42c1a850
zdeed3bc0c1b2c078a11504a0ff97bf4e7bc5a409cafe88d30bf2ea39cc257b247f614dd2768b02
ze905dcd8f56a104838ce4f5d207541b5e214b2130830204ad906b5d4bcbee5245eb67f0c71a86b
z25a80612fbc80a236bf4088a9cbe4ba6bda969dc1ce88e62c7ea6366594aab50347c9cfae0a7cf
z871b06202ff3701a6c69dfdee7bda466d1fbf9f19f0497cc522b3373577ccfcc28bfcc07f4d314
z7478bf8c23c3917511127f6ec00891150dc182f0c76afdfe78e367cf6b362bf2e7b773b89997c6
zaf7d7fe8b0741b7aec6d63997f9b58ae804a3abe1ef1223f2fb4c95ec15f317b393bee4e1e282d
zedd03d61b20d374d89607d189919879b5e31ec81d3e62f40f98a3a7499a6f3c584c94fc7d63331
zebf13c1690444f78b55829fd2a81129597924243f61a420d3e13504c2d9b1403dbdd836495eb07
z35d392c9efa1aee805f4bb716d58cee0df9454ac118d884aba9a69cc0bfc69072323215b97412b
z5bf6401fc1e12b85874669616cf8c7181374db26b0674f56eb6bf9c1c235d0794d5215a97629ff
z113fea6e030a594379715aa3e49615f522c8863afab597f3d386fea97954fffc37b7fe015127f5
zfc7cdc0bb35dd3110986fe00987e01b23956450ad576532b61eafe16cb4159edf631dc9ec783a7
za8b3d801e95865c7bed3481be703ec6ea1884a622994e3b07cb5f02f2fac940d75681dc3b0b62b
z8cf3543b177ea92cca02dc042b1f3152d34325fed147864a2514da8f4502b521961b77e58c6e19
z9774e21ca319c4b7b8b7bac42c49d13657ef54416c7a6df1080639d7c636bef96635cba63a5f95
za0fd2c4b192283dce5ab11425e1a4a8c8b41e39383f0e0b2835001c31f08e449396880dd7da953
z7ddda181ab264df06175a24edf01d55e8ca39199ef6a99fb8f484b6cd89702325a9068be0d66d8
ze09f5128940f3462e64e68ede11765ebacfda3a69762625456b796ae4f5865718f5f437030d3ed
zffbdfc6370afe91a8bb201e442d6b6582b329af6da76ca6e033e08580c36804385dee24c9016aa
za5f8b9d9274db07d85aefa08367cfd2417b3a911b73d1da031703a5c50ccbf5d35ec71dae515df
z7c28c8dba371fc5e650da96db976d48ebce8614cd8db682a85bb8ef255a145a91417f3215568eb
z4e70b1e39722a0393b226eefbdc50af59cdd8ed29868f6e27e34b30e789e2b873b4dac25b808ee
zfd63e6e0d9cf04cc9e58aeb950219c4feb5d976e69dede7f4fc284b97a5cffbb5e8c022becf8fd
zc6162bd34267f0da2b2feae7362144971905027f87ea9be53d7e83871f9242fdf219e463a6b033
z77315e26a8a1a19d8c491fdea36a44c7e747759dae8ebc99bcdd9591d496498e5047857eb69764
z39fb8f9c10d824db61925c4ab9c952a105c5c90d0de0fe8272165fc21d74e50974f51eae3b7375
z8eff9fb7731d1a8058a1188ab7dac5ab39415c7386977d781c3a8ebc34909bf5dcd17102a832e6
zd421d4341c138741b361b2b33d6805c82234596469f03336ab19e0f13425658a934169f53565c6
z176f61cd1661f5e8d48c401875af99d0e5367ed011f134018fba9973e425da82a8772c88fcc6bc
z1e43df3496ee52359c47e8dc2dbd1a8b1f956eb85ed5f68ec7f994da76ec355d6cedc0ce7f68d8
zbb2790c9c2d41afb02f8d39b493c55b7f3c97b77a000dffe515ee663af60cc69d40dd20be91f33
z0b1ced237684967219d426e3c63c966c8cf9781dfa2696632a93efa72cb3f9f8fa79d1cff5774c
zce266fd78970a5818c3d441725a0c7e5c8cc44ff0605fa306ba2a5c00ae85f0637ffd1c8749911
zb5058c482c8ab37e869459d38f8120cd769c618432a2bb2ae4f208d8caf8a813125e79e244e490
z3e9a17d1c37e8883dd744781bf8652e3a860c591523825d9ab78b327ea74458f09a91a3b94788d
zb58a86429d3b55107e57a0f4e7254d33b395886293a7acad76190d7b6fe18613644d177ac84a3c
z41fdee8906af9b23b587aab0289a603502004a51b3b0d81bc1d3708448a903dffa9f7fab08367e
z9586650d8c167af89b25d5ee84c806e26921422dedc5af9de2ffbf3b45352d7181d45845f042be
zbe8fef32a426015321fc6cbfbf7329d614596119f76facd7a29c1b98b0db19cb0ca0d1088fd486
zcb3e5c5f2e17aa0d4ff7327cdcbb4ac8dcee118bb72108b7b194c732ad92329ea7adac77d4e56e
zf97a9b756fc27e2aa7fd3be1306e596d65d5ef7af0315a820c0675063e396d452befd29bd445a0
z1c198b2da093825381478184be8cc9659c3d03b2e8b856e47b2f839fa80cb38bc47cfac1931907
za849e2057f15bdf67d0ccc0b434c79ae1aec5dab1cc535ae03a88da554ccd1753ef309f8e1733f
ze49d5dc2a3b536041b8d16499c7fe8a1bb9d1d2ed481871ae2eaf972aff91c3853f9060885e8ea
zebbf2ef7733624b9487af1cc6ca9d8c1f9051d4c6791246c2aab7440ee57a453c5739d195786cd
za9f8b31648553ba0a5d1739db9019f57a04962bbac780c685418b51425ce71a6c3fd0ff59f6e94
zeea4dd1b4dfc04868de92852293d0390b85a0b26587ae281f9aab11858509562914e5bfc505b19
zd6396407d6bbadbcb1ccafb7cfff53797cf01a2c7715c2402f365d85e786198d8cf4933d6b6a2f
zff161ab534a881a155a9859c4bf4ce2c613fa834a7a53b3ae20784e84a2edef1076b29892b8a45
zbc7eb1c5711c9947563398de44f2b217d7d848eea5e57059c60378535a74ab4241b7b1bfa80e67
z0c6f0921958366aadff88cca929e1c29a072e04a3b73ee9f5d608ca1ae05072008a1d496325e16
z24268efd70c202c900d117b9aa3d2c05d37ea6a4d4ef6b93db5214673638161c382e63d9b439bd
z4bed6aedcb1cb6edda3cc6402d977ef2b90a514974c8f30e0f477f11b8ef6916099f28d8b4051b
z4d89b17cff9c9809b3d14d69d772d294a3d3ba84d9c98870c5cf9afc15c01fbde55e656e186bff
zf3735b78fdf6831cee05ff440eaa1ec09e1eebc1ea1d174b0ad23c662c3dedfb67d2e9624e8c7e
zc5fe5323efeac6c7d9b6402eb7c9c9a2e85081f46b4b4cc0bccfb7644ff22e7aa15b754aca1b8d
zaf838ab66bad17c0943b3cb2baf328ce4ddb5bb3748510c9741cf96ef3ce2f97e0371c1b58b5a6
z45591c579d7cc34c5acc2d650e083302b99414f424aec97d6f31d8f9cbb3867792ef6ee8e8e11c
zccc4def1b26e3c75b3146fc9324f021574439cb704f60d938a0a13602b10feae989f658798edee
zc39d2e5f294fb32dcc085df66f9f0e6b34e1cbe5204f737ba85e61b52a6f9474047d4aaaccbe43
zf25afabb752187ef9294ccff3fe6452efebf7c052f14072586913f602f0d4e82bea4ada01afca3
z1847a193f0cadb5f4e59951b961e73f10bc834f82e7c2b15931fa0edca67b20ce64b58cbf90369
z4428970f06b1c93211788fff92f21b0a75427ca07b88e1601b448bd0bc0ddd11d63e068a56d53d
z5145c62d6d8f9d5f79aff40f47277162ab53633ceeb3cecbf06743a6c6500841d82c4e40feb12d
z1c44472943320541acc164df2fbb4812ae43e6a71452ad4c00630f4433a6ed449eea763d5569c5
z15d99c3a9fed9f23cbe46732bf7ef146084f6a90ef1df6bcc13fbad853ad09801d280d3996420a
z14fefd49ad4d225c8f29bb573b62a69ca919ecc11b04a9e7e1a1931b9f0903887bd61485a43b3c
z11b5d93cf0bf23ad29044a3f572b55843e7e2f13fe9cf4d05437a9357912ef8194ec1913e1cf25
z9de438deefcf5d97aa68c99451d028e62cb259b18c1dcde1e0a211f8db42baeb125884f8459a75
zd6fc9a0a2e58da2fbd61af7769147e820830fede93ada9c72b5dd5819e93650af4c2eda8d0d9ed
z93cb10f2a1bf99845010fa82233326402f7197644c3de2e6e1108a88de442b33f52a80a54a0b81
z361b760a7cbb5f90bf3fe3a3ab40a7fba57c832e82476e5c6224adce47e5a8940778cb2faa3445
z21493ac27719e2813edd11b483ab77aaa78cb75622167886f74629331807255c2ff833e8a1ad04
z06baf9e9ac9d7012101b98dc5f539dedc6902ef021ba5eeceb185b9f709015174164f93d4e9c4c
zcdac110d303ee8372811883f5dceab81626fdad8c2816f62253d22c90a47b06e986ee78f34b429
z2c58184304d3ed318674d4cb336c74d0d223f6790cb56e0624ae6d49e2e385e0e1bc866b3a6909
zeeed1ae0632913ed5c3c2d81ee2cb91f91411b5c692f1424910e239d16e30c28f9ea8302b3cf51
z350f6cade4f2dee965ec31059fd62e193c3f7bc7bbc63c5e3c1bb753821b1c53c8c4aab30b265c
z380e02a5211c69110c5a35ec077260aad7d1f3f4939322a28f78f8dccbf7ff35818b5ed8f1e803
zade96cfd4d0a0df666dd56d70d8daede438582e4a83b94b0bcef8c8d99c712812821a2bd102909
z8ee564ce7c34d1ab63e88c07c8719bf07436e1ced1a111ab469df85ca3af2d7b95fcb4db442dd3
za343953913c95d4e670dea500835d11f1d6d6ff6a93d50689af59abe3fd479d85f325c574b0a32
z6be31c369a70bc1396499bc1f85a96936b2c4740aab3f86925bb3b6f3b07eac6fc0bf3785ed6da
zb928b9c7204b9963dd45cbe618f64a2fd1fa4d98864d0c8f892ff92e20954999e6125c40131661
zad6e9e84d8a2518934c50c92ee91b82e000ac37d9069532d155083d425e4227f640ea14512cec2
z72362b924e82b758367649b360ed5fae59b84c8c31624e380e97120a7c45af8168df16bafc8c21
zc89f7d21adc3fcbee5b4bfc2b49b723c26ad9edacc94f0a7d6dc46ee88dd25383d1052394e26e6
z03a07a6e350dcfaaa1e49f44397c75b134e0174f1b9f8df10038e93bab790e74b3339be4a9edad
z024e5c47fa3d68e43fa764cbcbec51670820c794d8d3983c6531af91f862366798fce17e0b942f
zf9bf70c3f58c751b4a7161f2bb442e9bc5c8a93d9d1e1549ef45ff4d955bfdbb1384f09c5cd28b
z4461a7f13bbb325eb56bfc88623e46bd316fa4527fb115cb6c8bdf6f4568811db86381eba731dd
z2a36327afa706889ca3b2faf90a25ced6de9929f4504322f7aff956857142021e5c41c79ce13ea
zfc5ffaca27975025f306b0e71bfe1e50afa225d0ae088b8640162a43b427a2918b4e8428b739ac
zab162f9a531627b5194a9e5eb0fcd5c8eaa4fb933d92040592dd9fdc56415be71fb7a18ce630ab
z0cf28f325cf1aff496617a76185772eb21ecdb017caac202bc97d0325a0b78fcdda0acab1b5498
z3f97178e1615672b0b4af99a85c143dd3d7ff0dd2fd19b905f9db433b266c8e537e5db3667fa84
zf5863acaa0393ec1da871605274e5245a9aaa27550a14b45d2add14a75ea239c3eb10747c1697d
zb0e1c4c79bad4f496593170fbaa244af41c0b12963af308700d9aa747550aecdd1e4d0e7d5cdfd
z234d435747382a4980ad366b3936b3d3e76fa40ba711a414c9583b6afac025a353a8256e92121e
z3081f5dd524d7fe22866311ba8a53d17ef12c6c0e6d92cd8a97e0981dcde4be7669b42d4f6f5e9
z246e32f5d5e615fe27877f3f760001f0d5503e6a5431a6859ffbe260ab2f6ed5538e3796c558bd
z5f5fef7222e65785fccddd5d0f0d80ed1c34064c8e7db733b85c500e9a6b0052dcd44c7027635e
z9f429f33350552ccf00b568dce1d0471c85818d733e7c99a1107b4aff1798b353108469f0cfb85
z7a23737b2ec140ed0e45610af1a9c4bd150181273f2efe65abba50c9a1314fe4cf43dca98e3d2d
z30540c95576024dcd361d9ac4cf2ad3ed62e5c396959b004ccd18203460ca2db01be66a6c51bd8
za4fce99d0fee4a50398067f2959d966a3b3fb3c01ebffdf239935b16a6646b608b0aa17ba4c473
z2db50bd656f59574993f14200767ca7e2a6502de28ae238fa0b0b731c25b03dee4378e7acccd7c
zc9fc7ab46dd75c8ba1527943df8f35e00c776302104d48668f4824483ea8acc0801c361c7de42e
zed88d6a754323e2eef41e4686506321ca7991472fe263b71ad8d8d7687878a2a60846e1ba9a329
z15de668267fcfeb97f5660c11c217b4d2d20e8e686d00527e392fc03ac4677a548ed7a139f5b1c
z9e327a5c6ad1157e7670845614ec5595c15282ca3ae4a4e4c47fff6e8accb44f55a23831a5d5d7
z3a8967a6f150b59fb95ba2d0ad53f525500944c964d16a5e489c7051f688b208dfd769e81df464
z081b56d24834d0c32b1fdaf7552cb1a4839cbe65fba4f5e74d8065807ac4af6a109f61400acd5a
z1f69db6d6e8b2b91673a53f6b40ec1c9ce15915a78c54f921ebb7da92ba9387a37bb8d4e5e9b49
zbafaf27fb64fa40f21a48c546d761f455d42afd28734aa32de3f73905ada77c27f3767e9c2499a
z868e6312426f3c8a668a78100cac5f22d7d7d6e937858da2ead513f69a8ad4a9749ab3c4aa6846
zaf70ac69c9978ebc70ff3d92cdc348a8fdfe3dcc39b8d62b6a6b26e4e3e2cc28908be07584d696
za442e1edfd34499496250a088e3fbaea763d15a047ae6d7f4a32f575b7b63892e0bb43886f1266
z5d9e6babc644cc0d8d3c6b40b33dc7aee3bcdf06a2a170f0b4ea247b7c077e0cea6846042271ac
z3d478ad40d520b6be00a0ba3b5b311843e5775fdd892b6795b285c95c8167fb2b9830e303fa95f
zadeea82054d68779e53e1564ad8376579254dee20de5dcce40600c8301671e8f20a01dc47abc96
z9580eb52fc8024c1018359f85a2d29f0fd231a0e6995ef1b103e12a2d002e7411c7487aecf2c4f
z1504a264a8cae1961ca0ae49ea72bfb4857198c6529dcd272ebec341796fb1fd046b629438ed9d
zcd1d6408b5805c8e98e16cb0b3d0247a4c063b694205fa80c0b2048c3fcdc2cc7bd5355218892a
zc770313d1f60efdb1cd8249599ba47cc6716945ffd6d7496af61e364fd9ce9c89bf764516d697b
zfbf5a2d0fa6b95884d8b14d74ebb37456aa966dbae359ea22a2001ffe781629d6f3b8d5ec957b9
z4cb75d0ec4b48245d79d0f62100a50edd1aee98c2462b9adfd5c032c11b686e14da293baf5fd96
z62172da11ce96f52d972811616b407bab3114dce5eb9a1f46819ac2451c0026a47a6df0abbe0e5
z04ad358c93de20e98cef0d58917e03e97683710d17c681e2490fa16aa961942c25490a6b3a3e29
ze628d3c87a2ac28d82c4460c9fde3f7845696d1a3e4bd93d601fa3bde9813f7d4091fe152567b3
z48f9a8073b97f1f762acbbf75785284128ec893912bb7293c5139771f8b9dd25ed7575f4b81444
z3d9b1bcca1adb3ad90e56a60c9598347714e5784d266febcf10413b709326385174e22ec9ed5ea
z2afedf2967d7031ea13ba0d160bfaf37e27335237df408586b594ed64b1437b74c97f64c67eff8
z0ff3d47d98595d98811bc8659eb22fe3c837456ad7623aafcb5d1e6e1b290ba78be274347c2437
z64ac3bad969905720184fc0530e0024fe11346ea6887f45ac408723432ba1616800b02dc23d488
z0a609faa1a031db940f6d1a55f1f56dfd3e981a28171e9032fcf86d8c39ed5ccd23e161fdd1945
zf9b10ad8574df450611fbee6acd07bdf894ce53e7685a0cfccab9f9de3fd5200b3454e21325c55
z0c9b2edac614b1341c0cc6f7dce164e95a9f7724708e1539493b0383de5816def720288bf19a28
zcf98146567f0d27a6d5207a90eeff727b42c28a1fad92d476bc1819dc4d29d26f1ea27740c2ccc
z46a88a24f426843c047810e407bc5110d3465532772eaae08bba70feb75b7490677cee04e48924
z2924620aadda045776e57925a3c4978d0d013390b7d96c0ae15a9a0e2d49fb08dfb5a79293753b
z17ea22064894f485d09012d40e88b644b090173c3ac18c59e8c6b6ca320db879c88dbb41f26f94
z017d73257ca09b5de9a0da6389e4a02eb3cd5002cc7c94b21219a71a938f90fdc701c3487c467a
z9e61b10a930ce7ae1e5595e9c23ae1b2d7d79594837fbb80589dd2dd4b790bd253c7296a61e758
z3443305299e49dd064c48ec378fd439c0355663781d29b0985a9b6f36a64b2e14fa041c9d765f9
z77f321624587a3f745b2a99e264a4bfed013eb558f197a8ddf2cef5cbb481b0d4de2ae89207597
z717a7dbffba0d0de571fc35a10b673cf64e3cdfb9cda7004505c8ac681b7e693cb6ecc07a7080b
z37949e78da89715e33bd04e4fcdb3fa84a6a4615f5bd7de00d400246e335a81a449339321b7d15
z584095bcf212c2b47387cd762e20b2ffd575ed79d6d2ee4404230c442ea38ecfa95058aa7269eb
z7fa0f2a20ddf5b783d534922438f61237b2a2740fc7933cc5de12c638758d46623438b525c7637
z543bbfdc54b3023cb03bdfb616748caeeab44f273e29810f8e5840fcaa731c47eb4d406d1a473c
z1bbcc87ef663355a5eb2896df4d85018875b2f6f0bf64dce2d929c15819194305d1294f4b4f95d
z0bf46875beae9f8b8d4edda8dade821019518f56df5a16bbbae34aa8845561ed190287b2f70fe7
z0256bdba1d281f916106c54af26feb336c914b7fa4980a4aa7ebdc1672482cd1605d68fc953f95
zf2576996bec39bdda5198398b947ba4a868ddcbf57203caaf335688020dd7f91473903d0c52cbb
z708f88d0a9c9046bad5ad0b33c8c4ed087134cd605683748acab953383c5619413c5ad9b0b3a57
z6092115f51fe6f77812f04873429d4a2ef130e04ba6e71c50cc731d9a40a3a3029c2ffdb98e218
zc90e8e2ad897568640b5011b69eaecde52ffb9eb76ecb90080dd14a8f55e2a66091e09bd158ad2
z3cacdb03d236f2149edd813996343d858bfd219b424d44a9ed0f9e926f13e22a2e2c6281079357
zd0d3f483b3ebb6ca9ec0b667a7eb41cc7c46f01a42e1fb57165e2ac4b53cd9b4a157f33058ee34
zcbc30ec4859ab7559ac792bfb59fb85655fe64a20b0267e8b7a0f7a828553d32714bf63c4f26b8
z43ddb8b92570bba9a334ec3ff5093c4e791a2b9bf616a3260f755d2d06612886d3910b8e3daf17
zf21bf54d210551f216bfe7d2656d9d9dc900f91500e7828e61da405b73e6cf688643ac8cfc9a96
zcf687dfcf4e238e6e5f2968689bd81144673d2cff12cf4900a2007acf51c7f7a56d7b04c7115f3
z9c758503427f0658ed26691ff3c8089c36cbac1dad5254575380e205e5052bbb92cbb912f6ebe9
z4bc53d747f9d28b28418aab6cbc071b57d22771f9f4ab70fb36173ae16f945aefc167ccf8ac6cb
z76ec0cbd676f1947adda4f1be3a23b5658c436e4f252b65b21f3ed3b4a3f92da78e2c7563c37aa
z6118da3763d56a52b659a9a9bdc49d7ba6002c513715bd5bb9f27447245e76f1991ae993e06ba4
z0f0e9cad0ad122824656282c4492cb8f10c93c978a6812ea1b43dddec27fc437ae1d692042c094
zdb56992916f49a7168e670cf618d58e9712162312d8cb3b7b3b83f7204df58a74766f01fc079b8
zb0b7f757f722f7911b778f108512830a543fa882b727765940e7f54c27dc884738f6696872536f
z42fa258e8835e19ee608cd0c3868679400f42e5043a450ea5b10f50b3f8773b43732918ee61218
z9fbb5c3a7a5344ea4568235897d9d6895225024475e52ce7b4f8784d9c6737301b210abc356964
zd992f99d593b5cc9e0bb833d6e7fbe482231b477cf49dee3138ff0d8c509cbbe51f0b393d073a6
z2c77f0b6d5d94af47630c191e0fa1e150ea54eae4f2e2c71a38750bd315b36ec2190e50c5cb9b1
zfcc8b4f64002ea06bc5e30a262040a83451ad990149e4d2a770559086e1c2b289650df146f36a3
z545c9aacd0d07384fac7b5950201f7d16ed5ff5ffaee7d148cb97f638b7e7d1bb577dc6884bcc9
z7a56fc5d4615dc16cd600a491a31f7600e7f31d1dbd8df4d1f398b848414f65731bb6997932af3
z29bf0070520a8d6b5757a3658de61a13069d561dade6beb9443225556c2b03c640d1ad5e5173df
zd55d05e93bc831bc030a2fcf9aee63bd4714723f385b7eaeb79c43402694cfc4b110cb1a9f11d0
zb00c615042322f9a818b41b9a2cfa6f1c844a6d53530b50b1f170b076c214f0a737ce7e688b40c
z124daeac8c62e80a5057ef542c677a6a0c12f4c9bc6f8f7b43e21f86cd5223d0cc05d4c303ff5e
z3d14ef49aee72ab51cb7551e7b1bbeb5c95afcb6f3ad01a1a45ffd407eebee9f6a11bc99aa815e
z8cad07c9653828c0c3fb61c006d64410dca948f7625bc07511ec6d7a9dfeae6f31cd8777afbf0a
zb2fd8beab913555c73df514965bb04de8782a5550447ff956a273afaa6b3c3b01a0c1e1b57bc5f
z88b5667fbe477863829c62db25863d32690f35b82ad1e7a4f9c0c46b00fe5cba7f67756004ee92
z268c34c86d26b5feb32fee0796ef5c6ae1986d4461ea61b70c16a411eaa579bd2877c5a0cc6c97
zbc45c3c3adea34c9d3d4fed5bb08c4e359f286a482ddae256c0c0b5a0949faee7e0032672e391a
z2e5fe4cffadf99abc59494bcf6a97af5b392f972bdea529db1fa8cf4fcd39abb1cf2c9eb217385
z9d912e6d60be84e998b74fb2ccc4422ea9dacbe0e45026ae717550d8d6873d0bde5664645cec00
z9c86c06949b1fd657ed14fc945ee201e8dec1773620883d9cd72cdf4598f23e01e7f7dc8f5a5cc
z7cfb6033e4189d5736ae9fd8db0e5621f4fa5596e1fe6bf4c172d2c174c0f82692d6a4d2bad6a9
zdcd94f1aae1ce6b50c9da89cf980d09cee6937eed29b06582afacd9ca921b29cce5faf7103f900
zf6e3c3cde8e26ab2d540cba799f8be0275fa423a8c6502a8caf06c8849a821896fbd5d9039da94
zd7041c616aa900ab257a245818586429d0a568ddf027765af3c4e5720cb50224221ed8de7cd414
z547fb572df0abd17773da9d057bd867c7c97bd08f1f444fec3b60200e6a1eb2cc7582737724698
z20f6d0bf841bb0f1f2bbb0bac7e5bf37b2f0686b4ded2e338c444be082c6c01262767a47cc678d
z5dd71be020a3d274fa1d748404484cf5ac7166a9f96fc3fad93079c1a8bdff400462a6d5bc43ca
zf24b9b2d1672cf368a2789915908d37dde5b28b2fe23f4c010acf3487650bb4ba07ac4c00a4e03
z9be7282eb9b16ed2c8a87c02c3b7ff8db418e2e29fa8d23bb5b7173eded970e13b3392653fae2a
zc437dca2ff17a801f3a9e1da637bb5842a06b8ddbb26c0dc8680002d720410da258dc3e29d6323
zf5888c27b41ed2d996a4aa5df028c32c5cda1faa08dbbd4f740dfbd1e900ff13f50cc3e6c3a7e6
z00fc3c3e5a8a0325f947d9c26afca45824aedf0f86a36f0ef4c05f8987f477dfe70d1fe684816b
z6dca88eab648757cc49266ea8b7a16749bd3a9dabd44c8ebff3aaef5e9fbdf9dda80c1f8f4fdeb
z87625e8f1ce718f906d228c67cf50bc062d447926cad641c5f5cd5bac73ff2f6cf210bdb21abf2
z5517e1bf7d284314d745c5b5295f37ed3143a908e3c4271cfca218f0b6e4343dea865ea386b987
z1e33ffc9938b6a71cef52227705ba84eb9ea0f43df96681c7eeb634e3c26fd75a1ee56f434af1e
z28be8d78e8ae253ef22ac44889c2f46ad8ed37ae71af7fdbecf8d801a0484b5ffc01475b20f497
zb849e3ba473eebccd2c68b520b77a9f780e7b7552969649d34f74920c3f871c08fa78790ab8308
z9eff489dc82a16818c0070dbcf466cf325ba5cd5b98226122b81f615a6511d0120b80c28356bbc
z183a68c478cc763820b46381f75e5642c1fd7dff517966c7c8ddc3200ff2b5893928fe7ffe6643
z633264f4648254337275cb8e89c800810a6d93c98654b1367003189d869e9b04b910239be71724
z64f900a694550c2d9dbfa04a605cb718d10974fdbd8f564410d196a5d95b10a2b24472b0c760e9
z8b163fa27c8386a0e029cf918e71e24b3e09242aa451819abf3ac0fdd6cdec34aabfbb149b9ec7
zab2edc9fc66cf94397d65862af0e11789900ee467c68392cb6feec0848aade8e2678e9abf95d89
ze115a01d46b649edb9f866d066bef7d5669ee8f75dff09963bfce0cb83c9163a4f2e28bbf4e987
za655a897a9dcc4409fd308ccd12ad1d8a0938c7e2239e3272037c765d3798144fd50955bebe99a
z28459918f2f985a1d20838f7e197f8b808e177df31d0c0914de937dd1a0df59f22ba647a2a1ed8
z7966e1747c1ef5e189e71f0ce00d546a5a54e13729689ac0cd92b685b656d18382c24a04571b74
z89d003c2eae6ee4d945900a8ec2c4c6756a1ccaa16773ccafbbb60151a1101fd8db89b97dba19e
z2e3055ab1627a1d72bfacaac9fb106d1bce91d21515f758ad28c49aaceea3e7dcdd38b36c291b5
za747c4540d619e0286c1597e759a8ec2bdd6db0e3436e66a400020e0b61482d5aefbc0e248bb09
z521f9f165f8a5184f6b200b3ebfef968e387c4b7f697b1e287442c55d54f5e7d1db9c78d886ff5
z130b9fbdc6487d7255a2620b74396bda7e7c87669cb9d7cd1fb9fa884a3fed4de6aea77598abbc
z5e6c7c9633b55db1bc8beff4832869af59f10cedda898a3e0434c1785521a1b3ebeb108ca692eb
z8655e76bc1982669281e364285135d7f96b85aef2e312959c51a1c0b5fe4ac574fbac73f33ed1e
ze06b94e0a5825d55e3623659c0b8ad44d34069768551e0baa23c6b5be7064174121067de42757c
zb48c5174f2d935287c090c49e9812282cbba49f3d69ec2688c14fe0cd68f811418033085a50990
z84c5252aa28e87109a8467da7daff0341e1a51d42dad29ebaae79de59a1bd8f2c47c016b8959aa
ze0509997820ed86530d5fc165b3e104fd6af2ef39b2974b5e8f441ae9c096021bc14556013d49f
z7d9422f956af30e75f339c0aa2bd3ee681f1391ee0f100f3168df21df771829a8e90d273fe5369
zccbab2070193cf1e95cd1808f60257b6d3cda293d8bfda02e84c31726a899402d4e25002a566d5
z0000802be3403059a936ee000c3c4bed654b37dc6db19f0fcc9d66ee561ce416c68715ec9b9c7d
z8251f157e969a41f441863d9c7f67412e020717e13d2f167b4d292803815399787a06b5414fac3
zd832d218c8c05c2b6d94fd45ae8b439172276c58ccddfa00ab303506df82306a8f9fd0993b8eff
z00592185de695518fdc18a43f849c1b6be9790b885ce89778979d79d8a1f86013a7139ac3559db
zfc4bbd41f3e552be84f3be601e696ce99eea84cce522188bbff95eee84e751f2c118d9990238be
z121222f86e00027a55c37d5e7422d6e2e4725e8ca63f30c3cebea7d8d9e83f5581411b3fd9388f
z054e9a221534793bfd0fa8f67225e64cac9879ff719eb7657bcb71a2f88998e43951356fe9e5be
z523fc350ef03ca3294919605193b18a7cb33ecfd83f4315e3c820cfa118365394d47dee44d0d9c
zf746321dc57b66072ee8b937c753b3a7fa4c239c671662a7127dd59a7d88aaf40c73ece2d25d51
zac675bd41137fe0a3c0dcf2161b690ddc79c27269abf15add155824d77f68da9512e4545e1ae1f
z6be86971c6b0765627efe025707ba578eed68a0e9c311cb0eff8e4ffb913d336e188014c6a2e8d
za0a48a41b3eb30f55ff38d09f3fedfabc352911118d0e45b6bc2f33fcb4a9d40be1067c580e994
zc9b6abba612b364f0993d09f5de2825b6e9e164f10223d9089b75b2ed507a7db3e672acf93c266
z3ba8c1f3314489d5e0cc63ee0f5693e1a152848e2fb2b127f9928f33ab6ff860d8918ab491e288
z111ce6a83e93a3266a787fcbbb0daaec0f9aa3966e63174c3b62800b55326062c3474304884923
z08d8279c63d206a1da7198c581c9ff9ee2f48062f9d37e482d952de59fce0059931cf93b8e37c8
zcbf58b39c622c76bf75d48edc79ac7ca25974082958bcf8489c54e871d444695959a7f872425bb
zc606d532220b82923c929b500017c469151c9bd8b6d6571cb8cd04b286989d760a7ebb09eac597
z4a1d0a481c197612dc42c4d9fe6dd2ba88589470b6f266df8f77243b8679ee16ddabc0d924c0b5
z0d5a53514f3b256ada1ba2ccfc42877be1ea44267bbffe8925c7892be3308e01c317db9a429785
zdd799c3b12b545bcb797a3292387ad6dedfb7545bb6c7f52f135176bbc11adddae5da79e4aa7d1
z033524b966bc7920a60ee75616b4e4bfcf472fd28b336245879b5553a97c73e0a4fac2c8017210
ze12d55e659486a6b0a67568f362c05baa79fe4346bf3c1a56597cf8a1d119290edcd337409040e
zf93cbf68aa52ffcf0e61e8fc2d20e19e1d18b3bd40ece9377fe4480108f1d1a393cff2b02c5a7b
z05ab8ea8b59136b9eb94476f7a7936f4f2c6db65aeb9c564963975b678c4024a903180cdde1794
z959816d5e029ce92ea7ca7a8f8ddf149ecd41100b76ea2adcdecc8f6cc2e70d3b64a71320e0afe
z1809fe4575d262f7a5f06733e84efc6daf750b4d80078ed271d2ded1634237f7c173438fb597c9
zf378e95175bb9153d40b0b3aa254373b42cc466e9461fd7f30575e90d71319a5b4e49bbda826ad
zf63c7b9f6970de8a701ed8cb82c296ad3477417399b07b3c8dd3e0ece06683b06ca1d851fa3ba6
zc35052a4a4c78eabcac01106f7ce1df4ff0803de01ba38145699fbc558fb0f4b5f37dacede377e
zc87edfbe05d2acccdc43280f2c9eac216892204b7fd7934e6a74dff6a74c8265277ed678da9132
z343856a7066e481e477bd65e8b8a7550080e568232c880b2b78b62d6c1d32af8c1f2146dd6e9b3
z7fd7aeca028f58f5ec8d8445ba612564a57ce7f627440132e047420737b60825fc0611ae4b2913
zf905f8173edeef67b45accfd1df16429e35df317856baab240f3d46147f1184e8b1b1f0aeb9802
z8da5e804be707ddcb0787aaf69fbd3eb339d220a31885e52520ea2ba6d9c87546a075c040afc8c
z31b1ec7d4d1db3e080e2c2a6be4e12f4f61defed22debb934b944625c249d1046ecc02bdd4be72
zc43d2bb6242a8f3ccfb729c93c09dcbb5e340417c8cda30a2f263fc4db9158c4d6c7b34807380f
z7638d27f7102a4c9558ce077fe52bbd915023c74d123af35050cf01ff23fbb8c488f5bae9edfb5
zfac47058d2addf18b3ba4affdd076cfa42f3a6a47b23fc37f353fc1f3678b25ed215bef5562afe
z7ff9d8ae3ad582aa2f51652c23b38c655077a0420e3c8411d9f55d86ffd845419902f19c9b0a43
z79e4263b5f285fd50c24d3446f1de71245cf70e2f6c571f3b3f2823e4a43c574de6afe1916b4fb
z7e8987bb7cb0fe87c983ab98a01275f00f544687018ae755954deecb7fe0f65664bc2a66c68b05
zdc084dbb7ec112ae8fadc1199f0eee4f82df2372b576dbe4c6967d5aec37dfc538c1107af6c92c
z5047f5d9603c0904126b01272328988ae0d2410c22054a52aa9731fc0019f1ba7f23e80abfbcd9
z90c164a6c29e21d3e075b823fdeed4da4299d2de5859eb885a817486f944a3a1bcd7d394b4c9c0
z7fd21cfdea7bec87ca809906f7410ff8f65a71f695072aabc099bec50146841bb7a21ac512ed15
z9d7103e574546519561d8ef2ea5bb0ccea17f6d42bea38a3d8459229252823454ebec156ae5412
z6c4c7947c5ac89bc8731f7ae8910889a1a3fb19a2509115e15b0f132f9ed8720f8b9dc604b936b
z0615c2f72c93aaf95e51c91305e4d0e9a4cefb1a34d44448757c2d4d6fe1ce707ed52d4428025d
z7e1408c5ba1281e01cf507869560ef3f72b8322e53a8c91cdc4f08387b96902eceadc580e620fe
z4337c5713d9c48d5dd8c09f282301504066f956ef9d98a0da560d28dc94f9a3e511248699c257c
z04ed5d528a4b047c19639ea1c5b10434b52cb1913ea2f0a8c06f564d520d9fcdb11dde71b6c4ca
z85394e2cc9d0acccfbd40c07eefdb95b8cda6f03239760a7579794388b330cd6d7e0fb2d6d5ba8
z80994f92135ca7f73e53b461ea94ed5cf93543a8d242a632e15e336ca892fd9e8d5349a2ec2291
z1ee9dbcc8097a4149c255c98f28ede616087dc9d195f5d93c7962f474a1695bd3b75d1cc9daf19
za730a5b09d34d023b9945dbb016b2979babbc64fedc70737b466f4e23724d72aca5adbb4be9419
z350f69708571a37f8d5396949b18e4939657ae6941cd1dc4cf19237dd135ac4c27fde28bd89928
z8ef6d2ed602e890e83e4cd21fc84d6d4a564c6c262af72198f08349e4e6d67b76f43958d9b3b02
z59fdd2fc6b83a9f8a890167d12543f6f1ef66b959099107fc0818695ef5a906439e8f5d642dff3
z96af129b91c19ce229715ab48f79d3502b0098af5028f6d57bb027798376616170647fdc125716
z108824931295b1afe8578eb537ae252d6e8dc053f4ffaa94577ed5a3abf45b57ea0a13cbde7816
z36e3f89f43b7267b7373728f91533b1516df01fc09fcdc10a8f10c2e50bc1fc52b9635e7ce9a3c
ze2d538f0cc807c00742b0ca784517ecfc033cdcf03798d6850dee705238a1f4a590ef1a6e9ae32
z022a92dcce3ea9bb99fc517188c6f4788762c7aefa139e2f86cf8a05550268728f06cc6f8ccbf7
z738b375b8ea0fd55b1cbb14188ad30815dd71fe6750e77b1867f569e10a53c1a97201b584100b2
zeceb054d35a493317263dcb66070afee53401df99b860f200e4a21899aaa410474800ce12e7770
zb7dbc38d7506cd5066a61152f05bf2e50b128a18aefe9a12e211928594e1678611c16080c35f77
zaa8f5616e7a25a80040a37113145c98b11819621cec6e4b00d6da67b4e9be1aabac5dd395db95d
zb56a9bcb1b98380e0415c4efae4bd4fdb142c6ef03780896e4dff0262f264e990ec2aab2500542
zdf5f5b85a9978f93ccc140e55f78ae319c90709913a6f4c1c7aa5e20d0938b7dbc2b55ba0e3a97
z5b5e8d913b459b23e686a31c999fde33f5fe8267549616db3a121a1e9f2af4297c2d6a403d0c84
z1fba38154ba47dac1d773d88037d78b93c132d0adcfeb526c28a1ce2d210477fa670f5dc198b19
zced6d7ae2be24efb9af0516495b72f6e658197259fffccf2e00ba0dd29118fa9e07cf785fbd34b
z506aff5d501c7c227889337140fb898fb852a998cc55937e3e24e2a0ab1c8ea0143b3a7254b9e3
ze51e47db2435deebfe9545c74809f45c6257f684c6fd902bb2ceba36e0ad2b072ab13052031184
z124c55a21df0fb48619e4117f2c08215f278496a2d9e3bee228f1635245742b69e3ae2f3b6aefd
zac8ab65a1313c39ee5654a06cdad499b0a3ff88a880e18dd1fe0a4f53c491bd4a8c551ce512163
zbf0f8490b127a03ec7c5773801f56438f608a226edd16abcf7fc6a01a2ede270b56c294ffb7210
zdb84c63fccf59fb2d28b65d7a6d0c71ef9b2a731decaac9f4f53f14bc4d0ef1ae08f301eca5f90
z6d96255a8766341be430b242308370ae5cddb270b444700b668e8696fb0e97863e9e9041a518d6
z4312052f9f113dc541f1e1c2ace36d567c66de450f48b8a4e11ea491a460d4e19989ae7a4ab19c
zcf844126d057fcc5f4eaec36ffc976fc9d6062a507809629e2186f21f694218a63c6ccc2de3df9
z781d92719fb71ed87b9b3f97445f335ea0e7a2365ce9ebdba8ccb033a464407404d8f78d6cecc4
z561a65f6d9360d75f55eca6ba119b72eb41c9d0fe22ee2b6c8842a64df89c71712c825851cccea
z88e39a69d792aa4863693099eb36860e286fe1c43e0982aa6d4309267ae0a2d3122ec1d2d11504
z8ca83ed09b40b2fd774bdebbcbc851a4a1748112d05b2ec6806d6fba10d4851a3a0d8adf251687
z92e1a51a039a211818afa46f0d3d56859ff8e820d3bf6abb76aea4c718250a5df5b1abcc2edc61
z86fa1e5a8f95477b77510f2711df990a1b32146d20f8619bb0cc5fe98d071ae294215f6a8105ce
z79ad80dccf7616ac2e26dfa220724c96b33a6105b895d749272d8b347001045ad24aed4391bf1a
z1172a8c7942372b8e4e2809cac560fa17601ae0efbaa757ef9a0a0969bb44f978f12cbf928067f
zb52c3b374d46ef8bf5b50d2e4b4e2321c2fc8c800d851ee059ab80ae5c902c847d5d610b14f3b8
zfab6664a7636713e53d4094412cf196bd8c54280866fec7651828d9dbd3a9fcf18adb67d686a7c
zd933910da840dc698cb791d2b38451d713325bf633d1b498f518f999cc5f89583d8f8dcf0b72a7
z5596d0629fbe4c5bc033901a724a22299a67d9a3553f0de7cb7444d7b8e8563658a837ec25dfdf
zda064b04b17dac2e1d70c2c5b1531fd445cbc2fa2da46371479326731f745ebabf222eeac3fb3f
z47151e3ee215889fe3ec89af4efd88d42ac87582651355e85d01bc1fd15579d4992222a345c8f8
ze4cfddec82f455077d8fea70fe991067425e57c040aa308d68799875b78ae3ea9d5cd1da3bf6d2
zd0fde7badce287d1c7701b2897398eeceb4c8dfeef48d4d4d85e9dbf24ec715f42f8131c9c78f9
z2e9479069594bc22539f2be8f77edf479e623a1f7b34336f5f78c147f7c695bad5d635e3dc4b54
z6efc8ace2322a69c3dcf1d5cd56806715f31b9b3d2071c629628ed77fa9b9b072447888e7127ad
z578e074d22226b93ec3a710112015dd60f1d1238677c758325e1b007136567dff1cf997edc7445
zf5a2eed6002492021cba2c6805b5b40efd4c275b517b818d1e3740b6d87f9a34e7ebaed0434175
zb7fd4a32cf42f0d7152633801d4c9deca11d3d76033ffad9f3debd82a1140c9f0be778f1b5a8dd
z7d262b2a4d5593e2572b818b2cd734ef7a20ada7985a7b7cd90aadc6e2caf327b6ca2fcc71cb6b
z6a24d6333e92be0a9f01882c5deef170ab21d73645ae98083a9f32f9eea9831c5ea59fca38dba0
z6a0ac45a6fadcbbd362088c0f28e69b5c20adc8cd1f5aae20d9d926f8f6002098d8cb33d72e2b1
z896ed8abe1c5495dbccfceea5ccfe0b9e67e7ea14acb6ce9b703a1e04b9c0cd2487bdca2c8ebf6
z87f5dae96286cc3fc9612212b44ce08ff35afef73046f5d826d5b01bb0fc31efe8754392987e4c
z8bc5282775723b5dc995ed4464c149601cb2124d4b4268c23a1f4ff105fcbb318ebfe74bb5b1d7
z9599611258d005b24aa54c4c5172ca275933cf705086e675acdccd170093c88b3fbbeae8854ca5
z061bb0b27aad89b6387d3ef94c8de71f3ef148dd53b83ac667154f2ff0ce6a36e234b32df9ccea
zc8b0905ab7c619b9875bb96ca77e97d0852eef35d098bdcb23bd8ed9f4d7509ab4496811473d7f
zef79bb9bfb49d570a09f9d9b89a4690d95eaa324a7132b5bd7cad252afb67983984ff6109a42d0
z6f89fce458e62b71a963ddca133fe445e3e27a6f3c552bce7b049dd71913bbe765c4a62fa23de8
z41676b85c27097f6c634c73d11e316668484ec540963c2129f33f16bc48e8b69468c92a1e2a018
zf516eb0c3a1e003f08e9aac0f3808c56633d1998c71d54bbe0743efde18bd14f2accd00ff39ac3
zc43cbd80a7faf1c011292670ad0a96541f10c8acb21c81dc0b81bcdeba1fe19e67d9a70f35f1d3
z6bef0f2d2315ea9a8c8f88f3119df60015687d1a2b9848824d210c85cc480d20b97d5f50592481
z580c20cc2fe917a7109c1c63e1e52ed334161dcef16f6570dad4ad3f28555f0be3a99498a1cff4
z2f4a0b1d9f27c284c64f5d65f769f9976486e9ed91d5894e5096b5552442d3963ef48ebf86c2d7
z291bd2e3feb5515b79131a49b1fc7317cfe52834b28ad3b3176eeb74c87883d3c6f5647c80f018
z437cf2cbbe35f7e3db2d05f234a2c5841e0bf28f95c158733f896e0bc65d3b61739bc880c7b60b
z4d8a72082f764b9c7b91dd4338a7590d41e3d66d4a79865891914613266c24e99179820a62b909
z48b20cf2c715ea7dec2cfebbdf9a371d0b4aa2b073930bc33c8b403b238785a100becd52e18f14
z6f19c8509ce063dbc1b2739399bfc9e4cd6593bbcaca2ab5f3c4eb3abf7f4f2e17060a159b4fe8
za7c89b8c2fac56444a1b8c79dfaa5027b49d9420f0ba791ab6bd2d7777f08bd0950a4c6801c794
z7c9e1d417267eebaf809ca4b57b8dfb3db2c04a1e953c2c9dc789ed96b5760c70edd18f7570463
z324729363c04757551bce5c42284aa072b73b9a57b893848bb76c3ff7ee305adc82d2e66ddaac1
z058da33a070b391f36a85c1036417789fc535cf867bd6e62b167101de8b9b3504cef81b9d6e062
z3c923cd46e53ec171c9c8d1f585f918a3ce98b6c0d2b6d37b45f5679ccb0c67e4040857cf680f9
za6c60dd93df6c4370a0379721e9950244448a8840b6ac90dae21c3428d2a7652c0bfd7143ab36d
z1e079f42b474efcf7a75a7f5ed2db6a4cd97d9d0bb4cf3e7bb22532a4b18ffa71a5fc9ba880571
z7f63b0539a5912ab940f25d857bfb961607f2ae68d41caba00cf38a5fd0e1e3557d0fc7c862304
z9f46c11fb5c949de060abf02ff0d05e2777f77d240c53d571cca5e7ff534cd6afc960bc2da1fd3
zf9e0c9658ae22ed2fde1609c7c98312dcb7d852c919d68a7f6f872567219792a0da48b74218a6e
zafd8743a92ef7e870f62963bd1764ad13273c1e4e6a182efa219b5027f77a68ec143c856b73557
zfd192a32728b109e6a48d3d4b9a0633384683a875258638eaec56ebc35be09ce0e7d3797905199
za15ae3fa04d69c2f4021286630406b6d85ef1c3f5c2b89255fdddbc2f7bbc36050c3cd16739a38
z37fa3844b305d917a046198f7b4a8cc513b186b57c00ad2bf60591871584be0eee5e71687b30f2
zef86e21734168239f5f032c665c35a4c501bff9d660fb9ea225fc2f8ddd6b4ea5853d3be00bf3c
zff022a2dda1e4c609efe63ea72c3d762b69e5d466d063251c61d103e7d09fcf8404e7d868c2da6
zbcaea0bc0b244ea7925d41e4ca3c1fb8b18f0f23549ba070e73ab7c241755b8081ba0e05ede37c
z8924d85db9afc241f8930cd40fec6b0ce2f31b1796e6139be33a5ba2935ec53cfd7861c9169c0f
z9c2af6b1d9edb4d7ca3a9a5bcd95f64da010dd81ae13e700e081906d10605639a9136f2e8eba4b
z25ab557be5a04d31acb436fb9a40b94fa961f3861f0f9b212e6944bb463ef1913263311a1ec671
z06848feac8ca50fb55ff96a43cf26f179a826bf05c873a9f57b292828ce2b347546d3343180060
z9eacff4d153b0cba6d4f45370d5c01cb3adedd1d97ed93e5d9b349d27d4bf34c2cf56f3f1906c4
z54f03c31fdadc229209ffad81c63be7ef93013ece758d9c56e60cb1d76a2eff630d4f5c8267481
z98c58c48f44a2f96afde60b00098f6e7ee6963bb7bd8387300b006c7191982e38244dbd52c392a
z0161cab39ebaac5c747e4bbeefb2176d70cdeb41f5f2d3de19fe03f3f2d3e9e59d32c8c4966a98
zab3aad4338a4f0ee293fda14ad8edb6b499fd90349e862c67e7d3a0397dbb0390afc5111a389da
zd9319952c734f1b58de555f8ea2ad3151184dc1c9de35ec866910f34a110b361dc74cd4608ac5d
z0eba4d1073a7cca5ead45fe624c4b2bc18d1f9eb2071cd0ebfde7079a6badf251dae39362772af
z7b183a8adf1224a0dd3083bbb9d174402c22330aff0809474b347964aee736bd3e1a6c8eeb3222
z07a82115562f29fbbf1a88985a99102eed10c074f57ef0e5e2cc7a07e9f80a0e43aa45c0aceec9
z723030674851114a325d895538b02e324754646f9bf68533747b5db7694d8bdfd59061a20b739d
z1f32d46b32b93d4c79c683ec4863da330e9a7a7677bc0c6e07677aed5d7a751b93b178d3cb5619
z54529a80167f86fcdd979ba04ad0ca698e52401f2e7c958892eb48ee86b95f4afaa98777358916
z39216e43881e80db12018e59ea23e7d499a55f85500fc9c1296ed915fc204c9b4df187f87ddb39
z8c4b5e664968cead03e89d4336f091b7125730ebee461d1a251ed76a557f5e01b4569f20f2c638
zcdce88fdb68da6af02f891da04755ad8ea9a530906a1c911068b5b68118388f0a60bbc34c4a0f0
zd3cf626ea48b73662e450576a9a19b45b758000f11d0429046f05fdc39f67d993ad7cb8ccfbc16
z0e4da3ccdbcb5d33f6998cb741afda09c1949262a87c36e08b23b68197ff41b57a7600e187ced0
zcfc0fa8e3d2a339d3c0fec6052c0bbff7978dee90f1575f573e136bb6ff2c44c332f0b5b30d166
z1d4e6dcb77d368298a62fd4f161f7957dd76376e025b5de9cc97663dbd6a026c6bb77ace70abac
z26cc8613b60784acf4f6a5327d32ce81193d736eaec521a694e43110491be2e06f4fe8bb7a40b8
zb0212ebee3f332d00de9768073021325cad44d239748be000397433a757287883f5c0e84ac9548
zfb9fa0e516e80873b03955686e3e7d1f5dce2b02b3ca95bcd98106fef2add3b6cfe8e9d3f400be
zd6e4334104fba64b317932c28048d81c054f81ee07ed624905f4e96dc1ec22b850e1670237c3fe
zfa0a3f76e38d7a53ec708c05a1c846876e2bfbb34fe2951deb5e4a15c94f7d718fbfd0ca00c4f1
zbdec651b71cd28c62c48a53018937b9f663468183c91709a7f5428ed2dbc8e4dd3512e44014ae6
zfb966cfb45d646720a9e3b54e0f1ec7810e33302ccfc8a792a581ff9059b239e052625f5fa4491
zed35a0b45575d33ec1b9eb8d8684fea8a4124f6e7b87eff61b29cceae958fdd848bd86b360ca66
z37400f9cc954a6dfa64094f40bc42344e73b2b81e2af593cdc3c83b6fd4fbf3e9ecc5b59b2eefb
zbc99af33232fc8511639ffb3c4567b98e86f0e0c2440a90ab8c044086f9255ba34f621c62d205b
z671cd27a0de33b4cd95eecd39c5260e95a8512173c954ca30f3cc544e876542e3dda19f53ec5c6
z532c7ccce0929a896d103d5561577f70da235b1f74c5b9eff2ff24d5761730ace1662f2e9d547a
z3212a77fff356ef17f50d34a1a5a1e16b52e667f9d3264bf23bfcadb2d8343be7ea788432c69e3
z747283468ab2efb7642bf8c717604f86854d8c6464d229e8777a606a18217e95c2ebebff178403
z742a3923640cdb84b7df06bf8a71da4e15924784adcb9c6b20d8683d5648d06fc99bc4c07b0639
z8c2bf1e4ae0b1534ab483af8262d5b9699423bc7f79541aaafaed0c26a0d6ddd01ef047d0bacbe
zbf198fc05de43d400cba6aab09403ffea7fffd19fa1aea579eeb36e7552133c1a17846a13f21c0
z5f298e79d0c368ce093d8acdc716681b6929f03684042adfe3e70fdabb0e6189a00e89c04e482b
z5eb6332e6138d14d26d9e1eac27fa2b45768026f928fcd4e92f79f2331417a9b918ceb1e438e46
z927e0c2ca3bcdc7178f091363d9194fd6182d7f720be26ef563b568414cd6a2d50e38d43a6f12e
z0d21f05f842e06a0702a8eb26b3b7c7556e69439598af39f7657d246d98aa8fe0a3a81a1cf60bc
ze1e584ad24a06f3140c2b752237be9007eaf11eb1a309d2939c655d98745024df49eb7be13e468
z9def2bd571ccfe06f875c662bf473da00ac59686c0622347a602a77e3bf0f1cfcdf7e145895dd8
z9efe5e2f484a8526aed3a6e5f6312b58843e972195aaec6b29c23275c6b7e745fad86198faaee9
zc4eae51d6b2fe9ae1b2accaf2b97e82e1b74647c7468f521b88e77a18efd190efa4b4ec51f3313
zd9d6c195fabe2ae2df8e59f5ccbf14fbd0b0c719827e0b6225b290efd51c6c8295b44cda1fc6fb
zc7dc56fea480185d4fdbc4c242900dbd5ad72e05c08943c28baf4dd3abeddc6f10f04007283764
z4770803a9878651721caf70944e50dcf5a99daa1055f34e70e60aa03a55d0bb825339656738d0b
ze468bb8815100ccc53f2d9a8a422e3d18615de23b0ef008a7bdcd18a78d3c23c6e577d35572116
ze1d05e608dcf9e2a68c88a7de863c31293c3d29f6b08923b70bdf3fa6badff3f5965f053bab551
z8f28c51ced9c0dc19e9f8596b4ebb39ec29602b89258d4e89873eb4b840fb091be5d763c3fa19a
z9623775018fb1882f936b14daf053e7c41dd649d5e8c2f4055dcea08e210be872a74844852aa25
z83285c4f8ae069b2f033986ae566129f77fc91473e11a6460c18aabde8688d4d9490e7deae431b
z1fb7d21f9ddea17553b863bec5ec0d0d8e1a467acf211134dee97f4eaa0e0ba46c8eb49555cfe6
z9a93ff9eb2cd89e6c788da72e42711b080b3e3c7313ddccc51ba2f6ef71db872831699093a3690
z4097aba21a613ac0fb1d9b56a14c3b4142397f9f04580d8e9203c521e1c11a962f71e071fe9904
ze4cf71d0ed579205740c88151b7c53b9ebc35431be7c7e03adc9ccaafdf882e4aa0e3bbc0aa8ae
z1f9c6777de23dddcac4f2baa6851aced8dac8baa57b12ef9ae6e15f3246ec64d8f72e59c8b2892
zc0f16497673825612fed0a1a79c83c393b0f6135bef2749ae5d196874f90955871879098c271ca
z5782c52d085a47022241a62512429c6873dfb7d171c33ae527451c3bde9be764073697fa856e17
z0eeba2ac00b7d2558f3dd72c4549edbbe849a0239d7c03e4321e64db9ffad3de7d0611203e6ccb
z23db20b8c03948266625c3a815a3589991717e6b0cc5f673d01c59a0cdeb3f13850ae2125636aa
z5552d9ffb7e532823e97656c4b11a747050283c05a8e653014119b998dd53969e524d9892d7671
z905bc0972bdd93a72602506a181eea6b43ce112daf6c7cbcc709249aeabe3f310d767173755e47
zc8a55572739391be547ccc1cfbe9c8f26eaa2b235c24e0ed7d51301329096b541bea03c8b4f84d
zd2d9a30ba69afeba5d433a50966bf63035531dd1ed28e494876911b2aaa2ced8c5b1d5b5ca61bd
z62787b3d1a88d7a9f42681831b0ecfe0b2b573cd67302915a6aa8f3fff75aff524626a80c8f0ae
z1ad58aa669ed96351e4f3cea2c549853c9a0cfd702b32b582e704448d37dd40b1b9a0f16854427
zd83a88b4d4f1ce0ed302835464cff255ae12a9767af9aaec122d7caeb8daac82b6c3ebc0d13d00
z66bfa8e1839ee9611e647033b2218d6d7950c2e0f436828ccf299b484a263fc40aa99e05ead707
zdf7709625df0b18ed608676f375216276873adec2f1fe19108b600211d2c2483b28e8c00984abd
z479148acd62418d1220bc0527b3e541745cf55276191d446bdeec45dbb6d74ee9995a023f4b53e
z485619da211d24f82d377338923c2537a8947d862f8dc2f7ff0bf15d49aeef439bb87cd95ae335
z3e266c29100e5daf7d4b05a8df79afb77941b3d3a4ae7accd73664d7885b9ecaf4aa8887ac4519
zf3c39ffdb115e7f737792f7c204e2cfa5ffdae9c4e607d73e98859fcc9dbe9863364e070469c3a
z30739fe8eebbc3e6cadf4a83c89c808357cb88ae8088c04a3033bff32f1eb5d08f1da855601602
z9d0b4919554616778c56477f51964555913ba7a8084355d1218a3c860451f8e6bf61a700e35233
zb9979906d23aeb582ca234dff61cbe5ad1312c40ae64f23d05719095af8f1aed6b15e558e245ca
z113e06ef18adb224d47144a8b071c01e69bbcea8a51fca43797047b10e9e332e17ea9e7aa28531
zeac757494d623225c645df19617f494358aeb8bd43a6aac3375123ccc80db791a52f2b3ad22171
z85b6cb25e3be9dc7fb2bb3258cf0d494f473f82d42a32e6cdad400574ba6d83d71eec2c00f674d
z585008cbec30a5571a2e091bf61923b8de65152502e8be03feaf3379264760d1435cf5f32a27f8
z099d37c002c1aa9b836e8208e99db70f7d4c34e52641e33c16a4424986fe3c0e6f403f2fdb2b24
z135d3c4292ec6db6ed76e042f23c74b60847bc29ba34c597381d97c05bdf60bfafa09d20e931ab
z9fb0c688369f277b3d92c573f5367c91873642265df73325facdca96f93e5f863579b42954184c
z517134aa09266ffde84a8bde84be42356aeef8ee16da5612a7be8adec8980b68d689f9e2c75075
z5d6872783e4415a0939b69e35866402806701b63cca844a882dc2a6da1bf3af40f89ef004aca3f
zbe86541572f89f70075467d09df6bfce6df19f437553d54112ad4421244c7c018d4a713a1d22a9
zfd51df52b28ae70a92b324376f8ac183249c25564701a2c6b246878dfeb46ca740984a7731e2f5
za0a8216cabd3b84a84af1211d830fd04fa4813fc6dee49d0c2626fe69e9b75492b88dbfd3bdcd2
zc14bf153e7b67e6397c08ca06aae006cd7ab1fa117afeeb3d8cb1a5f49fa6ddf20c0446d0f58a9
z87378a66314c32508803460c1fd247d672d90b9286be29231c0f34fbc5af9eeffb80f5e6343fd3
z9397900df43a9e1caddd3d144d81a0cb764281323ab8f19a1427346a9c7a4571afaa0a6b5fb06f
zb20f3216e3ef3caac436128c63ea2c5908d068bf7834b60bbf0a39a23cdf89f35681f3845d7fa4
zfc237ce43e84bb698c3c3dc6cd6cb4fa7e45753ffc2b70590d7ed10ec563a08293c0eb77fb294e
z6c5eee800d44a7890d7ac58af78b583867d743fef59331691b7c504fa8c27a928d320ec76f6965
za81929ffe2aa74e4fbfd430facad0a24b7e9610662ffec2818cc82fcf62882e93f19095c1e6c97
z83ab6ca6fb6de8756c277928238426b5cfb22d4f24b71668a56b354ecceb1ff0f07a7e9d2c6a21
z57f121d0ff06b85fe4976d0b1bf7bb91a8be183c94078574cad7d4427a6d53683e0bc8fe1e2a29
z95947a0806d3e063f2f8e1e388edfb3a92948a3638a946be91da272476d1c699a6ce3ff3cb3573
zfe0b11574570d9c1b73e37bfcb0acc175e44278d1572cf7dc406deed1158a35573b5afdcea58b4
z90b5c7bc71d5a58b2c0948d7c32c89cedfd8f8a9f3753fc5b4c8de1fff25577f8ac0e113640d8c
z4cccf388782eb213006e4bc95097b8d9f693d28fd73142c1b354db42856a34e1879b635e06ad29
zd5cdd7dca909c4f5ee83bc2bd7735627285848f09e3a2493ae9ecfbe44233bfa1cf8660926f318
z8ebae09f282d9551a3047ab769e251d0a256abc255199f978ffe256ab69f0475248b3afd0a3c30
z5069b010bda6956aae8ca43e868678949b30dae54f2acc8dfd28a3530ce368cbdbd43402c19033
zd5ccadc75a72fc962b745a45c9b53c96d54f0388877b164c398d7d4fe678af4e7bf951bbecc53a
zce72071fd061a1bb97420e7522c5f206985b78d4620b0e9ee47f6adf822c13a0b337ab5b38227d
z13f70296cf7addc41c5c001ba81a6c4c1b390a77ae267b2209da3625dab315accc86e6d8c97391
z9cfef2ac3be0dc35b99a9a49fce69b1deb4a7a23d9ae1fd7e78841c3ae5fcae2d49f11ab3dd33f
zb695845a9a19498f02a0f9befa822a8449f371cac5a0c8990c8bc950222074bfb31f6833d2dc7f
zbb8ac2b3b778ca6c2291c1c715f7054a8e1cc77bf3869250f0609365710af7f4690e182b245c68
zb0aee51115cf5b67644f9e217233fa8cd0eb73a66140ed9ffa51d221d028cddb76a2caa9c2ceef
z9cad6dbe5a6c2a13eda733847b375f84caa974b80d2b888fa4ef8e33ae4605e97e25d2ab0f3a2f
ze2f14ba1906640bbb1c889fa39b0fa891fb6be527583eccf3ac3d9c02dc8f85217d594bd0ca260
zfd8e09d73d4f33ad914de2200346f346383c861f50ea42f58382d216761e989b611d5b73a4ca20
z4e849b80fec8f586642dad3cf2193750f3ee54965e658455e45ba3fa29909e53280710e284bdef
zb72669f98b52d33e9a39deedbbd34dfe48a9ed4aa41e90d6fc945b8bf3808058ee5ee22baf0aeb
zce7e7743b74be7985a4698ed3ef62f75686f93d079d842a87c0505bf2aefc2f2162e524249a154
z44bd4c2e423693093a538c0ac94a64f4ee2acf7aefa16d0f5a885fd2e42c3ee89aae150fe10409
z6356ab6d4813355d81f2d9000ce1a133b7f153ea094681e75ec162611dffbb94ee2602222291ab
z0d3f43c2cffd780564d1e2867a01920d79b3d783a34b03bd618decc9609f1163e6147adf7fede3
z9d91e350e6f3c4d80ef50e186929525fa9e4ef2271b261502e68945262d95ceabc3a096160b3df
z69b1b6afe545acd423f0243ba8ec5df081a41a897e58797b4b665cad7312948f94a3e94ab788bd
ze1b56a6773b160e975bfc8e816c1b6be6eacaca35b39f9fba1b2c10a0320e5ed648cc747b809bb
zefc09f9d8d5dee60d67a3b5d405c98346c1dca028c380a7bb11763e6784a6a489f22e9c1562bf2
zb17b578a602f063f9e9ffca89144551f9391c866e2439e94b531d5adc1cce3d4b651e5b1e93a2d
z894a6ea0dad85d828490ccb19f7a0b91f4b2194584f1bea891783a4413f14549f4c5db90005b95
ze58f8b081f23509a8d02dfdfff4757062c55e77c3a1e860e8b74eec31a8aa16b03788fbb61388d
z900abb3da5da9172ca4f4cd775d4263d67bfdbdcc92b0226cfa0a9abc1873a61a611abd8bbe5c0
zaa114c95cc87c08ec033ddaa4e48d813c965740a68c5edd5394e1d049bd14b1c521ddb5c467c6f
z76dd56a30dc71ac3710940c554598a83ed88eaf0dce8c83d73c7e7510419f898809e46a16f14f2
zb420a2bca4fe81347af0ea5aa76f8a2e77423d167532c5efe1b143c792fbe05f4cac502432a0cb
z75f1e6f1ab1bd29e4ec9e9c246db96c5d978fe04535d82b71e50488ddad7c796f7b9925190e67d
z09985736551e4bea45e95a3cd1ab167520b1827a55b32ad138bd89ac7dade454b1d7dee5ad7978
z0d8481c5551a238d2deb35bdc277bfb088ade40795dd3b8f9f8fa3762af5fcf2b7d34d41ef2910
z6ee46ec524040a490611bb03e4786985c115ba15fe108eb851f8d6ed51203af35441a94c23168b
zdfcda4e7271976cbdb0397a1485d58c3063bc684bc41418004bec777670d701ef5458867839226
z76d986da48fbb51f1b000d964568e980cc7cb600ff09541ea57c86cafe74a1ef7861f325f3b972
z3b24b30e632ed3aa0d6deea8751985e0235b6fd61cdd665dcdea0d18321d255090024d5d378ebc
z61d9bb96c8ac614424bceaf4666aae114a43b07c33fe80862e59a17f5c078b08a02cd124d31764
zb5d6ca7842600b852bdba9525370d7beed40e006c65572e5f1570383383e9c76f42e847f001a9d
z1b30b14279d29a592fc7366a06aacf76873b87048c60867f52fa7e49d8403a20ac932acb444b7c
z17e159f786b0c393649a7e3856560f9d3ca787280b85d60aeef981ac5850f96ae845a6914a97c7
zf0a01e7d29ab7a0df64a96ebc186b90f07b24251ddf2da433a22cc1f50100da0ec9c086cd26fbf
zdc4deb1245b439f9d2003297b010eb609a2b3c9d7925a0d25d6886201f5b2232c928ab0857d828
zd1db8d9f97e51d4f2614f1660606ca4267cf2aaead4932887582e95b4c34b30cfd2a4eb7fdbe42
zab1ae16205d99daad80ee00dd195b5e9136c7bac1d4ddbdf5b99c499b30060142de8ea8fe093f2
z61082d8b96a8ce09d26e346d72544f8e1a27a24df47c8ae80a3121f4408e445b41e4c29585e110
za79dad30c13034e7b70f421a5c3972a6497eeaae0d49c549222782d536b692712dfa1e1a42d05e
z5ca8b7d773a280d3863d8fe44f725785164d612029f37e8f206321a5463888d7e590b843bcfc3d
zcf61390f911d40643fda6328d8a779bdaf8456233e3f34d596c799ab51460d20b401ca5b4f2330
zea37a41cb68296dc8c5ec914d9fcc5b2a4e36f62f31ec76ed4d8dd30d8a1fcf8c2b38a278b8c01
z71285d90c0f52417de1d700bb20313317ff16a809bdb21d8c2c3c015e77f40320ffb46c5496c9a
z96a1eeaa311b6226c6cb4b389b7832ab26852ab46470f6627a2a07c3e9612aee025a99ae2efbd4
z0281360df71f416b6cf3c9b77484d6615e7f46f5cab5dd2b0551885639fdd77551a528e4e5f610
zdd7ecc6dedfbbf790e7b706e65eb077cfbbced51f9f8ab0d51056a7a9ba2d85547412f466f5d83
z4025897bf9572857a3376486fe2b0e6ab4fb01ad357e36ea294da3df2cc0e7bce81679e35b33c5
zba88dbd27fd8d0f452f0f04e21c1c70b962984169ee28d2e93bfd9c2cbf8e7f4926fa393cce436
z837022fe3984fe2694ae57622e83ed4535729a3a6cbeb3fdbfb98d99188fc4bd558a3ae7f3b330
z9ad8bfc555e566c3b8a129d6e3f3b6275e3e5584459aba42e3ccc551e2bb19a88116b147996df8
z90ffc7c1cd5dc72c42da561f9699bf76d23c847b97d6f5c4b3c2d15eff7a4ef967fdaafc76f4c5
ze3e65e1d901fce85ddf922d6fb73e54ff3786861a5254ca8ed633873af05783f0361ec4ee40d4c
z08e5f51ab4259447dfe94c667ca8e2612cfd9ba913cb2ba22bda0cce49881925deba440244036a
zc7ffc533ce48dd6daad90f5a4c519958ff268669c45f81beb3f113d7bdfac6d216f3d55fbe500f
z73e9166eb55524ea06b2954051ad923c25dd58ee2dd3ef288922edb5e27de0d85084deee69fb33
z6d8f695c976617ae4783ee4f41e00051fdda546995c1f1250eb3791320306f948365e472a3de57
z80b6b415746d10439aace4f1d9848f3e693345e2856e861ed53bc7073556cb12261ecf76d8b773
z64704f6292cc7361f1fa21851f63d415fde43e84fd0d4e85ba6410b7653f271ab7e811ce3eb328
zbf546e64e5c12ad79ea4bb0f7402f4db4bcd523558d1d8dd880ff94a18e1a997698b59f84c4dae
zad6248848f84096620672b737006194e6754395912284752834ec35df32582e947f812376d1399
z631831f3215e927c0ec23e665e33b1ba855de8b899a887a21cf3d99716340ced1d83e8e668f458
z11e053f8dc26c3783e15ceaf68700bd46c3afefcc63191cd41ef8b48825ba729ef65a9fed0d0ab
ze97414e29124eb6b18f3439f207afcc6640262a70e0a1ad8bbd1efa33ad6e9606ade06f48a4d40
z040d97513a8f183f88307cdae2e445da7794666123a03f9d8068cfc0d96e293fcb7852c6a0d929
zacf998e7167de5df24b06356bf484f7c10bd2f9d48bd20d9460dc8d018ee390402f29339d49c61
z9aa6dd5e532fbcbea07d10bc4d0a602b15957c6ef5e5e6034115835eb90fb8373769104a5eac7d
zb34469d1e6f0a95174f604f6d8ca7e01fd77ce9d11956629f5bb536c12279de917cf0acff4454a
z602872d4034fdd8760c739da38d57eddce95cfa5f9082572134c88457f84961f5d92863073acda
zee586322b5dffef71857ce2f726db0f247d4b00d3f6edcc0e9659d04b2d1efcf36112868f4298d
zccc16affc90423f2ac80b571ab4e55012df51b1f29f2b0c111dfb8619afdb4256b3e48b27c5e3a
z4e0ca780579adc6f6ae83cc602a5a8f76bcef5ba85884b9e04d7702a75d02fe4341accb14f837c
zaed9c87d777f2f9e62d5a823cff82a570046a234adb3461b33523a5708ae8ff9b0dbac75852d44
z5147990f5bc861054a6182a44c029039fcc2897c0b281952749711b12d947483d41c89b179c042
z9b6ec3e27e90c864f15123d498507772a5cd8fcc028be4d7068e87d6043236ce04561a75497123
z32e11e7763fc52d8dbd1e827aba60476e0f39ebf9919d14cc470a0ef2c5958be0e411279fcb90d
z0f67b874281796a4be39fb8321b5c02623d91506a6aa547b13d70b02baad25537927c385e1c514
zbfcae258beda51fadaf204c05fb35f25ac304085458b340752f3486ebac15e18bf19da97578c57
z989891ed2407d348c0eb1e54ab378aaa4c67d1a51ed78e7034c615f76ea6e9397acb20be95df56
z6753bbdc20f344391a4d9e7320728c5f806d3d091524f9865b58f85e76676ceafe7b10e37ebd57
z1f9b9a4fda16ce7341f7c1e5a32a618a70f09a7e96d5111d8ea4e0b5b096a02a5b46b1e2d31f7b
zcbbbcd744bc7ca0e5508a237943a61c27cd42f7d0681f09467208df7f50cf6c255747f1863c94f
z009b81705d13c41541fc935c759adcd8f88d6356fabb2fc8af4bf979fe73b70e05f9912e4bdcbb
z8ad16e5ae22932a06a038e60e2bfe170b8112b110253c8bb3303c9b7d93a08c0dc51b720aca1b4
z536a4f90cd2fe0ea76261e69e4f534425f0559887fdc01c000c558f879b2f0f695326e2c1d36be
z8f82c118b84a94a174463c55201326716aad69bb6cf065e131c712686813e5fd95adef49ad68e1
zb3ee7ecb07f52ebd796949105bfd2bae11524544bc542c4f3ea586b488390889a63f764b3549b7
z5d979d28ecebd193087603fceb8c4fd3199a8c704b3f86bcb86d35ffa9879d62daf90751162d0f
zd13b29479f85afffd187fc1ad5bb03370c96db0757dfe28547823638c7edeba8af42181850c63c
z94bdf4260aa49a3006f75bfdbff140684309c3d5efd1ab3ca9954a5d834667fcc1b389bface804
z0817f3d7a3ba55a5629b6262cdc160d360dc8f9e0ad17ce283b7fd1a54c76bf23d91134ddb22c1
zb646fd807109cb31f94cfd8d1f410fdc78581691211eeb714db2f3b475c77b9277ac4907e55c00
zc6076f8835b4e71f8601ac732b086a47ac39979a38714689ae0b20ea6cb88e670e191bf75e7940
z4236c7bba62bb29b67cb37d9a5a657ea41d6e73b13332d5a020882229ddc40f41c96871ffc9cc2
za768b08b3482d895f345d1290939c47cdc6bd991f1b4135a9decfad5974ac91b49b096e4a1d4b8
z2389180ab1d1d2ae4fd527939104d376edf5a0760ac175ee71377d3918cfbc590611dffcc1e5a3
zcacd1cfe0fa41c2c8c182819cd03df898b39a57d60ea396b67ffdf0d01f19a31b498b5ab3a0178
z7c0e7cf3497b76fe32055a578ef7edb251ccecefbe69dccf1ed619b265b9aac32197b578a78b91
zffffea813d7b44e3690a3c1b15e4b1af4043d75768d6a3893dc4378d09e4f1bcbc9cf5cd9d1fa6
zcd4a929bbb5ed9c2c6728ace61b14fa7c42022ce5198a6b7df4a190f80f163ea2bdc326084fd6b
za5fae848d19c40c2df3275fe9b27392960bb24929b22e9faf49a84d657847a2b31f76a49917482
zdb45f2e5585282ff8ec5df5e1244c6de43e7b7ef1ef7492265dafa7e800e316a63d9d2d9ba2aa1
z085526819e1bd7af13eb727ff2bfe996c9fea85e5103afe51343207211db2e361a43fa0acd3467
zb13dbce83391736d45adbf3ed441807ab62063b1b805a6f10f9fe944b3275b9f7cc0fbc4eec37f
ze8400eea34ea2f5dae04fca6f015bde0d34bf28209dddbafb6e7dbc12ed817c90a4a57456753cb
zd9c963e83b10105fa6976b8aa4be0803225e2689db6920a293c6401d65e292d74a75b4f9c38229
z84215e5ff1c533ffba04b58a9821a2bf99ef8dc65cc14bfee719f40d31244221a39f79b560e11b
z49eb7a68264d3b0c720a3fcfa0a4bf66cbbde10125d980d2e0abe491734cdd9441c63e5c985bce
z79d51e1d160019b6715787bb4bd544aa7a0a1923a3738484b587d84d17c568cfd20e7677725654
z5bdfe4e0212b562d098fe2b976dc10faa27bfde5d9ee61bc4b30a7b8d52242ac8ba825bb3a86fd
z061b45ba5818e9c22e7ef791ecff2a0943b25e42df3fe484dd9e7e3a5d11743bf394db2e8c59ff
zf56a845932f494b20eb17d165ccc5440e4963d812ae81901f7adf39139846f71b387fe4a085233
z6bab1804da19af9525aacbbc18b3e0ba06973c0c43c9e9172fe212cfda2f9ad1a3ecd97687e7c4
zbb0b942799951453ea79e7601c03a9be8451c524c0f784f13e5b746241b5d03cbfc9a7f0fdc6db
z39b3526969544e03bcc1dd27d6b5560a4a9b6425d34f6c1bf14df25406ed3ffa721e878903aee4
zcca0fe4c0a9890ae61818364e66338ed7278fbab5accbb47939096f6658e90af5d32d952b9a12a
z123efed9607724371639436639af5a7380c24f123fb74efd4b1a064e0502a1b57dc6f270ad1df1
z53bffac8c6dd3d808994546e2cbbaa38af3a55275f6591c2d859bf16ce8c24c09eff18970cc9c0
z310a0d695e34dfe6362e6e612d47ac4a22033a4a1a0c1b219c44a480c8b43e4dc27ca6ff149501
z8246de9d868800b4e191805c0fcc12e561bb145a7b5ad975a88bb291818bf05a2ad482e3e12bbc
z8d60061cf384bab3544bc50d7d0973e7a1361c32d19e0c074f1fcf897b66e9f411fc63810fedde
zfa7df846b4c00bbb1a7982d245bada019f2d5826afb2f69e0f462725c7ac7a79c380b988295b79
zf86781f1e7ca4978a6a04d4eaaa286bfa099f7988ab1707a941ddcce8d062797e9426bb8e78d32
z6fe092e5e2a2168bc50db7755cd2cb293652b8ea5cf94194bb72af9dae3a27727de9d346589669
z96b9ac50b4ec37404878b860496cb4217cdefaf94bb9699f9cf7f236f49ecd1d5b1f4613d3005c
z0a17bbf6a79bfa88857f98eae95987a5cfa894bacfcbb83de8cfa5a811b672aafd004e8ee61418
z7d1f2424befd24ed66942f123ff6c6f308d1699b2f9705682478955bdb8f037f9547a98cb216ac
zb226ad7cba67d84492cd97937bc9a3c454439c86dad8228457d0128c55bc28ca778fec3091025f
zecccb8d46de49f0adaa2c22b108d4a2ed9af991bd838003eb2d2c5586556d9da4c4476595d1510
z3eb3cfd90b06eee56db1b1241258e85678cc769c28c9d717cb60dfd900183320198cb3557c58a3
zf7b6b4a9afe0dd4ca265fe8b11f95988262dbf6a35dab04e8c17567eb4c574ba8831ae194d6e72
z1f6aab9b2dcbd6793cacfe4c3df4badbbd26c283d13ff3d5184c548285e07984893704e34033bd
zad38f728f3ddaa9efcf6aa6131ea488147e19cab28d747be3f02e14547596b71177d1cdbcdb9d9
z75f3f8a1a680ff7c43ec6c1a4cacb0b16092bdf90b41bd5a020f4105c5c50aa18ce62fb25f7f2a
z734fe91720d59f25fb0d97e11547a3a1ca2e944c9ede4553b9b21acb8e62faaba7b190d7fb173f
zf6e92a56115e77c8ea34a6c14582e2a5ca16d84d40918a7d0aa167f3d03ef981520de49cd852aa
za1a4895674ea002b98ab8830e494fcebfc54e7b6bbe7afc06dd04c36769e9a6a81fcc9b828c1c4
z6a12fd4cf2c3f8bd8cf196e620c0bb3a22d70c4fbd86681a937ee8fe27b3906e0e676f716b7acc
z2755ab9360d6014f248760d82a4ccee557392880e5558309bf14a18b18a770f0089f8869cf2334
z7c1b14d4c5c0172280ecacdadbc5711505493d6eb4dbd5879bee83707f986471fdc528be21cf9e
z9250f7365d76339b71f9bf929a8a047e0869081838d19dea0c2e88e7c38375f3f3bce5de92e655
z33970c9a614597c0af94c049675fbe66ebb556e51bf7e9bbe7a0d61347a0c22dcb34a66b2beaca
z3f4c352384047da60d8195cd3a1063f3113e80c88dca338a1fedbc932209aa48228065e0322436
zb69a90e86dd963ba107b48af28ec70441ebe104064a7b04e7f7c88d7f3e3eb0a25cc61379ce2c6
z86d54e3b3d0e7e107fc9da952c2f7a490b1816feea3e34cc2726d5fef2e3439a5420bb17f27d1f
zaab54b2524fa5201aa7293c0dcce916f0fae2ae15dc64ca5ea943a771347fad420fa242985640c
z315307673a20fd8c6ba57c39282d34358abb6152294a380d066c3380b2de6ed9b04b620e65d0cb
z621e4e24bfe7885300c5a69de139bf9f754053f9b270fb8c7f4f1a038a1871e1059146981b07ae
z825cfd9d2ef33566c611334645d538797a5ef534aaba022eaa78e2b054735211b1e7eb2240c448
z0785cb752a8988cec13e5e9770ac5e986e008105000445a9f8d7fef52693f57a4736fe387bb7a9
z77b42c87c8b566d84d3a97860eaf4ad2913fb3b822ecb44d76c11decaaf232439557b4f743083e
z44b6c23ca3e3e33eaae47b9747429ca61debc94c9b02eaf376c6445ca38c189db83183244af688
z2e58b2f3c68040e93ae14c6b5392eca55ad9074ce86ca6280eb3023010afd1fc0ed89d0f4aff5d
z39165f96d3c67097d495782a105cb3aaa78fd5951e2b615e1fbc6676b437ea6a01a2e62afd1e81
zaa1e7cf8cb8f83cc858d573aff61bac2dbd5282d45bc44492b4013039837084433e1a6f5418f91
zb3bc346c836bfa47ac9065cb5b7465ff4aa6fdb64b2ba004390e1b491bf7ab0300c35d26792a3f
z5c8d55fcc24677eb8c8e20472e52d4a82af052c346b4089554b6610de182f369855ac546f4b0c2
z02cbc60f55ceb62ff77a247b7dbf8dd25a815d15229500b13719819d5016b0873b5d36054c390a
z60af4dce8fb27ebb1efdd1ed449efa2966f2ab1c1ccdbbc93f1e8e9b4a198c9564bfc03d3bf310
zf18d7a353f60eeb63239f7222b3becb3dbce1fa17c5c1dc76625de6ed029e5fcddc04b4d4d076f
z1a0167d5b2451fcabf9ea26a7d4016f05d2ef7f69e848f6fa80eceb91c6c16fb12f4bdc5b9d536
z124f073a6553049cd73f45390d23e60e6b522575fbe92b9edcdc1b5cbe66f772900d663874a414
z9979cc52020e3727936888d954ee022ecb4c5a1c5c919f8bb1cbc880585914f0db8d1e7e9cd79b
zb8b46c458a3aeaee1d408c7d8f813a03cc3c050eff6218d2aedcb54d5e3bf1226523b70e64a965
zad0001061ad9c044de0d8e1741f60b0ba6190f6b49ef8a7dcc9e162c7338019e14481104790287
z4c3bd474fa836fd81907da52538750cd52cbd4bafcc8a741d455ad5e3d87b4246d80c803b9af73
z07f9d82f3aa737bbe7e08739b660dc8451fc6e81594545620c499cbf8a3db362b4f75d938f9d7f
z74c8e1bb103e4b6121834e9a17a41ac9890695ce26ac838c6298e049ecb716f6d1f00b13114309
z5aa6ed594ea5cb4333d76c0f0aaaa861b9e3740960d1d0419794a490da3bff540d6b71fd424a89
zd0a17ffd24ead36a6b5ac4784caa8d092c3a5c20733ae02d0f17087b7a4a80b3a3db525ac0dc17
z0d7a3230b05d04720fadd4e4159786deff2682ec0e8d28d12974f89b463c5ffb15dfc64d7833db
z1ecbb8ef32b558c207e552438efe6668f8024c95a59c04088870d4a6a1de18089d2a61043e543a
za9ea0386c87fb4919786978bac61d71e2273cce87f0346b52e75ada45691231159e2b3d4702996
z881182c3130f938cab4f8752ffc78fce99bafea229e91724afe8ec1d68ec5d97bbcc846eda164a
z7f75d01a6fafff937dc6a06ca04af7445f97bccd90c1d18316f4a0dfe9f8b913403297e62f2c61
zc92a300702bb4fecaf01b22c981c8851b98385d00aaa7c1dbdd5fbad5299b2f1083a37611ced3e
z20f19f2b0025c5217078fc8322737e4081701d7452366da16de574f7df166d41f70cf9112c59d5
z7e8ad57bee5d8c7659be72db6bcce9666178b874d1d6383d147e1727a69935c4056ec924905eb4
zba14ebfb3718198bbe00de19eb7a0b74146299b276e62803e61df3a9d67886e306a4402434cf91
z5da4752ed5e6f88cfa84642b36713598f1d5a2ff68984a83988cfd68a59b4230cfa99f9b444bb8
zbef2fbbd5017f6f9b3f81e3eefc0e7fde62b927ba36c71565c9d7258230f5b39fa9c1f3f37491c
z931663bb4b8a33f0acf0f2aa89033ae7919788d612dffa6f469354f857752a280f37168afc0d05
zc2997d4ec1c688d29663511228ff987512360a30c62e4192ee6e2b152b58941d0c003e98919a32
zab30525260489a232e68228db1ceb7146c1964bcaf2cd23b80796997eca8b00c77deafe2284c8f
z6bb6381071d86f6fca62138bc3f07683308fbce77544cf402dfe7885d50bcf0ed563d0733cab01
zd689d8e06cf44131192d5e2f384cfa53cbc4452e7c316a5f4af5c0f6570194766f659c51346807
z7498ea6539e7fa6f76b8d43f51277438aed5cf055e1f241e29f2c89bbdb20ba87d24529b793678
z62b87ea8c0d34e26a8be0bd4d19e3a9bbfa03b4e20a167353d84fd0d00ca1b2e7570d412d9a22e
zd70fb805c12f5e9a703502aaf95bec742da0212e1786b9a39cf5d11adb22982ed6dd1a2e5f0e00
z86d8a91cd72ee140a2202f1d3ab2b47cef49ed40d38fdb7557426cac1bff49d16fed30d250774e
z9835e9184ef7439372ce6a00d5558c18f938bcd079a0a28ee924f7ef4e7659e5bdb9fa6f6b7b6d
z6839390f696391e987cc87c810a800fa425c01b55dd297a01ae550fc154e2882c4daa5fdf8b7dc
z673bf39e29c5d5d0e9d6d5648eea0d7d5676ac561031c8d81e72f33b2a87153ede2b99fc115f8c
z0ce397a1fc75b92f596e69c34e16b528a8241febf37d9e4573057d88a42639afd96c26efdafd92
z7df1193deca852debe3c80e8df4cb90939c1413fbdf208aa5a869b921342d0050ef65c242eaf6a
z381a2a123df8633b97afc79217a1bb8905959ec9f504e0c4b96f527753174f84cf734a87430cbc
zd1f47a9633832ac2bca8f0bc0854ffffda76c6d7e7df5eaf4f80576a0f72a25564d782505cb2d3
z9836c974c717d329a2614fb3925e6bdfea806a1197f98ba38e6a94ba3be46fa6fcd59b90e3091b
z45a1f0413f4363e1206fa52f6469e94d55fb1aef1e0fbdf1757567b3fab8ba9ae8f1154a8b2ca3
zcb40a0847370c408815ff3438bad52c03fa3fa40e553403dbce5a92d1962488318b1e3e2fedb61
z96ee664f1dd89f371dd037e0243faf353c0d7cb3608999f6f6df38fd67ae2d8b897a7fb09ee39d
z361b829ba79e0fcb351ef8a97b97ab750d0108d44a4d581aad3753f0dc7ba28eecdc0f13520aaf
zcf43bf1521aaab3717c2c8e112bf7b0512604a8a50604871e2e3746ac68d0a88d20465d1e0b0b7
zc88d4f1db258d97f548a975eb21793994cd301440404f09c7c11a237615724e7cc3687a3027d8e
z9963745437a510d28c78e850860e4775801bc6b76c2af6ae13717117822426fa6ba0cab41a9e56
z1cd2acb8f462e4557ab341e7faa153e63cc5b6740c53cdd92e31a7333517adb1bc2158c3f0afbf
ze63de3e1d7fbc398a636e7d344abc9618225979197794cd9d1e5a825620c48237087f7d894b31d
zb5646fc3392f9e2d8f5f74252758bb668393ee7696b7e15e772f4fa27533b43e5ec341964dce40
za9884765df5f0681a31b8a3aa2cc5c534d3133aebdf93cc337a23cd85fc612b5775aaaf25ea93d
zc71bc3d1b19dca9997df2c16c3c4ec1d64359926b543a345f7f8018343f3318dd422ae8d44dbfa
z006ef8839bf2f5b8eb4edf0420256ede9349c90e981b2ed912cef0c7b6276cd15f6c042efe519a
z11be726f54ff0616f5a1f866bd4eba7f96d4015c82cc7fce2751659ce81fe9c291c8fca7c3e989
zac10ded06572d0dad4adb62b784924a11562a5066612b682ea5e79004700883cea030866f2ec1c
zcb481b64aa71e91f9a4d19e130cb64635d04fd7b09c8d7bc9f0f4e877ee2149a43cd04a187b8c0
z56ff532cb62b245d7433494017fac9b29c150c8ff2013159ab050fc43c28278677885f3e1915a6
z66cf637a790867838d5734778848d90194c3aeab61fbeb5ee1952a0618ea10b195646bdbdb7005
zd9aed6ff5e63d8f9dbf94e6bdf775950557d5885192aea2a0c4843482debd1d18dcfc984bbff75
zf67935aa6a4cea7eb653b9bd9156ce57f9480d1f5f27e1433e6b8a9aeebc7225f495903353205c
z254ca32ec5243c59e571ef9c400cbbf4c4088d80d85202f96734d6f46272794b29a69018d1e9f8
z06c15ac580385777ee175eb76d1bbea30aa0b2794a460f45acf499b4fd225fd3c3ebe471c4fd71
z37f2ae2909e6b1a166a12701fed35ba90ab404dd68ed83c373ff177c3ec63de177ad5b56d998ce
z402cf9fd2c93015c2b1ccd3db5fbff8ee94ceefee39f4bfad8d7caab777b56dc803edb607ebc85
z61be37c199dd839cf9141e36f6aaf5a61892c7e487cf2edebb27ea4fcd5ad1df49ed36d9fde03c
zcebd949824f82f18cdd84f88ce14967b68e7530d3f340477741c978e5a946a53db5f982cc7724d
z34f0e6773faf10c236748aa53bea5036a04602b50b169c36c1d3e244db632aef8a39d8ef3afd98
zd3a4016ebb308e71f5f64a456fb11458fe31cc754b6e1b66f600150339b2d682181d47aaf44260
z93d5f20de02fac57c64b885463bbd0f349b5535a13fd026fbafbd4682fee531e892279b2bc426c
z46c227f2b11bb58f05bd7d564c4d5c3d157e51bfb6618d56a6d2e14047a7cc8395342779ebc1cf
z9dd98a8394140f42eca347ab920785da35e51ca06a0cecbbed412faeda70505d07ba36312c5cb3
zad0c6cf39e630e19bd9fd92943cdaec1c3e3331e85cbf9d20b143f175a08e0fe3823898eae76c2
z3cbd82056f0401de730e251886ab3d9db352e6f4f5ea3804ce6e931dc6a56c3406ad12a206384f
zc2f8f0dc1cc34f67edecbae13c22154aa84d7f799ebc2acfc4ec829460d18183282b8d491e4646
z6b1339550b017d6556527537e6c35f6db1e6f0cfffaae1e1c895b9ec6fb1847f4884a35f577f22
z020df9a4de7d43556f4794861ae5bfe2c156f17080e704fb8ea3ee0f38b71cc4a7ce2162237517
za3d211c08756ebbe62eb5b12e0d90e1e2c69096f4a6e806254e50c3b0649bfda51a912feba1d29
z655bcfad16717f0dc5094c7a4ee700a0835bf38dfee52b3a6018d509e70582b1d579bc09df9f5b
z9c8eec75950f2a9673cc59bacaa18c367f976c7405d994670d071ade65b2078687e78a6a8b1277
zc6b5abad6f6cdd81709fd87ae89f019973b5e4cfa134ba0c208073c297e670c164ac3e90865087
z2a2cf555a651a381b93a216ea207c6b514a5682448116063851dba7ae40acfad32ceecb91e8d97
zebae7552fd192aa3d8c22631650bcf94a16f06c2685ddb2b122401d71b8010bdf00ccf8cb7c4c2
zd3836209f3560bd800761f9cbe30a1ff35430c8f7d57f0499fb08716a8d8b129ed5a860bd59eda
z8df22e80cebe129e434411eac36e1da0923547a9d213e448b1da861cc9704661cf7bf4df967de5
zd6db1c9218e0845571a22b8a72525627b5dfaf8c86c034f6d6b4f2f8e851f20ca8915e6564dd50
z92477d82a6869bc3158761e09f50004ccd6023fe1dbab84fc2deec7b81c8a443051d7833eeb739
z52d71ba5037e46a94a282e7d02c546db95820e392738c785bc52c81eab6cf26cc3d449df587600
zaa0a94a993aec4fd6dcc6e7c62dbbb23e76cfd88587daee760c47a03c48147cc582a4efa0a2755
zea0f94493e760ed272fbbfd99d90ff9fc2e09a27c8f5536fda63a6cfdaa6fcaaa4c2a7aa812f62
zfffb18b76adfd8b68fe0ec6d56c6801e6433f32220cdb1a5b6685d20438d11e11230e1b2c3d797
z0e5f8de43a474ae5c1a9258a939e9a9559aa38bc9dc9066dff892785ffa14944d1d60e42f2402d
z5822341ba865e5437ffc22814b36728c6d8757b743e2e84c6a4fc0a908dc5ba0e7dc36ed1ccf78
z1ad10771b4e259d15ed530d8f3d2c7f7326e739f59627a59cc553768eff0985b129f62a53e8b2c
z2450b75de88765df10535679c0094239fc1e751c02ea5b3e1e9abaf8b4f562c2d088ae54543bad
z1b6a1515b52c26af3a5cbd28c44e0260f47a6a46ab66478f5b53e44f49337cd77b5a1e44d803e6
z8ec406f704631f6cfb07b41a772dfaf338ef80f5514625c6c15473d806ecd924fbd63aa99af961
z5ea196b482025d2a28e0564ed5cab58c317d13881257176fd2cc96be5d32876b34d52c3354a825
z5e77b3eaa45996f2e933a0b20fc591665ea82435ced2b9b33a6a52f63434fc291bd3850bcae8b1
zb73c1f0f507fa9c9b711d599f378a0e0d7ba85e96ea238d4259a7bd2857520fedce9f207f241d2
zfc043e322113269a8b27600f30f27c8ba86a64213ef90a19ef85d1dcea62d005a9a3b4974c5807
z05be8369a04641f748871c92cf14d9bdea59ef213ceef6d76536ca1fe5ee9ab201a281ecc66522
z5eb6480aec3b356898110cd822814a85f6d404485e67d36e8ec028e6d14356401aff51faad153a
zec3efbf6231f326d0b0685c5f7665e9970b057485e806158605defa345276491c978c80ab7abc4
zc33490d141b7f9d4331a210ef80d628393db66767917db2c274d27b8d3075c0d302d3a4e25e030
z4a55d3bb47591c447f0d9cf76a9b11b6502cce1a6c068fd06c7233debcda44437a416528a9a89a
z3e062e19616969f3c1bdeb89ea3080690ecdc4e87775c6d2081e618c9c62ffcd6ae18ff85233d4
zf971b90e37e459fa6b345099eeb7554e23f1bebd8c97cb21f84d3059d338b7e1a4abc2d8bb3933
z58f70780eb0106329acdf9377c2c8de6a811d5dbbc441e2386629e0d94f3feef2aac76d7e6dca8
z22a5c5d18f969ff4bab84b8db6474e45d72ab61f306edcc5177ab3b76aadd598a1a7f85e2fdb05
z7eff000d5908d224d6ebb968e1765ecbe347075e69bb43919aef42f6b99d6f6bd8be9334658a63
ze19ba1cf7afb6ae75e8a88748e90955b0986665ea59223d72bbb1c043b572f7d0c91a90043d5e8
z460b81d425d9c3c87d9d993814d60cab11389f7521765d62f3b876f5d52fe5619cd3bbe7a2a14a
zd55a0612bc55a1e2f0248487a38f5e4fa501a8f96e7be73611398472a85d279778e1b020f3650e
z3bfa8f3c819107a4a46c57c6dcc2d09388e53f3fdbf1ab6f68a2f1882b9dc52ee40cf969ba6fdd
z8c4877e739d3d44c0c95cd17a466c7bb39425343182384718c1d0aeeaa147d9a9ccf6841924b81
z2e14faeb40355b1341b8ea3721f3ae0cf6bef0ba703d3a76e75a03f460699c3382af59af0784be
z0a82232106d82ac934a2f100ea95e3dee2eb5c64047a548357506a83d56e80d7b788b730c2cc64
z7cc3c84e3af2108a407a663d9d126bc718103e4a97ab12d71ba8da04ce516ba586c35dfa267cfe
z6a2582722ac7f16f2f7d9e4b000a0e5cc6f0e4e0a4e87e15269469993a9111874b896463af5b09
zd763282b96a7cded28780675656bba5cc5bde6da51940b61af351e93ab0325c846c3d46ab6e96f
zda3b18fd8999585505ddc2e3c98ab4f69cd727ea302432f2d4ef04e106a2b85fb202770dd2bb57
z3314567c6ee12299ff84acaf927b0ae9b3ebcf075a8446ceb8e47aabd0c50fec173a865b69742a
z99e14abc3a1ba64d9a9fcef3404dbe20a642c96e90fe5972d9206bc3e8ff1347e2c022e16ebdb1
z8a92814789b68acbd991c65d7816c372838a9e2d7504460b82a1efa7472ce7d5cdf02064e4dd04
za65d0d9485802cbae66455840cbe554b3c22a10ebce0a29eb1980aaba2ca63c530f57101d00c84
z826dd540421af9d392b87583de69a05aa043b597051ceedb39c93cc60b1d09bcce49bdd8538cad
zd744d2dc3a607dbd4ec60e3168a7eb0a1dd8ab90a1c0f0a8b7cb4186713d9457bc379a4154deb2
za4d8c2d980f749fca8708fa94648d3ea2a0cdc2b837ad4049dfce765675549774c89d9d37157c5
z2a25d09cef1ddd5e1460ffe6e543c23e95d28e9a8206cf7482cc8147a625599776ce8043f8bd3f
zf5d99b7b82f8a769ec8fc3ef851a055f91898dc5376549cddf71075d88d5fd05fd83d6ee17a004
z430d6a8c513efe17de108b5bf44117ad6209361786121e59dafbcc4e665805115669e4be1ce49b
z3b1a8fd3302fbc67d960a586f5a5a13884226bade742a2485e1fcd1d014a1c216f9c329983799c
ze7c6cb79aa215ebe0b2db62378aa71af2ad517a711c18e0a714d6f026bce93ff3d0d45ca62574a
zf920e7f89dfa274f06be129a2034e23ac6803bb595f4dc15b58e6b46a87a6a327844d6f35f7363
z1af5ac393f8b14e17e1e9f2bea5f8979dfb51ea5e5facf701ca0a36b25444deca9049e7e6857d5
zcd6bab4e581a28b92b583647e190e1924a1f138070c4556df24faad21a1913809553119f3bf5db
z17508cfde852a5aa4d5cb02e3fc4414cbba18cf1aabecb960d8b953b4f421a27e56839c669e6c4
zde8f4f53de2c0040a694a1e30f6a77042e6902164097ec3d3ff2d60c5214d216fe2cda63ada4ec
zc1c71117ffb35e1c7e773f34a0771cb9d32e2d5b11b45bb32b205be81ebfd4c786f3e671cb5f61
zc264022b5df5296a9f98f3930a49d5d21633ec4ce9b173c4479c34b05090f011a0bf7e44aa4fb2
z133aa32309ac43ab79a3cb4f85cbe2b49642ba89ecbd95944296bed494e60052ca6e47c4757f56
z2c45f0eaae70884e570832d24d1fb44ca31d15fe611cc8c637a8e253fe46517400af4430bb62e5
z5539f564c90edc01f76dfd6ce1b78941ba3017a2e6b76c3e778dc5c8bb09f7033c4aed6ce9e1ee
zab3ec1af250e7f3466f59d24f09875d9eccd0748ca74281339784644b04cff6fdd0dd83f03a024
z9760ffd80929b27b0cc9b6c73a26da6c4b2bd815755268486cffd61ae56e90eb0c61450c5dbe75
z61a991c35c340452635c64a24554db420af60cd72894caa4fea528c1e658d3f1c4d73424b0d0c6
z7045e6e04be5ab4645ad76825b84aa8df2093d1a096da31c00171f99b59782b5fc16d066d29b1f
zd9b81bd7756b5dbb1bb3761690ad995ec533accc82ee5fb976314e914d37ff2a99ffff40d78a3e
z9cc2463a6bc15f339c93101c7ca4edc28e5e7c8f3a0c09c844c0bf755225f8a30c52453eb7914d
z66e50fbcb4cd268684f0b71c713b5e2506bd0cea44368cf716b3447798860fc963e1bae28fbc25
z1a701a5ad845b4b01b910b1ea51394d0873ddb5684e73919334f19fbd3ca0bebd657c7d26a180b
zb075a8fd494680e84de51070f957daefa02e559e267ccccc25d00ed4d7d020743bbe59ec394bb7
z1d6e3b1afa39037c1814a6ac78de5289f29e9fd8dc3ee5c2104fa45592e4763b5e8a641d9e593d
zc86eab02363ca2f7b3d26eaca2af7222f362e673269b11884499e75f822fe0a1ea789c205da589
zdf878bd1a36535a82b32d8f55964cbce0c376420a77e317762d567d75337d81b7e80b41326abcd
z886974df10971f6a4d237c3120346fac5c7c43ba24db6d2d3d11842068fdb17f903018d4b27d83
z74a978c712fd0b26e889fe774152138367d28bce0a1547d9338a34befb6d8176672197a0470a3d
za3d48970c8f52339d4f67f9337e85050c12cdeb57a3b6c9672972f51814571e8396c3318e7ee4d
zf60004b5bb2a6a0efed6e22f0e1ad48b0e6d9e2bcc1115ef8c111814880029cadaf5f560f76b28
zbcd17621df44ef8c81e16fd420c3c7663038d6dd129bafcfb2de56a8802c8a841bf2157758934b
z39115bb29323ebe1d9ced32b396e4f5d155ee8db54c34d58999f721bbc9ec341b3a1b6365137d2
z10fe327e8ced463ca9f4a2d15cbb62169532d524ad02df1f7bf8c72047f92c414bf72d235d5de1
z7ece621f13b24dbfce03cfefcbee4d407b978ff93a19057f374d2489b01ab046370cfebbf9bc48
zf6a7bb90c9e7c9eb2e31f9ceba1a270b9fb5a00a5fcd53728b02ece58b52d19f77b1c21c3caae8
zebc1233da91ce0cff08147a84ddf0d5d8020932bebb0d962eee2c529c6b3ad2d3ba4926f712f36
zf0d7883dc317f0ac381d8adbd4523bcb44ee5e30b369f6ae8329d38fb03fb690fc68736003bb0c
z0b04d0c12087374cee890f8b53acc6002eaa68debb106a02b61a4d75dae8ffb0cb6988c8e62f07
z6a0a97f638c35953e49c44f750caf2d19d1a3bdc1f2cdadb09f2d6c9e2f09e6bb10c48c5c7adcf
z93cd06227b8348fa2f55a743850b954a57ae10dbd448494408e9debcc778a296ad8eeadd3e5153
zae734de9a260dc28d312dd17fbfb12e6997d73a0007636813146f06a46f603929aafcb4d6f2218
zb567d17fbda761c9c7b8e6bbf5cf4d59e3aa7104d02d7e6669f0180f609bb2f513e6901071aeec
z60500606ff04a1b7010462fcc1c2bf489570e2fbbd65517e6fd198c5c08641a9c5dfd515faa31c
z1bc1d392e54a5cc55ff8ce342cf405b04366abf429421ba51d18837e0f2459eebd8adafc809b2d
zceb91f40696caaf690b7aeaf32db85941e4aed73fd7e2a7c367f87f8d864c0eff958afb9f7f706
z45a15ff99199bf5fcbf9ad53e8c559499e478c624fe6ff98c1a7131fc529a8fadb18f99662a1fd
z305f9ee46acc429dda7f432f8a102d961ae3925f3bc96b1d43a572747a84e0301a0f8534b4a92b
z48581933c1f15a16b713d78a6c8de8bdc017a4ca9eb83814b5356f88cbab51b6f1e1cb84bb63bf
z40b173d32f4c899dc2446e874aaa45e8f1bff6441ff30e2794fddefc712ce08c4e89e0fba1dc3c
zcf92639c72e2778a6fb45b53055540496af0c98a0def642b1a08543b64badeed3f81e362b2d326
z435e9d26210c9fded6aabb314a351cd81a0e019ea31106ddd0aaeac367f7cc371d2f0670177768
z71d5b6fce71429e90d4a7a435f76e3548f2788a6800c4873c1cbea1540851a0f62e06e5ae28f58
z6f48edaf938a3c8ff2c21e5b750bd3a516702b7a3a4cf749abb51ddc6e176e5065b727b061d922
zce5ad38852ba41aaaeb31c5989251884d814a68ab7c559bfd19ec2e7fa9ed3648cc6d9826dee82
z130dfd898576218c8d10a5eb16fce1b6f7a70f55a93d76173d397ad142c32d9630b710591c8046
z0c51ed90289befffab70341371d41cb2248f4e6b04c76162f02a9466f2bc14f21c65607482e507
z03700ce7fd851fe917d63a193ab7d39f1dbd9ce415c2166ef60027d678ffad287c0882253e3a47
z3d5b12c395e4cf4004726c5fc9f807f335069007010cf276b36f59153ffb7190d4a8db75af0c8a
z0835378802fa97f3cfcc17347742212b58eaa0508b9e91cffb168106ceea9cdc34b07d0bab8439
z87896d834d5beba4f84d052606ab7ebd35a4a22f9469ac7d592e763f561fe90f44c2e6df01fefc
z47a5599e7a9f0266f337942be8244b8033082928c54b960d1fa20652d7f4bbb2d6f5e28dbf1822
z1d8378f2ff535f4ccb2b81189f9e5695442a5df10d6316e1d8846f364abd9b04755cf901bcf5b7
z6f42d06d14270667cba6c634a22e732387c0aa749a9880e19288f55e7c937ce8a81d19efe0d9e3
z8a0d0a3c43bdaceb10a6369205dfffc21c4e501c3a8c2ffb00ff013ece8069da79312af167d957
z7eff71b6523c871f108cdfb9f28403e8f7d62ec5f32eaf4f8845300f905b30f413660ce8d6e0c7
z6811e07f52f4fecde06c6cce2325e82b915af3ff1490551f782f7ea483b18d027a93a736e57efc
z1a5216e7bcd9b461750f787480a4c175f4198f9c58f7f4e4f46cc5bfc14b30e45f6a4a319214b9
zf0d9ffe1b0aaebff472671054c33ac646850635f245b08e72d25aa53ffa648329e4a80933d2417
zd0da764fef35b2cc8f8c1b4b7ffe534472733bb257a9cb3f92fbf990bb463f05f0f05e2f4d6316
z01018e0268d84ee2128bbf7c2e2d93c201aa6651e03a050f0ad9fd231ba04aa1201dd4c4b9df70
z909b7561617e7b9f5cb5dbb8064866386182477570573f9a0441af93ba438408c2867d4e1c0e27
zc7d341c916cdc896efedfb61f9924e9079431225318b31495155e6c929285f509e336b2fe317bb
ze8ea1e1c06fcd59d085c80811bbf5de3c1ec98c517219d68bf80ad00001c36bb1b14abe28339e8
z79e2de18fcec26cc9fb008ead03c7e5c2214281a402bc65fe400497df5b97bc31229ca946f169a
z2758a2f07d8f0f6e26dd1e8d3105dc13360dcfb08b48bf9102b1438a74e930d4ac91f17210861c
z7def70b161c0097bd74b219dd59eb4fe9492cc317bfea746bab35fd72e49a27bc04d1792d4e9b0
z744da79f434f84a7d3af3b1431147ec5be900bb3e664bc379ba72e5a9cbb6bf470e581a6f74382
ze20d9cd27b63f2b8fe506e05c957400730efdb225ad44b8a3a8dcb7f85ef081e726097f4c12621
z23369a0f415750836b263744d70af845800a4c9e18d9e9e23257bae6e4b72ea0ba6cde49cc71e3
z8be4017ff54aa3e04e6449b1d05ebdaf411b7262a2208ccdebeb202b15506900bb2710f4bb2271
z95dc0c56023c12324d2d2140cdd95cf682133381f734bcf25166ac59818a3a9a680df02223d68f
z9219c8b900c40fa4da4033f516b5c2fca1d34df85a2a69d8cbff7ce1db11758012cca5f4c8a6e4
z2b34108834e4716a114ee8270acecf4e121e321ca00131419c5bb787be30e17cc41ec5a14c0dae
zbdc9ddbc03636d158c4ef89f5c4ce3f3d0665263fb5b62d6be6bced6a54392f471de7372750f9c
z3656d628312aff940a3870bd18a8f19f0656d28e0aa1a794a94329be7da2c861c5165d8406001a
zeed66da4e6316d313e9581d4fe1822fe2b6d41929cd6f988c77da3a957447ae35899367b4152ff
ze4883a379d385bf8c628ea137f2e7436e457373f3135849ba06553fff050e1ebb4c6ea6e4ed931
z9c985c4a832e44c9d4c2266ab71e7d2e3941efee06a5af8397abe80b39d2c6dd9fd58cc805f0d7
z4fc52a662bcbd95cdc2e035007caa5141b31d63129fbb33b1a3ed15ff65786200df511ab53faa3
z511e4bbdf2796cbe812dcab54e44f79169e5beff8d8e3eedfd85334a640cc594afb236cf29c29e
z3212f7bcfb7929f140e84e02672e2b58a5db75cd00cb928723c0c290e644f834184e67ead8425a
z7b7296b70528822a345c4e3de22e6a686a25bd358cd85ff26ce8fca4440a1dc3801770e89f6e71
z96bd673f1ff02754ecaf7d1ef1d69e81e76d1f1a8c486ce6e22e0ecef4af4b912836cfcd963ac6
zd2baf1597194175a441b08e0fe2302cccf12fecb2df014f8e536819a91e1c24138ac01212301ac
z281fe6209d5b1df1dda90c217cf1176f30cf085c01f49ab94b090333383db5a9b261cc5d186a84
zd50af2d5c9d6342e6a7a35eb2a40bebfe99277bdf4039491b7b64a657af3ce67549a6237437cdb
z4056e424cf298152999ce23ceb10a5506203645bcb0bceee298cf358dd9ac5f2f80cf7414d11fa
z465519dc70e4fc5d3b8b8bdf5ee367fd82d77befd64e3330009c274ae374de4477ceaf0bf9c8bd
z8b3930f833c097680acbf9a80122c801e569e015b35431122dbc36f181cf54db19ddc434d521f5
z31890a452f86d00f33fa6a42b19914a562be26af30ff77e652b8f2203ac0f9470bc82cedb990c3
zadb0c9aa4a76ccde5bfa46f6c1a35e0480631a1ff668706f707d2a125508e12eb2093e9093b90a
z49d7b5964ffeb8f552e84f5064af8bf33b0b61e36f9c2a9b427aa56816179a307fccd83bdd39b8
z91ce151259eea5d5eeb84e9cb50260d9e1b6621cbf758e4b76671a3471162164b610e4ca77e0d9
z9a8581c5e679b56d1ba91fece418d177362f1b23fadb48918d365b7629064a50abb86188375cc8
z9db3abc3393f8c27cd5874538815a99b995e798846ab3bd35935d49514c1716d8e963f9e8d82f9
z06cf010d52ef46ee103d7da6850c911f6f594b70df06bd753b2081cde5a48b930f220571cc6e62
zdaf34d54fecdcf71ac15e949f98dd5153fa782d7984c117f66015d2bb21e7eb84e990fc36c1d59
z8c7690aa2fe687f9f372b61e27d7c44b9e1ba8c4359260a95a1e175f9cc876b00e2b1027bb6d33
z81ce621fc11ff3468f6ae4ba8735e229b038852bbb7204bcf70e1648a7e13db721a1e058b0ea0c
zb649ba70893da70fc10e4be71d473e66140e47131651c86278cc11043e87c59d99b5c1de2244bd
z066080dd77c542f763c872feaecaa661d2fecc6fb6ee018fb3f8b946388e1a30cff939e83f0926
zd99f8c87776997693363a839c5c6a801506d0c209f8c2f05f30687ad20090fb2ebdf7421140fab
za4342ffca22b3d393a67cbd73c7de00880d429b9bf68511edcc30fe025c01d1401fbc0007dd074
z48759f699499185ea67c8b9c1d6aee862901a537065021db7dc5d9efaad6ac5a503893b81b723e
zd8fb7811f871f3ef83e08767049b9d64fc932b39aeac7dd716d05d1136e1463227f03c65cb4372
z147331bef206dfc5208ed17c388fb7b2458f3b1dc13f7b76b1858011687ea460efc4b2ddddd8c7
zcf0ad5831a3fedcf725be7ba27592194b9e9fe0d4cc476560d2b2114ec0a7b75cac70907a3ffa2
z88ca31129456174359a49e26039fb29819591e246cbd02729ca3b1b381d525b3e064fb0a211c50
za7ba216ecf8aef7db1abe90c9b68121b985dfbbe642e299a4eae5b4b799f3e63d61524dd4bd65b
za3ec25f2f706e8078f2759b39268de3bef859c88c99c73160e2665545d471356949e1acefcd128
zd9fae41888b535243143159c62323cb463527aa757586bb577a89e9492694aeed19ac7edf77a40
z17e0d48d333ba43e08118da4c8f9516a38f947f3d187f65d26ebc2a2f976e554406d2ad9d643d5
ze3a84b6e2f5309ab540a3feadc88afbfb22020cd2438888eb5cf561fe993edb5e7097161611eeb
zd20640d6bce83e887390d57e74e8f7d1c5d9bb19f1eaddf340e063d0bf597276950e5daa01f46d
ze04179d99788ca2fc7a59d806d9d16ebb8a237aed09f6076d304b83fbae661e19b361488527fc6
z9d989d44a8b0cf93da3adbe5a3605b29e90f5605376e5aba2de8118c301c94cdd4f12ab6da7ab2
zc59f6a73c8117eee88127c36a825550f5618fc5b655360021ffd6df4952a6c832a96d14ea6608e
zbafa8ed62259759f6e2fc5cc1e93bd30f38aa6df40f12d5137c93cfcc40816b9197a197825a028
z04b7af4944aa20379758da66817c731a4c7b3e3a3cc6d7576cb384a7e2b1b7540ce3b6f16dbe1c
z4f7d754f1ab2c26845ab0be9a6a1ace9436aab1328d27bf1ae103054951511e2eeee3013c8f8ec
z6ee71a028921cae63f5282ab998c034395044cf9680a4db869f2e249dca0d905defe6aace3d515
zbb354bda37547845adfc05886012e9bb44aa2183b0316331dc46b446e7843e2172d8fa459005b5
zd825c43c013a6469a47e71da75ff86a02970285bdbbdcbb1533ef5d0083948d76dfd971a17cd31
z5702a8a697831c277d8bb0361b778bc935931dfd9cde3b04ce3dd8de2a0f131c039358ecfbbbe9
zfe4558ca6242b40ae2f7cba047e429fc99da57a66139cf04f5591584872151439e7589c29bf623
z5eb3f216f1d9995899d9fe81e4ebb628b06061caf3b8685189ba7cf3091c28b6db2d0548361d95
z59ad5146d61e0c5b50b425defd1ecc146f7a509f874bfc84ae6c854f13fcbaa7f1701d7cc3608e
z9605dbfe211ac305c08c39924958584c3e9a34c4a945277dd5f427b27e2b1096066838c84fad05
z603e73400c8e40d091a3c3b88f4f1c5c5ff30fa71d78097b02eda6c4d9dc14842b0f42dfe6f50c
z2d45dbdfde10a2c3fa6a0bf8fce732f5d2d35725bdb3070252e59be9265864106dc658eb850b30
zbd42df2264e7244bb888a8305f2a8cf645d683fb31259d4d959456bddec494d78d65b9e4722da1
z296aed55ac62d4fa02fd7b358392bdca2ba4347e0b7504d9d5f48c9887976fb0a181c29dd10c4f
zf4f1d3a0a7fca4ffb355eebe378b4e353b072e539dd5c494a63c3a2080661071c2de5f00e038af
zfbe1158b22f1624e8c72cd8235b8985bf30b0e53e4410c925dc47f6a8d2bb24846d6f95f281161
z63d99f8515e2b6e3a12e7c2ef5b99e850f275b5d5af4f76f8a10d4338f7b2ab15ce8bd6776057a
zc3025305b50f7fccd995abb6f216f1a92bbeac08622436088ccabbf191d3048d65897a2085ae8b
zaa4b5886201781950ab3c18e7d1afefb4beec508bd3d59604df62f86bbf24a76ea2c4f91bf7248
zed1bc7b8741ff643cbfb87542dbf4a57b14082a06beba863ba04dc7e1630aefb07e552d64f0e15
z15f7f0302ec6042bf1c0cddc9a884a626f5407760e7ca6b073933d58b83c3aca0361263c38a04b
z715bb4fbea369288eb6e4747c166b127a638bead3c1f71d293147e555da95f7fc1fe7d76550bf3
zad1eb75a79170d784ecf9c12258651b855d824e013413b85fb5cc8a7ad98756f0c9823edff717e
zedcf2fba0217b505cdcd12d2c7ae8a1ec7be76a647d3b803252cfe2d0d93f2a7be1154d2cdd1d9
z3687e0ed577c67f75ac0cb60374e30c2726f8670547cc965d5b2793e1a21edd48a289987f53612
z145a2a89438dcdfbc24e3841e8ee82174c982325736f55a0182eee25f9e77f0717f7dcade9bf9f
z68a449075a788c8bb710740392fce33ba28361f63c9c076932f09dfefa64ee436ea824e77c8896
z232383d1288ab1f08017430a1e803ec11caf76a222bcb0092ca7ac3f02b14a21f4d99ba3484f80
zee16decd68b9c8a92ebfb6b4baa0ed8391a4f70fdfef85dcc2ec7b5647ddcd8a8b425523e1f1e6
zcb01fa36b1dc55b09e5b57d09b13dea373ac4c627c0eecad51060092788fe26adac1e985359bb6
zabba1b34f9797e06b858efebcaca0a043b4c9e991a1a59ce8ae9eb337fefe7c9f1d809c8df2176
zf936e15656bd62dab1e5eb3da72091ce3e3604bb31f528d9bff3132b6a6c78218f2466efee39d1
zd356a2b2352414f28973dfdcedd1636776c683a9704afa9b63ffd9142a8cee31b29cff2e2d636e
z9efc2252849d46e755303e8686094c034d10989b08385b5f965c7ecde04efb6c76343cdf704000
z7cdca72c65cff4ce8d270f5a7e76c27592a1da64ebee63a74ac5a718c2ec014835890a6cdd28f8
z832119d63a531a8a4355c2de3569047a3c989d3c56c4495408a89e1e02d58d7e1419da42010fd7
zc95b19fde8353e3611570d999eaf65038f42dd1eac572fc4496fbf3a0ccb491f3920036f7c2cb5
zdab4453e6dd4035581daf537facd439fd8122f2b1675e5803d4b2db3041b741e9c5c591643b74e
z22d9efb15f5dfe5931e24dc351eebcba8cca147d10cae4c24ee854338de3265a8e98941419dd99
zea04d8c9d3dbce41a5ec60c97ceaf347ec4e94e92209add7066eb5f2033df917145ef09ed5bc5f
z6d99520115879a16e96b6778a4a68fd79c8706c7f1678cfcb1190692c100cc5f7671121d53aed0
z5363c8421ba4e79e3e2f9890d4a04e2615974973d202930e58dd17d7d161a93e56206ec3b0e662
zf947e892ac3fbd7e7848337b5b7c36aa7f42fba6d6bb5f879c927b97bea5ff20d579dc383bd7c3
z3018fbcc8c7ff3cfd520c62ed31619188503dee642f58b50dc368d28701030e91f385d0dd95cc7
z6eee3b0d12e646607656f1823a2eae04ec0dec170cace054da4aedbf43e46d518f4fd2fdedbb06
zbc128885ccb75111d8f65745e441ddfee6637ee9bbc7fca14a9a9e890d9c738d410559575362c1
zcabceb9dce4891f0962eb66b815d9722fc2dcbcbf79aab2137cd063536f6efc933feae8aa25cd7
z8a7d2be7ae4b820b60a3ff5b588b0cdd2f02d4f8e99807fefa7a95d68beacefc5e41647aec8e51
zc5c6d0262544688e0f971e39d80461fcd4fae367078ca9d91bdbf82fb58dcfdd0180102a0f5724
zed50803b721182c97e449eb5292ba9bc212cee13dcb4ee13661cdf33bc1d04b4b7e18da39eec68
z6ca0d42233948d7720f9c6ae02476b58a911ebdc54bb0912e8a74420879f3adb26f6e09cfd04f0
z22a10b9947c370125280aabf81ceb27542f043e92d43db0a03628d4914b67392379dd5fc956445
z721bd9e553f6ba4daa32a565ae935ea4bcade07f46784314b39c2398bb45360fef77a19a91ffc9
z70ac6399f82c7d4787d602cf8eb89b157788e789b299e512980734841ea61d4a
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_fifo_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
