`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff98478405cb2c034d92a13b0536cf592c53efa2bc42b272
z5c52ed0dbbbf085eaf8efe097f8c883c462180ba59d4c6ed9946d2ecd2f7e48dae4f0b7e0f032c
z999d801d1c8e430c47c67962b0990dbedd8d823d21397c50d50f02b47eecdfa92812e746860485
z2dbf6f2f01db1ff3b6d1100da4c75eb1267d3b9978696b9eefabeed59c314f1d2e239b41699cb0
zd8a2c58b1960232c29af39617d93b134c86759c12955c49d526ef01e3f36b74b4a4db0d501dd21
zdbe0d3f3fe86b1b61647412119b39ea02237a0503cd73cf608443bf282b7986fdc42fa87999978
zaa252f48256e23a64287a631616a42d8e6adda0c9081a7b0056a8b8760018c8aa165aa83c661a6
z30d999f1f73f1556f87fb1809a20f960a226a52c7bfcd979a276e3f996ca2cce751151eec09ce3
zf42d11cffa09cbfb28a0b8bae9d8b511fd47829d2377aea8e8b99a2e8cba00e656245f16d32dab
zad4c2fc92ad8ab5c85b59c0917a1f89b1f8ee853b0941433096723d7992251d53cb7ad44ef1133
z5a46dfdadc67b3c338b6ce718760f468767f26705a43c25b97aa024d5c7cdf5ee26b740d3e2b91
z226891fe060a776c478544d5c7c50cf9b1750f771f018bd2e71394241ffd798dfe7ca765ca5627
z0a28ded5437f38586db042f50e21c9dfbb7f13202556b112e7210ca07a7745bdd49cd3987d8c29
z9d64da53f09bbff15cae7232ca1f91c00281b8568712a06c26c1d4fa2e5302998d1a9c07360814
z77498845284a78722340cc67b908ad857026b4c14d412a4fed4e3d4b3d899a4b55dad3696c4980
z26722bbdc7509e3db416efc5973d4d2a38f7d53ae630cbe66bb937c632c46441c0884e4603d0e4
z736c521a22b8cdaf4664fc72481782325f86b986c978b7029b705e9c287790952a87d86a98afb2
z8c272d15cfa78a27e5a7742935b2f63920f48bc18ef527c06e445d75cc431934ca873ab0482a9e
za1fc6092dd66e092794a9ef30e26f8ee31f194cda3e429c142cd18b78ab59a4a1289912596b062
ze402b5ef158506a87561e5e61a3ba703791c907c58694604d454a6ffd1fff0b116b09add4f4876
z97d912116bf4852bb8e6212e3a51e7d6fd9f29d66bd8ec279f6a4f1d8ff79ba473ff1636666513
zd0bde03f0fa3827a952a49e6f790e228666227200ec35bbe3dccf1999625a3e2d82bf502e8d324
z6a1c7a6f65bbe8cac6aa02a69ba241581dab00d3adaa14f78e2ce971f76eaf5f334c1fafc8cb15
z0e5b69d6385cd5c660230b1828ef05bafd605323318744f26b267dc7fe4be956e2ca3c2b0b0947
z9e3f845d4ef84d052026f0c99d83df6ab649cbdcd7afff1c882394b273e590614b23d9403efd46
z627649d2fe74454d0ffa15e82053900282928f95a93a5fb053407dc9c24543ade3852b64926e75
z48ba86b4d0d8bc729840a4daf454db72f58776fdc4d1649eda3832a75f6cc037497e1d0442e4e7
z446ccbdf76e732cf7d2a23461261e3805a3f626d48409b28b254e9805c9f67af188cc96c97f707
za4907ac21ebcb8aa0f2559b42ff6b27618dfaa4931745fe28a1463c6cae86c5f4ca66d60891e83
zc472e5d6d5c1f4e1fbdb3d2548acb4dc108c0e0dfaa6f6cd2e14b8bfdde57294e75e30e51030e5
z712b7330ec28c3241d7ece7b3614058410380b6386d06d6316caa80111f661b9544c9985d9577f
za1cbb46f3915c219a43e57a283ac0cb02bd84b17ac2b088da8f12d7984926e4bde566378ef7dd3
ze51b17d151ee20fbdc03f3638ee4582874944e3488674e87e0fd3a53caa9090abf8d67b873980b
zaac7ec01a7e964c6f0d7540008f8c9e4ebeaf9d67902af088da29d83a01039e0956099f6bca432
z3923a5db82b76dd30f445e4a58d6190416b025c6adaf57cda9c3876c154b55169b952ad0076708
z82015234b017fec39a667d2cc36beb44ebecffeaf79f8ae569ea107b8f075187f3f8d1f592249b
z0efc8c5530f5310052932f7abc956b7821514952074902d17afc4c1caaae95bf9e94dee35da21f
z76ac91506f6a76f009fbf80b00c991f612238184ad2d66991d99d1a9337fdd6a1a9c1034c3d6f4
z8072032d2216af48b79fbc6c61ba0a4fa2a4cc4b08c78c558e6c3508526a7725cd83cd1e741345
z12c0e2ddb3882d71419b7733d86ee1b1256240ad19e52ca09b4304d3cf1ca261f8f16b01a8d3ad
z93fee5b5e39e92153504a2b393564efc53878c306d9692479c3916fcb107cf1db54c2eda15c7f5
z0099ff01fa3c303558f00a4c4753095eb851ebb7a12589c284e69eb7605512e677a62d08f5666f
z198253829d5d87ed81862148502c6e65709c7c8810537a5f53948b52d3a01e12fceb8c5de3086e
z7a8cd16b85a1fe9ba198d9656f04f3dae60af45227a0f02df29e60288e563b8460abfef550f8fa
z4ef13a7613b6ccce59cf889400c2f6b8156b6fca572c564fa7ad1c50ef19aa666b07ac6aafc9a7
z1ef8ce6726850487ad123a134b7094af36a8033dce957aa038a2c858b3b65a5a489419f1b6f6c2
z3644ab6409a4858509e69f2af32260f33ea17bd2eab90439acbd2df0130423704d22e6dd42b79e
z0674f686fb79a29006d97badffd852323eca9827a3c39b73fa8c167004b2117e6303eb19b3b258
zd0fcd5bf9ede4f6266029298d33e2905a9925514b66b4d6e7857d33e9d8e6cc5dc3405691a548d
z773884e4a7a5b3b07cfe61b2b10b61cc3e70bc642f1b496008a7c1f9a385dd559799d46b8bcf53
z67531e65d8708f2aed4317a5b1a6708d716b11ef00faa414380bfa1ce93dfd2c863e2b4105d243
za839639fb393e4849f2233efeaffc5500a5abb2c75253d6bfaaeed1d711caf513ffecdcc3a439f
zf8f6fc26c46d8241c67273151c7d1cb1cff24991ff5bcf7adca92e3183beddfca648117e8b3cc2
ze4e61341638b07316a6c0ea5639c8b46c03a3eb46decb3f50de7d11626c0d8e4429270a8427f4c
zdcbf2c2c050a7d245c0aac6e1b316e0eb6585ba64ea7aa927cadfef703b3afed5b4c61189590c5
z75bd7ef269ecc19372eb3fde1fe5fd2a361612299fa2e535a4abfeefa065b36406982bc31d00d0
zeef29c6611c2b63c44732f0be944e05bbfb8eb125cd2ce9b8dc17d7d74901bca60ae1f861e02b2
zc40b0d539083773803b377a6ba94cabc3b03fa96f58ca4dc660f3c5e0b4d9d78208fc71efc69f0
z2f72657f1193768321d928fd3627b9332714fd3298876566f4c879ee5488d58ceb6fbc4b24752c
z52b1d4bd55605e819462fe71a5ffa8dabea231ce1d8e411d24acd07b205ea54711d04d9a9a7d23
z572c695567880a5ed5952226dee55fdfc464b44c4d80de7b58da49a5c9a404173fbf8a8e416251
z9aca7c10d8c2f6f76f01eee93896fc8d5c13c804a556d9761c35fb3b30a6f1ec820bfe9d13c647
z9a8d236769b53a08e8c17d489f436361b94184c9d9a94ad1929d3d040c93ed56b4afef8611fecf
zf8227c038a26a4f7cf8c52aac6c3e03d4701869b723aca6e2a47c5fea93e7f67f6e02af75b57bf
z0e38bebff8cdaa1a7d7c71118548e6304133051bfc7ba9603c733ba924d7ea5e19fb75c890daec
z33444463ce05ae220297b96601dbfb00d61aaa3a93565757a2ea5ab7804676a141d7ef594c8ddc
z078d502d0bfef7050fd7fc99939f1b04d95dbeba43ec5804ebb36f54ba8a077b4f2cdb35c0cfa3
z89d0e091c91e977e8d4d9529cde46cd8215aeae95f0892916eaeef44205a1954e0658131fc803b
z66abaaba35d9ff4f9ed025e4f7086643906ce8741525814e88d0fdf8d52a7255d9d67eb38ef39d
z5c63424ac5ee3d53e0699c00a13fd3a3cb54ab51207d0d1748189aeb512a9dc6ee80288a48917e
z506cf1a80ab9eaa4f71e450059f192cd95d80333a34ed91f186820a9b607a75b845ea2f12672b9
z9d919d02d0785329025111aae6922cb177c9d49a6c0ca0b13051b4e954fa9afd6ccf031b6a4bf0
zfdf85b0fe5f07d80475a418575eb3ae3603cf3b38da93dfe1ca87a78b84008bfc9d4f44d8796fc
zcba8ccfb65c048cbdf09a032ec32fc940dea0943108e0853d18c951cc26e58c29077a531a83729
z88d64e1e69bbdd93836d007bc5335e0ba0986069a3c6b4cc6d01958a6dc8d8f52102aef0ba6fe6
z165ad75c56fd9dda47e77569050d9f7137043b8e31ff28d8a6acd11140d1e1fe7009587c533d8d
z12b1215c0c2f152bc6cc482dd9a3697ae74b5527da02edc3dd8845dfe240530c10c75176b75002
z00dba7297f76878025796eaea5787ec931606f0d4291b4e4ba7e0973e6ff0d1eae7a945b9e14dc
z4439f78274599661de70b23f8396c41f27243a2e0f80c61be69a73df9633519ac076e2cf34661a
ze9ec374c79e0c624b552b99d5754fc88519abd2a7ae817d3dc933eb68e1abc40873956039863d3
z94055b0852ba830f089ca8682aac92366a7dd5dfec0743fe9bbf96ea7ec94a1bf526361f19f958
z4bd3381f312337e2c044fed6f6004fc52935c4aefd8f66f7b1fb649f0f4f794eff57b47946fc1b
zb45d945cca0d70d1b311b222625b33a7b4fed3edf09479c464d77a0c2b37187e9eb0d0730c04f7
z874fd5aa8040719f1761f0cdd5825c66bb6d20db1ff4b00f734b1db3cc1a3812704660f1db62a0
zd27ebb051b710521d30ec06b9ed7345eae67a3563ad3403e6bb8ab4f4728361f7a11e25ea13f58
z93755d4cbc826f9bfcd7f67e698da67bbc89278b96813ad66a544e6cfe8708e9392d21d70ba9f8
z05c31bd500357797425f95f5f7d2858ad98a5b95cf58d5a6d7c47f89b99d5985a3d2ea14674340
z7e13e247fecca27ab5a6696336fdd0e3babe5bd4d5b7439c08b8357e628215c9f348ac4e579ea7
z636635142730f615cf18595ebe937a3bf73957d3298a301487c65d6cbf6624534399e94f623795
zbfe2f738ec0ce3dd7432b97d8b2b1547beb56baf53339244bfe53068588b55ac04bda85d126e4b
z78d88ccdcf8460dbe06099fbaddf41912dd942233ed51228db40d857711a53265df1c6ab32bbce
zdccdce88866acef4951ee87e8a5663d0ed0b548f3cee2133163bfe90dbd440914208cb12493034
z82a5a817a8f4789015f73a0e58c80732ee97fef6addb2a39cfb7a01c8490df91fb20e16a7ef117
z77ea098dc1f213ba457224ca487fdc26f7cf88a3266bdbd79b753980652663c80389038d603470
z77e9d468a36535a0ba9f5a68399cc3c2ca492e093a9137bf9eca8f9895e366e2ec18537087e6b9
z7e248b705d50c68cd70557951fa35ea3187507094cde1e59b35cb17d5663bf751ac24975fd19ef
z90e3e307e0512a82377549f33d29afe8ae5ad6e6e147eb1c47d9f5dbaa26b5f5b358a32ff265f5
zacb6d7181b115d25eaca5137eef9fe4355e34a266618a5ee5b4e50ed5da478a4d82caf47013bfc
z964ce104b256f3d06e6c2e9556cd0efc786fd6e0394064102e22e3df47b63ce539b1d642acf131
zf03245d16bf7ba979889210443063dd5c24c19e17abe3581f2c0001edf6d45e638f4875416ff27
zb9bcbba14627ae9ae706abcc1b05273293899f60065eb5e850a7b02fd570f9e19dfb3af54c8b95
za9d8de6dc383cbca185a9574d474384b473354179cea3bf619b77762dba3f98bda3f8837e15752
z646a069ba5e9c5fafac03ec1edf32b8daedb84bb9403fd301f60d12538e2b870156eed8fb335bc
zb741edd3f38a75ddff0e70dcf443a7b6de58b4dea4e027de680459c00512fa21648c5578bd61d3
z338102bb22f18f73784ad8aa76198d16fb85615184ac5e5b356a8f6d4351472be17de184a42bb2
z668f59eb3b187f562a4066530656cb8a1db29581357f3b9fc4572f0a184266f06c0893277f80c5
zf8ed6425ae94bf44b046d2867651307bb86dd840bb4584ca3c31b3b823dbd0f13ac50e29dcfe4f
z1faa0e7d8079e3e2cd20a7f5ceb3e4cbf5d46959cf620226c188a81d0c7b6a8111338e98399e68
zc2a0974946312160358221859bde01f41ccefba143960629e6e33cfca6e338b28b8d32eca441c2
z1c765c6dcd8ac0983aa26250c0e33e8c32bedabef7a1b13dd9374f27b2e0cd6153add7a5c21f3a
z7fac1c8277973706b19143a14398dfff6f70357b17e4d63eff3fab635aa22adec7dfd7b9647ecd
z8f7314d3f3d0b83bf0e1387d8518715ed41b5ab5e5815de88918011b0a90138ecae7c3de593f04
zca03d9fdde6cef296b0e34a6af709c0bc6e2fbd04c63353e488c76e2f34555d023c961b365d71b
z078a359f316ccab73b2eb5f756cf8c9ade2376411c98356cccad255c0136b1a7143a84c444e425
z4831271744fc81c07fd2b9a8f769b89524c2a46b80229f3d109cd9e964c0ecfefc96e94d9f41fc
z7f27bda0e0bed8a7bad6458fa11e792aecf0626c709c584688b8aad3c2a3fbec9fcbaec7d27e24
z0ec5763afa321ffa0b76d6a50358d5212b2356608815084791cf62fe17d1ad753562fdd96ceb66
z07618e745dd5566afd6ceba0b2c5f0938f277d5be79ef36e9d6f58653382420e8f6a6b619881a1
z6e849ecf45383db45cea87c1ca34bf940d691cfe86bb46210afa0c59d850120600e98d6993556c
z83674c72d44ded4f5eb71c856deec370a834528e33fd1ddaf1a5477f2ce0efe108bc88a1bc076c
z9aecc3f2ab9f53832491aa461b1ef573fec2440845e697c96f30547b7f9b2220c1cc011e2e7baf
z716c83c4882f05d99864eb8bc1f4b1b591602f86de918ecd1842615c1cbcfab8b1ca41cdcd59d7
zd541697fc8ad00331a2c28b2c3af9eeecff04017a83789fd6e08b0e3d887dbf3a7a0e17282ec7a
z21ed88e52b1783d807b27bd39aec46416b88b5379af68c593fb629988c70b367a1026a1fa12fec
z89514d87b1259dca9d94b4b33e0210f8f312fee2af04134090d5f1b789f2bde7f17c2a03f9d5c0
z41b9cd3d8a516a3e28a8c2c8f17e9da92cd99856cf4e89d4c30cc45d3b61dfd12085bff56826b1
z5fa46563079ce9bf08440d02149b0e50f6bd6d94f57bca370e0544274fc1d97be4259b15950a72
zb7eae482a62e278ff23ae7c3b93dc2ba3b5afb047db4100f052d69d2992852ba2f9d2389e23290
z09a4c6a2267cbc1a4989d62e60074cee52a821120415dd46960b005a59f4b43a48e13a0ddd4b65
zf84c54e522205710c52d68cef9b35698b0316cc11bf53961a4d4535e40f1d476654d7e07f7ef17
z93095500270637dedba377cc267b7eeeb3e3c57a94b82064400304f328d8402b7ed9622f050f49
z53f227d9ae7addd4a514ff90813abd78b47804c6ae508123830fbffa8b7acb649ed9c6f71a5893
z959c9ec41a9dbae4732e39f304078d5a7a7512a1c64d237f78b9a499ae2e38d9e40b0801a52297
z00ee95ea97fd3290a862e6f6939d07aae85c852af6f1069e3a6a1059fe99e4c06766d753aedd59
zec7bf41e6b5785e9d5625fa56386bd5e6419dcfb4c061d5bbc5f36156b75dca2b9bb79dc64e594
za2fbeb682ecf1c7590419774d5afca3ac5b765563056886fba599d5bb1516ae85ac71c5936e9b8
zff84b455e1fe583a6b694bcb4bcca01700143a8d1f890c29d4e9b025ed9d9deaf0cc0bcc8953e8
z320fbfbabb2b4d2fbf758a9726f7fc6b1c6a9f182ecb5ae1b3e1ca0a12ba6f068eba110a935d11
z45f6f9fbaf4c3936c9085f64852a24b09b1607ec1a4bc0ef0e5cbf0be004b24082446705e8cc73
zc54ad5eeec070a76db96ff523ad2f4d8f50e7b38244f5e6eae0cd513746faca0d7abffdf973184
za48071885868d65c87ab8bd9a19bb1f6ebc7d064fa2910b1a125419751842906a9d91210913e5c
z081738dc3284762606f20ceb638dc45ad20ad66d74f43b228aadeb90433b59335eb37b88f29348
ze1e58b5d02280c8178af447ba4b18499d7b56dd3c82f5e751a72c094233c034aeeb03837c9d24a
z16b705f875e295c47b8720f60450e6a13e9a1e7d6c78ad41a4b82604937dba0efd976e2b0f19c8
z11f7c902f20a6cbf5728401b9af3885c1b2beb25185e7cb943587c5b0058917f2139acbb41ff07
z0ebaa3f2507a99d271e12165376f2ba84a28228b14cb2b631495756f64a0b3080c8a78b67c1598
z8871a22d6e1b625db0d0759e1b3fa5a665dc9ccb58256c039c571cfbbced84ce8ea047e5c3f9ad
zf545465048b475b04b0d7dcca6a6c1c43c633044657a96ee6ff0384b38d6e3d1b974784675d201
z4d2c0ff8765585b759bf391d58e366caca39218f963f0ef6ddf8769ae68f9d7ff1a61d84bbceee
z1f1bdd7b243b5092127103fac81739649cce4f47ea9cee8b42ac762929ad36c9c33f8687303167
z9bb6e198a50b0260c2e420c32b7c4b4ecaba957c191d12a1779de29424916a1204955132232f0f
zbd3ca6c49f86081b11b924b0f811faddea5f6c5d082e15734058e477e88a2570a4c76eb359c660
ze48a9f5cc724f0f43246519a1b204c1bf5543efc4e73e398e5f15571eae8aa138cae988382508d
z59f72226c06aac3d7050cf19627edf56fdcb7bd4700ceadc3e5f4e0212b1b402187ddee4353e74
z937518e7c53266c89110cc71b06327a69705695fe316859c5d8ad1e924ac044b0fb6b0c52208fb
zf22bf59b4c595d6cd9448b5262ae5259f0439d5fb4e86811bfaf0c7fc039291fd32f031a088d4f
z9f40c18be1a4d87ae9540f313871b32274987d214d06ec4cacd2e533e944118631f70757e0e737
zb17b7a17f6f5a2be1408f5184eae1908e4e18314a70f56004131dcbefbc006c2ddb25930f27357
z80421b4a47f5689fcf9919e8bba8d7b6c37c96bbc4a4c4f8b7a0c8842bc9ff5a5eb58228335a35
zc75909cf4a34426e1db1a41d712d1ec9cd2e084a23ad68b390772cd64ada630109596481be23f2
za2bc57be5bca387d44c8fe00bb15382dbe27334dc635ce0295b22358528ed7c93f329ac3f9628f
z958cf43a3ac3dfc72e86daa100b32226364fe8803a59a2d26910c553dc1a6bd098e08a6ed0a0a1
z067efa533db2080070e0ceb978bdd9278441e94b16bf40d2fdcfc721a06decb5f4182d9e70f0a8
z7b41db139ec1e8864f1e242f095c4232004ab7ef8d4c0eb726abc14b11bd2dc758bafd8eae3067
zf859adfbc6560847763ddaeac3eabaa5614e876fb56c7f079a954c7dd60317196d199b6714bec8
z87b7995a1796e304c81707f6ace3e7630c9d3063b8b0ccfbddeaf503553d38f3a9f1ea417cb453
za4f2829b6a9852cb5ba4882fbacf5ca83d803811d4ca2001d01a37b5aae10af0fd25cdb2c55e0e
z066ff6bb2c2895c7c57e9a7ea45c0ab3354b69154c750241157a64032a0143a8d9f58aa6afdfc9
ze630659999245eaad731228bf1e6571dc5c06c8ab6666a78e6205e6adcf6926277f9708bcf5228
z6a64c1ff6577a4e103b45cbe70cc22157eb00d39ef2394c606072507755d30aeb621f913465d04
zf28611bc699d9527610b6ec1478a19cc0715f3b2f16b8b21b4d7991a4fef678ac3e18f1df28f39
ze55f3b0cff58f99a019204440637b20c4c0c62560f4643faa1fc119eb078f735c07085e11cf3f9
z21d28acd9ad191548aea910e42e26dec20314e664ee28c215730db64de516499f323d70e97cda9
za48e5faa6ded7419813552bd7492856c9b570171dfbce3e41ea394dcf413d95ff38cb4f81e1455
z866eb358f38f85fe5886defdde9f8caccca5cd1c827d1b7c76e6aee23b907c6db04ce9b5d50405
zdee104564c5bacb39cdfc1981ea53141b458722acfe2bb67b750d32d2ffe4bbe6bf66a414e3f29
z15cc5df6227ab09ce5894a45862ed161cd8bccf3a8b593b65d24f579d3f025d50e4617b54f7f6a
zfc589a68df06b85555ddddf4eb28093a5bc04c1464d1a90d01066f6b556ce1e039124d4ac841bd
z33ee779c0ee5b219d32431f9e3e54fcf25d74bc3e2b7889944f522ad7699a9672e48baa7e7e284
zea156dfd3c6f51e2a969d258509047e3866b092a535592051944d065fd3448fb86c883dee6758a
z514a5875a01765f886bb6c07c6b04114035a657d43969e16d2cbf3eff484d9b2ceb7c500e2a133
zf4557f9419ecc306ee335214dab5cb3eaf63121d31f861e73ee0232c2ea5f534488870954fb13b
z8c2a824ce13c2d7c0f2e36e853780c89578229054f16b47b9e66ea329bf007df1d876eafe4ad0e
z3ce27664afe868409b5bdb51874326efe2a43cff573d95ef5aba84c628aba9bfb9beb928ee4ce6
z6b1bf1e7c29d15e9d39be45f7f53f7cf95add0e3013145ac44f9b183f21996546351834354cedb
za5610260664e8e19387bffcb1e752525af1be3f2e158b0df4c39e617933be01df584cbf94bdfc7
z5e0ec0e6727fcf4a2ca42fcb28d114aa0708434892115f7d375a18f334b09ea1f84836e4466703
z252d2b563e516d5167b609915003cb4400e2bbfc2d19712ce0551f565d37802d033e974976f609
ze355b26078b574718377263fe4a7e17f99dcb3c0e54740b531d11489b581d383901b0db2459e7a
ze279aaf0308e5f31cf6cb0a0befdf789ae17f8430b4868a5076bffda082de875bbc3c55ec913fa
ze1675e468997b04e91875098b937cb86ff88336455df252ebd848738ecdd002b385000a7f59550
z58e48bc3c2cae0f95d7ec6dbf4d4e22ff569dc624d4ecd2fea0068907ce97bb032fdd11ca5d08d
z0ca21e3acfe687d399d5ef2a8c35de788c32d76f3fa08ae4bf0c25c3131377acdb98c71a5f0140
z6b55e6b812ea1e4ca75db9205982db6b47c7b3cdb539827cf337de2c3559af7a9df4c903006914
zed26367f2bd58811a4b2d534771ab1173b13ef9ca7a37367970854170b2cd41b187bd2fb8b51c2
z5ddebc399e2b327e0df074a2f7be4c5a61ddae6c52e85ac06a3004a0e5aeb685757c9c6e9b931e
z6ca3d2f42aa473a54a6bcd568af155ed30e1718bbeb30de7eb7de1ca5a4e2e19c7a23f0ec0dd34
z6fcfb6e35fa69c77dc5739f9957e25272dda9464bf365ebb9d5d99b528de68dac6c4a842dcb3bc
zabe98af64f58447934294bb2736541a456d19f5df1ab22190ba704c2dd6f1ba24ffe3920b843d3
z0c9d8ab98c0c080fd88a6f18fb9cfeb9064d5b3d605898dbcb99af6fb19ffe44db861036f7481f
zd452ff54d173e95dc3547592675197e065c5bfa531503c6d641997e52706bbd546de65dc7313a1
z0109a095c41147d6e611444d653e833b5f4ff2d30a13e78fafcae1bc5e4f79552670e759d5beeb
z0f0c9d6beb1d8f1f5faae543c66fedf345b9a083b007a582aa7b03c94023ed6a0924ebb77e40f7
z786158c9937bfa5f72036fd2665bc36237521334902017e17f8f4f465fc1137543c0e0246cea17
z67cdf8ac682e976b8996e172fc2347c03c568ede31e941245d78a129085d7b516d0b04e47c4749
z4e9b585508f2bb6e7872aa8d9d56998386bf53f2953d24f18fe4420dab5e91e844bb14df3eb486
zb37a06c606982a095f88711eed7f46fa2284d5c33497d267e5a8ff6e1ed3dcba9419e4192bf80f
z679cb6e8502800960e8536721fa0163e9ce21d7597bd550c9c062df90182e471acf02fab965069
z3d60a706bddfbd6e7037c2a0380362f195c907d088269b1a661091e857435bb5297a9e81f3302c
zdeea89dc8b00187bf6e2088450b934b90ea7ae17f2598dc7a87e6613f56476f0faa7b30391312e
z157e180d287a3d028c598549455d740b63ba07137eeed70f65adc7ffcc7b29eda3182143bcbc59
za8a6744f555a121bbf2494750e86d384a0142df200378866b3005487c1da06f97f6e67d1635799
zdcd0f5243d3a596be2fcab839df157656673e36c039088b2702bc1dccabe1c093f7dc04830c4ae
z817c821a1454a6dcd6013ac1ac67284cea0282b0f47d84e0b558d62b6d9d8b93ef4893d240d8d6
z94ca05c236abf3ea1bae2ac79c23a7962875e92005ee68c783805dcaf81eb806bcdbaa83805fa1
z27fe5651a42d290a27f683d63df0aab0d6f56e1b1e27559519213f0301454650c4466061d19c22
z3de62840ff87a51da09214cc5ef4995468b0d8ff21e8ef7c3d8328d97226c2cd93aa0b9e2727f6
z4dfd3b1facb08eac1daf1299d23d7506e8f46188e509403e04efe41d933dd8c2576f48efd890da
z0c6e4a399e64b1540c38a690b13b122d7a85c9e3d3f9d4ea6df0ed816c05f5af90f835c9f017af
z68b0c603d8a1267390033bba3bcb51e7d3f56c82a27a5cfbe6cb64d12632290716f9a732d6e162
ze9b103537b51466c72ed782f0b118a4da0f27e1e3bacef83f7d748462f46961abcb6ba4e6ada24
z4e8f533fe09f1ddd8ba1c60597bdf1f7cf3f0643e1dc8f2b6e31bd86102373cfc810f3cd382063
z1c121c7e19bd61610efaeda9d1c9fccc32135efd44fd173f4dc3aa038621e4138c53c245f4603e
zbd99ac134e6fa0c5d610d656ae908676e7bac93c6291833f68feb78ca6ff54a8896da9b394353a
z9223e69432de7fc4cc409302df5e324d9142135efa211e07a562fb842d94866ad20165425a3be9
z6db0c73fe0b9c07392c27f02acfe145a7c4b96f39a91b0e145882976eab55ae562b6a83f38e9e9
z6f5730e8f835dc5e400c7eb8217cb982d8b5fb6bd2051e20ddf87c99c802e8c138d087bae33d9c
z6b5f85cf0d2b4084e1071fcfc64ce86ea5120faae5c5d163e01a31cbbfc35a44c405675546199c
zbec5706ee83f05fa3ff3aa3df22397333508948ea926881c203b9d9619b71a4d633eab4bc293b1
z12088b553c9fee2043f2a298546043d65797ddf7c92f1f8f28e9cadca8b91fcbbc543444290155
zc6e17947f5aa6bef8980c825fe4783778768adba59a14e2af7b88040480d7105ab6fa9dd7751d0
z04439e9e976101065f729de09ab09d750104a6c43de74f94173c62fa3556532c0ebf5c8564517e
zfdf44a03032ddc46e7044d6cf9a766302adead2d0341e6be1c367d45c60520bf1496a0f7caf5b2
zfa23e99e68809126d5e2dc5bfb4ffc1b8a12963b4e620bae8849e4fa943a7eef0028a7735478f7
z653f65a21be38e370d091f1befdaae0bcf9e9ab2b5187167e1031b2b5e1059e5f47e8f8d5a4e62
z826f88d68f24894490409f67d77958914423efecb8d6eeba61fe6794da98e8ab5c0a988bb8f46a
ze0107e197bbe574d190b14ac096b6c86aaea9562d495ccf6a7d45f19bd227261051842119bf8c9
z5f89214e0ac6ef2ecaab4be0e7e7db12fd2397f692f2b977a12724de5b9b58f726ec91d28ba1c2
z4ce0498d388d9a7322ebad0c68b185ae60a58b9fe73bc1c37493795e91f55bbcaf0b46367ea5bc
z66d7d17cf955eb7ef0d55e17f424ab2be32975f61b2132ac1c2bb5660f2c5e87fa539cd34618b4
z97995415e3f7603decf261703fa6c88ef299e5bf99244384ec8dab7365cf6afe235fde589cd6fc
z714f94895ee922fb4ddcbd59d139819302c243ff077eda5346605c10beb22369e96b1b6ecb502b
z804ec6c5500530fa3a9ea3ae2205b4dbac779fcd08530e7d6cabacd78d0d5eb220ab4f2d199f00
zc7bcfddd6b217a82c5d7098abe6f3694c374daa5b576d9e40d4af07e95a039afb749eddc15fa04
z5f9e76ff7daad7b1433d0a894b7fd2a7ea8a5e25fd65f4660545efa1e6f1cda4e1e06225e3909d
zf1235482453a222025c5670a4379290a932aafcea053fb697e3ccdb097bc6d194cb6c43b49f340
zc92157ff6c0bea17d5159085f6b7d051f89489dc92aab76fa83a135edcb4965c42636b13e5ef22
z08e7b38557e3251ab6f0d4324a8608dabdf2fb0ff2e8700453e6f8888fb2d1eeea902bbfd81896
z0ff066a2080418be94ec4b560aac006e7a11dd66cbdf07fc24b472563689c2f4ceac0290455ea0
z4a8e5d2b6f4a0b7374129296ca229a1541f587b38486af56dd7c4fc2999a766ef490bb8f429a77
zaed615f9fe39dc1eea27a07f1e5a168ec429abf261b1dad8dd46a2b9c4d6c5bf07810a11088587
z17414a1b7a161d7bb93f852eb995344c05f488f4838a641a48a34b9cbb0b33d3bd56a51bfcd124
zef815230dbeb26e4e4d62b1d0a92a69c1fff3d198f76d5f4471e1c209692ef56626b8d0e1753a3
z9e514aeb6c609a6543099019b6c723fec2660f64bd7682f09105db26fcc37dbb8638f343fb9be0
z1ff8acd819862d032c02e530b3603a103f2a7f6b6c1949ec1efc2493e3fa18519bb96b950f4cde
z0f2ad5484b44481460cc4687f5077a9f480a93a48e97e1f1be5522e7ae05249f1268b3289bc216
z067932735f647fbbdd076db9370e0633e445093de165ba4f70f237579402f3b4d95fccbe07829f
z0a9f26a23c86dd9beac6a26a2fadb0b5b8dd3573db717a7943f7205d67171fb07f510b1db5d953
z5bfb2ee2e7928ce975ac7e32ca07067cd259438ab53c81f2a6fa915e56a7eada563d73ba1cb741
z56f55219d1a8827a573151bd821662cc25a8cc159c8fac6c9474378e65110410db13fb39a2fd79
z1eaa51504b98ea1026d976ee7311bb4a4845f7b1736efeedac158107be06be01751c9f71270b12
z53a7d5dc921c39a34296cb766ebea7f1227d06b2bb85cab3fbff897007b16be34c11ab519da209
z10ac0e5cee61e840a0cc103b4ef2494a19f31f4fc08aab43ed605924e4181602b19877d173058f
zf5e47775b709b453e636108b93b4d8e23372a5ef58d7f15a4a5b69907dda1d6d8fb9a6ded442cd
z985da6b7047af9087cf22c50179cc7bdec9abe60ab286d0d6aa56db455a363ca9871d0dc6670b0
z2864789f03eb940a668cd5edf710602a3224f82aff25f83616395c24ada89ae47ce964cf8a225a
z78ead8b5d8326d76cba12de507018955dd7a15cd54167962ac5e015a3134fcf9ad410795de853a
z0e3f55c3241c6643d686a04174a4a1451d6242290a89fcc36ee4acf9dfc5415b96c74d68235d43
z20d21d288e4ddf6101d87bc53cef5709affa325736d302e106475470f845d77b5255831d17c660
z13a63ac4c30c0318bb1b4ebab23b8142ab9f2b040fc62071080000a9dee537720ffa299e25421d
z9a2b838c849a6bcfc703d6d2186522db8904c699785b625c585f0880361c085768b899c14786c0
z835377ca0f0ed73d4058620365a4f4fd199648b99c846295138c6891452f67379d6b0aced7f55f
zbac807fd39ce01e054e16ecf55c787e3cd2cc0bab0094c55d68eb01d64545b03a27634326098ec
za05e590f538fa3bc0ddc71f8b286cc8db1b77e9d60c2845e8bc3c3ebac3c5978a44f7d78a553f6
z54850e9d762dc3fa116a18ba6bfb1ce4d6aeb89190b49c4b129cd4bda22f8b9a09c44906ab5659
zd05f57b0efdd088e81c36d931478b54f3328a03f6901c556e32ea4a08f145e36034fd847d1b2e9
za63d9cf76140552af53dcc3a1833fb582b362db79b0431ef7e6f8a9f3e74e22d2c478afb567af1
z97b5937fe38df14276139692e64ae740ae008e0cbec7bda28277a8c61c3a3cfc92621da53946ff
z7f1234f4a57b41a9f65aa3eab968509f6f7d4e50d7eee4ca3b507e4209f81fb8ee981a3fcfec9c
zff51c675159db1e9e961b05fb44ba0d29b05d13731cbd61d44a40f6b0761dae01ea42aeffe56b5
z4a4ad9c51d2bdf409277454f95f8ecc969871afd791bf15785f16d19393d2befb1e3c1e4c73759
z6a6780898230a5c961e95d4972330edc3c59e9d4aacc69853d2bd5033c58d946c71ddd1b1e3bb2
zd3cbf225c141e21f8e662c3d473d940e46a46df87fc52536b5e574cc0164c9e03d5f2a3a1b41b0
z4e53f7531e46921430f981956508f88ee14f10c3b819dd7ae0480a49ffef1f4f49a877a0e2f566
z8a9ee479febdcf285748873c25a9a743ff9dbba5a5ec5f3fdfb09be7dac08a4d7061c7a6f2e4b9
z12f9fc493fc4bfb9fa5869c7e3a9baf43395a45f88ec6e02f264d94664f4bf7db98f227be5728b
z42a342ca387906e2f11df62abd9fe20868344a496c66cda3ff11a80b4bf05f4acd0bbd764cff3d
z3df6640a4c2ab9248f7494edc1396e6876e83a63c284e6f7b705d9e418c4b9a43968e957786c6c
z630d5dbefcf92d3f516794fdc470c971251fac546a28d1fa10ff217574ce7ac69298b821a03035
z9b07ea86ee9b0fa30cea33de031a2166d8d9de5f7644717aa3301f415ae71e739dd0de35834d41
z7759f4af7a976f967485352fbd83dbc52c9f03d3412f033b95ef3bbc799581f2d42397af5c285e
z4b26b31a2334b560e4cf2aa4581d7756a8c06bc4919d6715aceaf8e8510dd356372c32897bcb57
z4c510335e6d61051ffd5956eae76b31903770a8d70feefda6726fd4d1e59c393a3634edfa75e35
zb5f693e50c7df69f172ae2b747e3a054216ac7133c9099ea0f73eea6f5d2a64eb3ae9dbf7a3591
z96c74b038f00d9723dafb247851b5badcbdeb05418d125cc00ad605cf73d67423a144f8f90ec04
zc02cd8ee085b0f21a18c0c5524e9cb96cb41a951708cb3296b9754d0dd67e54587e9e5371d9366
z853c667cf34c0c36705c66fc81bbe44da99c587faf93822c2218a22534bf8ab0d529240057e9c1
z5c340ea981e3231849c60da80e4cfca35ce0652e71fc4a05426c930daf3b8236d09f05d80b8742
z5223c42eda08eb02671f31cb93902fc7f28a1f8ad4abb5dca9272ba9fc5e7bc099b75638889dda
zc1b5a1b930795a9688b7af40794b4c2f8775adefd66981412ef432ce5bad0ad943c3f9c277f1e6
z9cc6b8dc0c2111326d6bbef51dbae24478c8bca7b90fdc6be8b19b1c690b71ce21e5aa86fff624
z7c5c8daa13ff3f6faadc6b8477107873f6e1821876f9669fa76f68b1edc14e931dd71fbcfc4fab
z97e0be131ccc794ca9df2dbaff2cf576197a32d3567d30b011ab7d18e59da5ae8bfa6c8de4a0c9
z9433c10da0b90e1f0a0bde6b54f28ef492bb9131652aae56a47eda9c6d962cc5f3b992219c9e44
za7727bfee31bcf382e548395f9c4badb2b6a1d7d79d09dd6e95289138baa12a634c32db79e8990
z97ddecbce3979ac5153717bf9e2c9f507c41b0632e9dffee392d8da4f421916a8c669ef5b27eb0
zecb6b9df68071969fea95ea9ca5f6969fbedbe7f75b2db44ad2e4c0b883a4544303d1e037ea7e9
zf0ae6ff2837e0bb0287b826cef3445707a4bf4d3526c6afda6990c16ceae5017a98812b109c2e3
z10decdb850ef3d2897a4874bdcc1963b8a96c49446b0cbb6621d6091fd20db4bb18c5fd353e938
z6d19ec494d4aceea76b909e309d5819bae9543c7f750e40d8abb2979751a0da57b957f4ed8867f
z1b37718a277e9a9beaf33cb6a037dfca5c819e4231dec75e72066e2a5963fcbb9b4b18b4f79867
z550372d97b853c0a14effc5c56038123aab5e528c283603a2fd61bf1b838dd2ca114e062428193
z3e51943d09d605d0dada5b5b0657786c25ecc28f2f9ca33946ad2f280ba0ad684e4491b1020a03
zafe8d4d16550cb3af9d9554a5db977ce09820577e578940c1d41af8ca783f035d978a47539a52a
z35fba76be5c5c95875e933d5e2b65342ad964094dc16da005e365bd735867e81d1a2338a3a0780
z0d15fab93de747dafbf3bdbcd60a109dabadfa14015e62450518a84d6b90e284ed514328b9d318
za23b080d126d02ef31818e796d8b9ace5e8d534f73da4c5cb19097cb9b17ebd6f820b200a2a7d1
z594166215046091286209710bc9114761be81e2199b56ab955638599015fc735cdacaf12b5a883
z69ad6c9a74ea705d02ffa2b464f67588108ff803a3cdfefae1b39312a95cc79101bfebbe9a6c8f
zae05319077d9bd73ff8d775e7721faff56af1386cb82fd47a09791599afe7cd6e59b192a995dc3
zc18d1f6784696b21f41d132008eb0df8792dda1e1d0f3dc89437eb1772c140a21891dd4058a1cf
z320373742ffcb3f3fc4304ef7901a4d23ee784529995bf606095eab23ed92b1bd9b20957faf57f
zd2689aa7f95edee710aeffe7fe9897c292c1453cc6c7fd1c9090e4bcee0f60b70e9d0546e34df3
z6c1ca2c1b1bfd26a1f849a3cf0b3f5c65a56ee205dc8f15b644aa10730b97dcdb14853dc969cf0
z16233250d45b5211eeab421b3334b502ff8b0d5176fc42f04d9100a1797e5c09482997450e2f7c
zc6c688f9dcd777706c8959ff300efb873358448f33ad04a1c1c6e52360049f2514c3c7ba6bb9e0
zaab59f811fad8a52bf4d186cead9284baf7e35def590eed3e1f7b324d9d015e9f131c360ed08e1
z7350bacad15662d770a9b58209605389c955b25dbd648f7906ce19e1d7a0158706ce632609c834
z70ddb35e773b240685cdd2ae1bedd52c7235aee163d6f799803762271ffe393a1fcb5ae3b9b9b7
zbca06d85d2d99689ee07c59a7c4bb7f9f7829843c881f05ade000c9d45de40410b56c5938b0572
ze2ced137a85e9e7bf07758824dae5d0b98ff5b14571c9e79ce89dfc58f1549999d2155ce8630df
z155cdf30077a7e50a4989ea69418d21a0a57b2dbf249eafd610268c298fefecf2d9f5c777f5c26
z35d19c9a26238ca58ffde50935950109e720d823c5e0f0ffa19e4918048b9362375d4a67fa2979
z7760b15410bbbdf8f47a465bc5a565e48b8b1b1629abe083c5aa7db1d2079e0fabcbc36f2bdd6e
z6f37a16ad22825b1b43782a3ed874cfff5e248a5a6aa2cff568c76dd4e4fad001418acd22a1868
zc2464db8914db82d8525225644810e371f18a28c6802e16c0a7bd2f2cfe2ff24ab87a7c59e68e8
za428e0fc3d9bb6fef08e4ebf5a2df23971925f13f811957c7d831d2ddd89e4c8f98229f1e0cf86
z9ae51228621823b52bd5293e8940cd23f020af162f9983753f2d6af319d8f202415a5b18b3be1a
zdac60d703ca5ecf37a21ebd367f64f53fb3b0707348133e9ff8e05e2527d8ebdb99fa3874dd62e
z92c3ee08f25453d2f51ddcdeda7487afb1aa73e25b96a27b733f986ef22c6640999be3c57bfee8
z93e7f215191887160c2011c9693887df8108850766749ec223bf6f0b5f2429f28d330c9a953b40
zbcafca5d80446ae0b85ce83f91cc773dc1180ab6ee7c7f93cebf54eb41a662bb21f0448e30d871
z39ce1eb13bda07ecccb39691c3563829a7e9a04244ddafbac849c1477ede34342134b8fcfc05fe
z37642504d1613559e3c3f7832553c2b55f9f93aba3738e0b92e4e6e22233857271b258819fe8ca
z5f4986363884075078bb3c87d678d6ae1aef48f1a74b64f77b8054f7ad4b89f12d14f5dd819683
zd3b9dd090a714176b87893322a413d538b0797b467eccf9b42dcd5bc80f2793c56f8146c973764
z09424a7f0398a0968b5ba84822328ad59bd92f294d7e324ba24947b68e87ec5c4b3fbb01092bd3
z26afc648ae6e8f11e6f9fd70e479c5a42b6d9271b82da36255db3c6a4f06f867232669911ae718
z939be0dc3505423cfbdc8cbd1362b2aee629627bffcbb3c6b54aae1d1663acd4299a2500df1be3
z75e49a7cf8785a456cc6c6f886b5d4a4eb3f42bb1fb26dea7576409f1bc1d26d9667a67f5a5dcb
zca631b172887b9076cc6ef819e36500025dae2c8306fab151fc25fb8ecb79e834fe62bd8c76b99
z3633feebc62f43f713a9d2ee5f6aef99931a4c86dd3cd2eba62ae95b42fcc5f8ac569724229eaa
z0476104cf94c6cbcd9c1e3f2fa5e750b7a878b87d1d8aff9299fcc1836d32db815d0a7543881da
zb7e97909f558077786903ae8a431ad29424fa3ffbebbc1e4fba8c7e0b0350a20ad3606fe3023e2
zdeb8e338f8fedfcba566d494f79aee0cdd63342731f0dd2bf6389ed18fa080bef38b9d3da862b0
zb33d35d1a28caeeab71c66995c88313f5e2d84ef80d5dbe6eaa3d135e30805b6e9cf0e43336a89
z2caba1e0ea060cbf947019e9f9b1fe31c5b864007cf053eea70832d35cad3f6fbd5d9a97c6c2cb
zf38fcdf327dc9b6e4ec1991aad93de400ff25f9cf0b2f2b27b71f73181b9e72a93b5a010052f4d
z88687ee77a697d9c325c50ef81b3c276799421ab29e11c12729cf3cfbd8611fc43653dbc6bc534
z0fb77ad71f30bec492fca6681403a5b39aec7faee3bbd3365f9edf55d3246ae66f6d684f8c7aac
zc684e755b6fac8478c17ee534edf0617fc6f4a0ab5311363a9b6c95136f03bfc86a9d5b15ee32b
zc1cbb76aafc87b7f6f555920386eb81721449de309dd758628166e64b67bc73c2f6791be1e05fb
z54be32b42c02ba9e56969689cbb879e1bb8e148af58b2963fcc84a17b3bc0269875a403159be44
z340d642a4130f837ca37b917e526217f981293be368390ffe22e76f3dbe2adb79640810df32905
zbc3d35289a0a691c35760783bbe1a81a8670b2f6057223679ddf2d75e6fe2cb49f385da7995e94
z2012abb297bf820f0a7ebd2b258136a7dc0ba1a4da5ee49661957725aac4cfb7896bc0c0a22161
zfcd203a4ceb81a6ac1dd2264cd227126349b05cdb39ace055030d1eaf9c61f1bb47b0eecf7ac61
z4da4541d3e7ae92d162dd208f28fc2d75f81e030e6c16b6e66c4437c9f1b92512ad486db72a7b0
z52341e7bd6ada6919f635c538a851d00bde577c3c81b7e825007c29034212c8a9ba58a614df0ab
z37c176543d027f25c22c0dbe32d74d48d2f8acd564495a447e40ba2490c22a5515f685ad68ac44
zec5664a4011cbf5172dcb29bddcf9a7fcff18efa02a2b535595d7fe298429d11396f17a04063c0
z171c7ec88a4a54949fe8bc10d6e8ce4bf121fadb57a2c6a66d20ad64c718b057d48e9d038a4ae9
z2a76c2f3f86dce27c05f11fec53422f662afb0f0736faa10b88dbcb4850d99b05a50b3151ca62d
z10543482573b94d1990a90307eb824874e4914a1ee80c0f5d984b2e32bbf309d5d56d338032630
z80ffa3170484dabfa9766d507cfb8e64bb1a6746e0e9cd7f8e97055bc69c1e72fa01559175c77d
z233fb3db07700d4227942b1fbd0ef6531b489ac6f729e04aea790ae5904471d463e8563c8ef1a8
z6616ba06da46bf93f0659cd397c59ac1ddc8bb1309e27d5ae39a40784509dbd6c37bc28e2850c0
zf20ed5d444e25160a5e19428cee4cc014b2dc9a652bc5f506d9e93fe54207ebdcc432fbd15a367
zc17ddcbe66b377d0927f6d7962cc2cca687e74b0ad6efbd478060f695193e11b7b4d2d920d96b7
z0cddb80d109ed63c81ddd6209039973e1f854eeb0b8e5174d16c10f4f0a5adf9a21c1fb2d50fc8
z06c4ba6f7615f6d72e7ee10968afa6781d55bb11433bc77e564acd3dc93d3e35835316611afdaa
z540b820051b9a7680a18fa2ab0c807d6b856d1a9d792551b7a24b622f2472f8ffd43d512602e2b
zfbf7de7f419d5ee36fdbd62cb17f49e3c9fa5b90bc23f9097c84f817a72493cfaba6b7a6bddfbc
zcf45aabfe78dd86204e6c999474a731d46d829427bb6ed4c6b228e53339d7829fe885b0297180a
za52bb4cee42bf2517f775a303c25f1bd855c6617606122528a1d7de739939784c8ddedb28cd6b6
zbf4c4a5c7857fe5e675a62ac1c55b63aae2788f34a1c4a5a8d270b585ae5bc73e77e1556acadbe
z58cac371ee84919eee3778c34dbd21eef1dc86a3b28aabacb0593f14b73b9ca990268ff738e795
z67860a1114dcfce16a3e9a8eeefab628ff7b3b0e21b59f9d4bd8a3a1b5f26893701da0f7c67920
z98c3c8bb1931b1cd086276add2c406cb09f68f7b04b3a2a8a6ae084bfad9918b6261ddd556052b
z1631ea32ee25f7ab89bfef49827d1eccbab641c33c13a9d52934cad08e0566831c849c1c9db449
z3c8e1a32e0b2679de665bbc48d504a8f40e467f42dc5f2508f117f78f4382a26c246ee81876914
z2b2511a311a91f39f493de1935964f185bc7fd771b467ce4c0e407409b6bc2fde625fbc69e1979
zeca8ad2afc6846d9d76716fbc3beefb9c97ccff21c433e7012ed5b33b0de8b5c20a717890deea0
z68bdc6ee4a560daed3b57018ef5cda5d3d6338b3589c2ab01fc20aeae351c38a1c748c9eb3e0d9
z0fdf9a4be85fb47dbde1777cd09d11aef39ce949105531ad7ce99d8e0fe2411b6ce35ba3703a2d
z52edb20d6809fd826eb12296d269de8cc906030d55650bdfb5e0a11c4fca72c0d79eb6dd8a9cf7
z051413f363dd2f37c87d1c895f74182f0035e7b9fd36be9d0cff845a681759f2aabfff1c54c672
z09f971ccba463b999d32c8aae6413838a81e9800301ae40255ad8efeeb8007323cdf1e5432c57f
z2bd3a944dd1078e0dc74f409f3d7ef2ec578c978b5b4284c17a465dee536655d0b6d82a413a5ad
zcd21328f2d7cfc3e86306e34a56e9fde7818d5c99715a80069be2d8e9163bf8ed5baffdea4ab02
zbf27420aaaf13ab33d6fc865f5b7006a505b286473fe3584d39bfa4cd8c8943ac7461a9064e39f
z892373cb9d86682ab5a55e9816cd462d34b1bc64b346917a575c10bade7ad4517a751143e6350d
zc26ef28080f3f420b5f88ab0130875b0b70204f565efd82e55b3df9b161879511918b1287d0a07
z2bd99f4ddb8911ca66698be24a1830859a098d9de5f9b40aca1aaef2cb247e542513f29cbd0e95
z9878083144c35e7d759b05e5fa6adbb2effd5a72af340a702502fcde0eadd280b67bb54cc3388a
z44a2a69b20bfe12ade35eb92ff53f094e985aa4c7e0200639cb01c455b7614bcf8292a06860e5f
zd8a00f8d4671ae07cffecbb3245c7841bf098a23f98f8401e06c1bbacd10e39bbf0c30ba1c42e1
zc8526b29fce4b636d3c694a4113a467bba8b5f087e9ad844e7e8eb7c3d40b64f09bfcc0207a2fa
z61fc16456a2338e2adc7ebc34557056c8dedca571c9cd9a0bae25e09eee7f0e925bbf4d18a3882
z7163843df425859dd28a2ea923e074b5ec30b6ac4b2f1d2eeb3c8709344047bb7e76b641c93390
zb655c09b3e8f35adf910cd01407db497398fe1090d6ee8b50582d3329ef633253e63e3bd4c23a4
z7e40cd35b5fb2f369bb1044b877bbcfb2146fcf9944a5699988be011de7b2795bfc8accce3f9ee
z793eadd35466949efb2a33a9afc05591a393c09f7a84fe4fba703bf527a5fc972eb4845e62fefb
ze63f0af51351e8b6e1119740e951a438cafa49cd3371469f454a2e0a072a7afcf65d72192c978f
zefdd3b3efdfdfc604a609fceed7c33c254e69fea1bdecf359ddcf7d3ec435d7112cdd7f8353502
zbb6a059d128a637cf19fe3acc1b112b19820fa184028bf6e2eefae7f922a388246dacee8233b81
zef5885012e37dc98da0ea899de26738d266a7c7137c329875be376def2c4880955647af6c77cc5
za58045ccc9f45914528608aa23bf35f14b922fc62ee57cdf25d20e5210b2003d3a06d4920092ad
z2e49198903a919017e4a138e464a683b3663a145e6ac2531ad02ed889fe8f75af4bac56f3ecae5
zb59554695ef743501859c6dffff85463f0d1b47ff432720548b0c41e56398ece0993beaa540d47
z7cced13c3881959e236e55c5e2726447c08ab23f69d03c1c85a0bb85741e30b36cb4975f656398
z34269283afe37ad6aed322cb1befbde678f1e8339c2e8355ce4d8bc8233f3a2369de97ac9017bc
z140be8f929238ca7cd3d546af652c08c94de7229c883c0970102fdc3debdce56a22502c3cb2c48
ze84e1de97ea8ccdf239fe3b0ad69d62a7234e01a00557baa79fa41c846e0c4d064a7635642d3f7
z55240b467b68bf81d78497f9a0d827070ea142ede01ffc604e223e899ba74e1348a156c946dc48
z0660128fa791c375321ee0f46e3f88f0874cde1f73232dd6c8d154c042097a093518ccc0fe9b4e
z2ab2ed8c478e9368edcb5f5384548150b103b23beaea8fe3386a164f6e6537f8b81f2a1f75e1b9
zb82308893677cf72f88472d6b6053dff5b8b022d6a550b8b12f01dd2d4a87ac2c0736c8b57dd3e
z79ed76611c67aed475c02138ab26f5f6f4e3cfa41fd8da88e28c47797c2bfb32a70877801594da
z653936ec44df0d0bbd461ab7ef48df2f7fc4cbc55919e4da8d39915bfdcbce0c50b74cdedda15e
z2235546da9a7ef36e20d0385d799a62aa5a7666d586803a814139457130704c3a6f7f4315cf0c9
z4e2ae1c996fa6a5f8114ad47249e7664d97d0e9857d90ca0f1ff6fcd160b136cd1cc30f4124822
z790d82b3f58f8a6bd715fd5aa9fa97160e0e16ec4f58337fe93870486016438c8e13485ec24938
zb124fd794786ebc092a97159c52c89653d818b468da795542b29d165bec090f882f8cc150da1b8
z77e9846f3c3ecaa1d34ce01660f6bd48fc47437a2790f49af029b590ff5abcbe1a80690c403cde
zaa256cd273199d18c09470743d472d25d9681d87e4dfe1a9ee3a2730a797cca8ec400cb0eb03be
z9f3cbcf626aa5bae26f447e036e260ecaa8b313eaaa81e7e18f4cadb45397f527a9e18af681003
zfb6474b369d1842f6a78d234aa5aa446ed053bacf1ae30e7238d1bb5a290abc73050f5fbe8528a
zfce05332c35e7ad463bfdd81748c46945594cab7d23d76e34a528061b38c49c6160e1f83eb9e02
z4d7771e4090a18366c4d334ee9e6d8c9440a4e6da16d1d30405d9e61d1cd2604bd10432bb89ee7
z36feea7d1659bad107146a0beffae0566d8cb05d7639d2630ecde70c456f4671cb28399176b765
zf66695aa84700c706e3a714c1385f0a6770d013ca424c5693983e95a36b3027c47a245d8e1ad1a
z930bd94c2503030db8a0d108c821e2b51414e9f1aff16994a52705f91a8cd75753c1c4f635cbc6
z4734ffcbd304442567c36e1af4d6b0a5fd999c504729ba8311bb3a9ae4b97321e9baec25256609
ze89bc573a72d456c54c0c31568e019ba723cdd1417680b1a2234caa68f9a2c2dcdc0aa46a2ff11
z457d77349376161697e588ecde4b58af7e2a90e2a7bcc02c53bc8f624c164237a528926b717a3e
z8d905bb40fb290ab9c1ea66f43ee2f0341b388f9d668c14455c158df13301d9522c0c3333ff3d3
z75a0da7e9f2758dcfbb40dfb2a5a8eff1a02b996f01d13297b36f0302bdde760ac78ee5bfe5c96
zdcfaccfdfdf8705d0b7803ce4b5712407e1fcf61ce36cccb6f42330534e92858d1cc510cfb7969
zc631bf89127ea620942fd3584b46c8bc196c65c5b0ab235fac703ddffbd8bb5cf90a8cfcaf8dc8
zc7327952641cffa543bf54073cddf4c2303b159afba06c5f56a9a0a6062a9287372ee6967f19eb
z6006e44e528dcb975625896a63b3c58e6ad6c45edefd494ada6f2b09cea19686cdadaf7b13877c
z0bdd4e3f417071f40558fd7213a30a7829f7d1ab21dd193d9ae9ed8a6f8325384dcce93c85db8d
z0835ece9d6521650c29d93f0f6832fb3c268e4f7366b858cb2d60c3070a0e10b3c9e4e246031ce
zbe4c7ad0bdf328e3d6caa151685b68629ef7010833c3edb6c4fc326cc785b45d39b434ccd2c968
z2f01702b21f1cb221e7234a43b44198c52759dd3e7d70a089022ba2b792b59af9e2b54c634847e
zf4c741ca46af4cce50f41993a314a914b2b2e6e14d252246895d81efead3083025249b0c97478b
z90c6926af15a8f6675ad9b08f76d5695534786fbbd4afd4fe83d485282bed9d885edd84c5b2932
z7ef5f5a2827c410677f0e0fb409196d936b7159de8d3366d016b45461dcb2d0a38a0f48f3ffc1c
z4cf6d05b3a540db559b50c9db8e88f0ce781ee887bd07394bcc71c7970cf413ec8ffa9737a6e77
z422559cde47de33259f51ea46ac647462578056fbe287a17bb923360263fc9dc2712ff90f7822b
z578fe2ef1f22e73b8604fe66e3d8ca9f945e9150c6236b6b68448fd18efd0349e20da8a94b059e
zad5a15eeb16c785a32e626a9134cae0022f2279839167263e07c7e7ebcbe1109f4ba768567eed4
zfae5d75c0b90e1e5737bcb7734765cf3d8909da9e8f16e221562d98117523743535a111270a523
zc2d245f10a59676647b152b3faf185630e3544c599a5a9039cce9ccdaa16419bcaf188aaf8aba3
z24e78a2aeb8a90808b4ed624fb7cdd2096f396a70c27ae6f119d5b5bd334e3506008d7b595a36d
zbca09fcdca2fcddf1b7a107b5f0e929279b82bda7acf31c57bf245612393f058863edb96be10b5
z4aa6b746edb1d14e0c0cc113daa73b63fe816638aa583fe33b1cc8e94e1564c7eeab37e366f180
z7f9bda5bcad695d9c51ab5c4b04b01a7c25f7affd71c5d312dc9347ad9e7c02fdb570ecf286040
z3094771826d04bff4caf2da50b1bc22ccc46cf95ef631c4d94649f15c8997ff26856ae024e39fa
z6b07169af73e9d2f5442cdcf6bbf9624792d1aa8bd412efaf9521a1ac697ce4653596877c14ff6
zf9ccab8167eab9c2b86dd9e01a6af3c471aa3b90c35fa619ebb6343782218ddde486315350e3e4
z786b2574801ac993218631a3e5e94d1278bcf0275497005f8e14f8af5a50c6f2a7e1ab77459051
zc8320df98a5b29b55b528ee8e40af3d8b4e4ecc2db3e2d5815748c5d7ba5ed8fdb799890cd0f46
z432784f6f140099872908da6e7b5d21071d67b5c18a13afa9aa867f23ef19902723c149747e073
zc3ddb2f7deb1a417310686337ab41ba183525eba3b39fac9b0b4cb57a1045c9b299f64989b26c1
z593fd1627eeea54786be16f2b01670b2ca7457c0a2648f63e2d2c8a4d9b1849e4dbf56f2e485cc
zba558d2f4d6cd9183473cbb0af00f266e8f6e83512d297968536fe943e318c37f38c7fb53c4662
z522a470715f4be88bf845ae3b721f6100f0cdfa48c6de35994ffdc5c19685f1aa3e8d3a73a1ce8
z27c66e3b9fcc9ef14eb0e5b3a0c2348d707b3eb5a9c4b37a706d74d970801362b2ffaa0de91d31
z55cf56e2093cb24fd29417e3fbefdddfc0390126609b58a47c01ffcbb863bd6b23451d34df3413
z120ed4f0ab583f6ec97d53aaf8fb7d7d77deb2e6d2f7c20b71c2358d04488a5153112cde94416f
z11eb238c46c6c9c45691970f84b20456b0a835e1760125da2cda9d8af70f29db1108a8ec563306
zbcfaa08f46caeed9dd6a3aea73cd59b2943dc29fb8e368b5c172bfe27d693d4b8dd08f3788f2c1
z9b5ea58de575878af2593010bee48b845417b909a1d828fe414d4054d884ba7812a138ead60e3b
ze8c39ae1351bba7feb70c6f886a93674088612ccb2dc096d89cee07291a89a25b8d841346df795
z8d6d3a165d0fe22e95817e36f917e593e9d14e172ab87b02d03d0bb3b10858347e60bd243ba56f
z40837e55ce6202a192e6fca10e7e10943399bf7c00ec362fbd6a19458c842ad47f15a4e0b70ed8
zf50cf300837c29801023d466336d9c4857d1c8f01da059f81e353663df064906468e2ed445f36c
ze107d3c2dc13e3c75916a1d9a686bd105bed154fb7128014657b8736ed5b5e0cba5ef9fa938051
z6e1ae2ff449b264ec5126c989214f13051cadfc09ad9c27e724722d6cb6389276426e3d5de018b
z039dc2d7e146f552d58a425bec317117c0cf6473ab2bca8b5733a7a5967e47c000526ba6b73388
z7bb7b86a3e74d7ca0505895eb70a92e111b3f283c2cb94620d7acfa0afbcfab3113c1f577f9cf7
zfbe6e3c4289bed8ffd4ab96a8e41c6f09a5a40f80e278b70a983cf289e98ff1e7ad02f95658316
z3e691e7543d66f0ced7c5c16c126e671a84c8ab2c93222330885d2fb4d982d21f908776ea860f4
z3e4728ccfaedf5893919131d6ab17c449026fde4bbd8aa7e2b5bf3b6cf1cafa52abae92bd2f251
z460e138cdc39c2cab9e24ef22c0c942ff228a8e3d3a0f17e7bbba852e869fa1114f2198d0726f4
zd74e5332264f881ac22943d3572bd3dce23775acf328d0f012aaddad12a5e984c0b8609ef4a718
za0ca81a700a9752098c038f4e1087fe25b046edeaf460f4d8b92523b4aba8cf72bf9bf33c4f450
z741e7204d3cafc04ef9074f1c8abfafb57f2fce5ef3fd5a856d681bfd87345d661d339d917578c
z9f0df548d0cb9850c5338b4c952f5bd1bf43d90a66f6e913547cf7559022b3f0c48f3ed94a5d0d
z01c5734c94fab0d9d2668cf3db869119883239e04357f7cd8b4cb3028abba476295d0c2ba9d559
z5abe576aa2e2b4c6113b85532030c0bd839854631f009aeb96dc40b905f09b7a673ea19387ad1e
z7de4620f1f9c0965ca3498eb0888fd8677c71ab5b5845d185a02ba44233e0491f2a5a8be228a14
z776d101a548f1e115676f74a5a91a3191aa0e5b0f19fb9517cb6bc21e44f8a7741fab81b35ff8e
z93eb6b2b17c10781ed49941ed7de0f524f0b112c746e6b77522abdb63118318ddba1f1a1ba370a
z059b1065e60515bf132b619be4389b3dc53d64f3a89f47973ca77ea1c7f2b340062fd87be56f50
z4016001011a7c6c1bb8929e18e17bb53523217ed4b5a9ad855df433d1357794eebeccbda158138
z3050b66a763bf78887254b531f684e4cf39afd3c40f4e6126c91f0d6035c4b6239c7dae9c473c1
zf1b5501b065df78406066ee59455dced9968c46db24b9aa4be96cfc35a0dc6636e6cb4116bd49d
z4ead25ef79da86a574fe5e93a52aec40f83975bca8aaf4063112ba0bc0b44c9048289902ccd7a0
z5a135d113163b2fe32823899c68e0b661cabe782de1cf33bf9afae07efaf9dc46f868ae489b432
z98e388663700697496d10ceb733889d34f09fa881fbd6e42f473d7c2824e1bdac167d429496329
zb03fb2f15e56593d95f8216ba4f986f5ee5ebeec1827f53757f6e505685aa2a60aaa34474e6d4d
z473539c9c7101b28a1292d250eff3f7a858957db6a49a0752c11a343a978023bc4947a67e16f3f
zc358cea86e9b7bb88c871f7de77e3b1555ad0aa8146672af46f176c3ad3d3022df2ca1c9510414
z1c0a846a4ae99dd8101b5d62906f6b10ef4babe394e3df9885ab2a2c0c04e6c28806c8a166833d
zed54012a61835a5934ac82564f771f4ef77a5f5eae5403936fbb98a9c5a61e3a4f2333bf5da5ed
z7e6de6421e9b859d5c8e6b5eee645b9f0e77747b7b9cffd61fbe979a07e32fbccbae96573b439c
za2faebc5a04fb08b97daf32868d4d4a77cc2282c9acf7d56bbce3157f22afa14df52e4cc722d44
z0e85cfc7ca446a79a850b67cb781ba7a4b1c1631cff4a5e453f1e02a7f16ee74e4757b675e4435
z2a65b87243a83761e05a8d30cb113cf9fdc8cdc5a20e86be58b2d14886523911ec0644d67c94e7
z8ec16a73491bc9df59f221b0f4da8f086bc6ec284949978b2bc9f6b703523f48b4356fd74c2e16
z5ff3ef0febedc62de5dc2ba1bcb251ed6ac220a5c83fc3ecb82d86ccdd5f75c9ec3dfb6d8231e2
z20e5359e8ad8bbeddd955a7a2f9dbeac5d24e664ee719c18e6a33130adf8df0ca92833b37de9c3
z00ad8b897a494abfba66912c4473db09f6af04b40b6f3afa7337f8a26d03d071deed6b9189395a
z030aba492101a2ef796849f54b40f3ef2449e51a46a71e9ea8d2aa6b4e0202981164d14ebc309b
zbb718f3b61c238e341ca231c0640998c90751a35923dbeea40f331864dc78b27f5353507e46eb5
z677172e08db3457f4fff7d88f5857f2aa4e478a2a2f9195ebc919a59e48c096088fb9a326abb6f
zc26abcc31e47b903dd5a0602c6615d554b815e60bb8a63aa55f93fb0804b8c14f4ea96880a024e
zdcec79997b410056d41f92a152ef8da50631943b965bbc86407577363acee75ed9e2e2e100b081
z3d29a9ca7704b3ab270729dde9a43e2e9301ed3d046e13cce62aee2dd509768dc45a75c3c228c0
z4a256c36019bda280ca029728263d550bbe578462b5f2248863537a8971d1d30393cb43807b0d1
z153ee878301900a26bfc42412597131e3626afce7820177a0cd2d4805f38ae2b08de24a91120de
z97477d6c65c854f13bdf9b70db13595abd860cfa9413b430b4f4e482a0a14f7a45a13af899bea9
zdc91f4f7bbd2a47ecd61fd0acb889729a640be5dafa7d00395720afecc4e2deed28b8ac1583d6a
zdeae5c378d68547fdd371cf8fa09b16f3c6d18995e69df8903f8328ed10e207ddd3f2af909a634
za2c612d176ff77ab152501c3db412bad1bd09942b29b36c2b4c69079523d56e22df6ab28f1d14c
zaa2454de3a63b4c7562bef1ca39d8571210cf1d620fbd788dccf5531cce66b833e0a6f65643004
z1be2f0b14f80cd6c721daa0bb049ba77954e5c5f49041509971eec9832c0fcf9adda2857b25384
zc1fc595dfdbfbf23f935bc6074d0dfdafe12ba70c2a19721c9c1f2c148a3cbc69d167e4a1adc59
z731bf2eba9bff17c71cc30efbb67388e471ee45090850faf59cf55fdaf9c64de1cb6b39c8e9a4d
z135d3835efb86152732287fe9f6ae2417ea89284c3331cccedb5d4d05be75b91b8da660b331e2e
z145f9482b31cba2436493c719c870eb90fcd750f63446d41297994047d6dedeae0c81519884fd5
zce608afb182564a45a1430f6731f4de68e1d244068cefb069440c89789d304d334a0c8af941a05
z42c915067d68fc2924e31aa500cfae4afa3fad73d107f9364401806fda03230ac6c148f4915bc0
z578f045f7f145ae96b5df62f0a4276cd09decefd68cb95e9b02c489b6dc49e4d7ac538078e190c
zc1c12c2ac43f2d90ad05218f8974f24b64bd8cea5c5685a213d4fe3f9b38422ad0baa50b169e27
z0b6b8243215959dc229960baaa1d7cdc5884d00e89916c8c82f077a77e8fb0d270ffd7dafb0f5a
za1bbe1d5ddc2970bef3822573d39e00f276f146ebe0b20899efd8e6959fb21c3c37c3086eabb46
z36518174cd0fa34054dbcc26097b0b62e3aa67efe5e4ffe4c0c7fec9eef1000ffe246cf7db5c0a
z310454089eb54b5adcd9851562e0b793d338530a014b9eb0f96ef39b122f566900f43fce3b5f59
zd9b91f0ea1290c8a6e3b28d918172ed9f4651e972a5f3c3a48893df9c812be2af8ce823cedd81a
zc64011a2984905964fe74ebd7a5bef2cb16381ddab5735390adbe221787d39cb2eafbf2cbd6049
zc58f7be1451462066a87f59bcc0906eaff159919ffdc1b6f83dbe882b8c39f2f6de1d467182462
z18ba801be5d6e2d305b0341d611e7d3b2aae83a9dbc40f73b87c13d0a846a5d5389aaea3f1073f
zcec7fd1606d4d4e5a2eab5dc929ec8c84a8507d817cd4b51d870e7b767c8fe56905720099faa73
zf1548b9a9a705395790d3c90b6cdf58a6c9b925306830c5e917aecc00cd2861c3776dd3b0864f9
zbed3634ca3ed1f5c1f4a777b7fdf6ac0ceec9599096c27fa3a81335531eff8c85520d26eb4a810
z9297f90c14f68816ac8bda261937cb5c5188152d6254b54c899b75e89fe17a283dea9fe6e26648
zf2706615fd359d6e8e3babdedef623c7f7d1d5217c00187ecbdb656819969fddc1cbceb98ed641
za9e579f91becee30f980233522c1db9f6926725432787cef816a0c09962259e39c1d0f0870f722
z679738973eadbadac43df4c0bb8a73e60b59932c4e9eee215be2c58b837a82930ad2ce78706200
z1dff4e761e188ac8ef8578140a1f07819c2b1c861736d7fce5a5c7cb09517b707c26bee5b433f3
z6ee94646486fcb67b5db3aef2b546876318902188f39b746d52d2288dbb12076dcddd34eb3321f
z70c129e1728b73165b60eecd6eed464ce9671301bb90cc4f080689060cc4c82a91883f4594b8c5
z9ae70c057f1ada36d6c8b975f1748988b11d8d8a3e9ad3015cac1bb50bc5adfbc02f465af4fce7
z283a9b9cce50fbff77220b64e9722c3858c62729c26d7653499e1ec5cf945e8174941cca5dfd4c
z08eecc92262041cee9293ad24822e2c504086d23645668d11980d515fc2c8bd1c299646da8eeb9
z45a36af856dc5366ea80456aa696b8ad11e9a142ee5d18524baf439da2277b874d7fc23187db66
z6066ff45f5547b5f2a87718a2860c3f1d2d1ccb0d30cc021e974df74973bc77d81ac2c57f4ff44
zbc5349628c981a86c68f8200da4937df887329fa1bf826bbc4247f596a0f389f39151a624a5487
zf00f166b86fbbbfdc86dd1407e163af8817726dabb2c9817c222dedde701d685363ca3f1890378
za7b8c3eba191b49ecc1a4797f9eb6d1776d45316b57b4296fc0b723e4f09b45cf421eed6d216d1
zfa2f6cc806495fa9174b8df1d0af046c7e168fb61ad63666681fb5b101cf024b4fbf96c959ea49
z8c8747249d1e2e70c6262085d9cefb15c6456fce7e5c77914b625eb4c017a294ec1c8cde73004e
z8801f6e4190c163be905f97549c0f4d142ff79e01da858a6a37d7a5b5d0a6beed235cba20834da
z2afc9eebf5edd89216b56434a9c0cdb01a1d7d39a18f3d8b89901866d1c4a089b9a60131a8c54e
z2a01adf6726d2af254e1adf00b46eeebb17e673a17076a79d352233f9b5da7fc6f74cf22a8ce3d
za27450b664f1f9bf4e11540a8efe1c1c026135537ce6a1361a14f6bcc33f8fabf8af8d2aa505ec
z56a926d99d6a850613ce7efe1a7adcb219ceb7bce2a5bbc8e9d56d6b1a0707828a8b275d275626
z1de3e6dcd8ff85a5e76a316e00f4018d12004cdaf3ded9ce12c6286b9fdb7062ffc118866965fd
ze6c3a3135055820d8b35503b360c2e95ef6aa650305cdd2b88e9a85e3132b88cc60b23e57fe06a
ze1e034172d299242c7e3ddc0cfeb6341ab6f0b53544b0bc393f052b08e6e744eac41ac7a1ef54e
z97b12e47e8dce48d44db8261a20f4dbed4608fadee4b0a370c42587a954834e507ef837e3eb5bb
za7e63245948cd4816458f4bde3937e67106df4563e5e58ade64b5cb8c4e86878f100f0e5b8e027
z852d949db05ca45ec079db995204eb847dd2650ec26a3b965c96cd81750e0236fba00c6e49f52e
z9c7ea8e6588fe1f76d1a39b012cbee301ac28d9667f21589d3f23a91b46985f06bf416d040379e
z8b117a1c68992d9ecda5df1e9f0777e5c8b01687323c55b5524936ff7ac0d3de17dc16b6f0c5ef
z69456a702018b86499e8b1c42b33a5ca23b645fcbc1c5a50603f6c271f80602c30e7b7bc13bebd
zec34feb7b330f4e36c59b20431e70e39ce3a3647fd4ffc7c68bb8f05143c4886026f187309c11a
z3fb8f2e37e69dcdcb810e4f1834a439341ef6a1800d3898888abd61967939c8a4db116bced0d3f
z0e58a7290da10d199bee0e0cad9d6b5ab31caf8438155c911266cd02799fc3dfcb987df91df116
z50201392fbb3081981f24ed4ff741df7af91460b65904408e4aa7a33f2409f682684b45c7d3088
zc0ee1c330c7b3aea6e036d0c263ff947e6d7b4139ecbdf884754768314681c9f7fee51dcdf6cc7
zb82902c2eb6ccdb6ab9f073347656b08d99fd95db8db085c0e08928cd8b73455945bf9990104b3
za1537f22756b7bc84ef42bd98124b25863789e19266c6548f0eb823c6887b58e3d7c3973808f61
zff441ac19ead49d01f7d8366789ab8c1bad03d231e54a5ad3df8d2792fa9682bc809a6719678ae
z7812b061da43a48e3b5ba6873ab62e3feece2735fe701ae6a3cf8bda0da6ee99c5350f01c8adbb
z3d54d9ac7459cb3248076db93d8f0d69ad514d554504cfe4b0990943ce3f61f0951348811a11f2
zf7e1710cb47891b5f6a2f3363b27afee3a27448020109e08c924c97f12fdb7625fb8a91d8cb63a
z139d81134e380409864e3d8c15e1d929d0077323140137331debf9cd4f8da660c6539686acb112
z594e89e2d87b72c9495b59e665f1a4df8e87136d9c5d648943902dd8588d3ec0dba694dd930bd0
z6d063fce838b43f009c5538867d021e75c67f6433b941f70193735d672c89f621fbd7baaedb431
z6fbbc848bb6e1c8ec22856810e0faae7e221df1ce5f543b8158d8e4618cf640c314348cdb843f9
z3c34e6e58c84f0c03ff5a608418e396981482842b71f6d98a43659941cced8c2523f3903996f59
zbc1ff26e04b3c927c226473c1f6640febfc017a17543f3e01e97ddc20b9b2b52fd3fbd160658ff
zc241342f07f677c9a28bad893b3a9d2b9f5b4a05aab76c9172d99bb2ea5bf04348db705747fcd1
zeb0ef81373c186def065ecc61e532c2d64c773c6278d2635051822190bdf82750c02a1026428be
z9a18159a1e52ab72f2b60b61a8db4f6f4b74f9bed4e5ec8e883f8b48523b936ba54914bc891491
z1b6f65eec47f4e3eb97c7a73228a2dcff5bb95d65c8cd12da758f67c32092404cf1946b7409283
zfd7f149b8191c8cc9e94153ffeb827d18f5802f507872e344c2385a1bbf737bb934f1e6354b720
z9b316d595b0330dd87081adb64a76b7439a0e66f3ea7c8802c9b18a64e0b7e282b90f49bc838b9
zd5be3bfd3cc86e24095c74784073c0e8894d00cb3efeadefdd9339f103604d3adc3ec92e550d13
z855ee83c8505d32c83d74b93de549e216c954c5f7120d01698a5de70fe9048846f46e4b5f42fce
z5569b655b4e420c527bdad64d3fe38a8f5d25b99719674001ad94a673a8328b5eec8f540a229cf
zc194b3cc246e32221059a9f91a6a7c607974c7851ffdeeee97fa96ef389c5fa092309f26598a77
z326362cdb2f78ceda4c25624769561a007036746b8a480c57ecd3f231d16426edd3f82bda81df2
zfb9a15f392c0a259c885fddf38686b7ce5cdc4d829d95fcdf28b216682855011611367cc24de46
z6b4ad470edd9b15a1f84f8fef052c0b579b5ba1da236a668befa8e444781259a994b16fe7585d4
z27fc736f0a6aa7c3972fd80f6c7668165c82281ef805c4d6546ec4cf3c5ba2e6bf5c685415f61c
zc31c529414d3420d44c9ae7a7f988f73e695dbcfa2654641480c9d93c1acf35c02fc0345becc6c
zbb366049a65d3ad1ff723b4b58a9b5f10c3f668aadccabcbc1bd195577a13eeae517d20507220a
ze368fddab34baafbae5d1259a370a6a5bc6253cf213cb880c0fbd4c651c7633e06b9ad7d220c85
zbd8d67a950344d9172a00ac031278859948977dae34416662dc61ece66c0f1a4681f23f1372572
zf8a9018f31046fabad6ae8392dc61767be526b4addf3036a2c47fd92725fcc901bfa08713405ba
z2840883f01460363836f7fdd8b93ab77f9f5e80cfe5dd693951cf10ab2bf69b628153eda03b8e3
z70931aaec4486583b90baaa200f786fa850d0dabd7de11f432f2181dd6dc4226f1c6026bb92505
z26de4e76ada0acb9f2b026830b61c26a138fd5f69d26e885add0ed3fddefb521ffa129965f4e7e
zf2a3c0e9777f93b21a6a2ac1dc1318dceb0b06fbd10cf3c1774b8327d111eaa733288dcfdd3d81
z448b7a5aaa79b9efac1db38b22277fe1b3c2f4203b75b92dc3692b78762d95ce00fbf751cbaad5
zd31317e69f624fe123524c953b100f3b69712e2d17d3352a552802de3f5a67dbbe27687cb1a188
zfebb871f2b5e194cbe2aa0398aa02908de3343282ef7441b97b62e64722e3fa55a2784929c1d46
z77a14de4bfd898910b43b9709b67d3ee27ac1548256217c370c479b8060b8ae1431f135826dbf8
z60be2eec5e846e8468ccbbec4c1d438553bd5150667303736b1a1e3109558466cb4a29acbb4d8e
z497dbbe1aa362adf0f7261c0e87056fdf7b81270c25b48724c4291784f1ae2fe9c24943268cbac
z1815f9c2ce94af09ece393e9c3c88288e44659ce72cc13fa380425189281fd586cbc8a73c4c8c6
ze077c6ee33e20b08bc00d22721385201a7ad9fe04e2223b9b93b7ef535836a95558221900a982d
ze03790bbdcb42466ec36905dbef41e67ea26903476f422993a04a133c6cf2faf678ba7ecab57c2
zce537ecb5f1d5f50b7594cfd3ad2ffb647af46feecc06244d2e49c4a3743fe91c81511097b24a6
zfa15a8ff8e34c44a254a98b9ad3c0e1a00ed0b214e8d1a175459cb603c7839d1d022fab749cdf4
zc68f28bdec682bab0d6ca09c3aa4195dcb2a3142039b2256495acc401e705de14ee78519cb32f2
z9a83eca4691b6ed2a607579b05b0419da84119f8bce4e0b53c6633bb6bff88b12400cfe7ed8890
za9b75dba8a83f5361974d1a8f7d16db402975750291e7ece6c2928d5ba0a43a5d931cc2e68ed69
zcb2413286d424beaca352f8c32cd1e1ce161a65b870ad06b17c1d06eb0a853805fed5b722e0de5
zc51ae62f285e178140826174b8155c42a5469e18b40e53663b5abdd0990638afaae91f2dc92d93
z981c2e9ea6a9a41288b499c231f60dae533dbb4ac383a21baee2341a6162b4bc48871357ef106d
z59fc1d6446d5899723e49d1b85760148d82d875c00ba08a88b9ce9b3aaca7e1feff74bab67d4b9
zdd8bea8661cc1f99f2a408cd70b15b802ca97c3a70670448bc85b82ddeb713ca5dd482d6e699c6
z7e8585b7ddc9e394b7caa14cb797d3674ec07bae7215b2da43d8495ceaee47561af4b8ad2e25c0
z89683282ba394efa23c80bebeebb992b7aeeaf3e94e27512d1267e4ddedf0af73383a5115e83ee
z7cdfed1d878fc9c0e6ecbab34acabc0bf28a160ce88503bba17620bd88db2002cb3e3786b69fee
z994f2ff62179df3637b462d659fa2e6496f16424f540da067ed3f93de6d2d9cf05c3d57dfe4c90
z3875072c2be7a0e43726c1c602756402f9284c3e2a1a449284fb5484a0db59a4164e474fed43c0
z5742cd5df8adbefed30f44adcbbed2cdbd56be096d2b30f7593ae73ddc8c1f3e5d6c15287f6af9
z6e224f64aec7e2c93e3f2da87fadf6087a118ec51396f4d570a00bd6facba66e1daccb00978084
z26c8d2a8da129a0fe4ab4a2748724ad766d651bcb6b671912954c1c28dbd64b5aa946c8f26c9cf
z47c715c60c811b9c2301d2fe8d4117cba61f90edd46a4578359813fc4b854098fcde5e5108cd5b
zb8656cc0b3dfd4ca20bc27f36579bea2bbfa483dccc10e32f84de51f142cd9d266233f21fd58c6
zb8c10b6503ca61bf2f5295b369cbf98b5487b22c860f36c1195d8d5cdc5281beb99957f3fb759b
zef3432479b0a764c548641f38207be519aae40ae9467d8e956bb851fab4e27bab4a3b5267822d3
z9b12be7c005d26245e2514547e33f8daa68a32e56ef98a7a0fc80239a73604aa6d1c5600737053
z9cd1e89ada2c0b9e8bd0a85e467b172b8ee5e6170e4d06064e046948c7d4a8bdf28f68df1ac85d
z96e701eb2ac690e22351c5eec3ba5e6bc688e90406e0ab000ef1d767f862df5ead0adadf794183
z3255ef2d7e2b1d53a84c1508a5d83ca39fcaeff59d58979223f24adc3e5bbfc93e00a2612aaeca
zd3418a85d096f06961d10b2faa403ab4ad083bc0efcaa1a6335bd505d132ca7db2dd43e8d67b7e
z0c8eef55847c580866e4dd61bd0fb17cf47a5188aaeba37213f7cee58a7ed32c70e482276539b4
zb7ce4e1725e999e8861b903c7f710e07b9b0bc60ec50fbfedbc1b63dcc0330ba09a65d50ae1494
ze95d08aca5e076f46bda234866fac928689f4abfcebd3cc74e0876d7e55754e2a9b9ae9f479a65
ze2d7bbaaec358302b2cf2470b41f7ed95209c9f701addad660496c29ccbd3d748e87ad416b3d53
ze15878d76c1458e583b0fbcdd1fa20bb5dc9db39f11efe98115824b675ca86442ae4465badcb6c
zf6102d212afbc3e6179300c9e1aa4bb12c5ecf5225285024689b74be4feb7660baa84a84a9ebc7
z7db09f6eac07142f48a65a6ed7b18c32c944224a088491875874574af1eb229d503b7424a61181
z3e2bd81d595d362b135895802b2d5ed979dca61ca9a81454b76e078ce0a3f1da1ef0cf1431c65c
z5e35b07b5ddf89d159fe9b2c4d30f324a5227f0123b3533ad7537d5b61f0a57e786141aa1d3d90
za2fef6d122d9371bdbcabcb81887b10df548d28bbecbcd23daa13fc6cd8e5567a1bb016e7dd42b
za8555575574f122433a4387a9cd6e15de923200b78c2e45a82eb972d0a59dae53589b334adc471
zedf66be4e8f9d04b60d00815a68bd1cb0800c86f49b507a0c32686873b9aa20a540083d7c41ef4
za54b050543f7876897dbe5e49c9dce3b0e01c4db8e00bd6d0ff97cb54c61418468794ba3c3357c
zab079502aec55a02767d8f7da1e93ff6f442c5b624d54324295ca950b69f63461bf71fc4e67bc8
zf2820350e72defd19900994931e913fb4a1441965bcf378196bc5f2b1e9897033c15b2afd0dfc7
z8c24de609459b944100f35b9e895a43128696277eb8153746cb3979f2b308b5ca57f2008570c46
z4f8d750b0d6597de18fca309ade0cc06300f75d40a71bf82b60428998d722a3f1df55c46f71fd4
zdc759d468b67e04a653bdb76f04496cee075f73f9089589dbea77415c52a3c0fbcf5142fc0ed5a
z63ddfbd6f42a91faa907af136341c36c2186373213b0d94c8785855a8f1824ec268b74dc505d27
z5efe6a5cb2f769f6fdfe596a29e0eb4f53a8bc64254878142bda6bb97cf4d7f35e1b788110b850
za6df2f73dc79324ceda4d44d732a13d097c0e38e72fd9ad6031fbbabac6663df12253f1222a221
z9296580167b07d4133f66badd44d7831ebef732918521229a67542af045454e5d3b421d9a10464
z163985965ab9b6ca5cc76e6a835fc45162a08cbfa5bbb53b536162fd5d4ccb9dc279d47b9eaad3
z1e57f3c577072be7b80e492d581a818b0d9e37840a6bc20f1b6e735e23813565712c69b6776d8f
zf46e3474b58c33e9c25cfb24571cd85af56eaf865e15fda99a61f5421ed854209a26f8d4f4c8c5
zca184edfe1384bed2df3a610b70604e61a94afd7edf4624312a17e48a94048e8a8765f309126aa
zcc97825d6f4a597d5db9386596c279993803f087051f40c7f12d42b42e042167cb9d5a9c90387c
z6b2fb79fd365d48b83569e3606f189eaed02103229c53db933f37b529abccee2e8c1783792fa21
z1059ff778b5ff86e0c1c9feb1176b5c8d74091bb6259ebf19a246acb83ba00877f249764a0a3ff
zb079ebd486d613c0808e714cfbf38ec389e41c6e0aaa32d15b279c5554d2b27e320fb31d140352
zdcc9a02e9ae2bbc780f5bbdb9e5a3ffac127491493ade9599954093861b7e5f45ee74d8b36fe37
zb1b3e46985bbfdfb82b5aab5a1999b3a0dd19eee1a495e59260b474c038b5da28e4257ecf3953f
zf25a04d214850344f6184907d98fafab7a0009efc483dbc7b4f24bb52c3a9dd2f2277697a1be26
zdc1eecbb81a67aa54c9b847f1d8dfaa9933444607553781f1aebb5896f3c74facf8af708ac286c
z231f405e0baaaf15aed88df20de7840b9badcddeb66244e6baf9b9181e74427ae81970a42e93c4
z8a5bebb2bc5eb515e4a71eebd4a40ee434463eee529b3126f0dd6c5fac3412f2f02f789f1626d6
z194673717e0623320f58bec5c4728a6001e666ec185b6cceaa54dc1c3f4da90c712db64bf3dbf1
z0992543a68c68e5e9a7993f0ce488f488258a2b4324597a1921337ab8cc043f3ff459b5871ccab
zf1c7dd87e082b075f746075a9763484be4f8c9ee4481270b94f0db8726facc6795c0610699eaeb
z3fdb7e35f90f80127825a1ff4ba741ea7b181327d6a80815e6cbdc56116abf9fb5fa7ac5518471
zc53300cd3f44b891fc1e860cb00a5e610c3ddba2c81026d629a754188fa6d2fda8389d313892d3
za11eb6bd68960c538417bc6b300ad1203c6520691b0583f64a8b54456db316cb01fad3a6128b8b
zd5c2d6808aa0a5f7b7671a5257dc09c3a9b7b612696b9641dace57e4850811fb0780d8a88c9f0a
z5b7a240f5dc98cde4e7c7c9e9b3afc1dbd24ae33f6f8727a7527214edaf1dc0185699ab3793fe1
z4af09f3abe55c81a99103339ec1c4c8b6381dfb8f50a886b146dc9540015d6d1aedd0d702fe8db
zf09125965e9d8f808f01c9ecba0d9a57c34372171382bf2fcbd9db278f1f9798bbd46e739b0147
zb00c0513e4180010b199c166df0ecb246e7398b6af6e6ff75d900eb22bcd9ed34f53286af36310
z67d089c6c28eaefce14cb38e9a0e58a9284f433c071788133638bc88c68a9a5fb4c4a80d436be7
z37e84e0c477dcf263c26cfe8b4a6976748aa195b222e4582bad81437f38d054429fa22fe466442
zc4599861e219783d064c047ecfefd1051297bf21903db98d345784ed7a7c21d3936d457d393edb
z206ceaa3b38a97efa0fa5a326100bf1a006e1356c322e57354f883c39a9ef7f9673c696edefaea
z64c2defc8383eee332ad121fcd1e214289f1ceaac6b76539e9e9a999338816fe514c45c3dc7fe3
zf66f3d12b9451057d7444b53c7268c5c0c23309cfee043f6fb78571ba8eb0e8a6da37e78822ecc
zfeaa1d4f5289d0f021c19131f8dff6601b4fc389330f5ea232317c2bc9e069aa7e611b2e953968
z9f86f84cc2e979f89b81f2fb45cfd6482af99fcee71a8c0f1fd745a9b20543ac8c070e2e984c75
zf3e0320e0d48a0efc74df0f7c8d61ff38a694bd9ea3b62dcb1a9d6468443ee4a4a6fc7002a6b35
z7baa0c5c0269a4238a275bc3e3d8eb6b8e332695b34cba19668ca2bc6ca554048bd9ad224bf623
z41b4e881f8782f28a0b960e888b4300c70292d38156cdafde825acfb4aca9080d20cf960a0bf62
zbfa42207313f81154f7caf532e6096e207f4d3663267b4c66a651d5fc933a628676061eb297a79
z92f9b1925003f1e407384a4463a788fcc80537531198d8f3b6a408230e573948473fa3cc9422a8
z570ba1de55b23b2dcc3877e88e45d2f582aac4d06a2f5e5bedd0416d9e33151344e4381415917e
zbea63accd98742402f53d156d4bc9f66d4599c4cb272e429b91e3e5a245b88baf9e837acc6d533
zd79f953e7481d07501a0dced808b972fb22c00e0abe057f3402b0bc327696780ee8ee63e5ebd93
zc4342f2b499f17190aaf9607a9e7b6f28dd5a3381a1c69c28ce70d7ac7c746526b4ddcceaf428a
z51ab6f3f9b1ff417c1d5b6ede99187069a2bc4d08dad3ee5e6336c7a904d7f8eea9f14b05cd1d1
z5b7464fef4c183670014f80ced1cfad89d71725e3e2d24baad218f1109db4d152190a3236148ea
z00637a320b85aa4070394093fc5be48d4eb58e4c7bc04fa99715899a07ff9cb64263b96c608f58
z6aa0ac92616c7520cf9b3ebe33d414612c8d62988019db0c08ecefeedb977be767f4ec85e68e0e
z900bc790fc018847e23eaf41dede597dfea918100949ad80f473ec3ff23007f95dfacf3117f34a
z274b9886cae11a7754b21cdcffeac291231e75643eb8cb5e51d9f5389337bb4699ff805d833222
zff5ba16971f6222236c738226ba261bf737e00283332c0a6da8849b4cf96797e7cc0e4bdc2c6de
z45b409fad94899ee1828f28437601532a709055d51a0b31d3bb94b63c0a91e762fdb0c155e3f6b
z0f189cad753353744a12dff9581874bcffde5ada6e59a85711306984b99a73824fa73759ffc04c
z069b0bf5e7686af372d19771d3f483087cf2f7a3eeb4f4f1fe56610b68c03943bada1eb51b11cb
ze8939f030267a020af150381e3295736466b0cfc30f17a7baa23e29dcf8474d570c4aef2962dd9
zcef55bb160ec916f1bc48244cfa029b2efe4990bf4c871b3cb4bacd49ed487af7d1b355ce79774
ze049904799d0bb56f2e4a63a694a67dbb831d1a6da6a07feb0501066570daa0feaf8c770951db7
zb7cce1e77be365f9fdc3d5ce95b9bffb830976f1f6e369fc7cbc1e532e1fc2fc0fe8204694e266
zc12cc0e48bc412ae2a2c30375aa612d6fb7e5f9b8896525b0629684445cd992ee3deb59da72fcb
zb37d21957879cdbb89552da9c07c5e6454fdfdfe0463645e1104d4261edf140f28e105bc5b84cb
z88582ce93b6c77ab8fd8c6538ff3bd1fb9f93625cbc37084934cad0d82b0b2fdf68a9737b31256
zef42d52d04adb99eee4034ae2b326f62850e30c0dff412cbbd49e02da81691c70d354b0b88618c
z1a364d5591ebfa6ed15e9e38c9d747c5a4fa7ca9c368decac4c4c9464ae265e313bea9a263e4af
z00a2abd5bc319c9742966f6c978334210ec80b1e1747f092526aa0ff76ef05f89d94691f28df04
z7dd80d43cbe4a40dc5bc50f46831d9c201eed8dcb68a68b659ed839c073d19741a6dd6104d003c
zf0bba28c89df0826d991bbbea040c38904290dc2d448f68cd8f22e1fcc8329b62bef025b248810
z6e9041657b1794c26bba15977885612cfba2519b314c830dcd96e478fc5cb620def33198d034d9
z1649485569c9d0064fd81ddc2c7fe51e980afc9214e34801e3085e8158c5c983230e68682bb1c1
zed6dff8496d909b38c1452b79dd7aae04628f41c45711214664c2c1dd3a9970482220ee0c2c4c0
zf9a67b5a10da81ec0e60e797749f00303c4a1f3597b11f68c73a53cc76f47541eedd181ad7db28
zd8acb500d607794ed9012ee4a3b5ab91b5ba4617137010b477a45e29e87543812900002c42c606
zb1070457bb9d668d8c2f6f3dc6df242acb685d1e4dbcdec826ce3425bc0a0910adce46386ae521
zd228f205a5854aab44b56c6e0c50d4a3e64fb26e36ecf0f1afe9ddcc0ed8c09cc4e3d2b7cb8674
zae0dfb54d4d34fd2a315c2b887cbee269a663e7f153ab9a8e14807381db775b6f5f94170373dfe
z0c4a602f05124fb4ed2d27bf93659124bf02e37be1824ecc9df7dc755baa61a5118a33b83aa6bb
z1ad82a1786b02f745ca1722e492f27c5263183402db8efc568c16cdae106927b60ea9614041cd5
za4c89c34cb8cb5654c56aefc48eef21aaa7fadf92c1d0665a34c94d44f396276e4f5ada3280d97
z9bebf47108668be82027918b72dbc9b1158ccd49d77931d1673f3f645915314323ba8b64cf58f6
zef4c0ee3245937dcfb06e22efc58f5977ddae57b5e3a5859e921f6bf2977939f3d2e5ca1a94d91
z9d2ece93cdb4ec20984dd701ac8641c5abaa08fb5a5310dfb04b5b131c07c95664906a1b246e18
ze3dcfb6992321bb250d89e587cfdd0ec84fb9af55f8c1134d46ea508b6c30d6ce721b4f624011c
zc5c0cf160c343943ec273766f22eba51fdedee727b0aae966675e63a12b2bed4a742498a58e844
zf70920745488f3bd8711a88e5f9071fd8bf7e7ae37a06db5af242ec725a4a1d0da8f0732f9e552
zed49e407c578ac30fbcca4da687609cc392db2bb9c3c1d2ed119d45f5e5828bf4f7b6c45e4da5a
z0e886d9ba933bd063f210caeb5aad3b734c386b82a63ea7f3915c182dab6eacdeef6780b76c9aa
z63f20a5e4e3c02999923e5c289ba27dfec7c265b9ebc9f9f3601ee495c18daa271f075226bb339
z6d2f788bb0c0125ea57a5ff2ded5712e123866d21f6c82c197155509671739076e928e33f7df10
z4b9d8a2bd2aa12c4391cb090702d5a3a3d05eeacb11a6169ad1014e87ddbf2f983b7261f5810eb
z4cda9f032597cd4bb6c4b36b905a0019fb8337826be0eb8c19dab47a448c2a8ad11ea6a507df8f
z743fb93333084e2bf7d1bcfcf6f824ba5fe718e0f1264569ed8b192b20dd5711783683bab59658
zb43bdeb6ba896c7ef575105de9b286cd648e1004055a268b5e313de4f8e9db8af27c38b431748e
z24779c6ee1128bd7f6a89735cbaf3f1360c4ce0f6eeffea1128b63a37688a52638d0d26360f00f
z67c4ef911fb1d98ad2f094ad4397493f08b53e6bf1fcb77b0bc14a6cd3d3ecb3fe5b87c3185725
z966f0cc4580ea70b3d086ab607050b708a59718ea2ebf4670a518dbcbaa148a3964aaa117e534b
zdfed9e7b0723ec387461e8b31279ee4acd360c42003037a1fe69383fb9d92015fcaa8681c55733
z8fe91b6d9f7de669c72c60a02a4058cba8aff34df54763731caf22d3c32eee8c1a0fad8e11eddd
zcb53b24d9faa1207b7f4b79c3f587bac6b35c15880bde77e873f7d9d29c9a2a25cae3d02c9a187
zec1bc46f4c411339084ad4d13b7c25ee9cc4a8a7922edbadd7df362b11e111c496b6a7a3a619c7
zcc68e45f9747a5120ee41a2764b78f2da8f8e2b484c752e9479b5237a06b473e2d489849fc2a82
z036ef0edb989aceb44c60ba4e0b38f108bfaf8b0321096109a90a0fb8671fd50d06cd3bd66ba5a
zd003bd816deb1511f24ddc42081fe8c6239ce921000260b7e01a632650f6d7f4cf68ea560f3962
z3779b20dac0e5891791453417cdc5b253ea70353dd0b0fb56392bd2706915952d13ea49111fc77
z40e64b3b66d18180afa1c983254fc382621bd16cc5fa7a6fdf1b2e0432e95ceb2ff767c915603a
za3cc2192fef95c224ba173e3593bd5e338876c08bfb4673500e945c35b0d6920a8543b6ec6b7e0
z855b1060742dc6cbe1975cf579630d1d59f05a8f4c55df47219c68a3bb37c71ae3bd7fb17bb90c
z256ecf0cc02c9404f903c674da4ebe373ce3275ef2785c48b2f23eee61166f1fdba426b9324194
zaad9e0612b0e3fa7c7be4f3ff00c4eb389a4566eb630d30598202596ff21aecc447f89d709f02c
z247d8ced9ee47220f86259cb94fa04c29a5d4743f5a0c24afec7f952a7085e8b16d88bc835e211
z13519ddc74b5cf34a30882fb9e566d8b6e20da7b2f54a6c77af33e9b5e6e6f2231cae7c16d6dc0
z6611858a1d1adac6402a413c723c3e266864d3917a21e569fca1a97aa4877ce20f24124d2f2f48
z2b07df3e137c8731eea699ed9467a821b5b08ea05cb0b7fa4f3b8ef484eceecefcabc37c763b06
ze33339e37f0a5d5a342ae6a8d90e521e81d43528bcd1111f872c582ac1647f89b659bfe4509b59
z6984a95d26a8c8463a484e6dbe5643876aa742a6fdebfebebe3a34692b90e24b87f95ff269dea9
z6204cd0c549b43e805b6436095834beb954e7517bd0bc9aded8a4b2dff432a52866cadabaad61d
ze893774b8bb62391cec573321f331aa817fe9846949a23380b1306597d9b479d0cb7cfd948085b
z84e2078b399863bb0806692922e143c94a9b5d36c51498f605f1dcec4296124a8494ca87fbbd7a
z32576c298e4f1d9365abb36c3d74c7e2709e8f23546544f4a784bc0a3e075e2e351e7f841a163b
zdc15ecc1c3459c7666096ac64cd322359de448d3c20a5ba1b7df9176ddb96057c74358ea22fde5
z2980c9a003a2da4eca411ea75b48501d5b1b6523c30a09775cf9c8e40b24db81db7ba9c0837145
zdcb2d11326d141011dd69c2f31bf5d9ef767f278c8f55f180f90c025eb1249aab3cbfa2fd77a1a
zf554dfaad12228d5eaef4e7b124420c7fb60a1e6217f17131ae14d32cac6131505db89aafa5ba4
zf66af27fe3753822320222be866bb1554a682f7daf9a0ec9307c9887cb09d5406d10446d1e2b7a
z6e21abdb24dc90093defc27e8e5169a55fde253ce45e8578193466154036401b127c02f6a9a0a1
zd2e0248c3b98924b23f8c0a1643ce0040bed39fe4705f07a61af3eb3be01200bd87d45d62862ef
ze8f35d77a3d6c77eade9afdb0fc7288a8b31b71c6141f26c2daec114bcdd208ca02bbec9616a44
zbc5a90edd350d51bcec128ef3c5cbb795b964e3805e08d89dc462d68b851c3efa5d13f626c345f
z90fdab1c5c72598737a3f4f781a77211d85ac7af299e455c9e5e8ae06314c3e2d0a1b34199ecc3
z1c2b43188765747ef1d8843bff779bb96c098611f8c0939eec5627059bf92abadbc2f8d1200780
zfa4512aa529fd6bb57cebcadfa4b37573441c63700789cb7b9e41904910f0e949f06ba09b1fb3b
zbeca308930a83ce7dba599aaf6f39854e62879d6052a7d990a2d7553770654d5d86a633d7baa54
z8a3c614282e8a07d6a997cb9007c7d84f0f71742ef73dd4c0c8f5f911fb8c0dd84ceed2d3d4cf1
z9cea139a59b63a5fe562edeae93839ab4b32e7247a9cec658b5a3a1710c470f6265178e0ae86a9
za9f031ac2f17521b1eb935253be405d3fb7ad06c0562bdfd13d7d256d9256e2034937b49a83312
z7cbefa1fac849c6ce8d888b0894788f507d99470fc0cd404db9da581faf1d6fc3fd0bdbad7827b
z6b8c4c75410f7268c07690407412d8e69f2bc7d889c3c14e6262cd405f84da1af39acf0d959357
zede55acd9b7f52f1b4cf36e04c65244d28889fea04004024f8aeab1bff84ba0bdce616651f6899
zec9a333ced79f8f0873368cc8dea617f0dae224dcf02f22fde9049be8020905915645b6ff0a4c5
zf5572f954835fac49637b97815bcbb408a994dc6b33b39e064279abd8c8bd10dbd2023083ed213
z814363793c884c235cf102e0fff5382d95a9d7b8d7c46ed5085790545b5c976ee8a818d1b3b300
z0a3d417e6664ec84f0d72173e029ef183995b9100d9c9d3d27c37e9a24a815780f448a6548d033
z744d39f41b4cfd51085df53bb483d6f77db679af4d8e553add8143f0fd62138495724a21bc45ce
z4df827f777f5e853486246d406615c716e6e408bb5843c78426db567269f3612460fc480b5e5f7
z4315a56fb5bc1888ba364a33b933b51926c2f42c6b801f723189fba02b8afae3bea9ac7770af8e
z87b9c61533b86d9dcfc2648ac2af8f438dbb49b0c50815f957c776e5a8abbf5b20e4f1fd3912ae
z9e940c20d7ec7304481f148c5c57bb768396cf3c7b853032074ce43df8daf08f8964466b137648
z050cac71670f8eb2328f687c11474971b0037e74eb52337cfb647aa99ec49548c361dc2c48a93a
zb33030e8674cf29731bcd3910d84dc90ad4355ce2cd558c5bd05cbd96a217fb8ce50444efaf687
zabbbbf1ef48b61a936245a4543fc1ba29dd0b70c88694c07f4ce62640e7104337e47e654f5cfc9
z1dd02b4400e85a15e9f66cf43bd168f7258fe57b957b0caeba7810bb18412c0e894810a4fd5aa8
z79b9d799c3e31ebfb22ba8d6dcf6d0fa339266d9f0e7ff674ac1da2dff1cc6626dfea7dc59a391
zef4c049acbe5f477646ba9b9c6a40a42247ca44b6e4cdc527d5651bd3367450704dd0edef6ca24
z9932376b819ec0e6e1d1a2c343df742d4aa975b8193268cd90a5256687bafca24b3c373692bde8
z492b863bb50b52322cb6474d08fdda9497a72cad2a4425ff4732bd28ee85d18d6281d85b4a19a5
z5a5f36e36e4be96e5e1bb3ae08755242cf26269e614767214b82e01c3485292f4f90cc18b07445
z0a4539cc90bf690699aee078fef830348b8b62b449968e7e5ba4e39a02520b23c0c8d1125b47d9
zbfe56ae676160e69b2cd57bf947e1b320356330c33eebdac66390127e6b9d00dc09788bcd72370
z88fd1b1482719b9c5ebf92e0d0795e91377e379d3c2ee0fa23e318428d1878dac331f60ff85f45
z386d742ea56792c93634904f12dc250cf6831a25a10d852681f741422ea45650693c23efdcec4c
z477e569a309c4e825bc9dcb50f04caf6f10b1a7b1965401f7ab1d84cc7f3df184831cd931753f1
zd583966ff2b5079b3c3709b7eb9510e2f6d9f04e6a420d6f2d8d6cdb668adda56b381ee293abb1
z8a924310e233f9ba44bedacd2990ebc20936868acce23dc35abcdfafee8566c38eebca6e674bad
z2ede7e629b5604227d71edba2fcebade26a9a4e4adf12931257cf34dd68536c783443562d0ec34
zef7747b06f257976904c8c6227a054b0a15ddb4ee80ebca9a2318f2278d27a545d5bf6583a0033
zbc76233b09a54f120f02443fd9a15095987d039ae10c860de32e4088cfddc045874e1309e2f320
z13c74f307f4c934b083231a79267ea04afd95f9c1ade32f59aa729d0c988f89674dc0395a4fd4b
zbec9a6ab84ec5100162f65dfff54fb57f3c471a6889f82f3a374758fbffdef809ca1c119f657e0
z32322e706ffd8c226480e9b281aba380c5b723729617288b24798c44a8f7d2e1f73eaf1f247bee
zfe3254ea3d74bbbde86798fab2dfe82476cb48ffa452b2e9669979db7ad388d71dedca78846718
zf87e66b1bbf2d18ad0e1d1bee8a187aba36b0c30b3e5f33b7f50b5564604e094225ae26c94a6de
zab61837dc3d35898f45efb26c42a40b7ac55019563f5816cbc1fcf94adf4e63d71ee33371319cc
za343ec4c3b23ec82721d10477975fbfe3adcd6dd9b517dbbf7e3fc0bd643ba82d2fafeb2462c24
zcd635fc7326f312e726e81d142af9fa2ebf3993727ebc810970e9f1cd8a170c53d93ac39d25bf0
zc17e6093d8a9d52d6d3dedc82e3eebe619810c1d5be8c73a76916fb9ff76ff01cb458b9db196b0
z7f46f10706e7ed7e1431d873e22bbd7fffd08e9784c409b4a0dcda95d12e818c7f492aaf10b5b0
zf0d8df5de9e34d11d38110e483960b49bb225d6547a54b3d3c8a26d26fe57b4ee8a470f44f3a31
z62b096709a3b0191d0ff5b8a7ab962e60a5bec206db44968db7f0ac7cab758174df89b44a50ff4
z8d58d2c440f3ace2cfd223f18a30aca5333bf464dc268adb0a00e9ff94cc063a656229bb8037ed
zb554342d272854e3e17b5653525c0fb75593a0e9cfd9a22ff9fadb2b29981a95c095d2394ca483
z6a6ddd3e35ff32cda2bded6cbba94b031ea99d93f372138937f4c3ce80f0ed1e35cf1d848d3839
z4c2a44d364ad6b5eb9533f2292ded95f06262b6914bf7e2b0dbae10de4d7e696bed5acff6d1047
z651cf9ebda098375d6791a347efde90a20a5896771ed2b43e8ca704a52ed06f1a0686ac3d52af0
zc13ef398fceb16942daa34de1db903ee4c2f8b763d52571e30283a5dde820c2742633ccaaed42b
z15a61328d4a77201e01dfb3fca452817fbf743a88f45a77ca8993c36e5ec61ec05987a07636d87
z813662a15f7cfde045ca982c1341805d5e1466098786723d9850cd997e2ad403f4e02bffd1f68b
z2d8d3d52b9f864d42fb94c67f852658a3cd6b51d8ad421888ce6ae13744a495ce4c327b4856611
z0b2d4274ccb48260b12c2fefd1b670e8089b7ea6a39c1a63a3c40a943c8d45c95658d425a8f28a
z7b93357184f3a57466a14e433bbbf60e1a0979ebd08ec44fbcd5674ab634086d1f719796853d0a
zf85a55890316d6ff8ac06fb3993212a5e57f6b95e59ca5cca85980fdb573c803e638155171652a
zf894a91f3b400a103a71f68f5428843bb044b379628c5e9b6182c0ab9facddae62fbfcd311af41
z36395a87e6dca3bb9bcc50c73ffef371e5d69c7f1ad4dd46af0bbf0c43c2b28ac2894efe5edf1c
z151de3aa0e2c8e28cc05973c21aee8641de9616378822152bce89386a863418ee6ab16d1dfcdf9
zd726899e88b3efdd62526fcb18d3d5271021251d865055df5ee7c0536194a13af18e0b4071bce3
zcaf9ddc112678c53681bccbde359db9268a039285e99f63dd93f40a0cd7367805a0643bac4c17a
zd7c52fbf5028b71e8a7caf0fd1ccb112f026e11b4604d6cd1efd0043a400d655574e1a80567b11
z8bb89b7bf891835c33654cf9f8624fbd986d79f25de67db30f4cb918be9f605846f1095effd370
z9f1f9568fe19e1e7318012ecb4e21b6f580621f55a6ea28ff9db2573f0a0681d65f59bf0989fa5
z563bb0b26ae42f8fb39643b43ff2e92ef19da57cd5317c06940068c9779d8a3c27a3751cb2911d
z03d960fe523895a6b9825538941b606e3d6aabea69b1b777ddb7579717029625c2c1a88ee00997
zbeea13fed8d14aa062eadf9ce23fe3cc20edfbb1f09e99482b4fd7285c80884ebda8e2b3290a67
zd3978587b793f904e56d02db1cc196f01ce689a2103c6bd6532360f3fc536f73545e5a1f4e0577
z60e83d75243224705b27bb7d42b01de6f73d40c5ed706ef3fc87250ebc68fca1e4895c2de410dd
z707c85d45a099b5807a6c4b1e330a1267420d661b36de74581621f080b36da2ee5b4b8b53b0a9c
z405d8f09faa80ca78c6fa97f21619df5de6113027ed96be9d35dda6379e0120a4bf091857b6b97
za71cce11587ccd42698c52fb7c8af07922c010a4983aca732717358b4d5b6f0d3ca3570961e2ff
zd7164309514469f4c0e52c0df1af710d83993861ff77b259c23aa9933d45476b811f29f4ee1729
zd8fdcd1e18757ec6edf68b896a57e59fe8b5638caf8ed20c987db2a7ed0e8957a10df971ca4003
z55126cde5c8553b3765c04789e7f075935a014896a7b73d0268c292e8ea6dce03eb67c00971c32
zaea91f8462033203404aaea28f8a87b8b1939f82cdb565be32d527df7e05237bfd8fc316f72480
za8459581d862e0336a235308e030e180a3fc3f7181aeee27b034bcdd5548a137bce4ffd2cf0871
z3c57697bb5c53260e6f037d4be673e7e7cc718f7784cb9026e43f736cba36fbda595c78cf3bb6d
z2440880b9e13e087258dcef754a873c4e52514e977f9632e0afbf25ff02e5ada196b986679c24e
z64ec9254b714a9eb5e0a2668f17e2c4a9d22d6d9e231ee65e5b64005d3e1d68f99a0e0d78bd2de
z3104a9b9d1205bb7e4cf531c8ba0444a7375f9c20fbdb6b86f64b1472cb9121106a035fe16f72f
z79b2cc7e5521b3af1402d6ca55802116d7ef8327281d4afc211f0495115c8243ec9b7c2c4c1197
z022a17988ecf4f8c36f834340d3c6ddc828e990be94f080f6d9f0c535a9adc229522f73ac501b5
z4e88b6a92ae417acdc659d2df857a8d558409016b24872d6e5700c430f746e54288d344d47f0f0
z981ba405f9948369b07612f5307b6ff4a14193732a978f7dbf09648c2452e25644535904ecb093
zcd009dffbe1764aa70a8c7e93b4a4f60f223c2070cecef82aecd7a83da7d0c4b7620c5a499158e
z2554d08af7ef8b8426bf7fd9f2e4e7d111502dbdd48828d5117c48320a8172633f72b08bea759e
z76495838fab2c73db862a50197a383b7cae65ecd8c72e218cde7cf9be4da43c2370994e723ff7a
z08d4132ec1e4d4bb699968d0ac623970952735dce813036273a04ce4a037cf7b4e265506c8dbfb
za607cca98e67a19f50b061d2c4ff6a7dbf69cf5530682a7da19e637a633e370371d1afe354ac27
zc74aa95fa1354449c7fe35d0073b7efdd07dfcfc915de1c05b81d902625da766935ee9aa9c6e30
ze0f8b443cc7c0d9eee97692b46c7195996e728b37e722d3f1cf285c49483fe8acaa33815e01fe0
zebd61c90e70f35270026c3de364cbb3902d8c96296587112fed53c4fa6c128463e1774023fe74e
z2fa968b7d936e72909a31f5fdce38bc8440810aa477965b65f100a59ab324c6cbc528e6cfb0b72
zbe2d7cba46aae7e0a3efb692b9e308c1b08eedb28ab5b8484f01c71b506d2a40053bdd41815c54
z35af0b66d107ed1e724aee4da6c28fca0d48a9a4cc13b3a9ae56f16cc701eabb96d04061143f04
zfddd3cc9624e089997a03185348bfb0f0dd46032a2d11741f63e2825a4ce8ccbecc591191d6073
zfcb6923fededccc5ebff9089bc72b6805c7bc83091526dd0467d1fb332e0e145ee47de52080788
z3dd0538b33e72b3e115c18900d3f7dba8eedbec188133cf011fea15183abb0318b20eeffc1cdec
z2f31ecade2eeeb617168d4d23fa5ddacbdc0424044ebef5a18ed8b533e7879bf19a7bd67c45e02
z4b9a1a46576997a7ee02c7830a2c1997fb11375f3c114cc631762678e2a0c65c5fddbe2ad5b7d3
zc34cec61750d869d2c56b2688c849c9ff947254af37442efa2b87438aed452bec526e0b89de625
z6f4cbd498e23ed3256143d3e09642fbe8f9a53b79e9e3e765223c8e456155a08ca086103eb47e3
z0d4a197e8b789131eec71d4f56122a134cf7f82130dbf3acc6455e0bbbf918444bea5473745d62
z024a236f953a2da8cf3c6b2ce786da583e7352f80f63bc71d814342e5f6b8021c8eac6c51e84e1
z6351c40c22a1ef0c14a98c4c27c5cf2e316a3d3ece2a6f842bba7e939c4d66e165b42cdcffb2a7
zc926cc0db77b47d6060cd02e0373305eff8db2097edfccadca2ba561e7379f91bfebb3c1d5052d
z10c284bf2b02344d3cc6bfb4689331d1d4080053fe4018878428a3e0a3fc847a8b9c5b57b884d2
zd98a6ceb9e1c9fb6c95e05a4330d110d3103af21e7cae5adc7eabce4637ab525386d9d0efd6d38
z4038f2a4dd3bee4d98ab8d9c087390285e40bd847e338c63b08f6476202c96dca0197ddf5bd4ef
z85c5051dc6dce37a65619f98418f18faf1bc1d0c91501435d44689c29af13c32478e5b6d49b1b3
z40cd4510df44b6e03c7992d0445863b90fd631100313e5075aaecdd220a28178b6434efee8fb7c
z374815be75acecd7aca50d4ba43b84b2ff26a040bdeb8d1c1c570f7722cb2210d01c1f6241788b
z4230a30c42f76b496e174790d20ce03d9ea0c69c1ac9428285a5608c429e143f33587aa1eff3d6
z5d3b1e573546e6c2f086796d2604b74f36685123a7d0c13e153b5bf3b3a6634c85e51cffa907b7
z714569b5d92c9ac58cb42fca0eb61703f88d88b23d6b6a9983bbdd34ab9dbabc21b4d067455ed6
zfcf87374d1496cceb53015fd5f7eb856fec121dd14287d3d990d91061f2a87dd7ea8db9daf9703
ze742a2c644dc3edde88120eb5fe23a2e51936c9a8aa314060b8a44eb851c236236880f6bc1a359
zdbcc05522a5308ac6ee5d3e03e95afea6dd92b71e7df209967ad9d9cb5da41cbf729d57827fe49
zc7f5a90e78e8b95f418183677cdc46fadad744319bf05f1ab6fb0510f2b6a607c093a9c7a18b74
z559a6cdfdf9cda50350565445ad5390d9127e2ac0d0c4655421c93045b8acdf0ddba7a21c69753
zd3f5e9fc9245fbeb47d8b380b8963cc58a1b98588aea93cfcf0e8ebaa87f4b3278ff9ecea40f2f
ze5fad591b9ca9c3ec1d99c58f9885b6d423567d8c6c3e2481d9a573669ab6be9f9fa841b495776
zeb0470e71a9523a87c63f04d719fedb972ed25c7d5fc1e1d51bda7ea64fd1702ed6bf7ecd1c4d0
zf89ba9db9e61eaf60ee6be3d1b155a220ff5dee18b6a7ef644fb22651620a35a6490d2c0dd1c04
za2efeec300bbf9786e098f170a50e347a07fc143619c7d2b6040781cad7337a7f783d302bb4b8b
z25dcd16475116c5d69c9b39a663b3cf9841bc07d25e235693709a02c57fc788e2311ef38a22e0e
za8fb857aa0fe4c57dbbced592343a04fcf9360918dd83434d3ec907d410dc411ca03fb73089f02
z7e807cb7a5e7554478f7ac0d4fa194f5b37b7a1d0f134421987fa9e0fe2f9e725ea1eee388dff9
z1bb7604bbf3a395b4286539871a9979a7cfc888d30c2293c5a050842801b53d7202155dc31a7a5
z9c10beb197e81372ec5a36e89905614748a3d71a8861cd713ee3a81cf1bd8deeca2285fb8bd2f1
zc78f6d442d7484d1917f10e3831100269af982c528d69a47542d964ba777a832ff44dd09f8ed9b
z2a48a59411704e1a061e7e3265c130999ecde62a4f2febf211d763287bebc60d267f4588c7f0f9
z775443cdd7ef13851500de1ecd74a4ada347c1513ea414794dba5f5e263e3bd2c85f4485b31bd4
z78c2cb9e7ceb302bf6c5211f1d4acb89033a65d612dd3f52e8f4e4cbfdb9789a408d291ada7672
z82142139cff0c28fa7f9b7f6217d1660a638211b6591fa7542eeecd4bbdb26620dcd4af0f0236a
za9670926e9059f53cf1ba287de225e08ea2464abf58b12a1137ed660fa192e2d984f60276e29e3
za0babc120427957549c9146cde181415ea3d4256f54375f05911630032bb62f6d5ecdb5fcd7819
z6cadf1c0af875fbfd4c5709ca9a3e982b997af0cada7b0cbb5769c7cd669714d4e1a8949a3aa84
zc6d3e11e89a353dd692a06c7c5d7f5328c8ba8ec6f318a4620d63011c1839f1b4850f53a94394d
z765b4c316b6c28cb0b01003a3a66ce55d44f01ad2b47a99b0bce1500fb98ee7ebe59aeb5802e1e
z889548bfcb61bbffbef31cccc9d3864ba6c00adab59143ac9de2ea0e6994b94166841e02b28687
z7647eb4683effcc70d5867a415c100f2d11e6cba51b76c5cc056f89201405cc50949aed21677b5
z63c3c1831dd0efb1156525172444c5417288a8752941d703f2736a08ff8589a07b9df2782d61d4
zff2b821cd89c0e0fbdb82c3fbf15de6b87f415cd026fa2d6874b1264f5e4a3ca31ffaf69e434cf
z3825a7788f4bfba888fb16a508b8142647063642f20def5cbe99f825abe33f6f1f792f135b6eaa
zc4d6fed8264e75e54450b119408d55a3b78c5d00e9520c2fad9d345d480fd7a96405980286eca7
ze470f49ab41631de365edb3d67659dd5dabfc865b7bb82f1e2ed619f30f8abbd8d883720f4f585
z9057c1255ad725a9084d5b48dbebbd2f2998c04c65f37fd9c4e4810ee392fb1eae443e63d42c81
z80eab197af72d6bf15a49ab2a325aa0a7a975fc857855c4c668b36abc138913ab85109552d61cd
z9a14adcec459866af97adcfc17d7c74a872969c6cdd691969e97a3730bbf6362e749c90bca03a4
z30ca480efc3724de374dd975a14c2fbc74d11a04186a578ffc20a8bced031ac3a88826a3c5dc69
z508b408fac0c0fa661dbb5f675c5849385f672e9357241311656ac935e8de81da1d9ab7ce39ae6
ze5ccd555bef01c20965a2f45176ddb26cc033b2c2f278f82114663878f891f47c593cde85521ad
z956952277eb8695652d1c358a484acd22949683f598889b7e0b998a36b4ebee67e3d5e5df7138c
za631a6f4dc055a63fc091c6f80d4ab655d5089f31886ec30e866c5c088edef538c2ae0b1849c33
zd62dca73b9ba54d57f6f6508117f28feb128ba1827f2700990abfb1a3950275aa9036878a54732
z2935cac54c2895a10187bab956bd4148c5f203662d798e5ee506e32113542df2d7231c2dcdbbf7
zce07a47bb093c8d2018da5c52b91c806d93bdc4ee962cc5a3d53113d354cf17fd55292353b3345
z49cbe08ae49dff5b8ca26af805a4ff53b3347be0603329bffa85e527c74a4a4771ebfb1fd92dc2
z3382344c1209a68057380c42ae1409a9afbe85481d413a448e4f4bd934d6dd85c09a2c923ab407
zbeab5a419900ebd25063bdf5b67bcc56f7bebc1ba6748e64e3407bbff6d727fe5c65e42c17052c
zc007854abd2854b0a04593d0c824a0d70adceb36a5d68a8867edf7f89567fb739ac9b6c9adb230
za656cd03b3910ba17857cd8d891ea941b7d274550486f6c955e5b7467a90300df4e6ad15944e62
z7d70535b3ac29940b314a47887624bd8abf59528ecf506a417ae65a99f0c07b37b6b0f33c818c9
z168870c6f08056a24b728ed7361022ab550c8ffda97498e99d459486c52bf9baf7cc93f445357f
z5c059dd1993712f598f220e24cb2a7026c205ec8dacd61edf23c315ba96cc2635ac798357d1e2f
zc7540b0c501c69f08e855dd5900329ee025b57e2265452683113c821a9eb9705e55d11a8c1f314
z7ba161f05c11329dfb3921b3ec8c6e0a98358bfca8672dbbbe95de9ab573c443bfa795a3497ba9
z6be1ad9efa5a55a00443472a5693b7bb98fb05a54ff44e1c10171468f28da5365563c945de4f30
z5d7c4bad4478cfba1ece301907d2f16678c14b4e0d1c5775011e46751fa4bb9dc74e6c70291e5b
z8ef66521ae32aeed13baac2f28c532d7f2704f99fb2c854a19aba51a45b75f9f15d78a987f09cd
zdb03e70783afe8c906f3a113367aff812982cb50975ae7f686e2ee3a969a7fca68ebb1ec14b4fc
z9c51d9b3f69ff6bb14feb4b57f9a1f41acf9a06448497889a42689ec66ec6d95bd58e71a3d3c43
zff7b60410701d392ba0cc47e3173d5529636da7e296a7565a6fbca504a01b1b105369f49b57281
z1cb445e9b874a35f49ad553c3c28c32f705761edc8c2b36917fb90bd9116e0d8941cf7e6505e7d
za80942f435082935091682fb446e2781fe00df2ccd0e28e3594e0d01a7edcfea056ca189853192
zfb9fad514b4ddb0c8047a55b396ad8a96381ffadc0709556462ad2f0076435d93421e10c33bf4e
zbeb42da4da0e81b506c2d6433e63ca062ed4a59388343d9e326e463bf304ed8aa024d033a1f4dd
z35d3737d372ef293a636c8f89795623cbee1d350d58335e94c004ec6357760a69dc01912e2d68e
ze5592722f715db6b046b346ee75d035f7600fbe1fd28a40daeac77adeac8465e12f4e79004c671
zdba28a41c568aa25e582fd6c1fb73a5bbf7edbbb531baa5406bb4235b6031e15be10314ca17400
zce1d8a990d037c77c594f1e1c76db78de87d5940d94a8abfb9ece9fe01a3018809918aa7b76860
ze3767861d042c1971923e01b7ca9f349f0ecf3a514375baf5fd50de89a212ef6eac47627538bf0
ze4c40779c7a25ed04d79d0e6e27fd4045bca597a1c0287155927f5800394f6f0da663a4754b1f1
z978377a8c090c8d620f293466241a97c82f819ce9ea28bec2d1dfdb69cc96e922c78345fb34bb3
za5a74c1a84396b9025d12961c5f9ce070e3b9c53fac955bf33673c1920a172137c062a6f810042
z1aab247eb6b678b01eb1506aa0e88520ed5681283be5dd2c20452bc7a799a864af3c49423d1b99
z49ae0be42dff5f3f4d61da71115c169b7486ed5738d094971bd44f6a8b04667ea10bde2c79a6a4
z2143a5c7ee4704d0be962fd0d1833e8086b92b6e518e32f8a87a28e43faf935cd50a4b847ee337
z664087b6e52d15a5c3c205115792b1a7912798b0c0c5a52c8f0c4b1ec3fd2fe508d20f5f88c428
zab57ee1e352baf3a6b197cb9043d150c5161c53114ca59b5e2f2c5586fd2ec71f655616d91b76b
z29c2245b61c3657989b15fb77763318d73f60ed1066cbb724aae21ef1c3ada0a40159317d9481d
zce2ecdc5aa9cca8dc3ec940d594c2818fb809fa1c56b54fda20cc4dd47bafec6d53e7f28438632
z267a29cdadff6423ea0b29ebb714a31b8e467574d82ef9a8c7868a86fbbb0908fe54fb86575a1b
z9a274c273212d8f7e432cce5cf0be28cc04de06de6dfd61e58035758a408902a3311ce566152e2
z1b5779e7acf8a46e22ed57cfc78a707ead37aca74f1c0ade337b5142041fbfe6cb5965e0603a73
z269fb7f012d3c9caf8f981c0093dc3d9cb4fa4ae629d2a2423ce2047a80f6af97654b3665e7e18
zca76afb42aaecbdcffcef268dc6b5022013ccb6183946a92e3dc44d66975a5803554a3982b579f
zc38852f524a28a0a8f3e3d91d8a6d077363c6d07ba231c116f5a1f099795043b310ee79e4b3754
z720783550df9bca66aa57e086a240fb2dc99f4b229733751923e0eed2efe9783aceac91f818694
zc247d5dc75471f3f0112145dc5486514114d838777d7cc8b763faff0078909fe0f85bf9b476f0b
z74d9d24dd1d368437e1560c9cb7ad04cf4142b4426d37cd2696edb6e0e61ba94f609f2a94b704f
zd0bc272414df0e37b741a8b06254440db2e12dd0bea4424b642d34c101bc4c9cda12b238fd0492
z9c6b46b1af7ad55a1499ae50ed1b47274daa6ed776c7918123fa73d6152bae372df5a31c4ea77f
ze4fc41a4ce9c9a0e85e7e559539ea19bafd5facd555854c51e432c9bb2bd2f85d3be02b8b25df0
z6f6913cded193bc5f75779829f3c024828aa396eebbf521f3ae7077474bd5432aa348e191e0cbe
z7861cc0bb04ddaa95e04909d307667e433768986740d4c267ee75636dc5da13c1f8a71ff3b3b02
z4ed3cf1d9cc4238d72325f8f38a18a1b1af3a3d23df48a69fd37c14872ac5987e004664d3719e8
z099cd38820f9aed09dce33abb3c1840434a15c9aa24c66a6feb60b9dc1f21d665dc2b29fd7294b
z34807a64431a36221d9a63a9306c148bbf3d4a809ebfcda5da6cbf51a296b2fcd7a6d326bdb672
za1eea76edac80c4026df826ad1e056e716c2c022951e31c8bafcc8386e5f3de10d42eb131b0473
z8f4bca9c5273f83080401e16ca1ee879d21a5acaf97f11ba1aa72e0416966527c3929bc2f4abdb
zb2e0e8f1df4a6ef558c7826c2c923227c4ced375ce42d9289ab0f371d2a48974f3791749a2d422
z0c0e412b23640cabe68df353ca5d3c4bac11ea9a32a41bbaebc01963464c4b3ccda9fa8047f0e5
z97c10d18cc9fc02fb503a0e68e29540a3a23f10827fce269f2ab90140cf9ce0ffa61926b6846ee
zc05bd1e70c499ac1b936d39e3089920f6f63fe53414223481ada710c6960ea035fc51783f48674
z65e2b1e7b913f700dd0a5df0a39abfb2d0a7c755659f4678eb2017815c6e9d5a0cf097f65f2504
z2724d880a5aa24a406140e410446e7844517604931b53ca03b64cc54ed55653aeee8d3293f206b
z84ca63d4ef0ae182d9d24d653fd62daa302e3585829122d030c254933628aa3a70338f5c7998e2
z398707efb640e99ac6fe3669de8a3c30d882ff92253e8e4016458580fcbd8f835735f5b262e701
z242f003d3f1a526e3f36f1fa8ac5da7ac411de1f9651572cc628ca4889b86770a8b9d5051c3d92
z3dcf3ec6babd19a0ad39bbfc3f794b5d0275c56054d49afeb1dde112c63dd0d442ad9808361ed0
zbebd3a3d69ad5d3d997d65ee4c82daddfdbeb0b114f095192e6ad49957f7ff02ff859596e9f624
ze0d2fcfb1c081bb01e87dc5adfef350097811cca9b69c34dccc3e69e5b840e5faf7feea583f913
z7ce1421c2b0ceec40cf77bc4ac6fdf23027559170734291ee40814a61c0dac1c4530e87e92a5f7
zc01d8a98ded151f0bf9bf05348b5323fa0e369ce5b216bf537d6547c88486944d5843ba333cb28
z6348d796b5db2b679ea3f016db3fae7607a140f0c2e512c3308121ae93c528e98f6de9a2b578ea
z79fc506e0add10c3c982ecc2e1167e520cd7850a5f87aa8a55acea24449c54aadfa903f728b961
z03f41b5ea7fe6a9558cb542e43cb86ec9131f68749d35f1fe880fc2d7be0f08857c91a3741bb7c
z5d7ac99270d1ae592de88b36307703a585dad81522b8d710d04d52bfbad8aff1d6c73345b6eb18
z3a7df68b61fcd4aaa4b57d4ea6be5e303791a2344c706b38f9fe138605f02ce4c62926d05e3513
z1a4d72c31c85c21399aeb81f7251a25540f5e9c79aa187d3fc48b57710bb16d149d9767f32fedd
z3403004db2d775207d2817cd1b7f468250d0401479a57ed3e9dbe4e1f4c1a4af4e067ed7f6be44
zf8efd2daf764fd9711b0cdd8d82e8e4869a7ec9442ed0746fdf402b7827e24c1815ea8f6bd4825
z07e25ec76a6b80151426453460f759fdbcce9b6e782cf79491cddc52976a584b71a07a9ac0a67a
z9266a78def26c05f5697a2cbcfe7d587bc76197403fc116ea1aff0c09eb35f3c2f0b45f91c0e01
zfddd1fcd2fb1f42e6348eec9fe980fd3ac1b51f5aa43bf4c44fe75fcf71fc241dc5c0703820883
z4e87f053f3893a613ab5c62afffc675c23ee9726a2dc88ddf8c814d9d1307d872b03b77b07b4f3
zd7232bbd5ce98dc748d8e14abc8c571ff0cbecf018e9fac050e6f5d4ea8479bda17f6a9e1a55b0
z933358a4de1bb8a00fe9ab789eb3e7ab4024dd563161e501c50bb470ce4102ac6cd8d05f64e1fa
zceee72258f842b20d5778d0849fbe7adaf60357e0c05863844795c5e0cacc6296010e29b7ca4fc
zc9c112586ae9a4ca54a3433192d2ef8d70f7f741e23152877e8cae4d9e3cc146a6b57919d60ddc
za7493a7f82ab7527c84adcf580e3c5929203942a39a157886292679b7d3c5baadc1e56b6a8134a
z73577ff90c0964e67ac50d776a5708cd3c9d4f01a9f161d0dc37fab0db7dcda65a66cd82375bce
z7fcfebf4e370ecf04c9098b1f005bd9365980b1232b4b89c85a9f03c48305759ea4b2778ba3b5a
zf5068bb82fb64a2212751cd66a120f542d117c1bb2d336231c821913b62589b76eb99f770f7e73
z77905a2c7f248ec5b35c48440cf983403d833daa61eb8e6bb18810a9ce52ccc799eadcbe5844bd
z3c730bc8af238e8b85291f997ae021ad4ffc73fc96ac547d2edaa2a4691703a8c4e8d9d8aa3cb0
z395b6296db2f17c1942c0adba576b61eef0a57fc8a515e81691e610fdfe35410f2e0bf030dc27c
z02647434b5e5331fbab3835ab4df35153f78c126e082ea107358c08fdc7283258eaf2387e440f5
z49c6b49c238f669a76ae499b123af0a0302a47f01f4418c52fe8ce08a16bc8328a863e3185291b
zdc113995edd06fd096747a509667510edc63cf062fc8527ee36688ebd1b18c489bbbd55828f91c
zb665e10b55a75396660d8c00475318c23ed290502b0edd799d87a548723eff837d10940e6609aa
z3223a14301ecf3bef02008aa0be2eed9d04d27a7b28ca67d183b22cdbb59f64f5cfd7c9285406e
z3b68fc133b54b26fbbbd2dac2e585fa22ed690c76f9ba8bddc529ef6549ed5e2e0bf0a2b4f537d
za8f54fe03091d88f4687f502e0fa6be64dc2ab3f4c8c67c3ebb989975edc29ade25b8e8b3fa1f4
zcf6841567f93f862f72ff6ad9db99bd1222d9e52623b8db305cf82d74e58dacfb2c90be7a66a37
zb21c5431e6769be40a64f8921906228e00e7f5900d5a31ea5c344e5f13a59e392ec3d4cb771949
z0483915115f29174de8caf9f15fe5f6d9bc98c44b3043b467f6298edb5d4eb765e5cbde7114055
z54434398c1b940d93e94445b94fccdd5320bbb5dc9416301df5b354d7cadf6035e1dd518c3f791
z716caa996ee606a2c45442a1161d0e98c5d2334164867baeff13b330c7825c198494c7a0868709
z3aa59cb1661324387d1e5e79e80d5c92ab6e1bc220b95c35a5371880deea9741315c5deb1704e2
z4cb73b6c306e0692c9d82fe2f7f0262781d2c0781bc25fa7f8333fa3e7b54af7a8d9d4c42ef0c1
z33cf21fcdc4293a06f703239e971de2160547ba37e067cf90a7279a629879ea3bf3dc5be9a964c
z06ce2c505e8ab83e5e8e4f242af633422f0fe459e32495980cee2f9ef7fe4f083a032efd54ed22
z48b84afb01c4187469067a9045178abc127c2081fb4c413fb9a2730023e5cfbd7b5642bf1f79fa
z23865891e5a6d7b4d6f1ecaf4e6b2c691e105b94c7363cc4ae963a0ded303b4787e67522f7b197
z59beb9e3f188351b0ab428beab6331bbe7f282c4b4a3408a81b014a3ac9ae3b8dffa58a7adccc0
zab1a93b18f84e61525c370fd867e2f8ac839e948b5b17bc7f359a1062c2089b712a4bf49960b9b
z957748ba1267887781efe5050c0fcd9bc03bc63bb2b4d3030268c2ed6c4a57956281a6a45d49d1
z77ef9be1cdce03c31709c7f69f776ec580cce3c421826001c47f537c5c40ffcdd70ac60f746a26
z89df82a6a01196f1c9f2940142f6d3dfd17d9023df271dddecc0d55325eaaeff2d5717da703ba5
zc39c8acdc1ca25d262e8e874ccb52e51e8ac9f3478d5abd690607db71ee3d11d7e477d23ba8030
ze5ca31caca3496260d1c66c0a6adc6513443ff6efebfc2d2550d457ebc938d25db0e65d4ec9d9f
z843535080f3fce28fd104aca09550588aa0d62a3d7fec888c7cfebbb403ac3079db9153c7b7543
z0f76166e9bb265a767bf89609e4be6366e3d30795d4101278569ccac29af8c179c3981ed0de8cc
zf027cc6971feb94847141532fccc49f254937e9dbe9b421924aeda3120ab3c84523ce9ddbec64e
ze8552e2f4f510ee7203d67c86a8ae7fdfaedd36c8c1e4901d9f3e76cdd53d8f7e7e4e051a29323
z22eaaded681a6996775b4b4db0ca7680f171537eb0c7365c57ec9d3651e5717c6979f0312c8d4c
z0ed6ccc62b8168933e5c0719abd6d494191195a829dcec1e9e749a066631c0a074074394e2c049
z95c9e2a6f82dc485dd6cd7503918ee7d59fa6d1e05abed1f4b007a4a4ee0f2ce3424b3aedb2250
z0167af4fe8bab2e1a8ce2a78e6bf6ae3dc27f3c878d63575d5ac201fb24f0e562e2c6b3098984d
z458d9de7bf495b233d2fa09d39c48edd4039a3d37312787584c2e29ac60cb27184acce0ea753bc
z2660c3de823d0e26bb906daa2b1e46d1276d6aaeb1886f4afd22c98b449207141be095822af79c
z39f63527dee8b599965baceb664beec1fd7775f3cc2a2c755e3035366aeebdb9c85e8cc07c3878
z8e107f9548dcc8f8348a5a2efbb5a0f36d25aa1ed35853702572cf7006c2bfdc55be6c4e36f768
zfb6a9cb80ceba394ea3f360ca4b012b0af0019bfaba917aead5c742d221711fa4938ed9c5c3ee5
z40050e36ac1b98fd9ce9ea6812499277c3c7f3cd714f3177aa5ac634f16c4a8d2b9ddfa0b1c91d
z7b9b8d8848109419764be16b09e58ce489d7806b15eb09c33f3e706f4ac945042eb02a9263bcc5
z3a224bff9116e47f3cd1e4d4348c581f4d1acd93c391dd160ac693e1f4cc1d9d3335b65d5f0d2c
zb963f2cfc50d2490ff509c96fe57d3279bdb5eac3f4c7aa83b698c4d140e470a3e78cff775751c
z444c7843365a57981064f85d40220eda516b9ce0de49e900deaac882691bde80c71570075799df
z52f56e5195013e2ebf59da4b28e1e6444b2773e89a10b5e8bcc98626ff10888c237865f4b2bb37
z08beb869e5ba427c4f15580cd238840cda419f17b465d5bdc0b97f18ba5e7beadcf92b10529602
z9415df15fe28a4bfbedca50a3329c2134b2a21d0a1acbfd880c4d0066605d0cc105495cee28071
za2fe08dc75fa7093b71b6814bc4ef98632e50c3acca3e4ccaad4bda048b905888ec1354ffb2b14
zc0af62980410ae1f2bdb299b4b6ba8817f37fc9d9773e1adadafc98017c034b16405f1b4a9c912
zeaaf8b599ef26581872e153553678a60d91770cc42611fc9f610eed615fb7605c34e5d775b7379
z2e1935d45f5760cf45e1cd9c498da6bc54d6f92dc5f002fdb87a94f12ff61fdcc7b327fc4041b4
zb7e36c46140edb0e728ce72eaed7c8cfc50eaaf8bfca847d390259dc8d9df69c76d40a318b3e84
za2f41e59badeeeda337445c642e18784755de545cc0a8d87e30826585dc05af793621af08174d2
z3085fcc802b7637ccb300aec40b94a8b9a90bcaf7a08c7ce945982fa5f6c401901e58e48aa31d8
zce7c36de7f9a848bc770ee6977c1ef3fe75548be0c69945e776a8b7fb65855afb832c0f9939fe0
z27d3d130d3339a684717a1e5c8205404428567a3019af49c5109a2ea0d9d7469dba9a1796e2a95
z800b3dd16da90a105395b7cb7ca1375d83a66c9347718a71b3e9f1594c085774d51ff6097be3b5
zee1f253431fd7636dab39b97def1010605340193f2fe9555d6592c186cbd5a7f948969663feb38
z498683491e2b2ccd82674f61c74dcfe90ca7d9d1f77aeed6fc752347151f67d1900715ffec2063
z0e723df2f8ee27e79e666686ff992c99798a4e68536dbaae812f5ef8be36234a7232e99503369f
zafc644cc05b5f309281176679bc4e18a66a3acf125c749beaa9254d52e6a312e92e30be1425cf1
z439f7abff792d7ad0b6b154e163204af0a8793c8f561ed6fd3b9b6577ed3c857c271b1d6a104d5
z937d011ca96d9b339a2fbdcde2b8b081004d213bd2fa5fed2f3b57d130f8aa198deaa70a98c4a6
zb8664e52e0b5f2de83bdac31a942748ba045d0b18ba222c7a33abc0a644333de9abeffe07dd5b9
z269038880c748d5f421d7106c070e32213f5d174ae83ae69b1745309eb217b945af9dcda273b50
zac5788a8592d61b331f6b7d83e01a2ecd8b67f1e89298adf1ad1c104a496fbec47cba33cdb8a14
z358b80f58b7097178ac6c9129e01c218639e90873b281640c906154a22fcfd54b914628250e077
zf0b147d0041f97d82c0e078363e723770b9794d600b9c574d22af08e353bea6677ea16b30da3d2
zf7af552f3e6ce292e22b16963025463c6fda9e3ef6f103ec5d52d8d3e7545c546c3ac7ab5d85bf
z6e6f7f0b795ae06a9b8f6ee45f0fe2bb88c02a3891a67265bcf48f70dd2e25ba238773eda60678
z609065d424fd6a05fd2f7444748ba276466788348e22fa2e68f5a64187d274f9981c333cac9863
zca4439470effa7eae051d05e0302eb5baa7dbe038b419e734564bb0213549b914331921f696fa2
zd5500469f14b2f6aa814ae07910cf785f6a2dbdde162b26e2aee11e7fee5aba93062add9e384c0
ze3925a785c01473fff9710a8bc501083c505dc4fc012c259cf623d09a8fc3f172c27c2bb9cdab9
zbcd673d1bf451767195939fa3f38c2c7f46f744db7a198a64c71648485326f35b58395f5cf27c3
zf2226b62f1d59d921e87a6bb15a064c0b93eb85cefa20937e460a7e27c1ebac6b93514a6bd9d7f
z8abe045e31eef3738108625a1518315278b7786a302342b91481bc8a80dfb95c59a78603336c82
zfe123eced154b6456123308d706bfac9821763acb1582929d4e04c059d7ae2c1393b0e95928c42
z99bd17a7c6c6ac671f6707888304df70797fb2caf9f94b89497929df7f66bb6da4a1272f040f4a
z0f0720c48ba808d17315afd69c19538225dd8f6c0f0e297fab35243f800ed88ca28ab4b53cfd93
zea7fe29378b1dff59e68ac7797ff583dd3060a7851c0c2ff773890ab05563b7b7c00a6b399da5e
zcfd5e21aa4764a8dd2af3ffd411d0ae2a4f565b2c17feb64677171c8c09c54acaef6a3f675b830
z73f8078e4b14837404983ac21076151d8549ffb62e9eb0ed333e2efc892c063bce0cb1ce301d7a
z9211b92492f8cd7a718480e08e13b2f82f3dfcbddfcb59a1b5378a8956536bb7ab2b73954711ec
z164f6ea675b1540aa15fae05cba654a06e0a94f130cadc3364ce164178bf53e00fcc1918e06ecc
z2cdce5fdee0a3363e1981a91830a1d1669bdaf384bb718150aee409a703812b20330d03bd3b924
z449a56382354ef37e55a92b2dd9ae27ef2169cbb1286d187ae8ef5d9ab3e759d0a5a9d533bbbca
ze1a9c4270a55dd39cede18c294e6f7f4d012f7a076a3790a8a0012279588892ce5c995dfe60e2e
zfd5d3c933ffd8743152dd91c00e57b8a71bfcd832dc890ac61596028cb939af4ea4f6658b7a327
z5de6569794cfeaaf60c2240bc81ea23edb3d7d468424a469fdf3f3d1c612c3ca055788d6d4be29
z163892830bf1f0adb4720487e33c04d0418ce3b309d88ace5e4622687a1e202897aa22135ed558
z984e4b6f453dc9d85c69df07d5fe4f72d0571a3d10bba56e09b27c902588f67bb5c668c557f18d
ze746c3fda7422f864eaf6b7f1d9e19630e7bbd84c1c086a90ea06cad95e015b52525ac7b29ec28
z6d47a3c5fa5ae512611ad64bf3ce0744e2ec00cb570a1f89af99db1b7ae2059d442db763e45266
z76a41e85c7546e8a684c0dcb0cb59db4f139939fd5be2bf23482a2b47a626fe484cdd836f9c7b4
zbd2a8305682c346e72f989fc948b95c37a029601cb543265e88dad183a2dc497e60dcc7fa9ddf3
z728c56b16b0e36cd29cafed8a78fe2a7b6ed1d34e99c31e27a640507b7cc9b705e634de402d684
z4f2cd58562127ace9c1768b893af0dbaa1959364cf787cf79f5da96d91311e0ea85e98f1ca90ea
z71e0cbead1423d9f739b4d4928ccff3154263525dea8adcbe2ac94db2e00b13e4a464df5557a64
zab83ed3a495dd0849711095de55052ca380bca1b835b4f5853fe54f281206a5297238e0ed07f16
z1101481b88411460c06b192965cf89f22f49385bd0efbf0faef79706a4b9afd986bd099132da6c
ze3ed06c0c1d18dd75bb3eb86b163a673e371669f830cd17e5bd917e7323251d5d39ffd94a241b7
z7ba5e108997e7755a027754fc9cc7644248c416f8ee0dc901293784889faab3fafbc05b0df2530
zad4ebbd203d5f2bc13b2aae5ee432ab145c89afebb72a12707f327366e1b0a54f7173a7becb24d
z8e4f9c086542d8d3a85d160932e7a509fef9ddf7b5047c231c939d2c2355dc04aa88fd50f3d3ea
ze0f7754a0ae201b8f42844fd094d2f6b9bb15055468f27cef7d2fe45f8a8ac0caf16208a8bffd1
z21edd4c43e10b23b5753ac7fa209e0902047152cd0a154043d57ebbfef5a7c822145f2ff5bf10f
z6ee2a38df020555e5ec0bc8f1a4be466a09366f64fffce24bfb6a8886b6200bdeb40f91deb6777
zc157da1da38bd5b4e419c56821f8d32f96c7ddfd5b33a3d1ef9d97c3cc9c6bfd490653cbf3133d
z63fe4c4439b678fb7561dcbc1bc13c851aef4bc40b12b86145a56ee8169b5c714576bf0e03f4ab
zd03a2da2b62ec03ea8fcecf72134899eccab02f5d9a2a93817a5d90f86e94f680734cd49cbe221
z833f5bf1897ee3a3be92b8b2d5a45a196b5236f138e7aee8c4051f53d8c40d409bbe65311f9fa8
zb701cac1a7e77067d4c7f6eddc3c194057dba4eba28d01ee0a268178fad0a771b42156355e067e
zd4823ba5bff4e18bcab846fb76246da511059f4342eedb6d750170fc7567ac7b07d915f142a8b5
zf5bce6eda07c91e8df7b2386ea90040df4dcef92477dbcfdb0ec4ea09d1df1e8aac2682d01ffd2
zb9bc6c35cad83292535e48ad6eac5279db55fe20597b9cb845f79c9ec4b08a21a01c954ff8e8cd
z0803dee03b3fdd430989f3deb45761a8ac4c2ae7f255b2df30322a7a60cdcad8392108b1aef351
zb1ae571c7f4ba4b1f017ac42d8a45ec6c94b643ec1fa082ba5ba96d3d89fa8f3fb46838f4fd3eb
z4a2f47c773b3b27504a04e8b480605d0bc4ea03ec03eaa2c8df930cd0f3dc1f78aa118f5f65215
zed74f6b8145b0fa634fd4228eea7f8a5f7f1a346e1370040096f093b8101e55b7dbd660bba7730
z64f0ce42343dd600d56c81c85981dc772f798f9d13199e27ca98d3d8b484a8d0abbf62410e2797
zb424639b808f1af1c9546ee79e444299982585b90a1bff154092a49d24bfec0736850aac4645cf
z62b3ff2955d72f951c7abb6b9eecfec7aeed351f68889560bc275a3e0f95207a08e15397b00247
z41c3e2e5fc253a1ff622a38c13ce435bed316b5d379e9b13788ec1930cdb5c9310d4a624b2e613
zacf3a74a6355305424b97191a3685032b47fe1d59835d4a72a2192ef4c52c0a81e9c872be7f449
z29ce8ac0d7ebb9e9f3dfddb7ead5881a5a6ec22ea1eb43681870aa50de60b229c61846429e5497
z6dba8689680a711f8e535a00e200f0e9a07d2d5d8c92e7b96ee49aa243b90f4ae02731e8bb2739
zc9eb9e7a6495251e26975855a806748fdc2efdeccdb2e133f016d802a24bf8642777c5621e44fc
zc78277d1a5a460e0405fcdadf49ef7f236f7cc735a7635fca581f9436349550e24783acc428f90
zb144415a3e2ee2ceed7765cd58af3c9f930137861017866f048622fe2e71f4c178a897146771dc
zbcc1c006ee1752ed86248ebdce5d5ccca1f6ca6ea1775e7919ba02459c66e4df3467cbe4b3fd7e
zd9594aa439c96604962f5f30d2e56df178360f216ae4865807b592f1c6972ac0325a9bc563084b
z699f7bdde6c971fa278146737b72be28502ca72a29fbdddb5e259521b4c234668fa01bfb299f69
zf36133b3cf0b766388655edee6e8171da6383b61970759e3c98c48f86c77fe6c1d284a7950eb25
z5aec89b603bf09a92733f127fbf5d556a4253ca0891eb05757574a3b310ebe102a0385af6bac1c
zc6330f25dfa8c83950a93bc01ecf41c719107ec31d89c83c4e00c4968693db29754504a2a5cfb4
z30a2afa401c1d74dfa5da6dd903ab3d5a91f4c127847c6db4b1f3330c89a742e3c5846e2af0138
z73fcd7bfb42f5dac6a4564d7b5e198ac01e3018c4c1518f1e6b2bcdd1fd96f0d4eb06a4f5a0614
z8cae1025cf9f83a13a11a2c67cfcc64b39acee3ec37122a3369fd73f312347dca6ad5451ca7ceb
z3237c984ce2b7c82c37d047050c9b55e9c4a0a5191e459156392243132d01ab9e214a25595c2ff
z35aad5c678082a094a9bc24dec410c84cac62a0bc1edd10cda1877aafc709b0af6c675a590ada5
za6528a15955c02617828540d1491e17eee06d2d15188aae363d55f3f68e8f112ed34f8f22ca2f9
z057dcafb38d6805d9c85e8eeee7996cd956291282c03248e6497b7187a7793450889b95b4fa6c0
z5e2fe8dc2516c745946819d4b5a066b5ae5fc34fdacc6cd59afc3a7d1d2a30851efc9264230bb8
z5bc0c65cdf2d653951e20c888b9c92cf7b0874424741fc3659832e254068fa767e8ea11c9842ba
z5d225306392d56b11f1b20ccc55556fbf81fce844b3573c3d289352594382e69d57037239356b8
z4037931d41f7d3541e1adeee3174d6b63b9310a1a1822a3e40e83267ce84fafe73a9d9a5b64609
ze19864d5ac64b50c2074168c51bb75d26a30b354ccdf37b9e8fedb78895c2ea9679baec8d9589e
zc64015fab52df160500c3b1409b04d5182892c19c1d62ce6c00a0a0c3e5f757ab27455564c9b1f
zc3ac447c507077c9a64b8370cdfb46faf78b340f4b98d404470daf50d9a3313c12510758357650
zbcebeb38bd971b44af662a9ff5951b75b8a2d69ef9c355356cf05902f0e4e5c62a1611f936c03a
ze42407a8dd099f603e63bf2f5ab3354abbd5f2cb533594cd9b0cc8fca070c82e60085c4be9351a
zb0056264badd6bcab5c1ea295ad6a4cc4f06bc31d351dfc73f492cf85c17656cbd026ecb0ff3bf
zdd57ab28f7e7ae09c082a1dea2c6dbe4a13b58c58360b467c266bdf4952583ca09af6f5263648e
zd0f1e56934c6364b733b259421d2ab0351952a56c47840275148937af3cba31bccbce8e2e6bfed
z238c916a7928ea0116188054c3485101d6207fdb498587e72d26c9b9c9a74aec2dc21b55e97239
z33e9cb19c0c45be43cd220bc7735caa2709728d1956eb060296926d5b0752851a7c2863d60df35
z45c1bc96b4f355b3fedfbecedc92bf68777cbf5950290c0fc3f400f43f4807c2f9316e4e0febac
z1802d7706ebbf367eea9bb879f678b4c4f76f634155441540e4773ccc3bc31bbed9d0d7a73e1a9
z897c930737e6af141c394a61f366634b9d7218af934f458c841a807cebe9f84a2e2fdc1ac8e2e7
z80a9d2c772544346e704425e0d449f46962b594ae779141398f2aaea52e1e0d8d1ee9ab33ac0fe
zf7c483721dcac92bb0f4b2087ddf1f9b60284a0b342a7bf684d3b8ae4bf07e89afefbfe32b340e
ze49792a8f74831d2d8f846bb474b2d0a5c91b2ef2c3390aa6ba5fb67b3883edd27370cc56cafd4
z0868e0a677dcf4f15f5c69fd8d8e4b41cd172950049042f693cc12245b5fb8b682904901204bfd
z1649bb8cd35b5f4290bff85ef1ad2f8ec4eefba9ac8b6236d2da6ee5969087a7f6c61095db6297
zc828ee5b73e9f03a5fce3f2fbebbf19fcb31795efe3bb6929fd92b9ca962f4f45ac784ed624d90
z71ae0874773d1c27f2131e1be5416662a24a8fc35324800bb0698b77e160e7ab6f6b5dca3784c7
z1a58fd657c568384a9078a1464535e0984934b29c07663948a94d285e29c8bbc3169a694e91e2b
z86017752e9fcf5cf554bd4adb4ce9ca7363fda707b63ddcb864ab12a2676a68d9af012c33ef036
zbda67ed27c7f537c8106444c307f07c101a5c0bf86e38f957ab42044b37fb2294169775730de92
zcc0bf9ac1c35ae7e1686395af9c70af22d539f93949ee31a0a1671af42f4d51c6ff1e2d66e2202
z4b2769ae25a5f6f2a27f86bcb86bd808b849545bcc129746200a45f1501618ed10e6ceabbd7f73
ze1e1df012055dec02e5c2331f782f2d9ccef3fca680e7ccc13e76b67f63d26afb6028daf251dec
z232f5e82faed0499f801c2421543381ecf477d79a7f885df44b5ec50e989c3534f87b84c01bd16
zc5ef6a0949d7f02c92deb3c439ceb7bb9b5a6c305e7ed476161f273f9d7d1d833ccc9c1337cc59
z133f86805453ead09b2a01ec2d5ac3399cfdc63c572e58c90a10f459b86efefdcd182162647387
z1a1b9f5278d0df9ec88fdb96ec64aa97f166a239a51d243995f94bc0a1851783fd2cad2148238d
z428b9d25f86d951ccfce40c5569c11eeea57cb777a78972ccba5ddeadd7694e2de0a31666cc2e8
zf944d14194325030e7b66ee625eb0a849cd7fa0eeaeede4f258051952d9dea6c7764db46877ffe
z3f08a3e1ab3215b76dbb441ad5397013b01c5f6fc81a893f90d93f3526b0d47fe6609632eb1278
z4412043bbc2e5f5d3ff8d9afdf8868ed37fcfddad5dea8eb45a17816592fdfd2b6af8e49ecef67
z8645fdaa46b6047c9679f6d0a84ea7efd3d2c0ba5dbd5f4f4fba1e725c0d53ac9b5c90e7ade29b
z6df782e7d43bca7552591222d66ed846fa407febb134353c946513783f554a1544a18ed630d7b9
zae0981827492dae4b7e9d395ba3198564cda42b5c79c19825290698e176a03b95000c652c77a82
z59e4479185b407194fa06a57864973d7acad314f13af78c545f673b5571cfdf81aee4577b9bda1
z66d5fde127ba39e25dc7bd4015d164fff4b485a7a03e39d5cbd3c225b6e863460ce48ae670b8ea
z3efc4df65a2f0ca37c0aeafaaa221a01316a20a7c757d0cb9c11e3ec2c11a7f8fe5f0a350af78a
zfa485a8d1a03cf775f13d1b05ebaee8c76be6af6fa8c31abaa04f81f215240035e5efc7c395ec6
z0db759f509d30b9004e8bf31b17d627eb98dc724ddc51f3579b838b47bab0a4e3e8ce2fa8019e6
zdcd3d3c1c7ba50a5c9529348cd0c47a53edda9278f913ff66f3811b0bb7efea256522f050dd963
zf7a12c006416b835673ea43ccc054eeffd179feb89fcee71c6b45579db8074a0be76b29e584eb8
z78a6b8ce43b1ba5defc931764f73d962addd95e2f6472d987a1e20940411852e1d1214e9480055
z8a4065f28ea5d43cc8aa8886c438e642453b26da01b2d1301f56f162a0418f25cd66bfd94a13d9
z070501e6a49d769e27ecdc721c06895b75cfb84b98651bc0f256b624f071b5536ef38c9320932d
zd06159b061ac8f4f17fbbb7f456cb12d301abfda7d644bb3a743eba130c34d6442d822f3481437
z9b515389bf109eded7236102df4139df7342d40b705875cfc0bab0baf3df090569651d6cb71c9f
za6af3003c4d7f6b4485b583569880a4eb3386a5f80d652d8925b5035e54b187c4470a3cb2dd57f
ze7a876c55f0c3018c92259ccd4e6318046eb158030c3da3d05d7541f3f3895d14a848ac91fdf03
zffe2718706c9a2eb07b7ae4c179b19b92e14a610f64ac2f8cd42f164217eb2d2cb42eb21235869
z894d6919f97dce124639d7c427a3f06b1bde8b796d1b84d046a53a43754bec1a0b1c9012ee6b7e
z4935d2097675cf53fc470496c6d2404476afb447887c45a66c75972c5ecaa0b7052bc9e04c9aa7
z4765e44e0cf7f9623bee7899e143f1c6573b500947e4b0394b765ddb4487f6a417e9e15b3aa095
z5c4e03fd2de4aa1ae64a6e8430db668478c70923552db67bda17f2e66a318bdf4bc11461554569
zb16ce17992e93ae9f8615030bc968ef8ca1893b1d2fff3d6f903059277039dc85346f8d528b427
ze26bf07edace3efc0404b34257574ef491af734395f8ebea2411a8d3aab2f610c31fa783c23128
z63213d4692cb59839d49ce2d0dd1f8f2478fd07ce2bb8f6e4b7496fd05199577aab123acce360c
z6419a701fa930d519836af87dd00aa1928926036515429007895122a1d5b55a9416f6be41456c2
z9be40401dce4ea5f56a2daf1f51b3368cd3d626d745eda038a348a8e57dbbd29e81bd6fd91d082
zcc7323459cac4f0b7191a60cd52b8bb18b57fef2e9914d3a105758fe46e3b54452b07a4eaace58
zc66bd5bc4cfc887a920218cc763aec2cd30e5fdb524d2c6147a3bf4d7e9ebf443d98092f81e80c
z54d4c39edab14d522d9a6fb0823ea068acec84f32408cac8100a63ecfcd8d98030287b71516988
z2493da32c4d6a563ca2752fe2bda4528d02f7af6b5f1a4a4cdac6d1b0a5a987b17c7928d43ef0b
zc5eab634667672124bee466c225a35bed0da01edb554525850a23d749c64eaba86959c0e475252
zae6cfd40cb8c2012895aee9bf5a8bfb601fdb767392003d07f19e08c909996a9da9dbd7b20ba05
zc05a3af1c8d35890c8d9251ba7131447d5da5f32b97a9b1e8a143492598040c8819d516e7c35de
zcb1fd4322814799e6dd747957273e3e76fa98e3b52d358eb6a94ad683ee6af1ecff9a0f2e092af
zc8e2c6e862e2ac8431d6ce9dbc023603f6e6a314e6fae375765ceb2d9af93cde263a070d8444b4
z56e414670ceeea1cc080c27cd8babb31bfd5c26a80366e9f23240f81061636365bf44a5c63b831
za8021200a7075552abcd57be2e1499961209bb6cb1755ad423c76e4f87f816543a4598e4adbdff
z03b6e5c6f5260b5c552fea0c572b56d0b3c0405153a6ce65d1abeac541ca8ca43b75cbf7b7cea0
z8e6af65e915d60e39af3aa557e9999c672ad8e00b3794c102aee6878d25bb36c2b1f97c5346fdf
zd203ffceeec5a7b879ca2782094a062ac28982e39160b2e20e6942bfd69c3229ba9a2d5a3faece
z4517195d1fa152c9d1ecb6be0e94f405f23db789d13f29bb33f2d71b84091fd9f1ee27c920e34f
zcaacf4b5f75a9df9ad5da824600def91da534943baeeef3277aa3b1d75746363d15a32e3c6c249
z0f2928f27a412ab1c83d1712d1b0563404418d32c6d910f2bebdccaf8dcc3cc38bf2d3ec7edf1f
ze2751b09b832e47d2185d8b80b67d008640582875bd372074b73caa5bc4fb3e3f72ec90d86bf5a
z73952fe17f34d2c4e1bf38eabe9bdfb614e227425d3adef4bdefa1069d1684e7b6299d5ae17ece
z16fb147df1c07da277fac0a2b484269d8068e9335108ebc99143a42049eed08504ef83fab045f4
zc47d1ab5199b7af47451601608f0ce2f111d8955277d31919aa92e8b64caef4a25e94a13eddb19
z81764e9e05de8ebac4356e93209a9296464ec32a0adffeb1ff82bd8e43355886fe82cc2c5cb069
z47a7201b41e7673052fb6732e57032ba84a88dd1647c7415cdaa1b04078797fb99bfab041d886f
z600abb200572b723a5757a8e54a51f762cb20bc1e4563e6c11a201cfbe37a43d84ec166ce24fed
z7d685c8a94a66c6c0bab529ab04f3bfcb27092ac9a12426bdae6e3b04660b5465955556885a171
zb3442106f9c7281bbb5ee135641b957169947be2b2c660af814639715e158a5f64182041bd57e7
ze0cabd6b78eb3e9b5b5949444bb177c2eb285f32082f9d07b977839439f9296fe861b64a3ef3a3
z81de63c049ec45dbdc5aba4bfca85b87e026d5951f0f283a368d3f5c53580cd0ba04ef8a85e866
zf1d337c5c1b1ac3e499df264055e76d9f000cffe6705ca3d659927a9e962abbf1fabf584ac7b3e
z3670cef5650a5a14e6ef205251646fd6757167738c34db9cc8ae4c69d33694b736b9e097443262
zf85f3014243ecd26f99ff63f062a1219c8e4acc58fc6b8aa7f8fb0cfdbbcdbcf0791fb2771f427
z431f94020f3fd2e7a3a72bdb9177f772894751f5a0537186b5a10708ed68cb680a49235404ab48
z1868c768c77e4a40b8219e9ae2d580d17978a16f6178023bbb730210acf4f203bafc384376af05
z90901bafb1517fdac479820ea78f68fce9d8515d6dd1e331129f294ed3adef00c3bc2ef9abc5eb
z050a47fc87cc385dc735fe93a8995f365091fcbda1172311be122c42b519ed020ae40e3d9d800f
z9579ab913fabda1f616ee0d20a4b2d237324c33697b45ae45d0a1980fa8a9da900be47ae9b9529
z0f0726745ef339f98d4b06ef52915902aef7a8bb1b9bdae8998c8b2e6ee32b2355a46d39eea19b
z187bac0f32ff7b82a6bf8819349e2fdcc17331264c90d28c8fb8422beee615c19c4df4d7f0256b
z7e7653cc29a446a5fca4a35f8119b818c8b10d54ff987ff7527184371875cdb1e6f428a1bd5fb7
z001f8716cac2cf621d7bff4ac72222b942a08aff01567ecf1d1832b3fa5836cbd6f0d365745982
zeb891974dea14cab03fe9670f9a16b724196d4d94745f8f62529a82f184eac5f44672a9085c1e0
zbc2fe7c10df3b2fe41bf5e0313ab19c4896b56186002a0c235cbabbcec50660eee7e3e78ec3613
zd69efac2be697866618433accf82ec806b2d427780b01de28c7a1f6bb54a49d741c35dd0c457c5
z3fedcba790349fabfb327bbd85a27e15adf6af573ba82d4873c5e8c152d1a959d0e9e72c2564dd
zf672a6496849ed337053c8f10269e577382c8c72a419e41d9b47b8d80ade34083f8e2271a70f49
zc0ba8670564b42882bb6ead4587d802432edb1eca393a3bc52ad6b1e07790bde5a154bc0288be2
z3332ba0529b4567acbe343d143c284a7fde191945a9b94f425570660934498c9f188bc91e1f611
z59bffcaec4161857eed0cd08508760ad7cdb2f28951d5c0b83a7e0512c90cd42b70453762bd2d9
zdf9b18d52ab3b3ae4571ffcba6ab28f789e234dd40ff285534a6b9edb4ba38804bcb1364d64ba3
zd182799462d41e9817547d499f7471715e48a78caa1d552b6fc6d1f28ebed8ee183f7692145c12
zcb580200a2919d991386686911b3b643e71f3958b198abf689702615c1ba8b6dc1c40fdecab7f2
z055b96902c8a54e4d2dbb5e04455d8a2189bf79b1bb993cfed3fb3a2447f6db321cc8a3eb0f15d
zb5b805b49213f14e3b4be762b80f5d378842c85dec4f77cdb8d818ea6265d80651776175f2a2c3
zcb867b9491c80904b36dee3ffdbb066ca98aea60155e2237ed32a31eb065c3fe6a2d6e2783a71f
z1eb716d2d45a2f625522388e3f76799b7c0ce97fc9f7701d26a965c458fff7cd8d7523b4c9b6be
z86f7352c9ce27185654142e1f8f35e3129ca3790f3c571173e1123126b71ba42349e4387daa95a
z41014743f856967645c94037672edb27e843de959770a1bbab261dc76b62bdd64ffc77696382fa
z47e66d5c81bfb9e27c06c0e1261625ee00251ed489588e93503a4bdf16c45b78baa2ee989d4e30
z7fcfa334262e0095d87673e69885c540025779a0e9e68e3f533b4f78d1e82de13d3a00404116c8
z87a4a192ca6f96934bbe4d013d7fd5b6baf5f518474f54af0257c4cc0a7b643e4ef0a27b1cdacf
zd65946b7ce6e485d63183e6852e651234dbbce922b6ed4c1c723187e08633ce3e5576ddd5a2a30
zccc7ed97b6730e6a8defa2b568ef9ce0ad5d367e1b7889cfa843c066ffe2dfb3de03916147b894
z28e77b8872a75ef68237755f1e64c362dbdaf7d275b852de94ad71ab4ce3669b5ff479415ad6ba
z7502597e944f6e2cf9c60af15324cb3e7b9d85d0b1325bc2a6cb5857e76b2f627baa3ffe2de916
zfa96b49121c98c92e9543c7afa2bbbad35c8ebea9c0f7242b99d6136f4d8616310670b870c6a62
z02543afd2fc23f9ccdccbc60ba96005af53532bc40486af5044980dca53832ff5fb4d82cd42593
z5edca5468eb2f36f042a7849fef8a99614389c64ba741c7910a8ae1b2ac8313724f31e25933061
zf7611b609f32778772f426a1ff2837caf1f73132c275230be9a9dd3529c172efc962eee7dcc74a
z69d744fc58e98d7708b25a51b0f5a2ea645ae08917bf88d2a69335196976c794b2277903d934b5
ze013259b4d40c2196b38d835e79ab409f1024da4ae3e77adbf2706d72c735cb238c6ff40a09038
z9630b209945de59afc2f738faaccc6bd02a53daf339721b63633bd18aa5f00c92efd5b4b694981
z5728cc9e0c89ee80b704e49acfea085052b6c3e9f880530848a9b4a27a08b521d71f9cca525dda
z23d0ed256507731a12b296fe295b2a2a7bdedac167162b687e77fe239f4efc40457411455295b6
z244640913bf6b115f35a9c7d3d1654c1d430d89c916f898f1f579a738410d1fd82ff3a44539224
za677ef4fdd9e7c8b11a8bd9e35d5689e2e25da2a427232d86bef1e3e2b2a065f181686a04594ef
z290428ca5d4b9e9f844ee1b6bd385c6091c4af2e3004dc07275108c9366ed221b317fcfb2aa585
z979d0851e36d4acc1afa549ad022b436ee920b9c9c002de773381dfe8f1b321e3d5479c31f151a
z6db83f905d7406051e15be667df7af3be2c9f5462713e162faed6a240bb196d8fbd069b37d1f82
zc7fd9b34657dcd7641e6a98ebfade3080a003342b51b6d4c889870a2af0728a98857bd2ac05efe
zd99b8ebdd60c74c664e00aa49ebde9b547fd801987afee74aa19c8b5245f8048389654840c1f02
z19f16f9159b2c975ebae4c48edafa1cddcd6e2404c7d7725d56ea0915ec7db981ad25cb5a7206d
zb151f9ab42853dcab15db179923a12c33c0de0b307b10d8fa9c30d4a9145f36293349b68547e9d
zb2f540bb0a38b583ac07bd4922eff3236d91c84948bb3dabc1e0f44f7b10051f5f3e9ab11ddcf0
z326605ed47f64a76962b1a065dbe5229521e48d195103ac95c973f3232fd40502cc4fe0a6c39d3
zb46a475ef6cdc9787343d34aa7e0d07d341273f01701a94db4adba2071418886f748b73fd26fa7
z76eed4704627d9312eef67c01e90c1750ca246bcd29dfe6f0a543f94637f4527cbaea88b07dd03
z5d7127a49b77679147aeef0e621d46238881aa16d9a60afc2ad8d93ee188afeed2c8828d2aef9e
z3e3fb7413895f74a46b8439792d1ef914fddb0c99690d6b58e6f95142e098b91586aa92228f4d9
z43fbc94e538de133765e5a67dd3518a871b46bfce3699cc3bd1b1002d56c3a1c7c1c175a3ed3a6
za0ee0695aa2fa54597fc8cc812b5b445419754c0681b3de929c5efbc4964bd60a7d7ab6e622622
z2d13c4f1265ec9f3b00041522a6907a8c889a360eafd0d53c64fc14cdc1c15f213fe13149e1b49
z6267e16146ad0fc8210353d5a2d12335b399ab68a307bd841d56d50ba40e14333bf68913ddcddd
z05d73303e9bdcf739d0447643ce244f037e9178a3d04ea86a7d6f2fedd118570b6e44def4bee82
z8c5933bc3b5b97604d1eba03c274fdd2d88c492a6601e01fbba73dbe2721b0aae714a779a88d2b
z45867b384ba32f25608f6eca61725ed3fe423e13973114c913eaf94755f5a15ede5ea810b97e52
zc1e3322d95400fdac6bfcae4571c0326de40a6f1942a12711c6a44a90d28e58990e56529f286a5
za4bb3d04a699a7a8b8e35c5fbf7dee07b065cda9115f4a81c71b3784abdbc910e568cfb2f83898
ze4fe8368a53b652499b89260e79017e7ef15ee50a139eda97eea37479efd67c41a9b58220b9339
zaf7bb17a9c7982418d27bc2347dea89e8f3f1da9d464924df1a6b7fb8d7825f74e0a2b4d950440
z08a1add2a6e80dff729edc7992af3f4e2cf6b1547eb0c881d86b2da1fde8fdec915d132ce87963
z98981273fa00d0c7f4ad792da80d358bf5dc7753bf8ecfefe3c3d724bf4148efc3a17e61d5df8f
z28f4304d0f61aae42f07611ad1e9ae503c697e1c218f395a73fe489a29b882fea8cf62a471509c
z2a10c402eec4770d44ac7dae080d9c74d16024307f5e2055717ecd51abd51db1da6114d2f295b8
z58fbe11bcd8c076ac5231e730f2d82a0248875df38d310595444e65c2bed8ca2742bacc8a6faa4
zdf325082741f66c724a62fadaab00d69a70cfa3bbe351e423c1c006bab4935e0eb75bd65762784
ze858ea870346a2199ba1613150c9780f168e59e7cbd349881746e7b8f73199905ce915607e08e6
z549b0b19ff136b4730257fe089e7c7852ae3f9c76ddf23098d59703c83c0739d2e63404ac4f9a9
za3691134b67f4c450b227eb20521762be8f0fa46a811890bad358c176945917d4ed5ec54b79706
z8a696892c91a3069f8b104e45ac48640b45bf99031ca2f40eea42c342fc8ca35d258feac34aabe
zb450ebf5ce624dee75829eefec840bc6b3a3194cf532421ee1fa0d80d90580a3538a3a4c7a6a31
z074c1f5d59ffa80bf55f63a86cc104e78cc726fb97b8505d2be7089b2adf01f2e9c897a04acce4
zd04458c4185f629057d4dd71d6c728132693ea5b268a12018fdcbd8eb19fc4e57b5fb601a77e9d
zf59e90f87bf9c171d5d455509f3596c42c780f3f8c1d8a52221429f34c1884452b275d50a65cd8
z419a3f10a9e35f09aab70b4aba005f3154cf5bf852650875f5bc5c02af3707a64fa4886e211aa5
za0f89f12f05767418057c23c767d6498c66033b7b57242a84b937a830806cf83c0801edb85cf77
zcf2e897e19a88bd54e6c53169c2a5fa022847a1efa14a90622e38ac76f2ca229e4b44a8220a6af
z5d063bb5feb0b9d2365173f62cf747aaae3ce33dc04d7520bb6e02fc445ae58ce12a27703f1b1c
zff02256b7d358bd9564d9a9911f96d2fdf983e1b89b58a1f1bafafc712ed69f6ea55a75b697497
z9703bda362069709cfcb3093a2272fd39a9b5ae6109274b5dda20031ef869fbb9f10254eefa76b
z5d6c77c1c0da00f266b5e06b632f68900b4a584fc2d7974ac5c5e1d62c23fc51069dee0a92f73d
zea9afb31d1858dbb00c2835305d4bfaecd4772d2bc06b1223dd9fa852f6250b63766438c806bf3
z5c18abc077501605791642a3e38ad3cbea5cbf3cb41fd326cdb9ba79750d20fe9a19da096679fb
z6743e3ce6f4fb14fb59c3b631780d4c6b70e6c55a0654e0937a13f3fd8cbff42eb022c40114238
za6209e92ecf17678bea0a4831cd28de20c99048ab7a4048231fdaaefd11bc855a44966b5cd1a4b
z4c1de856d769f68771f2c6ebac22801357c9f72fc94b2769bb9e0844928911540d4847c537b529
z0cad14a3f63a11aceffa435987edf03937135edc05862ec714839f9ae262148f4b17e62c292162
z9b072e4caa7e2e14ae4807845bdb6f3cfad95e7ca133d5a5b925d6fd40a04cf170b7f707192d2b
zea74b870121c388c50dd341254403b2d622df6c163825a21cd2fba8efe9344418fd126b45fa56e
z54aeb7c883279d4f4c28a07ce0f29de82dae2be0e2e49cba2d5d436b54ec88b8cbf855d2d4897b
ze5f4e18bb872fc77a104c75d498735d8f676607bef2ab396c949d14031185dce455148dc57a3b5
zf8f3f19e3e3e18669d4e6c0d41a77a4a7ab02d7f7ce109fcf7639046bcebc7fe3b902ecee4edfd
z143104d3a5d97d77267b0010870039894544b31465ca66d60535c283b17feba8a6f39e791eabb3
za73ebf9675902e87c5449027759dfabdf813d97065f5d7e8b3a82eb0a7216e846c8e5b27687cb6
zd10b874973ad37d4fda5781f8eeb00525cfe74f03f2e4bc7337ee462c4cf293e822200b45067af
zb18b49434b5d55845c1e10680f2ecafba10a12767880f54d29b025e9310eecfc52302c1f8d4287
zf9cd5b83879c30d20fa828cd6f13d52ef9229c6f61872cb6b261663787649ccabf0b74c2cf8de2
zb783def7233dec299701d56b7b35ed56a59986dbbdd87e2352b80bcedf58268f8d9b7bc397dcbf
z20b9fdd3adcaf01b2daf444a765f52fecdae14b9a4ed4084e28579d86bc6967ba3e3a96f06e06e
ze1764d51add2ec71011f761d83958b250a7328a81a4fcbc7b1de1904943cde910f79c74c4a4c0e
zc7492883ec18c3955095abe86dfe494be953ee9b8248f91689adf6305ee2ccb08ed644cf530ebf
z22e56a891b133197fddeda5522ea4af79be64b7bbde108d67665fd9a2b2841a7a69eeb66d80465
z4771293b3cb56cd05434a683b708672b322c5b189ae89b3525d033d1987bfe17613787781592e9
zd73ffaba24dc2e0ba7b6201b3a2a5161a25509a6aae7fb28ad676fe7d7eddadb86a71a2eb76ae4
z2a8997844cfccf0589bc61cd6a5e2db1ef2fcaa96e4b6ca367457c58a16a6071b0edecd2cd36ee
z97cfe9147c9234c5ca28c8c1186fbb4137e3f1ae002846fed5f6765665d9505fe7449d44f6b16e
zd200ee0eb49e926d9c6e1d5ba7e8a7f0e5a5e36dd6c83e49930ebbcc89d9446d2444a59004cbe2
zd5804fe3cf9a365e1ded2c017611ed06c01d1fee86701b9d13906fc4ccac558d375b9c96389dc6
z96154bd6022264d8efa63f01f28f7d6aa5b208548e251396d401d5df4b0b923e79c9e3e0f6f736
zc999fbf399c49ff44da05152d1369af95a19b96b5a5f6b5e09f9e07905676c256b2f2a737b2b2b
z37d21cb616d8e491158bb850ba3c64250a5a133bcfeaa770f1b5f9fbf277b6f7d3f82795a2eb8b
z901660776f2b0a66d9c85205c70c0adb27f55b5fc1f6cd6d1d77c0995146917b0745d3deee46a8
z3ffadcc9dcaa8b72064afc2b7224fdc7462d19207bdd5f61735895f09a2e056c35131b93aba2a5
z269751607a4d4a49b74f4c0b63af0dbacd0563f8ca36c8612a740488731e8f3c745bd02cad3161
z318b02770ab561f1fe2496fd936d6cb48cb8d83384f426d419090b30727e93fe256bb6aebcb14d
z193427aed29988567af6c3cff7cb57ad0a490433c9b178e77e65c2ae3ef46b40355df6dfff2a6c
z3454bf6713578603406b0e6a7c14c1377101ab3293cc46e1d2e26002686c140b0ee9341c5c480d
z567b5d5d6004d83273a33d7359994159dcb514ca27d59ded01c365359e744d2738dde9ed1b366b
zddef0882fde81648389c85efd22f47119cec8e544fb30062be69f6d8ebdbe51d2d05c5d0541cba
z2c202391153fc276319c5f5f27e9d52d292ce420408b55170f210525dcf14c2df78dca4a1526be
z45beb3cd73f28a9b4fd3c3e2b72f1fac576a48d6f84bcddd565d9681e8382b0b44f45edc20bf2e
z399735fce576ad62aea2c0e30bd9960a3a1cf2940180b7800b5a6688d54d7af89005b45c0b4d55
ze6763c42b7d326b3b6dbcf5e5f4ad5ef58ca77ef49290b3ea4834a8ccdc57293ecf17fc7aa90df
z558319121a1e5a89c5f23c6847a151f9690daa05427f2d91b7581b65afd4a3243f5c8808e8d586
z4abd532a30870bd7794f477f924ea3f570a2b9b649d7ea891cc71432fc1d0a996adc2748fb1c48
z74645043299a4985e2cfb5ea9e74100d541ce58b1e8df710393b71dfca4e25829525adb31bbca0
z78dca67fd4f78f6aa36d1908151db2413d9efbb91d43eae71683595e734fe2e3f8986352e55e1b
z08e58d4cfd439227a35bc5a10f0c176da00a014373a6f2252063cb828c463e470a447d4693b0ed
z5747296b847ef33b4e2ac09c7e41e86852675e7ec6f13aef75f5d535e7cefe5d4d2a1ecd469ba8
z58f7a76241469edfa1df3e1027e3b8484e608875bdf5b1157378c284e66335f6656d525ecf4a42
z976b9745a9d7d5ca9c0c6f6b0200f5d9bcd5c90ed2dfedd9bcd0dc4773f4457acdf745d2b1a027
zb7986d705ae431916ba158350580d612ea9e55b0713301f6f0754ec72fd188fd8cf767a957cf24
z5e383fa76fd7f60a219834f1e3a16cd732b1515a8f12130b1de5bd5cf7005cc4f48a8e430e4c7d
zbb651914a550332e825b942857b52cbf290ac046aaab123bc3ea4b17a1ca5be538203bffb224e8
z56762351075632a3703488fbad746266998ec3e8ba5ef0e72bec17a202b5474f8fd2018c3d1532
zfd4d1d70990949afffaf90eb24e07cf2fa5d3c703a5a7bfee612b6c28da8dc2ba7e6a3456c6e01
z6e19009eaa948f01185e2708503ad2697c5cf7b79523931a2dcd7472c444c2546af4e5abc6069f
zb8abfd5b3a7e451d1b7372d387a529a42bad52236e575c12442c347d1d459998a5ef12defcf04f
z2336cd266abd390c70880ed327bbca2628ab930a932e5f52cdbb8c219b33abe1feba9e726b359f
z3dee13e399cd938b38d2cdb342ab0240a08e3dacd686167a600028932fca5a9cf35586b766036b
zbc18493f676e0062fbcd8d46d46abc7cb26d10c7d928d6f237e94da38be98e87c1ce40de4e8139
z9ee72e908ba700dbce681d7600a487dc9d0ac91a04a781f252e8444158e17aff1a6d91e25821dd
z7ce3a9fa2960b0e8ea6b5eff747a6e8ed7c63a5a76253235a3dd2edb9d1eadf072ce720552f206
zaec165657ddf962756bf9bc9f10fcbb5d4ee3cacf2d07997db63ca3a1bd18c0dcd0adb6fd60059
zddbee394af8f20657462ea64c2cd00f95ad50da4a6461e3fd81f2792cc48d27667bbcdef9497d7
zd5b1d0ef148a56957fd3d793f1dcb3384baedb0f20d9a6725a5855a7630ca44244fae7746fd4cb
z99d2c98832adef76ae32d53716a60cd90fb1bbe192b7a9b1bae80cd16907a7acfec04852379780
zefb01db4e743003e6813daa40da1418e6db74a7b6e7b615c2d8f691a9403358c5c5fabea6966a8
z63535594d344778e5b73628532b535fe1498ec69e0438292f61a705a82859e32105ab5d349ccc4
za420ca6ae65d67f69113e110578b8f6b614a495518231d891214c396e9140ff0f29194b32fea5f
z37db155100168c1c4f257829fafafbacf4b34bd3aa449e74a314ac35cc36de2fbb56552555e013
z598d654cb77140f0a2732b80f48f212621937083f7d146fbcb36a4f38ba14ac94065e91f1574e2
zfa2bb780fc1fe5a6dc0d7032f2118243fc83065d8c6631f6fb9b43fe06ce43b99c9e7119813c94
z00b23a97b4327a5343ae9f88b9cf5384bf24986c6a97e0b256f884daa060fbb81ac921bb9fb32e
zd5008ff43986a288c9843da155c07ba325a2d7cf578d72b47861fd1cc6e529565c67d8e7eb0ee2
z2338fb5620f5ac3c71f1f5606457ab0030b930f10623742328e98ee1b651a7741f7c4f441d1b2e
z273c28e175ac5bd7c37a255ba9285685152705a453e37620286b582d8ef6d462163cd321cc26f8
zb5db9747160afd52a088cd0107630bd3f508dfd69d6f023cdcb243de6ff75b2be2a010d11b4a88
zf4340e87d8f84b52fe89ba9eb6dcbb6b2cf13d576021bbad3b8c6831d600441451e0b7d286dd84
zfed8abc53f7aff2e3f1618ffebd7ee2ad27d2e1867014fad739d4f5cf30169389a01119ca539b9
z373d7286e7b3a657c13b4d753cdb72684a9915a96495e4b086ec68161cfecc0d6ec8a637254acd
z1647bcad8641e70df0482834bc9f12afdcd77d562a26173b1f1ea1b18eb102e82bf2ed3d55909e
z05d9f967decadee1efe48462fa79760158bcfb9e83671a565da8e602aadc0842ca5f29a8cf083b
z7a762735e4b30136aee87480c254b0c56e20bb62e86bec7b099889bfe7da293ee3807a1043962e
z91c584446d7562a261cd55e78a8cbf8337f161453060a940b1a2d32fa7f3d37e8902753994f4ba
z012ddfd059c9d7801e38fe44f6f4900f034b65f3f17d28239ceaf287048c07c4549a67746e7996
zada6bed3f31ca62b4461e903715e6a26655937389e113f1c9578b31d88b6c3d62c3b7b7534a77a
z99fb00c7bf7613631ca0c450472c55543ab113d55572984060c6036c07f7f99b3116e539c55604
zf2121862ed3d4f3bdc5847dc6bc6a610adbedc38f1c3c8feab6490ecd9ebb2b34e612def6a12a1
zde3cc7b0f8812401c9411fbcba4aa41471b1da80964c87f1258a1e1e8ff39ccf68552cbff93252
z8d3b7e498b4d84e3fc4aebfa5d753466f66784f1934fc13c2fb5386b9998fe13e9039c531b2333
z2d4b25873aeb4f06fdb0e4cd1a3959b7471eb7d07d12f289d1bf11ee5453631050553696f585de
zc9d904ebd25e0c1a38e71b359ed0833985603dff460b76f7ae98d02d0784a46802a5f6f77b8be0
ze4a35253b3eb0dbdeb19a579eb2831b6c90f552d522bd1b9c7004d5c2625027ded34d2522d9430
zad63c515d99c9f9ca1e14d35a52458aac040b470d7006d97ead22ae553235979d37f0f021dd66d
z084605bfeb2a5ccb2bd056c440b2e439da4d03ce6cf4b65e61c69a6c0428faa36b436257a4f2c0
z521472b5543a261cfa4b48c7edee94bfe39c03d533412919d7dc817a63274ffd79486f9f84fdc3
z516a523a0167235397592c622124942caa3488e1df04703baf5de85b16ba32310486b6378cd7c7
z6ae2f791b7e9ba11a992b6990f1bf848b52d2d27edc3645523ea4373dcae9cd3e512b2ebaa2b09
zd990797a72923fcd90ea8cc4a18531077197a66f14fd1feb3dbefaf69accda3e9c27b1f42ec988
ze0827f5f03863f9f7832d399d115d1a3ccf36c0a39d2591f3be8300f9a1488496427d58dcd4e3c
z80c96c507410aba4ddb27c42713034d4f9d31526c6f41997552540a1a6203393b37f0b852f79f2
zbc3de517e861ec39edf2d15273a97493982cfefd519f2fe30e07742973488406bd8d5e843f1848
zbbb2b906850a8a6b0bee7474a324b45b02dcdc435b031da52421d36fa0e7e6211608c0f88894e3
zafe0d10aa7e80bfe36db27e48510e07bdd632d0c1c241629cd11d8c8d8972309a1ce6c606b3c57
z31fcbf4c149a9d496233f4924a19e20eaced0dd8c5aee7d3af9d143984f5b34b208592b58e88d8
z8f0cd71aa3b71569dfc3f59cd4cb3b9231817424eeb0be77202848b589faa0d0feea0e907115dd
zb0982447966599ba201334ad49b76f34fb675d355aa251ba46a9c3938c0086919f1e78ab62b681
z8052be04e84127e387f7735b2f8e7d6c914d8a71f38cd473aaa7e0c8ef90e527109dfdfb441677
z1091b25daadcdd44595f72c4e17ae05870be99487cd81dc8ee841842b3458c38613cb5cd18c376
z1b50dfe1e2bd0d2a63fcb8075828b841efc09240bbaa9b1b0a7ba3b37070c7d6ab777e72842858
ze0e3e23ae2e06143b1b10a3f465e65ec9652f548668ac76c4221b3c307a6dbc40b11c2fac10d6a
z511ca4e56bed1a5a8ee19cab8a5addde8452652e194df01f07af8d65a8cfda5475d32b3f0f154c
z23e0520bb4a9b6c91ff726e057d216bf7c704201d1962447ed47b480b6f8401f5bb6b12ae24320
z546bebab35820b5b843ff6fd66f4fafaca5947663a63a3696b58ff882f464b5282b09b961a4826
zc0eb0c3f781305216ff2b3ae03c565ef11a3b8d3cbef72ef5a3c384f9a9f521d4d06535af6b7cc
zda4704a00141e8eaf6d7892c93bc05432cfe939ad4e87eafb16b51bf35f5175b949c6f0486029c
z605eec9e86ffa982af043c2027d9aed383fd7279cddaee3d199fa00dc61241f7834412bcb69d25
zc26d12361726f3f2743a015a266a225840c6315a1e87ca32104121b45d1d30da2574355d133c8a
z5939b323c1288e65a49199b63a89d3f492a2bfe233be3106390080a6d9001a2a68ed17a6030eaf
zedb0704f2e0449030f2f0bd8c8b99b180c74e5927e44b07fa2daf0fdba616248630f3c8f9a0f50
z4aaf5633c4beacecfdd8c0c0d8920eb0411d270b622b6662bbd549c5fc5ac35eea14e046667760
z4f10bf364d939e375ecfec993ac3d85a2b2963fec93632f15a6550b9cfb3031b045ae600304cc5
zba2d52ac99a901caca455fe1dfc0f20e85211ecf1bd0ac5e9d271f89be93511963a291a4dc555e
zf317d1e4a99dfbdc920f76531829ebf4afaf0c5b957240af532c03db86f22611a46f66510f1e4c
z4fc3a6ea42c07fc55ddd5d3b3b22aa75cb3adaa72f4be14a3d24a29b0db3b08c1109ca7ca5b6ff
z455ce6362caaf317144dc50d21ac785254d21f7c2016012aa1cd640309a85ae77a710327582184
zb49181a917ca5297abb33fdf30288f95922fa13e15bfaac4f9268769e8b05ca74406620a7745a3
z32a820593e23ecc03019703f0171066a3dcab302784e284beab1b9867d4e8389adebd71273e31d
z064c72253c84ab11f4399f04a03e420043ab7e01b9622560e24820e8eba73c309e28cd3c90155c
z596566747aa96b33145656c22ea596b1c20388a63ccc9f91c2854f56f4345964330da1081d7853
z4b5a8a5bafd2a931f267d5299b4ddfcf7e4e785cb5c3485506daaf461f8c66c6367736291c8df9
z58cb4964fd09624371aa50a27700e9cff417faf9f54d9d5000b2c8617ed77fdd773f2be7e1cfbe
zd28bb8a2c9da7495b4e85e6488959020a20c97485fb91978f4e3408f21a6c620c7fca821703190
z127412d44874fe8426cb2fdea6fb2f82011fdf231a0589a43664602641101dc18d89989b8cbbf5
z55c07cd7a06310f3de042c097488e19eb722fe8fe5066f23ff26192c48bff5eb7e2b9c62ecf5c6
z84f780e1e2997bff7f536b9ab00ec933a62e4f3a65879f0ee5c9fb14c263d272bc054be263d323
zd61e8432bc866eab6bdce4ade527f69f9bddba2b37cf9cb3be96204e2eeb6103c9b9c2d6222013
za859dac27135b266383672125789b7a29c8740c69c40be281d559922861384926d0c433c72c252
z6f830b6fcada1d6914af152faa9f4af4b1170457dc3036877886a02f1c67a23da65892e3c471a6
z932670b9d6c3d12bbc9ca861fd683ecbcfa19d1ab96a8fb5aea5e8610227ff7049c576d6e1ca29
z7f9cf9256f2b250ba201b9354d3cd5dbf26e15c2977815734f79ca997a044c94f4a7e381e3551a
z7976922f2698eda846afad1c084649edccc28b14fa8bcd0b437354f08924e394025dfbc915c7eb
zcac7d325239b8059b41e1c8570eadfc8fae4fbaf7da0318a081ca6970fbb672e32bc7095957779
z2be6dcf81d70fd5c55aebffb145ee172712b341be393346a259dd56704bc7d9b1fcbb840b302e3
z2b54670cb8a88e8aa3aef43af86ea49cacee977febc27663168cca1f20da1f9ee17af3d4e437ff
z1ea07dc2f8def3caa05ba502413242a00e6a8aa65a0a6ee0c972230ed9de50febb8df72747d5d1
z9f1498ec4f7bc1c44fca34660f29f5a718a515bc3f4b62be2c671d6ef975007b2b9bcff23f59c9
z5b16275bbe21bfdcab3e9fcedf81ba0635b0f0f662bf092bf51be84553bfa69ffc79b38fb64855
z0f51cd9b85c783832ff0bd9c92bec22837e5e486a0f4cd41fea6aeb7c38e045af0aa0d9ea648b2
z1097bcfbe129c79ce26b3717689f213cd77e27f7fc62e3c85af98d28efaacdd8b52a41073342f7
z2613b96708cef3ce74a8913e2cdea3542b4e45e1863e86e911873280c4ba4aa6e8e58c8a838297
z485ffc91bcae94a7fa8917200f814d5e0d27e2b124548eec2265183f7366232df75f8da2ab3ebc
z56409d46c5897c8795ae81d0a75553e5bed049d8ac21d71616699462fcca41d5e9a85f071190e3
za2b19296be2055608fa914005ccd43df32905010e51949c23abb9f615b7e20ae34b3f8e434f2fc
z6b2c17c0b55c5e9969abc3434bbd150ea493219804f9a2031e6c36d4039b2387dff2c4ed1fc568
z37d92e9e0fe6d97b85ed23699c8909d1bad1f6c19713bb5cbed1aad0532edac8b39a1db3f87a6c
z2814f0c3b9e31c14bf9b75261e25bab372f730a174f1e3610e3131d2c83467522e3b6d504edc2e
zc9381c9069c0fc5f1961630a38580eb02d94944f51b772d22bcdb80eded3e3a21ecb370d919950
z83884f67b5dc95323f8e371259e852519d3111e9d589d18d8319ad23cf51b9429513c289353b2e
z0d316174caa1c2e66606c29c8a7b03f7d780d0136b66e4a2273435fc211bd2963d8b02f983b6b0
z5b6406aba788ee8193cfcbd4baff7e34779c1896f7381017c223a62286072565902c7696be8c29
z14e058e22b94b3fb8d7fd69744519cd8367b23bf05aca6d88bb528bfd826d53192676cfe03f9c3
z4e493f7cb4d48a0738c5f02ee8938cfc570fbd174fe250eccf869a7f0bbccd12f95979d1bf1339
zc48f72350cd2e71800f285674e6fd47340f24d1306971e50c6787f7a52cbf0443ddc8a435dd194
z0ab84feb1f6e341d32765633cb4638da33bec927ea8d2c09513f1a108090e0bf21aa4ef11e8b2c
z8239124a8383a60a66216811e5a68f6de1cf3e1217244aedbc1d10ae434ba53471a3978e2fd844
z2c938377e66a4c0f277d1d153db6a1563a01515dc634e67baf5d5c80e32d2ce588c40ad7634905
zf2e90a2e2560566453e7f66183e1638209e7a888c13906f195b86c802f89e8b66f4c9d79cc7b4b
z6a267ac673e469e5fcb9f2c955af9936596d95dc27647bf402586705d0795e47d477fc6ac92e2c
z395b5d335316cb45f317d98a012337a8b731709a0b0be9a22239624212aa3efe46b20ab9949cc4
z5ec0fbb7423199a09c20085b8d3b95d78699413b8b706acf01356cb6a7e1c907787f1d8b1aa8cb
z5cd76ca873bd17a6999d03adb6cbee14de17765c4145847d0abbf71b8430608609421cf542f441
z3aa030c77a28c8672a905a948dee82a305ee2c20faebe9f4413a44871e8786140c450715ac1cca
z27b6ff96d5ed2a4c7365e123b61c0862d2eb00fa790225389188f46ced54d6dab6363d2612646e
z97746d7b6b03996b949a1b79a873bb2388bee593b9f63637282655923bcd761952e3a3d8d90e2f
za8d2102ff5c1f0023ec5810ced86bed26694529fdc06ff91b54b53d2e5746b3616472d05a7ce89
za4973971360fcb48b0e34ef53906a933dee6c056344d6a38a4e55166c29fc6cab22a0e211c5c8f
z36757f6f0f3f2b4861855a98acc132d0c4ef5c68989c21bf7d64eb0f48bc5cbea02136ed3fee0e
z70c37b263b9efbd6b990cd85491a48db4c4d201084b372b4821b53a3d51496d0604d2b2d8ef63f
zd349f280eae1fbcb85c53b4155b0d9b18409a6b3c0a7032a89de00f5a18cc7302d6ba8cbb0889c
z490ca281241ac3a26d06dd18dd3ac6af3534740dcfd8ec09a13d32793fe1fc373a5ef99ee71c1b
z9c7e5b7161f1ae17d02ca2f5ff099e6cb5c07d4671335436bd1d689df80e8d0fb1a4845a4af588
z365267f1521f5b532958d251df67469c1f4d91a1cc46cf3507b38c69546567abd064e7b447035a
z57e5dabce6a6d8c095155016fb5bfa59845621c883cbfff084bb5f138e3387b5968774f11f7d69
zc94ab8aba11f3d8b1314a94bb50d55e56362cd5cee3ac3ff4e1fb1fe13ceff5f59c57a84ab5691
z3d1ebbf238ea7895232fd5773e6414fdc1a47dca7c23e236f6ad8695ccdc47b8f40b408625af5b
ze35ad37b987c717ba7b2209656f8f7293050bc778196672ae14d1581da4d4dcf1f20a0e02e6673
z395f6ec0304a12e3722d0e6d33d06bcaf4cfb6249531ffe5718247cdf8d5e61d4552f5084912c2
zf2871a8fafb09d486b9b7beebecfaf9a762e78132553436b656d37267fcdd4a118ba0c5d62ff4a
zdf0e959616f8cdcd8f409b88cbbc12215fe049c822912a2096c6e02c4a8286267c7ab15998d99a
z5007f1cf0162ad99b3c97f9feb3c6ef227dfa7ad7b8df35e97a8d6d476b6f0841848668e998e9d
zee0c2972a5f9f388dc68cebaed6755011b7733a6109f82cc44415fc879020c5906ec34bd1ae9e5
z1293b017ac7091f16987aa2227a246900b8a245832d2f1d137e5cbcdeeb3f1379ea57db570bb97
z55293370f08faee49c8457789e3af8562846860206495fd26cb8f96e78df124e6d11991093adeb
z9cbfb003959f67afc840e2dade718877bc5f9af130bc385ae9b023fc6deee9b4b88e49dc4a2102
zd84fd07289d1aed6e0c2242364a178e2b29a0d00558839dbd46e55bd9a6ca41387f8b93e623047
z4b074b9f2002babca36e2fc0550402912459f7769cf413082cb61f3f82a7d6678f2cac3be3f5b6
ze55520aec5ed4c5083d776b4b16a40966cae27df8ff10279a4ba01e3761c27134de1158cf3f7de
z7538d2b2e7076c3780584eb615fe2c17e9cdd38f0d31c67aec84e94484c9edde3a70a76922ed2d
z20057852daf005493f2f77463f12c5894af4c6a6dffb8fa2e78a232f31681c5138c26d11ce8bb7
z5dfa0eb300dea62c8eeecb8a5811261032c327fd4386dd17b7e365e015c1f5d4978c22f51fc760
z44df57668c326ed1c10f550888aa49bb096076486b95c594bc8733c8bfb21ea0121e24727ee882
z643bc9c06b436480cede820d7193b029cfda1185b63e909ada035088868cc3ac99e1107bc838e8
z7105085840cf4bea2ab8254dc25306084cc0a5027089891f798699c264f221014c05337019e46c
zb6c7c980aadf2b344e1ba118efc77e7e590e5205bae06855ae79f4073e418904f99b63f32ea9e3
zf25d32f818dbc173ab6a6c82dbd3f507a403556b56fadba1623da9c155e3a7e4871e3ca5b9f8a9
z7f52cb960ca9d51f8a66d49043cd949f7ba3d9a94c3003034eac778b6488b7a349ed86074a7320
z14108f4e96375748d6241641d3ca52426bbdbe956fe8256b8dddca019ee9e4098ba145485f0c55
zc7791ce0acc93e7c3d7ad3e71b631dcdc71ec3bbdc98e3cfd403558e4d460f3b299c45c5f9e306
z7b017ccd7273f633517cab5b98efd363e3a821bc4b1237ba921b75d1b956fb6d506631f7f56e69
z1376bc0aebe318c34ed2b3dbedc3b9f92255730704daf1653f259db299df4fca6364fa5c569c78
z17cfb905747cc21a6c252521dd8e3f9643b14113b5ed702561c7edf34a7f8ce8da3d051061493f
z187b5c05fc9541b8ff2e2ce661d160006145e7422f56ff3ac144397688e4aab54df67c02a7a8e3
z5eec22424e23d1c1a8bc9e7c506535a09634081f0e7030ff093b7f627722954498c33010c528e6
zd0e2076298269da74fb3e41d8e5dc4dc38e5ad5f79d7276a95ee712fc626940bc909f72364bd00
z7a1b90fcc85fd52c06fc5e4d9f41dfc279d3b30a3cb8b5394a9a246765fa438494d2feafe3d8bb
z82fa3e78936dd4941c2a1072c164d3bf09235ae63faac72d1fb262a75dd451b34411fc3b3c98c5
z0820c2b58a4625cf06ea13a8075668f2237757f09c378a8c64c0aa50da0fa7e63ae22851fc82af
z2aad0b39707a191f14c86e089d726e02613a4e5d3f9070e46cd140a07de03dea5d71c6e34557e7
z438169a11827fcff49112e24f55c4ed084147a2f7c484377c606cf044a80dd12d6ef96a66da2d8
z7faf253657454be617384c608d1c9eacadd6305ba3a4af93f86a3488e1c24dffdcb44ca17b4795
zdb37eab7368ae6f0c1c626322e81683d20148b84088a5d1bacaff549546f27957fcf32033960c5
z61c282ec4c6564572b2869e7c7a3f52c45f1f3b72e8394922e83d7cb42f9f34ca8fa52e2907e00
z56a9878f34e77442c363a9b3ba84b4b5216ef696f6ff7376f5861e51f32bb738f9e03bcffc2af2
z57dfe72aba4f19c25a079ff292950486dcf0af9054e4721b1e0a70d7b6045cbcf1faffe25ee62b
zeb8e993a32ddfe8bb570cc76aeb5715a0cf2a953826bc1c464dacdf451df5c198991cd6cde1229
z2eec781053c16e5f74ed1131f0f060bcdb303fe4551c4e782ded3f2e660b488034e3c28752ad6d
zf66bf5fe73d1fc10abe4ea2097aaf270e5f017262566f41400ff05da911ee75e89fdacee7dbdb1
ze24e66beea3250938e2352389511efbeae1f0c292b9ae35ef1ad182af501a1f550af86c5c6d071
z61de143a501f04c19ef201ab94ab6691a0d0ed352757a9a56eb4ac72e40fa6fffe068a75a346a1
z3eb72e0cc36ef735742e5ca81b22f4c79781738de2e21fb8ead84495f40f5152b75c4e13841dcd
z9d00fa8b729476e94a6d420e53d2b6b7a6c8678cd87e6bde32f6fd984950824ec04fdf887475bf
zc070128f563726cc972f924154fe8377a262d8637af762f39e0108809bebe30cae62f282faecc5
zabf1d01584de4c62257684517328bd96b0e66e856806356a9f77e56132c2582745de9026488010
z6715e2f4ee2e336dcc4c01f390f8acc8ba0814d23731a4887addc86db6a908ceb0ec096cfdaac1
z284ad39c2f0c2ac26a4fc41c2b2019001fe3b97ebb2d7b511c3ab62c4016d062b86135c8d4f733
z71f60e2a2cd8a6bf1b2d742342f100f94304c58232abe0050945125caa34e50e808b2ee1571171
z2ab132549cdc0796d0a59aaadb01a5ce421f1ace25fe2cd7fb9b695e6e993eb6e83b6c6d237bac
z761c9c0054b12ac4722c269884f916c484e6a8a939650b195a196538fd052c1a23d50678819089
zffa7482a058e78b1c65d9a428acadbfd3c3877729a7fcdcf99b0402d2b4de42971be1bf3328986
z3f2595194454b8f4170669cebbe4771098af6a1e979876bce8939f5a0cae9d6b788344de3f4aa8
z28a8d134542814f8ae82670328825af65172c046770d04f0cde5c56163aa3f321fb33d2952a377
zce23ed5b8a425d240b1c94e41ba7d29b9388c3587e21be291f4ce6a9de9d8646ba4b9c44460353
z314a4d16d2843bc0f8e44432fc92a9470508d2677ae87ee15fa8e459758c437df6d1172da12fdb
z8b203a8b254a424dee8237d135262333f8ade162d5f8a1bcc64d917ca426d9248f4b71ee5fd93c
z0ebd7860adf2456e7a9d54dbcf4d1a739c88b528ab623f539c8139d2dc8ae4a491063a547353c2
zeb1f51c2042b83a868b99784df1059d1c01a4bd8b61bd949b46f5923d35e662bc382dd36d02876
z0405e3bad86ff9961365d314989c6cb194b72996af13237a3707c2e14f40dad18f53769b949f6c
z4c13bff3e0bdbff5eb5ff7f2862b4470b0ce980f8e1a1a9edccafd59cec17bdda5be445c90ff9f
z660b170cbc01f2d7b0a55f3f16966e354125596af52691dc797f0004de6bded1230a43cbe2165a
z58066cfdb4ca5a00b387993f390c18f99c3264b136e231c7e82477a350fca72a5d1cfd0a40d1d8
z30dc4789817f423f364111449b8dc382c1cc1037661cb8d3e79ff35d5168795d021cdfc445645f
z6fa89ecad59137bb8ab8897f78926bdd22d10ea5f01b324cec3c0d492b5ad230392c212cb9f7b1
z3d6d8298e36c837a7a7d3eaf9c0932c5c04f4b9bd8595dcddb920b0a88a7ca4bf655aadf0fac44
za45d79a11c08dc505ce04994887f5494e5aecc896f09f7ad12674e32999ca94b492e0b692900dc
z1f1b806675d657a1ea591b2226cc04a8ffd3230bf31ab35e0119dbcf2f5abb47878ad7ff68b792
z57744d81916e3159476e878498c0bdb2175b653a5251aa84343113754e6d7fef7c6b6bea62237b
zb4801c6a157821cd58e60df737c096907219b693a3f1aae6b2d5dbc32fed5f4eea83fbb9916c28
z7b7e5666297ead1d71579c43a1f22019681524556a903ebbadd8cb47f3d43a876b5dcc1eb8f4b0
z07327a04f35ae912cb3639e307355670b9cd2c1f91f5c4aedc59335d442a889a1ae4ad9b179575
z25cf55f138e025a575234c7bddf5ab39cf895d6df4b39b6793a04e1f7b8d8fff78def86181bd3f
z8fab4da0d92550b83149b62846a2bd5703f65513aabf935b2a2c52559fef9089e7bbb6821ef768
zdffc70dd2c5f7737b0e524e2a890b0237fa55f8500a4e211135b14abc2fe7073fff253b5e90245
z4d59998781e56c41a33f990ec57a9123c080c41ac5feca0f212a2170feed25ff9f50cfce98d535
ze85eb035d7841d9f90e88784b7f4b09ec24ff742ff62ddbb93e7c15fc3319b6b68a6f3a2c25dc2
z0a3c50af4bd00619c00784be7e5f2b5de067ee0045047b89aadeeff7d1399310ee6d9c1e068a98
zed49daa6a5ba1657a295f39057acdd65d1673ab2e641ee3dfd44001d74501d476a6081f6944c84
z9ad0950bac07785286ffb7179784f53ab6df02201248a15c7d5ed171989b3dfb16b4f454c0266a
zf6c623a7984c76a62e6c195b587d64497e8c4133d1d19cf2447ec42eb1cc1927ced3d357bfc0ce
ze6bd12103dbc4a2240f4ba1af446d4435b21b6fbf2f93f405b754151c3209fe35c0f0628cb314c
zfa31b154bffe429c86c196aca4c571c99bac3a14d621888346cbef01e8a9c2fc4e8d16a1527f7b
z3f54b3499342b3952202fb21afb0afe23a3de0c52bb4966fdeb17775017273b1e03875e6a85c2d
zfdc00629ce377be4dbd85737a82980a80055559ea3b397aa691fa638b63e78030ab8913ed577bf
zb771433bebba79fb1925bb3d681eab6568a97e9c2454859b70ffdaa9f01f135ad98f14516fce72
zdb077ea76de9163bfea7a8f25580fce429b37286b8c6aeef5a8b6d993cb3df5258287b7792a308
z3c4e3fdf34b14784216a0b6709d53f2dc6738cfd0f38085a106046fb1059e7a2bc12cd57573b81
z64129643dab3c8ee94126c40cd5dc807842aa3d75bb6fc6c645b1c0bc93bfd8f4e9b49a827129d
z98acaff95812152fc68759dac64a4203930442601703a58c55c37ebaec9d2d0177c6e29b23876c
zaeb3f9dfc3fc6a129bae1c98d137e57ebadf4a8ed09dd1d96b2afa89c9abe73cf1454a2a8c71f0
ze144f33d99873279f7bf0080d4e6df43fed85d083f4061b4226a459d2175ef4873f7067574ff07
z4c89403066f0c5b86634934d55e7ea97bd887ff1276a8b0c2c5146079196df7eae38081b54ebcc
z0e4b566e6daf0a5584e61641b32cc2921d10f5ac5423a4b3d7126c90eda8ac02a203d99c192c6e
z9f3314587e449ae80137e126e42749504234ca245118fa81328fcfc15241eb78975487504ffc2f
ze67237c07b129feecfa15450d227ebc5378617b83607b478c9a35a914596b4a1409c5a42981db2
z6c3eebcb762e80f3eb8888adc30f580cb29e477c5680fb5946a36d0cfb2467dde284ce79649bce
z29f97ca41d3b16d03d140547a73b693f287842c6949451fa3a377fa4cf529f140414068d7d4bda
z99d8a7d88be3e3abaf152a390caef22417d7b63335004d9c312a7c7f97d1897c5da0e4e7fda7dc
z9e0b0911ec022e7909c8be3e5bb48b9690fd19c5055e346e38e7aa78429a57f1cce7000b094594
z01cff6959c7fcda072716e56cfc6b5f9c1d9151515b3e254c7aea7f7112c9e72dd97873b92b98d
z516e69525556b53a4bf816e6e9188d118cca5559a7107a0852dca3f26e48ef87e4aab863013b4f
z7b397be92596f71d59213ea40d9e8529ea225f0afcf7faede246c0fbecbff92a8470b7c3e71947
z6c5b7f981987429c3da8778f99b9fe22fd1d027e5dc22f97736e8ae685abec57db28e00bf8f06d
z85d06e970af32465eedd3c2be6e47491d77da668adab86291c7cc0e18c7a22b6d9e7939f29d328
z54074069b9916e2257054944ae4c00654ac419790d85854f78177aab8f88b2a823cf05cf807f81
z3d512d630d1a9d5b36dc43e55c62c8225e010d1663a7d9537cbfb0732a3ba2093c6e7c311a5006
zf358ca233028f68c0fa287498ff55e4ad33de7fc586cb6e077478401dc916619460cb490f9f5a0
z453708177668706f8aaceebd57674a3a2891909e87f60d6dc955beaf49eda7b96eeea3d8b41aa6
z9585e97d91428c2e57163206c2fc97a288c4b378a273d9ac36980414df0d6b988d64fe853e35a3
z2d788535444455edf678a6f55d1fd079c14ff4c90245a85d1388d0db82951694c5e45d825e2147
z1210c72c937fe2b359482f9299c4f741432590d3c3afad26cd03bf4e63aa88665eb6a948e59839
z1d229655aa4354dd1207622f87d085a2066fefdac1965de1fed4b1ea0fe72d7817017f3cc49a97
z7cce6e800aa31427f83adbe3678b65be4c45b8238a01c9370b4693095205d0c5284f61ce23cf0a
z593a612c9b5ce4e8d8e2e4b5df9b35d09e8e976dbcc2d3d1463058a741809ce946f72a98af865c
z330c8f79cfbdc07a997fe11e2e7dc009e43067332db57bb0a0840b8cb28fc5dcadf9d42cdc3962
z2c59aa53c39dfca0686f78cb1f65a0eec1bc682933238bf2d27c5f3152a1a033baa5285adcbc20
zf71e610b38ca6e85ccb88a92a41fdeec1b9b22a01173841ba2bc69ba318c2b3cc5fbe9ef311acc
zdc56efa98e0c330f8ad1dd77d6941c7346503cac83623996850dc3cf4255633fc45b0eaa65ba2c
z57db6b1d20bd3ff3ec8f63f661146ff7b68e5f4ac612a2f1f027d2c37583df605b1d463fd323be
zff51d0c0afb6836d8c642f939a5a6e11e2027fba3545f57f7cfd1c278a360b8b8a162e5279e8aa
z6c591744f7de320cdb8d7bb20e27558c72681134a64edbc945b01035ad925607750a2991a87d94
z20e993990fc708f2aa903f1f729705733d98bae436da45f5c9001d69c5f1a5bd94592b73595418
za643ad9240b6dd4fea01ad092a230827236400dc9cad7f2cd653aea1d1054af8f9d2f2296d9dbb
z5c85f8163d3047a4648dd5867b4dccd66bb20c74acfa167a2b2fca1b49379fccacefa1f60a39b4
zf0a60dd1aa9c5ae527811a97cea14155293798356e213cd1733e1fa1a6164603fd528c91faa5eb
z71f07fe879d89c4e1bc20afe828e5893c520f678756a673124f6dad2a06bdd78e8afb21b1acd1c
z3b03c94b68c9d36518bcc175ac1cb0e819cf25e4f2ac095e8a1904e27229c96e4a14c99911f448
z8b57e3ae1cb96ea2ffc9b60461264fce9c3167af7c1b2417c2b1b639dfab84630ea9250d287d1a
z1b21da889bed51f3e2ab9194cb9e63acbdcc98c29b9ae4ec5b934de6a82a3258b818c93ee45116
z4a58a9fc698946a25052afd8e031d0e9b5747b8e038c0a9ccc881a79fcf263eb76733e76059413
z520e938e0775a2d73d6e92a423b8dab122463b9f50e6dc4e93a7a16f29f918ff4c277d4c536c06
zadb311d2a942521f9999980e0cb6bd7e3020e09ee8426c032ff40c56929f0dc7c134950ae8a6ad
zd28a00812f859fd054ed810d19a83ee82e106d34206556b88ed2a0891e01a153abb27402c13714
ze5ff6ab9141a760a7ce698439971ab2ba731b0a12f01cc260e33855a4ae44979153b45576d02df
zda57a4be4c3d319cdd2adf6113f5976a0b1af2d4362691fd15b41a1b5857a8c66b22619d3884a1
zf5e12965f422b598870bfeb223d68d32d821b9c10a221313f8c811611c2119f6a13cd5e57af0e5
z972ed857da659c7e1fc141d3db7e96484f9f8c0f71d8afa396737e5bd498513f0f05ba5378f05f
z365339d6cf2bd6447e1503a8999077ea628b507052039a6b903014148736c9654f3a5cce08d89d
z5392e5d37287f0e8d0eb95eac540706434cc41b816d9fb86010c6244a01ccb2bc6ba1029348c29
zf5b0265de879f6e97dd1ab2a88080a82f813f57c781a46b207acfcd8a1b74f1ac7102a60b62217
zec83f20a20fdcf78850ea1bb4111701e62f38f9354e36f8768eba4d919b6793618f1d9f560cf89
ze7f178e013a0b68e4ca9404ac96e396f0c44ba5a853b4296c6f2011ba9e76c0760ca99d80a350b
z6da92021ec3e711fb25c20225efed8e11170891395b81cf276f0d75e6f01fb234f3b895ffe37e8
z94b8db65a25dfea24c78cb4ffdb8803d9ae00aa7c8e79b095fa023d95f794fb8aae54434e2bfe2
z9de70bf5db376d63f44fdfd713d5e1e3313ce78554714ac804dc88f90d444a1b5b694507e42bfb
z63bf974459b18d5f14546dcd8592379595783ccf1e435ca84c4139ed9c03f1fadab364eae1f404
ze38ef836c84bcd9fc6d283197739ea8fe3518a5b923f9f0a5b7ae7b77f07f6ddc7f96e08daf387
z2cd6b46b286693bc20f13bd63172bdbfad850f212a21c9027d9f31c14e9af3d564b8a71d9945ae
zd26d12f9be40ac8eda1d72dbdae9315cfc99712edc2b1cfbc96a6a81a3f3bb675b99f47312f7ae
ze5f63a7d9ef771096c354ed006ca2ef06d316c00d1f62164f8b6050349a310a25aafc894b24fd6
zb5fd0fe0cbf5aa4b3fdb58b744c492e9d24489d45595d82a2c1b37663773cf80e780147c3522c0
z7f01bc075db04dbf48058cb5786dad9695370c2b912f16491f5489a9809fbb7967c9e54da4c566
z35b02e1ba43ca8348e387b2f34b6f43a00b8c0136583aff01c625e5700fe2c02f672065f855043
z5ffa6653fcef631b3d043444806c3169d1fe987dd22c043aba584c15f5cb9d9f93e5fb017fd6d3
z84a65fa59d47752c9d3f0dc00abf76041d407a87ab81a5a3800035b831b2ddecfbe50a2b42ec41
zbb1c062a8c76696e1235c6536327347bfd2bb6f7fcd7877a2796f4cda9b46e8e3782d429251e85
z27ec548b649aaf2b6a14bcfa4a935ef1fdb9144b985d65aaf8252da773172b4ce71077c20aef5d
z923bd3928f96e0d2095cd118b56ba410620997e8519b6b021341da963fca0610006b08f05d56da
z3912a123ae4b6652695c8a78d8e2f114bb9600be25e3706ffa2f038e1db403e89436dacffa58e2
ze216a3657b607f042b7910b4d8a07c6449b2da424803afea63b3e274653a89cce4f01318209117
z95f9994d891a35d485a47c01397e629ccf66caa715637e61e9c0676a7d146a9d3fe30cd26d4d15
z2c37a258821044dd0e1a10a2209920201e2ee89908ae7a637c6036f417d006e9559d388f6331ad
zb3756c9fa71fa048b2529efd462c7b427065ee6cb5f4a21f502b0ff03e0f8d4e50869d9fe15c7c
zcab2669f2ba4fc90df60a215149c1d04330f7ab91186cf445e3801f445c15cc5c8d0ee5fe4ba68
zdf90429b287b4b2b6ac2e46c0289cc5ee4d4e9b4d377bf5f44f4023e2dffc33767741154e8c2fd
z11dbd61ff11f61915078b3ecbd30e914f552ac069900ed16cce2bfa4de83f726e3b6446991656a
zf9c7374b634c16175a7e5f73362d10ed61afb2bbe9de2dcad9a1f017d1820b20c44fe885f8ff0c
zdc9b666bb3a54f03479579106cc31710fb708d93034c68727ebaa75c9400243a7101f2539e4c5d
zad1cd94ee5970081795e0ec7db86dad7fcb1d90ca26a35c634a52dd5be45fe70557fbfbfe5c983
z6b3349220162a7b12af8d755903126aeb393de27cc94ec2e3d4b48c0c273977b7d2cfac217a115
ze752936592d874ba71f68ad0cc9b26d9e65c75fc68654669bf0eca30c5e8c977c473c7953a4468
z192eb46f4d7e111c590b60576aaaa3876a8c1ed757ffe00c0b37ebbe188a5768e261350b5d84bd
z38a0df5741a3b3e9ec32bf1de45897b6509e61048c7f2ec35cf789364d848e9ce9896e196e6cb7
zb28838816f8756de04abb4e7fc2db62aa90df77af496ffe0b04a56297a58a20371bfbf3e1db908
ze5a9b9a03828304d6c69621f9dbd166d62d18f23f9f371c95588ce97528e6d7104b1bc0dc02f5e
z96cad8ec36dfacd29ac23481875fcebe0308ae5c6f3a0d4cc99b691c6ac66a0261c546a01e8647
zd11ec0eab2dc7344af8c5e0d1855b5fdda08b5c8cdbb221824cc075e34d0dae55c0ff5b63509da
z682e9e39382e904431778d35ba2dd82ede21591c3132b06aa22e402511f18c60ab7f6b57205889
z4823e0ac666bbed671aadfc92303f7707d2aeb6f9383acb85a5192d56525f7114f64bcf506c9f2
z8502bb1f10322ff280c240fe5c02a5868bbd6a181365febed954ee9a20324a323104e9b0699e6e
z72048078f420b75768e52b1437007b01db6ec65850c8552a2627ba317db79951a7bd668b04ba09
za32d1e05a6153f0559459d6a97b68234453858d3260786b852d51b10422ba15ea506bdbcdaa901
z59db6158f07987afabc39db7eadf8ad1efb79d7d3c2bdea7a4f528254706884dbad460ece0cc3f
z8ef396c9444320cd208adaa869b135405cba3ae0bcb216ae47aa77b34df70432d1c6f88e8b327a
z90bb7fd4ee4ba592b6d3907a6a8ecf13037b373c5b71a519746fc6eb73e4f86a909ddd93756c8a
zec9227efb2a439d1076102d1d1903ab19733060d092ac7f3ce6f7b52ea37c3d7179b7d7e2ca118
zbfd931813d8391a8da7b72d2e6ed513e24ecccb71b795cbeb1e210624bf71f3581e0e2455d8af9
z4209cb84b54d8027ea7e769dd4113bb0adfbfc73bb2252adb146efcf459a67ced352cd2da0df88
z31fdecac9b85e2c6ebe09232ffd4b087529822fb6fe94905a12c2e4e717e419c4395b1a23cb81c
zfbc9d32ee0a810fcb71e60ac3ac05994efddabe4d64af42c1938d6e965752ac2ae7b3068487075
zacc6ee02f241d026f7c674ab76c9f4e62550524e90349c9b545718b853d28c034b50e101f22c66
zf9952b1eed16969cd48ade3b6a358e41585b77ccfea374ec64ef6e58cf3e3adea74f2cab5190f8
z8425617b41a1924b6a7a7781ac4922b0e4625bd10a937c10f8ab8a9d6f0571d48731ef8a961db4
z395ac17938e2ca188f11fa0089d67b797a297f6fc271f1b397a8a4329d1d1bc31c5c2cbfc913cc
zdacfd586d9ef134964a495558ae5bf5e90d959e91cb867f4a2e25e352ce6376f69ec99caf9597d
z741d09a93c2cf6de2074d40656933d6469ef692e15f3e3a2d4094e8a4e06b9d93d0d9c164a4078
zec05b791cc410d0ab906a197a8601397f1c0b6fe9738318f0e4549895fd2131745f96c95d7a312
z045a85aec8707e978f291a5be2bfd9d6484e9146e92e31b8cb6baea67efe673bfb3ff44b8fc14f
ze9eee79581ea227f574529ab8ba2482c3b9925bcea3a2b16ef5bedbec8afa49bf1ce81dbd7123d
zff8ab027603ecff6cb504b1f49832701d6bc2376e413ebfd3e5fabbadb190e83871d86feee1aef
z02bc3f9c0375a748ac190736e67d53be4819ea59e8d2da32e70b5ccabbb91b071250639503861b
z0ce997b3dfbd4beae040c1e0e3ef6c636a55c37fb42c47beb91ebe8bfe772e6613582f20a69024
ze4a74ed9bc292cb2c8be1cf935a4523de336160fcf4010ba94ad6c93f0c5ed48b4384e7002436d
zce9d64cf14fcfa8cfff6f79c3ec43c39b0878fb3330675661b9d6ecea438219d316a7d334d6b7b
zae27dd619e20fe1c082e1aad870efd25daf84194c36e71fe61d6d5461a0be5b934d0f8891f0604
zf9b2fd93787ae9a662b612557a0b3d9923818801c491b557d0d6e1836b2c07e2a867c9747cb05c
zc5392a770d47053ec6b1643761babe1a2b0e1c5d0a196e891bac7dabf821209730de9eaebb4ac7
z4170cf7db57126f15664b32899fb8aeae8f2d4d8034cefe84383ae639955decd56b8607bc3d12c
z224ca8f405543b7ca3be3a1abbec00b3035aa88fda2723612bfd1987ea862500571d26704cacda
z78a834924d7861a9012c0260d7d510d9dd7b12aabdd58c43f6306bc4b02ea1f60bb34adca38e8d
z13c318f385d2942066e820796360d636a8d2a4fc91d77716de28e0bb882a0e00f04ad19f000af5
z3478bb380bd9d2e31ecaea5ce7964b97d0eb9781e3badab5c03c778eff33b6992420afd9473022
z76887263e3466e42cb32303653fbd94eaf09e0749323ae37067ecd07cec78305670d95ad15529f
zfb791d179a0dbbff72fc245c38b692323021a2cdaac6789cadd885e81e6a3b80e42d12a8be2989
z843e116d94bad606ec42d7f4723489e28977b08675a9bc74166bce1b21821a193e94781d6b9b9c
z60ea0eee2947afbf97a7162ff35903ad465520d0538cec73cd6affba291ce559147030ac47392f
z4e8782d63570364f4d9a5e947d0fbf8dc39d5bae3e27df517d089c5dbd5e7624821727d7295ecd
z0d832978bdab933f475e8ffb8c9f92a17a4d71dec579a16c274597b966fe3484a2cb2e0ca63db4
za555f45cef661234e50b58023fd5cd8ea3d567b9f9cbe3767b740575a4815b2356eb79afb80a4a
z0353a7edf36c28d909fc6f25fdb079ae13a81e6ad30defb9505775952c113d7d35b0e866959843
za206139834c153531d503f63607c5e436e0f860cd4b96d8a7c302b3f475974e4c9c5fa541d0616
z1594ffe7fff51cc4129f4e1b30b15f20eb786a07238206e3ea666b0a0eb1da64032bb586caad4d
zad29ca6d3c4f4e6b42e62ed86f1cd58c6e49b5b925cf125dc79fbd9be6df31f9ac02f918980e3a
z65598e442aea3ecf13fcc4ebe0c93da1ff3aa0ffca1fbec1202b1add00b89ac36a0aebcf17ccc3
zd5c5c73bc8c1950c3eb93ad33b2ee73e4a5d885098543fa1f8f534f6bbce68821dd9dbd5fe1e39
z866bdb3f7b3986dcd22d2898ff3855d27373b92eb69c804f39a7735108d603f60a8d4724f19bd5
z9f6e0ea648f60cf16ed5bd24bc9bd4dec5f8e85ca28d4fbf6592b5acabe30fa0927af2cda9d811
z48861ff74bb6cb5ae74561ad7c30f7aa63d45047703615b0303d4975ec3a17f16bfdc38d0b44e0
z53ef75b0bac20036ff6d8d8e9a1b50e6ecbf2b9940ee37bb80a6615bc012ec37d676a72381e518
zb05a0c4e50ae1136049baf0f76e8a190979e102958684d569bfa9b6da5332e3c9c707829eef546
zfe4f5afbd671a39cef9fa6d580d13d0e38b58b9a31e24a1632d29ba28bdd3ce4af803c8a13af89
z331d680eb2cad8bf24194fd8a4f423096de6ad28d6a6c7252a7e8f939284071d498e5135196dfb
ze15ae2fbb50e0fb934ad1257430ea43e66c655d668377b84f16ad8dfae9404a99cb807d47de83f
z320e909b2c68067497e8b04d38b384a8446cab25e9049132a8ed0eaddcf427bc677bdb53dbf2c8
zcd4ed20693cc9f8c14a81f5b7ebc5a0b4313fb7596f7700c75f45d18abb6f946a7304acf4c9bef
z1116bd0f67bdba0e62adc04d1f9fc9e026e93b778d000fbbb517c996f9bfca6f50c6c68328a359
zbecfb6deb2b2b5255e72e6394dd10a8564550094fb9da8ba27996e8cebd8b85e40e0c1a45f287e
z1aca04973e361aabefded05d694550708c64fc4c439056aff8931098c7cb153e295a46e11b31d8
z2d3e9d949d01e6dea9dc81d7968734b36bc019cda761c4d58c0b12181102c5af13193fc7050ef5
z3bbd7b76caadc77dc54c644583219d8bee7a694d46b9c620f088a4832c477b891748412691eaaa
z22996cf8c492f88975900c9fb704889dad252fc1f50ca363262bc244b67b9d5a98f9e25ba34145
z06ef811bc567b8e5fdc88fac8028ac6f9cf0672b7d3eabc2994b1afcc12d371abcd6e5ed47d630
z5b1f7d57c2daf3537dbba6ae49e71c569e18a1db7903173ffcca13c40ed4b96ac4211f76e5024f
z0d055fea0fb4e2faf1b7a054cc02cf7f0f17ebf8da2fab6bdc617b50250cbe1cac5f3a53cfa42f
zd0dbf4de72b7ad8288e3385a098f35a7cb0720d9bf2d4ce955eae7f98cb13498f4fb12ff034ba7
zc692b70b9f7f6864d430e16ce98e8c0c4875a8c2cdac0c5ccd8bddbab86238b125f3211bc79042
z0acdd5ee309ce58a7d33c84825f1c71790057a81bd7f043db21afc25cd505d198fe3b19778eff6
z44db96a2197b8f46940eba533bed1414cef5b81e7c5c0c32271823e3eaf2fe75bddb1f6ddcb7df
z15f4ae8674ed06a8260f8514a1c6d248a4d85aa7b98e7a5901b53444028c5e16722c9b04b45d6a
z12ba1c8dfbed64797c3fcdec72e6d697eaf790a840003f51b71ba8c2cd1accc2769df52fd8d396
z902f5b2f8a1af1138fab44ad1f33b484b7bba0f0d915365469e9bf90c376e2b67fa05732f02816
z50ab8e68f6f3a423f1105b266cc24320d0ea8bf8b82c50ae3f0fca7b1fc132a0ff1abf2a1a2f43
ze883631cfa8f42e4df44e896e1e865d5fd44cc913b687efe725d66f7b4ad1ebb6d2a8279b20b04
z9168014878b322680f014d3a47b0bf56fc82462ec6529d62410474252b4c19f8d023d3c4b2683d
z55b81ae7f785c7d0084deb3566742661e70ad98b0297fb7bca709beedbe6441edebf34cbeb4fce
ze54876da18ceca726815c704793ec27c33cd09fcd732e436c62e6fdcd6db8b1060f23d3c93a639
z21469bc0bb580ee8aee8b5a24383d8cc81d5813c2996c11208ceb84ce7a301976388d7a11f46bb
z51080ce424321a037dbc59736ddacf23c6f55e50aed243cba291d8d60e24c155bfd5574c4ea447
zf1711556555007149859a0987503da7c34700096d1d5fb6ddd9beffc60396bcfad77d9add85cef
z17fbc4d869dad93b4c26f06eebb0546b043909416d0329cad1fbaac2b1886d1013eb7034da625f
zcd9cf0a2b4103a6ec236b0ebff5c2b6f3ef1f8471a45a1d16b9b97c575ada72ab90e2f4a72126e
z50ddea1d826eca230f60a3a029b487a987829871880fb2dc5d5a5d5789eccb537ebd6e65f2e7bc
z5dd154fd24c5e8457ee24ac7c4b956876bada6fba4f6ee33e3e52f6c1b1a6583783be37719156b
zccad418406dd9afcacc36a5ad3b2c990fd70218a71d5c733cdce9306b614e46390d623cec1d3aa
z1dab9189eae0dee4294a33ebfdcaa6b0efe630d375e34d71330fd0d36b76e1ef91a32d9933e810
z06fa5c900da14fbc5281054681faa3993e7402a17da74898f8267b736e64f52a4739464ed30e75
z87737a3c94140e10792e1712077aa3f1249f0c32e69731aa98251e3081fba9e4bc90e5436e21e1
z61cd928c1d6f3066d5bfb8bc79a246e63a61896381806b01aa959981e51456c1e5fa98df63d5ec
z1fd002664005176a4f3dc96a38470dddee44281d63076dc911bbcf1e818388160b2b09a90d48ba
za2e6eeb8d247da0b4d5ab35ce34a5cc72c07ca920337b938cb0a7da42bf93b212a4e1986ac9698
z340dda588427f3f674c561cb56ffa033153e2239638770d65832515424dad0d92c28c32759b33f
z87df3b7079305e1da5c58b9af2010cbafc007c862f7a671d51f793b9f9dfbf7a9ba52ad81a4c8f
za42b48da4c6eb939ba9ff6019e91496adad45a82e623fd754bc455bb0ba6bfbfec4dca5f36370e
za400fbd2cb58fa81a4e7de9b0b9b50b12ea92a67e2f37dddc1ed19ce393452232714a8dccfe09e
z571391378c61c1af12e23d87300032c4924ead456a09c0afba3a6fd6798570a112ac29bdf7acb6
z37b83c64a1d0dae97f58480c8c8fc71f9e8672fb8977a252fa3b10013d67fb94be48d26bee60be
z76b6ce68c378bf00e9f7be80ff213d1eafcb832b9871c4881ac1609d64a57d968ffee51cdd8d52
z4da7c7bb328bc300c4cf6bac64462964f3c660f763e346856fdeb4eee5cf1287d8def50b35df67
z978b9e4b43da49ba4292d2d83db278a229d1dedfeaa106dec53a56a9a257e492a357a9467c8609
z833f4e4b494f9daf1667da8898a20a2497ab946850f9ae7ac4e5f637d0f3b14e5ff1739d2e76bc
za05de8830922b9f9d5dccb0b1fae56cde4b0ab36c388ec6ceb5f35d53b9f381f1209ec3472d2b7
ze1ed42dd40cd4acd082d6552d08808e392febc422acd8a18a28bd2735436cc633fa73ce91faaed
zc710172452b0cf211294d3b519e75690ee77931a0749892a5f812d8f834822ae2779aa167df889
zb005c0b031faa4ac960401d46e7816c5168620eee60d3232082c4ff9039f9be44acd59dcafd2a8
z2303738639a353d848be66200be397d95d2a53c09943f5ecd34336a51736ab6b5ef17b9ee93c44
z4efd4af44e31da4a175a47e2c307e045735687860ded81d140f6c88adfbf56a2e1852df11314e3
z66cdb1f4fbd16c1454717b3dd2aa162efdf91cfdccb7f46582a9a904d61d79b348f89c4f0da94d
z4c64cf63935eaedb2457bb143f0d69321da6c8151549b29a37b35ad8fd735d38cd66ee0bdcbc9e
z10272bb302d1fc2d9bcbd0d4829bdcdb65d860c12540852c1f52e55b920a5ca10b016370edb8dc
z22cd9c9f830e17e1e8798a3252bb6f28c75c54f63e9883e48a511e21366a4a33cf2e50ca248265
zec3e53a7ba5b5c38158f93080dfa2b8321672305f67f73833a8454698c30d95f321738e46120a4
zb74ff07053c9aa90d8d7d37c159ad06f36cf7dc6c1bde457a954009ce1af5513a14e3c2213dfaf
z599b2c6a8f12be4d748c08fca2cac02ae0690ad9f00de36a13e43b355712c3f91856844a6cc26a
z1010f615989485f5ad836b7735e2b4b7d5a55c0265423ed80b83bfeb0a3a1c968568299d5ed2aa
z88e5a5e34ccefccd7c066b8f26f2087ced612fb5bbea14ff9c82e515e2b0ba59add037898aefbf
zd9a4668a940e4afef463df67ac3bdbf75023ed33ed0d29795c271da5d723f39f4abc25fbcce098
z12fa3bd01c78132ad85521acfc0b77f0755607b1c4c18bfb1678f6e5870e773be9ac8c2256d51a
z9085d1d9cd18eaa9f1b64fd78c7fe34e1e99c0e964aa1682b8eef6c08150976ff1fe0657d48261
z02d62462f7e6872b2d25626356d4b3b20e38ce6f261ae517f732fc97d88f8d618449255d66b697
zc0ecaf3bc61041123a8f5c79fb54c1209a2b4e47adc8af8109ca6f9f5bcb526224682863ea580f
zb9b40aa695327e49c9af96931c753a7115ca8b6c0c3ee56b293cc6a407bd0f31457408ae2ceece
zdfffc902216e7c5f126a33e03f4c94d6666379488de716fed018bbee6d604922e20c9853276e82
zc0b25e8bfee2bcf28587c7018aa8f1d9cd901952f92f16b281ca0d6b7a907bfa906dbd250e3848
zf5d12211e9be407f281912755e3e31ea710576da34dc8e60f3bf8569ec3fc34544b27d395c5760
z22f3e1c8b694fcd89590853b3d8818c48c7e0beb9e0fe2f644cbc1d6b58f6bad314399bded4776
ze9fb96524ef7da46f10106593f3913acff48eea4f859fae8f7ad18cb08aa4fcfae80e63f566c43
ze4238428ffabcc09f4331333dc5afd201dde9f3d2c773cf2b1be901834ab94ce1e96e04bf0eb04
zac2b900644861de5eecafb653507a497ddab0ab44b5c5b930e33a5847cc30c56bf839ae6296c8d
zb7eb99a0456ba8dbb7ed40723487b16207368cb58ce5c8d74212ddd71dc8b7eacb617c71702755
zeb64d070f5acb7719fb229d685b09c9b04affd31adf0ea9645409375b127220fb3d3a485328583
ze3f510e96c7f3fd8c6b5cc9315e4e537480fb1318c3e2f32371bd6530058c7a3b30a1eb94b2fe6
z6d82e89ba4ab1c1c2a25ad27a2d17fe7e728c1269118aa17db5c88d89375ae9a3a56a8e2e311af
zbd3fac60ad9572e9956263ef4a8c144e30f404f3359fa33ceb92f0d471b33449835c08a59686da
z58bc7ec87bb2fac87e8106f6833206bebba9e95b8b80b5eebd148dcd0833fd5dd0a17a712b7e10
zd4afc839a69ddc3581f048cc592ccdac12ff5f4b469645eb0fde0a1d5862f4407759f860bc3f51
z51d534a9ce17ccc8765bab79877d4f81136e59967044b88ab8535ca70ce701c6953b87cc002b19
zde92992c4c98faf7131c26821eca7abaa5e8581e739ec017ca7fc716c67b56449b0c82f4736b8b
z34001e9bd7864127d1976c444d5b5666bef66ba1753f54fb4ae3661030a79e023b2ad2bd22ea07
z195804d804fa8a87d4bcd6d029079c5b09ca68be10c85178d183d08753ca06c277404edc1496f4
zedf2d1b0f14355774b707880ca9a6947fd885d0dfda5a2c494ed9513bdb4812f8975cd4a381846
z41662eee00f63a5d8322bea6e2daae52188c709b7b73c7ab6fe1b62e982689d648b521f7451a04
z3ce79981c38ed91896b1e4144ec748943f2eff8c20184a6db84585de2bbfe0744f8cb5cde441e8
z2ce2ef30d7e0bf2c4353bb4a8eadedcde1996271bea11de5213fe33eb4ffb58fc62d3d346e2fa5
z79f8bbea045149c326e5781772d70ef889128986f49017921273f8a11caedd40ad2a02e39f2889
za31fa62d42bbdba8231dd7cb90d96c9fe26c88ed7f5c9788c31cb06d30a062ceee033a9c2133f7
zc56c33db62485594806f7a897ceac4033421f6a7fbad1392e309c9a07d5b4bb13ae5bfbf0ec42f
z77d2e26fabce25c4021a538611378a124d3d45896b1099e41fb279eed6040c343389346b57f917
zff079dae9e965e08dbf808dfa3a066985e616453cc28371f24dc6f6532e16368618207838dd2c9
zd2fd1e58adb14bf26997db5501d4f6b02eaee5f060781cd7257cd3fddf9e6273bd2459ac0e92e1
z9e4b147384e58517b373b5e084aef58f187da67c2ff144fa87c4fdacd8fab4755e14a3371a36b6
zcf2d74258280b9e55cfee026412eaac623a414ef275698f6b506577f7daa37607d9ce4e7ae9b6b
zaece4f07fd8009bbd363c8a6bfe05f349d103e26456a7099c3352d82a59573fcd8225d9d9aa783
ze4562598101dea75c0374ec72de8a03aa69970dacd5166b2063531ed7db9fd676dbb9c1381c907
zeee66d6445c8f288f786a19900072633194eb0acb15b5200a370afd4be8ee858838cac50efb7cf
zdc5c09d4306fed43fd8d27924d6e85003b26d2b44f1f48f56c2d8ba01096f930b51f4910f82ca8
z81422850501f10642c3de8485ced17d1d3c1c5ae031f52edbec276e8cdb66ad3ec10fa390229d1
z7a6e9002f27f712be237c61a4fb79007f4c84d897532d737ca9753333d1a70ad95df888aeed4f8
ze410114e96b190ee134c9528575515441de4899f2b03dbf9d02b98713256c78ae77edfac352a4f
zf12e9a25e759c4832bc4d330679a88c86f8ab352b8d585bbe44a7d696f9f599543a3209643c8ee
z76e9840063617b758dcb3b4eeb76ccb5d948a173491a62dd16af8fbbec835bf0e0af76b469988a
zd2a627083e605f92e69c9c318c74f9ffbf500782962652d2652ca56d33ef1c367d2e98ce3cf39b
z93ea74d7ae242c61bb53f2f8046fe2aeec823d9778c23b3c47a40d7b0bc802648a662af4031046
z9ef08fe69bd754cad9f950968645e51ebb723fb04652e8f4daf6a969c818878273a6606bba9241
za165a7aebdc24c9169526527570452cdd43d57287b3c02ea679b7a48745027865a1fedeecedaf6
zfd54b273c4e2e8ceefec48538ad55eedbb6de2f6416954af789019aead07ae9a940655f7cf8193
z738f11bec7ba32c653b7382027e1266063249a545508898900d2bcdb6af97e01cf21756e2abdb6
z3a36a0c75296f2ed5ddbd24a5ba8b83ecae6d985910e53431c4722f275fe0f68d2d2acf194b2ec
z9e08ce9501c91092374f379a70cd4070943bf80bef26a2a02e95a5848e7b167817343c67d713b5
z071ae1c3d1f7e72ffc4e71a444264c6d02ddcde42b8ad0c0dc473c9f9f1a056ea7b86ac885a48d
z5b27e3640c857c136c66f77d5ab3d3aea2a058f8c2d245ba8ef31ca80f2e627e4bf7b2618c7f66
ze297b7bb9d0f56d6d0ab427df47f08a44678d254177d6280dde7aefbca7fcffbb79e582d6e2f5f
z1dfd8bdb2b8c0a0693117da8beab6efa8ef11eb64cda94a08815d890416e52b8c77d7c181e7c11
z8b88120659baadaf488ba47cc154925bfa0a1c7757aa181fd8b1d3df72e35306c24615ca80d482
z82888e945d63e0cf20706467d5cb71c64f54ac28959659f2723931d532728ad8a5ab016b510ec6
za6529232f505fc03a9791316ded347172872b771e8e289bfb803445182c5416c04dde7a58b65df
z5029cce806eae1a7a336829dca6a9918c696aeac002bfa2c5b79d983f0086f64e1f2c488a462cf
z384187dbc26633e214d515716712c2ae958b5624744f8ea5c0d4deb064794305be5fc2d0af82e7
z55c1fd7554f6dc186aa8d1abc0b77806c15289b17d1c45e8c71a980e10541467848a684a308439
z46f35bdb9d2a0541192317e3fb697b3eb0c051792b63a1e7338a9942c02003208da0f69a89efee
z890417fb472b99268a0304dc7a81fd21f649710b0c0ee1328cb34b1e52ffa74c64f339436c7e8e
z2f035f5d74160cc362ff4d999f97418b0cea0212d942436b5f1f3e96a06d4156491c7fad6ec779
zcfadf0d3b23faca02a68b94e89a2d5f2f2c3eabb35dee51f761f65299b5d2abb47ebd1cdcf1fae
z57bf92f1b539539532eccf1cd5a49c0b8f54bdc5ccef96ce539c6838d000e319cebae9c9feb9cd
z01ee70748bce4791407332532fb26b60f9ddc2fe10d65642e92b343392b6cc29653b1d836605a8
z92b0941a274756e018fc64dca665e846773744a089f575c35f4562dff6d48ea77a716e8077c2e3
z25e05a4888de70da9921ffddb0c862046b5e9f4f33fa15d859aa36cd13ae4988c481276c5e11b9
z91db56f9c2c495c827f85dcd7d5e2684d66780b40956a737650f53242c29aa606f350ac284d948
z49427d912bc9b21dd72a9820c657e1006f640d8e74aa314bf9a5aeb85c30b3bba158d4c7d58e7c
zb8e837ee9b7e4196c978961b44d6b8b7b14d340ea2eb2ad9a0014551a32c9256485e2f80db70ea
z60d2b134ce06b820f41a71ec8a57b0ba86117d7ab59774017929298306b7328f4b6237da8ebcc6
z8c6856b299d9f209275405d866630cbec91e27a6d0df9de6cb097caa07daef1deba081b6ae32ca
ze9c703a129278e64aefcab04872b7d235e03829313f46952fce60d7910c0b41038531097850cef
z11cc90300c40b41736102cd5918d565d1057bd8c62f91746cc635440bf89e984ceda8eae73c95b
z3ca6c09cbc4943950accef47bc7a8ab7364aa7e82141477571a70d77f4bb4d175e65c13692198b
z6b926ae46882de8290ad0f68326f19220ad38afcaf2f6ece0b92a0fde80e5d79c6393688bf31a4
z3e87361624f4dcb4528c9680f75499dcfa36a89b4c001493fabccf7302744da26b8b166f05a10b
zd1997729d4d262b258c28f9be9acd3d0a44212a8f5559f4816c200dd081b039fb92b91443fd54d
zd269589273318112541f6c630f0c91941529128b1e44cc7a4bc1341eef9d3f1809e3859e5aa685
zd3b123eacea8bcd1ec58913276b3390b864ed21dc5214445031689b46a969c56113e32b077791f
z49c5e17ec4f16b91f3092bf0387a94729438505c971ed074bcd7f0bdb635d8640e03cd682d4927
z888783d2bc3d3f1408c886c5b737805e8a934ec60fb91c2d9a65399f09cd3a3c39862b9373b428
zc18aff3c293a32ab1cd7bb0ad2d4cd141702d564f5569d9126c00e023f026481ffadeb93d780f3
z10acc5a9fc571ac7cd63944b31b287b9beb1ef00f20771ebb33a04ef09cf960e40dc5b08f10c53
z608f8cae852d5194513e0d930f97e1d640a61141ea601938ce402a587dc3b8c9d8c54083a55ceb
z85897633ac0d68bbf8c72c0a99aa3700bbc3c366a9c527a7b9255546924730a8b3c967dc0d8f69
ze6e3ca05aea79ca80e68b27238010680b591789033087a17d4ab1622773ab89e3d6d0d4823cd33
z82da1ba9a95e82cd6ae2d43832d4e006ff5da923b0ca60721819f9b82a175e64e0ac809b70c217
zb465413214a249884868f839c7115ea47cdcd408d28fd57807d6cf1beddf3d8d839fd219558f11
z40d7926283409ab23d5c3d83a386d7aad695acd8198bdfa8607f6f710c376081416937296c8453
z17aba8e376093e78734f8a2576bd0203d21ec11a925040427260bbb5f20ba0459e45848294f868
zcfc074ca2edb8baa9a654074645478d50cbd4e406de4aac1dc469b36a698b602c23e496375c4ed
z9caa07bebca331b2f948b2ecea6126d3e7e8b2a1a43107bef5033066bda7bf6ff6e4ec2e6b1c4f
z4cc71d3a248f82bfe5faab715e3552adf56f32bfa2d8283600a29415772172339ffc23ed50854f
z6d67d62b75fee6cbddbe4a4e7dc25ccbfcc8eb3740b0b551b40c7c9cd5035578021cea1f1147a3
z9afa134a9a1071d5956174eb4183fd55a77d80e31309e0c9da78e2ae3917aaefe4c9ab19f8f0af
zec47f4b266e55e4ce42877a56ffa6ad46597ddc578894a6ef2ebe28c685d466d941e2ceb0d9745
zde72aeac14990ca9ba46a9a1212c1b5121f6ebf0d28cb35a96482e118afd9eefa1e0bf2b84fbb5
zda13f4b202554579246e322b0c5c5f2d51d16ffe528d769188a2b236fb770ccd17181c6b927ea3
zc6c8c98cde1e9af4101b24426451d74ad8636d1fe574a742d7a1001cba491f3a9ddc316b3f7a5c
z89630a86f6b7a42e0f1995a2e7c46a485ab4a6be16b6b343126c577ff9c94d58845bcdadc50a54
zedd20120c50aa62db23e810a8f2af997c30568c413df8454f23de5c842552cb96469b3ce689482
zacf7677c5645cd22c731d31615a221005165127446d8d224ddcb5e2f391b4320ed6d7cb25609f1
z927917bf6583fe7107a3ee46423c8e71712fd8d0b562630fc0d0cbff909c72a3be012e50377cbe
z0a454fc1d853955181d07ebaca72c4ed09a8b549abb769c159614706f70876a0700b2dd4be574d
z4db3e39d8cafe2107f01836826cab9fb0cdbf62d663358e839392fe814b86317b72c2788749860
zd016db5ec33e2312df534e75ddb662f0acd953b8bb6579c95db011fa367c0da26442fa53ce028f
zc1b39b4e64665ef048c0d2045099c8156b8d78efc586dd4dbf50d4b8fa3d8453b8c135b26209c8
zcdf5289aabf0c90be05b0d1632fb2f5e86e0c705b9b0a9b06adafe8d263c2a7b6750efd97c12d4
z75448b950c246356b53e2574dde14a91bf5cda5a0998cbacb348a97e41e6b43f291ff9701d7540
z10fd4835264f72c3ae52041a8f9fa77b2456fc3e6cb2a81e517dae6c4f4552bbf4b712e9692e7f
z56fc640aceeaa41eed9dd8eaf8dbe70a6bfa941d77b611baef47a707fbe2dc12522a14e414df1e
z69beb0546ed979d27013fdcc92713e3edb29b5f6eab1d6429145cdb251bbef53f5bb184417dd02
zbd5985deff43b798b9ca9bad3a2fcffab07185447fe8882f74ed7fb086959a3357463a1e21fd1b
zddfd9c66b45dba3648f8d49ef43ce419076be1ab0b8e5b8aca4df446790387475cfba5a10e0172
zba733fdcf247cadbb906433a4c1faa7e68bce3f14160dbccd7cc1db05bdcd00d688ffdcdea9624
zdef78bb17b15993a70bb915386ade5de6ff2daae74a80d89100186381ba9dd7e3a5aac06e60dc6
z9fb445b91da4a32848125c627b6f7ddd47bebfba3f9629ca1b0b56cb8da434e4c851edafe46e40
zc91d67fb0396e36280925e66f2ca36c6ed713305d8580bd9303be8a02afe3ff0c91ea0a3155cb3
z4393f252d6fe07d026d86f68cec9b32b8a90226c5ea2c99620c4695b3e3550349ff73728714e75
zed2c4cf3b7183927167c94f47a8b58062f9aac7fb821e7efb0df13a47aa94a33d4bc952c3e3d58
zab81572733bc7cc9ea40c481dafe74087178789b52c31929dba1456f2b579996cd0c3dae43e911
zb55aa121b27cbb8458008a6cfa881eba8e50b060fd74b60923e8953e6a99c49ab4c89246756063
zed466a9eb7980bc938c9d7a5216b37faf45f371390d3b98186865ba3a7871cda119e575ed3e9db
z635cb1e4fe86b3e170edb511e812381c204d91e231ecba6a5d09a804476ec412cfe5c067d3ff0c
z16bed20c0061e5a98d7d673993f2612c926c2a9cfbdd2850c4a3d21623a35351be066b76fb3fd0
zde00b51a821df100ab00e8ee69014c7363b939618bc45a458ec3352aad24c522316fcf772a6f2b
z3dd106fd19794e8d286e6dbdbbddcdb1f5e2b50a76831917a44ea71d537da153b87009f6a6027b
z72527ad8f477884057d8b4d1bcaebeca0dd7d9ef31139cdce215824b405eb93f94d3bcaeeb62a1
z8a78defc9bbf681b77be41023e3216818c3c8d32098099164c5e8dbda6c8167363f1ce5a314b1c
z92ec9c8c3c85a7c1dd749f44904afd42f41ea72b81bf9277ae1a91695d3dcee79ee425b910ff42
za955bd7c35b24379c8bd116cbc93c526fb46cdeca0949f5479ccb98c212a077a34e89bd06c85a3
z248ee2d802a81e72969bbf456e18dd83987f20459b6e5e96c6b92664575203a719789ecf90bfc3
zb45d381191738ee36fdab33c0c3615a4f2ae18e3fdbd7bd486135dfa68b58ab12322bee04f47dd
z82ab238dd5a0f815ca77251b9f2b3155926ae3727c1b8e6ca26218fa9a03983b9d70683c914640
z26d12ba7e5f9c6a230ccbd518aa47c7d4279ad5bee107ecd7911429e7657c2acc55204118f14d3
z740767af623773dc2915ed030233aadb488f23582de1cd68234ada68685189b6ebc8d6f697a837
zd514447918f26882e5190eda8234b9ec8ee97b5fe1a08fcc10f42d9bb386e7c1dff0ed24345a60
z5cfa1b786d48f82b75864702026b06b0f5911780bcdaf37496841c3ded7582921749c280cfc6b8
zf7a7d219f4a8af574fde81f29253b0faf5ae3d35b4522de919e8e60b1c4dd7a71eba06140ae9e4
z3bde355ed4345c4ff431e58b94085e57344d8f89094d1e3a943e9f81453fc64952e6c6683f84aa
z05090d6fff87eb4ca8142d7b93439c91c098202320f39d803b0c0adf5eb62d357b232819f4ca26
zaeaccc1ccfbea2881976405ebf111199c6a0ea43f2bb02b2e68ff9d5fa264fceb10e9649cb22cb
z0dd4bfc640f29ccb509ddec3540f56979ab9960c32dd2a5b9077d728358a2afdccd6383f31da54
z850decad7a50d4e5021547b18988cddabc78d816d31e12f6d665b13e2ad619ee3b3dab2c979439
z4adac7d973d6df9d741fc6a931ab81545a2ed27154b8b672bc80c6e2918e1b52f82bf8a8bff69c
zcb50567d56f2ba4a90b752495196276c92441fd3948f4200c721b73407867bff0de307f04fc491
zfd637647caae48bcab9131240f29f84bd0cc5f36725abfcde7c88f0f95376bebb1e61e4100988d
ze2ce13e335dec0149f9247b7a41a63f41bc653c813bb04f144573187ab729ef48ceef6f87596e9
z1b5935580627a4d03ecb8f056c455fdc48d3b0199f14093f4114ff47e755475275fff21a6b16de
z42da2cec3e4d508379192e80e8a6420697095ea9a646100b5346124fd2c46bf2f91c88f0b51c09
z5e266e25b8531f250e889a737a5f3515d36720dd1642cd91fcfa0ebe7ef92e2f59c4e8845ca75f
z8de9194a42fcc812c2c278fd4912625db3a72fc00c3a8ac2e76973465230ab30d96e145d749f5d
z4a7dd40866f768d00ce678e8b97b077973f485752d94ddddcf3c15d7d25f86890763bbb8398c5e
z1e9a3162eefcbfb48ead946ba17e5c569510d8809b4ac45cbd3121d630640d6ff158b8c3cf268e
zef443aef194debe86c79ec5e3ae595be57f30d5a07bbc21336e76236c8f7acb5afbfa5b418c1a0
z99a036c6d1efa345b827e4db60fdc844a3f9bc0fdaedd084c1742a5bf2ac3332f5f0fa78823e25
ze9e34c7dcf93c2c48f6cb875c36299c2250b89f22f879efac804138df77824b70b326e4943fa84
zccc93d9652fe07b9eebe9f9561b4a5e508f4077acc23479b629e83d862e3248bffd91878fdf00e
z75c8ff6ab48a521973bee20bdc35e751aae2deeadd0749871ca17023ae14cd8a417c5ce40c704b
z9eb532a46712b336d248f24234959293cbcaa0c978ba7218a73f3b2930f019cc160e82a0550855
zfaa901b3689224ac4a99f9cdf43e5261276157958dc70a841c33c36ed5b9aad47acf29fe217a5a
z06b99a59933069eea6b60894e39a25d11f546ae8ceca1ca3a794350cd1e2fb8871530c6880339b
z834c11e819e507f0c360a40d4d3ddb4b1a9f45fe894fc58d25f4b4499849cd4fc1138e5aec33d7
z5fd3b30a708544756b51dd181bada96fcc8e4a88f322af0bb8f1530034ebab8d13197ae23484cf
z9837d2a7fc78a624de22e32647553cbbdae11d0abdd10c0421393ceface18a1d9ecec385915559
zc6d1925e1809ea891190a1dcf496013c46f1f0cda453f5a678fd80b49d8a3062ccb4b584bfc86d
z8305e33433016bc82e53a6ca60dcb7e54b930d6441e0762af9bef18598107df4b88a6d6e4e1254
z835f2b39d8258abc259178bcf888c484f16b5368c81f89e60179d7497aa24bd457080147171846
z5739b0603ae94609c69cfb73a2d7b29045cea1360678dceacd1d2b2af4e3f1953c6a2b8c7e73f6
z3e83c4b6286568d4645e63c03d0b19471382ffda27173346c424cdbe277eac098fe388cd807874
zdb37d116d489cacd6ea4eafa1723ba682e5c021745c43bd31039452c6118634a80e451705252ec
zb9bf327dc0c1aea00a71f5160d5651251c64a7af3f79a98621db57acafe0f52d827d029ce910f8
z878734c901d105931d1c8a2a20efab4b52f109b06779324a20abfa313ed6d0dbaeacb956516eae
zff99405d9fb68d8cfcc8e7fae0d5bdaadfefd1d1f5b01eae5b940b02a819c2d20b006d86bdb2ab
z9b6a96cf8d1adf92c8596d8dcdc36966e0e5258b8e7955334a101c0d199e521ae4f90db3eb118d
z9bffb3ba47ef592e4126675a596d771cc9215b4dbe8f171e30b528d16f1aed0743496d9f9ea6ca
zc0dec5c2aca849ea7b99a67899549ce0ecff9e453cbb4a0871c568a5b0b2e92f07d724b285f13d
z4ce37ed4f13d64d2b2dec36357d230fcfcf8a99c52ed3458d21852b0a93794e7a3c800879874bc
z114bce40851bfd439585f3d46ee06903bb9bef98528bfa2dc8a1126ac7d401775498ae0e097496
zdc8eff4c54c1aea10ebd14840c6e2d0a8c2eca8a7fbc8cf96827cd6d8578db85571469ffd3814e
ze9a3e010ec0919ba0caa0f1a1314b5d34ee7afdd6f59d13f9553c9bcb63297905fdd2ab142b130
z25b5c42c3eed3e551861d94b250d0509e1000140eedd1ec6e623659115633532d9a0f780adacc3
zfc3bd232e4c9161cedc9b416e931c72efc030370826e1f72f0f729ddae09d6677797f71784fca2
z485afe67c32658c9c525a282ce9363c0a4900722ed83c25dee76bc0599fc8562a268e05e5aebd3
zbb2ff360ab6c271bfd76fae49b3ecc961acee3f111f4a5bdb9ec1404ad21bf3c39afa3edba5774
z0bdd4c5e74881613345026394157c6651b9c21dfa833d4a48aa6953e732590a5ce469907e9a78d
zaf249c37b0a2d0e977f4d786ecb7d0fdca9ea964289363a02fceadc3d27f29d27e2f78cb2e467b
z828251974000ddc3c449caa11a73d356e6fa14ce823b25b9acaf9207af2bdca42d305e6185e222
z93d04a4a4a6854c035c5b97b56c8f5cf0adaae2ec6bbf00b7b1f06917c3f6278e98812789dd95d
z5cc7bf297493c0c6333d8774fec24a7ee014c0f1c154a6261514f863ba03dc15cf2880117fc5aa
z9eae276de4a036a38ac3d57d98efc8bd79182d9d5073ff64c8cd393f5a2eba02483a7ca8eb1553
zda706f997bdb4453c55e298b8efaf1e4da238cf3ae8dc7f17dd817f367997a5340b241c7064f27
ze73ee0041d89ba736ba72e36748f5d7aecf7016b11be288a4d507507b662d8aaf28c5c73288aaa
z5e4d87423a83851e0118d12210664dc5c78cd65f1e1c8ecbf37926ff3aeb93768b870a7fa56682
zeec395d2a62cd6ae255e21507cbb29c57e80a0e7b31b254442a810ac1347270f0a264bc5b33be9
zcd4719b32e16a9f5dda11a815b273fb7e74d28a08fb6784509ca3fb686f339c46c5a08ed032655
z9bddc70deb6cbdf3a248a115a1821315e03a4474b0eae4932438f622d984e894f61b809ff27790
za5d9fa8312b9c0d82e5d4257fa3cd505d7faf275bf05205ddd4de2ec24c9183ae3ae8826197572
z04a0d2c7a3d54849e302dc415844d8cae15755ca203e2f414a5896f31706cf564c37ebe78b67a8
z45f5ca2b4c00dcb6024e5197b3cb79728760fb2546ca466d7903e40db9724ab7ffe94193d1460d
z846dcd8d2214d15623f4848c5390ec2a32876858810772bd8a4139d41fff6f2080a5cfb1acf734
zbcd6eaa91924bfbbb1cc203fc4b6b4a31420e6b1042b02179233d2abed487e75a0df0bfe3d203a
zc73a8ba436cb8fe4f31ea822f22f665b69efbf9ef08ee295714b0a262a9010b1472af4a53a5efc
z5db099bd93fcac6c32896b5c857795ee97d487e6051e35a9850b7c528eced447eb81f9ae198b0d
zd654e62536af7fbe708136c7c5656f573867b2760ee0cd6646e077f1050e84715d90f47c8113b1
zfb87647bb17471f6530cbc8f1af9e316f0ea7d24db6216f6d590c53740d428ebe81628c3402496
zb36ca25e89a237edb5bc96ff58c4f9ea5e3f87e9b81ddc9c84c4a0186d6a03fa390970be0ae296
z743bb3b51108002c0a26dce1138d66131b35fc1fe1e06709253df671f9150c21efe6715f17b7af
zce634ec1217a11139094177f3e833df0ef349b3e3d0f43a10a9c6600d2aa91524450397c061a62
ze4158f7253c65c98f06a55097cc33366a67a3dbe696c50bd26796cb824266407cf69fcc40bd57a
z8cef0b2b8fed99f072fdb0cd149497f3f0d293d82685c93c073106c14c49e93e49a64a9a308277
z074695b7877abf0c1acddd0bfccae4dbc598f5c19905c57dcb732e0f57d472727af447b7d90e24
z965ddc16cb1cf4ba8f2cf9fa69b0eadd00d9022d64faff0230c3de33cfb8edaacab5bc3477a4d6
z9dacb9262ee6552c64a85a2191e087b9704039149efb5755827611c7737fc3b419474514a8eeba
z68ec1df4c84c0cc2ce3e632300caa2e52e3797c2b75df8db1a1be6033a9863f2490897baab6f70
z142048d18ca6b77dc84dbbe9d01dbb11697d430bf32ad2da7a4c63bbe3082df76564cb9acf09ce
z6acb72468f68b3f05f4de9e876da9a75684a59fa29763606865e802b36a80966f7bf8fa00cccdd
za197b614d0ce6b4626a228bb68722fa509d76c2535bc7f3226ddeae91325b04d0b6523056010d0
z0d8128c4cdc38ddd54276b69632e4ed9ff71ae4ee507fa9993bb475151fbca1b03416349d8b8ba
z8868078d44a826c5b5296865ff74f76cdb8be64a0a59ea6f0ff63e7129e44ddb9930d52ef61c9f
zbacf4730305aec5b0f382bf86404245095aec6b97beca20310a524a1bc1ae25ac244745e5e9956
z81946aec58bf0975504f8e86e34d18084d60a3f710d6126c1787cc4e66ad99cfdaf54753530dda
z8f3f0e6e053715b618e83e499d8a0b74116ff0e40f1f741eec210c3bd54e557dd065a47dea5f6b
z89a20d82c0c986d63f1edaf0702c7e819e588edfddcdf6a469c1524c75c2389042295b5138fc1d
z8f0efaa5c3d5f03efc37f680b23f2fad9bca01eb51afad55a1a57d13f1166eac1cad890bd8db53
zd8938b13e7f5e0e625882d5cb2798238273299d67fb3b2d6bcb9cb6776ebab207abc164dd757b4
z231bc1c3d7676c58df5edeb33d06ecc674377b2d621c819124a6eacaa5b713ff3c2eb3b9c9e2a3
zfa273857859be1533c88a1bc8643419f6d11cd958c07aeaeec0abf051beb62cb7dd73972617e5d
z697772cf82d6be48644ee3584d3746a00f80453dc2ebd00ae354cd605aa66e64178045f2ccb653
zb255e3225661c3f62a46c2d670936e5fe55bafcf9813a761e160207f1b63ba75877d89b0a3893d
za35a97595e5922fe6cf2f8ae23ce802751482651ad71d997bce5a34b484f04318ebfc396e525e6
z3e7c6b5f1831e3358479db6a2082bad05d76cc7ea45ba29abf390d997b12e1475a63a900bf6df4
z334b40eaa8a3572fc9166f091141deadc800cf4d74b66fef726432e85c79ac351b9849dcd32a55
z92eb8f98ff44691ba65971ff72d2d70f4f99b8abec0e581398b3d0c90692f94076c525f8d0e75a
z8ccbc180878dd91a731f65a8d096868c86a64fb38abd3d30897ddd18d5302f9981c9fdff530bef
z0b02f2527e04d54bcc2c359aff17baaa2d9bfb93100ef5a1d90741ef0405cf4d24fad0f60a9931
z9f8a927dfdb91b3abd123c6f9c65825a156ba5faaf4be3125950e8974497b78028c8d586e9bca2
z5f4f2f0d86956c18c50150670960a6d6553cbde1f6f52fa8102408212508a0e473ca0c5f00bfe3
z4b481edd9751ab874fb03900c60f148992c44417025299a25a9fed25df4ed8720c0f7a53410614
z1f1d737590c585ed60fa44b5c9902888f1e50b28ee5ac5c89c507d3631dca8fefc81b944feb8d9
z2ab3987cdd19ae657827b2a74cdb49ff3d836cf59c8e6b1cd415b1383eca4b54a484c96108151a
z32f008f399dd909703c2d85ec6ff9ab2c5b7e2164570ef27124ddad475b672e876f5666b4dc06b
zcc919b2680f87ef679e77b70a8c166eb1ce5e318f84330282447dc5f60653826cc4b31e05e7071
zc8644825a7bfd4caf0ab3495367b939fb3e2d20e8a7eaa977d4dc1cec50a588ded29995ee2ae5e
zd63b1c8e77a66990d627a57a8fb495bc82fbede2799e2a033ba485b666316f4191a0f5da8d9a13
z731107a9317077fd0ab2684774dd015768e37c77c71f4623d2267b9a76b33afdc82fd5be7f0c8c
z3df79d3a7be5cd2ebe8d65ae7f87a4830ffb073b715847aa8b5825d4f9f51bca9ef3e13f9a0ca7
z303102a46e72032fafe68df40fca881930b2cc1f10af504cc5def41e63b3481b3fd7c625ceda96
z632e0a870a3176f6827e458311b3bf3ea6c54a1e532c540a22e02d1fa7aee34ea89b6d42155ea5
z1f68d8b731dd8a032b12525da6760a6785d29ccfb25f69bf563bcf086e4eef5993339eb72a8278
z89fcc8351635e5b62bceee064a580c5b9bb2d53abe0517946684c143f9e69fa8f9d1d707c5ea26
za7fb8a010dd7b26eb3e3c193240475aee9d8f9fcd71273438668e156477f9013b3f5d7813c6af7
z50c43526da8d34ccdbb4f4dd073ac227cb925f44ccbda8bd67d9bcd788b0484e0145d899f70278
z15a47a0c2a20b8bce21450708e42ee52dbacb4b8bf75d253eae53efdc8f8689ac75c3ab9099898
z9c1b2e4470efd2106cd6b56ef75a44a00e4c09f52edaefd8b5e8a2aa6e681db4a4ea5ff356acb3
z50a3372730f63d33adfe9d32b8cace6358f89584032be42dbef6358a210615469019d00f3b3bd4
zed41514a97bfa559733a54c9184c833334165bbf8117c0f8aed4bae4ea91a4bb1e23ffff9cd979
ze6ad557453651892b841996077cfe6c9b3e7df3834f2ca3ef5d91ef6ceb79acece200a0f7835b0
zeea2dd322ce8e3017bca1183ea6a3f26af89435d3144701a64e8adb133255cccebb28680a0c78d
z76c3f293f4a8def2f43d26faca7f0019049d15880da6642e6c566424eb6b4caeed9637b6f36646
z7f28438affa520e5643147bee8e235e8477a4cc0b86e82febac74ac30c633ce82aee74b0a207f6
z1da60f579be21e385eee314c2bcef7b38b2e6d8450469b882d729c4577b2f115df6be2023e5f4d
z9605bdd4af0da74e3e62eb5f36f72eac098d6a324dd930b9f7b35933e3a72e6fd61ebbe2189ce5
z6d9b83b9af98cf1117bc897ade75f8ef678c6be945c84df6341f787fc92609973b4c2fac2d749e
z9f5070d480763f6810ec05c659ce61c628ab8a388669d7f01e3bac393c0e1f023e8cb6648c6050
z122e074c773982487cef17975cf39bf9fdb0d6db41ce58cbb0fbb53a8b87b6600765297b0dceda
z2e50bebe11e0ea702afbace2dc463e0e9e7f8c2508b6c4f825c7639d4e2331885749686a71b3bb
z65416488d0afa15364f0f8792f1ddce097ace05fb9108accb5a7e036b3fe98223fcda8d32bb193
za6a22659dd3792c57c029974b5665840d323ba7d7268ed4ab7052f418e031b003e115566e12d29
z180df3088d0ba80137c4337b6866dec9fccd8e6104bfd83a2fdca4bd81e0f97c9e52fb54650ca2
z876d0f5fe6dc3093f0da304c0e23e1ba7b45d56cbfcb7f8db6683dac6face207b7aaae7edfc2b2
z59aabe149e800ce539465c63e97639c93cb8dd79fe7ffeda7f60bb6bf4ca432dcaea7ae0428bee
zd504e7bbbd904b7aae5c49d87d345d5ac75160a34cbc103160141425967040710a77b3d7485b11
zc11e2939eb22e3a729897cf415448ce40b25c98132f897ae33f0033e5603a5c2e1dd027c003b70
zd90aee7621ebe8952ca39a4887ca07d46ad0eda33283ff664a048f4323e47970e58cdaa3e94330
z5342feacd565c68e4e1b7b85d93f7691b27b90f063c00548684105cdc35e801ea4448b39eee323
zd6bffd424827854e5dc37d01e258fda79153b491892fdead76d5990643897afd7bf8be75494367
z91cc73eeb1bd87da01555ddbfded96965da3dfc333ebcd027d20167e1642d6038a75a4dba0f46e
z7f16963f8d4b37f95f804d72a3691c91c17ce472754ecbb8de5eca1969859499cfbfd96dd9b9f6
zcc0b49f4ae51f7d8de74605b054ab856da525947c400a5adb711111b955a4006f54609eb0de8e1
z209d902c321397f46fe5d9a16b4741c65f24cdd7e9e34dee3d3a306523be553ad97a3a2f39181c
z750180b372dba7ad1c649475a6ca4d615c630c73d01ce65c87741beeafb01e185f4779c8d47096
ze871f0c914ce8a2c4ad36aee5eb3d8c1d95782cbbf09368bafe8851d2ebedc85d317ea774ee1df
zc5d8344a4f7a35fffa790d6cca2d97e871831a6514f0788dcfe96d75f036122820733f377aa40d
z0d9c56eb3a7beeec040b31cba809942e01d764ca6c4859042dfbb96931136d138bb44a8b8cbacf
zea91f202f5dc8a9d192394e98ec0877f44eeab33cc1d69cd58293d4c4bc27ed3741456d8c90b9d
z20715f3bd126d9a8064e8049b307118d84339f5f9d78881f2db39d91b8bb9c9eb3e71a7fcd7b61
z8219314850cc6c0de5e0ff4ad75d515921338226b599bbf6bcd8116327e78b19c31bba2fcff405
z9de2e7e9204e2c87cc396cc8f1c98efee69a61e0ad242231cfd0d6534667a924433018d8d64e6f
z0b40730e32eb6517003f445158ac984a31c6e945c745e04a3f13ae75219b8e671e8a3427d2ea31
z0f3fc90bb98e4175074eb7378382f46fdd60b5b7efbd68a5b96fcb38466bbc76b88de919abb313
z52358f4d557580b0269f9edfa7daa794b5920b27be3e3341e965f87aab71cd6629d32ba82150a0
ze4c0451697abd5e5c70760867585c5f1b18185da866977cba20af52961fb61b9738e641a68d5d9
zba1890d9ede84d00f4523addcebe347b1b7ccd751f55f5e980b47c62a72293b8123e7471cac4d3
z0d05a2859f28a49f26a489bd0855c847a3bc25bfa9a2075f23a727ad6a786c95fe7d504ec0c65a
z50693f73c7979aeb82cf6317d6de544d1d50823bf06130b0eb984f36c7100cbee60002bcf0459f
zc5dc48edc15b10ca281dfaf53ac74eeb242e71e007fb0a38698b0a9cd86aeae2a7aaa5529daa76
zb7157df9b94ac12a99d9573804d827dee7b8145a55c1de24f3328e8ccc5977ad93febf3c852b1a
zdcb935222f6325d4d248939d4d9773dc012d7c65a456fe9bbd611ce4b2b41a77428215ac2dc45e
zcb4ca85679f62aad64df50ce775ff7455490aec831bb603a0b5e6a4d05b4dd85e3b2bd672b9def
z34952cb951df667216375bb46f3d2874598daf158a09706deeefbd8c8183ab8dd8940b5cfc3d3d
ze816b6afc7e81df4350de225050886159fceee8ff0ec09e3ef0bc4c23091fa0b33340e0ea6a45c
z7b3e950ec18c1313d68600fabf3bd09e226c09adf3114f0e1f524ea9cebd498e62e5178519a1c2
z63a249ef68febc636c3b0f581e9e9ca64367268552159806985ec3f73d9d88889bf5eb6796cd59
zc258bba995e0eca8c220394678c68feadcd9636232daff0a2809ec03da49ada2d622fa0c9e8b8d
zfa04a6034bb09126f8bc803db7358e968320c17b2d61cf06b5d404b4ac762c37801e5b0457952f
zaa5539f6ac1e757358ca1d359c3489ad581e105dfa85cfed5fc12c3523ccc3104a72d6d4519832
zc458dc9bc9298a7ba92cd07597b930e543f06e888c2aaf6fab28240ffd7c1a93c8b52b142b218a
zabc3bdfa3a9cad88348190bbfd816b78978f5674d5ddf8ac4bbc8427fe0378a45fd692f504d465
z4d1f8f4de0d6dcc418ce9cbbda0290c255860efdb8fca44137ae51617eb81eee1e5cbae0c8dd90
z23179a7a08842dcaa4d45d61ffdc580c63839f409b31fd8f17af0e8ea7ae590d5061d20956cb83
z9751c8b04dc314383d4dfea986188fcc525250903dd396fb8fc19154ca1e78436de45c82a05e83
ze1f38785e10fe064577c9baf08ba357f2d7ff3898f3d34acc641991ad80deebac5d40a157423f2
z214aa18364f627b52408709fbe986c3af79a6dcd1e6c4d53ce4b279f667a3a872874b16a40d17c
z2280b175a7ad3c5d17b559f1615d96e9358ced9f48339078ba0cafd3eb5ff97e1a5b15c95c68f6
z8e0a6411243c2262f1fd9ea4d862865a0043e4ce4fbeca963cad8612587f78955bd6ab99e7b35c
z6e69df69e42917630e7fcab1e040177fb9aecc565e9a642b5ca5fad953acc4e3a66606e5540b57
z2f60086a2ac43585d985afaaaf90fe9cb4650173c6f3e1440c766d27c3e903879c628311189965
z4aaec41dd420b28f255544d8547a5a5c460bd8d62d0c85de704ea88d713078397cf89ebba28d8e
z7576ba0c53623953830f0c3f1d5ea27eb4fc10e9e74dcda1b8570ff16042e450697458474049f4
z61c26f8dd12a5d0336b776a5a4bc3abeb261a4aeb1ee213a8cf130a6de76d708bfde9a1074263e
z87bc8664a4a922fb5e0ccfe81aaf8064a79f7859662db06acd8631f1c0aa3544204958d54b3a44
za2d271db9599721b799dd4ac6743a505a6cf377070be4c587c5a2b6f52e03242304e4354ef7eba
za8c819fb921be109d7e034ddab60203d077201a98a37f47bd50b3bda80308c9f1d466fbf894cfc
zbda9716acf4311ce9a25665988885a3e44308aef35e99c32d8f79d6f49d177888d5f7f335e4699
zdbf4b9114a4265019f004a72753290a531610f72f7c24f35510b687848ac9b623576832b8779e2
ze51065f546c3e69faef2cbf3fdb0d41889ec8785e93e7c91d899bc11e8df717e544dab9c2c11b5
z9f8f18496303017aa4642798b22afdf0d828d7c63d3766ad11f0511840942f6d4e7d01585d3c2d
z96374dbe962ce3726f30a5a67fadb0c6a70606bc8cf3fceeb10191eb99e0da0a3c32cab65bab5b
z2b433292bb8fc85b84c2f96ef6dccab308308e7f51b98ba2d3612cf65bdbb754d77e01f88d4a61
z4e36dd1d9188e42bd4ccd3bb8829809f7ce4597b24a5d295ddf8535c1c1ab6bc500af13a75e3c4
z247188fabf306efd3ec98a792ca0233bb330847a7b079f4147e3151579014c4b54056e910073f0
z21e08f8d50bb28e1b06e001b0f78bbfe257a3c36a9c648cb28c4bed42fd482eac5d44f0f11abb1
z62a28999076d2da0cba6e96053cdaa7c1c5a20dd324d7d4122bf6f06de2b66eb4060f8ef635063
z2d75fe28f2179a974f98c30d3d0d9258673b4ee72a0d15d6c3aa474097a097cc5cd32624b37716
z2dfa4ffce5b6a904b224ebc15442d847b5af21160c830846f1ccb26961d844432a6ddcde0cdd62
zd2438e99ce46cdb7e0e73bac0a679cca2949c3facf26cedee92f8b2aebdfe168e336c3bcdca0d3
z5c9cb864618f3eb43ac6d05cc5812a0cdcabc9c256027ebc925109b3e2b34d99eef1f70f5fb801
z3b4ee36109bc66a046c9f1af6662acfedfb746a0e04f859b0e01aef2aed5142f48b77069e55e52
z855649aeafffe8f2ff0a09eb9b613bee511508757697d53dd346d45bf10d21bbb128433c98d106
z9768d87af1e742cd70734be6ed96fa71bb357277656a605932126837c7381601c92719792acbb2
z72db959ba181e0f5d01c7cf4d8b2fe0fe705afe189be4c8d681293d6fdf611bb9371f10a3c7fac
z00ed5e3c6110e0b1c2d7d0fd76388c9a3b8900b2904705b09a103c5f1cc93fdd8e7e5f4d6fd572
z672f19908c5d647e6a02d7146f28bbb82dfead23a9f74a60e53ae0c5126a78be6db337da0d833c
ze9529b95700826ac6edc5f27d52289130653de936bfed7afafaff1a69fc837fae4c2735e651804
z4d7b287b9432e368d43208e8a0b202ce39770f317d0fb362863cdc9dbdf907c7b16480e117152c
z49206dabd7621d6e77f3d8839a714577fd1b508ab75aa37d5d624bb98f982159b31f93fcaa43a7
z80856359aa906f1116efeea4ff047f72b84421f8ab3b886baa20dbe6a4ec4b89e5eac24da0b29d
z30e58f439498e88bea89836bf4b66421247f46890286b1067414bb7f98ff3869e80d054937824f
z573a7c1240fccf6e9526f664ac4ca64b4eb7eb011e6eb8bfd8bf4571ce8ae38c1e08fa1530a57b
z2f28db52f33b526ef257b0c129250a041264829652e4504ad003254b4d1a3810840d93cf3e4e97
zacd7c7ff49eb4772b478a55855c977b516801617361c8c4302f86ac99e2f5d0b5bee69923776c5
zf02738534a13429edb7aa62b6655817a59b169201c65d0b5a23f09794ad39400988e48c1af6379
z90d6d11a6a74b03d15b06fc0791c3551bb64e52bd1096f0f545154240a0ee4a470ab973b716da1
ze6099eb816aa5c8c2478af94b613983e32b68760c3e89185d62131b536a6f5bfc89230daa99fed
z63714818a1a6d64790e8ac4ef10050d97f95af9876cb455fa152f8cb94b67b113bc22a3f0efe23
z2774cd7cfc7e41bf0cc1ba3171173022919b53d581f9cf9c92f98c1f9e4d2a5b24bea66a8f265f
zf4fa4d515931d23a6e4ca52b405a93814c861c9118b683e5391f1b301165c365fc0eced966031b
z5cdb330ed9c3ba7557e489d484ba55772a4ecfe045d0f25785bbf12c0c5f52b18e3a747dc967dc
z3f6004d9d769a5011362d939a81d4aee6782500af2c667a82f02f6f7c5b71b76e66ed98f97032c
z684daba1d90d9292b39055e781aea986dec2b399fd09cfbabb6e39e47f9857233ea56ffeeaba9e
z663e01f0d5c0f532d9e97b351c4c3aaa4691b76ed5f8065d2517c1bb683fed25e2a8d559692341
zf2d5240a7cac19aeef3414fa60f3134ded848fb8536810a554edf4386e994c7a55beb6714377e3
z0c9ac4a5442937018ef6a05a6190f717f9d17d95f7ab2a493412d10dbad6ad07e782cdba2c75ef
z1156c85ca860fd9583911cd01df9dfa44e3e94be4ea461db2efdf35f5fd1687ebb5ea685845a72
zbe62c682e595c6c6780856886e8623b9a9184db20657f5b6d192709517ad99689ceda7da88e578
zbafe372fc56b3d08b6aad3ee741b1ab74c690c943935c225a333a4900f0515803c14198f43b77e
z8b84fd1c6536e75f28c2550f5ae5d3f2e4b29ead2a7d62c544d9339bbbf58a9e35da1e603e50e5
zf7f322b3d843d435c90650387b73b4e8a54fe11c0c886d4bc24431b50c0654963b08666a49fae3
ze42fadc6090ec45cd6ab62f09fb9a3d28deee5eedd798c1f17f64a0a1a2b7d260e9f20550d959c
z3d7df6e05bc7ee5eb372411d8122274962f077e0f10bdca93e149a64523d677d425bb654a903f4
zaff77121544fdd6209713736ceb4786f76e7872f1a4d91855c5f367f26a97652115187b658a98d
z3e1bd3c8cea8036fa84f6fd8936839909ed61217464bfb2b3d1b283518b341ad2a7dd24317119d
z11296306ae79d235002eb27482610a3fa401346e598698db0263a39499ef2d1324a88dfa339f95
z16b9ba12bbf6f8922526eda5631ff1d138fd450e6d76ec7351405942cdf2c7e76022ca0bb89ac3
z761d5f486798a990bbfdaf94cdd1cc6d9352603c02634d0775265a24f2874106f503ecfa7388f3
zbcb1da2e6f5f807410b6da8ecb9addc996d64deee020f6a2cd9b406bd9d9d99f4f0077c8dc62f2
zfdea55085e544f32e20214cb8b0de21d1f286694fd753b2992d9c07f32a9bc472ead9fe2575214
zab3b2792cf2503a6aae1d495dc779cfdeab7303d3acaef977a9c5fea1c37faed1fd85f60253a65
z22b2e07fbdb04b7910c33a638e29757a50db8a9da9f7be7727d8a19346cd5383613e04ebbe4793
z7f86c7ffdd8fdc1842023a2ecd31d14acea486962af80eed34a834e6e264e4b35987e4240f4f8c
z96ece019f034454495111f95cf0b215867ff151b78fd5eec1855a699f3af075e0a21e140b64e27
z949fd200293f9a14e6475989b2322b2729d10c4656605e2ae4ebc7444deca3892ae09469fe9f77
z956d0f1ed913ed1e15581dd4ef5fcc27c489da8ff6bea18155f3716f5b3a42844e2f6939e9384b
z981478dd34b8cedc70d0af3d8135137fdd335e530af0fb92a22950410eff0b43c6e42b27a54c17
ze7ef7509d89b8298291aef257d53c6584fb35cc7287b3bebed62a6c33da3d0131313f08155486a
z89f5106c609cf896a566cf35f625cffde0ca60bb8052b8a5f7be0a3f56d3f2d24ab3f5bf55711f
z72c3045f44698da8867f8c12cd90f97a2b486d9f1d3a28e63af7526f20e2786d14f9f8b50ba107
z1df3348e2abca3385246ffc615c17341d9c2506b08d729fc35441f49e8bdaf970fe026d730b285
z5f7db14ced46c5316b4e6a9a767c48f27a09addd32858c90ba0d7d74dfcdda747717f4624d9d9b
zccc2084350e55e2bfd32a1ecfd5fffee06ffce241b7b72bdeea0fb4dbfc0d3bac008458aa78af1
zb97a724296e20571cb7814cb3f80f139323a78dfc11b049f8851498d68365c305c011a67c89b35
z551b808ae36e5348357c3dab558eb7e8b56a9bb6384b46150d17dc19e4cd19ce447950c563e8e4
z4e022588831fdb2c7dc7a797adecaf72805c0afd7020833257418212c62f5f80cba9990bef9249
z8fb714c0ae9b4280afaa008b3aba64c83f6f077971d08bcb9ac6f61fbd32cc484e53bbbce73f5b
z1b7b74096db71d0a37e65a020357a4b5eb4ca8ff0825701ab2a469ac69f3095c372a87dc09dcef
z72e00dfdf4ca806a7e66d1ca2a26f8396f19820685add80c0ed93d383ee47252b0d12e5dfead27
zcb772cfeaefc0d0b74e9d1afaf49c0c80fad0cd5532f402599b46c0eb47f6565b94d348ec57d67
z05f129c91db99ab58829728874d80dc9ccec605d0925310610fabed8d63a26dab1e825a1d8a377
z84d1567e700c2c5f34bd56e64c82fabdd5c6a657960cd7d317f0d2423634b4a68d8427e5681eb3
z460cc9005573f27f83c5db36fd30a0ecc439aca5f0f89f3fc4d9111830349950a43341d5f36a48
zb43dcb9c89a85ceb7817ec57bc5777d2f9f3b65a0aa547d87ef5728ba2e6d75fe184829b92d366
z628ea769430207c51c3b177840a0204dcab0b3a281161d94800fbbcdc338b1875c137d8a677ae4
z19a330000e8f8f97323d963593638eee218e1e99e2e7749bfb32f2ffb88fd07416c129b0b8a6eb
zd49eca516f736a936c55c7b8ed868feaab7ccd11ff7978f2364b62e70ae2b154e86ddf56715448
za8b1771515ed99dc84aedb39fcdc83d141f57a7870d0dff1aad1eb2b5f7674e964477d4a5ec514
zba127bcf2506bc70ecaa68b4ed09fb54deb2efb10e8a97df0b067f4ee8795a24bbb5ddd93bc97f
z9bd9a6c9ebc8ba97de7c2ada440cce51c53f865806338da0edb09d17562f8ed3a32cdc7796464f
z74dd0c9116f28ce5f6d5f1f1f68b38c7e9a41dec55c539d251618b9552fcd1e1358b73821356f9
z7de82e9e2a1cd1bb0d6a0b26d546f9914b79eb410d0c4c5d87e9dfc4d877a0832b520cc32e00e3
ze3477b4d3c8afc77567e8ba23005c9c1d9d2a369325b30ee595747b533359886b337827934a17c
z3b69f355da4de4151c870fb532e3cbd458bf19711c0731b83558d896d5f10ebb5eef9748bc1e03
z1d2d50869692362dac557307bd06d4f4ccd7ebb4d1272e225a174ff7cd7d7ae8604ccb20fca8cb
z2b01484ff419dd51dd05e05f9d18e3df5b9ebcf6daabe9e9723d7feec1803755bddd8261a5aba1
z410203535c6d346c29d09b150dd465f86c41c69c3e682875ab5d2cee38e1615b1fe68a51b500bb
z7ef276fcdfb41039f9edefd88c02dbf4ec8ac7eb5b11b64649d25dc1ce0bef52b0de95615dc659
z5b7165ed051e23e6ea9ddfc262eba5bfb71cf52929643789efb399a9e34fecb3de61958f6dbdc4
z2b470d2cb9e554473283bda9df120e059eeb1bab1cd70744ebe1a1bb4723e378b8bbf8f247e66e
zd7296fd4f29b1c6863812fd14504d20dfe7b82427f89269cb71f291b4c65fb94ea53f948953777
zb80c5d9c2ab636eab1efaaaea47d0229ba664e9a99267a29c184e8db1cea64e1756dcf19e8bc8c
z669636836d54222ffdf5873e235bf4a3628d9a36
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_express_link_retry_mgmt.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
