`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc94254008
z852a47c12c9670712b4cf92255dfa2c226052261139d0d5a2f27a39bde6d7c3c2a7a36efa6c1a7
ze784bafc2883e5cb6ed9fbba690afda2f8f67125e033f1ce96fd0e6f25974f49edadf5ff78bdbe
zfc52aac4520156816e11199f0bbfcef9df89c560353153ebf74d0985a3bcbf3b8dc385eebf3793
z4f73a92fe8f63acbe7987e48d913e0776345e747e52774fe146a792fa01c75d78f1de8b0a25186
z4f7c5915e377a253e2c4768f7f8ed05368299c3f4f10360d6ac3028e3da8e67e2dd5e38105829c
zf373a3ed5f2e9895e28a987bf6ac27e08a2e628ad02c54d989ea4671c80c3ca0e4251636598d2d
z44668c7f37145f02a35543fd907901c12826bbf928194aca8325012e606c2622ad6d4f2d603de7
za4e4ed13111d3ae3b820cf1bd3195d081542fb4ea0b8187263a2b7ede95a3cd4efeee718d17e2b
z3612086df976d5faf134e95d41f96aef6aaab33b8332ea37ef2bafc5602df9d998ce8fe23ffb2f
zcf7565a80c9b572d8701576f0b6015da2d6044f7384148e081da686bfc46b5ec605106031f3c31
z5f1c8ff88816de71c100af313a5ef6e312f17b71e707085c7460abd427140a3aacc88ae1c6a51f
zb3d2f68ae5849f72824519abcf297f74ab2b45d9f454802190e7567067ce4465c5f5031370cf29
z90ad42633a4d7b9feef3df21672a13c6761f3859de2a236ffa7ef32e50d599753ab36d56de77e9
za804ed5a3d9ecae47d3c9374c447586bf0717ac257adf509c788dbe31bb056297bec2cadb8415f
za4e3e907106846bfdab5eed145af6f0f4206cd230f9a7536bf7ee7902725ddafa862c932d0d7b8
za6bfb037fd2d57e96748ab415e1d01181c8ca27f077c72891caef59bcffe55dab5896233ab2090
zab74954e51c9ac845d7493b7462972e3c9f592ad4f532a101699ec47af709059575d95cb3fdf0f
zcf22708787bd5a8f5538d50229bfd89529491d6ccc5e40b311ae30541337217b4cad56362b9860
z59a70bc8935f84b8a5085a6b1b2f621e7b3c1de80da16bddd10e5064359c71f3cb35d752c8f877
zbb4f39c9f58cfb8be6d70de9c6bbbb08ad3cb222946c2cc95842d176a3262c038448c7395aed4b
za95780dfe309be36ec0a78e126ce117eb1484ff3bbcb38cd5c29523a0245edd81e0aea1b5c480f
zc2f99802f668b41304016a7d846f1e695d015407c91409ead05e43e487337d3c72b84df981f25c
ze6b2e07d91887533549183ef51cbdcc4e3b9d3175a63fe86a8b685ac8d5e7bc3ecd2af74fbd893
z0dfe242bf3efa91269b7e4a047c3132310b19cf9a3703cd774df0c0252837989e18b089718879e
ze2e687f14bc726a41d01b29b9457d312bbf5e894ea218390d4e2ec0d76c87a803c1173ddcaf115
za563ec56f4906c6e76c8a43ad535dc736afa385a7a6e52e3313ae4e59e8cdd0012aa3517da56a9
z751b94b0c5801dfe01637230e6d4b0b8941224c52dd14cedcd2a4d5e72da0abe5c94ab9eef03d2
z2820b4970fa760aeae3aad86d3bfd02daa1141416c5820e68421d1de714af1c93dd28e4df1b620
z359a6c641cca873ccd9ff40f69c90de10e509e58d6888b2e6d785b3c61f71315dae321992118f6
z5d2d3d65c1fca54970b1d22b6163e96c151d7d5291baa10885b727e5c7835131c9df2137dc78eb
z82e07e358cde30e6e0fba4085acb90cca00fd65fe43d5ce756ca117b1f12feb73425cfd7118085
zd5e35b05892ba0fd27aed80553f042a780ef6c29173e34ce182bfde2e8b0caba526c1124f96e16
z32f6aba34f50bc23e4eb8b7515320cb58c119732f48d46903e23d9c048fc6422d3843d06881418
z51b0bee695300c0363ce68b2844bf28bdad136321999ca4c6fc845dd211bff366846d1d86d4261
z3622c86b5cfc1823dfd0f5914d77656cb272fbadf9fadec77f5e22a311a332a2029ade178b0fc3
zd1501851e3350eaa4a3a4e14bd353db898f6bd7178740bbc0b0768762a76c9360ad42ec0d946c2
z883cc4c16017b8691758634e22068fecc02e5551ed2cc957d81d5da647d86dad20d38a468246fa
za7be8b6706acb6b92cc7941acf451d453a37fb6f7dd8dc56196126a21e65b361db7ace9273669a
z0027605c86d8fb433290b2453efb20961c2fde0c65bcec96b5db433a197fd24d01ef64a5ed5874
z90e7a2c402b90e8f23115875b739b01927a339c5a3771bdaff2b764d1439886449a7bb98336eed
z21e43e4de293edc3131801c1142dc635e65c5170b693f3f613f99d8d2beb0fa84566fd7f27901e
zfa238d5f802285cf34d76f41b0e4bf74bcbbca5235725dba7d1d5d05868898b990fe30ab899b77
zbdfbcb50dc2af9df5702c277e40972ae60e50679e8d616b38a0a4da7e374555253f4bee03c4e8e
zdb9ea2ca62c7767674be689e10be085683f179037daaf4a5d2bece5c8e290849772afcf82bccbd
z67fa0d945e33e2d8c59d9f70521e8b632c68a4ddc9fe0ced2aa79295a95762538182563a15212b
zf4b3869e8151ab989ed35d9243337188329e4668eeeaa8d28289dabb7f0267978bdcc3393d1fbb
zf2756b4badc4d213e8039d47e0b83d367c19cf20e82965fbe9b78b4c2d03ef024f3548dd692bb7
z5ae4ec97120d9d08505b8c786b3620713a120a2db2897274e07f553d1c09d0d0e2f2174d5e8204
z44b31d6a799b55208563717a783a761efa294e7087ce6f651c724c2cd3cabd1b181df387fa1767
z18ff4016878d967f373778d514a7353679e7d0a7f161140373d518c25b0169d5ea7d744cf735ce
z0cfd849485100f1f2926b3b5eebbeb4626f16da00cc604b17555f7117bf7780779a967e51d69dc
z812d149a44817f2d46a2f7ed0999193a79f3423de6b338010e24b4c554e24f1d5c2df7ec0dc323
z6d3c2113942238898ad371ce639460c5631462b3f5f8a3bb8c5cfbf71385cf0d9340f7f9c27b53
z02f02275d78ff0c3c3cccb76fd2d17d12577d13cdad8f002ea7acbe6fe905169812a3bd944d421
zdd52996e41c3f1d86fe69a7f785e61467e4c841ab5d31e8055e4d8761b49c21d40fc946ec8fe5c
zc61229f6df67f20e6103d03edda77c3b2b19c149df86d9bf557b1e11539a11c9a5c8f6c1282701
z5b0ed893b376954cd62daa576e8f03d95ce210b5933e31ec328a93bf9416b5acb3c97188dd2603
z08c9f801488dc88bff2b3f87629d30f9a691c3428ef681c0c902f88d0832bdbdd4e5a6b44b425f
zb293ef267feb952699d13f9c30d025a6c23afb05c5af2f1cffc9acc2dba419207977f72a248abc
z1c71cd2a59337219fd81490a990f598b91f0d10e69b58ffe9691c4825bef5d4c0fff9e570a6df2
zc170c41a56ec0f543b04b955b5ce9d612b4b68ab4ae774f9a49775e2e9798b28edd3dc2de2d018
z2edff202cda6ab0811a4e11c46bbb0381f843f8a697af79a5d444a03ad7e0c56f5d7166e4d737a
z87c360bc93f8f0da7de95d869f3065d7c7d9b13f6e873706c01bcfcf8ca5f78485c65104bd0843
ze59aa6105d629284891b06aea7bd9f726d5c9042b47384dc39409c63ff6210ac3685cac0365883
zeef7367c34ed81157844ce1278e3aff88bb8fa26642e262a11b87541a5f58950937f4597514143
zc97c467e9f53518bc6ef1a8642fd97ec87036003cf389d3c1fff080012b0a208d12902ca3246bd
z8c0b7ad8d593cc10d64ad5980509306cc711b5b076e7cb3fa4b212efc217de8121af352ab5e794
zea7faf364fac53f3ebe6bc0c6347ecc0526fd8b8d46dfb3db36a970ed82754225b3e11b58ea1c2
z163ec5631a97be62879e04a50b359c3f73b4fafd41b5d3f3a19c6962e7837d6944868089528112
zde91d5db956fe3c9da3c1440a624ebefba661077aa434c4036acc009c5cca371d59a76967d1b39
zfa9ee19cb17317786b08ae2dfc7ab69459fd3093083663c54e6e38e5800085d197a415cb1ab504
zcd29b87a5ebb4c048142d72ecf56a21816ab491e571677bad6dc7cf24dbdaad02e2089353a6a77
z1e87450590367f3344207615dd4b97b0d117b16d242b7558f07cb7e5a6f9f1dea75201f89539cd
z9657e86bcf2fc51f7c219207b14cf261130b23b414de8a9e11945902aa210c147666820f89da5e
zf5daba6661f12c40b8b583f527b5971270a3744e7dd2d4d7fb327d34421e4469a32cf76e236e38
za03f0c1420db04e56e069ba7c1878ba2fc53e4074c7281cf6d9e1ca49ce20d63ada1dfe4649c83
z1fa16d3bc60a0a5def4c4349e29898a6a6b96ec2ed3b5c5e6ff3f29821f73d64e0102c16fcd151
z30a54dfeff90671a8faa2c2c0eed5c1b0d1f4ac12e457fddfa174fc7d6ef46d0dfd6e9d8c2b2b8
z503a498597f4a65bbaa3a015e3ff86f9eaa3175fae4a04d29172d94b4e4e268f3f8894588e68b5
z47e430b5546293569206e7ebb6e673737b4f241cc8fc88025954c9278f0865b0a96f726cffd732
zbaeabb1c7b3349407292d65ca17c34992fd1278dc49b1c2eda2dda4791788d6d6b891e8d462aac
zec855445314db6ab4cf136ceb6c93055670254ded0f0893f84a35d70b62a7a08d0d690741f8d92
zffef662d11484e909bc83e8a916334bcb56297b0b6d715efc231d5654a633fda9276cbaacddf0c
z5eafc5a099eabaa9a5ae1566a002c6ac21e8ec4fee5fd4d10da14930b13f29c579d91574bc7062
zc0b9c317dfc7d01253c77480642d9f894cd76b385260baf81e440b8e95cc2079a2d0bd8978b07a
z681cc3470d56b2d65853221dc391a33161c6b9fdcf54e66838d76d8c8e54840e5727adffd078f0
zb83586e24cebb58d3f5ddafd64542bd921a0f62b8e316711005ceecaf594102ba75806704e981f
z4bbc94e715652b2e04b1cd60e2466b9941d6a81589ac021d08d449378e33d8b10243c3b18587c1
z873cb043710e8bfe67709880455aaf7f174841e76e71e3066a7c258e68c6d041702c4378d4b1f8
z6a515dbd590de0d9ed9d77b160a1e3ea3c473fd14edc487ea77f2cf266670e70bfbad4860cbd1f
z83f8bb7bc8da3518ad372b8e0c09dd2b96e1aeff1ad9d0733377c034bf57aebdefdc474f4e8cb6
z0196511de2b12b023827651e45e3b02a4817b83b6e4a74ad2976c53199a1a4bcc2d2bdc11608cc
z0e3a7e7cd4b5938b9aefab7aeb87067f67a0094fafbb17fc7059a907cb9f43f19599f48cb33390
z2365b5fea1e141a5ebf71c7a708e8da4d1ec21b5ed5ec1f8fde4adec19e277c25fe465fefa768c
ze3f8ee1d03d6f259cb6933afd39b88f84eb1057fe2d27aeec448c46c95f30324fa77f4ffcf1de2
zcc8e10053f14c62bb4275fba76ab9eadbb69394ea4a5134e7eaef6c1c4432d4a9ce85b42e5ef93
zffcd8f5f9766f50eff504b483b3dc6130001ca73c9d2cc5d965326ed615ce5bd334f271d25e77c
z4c321994a87eb41d11e8893f7e9a705d106d687b820e85c423ec30aeb624dd5d16d737adb95d2e
z4bed0c01dbaf11fccc131d194f24d1046d8e56931aaca061b5060d4445010fc7913fcdb2e80f58
z24d0e0691c8e3a1b82d79507e815683f2a9a8ea97e23ea7d298b6545986a41d629e9a7731a61bd
z89cd11049ceb2b7ae370dae714a96c276339918f0cc08f3e7a7f2ea3c2e17f45262fe2a933756b
z8a87b891066154fc14eee231883fccbd0953172ccac2ea7e15674f8cb3519c86ab85b06ae21f62
z3cfd5c9dc6d8943eb8129fc01197233453368cb48912b197de1730408163e373520b1d84adaf6f
z2e37976612bad03f8f546201c236c3817b73aef0ed4659f88145bb889b7b1d98538f85318229af
zec5e24f57d62023b8f579022a65f0f4e0aa97e9932a9a55d64035911868cdfa61b0b2a1f750b79
zc68915da022c340591522bae1a26a815ee11b5bb5ff3c85b2eba15891b61e35d6f8f5bf45a76e5
z43d3118fb3737be65b8d3a457f4f9a43c6ac89931e27a63b574b5ba9903ff2b37c0ffeebebf3dd
z7fbc3c43d8ec87b7295ec38a8113baa9b8a27133f08146e39ed4d71ffa9a9d337db1ccac18875a
z037870fe5313b1ed30eab2886778e08fce723697517da7dc616305eb51ef9906fd919fdc83be03
zf920c56703b5a4ac2a9f93119dfb31f4fbc5216c8a8bb1925ac7c298b3baf397ef21d391ac7a17
zeeb4f067f5d482e2066a2bb2fbe7bffb76c26c59e931cffa4cac81b1be2d787ae538d25bcce5ee
z69e1b6788727970b796853d9b9096ba81510dc80b1738344b2a3858471b7e9f8ad77665fc35fb2
zf001013c620b0ef24ee52d106d341e48a34223cf09fc2982b5f4108c0aaadf1a5042981c56d706
zeffd9bca52be4e069531bda088acd6bd97a123cce49f32a955540a438d000b76e0ee0cd0b00e21
zfa512ed725899bdbcef71c36c66048ae7b8fda9ff11833c031b08beb2c7d4909b49c12fb5278a2
z0faef1c5ff121b834a7eaffe9ad8fa17a0f2a5f64681688f2c3b4a017754944d1a89571e50a848
z1f1bcefc77487b5a554da96007e0b81e829d82ce3ded72807c98ec82e9cc5310ba494a9129d3a1
zbff5324be5cf7ec20ab9c14f67fbd485a549ae7a50d5d5cee724d04532ec59918cb00cf1e9e083
z2b90634cd5543e9fcbd324fc5ce248f48b5193c378ff7b10b8f7c01cde693e9429a8b92df3c516
z7d3a497167769d7c99684af57333511befff1dfd6507e6d8cc3ade9e4a800e34ab758517a54035
zb213b2fb763321a04943c03fe1eaf9eecd51aff87ed86ecab0ca2c7c7a9582813694992a274c54
z1aa2b1c5d7d1fe2c16ce7449f7948c5e6b9d487588add4a5377ce26405d8e998652cf3cdebe275
zdf4fc6696cfe7f2eb1e7d24925a376c78ddaf74746a92c65129d2d7caf00519e5b411ad5c4264c
zb76c7bd21f873fdcd576f9e1fa4dc00a3ca991d66c5b3430b94cbac2e2b531f7b6635e5bab5aa4
z9ec578da8f2e8986e3def40b0fef096520a3a6c0b9953b23972e64eb688ed7f2a6f8aeaa8db04b
zbb64052483c3755667874aa3a2f17b39936905ae907525c9046ca7a5ebfc0eb31ea1afae969538
zd613a166c088a2448a9d4bb8b1fc2a53d10733ed56f9d1586a853632248095eed97608cd008763
zdd2750ac34cdb605f178b5cdb433badbe40f72c81101f055220e282ad55486cde8e7dcb99d5a51
zc5e52c8f429bf47f0d7f265ab764361be92b42e4eb266189ff8a5cfe1ec6912399d0c6438586e9
z7a98db0697a06528a2ae8758583e2eb7aa555ad0ef0cd1a714388960a3552b8482a5b92ba92211
zfc70de64542f52115ffc7f0c3d8aa22c1b881cbaaa1084d9f364a63a9a21f6b25bc8192aedb9cc
zeaca9d7ae8e0ec3bb64651d9aa0d140e42775c47aff4833efac504ee89f9fe85e96530d9265813
ze434a83a7e7b73545c25803c168439825fb1fe5b7f90c411623e835a0aef9790253165eee6d4c5
z811a3276538c6ed2015ff44437a1a0227c7740da92ff4fda64b9051d465e99a8cf708d057c646d
zde091abac5b145e2fb1e9438c25f1299ffc3b324f4848c92be4eedd4ee1dac64c7680a160c11ac
z4bda7d8dea16fe9f676187c4d8d56d94cc8fce5263bfbe7c53f693a8c8af503dec36bb919f0faf
ze64709458bd6f10f6f98b721b3053fb4026c6b14f12a6c35da504d9f257b98f6191091a5d926de
zb580589fb83cadd4a82b4aa1f20a46c4122face9abcfd6a4eb04a810296d528689ce1fff52f364
zf413019d6dad0b593d1bde5c1238a17c244c694acda8642365d622718bc4b095f1f561cd351b88
z440a9fe852efe625b6e2a4593736383bea860f16e7002785d1ee8795662c387dcb2837f4c0a420
zaaf3a8b2a304f335f5bc24badf72c3d4f45b6861b988b677b4cef34903499da5762cfd74298ce9
za82af5fd8fa6b9ffb773197db736184a23ff27aa6e082bfd695e283670f80c44dc17c0ea182cd3
z16b4595eb15c263c38b3b9b45281c1c60590b754cc47434c316fdab742f11d4d8e007182234c58
zacc73b21e20a1fc6a55ed1ecdcd851560f7e8481ecb864934035d0b61782270f94a55d9f3c29e4
zb599e8d6778bd78a7f7342d91243875d0d63f29c040b85f4a66ba07bfab58a7658f670eb26b736
z775f374a575d5a4de311153db1dff3fcc3e417c4f3b22a019e0e4ef9f053dd08d0f2d182056d21
z9700f5f0ecd388464c10a6233ee3b6800ad3eeae6fb383b92dd1148d8760f7e2eeb82f4113585d
z643935be5cd9904b53fb17f81449efa008bb5d10cbc4e157e2dc15d68b0eba6fd8b1de99d907c2
zd070d732fdc5663e7919a16de6bfe682a483a5f1241b2752b2463db824e8aa8b66395c63b9aaa9
z5d48a023526470f5d0b6762cb6c59cc97b564cdf697feafa6bd05ec4562e9d5ccfa4241ca0e0c6
z00262d298064f6b334ebe099777a1b81c05a02f6ce366b4a1efc5e9da59f77775d5781ba36c72f
z7890248d78ea4469c5e3ea0b398bfa36abd8ef57573c9509b313020600c29ebfc95ecda9871422
zadadbd5ae4330f646366d07f9bc36b8ee4f766adf98f84fe6e568906d086c7e9e89aa2f46e1bc6
zb1e46b795e0cd67e1eb282928a86e6deabbc456cd56aaa8cd6cb98815c08796cde8f859497fb33
z5a0a9b0775f3f30b47e8e09f7026d36610db7fa33e0896fb76ced749c92a4e8619d1d8c4ed01a7
zf83e464c958460bfb2df8ea4218f28ea0fc7aa9767e1ab612ddd1cda344ef96088ab7dee68703a
za1c225d247f706df2796ee8be304a86e95ccc75feb12fa91d05ac84d300cc1491dd7a55aff018d
zba288c9676bceb2dadc1b15a5b899ed414a3d97ed2999360552f6a46d578d26f69f7e5aec97582
zcb0938afe4bfee3c06c74cf6848b76b22f9fa5e278551993252a655b1fc9b3c9a3298b2826e33f
z446b1691cb2673e5812ba146fe4716987c5c7c07686128d3899a66a4b96526b87b3639ee52eec8
z39e9329f0df0913afa67674fbc0746af2e18b07fde63b3b6299231750973f70da54be28c728506
z0f8fb1987b5352e7e501eadbe6c24841d2f891f62424e9eb5cff213f75366444736ef1a4804712
z39ebf40a0867e8536316f20c5e2738eba6ef747fd383baa3eb67cbff378065df5436cf03512312
za9236defc2de51291abc7ccfc5af63ed83abf25ac6e9c2dcb0d0bcc7c3e277c33adffd80219565
zabf2c6550b99d403575d6cd825caefbe8194a9469fc578538a4f3f994ea910bf3874f96056fb59
z443df1ebc4843d41d1ee424ca343458dde7fb046df33f4b4f07368981e5b8c46ea29b65d374b85
z8d2f9d53db12354980d1acd68b2f99411480e44148b6657882e382fdfb53032c74d1c9c472b8df
z9b799e421ebeeb9c9d22f0b92bf2b53083f1e88fbd190f663f01965d0be4a00c065643604b004a
z1c4d732968ecaf5e68c61f1f57375c42c9521b14aceef5a359e3cc122c276677be359e0f1400b8
zd381886468375325a3a2a17f24c19d04aa63f7a890c73395e47eba4671151c45aff9e5962d1437
zf973a6a20ba266bca6839e38734ee8acd6c8c41dc0f7c8996141478f0287126a70e61d5d92ac29
z5709da67f31eea00a85a56e4826b942ae48adedcb7c47f724462d995372f61efd3e7a5701877a6
zdfc505eeca8e6dc05dc8491004923c0b662b3be25a159752e3703ee6dbfdf52d15640ee8c22b86
za3ab3294f6d94307579d4d262ca61f71ebcd301e5b18c9e7745c0d4d9a8b5797bb77bfdda5858f
z09fa9e83d641d45d5bdcff51057a41caf8298352db4920c797b7b42b9df418274d426973bbfacf
z8e86fdd1afec1fe7d5b8a9f7da2795437b79592a18c6a4df9670116c463585a998492b4d5640e1
z2d4b9ea76e51d13e28cc128502d371332c5b2b112a70ca92f7efa6359055a32e42adec46f17912
z97c936954af49d2b23d1f305eaf71a36724f0a91f784074f920cc39f14f935d3f9b801874d8e61
z20e71024691af3f636da5b06bd3f4877189ba53e0f5afe18cba6e93f8b2d80aa5904caf9ca148f
z8cca820dd3ff6c11146831b6a885ec4b1368bb276af81130dec35bb87f0230f2427b406354c718
zb51a8d3933ae7cd48ba6b7a06d39c43917d2708524af3aa830b50984c7a1650a0aaa6e9ad90ccb
z11e4eecd97bb14ed308fc0443dc47e0ee2eef667b1acf9de6a14af07945cdb88370586a6d9ea2e
z9c734610c372e5ebd961f10946bc6b3d0e914bd8ebce171efb6b0fa089b73a05b438b08e9fea9a
z07fb51ab36fbbe4a863a70d68221dfa06b40fbde9b274438cad3ea66f95b7efc401ed458394c90
zf95d11f2221943146dd7c90379d7bd830f3a5f7c2bad52b05e64b2284803a47f5aa5f24fde1dc5
z05aacd456200465ea0e3883a0dad022b9f3fba4298774ecba835ac0ff7b6fb9a7d0bbb63d612ba
zb3a423dcbea673070ec267e82f1e2b6af25f267c2bc43faac9cd8a266b44410c184fb5fd840b94
z859dfcf863899369bbb86d0d67186521917f377ef0e8655826ac802afebd1e27f35254916f8ea3
zc1262931815c00783729653216418f4111854ce634e3bfbb97671e5fc826655a194c166d56da6a
z5e13f636daac8bc0d9e86c944db42f802b510edf0daa8603d2ac9031056b93a89d2a432c3fca0e
z82000029347a929a6757d6f1bd5c73076df4cecfd7ce9e8fcdf66ba46f7820c8b796f7b4f56968
zcf5a44ef863ba93091ddb74786d26625d1e6b748ca78ec9170860b7290be428a77c08527d3a3b8
z26a933ee49b68d19d0a7c62a20ac3573cb51572346b8ac98538ba0fed7a4ebb839181e168c5ea7
z34b054a58251fe978fb6663e46b51187369fd09fecea137803ce7c63192a45de5b3ef4ee58eb60
zb9771ebdc374e3d8b5d16398efbfcdff01d423c907a4011879f1b4b3774db638c94deaa557399f
za495d0ccbb83b374decdc3bb6ff065bbdc48d51c189817cda9d93f3ee4b4856844bb787b544f17
z967d1679765d89a7daf522224f77297685f93e27cccca5e8adc171588d6a3ddde4cb3ba21ff2db
z7e8404f07569a4fd8cca5572e115ab28900f3744ae1d5d15dc51886e4ca1f97583ed37ca60d8d4
z782691fdd594ddd720c477aeb5554a8582676dd9fdf565671615fb18e8710cef916afc7d09e8cb
z650e58d3be35c12581434021e3d3678000269d0c72dd464e68fa7a040028a91eb7b38ff07efe10
z5f9b2f9fffdc874c41286cad1c3fd18a54a57c8f57f956b2a2a13ded1b1389b58fb5a197
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_mutex_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
