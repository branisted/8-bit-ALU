`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab30857016fc53a
za25afc8341302f0c829d94450c399b8ff9b0386c187cb854ee330605b7b59da379b1f26f488e1d
z36e675f0b1336408b3a1ad87d0723054f952fbefc8d5a33eaca6ef5be8f42bc59870a29a5cc9dd
z4fec09ce6e44cac279651402e7e1f590df88ce49ec26ab39f12b4a02855703c6f03b1e85c797d7
za357087d98e5b1f45502e45892e5823d6fa4b762932009620038c05d74efcea7c3fdb38901d620
z36515d0824367e48d1bc182335f158c262d396cada6b0ad58add4f945eee634c2dceadbfb5118e
z14969c29a743830a07124bfa78707f3952b96b0db7af7c9ff36f77137d8c490c4f79328328069e
zd7d5280e4f95742c9841340368b9764f0f80413adb175ecfbdf3c40716abca7b8cef6f7fe92ab9
z6bd2453f1aef7f7899c5365c5c83793cacc7795c269413f6cf0dabad14d40e9285afde8c01a47e
zb61893788ec5060288cabde8fb553f21b02eac61ab0b48ad3d54f4d1d76508b22f0c600861b5ce
zcb30ba708be817b1f50f59c0f6fce449203e7355c1be55b662fef3f92ba58243d81537761af8d6
ze27d7864d2dae99372b2b75bacdc0437a4f7e011d68c3487a89759e3625548fcc920ad06471ee7
z2d701aabf726859343208b0a543c73eeff8406febf277e3babff437ec820fb49d6b78e73bc2353
z884917487d35a6cd06d7d73ccff5f05355122888b886d1b7ae29679db6c9d2d7f218ac9728369e
z0ba3297b105b1781345d5dadc1077db50a0833d4730649f7637b2138ee147e4486fe0551f541b8
z43cb1f566ce4a86a39651786521e6c831c0a7a8984a034633d4209a41890c86668029516983a5a
z2a2918caecb85c3a38d21805a4b7e2da92879621bc299fa7b4555f7e1319c222d5509f48164b83
z9f45f9b9fd8b57ff2290408ba1dbf726ff7b13b8cbfde6de453a22cf49001d87d40be9d1294fea
zf8a4e779eeb3a77fd351f4e30844995b607c86e83ed23c87f1e3e643cd626a797a57229093c8a8
zb49b28c85dc6a1ed8378a68ece4f75f7bc8bb425df5a97e4918abebe960a92a0cf021afadd210d
z740e80f431452ce69f128befc87baa75ec9d83b23a4686f48b2cf323daa0a59a3e38084755a6fb
z23946e25fefddc4658c4a11c7e7e0fb4a5c97e53a82d71eac3976e5bf8f2ba284afbf2db6b6670
z8591ebc96dbf81f6c472563caae025b629214a41c49dfe44355a2a0e413d7f3eb61987e524abfa
zfbe09d96faa13efa9a26c93e069b7718b32c51ee39455cb30ea1b434377cda63d50ce713f29cb0
z10f5e5003341f38645727fd0e7212799edd900d19a8309b8cb15d3bda32e6247e4d9bffd062d0e
z110a039f6d797738d528fbcc7f1fb1914e7b324417bef00b0ee9a2fee173a5bb898defdbd380c5
zbde4ecc5f4d2843e2a407d7f35ce3cd0cfe7b5a392c43c70ee96b7b36b3427ec657d86fed6ed46
z39109932d39e895aa0a2c59a8f68184c5689c3d46df4fdec1943af5fc97bbf6d9078bd35d883b8
zf1430630f3021e8e45d34f63761e0e694b3cda21eb35e435e3e4c1e4797ab7af65831076702d7b
z1758800365ea172ab7553255da7f589bcb772be00ad75a9729734f24a659c442376a5e68a8020b
za0d88d4d5e1127c25fff24d05ae79ea47bc8abb6fd636265249815c7a65b0b7a3a65a14afe17d7
z98ef599bb9a3e27c01bf916d196bba576883b3fc73e5d604530a16fe290e470f9f738daca94dd8
z89e7c8107675b6d403082267e1a5851d2c56a2afa97ad8cc5844c9a9dc90def92f95c9c5f0a26d
zdad1e2f02db80b9efef189e9fffc7c528dde6eebb378fefbabfd4dc3ba441025042cb2f8ace984
z8e15cf0113890b3f97b1ecf464416b3eeb1ac71d356755488fbe9a6a29a2bd5a6ab6f0c3ecc91f
z9eba9cac3ba566aabadc3287caa7d60d2d82a7df7a3fc92f8392ddb0618ed4595a4dd66fdceb7c
z1ef16c8b545d36675c7292fd602cb9ad6080404b3d08616ae1aa357915590b3b385b9b06140057
z92cf52f4760ddfc1a69d8665f490b10b4e1cd9b048e5911e37dad9cb116298d3b7127921bc6120
zf394cfd191b44282f9e8d834da37648b0178fa8c13fbd1a4434e12f047eb1969b887b0232a2533
z921ce87469b85e6ce3e0160b5ac525f7c3e190b11030d27581914e982fb7c03b2e9210310cd4f9
z574a921b3b75c115cbb5265b3bdd1ccf07b5a0a63c2bfecf9bc01467c6d432f30338df65c840fe
zbd246dd6b6b866ac3591fdbd6166de31c59e94cb5db6130bcf72a40592ee76b3182cdd416fbae7
z9022841deacd9acc63161152a9bd97eb261b66961c99e4abb7b1c2f16dc6558d682f775e4a6f17
z8cec98721edf6bca989785faca7d35cfb696724a4868e247bc0ed77031f772a1b698718c76a7ad
z73feb8958164a954dd5318884a839be3e256c78cfaff18d19c07693afdf96bfa2d3ed1bf7fcdf5
z48c46fa88b3581d36db87e1e2df5aae0811edfacd04b5ffa2ac4757d9703166d17bf7a35d6572b
z4f6ca57aa50fa76456f239f5311198a5d389fb8b20625798a3b2664325ce29044a18795a5d9530
z67a71adf8ac6a397f0722400feb5de0dcb5f5ca225d019c2110ba8094c9e7a89f6de46883508fd
z2edebe4e9cf0e0f6f769718ebcd2b963a089787b945f9179f3b4fdf1b74510708b4fb92294aa5a
z5e4692ef163bc501f42277af0068f42f397da922ebc5e8559f117b2fedb3134d8da99841863b13
zd30ca98ba5c0475fd772adda0b0e6322cbe56f53907c2f980945a4c59dc1737b75acbfab4af9eb
z03ef996d2aa6bf0404cac2458531655576aafe1dc3fe9d389a282f8eac61c36b6c9e17d0b8e5ba
z47f65386b2606339499444a919d64385d07e2a2e865470b38d365d25729a7395c8594704435aea
zbcd5fd23b3d936b68a03fcef955a5dde0370374e89623ecb73f8f2d794f1929aa05507e5ed0e48
z621a06dfad0e716af6992210348adc36e344f9ac0fabd777055c15c9399a6376d41f170504be21
zbebc5ea1ab43a3d7d6a79483a871b1486a9649c0a9dbd6564573c1c4d4243d062c068ee70313b2
z66f03538df04042a53a5e65bd51d3e9003ed8f8b8c30f79a52c8099cd9d604d8d5582671fb5ede
z9c87f11f96fe77094281bddd881f35479c46ded83e36848084dccc734e7c951485fa795409ee3f
z877310a25faf24a333e26bcb7b5d6a267f6b0aa7740d3b09b64112b56d8374afb542aa59817f2d
z3fa7f7a42efa50afe444449c7059e931bb71ad2ccd8cfac38ce9cf8498922b9078e69c06746156
z309ec37236a76ad9737a8afb220a0d12a23d730dab949968a6f512dd21085de641351533d184d3
z4234b934dce04890e8bd0d8ea6f4238044bbfa311df8653af7addd85dcf31b4820f5e549512ec7
z5a8f3c12bd80aaade03f3c063694231e89b76522f25a8c51ecb002cdb250d170d56a37652f1316
ze9a738205e8114ba6e85d408dc5ebd18a32af4629aa281e7fb20f37188bdd122f8dd84940921d5
zd7a7b162ca39c5d3590c3198f5e6828311b37800b8ddb76a50d0122f42157306c49b4fa06f3d03
z8d35fc87f706ae0b189d943b2a062a0ecfd03953df8538817008dc2f5f7e86601aa96dba91ac71
z32ec90446f81f21a4e05d772c57a595d8f2db50e3da280c5c0de72ac22cec9eda9a4949a5566dd
z7bed8393581e29360ccf5c2c972425bd74ce914842fabc50d7703835f51843f8549477afa13c86
ze40b2bc59f60ec09bc42722218358577bfb43998e4a5bc83fa0e613db95b27e773fac210ecaf13
zc3ca407d963b52356ed4df9102329d1a4bdb74ccd2694eb2e1236390b46803c552818578154a7d
z538817bfb7fa89d3608d1d153f27c8c0100dad6f3842272fe3320305ce92f65618cda6a9f60029
z872f1c8255084d63d308ead523ba9749951a6c63adf572f5a3759b0d35cbadd3a57678b3aa28e0
z8b4ce15b29118d1506d0020a3bd2aa9a514145271236a167af82d7d5a6cdcca12979cf93f4f9ed
zbc5ce5694edfca51ec4f6780e6677044458fe67afc57e3ed6356b3b4118e7007b85a735e054abb
ze58eea09b827bd7c4ff549f8b97d61bcd41bc8389e5ff099b2bc1953977219a683c1b7884b326b
zcf88a679add1bfc8ce63b383691380c1e64c45d210bdc5a4b247407babfb91dee562e966ef54d5
z59014d883c27ad2c18d000c59e3207158f8de9b2efac1867d27ee60ae55e9b8cdbd35ff9c8c4e8
zf96029af42e4082ab117bde105b7dde6db35c0a3f3783a6d46c22dce152f57277480dec1c6e829
z8b3674416165a842a56ef0d739b2f00a010da10f50c2fa9ebaadf2acd10cc2afad7342d284fb98
z0cf14e23b9b04ef11f883187ed7e7f5797626b3d0d47f7763e766e8ca4e396f1aa819016f20c49
z3c58ce73af20d53c0572c226c2b084ffb68212f7e62eddf21033951d10a26b30b03a84912e9a34
zab0de6018c9d7868817feeb5624970f1b16ce0bdacf702510ae432d3cb114e9a0f0e11ae24bbc3
z77f01b6aacee2be15d94584ebe67cc71a7c150125763220d041fc11ba67bc41a4815cd1cd455c9
zbc3d5896ad6cd829f3bc8e1b09c0812698a77f577e839f82767a1d1d84552c34671ba41841d726
z3f02555c4c7f9f6ab1a130e922c23ed1878275fbed0962b6a49560cc0c5f9902cc64bd1f79e195
zd5ffae60fd03e6db9a6e7e299ee1af0728c9f6baecdd7104768fb5e27aacdc9250a1ca620f11e4
z42539259e828140b3844a2640d490c545cf3927153ab5ed2ded70250b7499c71cd4c19fca69c65
z223909e347715dce320e45bacce845e5b1bcef574de3ff8ec9e160b5d4d53891ed79698f64a909
z07fce4f3341b183cbab34c81e01c34b554546b5e6224de16474df42153986353c5c3e6c23b9f32
z79abed4d54bbe81681e98ef4c9145170937b73bbbe983627c0fcac7d8ffe5f003090f459e31120
z3b08e944ae802af50746ecc2a096ca64e7f4933a7a221e20d173702fec167339299aaa42120b01
z7d509ef017bab3276220adf28812dcc8f73d60dd77f8f2e4ee2e499978599c3e4a58834d56652f
zab944d17d19bf15a37b88ddc8f5bceeedeb97c2fb11201ce294d4f57280ed5632f62ea0a5b1181
z34b742928a0f6cb360a4fa95f163dd2b7b8fb04f4b0cdee6bed74d3bac03cf8345203aed5b09a6
z1fc7e06993f5f6afd70b179a8859d38da51228fab0656ac2a1db98e571ed2134183bdc613f0157
zace1928ec4cd7da9379442f5053f3a58cdeea602189583465cd553e07446531ea4590feb9b73b6
z91fc573e449799252e8abbddbf81614ae64c512519a2e5680195206aff3bcd5ffc877bdd6e93f2
zde878e1b11340f9f284b9544531301f80490558456dd25d10d6ab36931d33602dc5285d840a7f9
z5c0c77e249e17adb1dd075cc3facfb263ee83379c8eb95fd77ad8750a9a4559f372a8854bef92a
zf23beee5d79bfef09dfff39c89f82b0d0b038fd103c70ae88b9537434f4f711e94dc943b90da50
z7031be224d29555b0fd72611af53a0ae5ab731178d18076780bfee3c183fcd2fc5f270978de64c
z7064987d3e877115ceff9bd781b467ef538722aee3ca5e828e2c1f187ff3ad20d6e24cb0336c5e
za719bf1af39f10bcc12e290f0258db4b7d5bd7248751a7612e402bafb4541e7b2de4c509b76a81
z73fb0f097cc5a31c8e1431f3d0c02515fe83c34c20c0a3a4e23bed81f91bf6fb3ee036a1bbc011
z854c3a14dc64e0b707a4bebbb6d30e777d26001162c9324aae98603cb08d1f1e2b685e94cbe530
z27c917b0f6ddde2c34e7ec452ba2f2731a20c93c09848eefc41fd277f164acbe865d26d2e109fd
z49c0fc7b66372719379ad68c45375d32238c08016d2399986092940349b4553c3fcc46993d27fe
z31bfc7dedf833278f07245606012636346bc29dc70a014f150166a728f17da215ecf3f025aca23
z5ed7b07ab4912e7cc410bc1cd487c4f877d21065207fd079fe6bdc495eb1b14bcc3d22f53dfed3
zd97dc419754dad876d846f15f1043efd6a746224a48202f3b80cf5c6f27ce1c2920ab8dffb8ea6
z77bae36a4e110c95c05dae2cb9a2daeee6c1df9e4f1937bcc41320750447a4ea09c569f7f5fa6f
z36e9d0971c146ed12a7c7d8fc6758dbebc8c064ba85bfc0957a122999b465695e8c61dd963e74f
zcfc446a3e41bd33f8b84209aa33c772038ec8a8123eeeb5687cb58eb0eb3ba8c8d52502dc68895
z195d87b364f2509095927f90a68f9432c49f3672e8e730f22c073eca2927a74e42ae302bef67ce
zcf9dc961195340939033b2e2eadf12fdb1044fbc1658d6b645cf16314d71720a88a06c7f77d791
zc5d2a2edff89f2a8baec3a07c84936eb5ad9256e700556f596678aad3780a7decc204e93fdaba5
z5878954dcc5f829d865043cbb801d7bb949f04b7afd34d12fc75a0a817dd5e470446eb8b326ae4
z97a9e3e233c24439032a0a3b137f52e473867d5f1f11f46c90fc0fe9ba0764d6325330965213c9
z98fdb58b9fb3fee9f8152953dac8700d4db3dfbd38080553a04e94ad41e8ed788523a84f94c9bf
z4849a30cf6f1eea34b92a04148c39142a6bce81230452d56f563c59826f36693228e27a1fffa89
z5346b15bda33b365a649972442c87f2e779bffb480568daac895a9d4a9e9251fcd3362c88eabf3
z5d33c9b4de4bae0e1aca6aba4e8395980efc272f2563dfdb6b862f3fd2596fc46b8dbec6420704
zb82ce801dae7e2887ee0e7e794f4fe9d1612411d251e543e3eccc86020a520cda78654f5868948
z84062f05941ad12f6945bd86ca2569e2db87cf20a7c8dcbc363b397ae112b92dc8c5eb03bcf8b3
z822b5953347ff09c0455dab2d92a49dd7be8f92c1332f167845bee2edafb93ea2be39fae273937
z11f921f1815cee691c08585a379ee5815686db44a2b05365aec88a22ca4374ddfdca9a17a62243
z5c2875418e1f2353137e8f903630eb3fc0973e6d257ba9a2a0c23b5908b80bd082bd875fd775ac
z2f5e17467be9bdc0c9da2bc164fef775b7ed872fc8d1841e6dcdcd74260ed6171bf1fba21b5d6f
z536b3d4c533a2547a299626bf62e7d3cfd5544e39f9332795d0c0878609ee16ca1874646534166
z8854594b98ab5883bae2a72749c244fc731c38aba9a05714e2843ab0a227bb29009437f4a2455e
zd04e750b57ca9e5ce498053f2a44082a5d69d62a09ed8f01fc4ca9510c3472c68c573473b33a9c
zcccfe04cad9f376b54bf050ade3bbf38ad9dbac209fff99c02e3532efb935964bf655ed0fbfff1
zb14e56bb8c7d24d868846ea46b7810f8317441819801eeef1e5bc29c5046e90fb7f5f6eb5945a7
z9fc1557393265a435d49cd17d15698f67111d75561cc7c4d933f4eb13e19fc4fdb48490cc4517f
z46fa8de4297724145824fe041f156939ca37ecc66614f154915062fcb9d2b64b0ddf8a42efa81e
z243f4a8c9bf9846ba38c8426408d4d8e6d9f26d881c24fd97bef13e5c225d338e29f41639925e5
z20261dc703e460f894ba6b05158f040a41a7742ab9d52c0ca9a530c18d9c69f47f1d04651002ad
zd474816e51cec43850ecbad1684bb758e008e741f7e1f3ea04bf9f259e7c574bd52b33199ec1cb
z8922e27d51e4f99262f90627314633dfdba420d38b64a46eded6ff50f2af8f040b4d1480bf612d
zc5b5fd7b7eba603891b3a3edf3259abbc41c696d0aa415619a340aa11d73504dc1e8c90ce7b05f
z5da1b790a2d825d815badb1a4016b52e1f1a6180f9d9c3a9a10a48ee3f16c55be90603668b3934
zc9c80021669a1baae619bf22e50739ff2f20e4b594959272af1b7446adf82b6a184b04d2f68e08
z5343fc637475462c60c726abafbe358952c9def60d406a8c1a72290b2c19e4fcf8b66bbac77d37
z6dde02454ba042739040906e1cc9b686c4d3367c25c81df05b27b9931f9d8aa045ce9a66a20ce2
z62ea56f0a107d1e3feb88aa637d53ef95363981d7cf6f002b69fe4dd297c2d6a6b58776ff01181
z1963cb5fd86caa7748a2100d866a950bb31d1a794dc5a17847365848b79817e75cfff5621d5c83
z7f88b71f5efeb1f2731a78f66cf096095d6c2121d85b16fbd4430e907c5f5e6d14e4e05ec3160f
z7a2da27a8eadaad7a4e31db45072eb997b384478f5b87102c9a80ef1dc3895c93d752075a5133f
z329af6c461cf3ffb6c186ec6f567f11b1e1c094c586002416231c72cfa9d6b1037e9eba039bbc5
z376823a02b3b89191b6451d363eea5ee85c968fc159a79cbfc98a77b7650668774ebb5301e8e06
z6d7c41f31c9935c359257e8e164936db3dfbbbc60d47a80c168bd896e9732371dcd10c205a0676
z972d7d0fd49661c3bdd7e761e444f3f4a578c82b38a0a719f1124434b57d1c0234181c7543db2d
z1db563105e024eb8e9d23f375fde263c2bf0f5943524d198edf10b668af532433dd86a92b94a5a
zed71be8a88f5203aecbba67dbde19fbd56456bd4ed26d4caedacaca5289b69f90bb5fcd2fdf909
z76dbb6720ff644d35ad1762488bc0199d9f7290de4a33f206217b0ab3c2f9321774270685f2594
z45faca5e859058ebc48c43d5f66ee6649eb11be8a32814734316f657fe0ca3b21e4ece67c5f81d
zb6bfd6a2eb40815ca659d5122dde5bac00eebf6a203d7737112dba03462503c90f87adb8d37c04
zfb19caa9593b428656ed2bca91b3523e1b3b6469fb27a35d55fc57416fe2d44e9f79c2d2d35663
z9da6ce5d019db859d153408211d3fbc21a9d2b94c40548e1c18113b9f8f13e71acb5db4a421d93
z62b985e2c6e3315d154aecc19b613ed7d76a31be01483c9b3582f0929c019bc2453eb4918e090d
z24dab4d6e8805cf652a93675698ffe7881761d57045f0b62d97d38c25c7e799506eab3e4ebdc94
z24a354ee69ed740b8668cc0b893884593a1ce7aacfb73e43deb2cc7a7fac8283faa5db3a61ef6c
z14fc4f57d5cd4f11d951b56deb357605d95f86cb38089024190b29391c30426e4eb82650a8d029
zfb5cab176d681a66e4606206e1e35719d29c2079401cb498ce5f880a10ac670bdfa69a241c78ba
zfdf8b172084ea4ba715f13ba1ad21435869fd1bfdf0cd72abdd4514c38268b8b7f6fa2c872b1dc
z29e2804a9951ed2bf47794ee0542c3435dfd98eb1c3b41d010fc22f51261e4ce2568dcb72a8872
zf10bbd97536ab508f71c4ae40b50d146c9bf8006729d47e1aa0b84c93d6e855224dc2a703b0629
ze759c77e5ae57f977f1b86888a29f0a618f504e1eb39e28422310e8729fbdbf05f46ab8c64c199
z2c7070c94514a800afc2344e6ed62267c457ade3ffd1f8577d7e55bdd9664d943f0698e8e0d212
z7a2a12edffb9e699cb002d4b3cb540b51aa5f0a067bfb53a77022275daac9049812e72f1d3820e
z44b5d8af556a0ed8536b59da1e36acbcaf3d5df40e0b8e8fd46250eaf5a12f6ec4e5a90ef4872a
zfa89da1f57fd2e6f8e4231bcf046f2aa648702c33c79f54c0e123de3b173edb5f0ec7560068647
z052dd54118bed581a05ce9990aec7ced00ac6e027677e4b46a3f3bf31ba6b06b5a12219f91ecfe
z67bb47968d8a62a8f9099df8399c54cce85581048b1307422954c7229226f80091958ca5bc3b27
z1e4a53797f6315a0cdd3d038f57131f6b04988fd997bf4ba5a809a391304ceeab0a2d2ee3a08ac
z390f856e094767c914e94acb71c22273de05a063bd263bc657d9e2412c9b5c96a9cffc5f0ec56a
z1850405871f4131f223d696c9b470265425f588ab8b6eea9fcdb953ccacaa730ab36c9dcf91f0f
z1424806be86270e9e87bf6af1de0e1c7776752de7173d260fe3496f02b2b8abbe040da140f2126
zdec68f1d4c73a3c5a1277c75490fafc77784ce6b0dcc85ede0310eec54dbbd8a36175cbb3abcb5
zaa0902576c72e588aaaac616cfa5eb64ab6bb9d820cb05f346dd10bbf223ac242d2d6e8d4e69df
z362ef758d38759a140cc5fdc4bcc567a53eeec4a5bccd0fe64a180b6ea13c1e8afd63e61ecc923
z556f34804ea024e5da15a7039219ce486c8ba374cae887feb3db6b521d115cea752f71ee453984
zeff8fbb2d3779bb5fec6d9a6dd13b9b7a0e840eecfea834e4e45481fb34ece9cce8baf360ed278
z90bae6563dcaf6c78df3217974d2d72afe71fbc853bbc6834a17c2bec6b915da2a68961f83f2b8
z4910239c0a0007e0047ac06d7eec2c4d1ffaa4cf8e9b7406b08018c30758c93a90eee5b8f31b61
za794a6a886d982f365a6195ae6c44a0b45f66c1a3ed3bdab92f82417502120e10f36b398d4fb0e
z0033c1c7900c9cbd5055e12e4d46e7dc1da60fc29e0627bae2962138c5fe18580e4c631f174f0f
z6fccb8ba7b67dcefbd0a4e673df459286bcd6f8d383fb20c5297f7ec217fcb471f72252ed5de61
ze759c48f8e982b1efe005e967d25ac39d05ff71ad78dce39fecd7267751f3362b05d6e28c401e1
zb028bbaf3b39a3b9b08b4034fcecd95fe56fbb1e68aa66078e891ac45402e0295b72cb60b075af
zda5c48f8bc6d960daa4b53620526a9d10616e7f6a7dea48c0229e804af379f675789e726772c16
z4c270e11fe56f5c03906535924daf231ac37fdc301adf2f7752981c5dddcd27782d9499f9847be
z1e4d1937c8b68453be7770d97b2348af1739c0d256133d75f8ac398c3533b99ab1c3169d10afec
z2255b1016d518d17a5cb2fdc2048ddae9494ee2c55d8a5d931988313264b16cbbf8f4d272ca364
za7a3897f39a8bdae40e000d22908bd4a8331a6f06235ebe973cb4e7556abb6e83433c28654b857
z93997ad4f0fc7c5bba238c09b3400d79f466332279fd2a6f0f48b465c16a034238f0696fcdc9b7
ze4532c5279e4acc2ab7557192a83c13f9eae9bbad5136b2a471c75d8fdd210a8f7abfbf3fa8b0c
za64afe74213751a62cdb92272a40b378a1241fa9ada879a1db34ee60e18c1791df88e8386de04e
zc8e0dd4e5b3824a06c6790bc29feabe25aa6ceee7d1e116f77c4fe97ad9884ad0373c652a194cc
z2b235cd000c501e2b49a8ec848713fedfda543e494be8e8655d511d88bfe2531d17857ce62934b
z3dc137fa5db3af79c4194facf2213757dd1e32e26636c6cef59a3326c473f49bfaa683742e4773
z26cf254ab2e80cb75e9c85eebc997e5a12a86193226433176be3b6ca9d45cd62b0fe9599481c76
z1b69e047138e619e7b5e92cfd96a99aedb911fcbd2a99778619f9af5f09719b116aca2ade0ecf0
zbf946208f6fa355db552e97896980a16baa9663fc526acd14eadf6f4ab99d373baa5ef09daca04
zb374bff2d8dc3f7b1b38096d1b080a181fa506552a49807ad4770d0f303232a3f99d584db0af1f
z65c08a0ca75b4bc99bd40eb23d026f35b74ef0925ab01faea1c48c77b1c9bb50b688e1b8e1142e
z4fceb74ea0a5577118fb372790f2d8b165a5aa7c09892d8df670ec138d87a6731cc6273135cfd9
z2b2f5094ab4de5d6de07998109b4185dfef16c4ec9bbd298e1c40c9f9f882883497461ea14ad34
ze3aa1eafb982bdc8da884d1252c64b5fafd877ea74da86ebfec6febbe13e2f88ab3a780c47a93a
z411ddb010117a56384fdf5220de12c7d6a98443525145e21dba93c191d61a15737a90801a1438f
ze66fa46f86087b83ed343fa260f1325ca440c99e292a432ddb9500ca8ee98e115a31e1c286c70a
ze5ec680557142b9052b8e974bf32b6a3cc5b9911f326ba90f5974c022b8f372a916e9623b50c51
z5afc8344715cb1dfdc56063cfcad1cf2fe1039d4eb61027566c5f20e16e4fc8bc828aba4d21c5a
za612549dcaebdaa28069d315bc52f4cf6cc66469fda2e3955655e1a46b53b482b696fe4e8a3cff
zf7f2f0128e61d3dadf68275c97bf4f43ca15e8967da9a52f721da820b5dfdc11b74badd280a52e
z888905636bb1e088d9b35d76c77ff92c8274f07ba9c1f935b7e862b628a99f4fb4006faed51fe6
z6d577855eb2e90b38c2a55e25eba7b0e981282741952ceb4dad20de127d1ec624e6a65d30b4bb3
z06506986ca5d8e2607c09ded829885eda86f362a01889239de899d5fc79549afb039660d5c8547
z7317e91f793f243d0b0a2c69efb15152926694c030386252fe8f2191b6615fbad40f4f345bb35d
z85c9e3dc2a601a1a6462b0271799257cf342803e596d5227b77ebefaa198848c992b97654f2155
z94934bd4c4b0f08131cfa690991a8627c0edd429ba8814b091f47ec2118fceca8af22a279fa174
z6ff28d0832faae6fe238fe7549a6d428d8944189e73457e9c55de3e86f4e9a9f0f4335e7f2668d
z2f91cee5efbdcef4837ac6e0f577c2e82ecad1ccea72fed320e139171cbecdcfc4706e84743b4d
z4989c969f9680631c831ed1908166e1282d0c22ed0b44f3ea4ae0295b8ee06cc94dc92f4f7f37e
z46b59ad3fb0954ce363b788d95942e7ab5f298f7395292c3c16b5bd926b94744b10fe6af8ede75
zb51e199a21c3d5ef8f0bc6ab3ee7032748b49568d5f2b5e4317333d1364f6d440ec1c9b83d94ef
za22add8a131b6a2dc61aa97edad54ff94e3956022622bffc336a47f115a916bf93efced2bb4bf8
z38789c4cf0c47b2293ed32c937540ee8070cef208bd065d82788385a15f0959e3d48a433599b63
z0088b6b9fdcdab0cd314cf4a20b9a6285d1b97b22ffcd06a327c06b5dcad4a249df18bf1bfef24
zf0102781ceebd8882497842e75773cf11a468ddaf1bda5877e7332ef18692c26ec78c5208d62fe
z7e05c9c8a296f99bf707b1b04b86d2e13405f007c61d7e4690ac9a5fabed8cc1e2bae78a9ec49b
zf930dd3142141ddd5579d8ca941a119c16886e42cd518d80a412e4a36fc56d3f0e517fd2df402a
z90700a470ae2f9831dc4136b31280d83e880685d537156e5f82bf3ef4993541dc31b50e8b81f48
zef92fed8e0253593b0248d1427f881e17daf39ea36e9a140f7a7c4ff348416987d69f841576557
z95d24abba583af6b1153f928aabfb2aaeda9898ea2c25d1b7a179ce40df84a4a2fad28db5d79aa
za1fabea9140e53814f7be2b52f9c2ecf0fa532c58393c9d37ef70a55d04282a9e4eb3037032c7a
z8393a31efae0e7d6d9658e12f34a3baf98a12d3b829704d667fe201e4df7d5292fae4fe1e545c5
zc884a991d78f354c5e9dbc97d790b7663c7e371e134b8db48576a1f91b51f945c3820659612ee6
z96184550933ba0474545eef165073ea7ee68ef48d0ab7e429fe8086e3be7901fbad0843fd9bc01
z2773fa72b40840330663c26b88c03069235eca7233507c3fba599aa25d676c4234a90202eba4ff
zf974c19427abe6968cc409b6c29b44032dc427a9e9b6f80ac05c0698c4ca11395bb42940b6480f
z1051ee406f5b58721bb631c5b22f803d004cc072375cf19ad34b563d8f3e70e40da22e9d92c9b5
z0db0923760e377e3bbda3e996ebbf5fc397a39b0f2b3781069d8e30b1168105d58528c7754eb02
z34c3499390afa28273c0ab7ca5ed6fcf90d750dd1da46b47580846b447815c5633eee7fffcf2aa
z1d643d0df1987115961b15ef7bf40f390e85b1b5537eee34df133e251b7c0169f8ab3d6c271c37
zd165adadcf2f01ed1cf4e2c74ca672348ff58428a844ff15dc45c2e0ac55de910cca5bb77dcd41
z88b595253be00b451bf27c9837d5002f921c01570ae09a899aedb1518d2ce2fcf67411cde68582
zfeecf0e655da0ebe654a4f99976cf9a7ee16eb524266b565a26b7c9d85ec140dcdf9f6d55a3077
z9d6b9fcc86bbeacf750062f9c484939f3aefb908061629dba54fadcea74a5fcc51c3ff416dfaa5
zb309648d928eb3de087859e79d5cf6ed8d7b4c50e8dd488cd0df489eb25a1b9a25b2ea15e3c0e6
z2fb084bd077b8dd72cd41f3005362d251e1d900bdafd9b96778e3773df67fe36d60ae8dae7b7f1
z0d66352524f78f9886e9ddc89f0d9e8c830a216078e460a34246edc9fa68a061411c6262a24e3a
z0d80f273ad34259ecd4f920dea0ae0506f31489f194e3262f99e82b999260b61078a7deaa34894
z802bae80df479c4d979849631f267b08e67d59a6e85c46b6e57dc5f4e1c4d280031bc350b0df89
z4b5e8a278c94e733b063ad3553ec2f2c406c7b4e13e06ca8c25ffacc7519279975b15982111123
zd1607afdf80364109ba0f45ad6d17ace91b94909cd118e1b622dae649d6b19d058d8e8642cd401
z058dee12827e7fd01cf7944e52a4385d9ed7d2a074a45d43129605cceecbd9ac78c0b0f429c7d2
z367d2c143db67a3a1733765a8dc4703ded95bc4980cb43b2b25781de133c742c27300eda0df4e9
z1f8173427b06d35949bd9aeceb7f3ca39e91885b9ecdb7cbf9341832c4cb848667296a5ee79259
z93ae1f7071cefb5d92eeaf906ffac8eb02c2e4136d7a0af4499624e266a0b494bbe989b7e6d459
zd2d335e2a4a3f2e41fc6245ee5aa2b215769adaea6248d33da7962ab70d962f68dbb6fefbd5eb8
z716ce74e523883370cf7ff93e8b63c306b09b8f3a3724b0f4892e975821518c20496d3ec8bff2e
zff95645a94ebeb89fbbeb02fe916d40fa777816918f4fe63c10bc91a5c64e3848f066a62da6fe2
z530a60ffbd2db3169d040ca9658387a59c82e2053383fc6a072b2c947a07b2724a1c6c85f04229
zc6b0bff96c7f86091b9851057697d06698d658ab894b279f948b4db0bc94c9b18fe7914f6d738e
z1ccc8d74d2abfd1b0737e6809aa023b165d7cc8c12e939d7d18327f13de722bc79d38d8181f8bb
z2c4c54a001050dd2e4e883b1a142050c52c62ddf351fa1bfa41fff961009385c0ce8930f23f909
zaa19bec54d68fef486b50bd0a478def376429088b498590a7fb49773b62720ec585fd09049d58e
zb8ad6b9445401c7f2fd6912c5af144c9815a72f6d1d6192d85197090168a914d77f986e96aa3ee
z311feeb4ea0c4045628afdec346a4ef727945d9af0b26fc15674ab8f5783c1f8364878be54e83d
z71a5b518c809175e46979c10ff67ec36c45d14510944a342866b2f4583d4ba74f9976c06fcad8b
za8621d1cdccf0756b029b58bbb24c0a952f05a5fc0b6e86f820477aa5d0753dcb451ce5db64e44
z807f9a367b18ad401a8f1540feb2ea1ad0758dc126eca4992357623ba0bca97429f0596bffd0dc
z7550dcc28672c61988b10d08653b09d27e33e77ecf514b2d418cab115b55104f7a2d9194687e22
zb84e69cafeec08eaf7125353a33358941249adb8dd35a24999982ac26231bc16d467f48730ab64
z5eb7e93ddfe382d5cacac838123635a1b66c106e529b465555c019cf2fd7964bb90c85364b791d
za9e7cdf34ad862c9c9a9befaab02852e6f742bc7ad513e546ed817d9fd9f1a2ae24223a89b09e5
zabd642fb1e65e61095f88578348fb44a7df9733f4398258be67edf7f5819c8a94b73d13685773f
ze52552e29386de0af79f25e2a4b7f7fc249f4c039a13676563e848ace48522782116d0e6e354b7
zc8ca68933db46700cf5c9f126ae710407a932c64df0dbf16ed79b569a3fadc1180ecd033c7cd32
z3378df5831a9ff562e3326c0ffa665f36a0dbfcfc918d9e1f58b9e3e6e116951b84e9fdce80872
z7f900d3e90698d4bce34e89ab94d88eb4e00f7c6fe4943d67bd1aad20049422ec11ab071e3cd04
z15ef701600bc1a99cc2b46e8b413f9d5204e779d8992c0c62cbfcb276a10b3e3f388f4db9c6066
ze91b0adddf7b8058a7f135759b304dc8d030decca8d47647712f96812059c989e02dd3f61d9a3a
z67ed8f102cc5097cc979f447dd361303c7e598f2a5acd65cfd4ed9a1a9952717960b113350c4d6
z73b09be4c9202889a8ce83a37d577eab69009b1d7a5377a72e14943ea0cd9a3dd6011865681605
z540df7d96f04a8ec6f9a4ad7be9dc9e3c298e24e8b896c5c3fa155db232649ee78c2df6afc7f95
z55d3a8afb79fb8ca17beda1116c0fc2b6d65655e7084507e04d119c79798abb5852558f6e5fab2
z6616ad1a0f712f3594283ea79c5a12d2df504f5caa68c7b92464613cfeff460e19320486e86e56
z73010c2dfbb9973ff2f26f71dcc3c8a7d2dbbb1ae0c578251b9275797b78de486db79ca25ade4a
zb515b1388c392146b249dce4b328ddfba42ccddd640b27b6dbd930ab69b50819841ea9cf4949aa
z65c6d6f7a04171709315802bf2010441c6b48d3734be375b7090e18805b696e07d9543cb2c3178
z96d416a8e1119063669412c95456196fd058f7fc667e6755927355cd18b3947efa5ceae1b2f9c5
z4910ff0003af60c28fed57e752339db7eec40c59035dc7592af1b74e9a080423b717eb24aaed34
z9e58cfe3c93111f44478612ba1e267c64b436bb33ae1d41325543365d1c45758960d58199d4d0b
zac809822eb1c45bc4a5a4a28c619c0f31044af54302bf275abbc6678e1f485c8b7c1abae30555d
z4ea77f1eaf4c3a4c5c037e8a705202a9b2e4fc25fe3af676ce761239a115a7a5eac53af3641546
z1af7336b96eabc25a2d0cf5737945ea8354becc28b7d90a0b8b38ce89835e57e9da8394c075ae3
z690ef4cac3727f6f694f388c42c7e0e14556e59070b66de984fd58710caa237d676ba85647c1a4
zeb4953f5664f124feb032f4ed73368ee4879a43b42a687d177d861315eda23e2067ef55337b5d5
z3536bb296097cb7d38006ff28d6dc22d168491f9535f811bc53cff1cfe245235710b6910bd440d
z68e23c36ed5f4fc870c09d8d14c90997be20297073c670fb45d128114bfb350f98e58372a2df0e
z35186753f0e09dc167bd857183c4f1529be6dbafecbc0a02bba769463dfce9cf2f7de7d82c7830
zb4a803343f871e14b8438e3ba11efcb577db5a5ec5a1bb9697fb31f0d0d84ee11ea1ca6a9fb1e5
z13d371ab4cffa338c9f78e9c9313b8368beeda7f358085c9ba943a17c72a70297dada14a27184c
z32b3cb73a8a162d2225e5aebfb4f1fdf55b588003a6182aa30df0df577150d7e03fb7d275628d2
z86580b857e2cfb3fa5c5b73ca467dcdfd7f358033bb846f7a0dc283299b01ef50306a9eeaf21b6
z970be5dd9ff66475735795763708bc5d62944b7015ff357a798357d438df3ccd42362e541ff8c5
z9506359703504c44f036d004a68558632fb82e09ac28cdb18284a8ceb4e9efdf1668f2ea9d6340
z20c9bf8eadfc7037440d06511a118e05134debe0387bb3b3114c54a455559589c5bc1cdfd3b456
z8e877f22898f4ecfe44b8d867f31dea2a357167661b68f6ac3dcb6e187308a0dec1a485b9d9a94
z5bb74b3764116c3c4a7df8d2825b790137b42d026c0e5535588ab8a036aa114135d42b45251395
z5332bc315ea630477dcc70d5425741138bfed98d1f602ad32b1664cbce84274267396cc4162ce4
z4a7cf4a4a5e004a90e97f9f6187d89a5118e72c9e3b421a37b64028ce496ade2e12b9433deecb1
z9ffbd0f60743e61a1a6f739737a692274a6931d2e69782f1c5975e59e1aa9e848b0057ecc8b4bf
z1e57c1e3442fd9230c0d921291b23e85eedee1f298c5cccbe6930926fbe3700c4908d36fde4840
z5624e6498d0e6f4ebebd7d095954e95d0d1090ed16f2e534c617a4c0a85c7ca3056ae04bd5b69c
z9a0ce26570be1f359b9bf523ff18c94df54ae9adf9b0da4746e179b8f82fc7f3b376bd0069f007
zd81be5eb4c5f0d80d7f007ea8792d7159609059619a0c730a7f1a417225372c0de051b412b77f0
z979e0e332725e13066aa197e29e9c54ed1093c1645c6bae318457f65fbcd59fc2b01b35ec113be
zfebf051d355164b6c745bc0d658dfa7206473171ef00d096645f7e14a98c9205c3a60846c7f9f9
z044266a097aa3870fa6de4b5404fcf1cde49ba6de372c04f8774a3e3282fd70e40ba16e7dd1bbe
z7e38a464601f1100dc6f2a556b6832806129235ba45ad69880322f1920afbe160cd7d705512d8e
z3d2ea3e1ed74efc32b94670496407a0afead6060ae049df697d0eb3556a6dccf179b69eacb5d4e
z1b8748ce8af040712e81d218f29b87d80cfbc268a54a7ef8e54bebbbc72808ed95d0f237629920
z5000c6a5a268765e2c647abb90d18614f3d933a571e6dca68b9aa9fa0b9ad1fbddd3fc500b7ec7
z063f7079a3525f17ccc88905b06ea65535c4dc39b965139414055a770182141be88feb4c264a1d
z28b94bbbe5d3370a9458f1a4ed63393422c4f7ca204e3253d0ec0166b996d61e829fb5955836ef
ze840e95db7f5af35362794fb3aa961ff3e65ebc421eb55a61656189281d4cf218b548db2cb470b
zf2adc4145687af57e6c10cd930ea6009787ce005ca44621a05dab3e7bf7ac6341222f4b191e354
z71b99613aa86884efc45074cc9bcf2830e8e97dc15e9c67a6cf7e36a660e50eee359de6e5fc527
z02fc997c169e1306bc736095942710271ff828bfdfb7ebdc0635fcb1281551c6c7a57be8300138
z3e6d734d6cec34fd549fb57d26b31017fe1705fd9df9b7af73c8f87a2083a732419d35fc2af5b5
z6b5fd0907cd26cbfc0355b8b26f1bff2f637bc0a93c0cf784e5f10f0bfb6c3578cf93b4805c473
zf9324a5704b767d864b026cf842d365f568d4b473fe24d4c6e71206405006e1e793f16fd975f65
z43160690954aa50b16decfbd9cd77c28cf71f3a0b7458e085ecfe9534c711549dae9a904cd8ea2
za81186d9eef981820bd3b08320eeb05ff544465df9b7d11637bd87dd75e0f8c6fa3e100e6aadd1
zd4717d721d90c5ff4249a1f5da3af77ceef65ebc4f15448f595d81377ca9830c01225c883d156f
z05e534fc6bd3b872e7533db6c786379c6468b7f4678f8998e2c4a002a9cb3dbfb35efb90440618
zfb0d82fe1b26fde26bf10ecbea9e743f1459bcd49f624cd87abc8264e4df7616f10b326593950e
z472838c3c9d2e5c1a74d6a3c4f3cacdfd4ef035558b9a556bf0c1eaf65a4e997194f76f6a29b0c
zda0d23166e2f6a145eb0141572fac151b2c95903f4d9d0211cbda0ff68c810a03462e4146591fe
z30d4977adaee26815fa6dcab6391d7dd6c0b16bc5d8994ebe05e36bc443c86de3b0d9cfae08441
zb0822c1bdc027c67b0d1e91c6a7930a45e2798b9c2db9cbf96852bf5406e4763b4b5b684045f41
z4ee12983b66f8ffb803ef44a6baac8e313f5252ae0002be4601d30eb716ad04d65bd1c50767c8d
zd7d7db34af665ec3aeb950bb84d1313bf32e81ee6d9433e1a1386cdf7cff2703b840509fb89fb6
z5c99c860d3717a810e511fb4075d055a33d9526e823bd129231f2cab063556068c91f63419768f
zadd2de55ef7e270e1104ec55121fd2641f3d688be8f4ac82c8eb4a25314cf76681a0d3ad4a39d0
z2987bb330a64da175461684904ea05094030095899a9ab183c782575a37f61ce11160706ac3e38
z43d51c77b0e0079f381c253a0ab2be22ff3230df365430645baefcb900ffdd7527ed5b388c1dbf
z0a36c61e83043ad434bbd880d6d2562a150b0ddd03edb4552d33efff65fe55d9a53114fbd19bb3
z13f21f9d6a8a56953ad9350c75e3126c42104c8447a01c164fe6dfdf6c7f0e342161ff7612f0df
zd058c93001b5f188a4d6c06cb913d0e58af24ffb9e59ea10848d5891e1a9703ea3d46b5a9eef6f
zc7c319a510e674646269c007da84aa31d523f41c4ef7adc351e61367adcfe9535e54a49ea6d1dc
zff2bfdec3d6bf9aa10a7816fc981e3d8f890e7bd45eca16a994bd7299f812a7576db4b8924c640
zc92820cc77fe3bb9df2d7c3662b33c061668adb01e232eee563417ac5701674647769a8ab24c2e
z26a2b8da6c364d832cfca54f50a9f1cabf94456220eea578c94758c61ea3656ae991e55e330bc0
z399a9dee1089a6f6a1c9d330315937541a576f72d6a835d82678c1e2f13276a890b5790cd1ba6e
z81c08405e8151bec091090fab8a49e66cd8fe3e47684c9d508eee6b46c21526a2048bc3868b142
z3bdd36b46d99ac8752348881dd4146fe01170d384fe851ffdfa3610650646d634f205a7e005751
z3bdc2be200ad4ee90498aa614be0cfc78ec19206148a05582317225ced8bdd595f068b8441df0b
z798ebe74f322dc299f0e48b8b340d993d00ef8775d82ff3c4b305bbc2b0f0c70624f0c9db52788
z703dc3b2c34d7a507f8882dc6b8fdccf67483a0b4b2831b3af66e128b3d218d5f03309c9e961a3
z1befcd3c69f5e6269161b62ccfb7a66b33d899c96ba40eb721c2928fce8fc525765819ebc5860b
z764d7dfa943e2579e9a509520565adc405be114e0f106de2163eba560680f2d490f435b6f21fc3
z741c4d0da8fb7fe0d915868ccb83d04c8ab608be99b1c19f29b1b549448c762e795d921cd0e719
zfaf5c1ccd4bb1e6218793a74473662ccc7b55915528f6ef183011d4da58ae71e74cdd3739838c5
za62033aac1ce817da85430f78af69e601ee12dd33946d074a3e55d6f4a2385b6fec75f8275fda5
zb751099bca560b8267115f99de66be540699a04b8009793853cf68e5ab08af6b198739bf33c550
ze1eff5af1415b768ddf9b2977899e3db4fe111440f43978e943b9b51b4c9c292dc8f44c29a39b5
z5f07f9a61e0ac3e9c716133b5b10e0c517868ff5edc8414f8211c8797a5a5b5e4ebf5b5192bcc8
z22b8814ea40a01d78f4cdb7765df2fc553aac15f6f697812b892537af6baf5465b45d4aa52c75d
z494aa7283dcac2d6cde1a5ba56b9e2e4d49efc2ce3b21731509fe81ee75d5fc6fb095500ebad75
zd13dc8eff615ccc09218e93457671e0590fbb7d339a22862cb9499beb03bf021d596b635f95523
zcb58e159eec0c94e4e63104db605d2547e61bb38402489622aeae000ca9b11fc3cbddac8c47ae6
z90adec3ee24f1d72e68009e51bfd035c76052882cc8b0120159f1545654afaa09707f0d79f184d
z40a20766435acfcef6e85afc7ece40c02968d399b3c6c5875e504d1bdc6bb894631ec611db976e
z2e71d40934f214d914bc7332f5009c4bed0b01e1aab6d98a49f0c3ad91ec16cdd2a2d87dd49892
zb2fccc700a254f1a9123162989f79b375dd905539c6b43ec0b0b2c8fa46874369dcdd99d11ebf8
z14c1d791133046f92aabc4f0ce62e6b163d5d8fb1169d344b690228c196de0a47c3570d82cb690
ze47eceed315de892c44aea7b49e934d55dd309e07507b25b7ef4818baf601e8482785e29d1d185
z74cf3311a838d6bec58d2de35c63b2967d9a07454949ab45ff9506b2ba20a80a778ca05d125055
zeacba01970f7387d852344cf0338b795157c0fe5817aa2b684d9dbb4d6bc6e3d37761b27221084
z7c3568fc4eaae303a14ef967721e76083cebed99421a554ef4572154fcbbb84211d958a6b37aeb
zc89c56bc813052314b67c03c91b7a67538806df747553360d30309b74cc0060fab2e989fbeaf41
z3ab38e4db5402a183da2196e01a98c02f8e009d70e1880b9595e4a2b0ba76a01513708660a1961
zc37ee0bcd055a3d166c39f6b1fd35519dd666624f6972ce84ac1c209d747a7f798476f215c30d2
z4b57beddceb9d6d16f2e765fd227457ade0df01edb6b0834f62102ee87c74abd0854fe566edd50
z003f204c58e08d34a29081ac9c3a5a449f0b10a2f464f3a4781359a5485e819d5d88315ef3ca9a
z9a13c4188be83dabbf7b58e7958ee6089ab0c2367d8cfaad2dbd1de005e866ca0ca23d6358926e
zde62a328d58adf1b32f9000ca7dc464c6d9f2afb159c7160f2f1183e2543b726df1b34b55f333c
z8d79534210bf2ca4c1cf6624fbffb14c99b3165475fb2f08fb13d522bf09bf3c6e4903798c555a
zd07ea5c7a5ead98241702443e6f905687864d436d4fb1f38e6ecee04d00e1b54551e12dadadfbc
z7c1ae4d98fadeb2e61ca2c20efa5b65e57ea84e9467d31b6995c01f9795736876849791559fe81
z027a9d85a634470c67ac96a470e8a0fa9c7540d148a0fac6478e624200a4166b4cc16ba3f52ee5
z69cb8a15ddce4fc7f4ca98fa2b5ed9cdac36a5c7133a9cbd1ef2d5b17e5cd9919bbd331191541b
zaeef84f0c10287c07a90fca97a908567cd244f9c4453d63455c1bd37d5975b994008fd50359132
z5117302be3fc4e5bbcf31081f8ab74e85009c0ad2875259a51207968e8249ba51328368f419939
z1c132f46861f7d77e169f5bca8a15b84ee964c47d6db9d9fe6a0fb95b0a04f202a6a8c6da6103d
z0c3703e833df6fb2b1c41b4d23d0f38e445c0f5427460c39231b3ed7dec7167eebfba4104200a3
zb5093d3e37a246b840181d6983104744100805d480a039ec81e633cc80b56a01b152638f6bfada
z53f6e75712549ad084cad5def92b9b35205b612f4a3a510e92fc0a29e0e3061cfa78acc3b617fc
zf1325f3c03f23d92284f9896055998c8b13b9f414f83a92bcc6f910cdd440534be7c092c2cca69
z1e474a3ff23f7dcf907e91e7540a1239580971f75ae4f5ef373f8d811b42006435484559e1dd19
zc49f7a10ca12587d8ce7ee51a0849f605ccb8a0d67e2402d7fe21c4e7f354c3e33bcec900a5617
z413f902cf7a361b3698292c3c864d19f68ccbaf32e201165a9325cb22cff9847a9fbaea0374666
z86ed4270c3f2c496f7aef4ee3eeaaaf999f6403fa2cb4e5b0c7c0af632e25e92f1ae4b10a045f4
z1ff717975da9802e78b2d7d63a6e437485ec7e0823e1b7cba6a807baeb9d4686ad1bae68356bf0
z3ef80a382fed208b88ba72baecd01dd38da2977a06eb93c81f137e7e205f48593df45651157a12
z5f37673e4ce9f15e7d9e14e6acb369fd4c7b81c854dfb275f17466476aefee2301efdc1644686f
z62de252a6d369a3f352e064d69565f2ff98929c79798f379052ef2e4a6ddd5486dcbf4ddc10601
zb3e497b179b25de536ce0bd444d801a90226aa879f8285c0e201b87ca8b81ef7f80949a1ac3baf
z86f0860f2adfb89bcb35b5146e15d781db9e17ea0745e0332cb8c19930f33ed71f283d1e6922ca
z543ed6b0069379370e2d43a3f698c80843b2c75e981a768ce6cbc60ef2a91d2fa3eaf9cf5befca
z23f7c2fcae737c3f9dd783fc8afd2935e892154f850819732c38babdfa5d0cd0b048cc7aba8da7
zbcf06b8fff8a3cc26dc1534a488eb82c9cd05693f5ceef4227853fd500924d581a5869069e5789
z492eb41a6cbee31c410bdc1becc73ca9b45797e952af44e507eb6f47b21ac974b33a52bb5f18b8
z4b2bc7024245ea733dd15a8b9f587b26a4dd469974468d1ea1ed6dc7ba198d65c9a3e7ab7d0c04
z626c79e0994eed6f33a188872009d59032704c94f2ada2a80a540ead7e69407732ce0cd38aad6a
ze7c7634414ad27695a41e6f9871b8b31a8db342780f6cd1eb6b33f08c76220dc341a22b95b9cc3
za42309dd5398887de99e79021e4e42bb026eb12397b03a2755b0c9e373e590ac31c05dc45e3e57
z1a19e4f983bc5c0218edccd8d83946037d3fb52f592ad09c32befa4f4b32f9dc028ee66ee80150
ze85c15da0632c0ae3b8c6928ea52408a8381ed9d514778541a350bbf771ed1e1d6f309ecdb550a
zfe04c3fff80e7be702070b59be229559fe2c73660b27a231cd5a3591e05d25a523f93f166cdfb8
z7a0c74250ac1088c66341a844eb29371e74febe30ff83ad9895e6c2414153ce9851ceb70e73125
z51a47659093b4ec083a6f64a807d73cef10428101347659aabe2ffd1a092d901a00aca8eead613
z8d5300ae43bf78ab75d974bae2cf0b304384b33049a1dd4e7fcd915b86bd47fd02d866b6c73446
zf36bebc2c7ab311db742116f6a41efa11dca148ea744391ee2c283a486233d04a3407eba9a3165
z3fc78da71d4f057bb61f0fe820d51a91629ac39a2543d5d0dc63229dd861b76044b2f54f58e37e
z883ff7bf914f360db3d19f8b6511f1d1ef685380a9b3566c33056d6d1e7817c2a28b166443a666
z28ee221632ca9a526be48cdd97890f5805dcbdd6bc9f3f50777b796f86ce54d9e4a544e8ff47bb
zaeff444060ad4f3646708855e57b5c1ab0e27f5d3186f92d0bb105b839cbd8766b887c1f2140cd
zc3463334aaa15463130ba360d9c2445790d46812736178353de67dbf84c85e3fb17d83cb383cae
z724fe0b3e7b9d4feb191822e37b46039de7989663dce7b709b602ce331648cb8cd66e31c991c88
z037ed9f50f6786dc9361055b4a7398b7e5b9dbf3c7d6760487d9c968bedb540ba236aed848f0b2
zfbe97b12e06c448856d22fc4d64077d0d05729a1dd13c51dfc19622b192e3cb5fad512a97b23d8
z6f48f77943bc0dbf6b7b79b39d20b0f3b983ccda6be7b9a39cdf367d72b1cddf57bc94c8be6e94
z32cd9e6c90c3871407d440829451452e8bbef3b0286b7ddcf9698cb172d34ce7a5fe7f2d7cf64d
z2969fdf800619b3c40b47d0cd5a8b66dbdcb1bbf5ca0b2db6d3a15c09e7aaa2194321dcca1af8e
z930d525019c8c61b74f28e3d39026839e978f5ac806a08e214e537b32cc3552adaf4beb5adebf9
z14619888bd4d063d359bbf01d1ddb325b71712db503f30258e2402e57afea7c17f975e9aaa1fe2
z9ab9e40b580bc19cb5f2cf2f2ff95e58523311dd330179ac39a7862d288f413a1e1d5daab00e27
z98c3c9631b01d73732593e73f55ce6aec8f8fa55b2128f87205e8b69e0f7e0ea46cc00d062d442
zd47e0b15367e99c233be05dd584df48c97356bc3ad25aba774311e9b51c02bdf53d6631899ca20
zc870bbfa8f227c789cf99fd8556afc6ceb970e8e7ec4df638cb01d70f29299dd8bb30273d7d896
z3f0fb2bd3a035f94eba82379e4869982160d93be0442c39c52e202b8101c91c850e61f967c1802
za17c5eed414fb4d2bbf8e82fa869eee1793fe1e7599ed9044c2cd212225e83e2312777adb7db99
zdeaa8ff3f79634f5022e4771d91cfb4c59559be8da741cefce422381ad8a8bd7523dc0e5342bcc
z49b021c645daa0365a01702d7169b0f0a1510880b5145ebca8c68591c13282c5232b8f00d02fcc
z4796ae0a71041b48d8262faf3295ff2b4a0ef4f0adbd16c16f9e216012e1ff14eaf16f5955d292
zf3f8988b9ad7759a030e7eb8e068bf218e49c4a33c6835ede786a3135977f74037ba3be7db8c0c
z27be61ef6ee034713cee1d9dc2ada7f47ca732c8223b8c6d8ddda297ee7e91a93f56582f24fab9
z13e35cf7ada0a93505d45785cc81f1a6fdb7c5978069fd7eaca15b63c397147de78090921d693a
zc524ea575289d877ec39e534b76325fb344d3110589d4bd576c974dc5dd4cfaed24c3835110cda
z97313bb14f642596f7bc766e45ee9c8c25350461fe71c1eead6127ca5e3f8e39ba81c2ce823f7d
zaca1a4fb593926e989b28847a068323ba2580bde68f337a5f9b854356f7663b1d8031d3abd1bcf
z1b5b9c52065d8be56104589381793d5febacc2040b47783ac12a665489ff43643a2105cff307ce
z79c8914d49ba2318104acca1afd8106dbdf48dbc3f1bb65e876b4b8c57d728734a1ccb396a12d0
z2f752f8b29be780e4824495283dd34694a7bfb250b9ed6dcb4044c92ab289fc9db30e05a0f3554
zae91a6a463d56763e17caf04dadfa4a88b30c899a92cc4d7ade86966633b037be1a5aeba19d793
z442e99cbfd3be235cf4159e3a354d016fdb2f99a2aa77569cfb284b71125be7f369268bb359ac6
z7ac052f89e247ea9c57abc52b771b0a095ed4a77e6e210bd91b0a3f246c43cc729abc3c2c0e3d3
zb5d4032ea05e652310a4fe9bc63b4fbd00c18b648b142e2eec1baa039439e25575d2c4852ed3a3
zbc75519471d2e77d96c1ea278905abdcabe407ff7eb438ea6c2081b4620b5bf5353f3d6f01b4ad
z88b5df021ce0ae02f9c0592e7a06b31fc176417e263dee20829a1ae969ce14e9fe9dc2a02fca18
z468c6068111a2f5b52d42420ac68053c3f69e518d425d98b0e0070215a54770ff22be5e0ca04e6
z765452a5d083eb3eeb6732bf24be65987fbe4bf436aca74bbca8020d5556ee7f985f7c5370248a
z46f1bd4e1df9560ef5a4b66c37f0fdbf2eaa11b106fe7f1e88fe6e526a185f3e5b08738b1e1d13
z334bbd4b5c0627f069d265f852f6f22ba01529f847d0c33116fd7030f10802b33ab65a13f1d297
zfab23db452ce4f8f41cc31b376f2fc13d57118031c75f3d6ea805c600c6e3b23ccc5ab275e93a0
zcba04f41b257d0de28971fb86c443572921da7e96db4f99a38cc665a5ce66a207240ac9821305b
zc2aca3a725e8a6515a2e74cbeaec6e0a8644a6fa11369f3913acca4d34052bbf12baeb22aa9ecc
z939f307d7d85e2b891765bbeebfa2d12bc17ae0ed0c65dc2193c5ea4db70a78e5a9a3c43bc4efd
zd8b8a6694cc6f74653eb20d699cb404aaf01c50a57b8d294ff456f6d901530e02aa69805755182
z9ca1f0dda75b1107bba12d1f34d9125648d38bc5419d4e720da93c711dc9824578385180452c00
zbaf21757753f54b053b974635784d5b39d9f9e4e08171f8fa74f23ab0c8907ac545a6cc1d966fb
z68229f3aec6c0f3b3bdb913e84ace3a287bab456b7a3c1a42cc659256933aaf41ca1ceb766e89d
z5b4c008d311ba0fa6e2d7a704d4655489db6360acbdc34686fe8b285d18b369a2d62d352566108
z633479bb564c81bd2ef305773ee40b39333e75bdf8722fd987ca3ae167e3c2a018e0b6950c2a5d
zeb312046bce9a345395b28498457e89bef5d0b4d991f969de36582335e684df9bb9080b5fea0b0
z8987f7e79626c8e6f14c0bd0856694b103287f5a168260b73e413914d8462a4f4cebd23873c267
z25e671dd90925fd572a037f995d6d4b70d0f43b050a431f4d389a7f87a8ba57a35403b8eb92806
z10d369cddbbddade0986c5c9cdd16430cd0194e4d6278e16f9490ed4392f910acd4ae31568f75d
zbf549a64641bd7c55472af7928006e57bf772e67b3ffd2693181f7dbde085c21ba18a4b0569aeb
z1eac2e799b2992ccae6e0bda11c6c9d859007f01ceb035e3deb63895baeb1759c430ca30374108
z491f856b35faf2538985788e7d62838761df3819f554a2718caa9d1d348d3aa670f6b4e60008aa
z8dffa4d9ce8b72507a368826173cb364c91fa9b44ce7f1fa5de7945362a97d7ded77301cb0a1d2
z27cd30a44f4d3cf0461fa1ca0e9fcd98ee8cabf027c303bb78f10baa434ea0c4ca00deef5b8a3f
z5366ccb77da317754088efca4741fe1af70f934459d45a332751441f21441c79c3b21f136b609a
zb2d39a01c604ffde24dec0561f6764b87bf0a9325ca378f6f3c9974341b29285b96fb47d058ae1
zbdc04506fc617a0eac149093698f43cfcce23bce22ba2f5549404cab7f6beda72b472095430357
zc382ae2a84d9575eddcfb767e7eed8d71c8559303e8d571f8d2c6d5f0ee2cafc06abc83b4bec5e
z548a087034b0dbeffdbaf6df312c7662ff8ebee7ae3f1a73f81fa242ba5a28bfbac8a5c5d571d4
z9d30fc636aa2c380f42d070c7754ba8d1a528bfb31000864a6c5a9811cb0b0642ce291e1344f9d
z411b7bba4c11b4b99363595eab3dc03be935057b4ec4eb2758432cf77c9a4f9048c7b0f923783f
z866eb013980dadda17b5c86f2ad464c5011ac94d197a2fb17cfb741445ca493bb530446349ba86
z826deb244e93c8cf1c06318dc7e1392f18a3bdefb8affc626480a312f7126f543eb59867ca543e
z90f5baa2c7c0c5a9c5fb2f0c6c09606b595b1ca7f9962169bed3eda8012463ecc83d7c13e2396f
zb4a85fc0680fee2eaefa00d0ef703098b100211d185e509c2cc86b8d28cd704f256d69a806a90f
z00ae721a552e7bb097829bbad53a33ecc3a65ec4e8ef79bbdcaf35d3dda4267f65ac6a42a6635e
zcdd8f915bf4e4862bc99906039f3cdffd96570091a259f555ca1f9edeb8b0b24b3eeead93feba7
z4681f02e7e48f34d8fd5fef91472e4954d0f345c563c868e6eb7b20fac489d08e5e98efac36102
z67e3f72d5c22722c1a5bf0cd0c71a8e29dca629762a78055936c10862eb69929d5344edd96cbb3
ze315748db4f590e3e5b6a9a5a4600c45a8065abc00d99cdf8e9f224a0cb210821e950599b3bb40
z5e5b141b42cb494b29e64a1fc4ff6b24c26c8d1f70ab41c90b3b2c34591e4d1612c967d300fd64
zf50d83b1583a9092b922aa5903e7504ce8b5628598fbf03d0f7ba6fcc105a1c7ee906a6556a223
z8d46b07cafc54cc05fdcc5285ad6677d369ed42b08f3b1f0ba0294f5d410d63cbccb0420a8c35d
zeb61c6d376b7b4283688f068f056e8aca144400b394ef099788a5e88680d27c874b4ec1899837f
za5c7de9887e9598909a4887e37ec0370a680c05d15d59d22d10241152a58fe3065b50778787e7a
z422759b922621884dcc32da4144d5f0a7dad8fa33a4073e98a5fcfe9c0d35bcbb0fe2245df30cc
zfb26c7ea0be51f24cc4bc66a290e0d61c00ecd927d080a3cb118e6e68ab014cd2203df6daa6d45
z559cde128012271e8ae9cfbed20d76a0eee68b23a0e55ad0a9f134dee836055e588c3f446159e0
z3c1a16ef3e5964dbd27066af33cebe9d859607af28a3845d120fcd859c55072ad058aba1787a23
z584cd0fd99bba5126f40717046bb4ba5de2cfe26417dad107dd42caed738b183e9c1c242e4c73a
ze975a53b43ee8da3316485120a9f59ae468ca4459d6f5d97df1ceffc9e8b304b0d7aa8440475f4
zc43ba0ba017835411073eec32b2b81ce0b1aed79cb491d5a5aa64fd90d3f1acb64a9031e402eeb
zd5ec44b6dc4ff7937608e9f500c24db1aaa5f11d791fdd54f6b2139f49212011dce3a86cf8378a
z1b201dbbe01bb10025cec07eea70355f783c62c87479506f7bd74ecd495ad191e96dd756ebc7fb
z34ad1e3fc9ced758adadffe846de1dd595e1535c4784479e8534d7d643c5bfa2c690d3a31c2389
z3a35fb5453405373d2fdf8553c970eebc4c63b05c4837bdf3b5ad30ce134e41c371c192604f7fe
z7947d2a4770ccdbfa3dd844ee4daa77a00ba538b7cb66ff5971aa21482e5c5c910584cf13cbff5
z61063e8f4ecbb1286af6c56a56f38b9378d07824fd01a65ed7d418e21e7373c62f0a5bb7203472
zc4a9e9e3eb345e13224a037745d0cba8f371b0fb86fa4e6d912691a3f46d9b272a215bfab19d6d
z6e4ff1563e47750f7bcfeb1573ffe52c17c66d2c267585745bd4acd798e6d95b339eecca85a284
zf998afd2708559d018be9e1a379c55d9e944eafcd344de867ca21a97c98f51b15ca216c00bbcba
z77928227bc99e3feee80ba64fb4a3810b2ce74b77f374b7a469f7ef5d2e7dd35c9bb06ea07b365
zef9f63220e0c90aebcf8de7e67644a4afb1c0438835f8887400217be58db1057a6eeeac04b1344
zfb3bdf754d8ef5f26f5483dc99c945a70293eb982a0a1b62d49c5983b69b09542375510043f88f
z5265b4a2f18c742aefd06d87644a15e1911546cc530a539522574102f3b53ea76e4a13366b4255
z900bb49db2f0a2e2c372c50cece82d8bdca5b37b9c82a556c7324563e2314416ba378b2e2ee9ce
zd3f9300ba9a39d27a2bec9612e1f3d8b86f75cb69f59c4666e5f33afa883f715c36ae9b095ee98
z4853ec8b644d67ff6200f4a8aa8586cd1868a968c96ea7ae92cd8e66aaab1ff658cf15d5721d11
z5e197c949ea4d1665487cb3c49070495c68486fe8c4d97a73ece38958a300642f82875f3b8f646
z2b4d8599cbdd1b25ecda7534bf8aa5450b35cfc668b7d3082a4ac47f03176be8404e9fb4a53751
z604b8c08062bc96918b7786b93e89db719b2e5ef095b1ceff2234263468345bfdfb0bf305a64e4
z2b10ddcd43c95b1973a33505b79210f318f18f6d8dc2a68240fe66edffe4e237abd7f15f903127
z28bc390e6ac7ee94320d05c51f95626ebd2ba6f9804c44a840719a850a4aae090224dad8be5093
z2e5bea1355d858604f61ec6e792ef739f314ca77ab677ebf378f05aae6c8d41310811e58f82b00
z15125d0adf0d73344821841231cc6dc98ff2d379276e0a9ec753cdf7385ed1645ec9f09bcd783b
z447e6b6c3e793edf0756e20df303700514d4c7c7d6433fe4fb6ee56fa54c76507d19c2fe026455
z2ed806bfe7855c45ae0af95adcf478864cd105825dcf0d3b8f78c820ec746de63f9bae4087e399
zab57d63a9767967bcdabbac2a40cd16d6860575793471147e1293046927972c1b958da116e3841
z053dbb22a5072be236702222748ab1cc037d4cdd44e4aa1512704dfbb9386d0ebf246f76724c46
z196f61c8c6082b64929e49ae971f4968d859e6f54a39a109543b45d9cea53a52d3898e1e71be29
zbc08564718273771d26dd0cdb4231cea09cd4ce1c82670aa00c5d4048cc27a30f541cc56c60746
z2d1a98ba247da446524b055eb55c8eb6fcf66e127dd459b158724dab0502b3ed069bc08200eaf2
z69f233995a456401bf79442b233e653c3881f059ec215f400aeff3a40a8f2c0d7805aee5269f57
zd50c02f7ddc6623e468479c47fd34ec5c5203a6a4f6e0114e2a2c2808451d2a4e6f66430cf4d1e
zef31656376dec6710d20a6f2505ee666b6018935a7159c0d195d597619cd1c7845ea234a1e0095
zb3aebeae0f9bc85f1101c9cf871f9efb3bec762219f6352d75134f8d001920388231cfbdb987c7
z01f50f7f89647167ee27eefb3b62daf7309e72ddbee4277d8de84b7b2bcf1f9109b0eeef2126c6
z57d98d5d305f0720484c8a4af975ac3964ee12a436f01a8b7b4e8e0a7b0713868b32b58514e68b
z81d18a89c0b08177e6b377da4bdcd93b529258bafa30644ad3ab0b678c1570a1630e73a0215338
z95f8610beaef3da5de0151a183f9e59fe394b9bb6ef766d33a3ced281d11d1597e208c36f910dc
z075f6a0725eea5269f83d01b08c4b496152be8adfd8f1d19371db898bf08ed5d1c5fd7bde302e9
zaa5c269583b54358fabcd5b62dfebaca7c6aebed5fddc9f4205dd79b82eb1fe81646db4619fd25
z2a18f63ec6e5350312f982337a6b832b9093b62bc4793dbe4cd745038016164dda60cc0b12450c
zfa9e4fabf2c5bad060e1ba773d0fbe94b7718c5e8a499547161909cfc885bf8f39e91b31742678
z663d403ca48e6a95ad7e01935486a156bc220d05d0954c634ba4228b36864b55d22c663835b74a
z1ca51fbd35021cabe48bb370facdc34bb764bf1407d5c4ec40b7ba00eb95d61b8a28e432ba0d18
zb5226e495543054ff7c63e197d6abf52299f5b982eb3ca55c6a589527de59b39b5160cbcf59721
z019021266b844d363686d7a1b9c2773cfe373e91d4b41ae698b9a63bf198c44adb5e96bfadeeb2
ze7fe1d170195ac5f1abbd6485fdeab2082b10db33d7c0e471b2d23c36c3c5348d838e4925d7028
z170f35a816fd86961f7188e401976c145ddae046ff97c87f6e76c23b6859123d18488c5486009c
z34e160802e05e29113bd1a55f9f91faae7a33d83334acb16590f27066b76b4b5b319fc82198321
z6369b3a243ad53494d08240460680d339b512c54b06f4fb6fe618c57728169b85957044d8d482b
zcd2a9cabec94520f7b6bededfd4009d958974a23bd1d360e93fca2f47e5f41aaba27473cc782ff
z2c3ffefdf0e084fdeabca28f85bcb40e2faed0ca4ddfb5f7312732103192b89ae6f3aec40a913b
zee98f149a7bd2736278d5261214206d2b8d35c30c7626c2a42cd66f263d930f44bdd2f9dd8d266
z20b2adce186d2161657714494884b95561352c2bca41ee6f0bc6320f446ec22ff4b478d148b9e8
z7c711a17ecf7dc5a36280c6ac1a91b6f385586ac825039b3006059eeb1592109cf0d7342aec8b4
z7f4ee9842a6be40dc88b8a78bc85a69e0340e94d772cec26f751e0631555b6912e6f48bd40d892
z434e76bc7c6ce29d5b6d956ce42986df3117560a043130d12044387526c2efb698dc7de59be241
z55c62243fb8edb7e1d8040b0959731e463f75b6f9b5551604675d424ea5f7fe88f5d444edee326
z14518bfe4d5ded6e6cfabfd87da69703c296a750676d2cf15ee3b5834ad6c88db1877470f2adc3
zce641dd343c220705a288ca1a0d7a8fcfae8414872f3b18bb3ac8b20d3116ce745e38204fdd897
za0f51840a84473a73d2f900119946147fd945a4b093e4d9752af952ecd6b95b2675bad55583794
z8033307c64e7bd9e64eb01e76b8c1119ef77352453e01d6e0c411afae166a4cc63d9c98ceb0f2f
z0ca9441b7b37ad7dc517be27508538a3ac7d95fae68b3139cd86ec820832f233ba7efbb4e3b671
zb0eef10bf30d14cbe9c76d8a413417961385145f018199cc5b66378a6b41eb1a98df17a9446a25
z8a2de2b79f846e001a5a8ce9fe9ec904ed2c4f468fcc6aef74795a33989165ce26d5f7a8431204
ze3446534df9a9e248c9e0b82d1bdd8d1c58bcea31afbf5ef7a275fc5de7acb22255766730d3223
zf54ffa062a051db8b55837d7c370e36372c49f53c86a8d8ef3812c68ed99d3d742f5d9a4637eed
zc9e48313dadd62be18afd72caa911c5d568052afa9df592b44c3c31b12b5d04e381a1a60ffd978
z45061c270443234f3ee068797b7cf44650dc865e1593a528a028629eccc9518423186bda968972
z9a6a87ef4e6c7995c87ebdc4c40e3872a5bb2ca6bd6bb767ea626200ee85b5c633e277b51210de
zf385eb5add4a92e6ccd4779026e99f7c07ccd9a576409ec7c2d96adb6d60d7944df9cb693d1483
z9e9ac6a01db042f44a5c483fa003b1bfa1a017b80950956f1fb7971d681a708686bc131b616e15
z305ccbbcfbee2812675226056670e4e6500831e5333dd847304e57733934a6a92d0162e6cedd1c
zab8364286db4e4385d390e9079048fadc7c07befe781f985348d87e556725093590bbe0a18d964
z00b9ec2279f2dd78e3b14d56306639287e03b363f73815ddd113f170614187200e17ce60a9d449
z5aa3ffa20b820f4eb73f5d4d06d1e58d306f7043fd853665297a1739ed61168e3c2631549f36ea
z3e414d20801da14d39fa3bcf292d9b815b817e2a3a6b81241ef2db07153ada6b3739bdf9b52ea0
z227e3d4961a6621314a592894b6abd7dc3cfab5f896dba1cf1cf0f3a2cda04682be2884d0633eb
z7025833af13d087c1b0a882b596e8fc2322f9ae78df6f5b704a768d8f0b4d71d3c66558e3fc762
zfd7445f196891ad2a97c60a61479551300f0263d6826b7c860ff5c2417c643b523322f57dc1780
z37313f618ac92200e854ccbaae2c16a93b8bb150323988429758e9f5fa4c22c57e4cb19674c542
ze7768507224d7f68085c34afcc66b57503f4914446d5ee4d059a534a3f1427d7f19c12dc49553b
z24592b6a362d227e4adc90e9209a90dda321f9805a34c9ce235db20b3c5155821b95b3ea486959
ze55ae5c252fb60f391237674378d81d70185f84fad7cc890607d83533d3fb8fc6bc2d52debfb7a
z23175f283dd81630ea093e2091827c68ade72a73766e59887887f50d6115cf35375be7157ef660
zda85c1106357fe12231f34253f39454be4894203c45cb15c1f0cefabcedd9fba0daf2a9b35de66
z15d9da06583ba7ed4448fd1b79677cab7e2f70cca9e673ad835d10dea8840b3146ccdbcb0ca2d7
zdc223db649a00ea4030f7fbfc33217140ac028732fba23ba75d4b517988960ae3213823da61c32
z24dd2d34a95621ffd66e7092d9816ce53d2b9afcb7267fe9934c17d8501a69eda87bcf7e21bfcf
z9f5a4807a07896e7ceef0f39a566dd2ddd01f64193076c3bdef8f1a70ead79b90dd4c2a784909f
z329c95ba6a464eb7cfa30d7891ff35d3bed2973491e9ec2278b1373f5ca4c765e9e66c22068104
za39f628742285a2e7541d71a91cfa3f5854339da1e844a75868ec7af2046c9337c0f2cf9c7f9b9
z0a39872c2577cc005ed6bfccc5a7844a9bd484be2f58166c03e3534baf5e982c2691abea7994b2
z3215386ab1ac7e4ec60663a1e4373fcab3e10bb878b1d140d3c0cedb966438b7014e1e4a82845d
z15a74fa21725baf97d17c9f05051333431ea5bf7c1e893b928b2d343d37236d3e27bc2a39b5998
z1737e0975decf9aa09c4e872778a49ce8e05dda28d82a6b61b23b03d756153ab05a6ae3c37cca6
z2cc4d7294c2cfc85e78d4d8d850ca87d43c4c32c0aabc5c0325786f17c05ea7b7798575ec8329d
z81f958c74ccd8ab4aa4bc11c44f72ff6c04d92f11612b9467b71b726a587d1ac60e93691ddbed5
z633f18b5ca30782cfe1c107d036928075f8a6b85b5253a19df0ebdcb0a37c33cc2d9d56e9e31fb
zc02295756885a9633ecd3c9a1b96a1fa4ec320be95df298c983179e54e8ca77a952f466c80c472
zc50ae5cb4cb9713dfcafe8c18965237ba1909421d64f31c366ca887c6038248b7899d1d0ca162f
z7842400da6d8e81847c1b73449b8460109679127e225a3b50d8555ec9689911577076df6ea7ef0
zf262c1183f7edcf63c98ae1ab4105e8c98ea2ab9242874db9f8834d0fd840d1d2f607933462c23
zd0813f6304f0f2ca4ac7a3712f0203885329c2a83f3c9762ae69f64a83e175fd665e1b2fdef2a3
z54ace8d03c84f80d1c4147a14d7836df832fd619eedab2162fff7f3181b6eb11b0488d9a9fe206
z0179e17b02d580f0041af03ac69b95d5ee8a035d3c66305a2e4b92d86a5e8c7b08d31c317868c0
zd9193780fe56785cb3adc04069974c2a9ff1cac6259f1ca7d02d340480bd7ae99535151fb7dac8
zeb2976b3c41894de8317abc1e1a5bc28295c520c896ab153739b21de3218a44fa6040e2eae5246
zfbf0603e333c0279fc28b035a1def0c34b1b9e4f1af8be0937d680113b2466ff52da54e2ca8582
ze4a866762019b0ee67a0f50bb66b823772f1e0e760015759ed2f232f24cfe95470bdbd6bf570d0
zd3eb2261fd8f1feb0618e7612bc923a95dd402b93e1cf0618b5d4965109de13894e733bcd076ae
z7f9df261368e3ccd26501d3e82709c4e5880e06efe4bb6db9d0b2e4f2899a615d07fe9dfb3b517
z440df5165ae005693126a599018a72184befcc2268989a943298a9addb82763e3a0118928c91f0
z134b6489463bcb570dbc6e85bc5339b3b765aeb242ddaf6e75d391346e19e8ec0dd2476eefc374
z013bbdd2d99fd39798673293d5babab264375028f3ea0b103976264892926c749b6bada655c72a
z000e66a33d4dff171663b0ec4ba7ce21b59915db2a28f66f05d734a04f67ec08dd0f2c0d0e025b
z32616efb8bfcc8be4fd8141a4e82673d140e9f18115de0b287707639e99f033aa023c1d4f59778
z73ead58c05496346d0a4f0f426fd3d97b55ea528323506af6667d4358c270557ce12583df970fb
z77384a00f0d569f6b22943244cf2af6530730b80a927f593a31c9292b5a99eb28b3e7557880b73
z20b273050680536759d6a357d9ec9c9be1e683b7e15eea66d45e07b19ab6c7cb46262216b0f53f
zd14da269902677cf5635d9ceb75a0a85de84e1e1f8bf45f3c9a94e2783e0e822ef94bcf65df1ef
z0441a308b5dcc49e7eb11250d05657dcf33002a159d34e059579e65f3fabe240ae6216a6471e80
zfec2ba647917fa01ef02ee72708261dcda3e9cc7ace70ac6675216d49fcab89e9fd4684c229642
z2a1cee2ef349356844cccf88d449b013521821a1797951cb466dbff3e98aa7b5cd6d4a6eebccc4
zc5ee1bf7ed7f426d240cefedc10f18b25bab252936e1fa64d203c4c3d52ed64e8aac4d046a7830
z21e27ee8756c27fda57a72df85fa82f5bb82280397a6c3ba8728ddd2f420248893e7a217453c09
zee01a809c726fe1ae2b1af27eac77a0e57d7373e9f82bf212646c62f866ac4bd57ae677bc5097f
z0d0f74a96bfd0956a65f44c24212e07b3a7ad0e79e0e362c59af0e491733f5ac50466001428abf
za694d690ee97bb1ecf5acf524e3eba72f01d4bc825661cc46d65e6871a2c710837c0fb2b4d2a64
ze076f7b088168795ab7c025e8460e8c898c5b604405b5089ddea5d730633237a5d3d2d5e02e574
zba464450d50585349d9b246d30366a30fd145c312459bda94074fbc11abb462b0cfec0827707fd
z749217293f173dd8a254f4c885bc6906be56662a7a49bfa3535fdfb61b7e56e6fe2923c0c2f7eb
ze8e4caca5efcb85bcfae630792ecaf5a13316b248a3c2e8d9ee944ec33172e98befd7b48a35c62
z05d973a9312b32c5b500721c5481359f20a33ff9a2043e667bfacd836e21e0243a82857a4be586
z4678c5d776804cb42ef280354d8fd08d8a6d73c8380de2dbe1d090bcbad7d89ee56aeffff12be5
zf6f3baf312c645645ab006094a8c58052877508ba733c09466c2872fa791394d55c53a4fd924d8
z69e693d88935b5cbdc419b3ffab0048d9a0eecdcf06d65b9a4a84d5adb37cc230f4f755ffcac30
z355622f5631529b9a3d87a2e65eae849f091be1d8e6ab0e6a65dfe6b98434da6679e83670957d3
zab2329801c0b2d5b7e642ca93b465125e02395d06a2e2c3bc531d68ec5f7d153e63dc13921300b
z98b6bff3a1c434a9f3c17cf9978d2f6372bb8ce08d6fca5282f39f1cf14bc0185dff8769faf612
zd550226aed7766571d67788bdb73b7b06d617124f6d85664a2e0f027ae24ef9d2512a58f8d11bc
z6eccd1785d234030970490f69e3baec0b2c74b36517db92093db0e16253108f53031cec8f97eae
zdf93f2c16303488fd939b068cc49bff8dd7bc5f69c93a1bb8a6162a9ef32aab0485c2b56d7e25a
z23ccb0c730228942edadbc7d19312f2bd706317f54e5f1cd8427bd6200898cae7fb9cc73de015d
z17d96ba3e1895a761ea16df206bd214f9f66140d54230c9800da513437bda642585f9eed4ebfd4
z1a50615d1b0ce81ae90eaac1c40366ed0a21f7eb5c818c15d9b08ada970c902bac565ee38a5123
z764dcc5497b29300881c209cefa09987fba41faa7b8abc30e60406ea255268d3e502613db51a4e
z114f3824e2e8a73e16ebe1aa134586d512ac075532456113e4a4f5808bb9d22c00e76ac0f4d32f
za591157c1929895ae95deccba33617c8db6ee358d88626391d5ae5e8d06d81dad42c9fab96a8e4
z8d1fa59927e19963b7e2d5200dff4c2c8e05c240fb6084e56a1c346a2fe8a3bfa4ecf4cb47d617
z94d6b0e1121d40ac2bd298071d74325123e3eb6d2098c9f17ac2f1cfc1ab688278ba2fdd87f6d9
z2f92da61c91944d9caebac227567d000fce410f5ff94c1aecf984ecaa5ae9cdaffeae6548f54c0
z0234174b75e614dba173f061359ade17fe23141180d3b61b34700165cabee98cbfb559c975120b
z8e176d656686090b1b536ba257610ecdb188fc8a5272b92834775fca523aab48d6a31ddae314de
z51efa40795c6592ddaad18e637e27f8205a85494a509363d4704fefbd697a6c1010a26f223f791
z5a285f172cbbfae4e930522a801fc4e1b055839e244d848665a5b1bf39390b212ac6194081a7b2
z3c9da89862c9e67ef0c441e5c3d6d043ece7c183fab3071c48de0bb2505352d43f15666e3f1dc3
z3b234368c1bcfe9ca769b1a9e34f9dd7364d027fb173c9b3b26a40214ba810717cf2a85602024d
z325337aff8c904270347ba8d1d265c6cb627fcb654c4d65b84bc946748535cd837ca2067bab881
z84fa8709303964494e7558c2e9264c814bc851d2c4edeb584e85e9b9626b03a3b584b001a2e244
z1e307a5f2e9548cd3a4dee9f5feb6cab1ff87e4a7aadd3147446b21dda6d3e12b52275517ed9ed
z73e291aad17d0bfe697379f945fe4f89edfad84d42b673727527dd8bd23616dbfed466f1ece20a
z81ee69412e14909564c931bcc93deb0b194b932add315be8678deb45c96469097195bdb86c6cc1
zc1930b6f2b7a2aa3449d07810ddefba38d4cc1ceec0a80df44aac5b462d2608b1cfade8d7433d1
z18b9794a0d7347306ef6c91f1813179d844c62405392106161d1c3443318ae4aac15c3d0512234
z81e18b12d96de9475a7bcbda99c786d00b0bed82f715d3bc98598650f86b6026a4a3589715a9fd
zfb1c12668c9a911fba64e056bbae523ad64d52a631044f9472a58a4dd4311f1f70e52ba90360f2
zce5ec5a2522a1b182a75f801ce20d40958dc41e11481b26b4299eefa5b5ece2c332377ff3f4f57
za8993fc79d98721757e45f9b87234a4e39d5776f7851e461e2f7c35254bc49f2735666438add69
z27aac6cdc32320277b8bf43874cc7179f47bb93e8d4f69eecca32d4d20104fad64f923e6f62437
zaab5162e25e92bac2d52a28f4184fdc91560437d034b3ecc7a0ea1a02ff87a6a7b646187363766
z14fd2151e4ef90f811afc739cd112cc995fa64572b49e74adcfaba4415fcf78ca322b57768c26f
z6d3329066306fd0c525e03f1543371308ca233de6a5d588826985d1216f27303eb2eaafad85a7d
z46a038917e649af599cc47ba5fadd96379ba523e7af44f087979757e62500a33e1822526e8f7c9
za0988c2cc72a6f8d724956f40212ee700c44c30a7d0a05d466487941c9f89d3020fa69161f57c7
z46156079e9f054dffaace6cf53881d04db0950fe5f6e790dacb2c1f1a3bbb3258006c7fd9aebf8
z30f3151e10281b4a78b35943b10fca980aba57cb0cdca33a8dd5f3c7cd7f5a8ebedef6fc0da839
z9e52d610c9069525fffd3be4b5689ccc6ffdbc565f32a8e2602ce328b34f288477a3ac09e75e15
z2ac53c23ef5088996ee53466e589f20176f5714d202ac29b4549a20a0b22c06d7b0674baf4db1d
z8fa6a5402127901eb7594415f0a4e9510276a172e8580993e4617908b69954adae230c39563972
z71c2f7d44053484ca3dd48dbf91b7b255f9de721ef43a288dca9a98862c4d96f2e8afd7388cd1b
z5b613954509ff14adec0a927f5638f558bb6c206549c83429854746893f6fcded8bc736902dcd9
za396e5617ec659dcbf919824359bf92041dff0ddfb145b4f90f6a18a2fec2c798ca5cccc4ca5f7
z2a88f4d615dd4b5e83062a41f0f5fc435ea264aa5a04c7e246a0d1c181821ca703fbea3c9630fd
zc4af0b9ab383bab0011da6ecacd4f5de061ef2612c44ba36b04ef9283e6ca35deab88e9a41dcf9
z5891c307c55c80085afafd27d4254ef79d338280880189356e0d00d583541701e2b4c0a1524301
z1e921191bb2c317d038f7d288fe245eeeec80de254c5387fdb43e9cc20d268830dddc9c4aca979
z86a9f65497a45eb79220c5a8e22c7bd891645b2f9bb0699a9025a303acabdb225757c08a2b4eaa
z0b668fb437fa96255b8d19804a4ac30b5f44fef59a7c7c6d04edf64e3aac917e14f39523129bd7
zeae51c32ac33e0e0279b5a17038df956a7c67cd2586ad531eea4c1fbdca1d3cc9e2e009c6924b2
z7aa7e042cc010f51ca22b62e548a57d05693b46ec7a724371e83ae65046f6946130bd94807cc42
zea6ad71ab1e6bddbc744af2f87e36f0e57be627fbd30b0b0d93e0e2d13236e43b4d8f581302670
zb3bda913619262ee184f5c7c626fa45772a2e4d29e246971054c0827135161a3c159efc987154d
zafdb5f1c9432d78564492d875e2b4367119a23d489e4056d38b380aa6c4f754543b019da715fce
z54f15acd2c678773530a616c085fd4aebefbd7d6aa7a4f9f6a6802e991bfb3029d6a127e532295
z7855dde742d289340a583b852bc090e4c32ec075501911fc58fda2ee6f8249c08d3e6e735e2b13
zd61a1a14248060b25c03e92abe190143dcb5de0778323d6ecfea63bb5266e6275d06bc5e19b0dc
zd78eb923b7c1215c6714611e88ab4662d23a5042a25bf0fcb75ddd7334f7c18d268c26c9102e76
zfd55766559379eeb6ed8181b609ec745ed166bd9a5090d565d90af380358365f505896ecae95b5
z167c6ef8598d7d2942407e8658765e6f4ede4ceb24cad9123029d5bcd28d163284b9866a41df9e
z31c194871bb4c84f0ff3a9a337cc6031fa2d82dedc73f885805601e01249d507686b44544bf74b
za480b9b32e493540a95a574ee9dda49485f1985dc53f199e9f2bf7492893bd8c6932556f42b5ea
z4cb4aa7578bc142bc46d424b0ca7f56615534740e9172556ce15cd13d6be1fc65ce63295c1d61e
z1ebc3896fbb99e2aef74ce68537967156ec70ad5d114b6422d56d9c8606e76e63f8cdfab92fdb3
z3236ba40d0474652e473748982e04bb5abb90092ae2aa5a021e3892f85e8e7de27b1fbdfcd2a31
ze29168fe3a4d8a4ebc68f47cc55b4a1a4f4f6e63595de3c58701f879057b2089ed40e2cdc5dbb5
z499d32447b708fb56da37aa3d00f3f971ccd4447ec6c960c93cd525321b1cf7c512ad455e6b8cc
z6ed81e3d5a414499b04029535a785a966100a20db9a056457a65d0f4e6d531798356c83b06b9f9
z89bac97786b1ab7a3d3f648cf76da701a1bc2cf0ec99b8c392cd613db515acaf0fe2eff402e251
z640455f7072689f93141ff2069be1a965761dcbd0acafead4a6f693cba3f4b51781f2a055ac439
z586686ff9c43c43de671d91654d7bbd385922bba7c9f5b1f92278cfdca34b9713bf17085d8b6b8
z91b50ffe5c309a3de6518c7e90be47848198897261d99c438c522738bc38de8957c1ea3ed0216b
z5487ebed61e04936037132dc2295138d91dbe57dabad4298618d62c173ff3edf7b848cb0fc42c3
z95f15e827c176ce94b3514218615dee697cb3de2cbce3dbb55d789889b7fdd64e8573b2bf050d0
z9f691612eb53ea425ea62c836c58586602f807a89208cfdd322f1cb75f4121c578c91c77b662ef
z25c517e1b9f403f216ab8c6235d9e0c388a44dfa72dc09397fa1bec0942612038347283373c439
z93959eb221e9c438d81f7112c819167eb79a45b83a1d96eaeef588bffb309ad53bbec0ea63a303
z2ddf2589afb9c25eedae259c934646a4b8a4fefcd08d095a7c6bdf467233da58afee671347afcc
zf20bfa073389d3ef4609a61149c293bf2bdba29498c141d36cf0d16ed13c5254152ee0fff5b321
z26c199197b9f6f248f88a804e0407d48961fcc923d210caccff989a75aed095ab2807d86f2a29b
zf0ecf04e888f2bc8e7f234fdc1ef25bea5860327a3352397a90250be0fec12b7fbc45f5cf445d4
zf9c67e64574e8b3563e374752f8cc6eaa27db9037ae3e49d742837c36969e98bc5d5ff52954cf2
z8f374e2e2c36915c483669abb4d19ecf76bdd87f6d4ea9defac77c51f60d0954b94a3f43865168
z55a283162eec706d42fda06425a2bf0b3cfc84360906953a0a065b68a74c4446be6ecb2e2b0005
z725d534b6b163c667325e5fa1b1c79bd230ddb4bf76f94bff55a196a46a00c91656c89e7ffdf82
z6bd21e27a342dfffe3dba26a6badfe5076a9a7cf8d63fbe9fe706508fe96f09e72885e81c8a2d8
z73883b98d3e0f28ccca963f4cd2e7b747f28f8a946e6cc80a4d15221d9a7c4eafd4034b864c9f9
z6d6b1fdefc4f11e2553d567476bd6aba363a75997954ffd2d6de8f710fd6e85f1802bdab9b4d23
z8dd9f61022493cf9d9cbb776e150f816feae733d9a0f68dd3b2347471e045db0d0f4b84daa71ae
z67a4073d624096b4de1a1deea20213f08b59d6e9b3e845b6cce7d81a1d04e118494b9d1de38c16
z4727eb79b98e8f55815bfc968d9afabe0be1d51216742776646003cdb988c1b9c7d6c4b0f7e8b5
zc12e27e0cdb6e0a971e59c46a5ebf1605c709989fc06c012f8b39b5d87e0a4258a26ecf58b5ea0
z676001628231d11a00ae5ba152d20b653ca008c387a5a5889c829b1100c3844982b6d4d7352b02
z6d34634e896d27163d0059746e7a37b891fd15fb4c649705676f15b93caf442dd52bbd532d6aef
z67b4894ccdc3530967e81f669afb35f3acaab83fee08d95284b96292a34193f1c33beed692b096
z1ad64fced467ff219e39ebb12de279ccb3c6decc4c8494471e5e48ea4181c915a29a49ac62ab09
z25be4177f02dbe0f663a5ea0aaf821239612d07e47f68d794d85004dcb2128b370b70f5ecf248c
z2505ea94f27fbb40b0e19ce1e6cdffa1363678880bfdf828a78438422c598aa9398819c18fa4d9
z40c13c6203efab9c4e132810ffa592e345ec02bf98191686d81d079e3e1bd535f21a3a5eb77aab
zc2403d7d41759b3d68dadccdaeaf75beaf782e030b0a51341ebd85c211a27955e492cfe1a2a1fc
z07e4ec3877d5c1c02b54d8f2f74103815e50ee0497e831158e6ddb380e1d70d67c733603fa2c12
z8cf2659473d46cdf3c512513fd44a81eb72acf1ba57b468b5689c5041a7b596ab40fe23d8fc9f8
ze57632c676017d78047b95189f34abbcf017b879daa4be012137e4e53bc5bcb63a52d1d2493976
z738a70a682d1117e884ac4719bdeb23b3a81c55f214c569ea38e97dd7eda8d1c5a0fd08af65a5f
zaa575083d7d94a711df13d12cae0fdc668eba677c218e14195fe6f0d28c921e4ab97057e078059
z6ecb32ee5174b66f7e73ba973ad334993a682b3585286e7987d257fedb603e0055ab8f51ffd9f7
z5ce3a5d3aca64ee5d77d0ef546b97ce4bd0f8fc7ffafe7a2712b49121283de4b030378c714d064
z5a1ce610d56d07ca463a4d2d2474c6f45bb50868370d8ee7d5f7b8bc96c5ea14995352cd3df316
z27d810510220e7b4474b9467cb0c74eed694be579886062cfe57ac316ecf9e9792a9b520b400b6
z8f00320be5cb195054fd07ccdd9d724c9552a860a9d12c1f9a47a41d08ccaff9ce6a550adf92c8
zee06a192a2abf911c788207e795bcf1b195493d9ad6e0072152a7b24e457599c631d7e175d1604
z013036bdeda524d77e81b7b8a6ed092d3334c44e9c583e8db7b497ffd2b9ccbc59b687369f70f0
zaa386fec19e108dfdc0edce6c52f364477153eeae451bd9e93ded2e03bad228b9378f1b5a259cd
z8a9af07b4c4eb32a68ab47bf1a4690440752f5e34ca60605ffe0e421ea8c30ce390b72a1ce5442
z91372f91a0fb21af58960bdd5c6b35a97c1851dfa751897dece742bf2cc88c6ad0c780649c7422
zc2c43f8567bf2406f5d2873dc15c5184ef8ce03e63892bca8d3dc5ce9b48cea5d0859df99c4da5
z47c0e613f433f36e0373618a04a7ded0cf6212f8f07ac45a6f5f9c6dd2b6e02eaa5fea19658881
z57779074317907e251d507c130afd66d8c8e03bc958653d4dd4be0feaf00aaf0a36d813c3650c5
z5666a548374781d0086158ff433323678cd03548a32e4243a11415bb92b7a4aa98bf4e474fbbfc
z8461630c818200478ead47055167ecf9ac26d10d49f13a36f77b5b3404fc9703b3fafb54b65ef6
z026cf5293edb16b4c6fd65e3766b626c462c358bac2498007e952c39d2e65023f7d90163cf1628
z300d52ec1129bd14b944e4881f62b30b9e5a08799682a85533ae36d09a9e6d37e42265825e7fb4
z0a4c5770b395e44eeee572a69d5f53be3bdafe3a8bb9036a3a7c89155095757591e7174db7a2bd
z230d92e8c20ba6a51b01b48ba4ee8c77c2ca71be4dbd2397cb2a0b70539e0ea967a51becda2154
zeecff38fd7f696d634077fb666befd82583e7289b19232c295f4927ed29e5bf651cd25fa45c222
za97c0d4434ec1bec64df8e661f247b3385b5d235a162028c73b90e70ee9ee0b288c64822a481de
z8c9abf4862fbd6b1782804400866ec467aa454f33ea79d998604553d282c8462cfe37f66f48529
zb662acd48222022808cae4b0c4c06cb75981cb1abcb7f5afbd1aa6761e6713c7495874579424f1
z0a0829a99eb0de2624fd324cfe643b1cf7db1329f56f15e1483532be4fe5144e789e90e74b7371
z1f0e6a63b9832a9ebf782c40c4573736ce34b0786e4e1b91cc321a5f1091065739a08091518241
z3ef2041c62dfeebced8a50a5bf3a85cfb07e81b488f5c6a5c041f09882066b6a82b7285d6c46cb
z4bf438c524933853d4722da466906be3aa52db5f994753876be5bec978850115d3a6d9c854e993
z948163c58f8b4c9ecfd97a82003fd6cde3aa683d1e91f881c8a1262f7dc90bd71374b3bd4b22e1
zf5993f303bd8fdd07f2acf5723f2e3e45b7649ba7ddd752e12b2af32dc9d070bd0f4e79fafa212
zc8384d9be4751a581fbb3bf97876adf638f352b510de8fb5535c6d76f3c9809a5d1c4fead1a71d
z4793d2c74f0b621b09598565a83d2f6d6034bdc138ec7ae8758d306ee7d759a73e1fc21eeb5fd6
z2d6c82988911cba2e44f8e474dd9082f3bf6e09114c9364bc83fdb198be3a1de8f0f863adabf5c
z020efd654f24fa3532b398ed4f5f37fe400b6ccd49fa8d44a272709a351353fd99dc9a08035195
z04a6e37e5270507891170791e4f99c5c18a96e85f19a33b049b567bf251ac3db2dfcd255c029dc
z33237e0618d4429dfb090c417bd835a845212824ad9dea04819fdd010c461aed0dad4e65fa29eb
z7d662738cce3e847c21fa999a5592067b0dc453d149e219b22b20b2a474739595f64542e6fa9f1
z51f1c895c2f2ef962ad0da3770b05b2b05c938c87425b4b1679b599348510e97baa414e5cd26a4
z5be00ce087f455393d2a2b1c4fe1b904846771ea783d567d09237460153dfc39372dfc2494ecf5
z370ff6c0a3823e782bd00976296f629c5857fbf8630ef504e7d265602fa90e76be1136f9995c0f
z144493620e38b6f01a44747974ba8bdfc2b42afab165a80f648d5c630926ccf350e7df9063295c
z4f0cd062cb388d4a3f360f520463ece14a78932c222880efa0721bbfd8d1c170fae335fa1eb500
za061d929c2bdd37ff6968d3832b94fe2aa5346e394a602a80a01b424bd543fa244e4018e2a99a1
z3f2918ace7f7fbc2de2660937613809a54299678caf30f02ad312a8ad07d25b38a577ed9c96ab5
z70ff6461c325272f0c88d7beb29e7c49120b392ec23650fa0750d4099cace47e506664daf8b81b
zf8441285add7e67caba30b73caba71f4f526e44bc05426a31fa2a880029546ac798ce9149ef0e8
zb2ebd5378e9d74060b484f7a5cf0a8f109484738624b9b67bd54fb596a9d222b1d575be9bbca18
z27dd6adbd37a8c9f913f2721a12ce249811f500297e50b58d51dbf0da1d8acd7dc5123c2763948
z4448e6a9ada88c70d0089cf581321679fac745e3a34bf6983df8674397d1114a8706316bdf86e1
zad80ecc5691cb206233eb7066239ea95a6dc44d8d16cf019cba52073a592b37d54df4a1bb6bcb7
z135c9432670bad682b0cee646ce5f954a93e86b686cc59e9a6ac1e92cee8d1136df098edd72212
ze540a4d7f72487b7b533d882399840aea2442430cf1adae3891475cab044fb966f2945dc0d3858
z85cf9035c140173188ea08a8232d06c29420d4e83354596247f1f1774fe34a67253a50983e38f3
z48878f9dabd7b0fa55ef0d062c279a06924163169ae02ebb6f22b824e0af435b1a34b42ec5347b
z1e653331c9112c12ed4002cf3502de2df5d079d4dff14b34ae6a00c1129fb816162e717b7fe32c
zdf272f8ca5a5a02446c318cfca48f2fc718527afd461ac81e176050e1f1ca4f245730b713693e0
z0ffe05934d8bee5da994715d279fe9e51273dbcefeccfb0a3e49ad7562c7dc3d62e35c99aa8a1a
zb4fa9f61bbaa82a1e175d161e57301a0475651a578bff069f6b97a9dd7a40b6251be57098b4fdb
z89711a44ea86b6fa51db3a49a8930d424d8ec9f0daae3d2655f75c061a4c09fa1b34f7b2bc8e30
z294f750bcb4cf3183f2dae3d6d7083df5565466b2e570444bb426d37d138d4bc316f1d522b8abc
zc3f1424313a6c583922c52db480e0ea041e0c4b7e65d2070d8350d666bce56e94a3b4446c73b7d
z65acf06165f99e7e4b7bbbbbafd3420e82f16f6d9e73bf16bbd244ec25b2a2076de25e598e36d3
z5b1b1908317f1bac21b5d54d5eea525a5270cf18ed25149c1b4c36e9ff866511b1925b832b90ce
z2f2da20b739b0a4a647a4f51e264d4dbc2279310913e351d791dcfaeabb9f1266aa62bf8cae88a
zb0772b5d2a0687c0c509cafd8afb35bf0e221a118453077ab84a33d7da61d8c3765564a65bdcf1
zcf4dbf23b35750e0fa22fea7479b205c012efffebee29da5277d0579b873d9e02909baf33a3655
za4c6bb67cfcd3a3a827db4fc4a8124fdf3bbca5268cb73dcba2bb7548e159cc18c4e479e05f9bf
z1a1477022c3bf82e7b0c003e29c098b095f44f57e59fe4b0ea5cf00d360299d27474efc2a8b0af
zd3dacbc6763e9d919fac91d8b3554895242ebfb13919055418d88a62ace3b9a9a5a46a2b64ba74
z93df22f73f4d8fe8bb1dc03f40507cab0b003067f948cbe1a3cc0451a379fab8272b51e3e4327e
z4792503184d6c5771e19726a2fe6af29bbc07d16925fe197392b2dda6cac84f207e5646d98a4aa
z37e545318e6674058f8343003f42cae9f75f08334ed1a2d3c138e9109ebce2157937afbd1f047a
z179d9476b5415beed79af307083a0d714ee840894d4ad74ad9505683d9402fe53f035bf07cc02c
z532619bb6c0171a8a39e73dc679a8952e23cc5bf424fc58e6e38e523a72621aec6551bb084283c
z6c78620ef8b4fc8c02f21cf395e0c640cce2e2372ca780db0481fd17b64830a8425a84624644a6
z5538509d4864e18b5129d0dcd6e7605bfc3a34c574694acf36d69f4888729db1170cd87cc5ead3
z49491be018aaa8d67fb47eb8d98d6c4c52668251a1f62ae7681353be745ae7ebf0a7c9139e38a8
z2ce84f088e36a6b00a2dc37bd7ef1ce4bba50fc7952606eb7d50cef85a26efd5ed38670010a9e8
za6eb9fcfe404d401cdfe9e91e89367ec100d392a24442cdd2c6e9eef1ed9002ea5e1dd3c69bac6
z8b20a1ff2c45c098ef514754d0c61079cff90bad890c4ff06b190eb0acd8de45fa7461baa9d917
zec953b48606e98fbe42bbbc2b2e22d4561dbc25d2141108fc42fd51ddbecc1bcd64d2b8ac7487a
zff47c40f5716c4c26a6ae3ef920972eb0c345902d9d93d048f31f164bea9b5cd4b201f5bd9f01f
z081cc04ff592b437eea6aa0209e58f7761d6b06df9a6395199d9170b5b37d1c17d71f1fc61a6a6
z5ae2783e5262952e7f8913b9d9478d00cdfd276fb40f4ac198393cb4259cb672bc3109f232c125
zac37f90b94c5584450b8a1a2d28f6709d4babbee078e14fe3b391b4e3cae2057e76170194b74da
z2ab62d565e647b3ca24ee3e7061babf646ebfbab045c4dbe65a6b932fce7d156993073c57aa17d
zec0636bc85848d9c04de4c3a6943372da21bf8654d2ee1c65df3652a1b02c7aa424cb1bb85442f
zbb194e810a21d87e0128fee25eea4f3a71d55d79aea5029d5e1704b63ae4b54cfd7fd1024ce913
z53d27c790d81f09249f566cea9c76d071967c84efea586b3f9b43c9ff5c88bc706673aa3639f72
zbbd5ba40493d4c7bfedd7d6edcf29234df31220f265ea519660f0de0ce1c76a5f7a4a2c191912f
z926ae93fc27c4a591c943b92c56b630e436be8e9aec903502814b003403bb44b6b3766258d821d
zb3cc1c26a226f43c1bc705aadbeebddeec9e48301b6f67fd92e61e03531187239d2e962551a6af
zc3890fa7a43ebb426e6684b17d268781752660d8316dc40fb71ef572d08fecff01e43fc87c7c40
zab02b0b002053115ba0713136505e71b297df716cc879380edf7ad4c4ddb3f274dc36003c01d10
z82366533b43bb2e7518ad9832365582b3c7bfcf03cfbe819d9b1edbf7aa43dfea62cd0aa58cc3c
z326b26baae01de50d17c414ab860eea13cb2f75a9130f2047a26697595015abc3c31d28372653e
zbdff61d0e7fab5dad0c383f4735fecd7b20e3dd94367f087f94eecc2a9d576044722a1e0c50a0b
z04b96541152a9b251775d663c470d591d28926f4d9585b9b06d47521b172186fbc428346c2366f
zb327ef44546261d5d9ee71e10d650888b331a5df8f914554067ceb1e67ee43f9c5dd475dffbeb0
zc4ab3668af9760e306f93c22e9fc22445e390b6f70b3d07f7629378202388357d08aae6589e6b5
z8e572540ef091fd77ae19212c058023b26968a787f677405ca2a830b033dd7f861ce682df5fa3c
za3658233aa9166dafd9b5067823502c99812cc29945ad056a8bcc13be2e75419f94c870f481e6a
z5c2b71821ad50c2cc2b4354213484f0687fdb41b4b327de7d27398bd299b5d17c9d660d021546e
z78046a66f545a7ec4607c6fae7d95cf8eff72d6b7e32e5f2177b471258bafc141f184bccf0273c
z6a117095f65b01ad6f7473bdcb3ca4d96e10e4f9166bf203d830db5711dc57230dfd8f257c4893
z5d7fe12ce4112d4cfc0951d1f001ae3ae9b581b380cfe3d5b0849961deda6202a5ed58dd7b4711
z4f407d7628c181985a3c77eb0df06cb1c63a07b736de08704f9791bb3b439b3ced32e5a27c62b5
z4c00b9efb6bd33df3ad34a7320fb4faddfd951788a9a90222743b733f31437fcba6e3f871423f3
z11817c8deb3f9ef3fb44ede2c557a2e50803c15cfec45d110a2629d8a6afb153e216817f978fe1
zdffa8fb74163afd502c876766d4ca932575e3e633503f652de6ca00b433148793c29e859de3059
z34e1bdf8e10a3f5d7c42b2d772ad87b60aadea646a266cd05eb5b0517e2f769985a5d016fdc28b
zd6a6a667328e98e4cd30af788848af57c76bb32753ee51cc241a278878dae7ec1fe03650849be8
zc7b8c243bd527641c76c3cc83d88006da00b435152eeae00aa1ac026ee55cc4b597345e3b4732f
z56661dafa3068b6ddb972c64d537bcbb1d23780e63f2e52622f8fa9d2cc0da2b8bdc84d5bfb964
ze9cd8faa00e840fff591b2291473fd41076d8cc439dcbff46d491fcb0213b6f771aa12f6739f81
z7a141cff5db8e3d7172e0dd42f18f26b051f18c03b986e4bc63b231b1baff830449c89097cd30e
z446abed0942032defc4f9b80b804c4dcb510e77d37bcbcd4c276d647cffe71d4330eb0434e0618
z4e9ac0f41bb291a45d49adb91ac71a211e212f66d776e47fc0a5c8229e4fcc1ec6b0dd28771253
zdd9225a7704d622f6b4e8eb7263b7303cfadf16dd3b17e3eed562bc2f873cb27acac9613a46770
zd44eb0b2a73674f6b37de19e21b3fe7fe779da181ff65604456667791cdc5a9edadb347d061992
zcd5037ec241783ac7a3a14b0c95ffbdc8180442158990858077ab9d9cd15d23cf441e3abe1bcab
z53c2ae0b07d922112eba4f011f17fbaa2c6290ca71dd97e83ec16f9520093863086ac9f0020a23
z24e223544065062a7035f7b1f543a00404426225cc9d9557c6d04eb7d8a1859ab73605207e1c0a
zd167e77ea4c3f1d0148740715489813668a7c91eafeb20f7e8237a2b7399a1fcf04bd1c35c60a7
za25d136254df14da65b4cd69201ebd1a7ddbf9c879aab93bf93269a35df44d843a21ed87b691d8
zc048c919055381b49f5e11655d21f42b6dc501e7fe1ff1a99d5e2c9110ef8e12f1739a282d268c
z788f10d23547dabadb280859711a201f7083a9a97b047dc22fc57a5331f1f389ab8e28654ed55d
zf69e6b1d549bcb443a684f0d51bc8a99499a94d54047d2637766600f7c3fd1e343d66261a7df03
z6bc2c18ffb54f86a84ba6e24399382d8dc6e32c198c5f5a50396e6ab5f9d6edadc542001840c30
zab93de9acda0c08a2066d923a760c6d355852268729fdfeb5ef6fd73baec05dde2b938e956b42b
z52ac82c6da033fc1d3c7860d1d04ae2526390db43f4ccfaf8aca1cdde13a28f559964bfe38e23c
zf4d5034295c38f15b2c21fa092482479f86f13ba9bdd699e255eea0f152a1ace12b3be4622e2c8
zaac380dd1ed198736ea28a8432981c1d72249d3ee2dd79a1305d34e2ffdb4c483cb32297446806
ze213b6c7961ce9817f73fbf0efcc7f09cf5717f7d08b0f220920600e6fef8bd6ff1aba50ed39f5
z0593fa7f81d3f66c4fcbd704a4baebb9f89629f607569d0fb2b4832da80e8d9b092cf4773444b5
zb013d20ab771387eb8919269ada1ea5a1f415d0da4f74c41ea3690adbb9e4e8db78e77aedc9f59
zd6c0a76772e94e01647e6b1ff12e580f6fea751a39ed9a04e5a08f7325e39a39c21773115204f7
z7e94180c43bc989891ab90b8e965daa29eb500763f52d7642c6cc5da4de2fc9b03a72b0b7a8fc5
z95795a73fe01d0b187893d570a21c30ff38a6d615cbea5da906b3a4f416cb35b3674b80b34f3f9
z27ec675ae185e07a4f216431a30dabe017f8a53e1d75b886602acef59a234b0c7866f3730c79a8
z68c6f0b31894df1d4de8cf86e3f4112780894c09792f9d848db7b7bb723a7ea296effbc3bab7c6
zd13809332378c27f7d929261ad793c75e74d618947830054eca013d19a3158f96fe8abb6e0ef99
z034ffd4813a8016c6fd9d7389436996b888db28fe2e8b6932ea5fbd38e8816e47938045d5572e0
z5d734fd97e333eb04beade2780867b787ba6c2251a3879cebcc7e4715d849c701566a4279f93eb
z1d45081c727f7b324917eb20f14f70782bfae0611aae0db303a07203ff9d6f2ba3f24bf451875f
za6046cf23d48160ee85c15c5fa786d591a077958546d2477b628d47f0ebbd5dc353522c87d32c7
z51dd7de52f92627a3b688173ab6e227ab9ecb8d7fd293ad9841d52a1faee7c2fb0371b1772ecb4
z892fcb434844038ce6aee690369fc6bdf09964775d557e5667a2d4eb1c22748c75ff123d023314
zb35208c58db8b0aab31a909803fbed3a3dc8611c9017bf32ca12431c786368eb9b4cf904d3fe9b
z9dd68c122f67bdd68fad70d8fcf4a7ba9941b412d41cc8463584f507c2fac4022445b082b7c3d9
za9569acdbfff2797587bf37ade7f0e142ca30a164fd0a23ab2c61b2f26ff3824285d834f9f571c
z6451133839c5ce0c8d43d3791081a4f2637895fcad18da5e10bd64b1d69578aec0651c7174730e
z6feccac7811d0aec42b0f1909f31cd46be8ee14fbd668039d7368acb8bac855fdbb3df76f79769
z9a99c903ee37004d71e0a14a55b21b4f09b10f496999ac7a6a51eed746018ea8c7813a5aff04e2
zae7839ce728c35220c5ecb9d67bf1e04190b8b7eb2def2439f2dbdaef5dccb75788b89e043e818
z027764fd046e478869b1f4dd9b8491ea73bb916556734e799eceddef8bcd3710ddac0d91457933
z09b6ac7f6e2bb47434a4a5b95fab3f0704e21d2cc1db07d829f9197abeccf0a5912344a103f412
z22bd8b266b892642014b15e8a3fb09414bc8662a0446936b726adc601178709403fccda00ad272
z59aa0878681a6fa39020f6623d6e41e008f465e0d7ffc89976c2162a22c643de9e60fbc84bd7fa
z5665c4840d131cae51befa288298161375f255decdca8429ce0e53fe3fade510aeb184910dac61
z33d03a76ca83dc0514b8aa2b42e26a4d548cfa7f6da5c76b9a21e8dd4d806209c2029b7b333a69
z1b70a4d9314819b4ef988709b5180c090be847fa533366a838538ac75eca623ea3b7bc6fc9cbc6
z96c03553aba4a7f1e6bca14cb6eb4b1198aec22d8b99c836e19561f62fe63b6fd259aaffb0e339
zc83447cbf5cbd4e6434cf1df9966c880a6a51c0029c3161c50cbb7ba00284b541e61876ad090cd
z7973ecbf6c0054d2555997e8096281eb7a8859d15a9343232f8045f7f5cd2dc8b5141fd3c6584c
zd98c08ecfdb35ec1a1992f779b2edd453c869d8a38d5bd7cb993ac24bd0fe1a4061576b47b6cea
z73868fc86a349d0ab02d60f86a084dffc2321f0ac080b43c48d2e7eecabf79881ddabb5a284273
z590f7d8e1ac16380b85d49db36f7743cac74b92282dafd73f6649755dc945b3cab5d32e67096a9
z3867bdc38473181560dfd08e1e4a905d17230a017f79d1a1cdb99f0b6635eaaca8816bdbf3a03f
z8777c7e8d60e2de41e9153d49c40f536584b6f81fe6b8069985ea56ed48340d0fe61235d1c0acc
z54dc39dc5889e7f5a728b92c6ffd0be48b89f1341e43093c685b20ffdaa28af793fbeb8d91a995
zacfd5525b305845dbbcb786d004fd7e1b27bc84b1937ca3f6cdc37374b94732ae6f22c70f1efcc
z49881350535c15e82e387614c23f01e2b4749fd72366bb3da809b618ceb936e484b3ec0a8d8ef6
z43db96a0b0a9e156b6075be344c1feb7bc0f551df2d5117e9d34d39621e7b501124cbde07a5485
z83d12fa218f9f843603bdfd17c61da211672d40bafb053594240c172713f745a2f5b2ff920352f
z1ab4b0516faf4c5851d7a1067113252564287f1ed3338e70dea9022da31e26bb3de4e2963818d4
zeb505f7777f5e72159425ef744426b2a9b4bf638e9c28e28e5d12ac9490b5efbf369ab66a0a59d
zffb3fb8c30e082b3254492f250703a0ab1f645273de677196491bb69454ea99db2868d57394adf
zb80b0fe512fb7bcab9ff784f1dcd3face2d2cebe2a9472d20396bac6298920adbd1e01b46147a2
zfa162d4d95a7e0ea86ec4f62a28a583ad33b20fd048da1d277c99067ecf600492ef98365e1fcfd
za01f572f9ce084f01ef58e404e04e4c13751b8699c500c69f770008e934f8d2fa0645a36f9012d
za2e37a631a428b5e8dc2746f9499305f9aff4ecf1469511edd912f43821b5c924daaee170849a6
z6fba8fe6b44459b4eed699889c5f423e8800ac739bca46da553a522bfd93ab7911ea64337c3da8
z917f1a9f3662780ab6688f25dc4c74bc36c7f610f87cfef3e26e4d126795f5bcdd41035e917b7f
zcc4b5284ccb561563d82a9bcca558cf4adf867e818dc626fbfd89ea00045887b80a3bfa10ea067
z4e56d8097f14b645c7b24b5083719e480d34a678b03acf1bf1cc982631877769fa73bbb692e00b
z8af1f5d11df50db8da00b836bf79aa9f3625a28806626b3d3a936da4318e54aaf0f2e92327edd6
z2083a3a838c8e5eb732986b8da25f08560d7fcf8dae4102269acda715bc4e96a31f5a972643e87
zf612d8934812c95016cd9c0a3c8d10fae93ee5d69e6d0dd9bedd6f8fd3b14d377e3e8ad449b442
zf643f83bc75d5095d81865df3a1fdd213920030942133b80e8847a308517003be6887a11a7a5c8
z0b945c08b3227e23048e064a89d4f0c5b144dba43c60bee1b4c84838b1582f274182b50857837b
z8f8bc3be34448b6b33b1f0e2305d30d9f8e7552f1b03325ad97b4441e565652a359c7f877b487e
z95b6bd60699bd3586a9d789e882f9aebb0528cc19a74062ae7eb2d30c2ee156f705904b88c5901
z3520c6f6a6f343e1a334522b534c1e7d68b85d6d952b83763111c98a934efefb4a43ff6fc7408f
zaf28ab49277d79a87cce0166b1411b75ce9cd87407e513010f28d8bc64b876480af16c6cd5aab3
zd2b0ef7faebe2e8a8ca77db1933a42050563adab77429a2331da58d71dad9a6055703f3164f0a5
z8c2aebeb9406fee984182b048e17f6a9869ae47a0a68a2aa0cc87dceb943b2a4b714e1b1beb92b
z991cafe78770f3e1080093c4abbdbc41f7f443212a54d06832ad3ed335a2d595d93dabe73b9c40
z15c7b5f1c05df7f5bcebc568370952b026051d8ddb86348f3965eb88eeba219d88acb568964a38
z98a6b536364be6b899b2cabcefecd07a0ac95f189dc14baf1c5411a8396cf4ccb8da1045b27ffd
z187cdd9ad78be109c4dacd231ca393a24a64ab8ac0b3420cac87495f9ede583b6627fb9c7ddaa6
z54cb56ecfbc7d63dcaf247414523c532e233ac7702910a9ef01771eb928d52e794ea4c10671822
zddec9815cf87ca3d31815085cd19541341b14bebf50dad9714a4db26d79ea308d8a5b5e80a6675
z4ecea3271cd6d11ccb03fa06cf7eaa22a1b5dae327f5b9a6bc1cd99590a4454d33bc59127f115d
z1f7ea05768233d5c3e83afb4ac65b6df03a5b86e03fd378f28b8e6e5c6f030c5651a6d9dbaeb55
z6f7a6242eebdd46d0e0483fb56f0661053a6ceed5bd9c024c083937585912ddc0da23f78324df4
z5e6d8f5159e9611b488f563f599b421048d9876b2d8cb5056af4ee1d2c60e53e498f1c64ee5364
zf384277cbff59bcf6c873934d2cc4f8c8452129edb633f8606398061c4cde5e02a0eb133551302
zc36e2d97f9f251161b4ea89c48a604d9ce42f827910a23a04e8a9773e52de28f993969cb6655cb
z125464527cca4a9b730c205f9c232c16b551d93149a0fa7d96efc53e087ad5791ab2a53ce12d64
za97ab605e2e5090597163128b4d670c2d4bf0a49d218e13e371e784321aa133038120cdf5e5945
ze355e7b7c8117627a3153852a18532f0c82137384333b8f6a72eccafccdef43d227b718a9975ca
z49582884fb5a39b1240ec548c68ed61c843ab4c2254189b28453e7e35eb25fdda3a34e774fc6a4
zc0af9f4a4d9f93919615e3ddc5b21c08178222903654d52029d25398fd7510fec2abe5246b8bd8
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_target_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
