`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc3904db24
zc5b0040322f5de9957e599cc6ff91e8e44935f0a5a0acf9d4bd50bb5681a15ee023b036c0ff87d
zd437147463f5c5bbe42de7b5ce2f24268118570f4fd53723f426e5dd3147a7e849fec8e8709b2c
z79df24d548592501f1b63aa2a90df111b468b329fc1e2e276ca5da4d71ece4625205df608ffe3e
zdf262418050e8ac492a51695bd1773d1c2911ffc50ddb16ca0cc95b867c3fa37087f03b5a91143
z02135f2212fab57548136fa411aeb3ebb25f0d1bc0290bb0fc55f15b53ac06bbb2eb04eaadd20f
z77831a2c3cfbd539ff67ee08bd2ffe894a5fdd7136992e0451946bddd7d173caa223cc9ef7afc4
z7a5080953e4a09f5805f1132f41f527f7f40600dac65fce9a87e6900b97470c34047afa2bc2034
z6d154b32dfed0cea6c2d08d5fb2e3a321a2b5645acc53a94bc9e032c44ba1638be78e3d7d3ec42
zda7b74e2422ba50f3978caf2955a2935b3fd9f534622265b20d0f236ad220d2e07f69a9b7a3bc5
zc3bb6a85f7e97ee3ac52b1619bfd5e3b85e5c7e312f97d494fe387fe4b6051a195ae74135a6d07
z41e9443fa00d87ce8b2715b724d16d337742830f7b800aa8e1c1eb7962a59ac42b64a9168911ca
z4939f61f22d282fcecd59cd20ffeba11a410a30625894a5a5ff2fc9d7dbd50eb0de235500d2e34
z764040a2ddcf250e3ac0e70423a5aacfbad36927234e73f8efa787335ec059c44866607ccdfaaf
z96a539c7d2cd42e0af0dd11ecf80e8ee36d7c4075ce8ab8e87833414e8e23eadeda447a4e07282
z225762b9541e3552f5eca029079dac028e2cdad25f451146fdc93b91a2ecdf5012015920d1b235
z8dcb6f6d6e5c665757c4a026396e44e92d6bc5e90bdd94402fb5630562ecc29620032447722d94
zb220d9fe76d599eacee40d69044f263fdbc07ac23135d06adff2de797ff7523d3e7e6ea1fc2143
za86df32b5b9b50e556aeb65f5b54c1407749a52e37ab3482e7fa415e510e86b1657a3cbca2deba
za466572d49757c1f4e47c44cae65373eb745fee4a366f31dfccc440a8f94518ceb04fcefdbe01b
z1de238856d30d42f7c83ce4f65aa6fd03ca5fb8cac34ddfb746be7aca5a00d69a2e6f4da862330
zda8dd64448e84a70900a602e21e58c7c74cc9aacba01b6c0d8f23273d7873c3cfa804469072f2e
z3cffdbc1b665ad898310d16b8b36c71d17262a7883a86b24e5184c7c05329a59cdfefbb48bb572
z7bd864fefc928a8ca092576a645b6eb2ab9785f699775e7dd8b5386319d23bf4960dd2f52215af
zc8582e41f4fc6fe729328d7069d2050f60c392986b5469ce9c6151580995b0d3a1617ff4d78254
zf6cbe88917b4bdce492c605fe69febc0066f8550a099b8ac0d0ef6b27603f871b650aeae32e1d9
z7fcdb526b472cc3a907d91e0552291115596ee0781ccb8f71193a73657ac0d0a6ec2552bebb239
z493fd2bc3e2613b9942ee6cb9e5011b1bc3ea240f65f370eb7425eee9743eef867a9e29f1bf188
zd0ab6ef86265bb38e49cb6b2e844edd089d1f6c2f6149f5287f0118a543577725ab4059bf5c404
z91c15f9e836b9d1c3747526e01d5dc8262738392d8074428af997beb02c3ac8651a75cdd7692ef
z143e7a56341ccfac6505d53d3fa9799763135bf56bb80ee09c37a3d2840a0f23b6f9deb5b12d8d
zd95d232392664dde85f99ef88b115bd542bba959a7f67d466d4d5dae48464a8e984d197b97e30b
z361a1f45143bc629f73c2b23630dd87d7277307aa367a85aa3a3ca7ab90c28267c39f61dd68739
z9d22fffe6a5c845031a1fc99108dd07d7e37229b8d0a297de6f1a9b11a9fb2a2ded5e266f582ec
zeac560c75269c4ce22bdfd28f11263aebb13cc23057b4edb6fa30fcc3bc20a1649a4249e505859
z0fbb52563032dd812d0a0d4c00ef5a903e7f14d8fe9e8e94aa06e547522ce38f4f1518826e8716
zc87acf9844072ffa9d8ab7559788e4b6954035018ffa714baacd39dfbefc892192d8cfefac7441
zf72f0042e676b2e7d569647b90fafb0c9598d6f02be84d36fe3ad250510240293562704999c6fa
z8a5f1e8b0c4e0bf0bb916efc528c4b21d45c8a846e0608e1375c9cc0a20b5c3dcc7d31a97d7d8a
z829b5914823c5122a30a778844ca0fd53743508a2ca25b99ef8ccd7c9b8275702d80f4a41f4cb0
zf3a6cb42bfd8f82663d413e3e35b2bc23d29f70bec6fc43c6c970e60ea7b1e3d1072cdcadacc2c
zea543e3906f028dd31218b872cca03f38b9061b1690ac6b3f460db40d32e594fdcf363d39be120
z68b8d939d75877936e19406eabda1562f239f51abf223cb00b4c3636bf544d1c89b29d2f66eb79
z1ced6a1f529c8dc00c2a8eb27d25d99c5dd5c1e27d5a3e1666f7286c69185dadd4f17a3299e2f6
zce416b28e9fcb53a6faa1132495b0da2e0ca1e29657bdf91d8a0b6ceedb7ab481f82e1aaf268ad
zf338e2e06d006126017bcd9cdfc1a02636abbe68e558559d0a06ee9c96089b57b1b7e92d2aafa1
z60c246ba658058a9ddbc7aef71c9170942aa557e3560ce15e9187d3aa84329117ce8aecc3eed58
ze50805ad5424e40d34338d0cb8ed9c057f11ddb2464b6ea1f877a73c2efaa88670ef8e4407a97a
zcdc027004cfd7e0eea4ccbc141b92ccb225eb6aa5b744eef4e40f650c6a891cb38fa58c7e346c2
zc6527a762d3f64bd9cedb0ad9ceb3dc3ed3e2e2945474b753dbe7bce9b67c6d562acb778ce7f08
z9a46b4afed2d31aaed793a23c8e7b5d543a3260f3fb9e0f9dd69070d48662f41bfe9ce2828afdb
ze866ada6385a8e8144637081184b377605a2d42d0b44b708397858d39ad16f49fd63e062617c4b
zeb78c136a5dd47d33129ed3618ca8f2aea0b5f0d3c6a83032a01cb75a0a3d947f3442036574015
z8c6909edeaaf16cd44a9c51b4537ccaf9ed20dae178b73668f3ec0d962db79031595f08679798d
z7c9c82c7109fdd8b88a7cc294615d187ac537cdb601c77c4cc2311cccebcf9c00d06670cd6cafa
zd2b387ce65aa7e541b00a42c6a5f7a806575fd84a0bdcddada3c973a9e32875d9d55d40d8a4e3a
zf7f6b8d0a337f05fe74de8b2a7bcb784ce5941ef130b909b39af92783b25343321bf03f8db6c41
z2cd595265ce4b5085ee5a52af609dc795e26606460b6d5fde3f242dd4a0ef8d57843b676a72ee2
zc855d902fc0079b451211c4153f6c9a7f41e19acf89a1ebdac94acc60f7d32819495f75e2ba593
z805e360d0b1cb7a56750428fe4e7f5cb22b1c780fdbc4acd75bb47b1bb3f1bdf2076e478f7139f
ze00e10f865b399ad073c069b9490557cf605b862bd419124c3d0c5bfaaded1c5f40fcaec59fb97
za8a4638757a04663719a2f1207ed2c196869d038759f19c7192cdf87c9acf9e10d02bb0ea44cfa
zbd979161b794dcf4e83a68bb025e557bdc2626766fb16839b0177d5e327fc56dba27febcc99e65
z473a899ca1fc277f460b5a3e71d1ab44294b76e69493bc02fc8342fd986d25f2d639e597e6a760
z8e77972d50e3313d2ebcc612c80f697ee3d6d68224dd2bb6b98eba6ad99923878b734118bdc39e
z55089029b3dc8b7f39a9a7db2af395351c8208bd00895ba4947ca8ec5e96df7f694bf100ed01a1
za091416c652d85903474f355836dbe67ca5628cb429b8abae0b2d6c941c6cab5c9ea87e714e58d
zbbf52a1549005b15e8c414f11db90f9b3f82ca8b9875d57a2a0639347a05e70d294f021ecf5ceb
zc3ca1df019fcf9a5bf78f9f863ddb831f5fde62f4662df03febc6ca3419188dc92715789d643aa
z87b929cdd6b050733b95d4745ef64dbc89bf40f5e765a8973eea47552e3c9c852789ead33251b9
z06d4dc3c291190478da54c76b639854dab722153519e3abe01bafe1e88df42b937f1e50ce0df26
z09ee40f612fb6506c1205d90c468bcff591eeb065d3c79123bc2a31115064f1b825f8235daf8d3
zfb886cbbbad3d3a93edae971b486860e42b2ac8e4c25fde998bd533163be68c1de0bc49dc2ae3c
zbeb066f6f5e4761cca75c8acde99402b483ef250ab83392992a944e9a06ae9ac622881162a1953
zd191fa20ff4e23330fd2bca1603a4daf66e5f44897521690f3ec45fdc0c42891ace9a38ea472b2
z7c8267e52eb721eadadb817217dc2eebb6ab74adfb252d7fc137f135a16917f7f7cd2478a83cbc
ze9d5fb050a7af4dfbbcdf320f93a63290ed62acbc5fb76aa116e15779f2bcf5502ba3f6024d9cc
zf59c8977bfe2c74cf746e821aa17a710a2be190a2d5139d057255b3004effdf5e1772d46f570dd
z0ae06df043eb6ed90a6d14c2b802c19e1a6adda6e18bd0843117724dbcdfc3a31bd517603447c4
z6b930e2345d66935ed5851c2daade7f17f80b035c69b3d64b6be57c6878d065760e7e31b49ad42
zfcccc67d5d90687ad865fd389e67bf52f5c1319f26dc2e93aab5a2e3fdd41f5e4b7667509ee544
zb05c0b610472b4efc4df0deb84e35d7df88c75989ed33f3ca43a14b4761cc1fb1f8e6eec1e1b9c
z000ef8a876ac9a683e0c17d04424c01fdf1ef351de7c6d5648a6c0d02819c339f4205fbc02516c
z03a9c2853d639caea5af47e48f75523350f494edf138b6feffda09ff3078093f80bce835ef485a
z20808d6dd20d3bb3a33131c6479b4e82b8520720205d047e27ae377d4d20f42034ff4fcb542bfa
z535147b9a59db1f967b9f42b166be1f659695bd1ac82dbcd462854ff9d3c58ff7b6b6a05c517ba
z465fde5b89e986659ae35888f0e9bbbec67bf3d8a857f8dfb1b38914b3c210878f58a13a0ef906
zf61a8ee0c80bde7caa0a1659510440ccc6fea9ee8fc64c60a6ae35945b9d3574c975f091b1f2ac
zda02463fbe43d3c657d8e7e19ebd3965e9eb0b0604c3a9b0ee10f43c44ca6c7373d841a49562e8
za8b1490d287f2604d0270781160348406ab6110c29ca962f91a574a412ef895cd911d57d79dad9
za379626db6ce3a97e3d5d5cb4d3b540d6ef20539465bf872d3dddf6374f4f10db725945a539d31
ze580556ccfde601d36b779be4f76c773cca873f735ea1c21ad92d46b3be021c0e6e3a2c1af8fb6
zbd295aeb481a115b827e3d81f54c6c6a032efdc47bd2550f3657e9a622ad3189d4f23b422ddf5a
z2e761ac4db336bacab2b3453362ee276e89c42231cd3622e4f71601c496348defd2ec5413215d2
z023e630da17d9a2245a6012e41bbe7da6804c25676a64c0f219d80ffe43dbecbf6ebe484d9d803
z01381516fada6b83c83060cdf586e9a8d099e731df7833985ff4a21a08d5ef322158ebc29a93e5
zcf8f3803da02eb9cf222a875ac1dd0709f2fbe9b4622246d3e05048406c47d3a22611fb801196e
zb95536459e7bf97fd0b8af8a72063187fe85efff1db95b90cea290ee584b3305688d6f320baef9
z29c9a8afd344a9db62102fe4230e42799d66fe47834641c77e6422bf2b06d602c21f51e3e1b96b
zf1d1fdf159c34fa461263c3f9c3d2a5ab4b587cc73e988bdaff6ff90aab5c5d32d29fd790eb2f2
z9ceb4d0cb9c214e49d38d5bcc8745d948defdd02828db3365e75e2e53394ac77859b7f7aefae5a
zf2e4c0991641d5a7e06ac68de61bbdeb958a0278aa6e825c14c7e6f72d64b01f0cf611add4fdab
z48c63e2d87b868c4be5189f89fb79e9ba76e197ea994c89e9506aaa2ee9cfc66a2a24ee068d1dd
z297bb47da6851d558979d1d6b8347cba2f579631ed01f2260a57ccad7f7f8a03ca32e498da547d
z5181d0fdc89ed6875890daa0d35220fe9747fea81263a70310cb2206e103d2f9898a8245468aa3
za93ce37a28251618472a7aca88c5af1abc2f934b36f861f85aef68765eb6d12e378101e00255a1
zcad3081adacf114a7660524cba509bb973b35916e0a1d8d01a2a49c08466f3eb7ed990f2188ded
za730933e0cd34995c5bfd6c183fbf0392743da725f82557404197a702c4263639ed891e79c0563
zcc55dbd4958265e0f031c1fc406a6d4f2e414a38a612f216fcbc837808a60baad720aaa60bdf88
za2b8e4b22959fa016e2b31f6e9fff095b7e777f62585dd1ac36752b4b5d802f6073339d1099fca
z4106bbb1ae3eac08fc9671dbcc07354d20dd6b8732282c0c4afc3b990c15cdc8cfa4c0d05872b1
z7539fc63d67ae4281189357877d9df9b7ca7c7947e5c7a965f218bd8a593a13e754faecf345059
zedefd1617afe7dbc851a9be132071b734f070a59fda5937df54e136fcbbc5e6d4a2a7d21a448c0
z32349eb27371fce054d935b4fab2e2768e8b45f9101ae241dfb69cf28f6925a460e7be7347014b
zf651b326312ab26a37def999be4c14a2c35eda6a65045fe111a926105007c589f76375453c10f6
z790f82b92a131bd62303a51b061e40781610842b82f9b81fe4e15e72f8c1f302729186aa6ef1be
z6731c2f7610a96d550c913444a3ddd04b087c8018f99c43d2166762d563380ce1a7d43fc0b78d3
z03f7782cba22890b460b5fce4c61c624580b47353ff48763ca68ae0f46b0fff30f3d88a581ea32
ze79696df2acd138ede4a92a6bc821607c8a2df3ff1f7ca5a34e4a0111586ead6cf04aea9775d7f
zcfb9458c007d1519dc22c4141aa95433ae754cd291e7b0cafc8a5490d372967482c2a51e79a276
z85d3ec1867a899e384fcb86f98f18693c7ddd7319a03d9e4c0ca4c592455b7a097ee308e4fda98
z10691ab5dc198f7eb756d8c91cb9480609da66e771f0860741c2af938dfd764455064d01972ed7
zd5f4db31f6d7223170db2bb014509899f180ad3238568ec5bc5ff16da4e743ba702bc3c950da11
z10b23a87991f61da1dcc7ad981327187355bb8fa4fe53f5fde34df9fb717323401e81af6a45aef
ze9c0b5c700b3ac554a011be97be663b1068457f3f3e408b3270fcc990a4f78be85cf7121c965e7
zc886c8748c7fa4df7f395ba62b457cb68023ed7fa9b85b4f173dfef7d905033bb0be36401d46c4
z32001747df5d57bed620502704321631d68173987a1affff7af1604712bf111826227081c6b718
z2aa20d40966b4a13bc6d4b3ac93720b5bba1d6f5e50f84d2612c27a781b98082f99919593154ff
z4094331aacf3a643e82725582e05673a4b8fd88d7a1455294b00899bccde13e965ebcdafc8aed9
z4c22838f9ac126911300c4dbd0ebd1bfca3411c638bf0d7f067b94eb37ad11655acaa586cdfd07
z66d9a3788529539edbc896b8b6e81e6ea0ee78e761baf2a951c4bf958d5301288b45d185ec2150
z2bf929dc989aeedf885dc6e5c53ad7145f9638c7b3cf3957052e1e9d0723c3f66a00bfc1f7cbed
zaf4c07675926a48b42b94e869444eb16a264f286c80b9d0c98af002b7f28f8e62b4134e8485045
z0e9237e8147c54cf4e88e7bf299e98f7ed1f7020360c78261e2e0ca4eeee25b24be0cdcf362eca
z56487b0e53b7c493e5fe52a95eac33190ada8e00047a492a62963d37f0e8471d54958fe3fcd694
ze83c3de7f8e40362dc9f8d85f3cc37c711c872a5595588dbafa598d396b3d9f680700d4f6a0dc8
ze461a963a35c2d826bf5bee3dab29285f8995869c3e54b0b248e776089baeeeb00c4c04271db4d
z16ff46941a56c452ff318ae7a25a7611d5ac997942cb68a86175b7c250c1530fb91f184876ffa7
zc5ee74ab07081da445d45fe38470c8a957621b110fb6afbff7bea076cdace4638e14345dadd828
z36cfb9d2e6adf6fd80f17ed9601deaf4f0d6ca0ef06bd1bb42c7393427e10d18088e436813b017
zb8324f69a8f04fd877948f8fe95d747676b99512325178076f807d7917b82e2f213efd8f15c327
za7de6e1994325a5ecb3f3d0f5c33ff93707dbd06bbbe73f68a8abff60c65f14f190da2e3ddb719
z076b8c8d74c3b02450a8318c5956ebfe21569d90cc7a646281b93c9d53abee2d1caa91b5cb6781
z46c0b54e9d437454023b67e21c1f9accb0e46c8da1917cddc9dbf7bb9e9babd7e35a0be2ffec04
z3049fabb1797ca5174d512896b7103c22a64d512bfa0792e14b4da4b5c407980a5499b4134d0e2
zc0c3d76b0b697e30cfd7d8174ffa555f1a478897d6adf4f1cf85ec9c48af7bf819ce35f4e05b4c
ze5083ddd8fd5f3ed92950e053285f45ec0e3048c791e4f2ffd3e40e215716bc0fcf9f8df4e853d
z6f5c3bfc9ab88b279cb2f5d248c314ac29b007aad9fb7e6ba4fae5c2562a8340d8533301451939
z3c5e624eafef7995ed76cbaa7be5051ae1d631302028979541e8f3beaa825e54b3fffb0209cc2b
z2fedff6220cbc6389e81b5ce476963c9f8ac7f09b14d81a8ff56a8f345d18d8777c811b1f45f26
z1c6f3fd1404cefe334f300d7c6b794a67c5bc208f2c85a561fab98926c04e62490cb3bddfba330
z221e6706f796fd0d21ebaac69ab373c0da6ed74f0d48079a06d4590dfe629d6250b8cb669476dc
za01555c6dfca462adf86f1bc5ca1ece593dd38036c7a2757d2745a9a2e38b835c782053d8fe330
zd972866cbbedc12a33d3c75db65ed226a6ae0661a8517a7c7211242b15a61269b10ae118202576
z89d958d6d589eee6732573429d9fb615968333324e5837442a1c2d07d2cb4b399022a34691de22
z4251f6c98d9b0c5decc9647aa2d13a6bc543067c8c3ad5f871c2113b7ded786c5a83ddcb511de9
z18155f9aad55b853e00a2c5b1c2869038214c0f6079645e9b3c0fe79c441dad49f406cb2cd4b87
z3e7242ae06efc39bb12591f218748797388ca61f5509328c3ff9e026f397f46911f60f192894bf
z510ac201293943552b34e102e7cbd68c11df7d32552a814206792deb0a2fe7a7a0a3567d2ecb09
zb266497a25268586bd7198b55206b57c1c5d1074c1f38eeabc650316a291a3835345f94b60cbb9
z23e4b729d94940e1c27e649fa17cc20379f49c64e79777bae624cfe935a8ef393dcf61c1a93da0
zcc246dd8ac5fc75bd8481cb8ad0b556564083d38b551cceeeedf37ae07bc9b21289660713496ba
za1503c7bda55e8e2e7f2033825b399884fdb0cbbcec223de2033ad2567c58de6426bedebb8765d
z3c4e45a80a2a1a1fe98d82cc87f3159ba521049d9bb6831347971a6186ede14b1955f3b5bd24cb
zfb2ff22106e33c6fccbfea496180758767bc30b4aa6d946906e1c0dd6eb23255bd900bee510d1f
z8026b84a39330a505733666d1b88a75c662883be59e53efc57c5492bf7eca350449efff3c1128f
z10cbd7dc8ef90c50b2b755ab1805d8f71f5b36ad78c18c5a749c75e218974ab5f86712475e2c74
z0774f0eeb0674ed5ea7aa1c456d60159b95ab2d69429271926e6c27ab2f76d015d2d7ec7166852
zef10e47a2bf897e2640201f5c381ec4ff9a714dce8221b3172d561e9b8c4341c33609064a16da2
z261ce649fc89986b76aa1fdd544ffa1ea4685059724ccbd500a14b801df0e51107634d59b207c9
z9afa8a8cfb6722a13be645d4b15a7b6aff94f84fcf4c689213b0d55e91a86c0e104e7e76b425e7
z5f5e3c2e8004446c7aef9bbd7a293627e4469b7fcd59343a50d96f6d3d5ca0bf08a64c9287a10c
zc656593c3efb45dbbfb6c38fc89fb46ec63edd88c7f13a2540be8bf8f2797201c6be4079c6973d
z626d5a4c7b4a7c0a30ab96de80860e8565e26cce5f736cb11226c860a161d878b1af93db47331e
z4928b0dcff137f12b40d25f2ed7b992ba2e5b6446c8b7bea26bb9bc869cf75eab9b926a14d324b
zbebd4652cddd644a8137eed9f874a1e986daa5a52130b6d4f1f8305f23e0f3cb08e820048c15c0
z6cfb300e1fbccabdbd6f5bd30e96a416d3249b39ddfc787d96e4165aab955d172d25f4287ca0f0
zcfa070d764fdc267ac70c4d34e6456449b3ba8ad6b34c79f46b2cf205dfd19494d3b1d18876aba
ze8e6fee892ea3d60886d34917f32cbaaf859cc98b6e7710bd5ee9e7ab90f9318d80902844589f4
z0da060dfcbcfb2ed837decebc4734bb47ec99e07c759516b7392aa4e8351893a548e176fa1ea9e
zaf380c12ec657596c4a083235388b2d5487e58c6185fb33a4fc18747cd2657e088a94d34b8556a
z1e655aad75a27c5887b041335480b0940229b6acc25462366969bb43f1aeca3845c79abb3a448f
z62256d10b3da11f3d726b8c37bbab2709c3f51690432b111e3c05ccd0ba6b62d2a2bbcbdfcde07
z224726b09d725c5cf64f82d53e8b57d24f6a15c3ae3ccebb0a4ff770ac231014fe166c88a8aec5
zadc7a11318bfe46e15f87e51e2cb83b8b96f798baebe1ac4a11525fb025176b782dd10ed1dfbe1
z7cbc3ea56acf1501ba6b4443b5bceb9ec3701ad78073d3e1a0c4b835f677e422a5e807ecfed608
zc356db0231bc77e3d83222d997d4a45e1ad894980046ee2d82830e80c00feb7ef93a4f733dd2d5
z160b0bffa4815400c3011064befb13792ac848be09e660fea5b41165ffdb178c9cd2c83cdc66f5
ze6ad889f41d8d29504fa0c4eedbe39f31f06a312a4f15e6dae997301d4f342eef66b003aa61041
z7c8a4687f09e4aac58f08dba3e05280fafe4537281c8d2aadeb267fba88a87ae920bf46930d310
z78d90a3c6f1b2c337a0ed71e330cbe0a77dadab43566f4cc055d889f65d10a20246fba191d676f
z8103c536ee43c44f823eaad2eccc849c980d150f45b62a78b84aef6feac5d55da3c909315bc53e
z3ab6ecd0d134a4388face96b746f6300b6f43e10e46ce4cdb77f6b45b9e1fd74984614d3bc4ef3
zb14c277bf52df2d9a06bb9376177c9de70ecd8696cb76e670aeefcbe339d2661054232c7529e1e
z19a4fcfe4fd87aec604be889e025d855a2676f160040ff89b899e0f630ec79d8b3e219b962e561
zde60b46ae3a911f4e7cbe9b11e42fbbb286057abf2343d4e52b4dbce093a1eb023dacb5c2c5666
ze88bd360840af43683e8c241054f8f2ec817f205701dd63b14f269122bed8e57b115d550ae0c15
z03ec0c624d22007cfb57055d46c618cf40e97c63adffa4577e976f37b6a0e0ee2faf19df3cd206
z4aa732dad6fdd6fe19c5d230e8b85050f6fca2c72874642022e8d51e8a817881d90a9346e5cb40
z39cc76963e4326ab9975fc1ac12f602cf5a92f7717d9fdc13753ba7d427301fa27ab2b7aeb32fa
z72eeeaeb74672f0505766535d89736f6cbe0221850d14bb96e27e3596146e6bd3f377f1e14a159
zfb59d717f081a29007b48ee885df83c0d3e3f1be197ddb095153586fe1453b95576e426f5a25f5
ze427d440eb760733bf6fecd30071ac31e0b7a87ff0cc2d85ba1e153beb17f9ab3d61cbfa6157b9
za02882537810b1498ba9b7083b501b4d834a086dd7183a7ab3070291970a6f579b7b69364b8120
z0841946d61bee85b87525d396f3887c9c03bfd9c522380048f63d5741b14515ff8a5380994ad1c
zb5507968b8801bc4412b43de2a750bfd9fa470403e585b9a19cd78585550c72346284201769da2
z7a64954681b96ef954ef136c52b185d82fdcd6450196f4d1c289ada8871933d148ad287f592785
z1084562b6c80705508434fb2609304ac1ede24e282289846b9415077d58936663e022122e3015f
zeb61d10bf011a4cbffccf8580da67027449c2546c6d8af802a145e34285a179f4807e6b8a1a112
z0089b03f00a7ed02b2f4337b4b45a753b4b916efe11d40f3d504ac2a14e06934b5661c172e678b
z298a6f0c2eeb15f6bb8e7890e11e769bba91daf44ce36b2134033ad48b12b1ad8daf09a3033e09
ze2abc25cad190266305853dc08d534811eb7fc3abffb09acd886266875dcce0b71aace30dec8ff
z4da9afdc605c3de79cb3f679d5c9cac79ae996665e30eea9b8dc08a7179e73b1d98ec27db1ab5e
z0101667597040c3f49bc993922eae8ddb3f59341e37c03a98eeed165891ed76aaad190280062a9
z001d307cc9726356e5e72b59d6a40802bcd38459d66f5bab0dc23bc02f9ea6cf5ab90ad6beb49e
z35f7bcf9eecc48d5b924a14d9a9796becfa521c716a85a9f61f1a5de2ccb35e263659e993b01f5
zd4866d4286ce98ffbe5b559f6ca4eaf1dcaebaec6cf3b3d1d7684307b8f8837183d259afa105d3
z7e3e7d2b707ff70c1456078085a767abd44765744affb5fa0791ad66372fc1d3c2d613df53cae0
z640416c7c48bb174775c51ed792389c6f30b3268a6b262db1fb6eb384b8c73a88e097860217c94
z3dc1474cc5a838e7c71cb44ee2c528ff1f5c09612e4cb1120bd145258a2a8ccd836b65a76145de
z2509f3c13a26895f267064c855f34fd8f0b13eea15d3b98375613022edd4b5b1f5309ad50e4839
z5f11ffe624e274b667f494c9b5ff3946b1fb044b681d709a07edc9b26017a0fbf5bed3f4c2d967
zb912b898566d9f47fb2f10d2d7d45ec56bdb5253fac7a65a96acc6d2367848dda824adad3e09f8
z533be9589ab4e3974901cdf94a1a4b7e23a7dc9098991c44a209bc5651996f03c82fa45b0595af
z91751dc4ebb5db2d339b22bbc82c0b26ff4e6d75874bfcb32fbc2c460404b1fd0ef6f6b227a0d5
zefcf2e8fc0f6a127231fad7b2ccef570ea8595f7e5214ea2b02fba21e20a59f1f3ceade1be7887
z725c1d0a1bbbe394d2e005c1c11aeb06a18002da62552d421559f1b35d25f7b5fe947a60951919
z5f6f781be11185298cf9fd4e9ad8e69ee1f5288b3fa31bb27f81fbb854a0cd078749c6b6d7242f
zb8ba6bee5f07c00d78b8cfa8ee70fabd0c6feee3c2ec94ff7f2fcef24654d185f436c74faa656c
z041788498933a966a082018ef64c34918013a5a773ae1fa20942b3c5a673b65e5e432b374f1634
zb440c776e108e29bd08a55b1d020376731f726cacba20ce4e3ace215ec5090aafd8e18d200e07f
z506ab326109f85deac08e36b12e60a985a9a3bff974b9e2c83d6bf5426a4c0d51f2a9b8f7ce166
z61f1342df5fdcaf4d61a3a13330df19b57a3179b6507b4c82fc50e99c632c6b5103d4936338957
z58df1afc7aec74ac7ec9120ec3127be4290ce6707814750d6f9454d9fc47fb1689f155089e3af3
z2e822cc07143465ecd0a58012ed9c4eed60b535af648f3d9d70694b16db8ea72875d987f52c381
zc925408c68c355264588430f3bbb1a9eee649efa834c322b2875ccf9bd97ac2b394fbd48f4ea45
z2c857de6d0cf3773e90881c0ccea3e4aa002d84af968d440ce986c1a95cca8c00899a345fe6211
z486bd2e8d31005f4cd31a9af4b2ce7b0715ef88182a97402e16c02ed966e63c6b91915362f1600
zbdbd58732a0461f8ea036f2cf4d9905841742db63f6da16c3867772b79158aacff1d5053213679
zd34463fa2d18c0df8a1855fb9ba56e41225508cc61e65c77e65f19c559d735dbb17f55c11e6c18
z612e8053e89c675d3bc4ab3206c94845f1b16a9cc8a280b78cf869dea01825ea1b5ce37ba4ff3c
z6d266557beacf9cb2b29c8cf6a0757857729b1049340ec455e38fd837b06e58e2139aba99b26b5
z4acad9676fba416902c02b5fe1d868d0c7bf1296bfc8686f378b2e11152d1343ee8f213d53ee97
z9c9b5d541865364716dd3459738fef803c5ae58daa135ddb2fe8c6e3da5e2315bf692f390f65a9
zd4e431274e22f749ab2b9639ad563711ec532a05f32dd4794ae8648d76526e076259a9313983e0
z039f504c67348d962838d5ddec45971db5693cb03e618d20d7eb8e9fa074aceb47c9e2cd787584
zda0985199aafa4770587131bf38051a623b95ef6002a61a990ac639178b12bff786fc72c2726e8
z5ebad2e1994f93394d51fdd454698b8880b54e120994c5b3d7299a45dcc162683042dfbe35a103
z61935400204e15588074d1fa7e4155d9cdc067ea4a30c98b2e7ca86b5feac8d6bab9b4f1983390
zf1f2748e90556a40a7c12f9ff9103408e15b2fe5a9071dda6e12bc6e083fa80389ef948a19f57d
zacb6a291142110e0c09074cf509e76b9f5ebf45e04e4e0bbe68cc8f2d747a9580884ad1551fcb0
ze98a4cc2dc9843dc03d99832bf38bcf91db3788b9468c020a010f9c44469626a7449d1b8415e35
z63f427a437a87bec8ccfd43a552eb4b644b73480fb137d35fec7a6c37014b7344b05cbf0a4d2d9
z8eccc97eb68e5905eb727db07b906a21192810a2e8d63a6ba26eeaac61492a968a7fdd547f2a33
zd0bb043f21e9f96551be415caa9efe97911ebf186104c62e25941508002f8a0cfeec91d926ed5b
z855282c5801715f60e9df57ceed42da8f278df0411349f630186f95e739555aad666f7dd1dd405
z0de351118ef867e89f391c0a8c0620af7ee4865d579f911e7f51b1c75c03ae230c38b4786287b3
z38b9707a13e5073cb8f9dd12c4c81a7a21419c266181b57aa65ae520adab83ff7851924c9eb8f9
zabdf1d7c1258f43ae2e34b4f1d5105dc2d0238a09371f886a4dfccc4102f930ede05aed868fcaf
z74da36b199eda25b00212c3c1fd85bd76ff5b61af1d93be974ad344a345fea674714043c5a2c01
zc395b6d57085d3fe5bd83f6ae6c69aa36fd18408eee03bfbe8423032439f631c49a143847df12f
zb723871b5838aefd76cc755ed1dfd14dc2a0afbfa2ce21030973a049c0a68005c5aca522fad936
zdecb769abeca570d0f4235344c542e5277c7f13cbe37e3d6a2a4e6fa90652c25194b38a9f83810
z6842a2091d2b1029b59657c634059feaa1d866239e6cddb36fd69a70d0c52ad8f434993e4a9542
z27d8a04bcbc186c6ddac108958474ed8e9ede93846e327e62c56bd9fc33169f9109db78b17ed99
z0b65f7269e8bd676e5d04c5712ff925e97b6bc95a44269f1415d4e99f8e383fb190f25dd4e905f
z52a650b4cef892d31f0d2506e59821e9b67b6fb29427990222124931a434bb91a9d9a96f98a7aa
za4c7da7b873a57f9b0ac075dd2d8ff8ee698e22423e0bd9a94b77d35f97661cabfa4e14dfe0631
z8c915cd3005193563f39f89ce1983fbd484d14814687b05d1077b356b9a8460675456df65a8b68
z4766fed624786c0ed9b9eec41f3ec3b4af180835dfda637da057f023a43a1689304dc39be0f7f4
zd91128f92133245b23e709d90ab18a4a26fa3937e11b1c4b6e32e7ba7e6b4fef813b8e9f6bd227
zb8c1ffe391f2db0c082f9469eefaee9a378c3268576415ca27b7053acf392ad43e35419ec6ace4
zca76f5122777507eeade0d900a602be3badd8163beaddc2d6d9b8e8013fa1b08fab16acc14b004
z3fa1119b8c499fec42e3e4d97102fd8459124722896cd4be4ab1fa1b759f6bddcef60cc90cb062
z9cfc73fd40b2d19bbe52c6a02e3e34856bf55b3755772f878ac87ee7dcf50d5dab1d21848c5b97
z6bf2c7ff32d38e755253c5d76c1b73c074ac2f7418b08e446ae43d577bca4e978039b9313370a2
z57dca120d88a74ce4f377a540f2002923e8e3379ecd57f887d821ff5e6cdc712b263aa231c2b30
z697e2d3c654290e9afd5785076e91c79032fee74a6eb20969e066382f712a5554f8b0a94571c6e
z52f2285a83a2f6f9e517abddce6a5c980065f9def3133daad6c2541990026a0daf7c6e8b7541df
zc0821e6d6ebec4c5f14954a9b0eddf4efbfa04388aba2c8b5a656b44dcb7256dadb62dccccedc8
zbfc8fbbeb5a184e435acd14a446207a5f7bf0606dc387c8a6808137819c5564297b5beb2426e56
z0e15b91dcf2faa09ae796ae97eaf5916eae30f9cddd039f2ffe304d30eb8380116847a3c35bb54
zdb24b681153321958f230b313ba87c50415ba18fd27b515be5153ec03555e716383b90a132e12b
z9ee8096b635facaca6f517571850eb5de4b0922bff9469050198bdd27839885164c9c453c9404a
z72ed2d78845e1bc960d85cc9b630fe35a952fb9981cf29c28ac896dc11cefa10afc74066855cbd
zac9763198e0d57f43512c724df49bc5e0746998aa4c3721fc87447ea0116541649689257ef1263
zcfde36c0c025ee75cec4127a2e5699a9cd8528870b186a39a8410f28ef32dc43108996bb7971b9
z7c68d744289cec5e98fb775b583fa73eebc66475024c6c6f7bd4e69352116799b11faa5fcb7676
z73b99405ef1ea31d16d82bd5954f5e81324f003182c9146d17a8562eb9a56739ef1cb3a0e14b5e
z8b353fb545aa2c65d5cbb5a623e192ca686d106a090dfd72d453b43edff012a58de4bc42b0e611
z24c6b30efbc3b11975cffea1d2a055b95d685d2321c2175bfa9e298f1bef7df4136acf8d3770c5
z27d264d7336d075fee1039009516c401f251533bfc7a49366c5be83e6a9fb042a76f1351d576a7
zc1d7cd456db34a0b8bc376c670bf796c4973bbd55afae25222fcfdb12cd9260289c2788bcc667a
z6b1e258e7e4214c42c602b74b37ce14f269c3365ba4c42c6d70449df6cf7cd0fd1b1d1bcf2b297
za60b6234cddbd8633605f71ec94f4dd6f3cb67028b0fba4a8958ab1f367b61f50cc868db7cde4f
za4889954c97708e4d32a81efd6c50cebf7760d66e2358bce1abc5396de17de7836f8b06461406f
z82b0b61b4c92e0b069f9ce3eba200d7978018b258e9b420cfd1b246295bb9751990c10b750378b
zc43940e694e21aeccf80e49e6713490318d3e4e19adae93f624cfb652ea570c3a57abdbeaedcfc
z63b90e2454b6152c7db41d607477aeeb2196be510e1fe231480290720bda7a9219ca66eb5c1ad0
z9e707cd23f340fb5fd3d4c523d1cbb16d961a3b1ec9497ceaf06d6995ae50ecb2fc137e3fde5a3
zbe25c14715e1ae8b3bee5872910118a9e8b582da71de753021408d40252baaaf9adf00f13fd1be
z040fd106a61fa78a226264ce8d16c8e55050c6033ed56625bb0beb9f15d0137099d8fc5bc1160b
z392608622c860659aec00eb4d3017026e4742782a67723a9a6400aab8c06361e6186fef480d5ea
zd04e06b48050e0c95e679ea0cc633a7d3e3bb924e15ce9e7c022456761ecc6aad28c1451cb9137
zfbe38bd5241660dfec4c855dc279aa5e4cf094741e0cbbfc087c5faeae60b13044843847a8f9fd
z7c0f86ef2f65e6a1881000e43e42b3f04dff1b4afd76df015d9fcce3097ba9495eaa815936e82b
ze752760a95a0ba7bfa6d23657f39c8bec72612836930d3fd3548edac859a212647bd6cbdd3d6bc
ze87e9784c0461ac862d4d64f9e44e10384b5a37f1ae6d9925541cf6ddf666fbb689cbec314af4c
z3c04aa8f331e943ce23953f3f9a5f9430de34253337a17b7dd9f4ecfe564ba6249686528dc0a24
zf0ea7e6bcfd305d175fd5e45245fdf034c54e875b3bd6ef9c13bcbc379dadbb944cd2035146ac0
z90ba4a04869987b47056f293ce08f1c7d1f654054b4b08d641831199271eec0014fc93ed9aeadd
zc19c8b79d77eb807d19997f91040ec9d83966072fce88c0d404e6927ce0e3fb937be6502e8a346
z5402d1da2804e52b77892d76ebeba10b24078fdbb9d75ff4b1abbb2dc30f6a91fa8124f48699ba
z4039aaaa026f147e3be2771ebab6af0933172aa317380150bae711229954a6ce74364d6b0f6bf0
ze650dba1d3d47c139404d841a315a92433062bd4ea867916d3325926e8f8873f1255569dc4f4ab
zc32263563b97e92dbf4ba214ac807afdcd3ac85c91d651998f853cb29b44d057b03bbee0f02150
zc21859165edc9e84bb5131292d28d3ddc6c20236fdd95d36ef65cbc6616ecd1563a17893a7f335
z554bcbc4a4fd757983adc4e30ec0e5fc0dc58bf876c3c654d858501cb149bc9da50e627fd25b5d
z010307c8c5bf15b81eae50a88ded245b3d36d9ac9acc49c4c39365b96e5c8c0ad8dccc6c2ecdb4
zcefb1d8e0395a50b6f1621e5b0be7435920caec5708caad9b9007f2729ec625076a2d1f1523ef5
z21902206be2668b0207e56aee52e2734aab343fe98cddbc598d85901587da6109b03a59bd2c16b
z56c26681768c324794cc7f0c41d1f54a49f75016a1d7b882a6a0e2bbaa358e95f58684eb37c918
z98f8f8b60bb7b5028a66216e9015593e0135d4f89fcf44adbb4fae866d1feb6abbcf4d5b51f287
zec72046fe3f1cc7fe8fb84064b95ae5af5179283335895d76d5b9232915d4150affbba028df3df
zc486655a4412ea058617f57b0816f29abe7e2dddbaf2fe7733df44949aaa530d834258137e50c5
z0859ef8cd1e702fee55cafd96dff1924b1956f04caf76d0512d88213ba07b71fbee5863331363d
zb26b6aa5cc006d0dfe4453e7a9c5b8e01fd328851a798d3776f35679e2beac287d7ad33c264e99
z66de4c3477e1a992665c2d8004e63dfc216196dc20304f8bd4c0da10b63d2d41c6c8a09d318418
z9bba67b65e15c88086df6c41f9bb6394bb634a5182e59777e3d175b2122a7b70cb8c4bc577690f
z111681cdb2919d02de3752c2c115aee8d502184ae0f283ef6d60ee9aa5d2db72822587f9870a0a
z8df0d8c3e928e59bd904e404c95aa43b4c9e47c34f15e4010a18ef056f02b353cb18002b844db5
z111d5a12699ac03cade388c5f095d5701e0585ecfae16c0518a0e743a24424146a0bc385c9dd20
z6cbeed5f218f3ad9f5c6a1be6016d30a07866ee34aca42334e3d24f802470747e45ee38adfa08e
z5497e500ff44be955ebc0c64612374dadcc8e9f553bc2f71d40df8df376152c7df7131f0155958
ze7cd9c435e7250716b8b6563f358b6b02d47443d1a2d6b7d8bfc013a28fa15a4c149af3b72e817
z2fff79b05699fdf6eb74a99a34736db8755302d9fa44697ec5ddad2f5d8ef348a566c56283ce5f
zbdc9b2d4ea760ea609255fbc017a72cb3c14226acb884d1dc130204bae7982ca7be3aa1a7bb286
z321ac1f60182290ef621991e6fd54060b96119d69eede8ba90b497342b59beadaba1d8d88fc471
z72fcdd74f63cfb9bea6f9def09829c771e06912b1e431090a24c54efbe0435bcefb4bd84afcd55
zff925ac1c41a12610e7d3f674ac77e65825ebe2d6705610683fce02cd6adeb9b3ed0e441e4cff0
z0a651aaf83f0fbedf9d705a58b77a3f49e22935eba297638e2d7308f0143c5cac90b1367f3b103
zc1caaa1665adf5f281c416d9c1d40617248ff7c343a39e1c2a344e46ec0f8034771764c9b92807
z95cfbb564f86ae847eb1d4b1efe3b940b3738bd7719cfe1d85e8146b65b020e691230bc950980c
z3d148af477b6c11e1a94fb4aae567c6cca4fb343de8d1106cde6e24f36cabc1d424e6aac8b4bd1
z896e6fb5e429fc99ded13e9beca78fc45f295c323ad73c157876cc3fb7416af32753ab2e751be2
z5bce4cc49f3e84bc19deeb25a04c5bc1abb938a1095c78aaa8a95242461a65e1677f7fbbd1304c
zd29f41a6c3df5171a27fbe4bf95b09171ada08a17579eba663b60a174bc327b0445caf51ad0c2c
z36be6f9180e485512ee5deaf92515f5b6a992e04823a5e9db7b2cb97e0ad99f0f1ce794320056b
zc65ef2aa68d67f562258661cf9d49429a945445dbe48c3587846855c94d98ee82119f27e881299
z44c0e7a8ac235c4f0e165646a62d68e6110757e8698f215aec025eb6445328b472c8126be7f5dd
z7408a1cfddd9eb9c68f55205349accad70beafa8a58a1f218e75f93b95f854973fea49b7b580da
z37324143b795ade35c5d3688ec49c891dcd75d249a3e7b09ff94afb7bdad874a3c819fa4e57be0
z84c5784c3ed8c16916195b3749e54ddede2dffc1810002c40af0c1515e42b3f76f730133ea9186
z582a4a69c6d6fd44ff3b465bc8fb07123ed5e1187b0c8641314e163a5c7697c5382e6a64775c5e
zc426d536ae88ffd383117e29776f4c5fbc0812740ac209cc4916c3e28e7905d489e18306f22144
ze983db6937bf0480f82ac3b21bda745464383a88409da47a74656d42dab297204505deafa84393
z94a655e6be88155c0d4648e02514752d23c04dabdfcb2087e590c635f5e8b5d73295df4aa631e4
z5ecb45aae873fd9a948e86523821593aa4adf1da31b4d3c687cc3589bb05918cd63876673420cb
zd0ffaf122b3693f506a107e622f0a651e7654558c8e6669c874af40fa626558172d2b4b576791a
zb2add63b9bdf059ea96d9650f810c537188b58667db6f3bba1987f9aa66002bfb40c421bd21b00
z19d7464b95a4352d67717b562dc8ab47cad9d53c6fabbfa2299f7a152ddf8f174cacd9796eecce
z5bc0fe39347d1ec035ba2322dc160a3e4bc97680a652c066c7bb2aac490f5b1686ecc7ef776d44
z5e108299e10d3cf1f8547c01041dc784699ba740cca839960e26da4bebc36c1746e1c51105a9eb
zc031e513726fa6be1308e94d1eab3ab7bbf5d4bbf4afefddb94936355a565a6858af3cd28db854
zcaa617aee6c7b069170f591be09a951565e1cf2af222cab84ef4805a988a27924862a7fad52179
z5768c64f45c0e2f7a78141d519cf501f8ab29e785db22afa796cbbe22feead4c8efcac501a8cfd
z95ae5ad5f42992ff0c836fb58d9e4d13aec5e0c0581cec678b9e3be57d3534e02c5f89724b0e35
z6eaed45c29fc66900e70a941b3bd0fbd25c04d2c6ae88538cf83e11ec37b94472a2bd9566b7d57
z1fe9677566f790b1e7bf690ccb2b6cca802bee08f6ca0c9de33fc0ac5dd16dfa87c646338b77f6
za5d1a4dfbe9568689d1b66ecba9bdb00d3891a4a3796a9ea298c3cbad468497aaf755769114a04
z8b59526c95f98a57f983a170b3b46deea10a8454ac060fe1918e87d11428adcc00c91d5136912a
zb0f45d51a10cc17df0b2421ac56aec74854ec1715e1b6e7eda0ccb431cef94f83a7cdf45bf81cc
zdb4a5d9f303ac07eea8af55858211751c8cf37f22c6cfd3b665a1ef0ec644e45ce6a7b65a1a99b
zfe38c2d577c122945f6f84c46b321f5100de1de047afb79ec6cee08574662a3f7cadccfa94684b
z2b64c8f6b213368cb25f12a5f867565dc42d5e17d34c1dbe5851fc4518b773971da116a627750a
zdf0b67f1853432489a87d950677321f4baba83c8854df2465498ec2fa9d905aa2d882e50d16d29
z5d0058ea8526dcfbac0a657c138887e2ddcc52b3b678380d6a6aaf1995bae8f13e61b210b7231a
zd855f8474a458f71bad4a74d3e8d61c9271841b1b1385baa3b51711a6705660172ae51794b497f
zc989fd281d9e3fe3c0bf039d1e57effb28640455132436940a9750f60f9bcd5f1d690b1849d087
zcd28ab88cb88e5a33edc41f09182c990a14603265f4181819ba8e7705ba7c5effd2e0c0c8783aa
zdd24639e50076b266128fa98071059407ae9340811b8d12828aaf6eb0bb4a3c9fb19bd0e8f8351
ze7eaafc0e602050a2db09a9c0a0450abe46b08591d02624dab85e36b81e38eaacd4625e3d3de02
zce55d8e82cabdb0a0c159669090e674e3f5101c9ca6190229ed7862bb0f306bb1f05982b19628e
z762f3ceaaf1dbe6ebd70dd425609cc9f7c8c46eedd063b10226997821c72e688f28f94422d9726
z5352211b31021a71e9248c1a126a8fc368ec080473afdaaac7909ea3cb87e05fce688b01a342de
z49ff567b6d1d023b980fec283f35b754da4d56efc7be2434ceba8f172a672b02da10a9a9cb3de5
zdf0914d5e4f44a1f3fd37dea79e3ef1700195bd1629da0ed2aecf43ef3c36d7985878144484219
z69197110d60baf3760e9c59452a222e9d8b303ea2e6ca2d34a5424fd2c76c290336535161b9e80
z887094a48ef163ad5da0f8bac8b1c4cd4f812fa45eae5ac0bd53120c987223ad11dcf8e7e456b5
z2b27bb39fd3841a8edc8920acf7a0ce35f791e7caf12795548bec63b8f2b399a8bdac277638404
z9fbe0f131a85b3bb4b7a221008869aeececb40a093fe0f74844c20310c742c99fc6ae66f9e1e8e
z54dd2144433a69a9d0382bc082e130ccba11cb157487e4ee9d3497207062aad25259097336e212
z4f54a7d7d73b4bb8b6c0b3ebd794d2be0a1d1e14879db87c7a001d52c4d4516b18631cde6dbdb3
zf85af920432e5806e24e29846ef7e8c6a984e29fe7672637e48ee41776ae8378e81dab17f15a54
z787505557c5c9fa36380560c6c738e53629c02cc2923d0ae75b95fa213035ac956eded4d9ffe26
z3fc577ebafedf59260c5a574c53a9aede18c87fd0a663ecc142eb4fb323f6c1ab43ee9cd60a9fc
za6a873994270a04be3ef28bf44de996892423749d1b9f64a571ac2e8ffc05b608cf96516fd91cc
z215860e3d101e544a3802ae708b7e2be259a93b266fbc2674e74577cca1148c36ae501f7210c31
z7806b628c2fefca745a38ebb5c7f6fc75386a46421a430c738395c5072d9a7c13456431d787941
za737ff2d45b0d6f0527147146e06637442eb331983887b8fbb3a8a2a34f517389ce46e455ce5c0
z169e2fc7950714a4ef5016be225552b6cf2635bf5b6a1e9c3de52e5d606a5f95735189c56d135a
z0fb50bd1511341bf021cdf58591e276e67146c6e66e149c5a2bee33de8b3d76620edfeb7949363
z13973b6cbec68e26b492bded7ec64847336f7856eb7ff06174f9dada576901657736fc78c18e3b
z0e09cd806c49e4f7bc6e47eeba5f4374a6d330b36a92b67422f75f9b2b7f79760e310c0cbae52a
zf569a99d52cb16025e65c10160b4c752897f647880cb8d4fe77ef162a1c006201f22d1f0ffcc1f
z5d08f8535e967ddc490f33fe21c77fd79446b0e8b0477ad7c7216f37d38047a598072f0d2175e4
z45f99317704fabad89ea2001bfc0236d0aa7cc3c2c32df672c906b5fd8225b8774eb38586dc81b
z7e6a8781614a7a2db234de10ef28c37313e9255b64d342b15c6cdb951cdeb7668ec09c06543b51
z61d1c6fbabbd9c0bff4ee0755580f01ac6f75ce2b3762ba5824b7c3f73249ffc7c066de1d473e5
z9c242e2d35145e72a9f5aeb96061d0890027f7e1d6333582736849ebdfb1216942e3793240fc5e
zebaf2b228474fb1fa15a9fc6760285adebf178b89e5f701ad8e51dba88b09bac5150862d7dfc33
zd49a521874e04ad79cd779fa98e6e442c4b9f0a6b2e89b42861015e4f9bcb43632f280c38e6b32
z2455e9f50f62093b1a6b23554087967fe21f59e581a0ba80e326500ccd32818f508775f17b7cfa
za17e0896cf18b56896c77d5d8b02fde43413b9f0af983cc6c64dfbef2287bd0298f165a130fd11
z2fd98b0968553afcbc91cd8219d79a0b9bc2c4e9f8b14b864b748f67d99ddcd12920bb0049df53
z7b16854018040f6a309ce1f090dd5c4b9615a169d00a61e8554a40a93001cd8218e378dfa403fc
zea9a682be5a17d2b2f29582d495af5b87c278321e3ffce5a7ee962ea5ec09ec60b8c58de6d123a
z5a5f5f4ff10aeee9baeddedb8293f800923f815d4fa91e8db03e05b764c6baac670b4eb3bc7fe2
z58dbbe0652c85dcc0a89c9742ec4a80f5cbc771c52f9ccef7b01b97f71010c1da51eb560f5de5f
zc9e0694fce87479867b42bb3fb511a40b0912ccf221517fe7e9cce2ccdf6673382b49f48d4a1c8
zfda1ee26dbf733f27f9596fe07f660e9ae404918cdb4c30a26255a43f21c52a5f97d0f89ceafe8
zdbf58145ec17c9d91ea6ef3bb10adec3bedfff14996043302573ef65ba1ecc99c162a130c5abb8
zc56a7d7af603ab04ca53577f4638db9d0b551bf07508ea60b4d1fece5a3dcb76e5ff77f6c986b4
za204ca5386f5ce830cab66ddb9b80ff2cd020898ef36e8df59be8a9027b0bef4c13043bb4ba37d
zfe9246a55cf8afe87a84b81c2f9d66afeb5daca388521bbb2b3732309bf23aace4b3cc16b47e30
z973f2f7fef6f4747a75a5eb5a96170a87e69390c28dc07e2d4c5bdfe99c7a82b1d945102bbc7c9
z994bd7423b1921e4c0ff9af11ebdc67f5f02c6ea2dbb7b020ecd6e157437e35cf5074fcab6ca37
z5a72fd057fe65c3ecb56e0556ded0bb6864b47852aea19eb79c7930b09b62e8e1af2aca769f2ec
zbcc1d71c2c6f7818421a66e31a578811ec0233910ac9e9b951903b4786704d8b99c303648bfa6a
z4b259a3732fd89699e639a4bde3b1b39cb550e39d524883274c95c96445104d0823c397db95c0e
zb2c48520b6cd4c347dfcda9fb3563d2b9512d3c8fe4acd1b31a1934f18aacb32709bb44b75f476
z3de881fcb785ff4633461f6e8fe0a2645c231099eef1fbe2f9eacd93ff7c6bc7ff46cdde3934c0
zbe4c9f7fca57ea486de4d3050f7d26c396360cd3ff1337890562ac53121df747a407f79d01a1df
zfb6ddcf5e2955b28db31ab9f1e49442a9a5485891c677ac0549a5a9a8675627768547400a4fdd0
zdabe58ca161a17e4989b92455ee094ac283876390e396d4a0c19ec7e3f227863572580c1c34ecb
z04bc5a6ac1ac10e519e5b1c339bf50dbdd5d574636b9471618aa98c2e262f93c8d7089f4969a72
z4754bd2911f816ab5066225856159daab81faa3ef6e546655737b269c66879b31704d8882e541c
zc5565c1a9e0d180dcadfce53c15629ba90807d4ac3205635215373e8ad0c89f147148df23d4bdb
z82504b7e0319bcb09caaf6e15f71f3fd99ae5b89960fb7e0a76a1c780502ce11c2d9fadba4c886
zcd1a097997595876283364289df440c988b74562ed8ae973c0a4d8410cfa41f406206da43313ac
zfbbd867a4ae5a935fc97b47eed52b658f8d88deaeceaa5d232b70bedd3499bc9253e8a1ed68f9b
z3ae99c5c9c25bcdc2686daecd2f91c64db191787c4a6cb61c6da240c5804267e125720f9a2eec6
z17cc8a024dbded9fed66a8eda5d32b381d17943853644262f87afe1753ec98b77f52525b5a4b28
z2f03ee90f67a4a9542711e28cc08d7abec036161f4a7b41355f195e89115ca29c6b355645d9f97
z036f136cb648ad3110c0db9f25bae8e25978be81da5e96459c1d5f720ab163783df8e8569878df
zd1284ccb98653fb81fe67a001743f5cf34d6f681cb740330fec4cc68c090e50985e143ea0c250f
z1bc7042115b376da71ece72d29f0d4038237ff2fdf4aa690069ee1d300d702ddf350b01a04b412
zd91dbcd8917108bc93ef0a73d734dd68282f5798023f86d4a5ccf30300b032d2cebd0e379a4db2
zba58318a74009948bcc423cc2af0be1da02a66f06ed10badf48199ee5f37ed873f6ab832e2f5a8
z43fe23e6d29269370e2b0304c59ae4c33f6a488840a910b70b5413991915d0b16df811c0d9f343
z6e6b50722a146bffe60208cd328819e623b63c3203159ba1218151db218708ee105d3cc8480729
zd091b3b1212baa01f9fbba69671df8589552442d948cb1af80b205206acd08b4c872d7d006a0b2
z1b901fd5cb0b40b757f45f569cf3089a4c5807399195810bce3e007b971aa27458cde25600008e
z84e044afd6338b4841a59ae251847c639520e80d567f255fe91a53701ca164ffd58fbcd888093a
z5d8be564b0d1747679894db336cc52f4359a1f56837de2288beef923f89f798af1d3a1ae5e155e
zb27c6aa5dbe4de200f2a2e5d3b6775160aff08a0a7d7c80a25e793287e1d958a2e95d71f670ca1
z58e21f47e6042a1d48b44d98fd0f39d54ab19e4d9065d509731fdef2a29870fe88c7027e7da74b
z6a6d9e4aefccdc56fd724f88f627076d19c9bd2609d63b7992edee8035864649fd956b1cbea5c8
zae592f89c3c109576c079cd7fda746d9c336808ebd97ce805a525944f1ad62f57cbc91045ad9a4
z31a46d55da0d9b8ea8992ea1e00beaefa809c196da53d867bb6302157f49f9f90b5d391bcfdcdb
z60d091ed3379c0b4fbbc588d550602889d153f5ca252d3bfd61d09e923a0ece451a113136ae3c1
z82369ca636c8b0f0b161bd796def83b8fabd4719bf637019671fe8cc4b503d1d4312ad7d5cf3b4
z8296c68f924266546bb88fe0607d1d4accd055fd3979c098dc87e6f4d88a52a926a1f21adcf9cc
z4c05926ae1faabb96e0e4ea77829650aa9e52111ab8864a6d52be0c2b39096ba5fa8d111b849bd
z6ce21572bb7e414c27461107b83392af7519c5e21de4e93b319362b931c072826a519e99b6a194
zb45008bede957722d0366aa62aa1e98fca1563a672bc49a90dc358669181c2848e2c27ec13d396
z84a5b2e13bf5526d796d6a0ac2199ab52919c1137459055bf0d338b1bef5dffb70b56e1811c2d3
za8871e6e8331217b9397d4f7243e43091c7127e5f66aae898e16b139b1f892e231d4ccf59b1003
ze3c56f73e533801a7406d8bc57fb59a69d65eee748fe3b00042b191f718447c9a1e28e6f76cda0
z4c929eb0d189faa5ef1ba5092551f9eb1af712a8b34ccdefa32462708253e8318a909299a9cbff
z6083e55a5cd0c5ace8b80965123b59d4c35c76ee9f7362adb6cc1466514cc3b6dd7e8d0ad6136f
z3d153a3cb96a1b0a061599d7f3233de4860b52f55b4009d91bda63979b82e19d59cd146fcc9add
z0bd75db15dad827fee7245336bb545545a19276385393855b7092ae5af01249526c234d0c7128f
z80d672f03568aa9be48edb87e16299cc12f5e9231077892a7b0d6e92176ad3dd62bc2c99c5065b
z5494562dd4e5ce97285759db4734d3147482e3e81754f8b4835727d4318961428d0186e592c1a1
z8f24dfc598589b4853d7ddc7d982e6e544d29718c0d8e4b1d4fede143b57ad52de9a6c30b12973
z7af0c65305d9438b74694e3420d71f4a2f3e83ac931b069d4883a817d94b8086dba1640b11bb09
z4f2e904ce7e8755fdda654f6af433d3e29c259085ec13072965610e7e4c52553da32ddac6d70c5
ze636633babe8a6a41760eafa2c6e86d88d954d09ff910a2e1021c81311e67e710ac77ffc1ff1c2
z99307333878d83498c0b21661c5df20b804eefa5b356f6e55d5910056e24f2cc028986d4e1d74d
z06e21f5a593791611a607bb89335a04981f31f2ba39895c3a9f08e6cab682642b6d9a9e1249356
z7ec110a7942417f137d0ad3c07ebdf491a0f5b17bf30e8de0889af1a1dfe9b8a0fdf9a234d2712
zcd442a0e6a68b86f67e0808ea85bd0d6cc21c6bfac1346e15b5bb21c24322edcc540ffbf7adf19
zc85f46fa495ca34cf2551fe22e10c9efb0d1484dc5277e4e306f4927f9edcf58b4aad87c770375
z979222a451974971feb9640ed8e2889ce40fb0eba0e7e232f7ae1b8ffdba0fa2039f48e2b2bd09
za6e2a11b7099698c7c68617afe3dd08be948ff2cd93234bf7380e35e6192c7d81d2733937abbff
za0f4a1a9ef8a75ba4246df1fe56002c77e19e01fbf95c2053929121064eb00ab1c92961e4246a4
z6c8597be1a7a3a2a3eb4400f5e5bf2b1fa7c2e2becf751fe53a01837b4a5ba189d7ff53bb04a5a
z0614f77298f85a81b0c73045b2920077461955c03398b8fcd624f72efb7c449aef8c75be300fe4
z7a25457a1c4cc3279cbd717083619ad9beace7cc8d2a22be70a1ca4575abfa17b0a1e666a83483
z6fe9a1d5ba40070a8a68a0df548e02d76c49186878a09713895a72c4d5b1ddd4fdefd464d2470e
z85731d029525ee0e34b9be1d0494194d384cdf8fc0af0a3bfa43e85931fb2888a5f78727ce71e8
zddc0d7337e5750c55bd0eba9e688212205b2bc5b43bc3b75d8d30ef2434f611fca3f1c8e1d7097
ze9a9b0697bdbf3aa306e66b138aa4e31558b358b00828abb1c9eeacfa72a60e011387632415f1e
z8b0a7bf92d701b0c6db38ad2211e92483a65ce8aa755c779819a3eee8de891fc6fb3614129cede
z85f3427170c51f90b60cf2be43ed26aff1e53a616cd35f2e8872dc4af2509d80316e012da56722
z14539f386cfb7ae15b5dddc8ca699f438a87e1c08b806522ea431e5eebad151ab6ad8733911104
zc71732063666693ff06d9a8b9eecb374ef35e2513f5de47b6b673cee7a34eed890ac55a8fa1168
zd2ff7674f83a20e53aebcca8833d4a56d97a023c3c3ede5372c90500ae255223dac69a5d1b9081
zdebacf3c2c6a5ecf77a5e7bbe2a193bd94894f14962ac6ce00928a95c98e2357b50a43aca701ef
z767945fb9c60e0051b8264f6d806d52294786a60b042a4dacefce7dd83656dc83d2edc33f20e5b
z3506037d99bc4e783f72b61c0a3b4efdac6ca1ef2f6dea3365b9ae008aa8d13c34dc5476bd5abf
z7a46b62668856a5216f367b3519096e7683614c8a3d6287cf54bc74564a6fb8d34b4b260e364bb
zb9c8bea6071aecba445df046202b32c27efc296caf0286be65133721d9ce271862e484f2d3e674
z36bf27902084fd53ef07a4c452d73113d6e7644ae2fe68a0444879619a4175c92d3539ac7d3f23
z4c41b25fa2fbd9ae4135b42743b911defc63dc0a4dfefccb8175fae6c626cbccab9a0a2fa00590
z92ac69ef3c35ef47dbefe785175aa10e0b17a64fa6a7193cfe9737c95d7c246321a1310e51334f
ze6c030ecc6ed97fc0332d2a4f066f0c238bdb5b2364bd670252259294c61d00d5465fcf6e2665e
z18517a19a8a68b333c8fc21dc824868838544d40ed7ab1eb48a187d2fec1df3062e7861a1a3a19
z70d8baccab0aa0144281b04a3b653f771c1bcf005fa0c3108599f4e56061b6653fdc5fb35a4060
z39cde6d333b0cd43a6393d7d8177c60f61905fb8fef827657debffa89da1198be26acdd6016fba
z9386a1c5e58615428cccd10b05e8f4050313c19a46806cc6be7db576b81b47ab2379bfda6e3db9
zeef408da89febf81901e93cc5ccad3cc9bc1a4e0670511dc725317b7ac24a332ec467f542d1712
z1e5763532d4f3191fed9032e18bdfbc4ea6f59a23b3544711581958213fc22ed818207253752a1
za1ffd3a20ad73a94d971f09c893b05bdae9b67ec5bd655ab91c0a8c6d77ff43cc630caaa033b49
z3c3ee21116726a62c085ae77baa0fb521d75aa243a6dd5943f08b48aa895b656822bedecdb65ec
z2331a9fd1ef2442cf8221d2e01d7f5dda580b96273b2f9ec9864104c91108a770bbc4c4115a5e4
zc98e06fa79b7ce4448d769019a0b54867af361835e9b38c5c4a4f63d117fbec1c359a892e0921a
z830e8bfb5ecf0c7dd93600940721aac47d64d4e7e1e4004716f7a3b99edae41c0bd9254ae2febc
z1dad8311deeaaeffbc1613d7ee21d9a249a275b605723ae3142609aabba1a2b04b697d824e519e
zb8e5d16af6d259379ce876916efd536498b0ffa167a4a3c4c79e119ec0fe639907acd5b9c82fbd
z4875c7b40a97a02e1eab6ec76c883673e9106173bf88a861f41ca444036b8a46319d9b4334734c
z01718093e070db1c9c7638b9300fa57a6acd3f6edb62db6d23dea0f51c11ea24088a2f07ca6ed5
z75dde5930f8488ac306808398c886ca927e00379af4173f644d8da5cf9345eb8d2cd3846876804
z5e73a908624b6beb1126148d728a49b34344f3b8f7c69687fb8acd32352a875f028117aa9a825e
z124580ede76067c168390f3df2eecb1e4a6d108478f7bce67e7140a537e21616e448a68ed44e61
z2b3e12906f5f881f788431deffd611dd5edf1d155c835844d7e00564df23346db38d7b67badee8
z99bd0a9a6a2155b64c56014f84aa072811ffde4af5bc4048b8bab94e8719dc811288ab369a146f
z649b59acc5ddfee453129e2c78c8c87bd37df0fa262d312590d97ebabb560f2bc9e90e444d1c18
z518dc2034b284256613b16afdb248096712f4fc3dc5e0afe9ceaf069e27912b351a286f5cb7f76
z0027618c8d87956b19785842e64d2ac7398f1f5681e826a399abf1ff709c0e5c678bddc4fec82a
zb0126cff34d7a76355f8bf4e2e7967414e716bdfe45cfa78f6ac1ede65a7b072bf1c60086e29a1
z543212429754a5e8bbceb7c22a08c102cfe4a1a4602f7910cdd1bb453024703fbad2291f14478e
zc2139b22ca68d7e1a764399cb9916428f9315fae5ecdc93b92f30e35a0ee75ea0542c1ca70f9e6
zd2330f6797c43e7f150f4678917c0045b034ddf933ebdb6c73b0bfbed6d54ae7c1a0d0a18ec3f4
z50effc1af6f8d5bc67349290a300a820bc9e92e0d4b15234c3047f795a559eef5ad0797f565c52
zebe9d35d01697705653a3ef5869839c9d36783dbad4f81e39c21c12800b9aebc9240d3c0cff12d
z8ab991d5fb02e8a3610d7771093ce62379c9d2456f34aff1805a25fdb6e095734fda8204c5975b
z314f8c3f02c304de1c143089064acb565599528f8c07432a5b8317aff49aefa3059e4a30b694ce
z29cf589a3ef61b00d0208f1c01e38facf9ac6ef44140d6c7756611bb3d73becd93fc72a8b31a88
z142f48887a276311927029b768cbdfa2c3b7707c093c2f698cc12935be692ee1c593b77d2e2fb5
zdec1f0756b8f87c67bbe529bee3d77664847e470dd68426deb71bd25858e9630f73ac2cdbb13ef
zd9dc9cee37c81a35a73f07559ac341c2921951a3f5f3424816a621f2725030d028017f08196087
z7dcf60618e1ece418d1cf9b6d63b8733b95bb048e8c58406d73f84d64915dbf04c17d0d5cdfeb3
z52b29d9874edadd3af605ac3dbe1a08fe030375fd9cd251f28c7fcac1f8b4149af6eb8c0d05a89
z44912a14018097b57bd61180c866f321b5bda02d95af39c8197f174e3f166f754b35170958569e
ze2cf2380bf70e970ae7baa19954a96b11512d8fbc9e67017e84f116f65425fdb36cc1a96bf2748
z462cc7a43eca0f2e93045d576b9a79c9350286edd809372b0ac6701484968ba1da7096fb37ccbb
z29a72824c46b2d2c2fd6f4b6995b3aff551672783d6eb3c3f755f521f2d98131b15299c8ce81bf
z160f72f42353e8f1378a48d9407a3ce97462cc2e199cd74bba2ba6c8d910701b1e1628a895df6e
ze242ac2e46c4819638544245dc9e07b52643b3b30197c67aa5660a7d04c7da5f22d53edd06e950
z288a8ca68e5e72c31c6083ecdc82a3d7097ca39ebe2149acce9a6f15eed4f77ebe96c5f3da337b
z72e28ed5de12075e6acb7ca9ea888426b79a0028a9705f8b070655b85247bf47d7a4e36d7cb8b7
z9a12f051b3b796355fb61c05481439a1671cb1a743c3b36df79bd8f1c6c2fb32772abd5bf68150
zc8e868458f99fb41b2f6a019d81bc8d14814307523c406990f1671410257bba3606ff770956017
z056f7dcbd96aa0cbfb3ae628e498cd8a8c293336101ba7e36d6102577834b4c0d28e43c664aca5
z9f434496d916dbc3334377907cbf610ac3d54c54a26d302ed8e953e72a085e6d34ddd56c03338a
z362d5d050824b530a7839c95e886b9bcbc456fa73394588dacd044e741362cfccf3c0e3e4ff182
zd4f6e0c4e5087354b0f74560951aa95c01567b18e87296b6bbb25d5fff5d1315f61e332ddf15ff
zda880897f43230b4da9431966f0bb0b67056a13a7f67ae8c255a9f1dc8bab5ea3ff020924b22f3
z00157f4f6d7df0ff376456edc1b8472cb410a90255f8b8b5f353005af1e23c1b4895faa0fe965d
z3be56034e3d9581f4abaeed2faec5dc53d5ebc150c1d47b3c530a843a47576ad0fa1fde5f4f246
z209abd38dbbe621b1c7297b0678156e57045d49e3bf3950d1c5c862ae440cf60be79c5de8f361c
zdfec0a15cce520b7d82df79bca096dfc1ca550109850aea8c0ba17ef9170a2d5a9c0e6024ca9fc
zf9a129753fb13cc4bb7ca3338cc153c419ee19ce9c8e6aff35bd0a1edf34737e873352d5edcc39
z815da168b53ad49de7331831f562aa13b38b6e2ee156d82a04b97b9cc24f579904acd160551d06
zd64350ec9b8c47fe722c12ce0b82f5389d535917febac249364efac2ebc44f58232bc507c6c5b4
z4b1084fd61d8acc3fcfc42ed39dd941c03d6e9f9d8cfe2b1a31a349770b7293c0afefc9f8c96b0
zeab7a399d52ad45c2a0a55cd22306dcccff33e43caf7925656720407023bf2625aef949e987b38
z2001ff6dd3bf9d7af0a7023d6e6b69d2d887561316c282c02cbdad5bc0f7b7a79cd19ce1aedb67
za559b0399d64e1257d78bedad5a1bdc36f9b3bc734cce8d23689c37ed6c8a96025cdf1f39e8179
zf2539171b9a3093cef1e808bb2a6e75ec706391ce471deb88a650fd6ba75cd545e003b284e3ab9
z026a1de25157dcc3babf48322d7f1cd3575c41386ed42d1147f560980c85caf6f3459f216c2766
z247882e5a30fc48f3e244c997ea5c6e963f2e02be84f5baa66c9372be68b8d54280d023e6bf120
z54297bee20d3546de933b0ead869a9cd349a07e66a181b03c46ddc76b81c54af39f578e0125c77
z1f52d856e14f4c3f657857d96b32efc11bd6e24f4e66b85a6169b28fff36f113e2efef02b87c49
ze10e20a4d8cf44cf889522eb5dae0c5f11febf06869d2ab4d046b79446b471e2fff459f0705602
z5644bf42cf6e17babf8f9e24b7486a5fa31e32c45c52353340d09c37b3ebd713d60578c7912f08
z7667bee68529b53c3d6da5421f7b6db5db650448edb16e7209a62a0411b7cf87327d1fd995226a
z8cdcd33fa2e5864ab43162e377a49ba8912647677f1eed90f365fc075fe2ac961d0d5ba1f55ec6
z62a6d4d3ce3a040aae345dbfb29464fc1463867b2d910eb06c00cee92615e74cb82d98e629fd91
z7513c3343472c008a9dafa12719bb1fcb027323d03292399eb6664788331438cc3714252a41ed8
ze5035f269c4f4972039e197dc9794e9975699deca5cfba28465c2f985bee2d5780df5209ad1e0a
z8ac2579da197c44d842c6c959a620d26529a82f656a05fdc9c599999637428a4b53ec5bf6a159f
z667c67be2fafe1763f4d20ab2fc126373f38a23d16f68a7911e9230d025a211f0f2f716ad70a22
z48477cfce0f2cd8bf9db85dec680ba52be08c4d11e7263bf464193869b3c591d758dd2cda39496
z626852956a1a38d6483fe62717be93e981fb1f5ce347620a5fdf8153933cfa951e93d1dab3bc22
zde5f1d471b9de931ca904bb292287fba7c163c945148dacd22fb5844360aedf69852a80d0b8a64
zf6e70eee64f08f5ce1753d901a86584f9e1658a1fdf0bf48d8d76abc48942a90859e55d4ec74ea
z69ff963cc935b685b214c3bd887d3c29f7b8b3335a611f3596b534ff0d77870af408acf7612213
z7187d5716d3e8d8ee35319eb8ede54d6434991e1d02811857b4f37ded52a1b034e71497a74c465
z809277dedd5661fc46ccc9e04805245590593581a4f32cbfd7d9161e055a8641cce3b242a8cbc4
z8b9798ae72184894348eb21f51cbd1f809d7bce5a48d0eea8ce8df53a96797bf1363d5dd377cc2
z4b6ab9de5ac7186c9e8824fcd125a8da1eb66abb994ec8fc7911e9ec80978a80c69947f8d380cc
z53d5fcffe0ef7ef39ea20a95016f4d21a69228889aadb7aff57ee0f056f9d48009689202c68584
z54757876820b63d037d2752bd01dec2ce09bb484b1a6aec1a7c3057cbdffb22ad803a9c246f9ad
z15b5b7fd26654e9987b2309b769bda953383a63e7fc89ce8b156341e7e322f2a5b10f270e70595
z2d1bcd9f2338f83e19de48003134d7a7cf706714ae1065bb507d6a339d3cd5484b08f6972fafa6
z2c0ba9089dc9806ecac826ac69aa69668f3d97be265db94bb540479c7aef9feaa6b022d6abeb2b
z7657c8dcb0f4bad24645c07d8b7e8f44498dae465a373dd377e6ce15461f22a4270c4e1eab170e
z0381fd572f50aac065999a8375e4d5d20e959d86c09042cf0ce5cea422d56057480541027e77de
z43a625e5332fa45674efe58bb9ca384e8ccb97aa7027341f26c91eb31925c28bb9659dc93adea3
z14d3fb76be431d41a01c411813b45b18c707ba1db26b25d20868c4ce4b0cb4c28e0b425123a7c7
z5001fdb73749cadb047c70d6cb8bb80b82bbd3a473e589f6a63ca4fafe06cb2a97e8a7e7cebd0d
z7f001c808979641b6825f6a17dcef71901f7a5aaa566d201999a78a654b16fd751856bd1f0ba3e
zdf35db5783a979cc3809883075f45828f4baddcb8eeba5e796163e3ca7d5b76caec6d587f5ced6
z52b5e8ca8aa2063e83b70564331dfe8ebc92fb770a193f82da9b92a9855601e51133130de73c1b
zfdde18347b67410fe132d3ac5f0ee73e386f95c9b88649ac200fb9c0435dfb3a434134118b9413
zaa7a8fac4cc39637bb0836b541503bdc4c59bc3812eeb2d37ac98968ef0d5563035f0af78f2c41
ze39c23f35bf5c28ab4db2d6e1ef05a1b67d50cea71808cf73a8adbca41434fdd5958798489bb28
z5512bef0d1968d06a79a7f65059e6be4da3fe9bacb83a8db12c0cf19973b5dba7bcfe780e7f8cf
z25b60a3c2710f07ba5b46dc84d1e23427739a4d043489564b4c328ff1fe9b45feb8a1b91b0fb95
z98281a3b2f0f0125d361485b405dc67d54e2343bd8e231dd3d11e979c025c9859e75d04991e851
z4deaef34e8837dc61a738d2eaccddad04a488df67f31f6b6e30fa9abc93728fbf2c8e97a3c0b63
z8b96b80d75692195e497a02b29152bb33ebf857c5a548e7fcf2430917fdf2dbabc290d2ef95aaf
z771bb70709efe8dce8ae13e4eaec832eeb734cc70165d58bfe3f3493654af8d9c885a996b9aed1
z2f3a3291e7d4812368008d461d42f3c5e4cfa16819c044451cde55ee653ef5ec8a429a5b60b9db
z0b39fe7c60823d567808e852d1ec886970def65b69c4749e5385d819c70bad821a44db61151145
zf25abb99aebba50878a045a74222f5e44934f498b3673864e5302c2f9c0c8451c5436fdb8393fb
z082a0f38d71fd1385f187f8065fdb3247a6e070a19572856947468a89d8099b19d95b523f3df66
ze936857129938991f5106ffd6680492d846e62d2d2416042d341fba0c25ec9c40bfc6a705b0ae6
zf38b5aa6d4318db18ac6b9983f7ed60a4c333f290c7c6d000594464b814d64f9a97ba46b3d1228
z4a7727d02012b12e567c2e21dc6e7612166abc9b295e5d273b1f6096e876394746e18cab13c50c
zd584c48e9eeb0b328c93c75022321b3f589b371911a96e499b139994f444b7d6878ea73ab8a158
za676718fec3e13f187263fcbfb38d0ed4f8b7b2428257f57d7b62396ec697511b1b2730b468a3f
z4eddb0a7aed50bc7d928a427b2da99fa960921c39628c8f6edc2c02c40f57c4f061e90b09df7fa
z35e496ca255ccffe10d8123ef43979b60744048f92094f71b3f9f8cb7e4a9b2850062968005c00
zfe04a8cc8191c1d0f05e7e3d31e85a38df9a3f341cc50528ea43ed28628c0847cff4df73ea5563
z03fba0db9492a94cf29161d04aab30788c1f500ccdfaf635ffe5e2190ec395d9f1f1e62bf7d60c
z3423f4cd5039e508ede50710516ec026b8b7e44cf5bc1810ca9b21d6cd6be9af19402e407547ec
z31de37f4bc1370020e13ad8c26095a8ddc9cd366966e396f16ab42b22231ee0f4c2dd37e4aa48f
z334feaf755ea455ac6bf7ee1296425b9135f94fc0a82937697d9fee9b1ea268a3c5fcadbcc39ad
z3cc971d679a4b61c41070c6713b5e5583213c294011e1928c807c3f12f3f144229f51c22204e30
z9f9dbad998e68fb7075c575cf30542f0b5c77ab0f71ac1f520465de5262c15c782281aeccd8ef1
z15d2ac041a6969d6dd9ed32d2742892cde9dfcf2a3829a6265520ce571240cb39f37d0c33a000a
z2dd602c82136f6644e9b9d0994f684dd4d31a34c6ac58ef84f41e5b1904ff6a2147722c196468e
zcccaed843283ed527305eeed6a1b4908a7beee08049c0bb5c2db2f2fc7ea2e3c36ecad54d9fa40
zbc13d98c37553bb669173702afd5034a3662eb7a566a8c283b9fce95ab740b1bc2452af8ca8da0
z74a57b5bd845c807793068d527e1d55b476bb345a8297c592330823627edc3c156c851ad048b5f
zb53e6eea0fe802f71cbd720fa072b2ab3f6c0555776c025d268c9d50e988c5a2b579ca30b94e0a
z3466b8464fe687448e5c8f8a1fd85bdc1343ace348f440620cefecead8aa7e37693762f1e996ba
zba1fa174cff2a3416a5549c6aa921a675df3583b2a9d457e307d8de9666164a2864da1aa03fac0
zca0bdbc4302d6ca65d40d1c95479cf617c6074f35485ace1a818b1ac394cd75dadb0b3855cc47a
zf6051c7ced95f39904018b4a9b7fdd7500cbba9bf313af7aa1fcd68984032aa9eb2ccac087332f
z7c91cb02cdcc05f70a3795dd87e6408963fa2f2c97b89f01dfabf96b87350da7acc498d1ef6000
z2905fa2d4289f28701a42e640319cc5a19e87c07bb924e26b1db105e48b6414de45a580e63280a
zadc8ab6259946c7a15d445b2c8dce90831a12acc5b80151c31fb0d13cd8eca85eda4eb01c13a18
z6fd4ef7d4655014f5b7fc0b63dacaf9c2e3f0955c5aed033282ff248d16b27c56944f0e683a161
z73784883c7b9c3a591f24b6470aa5117c86403ff1c4e798aeaa819bf20c84c0128215753a40ad8
z5570c1c50acbcc2c968111f50d449c2dabb08ba8b8afb8c09c0674b9a8169f9a1a644f89d27e01
zf07194adb1cbab411b4ba51d95e1f7b3811fdfb7b8f817a7f2af0f12999ca2d4057eeb74a15ec0
z1d08be16657406a9ecd03e2d396296a75e78041490499940c7728709cf7e11b283756cf9d27fe2
z627d0d03c4c58ee93eadcc0c5a5e3b2c41c3fee16c1523202f00a93bc7d911ae4a55a386d5d78b
z3567c682692b332aeb410fafb1535273bbfaca6397236c864428a29e0a4a672ff3f35cde3fdb12
z3dd79282a5b40047210abc6ec7ba741c92887a28f95667ba4242cf1254b4702c7b3a6e5abf65ee
zf79c035413815445ae19ce3bb64d5d8989b99a8da7cbb2c2318ff7a3528b9ba42b407dbe3a0159
zf0bd5d86d79aea8b2bf0183a3f9014394617a238f965bab7d3e0cd46f9fe14d93e2f28b8b87104
z5635d62185d977041c820b07fe760e5fb32d2fd707edb00f18342b07707719b64719b4be90596a
zbf2400e477908cae9bb42ab58c2cc5186ddc82e53206815807558c7db4d5a6f8414248b1da8ae3
z7316c966dfd74b1a4117d4e066dc4e8e1fcc98caf4187a2d8238ca8918f0ef665470d92cc3c864
z6000b1e37d3b1c73ed45240efd5cd16c9cd5a25db9c48b8de99554de4f25a05b81e05a6c665ba3
z829553b71afb90151d43c6da996bba55d443fe8c3eb67a1e1ffbd5a48ef2a758f65c3ba70fb556
z832a86b4de0b390cc4b5ee5511c4aa0238f76c7d8521cd6f0157f0f947cb0a4403ba7a5080bb08
z985f13b8adfa1c410a65946fb2d21f46f67a4232ca059970e010a2858eb34c5e55cae7131d7dc6
z25b0d3b06afe733fb4376e09f821339c4574647ec8b4254b97ebcfe7165e38933a1e768fb1dc65
zbfa96397f8c7d558591b9666f80bc0ccadf1c8a1e8f00e89ff5538e3491576cfebbeeac93eaa35
zb224ac1574e32f284e3ef9965e6dec39b814fa5d2d09235bd6b239ab8392e16c35e0abe1c5c972
z00a37677df4829febde2e7c029d30e82e1e88b39c342eb28f56ce69785da4bfaf3de52fd43c463
z714b1751a98250ade20a673fc84c0c8bea822626200e089c95ec1350ab12e477e14a25d02bbc41
zfe8dd568283590c0e10cf04487d98f8abfa3219e21e776f924efdfb1e1c683032966307cb849b2
zef25db0264a8a7f650801b76b64b4bbf77dfb6af3ef827db0487ff41b98e632afdfe073995fd70
z667afdfe0c15d8b2e37be1055044f76f86b6debc4791d95617c4c080c12bf9efba4b9ef3237470
zf2e0f20770071451a3179f3fa0a99a871426b469ba4997e9f3bd55a6b9b4c5f64f6270b268cf70
zcf2a27cb5f0e8a72d11895541914eb0716213cf908beb06be1a5c0274a01609747e5b7fdfd0837
z4d0e400bb88c549fee938ef14be4048b51af668b867bf0fb272be5b734a800db65ddc050a790e9
z5a2119e6bc5b455826fd8f633e28e85c238427c98a63c1b25666fca95742e0ffa96d04f4eb84d0
z1125b6f5d357f12a63cfc51a93dfae8635a6470dd0d8b678740b390dc0ad2725908a7fb5cb0bba
z5ed529325d26967d5c5198da536d571ef85705dce96a8309202e1370e48b7e189c29328c972306
zd42edfabb62eb244cd02edea9435c5865e29ee767f8da8678047f84b6e1ae3843308dd30666d2f
z0b577c4c5ea774c98b82a9b0fb4827ca83e5f2d95cba4d5af7d35dde9de9733a3219829eaef58e
z3eda0bdbef0170215023c187ed28d906fa1df31a98216adc853cb1f363dfc6ac3b7e43f66d9499
z2ffe2882b69794d1a78ea2a645add9bd6c28387e2cdba80f1f90ce3913807dc3fc98f76e606c22
z2df21bdacc31fcee2d494ac46846b4b2886b28af9bb1f0ee2bb96be60b8a73f34fc02dc27bef69
z4263c8482547eeca10d39b11bbf77bae14c5a1b0d9c43a41737cbe033da788c0d03d58b815c43a
z7b60e17317ebeaeeb36940738b74d4b98eaca6d2f7ef3cd25671c3841b2ed936a256dd83144ef5
z9389f56c5abd182b55550eb23219d65d1aee1b46cff4f00f663d833f1460eb44dbc1dbe6a5fb68
z50e5f278f58d954a273d2f5922935fa99d514ef3af78d5caf66ad254abfc062b8a291490300b35
zbbfd5f98fc9e4fc3a4ddf2980fc73bddf075df1d521e525e009bc5a600c2fc46625dd035f66f22
z1388c0bd5a555502c1b18d959e4595c1db88f6cfeb5301c831dc40d28b4465a7bbd64e5755c4d3
z50d776083525453e51cd0be6b919f27a696fd33f07a03f51fad4737b64b16cdfd890d4f37f0401
zbc2c037ec8099a00a1c7bb56aa4014d7a3bd820692a67aa2b996442510b4a1f2fc3576f103ae80
z799f841755c95ef403174d1b4b2c927425caf6f96bf9ebe460a6880a18d83776b64f8e5f6ed317
z1f56fe8d0bfab8f8c13fc2295e642de7a9ddd0b6d29d053f9abe75f80efd48c2b9be691a14a258
z4e874ed6baa7d137dc5084f35dfbec98e54f29a3ca552ae86e197924dae22bf5dc332b4f336b54
zaef5e03de77749bb1fed6a302efa0537524b8c5ce5b4d0ad165646be41f4635562445191f34c49
z88025423b2481c6a481a0b166ae8ded67e0c89f1fda1d8a59c7d84bdebde426fdd2173346d26bd
z4bb4bd574246327d9662568bc70b06026e8dad0eeccd3fca7d6cad687bd2ac896bb904ea0fab2b
z4f0653cde08d0759e505e40b434a3faef7b4f4357e97f90773d8026a08926a6a687f2516924220
z527afb08f2d582bca28cbcafb1d83bb30c0544149dafaa2cc56fa76309fa316bf6be3eae778cb3
z096d6eb5ff239fb2809d7edb6aefa4eff05e3d4eaf532385a6e9de82c8f942d51843f42e999277
z835d8b0bc2fe940558287e213f784ae10ee2dfd601fd393284ff3c6765c25f76d7789308f7bc24
z1d6295016edfe9ac09102d5b32400eb035064de543c7ac208827ece8f13bd1704acd74d2cde7d0
ze942e531ff3b68489eb9d677c2768505701fe6f2ed419fcecf089df9a5e019f873fde6490a209d
zd2886b7876dbffd086accb8340269520c0e6263b7e6dfb629278ee53981a66452d417c3ae4fafe
z28b8576d442479022c0d73a28bd22e3ed3210cde9a5e778b9908a0dc4760e230ce4e92491da826
zc2fa5b2bc83fbc7146b98baf009aa6e9fbc7d7f11ddceedf4169114e472f3ad041f9a6715e79fa
z558eedb9e73d26096766b84ab0de38fcf1ff5407becfc1e8277c8282874ab3e2e0f507f8188fea
z193d22e6c4555f1eed49321a935df88b571f4aadd8b65fa4ce1cc9ad18ed84be1d37e36fba4b96
zeab2ce81ff9f79fecd140c30af33570cad3df2316327c22287001d1e1f6e8ccbf5bde29a61cf79
zb926f92c0cdd822ad1c48f79ce9fa07daf5a46c8bacaab5e1656d287e5255852b7aa18a0891590
z483e00e33a86013d72138eb4abec98b7608638f2eaaebdb747f99c04cbc32fafe5e928b711aa1c
zea6c800297e0b9e4da5e6ec6cace050597f09e214fbccf547f55dfa7b9f1c6e09255083938b1b0
zdb064fbe43c8a60ef557c5e15de1f7faeee100bd92831d5b7e1197c8a2a41002f522c7292bebe5
z5d2271e42e8ca58c47cc4d9c477d7500d7efee10915f404d743b42ed9b98d96569df5a1ac08bd6
z626b641e543abdc24d14c37464cbb71eab05142ada3e64f514e228498ce66a0bfabff183bd2447
z25157ec980fa57232634d78d0d42677a2e692a9d95b0d782de4d244e9fef7deab043424cdda944
ze45ee0183f8d2b3f9e17891e3c8912b8fa7fee9e7690adc4c1e3fddef40f63151afee3bb069b7b
z08e50ddb02f35611dd205a9b1a3346926b074262a7f885f6e6c627c0291caec4b9795ee4b719bb
z32a4d2a09b2b98f58d04d16639a0f43d5e7688dec1028afa3cd89b9a3f8837bb0da27d911317fe
z242c737aadfcf9ce8206bef3c6fbc1ec7d4bfc385da17a3c9ac050c21b49646565b06121c380be
ze6b4a1fe7d36d3921cf7e018e270de5c022edae2d91e2ad7cc8870a733305aad64640e507b6999
zb5b68bb80d38ef21ebae6d9c0e8469819d57e03bd629eceec6070e062ede239d3d025025b15c96
z1a5498b4ccca8ee59aa90535b19b372de7345b0a1e49bd5c9d1bb16f3bd71bd20ce48eca740a7a
z0ee99bec2957ac196275b738347208f411428203206e2fd5cfe74babd6d5c9cc0ca30c1da37072
z30541cba1d058c0982484578ff4b9fad96f47a51e30573d5cf7f328761dbb91664020cea7398be
zb069e2be7e72e079b13512fe37dc8f6b887787a2b815145dce05cc3f29c81d875fb4f10a3005ac
za7c0e55a78c44565e0df3b31471b4bbf47bfe7d6f2c913e0d5c4a8abefc261d5eb55662c068cf0
z4b102fd92b313a10845903bc3b3b5dbe0027645fb03d6e12a7170dc953083fe15fd00da5906612
ze714d4eac4ddd4725938ab49fa24c7b188f2b2f87eb8a0f8b34aedc2a14189aaa6e62e2234be3b
zb47e3716b1da49497056598d96d28d6245a979497343e6567c10cbf0cc566c3d1979ff32596d3b
z716e46df449a76340d508d4e38c4e9ccef5619c795ed7347511f8985308fd6fce859394d27e6a3
zd86f2f58bdc4c494126b1ba4f88118fb033cb719374e7a309b7e74a33f3512405293b91a42c562
zd6ee7e3362299f270cb6bf0c290ed19e05814415cee5b5bb0187d350fe2bc955ee3b78e738468d
zf399f1f879cc0f4318d43adb69f1f6d5f1559cc6b6c1f127e96ba7e06addc5be6823614f589c55
z326ed65b4ef3705f524641f3d1b406348ceec9b3e4640e0c1f93d1fcd4b9417c601ca59b83dddf
z4c3ad9b31f72d5b733f25c729344a920011c1f221a1cc538070ec649bb4188e7faf4a951c07176
z5ae76401c27b5e1204b9c5c739a2311279299bdf0f4ceeb8af92936cb834081d58b3d420ca845e
z5ffa10a2c687177cc76a18e3866eaa2130c41f3d66448fcf7d458c6ac5b9e4a58bc4d14f9c7317
z71bb6be98ddbd79a694dc8ce196ba6f03f21d75d6c135208bc06ba27e02a9acc2ed325883000b0
z6c1142ae790a11fcd72482dddf68e5508bec344e196cd5b5dd4a428bdecfd93ec11d0f9386d70b
z34002157bbc1a959530713d3a254cd746f93745ab22024a747b705ecb0ead19020154242c17b48
z10dc46d269aaa16b86f19a465e9019cfaf8a7809d577a1486e1024ca0d5e19e9eca96c5a016bce
z439923f7d760ad7d7e16aa9cd895c8b226912c6836d5467abea7dcb933c08585ad08e6f17cda40
zcfcfe8df9f1e8926d016b9d03e258cd674e60cf06c60b43db5d0e7812707b571a2ba81e2f53dfe
z64d6623df9d430618c2515e3ecaf0349310c1de2c01dacf332ffd092d1dff0818b802480fbcd9e
z057ecd95be92a2f9a6977a1466feb336882eb77e7732fa497e5e38186efc37a77224cba12e1598
zcedd8765823088fcd58d22cbef3877fd3001be00008cfe684e20b95445f036a288fb9acbd028f3
zd7f8c43a5d8f0c2e93248d970324ed1e5a1121a2fe990a5f8504603d7fc1ee36ac9473d3f1ac27
ze41b74912681b12bdef498f285b4734ca1c61597b9c3cd08361c4ca2db37788eb9762912451b4b
z760a890c44d087e52de4abad70db50938ae808d573c40da8f62764c3c0e300931b4f30592834e3
zbf730d508ea3b9c7f031f0e936630022b943c69a359c9f95c23dc6b3c93414c4e323de1ef57604
z02c7ed345aedc5602eec2d03a05266e6fa4bf2fd037600450c5a0adf91f9ed8c927f27d511cefc
z3e7c3a3ca110a0ae8b50bb00400dd74663c9a584e6bc0577980634fbcfae5dd4e66ffa063e6dc2
zdfaf144d08846af8f40c909bfe2ac41a6e51bebd71e25b250b30d570992075107b07652d78a0c1
z75e67d2323bdc2006617734a62a4e3605d452925d0e43a6d03e0e8e141e878faf5ebf0a7ad5231
zf634fcde64658acd81295ad7fb1edc28bae79796d65ca68bb519c33c15abf1fcc2314ed81131d8
z947614454c8b3fba3bf6f1760a7de66ebb18a8f0a93aa01aa212e19dd0c06cb02884b1042f2821
z67f2b2da421bd40807ef3056795839ece39f972314d34dfc4dd05653cb08cf8ccc6eac3b922ab4
zddfe952e4c50895321ec873a049dffb2d7f24ac743eb8dccb24bf7e38e11e063f84015d6f5506e
zf12dcedc76f32139025c230492430606a11e4c245863a631b770abf2d3067708a9910f423c9b1e
z91002c6dcb0296df6c4ee972059dbf0ac726166f41e34660c83052c854425418557b2fca2f9b5f
z336972af59115068cbe21bf49f9afc8f83442bd657cb0946a3bf711299db30764ee042a18a3c0c
z9aef8f65484fd32c6ba85fc1694acba80ed6cc3fe24532366a02001597cc4da226c20229603415
z270b255c64a809eb0932c25159540ca110d18b46c4d2d956ea3b01139bf2fbadf9e7834e6444da
zf4ca4431edbb50316bf2e1d589f996489e0bcf2f74d7716703aeb3863df031021e1842ae57e599
ze76484a35132f1c53d381cebe58643e991b63e3da1b4b0f29738e746f8474f3b9593ba18deeea8
zfc9defc12b62a287844a25ae44bc3007f1b27204d81ed52de53c56152b8eb68cad452531a2bb3c
z47bf26b5e55c4b17b878a3a6e46d1a21d2785163c2ce6e18ba88c11122798f39fa4f017a6b9c2d
z2e1e4e09c4bee6b218befa3d80097bd3e3c79af7e098e481aa9b757a037bc4ae627c21484e2258
zc4ae87cbe4355356dd3c3281f5acc5d2aa81efa946e58e76ae10f00b95169e5cf479a858412b29
zddd8632668176d3fc4ede70a6b7708c3a3bb87bf403003ecc2c099633b3266cc156199404e5542
zd667d7e50753e0c1a3c68001b7acd99e586a95c85578f203f8c683a08a2567069d197861cbcc27
z97a24ef2ee6d72508d2fc3c74cfcd74c5d24d879346551fa717b8e7cee3fc68455d1868268e490
z35179d8b4b163066a9786eb5ddf911dc5e6ff5b88bb2d99204700ce44c9356551d7e3d6ee33005
z45f5e5adc6fa5d5f9fed66d40e87209afcbfb0e99c098b8f2fda11a08861a569661b563fae62c0
z2b81702334675c8232069940ab9e7ea638bed8c7f3ff7c6284c82a64b11810ef1ddf3c5e9a1b1c
ze17781e762fca682c8e261cf1a82834f94b40cd41366e8b7c2efc39d049c423e3e49bd78154b02
z77d594c02de046148301ce875cd917e5703affda04881913869872a55416fbc8e04d70bf3222cd
z43cf5cf2794139a1888a6239f505577f635781f3470ebec3ce1f8a5ebdc286efd329844168f26d
zf907b50b5cf182bc4c84b5ff9699bf7c7d500e5ac5c5b623d7b432c8ae4a9de1a991c5bca942ff
z85bf392881d70067221f57ff0d622f7d094c336ca0068f8ab80bd977e22fa2b3e1367fb3a4d7b4
ze55b93c7700465c394e5f8ed145f49cef005162ecc1e126892f4b34ffd7f81bd303663bb0fbaab
z03c65bc9ea9e04d3a2fc22fff189c8faed78989ce79efb076d3c8c953ffbf0f1caf1779d3d1735
z4a76f9a907aa240185a3c474a20b7da0c25d0e8a507ea2c78484a0a74b255e4608ed2415ac9a95
za5124384b5f1ded8631816bd3269bf1a667bb60ed0a2f7926706c9537ab9d10aba64c40f7b071e
z643b7eeb921609a95e7b4792d6e56a4871019b08f7ad3a992a00e6b0f3399838e16955f6833644
za82e6ac41d0e5b87ebd9cb03f797ed6ecfe6563a8065d24cefd354a06cb32b6725ff88b7bce74e
zf3709923d582aee1414e7f6b5b3fba66bb9b885eabb1ead3867c01aea95777afb8a74ce837e926
z84670ff6e1c370be4b6a7c9b3048a0c762043737ec8f017855bc2a45316a5cc3c3ce83cb4f3ed6
z3e9534cdeba1a7b6f800986048655320ab100e17716c8d53fc02b5946deb7a64a307d3b939428f
z02ff7eb6cbc2324dacbf9dd4baacef0bb6d6eabdba729936bb0cdf83ca0d1563e8935d378bef32
zab7c98ab88cb55e81c573722d6bc02189e2ad26207a843c1f0ab23de06734f8edc2b6b916367d9
zf776ec6081e96e5710f8008800406b36c2037b2e93855b47f60b3e3f68ac5907690c66755a0493
z0474b5af80073a686324635b65e5f4210801a2fcef2df0c69d47418bfaa1deb889f7cb61b373c9
zf9956c2a6b6dc5c40f6398c4106fe3d42e70716290b630896afca9c7e75b64a8d2222ed7854552
z81302d24137328e95f1bc953e8c15c5f57aa8a9f465dd74acdb2b29ea7c3a8d612b5fe875e0315
z0aa8572b14ff1f1d50ea7e2d7bcab6c53b8da6cc501078241361dbdc16c56e1c8c07b77f4bfe87
z76d6e389ecc304deb2c938a3e61e2753484521f16e9d0053d5d77cd8323e4025739fe11e592c6e
z3d65932e71e68887994f4ae20a38e9f688177d2abaf4fdba8d8588b55063b9db8cb0b11e83e0ff
zf8b2e7727364653f05d031095bac58bb8ccb01c7c58cf8221c55473a3fc04021fb78062da3377d
zf4a2685bb3ac1ee0cd902361862f9062117c3f6a624476f3afbbdddb19087c281fd62907ecfd8b
zc5155de5753c772b1ec6efb8002186e10d84bc668bbd9aebf64975ccaa3da61b1b20c21f9b58a5
z7f1f6cb6028b98e37280ccbadc69bb5631081a347b880fd65ad204b60efaa88960e17320062ec7
z65923b741bf0a68052fd8f55ae9a9e211f7224013b6b6136a437cb43800c4e512818c7e62389bb
z92952885f6e9f58941c8f836cabe76c3a21eda0f624e3e49c018790996fd2ac02e02e198f46a38
zed24d0b79e185c699f6700350bea21b402d915222b6bc0495a5decdfe7df44b993aecaac42ad97
za1242522519890325d13c7dd403bf02009feef4f283d1bb629c7256a759301a96f82686dc4c810
z3de24ce33faeeed5756913bdc4b60b4833fd6ae6af37446571103012a5ac2deef9779dfdfd4aef
z634ae31e9e6a6837ab9c34260a4045a7f85902a498a4637ed31cc268b42f037c7b4571392500e4
z289926e2b843eb49f391b0c6a378caa2e2c758261e09d4ddfdb00c33d35505ed8686856f38106c
zc20c69633c82ddbc966a74cf838cf6910869b80e573a2c3194c8e641595b6f0e7daf69a88c9c76
za80ba7ff12430f7b4c57da26e401f185aafe05553bc6b680ded641c1fcb97cbf689c63faa74f76
zbbeb14718df8e4610cc725746d5ad061b49b4e1c52399f5156da6ffc9b28ade0ebe9ef08a239fa
z01d04d9ef7e2e63cf23fc03b2a3a95e430c3b75cabbbbd761cc6f08ba20a74d0b5883f27abe5c6
z30daf408351f2850b5a5df76e29b2a2930dc51f6ef38596849dfa827f68238444237e9b4162c16
zcb3aefc6157fa8954031401a011f4abb7fd3f160c468d2d5a3c8aa26ee771205fb8550d86e6613
ze66607e6f9d15a3906d79eb35549d2d3bfc82df9bbebd4a3d08dcc9797a1865603dcf49fc2c6a1
za41d6c3839991306b46bd512f58015bf8e46ed51685cc1646a1dfe94da5649af62d9c1dda3c6db
zd56b1ca6636da7ef808712ab675e3e414677d9aa8e74712f9b0bc5c8ee2b120bed4085f5d91f41
z1d8a45ed2a842e3e9c6d04b5fe08318ad6658828f1dd47c8af38d35c71bc08025b630e3f618a04
z728e2512479a8ec38752657cd387fb9c025bb618a094f0e2a91c3cface24068891c68ff8dd98e6
zfc971203f036961359915a851c2f4105ebf5636dd183eb7205ee5ae1fceba8e068f94f68b9d56f
zcbdf83cdadc058b67cfd34312efb86553ce7630ab3ce79851dea9a3b25edf8d90d824e220093c5
za8e15f894569324697eddbb96d15c0f14e6db94c2d542a32468f605e3e8ca29d9868506b5fd579
z9cbc55270f030ad8b5e4b38201de26fa92effc1afd69ee10563cd6811fedb88db444939cd7043a
zcea5ae0f4cc8c86da616c6da9c753355fa6e54df046c2b5ceb27f4c73116f230845e981a655d36
z3276b886c7516ceb55030aef91ae5032a353bb5d9e253115fd19a318e709a4528e872552dc6a20
zd61e850befa95c5067e99e1f1b2bbcf1a086e4f8428fc118bca4a4c618ad3f60b1b697f529eb8a
zcea3164b3ef0261ae3ec7a1be22fbc5d80885f5afefd5b4e105f723813d02b79111e925a2a7e60
z9b6e2b637e51b135bb0dd05eb672659403a06bc64f58d38001b403c89c99e12f24de083cc8af52
z3a12c47cefdc01ab17e01a94b70c34125019e49c38a744a9167ad225f6af9d758a17097ef96c2d
z2bae14402a14792ff67c3b4d7a120a0194f1a75f233eeb0dcb8167aac7d0844b5f25f2f486d967
z4e7f986a3a31b05ea4fc43c71ff02e2efaad2de1de319c7cbc6801461ed1958ce0203110be12ea
zb0af67b3b404f9f0a094b0d37afbe63783277e36245f5502183005c4520bef94738fa2b921228d
zac25840a00bfa08fd948c55d5fae8c708a62f509c9552a0431e6c0611f735ad2e9622486b2ac4f
zbac9951924ffc22f1573ab1d5d0512eb8eb3a495e084d2cf66b0cb446b312e06e7bc51cba836ac
zc7b61e0f37b9c6f159e66c1c80c0c9f61999509a096c34e3e262894bfaedaed1a73f6165c802b5
zd9f4991cd101642d3a1a268c745455b0f3e2a8bb8e5d706637ca45071d9848938b6e2c1114591f
z607abee8455b18cde1ab3b36af8be7a775dd5702912857fccf6ccf1232daebb5f9e3d7aa6057cb
z2e1e299af5c2bb502ede89e33a88f174c44818d209d8427fcdf071665613ea9ec10032240e85d3
z4d8c407a3b9afdbd258359cf1fcd73d7f96026f330c8acc1c0e4bc25488e8f50f2127eea769c6d
za751fc334bf0ad3887a4ae91f794709220429c1fd97c409ff00643e0f26abf0e4a1e87ae281f49
z9db46f5f5ded11e3c2821710811224051035ba309383c82c64ccb9d7977a7d381aff122c08ef2f
zd4c781390eb5fba227134447c18f0ebc80271164c251e9111376348a1aa667e02433d5c067de65
zbc112a93184a671dc83f511d5b87ae19297d1d33ad9609c4dd408b9728b64747e1356eab5305a1
z9e50d0547e6f8407039057521abbe2f6cf0199a33cc671a0513f2565357bea682945cbaec0a5fc
z5f63e9b4cba38d0251e125bb8c3d61191fb8cdc1ee1b1753765d66b3f9d23aa6681a5dd70f9253
zd80239ed0fb79f5d805b4bbbb31370023667d60c5a24a0e844edd581e6637b990ebabf1229ecbe
z41f342009b23973c383047f8684f42b1310f440a123624fe9b5be167a46fbeaf52517fed6b1358
z2131d139b0d745588bbb5483a5f3a6bbf77c578ea4f5469d79b056708e017c56cf5d032dff29a4
ze9d9f573c562a1a5f52fb90977adc651936b2c58340079a54126cadd43924f8165e7cce307e064
z5e417d035f46249ee7b102bdba3ba7efe141fb08aecc2dfb9347e3c65725871ca7d47c14692cf7
z4cfa185b3c564e6ef3178a4e7754d3bb30b0da4e84affeba8685c842fc25abe87af0c26a8beb14
z16a26667501f78af2d5694f8e7390b839ff309a3061453d5852608c241014b3f07f156d590f811
zbbb38f383a434058bdc4fd290c9ac012531c15b57767c58c94bc687b06ad339a2ae0b30bc3a115
z9012fb1b8b5c5cde497e57f1429a4d56473c0b463811e0453de3531a388e60eb2f6adc8fcadf65
z3f68e6a81dec8227c31f560b57aaa70586191c339f946110fb6c782d263b2fa0ee3b1993e36c2c
za835fc91531a0e3d97e4f3a7cdd11a55b888b80b1ece6e428c3a7c9a44042f6e9b371c5dfd29e5
z260e78cdf046de88c9e5d4b28a0636c098baa3aea7e3c8c428e5bf7ab7e0f29e769b4f348b029d
z0db210fe246ad41436710ec9ce43731f33e22e1f5f69141543ffe20c68f6b9cdfc0ee1201f3189
ze0abcf3f767ffb4a999eb5559cd77f9f057c704428c30e370d866606d52cc95e06b896e3c666b5
z5b0c8b5de880d01555a2f700bda54e54564ffe4f14617df5ee3379fc28785aa00a12eb68cca1e6
z2c67c5b304e218ae9a0b9e697190e374a6a5d9101fa9e3c5a4494dd9b4968e8699061f303de12c
z4524e674df2493889aadca2530e7d4097e5c6e9c9c86d0503e7a27dc0809633588f101f68d0616
zb053d64c080e307ba614b24fad90a8572d3d193e40cfa4db7fb8d6b95921635977c7013213659d
z2075d91961a8cff38ffd3e0f731072c018a6f0d475a2f635bae70b04c97d838e08f088c5631839
z8d75934e628c75c62ab3e0a385a0477f489ecced91a605ed7bb07ea95e3bc9dce7fbc82331eff0
za7c733c1496ba663f298163fb4d839334c463ea686f893053044e8c5d7b6be844354d2ebb13d2d
ze4e5026eb1e50f5855bc49caeb066998bbe87bff8aeb062b8b2b9eb68fa201c399133282a5e049
z4a3bc9ac20d41a2471437c6905659010cb7a843920e49fbc1e45a663d11f3b8c60f3376fab1675
zad0981843b08c05b44de3161e6b02b8e19f2f2ef9d32f1efe0780f86ff34f80292706e852c98ba
z65e080f36710a25d45acb5a07356c054e1d4a44b8e65088cc2da9b9b361e4c56c57c57aae639b8
zab588fc45edf88c1eefb439b9853e850e97c883bbb15b9e7cbb5dab78f164df576517774d0d443
zcc0ce5381dc2eb6325425196d01f17092b14bb95c6dea9632d53c6ba4a364e1d260b5aa84c2a76
z73f5a687fe4e836bda508fe9abcd13b777d2b12650d9181ec2355431d37aaf233bea91b217560f
zb98afe1276291f0d871cfde6fbdb1b212b075bf55b0ebb2f3e284df94acc9bff050cfacda80252
zeb4f152c4b41b45bb863b11282d40a5cbf522f6cec2f71174e5dd5a2f1144662d275ea505fb68e
z34a8717491c730b490d625479793617c80bb46981450c2228de847613e46a6407d3451869b745e
zdfb5e313c05696c102dedb6bfff5993553596830c249919427c2b18f488c7b477059953542e9cc
zdcdf02aaeac09d25494c7468470c2f835c7d5404046891697b345fec6ec868c339becff0b462ca
zc46f1acc4e5f1c5875064aa9cb7c601a300e1c958655aec8635385f33ec7e0ec3d829432da17bb
z99f033fcc7be0302f46f611e20730544e7f06f32b887189f347b67ea2990dba67d0476555237f2
zbd5ddce05ec35fc9233150808526daa871033f5c504cfbd5b95e083b5ab9f1a2a039f7a5f7718b
za7fbff74d82f05eb9fd3c0c03d1607134202b1c787fae23bb91309930895e8e7fe08e18f6631c2
z7d0c3031948469ed092b7feedf2f7529804ffb1b268b68cab7bfc04ae1d9de1439ad3bf3c67111
z7c733572a2e66cd673dff4d9405a721d19d239b88dfed467fe457773020b73b4f4bbf8558246a3
z2aae2b2cdc9d75910b9c9050ef2a269e387a7d2c86ce2c33dc8e955b6b9e8841a92712c4d275da
zc91d68367c2fbcef3e69b81b1036b5a4301240b9f9dd8c7e9badb97f18a923b9dc79018ed6a774
z25ebf126c67db1cb91d33d2f42589674a08574982d1cf8be926b83c544ded2476daa5c12ba7e82
zb80bb1f75659b9c12404c5ba616cb204daabe3953c7b7e58304fa9b0ec11324a8e8bd6c7e717fd
z2fdc64f8ae06b266963498d0e28682c179624a614db1d9f98043ab9a01d9f2261cb77e6ab83df2
z67e054d87e261be3473b671f28225ff5b56d299e78361e75eac97db09837da0484a17443f5b3b7
za1b0d93d4691dcabb69910afef8d3ffede31a102ae22c68e31e934b7a304b6e21dc0eb33dff35a
zb23b9d0248b4a9f17d82f49c0dcf28f91d39b230486578d93c46ea3241220d61763a341cecb5ab
z950de1a501cd35007192f94df4824aaf534110f1b7ba7f2ff441dab3dd0b86b4b30dad28d2ccfb
z2c68b311c8a8a81aae8cd42a4ecb0e38686bdd45b8ab8b8c385b7fb839265e9bcc75a2df43641d
za91fc741db9eb03f9e311b64871394e7001acede0285f07521a6d404f44a955f4c50663c517033
z031456215f6523c1d019864ef95edb5cad30fd45f86b3fc7dd881f8e70ade8c6df1887422f218a
z5a9828522bc371caa44b58424ba01cc4f3d985e4c5a6304b03726e1aae5eba520068b3fe451d34
z1fd0c28409e648cbc0ce46124bfa3bf13b1d4295545d9925e4b51dff5db0d0ee2359efa62d895a
zbe1c643f6df8d952998c8dc405b5df833766b80c5c6f72a265ce4e2c0cd47a3f231516816e8c84
zd674cc71aeb99f0e1ee04bbfb9b0abe2400c5251ffa97a42c0c68109afb76adcd2103975d55e7e
z375ed8981b3749db47940514b4b530007ffb5acca256804900001675b4b8ba20fbc4ac367cca03
zb8e0990fe6885020652ec47303889c2bdd757e3fbe0286a566e568bd30f382a988dca2a2fe2c71
z7295d9ffb06c9e4a703830f6f57f1a1d9d5941ec18aec22625868165de814b0bbc47e361ef1565
z50516206efaf4164f596e123653c089d0e85eade6973869865f7f54aa38d8d143d4978c24d6ab3
zb421b45173039cedcab5b2bfe1c285ed338dceac5cd691b80d7f02754f3caf66b329b8bbd751b5
zd22dfb50760d63e77fe6a097a8ce8bfe13e2517c671ce1100db25562568611928f060c9dba69cf
z312497fd394f0845dae0d1ec5e108b9e192a621b7b0c8ef15aad065929c70cc34d2581c4ef55c3
z123b1356f90c044b6726684f83e84e21a796a352f084702bdf8e3c1ba58966e0acfe8e782c4ce7
z60358ab4ef940ffb86a08552529e531b441b72b6bc09ade98d899acaf3c546c4512ef459497f00
zde79db404c509299fc229d3b7f648d866eac4c0bf5740aba383ac3dfc25029aa4048fd904d0aa4
z64ab228ea3654763a41ba34d21f3abb1cbe6fd83fdf05c8913ee74b8a7a598e1a014a437ea9908
zb43bd296ae406c09a43dcf5674b48695014073b474dffc677657451644a57494f1d783118162c6
z5a351be578a7330fecb0c06ca11ed37c14b772292c4fa660361b60230b23fb5bd714e61ca069d4
z58d41b737f525a388347c1758cd62b25876cba21895ab568d28e9dfa3d40d1e11debbed0ba6620
z282dff2e14d85e4eb087d606e0ccdf6b1672678cb6292c71cd6ad76f000c71cc179a184c98dc8d
zae28d4c2fd974f0a69945f41d3ad8593ec156cbf26fc817ad5cb729ea5373e044d53cc6a8be1e5
z6765655c44b6748490220a35fb708a0f272f4be3d21e72a799fb272029a38b62d7dc89427f0f3d
z0d980b7954b99375fdaa0f2cdff9541bdb2d51eb9cbd9acc3ae21046ade1c86de096f9b75bb5a7
zc2aa48d538b8360446b4d91077de78969ce82fbb90579322e9113ff667287422cf9588d2065865
zd6b9fe0fbb02f66d684d91528ea68bd2a258dd62e9f499edd930a628881d7539c5cdab86e70895
zc723afce84c513cc995474b53aa535528470b8eb4025c04e417762c6334c6f840d8f57e015fa2c
z328cd5d429aa75a5b297aa0110e6e71aa233199395440bd6e491ff7291cb4680a1fffa8425c942
za5b7e8c43cb000d67b3950b6a6c853731168036786fd559b6cbdc4d2abb9e6348bb669011bd6ff
zd4d948a281676542ffc5168f4dbf454a8886676b3768c98b79d125e67da59ffa34f8d6afe57282
z7f43957d7e0eff4b7052e1117407cfb43c5641a13cde5d2ebeb920891188e285b0d8112ef2ec38
z0525561bc35cdf2c2aebfc819289cfb706af50d02dac5fcea7fcfd9afac1c0393eb35016a28af1
z8ed54135282b156a28f4519e35a75ca6dc0efca64f8a718eb1b8db21e5ea89331bc28e54f661af
z8d57f3783388552bb2ee632b49fe27c862207fe6d1c4ee26cb1a89b551debf3f9153460af36dbd
zc53c9187fad9ade5c50e9faeff591eaa0d47fb6742cbfed39de90f31689f45d504b58710262822
z0339ad81b50b5756bc1e17ba1fbaa8938bbc8055cdc6bea0de3245329bc9a845047ca16bbbf5a7
zb1484f03a8bd42cc6a761acf8fde274f8c3e46ac84d7a9774bd0c17bbd8b067c0ad159ff2604c6
z76ecc7a4775eb338c33925c2615ea8bcd226b2245e2e51f9e81d716d9c11dbc9436877746f4cb4
z3ddffe156225f155041efe3d3e2b10497831e19e67107e3dd37a8f3b869322206a191922704a32
ze5c3001cdfe2ef3408ddfb31a3b4ce1ad6774eea570386919ccc65dab892a5f32269ecadbf0a82
z49b84faae863953618263fd70d62e4cc05c62d2e66b98db62c487b124dacd3618df348249407cb
z359a43ab99dea31a5ff88c06a04decfb697d1ec2abb1ac08c1ab8867d98e4b80c0c9d7664248f0
z1d3db84f328ea159b8550ac60b55527f651d08aeffb10de4719bf5da0cfa192b9337d9b1a0b1cd
zbd9a891fbc629bedc60e9a338c1921e9868d7bdbac5393b08aa11176e1aa5a13ae642e83aa8325
z3a8a3deeeb4cb0157830312b341cbf77fc5ab6c579b317720fce247af923964f4370e96fa4ab41
za79355470341c812f2cc89b76639d95d7384c765ce0626db679e25d3f49d4dec9782e535524c2c
z1c3aad2bc3306f7843a0f3b0c9f4ad74c666342f0380b0170a2486495cf0b4120ed83516c339d0
z0f094e05c41b7a471f97a4c25750acf6a1b4699a0869b463008642fdb76028a77ee8203f40e975
zf376f3657da410a2921bda2779c93832029d19dd80c05f7153c2825d04a0a2d2b8872f4ccc2d41
z221141eddcf4b33e5a7a41b2e9080f772d92ac4e7856e62d570824aa7cd5dcca9e054c6c397a83
ze6e0afd2ccb81bbbf745a58cca76771d12b845604eee97d461c42c7c9449b8dd6dd2deaa53cf8e
ze733f54e456d20975357b6a4a7dd5667665a6bcc8017504fc31b604785774ed75400925eebfc80
z59fa73147b904d7c69a9dc10d036288f4f2acc9732cec5a18ccac549e49ef7b5776daf4a9de45c
z93075554ae6bf15ea89c914b41f55d025d415ae028fca0cea5d71d6b2843505bb9dcf341f2ca53
z366cf7593cf402135aa4a0bf5f876d338e48f661e73b4038debbf193e5424fb2edde835b54dedc
zef0da0c1ea04ba24ec9d0377933022511b97c68ad16f8bfe60c959c89cb243861539d7f4464ef4
z0222d4764967cf55f8ff66d7c1039b7a5eb8e524a8eb571f97811c051cfba87f0c321972cbe005
z8a8f597ee7c6aaeb316f6020ee5439f33892bf8dadb4d29619a1f89f377bb6d9a59f4668f5625a
z722d4a049cbe3fbcc292832eba6426f91358d47c6e82716e48748397f68fdf82cd4e3f3b891bad
z58ae4e92a09c856036c553e4f098e5ab8759151a8c1bec9dd17c582c546379f205fe13202bb5f9
zefc41b8fb722ecdeeb23b63d80eb6d72e9af91c2e5be7e9ccafcf3f04be08c07e60ee389c9b328
za4253dad17ce8984a1c781f1dc26d80cbdec1db730552182b7292babbe69c250b812893747b78c
zbcc27a801bd2667f8f8a32b3bd35933f12d94c49d4e088fba022549f770f5637b9aebac8633e32
z3bcd8917796baab41dac574ea7e75b1daba3a419c801ad242abec3393a28d5eefafc382c2e11c4
z71407f65ea517d20b97d122aa50444d81891bbde6bb355b567bd09e3d62d251416ea746e48367f
ze3b3203a54c156fe480bd2a4a3ccf13415a9d065c5298d698f9456c5c72f23588b38c523bb5741
z04e967e3ef2bdb9efa261ed09b96e45f43c06f9f77cce59c7c8657ad0084f6e0248ed6291fe1ba
zb48d1e9ebbc10679ae8981e80751390374727e071a5883afc14a187de679c6662cca174f7dbfef
zb6076609d7542f6cbebf575afd9acd145f2cce475d030b76a435dd9c6d436d02215da1c22bd367
zb97d2c1be739c51d9e35b3425c53c1c48d8516b52a380a65580abce89e16eaeccf8fa10f9e1956
z39c4794858544c9a927ab571e4e0077bdf6016a547a9e961ce521caa3cdde5e3d467da11f00725
z044ecb33fa215e833b40b1f476f3fcede4805a9d2904fe022f012a500bcafc74e727cc962011e6
z10ce7c2e576283fc047a4cf6bf26aa318b83bbba572640675821b22bbffec60b5e11c9a6f6d7c9
zc55314a91aa87dddab31ac49d06da0e0ca0e86c1249b4876dbb55c8dfdaa00d6f34b59a9c473f4
z460bad52a4dae7f386838a9a40661d3ff53039daf9640ac399a8cf7aeb4fe98b64a6bd3c1b58c1
z77c2f8edb512738d8f607071e0d2959b58a906ba0ee379b02d05068fc5e1787da8c36a3fcaf093
z60c03f1bd975cb8da76c6138fcb4a0d7d0cec12de1cbd2db2e4713a01105d24b3975f2418f2d1a
z384d799e41672bacbbe2b686f946d071cecef89f3c98e26b74647b9a0af2d8f1ec9e8a77caea02
zc6b331f06c7584f496eba8adc908d2bc7da7c73559e1fd14c49330ed5c8a1ab0e5c7ef7ea6ade5
z36bcc7836b51feb4be8b48b515603e96e41733fae3c9459ad67e6667bf46feef5247479b7fc69a
zad34baa20abef780bc912789f0242896cbc7935bb9f8ea8728a1f604276377ae100e1b18f6a985
z8493770a8a952d7a4587c3bbb33bdc2b2759014f59e81cffccdd65894af4c13e9e352e24b4e0b6
z088af465a3ca273326c86618d89714bac563214bc6936dbfdaab5674847147da4d461882413be4
z1b8088e46f0bc2fdafd21577e71686ab7e6c7ba954700d9ee068ae4ca0b6eeab70bffa3882febb
za20ece3c21d7d0563cff28260f5daed6017e848718e761c57da699d2305f357f059f5501c1b4e7
za08ef91588dff4739bc566309597f809f470c92ae49a3e88ae12047fbd0f0a8397a284dfab6030
zaa7be83e344fda55dca0ebc342b05e24a5dc38dc1d7a5c38b8f455e151d7f19766f51559d5cd42
zd31b2f5f0252096ccf99c0cb3dcf779ff7409e5e159115c63a6deb7e64181ecf67dfa482b2c896
z05f18ea7ccf7388b6e578b5b629af9c0a0cd178f609a424b957fba9dc71abd1516e3d770b80044
z3680c574f1b0ed47899d49823ab81822632e7c171f24d230c3a2840cfbdc2676c561c624f5ee65
z02fb37574c510c1693e5db2e95a225ec4268a49b220b7c39a3e4e30bf5af6cc0464cf7649ffe0a
za754ed01908e5b3dfdc93252f5e98c756315ff21b83c046f61b8239cd5578a93f4227bc3b95587
z41e3069c1b7872c143916859a0ade773459ec63b861edba4f9c0797d16421d1132db1ffcf9d203
zbfa111f688d984fae28e6c31f9a8cd3bd78475aa41f6b50b323936387005b7926051d41e2e40fa
z735478db052782fe78cc46c3dd5ae6f8420e84a21a1ae30652dea564e91d0a4f12bf7dbd7ea917
z67efaa1dceccf26d49599fb66d63b1402f410bf6c1696b400eb3e95951538e5b2fc22c9ba821a3
z2b3f2acf3448adfe0a235885e95b9ff266fa866c1cf4972c161d4847227a76697a35d39c730a07
zb0da104d7be6ce35e02488a365f0e4a35579deb7ce06abb5733ba900dc276b10285f7b1cd3d044
ze56f75e284eda63a368e2be5e4427fc2dc4e92f1158646803297cbe148d1dff0fdbfdedbdaa9ff
z21b80d49c7a8cbf3a52d19117ab3a29caf5aeb6a4b238358965b2dbea4115e6d706eccc31b2e26
z06f24897e7c88a3515364569a3ace7db323aa31a7e485d9eacb4147d4a1411ae8d209aecebd11f
zfc82356e1089970c74e5ccdc927a0874b9eb3657839d320944377a468682f628d1abc0caa0a7c1
z97a8430a922793d5bc1b8c17e49d334482a80ebe8843669455e3b5099f1d8d9b5a41fbbb18029e
zd2a9068c9ceb31610123e024fa6e54de871294fb1f1b3a4e9c58b829585f0da8aa848c92eb4385
z7d20df6ebe3e149b88b9af27e4d5688435561a80a28e869de745ee59f85ebd74adf25d87f1c32b
z3504643eb38708cf20784465c0ef62c3b913ad406101a4ae55e099350ea5dda30beacf606b965f
z908d7a4aff4b437ac1e2632f36f29e2231bbb7c5de19e36f379c7bfb9d4ac8fa741c56f9127546
z8146eddb6406a11b7528218bd9dfd46a330668319e7fb42383b7e3232ae7f63bceb22afcdb6281
z36c00d8002bc325738095c07420f99e332b27583dbf43491b228251ee16bd043ba5f56ec4f5e29
z70ad3b594581e07a05b63bb79c15e4fadb1e4d4da696b789bb9344cbc870e4d8713df5bbd710af
z7666cccf545457b05aa2cb0fb57cdfb3c65d535bd75e8fedb8e687104867cc4aa5f07e39c90aca
z943d96c77bd16eb833d7147c2aba7f9579f266d84cf35cb3a9b5d75ab697571f8ade0dfcd3c533
z5d8b8f0afa23f7a99e0ce52bea4789173d5592e2258b96c4634459f40dc730c6f9b16eb5f5e872
z505d545dac90154988ad0e194d4ddffc4faded06ad5397610f488157f27fc3efc708ff711a62ea
zc73f6fffef83d0582da33f6aba4c9b1605eb4a819bc87bcf6c00f1de7e32ab0d6c9c70d7b811c2
z5f2d9e1831d9ca533d21f3eab97386807f4964b8d48a53b9afd1c81eab9dedfe64b37b724244b3
ze6e9e2c78db9ac808c31d0ce359e8959b4c1ded97dc2388a7e2e2dff57b64e8b9440c95f7e4be2
z94bf1f09741c4b6a3927f7e62b8176d6076800c470629bfeb2f8dd95bb0cfb9911b853973d62c3
zc800e5b9bfd76cdb39273277e1f265695a8e73b4707a88ac77e6abed2ca54c74f26384b1f862d2
z60e21b14a61d3be21ae8777118f98d4f9cce7e18a8055368dea585836fb08b20d0e5336cb64c37
zb15234b118bafcfc8bd46e6d25d2ae5ce4071f97d9fe56cde2466a5ffb13cc45a937096ea5f027
z6379c653b284c9f18ba8b3a4a14819984ab98d880a5dee10e7ffba40bead67c2b5a330c230b864
z97a42b01aee96c08209a3e6b07a38ebbd23fb036db88b4c82b12b311d60d01eca95f8390a89639
z214b9a63a1e6063a5cd2165b854e170550564fcc1595b17e95b0a0ff4b313fda8a530093a4fd05
zfed256ebc96fecd7c04c18c660a553c5574cc7dc35a5cb2e234234c2d23cbee2108a2a018cdc31
z4ccb3ba8b2092da5db8d5970823c698193300d1bb95fc07fa005561993c254c8fd84c234fe39e1
z8fa35831641421f5834479bbb24d68cc3378dcc509418e65f07ec1b0809516f157c26197de59ab
z2e38fbc54b4f421cbc9171fc575bc13c2200946e3fcf0a99621a49f1f379f5434ec6a8a278b845
z9e8a8b51c4dedfa5cbb4ffaad579bbe297464935f23a7a134f1876c878ab04c653e79fab158c4b
z5fc0cd649fa151cf35872dfac8c2fee8fc69632aa05319271e5df7a6d3c7c90552da7aeed1a700
z31a9f62697c08a03245e76a5b7f131be333a1d526cb47101807fe9ef57a793d76a5f682dcb87d1
z6f072dc32e3d563bd2807f9923bd95600de14aae5cd2e966b10cda975e789aa831c222402bd85f
zdfcccf897967bb02504f84e0a6c23818ec5f9fe845618a6793b196df34b450b4f31a80f9f9c66f
z74c794c45a87cd84eda44bc35ae0ff6a4814699046e9b3c284605084ed3aeebe09dff3d5523d3c
z41bfa96fe7610ffc15a3c53d99c215efa336feae1503e3dc11decd3c86bf60323963f5f93e878f
z024362d1b5b9b195b5d435b428f6f39b985189d8dc1b54e821401e66b88ee761fc8b9cf5d1b2ef
zbf02a9e27792537f6f40d9b073d2259abece5ce96c0b5d8699636c04283cdfb304d8f24822b6d6
z084a15baf15641f8b6b5a157a604360bac5497404cf089edda1a568788d5f1cb6844bd9c7779bc
z1bdd6843cf8aad392b0d3f8c6fcc1c8a35d99c85236f49572eb11d98e3fd3d56fd36b1b1d5c0b4
z57a56abcdcc58dc7931abf8d735da6a230c448124b8728caaba7170e617a73844548ea24d4df9b
z913b6efc8e88660266915e69b6e85d10ae529958f04c77c27a1cdac907d1a8bd9dfa0ef47c8417
z5081eb65f2539d96998d45a5eabebd0d2acc04ab10b3a08864f53b1e5b4945c9a4944e0034ffb9
zb2815b8820d75f8b73b9aa4517c9be7e80add5208b8973043dee32b272bbffd93beec920c33c44
z08e6aa41415a4f5fcab001de74b9d24053a2b5f964f13b7b3cc85419f72ccd498513992255cc0d
z1200fc98aee4d193ed168855cc18dae511a34b0cdeb7e6a7cf1b8c0db766c60a574f649395e98b
zc54d854af4274d54d731b867f127e39ad117337afaad3b34ac1b35f0f6356be08a0739681894dd
z77755d4cd862d05fae948442ff87ce1c1d293863bc0d568f72e9107a23a0f84ad30cdde57d5417
zc31798ddd1a315d95d9934d19e12470c01c32575f6b59a20da38fdbff184135f5355ffd9f1205a
z5406be32aa374ad8b9d1f5b32ca8022d14ce38c246db9aeab5590d66f3250d5a318cc0a7747d6c
z4ae61d72feea81061f7deb3c8ac60b925654fb30700fc3fdc227cd5062f99d1e1480b056289cf7
z50ab9ce950b98eb5d690e40f9719a99cf7afc33977e3fbb35214acc77434a2f8d43e92868414e9
z91b0d6920983c13910e69b1375be4f8b027803f7242ec9dea71cd587d1b281c8f9bf953db3b0b1
zb59403fd07740809639fa718c929ea4db99d48b1a5b18b6f12ca0179f4de4c5db0175c54759171
zc8bf429ef909b116b3b97bedaf363361da6f3a436c84949b46c43030f380a890b4671b6afba14b
ze353e785400a2fd9072f015a883f023a06f0011b8123b44b9ef827d6c7a6bda6605c2dfb1bccf9
z7f5c7f51bae3552a12712a622f81215d5ad519bd1ce43641a6ff71fb7c8586a63c2c88623e1904
zf08eba25cdec7b729502e9fe06104472924432068df0cab57e4adf7e6481dacf3f3e5c56f418e5
z759bfa3c726cb26839a2eac327b838c5da4a8d1087e92807101507d3678779892d73549a398fac
ze15778cc45b30dab93791048a94dce82693a09217b74ee284cd01791e3aa33e0f3ff72f806166e
z10ead9232b22558fa29be445c050b8d4c78d18e0526954f407dff1bd129deb5551513c279e01f7
z98019045212aa66579bc409e04419205237a9ff16831c0e2f9e6a2a82216f70f4e89a2b63a34df
z6da3294b230c0968ea9803ec08c005eb0a2501cbf1a89883301b6bf2b83075a33285c8ff911338
z26cdbda1623cc99ee12e0becf5977c51fb05f4ec82bf1fe40efadbd68a0dfc2f0777810fa6c6e0
zd38bbe4dd8dc5adc0218b84dc889b11bc77f4c7e26ebea232b42c51d051c0d9b33479d8e40cd38
z444ac0779ad0d353c88448cf42d44c9987e41bbb705a6224ae31587e22d6bf636f6963a3402b25
zef991913ba50f0d1d2e394b40b4301297e4c15bdba173c839c1d2a830306f6dfa3a24a19fee908
z701820fa536486dfdebe1e8fcc9d7c3ba7507f8217f303edd7d246f74beb21abf0fd03dd289155
z8a7f24b3225b37e6e4eb5888ec57838e42658a5b432616fe4422c37d6f2acfa159b30999982ee2
ze340fbf9acceb671246988f4ebb4c787067ba6e9511d6fe79fadf2b8122477a83cb0b9d64dab91
zcf77508f508add1cfc43bd0ac216a55cc65fcb66b3c5e2c78dd67a862d18ec668385bceba6062c
z41756a2860141b82a8662b1f5f84d8560d462b04fc9b18c107e5af3e3278e978b26eda177dec0d
zc669b01747234d6bc1b0e2992afab187419f75a7bed17cf36cb98d718e54415478c6aa3d489d9e
z84ccd74e8842f51d3fa00a25c16fef8255ab5cee212dc01f11b7b54d8093fa5918194ec93f6d79
z3ce4c9ed4d903e0795f58f78d99ac02e993a74da88f42def1bf601781e36bcaae7d7f666d9a46e
z91c5a4470e66b9ad73e10618f55cec904366c5555af0343ac65864c8ade111923a057a57eeb099
z4a44ff3b896482c116b24ed33f06b3f832a263e3ac1bd87cc19b5a25da1f70eee4d901ba9796bf
zea0b99519c5aac39465cc28f92addf7a0b4d2492192b298407788abcb99bfbfc7187ee5305ec0e
za23384ed66033cacf6c7c1da4c5a2b82ed9c97f7463c0d8620195060575d7cdebbbd5eff9ba336
z079b9fe47a8409a29059d8603de7cda7c0bb1241505b0f93736dc1f99a957271236de2abb8f123
zd0e7d00fc83d0737a75b5b98042bef5f787d68c2af88edd6cdf218b1def42f56a862cbb12b1fba
z1af517e26342f1114c5f07ab164b280c7f872dd96b37636c9651475a16a2b8b54652535ffb07f9
z23f431a385d3c87571c20ee43198874c7c0648c8bb05a06b71ff8d813da55b5b6707246c58ebe2
z89c89fddf3fe8b9ff745397139d735ccce5b865ca63cec9aef0ebe2d767abc07cd10e5108bd169
z54c103a0b581736b53071788ec90a8825f879e60172adaa7453f9e9c51e0c2777d7e4fa25a9b1e
z690e22e4805c65663474ce1d535c8689de6de006581e43a1b44108c0d394f9d16145d9f3443a62
zf1f48e30e071ff292a9513d5bb403075299281e9ef200e3321155a19596d67584fd243beea6232
z28259e9e9afd72f51804975b4f38041c989a12075412321a04570840fdf09fac64be138d1762ff
zae02abb68048c2b2ea99b28bf21edaba0e3f0d95525ad8d7edc674d36d354e3e6e15863f7b810c
z664cef54ec4f22c187f885be856e0daebaaa7e186c564e5dbbe9abe0b8f4efc69639171706406b
z4d409b138a79e398882c973176cf916c3e35dd69a5a009a5c579fba3f9ff1f670a0a131828bfd0
za6e06fc7a6796b3dcfea843d30a80fb039d862251a41122eb0f961cd641df73f6f54e55bfaf373
z25619ad84c2340d8cba59dec9c08ea3034e9cb3f3ee613b767601d10892161b906924887ea5a16
ze7d7bfcbae0f118894b92c7e2cdda952bf46c210cbeef11966ff70580df1bb28d40218ef6c90d9
zec31f23b92ccc3b5fcf09702f083388a9d2239a6b7269fbe9039c09ed191855e0a8e00c72c01f6
zc073d7dbb7de3047b8de646d040808060148bb9abd48e34dced724b53fcdc2c11f96d2cfb2f0b9
zd57b2a9c53d86811ffd4c438166ddea343aa941b7213769747467db5795c507ef65e9a6be47279
z1bbf5328d05b5b33780821df7b8ce2921159eff9fb81e6c896073fde1f848fad28dc09b0164c81
z6ad11b1154d39f9157bbf5b93c6eba1f
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_multi_clock_multi_enq_deq_fifo_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
