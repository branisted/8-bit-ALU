`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1bc235c2ceff4f6e3b1ebe72fceb7af9adc96a
z694b4bad7241bfbe775016041d7caaa74d9c0e7b507ce89e8b01980415bfa35a8e346f54c548f9
zda8767c02ea87d27eb7a843f4cada7dc3b575fb5cede69da7a4701b2d725c73f1f7375e85a74e2
zdeae70c30f1127407402c955b283d7b9512dbb3cc85aff97f613d57a4efe57b3c092e5ccc5b6dc
zd04e277cea6810165bcacbe3f515b3d75051fbe8fa4af7e932d60d2b2a6cbc14783b996db7f97f
z0df4e054ec07012afe312c7c27fe5855e396fca2df20ec96282aa187aefef584e73225c3183714
z599297effba6810dbfe57acb29d5b025ac9a8ebc73f537d2977dc34b086017b79e71d435e90724
z58f8859c47b62c6b1fbee0ff19f88a66a8afa79b5c1920e87193650fc0cd3c6ab3d109ee7dddc7
z162107ca701eaf77ce18df51d1be11c0dd907a4d1366d43e0990f506187b3d9bd054ff243db092
ze701807474479b37f0911dfeb69e92838265d0284967e78f0d2051699430d6e5af93353f8a4ae7
z1c7984e0af29da5cd55d0e97dfcb42d4a71e64e6191520cec069152d02ad57291a620e755a98df
z6fa6dc8485546bbd2af18bf3cfd459437fbf0fdf80856bb76e4134572651e5be5debc0ba0a422d
zb22a56d6375c212b53f403b92b101660c31f60ef55e0f523e3c42b1912d207d2847c2d5f589467
zb0564bd25382cf356e2b913bffb723d2a5947deb138b8f58e3164cf9c4536c5892ee1fad6f37c3
zf49e4fd11075ac2a1d575a56df2e5e3bf605f3625e5ac43ca6482dc39f676a2a3423c5e7391bde
z9690bf003218e83278a8be82fe7fcf4cae5fee70740bd187fd620d6dfac2aa24f24cad95bd9e5e
z088a29f4916d902e464213cb2f1ad49205218054572751f2619e5af3b88e679ce12c00a6049617
z9c306e21442cadcad36b02a1fac4e0c0c2709a15b97471f83f51fff4ff881e6d8fb15c8a58a2d9
zf91348a1697e8aa18a29da465a9fcb3eb5c51d5ec96abb403d41a5a5e9a7c78648b4ec38e66045
z5f25fd4b9ab757e5a46ea337d749261a185f7544e29a3f75f4cd3b5c1b70900611f2a85e25272c
z6dc056898d33c55f6dfa9a7b7d21957d9e1ffbb76234a66b9ae9ab6632b62c8f955026f30d8297
zb13b62bbfb4df785af504acf412d8939b80fa7cbd44bcbf56aec1e62eef66621fbb59a0284e037
z4d4be93e5c9b3f0fa93ce93038f6b7a45cd4f6450685f7a8a751047e0a4c997b14280426a96ca3
z93eb868325e14910a914aa837b3ba025fbafe1dfc8ab33587dd65012a6761159f439078d61d79e
za1d331ec25c209d0603be398a62e9ba8f47785841a7ea42a8587976d192b94edef4233532204de
z11d45d034ec0153935917efb5681854a9c141d4109e69bfaff182e4bebc368d51b647c1dfdbb04
zb13dac030430ffca0fa6d62c175dfd9c6a393f850c4e31864d6e62c67cf57903f98521f20d561f
ze1449b5b453d86bcda4bc3fa76455fb29a3b533d9ad83486650b35db1d6c684ff52e6ccce6fbe4
z741875146a7566b57c530f2d40af505b84fdf23d9ac0d4b77b892132e370c1ef6bc811a2942055
zb5d51fc658f1cfee7adf46c218f9332b44d5ef21e649162c96e85272f4f464a9ff9da92d25052e
z4068a8b8bea90b21a773e37ba41e337ce7d34f86ca73af9199360e9105c40d29ed3ea12d2ebd99
z0f3a34fd6c8507e336d4cd9cb50ae256f74745a4eb1397a4aa88f2fbd218020f25d18b6aabf826
z320511d253c1ea31c50904b832bbeb49beb38dd0f74d5eceddcf7bb8d473c2833ad6b60672586b
z56a523a02e0491b5319babb53dbce907abf1b9e59f96e8654e4bccc9135ec13ab425b762817a85
z59994e55dbab93b4e65558b9c17986de488853f92c5c74e8469c6624af39f462ed9a0223dd94cb
z0bbb0ab25073afc613285271c0c96f17f05c146e94a40ec60931712be6f70c801d0bf124bfe42c
z4fd672650582c4a6c9816b13ebf62415d7a2fc1e8bc55f06ef1e217866b06fe2611a6aa5568162
z3eca21e9fb831c87b01f8ab8e1ff9cf447096921c92c210593facf23fb0523b374151059d771c1
za437c7d3b3f92b9d50489513496a8a401d00e030db7c0655483460eeed9846f092a8d6841b5256
z5755a34c466695ea219fe0508f0dbe8692b4ae42686a6ce14cea5bc41d70a0e664f379a5be7e35
zd99aabda4654f240e02e2979a0147b8242b5dec2fa608c5dcff4974c9f68ac349dfcdf1bb64969
z1ce8776e23d4d96e34174e8474ecd9380df4f89767c6bc3052ff2201739ee6bac74016596b6107
z965fb1b211b97d3a4286460d74ba9fbb6ad26b85899710fa898988a56f498cbad2be78b2a78553
z91ff5c650ddaaf2545371ff8f6023d6f310a6da4adb308928e83615c913c2e2290da3c2bb04e99
zd4d38843a26261df9679fc8702d8efbbd33074a15af75e35288f9d757bf903ec5b953723b7b14b
z73db34ca4a7dc01f1233c75413ffe6b20a579df01ddc18e078316cdfd927288071b977a72e5888
z8eb7d849833920e1585e591d45c86efc2274d06b57542cbb18e15ae3718cff3f1105d633e9b557
zf4a95299fe97e0af1bd55b97fa3fdbfdade445d158b63cf022eb3a15eff7c0f628923d7aab9005
z9cfbe899145d2338fcfc44d7effa77f89a9f246c1f080d89dab9b5718f413821209937c49262ab
zaa6e77aa3015186f77eefdc115f9883605ce1284a8f8cafb49e9a134fc0e6bfb690d1eaedd807d
z41bf3c2fc52394b3addcb67fb4c50cb1746e212308d470cdcfefb1da148cf74044494f1e450bd6
z6f1b36fd18519db9afcab7da065b118eeebaf0991de42a0d1ffa0e54eb4006d2bd901732eedd5b
z0cb1e2ee275085136164ba3282dc637f403275a85e31d81e65f20969414a8f1973b8ed1d05142a
zaaec58c3a6a7aae24b6092a1fe9709805f98ca1fd39dd310b551f8ed4d2c1e7015cbfde03b7f8f
zdaf68c36397f607027b7a27554387d55546e22f805736814157919613b344e0e35d79fd5b1b4c3
z6628bb05a7663d45704832f1f054c26f53f8206812b216352517b785717b7b82772477ce99e3a0
z5ecbe7a6f896fa1d8ddde2c0c2ddff850c6179583a050449e7a2189f949415c02c8eeaa7c944dc
z718d59a76ae56b39301aae39762f0df7dda7fe305b4c91915ccbdc7f2f6538f5ff5e1ca4a220ce
z4dd375f0abab00bccaef3c46b517a9d6e7bb94a6cca2570cad378fdf1b861297b8204337efcb51
z1ed284acc138e89a56423adc43b31d9317b6dbd117125443cf2120bc88853e7c9b55095b7e5dea
z982352df0f849745c55ccbf884c457b198b71898fce541cf681b421498f41a2e0a070bb69910cb
zadea1e892c37c0f775a7ea83575e8968724f8e1a3cb7c2fb926c976bd95f3c5c7d0f576494dca3
z5351ba2bdf62ef8ea416736b96d6aa1d569fea4d5e45145bee0aba0b97f9980f2ffb81b6cfebcb
z6baaf34c1c2d80d6e99b110d9bab32c7cfcdaec3753123c5eb1525143cbac0bf620026963bf878
za2d0d1e9c1804875f6755e45819b5f64fcd80433b50be9234229583e009fc381ad396f5f354fc6
z6b84e43d5850b758857a864c2baa58dbc8e7c7ff1cb824d77646d7fb920e04789cede1e2911669
z6afa9a2174af77eba04c7f63c7bb81e7ad3a321f69db52e288e45ed011e77128b774dca9a840c5
zed91dfa90345a0b7bad5b4274aaa7e86ae655653bdd0f94b9ab096c431936e226c06ff84628784
z8c96e8255d3887f4f25b9decbfa7029ea0dbb3d5a2ffbfd0039a3378ce716f623cce0d0937d7ba
z115c8cdfda9d5ca115f5252202c3ba2143e166cd880dfacbeb30f9eccf2aac77f36df1b4951906
zeeeef5c580c9753321316c2b31875ca37456c63c0fda2f62f969dfb271a62e8da37932d20f15cd
zd45fd3b3714d02c21bbc5ef2c20e90baf07fad387bb07a582673f17e303c38331f0254adec12a9
z3845a1bd3e05378f22f0a9e5518e02ac65e22e63b9b5110c3e71a0a0707d955b47bf1385d9f78c
z80570ad0021646a266ef1024630a8c0f8739be4a609b731c9298dc11ee68745debde542a1a8a52
z3385435e3878ae6f354039e0d6e698fe01439d9809237d04f622d70b2f62d7f551d7932077c2d2
z919a39a56ccd3b8021d3b5ec5c5783f2c94ae19066557cc1b1ed860e6e2756f883e28d9b37a587
zd8d82201e4bc0cfde004de4a0bd6dfd604985a09d4973647d0985e1132f151054792d661718c19
z06aae07ff75de960f1a9fd63f1fb2b5a2b0eec1660cfc617202f7d7e2805fab61d6ac7a014f407
z21da10b8a12d09cf06f3c05e89bb22f0251fba78f18d384249d485fae257e6bb5acd9ec4319ff4
z921fd13a5147f442689693c74854f1154ebac7cff3ad0bf22a176e06e4dc59703725b63d48207c
zb5ee2d34b82cc03c47fcd87780b998521a3119ea4d9ed6923bbb9acabc2df1914ca0f6160522da
zbc8029f3128f6b0f5bf8988474564b6a969e3662525212ac1058521781b02606308ad8a274aeba
z7517e83175591d4bdbd2aa87dddce990368e8ec2da067075c5e567ff92ce816228f12ee949966e
zc76d1a0f870a08254ba22026496a741b78a8b056985086bb8e02337ead44ee0a01b8c8fa0c3bb4
zb85599394c6577ed775c207287f1d6bde798da1ca67f897521797f78bfc65ac21ed42c982fb184
z1c80b5091920930b51490ad36f04c033bc2b0ad800d9b74e235c2046a874f7ab89062755646f4e
z36942e23e8e1c257677a059eca3561e05019e6d1f9cf09619fdc7dfa5a371e9d3523c316ed8c34
z5f3601fe6d11ed5dc77278d3e7a2ca70fca7cd16985c343341de644f0bfb4e19e892dc230dd999
z52e9cb1faf0dfa16df3fc39e471d442af9b7b9de266195996845182cbbeb3ba6b63efb68972d65
z803fbbf33e2b809139281b856c27ff57fe6876d2d3d399e3d1171807b0b85e63c17c554514c6d9
z0bb54f76f833bc282e77fcf83c2ad945a4aeef818c0535610fb60f9ec817ef692be6368fa517fe
z86292e3dc23cd214391f8f04b631f194fee7d5df4f7cd75a4ef58154546ef32ea44a818aea19a1
zcaaf364cacd60b3b0fc128cdb4dd1ca4ef3cd837453064872e532303624b05aa588e05c672314d
z4abd5bf76db3a6478231be1f3921771d1e15b546309797d8e82fd080958538747882e1388c9ebf
z9d0ddbdccf9ef3a12cc57ed0739ed0340ac523dff00d15a404fc284c82e81bca81f11c44a43913
z3dda6eff3c7b0d48e4a0e75173fa72a1e0275e060c5eeea042181bea39212ad6b52c2b1091127f
zb5ce64e05c6dd4b318eaaf6e5187cc3ccb6a053e992ae262b3cb79e459d3856e6866dd4e5dc2a6
zccc11279d73526ad741b572d5f0e6dfd05ed70542bdfc5ba7915a6857ec4fb49e4e6339d88280a
ze4eecab4c9df628920b597d390709dd3ae75b2601c4f8337d43f81205d205b3ecd722283044fa3
zb92b3f1447522cfb6a5ddb0f7adcb02236930ce0286c675aadb32a7ff05c545ca6491337e4decf
z3043a6619309abf2584374447a847acba774339db94cbd82be6e00a66478290673c02de3b6b33e
z11015206628781a6b81ad81ab23d675365683048c22cb473b13afc6af5fb317f784e93061df780
z580c5083c1913cd430c3f6a72050cabb4b3618df30b12e06e32295a7cad2e7235c361a567c1a07
zb409bbb3e2db2e1aa3af460be4f74124e9b2aea43da4c18c82e38f8fe4b9d89b079e4daf932b43
zdd00bcbe4ffeca717b0a12f2488ab33c48d4c5f9cab8aa46cd84174ef5608491fd9deccb8c93d3
z948f8c6bc6de69919a3a1a443bcc7bced30b0291018dc99310045de29fc24f0e66249d7ffca09e
z0b107339eed3774ef6a542e7eef03986c594d914d8fda0e2555b693089b6ca0a1f49921149f1b8
zad662aba35450beb8ed04d9763f6a9d93ae279b984ed7efd8ce489324eceb1a4f5a6531e1ea150
z98362173581d4b07da14003d9c6c42517f9dc7bcf89be9c2c4b3665515780fc5e08491d1b90d90
z1cd04b21a6effd09e54c81883fcfd249b5a1f2bebddee2e2ba01cb08f9c1c4bdec48bfe81926c3
z023412f8f9504bb2ff539d1d9624748f38fe7dbc69467fe614a0204720392c09aedc3a87a741cc
z50286b87dded4c5e565c4bfed8e4a56dcb1f9caa284568c500828e1c089b1290a405a675b06cc5
z4466c1c75ecd210f000d80dbde63fa6297074af60642dabe096ea2e7ff7884ce0f70c856861e96
zcaaae76f31ee24eee9bcef4e40b8d0b7c7551b4415233dc019cc38b24e7f6bad228321722e82b3
zb5162a1af0c50f819856765c862cfd1695583539ae5eb8d62ad0c0bc7e4d05442ff48d01f36262
z57fc05e4f4d0bc496dbe39c75a505d75737bcc4bf2be7af2a7f898c96c09e743f7ba4b601600f2
zea5066b0a4032121cf379594f29ed793f3e3dbff70345f3229a25e175bb187aeb3e804b33287ff
z03e4387a04db5cdcf19901580562ae01a788d0a0788eecb6bd0e1270d4ce9337e62c4b31638a48
z3ad9de68e1db62706407d863de55aa03c8aee112cb5f7a4b09a8fd7099ca6abed808057d3c6456
z3959602aa8cacf886ed694b427069094d292103022be87c1e84db9b90cccf5bc30adf467d6114b
z6d18903438dfc9f04fd38b09c4faa3db21a05a8dfc4aecdf07d101f9fa9ce8cc63a8ba8b5b2efb
zef6d12f91dcb93f4c08d00c7e236a923b10f4cd799200f441fbddb05d57084164f197b600c0fa2
z45399b18823989bd0971c8ea0f235828d329c944bf1b23bac4a25d29172e56d3c2188ece9790f1
zbf99a79d4283b6d9879cd4a8b89ba099735cf7bc88bf1f87e596d84725165a84be59db8f0cdca6
z1dadedc31fc368da57868f42d55215e581da844acc9aa16544f1bbeae74e3c42b07e2da67ffab9
ze29e2f2734477d7b5121ab3baf638dca4b665a2dbb0abcaa801b6faa7036a5c9fe56199c7a1804
zf3b4e67be12a1b84cf5ecd320cb93ba7c3d26142d86173b5dca6c7da5dbec66ba4c80db1071bdc
zbc1fe19189cd8e112438d519c7d977d08631e1849b9a978fe0926bddcc4e4a84f61d3d2219f4ea
z931a350d52b9fe5c6dbe7b40232e7afc779f3011fa64de4568c0976f26277c1c522e3ecc500db5
z143b83ed8211c6ab03d3dc07600b142ab0589ebdcf6db022f43213ac1585a42b283333f72db390
z31988aa5ce6ab3cd25ce3f692eb6ff40fb5a79c1192522b1b32fab37cfd4f46902941c7a5f4f5e
ze9eb6c901afe994fef7c3faf7fb24ea34e0a22f14b829ae9f9cf7428f1f34ef70668a59a655f45
z43bf4d9aa198de538723a0244c2515b405a965d00896506954da2f8c7c29b97f4958ebbe47ccfb
z56f2c1dd235c83d50098ec6b50514ef8e6a76a0ef8a31e323cf00024ebffd3db55fac27c097613
zbe77e72bd7f27165253a6d3e57ed9300f00ad6ffa41276b0c145efd235f623c56e4d1ecaaa2122
z827cddb7a8070336780f3447662a0027aa42312572a3965b16568ccb8bb7ba076fcc988e33ae69
z0a134205c280ecb22ce7ef447ea849cbcb66b15479678e249a280c35bcab54a79584f4e601d436
za3639a78695597e0a079d2b5eaa0786d8ea21f0c50f495e96ff999ffed4de306efb2acfbd4a6ad
z193df657260e4c4c5b646eb489b5f3a9954ed83c05a13f82fcbecb775116fda5a387b25a16c13c
za4930e085be6589cb9b598749dff7bd0f0b274f738396ecda2c6328ae35e5c6f9fa8ccd2a8c935
z1800c667d8ea9925bd0cb461bffdbcdf673194dd8cfe415e4587fb7ded48db71bfcc4e3e45f924
z339ece52a4975ddb4a1350759c01510aba110b1eb2435eb76d887d6dca70e9d4041cb526c78d0c
z2f0567bb202bba4e0bb112509c76b853d2e20dba26ef6baac5b09ccb4c007d75def6baa2b6aded
z977ad02cc12ccc15dfa1c4799fc0f7634a05af9494232b20981d05a35588142454ca6b0045dd26
z64355425e39326b8461f39840b07a14dbfd542611f1d4fc4df948b271ede19700f541e74d2aff1
za1a049c5f6124a1ce7a9741c8b31d6d52fd5286b98b038687e43bfef09f0625c59034a3618a838
zc09977cbf68031dd480431d4ab8028469996188079c5f1313d18edf9bd0bb69ed98b2120a5a796
z68e64f6a0a2cc41cc9092a58079b0bd20d4083da1287f67904de248cb39d2689f00be9da146ead
z952ba3c0fed698b0e6918fd6ef8c14d9c8bbd3c13a392631a1b67bbcce6e9e6e51689a422305a2
z409d13eeadb9495c8ba84c0d5411e655c91fc6df0cac846949db9c4e77b930fba4f1b5f639e8b0
zcf3d7391c4909e7936725f0e8a8f0aeaaec162767e99ecf4f5e967e407c47ca1afc4c58edd3d12
z194b15de3165fc32d1b40d22d5ef59625d9c456d201767a508f69f032552598a8244a986b3cebb
zd32c45fee3d22cb440804827f54e298bba707f390cbf7effe6c1822a35abd0b012f0446e4fa6c2
z1bb9c3bf0f18fad878f444ad4a369809cfd46902add5adc462d0dab4e3f3b9fdb7fe7de3087317
zad0697f0159aca7c7022c9a98dc2a647acf9f29d51264f49965b34ce1e44e7ef2e73d695a57ed0
zf316d9bc66cf579cd5d2285a9d172ab0da97022f45a317e9be8d0a7a19ac3687c346808981c3c8
z3660c7bb196d810a9eaefab6357ac8dc6141e38445a7fbddfeeeeb863969c5c5f2c15aefb43e43
ze18a0f2f40b7a3924195de3b3c8463410bd941f960f36a8a9a3ed1162fad11ca8882e41137fe8a
z00e29613be308b29c2c6f0e1e048a9434ae1fe954a3f8b0d8ce3be3433477ad303f4844b68139a
zf48683cf0af975fe521eda9c3778e8d89fff90dce038b2c30afb29e190e0e8461f2e6d6decfad5
z2f7a2d8c54ff6211389aef0d447442582ce0fc95c31535bb64f3a1b05ee44b97c6a39e9003de55
z76b10822171cf03e4e4378be1636fc3b825ad4069861b5bd16b77cd8549e6227aded862ffb2141
zee93b7a6d3cd20b9d3bb2cae08b4cad35a3209f0dad1d3ff8d3e2c6b3c0585d15ebeacb3648fde
z5545a6b9c793a6c9239970c62647f74d8d76fb1d58c8675af127cdb03ce02f49fafef3fe350089
z9063cb84d9af364dc945f6ee174aa77dc7194f336c7c5a3653aafa3a8e3e5dbcd51c3fd8bb1be8
zebdafa9a713b7101725e27f236f0294f20431cb3f845e03e384184c66e9f97fb20737f4bae82ee
z856dd72d523e222497f2df53ef6c0086c0aa4351b282558ef1d77b3cb211792e292f4a0e2073e7
zaff9b60ff74d82d29e44540f35fe26544bd597dbc318b55fb027b81d723cf72dbb17e3acd497dc
zeb0f99c33b86b21c78e657d673c617429e52e8fd6d81705e336091e0e638cede61bac6ea5382d4
z4b69d6294064c4d57a1d594a6cc6bcbe5d7655dec4a5fbea00892a884836e8c43aefab432ff436
z41c953be59114f07bcb0e5832a702559ada851293ce8d9a97ff41d30f203888761236cbce353bc
ze879926ec2a06b610b5fed2898f196cf3e2884968467af1f3ecd3ac89ea1d9a66efab8dbcd4398
ze4d17c1310864b2bf957d95bdf7caf66cb495cadd88453eac352dce0591e8a41ce314aa55a5ffe
z6c8a457033e24b1f851c4c29bb8b2a46bbfb4c5aaecd9adafec55b296c8c894769d95f9634f46c
z72d4dfbacf873e0fa9994bee4668ade34c37d6243996fbd3eb32a5462beaac3035625d4acccb42
z009ebddef46ee88eaaab247345128535ccc044f24a0cf70179277164f3fd478b471164fb268850
zcb5d769e7dbebcf925d269f43d2429d43d536b1fed244b2ba600b618917dbee3c4ba8b25106076
zb84c44d3faa5fe1a19d803c16b8cae94fee68c0035c283c5131d9aeffe3c653578c8a4e6360277
zb92ec405041203229dc5483c4ed9830f889c2d3857a5536fffae8ce7406b88e7116cdbd88431fc
z56a8bcb3035e10594c9c5c318e6d360cf29b973a4542bbb0d7bec70eee78b95c232f23fc0df550
z86f355316e4db269f6f2854734d3e1032dfc4eed5ad3d568b42c47f643f85a99c74f26c35f945b
z3f176b05951c42385d161dec8a2511dc634332c1d528d463adc705df5b14c20fa49a13f3de60c5
z7153c3b5d38c2a02c435e7d8b888370a08211533966bdaf4b68e17d24b4a25327313a684d960be
z15fb35a6dffa099eded4a7dc645a31b4bb275a0529b4731b89cb30bb60db1fcba75c44c227957f
za48613366141d8db5dc1da8e1287ae79c4349915876d85e4a5d5930e03bea8d80bd527f2545445
zea6832710271679228bee69e571706f6c1764e21bfbfdc3908a5a311e56f523f16f155f874f4f4
zae854a199afac8ba720025a4d42b6857c56e0285efbb3142321fe7fa15e06b35d7f5a2edcdcd08
zecb7f4a668d79b01d0b6733226fc7db4889b1819aea1f13eb1039dad38d0e9e828dff600cdd314
za58aeb621153d729403058932dc97940a9e28a67acafd37989c24abeaef4dd38c9f17fe515f040
zc5ff589f3e662167b625c96d353704e132c4b54b0e85e6f3ba6194aa3e0722a2a0c854b6f647ca
z21fea8a4f939540a0063438a2bbec01fc3bbc02b3b0d44d45f4a9bd21650a4b58338b2bf90c97a
z65757fed13116a660d80ee57948c8817a685c41c89c11c2b3fe8eebd3c3179e35d863a9b3066dd
z4d9c60e15bf39420ee85ed13cf29360ecb9c8beb274c7a4cd32dac3b18fe35e61af6b02c13939a
z92150bfef8a41e9d40da1997b5d133b82110474b1b43f8272cf4ea69a99449f7b63c2acfc67eb4
zde3298d2c423702273c1558424ffd439fe582df47e43ebab2a3e3375378178bc659bdc8aeea32a
z99bee3910eee614bd1c096f513ba5740802fe0f0e314945c71a1e888da91078f3027dd36c632e4
zfde379c77632409ee0ae541ccbfc3795681ebab4fcdc481dadf35e73d9a0899af0235284faea8a
ze02de7018d6c0a666206eb53dd6e439b5a87351bc019d66521166de3afe2ada8dfe2729914c5f8
z6f94266761b1c7a462fdbe720fc6d0b2eadd4cefe787835b58de57ad2072f7886f5343fc42bb41
zedb6ee8eb92908b5612c8a72e5194f9e6c2359b17d40b85632c26d0b3a55402094dd35754901cb
z2e535e4ed61c289caef49a55bb594de449f9946892b116d4f28fd333db9e96534eca427dd481af
z547eb14afbdea97e257801328a97da72c695a3213487f13d675f4d9dc0a743947149e007cf7f80
zee7406de42e6b064a90ff94fe23f799c4c03a9f32df005eb68959ec76415d78f32b7d798bde4a7
za9aecd877d32aa093b87fe1fdd58c27191d970ad695892ebad52a8366338fc28c7df0cbe3f0ff1
z7ac0f030ee9aa473a8f32b2eb1ecbf770d967361babcaedd41f58c13f738c0deba990c225b5059
zddddb8ae20453449ad46f84891f103208c497d033c9e60c14116288616dc4ddad269716eece260
zdefaf7da1ca7a8815532f7f41e19478f41f25bfb33c41996e2cd1b403195220b3254ac282df395
z8c4110135b036deaee29f8c180df40b7beee979e21cd0eb4eb0dbf262ddb1510f0ac5e2951b4b7
z589947aba5767020f921926bd76d843c058203cdc56cb4edc86e340de2a7e3660fa7cecb8ebf37
z2c9f097db13d80248b8741945573002ab58b67a33371e61cd93ddfea5bb2fd11ea32e3f752a720
zccc99a75ac07c20200788a79c102bfc56c646f4557e0edc5fbe17e74e2ba79562c55b4509c7c9d
z158f04b0343e4a074dc969d29cd5693f0650cb9ce35da7f516372d6085b8af834692fcb658a5d7
z8f73aeb30a538990e6bed9f10685038fedc4c0137aef711c58053df4bdb5b556a4689a753f287c
z6aacdc46ba4e41afd1de55953cc780d103859b96b3aa362444aaceccc06e5b45ca7f2d7ab8870a
z7e98b0395d2dedb0d516ea25016129e6ca650552361dcdf9d646437c5bdb41cb1d54afa145946b
z57c176435274ba969becd44c3771357a5a9681cfe87d68e7588d937b589891ac7b30176e9014b1
z9307db001d706aac5076536c16ea6c91bb380da94cf6fc7e2cc03b5d5f9b605f682bde8226797c
z612dfcc8bf4440e92129ca7eb137b9c5dd3434fbfed9e66296fa320376eaebe2c7228c71c7fa1d
z2154959561c1763f2297fe7ac0b5c31b69f4f7b047ba87ed9bf7bb920bc3c9d4a785d7a7105114
z1d8174f71179a629caa8e524fe948ef1de7bf5d78e82a6fe7bb067443fc744e1edd33d44b05816
ze27574f065f604edf115f407c7a15fbd7f798bacbb060de884fb272bfd7ba6465d7c1b1c5fc55e
zd2e3d831c69cad7e57080fe218e95120e0862e47a475068f2e0f30b4924c2b3800aa72f0365bb1
zaa44cccba643d2dc1fd1334c799ba7dde23df5cf39ed3b8998ece780ed550f868e72061d6e9979
z716bc7ed30cd2fffe48cc05823d17b90a3708b0cbe2ec5bbe473be84bf0ff147f3c850064be13d
za9ed9009cb4374c26b1580a5d358db989e1786c6f0af5dbc1471a0201be5b92007515876c6ff98
z74a3f426ebaac757c092236f79b6d41be756cd45f8030a490e78ec7d33efceae067adbf168268c
z6b8fad94c035900d5ed0d00fe03953586f77da3816bd54a7bd1933def53a8067c2f56438d3cb71
z8ff68aad68601337ac976c9c046432c364e2f7d476bd2561359b10969f1c7b0ac7e85af172acb2
zb1456b18bc35990388eb7a7c88a66e47c31a1823eda5ebd13f499ee93ef63f0cd2cf5143ad35e0
ze4ac7adbdcce34218573320c8fc9a98ffe4ba22ea18ad4969204144eb2e93c17727cf02c341d89
z70c86d8677941b6f11f930fdadbe64c5e0f07ae68730fa6bddac3fcf86b193e1c138654ee04ddd
z6d1fc5b79b2f155c71f136f70ba0d99bb51b3da06bd183261df1a8369658a57f668f73b56f585f
z02ead203db15b5d1cf4e89b560657427ee8eff0aaf4e388373c434558920fe0a89e21240ce8423
zbc28d2b51bad1e144932ca43ef3e670bb6d03df90a73d94a71867955fa6a2dbfc3f8b72c932e90
zaf86f77af21dfc5d12b7ddb5fd37b5ea85881318e7290ed5cf46cef5bbf8ece93a6ba9d666c256
z68287006b66825493dd29dcee9d5a5510fe57a49ffecc626ceb138cfd64bee2e9a5b4838b784af
z254e9e2dc8fb2a943c8e62a8ea6f61ae115a73b6d08771e46077638e94ba2cf5ba9747c06b3950
zbc5a61cbd33012e998b732ca54de72ed123298f1702192bda2deb9c96f688a224db64794bf5604
z35999ef81da1a2d120949d0da637c6eab8fe734867f080694c45904a2dd2dd00888fc67ad9e836
za74b8dd7ed4a6e95f632087b7724da89398d49acef480cf04415951f7f4aec8d99ad98e64d4ef7
z2b0ffac9656f16f59eaf8e9572ca5eac29c0b587f5517f3776bfb2261cd85db1fff0b9e412a787
z6ee40f518f4249b1b014d3edd1a01e21b4bd5718aa4bf497d3d1e6f05df02151415fe6a8da39d4
z2255ec43a086075e7c0e5c6433ec2852c138fff4b8d220c904e1507452a00eec360d6fe018b150
zca38925c8f701c4c8a8646099e78c2b106b13b0814a3596d29597084940d06fcc98689b4315529
za997927b569d2067abc607339d0511456feab705c8ad7f22a600854b1fc069471276426404dbd3
zff93547f584629b28f19ad56fc4a414c1af04e721485a0b89dc60968ec33e2d05480de8acfa0e2
z0a7e993d16edd1a24ceb0d445674cd4e086195e050e75d0afe516de8d54e07397d192a2b9212aa
z5c39498ce124f6f5bee7f7a31a61f909f331cee0a70756b58b5115752e1fdbd5e013bfc85f5f9f
ze9db706331092f0187280d9d071c64135ed690ad766a8fcb237f269052f98df5e4bdd82ef33619
zca575d29bf516f5085cd9e74e04e45ccf2e506bfd6e98f62bbdea3d1582f48e76e6c9b4a2b1cec
z23c19a28fa1cf781b2b61672b88ae21ddd3eb7b347a03dbf829b2841265df6a28ecb4598ca9a23
za8fb31483f49e39c8b039438cc204c773222ca4d1d466b7eb98c4fe4f9eb49fb181ac19526663e
zeb1b122abff06a630ae79b20a9e3ce0a373370b9bc320cbb0ad397b371b7edee353f45b39d0718
z8c55b0ad2f9922e876f6e37a165841b5161587bd0e8d54af7531a5c8d23705d0d497031a5d721c
zf91772faf5fc0340ae33325572e1506ac46b793f600436c201ee671bed2dd931f932d19ff0c5ab
ze7436ce56346de6941fbf40088fc8a9cb339e58da166b5df193fe1bc7bbc9118f4dbe41265a406
zac811e55efd1a50fc451861306288f44e62c8deeb7443c297c83dd47e3b8b150701fcf27cbcc15
z61a4f7f520f138db6b6cc81d0efc1ee2c13eceb65d30ca35e60f16e755a47f2aa96d2b3f474e96
z34bdfe25e8323485d2b8cd55f031feec837e81cae1a70e5a8fec5471be4ddaec71cf4a98ecec0b
z3b03f51ce1974a637ca91d40b2f8578534d7a60791d7d58edd4f9027a6b93d7b4eb4f1a7b3661b
z68aa0575f0c1e3a8e2e2ddee0abf2436345e189bfaff05127c9c5e6050c3c4d2ec676269154187
zd27d49f5bc8545ca01c235dbb1e7eac0f1c770f992aee42220761b5aad74d4812f3ea5ad15459c
z3fc109b1b92abc6f870ce763a02771327905e2099bb02e5253358bb663bff03972dff2e4026da0
za72d1abd0b2157cd9ed46e80e484de0270e35aedbd369d15311f568490bf6e06f89a9010a3e68a
zc8a9cc506820bc16ace299b62da6323137e8217b8f2c46c9d74e77aacd395f4d4e820789a3040c
z902505cdc3a2dd16dab87cad1898d3a442ee2a68a1f6e075d9974711040580c28d620f235aaeaf
zed70036a3e8c6917473f9382fc8a160bc43e8eabef1951afd077b4d61c0c625a7583b307d6a77f
z2e0d599f47d6b0b14148fdba7e8933c8c42996e1827bbc6189c2528438bb2c494d85aa3d4d33f3
zdee30b30ab783896ba13d9aa6c3ab966308a79c9787835f7ecd0804c8bb4339bafb67fdac258ad
zc0b0940c5b7dcb14cb63e3cd30c79ce3eb42d0457719a50bc57a87f59f764649f461f9fc648905
z84df1990616222edb88f6a77e9c687ab69110f19fa994b3135178de89c29bac2b240040bd96d48
za3a4b855630866c96ffc1965b76d4728425e5b083676db65552e2c27ee2a87e5f8c992bf955511
z5783d52428d2f037c0fcce800bfdc1c7cc19ec3ed13a94256d349f2a0663e8602b490f21e467e3
z053a6c84bdbbd6cc0aefe5c67a0d9856cfe54f9eea7f7dc2197db775812b15c2403f1f864d743e
zd045da519f775fab2dd47b2e3eb205c5cfea552d3022c24e1f3b2fd977782f9dbea091a45dcbe2
zf345074a2fe96c64a0a73f32691ce522e59323ad4cbc0ba25fff2241566089e150cc4218bafced
zc7e44fab1675084a6fcbfb1af099bb3b98c88189abeddb160fff9b3f383c830ce3aed69e61a9e0
z5ee8d1ee0d7f381619efabff619b398e3740635131d16603df0f9243804ff36377a12a60f4c81f
z04241c5a30fd154b996554d8e3953766a8b1ce8c3a97a4bb306e585a2ebdbfc39320ccc53c7666
z194678db5dfd1b28f37b21feda1026165ef3806bd52b4a83dfe909557ee2a80965b5714417a33e
z2c7731f67b98ee63edfaf4d48c7681511f4456323b512599a1a48f8148f114e675548f3eb67e9d
zb3b8de2efea005aec4c8db1fa2408650a8842abcea72f4e7e895f03a814aa682617963ab859d3e
zce521e5f43666a1b65ac128b4ce3c32f822b35865d5886044d6896225bd416bfb7a1ff85e4fcbb
z18f84d0b3f38bcd6a0c326ff3173940986011a84b96c76fce72b3d8005596449bc5488fbc038d0
z32edc0a72f1889e85b39f5d2c7e7c5521dedd572f2362eccbc5d3317ed2997173bbb7b4992f555
zc2743f32fdbf6edf1f4a784a16461e994a7b24b55627f147b77b537f43fe7081fd26a43c44d9bf
z6e0eb578fce45d4775bb0ae9e2c6ba21f025617d19099c025678d0471fbbf3407764556dcac599
z419f8d6b79a168cb7c9e0909ba1138832fcdda9171c654bddc38dd2b2be3220948acf8d224a29c
zf8667d8b28f93164fd1efd41bdfb24670d1132da54239c26f3cac78a8435ebe08d49bc4ff2ed93
zaf1013c5d7ab4a8083da9d45bb8dd85f1e672f18f80667953e1ca72baf8c26dda9f20107868c74
z0aef5117f9fd2f614b2c47969f00f7c8f76c09317afbae4f2c2713c67c59fb6a599f91d3904f77
z322c1ddac15f48bd8417c693edcae181a85deb1ae6262758a785c870cf0d3ecd1dcc1b65639c99
za70e831641990f74d794a4e63f2358ad4fee164d45043b0bbbcf7851750ce170f912f3321a8574
z81c7bdf0e69dff85bb0f63462f15768d420c8a64cea7b027d39fd937a41f9a52b7a100086aa8a3
z6f470f28de3c82247125d33a49ad56a1ba058b5de37f33707747ac5ce045dbdfee1efb44db2775
zea65a2a6a8a23a27234555c5d9d638f1e48560793e9f6604b08d3de7b43bf3eb7b65b87abcfc83
zc6395b7988505f0d0e63584267d08aac68207fe95ec51f7a1faf077c3929bde9d99449326fd7d3
zd9021e3bc8f079a23340c4cc22961ec4e6ad12065093c67da283a28e4ff61dc328e7f46590342f
zd411105a65d4d30def863064eb7c4d164661331cb2b2ee93afe3810e304188ea763432234404e0
z00fa65e0d1a8c9beee0ef37a9f9656c270d1a09a28e00241da8a018db294f2baf6aea7d7778f1f
z8d66bc71764cf60b3daef5e801983c39f3ec89b3c800f3929e1099e484374d6dfa8e0ddf2077c5
z14e7f606140ba23c045a241da98118d910699bbe5b87ec7102c99559da2ae5903ec61eef28fca2
ze95a9e3959b46d690168526238d8073dd23fc39ef875b971f4bea3f6fb2ea2cc882cf4190ec7c0
z457066650bab6e93ee503e492cb2c57e6f944ee8f7c1ffd17b5992bbf212336a1d0124fedf9b24
zfc9baa71791b3dda44148717fe95c4f6023232570fee5c2ce61582151ead22bc34d0e5fea75207
z9ee84d532fe14e03e2e67e13c2e31065f5d99e609422399f2bac2338c29072b8768a796fe8cd83
zf9bad0364707ed3566a4c2098beb8bb2ca3564ff55b1d1ae158ac023026b187614ca5a1155c29c
zba10f55e97cbb1de80a1230b01d2120b366df1997f5f477d38e5a9f2b19f15a05a73a4d67d50cc
z542dd8dedc204c61c9e5a2e790e596862d9a8be61b36b0ea58f32f7867ff288cc929069e4a3b91
z5734ac1f32772bdb29fe01ef169f0a9580c61db92a3737ebc4b925d2c56ee1ff950f6fb40f776b
z2b4af7aa15dfa3b2a601fa40c1a02aa60b17ad96687ab79cc620e07e548882a96aac3243f6ca24
zb04ffba27d0686e3e01125217ad22f0dfb20f769b49ab57c1c0c3149d812d5281baa50eab70b2a
z41bf1914abdedb341a7e67a8e027671861d02d95c6076c61757483fa6ce96a9714c7c78b6691d2
z1a14cdbf2d2bc7df56b20856c63629257aa005114df7ca2c0fbfdcae2c00d200f2ebfc331fbc50
z8b5762a48d83d7b4f662e76e187e311b17216717c8b26340fe9c4cb517cf917ad61d6d9a484d8b
z83598b66438daaa788671d5df92afd8fd6efcf3f49f0fb53a7c28bae431b5b341e16e3196ea9c6
zac80e20e3a14dab43ebe60d72a5f98c409281010b6729625db6065091c63f53880c53d2bf93112
za3a3cbfadfc25ca558df1c271762a647bf225afe45bbc120ca438ac76e780b36a1229a3d8f0f62
z18ecadf54a0640e0f1bea460e334fe3f2c329e2fe0c498d4e59f65b116139eb8c2c7b79e05aae1
zf2318983f586e29730c2dced3a7eff8ee2d2dae4b3238da085e2b11a185d68d7ceffbb940b286a
z68719d264236b16c753725d57dde7d5257e9874e3606d0aceaf6ea8a8889c1b216cb7396e3c431
z307e69a22c380f14a49a94e249ea345b83526f8d36f85beeb72f883ed4164ec042e914976e6c28
z6aff5263d8693ee6a2e3698dd9a85c756be1fb516e12d17a60fe05a4ee142af0c727aa606d27b0
z0bdcfcc191318273e60bd5643bba42a697785b784431f49e7ed0be4aae8845afb1769fcd092b8a
z79d67be91e722a0b3ba40fe39dad14430d0fad4599b76acb36717af7df1eaedc4ecc4477c61760
zdaba957eb45637d6a89507e4cfaa125f28983cb647802ad4e5a94f4186005030c4bfb4c3dc9e07
z477dc5bb0d4afebf496cb4fd0904bf253c07c73ca5caeba0dc9008ed1bab3f7f08b7201ed77390
z79b0e6cec980bedc15402fb15b5153564297bc7c1777a528e9259deec83f27111f6b00e4097b51
ze69f1483374032c392886b89cc9b90d3c32d8d1af0654c465d9a52b421a83585e5dde1e4780c58
z51fbc2879bf2595e247ab9c178087418211f63f390c4e9b95f0d76ea80c560b6795759bac98a8d
z5aa80383828688b907ee731ed41dcc308c3b43be6b111edfb88cb33509adff100c77e2aa145575
z2ad424d6a0edab0fa2c2a50b352afcbeb64be36a87bb82ca2a401aae2991ab6185802cce228202
z6925c7ba2674380ba315ee16c6a5235a6c700f26ffea034123393b2adbb59384ddead8119cdfc8
z3461bb3f7d2cee0586db9119884bd0b805bf8972a577448e962072774188b986f095ce4107b74d
z369fec1cc8beb7c528ff49ec52d7aa90171fc3c8b54587e98b414d0ae7257d9e02bac9fd6dcd85
z8c2237208e9ea7aaeb382891e637167f8c6bb5e7d4f500ce2e118f254776c4a3cf039637be9ad8
zd6db3f0b8768ad10700cadee966eaefd993fa82515228df00e05719d5a0b5bf969d697336fbe41
z9dd628e73e7ff682efc0b65c88637504f1d07d512102373f65c2c2cce329fa8ba4f411cab5da80
za49dd2b89b32162f2918c0d14e6caf92588cbc74f32bcd13b8cef1a05ae9cdc138f5d39107cfe7
z8d7bce4a8ccbba5c5ebf0a036b1fd874794068e71f8b00d847147d8e30970e9e76c07f57098e68
za26fc5ee5c4394f48432002dff62aa643a52bf0ba8ed7c02b6764eee8a0d89f4c36068021c68d8
z9e7d8412f09e50f6de881ef8fc793d097b021ea0389737406f7381e39ffc6ce66798f294660db2
z179c7154c282712199c76f5cbed4a0adab02d888169f5ece82be06600a6da1cec94635f7045b7a
z2ea150fe9236baff954e1096307b2649b73d740c9da0a4c3ed644cc425b7888a44705234042a38
z9cce3381dc8674e199de4ea8bef3ba68a649e2831725ae10f90919e88245733b4e0c973c0ba97f
zf0774627d18f1b73ce497fdac978944c641116c340965e5a5c036831efd20a2e9d9014f51fc11c
z56fcc2c816af21bc96f4a3c67980e50e3bcab75ebdc292e764147776963f008829372c7e199ec5
zbe6215fcdcafaeac1ea92d1f2c5330eba58e9faa09c97d0c2efe01d28deae86137900e31d456ef
z3c8a74e919c8b6df9bbe62c1c33f5dd68fedb4444716c8114a76dc85f52058e28df48ba478c1c8
z27e548b071ec0bf426aa37d3be5e433db17a7b13b87d4f74861ed4f25bc58916fdfaeb9b55ecd4
z6ad47a32931dc6a0ce28eee8c85254034abd3eb75e4be6f836ca619df2bd1a5e74906074797fe0
ze30f257fd625eafceb5a8eb25ec040b7795e1f1b8940e640b96ef0eff88fd8cf2a9286ba717e6f
z8bf076954b9a4b049e9ff53b265a3e31f3eb4a006d90025935184976f61b19886de70f669c921e
zb164e83235189395991f82c772b0597ebc7ae273b5b37d42189e902e0272e844c7eefc17319545
za8e4f10b5dccd9a0e037bd4f34a2aef2545669363f7b628937bc1324f342d1fc165d6a4adaf2b1
z4b057d77c4a38cc720a968b1964e9341a31a5adb50d9dc3f78eb9efb6b33e121ca9e2a37133612
zfc2197dbdc1d0703e2396d7c1b9e99b9b13184baae9325044425fccc2b55346f3d616d73f16c08
z7376ed66d6dcabd2640925182241cfbdb27dda46fdfe6b9d83eacca0c39e8dc3929669c75f801c
zb4bc8ce8d71383ff13ae2e139373e911ea40254b17ec0a38fd510713a83775d3350760090cef8d
ze6ce044efaee4fb4506b381bcad3b352fe1f474646edcd8ac626e099c7f6c04d555f39db6a5f95
zde752cd36f24d68408cd15532c6d6653e5b942bd13a95c9b68bb54051659f1241632aca7382b81
z4b2137356d1b5834e878b206e6b15a0dac9ae05f6e9e742317501032e0f515184147f503e604c8
z0d463383d3b42ba5bba7031cf376d32b87d7e45ed9eadac5c5062c355174a88e1c86d10801c837
zbef499d73b9856b79ebd194d46161b9046289f40236c53de48f091ace34b3ccfdad1be2ea11b81
z4a3f893cd7f8322c96b43a613e7861928592ec9cc5e19a79a896621af113b0a4b6342db276a9e3
z42c267b94d0c9b02c2934f9aba4dfdc22634653f9e60267c85e7a5e00d03a60ce4382a771807a9
z0df966f89bd7627a983e45e8c7165faf486770f73babf795d43a9a4cec51649d343b042c0dd528
zb8b6cccf794f82cef26cc29f2fdb3d068756eb7658af5cc76cbcbc6d880d6435aca93a37a05b13
zc001f536cb070f173131219711182f552a14529b09b5c86652d4e89313b9398f53476756a7c127
zd11dbfec2e2941ca59a5a5f73a816132375a6e247f0d746c0ef6bc28368eb9d935d7b153e7dcaa
z2805630203ed6f437fec6cb62387e992dffc188816c6914ddcbb22763a7bb9b1cb45f0d8ec1200
z8b9debeb9205b1cc7bbed4db80c37a65050ccc54dc68acad7246ce1c745a467ba29de13600f6c1
zce3d3ef79a44cad8e6d1de7e9d0ea8842c2ef9f2cad29c6cca86970d2a3a90ca96b325a6d73fe2
z92b7764828c1fd6a30c1b330ce4eacd1845c43dc2c3e88700dc78735cd18413589dff4ce1c6bf1
zb1f0c43d0a6d7f31c3ec839c208108609c98e4ae58e0dc814e2de64b49f2bed862f02e0722d69d
zba695b33afa3d73a3803ebd65f0b409ed8c305b873f74f78d510c8d7f074bd1c707d7f09d05ea4
z5844fa9f2078e2b0eb1697cb40abab963bfc8a7656694fdcdb504c0c15244cca01897dd55818c4
zac052217b3e103d5c943c7976bfc9d4d483f871b7c93e4a00638519838401f4fe6e0cd718f5871
zbc5018b908dd17323aa55ea5ecff2983ca20aef9628be8f97d7d0d879e0ab3138de828a85c6596
za0f7dd5ad8e584d98d369ef4fd34a54c8a4485670dae5bfc7c5d98e1be61b025725db3e3ce0491
z6b81405c5608ab5be15e7586341ce3a4c33f6dc69785fefbb667dcd19eed1e024bf949fa79704a
z8847f9d2e4bd3d0fd76304b2685c021437384fd13b1bc159fab490709f840ff4ee81ab7d0bc10d
z8e978cecd233e84edb528fa5f5519a08d64eed23e869f59a18b79b96dcb7e3cd5a84c545057de5
ze21ee0102d15d61a391c1df676f5751a3f7438605a2c1ab0dd8edd5f5c061ca90df858c811ea9d
zc43e32f186eec5bc1c7b14f21524d1d524c99891808b63b7e4cf213218f772db34c88c0d688bca
z04882410dbeaaed19cb85c43026f5d43ce36fe531ad4c8047b1d0b98bd6a896ccfffabce111838
zffc2de19864fb3f429779e33e0d7a59ce9813b831e808536073797f5fe9b2fe01bb3c54b0384c9
zba82709137bae8bda766e8ec63cfcef91ca1538e0d8913049e79b6bdbbdcdc5e5b2087bf2c6da9
ze2bf02fc1058da9409e14000cc71bd37dd2be0041bed6f463b7bf25c8df35f7e2f665ae85b3b10
z17f16908718f84b387f581e77422950af0693b2006b8eb4b9d77c962a55d7cd08a8b03b1ee4121
z6146c00c45e002326cdf2f542936a1b5a06007bacad28f4e747ae3c39f8292a1a3c587f6409674
ze410c1a00630a1c66eb7562dfd36325942d158c7d9fd0856b108900536cbd7810a9bfc93a9c55a
zf2b7be38505acbc96f6dec9ae8de2d271df07f2f5c365ade477c983eccc5de0db7cfdca82f447d
z83b715463c79a2068f50665e6bd9adedf7c191a4be6dee1c86124c8cfc7accd2f7859f06fc80f9
za7fdf9e63cb8e3998a66afe0e4f3df049d099330f3b683127ae4d3e8f7ee61c26cf9ea017e9fa5
z7db5921bd1bfcc00bb868985e7e47a8c1bc14034f9f6d35e14812d715ff94d4b6f4d24d5b8c64f
z389b76b24d8b8a5c59c4d4e678d968f8230b60f91f232b80ec175725e00c1447b74a1f3c1c0664
z9147e93ee5d770ab05b080e5fbbaf3957daf926ee4c1d350f79e6bfdc9c38e5c9624e0f8d8a353
z33485e4ffb4d06f44f888d8db5255c94bb1845025b0d5ecd906a7a824d4b223e4588965ba20b9f
zc501df01975fb05ba8011f783f9bbbbb1f4bd049b64d657d7c38957e9e54f78f155aad4527a874
zeefdd3a6121cf24cd78cd43b77500058ac5bb4b034741edb47e5f2c56f15295cf99d9cbaedce0b
z98e83d21706223be551ef8ee4676fd78ef775560642471442e2a949ab73048cd7e6a4e8268bd73
z654057e0686f5aaf4e8eca423f292a693b40a738c7cd6e517f8e2d681361ca825d3f36fe1dd542
zb0c35b558df0def195a0644cfff6ce7ca546a8eeba63dd4868e8c0baec2c392ca18e4a9d1af879
zce1a0d8f796c0a581405cd80663ee95110b0b275a44fb8b031dc7ea4d71ef8528e67b4a1a71aec
zc208c580969976ef704bae823ff28d007575ad43326dbf9d2e3c648f169e1d2ccc6ac482a1b20a
z34193b0a163e41ee5d66bebb6480e758a6ee175ec02f54aa18e766edccc2aca176fb4e3999a815
z8c08e9953deaf270b398cb6fc07b20929115f6fe66c657285f97ad3b8901a5082670cb300407f1
z823bca09be0fe4a8a756ff6c9a390d5a73f3c8d814f052e8151d679986ce1907911a07078add82
zc0f7a505ed3d7671058169c567cb93b24de7ed9a44f707b6c05769ee3190efbc794a569adbc56e
z052cacdf7d05099e6eae75bcef2918948e66025ccfa607829fb4e025eb5beb01ebb1457b257f2d
ze2d4fad16196b9742d1f8937cb614ad486c20f8ed62cded0e183eaf4bf4429a0061eb6ee2ccf57
z072cfa918432fa86e4c7333aca0da90d80c6616702b0149bc9cbe555e8b1719e573f6d3c5dae42
zbf7146b5c8c15866cfbf5a1d6e46a2a0ca2b3920a3dcdb271756142f5cc56a2785f501eea57064
z77d36889dd3f6d424f2518401dae7c8883c40e14f41f7682a457eb4c49f31b87aa0aff9883ee37
z9a8704ebfd9d377e70baa380a7de4bb02986231dd10b8ac2225eda95ebd29993ff3068b8186365
ze560225c873b8e33283957992d46fab4170f4fa214d2a7799c8803ee9150c7ecdb1cf585dd3cd2
z1222bcf8c1571986000dd1b51ca5d1269dedbf8d4240ff77f1eb8af8dece904a214a815604e4dc
z5682f9a2607f52a74b7cbf676cfdef6a04b9583a8475b40ae8eb7004ff3662d09c5c76e925f069
z3f28582c6c5ff6f953f1fe3057c296519aebdc6bee9358bf3ba0e6eddd5aea2255077a32b69b50
zd04c7abd868d1a9dcbd021622d45af1d8bd83a3c76926687439f210c797ea64f4978810f27a173
z58df9cf3937ee916945bf2778947702a1a68635ca0e42b031dc2a3f349a207704a9a80de5e07ca
zd3813d7317a32344653f43e7ecc3cb62eef13d5e3851d17fa9d2a02d4062e45dd5105ba5d17d63
zee34804e66e5deddb1a8b404257887096665031caf833b5a6331188a315c3040816ed24ae9a2c0
z8c289097e1571cd22e89cbe440a9db1323f76887a202bd683783b10e212b878f1f044d5d340661
ze03f836af9d9961d0afa93f8fa2d23205522ff669ff36cfd9a99df706d2d56638b337982a05ed0
z16bd2cfcfdf9edbdb0e3c912289d7e98b23bd7f6358cfe6666e93832b940661fcdff8f405087e2
z66f356128f6ae83291d2cf026b0348f58fe5e8e3ff38e7be1e157fad6b190563161e835b59f2bc
z131c3a0e1f64a5b1057a7eea9f3547683381873246e79665b2fa8c70035383c35fd5b5314e1f71
z357d345bb4b7bd0f89e68208831cc2faa65259b4463ae494e996927330954865b2a9e09af13d72
za0393bcd62bfa697e4d116b47c71e38868b5378a069a3df50d759937f380063daafca3203a1024
z506a28e246d6fdf185cec0771470a548822e80e29218153298dcfcb880c927a4990959a6e1c10e
za5d2db8d31c413b4e79c932bad1bce1cb41376af176c0ac7bf89603d943f0526ca6bd59256462e
z73321a3dce381d6e1b268f4cfceaf04a9e7d0a46fe719623bb74fd3496b0f608bb8bf23e8434ec
zf966cd4761bb68b7d767eca8e48f71ca6d03b960f2d91dbe160b566b17c01c73ddc2a878ae1fe2
zddd8ce74aef16807f4be9449ee2bec8237991bdb003bcfd61cabc65c8e17fed622d9719da56030
zb73f7b979e094d670abfa7a78d24e99b0c30ddbf8a014dd40f54e63a25c3f562d0ac65b6339ff1
z5b4f26b9683cfd8a1241af5b2a74d610c28f4ff83bc125140a5bc8b0b2fbd3b5cbf5acbd19d9ef
z33f6a10d28211fbd70baaad6705f95a1dc82fe4412a706a3fdb302f80164fa9042afaa0f07df84
zf4e2f62cabaaa2215fb0f37557a0ae0e82a722d280b704a645df027192bfab74942c2f5deadec2
za1613a3ee858b976f8ca341537c2840ecb200c301b7a795fd931e3c766fe1dbe84a91c55349f96
za111158896177abce00a26fc095f667887ebd31cec513eb648a560883d263d6be18ea5d99902bf
z89a9202e89cc9c2d5e4df84d10e06605a9515aec6bec7b51990063155f91d686c781005e2a8088
zbb2bba24ec63abeb7198ee7426e09fa989f512888763b2c37335ba04edb08f51c0b44fcd4e3623
z4c87a97cd8717d9cbfbb4ac9100149931c18082c6c28d0149f55c301b85f705ac4c73b856c1bce
zb1e4542f4327a6eb18fe877b987d42e392f14c6a40ac09eacdabc030a4582929a87816190c02c8
z93c65a12c7693714c7671deb27348b31faa2ce509b9b48c5fd1ca8074ea4e1c3bd54e4b66fc5e8
zda1779788ebf2083c4bb6478149af99086b69ebacce666de560aad0e0cc1c73f235888ce4f748c
z5610e829813fd9fec0eeebb6c4d62ce73afd67e0fb9936fa787820f6ab9b753a5c5cc45088cdef
z60ef1dd106cc44042cd424a5134611b0cd4eaa43345815f0316ebede613080619edb5ae9d09061
zadc6f779280c64497bb05618eb3c68ae0be820fd3cb7cee0ae0c7576ef28aafe8feb00a84f78b8
ze0f6987e6bbea37497b9079f9764ea7a88bd82cfb176bad3a075ac265dca140f433a67f3888f1d
zc62bc0e664e057d1d58646471bd3efe916ab1ea09b17d62da5c12db24a7e44d93f4eb229da5d01
z23052dac2bc57c4e6c0496c4d9dd64f508cfb887cbd3e32e49c40ab640814f103cb5a7403d2871
zb0eb15ad81766ae98b8b9047ad80317e85b125c4aa083cda35e2d86628def6ba0b2602c7b2106c
z4e0812b74efbe5b8e850a80d94b7bacbc6796f1b4d5b3e3191cd815244bdedd7a715f2c8b53da4
z29420c15455e04a28b8e86aa78a281395f41c0b2f52bc565c7701b79ce580ab152c07cf0e41866
z2f98ae9bff3597d4c383fe7e70c1743a6d252672da3365e88e5dde5ac00379fdb6311eef752579
z1050be24956b62f920dbb2baacca243d36a6aaa0e3ebe8cb43545e19f9a0299db28bd039805b42
z542c0a426365b7702f85b90cda97ea189eef27075b83173fea11b55d35dce92967a16c63bcf9d2
z1cfe855a7427debb52ff16fb1fd196aeb7754654c9189e5f40079218d9d0a9e39f8176de521934
z172f3dac4ca73a50a339ac1ed8c5548ad6dc0428036d37e2b861315da43207c93da6609425fb8c
z5f8c8856aa7c039478ddb3b95a1f67c0a9212b6cc480f2fb3823e01ae22d76ca077f9bed4ecb48
zf36e463b8f3caa99a8946980a9eefa220779e3f43f4dd70fd34298e1773a7e9c973460725ca233
z9a0e3bd73a5b13b4dc23834a7cb6a16077b85d9e8901d52c32664cf18c80ff68b294bcd0e28109
z1506288356f130e9b6b98325bb0901916b4148cf73578f3b3ed6c2169cc033220a6b1c327ccd9b
z746a58db0b76104d0a7ba7eb669ab00eefcf2f7f73350bdc61502793ba718987483bfe13bfb640
ze318cc27f2cb735550cd7d46f4822b7dbe5eae2808321068fdf86c9e0547315b765df2472a5d46
z258c3bd885b8bfe38401c23676fe5bb9547fcff4d4ccaee7ec63a99f6b4945b4c9c805cf224837
z994337cdf8a874814c8891864395627eb3a0bf8485383212b987b682a25f29db8d64cbee1e6541
zedc4a05870ff9088ddcb517700b425619caa20708c318a85b9611b84ee6c3fe2ad485cc9825669
zc02c0e318f146c708ae09bd1cd31003080768883d9fab0e8c0b9ed90879329562a7e0088f87531
zf9014ccad663cbd7cf9634a02dd7c0e976c34d969efd3dcfa3e71fe47619622698369132970661
z6aa58dd2633b0178dc76f23185f0353fadc589b71b8c0b774bb35c07d6a765b9eb646367b41bfc
zfd40da1cd0880ec9373c242ee7c980b1b03feb8202c329689f1a31419fe5e51859ac0de63eda3c
z9b3f56ee3c79750830e9c9be4e241d9286cfca8b0cb20255f2319080363cff2066b721592c71b2
zd0202766a8a588b0d0e44b035db13c24e42f53392724f65bede087d627f9dc90d93fe6e8e47adc
z7ca5d4fa089c7fc47a5b1b6a5f3a6893cdf0e3715f8b932286bfc67adf179885831377c3492c1e
z377b5e0d0c74b9f60f7955e2bccb6b29fb41fd38fb47c39527a27fc3e5aa1e7466d0cf1e39733e
z654a360f8557bdb09f500f0b6d4ca3290c2cdf4f19e002d19657ce4bbb05c99257ec5dbd0b3565
z12ad0024dbe9763fbdd7bf976a1fd5329f363790174eecf9214a436a437cae536b612fb06eb161
z6ca6067772cd0966d42320d67c6ac7a9bc94880b95edebd9d8d16139b4d12c884c756d99ee037e
z006fc5ce4bbe3e600736c7fc3a3b4f218af2ec778eb87787ef4dc45d62ff13f19aab0a4e630706
z01032419e4db4a3a90bd8c462b56febbbc8dfbe7f8066a92e192283b85f28ae49069c4e482ab01
zac425a223d88ec746b46c1896048480f0907d41a6c2e381772d29ed349a42293f5669a074819ca
z266146d66321c3172b6cf3fe5278170a70c99d02d277a72ef32a5ccb6a4b614b7b4334500dab6d
zc7557f7b467aabbac2d82f72e8c5056cf177bf79053a3d49da5fae3d3765a924be9c2fb11d2dc7
z868a0c9f0cf1910ae8bc3dcd7be3ca5fd4902b1a1e2def7782c2ed15509385bf051f1d26f872ef
z51e0c6173dd5253d28449b1706fcfc4239ed7afb5e17fa4242973439aea556ed3c8c07017c75dd
z84067a248b65dfb73d99b74cd107e7019f0360cb6a6104c871d5aa0f4b504af437b5bff72d426d
za8e5909ec15b958f3f399a8b59aa9373305854436d02b1b361fd143f1857ab14756da69823f682
z1ef251e66725382c246efdf53420740d10ebc1c7cb3bc58da040599594c13eedf4dfbd8277ff79
z72437b052088798618c927073e4ad6365f56cf443519a3d424ae9e0aeabc86716702062a85ba00
zf3539932874ab144a607a7c62ace37a8db4e340af3de24fc41c969623c2e76ccd64b07ab132d17
z9405dc95fb43855e53b4240038f73910393d24305a8387de664b3aa960e58f6d50f15098eacd59
zab4957838661db69cf1b44d13dd92bc3fe448f951085a8c2cf2614679f7cd4b72cb4f03c1d1aab
zdfcd154cd8d8313016234d0eaaa8c10f453055fa7882cabcbd9b75fcd5192d8e06893bc83403d2
z99574739ac47655ddadf09abd0913dc66a78e70488289d982178058c7085fdf0db85a58146c018
z315272b86b01294046428f39b700e6bee648e78519219e1fadb39b9095580c4af5ecc7df1a77b1
zf2c5cd8c0d4671b1c61ae14a30f5166ea3aca3c493e474a8e1fe3e285d2780dfef54c5ca85111d
z5bb427deee3f929eb7887c43ecec6d54a3ceb4a990010552445f3deb06407eb2d54f2020851296
z0529399b8e703b8a7309b1fbf37bfb7fe265f6f56fe9461270ffd4a00a5380592751d3ffb2eefe
z16ef580581aa87e67a1cd3624ff08de91167449f9f946fdd03e62159d33e338106bebfe0a4f3d3
z2624593106526dc4878b7f525b47b60087222511e45dd9911ced1d130312675117caa38d2096f5
z39bf75a54c52cf062ea7cb23c83961639513876e45c6668c4d51dca40fe9b85dc2faa005c23823
z67ba7983958352bab5275b193829be2f4474da7d951fe978b7f8cb76d20d0f19e2ccf45b8f0ff6
zcc07b8038a34ece1e03e5bed3d3110c2491e827c54594ab192cc86255e8adfb1712ee7dfe6d554
z53519636cbae6ede3132b0c7d800968de5a2dda9d3de69b853588572f2c838875f3ec65914d137
z521c4970ac6cbbbfc74a1035e8453f8e8fb4313d86789f8b68ce2274ef390905559d1a34013fa6
z284c1fa9bf3001113ee7e1016f3053103a19bf98685216ff36cdbbaf3dd925d8c10f62e20ec310
zac43aa6e88b394de77b8902a248ac8be7d64fdd7582091b253154b8af8a3b62314f26b2023fe8f
zdd2a8d95119b95150132f4ef06eaafd0757aa30bf43fd8d8f88e915d18006cdec23498fa21a570
z4d301d5d40973227a431a634f37f91081d3ce756da188fa1f8ee292750769afe74940af1a9b5a1
z7d243216c224500c1b480a2351d0f11fc94a1ff0027eb70520b162f45b984a38c529e31d61fe5e
zefc0b726665cd59664a833c8c9468fc6154c148b299e59de5d23460f6a5a5395b8a3df6401fcaf
z53726e8aeacb255a2f3c6330d79c8ae8baf887dd11b85d9232ec25a93b453676d077867a3284a2
z61f62edfcec040e02acf25aabd7abbb6cb96ff0a26ceda5e3c4cd4a96cbed8c3efed1013491def
z5927b64953ca3ebd6deeef4a9ec5abb67b6e32e71b4ca9148141e91a6e31ceed0d3aee451625e0
z794485243ebd47d7e9637b272562d57c902c7f69144662cf698087e061a23fbcf6c242ff30b433
z7965d42ee42463bffc32dc57b2a70def28de59f982f375c3cb8a6d939014c22be582864e60cb46
ze4c6e732cc86154a66db74af63f4433cc99bb275e8e946d8415d43d74949bc858589456027ed67
zcb6d4a4b113fe7d85eac8ef8842f29e6489e35e67da491448babad9ed3fd32e78d054dfa39d6e7
zcc94ddcb326bb9abff67abe0bf6f7f5b0a855075550fe0d6277b3010e2244957f77350e8f93fb6
z106435f26113992281a9021baf958e944170ad9eaf177653d164d734ba8b66fe5ca33c9557fc84
z6bc6b06df37995c219df76d5b02a85997311f84dd872c2870a1bae4036f9a16b26790ac30e40d1
z38a05acdf9d3e2c251233a3a28e9e2a5adb18fda4bad8cc5416b51f5da5ba6c49d676e3602afee
z04be0fea97b78f13d275186f2241299258703ae1e611b2565e0dfa30b596beaf15685ca4a6a111
zb9719ce25df36dec17949c760edcf519bc98983f384f453787e1b92e428a58169c2dab215522e5
z95064435481cecb2c0dda373fa4bcd592020880f69d5d310a8218cc54fee36ab5d0c8a2d218997
z29de40344ec18862feaec5b9650a137d7bb8e05daa36cba98c59670e2ff950146dbdb5dbec93a1
zb6643041f1e6c99921642e7693e57361979150a93d5291c2ad7c5cd30a52f46a009afa3df68603
z56b26a420c6cdbb654973869ec0f1b652ae0bbdf2a3fb4595cb3429c08e1cac78ca340aeefbf01
z5db61807afec73958b1d138a5c6aa58988dea9ab4e77911f0609d20793bc7b72876ed7688d8857
z5ca4882cac58356d06b451fe4ba96632dc384a3e9855734845f6413b877d452291710fa97348bd
zbe456a44e0536bf37737fcb8204cfc70e3e4d0984bb5c0ab8320fc1544da85275278ada594c68d
z2a21e9b36a41a0d8514534512aa4bc7175e77ffdb595014bdcea7865335899fc985d30f9b139b9
z4d73bdebe0b832ec90d46cdaccc661d373e636e2d93a9b577c58dea57d88de1a7fc745699f1f2a
z1ef88d00ec250d6e9df3442acbaf6e41314e3b1ef141c42d2a6fbfa59542fcfcc86f1c752c746c
z12e5906bf323d6b578fc5857adc466e4a30591fd1a846a35d1aaf10d213f841fd3716f83c136db
zae929a38c0234c9dc28063f51e0021543a1f478d762dc55c337af3d054d7b50353686cf3a8d890
z31bd6533c842492ab899e11307edad64e77bd2e36169bd024ead7cf117dcd92b5befea56637d57
zdb013e69c14b6b2c773f5653a3f50949d1725094d802f4192d32fdc9a802f20cf35ca2f963ced2
ze1032200159f38e8333e6e802f4c47c0ba4b71bbf720ce36cdd5315ae2e1a37db2c5f6325ba1cd
z4211dc25daff320929459bc5f62a75c1aa9f62b20fa55fed5070510469ff93f42d1554960cf8c4
zbff7813d13e92e2d016e8fdc1e6bfcada7d2ff13fdc22f0a934d679633b42be7c7793972a0e99f
z537604a189bd7be196aa712b5ed89df42c755dd465e306eb741e898c7af91b12a3c5e351002b54
z5e29f9796a1c42a05f9a2dea272daf30ada74591454090c3f4aaa407c805ba93199806434bc70b
zaf49f7396d87b98bee746cee549eb6fc2426cc2e140c009542daf762bd24363a3430b6ef016084
z9848ce2eb66c6213ac498d74d42b615b6e09436a3d71925cc027fa59302b44457dbee38942c63f
zeee141627ee22361868cc2b3315eb3c4fc7d551dc48dd5ad0f4c1fbbf22cf49ded406db6304cfc
zbbf9c2794f7a061b27ced5b00e1919c765e5b055bdcf538183c46d145d73164c53e9b0894308f6
zc2bf9a4faef6590c6bc6240592ebeb144c7e2573bf7f5cb526bb2d47ebda703ed61e3b5b62cafd
zed9ca62e3151c26d6c8b43f53aa65874391e67daf9eb2d163a0d56be582bc9ffb9cb76a632e8a5
ze654dbe138905d7dc642b92252f9987f355d1a2398663e650c01a774f18b8ce99010c7c5f996a6
z6bd0df2b57ac25452a0c0b85a991ecc7a755f53b4936bc71ce98b6a5441cbb3d908154b8781ca3
z1f51e64c2c95022b7fbfa7768d5940c08db582c87b0165dfd3b0840d8a52aa029ec76cd0774cbe
z9bccbba2084ae32caf5155c7bedba84948fcc4b35cb8e08522d40d7ddf7422eebae8d0850ba541
za7b527a2ee55e1d0aeb068863bff0935a9016315ad12df91eda317bfb05abff4e575a056b74ecc
zb3cb7210f2aa36a5ba1bfbf434bdccc4635773d38c8a72819a05e36265a5a4471397a22f8aa8b7
z06ab930fd4546d83345106736bcabb141491d9a8dd3c6f202761e8125dc396d61af40745ce97f4
z26afac0f2079d449c422b42fc93bfee1f139ea8b5ca7e32d78d931987bd1260ad0c3f3ac2a8b84
za42f971d7200bd68e3efa6690d10964292135fdbb29513c91b732f4f48817210bd510cabea78ab
zc7787a7d599be9cce146dc76267a1608e86d06cd4e4b5197850f9d1aede0f62946e709f1d096ea
z0bb883e8d26063e5e814c249fb708cbd87fbf7e80e03f8e1e6cf974dec87e29e2ebdf24adc64cd
z5b13756c75f9143766da3f53c0d8986d26f7051746777eb7d3aa0c8d4bb157ec9b2d55315df574
z402622379e4f96b845b0664989e81b632d18f88a9bf22e515ea344df0022a0097f6d02963e7f4e
zcc655995f5032a05ef6d92ee846b5d21b85291d9af3e1916ac5cb5c29e8179de32939348c7ac67
z3bcf21652a5602e0c8ef6fad7c7eb5ee18c9ea500009521953840ed86fb5c90f1bebaa7de3d9a6
z56fbe9015ea67c4c3c1fe06dae01817357530f0225e6a1cd1a498628c88c520dfcf9590d3e9358
zb8030a27b5f78bd967c2c64ecc1473a6c8cdb8a976fca44fe5aebeeb1ac016f5978341fb0410f7
zf12496150254ec621ba7a6ddcd11d90ed27730993e08fa19c8d94948989477b130e4ef44c7178b
z0f6c1de75abd64f124154f5bdac5325228032a58945722476891ea1a2850177cef5d322d157ffb
zd50c479021f6350375c9314edc19af53a8707f0974d34864a1e82c0894768043f9380781473fb5
zefbb87bae612f84707ce3d71ba28b56961a5f355f1155e6289c7f060c7cae315fb0b07b461500f
zb854b758d50ca2de7d2ab7f387e1d3d576d2bde9daaa3dde6cbd853f7d486f6c3b1879366f594e
z69b9618dab8894e09d72369459a0e533efcfd625fc79c5e464d47780991a108fade71d834028df
z1b7924c8bd6a7cd0a77851552f96b9ac4a18804a50cb5423b569b802ae083e4a7821386f9afda5
ze5f4cb1723724c1196a26cc2ed5d3846d18a622dbc421ba42292b64c61e992f56ebdc5cebb56d6
zea77aaef297c023cfb6e93226d14320545e65ff4828c833b5143f14e64ca85b994fbcc0fd8d8f3
zed566d6c26459e9b56f1b729d293abafb847dcb6003ed994bf441d5ce9a1c91fa2b83464eb1507
z131a24e8023d4d673f6ce909e872ffddb8ddc96cb762296139d2ae261402f59be703f4d7fccfba
zeeb89afc3f7f27131f9effd31c72b2faf01873591161c41ba953d72cba9d1f0c349bac069f695a
z29ef62d5202094e269e0ecc88d147592f03aa2a58ea517924d94b38cd4e540bff1f01839b3c198
zff341e759e7ade4d0724ef7d1cb028b7d2658516e907efe3c5b250e767e5bab0bff37ce127ee9b
z60657f7b3dc219ee0394741c513282e35dc7f23533ce05c799e26d95404e8d89bbc09cc1c73f34
z485bb0d645a9bc0407c41e3de7fa5b967827fccb1d24fd9786c203fddc5392cb0aa92fb918b504
z081dd3af879a712e103edb530c3d1e908fb04391b80a4dc79dc0dd4767c942ba8444b43ad893da
z9179c220f45d73f4562844c35e4d87920dab52225934156fc487c6c34e6fc8cfc4ee8f6af29b6a
z6da16d493d5e9d2b2b69588d5dd455582857972567a763c620b76508e57b111e085cafa4ad1e42
z2efa4993f55f65ae4bea1317b6dd016a9cd848f64d0d258214f252543363c22d24db0ace7e4d7f
z66fabbd66bd085aa284872f3eba75fc1ffaa1d717b33861fa359abfc36913de5804c3f6b92bb6e
z736aa36bd4b495bae2131ca807904fce499a6b533361e9c7508ddc52d7d4eb4a9f53be20b8ecdd
ze768eb97066f8b35d552f1de71ee072ee74ef2f492541a59529ad08b7b517c88a9491ae981d9b4
zbc6da68d199bc934c56219d381e3d9cada3b6202938bd490729e08998d997825f7d5486b0c403c
z61e5df02ff62be702f7a1e022d0711c2082196b7c247d29eb3941d347ddc877ecf41012b3f0c22
ze78720930fe32944cb9ffc37acb73cef8d05afb3e3e088aa3496732b8bc3cba6d1e25ad056d9ce
z75ad3cdffcceb0fae9105cd16a145bfd4f5c88646d7dcf0d22484bcfbaaa29d1c0e48442bf3a53
ze898ff9b3d39e9f65f43841d5c665519822e89953d69a9d69ec190857f8ccb9f6b4d4ed210b359
z64e7b274e31c07ae47e24f0e1a199da9808e8d69eaf9bbbdcd990a508c7822f571ed3defbb4a58
zc57c97d88d019d33b3b67360b7ef40577269f70686f225de4572a8838ebbd0fdad2534257859fb
zeaf1a63f6d8bef1ac3ddfd9c32f7b43ed89b2192e6bf1ef14aad0b7ba81c2e6dda771a1516d52f
z13c360de2522695b1c61947085c56915134d4361fe56b93af1cc1f1f8f37a44fcedf6e4d21b926
za7d985f4db7faf9c01ec2468b3bfce3aeb06f5976d7a95f62c6f70d5bce741bc3570181f658c70
z6611e55c3a1c5b009f8d82599fd95266a6cd13299f2954b4af3d7860b37297fd6b50ae43d10704
z09ccb4c0479e49d06e57f47f705b77f2fd55031e67f407f7e966ffcd4c76b16c857b1298a0890d
za7c7e33811ba66fc23faf3128051929458c6af5fbbce614285bcc005f181bf2e2e2129f8543533
zb75f8485e7ffe0443bc584bfb23b5812774e9a80b0ca92e22588aaadb6d19c5077bdf4cc019fa0
z4df06addce358b10041d2a62270c422d847dd100df56c795df1d9d2bd19ae3d350f142baa4b5f9
z071f978549a09e5d942f8594642bd7c6ef8c3917988ff39b33baa9a43729dc3235269e602d6f47
zf9e7c3721decebb3d3eb5f895170dc0180670d5fd34534197e3e706a07f2b824c7c4f8d6a5abf7
zb779c8332315db5b3e5cb08df1bee5bd4e0cb3f8561347e1b3a86151312de8f8d9d80a7eb5de23
zcc90d868dc7fa87ca422cf015afc56060275e96d27341e9e639630aa88f0b634a9d19e40dc3faa
z9c43e9d1079fdf013d7bd0e77ef132f63d141200c2b2f01e909b2c1d233476b1194278e689a94d
z5057117f060f7885267df000f99e2f9895e711d39417f08f730a8ec19be7857d604dc3524afb46
z6305b2293b5409bc63e3d10fca8ef956b26ae28af06b4099aefd814df1ad61f904b57a99986b9d
z1ac67fbef17ae1665b1f29e47cf7d3043d4df5ec25785b770d742284743300d1e03ed7c144ed68
zd5d1d3a8ab833e9df70e3998001f23a45202057ecfd5124c0916706e8ba48112ff1e8b9348054b
z99d5c63430166f6358ac3eff69504de543e20f5ff934fdc031063656bb0558996fdb711e358e23
z86b63fe07bc32b49732ed729c3faadb591bca5bbfc30669852811d3a1a3ed50f82e7bb98ac96be
z630553e944c74ee542e484ff327234c4fbc0135372ea8e8dde500ceec53d7bee0d46cc915324c1
z04d2672167d22954ea89c3bba5b8b22b256f343303c8fd70fc4cac56f663f413fbdb810610dab9
z3b44f7a5df56a4b9f49c3c98785c955eea7f2e6f12fb2dd803c28268f2b6960e0e55254990056e
z0204dfc5317e4939dddbfc65329c78642da48ae091c3d618a96b0147a69227ff8bb027c503e077
z1fe5b396299e740fee077e9913d6e7358d68c2a867b50d712af93a67ce6c8825b1ef1a4eff1e7c
z3677db7b87a806739a4b9f9ec43903a6aac31cdf903c00bb4cf90fc483ba7b3d978d441ef2358d
z7e85c91e04e67141166e9c9266eb7c8e1223d49edeabfbb4d334615f24ea0e88149b1630e17135
z6c14cb8d5c769f87364390651fc444dc50b51389995c01bdf62abff30d7b6790a9842b6d870bb7
z224088cae97c3543977c35f0f30ce68544e35e1210d1b851f3bbe4277f1817dd6213828457c28c
z63d48f766a9e991deb93238044b84cf38fc5ea75c655cda3e11ff4331bcfa17f59747b360db0c8
zb578b336e577f6e467dbc67a4351ea63963f1f85cb1d61a4f0389318e816f3d1dc8c89d0469099
zff6fbe523e68d8f2791070a8bf6b34bad127661c30dd1d95aa707ec06fd7142f55823beb3d4fc5
zecaf8cdbe8b7146011fbade486d623ffb07ade74e640b5a74750d8fb4892dca80f5f1efeb610e5
zae6f65fa0e1b6ea8490d967b7cfcbb0ae6f3e7568785db212b9ed2e061fd03d9126102c80631f0
z8f43dd35156f38aca92afaf6224001318e6f529ac0d2a11c07023f14b13c07ec0ee9360eb76837
zcabb06f03421481e9b5ed86b8b976f9f8cec8e045a333c8b4c4d3e2f8dba552b9e541c4aaa7130
zd7d6a60e23c0f3daa0a7aaaaea2cec86864dfa7e79f9896402f5000bf69c5657379a943db18a6d
z4b8da821b193fd441bd2d76187aec7db1a047e9dc19cc2c68db2bb926f4c39816da96dd56b7944
z7b07d713828428b3a0964c15d2b00ea14dd1b0d110553784eaae6879c48402cdc19737c9ab1073
zab003fc732870628aa28493ed8c96eb773928f1d1e5c8cdd5443966a6199a5d1cd4ecbf0352ecb
z22eddebd1d9957917edaf9041171aa17dccfd2c22149c4e07c9ba475635ffd41b38b0f6e50ae2c
zf2bc66fb956277ea96a3ac89f930d1736d3edbb9384b920225138ee12bf42630d4e2e075a50f2d
z1380d98e6b629a45614eba75bada6ae1f5d529a59832a16290effa2ee50c04486826cb3f4f9402
zf422dfe279e659c14e6a9d557d3cee0bf524b68e61250fcfb1900d7ae7bfcb836aa948356c40a7
zf74c750591c3f8ed5ec0f94530b5c8aa1ca0b31dbd4c3730748ca401c8fec18ed12e0708342106
zd09b77f5ef0240a421098fdc5213729025a5bfec53eeafb67efdb0a0754b0469354d52bbc381a9
zc02d023d43b8cd609277a753f90badc327c663e8f085e6cf009614dda0bdaaf8124f0e34764144
z2e00e23e49ae59fcf11673651b37ec8cb1847ed7812b082642c0667c4c1e8f5dd81fe80f1b89ae
zd969e81294ebd595060f8781ddbde4f4f83a9c576216304f71ad8090208f752e9042a697f232e1
zdca86264963abd82bd94df330101806374af5c6fed7a180a7268f10a31d19be4689fe5aaffedc1
za07c2c57bdc40ac4a8d249d63f997367408eb744df6739ab1e5cf1f4c6c725476cbb238b34e2bc
ze2506f15755f54dcef01f2fafd26611a01ed97ecbbc9c1b61ba688c510d6a84a5354542ea992e9
z814d17529887e8426e29ae82791365968e880049d8c26da2c6e89e9abedcf2a8125c4a99eab2a9
za4ec2139882fef11e4f078b298bf1ce6772b058738ca9b7b4506cac0d0c5b8c9b18b5d89362d15
z99a98520aeec025124f135d3a0673f60752e7099891e84341fc886e92562db7832594125eb05b5
zf203907c42f4c25c7167c7399389184c3a8a42f7b133854a8eb44307d40f953967b0501592bfb6
zd07b6ee644ccb3df7966bcb86c17c2fe06c74f8a39c1155a6da01e27a51042316f40aaebcf3571
zaa91234dd113388bc708c76ea9d51fd3ee6c826575db28ee30226859e80310e951e7610b443a78
z0b07d79fb21003001b8d38f21e7a1dced5cce88abbf38f22b0a1ef746168239d77a07be07899aa
z9f3cc239f8ecbad2f3e0afdb82605fcfc58daf79cd16e90821e6f1323aade02c41ece55e7cb7a3
zbf5c1d0e73dcdd109f9c6525c1be4fbba1375c099e47209a20f3c08e519e798c0b3c0ffd74d517
z71e1e7deae364a3f3d536f9002ca75f228934b7beaee4f950408168ed792c870e3bbfebd241dfe
zc7a4cdc64c532d5e7c0db531874d95609dd878c5087fd46d36cddb110041ee1b81adeed03643dd
z37f3d3e704dd9a99472d13b87c276539def138ebb3bb035563a1d90ed9dcefba4c373a319d2875
z4b569e75fec0e3bcce863a051065bc461d850a456fa62d6c1d7b24333f8f3c0ae43759317b7c2e
z397d5d23df79d8bb1fd8d9afc3f5bb69147efaa467dc42379933aa1712bbc9349ec631218a88a9
z2b3cb751dcb61d0d0dfc3d4b4b64315ab5db5d832ff39a7b26198e5572386f1c7fa91797c8c9a0
z028fdeed2a86baade737023712aadbd40bed83b5b191f4bf1935fde40b7eb0086c42ea9c7287ce
z3dbaf544a3f91f9f63dad35ce46d50a03915a9c002e8290989bd0bcaa9ce63e4055c3e646d6dd3
ze97c93442bc06e4d3e632737cc8464bd25cd7e9ef8833d0fbf4dfe51f0b860a8416e9985941503
z1bb93798445957d8a8002475650e78f04fee310b01dccaf5ef85f742bc9ed4ae7389fe70390a69
z8abca77633a23ca0feb1d07412141f36394cdca385d614e0809b4e3bc2217a8c610d5384d8e8eb
zb0e6f0020911a30ef2a2955db81289314e11fa56f75b7ee770df6475cbba539a142913b68c81e5
z22a5a79c79c7b5a6a5669280065a6cf37a9cc410d9924e0c3fb4358d8e1365f4690a707698cf23
z111cdd85e3b05237a2946dfd6b8bc63d0dbdc5564a315003c762c8f6b8e3faf6d1c50d6f24044d
zba58752b8d7d54097112f6260af75a5b0ce7aa551b9576122e329f87b4688b6867a9914203135b
zc81701bcbe806623afa88a07dfe1048b3a2d0a10df6f6ebff9ab61989e1504322a7a7d08ea0008
zd9b285828f3124d660f990a654e5345714381ac36004729a2b3e41984913e6a15819d857ca0442
z759ac9d2c47d3764751a5d667878de219ecaa29ae23129f46f940b2ce7118f6464563c8e4f947e
z76108c3da061d13819931a05304510e4650e8b13de6723f52670ce02692ed1461793d37d84b607
z7940b5c908f88f03869b6a32d63b7ec13e9b0e04a16b75b652f1a27710c727f57da3e4a55daaac
zea5620532f8a32505113fb88709850b09ae34579a7e4050b51deb7f5834a65e89808cf170a454b
z21e888073485cb707737d8e5894114ca5f0fa3f75516cbc5b5d50dc8e5e436558813a30c43e3ff
z4453135662cf07012b44edd04d22497a03cd13ebf0cad8b70dc11e1f7894cd8da21507845c8699
zdb6e932154b4ad0266179e374a8f99a440ac24fa15bfeb2681de30ceefe62a4e0fd20d18d17e9b
za12f908be0101f2fd55f739ec0931fbbc7c76b175fe411c4b2fbf6e0c7d4ba07692aa1cb2c0ae1
z8aa33e995789ad5c3cb29e0ff77a36ad087ad7e5c5202ce660bb797b7a005f8a42d6aa13e48136
ze17e7513fe6110ef3322ebe3fce3e6dd1433ef4dd75cd8de1005ba4b2b407ffa869f9b1826dfaf
zaed650a3381b5c376e7aaa59e4c2baaf6647fa6c5b8bde16ae89f0ac692d50441dd3e08b990a41
zfa1fe3cdf2a880e357cbeb1c0c6ad99b7f67d60216f91a478d1b0fab5abe6f35a889532272eab3
z9679a4798bcbdb52129d3467e9c002dc6e7bd52d82b2fb431b9fb373d1f909eb4078056b942d40
zf3914e59fd2ffb79d3cba2e8fb3139c7fa8f626a34ea073689063b39756c9b043da7c70656e4d3
z1e28f6244648a477a9cf422aeb4720c782787831502c285b67b45f2a82f2f871c357d2a56c5171
ze316efb555108c6ddf30ef333e750a8c16d22f209ecd781ff8ac23297fd1f1eb9761c5d04e8430
z8b47fd25421012d51360ac966df2e48fabd991ba69841d3be046fa458658d3d6e15c3270b2a723
z0a9531e8f8ea624d7c7c2cc2da826a860699bc5edbd5d07b8704ae81737f5f946dd8409f77e2f2
z2b79930f2cce71635064fd08ded1fdd59f21adc68c5cf5152bce0d793e5b2f03f530dee4aa1f7e
zd73b9da5d9447d635eb425a27769002899a128173cc335c636290b6f001d0964b4585c8e58d5f8
z6f40a7b93bb35440c6dffa78e16b747910f19f764d56ba6deb98050197167f43ef98e08650b02d
z112a9d55488e1a5b0ea5aa9c8a0f39a22c949f99ab61e39d4d64714fcddb39d23030ec840f3877
z4b6c2d5edfbf65cc5f38cae6344dd7747c38665096500924e4f0ba03b2903b9dc374d193f27899
zecea4c32cf3d3980c51f3bbd367c7d10a5d3bd22dcba082e22bb00a53b06d4a57cea3f405b1926
z2b3161bb361b9afd04d0e3832dfbf5b8055ac2569567c5990f1300a50daf0f27a1216197b27824
z7d0462c64af8db29f2e3e527d36bbf754254ebb46fc43984268234d2df5947f276d2693e84937d
ze291ab41d2c537a3db41b895747f42797aa5cd6833c519d1a57b61ff5368967844abbd9fdc8407
z77d4a3284036c293a34906e5688f8743a20400170bd162ec50e2fd1197c04db256a5ae2eb848b3
zcaee65e15ccf4e622fa808d0ad9b910ca90fb3cfad07ec93826ece014da5ba55ba76e89439bcdc
zc3007911cd7a0a229580f38545ade4a2952530c52944309b2e1490f7309aa786d331ecce25d349
zf3b02190bfacaf66f8143ad4f424a490f2b08a11fe2c5b526ebdb0b76ca6908fc4c5985b6f2b37
zc2e511e6df4ec54ae1bcac81844047822a1f9cd8e59d40163a8c2ae98c478382069482baf946e6
z88e0d8e20deb2c812be56c22d54e25793df4af150599ee6e3932647c9bfa96f54820cf540f6245
zde2a9c73120563d9de7c60ed0751077a17860d1347b98c507721fa4ecb1f6f48bb4840a562329d
zc075915e26eba77fa950318b9f62c71766506357cdd4dc3ca45d2c39a150303ff559b76c3f44bc
z3e4e155a087ea4447cb301d0e4ed78f54e3cfa0cf1a9a1fce2e57693dfaba5b792c7a0c5879dfb
zfbf0dedb0d2ca8eeb2ad87791f15da106a96ebd4eee1a0b20d01a8c8f28e71f11080ccf0e63852
z73f8b6b36a3ea2f0d959594c9a7b6050ed65066137620391440b0dded069e525d5c8aba5355246
zbcb6ae98d428509a9f568632bd882000d27deee9f439b8c82decda3d80d76c5be5e017bae91078
zc19f106313f2cf4cc1860d68479be9ee1b0a23b9e5e505c61da07719a0d30f5f69d88e1ff70b82
z8d6972d6408781bb2708976f61017585d63fbc89fae0a1260bd3825ce8630c15f4ddcd2a7a01ad
zd2967061ce9a1597dd41fb09a72c8782d3fa26b1880cc5b70d660a60b5fe74a2904edb173aff72
z3133c5c4ac551ef8d94ff2bf607a722cad4a40444bc4e2246cb83d6bd03937a19613e38be6f4b8
zbbae7f32ae34760d76ee38ad6b0988b33a43e9ea60120e77d70c108ba4f07e2a3da886a3aed66d
zaee1267523d05f9cf6ebf7d204e847c15524a725d3de96c5044d7b0e0506764fec29ce6e7faf9a
z3a0f7158b412dd23cdc2268ae6ade152f1be0389cbb4a7644ed69d074499343e162d1db28fa2b0
za634eb002ede48a150516c8e2cb195b06ea8769e537db4617d6cc8966f14683dce8433630562ed
z0add0b660fd314accc88bef514666d84c16a5df118da56b6367349e48a8148e72edf78b0e72d88
ze119e4f4c3cf23123aedbed50c09c2cb26cc718713235c2ccec0d7caacc13e44be79c898c96948
zf96381e181ab2c0383df93067ba4b5dc0e559335c4a172dda7243dea092a157548044f2cc521ed
ze7b454df40d1e072489e2d1d37f7b29aac2d45a1abaaaf9d74fee201e9320a5ca0d60ff19754d5
ze8bb2f604a49225f00331f23bd001b6f944b810cf5a511dca5e1ee7d5a7e3066a46c5aee825a59
z6c65cc18efa9552413a57b2de96fb004a5afcecbc95eadb26281c2405f6c68898b675fbdffd849
z1da6885dc5dfcca23a61e516163a1e1c38c3c3ef8c11f5288c4763795edf83b9cbc843b5c932fb
z479b3b6956f803f181acdff42de2f231dad94328f468c0b32e621074ce0505f5ab3fb895e76ff6
z20f2102393911f01d5581453ad5832f76174e3faec9107db197fa131bf09f2c86310b325ae7b0a
zdf2a806473ab516980b92018173d0bb4a01a6649f2f31c212785c0e005b559712673f0064d4f7d
z91dcbe07f99b67470788de284d7f267a10a65a663241b6af879c4c4e29ebf87dae7af74c830acc
z1539d641709a02e26a1c9490872199515dcdff7ed58e6ca4d50498fe1046e9af852d62c215ec02
zc82b82c781423778350617ff956d4b1729dc0ceffe9d25495376321239855ab9755e607e3ed15b
zc541e7fcdc7d2a3aaea4be6bbf758af90fe52634bce729bb3d09540dd429e15d22a85f4a3755fd
zbea7341f95e11d5bd4e2476f9a0e203e2ff186737942354f06fb5e82d3ff57f1d0642bef979b3d
z6106569d87ee1e3cbd0fae12bfb24dc790a0a2f5cc048e9600c96677dedc9d9c979e7195d23279
zf7585c7add82aa82318eb2391bd17d13b69773a84865c94b25c08f873ce1b4a905133c5b0caaac
zfaa3fb5cdf68ef296463f67c9ce034f8e4bb493134348c5219cfdb8e3effacd3f9ccfd9415d8de
z24ad374e5065364ebf4eeb7d040c6e1dd4c8dedc66f273d4a866698636dd59ff40de14a2728dc2
zbe229a61c0950089eba01b10aa303b26f67e06b4bc70cc1bea31c48b30d124f998b894d5635bff
zb442c649a1ed45a8bdc8647043a19cc659d546a1cc76ce6ccf50761678eac61dd5e8e38be37fd6
z283bd4551e59df5f9d78a28dc488cfa7e61e58b81125e9f27e905dd83c1795187a412dfbdc26c5
z3329c742b6240b9ae2932347610aae662ab3af7a1990dfd47994fa24f7a9fa68833862c9290463
zabde717536f62c3aa3c0a89d0c5374df36887487d2dbaab2e9142e8b53cb6f3c63e8a8068ab7b8
zd33bbbe236dc3975268448f260834a95008746dfdd15720ee2a9e4982ebe0a815efd1478f81f74
z58c85a5882d04f4072651d298ce35a6aa027b3942f25dfc88984ed231b8fb945a80103d81e5cdc
zfcef4cb193b10255c08f5a9591c5eae1ed3518cb95f2c0d4e7c64f05bb3e8f50a652c79c059f14
zfed8e36aafab1f063fea8e5ee6a1d1a39d0846fcee858bc6b89b30e4f85154d13d9115e8a58c98
zb182cdf7cc5c318b67cf3d2152b2cd7e67b3ac899ce479b68f6676449e26e69aff6fd2a1d4fc3d
zba0a6583ba86ee3e6c2bda90a94eac524e68fe2d541502e87207d7d3c19b6965eb320dd1f43a57
z1f683179a98b31dae6c91d7d9e1bc9985794b01dd5959fc632210ed7f27d858c2e2fc6f6875a0d
zdb27e414585ff73bc1a053603b38f16e8604e9e0e185fcfe5965de50332c26292f2bef47acf72e
zf68cbe6c5b8f7b21d0c159e60cf2a0ab65485f6f5550b3b45f036501ddfec65d5dbb524d10d531
z2e9c5ff117a6b250e61f73e05fe8927177158793012cca6004ead5a4eabe9548e10f2ec2d7f821
z8a5b6b109d810a02615f093df8e8020570a97be710494e50db070c382f40d58bbc5b0820ba9568
z53d8843f3ac1c372f9b1c4a6f1e595e733a988be6117829b55dd45f2594cb590dd36bcde8d9900
zb1e1081bcd3ed33d66d03153b800c9626a6873eab908e77fd9a15ee3329b779786757772cba698
z3f188ebbdf30bb02171747988c113acd53fd9ac0398de436856bdd77c96012d54a1f2f75ec6f8d
ze50e5e5ba0f802ae774cfa7a39ed8680d09469c53dc959c9fdc479da0fa5bcd265bbcc8997c7a0
z2c7ac46af9ebaceb4ccf1616cbc37ebb299ed7f68d5b1014b4d14a12d757f82b2d346f3b53cafd
za9d8b73d8e019bf1422a8cfcd6ec64a34318eb0410ea8459e4d6a2e03d9a0dc5c17260c5625138
z4b85ff90dc84831dd447142e97fff6ed8b429fcdb6306dd02cbea1ba02263048dca37155ef6fb4
z640ed4247235f09bed850d1401c069f48c35519111e0d0504c3873345aedd9d084613cde09e69b
z8be3e86d1f217794fcd8c13905366926dd80db43caec3c2489079aea80eee70b2f34c5085b1681
z1e6d14455330ece8800d88fc9a6af21c088a57aaca3a8d95c013892b7cfaf2db99eba6ef2136fe
z68989d3262fc59940506adae0e20c046d00e3e4b6e5c3900fe6f19077de3b2a92f0b67594f84c3
z2fe38328626df47edaf63c9f9bd72909fd9393d972103843c3298e34ce1cf3eeb6b06e4627bfd5
zcd2afcc0cb737923ce0e9d6f9ed3b4571e8598d8d4aeecefe77561087fa8ae2d83c8193efafab1
zceaba031994579c51797fe57091febc614a569535843fcc9f8341dd85586276035399173cc27d7
z38f2147f524c7141567577a5da05247ec4885de297d94da94508301756471c4350d1c486a89296
zc6176858a1ccea05ac9830eba78f06b53698b619ec6a107139b5083f81450b12f0695ded01b45f
z0436fac5f08de562be700f880d348fd87cfe7c33e7086c7bdf58d5d3a375ae3682dbe937a655ef
zfa23bc325d54d1b6eeabb106bf04fff8d7f59c4c2429bf1f25ac0ef42490d6dddb8cfa7768ffa7
z39e035806f45ed03ac3252f877eb888734af3e488e104c666909d8c57661f2a015e35ec7f9cfb7
zc018435caa001b0a96bae6ca9df88b280268637795dd8058ea1b4e61295384367a67574c29dcd6
z64760b3cc99f05ec184493f8c3dd0d914a6b50d1cc0cc4adc5fc92cb4646f057663f7a98cc9f5d
z449cee0b478047ef03254ce2fca4e92434e06570a8546f0b9d3a3ac6db82a33796da97ec8cef1e
za4808c6e52008e162ec7fae89f72fc3b2c6c1773aa9d06ff04b1cd65043c32394a91b6757c9d32
z9b34b20611ab1a9914671694b500e70293830ac2c18b7a701a0d96d93136871c35542f00f34b10
z731c74acf92415149800b8d836cff34e6da51f8c4da55a195da08db185f1ff93b748c1263e77b2
z747f6d240ba964dcacf2b3390246e9de08324f74405b24e477bc1e13e78397fb7ee6054467e4cc
z677fa4f17fb9859a258b961a6de7c8fb09005f64f687ed9de66fb30106964bcf1c9361d8c267f4
z5c95da985fffc771664c28b65d5b1aa32d218b55fec543da573a3c3092b8b3d8c123a752dad335
zb8c8af54df718620fca4528efa5497c8710d5df514449dcead1240fa57e83977902a0371ec2a64
zf99eaa4b1c233fa3cd0e9667579f8eb03ce7edc5481a52d333b5d374e78767c30f8093cf290700
z36f414b9a854827004fda7c2f8d3b8c37f0701444597429b01269dfb29633fcdc0ef903bc9ee43
z0b8f07f70c90cb14a480974f7c5bd199c74e1bf3e4ae069046e9b53ae4dcf7b5851682c6ff82d6
z6d20531c732489e984abaea5220f57d743f41b15d89a3eb70a6bfffde7e045585e98ede41e3d4d
z393bd51b7287b0b6854f90d39fb5562cab3d14cee1bbadafd8748581b26e4799cc25d8816fab4e
zf471678ca1652e4fde1c64061bd4cde6ea1f9901eca2e3dc1c5f129087dd65d19f4eba26919ba2
z0a40f970ccb9d4329ffad902f22c885881ed10ecefab7781872a7eabe641bf93e557c2085c37cf
z24d189278eff026fb1557b5a0236f334f270b6be66fac6960d3d39ab81bf646d758dd41311a8e8
z85253921353fd11d6d3c0212ed4256f0d1678e758a50be946d135b6b995c3769f30fc332663bf8
z9a13648ed49fd7f79ed520e5672517af5b3bb6b586c5200e0763475198b2a732eb911581287ecf
z4cb8ca852708c817d4dfc66a1a8ef64c4c80f48f82131a20b4b0e418e79eebe326139e66cc22dd
z2adba5ec04042ee3749cbb678c97ccf5210a4fc737db9791cc11a0d71557b5928fe4f5689e924d
z8e5f947573a84aea8cef6092b880bb64a7ba6fb75c3c55f4741148d5e0a5130164e89ed70eceb0
zce2e208ff9723c6a5aeed2dc8991370e5ceac6d31677075a35f1e8917926e083e5f6b8eda02936
zeec0033821a0c7ebbc51ca9781a5235bbd741ddbfadcb8cd58a7b07a7f89cd55031fc00da39066
z0494d362c26c00cd373c20b39e842582da4b6a9ea04fd704863b7516e218eb998cf5054b47ff43
z55cbeb7da7f46c8791b9f8cbfe1293f8e319cc6901e42b7fd5c3c199d97c25d19f75fc7c1b443f
z24b4fe895766d831c693d910cbba581f835c1743487cf8b0e13ef0673c22a3a239a20f09d900b3
zde6824e485821cbc051febaa2aeca41e70d170744adc79331f0d8434f5acf90ab819ae2ddd6d4c
z4fb7f2ca57a76f8df5b9582b7ac9e55f87638d026dade40e19e622aeb02aad9605fce3d75dbd56
z4c24157c2bea2a44009d300ef60a7d19de0c1ed2021ed638051e844345a10d767f660f983b8abd
z78c8a50f59f961489fe7b1e8dd89fe8e0baae9afdddae141b06294f3943517c93e2a228b2a657f
z5193b262c3c844d47fb58402635bb5b38eec4c61e8e52328b501371d532ec02862701302da2156
z2e7d7ba5ae2fe6c0b0bf7e9bc49f16e94b8ea58ef0baee86694bae976a97a932ef2c8263453b22
zd48baf5b91a83d4889671c1f2acd6ead5e0bff79359c612d9f17e062398bc5147cdb712243e65f
z54a6b5b9798f107d5b5be73541eb94c3b812715cc714c36f1e3e3880515cef85c2f32a15f19a83
ze2bb21301015039093d92ae7af9fa3e240d291449d36d23da43ab5c9ff37716799352970153425
z82ab44244876208658fc87be2b0b01f0c525b6f0a8926bfd0c765009a65723badb98687886c3f8
z63a34e83f39f8f766cbb5cd83d50ade66eef7b6809cf582d2458663f517caffe0d5bb8be98d31e
zed92abcbba92a25b41c80d8ae9aa9da4215fa692de1617d22055e9f47fa9bd4c3b287e46617fea
z3b9bbb3798b03294ade573d84338f8e4a251935d86cecb72efc5a9bc93f4e362e07227b0178d05
z84b4e0d45fd6dec8cdb88c23a29675a5031e66039482916960daa536864dd82a29002e7ad61538
z44865600866f61a3002db8d98121a264768c96dcf69316b4be1c680bba2cd6b06c04e2de4528f1
z2caf29954a28d7fdb406953dfa65cb6aaa8e3df8cc71e46cd9ef346a58f079a2ffea58ae984e1e
z604ffaea2693a6cb388761cee416b52f0c06d8dddf1cbd817e996f34973f18a80f8503cf6f4813
z0ffa15823e5d49216c5452e3925b3ccf56b401e4f51e2eeca4114bf90796387a16eb4439789e81
z7ac38429084542600e1cc13ee62d36754f9a688816af0780e6f7b7fc592f6b5394cb4631a5f60a
z75066727d0afba55e49d5a7ea78584309eacc0cd76f768f93479cc108c6e246923d622defcfee2
zc1a15880d796d6fcec41ceb9118174a489702ea1345da6aae00c37b3e5964552a18f50eafe99a4
zba2eb8b9a1eaf74be22681a1aecf24e35ffeace05fa27a870d14635f9228a0c3810d9b3690ddd9
z63f4855322999eedffba8ea864e27fa70cc38b798fb0e18ee90e84651441300bd0b38415039cdb
zd57b6b09d6b3a3e26454edef6a5fa134ff46e122c73d882b4b29b142d7657bdeedb935c99e20ff
zc46cfea3b014ea8642e622e30a0027cce5b926f04d0a61178952a50c58e84d92ce33a78fea65ea
z86aab15d59fe68549c1a326bee4389e8ef75fcfa03afa044adef0c2ebe0b782981c15bcf82d62d
zd1b4cabf1427532974cc2db3cfd2757b5bc97d77fd1c31042976751c493a4c269a9fb2539b2d96
z0cc1c2465e552eec43f5e2e2efc0e9315412b2d42b66c05af185968cd53d1327dabfa9545028ac
z2737b6a33ea8bca04bc5e0f33ef043834ad2b62a8f9cb0894847cdb823e1b3f3ff38a39b09413c
zc197d71a87b52c286dd26e6fe317f6f1107f44422303b793ccf7619480d84e877775f4f7a40e30
z427453122fa2026af39202c5b982d9208ec2e14a2aaf0b61ad245f4b9038e9c15e85ca930c65c9
za8868724ea87979508891c8478c1199837bffb20184feebb56fdd2c438cf1d5d224b2f96c40273
zae68fcc3a2bef8ebf197da383e48233f084156b5418352a285d9c332dff45548b45ba86890e4f8
z2299385ddff9a874e569b2b8943dabd80ad8b4631991b79adfd50cd9f56a87ee63bed0ebb33ea3
zb1537703090cbe72c154d7a78cf6089c53edfae57dfc1f275a61996fff5625cf76aaed506b21b9
z11d4bdaf2cd3aee91520cab222b07420bfbe5b468317e299050b8f5736b5d6d0de0c8fbe7eae87
zd701c166f559c1523a1e3cf0b2f3a5747df86222f25aad1a26529cf03c1b49ace9c70ad351e244
z5388ea449ec3471a96ab49b8413716ebee3b3c16fa380dd82ba194a9e88ab90804398c96a86556
z93154e949096d95268e3bc05475f9715939875400c55767d2d4833b2a0ca163ccdd7eb84a6abd5
z8b57b1d3fc4e0675d82a8a4558f4521f9b7f69595245c76e5bb071a3127ae4fdc3259519a94802
z189c871e9bc21c1da4f9537de53b575e0e0c0fe1f6265d34d7c7e62b46e67356ab27d0dc866cb2
z9b8f834c150f6b2ade46906747d984568eea8dd45a004c62fe82aaa3c94d1c687a9399b38a4a1c
zb0a5ea6d26128e514b562f13b5858ed0a05f25df23cd22085850d6355b9ddcc1d39592ec9d8f3e
z225e9671b555d8144139a3cb6adc6c679bb193846bcb71ed17cd8ef7a043309ff53079cd12f8ce
z528f97585af8bd8f0f59c06745b0759fad6d8e7c0902ace2a57f2ed4d1259ff80c088a8b0309a3
zc4345709d1833bec5c68f915e27bcc56ca79cd7decb775236cdb71086de7d19b3d42bee40c790a
z675c2c258929b0ff931345e969ce25d59bf07ed83fa0ea93440e6c6e89ee7ee0a2234004c11429
ze4e078135c02984846d552f8c8106972f50343078e1d3e73466e76b2ecacae848eb90cc25b65f6
z922826ca9ae1b54a4d6ad46073b13018685bcd92aee00d79274391ed2fe98cfa5c7b2071baca2b
z3366853e439d79b49a2960b99071e08516d584be980288598a89bce286a93e4ea00c18e44ea8e6
z8a70040b1131b630dc0d10ea6325a1dbdc399895dac4084dcd6d9634be72898306905ed8277987
z8f54c14ca91aa5b439931b31e127a9e717b8bb002471b0329a958abb29006870865152117842e5
zea4d2874100d963ee07dbfe8696d19ef5745a9497e86b45457c0ea6bbc275c08539f62d6c81355
z710bc01f53bf9642f3334486102d34762dbe73d094f2e94420a35a0fffa17eedecf8b657205f82
z5a89e9ed8f2a7ca6723dd4a505c70f70682d8d9959742f0a6e71f9aa18d10612ec97a4df2156ba
z71a3638745a3c29238d644f225ff0ecb3a9bc95a45854cd0ad68a48b5ae3380180d9fff80d8a24
z975b2ff3141fd93754ef91c2eda4f6701b900acd999421d5e9447ebee5534ed5419ee79020c50b
z87eac843489b48ec738a5845292297116dc81a83f18bf5acaf51d99e1487a8c8a77cd091ce4a6f
z1fc0f944bef82f6a5b1683b7001cd973c723ab7063dad2ec0a052b45d99919169a3f104ba9683e
zcbb10f45853bd8d2305e661a577c3734d105977416006c4d9f1977eaae46baf3982215f26c46aa
z1049046b82be47d9a60bcae825cbf9b7c2097c410b9cc3e1c6a95cea86af0d16a6b08088cff623
z5ed02d6d5012466166abd7644e6858753804d425bbc6bb3fab017b1e03b75d979dcc5fe3955707
z48f2319ba3cacc997eb253a8a264fec05903d4bc0fa4a58b9640dd62b037d4df88f884c4c5b6f4
z9f6a76b916ccd7df9a99b05b314582d7cb31fde1b0898af6b3b39a0598fd5c5226a8fb6fe643b5
z74017945a3ee66cdee59932ed144e3bfae21c32b21ac6e13b339a99b00455505ef383c12bf1f65
z8ada81e553c40c916beab3952deff62d7dd21d1a910d49342d3963eec95c1c1beae245f2d27e4b
z99c7e6b5f2225cb4f74a110566a01ed8cd8a16d2cb58b6325eb7e3169317cfd97dcefd8bb0d442
za6c1a3ace6d949e7eed914d64634a78e0beb1c520e07933c4d9e440bd493af7b8606ec5c3e5247
z1635044e8bf3d6e978d926734e85881690c3d7838e40a8f310e762ada29699c9ce320e57d10f48
z433cae9390a8b28e1da3bcc96a2edc849174ecea8255b97fa1b6373d433ff7eb152c7ca6d33cbd
zc73d6cf5ba639152d4ef25c66d43cc30bbb7944b938b4c317ae3fe62c5c252bdcffdc0ba4adcc2
z95338a89dca3227edc87759972549d5db94e686f8ea379f6d8700bdbd71f22ef6c1bf5f010c95a
z5fe764afea9ca2b6fb98ea848c97ca51d572a7d657d9ec228514fdcdde209732c0804098a47b51
z05a32033b4e39d1a6ca0788b1cf2b0ca21c993eef89ff86a1729f961d70498a7ebf798d2a0192f
z5222e95a48a540032149e4ad57e3eaa131e89e4151f8f6433b9f19d54ecb8cef47093ca327c9fb
zf251e64c13a8a10109a98ef12e5428b519b4687484e0759f8bdf5f2ab6cda188ec1b4d9de5ad38
z74a500c5d9f8c9e1625e25ec9a9856ccf30b298f78549e115e3678e1b9176ca2cf668dd38bda76
za82cdc25a00b88ec099cf60ef382dbebdf5567f8ce295fd493c5bf1343f649b484298cd8ea5b73
ze112f0e301395ab9cd423909e8f0b6a60a5d95560a3b166ad4195eb2e40ac30c00969a2df4a8d9
z0e6f86d9e9441530ef6948b492cccd8a988dcacf5cc11392fdb2c924d30770254b12b362e360e2
z180ff538539664a040a89951d692e0762cfaef83a8ab69ff9723223483b0fea5771881e6cdc651
z5be95824d16a02d1787a8d4ba94439ce3d3cf2f4c2a25d7334040d23c0aa9a9a5c938ad9f012aa
z943085c00d20c69144dd45e3d7cf2c53192fa15a9cab4ef69230273e59eecf0fa847da378f9828
z865de29bb549a599e0e50a96bf90e74ffb48c112cf3695ed29b80912aed3cfa1d4724aea4206e9
zddf9d52919fa1d96eddc93aab305830c472f2d4a758b0c960d006e217bd44ae6e0337ec8f37330
ze5172698311314c3a09b1b2e173e0d383345f889ae6086aac8b878374184df64dda98d107fea7e
z8ea888d6662ab7c6e72c46999cbf773c9cabce113094bb2bd15139b69dda5581926b6ed66197b4
z771431dbb12a67faddf5958aa63f9b0a98c8a5d25b6aafb32fba7c0d26865d52cbfc2e648bc25b
zbfa33b039ea98ae1ecd1678db2c35c184be79264df77dc3902a194ac16f7e145314edfea0e0e91
z0d650fede65ec3434ea87f673a78fda1395b2b44818cfce244ef0a0b6838fd9c2fda3116a25dd9
z377203fd1ebb2b412f01dc2ac4244b68535d960783d9a133f4d918976b901b6d698554ed5a1512
z5cb4cdf5f41e4bc813059109539199c01647d76e39b88d415b7b32620189287c248f8b07ef0de8
zcf24657d7d0b7dfa36d1441e835a209f6196f8825740a77159958014f3371e339f93e0135961a3
z64ff78f87985bbfa2cb7f265f1c0ee021e18efbbdb1c7fcf61cc8b64f3866a7d6239038bdf0c78
z0ab9b86e7d15465637cdf012aef77baf4521ead09cab0979533c91c4e2f040c1171a8f212f2368
z08e89dac36925e4d11c92d07c4e885bc4bab446803efc1bc6811fddd456666e87724ba43ce901c
z1fc4c8e124a366089bb440de60cb8073bbcd2959c75709bfb27c34eb6ca0e4e72045188d1c1f11
z4ec337260d3e1900eade2d32c8b16ad9c6be70bcadc6afd40a9f3647b502fa3be820037cbfdfec
z6474f4400c1e7a58ad2e006e052628888e89f316f03ec001e800b7f0e4ce500b7e8fe74de79c33
z0923a02ccb2fd3a030ab22309f33d5dc1e10c8890d93f87cfb36fb56dd5206d8522abfd2fb4ff9
z4d62d36041438a28e11f7bf288781265fb780e73beea194b82db8f566aa8257a682f7e6696a36c
z01f998a58c4e06646ed446cb0c7444287b426245e553c89028110dd09dbc60c4812e0e9964c1a0
ze6181d06c5db01a5ca3ec310ec9d3c2e7cf479e3579194a60f4df950ceb6602b8f3f1bada693a1
z9767f15e0ba908b122affbcb8eca5f15c4e8d7576873bd0f6abd718d876518035b6c11334f50d4
zade3c7aba3eed419e55f67b6f85b61aadec6750cfdb8ffe0f55fa50f17f64206a7b47cffb2444e
zc6355d5ab06ebd7a10a58772ae04d7a5420d391f9c31c5c73fb337d89feb0aec64600331054215
zbfe971efa4d386410464ec568e4481a5d665919b181e6ae9a7e621d448a92ada89c1f1f089b72b
z66527a82fd934381d5fb182f75f9c5c890f8318f92c2792c6bb879849334d41935a3891b169275
zc9e500f854e7f89f5686f8a514711b7eadd138cf937e7594849324ee0a41979007160133fa34dc
z79720b2d60b29d27272c890700c8985f72a375cbd5985f82c190bca087e34bb3fbba71887537b8
zbe1c7528811dc7fd0b895eb0d82a7110cf41f1520dffd4390e49cc870b2d15ff1ee04a6913b729
z6eddb07afaf685fb3ce7c8db1d32ab373b1f22691f8b29ab969e951fab6c1e0a96adbe2cfafde8
zb5af524f5e6c35e63a689521d5f750e9cffa49aa7d36d942501f469b1bbfafa18ab75c0bd02e69
zb677ee0588ad0a49f74297c25b25223609ab8063cb6b5c8d84f6180675a040cf9efa50535ea814
zc592722a72734c08c0487ab46b532b4ab5bb7b5d0c3fc9aa9961dd43244ade9288f639e008e5ce
z9363865ded68a241f1712091b1dbc2a643fbc51d7341d53d9414e1827a81321702c1c1eb80a7e6
z427c292d85bf232af4d9d19cb5236a1700f274885584ba1cdd8b14ddbf03811b70198102753ca9
zc02454c2d29a1553ae04d95132c0aa1f188291b34b2ac354cc7413750ffad42bb3b5be6b082741
z54e4e8548caa859f7ff2a7d0f69a2675d1afb0a42f786d673ea2787ffd6eeff19db7b2d14a46a8
z09418a6b4e1f361715f914550920a5c43de3901b856e9e29beed5e2543ef65b184ac6d6531de71
zb0e0399db411833f8172e498e573b52aabedbe40a870594226b31e14945057de1d8e4c6de55248
z0e428d2f2c06ded9c8bd030724ce8f7643446df42873b85b38174fc831730912e2a03ed3fff4bd
z5d32ea9e0e911b7b86c8937ef804c267a3e6f6351abffeb06afa17520051a25b971f95ef07440f
zbf62bdcce277d0d3fe67dde9a0594db1bff9ee5d30bb94737735f0869d6fbc5fe4a4f0b480a75e
zae1fc0e5819fcc32ad21d84b0420850e26368d4fb6f92affb991cb8c5dc039dac7af40f0f86c98
z737b8840aee66115d385ebfa38507dde1d0a9bdbade77dd1b24ba9fc37bbaade9d990ade57f987
z2c83fe13558a805891a6b0cf4b27d4c768d66ec66cd908fa78987e7e1ac1de766916863007afad
zbe5c6403ea445e28195e94faf03b0706e3f00094a08a1eda3b62d64e39d2f3e78728490634e14a
ze0e9e424765e499cac1bc5a76d6353c1b63aeb5f25f0648e6c378482fe9dfa7b67e47441b3c8d0
zca1bb66276bc875b92a246143a10ab9d66a618770a17f12b3421d96103d8ac50c42c3875149f88
zd1a4e20701c7621350a4df3328539dd542b786ab63101a7cf451b5a0590f80d4d1bca23ec1b6ba
zba752b728ae949451625476e46342fe235c347756a0b42d491590578902388919d457195325c45
zfa3131a59983ac8e349f16849956b8f81a80d81d3438fa0b2e9031c4658c2c9fc47cfd93e3f091
z4df3fd711a578845b07da8a639c83af7eed1b04a842f42b70612776cc7ddd138f8fa6296c3390e
z952d7fd9de0ea4956314be0ff6a95988d80ea4bbc96e43f199e33131dcc36e7d80b921567ea669
z8bd35e8dcc26deb42b8ac1791fca98dd5d6aed7361c1d43f662b32e941456fd40f022990ec8c11
zdd7bb19cbc4a5b26326b0ce15d919a61c1353fec0599745071a55ec6250d19bd91df7914858166
z3a441623825b32c118850d022da22111791a51e96b403300c6d326d1e88dd406fe77bbe5b2d936
zf577f7d24b78bf32e10c2b1901cb068fce339200798c6ca7f098dfee45bf3111738384ef2bbf30
z117db0dd31ba7c4f6f93bf28ba0bb81d09808e2f0a20466f8936877ed89455694d0412d19205cf
z6967c63ce91fdb59590eed31e423d8867954ab2fac52362baff2a64dce7fdcc76786d9521f97ef
zfaa7d1ab4f19734b293c3dee14ab7e490d93c411b224cc38f3d95d8dda447e94ba6fd388dc0619
z5224f186db5f884b10c705ea6f72f20a87cb5fabfd859d2367ba3fe2da48ac25346e7c5ea93b0f
z41ee97eb0364c2d631587506ca091e39bd8927a433ae81ebc11129101d3410414143ecf518ca57
z6340cf751b28e0d3e4f2bd523a2cf9b866833ab0dc285d02ae532bdcfa4bb99fe3f374b7a6f9da
ze8fef1a44ced8f50b4916ddbe30065c309816ebd4255ce26614d715d167642cc949d7ce4646370
zaee132cc42045e2f1f9f84624129691f79b4c29cbe09115713911ea724cc6d8008b5af1e952f0e
z0fabc9192f7e6ed18fc2f1507c44562fd4e55ee41f7ea1b55ff438507d841524579f650f294462
ze65a1e7dd9bd53f81dfac8970e43a41ca29bd4d4a27319cf9be5589bc056c8d1f58046b35604cf
z07cdfa05cdc223e62b8b3157c9f303c5e32cc363444fcbfca061fb9b39b6402dd5cde6b0ae4ca2
z0ea6934ed8e9a9928082f280ccf39d169ac5ca38d729540dad66be3f6fe562abf2b9f9c3e62db7
z5808c05bbbd203629aa72ac7ec013df0608422fd83dd3c5f83f176042993672e78fa2b6d9e0654
z8653da0e64ec7f4ee1439e6858b6e65f0503ef06d66b4fdb7c1ae6cbd36b28beeb9353ccd86f9c
z6db50dd5ce960bb62bcf1c8af5a4954d991f34f704a3a9f27aa73d72cd8734908c17539fb03ad9
z51bacfb3fd015ee9ce9f6c1605315dd45c1f26067e28c6e01fdd1518a52e6a8a9dcc4ed686f65c
z57391037eb2b7e6abab9ba4055d699d5ab63744bebc672133c86e29eb69e4228b151acc8904421
z2a4c364deb22c28a8595606f8e3fe7eacdfc7b27f9e8fc70df68476e9ab60807fb735fc6213f22
zaf2713b20c3354f07c2cc96995f0e2cf081547a018116396290dedf1ebfabb38182112a37e965a
z349c0a0f4e9b5cfb3cb9bdab767199473ae407759d2957b17c86a1aa2a894eb2688bbcabe6de89
z080b81964510d76172f7553ca72dd999f496c27f21c3a683375d17306cc7ad00d31ecf80824a44
z544c055dd298bef010ce2ebbcd1b32ca643f5c2f0a236396082e605c6f7c384d09c83a901e0709
zc44df700a6a65633d96187101c2d060aaed888f582ef7f2933c62baab6e826eb0b1c5cc7b3c452
z290c1662fb88f59b5bbde0f50bde833d9889bb982b942226627eb2556cad1d3a9b9b5f88786474
z463772f221f1343ab81469734b2ff499df54c636e32a46da2ffb4a3c898613a36aa0fd35b457c8
zfa5bc9c8e3381a97e3b826f2bc330c96c898154d1ccd3b8c68763492ba8d4b261cf8621287598e
zbe572d18dae2c1417f7cf56eef94601934fbe353c69cb044ea112dda51236e85728ba973b76261
z673063c496091b1b2a112c3f6c20eec6dee617f380f61b1e21be1462f732df83770914275245b3
z110a2a8940fbcd434ae07ecee4e0797c489810407d9f9660682efc3a482afa1a3cd952b1f4ffee
zbe57de111c717c4b92f06d46c8e03360cd2dcec392379fd8df5eba32648e34938705fda28bebde
za77afcfecc19224736337e21223caafe3f7cb30e838e8c84e8692817388824a199fcb09f28f4b7
za260f6495214cc5a82e96aa74a816b086c02e8da0bf7f144caf80605301b4135cb15c711fe4776
z45093b6e1e6aa06144e1db3b98a926e9e3442ac3ade14fa2844d8c0e96545820ed96ecd8cd6d7f
zdd337c4f7073c6258415f7f22ce9986b668bf543e20abd74dcace4a37ba9a5f6e4800cbf2f232c
z23dbb81aa3900f289e39c8589be7a49d1f6a075549d6e83ae39e69c9efd6b9d33c0c0a55c082ed
z9426147ca8f3984bd70d2363f4236cb42b96784edb1e1c937b6a7783973d66750b004720c03b4d
z9ea816976df66fd100f63515171bd43d4f53ae59836e893f2f1c5c5427ada8877723677edff452
zb37f8c633a43711e16b63d9a230098be553813a3f32d25f64fb5f9b1b8c35cc2f5656e47d2b6bc
z2a50bd4288a7e6932cda29721f1dae0a9a1e79023c57a4a5c7430c14f73775e2389dbfdc918cab
z566b8be06806fab6bad04c435e3f538e39b495b2c221ce82e1cdf9d8e7b706040e77d02ac1551a
ze4699ee2fa7356d509f90f8ee0c0fe282991a9784bde336a193708ef42df7043069d4d2a183f82
zff401dfb60b26809c662faee8fbd9888d7841d00869d037c2c3d6b347afd03ad0c5f29ea2d736b
zca0228ac705f139fbbe998726bc42c579ea852caa5883ac05cc1b3455668c30f2da7c1c3227b6c
z4a81d65e834ddae26a6c7949d2c47d7e365fb16381393ec599dba2caffa1cc100275c2e9aff5fc
ze1e5a99621ae4adbdf7a8fc7e6fdf1cc4a382a645b0e398652ebd933e358a304b900a79c6324cc
z2df913922cfe29b9bc5da7eab8a43ddaf18bedf7f47f9283af0a0ca664d09f61db9a69e56944db
z9d1d23115bef337922ad3fa0771fc01a4f4c624aa915a5b4acd100097924012533d5ae0a4eff20
z48cf1fbc509bb0397a77b13cfdbfe51a1c8bf2174ff9e91ac5d0090b08185fd360afaca361066f
z7f5922b4e9a12a6bd36f66fc8dd6e6a7823aacd772b22f6264fd7b1163dd6042642e0f3d30c23f
z34206c27330f85001b53aabba6ec9de0066534087a679230bafa08535feef9a38c1921123f48f2
z97bcc1720dddc7230bde0427d797d0e00a483c376f33700f80550cc27f1daefbd8191ae23e2383
z910587b933c61ef9dd60d1f0e36173c4320a92485ac366d7a8ccb346915fd4f30d33b5997e70e6
ze60cd11fecf42a95d409f468b5196edc2ce0c6d03795acfb928f5b30eb533852cf5c81467126de
z1806a1ffc63f5b5d62dfea597c65bf21ed02f2f0d8be758ec4b67cfc62ed9fcfc56d3e6d44beeb
z6a5b12e6cd468ee9fcd8554feb2ff0cbbe2910c72e00a8a3b3a790c080ff0cff55b4cb649c029d
zbf96cfc30c0ce4ba186dcabd72a4e162b50d52c918d0485195b2ee27b851bf33b334712232fd32
za581e278d9b0f4ae6b1707e7afa945ea1f855346d3161a65460afd1e2f09383d071b1b5cce41e2
z3a2f15b3265c9af70210ff28208960e92d684039798d1d70f8e6013c589b01ae58b66c838e9aed
zb1e8bcc7a9c01f8f16cbc75eac763cfc468c4f7a15bbdd348491938c9f8c1332e04da5964595dc
z6458ea3746f75bab4c7d35e4ffede2c9d5e5fee4b455cd1bd2f9bc324f5d6e9966b96710c1eb6a
zdb38df1d8a6fe9a285a1d1c6d60d617bce47989ac10139fd050197aa8c6ecab0e39eda487d2714
z66b30b4b4a51147925985f056e026f138503d8603fa3e1d33609e2927f9ac124399c691b0c4a0d
z3fdb5f7017ac58eeee0e2cd5366b77b8cf526464eda7670c71ffee648b7f77ed3256d30bad9f74
z6f38ffb85af9c4d13a61d073e606024cfcaa6d02841747497f4b2ccc3d17b8b4be3e8dc2e07cf5
ze7638ca91c6e3fd7d58e9dd0b6541f709515a77894d7152f03dbf97367be2efefba920426bb2f2
z3ac734c16c3de794c7f84d4ad51a8040d3a07f16300a1625c4e0faec190b3fb4df7d70625e36de
z42f3bc4eaa1b793a510a726cf676a8cb64d9c17f3d3c56b3cdba8e82e72974892048099e803baf
z199545c5c21ae93c8183cc0261b94fb1a187ef23880d087fcb583d5455fc3f2e3832e8071ec96c
ze44679b919a729dcd6c8975bd2bb4198bb147e7be78205f2baf4a7a719fe7a9a754b3c1ca07cc1
zf76e98e08393252b5e51e793dead16491cbcfcd9670b6ecc3e394abd71a1a99f4f3a49e20cf67e
zf8a26e16755bf0bfcc5d2e030904e3c7fb80b62ea257cb88509793bfd644019c0c1f366058bfe2
z38885cadf9c7d2c88389aedb89f9cb9d7e7b519f6d45ebf09c60e4edd1f2d329117f831ecb0684
z89ec6f669e8976708307b8cdfb9129f1d815f9b26a8309bc6b28611c50aad569db12a017b801f8
zbae9478e2960e83219965133222138bf4ef56746b144584bd7dc2e25f4ccde97eedce257320d8e
zf9a8246eda892afc411771e1c86bf4ce2b9aa2ea039baed7e4b8c80115404464d1311396b50cb2
z22d5d7fc494f81ddc9ab652fa639f70a3c2c83a84efe6ec4617d61bbbb8a32c45c70e3001ff081
zd25bfb7fb0d2c092470875beaf6756a0622b15217af2e7b03d7bee9d159cb33516930fa3b354a1
z6aa674b59a03b927c66b4c416dde0707d6250c781c2209b9e2eb50164bc53e4b6117b086a71d19
zcfb5a9fcc0f5625f44059112fc4358a7249c76e4e0b8f49da6df00fe9ccaad22c4eb2a5f97909b
z49bcaf3787603dfaee5be9d1494dfbe06fbe316d45a3a2f9fd22f626970df456becb67137d81bb
z337a8ece1e32bf7c749a84ca214c6c51b9a5e5612b24381f79161c05a9d7b181993537151a1869
zeb8257500829c50f7bea0c9cca642363b063a79b69a0f3f71e588e2d4f26ecd15e6a9ea4e524c8
z1e43dc85d8c6339a51077aa010729a545bb2d402987ca26e5c4bf46e18707d48485e92e47370c6
z403925d10c4e0226e0ad36443bc2bca8fa8561ca2e8c5c321b731cb36f869cb1bc42b6baf911c6
z584b993225e85b959d8140eb21ca1c74778df67790d685e460c2b0abf127f60363dcb42700d7d1
z0cd33a977ff39f3b249eb2d8f6977f846d1a07d56dee920728ac5432ac939f5363038658db9aae
zeacf746f97b47983247bec5c035d1115de207fa8e8a8e30795a841a225789ab3268d762c108036
z28c95a0ae2f50776341fcc63adeefcd7d5dbe9a4f4a1f317796b004e340d7ae40db1f03163389a
z7e1ce25101f1f6085c3364afaeca016a52a725145cf2910c681af2107110f2247130f895634ff8
z66e643d001fa72b17fb0f37cd710b77a5bbefb6e889e27cbac99837e4edaaa73ac373951dc2728
z088008f58b734fb2d5a62694c1d7721e7cf817491e9d3713796dc4cd507dd1625440a21d85b50e
zdb00d053a7282960ac594a767f554dca2e77f811d091ae0da85bcab2b6f8efad1b6acf30df1840
za067457359b48e89f5eda4df9a9f4e01317b423d665ede4dd7a60d7136d5803de4c179a1120515
zca6aa2557ec77870e4bfded33a7e2e40b61252efef495969b820d51017464677bde0ca55688134
zdd10c9f85db615e741ad707eafb5f07f80a4a33ceec54413b76b9ea37bab78781b3df2c8255805
z0a026b560eadda63cabcf6409d3efe26b3e9d70ec911f39fcc5ddc371b61f0615d1a724e39490e
z1209e238e06b35699c3325396e3cdf0142604353e17bd1143d325d4aa8c4da067463979b320e51
z7055bf480d98da5a3753db227e8046b2f7e1849fa73b824e0648343262d40386ca7d72ac8adac8
z8aa0df1ef383c9d918e90d60c3d64920494448311d85944b9f35f942b676a235540b701dcc208b
z13eb9bc1064e2c0c8dee5a60f64eb1b2d34cf1879627e2c27d1f20079ecd0b7f40ea42018eac46
z0679d7ea088b6b80165aba770e3b5e9c9323a41c4a83a8bd6f942a3712c3d7d95084c0508cd92a
z8cad278ca2a537e717e908fae8941ed44908b7f551ee15c97b2e0a957f498df0ff4219cef4cb5c
z288bd53f2e62cb253fe9a2acac0d844c382c7e851c1092c715bc355fec666a298cbec605cf365f
ze5b1887fbce10061b130afcc8c9afc621cd125cc9e0e9db2920bb60e925f08e1dd5664a58532b2
za39173a3fb40b8ca3953460a6b2c50381e432d17265a91daeec56eb90c79367ed89787c9c46e9e
z75c521cad84e2a4d85e8ebe6af9531085bd10de494d340b5d2758458ccd5e2099c26a3f9f9af52
z626b2a5bdfc1aabe489e3836a04670a959bef05361b2b9f3db91fae5a095b7360d5fc8bdc29309
z8672e3b4ae76cd9e748cff3b798c4eda0d6668566e2ed10c9e99a1f4dc8ba64f17d34ff3626662
z3926ba7524e1106864c59c8ee2b18ff86c787cddbf6437249c66e18b298318fbbb4b242b36465f
ze3d22e09f3f4f316a8b25d40a04d0ba71454e746092cd966d4456a0466df7a7643c23fb51632a9
zbde6ebd8437a61c97e19cb47c0566f7229493d21b22c69bf1a38c02e007fb4493810a78f3e760c
zd9dc91ba47ca7f6464343a492480f0e15992124381ec2f4ceac8ef2b845a920b72c12aec55af8a
z18f78d9c181fdbd841d75b1b6f441048a6e5f5715a92af664144c08e0988ec311e97c361d8db07
zc867e1c4fdf42357306fa301fb2b5017be96297669716c8bed80c3673c908167e3ff0485760b70
z40929e01c295547bafa29a244cf5c598b82fab338f57f394a926408a5b8aa4b7c57645c86bc484
z2c48085e78e47021493a0149692af30858cd732d50ac86078020f09a35a756cd9067e44ff4f26d
zfa705249429364d1afcdbd65b4b556ef3f9deeaba311c66ec982d00e2767fbeca50a0fb52f8447
zc89e30655da6a9b07961cf5f3ed99338db1b559b4d2029bc157407c916413a191b51bd2a7ed313
zb9de6b1b86a5219be2dc947ed282125b8096877adf61aac90c1d6b270615d5ac0224939341a59e
zb51054a0a8d54c84845bdc8e6edd907e2c9b0051797589a31c42d5866b9121c0884329a9d25e69
zde305856467565a7f4e7c1db2a99fd329a7c961da505dfe83060634d43836ef64f1b75cd6fbd7f
z742903fc4994c01adf013ab7ec3995997cf5b049eccbf5cca4fa35fe952bb28eab1e771d348c91
zab6d4efa55db7693465d41c326191e35ab2b351f0b0a11804c9615e6be84e3168d32ff52c6cbbc
z43f27a8eab4d476a7b4c37b7e9c1c4756d58b6b231d24c90902f3a1c628ade22e885a56a869f38
z7c624e8b0220909a40e631d7039ea34d1e33591b0ec09896b8ef264d0e111c619f8fa6b553f9e6
z0275101d3d518ff8eff1c1db5eaab35ae33294f6948c25fa6f421e4245253e10ee25e9eb9ed7a6
z3e9915daf1348ba08bd749a4749d28852196baa22d35b765bd2fdb2d97017d2333b3bb1f954ec2
zf4741821615f4f592eab958470328d21f2977f8913fcda8731e1ddc36d506908db3c48ce6f6d9e
z138582a645d3b6860329f0a16d803654d61ef596d3e99aa32abb48c5f72949be99c2cd696d7805
zce9f8b82ef37b0cdcab49c4405dd289e65c12e77e6c9cb9f0c5d42d3eb150f7aaafa427f9ca7ff
z6c4f28d9ac72462d90bb8379e24572e5e687138b653aebe40538b6ae5af0d29fef2752fb63499e
zbdf565ff15dcfcaa265098d48068b39c4d34c5eea5563b029c1466a0cfa4b5a84848db82bd58b7
z9f3eecd6deec5c8db81e4c4156dec4404d495d45042aa12feeebd4c6c98c39f3996744d878156b
z36a2a2dd0d6a22de8c75b4e42484548e5d31104cc4645fb000f23c442df1cdf08294c7617608b2
z6cfd2ea2c870027538f28ac9270fc8c12b199323d29373144e63bcedd47c85bb29559044a998cb
zd91164e29c8bf973f4b9c39beb3bdbcb812322da594d22bc5efae4e70b43f31b561cae387e4568
z4896fea95e08e6b97dcc2712bc81491e6eb5b9ac54c94004bebd0c374c7286c188d139dfc424c5
zd992a77a04e80d72a192519a8d2f28780445b67383d4678adc0212c260bc69924ce5089e800cea
z207b8d7032bace07ae45ed65264891f7de95b3a11be13dd365302c4795b2795bc5667d7d529ba3
zac1549f06b82fe7bb36f66f158396e2c9272bca1a2d37bd547a50bf6f64f804622d277bcc2124a
zaaa5645dc352a17476e864dc19dce5f6ea83d187c0659542013b13aa81b1d617b864da3274b2f9
ze33bdec2e86aadc387826eb631a99a848df4f44cfa96d01a50e5f8409481edc76a8423841f60fe
zed2568b01bc254b5ac7676671248bb910df8ead2dd3d4b432e6bb59954bb75be9705b4478ba7b9
z4bd81eb548c4736bbb33b407218b26f1175e5849348830934010f1023bf618757aa97df4ef1776
z88406b3c9d40a3ca91d08e7f17aebf9df34d8c057a0029fede7c78ea21b63248fb5bc9557234fd
z5d83bc98c210bf59dc47d2df8b7c90f2bf886eae648cfe161d0381d637d8f54bca76bf191c48c6
zfe980f35192af6c3d59f9914d652f43f3be950fbef30e70eb34f101fc343eb4f84a55f48e8ff65
zc1aeb60ef81abf0d0cc7242f79c1872a6157131773e9a3b36a1505f045038c88afcb62115eba5a
z4b921fc610a7e15858555628bb5fa9d39e49d3feae7754caf30966f3997da5e04737ccfb30039c
zb943ba0cee0113f0036577d6a4d294e97b88d62c68ab28a819957c03379f14b19533d87c4c2122
zef983314eac78dc834b039505fb5b9577333c6102ec9c552ad7c9a1ffe2c73ea1f12b3ae6f1024
z8b86b561a5a519a6915bfe1d83a9b127219280cf2e570bc5317f3507a17fc95e8935e4032337f6
z175845acf1a1f79911b9c79316420eb445cefa3c89605d7cb70872c421b18b986cbea6004f65bf
zfe4503441a6d19bdbe5271515955cbdc0e5d7fe08943f212e7ab7f32ac24164bcd6bf3aad486e5
z18cd2c026e3b9150dd89b046c179a2cb5724758159c22fdfccb8b0204ca2196de6aa29ccebb451
zedfb8030cf8c641ed7f106da15daab9fd9b71699426cb4315ee48d013d09002a4b25a006d65383
zc897e99fc6a29c1a66b7b72cfdd7cd623d291494d1c40b2c485d2e3b68d252c20d507bb2e05503
z2731b31ddde9a01ec9c81939420e7fe3b2f3a52ac9ed357a36b3ac0434b8cf47ce2548625bab63
z6c2408c4e0926373aadf149fcb5cdb934fd4b0b37b08acbcf0fef3f2b1552cc9187bba309cb554
z406fbf6391c24c74ad8b6312c929db4f94300042d7202807cbcaa6a63892055742c43f64687866
z0ccdf4ea10643bee7983684bda0d8dabfe7c7cc665eb34cd096204992c2bd09f666d7ae8540b7f
z8a9c485a5b4a64cfb4d56c9d4be08d7c61cc6e0b001a82f8e2a3c165ba05e4068a57b421597fb1
z0327d96b1e2274eb93c645d9fb43443f8eaeb9ad4bb97fd67fd08db4c143e32116bd2f8bc516ee
z7e4515302166372e664928d54860d8efc72c4cc1c4d25ef48406ad7ef54bc7904247202c5e6c88
zbc50d3822790d29c461ca2721c19e417e2cd0123406a7258a05fcb6c8bf3246889ffbd05e6e2e9
z2934edf2b2d7a1aa4bec0db6249b29f742458a72c997c95925cac2fe8502096938d18c63956c8a
zdd69be675ebc38a403cc2a09615365dbf951bfeef48d4d055d6ce6e6a3a5883b8705fe3419a43d
z4d41431fac9f3c4afb752d644bc7c21ec0335eee41354900e2781d3ef790784b8d4fc82afb33c4
z31c83c4d59ea180cdbe860b7d09f52ee7c5f3429979b2761fe42caf6aa24874ca7689b511ae60b
zb07f797c4d0729937838ad6ac59dbe05f9acd4d8b324330310bba06ef52f7b3bca558669ed7cbe
z67c6482d55253c4503c525a77f7e00bb06249f31eedab23e55df613a287057626d071d306bf211
z0573c89c4b36d79e7a94cd71a19f4adfe52d0828c5de3148494d040f14f3637246e8f0664019bb
z5751b250b12aab2366ef54fa41b7f66519204c8a3fd05e38ca577ef2e5b90dc2c22b6db01ff181
z5828c527de2d223340285357c8a25ccb4525ba5df5a5eb837475dd7219d094e3015497caf6eb40
z620ad00a60ec671e25a1db592f834994a1a1c13559f62c2722dfbfb99cef7ee1070ba10cf615f5
zce1c55948ea810ce2096c217e5058bf54e49540394fb5e445696171fc89fd0b6fcf101bd35a857
z6964666a639d6f60cf1551f7307ab6a86c7ac906cddaba7848db9c0fe57e26db14daee855569b0
z685de886381cb069ffe638ecf8c46b45c68adf8746aa728ca790432dad3439df7ded66df6140ac
zf0992a3c88a994fd8755277d780f474adceb58e061718c0c4181f93c860738665f553b4e83b31b
z30ee128e2805150ee9f8c68e0393b23d1b555611bb550e9701b4f31ea744cf924d17b090474e5d
zf7ab25e1c27c42b9ea6af3464a45a5c9182f672736fd1d0d1a468d9cd2b440f6da0a5a29bd2a7d
zd275b9c3ad6074c1e234a553eb8e8c015acb89c2a27378256f6643995206e0996d99c03e3cde2d
z0646b7e523ab5c49abd781c34e58df17efbb5f1e1cd61831d6fe0a880df53d16d34eb68bf395ab
z6dbacc8f27dc1c07b56080014a678826e53e848318caaef25c7e85049369e060f98cc4ecbab170
z3adebc073eee5ca49fd3bb32da362d1675d15e09637b70422b1c495e39339282bda38d70e498be
z05d4e04919c4056ba7ffd25ce043f2c73ad9366e7d3e913e8b47070fad13b5a6719ddd00826df8
zd083fdc250671584fbdf4b38735f2f43100fa47958a67f97068f81f20c49f68c2de72c63040094
z9d1dfcb3ba140ddc0331b750cda7fd7c8a47b5ec6e422635e634f7c0388267204ae22262a3321e
ze73c4468c5e310e670d1584170455c245522cbd7d762fe0343551d9a01e8e1e7aa52c427c34bdc
z9be66f1eafb5db9dc91a0c7b410999fac1fe00bd0b2d8d6a8d6b4c5c577fbfae7cda2bbfab340e
zb07123b247036058283bdfc152be6112ea763b919ed08c53971997a24a808d36e8118e2ab76149
zc9497857adb629898745dbb3c9ffbd39c9df981d75978102a0de49f86fb0331fab52c50c1b512f
z5174b1e3d74c46452415960057abb3712b3d139ff26c7a880c95a7ddb025a31f2cd13fba1d3b20
z745c19a8dbc931bd9ab8f031b25fcf9b5f2d41f9347326cfb487c45d67316c65333479dc4a45dc
zbd05383da4490bdcc4b54208a23063869dbb8660fefaf9ef11779af55d1facab22c21c923103ec
z5e9f5e49a96558872c53f65b5a24bc321f93bb754fb39a25d04ab42c85c79ec4def00d39dbee26
z347aee30a9a06a7cda2c716e81a91f2a7bc1996e015e1f8c46f9df9312d78fd2e1260502f16110
z44f6c86b7e87d2576594e7249cf56cff9331bd1183d9ff1e0e8211787bae713cea1674587cf6fd
z34d5d1332c243c81a537a0ba08b4a420446745f737d602c764b79c8524cf0cdabadaea68262981
z755a99c75f12a141f584788d946e5784535e38d789cc793f3e8203e9e437413ea882a767f739c4
zb3065e67ccf870106d1bd054da234cfbe07624b4b59089a731c372b534abf19396eccb60b1d822
zc5f49a874a67365e9b2c16871b0764cbc738491103d8a47e72bb785cfcbd0117d0f9d3fb9c3ff0
zd1d6e564595bc543a73e4bf12944c043daea6127a883945871663d794684598a829bc30b5b3ede
zfdf55bcbe2615b6a186b98367c6051c034d30bb4be19af40f0c082dbba28d0cbffdbd664f66557
zc8cfd8b9320dc1359160a525f72ed2f1195995be9a58f1ea181c3c4cfc0c4bbc55c1e591d30f40
zc1623ee7f3416a018317232922d57c4bf5c16938d3530d2549e41d17178ec350de562d40b41a08
z37382fb3ebd35d5340e650b4f2e12628a8b8e99dd070c027d5de541664c75b9150075889a8f3e9
z9a281ca6bb3d0716ee9b7949467ada4070dd911ebbf85a36a158e066eecfe9cd1864bfb6a7139b
z0b71d669678e3d402c918df6b91a467ad8b34c933d1704aedfa8b19506805f77beb1dfa9bea2bf
z907e564cc351c8171455826ee47cd809a81dec2353ee36bdc739a314db00c08cc17223a6bcf1ab
z8be9a72fd070132b826f48abb3f8787386854204f4370dfc0e7b37056aeab5c551e5f61db2c574
z5523e637d6b33639017f44a5aa45b91671402ff2e7b0a2f80f3c56aea174ea84e0750ee944738a
z0d99bb8544578068264c4f342c91ef0bfb3902ad2da791cce77c88f1504620a9ee17407a6ac232
zfcc49d7a40bc102122b2547b5d4794bcc316fc55f44ab4679fe48372f6fd799ca2e0840d173bd9
z99091dc1c7c4ab7218ca9a7010130eddb0f55ff18646ec219427363147ec4688a681d62dedaf46
zda3cf1f0a6e4d2e20df2a581747a17938409c38290be332aafa7e7ebcac6f216847abc00317775
z33a2b770d367c6446f317a321117f82466d497874ea2b70f777297c7f6ce5206a94071615d3ce8
z9c272f0a6315a01d30c08349935ab04aead7e82fa58acdb7ed4d7fd3709889bc739023ecb2bc8b
z8f52998ef6588f3c594bd4060873b000d13e6f229605c339b5cb2a273d3c23c7fd97eb40fd42e5
zd4e1c221a71afc2eaa46f1217a1764384020d15b7365cce9a017b104594ceb25fd00b8c641416f
zdb2fabb28bc7727185a810d582b10706f12d2f36a6c303906d1756c756838f9dafce313a7671fc
zeb773e93fa92e20c5bd43ff8e6ab13f5ed38a4922e99b5ec97300f0aa4931f154f911730413999
z18dcf924fbc26b6462f40cd4a7c1f51a0e9677a76dfdd4ad23bec1fa7fc8c5f558042e863a3aaa
z6e4ff8056ae1f4ed092d77cc2a328afd864647407cc279a15619fbfdf32ffe4433691fb91c47dc
zd22bebbf12e41e7383bc7d2b83c8a60f98d11aecce802669db62ea4219726e4334144e089f0cd1
zd4f8f50d8e4baf8904d791874999f3e7474b89b82c3b105bc2d378e96d8388a1a4cdac15362d21
z00d6998989129d2066b178f6a92316a5831b69e9c213f39de32f3eeabc1f87b6755cace0daa9fa
z98ea7c6a64b29e1c6c1634362452ca75fae93ba11058e8eea9ecde9bd33a3f1ead46fe2afdda14
z1e35e2cfc071b0ca2dc529b4d6310845e292ddbc7d0e0826e82a974d10d56bdaa08774d550eff8
zc3a8e4f8c0e2e21d197b15aba4199f4f854a266de107a11a3d92337516aef5c46805c50afb9c0c
z5a7c560776ab9773de085b66cf19aa4c24a09b4dac57dc97a5a9997b6c4b65d6a71f4765af29dd
z0cebcc86b76c8c4052372f035ad46080fa440be0a9d008cda00ecc6f3781b5f74d982777d82dd1
z11ec4648a593665b27a71519a67c58bb8609857aad45fb2bae9e6f595f04c72245c3a9a5232594
z2a877cc56ba648dfa8ed32494fff47c52eb64918565ab4e018edd67af898b2ec4c1b0d7a9dbeda
z0c316393bbb112a43a93d30b566acf3b9cab934ee35bf0528edfe172c0d1f4f5db270094b289f1
zcdc08ac1252a48c7d6444ebafe0a5cf88e0b492cebc906dc6f1ba4417a992fd8f30823b67d417d
z35861f54739f97ec26e1c1955cc7acdd028037aa9c7b6526e2b4ed0b78a07e4bb06d368bdd75e8
z8a626d90c34ef71a276ff3c974311ec9fff174519d9033cfb8734111278bb56b09fd59ed18b1ed
z82363d49443250315c925f7a5cdc73f5184774d6f91f4cf20d0bbaa91c483aee6261b63420c966
zc889d6208fae50a3767d4a73681f9079870126279496377b62174d89ee114062a4f42617d6d26c
z56216fe644b30a6054459e6faf8dc6840e925593ba96b059c92a19d66122a2489a2f0bb2162e82
z089d2c7db67a8398104986c20d86c264b9029a77422ebafe2f22bd48e0f50f497674781d5a53b1
zf35d66be40c6873589cb5733439eaeda3ff9ee7217da6015c485e4e530cd247e38589a4dc69316
z391b82aebb83efc774e983d023ab820a09c100df2f2086047af210e82ef1a1fb2424d1284089f0
zc43086f9053ebb697b3c121c47b018e3832b2fb2663cc961c8df388abb1774f021db3b228c6bcf
ze4b945fbab010cdc43aaa2b5bb14b6a6883058e28af8e9f7d478781815a54f7e05d10e06833cc6
zf72d1bf1d52a31cea02740103228d65ca2ff992e64b35ca926aa0999065a23347a665419addd71
zed0b7c1690fa11aa7d12f8a3ef39591ed2d9485aa8531ee0fe3fc3063ac9e2edf95f4a42004174
zd28690330f921d1ec56b4968e26d62a9d2a74f046ef06cc97899d6b714267b085783f266a382c7
zf00777deb2d2a69a226d089d8fce018500cbdb42a856e1bafaa823d0456529dc96c550db7fdf31
z675491bfb96b8cccb3cdc1698eeac81278fa52295831ea02ae4350f709658f35311a400cf94913
ze3c11fca74dfdbbd68ea91884147aed08629fba6d7fae0d3b8c55d8107b3a0d2746d4ff485228e
zf51895c56373120549f41cf27ddfe1f9465c3432b631f1d096413ecff93c97820d8227888d6840
zd9d9e52fa8ed1a88bba0744347d2e58d090658bb227bfa427cb3f4822ae8471fa6bf8bdb988029
z56ba9cbecf5c95f8bfc4a4f2f6b61f11191ce898a6a3c7358ca4b19d99deb58c6b4a8b2c02e41c
zcade2f70088123f2e432c99f9b0c24f3148bb05bbc828081c759eccdd34d495dc9f3e12d0a886a
z697385e9dd126741cec7bc541f8767b736aadf8a57314dcb07a860ba8f691fdc0270a27951318f
z2e13b54b97d175e7449f3e3e0ecd2dac680c4ba64d485ffbc6404c4aada58c436eb060f53ead06
z43c853b6087cf17375f6d2cc22796a4fff1f9b819051218502776f9c12d4f9c6da78a61716ea4a
zccf57243b725d14201ae6462e2df69fcacb0e5260be79a8a93934cf36016b27dcd22c78832f0ac
z5eb18c7d5a5604674e91a95e2f5210c1de63c78148fa4e7d1b50a54bbb59bb8b4c1255801d3d76
zdd977c2f0cba6d9d2fc523f1b885297e98e9943f68403974e648df503dc21788aaa90966857433
z48b39f129f5bdeae1df6ee1346df03de2488f0246a2a3b4e87e420e57ba50690b30cd34f97ecd0
z68cc7645628d244841c7f9b4533625ee30b2eb46bc084cb90b563cb80ad3cecb183315f3cf8314
z10998b45e734e82c0d4c1e31bdf20383b186fca8e911bed419f662d74ed90e9671e5ac9b69159b
z83f04208ebe652f8fe5eb83496ea1484fcdafce0de0c4e989d1e49e1cb77b3d6549b046bcdad71
z47ec5bc7110b10cd4d4f73e2ff7b4612fc6a02b83dc96fc2a5053ece002839f729e46b429bda55
z14d72d4fef59616bc8482d3137e2d56731f4a124bd1a6ff27c66e55955b056b7a265595986fc25
zcc542238e61441877dc463e0eac64320be77ce149fa9ef6552b96593285928c5ec14205acd0e67
zf61679d8015b511b4c26fe920e1248c7480ec8363b94a6af2905b4edaecbfd15aac552c01fa965
z0a292758b6a13eba05e735e08bf9a5214939beb0f95eeb841966284ce4ba70a576b851364c6c17
z86f124e737d58bca9b3ae3ec1b4cf5b016c82d3b82e82338d6c7f93fda520997621cece8d9095f
zd25da889d0b689aaa1016a39b62f1fdcefdb4e8e11f1a308c71c424bcbe5c99c99d82c45406572
zde49de5f11b5087e710f72c78c278da4934397b455b019c1337951c8690c76284dbaac6f987b76
z27fc853edb31beb073220dda9c38a2267362ddbe1116df82122e9133d01630c66ac565d7d6275b
z6ab26601e20c0de7a5b21c04ff7a85b8e2a73773f4c054cb43b96a2a2e86a465342b033883b16b
z75815d3763e1077adf668a5f4c94aa5c97c275e7b208a3ff6ef257c772a0223154367383b58d21
z553366db4ba0983b7f152507a05724ad4510177c6aa74e98b4017c7df14276eb2ae846d45c2c54
zef0ba448cc59faf310c521535492303aead00c32c33339fa1ee2e88571f46242352072d0847cc3
zd60a9b29f5dfbd14a482b9e6801f3a64e23d31145ed9a173614f28bc1c7f1df5783508c984ef0d
z8d7ef948e488f28dce907d0459456f97bbbc21f230d58a635e423b39ce6a6a019720fc8e900c61
zf32a6ba388aef48507bdfab51a7c6d29cb07c57eedf6898012c48012fd15e264b6cb57ff50cb79
z4aaed8c5a7ced465fb48d194588d0e1664324836e0b5d2cc1740ade1cd53b47f7d1ba5e0c85a83
z416de79913a86937f4c45434ac9b1bea35d7057948c6455dec41d8088c16bab7e206c9940ad3b3
z2e94f10aabcf93fe99a7e6f494695810ead71e1cd448c41b6e171cfb281995366ba2dfd1046670
z020aed54de255c536dc2d6b5d377e0b5ee9a9e4d934e154ca10e2088acef52d0c6c75936615e80
z80bc42ac8d110457f0bc0dd4c62487e804e3ddf107641376fd3e2b93a89cc0c1f11336e492c8c1
z6cd98f33175f569c40ad07edb205a5ca1b250b830ac7b46ba7e89665376d0e8b3150e10afe1359
z949ca434f09d9a8b23da7638fd71ffb369fda065056d0544b8a389b4399fe8806b0917770f7e59
z869a9ae6cd8c9488647a54deb9b351a1d63110c2325d955963cd503b896df9a1d9892e02aa5119
z2bda161204abd91aa3d080aa6c062a1916ebf64319cbd17fb09efad7edf0f865fca9b4a7588d29
zc856730ad087af0d8f37f1fa5136c10584ca034dc4742e0192230e77ff92a7f14a274f0b481e7e
z7b2b45374d93ca8f6f02d07d1c4d4859b78e863983ea2f28bd0e5f21934f2646d0501e6e6613c5
z9dd25caabd9568e2759984b961442dfb8e6b1afb59de472e18fdfb9dfa1f73e1768b771990439d
za0157d5118dc9e66fce846f1947a925264883059d27780674ddf15464da00355be81ab51cd9ecf
z0c9b7f560ad8e887faaf013670ea8b3770e42dee5e6a94fa83266ede1db1aba54d8beff6fdbaad
z584b90482dbcaf597ffa1678a82296b3842fd593f71abf382a9c5217edbe4276c17876d135c69e
z669d5c6e69a2e2b97beaa7a482a09743b9ac53ca6e77790cb2b8904f42670b320133575c5d0e15
zd24e0b46fa2c0fb7859d022cf6e6207af35a261e3e6976716cb56ba66505ee35c615ada6d75edf
z8a983d93f92f6797088118a19dca947c3bc9b7b8c224726bb268270420bcfcf429007a554c3eb9
z383ba0c92dfb0f2b5022e9f5d61a08f22599f7a6e7135f62e8b76a20a1590c6897c42bfe83d79d
z82f10b4c5b86d6908daf5b390633eb22824da79d53f6eb07682fbf1503fb605d9ce95aef42eeb7
z1ed42265874fbe543afffc91babd68fa26fd3ed786f4d7337d388860899c948145d1abc1986d62
z07b2aa0d56d1e2f79702da37656bcce14aa763d173b7f8c36d143434bed433056812a1ca5b04e5
ze2068319f58fd7fa9aba3a809461cc8066f97294bd3c2e7db213c88f65c36aad802cbe67f945a1
z414ff56e203b22e039de529b8538444904b04bd091981a43f9c3075731a4c450baff769a6774e7
z23659f18225759753d508ff20ca8d6b5f0ebd9fcb4f5f7e985c0f27b2884745a1ec2003ea8c474
z8ab77d4b62040be1d57530dd457c90ede42c6979637645fd51dfd5bc5116b7d45424a7f187751f
z3605f80059fb9e4183ee813f3e36af2cb7f4aff5ec06e6fc0525980d666aaae4346621137d6420
z2fa8efd5bde44e58e1c16db4f670854a174599ebfa8a4b2a8cbd0ef6070ef7dde863af6884fe41
z58e0d1647e0e993f701087e1df6845ae8d9d87ce4414a716f90fe8e1bde6beb03cd0e41c6f00d2
z0114c04f6feb78e5dce24e0e9bce2f9aa9f7e73af2846833728214295e4a93230854b314bbe434
zbd7f1eb92416a41b92751399f19623b9b2edb8a7344220496a546950fc7528decbcefe21872a12
z0f3b4689bebd6d6c79f1eb6569c4dfa0bcb9018dea2dbbfff390cb9367d30fcb699e7c055be945
ze8909fa94fd63f0384fd7d090efa4a304eceda2671d3693a8937f9ef50718a7b12c70443b6d415
zbc4468c3d306065e05eee6ae8f0d9d44f9120da265122dc2b0e5de777a3addda237e2203b357bb
z1e08f5e9b27a6897a448cb54b120a4e99943771fb28a4210c40213cc5b5de4dd71014ab7e78120
zcde7658d01aac61df35bf6552732e4d8deb14cc7ce2af996c5de9e5423d78f08c76e2fbf17b850
zd5f0add22743163697fdf462f7b5d826d8c789722493879b8143f803d602d84b232d7d1b858720
z390e921af3626354d9e04274d286f5287b63c6eab0dd3bc5666c4c6112c3a9657b08d0bb4b0a62
zec3840288825c7e67f60e9694c0e9cbd079466ba77b157edb01aa5c12f8f5826b409f4a918050c
zad0d39d374dc78f02cc14f33bc33b06d37ecb964cfdb4f6e8d7aa781180fd7e80c11b937d9f1aa
zfe06719bd4ab38ace0a06f33c71d989af8e0601bd9347031e651ca69fc4e99c2f3fd3b6490216d
z259771f385d80fa7951499f60443f86537f5a36a98d52b322f94738508773599cca5f2c28692e4
z55fd9cf93e7c791835bb123d7a6c372adb2e6db10f9e5f3a5bec35f529f38f14f2733f5b5c27bb
ze33b2c415a8ec17e98cc58935b5fa437bf7a2c66d0f88ec248a49b16848eaa9d3a7d5b25d2b3d7
zf90281754d271e163e52ae81826570904450bd550bcd26184bef708474bdfdf4e56c94a735f225
zc87b7fed59be4618988558baaec51e2f4202f486a98e98323035b766aa636727cde2064ff0773b
z2642cecb3439af72d9bfa7c1dbc761dad308107705e3c0919110aa034a3ce75e598e2b651ef679
zfd7076a038a2757b979ca361f7a9fee62149cd4fa0336c3949499161a454af19f1877f0764c083
ze0525fe9c70b059e5ce0b6c47e70ab3c0dfc9c998c1b70438a85290771e713e1b89a76a0059429
z93c6441e136c3e6d9277f256b34d70f6a12e2f5963797a752ba5a4d989e18d3be2324dbf3d315d
ze9a9bf55e237eea7f3ca2e22d461312962b6d54d5ce801c3e551777e5bf98d01a01262526a1209
z6ff4861a9ca8993ebe1c6e6fd9ab8d2e9a1295d9e2013e086d82b23facd96f78f6bd9f9a1ecb56
z07a77fcdd6577762a0352e007cc3e3dfdfc6757dd6eaa2097e995ec6adfc0901b50d97df913b2e
zeb547a34c71e784627035072bd7cec37b485a0543e06545490b3fca7772e229a81e1e9565453fd
z40ec31e46ce50a30c19b95c4c2f15e13cfb5fdb59317c9712e15da1f16a2d7fc50ef08eae43d1c
z7924112d43d46c8d573e8bb80fb379dd14112db60a34fbdf509878a1db58313abf212e74881a38
zb8eceba38ed83d4dcaad9388173350ec49b49c68d283eebb13ebce5eab6d5640e584cb8364a59b
z9fdff98ce33c7e26ddd12cbaa5ed654d07052079387401246a4d22416b5e7dfc86a3cf1e5ad7f0
zaee0be87c968ae21c805940dc5c44dc387f4dd57f037a687c5e272155234c762be6a77134c8a44
z3657254da586ad035b7ff0c4a432a92c808256675ac1c8c302675e9fd246985734824773b11d5d
z7612ca7395353fc97a0d1de52059d98d279a270c357a9bba797bbf75fa9037d11047b1cd81866d
z4cc9a85c8f09fb3211a05f3862089a3df0fd4de19fc0f70abffba1c4e828492421712701aedb82
z1b8f0d34864855ac57c0fef0a00e46416806273de056447a95fb077836092fb58d9dca35d056e9
zd3cb5d1879bdedab1c1c85b7c15ba245d8c8558d52810735facd329f009fa07f81ffe0374cde9f
z85e03f2443a3c67356a1bf782ec74803f05d0a9f11563d9055e17f66255b5cb710d43c61793977
z0dca1f7fdf35dd4312ad389abdb8557c045f410936c5cb79741cc14b59287b1289eb192e8db225
z1f234fc49785fd2a01dd6fb56de052b9d6e4f225d878ba9b10161497505f9fed0e7b9c122ecb5c
z63f4a5f66366482982ac93de8de6d1193dbdae2fc1e39a1895fa767b2bd113d73b82f57e5e0145
zdec6a8020a65819f72f6b70c21c4bfb35ca713c5b5fd34dc2b58902759ef405b0b648f33f0597d
z6f07fff007b24cf59cddbf575d26daebf6b2849e3e50bbfea8441e67a24b330ac2c799233bc5d2
za82383f5b018e23ccc7f6fe5f07f3d3da72d468fb33a942a2cd8328d4afe68345dcd9e15e312ee
z68fd405d83d81c8e866859aadd6d9ab45211a3bf24143233d49fb3d195948c4a86372bb3b7c317
zb6033819ad32baf70d05fd3f350df47db2262dbaaf260fd5812617a24675cc161c8c0c8fd8a03f
zc050f1012fd3bc985f426011808fcb1f505359723c0c2d5c4ae513404b2925f3be61cc3fee1a74
zc3a08ad1c09f48048bdb74196d07672c40484f8541c6fb6a80482550ae8308157df5bffd2e589f
z7cd6d255011e39c703b4dd64fd8c92220208798017dc8ff41dc56d909d9581b3ad038be1c0b67a
z326991cf03090b3afe7d6e56d0985a9be3f7c8850afbdd84a93f5ffdf3824bce1b2ebbba9daf7d
z7876e5aa6bdbbc853a6e12c0f40b1e3fc7f91ac5b68ea0bb14bbd8b072404f4f8de9d275bf4147
za9abb389b9bc85c2b7639f2d10d65aaf05d68ff2124bd81eec050b4440339b4b134a3849b150e1
z8c48f3a852ada8bb9b3b6b99bc9dc11eb1b8044d98b3741be3b894dc49934193d488cd57423c53
z15fbf612645199e22f246055d1caf209bd4c9abae04582c11e95f15b9a4f5a8a65b96256a0e64b
zc41fb9abeb085e6f825a0151ee2fde30c1557c0e1dec510417e49a45f9e08374f9baa03faf2ba1
zba4e2f6022b8b4e6369d5eabd00838cef82898c484b10704992705e9b3664cfacd665c11d15196
z4aa88324e0f811261bcf41e9d48b77bf8d9b9b068980bfd9ea47ed9f63ad0f31bce0cdfe105013
zed45ecb380971248b58a01def7e239e1d8fdfb1e5e23e22952275f1915fe824cbd6a5aa6761f05
z0086b9c63ddc661cf18bc2fc2c7305211a93641b8cea97bf15ab7bc6a832dc2d14eeb940b52971
zcc9cc7bf8d9413ac8d45df1b9e080bd1abad67fa73f6450847444022f788159263a5518b62929a
zfd3ccf3dc059c2831c77d87a05cf96c1701d8b03fd0029ca4840ca377c4b1243b277c1eb423af3
zd90845bb5a1aad1253549fe83570e3ef9a2c530c930ebb473ff89d3d1c58fc07da824ffd3e6a58
z05a0937245f6c4fb701d13465445fc138cdde2f3891ed988677a08c32cedd0a300b87f988555a2
z9a1b8ab2bea52c640085bcf41b5e42d1ccdae37ec97295f144e15794c3a9e01023e15956aea5ac
z80f85c79b92e0724be931431d5eb69d4992ab80a156aba4140416ff772086c041aab4c8b80cff4
zb35ca90fc1eec7fbfdcacb44d98d30cfcd64e4fc134e41670e83d60651057d50138ae35c128a9a
z36acbc38cd78162094aff56e4bb226af83065f6edd4f629671a905475d553510aba53b8ba512fa
z0566adda2868ccb9424391f4a78d61d334c82fe5cf05ff524384cdddd49cef91825a3c328e28f6
zaa80525353805e89985f311a642e3071af538a9eb3850f5f602b9dd53881a4286ca3f50c44d2fc
zc62f404b19e1f4f59a68f610809cdc8bb9bfc252e3bd59b7a217dbcfef609d2e27a8de391ee6dd
z0698515b6e61b6104973924b5fa0cd566b829584858fd06c42f21a6b0694f016b679c805f19fd8
za0edc6e6e00bac713f62129a9f5c8c348784ab207264b8d5d5eed46fa31aee43b40b0fdd2c08ce
za4d6ac51d191abb87ef10885886415bc6084df683da24855bfa4555126ef124548ed437b72beed
zab5f2d1f6b3522b2a8c749ad43d6e77033f0ff0051f3805d108b9d755c129934c2035f1eba3314
zcdc24793f364c08e39498fb6e8bab920a8711422cef3bf58ddfd5720247fff0390a68c93fdb1d2
za28cf58ec1c3a1f965becb8e301fad37e2238ba783cb08a32392cfb59c9b18f3e927135cc1f174
ze5554a64ca3a89329dd86a54cbb48dcabe94f042399afddffa51f41336da01ce4ca4450d7f20e8
z0f4878c63cdb16052fcf840853a4c9e67363373799a973d5c61f2d1d4f085c50d05f259de5231e
z2745daaa37d4203519bfd88c3f0e25ec06283058bd9d448477a5787ed4f26fd3f5686f96aa067d
z9290afe90a9c28f5b605b495f3bd52a853cf76a42c672facbced34f9899b48da416b44476ccc2a
z8f3e337af7a0bf078eb4499cb480f8475ad18a5fa8d126dbf80ff01a89f41cf536bf7ef7e7e850
z0936e5502ed119872fba37100ad5a67bf54ac9f359ef0b2f42e3efff8505f4cbfbbf171e782f32
zddd62a8d730f0c220809bf75323c6ba0bc505cbd9479ce51546f1a4c98ec0f9b884b5e7ead7db0
z6cd8096cf80bfeefe600f3490c061f941d90b277f023bbef8446cf8051572ac4384e034a7b3fd6
z08f2ebd1a3c110c18442b35104ea0117260c99edd5174c8f897a634c31bceca042e5ded183fb5d
z473bf1bd8a0b1a2fcd54b64ed9094341f1e9b05229a57aee090418e0362195526eaa0a3d30dd0d
z45f8ceb22e05b84cec589ff0402fb459687197c602ff71747bf86ad0f6815ae24ead0679856bae
zf95fabfe4855e72a4f4614d2aa28561df5d51d84d0928ad466f4c90df2c2b2835c02669c3d8014
z552f23851aca7e519c9098a34c2ff44c07206fabb8281dc14b106c25d1cbc37f8e8fb12f487866
z852712e562d8e7b9c558c3fa0d7506d34cfa015f5f58c90bffe0a7121e0619e1f32c87884bd60f
zbf15bb023d0cea0c4eac1c151c752965e06146f6daa2afed36488a6a652b99198330941550006a
z726e07a422392b540075e95096f948ca4d08a91ffc68445157c5b6c881f66956efe085c97fb6cc
z74f235e0f2acb7ea2ad3d20a1cb7592f00b245ebe4d359cea174a60051074f170578a560b2ccb4
zcbe0a5e504d26431bc72ad8792d116c6a09653e27aa5382952082bdf51feac07d42ea359bbd606
z90e81fa0802aef45dc590eba31cea40f94e64848eeb48418502378d058e1c66adf4461451cccf1
z38e56302b77432c5ff610891081035f4fc983bbe6e0d3bd74b1c9b937d007fba111ce84e8959ea
z8e8f202467d867614654d98846daff650f18adb44d9b8d4e8555e7d3af459ac230435463d99b80
z34b3bcd75e127150d79b90b82bdaa963a1662e34523a8f5433f27a449baadda40072f288fc9d65
z1d38db1775964736ecc67fa9b2e1024a596a2e47b5964b053ff34650db969c66e25c811fb200e9
z8f66e2032f80f4c38ab4beb61023b9ba9476079b92282418bfd10e0d43f7d6d62d5f912ae35602
z5c746b2554a41ec6d274330f2302a40f022d10d34e84e08dd7f2a80e279cf217b854cd9af90a90
zd2e91ad41920743e351668eab5c27aa06523c070f42cac6210e680b9cd6ded993af78ac72e498f
z6a822b13c6f7096e20c7d6e363a5ea1e4d865081f1229e49de1ab5b0e8137ea186ea4041853e75
zda8d24213a1142d6a11de6e2e76c40f8bb5886589b010d2e866c8f20bcd0da855fffd0fe9b4400
z45c34903730e634bf8f0facaf7c2913e5cce1a013c2dfddbffb8ce493700951ca8d47e03bbd53c
zc1350883370c0e233f824f6d0a6b2316c0c4770bbbecfc7121dfb32b86df5c9b64e00d4d8170ba
z36843c8ae5102a352aa1f6b563007facc6fceb4e7b614c3c17eb45d4f51389b31c2befe91d8aa8
z7f160b6ef20a4842e4b563d8f49a3b02475630d98baab411068d6820340a4f414f6ff018279b3e
zdf879825aff1175a3e7d9c225e70ea8a7565d9542205703667d27be50544bf6da8b180e4f67ad6
z5d45edb85178fd9971d1a166a8eb5b3b0c626a592bce5657ec1ffd069a55128a7190615083cead
zd9f5f47be5761b3a609f3086a3ab6666970187ae318543ec03727b6e55e82171ac5ff26e672202
z4b48e5baee2e3948534693ad5c5631a4f8e237c71a9441f9ee32296768763a2396157cc74c794a
z7081618f8f66ee450df7cb8a9e8e497c1c42ae2ad4dfb0bbb2f9b475f50f58d7cf6020b60f0f5d
z7f6956b1c9e0b36004e1b5b71d0bc7cc7842ce131f95f55ea0cf8682a984cb74bfbc7bfde7bbe9
z0dbb93bc097d4243bb2f3e65d8cf0f4a6a6a5b4ff3a4417d4471fafa65fa2f6c915f9ad910dbee
z65111489531c086b36b797f8f8caa2c79d32d21acbccd49c04b5412f6d7872bd3b817c724a6717
z152bfe3b44680f7bdd3004d8828f91cd47c1faeb468374a5c838c30c3233b3da89b96c713da505
zf32f9cc26ddec0492f518852836398983f1ab391b2c3452ba3198d5aaa5cd2a7a9c73a65ec5bb8
z01b830d5687930e77c9423cb3abe8b79d00d212cf0fc9a54db5608e40ba68a0a0bdb6de8190f8f
z4cb80a01be3c9512cb4ef63b88c79ee16887d63a571c7b420a70a208672d117a52896bebe9731e
zfe9deda6f47bd608201f14b09e5c1954c0cbd9c4a2627d62ef482b4cd7fea893f23c2abe30b177
z6e93ee34e4ec9cc1356dac1129ab5e7acf78c8cfc1a2cff2cc911750388f0c9d6f41c206c08dd5
ze16b4dcc5649f7944d74b82ecb248b5c38d16d764edad1690f23be9468ad078ce2cf7542937c2b
zab208430fc9f4dbebb847fef9b44b1ac736c962d458bbc621a58292005ab75bff3a1272a5ffb6d
z6c763e5652888149c8128ede531ef328f52697d1a10dd1b30b3d3b887ce22ea707a4cf9e8a63e5
zc668f206cfeed4e49667a24681c1842e3e9587fe10295ca6c58757790d2aba7698c61213158bc0
zc37c7c8808227890156ad1c5b438bbd87e706362eb9eee1b706933ef4711af2ed25f3277a86b22
z76ccf4a41da9be147235febe1a53ea4fa012e15e99c226dd124404624cdaeb50abd6e3314d7409
zeea7486d72f98e3a048b322f163abdb18463a98f41c0b05b5ac4cf0777349cf7f5534a7c9a50a9
zf2dfcf2d1edade8589bb1d3c2185714e77a95b500a694c5cd7869ebb7097fb828fd6c3bbc663a9
z1280231de19e7051fd5ecdf2d615aa04ff2001f01f07f92070b89527a9304cf9cdfa04936375c7
z10307ee0745d8907f436a451538eacff7a87fe715e8c2e80ff669640c69b8d0614409f76feef0b
z472f69987c3609250e5b75d47452224f5cefa07a3005ac0de563d9fb12466ec8c15b674dd3686d
ze34852855edda8a01a63cd8b740175d2a1d08a98d052339d1358efb006e3307a0db1a73e80049f
z85dfd25d27346a5c64b29177519009a8255e73e93122921be0349177ac0bd8a9b75dc153bb1a62
z5d5f2e6ffc9028023a2774be31c6fbd5ee2b0a2c7ef645723b99771ff7571af6667225afc1d070
z54de5f0f873a5299c960b7a05bd808ae4a5d65a6540adc37c014e5d41946096127e17507e68b0d
z4f9375c071c2c8770a871176b3a29c292d84db8a12936a35e43b551892df9db9ebfde925598337
z219b225b9f1cdca325106ed470571782c206aeaafc1a7dcc06dc9684b7c63fd388cf2039682691
z1214b4a7cc812288f4314d3f4d877d521128421a2149cceea580740fd17e109825b7607564f47f
zb688c67f4d45d36db0505dd1ef2fdc3990d39ae62063f46c26209f35257060920f03030690310e
z9c9e928bd839d043dbdde214d7e11a13d6076c80c68ea2d40d21a1146798ec059684fcba542aff
z895f804561189d2844cd994438a138c5b9e06ebd689ba41d82333e7be51f517e19cb3c56992b8d
z466c2f4dfb1bf88f86c93ad335246ea91ecc7d4c4b4ff77f5990d068add7cc36d731733b3036b0
z2c468db61902fe64392aa5b69363d49d20383f63e4e925f4226fd107790c0daf0284cfde6c8d12
z1c0c3c44d450563965a25ccecdfef0341865dd9ffb34d87d5184bbc83c83b654deb3d0115a20d0
z017535508b5477708afe992dc8179f483b7746b676383dba282887740cba54e56cd18b13a31783
zd46190eb6d8a368d9c5f3f8d3bd7f6e4ef21a04e653fb016c9312fc764e080e0f8b370dd1dab5c
z511cc53ed7c05994837237d3cc5e9b05a87c9f18d0aa56174a489c3598685fab795e427ebcfa0c
z865baba7b5ed21cb73ab9f00226a0935614da2f6bba281d0c031620c0876da1d1a3159e3f24f69
z77b96e6ad2100ce992b049c51eb124796a98633b063dd20c755361f7d356bf2818e051d0d398ce
z044d5c6b4af4aed50257299298c5211d00ec1b3157c12bb27f444e5765daae0799ef085d354608
zbdfe1e919c1729316d3dbf2eee3f7e5a93211718149a6ede03e056dc4832adeac43e59ce9999e9
z239eea6da768ea0671aed827dbb243e9506e1b649399abf3d67196d45e747f2a5e7e52fdcf7fb6
zd929dca2cfcc13d960ca763a1a09d75da35b56dabed34fe2b69a47b32416e88abd8c929326e997
zaf2ae6c677ed54ae4d8587df58646eaad5fea4cea8e21ed33fc7b8c789a00c76dc998d2b2bd08e
ze6e69518aae71dcd4a2ec0d2ca66d12939ee7e5c706d838302aa6ad74279abfb94e7accfdee8a1
zde7e026c23e91f7d0b6165d7577624e308519d6da8b3e3b7a961c61679ccb90026deed653a548b
z26e9e4d5195b7cf2614b26b0cbebdc77f3e947a465ed5aaaf6caaafccaa85fa4d24e3d03e7df57
z2ccd05289eb00956235931f3f31e747eab848a94686dfa0f3efcbea63194644223c9c9309b98b9
z99f0490544d19487824a4cfbf7ac426e7024ff21d8f5e15b28a7ec4f95a4d5532ec1ce66c86c1f
z1a4867569568cf9dc851fb2d927da676cbd8010270d0a58054c3e4d14b9c10e2d88d716431317d
z10aba5326301c4f8219e4d4be86bc9429c15d0f73daff6df9b268a620aba123e837f474ed7f4db
z397a97519a9823cebf93caf462bdabd29559f46e363e643bf198b8a674ddbf3e4d51dbf83ac5ea
z43dcd3af8e85e63d743375922d3b251560e4bc58e67f00731ce4f9230b5b30ab3765c626206e00
z6deb927f2e25a1d3c6411444959e0cf08b125d048d184c49903263f4214566fbcbef119bd28b53
z86b84e928a153273f7e00f9da75e53494f55a8384ac2fb7efcbb56e10f3dc0504378f166a7fcce
z4703b82f337718b0cc5ff84058ca64256f317dc678d6f4154cd8242087cea121b60205ba2ca140
zcc184680aedec99cdf7aca442a6d2c309b2c4dcc3221ab5877cbe8cb876734f8d5879955b82486
z5b7c7640487787b71b913eade2699543feb10094704138693bc227d44c379c898cd2cdbb4e0af5
zfd0bcbe9b3b90267f11188d920fd5926934cc9b2098ba741f117cfded0689c7c937b961485511f
z57a68d0d0dc836f06b154fd82e5ec8ace480055dfe15b41c1d007e03aa93a776d68bb3192a4ba0
z2620a157f13710584479b1713015b6b6658c32c51bc006add73b26af1dfc6371752143b1aff8a7
z21faeeb588a47c1874814815b800329b696ecce70a52f18c33d727a67c8420f237d792e611c835
z7c9fec3ed359e7489c3a9172e3c0b7101756919d51256d92f2f1db32aa64aca286cfa8a19b7b75
z12c78e691e4af4423971099e04e8210719c0d930321b39a2930d6e6a4497bc81da1ea951c57483
zad06cd7189e38831145da22320f093db49764b3f6e8f84b3c0bd6ee8ee5599cfc68ce95e27bff3
z99c3c7f3c3cbf2501c26ada8ea3f15366bf735a911d142420a136077b63e748c5a56f5e8c9399a
za370271bb20a9ff4833fcc6a2e7957cc1329b4df9f7ecaa31da075628b058ba8b31c1abbdb471d
z2eb53102be5e4d319c96646421ae1653239e30567ddb12da6bad2ce3f07a8d43a34c0407eb9ba2
z489d7fc7c90d9dc2da2fde50b06db60913c928caf91f064ec1b77e188407782462441f5717a539
z0a77b766535aed904d4c4a2e9c36d93b51964c2742bacde9b6a3abdef7b231c1d368f06bd321e5
zec1e6768f6d4c19c710a2ebdfaf813cc7a86116a83ae3b223afab9368d7beab6c5edeb8964bec2
z575fcb74773d4663f4480b198e908e42923d3a9de0ceaf2645be9df83f3222c4f83a483d20a220
zd4a674b78affcdd84b97d5649e7537b3bb3faa0bd5ce0e247ebbab0d0c2bbe8d9a8397e82608a3
z50b65ed50f0d508fd90314482d5907f86d1cd2a1eaf35a185ce5b14a6303d04d19ffcc1fc6e919
z8925fda564a5631c2c3a3b0ebf0bcd8f9b84df29c320b555ec2274d0460cb8976e9ae2203c9a96
z03c6db332eb6284a584b816061fd43f7f7e9240511cdbd4791163ea750ef4e448bb13f62996235
z38196f898ad23e7703fa275652f26990336ddac40b457a0c8dc47915ba383e47363d7c2dd8d5cf
z80d54796d0021be3744b30d01d906c6b7ad7b18fd862fb3ae2957490dc0dcdf5838f8f613f88ee
z4156684e603182028808ed1ac9692551f6ee50e98904f352b6650994de5b0305649679b34adfe1
zd6a21c29d2b4398749a61f52b99815bbc7cf38d45d1cb7c91003c652692d5a353dd7a43e019d7b
z45f4dce928cddef9f924057cad78613631d68f76dbc3ac661848590eaf765440793de67eabccec
zc423fda7fa8c130682357a8b918fcf2526a8e4317e8ebe77425d73263818f585f2d4079345519f
zdf6b02ebc7751f9929610f18fc9c4c7e57e5262444fcf6a08cb3b33d1f679f8e5f3a129011a020
z13878f363ecfa255b94d4186499f8b4e5149cafe6873c5e1a557bc0d6c9cacfbacce4838285f40
zd18c71af1acfc0d4d77f1ce90f8bb46958c07dc20f634cc80686f1409a7e9f3c5752577d309f0b
zad0c289f4cd4e5ad276596db326333dc42028e2fa66b7bbef0066ee3b7b0444bcf66e43a3b79a9
zafb5b19d7279c53c7f7694c079e1039f25f7478da95791e491959567c6537b57912df28dd945e6
zb1f976a46886343f26c835095d26962ee6f835879079c1a64b12aece807b6ae4a3a2faedb23fe4
z888f2a7b0b881000c1c1874ce40cae94006c1db0d636dacdf873000ee1bee429ef2a5a82b9dbb2
z2f050a1fd107e07ff3b827a662fbf7f7f24269a6f7f93ae71da4c11899f43cf984f7be04745cc2
z2e034d0c556494abd6436c69acc091a9433c843b44cdc0b8509b7a6818a5e2d74edf160c66e64c
ze073866b8316435a009fa49b23aa8edbecca98adc61302fd5c6eafe50c6777da1f1bd516a5becb
z0fe06bba7faa604069d4ea4bc21b2027348e2e148609b174ff278a41c708b5fccc34792b4b1339
z105d0ad1a8490fbbde9a7ff4060fecbc053ecb875c85c6ccd7b0bff06f2614eefac026d48cc0e3
z529191a4728d09625e8429b32a36675a5d19329d970d70ea5d7656aa24eea361987705e5766ed5
z13684592ec743e236cfd9c29e1b87ec02068fc66aaef4243eb978602731be8f945cac528f98be9
z9bcf04a4f57451bef706c8db5b0176f349f44aed15aa1021d14cc6b8482feba6df7ef3b4a1de6e
zd3b6cf2cb2f89246ce87c6ec6e71b85f6c05c52a0aff38e87549f9deab28046c016b420b76251b
z39f80fc36e0617a91adcfec743de72c61eae125dc072df85bcd6b107f19bc6e45ca849463129ee
ze764380fcc8dfffbbaf5bcd0977c0046c03421ef97567731e1316cc8ea90a6b38634c583b6742f
z92d3950ea1d2f9c42205a79e1440fb95bd4bb2d52fe9a904148170f5f6bf166049cfe30f3ffbd4
za24ba75bc88dcf1d57f891689bc8c6bf80ea69f5f3f71d7702355163313d51777066f7b215a71b
zc37b53792768a2b57a5c3f01a281ba319248f7bccc022d5be4ffd72a8d6d670d03f2004799d5de
z2c4e202d2e648c0877dae472ce3cb1d37ec9c38fbe21e28e3be70f48b403b494da0f672d87d22b
z2d32d9b01925bb6124403ea6b139a0340bae5c0b9678d3d4c8f2a72d6831006b218cb23dd0003a
z06a8baeca45987181cc00c3e9091aa68195b5bc7fe516f9277b66c95b45ac4bbb04d90a1e4c3ab
z2ac458b545a7ac8b472a0c4f6c682be3ab20a2b34c212966fbbb1384d03db1b9efd8550c3b79a3
ze6f7430a5ef34dbcd2320bf855b45699c0caedd52246d246c28806af6ade72fbe235cda81ec935
zf34eec0f55de009f67ce048b3af56703b4f2daaf21e76c2bebc35c1434c62f826e96c6570b17b8
z6df8c209b423d6b40a7230529370679d80580e19a614bca1397f6b18aaf2bff2299b329a93c986
zacf900356e25f8b2ea08ac3d14d2460255d1910566d0b6ea713afbeadf308363dde6906c7fd577
ze93fac578e898f166162ce4e12a7b375ad5ccb0276dd03e94f8196f606c9de5915c9cc9b33f750
zdecffa6521755d6b9e1f32953801b46f42eae8af284e8a1aa3110115c4a865a8a7854c25bbeffc
zceaf6629a68b0b1d126dc087e6b137c329d833785cb71f455458abef97783189ff0d9726846e78
zed6efe54f019632fb3e52c0de7127fa6f2ffc74e107f91a4d291295762b8a8f1e46ffda07fe659
z97c2136d9ed2cdbf357b35e5eedf750c03549518df31583a6e17bd57cf2738947a862c453016b4
zeb70d99196d7bc5e9708288206f9ebeea2531e1846267f5b682ef4019bbb07b91025cbb5e84e2a
z137302d5d7907a7676c5d8f417d3eaa27b8a4297de9ca9b65f295842b1324a3b6b0e80565e0f2f
z1c0f82ce29c98c90ac2802899dabacb565c78f595350ff670736f432496dc6061c07a12f3549d6
z7205c54074ac94c6197d666b72c4a91815fdc502840142056fe39306d4026c81190e108d5ef51d
z3a29e2f048e9e2d02650aaab03de4016bf889d74606a4478f90691cd7c2a3c77132d20399032da
zb821e2f3afde1a4c1abfb702e4a6041e52ce382651dd325980910385464f12c3d7c1fbb6460823
z45a1a6b93aae617b7aae9028fa802d74e43c2290dbf2745c31a46bba83f27fb06f81604cf31988
z861c86e7b68d985765cbc90e6fe179a2ccba45a976e37cfeab62385f51db79254bc5ff4cb16123
z9a4a74edb9e49a3e8d997fc18ff39665c47df3d8c724d7047e818574d209faf68467f73ffd16d7
z7bf5db08d56760e9617031b60683bc0797e6f7989037d1a200cbf21172ee1a3c44735a2a623f1b
z41913f721ea30644220dcb280e376f64d52ebbe5b56293e2780e1ac534c6b1263f9db3c4ec2689
z698124fdd69793d1dff10ff0a9b1c1d386e372adc9ffdf4e93c62cf704a9da00e709acd6a101bc
z0b7ea975453861ef5f1365b37ad6fa4bcad308fd635ce57448d89afd864877582d8b14afe96ef4
z5d9bde9b3e39002a29442e3192e6e3a42e90a107f632335c68bc9cd3de6ec900b7abf4754434bd
z550364ecdd80bb6b9bbb4461666bad7cfeadf493f862be58e24c261f1e1a394ba5aa7a47d429de
z9f37f9555aa2c6f3e7f4aa1cde3fc8f03fd3e0147e9cb81ba5a10c50faac0104022991d9f58f37
z29dc462772b8fa757faf1b6885e535d817f4f6bf17b2165b024e44a2e0bf4df88269c44b140d1b
z91e04db24a945f02dbdd8ec660c3b51ea4b43e27bf4386d6e64794689cd5e3cb2ab563a12e9668
z9c1340148bc2d439381f28a5d67c23326461b17df77ca644537f84a02473cb9016c6f27399dacb
z19f7a29fed460f0a75439dcf09104a2ade650afa331a8aa2a081d9002cf4495113e034c2beca3b
z2bc07ca03be88fe65aca95f2e54377b1b3d9646ae0f9528b7073eb32e1f3a63383127d670db786
z8372d0aae1877c4f109422ee74a46a94c25f6d427c6a435239b07cc8b6c985d4296969ad3f42d5
z35723b43db05419ba90232879da5ca28d5ef0807bea79eb142f57bfb602df848c0d00d9f3fd036
ze95f1e24750662980de2c24680f9433c98bc312d6da33e95c6b73305ee85144a5897d85f3632fa
z1297a932596a9d5fc73d3cb5d206403cea93df07239de736df4c001cdb647bc7e7b61727a10f61
zd2b124b420b5e307ed33fab99332260df426b63784c928c438ac815c06c2c1862bb2b2bf1d2310
z7c17c43ba8ee8a5cc5503356a391d1db348995d2be12a142e870720aa7362146e6fe9d865002f1
z8ef4c7d01b0e96325a7220abef1119f945adeb1ee51838c44dea0eb7386924403ed62e9c474ab9
zb85d909344770a9f3d1cddc650d5d659b7d6cce1fdd8f0c173c682c609feb13e0b0a771f396ac0
z82fa478f22cd11d4e5647df78f5302554ca5dd9c49b83d51c8a11dc3b82f6411c421f0e239bb42
z04bd6c78bb8bef7f79f105825d39ce967b8d36e5b8e4edca32ffb75d0e9b102d38d65aa6edecea
za69fbcd6299796687b415666d352a5412370174b260ac9733a8578fc0035e4a1781538d2c8acb0
z66458f106021bdb18518c270262d45feda42b907253388d74e064a8fba9a3447d4b3564d64ad7d
ze867b42d0c3a916960457031ada73b4a0a64aa993c88e59a4e59c8452f45bd9ed2173bc91c49ff
zb03bf84f30bd226ae0ce325ede3ace61101da911e773d5f1d327b89cd19b9272ae3ea4615f7aeb
z7f59484447e0dc54917efe5846c02c46d9ea60e04b06227d58e073708d2870e0f576497db64b19
z89e5dd6bca8e314e516e432ce54ae983c664c98c729cef67318f921483c62b164127676684448c
z025109de954fc01ea5670a02e52803b841ffd05cc9df2eeb4e998f7935d8bb979b739ddb0894d8
zb3ecf46835f9ab230b1212b86729418ab1f5fbcad1078beefb8846aca02fcb97c59285e09b6cea
z00f68e49a00c9ac36be27e835aaa168dbd8a804cf948aaf4eb1ba6aef5227c60ef88a438cc5006
z638d615499052ef964fcc65e92c7218725469a704311fc0b45465ba1edd1fa12a45e537f978bda
zed2b665f268f07960f52945ce5993da7fb5fb5fd7fb126d6d61962d07df68fc7abf7d7d13f8588
z0af16a6dd07fb278869ec5974b24c48c5df13f2b33b15aaf3a955cef6b3502432b14b82b1b3dcc
z6881a44dcd32b0a843ad28b62fcbec6f62c800dba8df0d92cea9c30a0c77bb16cbd39fe8d22d49
z5603ff05815d16a3a30bfd1ffbd66a1d872a3f7397b60c4107a477d35df7258a8431b657615756
zfe43f634e30cba46c5ce6ba193855e7cd43001805af7515bfed97519c1188ba7f2dddfbc314fec
z3708b9963c9fdeddb4760a6ebf2cfd55c2e2253a77f7d7a581bf5b7d80a8c687e400f4e53ef2f9
z01122b3447314189e360776014169957a6e94062a950060a2c9fde57124072bac5a74ec9b8782f
zf526ebf198f3ae87292a04100b98f9e8103de257c12226afb98771c0e1403dece329b296b24892
z1e65e427005ae811dd28bb5f856db7a04e994817aab8a2c06324ba234afe127ae344d6d1a10614
zda86dfca868e766389521ee06c7721bf602f309e24e23c6d61aca54f52fc01bf33e584081eb8a8
z5606f5b240a7399ad169f3e091ab34150ceaec0bb2922236717790167f206faa3b930a065f6510
z10d10cf738842cbf9ebdf6e3a50b262685505d4a3bd31ffb6a4515235e157ee932f88c889ee236
z4f01ad8bd2d82151d3534529a604e06891297e2f857ea3cffa9700014318eb2bd655ec58f3f2e9
zf9929fc5047752bc12e4d654a7f4b1a77d864102020fb6ce3d7f043b5a1a146b4a667d8c0988b0
ze90dc7bf28ef7e498db416ccda6779fb7f9653572823ca1acf2a2fe09dfc9c9f7eb85d9bcc8179
zc7aae72698af8de393ca51785565e615e326b4778e054f37fac2a97aa8a79934aa01795c90c752
z92a3563f1b478e8ceaf9bc1b13852bb6a7485c765611b8de3ba74c295a883f4b409aa61d601f61
z563d696c6ec9896a975d0eb781e0b1179eceaefd5840cabe263a6b1ceb98a762b6adf1b4c18743
z5139741190204a226411f9dca3b6bcb9960c6ae34c8cf45bc0cfe708a184d81a0a27df7ea1911d
zd45df1162340f17e57154b76aec2e2c08308b3434df9804ec582d093c739da35e53eb877feb80b
z25fba696c964e79d83d807246921eea6624d8061089d5f60faa713b407c1526b81194a90928f29
ze3eb1d3734e44c8bf2df4ff8c3a1af9b896a7a108b321485ffed92fdab26683348d7efe20b7760
z55f27a7d4ffa4eb51e6306dbfdae3a0294d7b5f7c1d25e1a1d04a058d2e837384e4ed94570ba10
zb8a27e5d458b10a7e4a211a441bb5213421db9125eb8ccf825bbe28e8ce3b245d1bc1a5515dabb
z477f51f8bd5a11785c86216be38ce0b7a3ee74b594ef07be6c3b69bc55b3847136efbeec5907cd
z7ca401d74b06b0b2c9ad2ed8de07f55f7479ec594ec697c09fbab64f30e129fdec420e3d1fa22e
z5055426d9d8f1bd604c92431ebebe36ebc7efacfd86330ba6572fd639dc7b99238c6de4664ee6a
z8e2b937c5533939c5d77da827fa0ce217c2d5ec38728c74acd77789592a6e68b59a42a06c5111c
z63d898b73b4976f4604ae537c39d0a05675b6286ddcacef36994a93b092a3fcbb9600701b560fc
zcec949b6b77de5f4020355141700b6a8230324965532ef1531eaf498cd671a4f6664c7dc035d2e
z51c663f3f3206a6635d593e5299ba0702cc746fd12befbc40e577466bddc0670fb475217b3bb09
z07c3b6498e077c6e1512474feaa99c0be2446e894f45ed17a5cb4e7d7f938cfc28926de4612154
ze9e117136d93c51c3aaa413a5d3991a6756319b14c09ec94c23678e9113f1cc81c0244301cca5c
z8cc4de9969409c07a7cf1577ba9dc9c35d52fb37e62ac85603c8bb9d3ef46575b214cd06eb97be
zca69f0484590a5bbf9bfde5156bcae663bb17097fee3b751adad4abd4be0efc52b30687b34f220
z983010eee195865466e90522a082306b4f763356fbadba0f4b689352ea92415888b5734dafeb60
z762c19ff854ac6eb467a62b853f073af8ae129883d591c1ff7b396b2cfa5c8d9c044d345ed7f8f
z0e7912d4e2c58f069f6183a4da3132b00e9b54778ae4fc3dd42fe6bfd4685314a92bcc8805f354
zca71043d746e2e8d9077f4a5da9e08cd01c95bcd99f00854b41b6701b25ac99237938967f03d98
z87ee8a616f6e03a8d170e36ed261f1c226d3e7bf019c0d534e6d16b6a81a5bf508b64b7725467d
zec621e5a810e8f34a767f5e389863574491df08f815317ee4e2c556bfd82bc72493679753a8d9c
zf972a6dd69b6a928ad2a232ab29d8d5e54ad3eed98b2201e8f4282409eade129e360fda7a6b421
z4371e752c06c8ed4049ee1971e2d7072ed02982ca1ba73d2d94cfb1ba4925b6e3fa6d46344badf
zf7573fcd72439e169d2b3d6e76416af40f3b073668785ddf813e4f59325b5484b414d5a3e74294
z7449a73c1bdd1f244c2ecc6198581e3d265325d67febd49cbeb53f8555971ee68179c1f3d610f2
z7390cea0ffe0963e2985890ceff010ac1a6c11a94cef07bc866d69860a033cccd6f6e99b2d88c2
z454cc0a6045d90f2e3f7c6d28e57216f29358b1b4f6cbc02e4318edb46cfe0ec232ff1a8a671cd
z11a462877ebe5f9a0e53d79f1c21c9319e55cb46b2f1ce672931ad6bfe9407c28644c7f760bda8
z3b4c00cd205a8a801b0e1bc71cbe9a9197761caa7db7925a4c2b1fc9b3322b7073ba1cc9bf41ef
z955725607f256ff734b049e0f157dfd90a572102e6a2c51bb660736d755e1f14df7904421d0636
zbf52b2955ca46ab566bb0cf8e3ac997ae43d5286b893d84ba54aa51eb2cd9c5cd7bce3d862e843
zd0c90ac3ee7844a90413b95670eb2fa31fff2e8de28245bd1788ad18d24cce84f56d6081ba9f32
zeb928edf7113ab4af78cfee57aed2957c743929b531252fbee55c6c6829340076c495b589f97b5
z80faf836363904bd9ac8571721dd5561f791a103e942dda50591039a9ad1efc39e581e048d988f
zfc63c85c49a5b972870c62fb08aba2f2720fbadeef618fb8f54bb1b0c4789c0daff5b8c53babd2
z11da8b407dcebdce7ef1dd474a56b8494097b4e206c0b0806c12e2d7a9d7ea5eff4505800c44c6
z58abcb1dd1eed3a7b5f50ffabcc9b3e0fceb70aba4e30291061c3776a427a87199bd5deddfaf59
zc8af62fcf2bc1583e89e7051c2ce871583c7a4655a90ca8f85ab7d9b398fb2edcacfe1d7da77ba
z75f5a472662040567e7b73e2937ef7bcb56f161a345367c27d855b6c06dc0e282641ba652709d5
z1bb98fbad946b36da3f591c9660c4630416960ff1e81deab8f2e488e5ca9c5cebbd8c13cebb28f
zd98adbb0f96fb766bf5102e28c5b2038d177027f853f09be7ff13df988066a3e791f9b3109e312
z768447b50847df198301f6eec1b1374e4197ea0c6cb2701746d3530a7f77c5ca45dc419e03caf5
z72c6569fe0ad038cd8fc8b5ff3dfce6aaa741ed7edf61df1e12f01eee8a0a60b225d27f063fd7a
zcd1666bff0810372571d7b31d66a4ce55e917d864ad68fe7edbe15c789ed7a3cdda50668b5c803
z84ba9685ab52702ca68c0a7b75def8baa5a1ad8cb57e00eae78f12c378e67d31253af0b9108200
ze7d4d334bc359ffb6dca9131312d30c388551fa093ed8424ee6da1c0f5768cb45a1c2a033d0228
z2e8890e42617a9f1a02910f8197cffbbd3cc899c24f03a822998c5399c1a688256b3dc1c75669a
zc00000f87f1d204a81365645a3b1c36076479c7183ae26e87c662894046ba2bee7158a494cc719
zcfce454422930d8d535ef2f9468a68cf1f9201a23d10176c62c02cb8d4a157a79c902abfe7d5ad
ze2c3008e93422d12cdf1247757d1a1d18c89e054621c9d8cfde2c0b26392763a77fe9ba9921427
zeb4de131c55e9f04eaab45470ab40581f5fe9085de796c866f2636fdd255c5367c1b783a7136ef
z24b270dccf3af833f80102ef6cc040541ff738078fb82f4b2f79f1e4c22398c87023fb357e031c
zd9e46ab13f7add5d47cc29f12642917137ac90a38c40811d6316802e2217aa80385fe539a598b0
za89cf49500793e18b28a32a3748f45ab6e542b63c13254ebf541e9645b9271dc93ea7804ef99e7
z8c16803cae534b682132191540e8b644a4f886df25534af70b157e619d6ef42da51efb8967236d
zc38f6d30c2829f558963ff88fdca9298947816b4139790d7828af7c89eb7c014d1e398f23ff5c7
ze3ea47a13c08f6225a810967a238baa0c314accb3cb865dce7343e631904965bb5c578a5d00e78
zc03f863811201899fb56d0d306c64820d1fe1074807fcb5af1ca1c57d7285e7b6887040a40ef8d
z1b9b306dcec7eb26e2eefb6b262e208114b16140efea602bf2762ab9330d6f8799d87ec79946bd
z874a5585d0c2e1fa283706724ce6650ba6c009fae472f4b3bc92aee4a607c958c7b62e5eb27cda
zc9774bf3a427d7dd8121a7c487b975fd276b25859d8e2506d12b54c23d7735dd8d516d5fd2f6c0
z5b8f637aac07cffb9fa81a19db7f51136b78e55fbb49f89e8334d22a3d19e728bf51505677dde6
z03d2cd9f226f34f06ac21f33668c7b7e0b005144eb116b4100603bc91485a48183377892e61e5d
zdc205a338fd2d42e8cacfc86594316ea2e595574a341aeb4b1927605652d140b03a823f6b4bd1c
zb471b0bb5a69c4429db4d813d54d3e5f8ec9b1513a139af06ab568650af1c91da3ea259416a532
z18809d6dfd03383e7b2a05022a681bedcfcfb9af564e04b578f8a93693526b017a82fae493061e
z59e428b821bfc51f97ede33ff1fefdbeaeca5bb979a11f61d3fdaa8c7381aa75cfa1ff51f16a0d
zd4f125de328f88cbcacd2d540854c36dd4fef4b6d7962675cdbf0c120182195996d5c8581195af
zfd1e2d1f678e31b3cbb77216e2211b1d560e18e0d23034c91769675ce8196287f73484ba4d20bb
zab3ef5b0863f130810e29c2581ea7587359713b486b0867d0f80f50daac2426097f6e432d6702a
z98ff17ea365dbad3ec686049ec8f1af94f6ad96f2f94ec9b92537912f486586f82dc2c7efa32bb
z6f10c98b6de2b0a2e2c72dd913bca5cdd34f4cc2255773608d4ca0875fb1c1c20377f566ab8c81
zc2308bd3a6cbee88fa36d696994058fe166d68e218c9c2d13b5270296c0ce6412e2a0f0f7d2da1
z73b5138fcc8ba1cc3a8adda4a17dced959b3939adc9046e03546a3a2eaaef9e8dfc6194831ccaa
z851c25c2d241818173d8e0d99d09aaf0690cccff257ae81f6aade8cb64a2204dae2e7ca3896a65
zb4adc31b9a17cecbd4ae65226bbed32c6989dac8885538302c4fea84e2c22a4222230f55558e52
z26a45dcab2add99a99e6aeae4d0c8c9bf19a66d2a75a780ccb187f1a3bab14275c271346d66a83
z6823008986932313918ece9db62f3b39dea43d04caaeb9bb048f7e9c5fda68afbdb319d00c3484
z83293c02f073a0fc82694b785fa54d34e7e44da21ef10a3ad484b32521488ce8361b07585c1b50
z088729c6b2e485f537a92302056c062272571e276bf59944e9b2a8bbcce9dab1ed10c757dee22f
zdbb700f8e2dd3d94b9770ab7f77bb3d27e1b01e8c1ed6a39fcd04bd1b0d3f540c2804220825139
z97280a849b5d1ecee9a19db0c1ce2f05d4400579472e163849b07c8d146ca685b2d5854b7591fd
z86e0ec3053171242db26886e50adf0dc6f260212f60248b3c968e571c23d8f76e410d178e6498d
z73c6e2aabc609e2003dcd210ba1b36c3820bedfec31fd03d9477d205cf1edb865912f5ee609bbc
zb79235d110dfb7ca813a8bd81dc56094e2729277ec1bd59780d4f6c0ce6b5127dce1956cb0da1c
zcc98381ff265000813ca929ef8b15897297f2426a78bf1d22095b970025ebddfff002addc40d63
z74b1bd866661787691c32e664be42dfbe15fa30e0651e5bf354a79808fa6a0ff00823b731e946e
z1335f60328840e669e91361971110a95853c38e50da446b2e99ad31a4cfc0b77de21b33f66d5a0
z1acb13175d6a1889d5928b5a63b996f53ed8426307c86011b4758ccab6535e5be26750b3c4611e
z9e8f370d3c3fc2a611ac687cd2fe9f63999de3ef71a428f5e112d25d23925fac0182a398dbce1e
z881af4231afec427a5298ddb841c0d3484f301c163c0a9a1e9c32cc44f3b5cac3916e4ab6c0788
z4863a522b9399a446c78d46381cdfc0ed5d0a5cf653ab6561d9d02b12357300823c27c0806e83f
zc423bbb89a9f25b4d949619c0748e41e9f9cf36ce8792edad4b5fb865f7d5a42958cb7a30037ff
z194070252ea1ad62adabf3d1763625bcbfbfc70efb9eff51ed32543e7636cd4ced67cbed1f21cb
zede5af6cdbfc5a3740232f293b5be85e3ac66904181b6a7baeb3d726ec20620ee998c99503725b
zac7af8ba5f2ad6cc1c28b818ef70c26f2c890b3953ca0a65f2ee5f9a8a8066fb1fad4718f871ba
ze0b876f3b7758592e05bc72e9962badcff61161d83f83074d6ef71d60724ec34c39f6aff65a6d7
z21a00dde41de8250a6bb7b370f239a7284908f22ce3c2e72cb3a0db2d1765571c29279552c4652
z2048ccf18be047c1651f74d862e63ee38409367222b0c38a61a4da80158c2818ca39ac44c5e2c4
z650f73551a5268cd7d5b13ed47170395e60143667365c3644d1e9a8972b1d0ea0acf835c0f85a2
z8d51c0ffe5410ee2cb08ba3e2473d6e53295931ab19a3d437a5df68014ffc29bfb37688a61c4ee
z6e2c8cef036a3f7d92b565159830cd083509809f8d407f09baae3b91818619f150babf2d209c51
z2680df12f120c7939d2f83178057fccd33037081782cecb8d508c297d2180def2671cc128a60b6
z92453dbc4a1e8181ec04a29b867a4074f80f8d006153d081d7dcd35a9b4989d4255cdb70f0fc2c
z56e3bd66fd7b77dc8d1c3497b74efb8eeb98a43444d7c2bbfc21170544bfef05a4db60ea262796
z8d4502372547fd1ac3c72b533b80a98913e72ce4eb76b89e39dbb83a2b606685e7fe509e1619c7
z2104ec5c8a443bdc37de256d72c8fe087481f7f9f478957fa104fcc7af04c5912467ab8c2238c7
za5d08cc953dae6ce2d90f90b24d222f73ab0fcd1e713aa79458dbd00b94d20af0acc24c313da9e
z8d8ae69704a97e13a93ba4dc31d1a646100859c4db0414ac24c0d854ff53a4df039f802557d3e8
z5dfc31829731828543183184e1e919ef26dc26d0b00977be03e91a483af5a43bbd7135b9e813e1
z075b0fee0f829d88b8296460889debb34f01dc55ea9a8647a3b1df66699249ea3f46be90b54669
zc3ac5b457ac69ac9edc0433815b24b1c75fdb5acdb9775246d41305b3c986c052d0e96a6871d16
z0d117af8cc2ecf304be9e0e3571a57b0746c61b0651af83e67466d501de1ea8d36483ce8ecc051
z7aa71557286bb423876a27d0e13c2426de18a62ad488db5679e25418cf6721c685ff07f093274d
z345bb3d98c1b84db0a6e6407066cbb562aa12a1cac67b68c3cd97e8f0d08e26ba378645a9ed9d2
z6370f458fcd3127e291bc3595309a38353fff140b9849c64ba54a36338da4189be4ed600e9a77a
zf608f0a524bf3a8b1858cd733519866acf2b6ba185ccf470490088abc8b4148119d4ab2df7d4e4
zaae70ed5a625ada92bc1bdfaebb65b81dbbc355e0d2a01d0af44a82a9dfd7a20f6732cb3ddbf29
z2a17cf4c2bbaa8952795561ec017c7018ed6b78b077abb2397546209cdb25e99d982bcc1eda778
z573e89e0e56978f0b667cd564a76994428c629571dd283b66488c3f4f8a9fc2abbad7076a0a5a7
z285951e5796a4c869c75b8723bf8bff93a22097dff68c11145dca7b53105c7a63a6aaf8c73bbf1
z800a8260c5218d40c79c89c401a6edb13d1ff2faa571b8c467b9ebe0e01429c976994ac76df926
z1d3fcd7d47dac51fc2de758030782381dfb9523841814d2e9ff82c4296d1beeb5ff79f873319d7
zf54fd466f5b8c98f25b628d623a92da7c93f0a0c5751b59acf6296806d7cb3fa203c02c5bfa1fe
zb97b6d4ffadac8a84d7f2e520ac41383d8ddff2b3b24b884d78b7b7b17a39576a2c383316aff15
z685b4a630aa0abaa4e495564cc6fcea505ea56054b1b06411ceb9648efd1b3bfebaa2e2a4b8782
ze1cbb64424ede492eaae1d3c941bb5e463381e8a0d3278659ae828ee01ce89fb784814e338c2ba
z20125d7faaebf275793bef2cd870fb9b6e32d78c1c659f40d072ede8630996566a24a87f94120b
z8d5f2f2a85f45ef417a5ac68e522e6f0d09271d1085bca5592d5f9934c9ff5319873180613144b
z7954611a79159c53ff94c9adc876e1df1a80de3dc9fde6b02dc06530f7ef02294b9e5a9a0bf271
z309ef0cd9a79f7ce9dbb6e16cde18e01ec959a37be50db7128dfbb122c6b59c42657c4d6300e93
z47015197adaffc0e69ddf1537186676aaa5da6a9570e68e55a8d5f322663c78ac6dc9fd9cdd36c
z98e2fedd5415125fcedbf3b52658e33d8c9d092170f283b5251e068487b3e687c79cdd4976d071
z33e6eaba38c4520a20406bac2bd37a7f7f13c82b20fccaa322e760ec042ecee8339d3f609283a7
zf358d3a2bcd97d284ae569f3d77848c659df87bada667d6f16a253d2b752af0bcc0b6f9ff8a9e3
z3dc6e1aeab7f35edbcc10b5f377b7f62f8575eb2ad30fe09502426340d0aa92ed445bef08de537
z4d687146a746b885f4a7992b0c448baeff3b77f68c5ccefa206ad3ab9e0070c2f19b6977dc78ec
z1a930f1071d5a7048c4188c52cc1b01801ee08cc2892bb9de45890ae4464262d632b657a1f3f06
zebeaa18420f89769841aaf383ef18d4f4bd8e5e5bfc70a4f8f2dbab5e16f82d7b70492339be93d
z93bf868734b1181e285830b47f4a839e568b05248ffd1903caca2ff2fdcddcfe1c735c913eb453
z914b9b94fbee9efd32c96daa5643062a25d53fb76ebbe9687c2ba7a5c87f1c6134e645f246b4cb
zf6a3ae80ac3ddfe448e25daa5507c8a38535569d11fb41bf1d00e1e5e2dcf77807da853e531338
z560707a2966c7056367f53238bfaf526e52515a954ab4ebd8f8a48e4545468405b50aa28e4c283
zd1ba8a4b853da47e80de3f9e0f90c1e13a70e9577bf8c00dded0374e8383ab5756bc8acf428b6c
zec1ca8a519e9be204ae7c4a7f3bb4fddf440dc93aa60647c31bd61efc13e567825ed76a5bed5af
z375db8805d84d8e9da4c50b96d14aebb4c2af54571cc11af4a3eee8413752bf16dd41c44105fb4
z58e1dac8b2d30ee777d4962e8ee6e2d71e60785236df9c9dd34c5c5c08102b968fb499bfd3e70e
z0ce66aa6134f6695a713e038e4cd55edd77121b079c87ea2704bd5ce4fd4e4c0f2bea88cdaf18b
z60a2f08269cfe929866dacab619bc3f4490955fe1d77679869b04fae799b613055fa985c83a585
z084ed7612033e0a54341b99e704fac270f8249d564be86e4f85dea108c8ed1d80b4520c0d4a76a
z47c8624d803fcd5926add9dea796e7463f43d6ead21e97564c91cd5740bbefb9b7d1fee5699218
z00a6d7f4880de36c9ac1904bdd666c78b6bc43e8ac049519189b12ec78f09a0614d0b62e592dd1
za265ba2901dee3c53956f7de5f06c79b2dca3a5e2a6a00670e0b8c3cd3ef5c775264ff2cec4082
z0b8a016f68a3c82b0f0c31f61621a99aac786b09f5971cffb3df29c798660da16a281686602e03
zcc298c4a0137a40935842c17cd43efc0ef5e2fe23cc78e9b9fd5181ab871f2c28e6c4e8dbafcab
z483f15592bcf24c44173535205804c98906201d98b6e6c91ad2a5558f2f77c2ee37315ec80d4a3
zfe83fcfd494cfa92fded85e51d36fd94087ac110798aca1b589b717c3c3ecf87bae5cd72644007
z093defa15c6ad5063e4c6be4af80aa25bd96a85270dab24fb9245dae9dc11c3a95e60018c432fc
za2f5eee24372f38ff4938ea966fe5140c78fe4245217425212a1420146b0e3aba8b09f9c217e2c
z7a97270bc5df3994f3f9746e74edf44a77d0de453ecf4cc04d7a1e0b55cf27e5eb75c186d86909
z6dfe981c8c5c3b634172e00212ae4b9fe56cb0d895bb7161af7fbecb4fc5fca6f115fac4de5c00
z4608a6dd403b2031c8f33500d804cb6355e30610eecd0534176efa3dce3a38468eae64fe3198fa
z4b35db19aa67e9c42064bba4203365fd9e1dd453b37741cfefe1eaa8c2196debe691fa33929988
z786295c6f400b294238566a9b92a065e5038a0edd16a258375608278986a81c1537d747ae61946
zeb393d6c151952103ef21efe752b540fa48db5937013085e3d55c4f5e48c5a1137dce02db0a540
z8f0a332afaa6dd77ee89ce9ec349a63bc8b82e8c0e49be25ddcc7d346543cd1d5ebfe495c931c2
zf8a0ad97c88feece0af1eb8de2eb0e30e9531f35df896064be80bcdcf65d3db495677372791ed6
zcf27cdc1cf0554751bb02ca9d4e882f3c59313c9f1bfa70404e3a8a39c3be82a62d9a8fc21e7b2
z80ca9379a35b87c5b3643dc9ee6cc922579e5ec91423cd198f910e350667350b184de8a4ed2d48
z9fd60ce8f6003b0cef60af65b1adcf4e857bf5a591ae7033a1203c16619287303ed5d3a3538304
zf2798ee20f77b7db184740f7762cdcbfa35399b987696c0f197decb0ed083938d69e254ab94e71
z5d9e96da93df56fb3a1641cfd11019e755e35da18770ed51c73f99552d2518dd00b23e8596e395
z1c0c3619e7600183691128b15de3a74306d4d535cd52624496be83d086ba815b99972cb3c1daa3
z2f28caa1294daa087e082ec1251e2570441bfe9e47194d5735314034e590b997adb8bb5ec20c6f
z2762d5f1bcbfba7fea168166775939eec19dea33e4c970487983b35e58204a3b5f848cf4fa068d
z4868593f370affc9181a1c31b30ec43a4b14f6572222e1f330666c925d16ceedec2b979c7585bf
z046f7b5f03a89d7011765bb896ff7c8885ef9b083c7890ac35017a2ff1483519deb8edb7ffaf22
zd123fd10db52036eada06ac6eaad620aa55c7742c73d14ba003f762abe41a22822d61d47b2a4a2
za277025a26b8556cc816948ac3eeb4a3a87df2efd2b6e9cc1905296841abd7da490b2c62009e8e
ze2a3fef15a3982f5e1830c599d630be781b55d5efb15940e644ad3b8f817067b9140cf12a0bff7
z308934200140c96d80d47de575dc6fa31ab01e278dca05afc21a47f3e0ce6a1d62191577992ff3
z3c076bdaaa8ab2c085192429fbd360ed1af68b8d4ed84e61425abfdf2adf534d649e993706eb52
ze48aa37245175fe637ef60bc5d514df9665134269b41f9e9da7238cdd192219e7ad6fefef370c2
z49030898d7adb08753d99a9b4b96e173923480b12c8f8b15df3e8c562d895a89f1c4355a2b45d7
z9d2af6dd94c314e3bdd0f6c56f1c8aae327e473c3c1b07b8fb90929fd13c916870db1da3fd91c2
z877df6d485ccd7e0a39103393782b5d7a94fbfb1171da06a53e114714fa5c255ccdb0a3e7d2590
z597efd4eb1fb0f07b98e53f9813560111a856a8d8e19e0b808e21bcaad590b590b83926f7214a0
zd06bc4258e68bd6e85127e75ef8543a042891da3d8015aff25ac33e545e3c65c2661fbc2b4f780
z95eb232ae23d7f99002c3db6a1948516a1cc2c4b80339141827bcd15bdbfba03e9e40d5542b4dd
zd3638881e2ff5195e9022134e4a925c4149606d4b00312af9222035ca04e095d294ecb6a4b52e1
z19d074647c977b6e52c1eb908c16cb947f7cd2ffb70bc7cee4d7fba2afb4366a13e1ecd9cd8308
z039960a337cd40ee5d3b125d26ffa03e434071b4163d6b3b83d59eb70e3a92b827110cdab0830c
z7b7e2c772d4a433d951dcad51b2a35f153466c284785ff6b84dc5a09ad9dbbf420f2a15284cf8c
z8ff79b52cebe9c25c7d54a7273edd2aafbf208276522f9c00152a380655188e00e1feb4756dfb5
zbad032700bb9d7817f474e21d82475def73deb647e2e3ec1aa8e0ba34ff7783b6da175bc5a094d
z67cbd76a26377fd57f7a155edd985c4ec1eb970e61a710f361a79e444c08f9f2bcc634e8e18c4b
zd66e929dd3e0b058f9185ebe8524c789fe0b0efeb8c3bd6a9741cfd00ca24cba19fc755b63632a
z88cd2810f0ff2799cb6ee94fa5ef36e07e646d74be4bb33bc0b7496833557822b2d8e434b2946c
z34f1e20a411862898ff4b54e463a25b0adc2541cbdc0df42d73f8bcebb198c765a35217e840d50
z767e5578f9ad99fe8ae3a664b5b2ca82a71b7205e12c1b083e66a8cb380bf47c3bc0932db41deb
zbd9afee6a6e0f9a50c7aaaae3d829497fda604871ba4d7f20ef7c3091f2440c30e9f3631a2690f
zd1ed042ee0712a99aff4b96606efa103572ae5f10e1310403d8a0d62311f4d112be2925637a3bf
zbe676cf2568811351675f284a0d87fe5ba882940749eb2daec8359662586ee2dc54f5aeeace05b
zfe2b1d555687fce95b67e98e4b07d9083f0349bf164f14151884e2fab092e312ff109de78a0eb9
z56fcc5ae7ca405ce259936b42edde4257831f031090f183e4ce505e8ce52defb1e4ee085c8bf50
z2ab9c757580fbbdea209082b09652e7cd37e39defd73148a176a436787e68d073ae4d84ac68b9d
zc6a7b193edbab811e60a865d5830264da6b51bf4fc0c92dd23bb6b2431092069ef2ed65f41163e
z25923da55b6211705b93e606cb129bbf182cc57be3eef8ddde7ec5c529f5705fe2d10f30c824aa
z9c378493b75d6ecc2021befa41ada76572658849ce08ce63fe301b35d550e10334b159d5ce9677
zac32ac38375cd2b3a4cf79ebd4f1bdc6a8266f783a69280e0ec5c0c6ab5b28c4496e6a28940f61
z169b5727590b79a53b04bdc931e39032af7d0f90bc640dc2fdbae6b15dfd7e17fffcdd95e1895c
z9923ec841daedbe25b5a6fa73c4775ce6e56c7ab8dfbe5098c922088e5065c2d632f45948b2268
z2ecc7a91f683fc8bcc2d98bcc9182085d5da4a27ba5dce55b5f5373e2ae49614b2caba29c45e8c
z22d15406c539abc60a64cb9238ca6ae70b647579817a57c119c603af2dff3948ddb3c17608ce28
z33f76c847021988a2c4caa01d6433517097ed0343ee168a23702892d2a8593e0780923f2691a58
z8c7a6b06517e573fe86e0e7b71eb87cd769ca8a1cca2fcfd18869a2ca00c43274d4490439e2199
z0dd7b9a38e1febaeb759411ab5f0e1cc89403d52fb98befa451974ae7ab3e890354a4d76588b6e
zd7a45cbd90addb7578f4bad9137e65eb98ee9ed2d992987cea7bb9293969e7e9e3cda0f0373904
z80f4e36770ae0c0bd4e4230654584f34a7f4749f080defe2d7029f1e922d6c0cfc28c545b43fed
z419aa9fb735b2609005062f477c2da01a1b8d4711c3d55a70a44fc128bfcdcb9417ac5799632ff
z4aca8671433b75e3877aa830213688813e7410ee2ee1046244314fb50ca6b87e4f32a6567b0bb6
zd118314122b40f2c82ec782844f6a88f628f5ccb51fd0cf5351bdd209a45ede0e48b371435279e
zacd00881bbee7c76d1f6ff6884272707a59502dc37c69e5ee1a9857deb1e4c0a8759e6cfda4f41
zcab85ea928faedcfca08919db0326c77622c4909c8769a31c47751b4e50125d53efbe67880c52a
z657e6c6fbe21425fd9ace10be0369530460294aed9525d0eabc51cc920f167083cd6dbd3f8a6dd
za2a41080c3abba2c8c1b5bd75f2c3c609976e21bee75c26a1974d7d9017e555ba474d27aa71792
z8129cb5c0d6b672a7a2b291071332c22ef7fadf945b55ddb970fc0b1ee6a3c3cbdc768207b1c4a
z8426fbb1e4ef8a2b666a76fef05638e8b511152ff0ac26d56fb032ce2338257bd04071850b9e98
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_sata_core_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
