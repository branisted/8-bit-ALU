`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699166942afea5fb7101325e4e5ba2012b92a44b9405d74cc
z51f880028f37a4d99d3355d22f3ddb00acc38bc66e1ceb4cc6eb8315ee8483812567c5924cf8d6
z8d19f1b2af1b714aa25ec2731f136cf3342f40ee20528fe50fac4b8b6ed869837a5e29018d2fa5
z037ea29b80207c8ad5f6b0b063ee82b130d967e93d90797d1ea082ca735d18098c0d8245d9e843
ze9eec21b6dd35a1952fff2b761fbf332702575dd4d25b3dde0c8a70ca78ee95bd12edddbe4524a
ze7c0790dc29c8217048cdb296c175c356df9b93240a43970c671c2516fffbea626c7603d2d8157
z15353d575240e3a984092db6f88571e2bd7b5a82b34d7f96924707840e30ffcbe8d8ae7bc3a704
z722ed3149e9a1cda2fe6bfe96e90c535dea0fc4350407df9c21d11a3a86d6cc10c5b716d5ad043
z82a169fc8786a60bffcdc3c5fee6a4c8d924bd371b6eff878d08f4362f160c839a8f92befce8fd
z1b4d7de76d77ca37276d918abade48d1a0ac53751389e9d3f386b196c0beae213a5b20e625a8fb
z51ef218de17bc9b6e53e3b5ad24f435a052d265900c7c9f25a59237f1681eb717aae9769cf53cc
z0b4a95bf3fcf6e9795433f2a004c4dd5f6d3d641b5769cbfb330963c9dfdddf822d9bdb4c4c596
z6dbf92e87bffd540775466eb824b32bd4786775ee944b513a0cd504b223ba92db84a2389e4ecdf
z8e7d0ce2689961665be22d3f4b295aadf555f59093f70a85f278d9ef6b612e96162ed609e17ab2
z81fb668dc0fc6806e7030c1c76fa34a1726d2909e05d3c7b371151c3c505f44fd0722991051f8c
z2f62f8c9465aa57614a182daa804aaea74fe28da2298f66260fbdaac872d3f848d760b1803fa8c
zf6e3dc1bca87d7692a0a124036645a732d9b0857dc10edf8dfb86e377b80597fb83f121f76ad0e
z4abe0be5289d3acc1affa0c3b23287cf60c0fcff4d0bd46cad387383070fe18716db62f58e1aa6
z509dcad046782157134ef3160866742124046ec1dc697fb6fdfd602df41a7644c5c001cad6d14d
z6e041461142f66aa1e1a02baf2aa8e149ddca2f412c70075ddd9b5db011a82f5ea780092b3e218
z8098ae0e74e482c2b2a189635de2c3cd8849c3c069f9a16a9b3298ef733cb5d5519c38da126731
z72997a4ce59bc0c37ed7bc31a4691f8bcfffe04fd682ad60ba25181fe1b2dca296804b3ada8a42
z8f01a0f0ca2ffe90a0da918a253803c5183d1dc2fd452957f9666f95cb64421be989b87dfb26b6
z821b552be1411c6fe92b8753e91c738b63f792ce0d9bd8842cda93be5a2282f9bc22a5d93cdc62
ze8b66e1a3aec7014fb8361527f2b1e547bf09d8096c590a9394df8871dc61f7f361d8eba25b31a
z92fc4c9f73e58106c8d82106ff266a0638a03139ba259a29b7ce45e399d2aad482b93da387963f
z4e2989bf4bd22ceab9338c500e9fc6fe9cee59dab0c281ba7905f8a2175cb7513d75d5498b098e
za380810a7f3e2c2186156960732746741b7327d9054b2a4b0c631b10ec0b0f7f80e4d5c10ede2c
z8814a61f87ccc0c0c4e3f71b66a165fab19176681e000d72400fa77d3c531493afc99cc2dbad06
zdab5b1696312540054d7ac4ae422bda51307c7483b7b5e7a5dab1b5181bf3f47e6eef3f99cc9ca
z4d4e4a8a2c0cc9adce4753a276b99a0d20a5f179e7fcc1ca48807d3635544bfe0b0b1a879ebdee
z068551b4488f2d4d8dcd4eb966c3ea322d7c9961dd68530141b3c471d443ac85797bfc33f7ee12
zcfe9b2b3d5a28d78059ddec08e3866b65d5f923fef13be2d30110f4bbbd009f36473d2507c1d03
z5f6f1b8ae320690b3365741de9063b437744f884c2c33acbf751f08ddac4524ab799120b27fc4f
zcbb9415f0af37eaf1275d36ba5e30e4d4c3cf9bda6df47366d459c0d31bbd4c4ff6d769a9ac6d0
z85ac457e7575092e745f3bd984e8205a653f04ea4b9f41279803265af6f1ddbf6d91261eae5caf
za9334e85308be03562d453a1a4c02b9b4cd5f446737e69541afaa35f0814800cc41db3e8870145
zc68ba1b35ec9d09e7e64226105d04eab478762fbc14c94a21c7a2e3bec7f761b92cfa3cdd72335
z6ebadeef6552a28fbbbf9d3be51045c675076ad17a62ce4c7bd685442de7129bb65d6133fd254b
z6932b129108dc0113617f5de31a1bfd997583de6d8c13358e5a6bcd3582075a61658c68c58aaa4
ze096d3c2d44c77cd4a45ab7c97cae7d3a1f696c96bd7a1dabc67bdea399238cfaa987828ae648c
z3f20ddcfc96caef1b35b615d62185d308dfec51d89f0881f45c426c4394b7b61a2aec033158cda
zaa1600c8d9ff96efa7829b091514275bdb8e3d4b00cca0da8e521180f14cde60689b7be37f807d
z10eb71daf6437aa4693c5e08c813f83bf5582177597de66b8fe656c61aba460339665e78b334bd
z47673e60e99719060a289ee8baa7101d9b13f5b2d54bb3951f46de49b94ec3fe746249528a36fd
z66a90f40b53de9caada21a8f28f473f129309e305afa1a1c12e575b2d44015f61ece7c2d5c7b72
z67881bb4d191d517e3452976a942b7e698ef2283b9a61e973639f9dbb65058aeded176385f6961
zb6eaaff45e35eee6ad2ecb339839178d06a8798e8ca0745de3a84e0e4072ffafe57f21d0807230
z11902f674f4c3732cec0c6042da92a35be6a5e6e97c870d7a55935a7294cc3e8e86690c83bb71b
z7f2a89e514b4f0abb5bc8ff700c39b5962aea30bcc5d7f6b2d7340b4a55a57ae55424953be815a
zbc5763c6ff6790d7b75dfee0774e5da7a23aa7f75d7038aa02bebb1eab0ab9179138a80d88f282
z0b8835031c166abf6b051d93880e81795e255fcb1024793c771e4b623c9573834ce22cadee6be1
z178f859112ae50748127b01001ce5a294a2c61bb673e5338e7abef65756c410e320218c5f90fab
ze7d68e8e8fa11b5b1fe781ea407d9b495f061804bbe23314cfdc08329cf3850dae8f7e0c12a5ee
z7a49c44c22f578bce4e68dbb280207931cf2873b968a469b69f8b5eb17daf74d63dfb8b871b017
z21aa073bae5c1c2410d9ea1969458f557a3cd0eecfb2823d12dd0a9469a8c579c9f48f77f77bab
zc0e781022e53d7daad534848a450e56483f6fc15444ef920ccdcac9380102d19c689fe1854937c
z04684c75974c0cca37a76f1b9d5b07b3f23bf2ed6905f72124436005ad02583d85c5347cc51be3
z8156623b8b63aa21da9ea2cd7a94dfbf2591fd135048b4533728f3a13249275e82b93a1b4008c2
za8995173341f8fdb75d74af8a100b0efa98daabf352596ca8d1569ea5a8495e861aba62251eba0
z1d27470fe106669a97ee8b1c71378de06fabd8bed57ec6a1400a9c700729783d25b9c6d973a3a6
z0707d55c0d3fe69d025c565cb9d759ecbe0be22f5763801bb4b61f7ba6649f36ba810f572f7924
za74357a62d719f1f531d3581910a865fb54945234ea6fc686948757528109b6a0c6e6c4152946b
zd946fc707ffdd0fcf1e80b1b657a30c09def3bd8cebb772b4c5872e004b9ee5c28a2a4808fb682
zbc88fc0e4a97e50b5b8013b25bbdc450179d25c7d1cbc39bc28d52cd791bc37d350a23847de17a
z2dd204d7213c5d9d6c97fbaa904e4bffd12112399bcce2efce1924d4d8bd0dbb4a4c0e700c4ffd
z1a49bda59c61f49d76f77bfde7a8448301ec69c9ffdd08260da435d45540d134a88033e9547ee3
z507fd61adc10a7f0ce506cddf518341293de780c3a2e0235f52db253181dd47b22161029c90ca5
z521e5448a45da1544f268872c1c35448422bb914ac9540ebf588bbdbedeffd0579c8d4cdc607e4
z1dfa8dd5d82c689923567077dfbabcc14a1b4dc1b90826baa62226572e165079c295c23317aff3
z237d3f96cbdcd78e2fb3e75a7461836e82a093b7299abd9ee161c10b08a70a17ede1a9c82e96d8
z3d6df006d6f5f2d99140189bd3e16c626e643e00f3436b4caa3161d0f4e969c8f54f47e8a2e6c3
za11dd5ab417382eab30137ba2a27653e473a20fb6d60c2ffcee7bf1a1abbf45de246f116344eaa
zd043096b5957c303ea48041ea124d8974da83dd1e4054e1bfcb9a622160325c7e92570483656ad
z7ba8693741266a35166733c382cbdf14f9d59613a1f063697f117aeafdaff5a272b1ba6eb7312e
z31ae47b778b699bda9597456673dcc21c0a5dc82a218f4eedc4c1268f575c880115652441ea308
zc86ea1dcc71cb154ac246313bbf8608b3ab96aee70fb200477c8bc5946bf572fa887cdbacfb9a5
zd39e4e987a75c4efae7ae5630c6708cc710b638ed0cd6ca7365a8078fbb4729a220214b8101751
z76febf61ae3b0e888c76e3a3bd96b51163b723622dd409e6bdc7b803fc9a5cc8362b091bcd31bb
z05e9a80aab2c2d695fd522e4ee96612f14f2536b0eef01df61e8cb1f777df547cd8785ee2dc0b1
z79f03bffe5146caa1175879117aef23e9899b0ee17b90e2832a8c5f9eaab0805c2546fc35d8aa5
z10fe8e48887b1fc77c03da6722692ad1efd84f589e86ab6abb32206f6d7e2de4ad7739e0b09bec
z0445032c6ae84dc0abf9402ebeb61723b9207ea958d2207b73ce4983c568b4683b103c0bfbeca2
z37838955120e1ea527a532d230046c786615617e8385290607a66f70d708751028cd0050d8500c
zbfd2ead67365aa8f1287260152d23b61d047cd4985dd0a742140818a8d27d18321571ded1741f3
z94f8df5300da48d83d297bceaea3353bc2d43eadcf7864571787adfb24c79b6907b88b15846d03
z266960de4185ba4d7fb70324086fd52877cb9f75856c9d729274a443f27905431b1d32e2fb16f6
zc5afe8a2787816bcea07bfe5ca3512379dcea821e1466a2f10fe7f01edb6a9ec3f8edf89178bdb
z741bc1eb8e71adc6c6c880a38a10b288c0186a7436e16d2c7eaea7c11f414dc910f91883f54142
zadebf69e8658a1fbeb1981399f2421a612bb2f54b4111106fdcbf217657618f71da6c29c428e93
zb2e0f8980207cd8b1cdf5924c86be182eb4f489be070522bd92f2e94b71960ca2f5e4c8d8539cf
z90d469ccf43e74c264a4b8aa53a3f3205b459c49f611c9aec4accf677b469a1efa8197710c3c98
z6bfbe48793441065af2c784583041ae5f6b005f2cf50f1162ec095a29e59f9e105a8bb6a793f34
z88c92c2ee37defae9074441314da39871fc4467ec5a9fb0a60579cceae8e28ae77a657e42b2568
z60547128607b41257314402bb782a91d1a87ceddf038b570d2f66ea6e777f88f0da39227672f20
zbc3f4d5d2e35d6d9c3240c08f2d1d8800be2a0cdad728344e1a4ccf2d5afb24a18ebea551e98cd
za88e711f1b60630cb1821d865cd10847033b5f004138f4d88604704aff493ea6627d60fbedb6cd
zb7c77082c71071bfbfb231104f45ceed9cd8b8e006536b889d41d12c69308a661208883709d739
z99e236bf4aaf8a22258ee9d94eccec3cb3618dc877e1c93e9d2b2cf65f7d2d69530d275a185341
z2a29e05ee832bb8b2b499aa8ff65bc2d20ddf07e71d175972c1a7406bdcf2594199c6a7c1d6fd5
zeae5a7bb422d960cc549ae801d60330d44e92e905fa778c1d881c1f33f1588b01aeb4b74368550
z91fc626a32de940e1c89010ca9085f8807bf7955193c975155a8c922a14e5b8e6224c414a616b8
z2c190b1a21f178d6b5bd5afb8a8e012b743ed3eac5d45a5ae8e83231009fbbd2bb8fb46995c891
zf2708771e3d48dc3d717e3fdba5f88da4f997daeae3bab2adf7d00680cd895060d33fd6d6dd7dd
zda50ccee4184e67b5e52c7b3754f16ddf6f05636d48a1da6a8817aed89f68d1e79d493063c575a
z57a2841d5e2fc4f06321cd6dd5823c67888b74e125197529951fa680f1edeaf310a7506a74781f
z794585251830304082e104031e036f951664420d85756402b43e2bc4461b2e32cf5d88535200cd
zc6d6c86276cad5bd8cbae745556991d729be1bb011c2ab6ed4e55c8ebeed3a39f4b5e43be2b4b8
z5a85fff2bb066089d0ac86c25df183b3999350cb32f5311e4bde0685e9de4a9e23cab2c6539410
z3ab8967aa25a5ec07fe9187743e499c8449e0325e09368acb95b75daedf9ae2a306a5014d24b46
z71a4163c54882d0467736702572c954eafa421e278adbf5642334d9cb8400eb1393afc1bcbaa06
zd6c211a2a2ccffdd09b0f1c1f1e1caa7f4971338ad56b7c6d03e93ef5a76fa8b60760e2b47ee6a
z32f1731459af51721aee980f7d2c1150bb4d4cb653eb7188ab6285f7d757ed832fdd3cc72bbc7a
zaf324fc7202c666faa771805bc97efa58600366f343bf00fb9dfe3fef91f1b0431c134e60f2591
z5f8834deaeb7e25b48fa73cabdd7f0a983128319eae036f17400d5bbdb10ee6bb50105967d184f
zd4f966b8eb13edeb924677ca0fc00c52902cee02959c9c17a5f939217d604fd2c2b97047c55f0c
z143b6359a4c4424a80b1f4714a5b69d174a5006b2aa0cbe20f723fc1655fd8e5f08f4567dc2ee8
zf5e2182665d0bb63405e1eb868ef254993bf3cb11047f44a5dfa878dc5b977e62fe13cabc841c0
z4a54df50df850830ce9c91adb9007eb0dca91136d9e49f024abcea41aee6a5059da58e93cb1d57
z50ac69947e7401b95c785a4ab208c01ccc3b737160ae1041dae7965fa42b4e2f73fa47863da891
z02749f2d56db2e9886c659069b42e1a669919a3981177d7034c1697385822b7b608fec9366de56
z1e5c0b31a7d46b2d833db58892bad8c3dcce98786402e4db467bf89bff43da33adfbd1c7905369
zd48a5152253dda219f39c0be2be88f6993461b9ba8f15975e342e6ac87192da47780f89082eb4b
za4c39d73c9abed030ef86652b7d65e7d239f299f026589c3c11d96e673edff9d1aef68bd8dc774
z5c5bd504456d5cc9e59cf73bbfc7a4184bd8cd8984787fa259f79ebf721eb91207352a59ad1244
z2c41e813b67c8da39f798474d77043d0f356184cf9a35c89212f623b7d666d508971ddc07c55e4
z843f8a2a6e95b8d8ab5cd45c9f6cf4c67414ca7f2eab19f291052258533555356ae6e88515e221
z7a1c8f8d7d3284bb61bc7cbe26c260eb27e768f7f791bad980e5a3e423735001d0700c2574d8b0
zf509c199b9179b91d82729e89b71146060ba01967b0478561d5d3a71f456322228ab06831fd6d1
z2fe02e388a61c1a454f671aba24c35a82e4cf12544f783d8d9be84913eeb598f88a6899a8d9a85
zf8b350e1e7eb24fd163c1ee4701fbbb0aa5171972e3075d1162f744404062dc38a1346eb9ba91f
z9cc02216814fa323e3d71a1aefd800a66bf902b4b98b72b11eddd2a298b71c7e5618ba9ee4e226
ze67798289c258a1b351a7e217c80b5fbaada70483036ab673c7b974b0b2085b4bb28b9586f19d0
z0dc7b9a2a7d827f06a51193e36be350268a9311b75e0cb4fe470688af128d4a999606a9ac1eec7
ze418adb3d9252f62c6c42de6f2a4ee99a345162e1a7dd6f11f513699b2b0d656359c5d50119b25
z72baac6ba8143f6f789ab8cbc53fd573d6400a9a40d5a1171635da91ceb6fc198adf86e2def2be
z6981149df7abbf69d1424a5063675e5e47b87ff843f311eebab5150dc6e1a56f05bfa75c9c2485
z16b7bda31200e47da0279de4fa24a20f68023064fcc36ecdc6b9efde99c30a3b7eb34c1c8330ba
z9d27a6b5d3a49e09852394f58fea5965c77c9662bb7f14c929e129a7d51c3927c157d176e151bb
zdc3b6fea6802a067bf1c447f8272800af0a2c1aedc6368380cc2ba7ddc5dfbcc19b6161adf6bd7
ze21f98873d1e48697e62afc5c96818ac2e4eaa10d4cedc0a0f5d1bf9b568809829a0f93ae0678e
z75bc356f86b54649d378bd3a09b393af927f6f19545edc4e865131fad33751c2bf60a415eca965
zabecec0d0454a6f6d48a29b87336e4573b949daf23b2fc28f9a37fc071d000e88a6206c661ba90
z0b83757a8b96628617852010119106e75b4690cd9b4ba6540cd453a527e410219cbc8a6da471fa
z07d08086e14fc9f9805b0e1bdb6a6bd835c96f6ff57b4a0db7c53910c411fb22fbe9874cf03ded
z910458dc7f8534b8187dd027917d698be996d816ae16f81107eec95ee814c0df1840bb7ad5f837
zdf85b9915003ff64a312bbd2fdeb7b7de4948237e78b9f0185fd7ddc6f26ec1e45387c35880132
z7cecea46f0af3a7af8238ee72e72af4549f158b9556e663699bb6be937539cba32da0f68e28c8e
z046cb24fe3d0d3f755304297156769c9bc06af4623b6f71d854b3546c03495885cb5db047bbf1c
zdee2867fe14621827f05d42128810219b3d90c43103b9f7ec22ea1d5cd0b716e587b2442c01a20
zaca5d38dcb89d5c981797af7d405504d35accc66a789a6928f0b2a8bb572d207767279b0946f33
zdbf76931949f4e0cdb690ce0b051fcdaccdf27e48e56dbee4ae50b756a2848f480b182dc9c6563
z8324dcab125135841ffa0fa558fae3ff6f3fdea506370b5d5592d41e82a049bbfae122146fe181
z5f9904e52864b50f7e9275c99b9b1e1b0f4fc94ed203bccb9afd995744f5d7acfdd48e40a42b79
zffe22248744167d80988ea40a99a0baa9e3c9a17c78d8be8447ec0d534fc4d997b45d5d26d59cb
zafc77fb2b37460374a764e80d1c8bc76ad26da4aebdb3751c182bb4df223c3554f12b54494af8d
z278d88dd848157c90fa9031c6893cda7c7b83452f2291058decb5b8ba6896adbee17b5ec4a7aa1
z6e5a1e0b38145b54351ccdcdb88e12791a7232a55d941fc28a75f141bf92dcd95eff7e64fce08e
z660ba06e34dbf972a6a63e9236c6a215b5d89cba10e52713422030abc4f728189c0b44831f37b4
zbd515a6e21ba76593fd97cdea6f131264a4d788ff9c29cad693649f9db16feefd7c37ce60d0ce7
ze5604c3773d58f412b9ab1cccbfb54ba7d7d44d6f45189e2ba84942d7808463b7e9b21d2da2cab
z80231945ddbf245484c5ebecb99c85e472620bb22e49d638ff7538c26ea4dc617f3f85662692bc
zbe6468962d8026184a1174eee4ff01ccc06fca30abdf4233489c8b3b649f5340225ee1367d5961
zddc3fc7cc5c2c758f8510d4b2b0050f73cbd419a5bd01b364f5ebeea556aacc165720bbe9d5d2a
z2d78435f23b1c666a18bc3e7614e848fad4ae4ce2ce98b8167a03d2e7347a84eee5923624ca595
z7f11053ce780f0ad9c9e90f486c117a94b3d22710373c73a1e6ea6539ef88f29eac6d7e03a8503
zf3f0db77467a4abf835110a5ee5851c18033457814006fd2099719fea753db8497ca9b595c4da0
z377870910c9801322e99d0df0d4b579d7177a0aa57bf2bf1ab31a90430092b6c9d998a3c31e00c
z2680309f594437e84af1b0d6c1d40120890d483b84bded5d9ffe19c05f0fd66a57e4d6c5d9af4a
z12c141ffe4dae67873907093cbd2f3eb2f22847742c1f0eb3245612719e9c94a99830b9aacc336
z801ad00cc925c6273a77a431fd7dccbf0ee04edaf3d7bcd0d7f2bba5e83f5d1a55c5c05a1a2120
ze9e872862a455e860b3a087450277ab138873e56d1517d7538930158144e28a588acbe6b544b6b
z3eb4d48072788fb71bdf973528e173db9419915c3def4917a8969f517c1eb6025cf877527bdcf3
z94e3de21c8d4b8fd8e379a00517a94984d24b1035a0caf959d0a31c6001667b64c9b60e5d59638
z56cfd4e30d8cafbc1920bc4962c27d0a5cdfd9a8c98bf20a64cdea2e5cf6f848dc35e4b865ff76
z29d2c30e4c8f2532d30e921f57f673b94ab8f8ee9d01c9d349c80d377a5d5f501a4627fd7ac686
z6d5a61c0a0bf77b46815afd4cf056bb3b31ecb297de03d1c79709b26f267fc33ca29543333c385
zab4112d2ad0f71b1af70b1748fd4def7ecbbf9ce3c5cdbb77b4a1e84f343c4cd669634c72ead72
z55818462ebe8e12c29458e455264825e76c688e4cd22db9887626fbfcce5bd1ee3cdbe9e3e7d1f
ze44e2a56172b8767ef6fece9baf5c973be61202e65b061156b329328b53eb38d160325430c84bb
z7a8f5c7e530e01cd49a7f25406a69da63a491946ed7046768a6dd4aa9010f2f21547ff68e9390b
zc49f895eafc880925181159217c9554747f86f702a34d299cbd8fa25616b5da4a72c3be80fda6f
zbceb7bab17c6387615a7b88ab6395c88540efc402bedd71d5a7c16409843bee0132d4683eca0a9
z735a30940de0badfd4caac26d2e3e59612d05fd618ae7204d90f6227ee2f7084f06a78a3bae318
z53aa9a1b4533df589a31c29cc55a739a6e64154412e17b5c4cfbc06f12d027782d9d71568a6478
z268d595f9425185126248ce66326e6bdee9324a3ea62975f56b7da6948a2b72c3e4c9675806cce
z5835d79d9f9e0916609c8cee0ba8dc6b320aeb12238c8bcc2dbcd8223db980e996be4c50c25c87
z84dbf332f1d65c468afd93dfcbb9b272491fe78717649652e96d8a5738c657c7b9cac9da510daf
zccb9eeb135964a09b2c6b1983fd075ea3cf9ebd4c4c5c3b3daccadda0636fb128bd4c352058cb7
z14cc47af4b3c6fedf6e9c8ab5d6023ce779c5407316d94db71d785da2f43dc95aca3845e8301b4
zcf07da08e839b763b962117310f5f36611ba18d76069aae9110e85997e19e967b7e02fda164583
ze7c496c77fb9a92abdae3b5683360b4a3125f3ad486a9c079d7c47a1e81360b254445abe37e5c3
z78b86b83e491bf5c4bfa2987f9774ce489c3bb4ebdc52add63b249568d9bd241a12a3a136392db
z8efbd869dd2690723a3c46d5bc9b61000ea68555a94829bd2dff4e6bd059a87bfe04643943c69d
z57eae53892d4f47c8f412f3a05606f732ce593534247aac6c528e385439c3dac853ec739a3a5e2
z27f6004b3dcbf0706709f0051c8088455c81c38bc7fbcad5ae89d1d67b9475ef507cc55eff9e8d
z7c1e94877c31b187df30a56d2d910d4d20e1a9869a3e158a7254264b6ab425ea42c5f37863597a
ze5b45206837ca16e962a6693bf6da812255b6f0cc9716e649549526f08f64df17131dcb04c91c8
z06b7a1844a22adf1a51b4d573439ff0964603ce904cc9f2f018b728ccfd5a064ad3e916102778a
zbbae1de55c01b3e65401d6afd025b817ae5fcb1751b339ef038a3ac57865145413fe18d365b5ff
z3eaacaa896c8074059780759864a7a2f3d267d711046c1e43b61dae83ad19dc0cc0b6f69dc57ff
za3162f8b925fdfd8bf541384e726ea06bb61bf9d722418e3774b8b6c1cb1914011c6c68ffa35f9
zd3414b4bba24ac844b2f2c28326700860bf6ff4d18f375dd975a1aab26046c1543a2ed8a84515f
zc92e6eb4874683aae15fc5e3ed4dda7188afbfd73850e57010c903c7870e1517d5041ec18bfe57
zbd969f6f389a1b125acae56ac0397194643047567f7a492c93c5ff47eed4872ddcfab06d10fe52
zb6c2c98d077e903e765846623a2307fefb48bb7c46b24b5604cf13cf6f21af3300c34a71acda94
z37caea744351b206f0c6e5c844a81e21958df1b2d8b9bfc45fbb3be6a779d5aa7b3af1243a1c32
z018536f37bc2274c4a6f3b78861682ed7723e4c8f90dcd760e1027254b5cb759832dc2c1f53501
zd07a741d10cb1af992a6d3ffd5f55e8930740dc9ae605eda6fc3e3446a1bddefc0f3d36b359420
zc61d42b764a7c9270d9ba2f448e113d8b27e8c7a95b3719d130523e882c4970afbc534008fb954
z1ea1a8faf843dfeff3fda8e6a3bd6651847233529113db12d11467eac6a20e6e0e845489a9d69c
z6f276efb58718057178db68dbb798091ef9811143e15bcb0dbb027b1bcc68a958d835c67c249a6
zfdeab00f27631aa3a3b5468d83a2d414561dc6590698e294f513aac41295d8e9c2f404efa61115
z6bda5838bc16ae7a380dfce1f773736f66a23320e06a45b3e9969831e3a32e7ca4f468f9dfc2dc
zd7952a734187bd38192d024837395edb482e1bc1908016e58eec73d4ca818002fa14f434e9c3e5
zb0f15ede42d0074793c97ce1d2ee3b3da3efbfdfc059bd030a4a3938ff51d115eaae5759c405cf
z567574dcd7655a5a37c5e2f99cddef523483b1beecc42b30f5af4237a3fda39de7c29af79b108e
zdc73549f324fc8fb346b2b302b93bc783c42dfa2b2beaf2aae755561d05acf69f53c3cd651caa8
zf71eb857503f66c3d608fff4dac8abf9d357e2273f4f483b39f1f66945abc1bf9db64d68281fab
zcf9adc814bf279acc0cd510ccd6ffdedcd3e892452f3783d10bfc8dc6a74aff86a0a15a0fe971e
z11df4fe2e19076d31a040ace8ae9fe63a662c72ef2a8af7da19d73cbc7bdcad306426821fdef48
z530f94a2a6cd7700722b2d9f5863fd6b223b2a33bf6a21bb8eda28c601eed913581a7d93fb789d
zca6ca5dc8d560a4dffbad9a94af4a65af501d47f7ad824ee1b2b7cb0cf6c128ea75c6b6fe16cd8
z59a91b93f7942d5d2184a88fedd581f98bc72c4cc6808dd82a2e6856bc13d0d477959027ee0a15
z67716b4b6ff63d38f522db1cd9bfcf74ba68f8d20672c9e622bd478f8c764933ed910d27f18245
z5a50174045ba631c282dfa10e12235f42672b7464bba49b9eb168ed7edf4e2b5c7265aec7baa7e
zec044f17d676e7cadbc01e4d0a7569f3eea2ade13522bf743bf90fe50e898d5396c4863c26f838
z99223aa53cbee32c0d163671078ebd67512514cc99242ac9d0acaa3857ccabd39a494c04228bd6
z35428a2b48beff8f7d279e2af3873f5388c4a2a284ec78551e83bc96aeac213139fbbb0c9df7d5
z48424c1a7ce4e1874d2c38c0e0c37f3841f78e6a6564edfb34855d563285e23989b37b442d400d
za5f4c00b555471408bbc978e25d30a7ffd2e0d27cec6e6ae10f6baf350c7698d989aee0f354189
z070bc629999447532aac1c2ade468cb511fee82f6c5fb1d798d2f5eb18e65de11bc4539cd892ae
z59c0afb5373d813d97a0be1599f1f4c915fcc1879ffb1c002f535ff7c4d5394df1cf9d76a2467d
z6bb4aed274770d25059cce521df4c31a1b0b8524e0a915df8eb9a25294e2b2773b2e0ca4a25b73
z4bef546c003aa035914bded78cbf9e2a79e421b0c8b6578e26b607b5eb6a171bb7d4f40df8903e
z1c20173539e4d48092927575ab09e756f2260e0351818d63a18352619b389b3c7207feb830a0e2
z7c8969643a342374d03942a8f83e3db879c10df17e4f6f4518b3ede9ab7cb4479420f18e4b846c
zf6ba24b3c98b0252d32b276f73dbc816155b171d0b7c7131633ef334c0c7948d283d1804a5d084
z09f41a5e03c311175a62bbb5312de82f776e6845c057c88afa1cba1f15f9771fdcc65cd572d738
zb892e74bdd292ff8fff2bd87a6c1d8c45014537aa6b210c642d1d8adf61a8c897f08d1dba31828
z7fdf7119201fc51401dba36a0ff41ca0f122e9d1db4ce7407d8f0621c402f23416d82fd98a1c19
z6fa01a45ef7fd93a42eee617964a73fc8649aaa4cf3d9033081936f14ee20d539144bdda3e264f
zf5a498f7b8a630318e741c2fb393ae859639d95c66c7c597d4e1822183066e6d7dea2bdd92ff42
zbe7976036119415ffb2116317b6785322711e51fa9b2a32ad03967b099bd434b355a366f318a01
z4318e97642f0f7c0f06b131a97daed2e321e2cbccb39abb4044f4f08a5edfd8acdcfdd52889d3f
z2b3e81802767cd2c798fe74acef4077b347b6c37022ecafbddc49ed2d80259c46652c5956ff14c
z936aaac6b7bb16a7052402a8f6c33151ed2bd69d1d58c3a63db1f8f2b086d60ee0e5546074f4c1
z045ecee9cdd5eaffbe477bfbee3335e8fbd173436e7c2b06acfdfacecbf1b7f172710130fecc35
z14311110f073d0a9be702117bb8c6507fa809f27060ea67a366da90ea772dcdb6f0849c5f6f76c
ze921a4b25bee87e20fd0da52fff884f49bc7ecaf6c42b42bb43b2bd2601e74eec5faab432de971
z2e1d674f1eaaff4444b54ca553af579b8ba7dbca920c65833caa85d8868bc38b290b9073143e34
z22f97e1ee33b8350041152128a0e942e2d33d04c4950a703f88089bddf10ac162f233fb4236d18
z2e6ece0df21eb838b528660b529e7fde479a8cec18938ed9547bcc8580219830c8fab47f03d344
z45bd825443e86e27d3350c9b1485ef1c7df0fdd9e38528b169cc6aea30fd0d4e36ece399e7bc0d
zd5fb8bfdc41d35c018a24a7579b6f7282c2a68f7f0f42b923457f72ccbe4df4ea32c7f43286206
z4553ef614ad8efe5c013b8ad1f5924505d28120d529c02c45dc6a693b4968cfe3e654939b90c1c
z0e97c1adbbd8726176626c24c84afeea0766a5d9cf9449121ce9038615683699dd27c7ca73440b
z9862850f15bbe92d6d551fe6d0a9543d9ccc0c37586cd90845020e346fe9f3c05267692d7aaa12
zccf058027917dc45710f3177af674015e1a1afc40b97c4c721ef0fd72ee8db8933df7996ea4ed9
z90cee4bad92555786e6bfb3d8b3666746e61a0442e92dee3bda8317fa7e6f4d51b73b4ae02308e
zcfd464d1095eab5bfd790b52e51345e09b635fa490a8ea7aba7a34687e31d8d539049112290425
z5a02f9b50d2e2a94c92609b3717ea94dfd3f7e8fa40ad0946767fc2f569b2cc6cbd948b2e241ba
zb32138243bd53de420612f6cdd99c64ff62b2cf0caf2d99111354ff78cb749074b7709545794cf
z40189e6cf7dac57ed06a8ffda7be21e2eca51ff1b484eadf1d77c353560f8ec81a152784a15051
za1365d8e0e658e840a9d57f7c7a89f20ceb3f28bd68f7f042f3877c23a6dbfe7c3d666207d58bf
z7d7224a5d1b547e799bb26452871109562e82d0308910be6e37ca0c49696b81cbfe7e42f242937
z1803bfb7a3a863a446697aca3a79178126a778e7a7e6dcb6ac94f22697ec8d3e7cc03ded2a9e30
z6b9240d3ba255b17161f137ddece242777587df41298cec797a2bb4018a83b4fb1cf7cda9c1f47
z933ac154e0043b12d3173f4110055620fa7d2a235bc5a818a06d9d5d68a634419381061f627cf5
zde4176e5c7aa4622b629ce15411aaf10827b76183acba6272b6b8a66d1f5a868d557f2c97b06fe
z52ec11a6cd128594bd63105a89c6e70f66e4a4dd44c37d8907ffd1528fe72da40fdc873e875cf5
zf34110573aa945cade55bb00d70d586ab3c22395d727b17bb65e55bbf85dc82615dfd04d62fcbe
zb149004df003cadab0e34bd42ed000f07a44c3e7b40a999db5929ccbe9c30dc7c1dc34f4532d0c
z553f4dbc19b003c80ad6befc53cf370e80035f318eead52495d0d947ae9e80bd90d918f89bc7e9
za7d04635acffc92fcf93f71974e573042c79a51a28fbbc6fa75e286fe3b0631d8c09d3d3777095
z439fc9dc19d33120cb18c2d6de02c1d376c387bea74f83c52c6aa662aed4b47a58a90529664128
z9f267a669e3adb3880504a743e8ce39387b58309f4033450046062d3aebe3776d5b5c520f9ebe7
zfc9f9fc60e10f213b9d2f06c98f35f357921a9cce1fb9fd98e2f8e299e592ee458921d0d5c8d34
zfc984fe11887f39da6f0c427303ce98b3fccc2f9d34bbc04288ea0f7246f02a1e8bcc9254cd9e0
z81170b0d6082b5caad27ad555736f3fc047433c7b2e552a25d3e6861fff7b2dd2db917838d6306
z9f9ac909d8182f2aa39aed8254c626352c3db032357b1ee2ec9bbd6bb5b17fca0268d727c88740
z409da269e60e2f0f8a686b71defd26bcff54ee0aa2e869d023f7c80d6649d0339f3769d75a5c41
z779a2717d16716ebcc6db133e9fdca2b3c9b2c964db086ae473a37b4b3fccab79407150e711d7d
z81010310a94a5e70b1b24e350c60e1f83f6075651c153ac2e057e6d91b31330ed89b7b5528d7b0
z1d5c22af97a6ed422e924a098eafa3a2746b75b583ac020675b8569b711fd3284a4b355d9d96f8
z927e56cce3ab4827b75aa839aa0d27b9f3348c5fef9f6324c67312e697f9868db9b56cade408a6
zc3b253e79c4ecf39b7079faccf13187db81821b31debf704e8a79536f0b739034220a91433ec15
z05de9ac8e3f7c6e3c0aded9d48c5a1bf5222ce0ad9cf962a90ccd19b448ecab0d023ff57e18ae6
z88eb6e0c211da48b3fee12603ad37a1afabe92e30696a2dc67385283d37671414e61818b04a50d
z89067e79f89da687e28e23a446b1d525191e12244b1b9d72bf1a41772748a5a24edf2097c53e0b
zad45a696033ff35f69e780d99a380f8b7f5b7282db523fc05a69873fed152af1c55d86c72f4e08
zaaf58ffaffc28cd959dfbc44e737b391a9941c06c1de5e95e4faee2e625bcf58074ee78a65fa66
za552c5442be535e3c2b80658812dfe3bf84c8abf7f
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gigabit_ethernet_xaui_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
