`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026251e18d0ab5f991ae6977f59097
zfd09fdab6b6409e7e0a1b9964ed96e3c6b19e365696040da73432c85429c758c1172aaf0c46ce7
zfb0171592f7c53c8ea6f62a7ade6866a9a5c54e82001f0587f0edc24f4ec3d15c31985c4578973
zfc757ee295ad6967786147465457d534e14f9f9bc4947c3f00afa459fe8d7e34912040011c23ea
z356aa8494a105aebf21ffcd4f3c84c7d4003d5d04ef8009de8dba4223d2c15449eb6b288f42100
z55da01538391e2661ae096cc8bc4f049d0d919f25549280e3259f0d548f1bcf8dbda0f1d3c343b
zb65226e18b6e9d1a1c3fffc6e0ebf4aa96afaee8930f10de5fc4113b8edecd2cdf079e6ce0ffb5
zb6c98ff9c7155914fb03bee631cc174e4d59fbc2488b29bc97f9148efab050a77c4c14885ab50d
z54cbec68781acacc8db85c1a112c8d7271a8630194453b2e5b3e279249c4f1e40b7dc16d964664
z18f9139c5766e447ac6c394c41d2eca73b244323001e27d434054ad6ff80558316a6b407872c77
z20273fe97f93eb8df386b934628500e2c5cf7dd8b058f5b70392f5e79ea3eac2f11972cf516df1
z053c436bdfef5dc738fa8ebca344570d320bf3cb7d7d44d823063522da1f35537a96800be040fe
z1277109798d250f1e923f54ed56bb681019cfd31eb098c4719ead2ddfb9842a9febe0e35e3b97f
zc9b398c4b5a31595cb09a8cce33d4370b2698b4d95d0a751da8a665cb239649ac135d762ee0eb1
z69fef13ced1d297164bad3c3800c49c950ab07fe642c0e3d7d98fa84c65acff0179b2c51ec1a52
z8b529a9c69e4ad5c122fa79a41dd3a6e50ec694c9a1a8b955d8fed3b643ca515340316a6543ae1
zd4a4cb1732b99dbd8aefb12f55b5d7ba2d1610acac54f6b248c393ed273235dbc5d3787b37c97f
z20663c22b3ed0b44403ea82981e707c0290c1f2b1d90218949236c936d1913541ae3ee6611849d
z93d9a156204eb0b50ceda4a06bd7600c10fade545469f9e098322fd4191cc8b952ef6414886fb2
z548ba500c89d199d8b5b3517ade6af549ec7f283f1a3ee2540777f86d6bc84f17bcb849e2f4697
zbe8c2d840648d3a634cd06706865c18a22c32049093884d92ebd9ddb89d9e028b645c78a56d1b2
zedb9edf63ca34fdd76ba4f760953c7f1bd29591cd252d5307005b9f4ac194a2d62ae38bf27f13a
zc0a4919d6948f586c8c3873a376a58f01b20d60ece2121732608d90de5cb86514bc1ab30a65c15
zc414751dfdb126dc3170b8510b983ba4697466dd82e613d2b97cd3e6b2aa5bbd140ef23f0f17da
zf21c53c2e1406cbf740f9c223c670736796c4751eb74aee4417ed477bb286d455b969e2b5ffb37
zd71aab1b1a92f84b56b0950e0811fc6b35a4a6d2c09aef8499d98a583e92364660df4de798d1e6
z965639650acf33b18f97610dfdea182496948afd0404e4a7138ed95beec5a95ecfced9419dd9a3
z7e705c316b05e89b8570c8b0450dc3c529392d07d9c75346ae763bcb9dd1e1f98d5e90e77ae15e
z5a32d51743394b30bf56c65b6a35ee2304fd4e4f38acd9c5ecc547197d27903161020ef50fe603
ze76cbf1e85d925a0ac993c8f7913d9bdfb7c7305dde9f162cc2820ec90ac4dfe39f305d4f5cbe2
z9fc539550871d145e0d4082ec1c6973b95e0c82dcb44a174b045b1c81c8790ea2ea4a08c8ab39e
z9ebbe455974e979bf18fb3d7dbc145c87fa27a4efb8fd137da89eaaeeb6314ce1053301b51f8ee
zb35b1d31344657de09d635b558c3f96a7af88e5da19e75ea6851ef256660120bce41e521d5490f
zd9e5bb3b81f36a42a2598cdedfea7b69ded27d850ea1806ef830771a6f729d504cb56b44e7aadb
zb91e83b4a3732a2402a66186c40e11435b6d48fda2b4ed37553049d504e6b98530d181dd93cc99
zb59fe6e9ab19a23ec9a09b408a9620631602d420438f27443e5650c9dcd1c045bcc23fb7822f38
zc4cd218c2cff5421f243c3c87079b1a79df75e38fcbb1780f4d3605d977b5bde54eea06548afee
z19fa4ed482ffcab3ec1ff0590a59a4d27239b1790eab67c90b4cc0229c8f79664ca43a1ff9fd3a
z8242f4915c478f3d35642bb93a8bb17992a27dbd6c4c018dcae2f759cfdedfb3a553882b0e5c08
za9d9f740d9fe00fa976467fc8c4b5c41d3f1789a05bdbdec3a2263b643dd420c960ac3dbc8ac2a
z0f072884fa868f522c4386c12adaa21199611a3b94a98c9a56aec7208359a14259817bbc90ab9f
z239c69044226dcc0b2ed08173de09b41815595b4e8ce11bd2723353668cae6b3204b2ebf276fb0
z0cbe1a04aba72d590484a59093b4ed13c6767e244cc5cb0fc10db96d1b473d5706ffeb6839afd3
zbe10633ff798f233c5426dd1cd49f1ac5c4ea1b141ac54e0197d4ff3e231c15ccd5d910cbd1214
z636eabe3a7ca2034e704e8ca54aa499164d3cb81d51c02d8fc1f7582ba1e676fc3aafac9244b9d
zac87374a40045ae5e24395b1f5b57bad2c11cd8ed045a1d9e818123a6904b0e90c4170f7c99af9
zffe521e46750dbc393082009ea94cbf63209bc3c226639b2f9fb478bd1af8d460da33fcc93cc71
z64036feb78f5f43128092eaaa8943cc2b3a7aee4d8e07bd3f52b5f58b3e0bfcfc4c68e9f9301ad
zb69c2279e4f67901fd33f117db67141ae81fa3332b8386f35fecb313bdcb6dae3bbef711602c62
zfbad021f1aba67c61895ff38eeee0004a0d2573e3dbb85a0c6b968286b2f6e59303854669d9a5c
z5f7af53ca830e0955996f6f4fe22340e64b52851c7c29217853cb4b6dd709f39f4143731c315d3
zad982b8e11383598b2871f802823f08c3aef3820633d23c32d70a04d2594774549eb3007a7ff63
z5360b06503d74f973fd2fcfd2f92c47c7209b0e6fa3302bd68b182351dd2c52615b05996359207
z05392c8ef8181bf967de6a52c88066504ae84bf8c535356e8adb0759083c8d0995191137e50afb
z4db8ddaf07c590e7c75cac1aad9ddbfba98ee723b39e537d7335614edd3f88a0a74062a1730573
z266f458084892e8130ac7762d839a88ae17dffef5a586787864882a5780a8bf84e1d9d75576f5b
z79bb767f4f4445d5a2cad8863984cabc48f7a5c42d5fcd9c0b96091de4c2805f420258605163a4
z20308a1a627d276ec6d4b38c2ca086afb28c6b9475ac3c41c738f0cab5eeff0acd0cadc889959e
z925fb7bfb06e004472d7b0f7c6a78fde63c261a35d8d8d26c5652d23b348b90e605c97e8b9af1c
z52e35029e64ccf4ffb533502bd9ab5808e11ae21c6626d37208aee07ccdfd888f3c5d834af5c22
z90c8c3598d0998e570946f01d5e46b5dd1d3effa4d8adc4a8740a33fdb542139d046f30a35319d
zdefc9d928cceeca53adf6a6774bd9d85e89902dfbe51a5eb947738bccb7f99bf34316e0eff114c
zc30175108cc647ad0a480e50b44f5a48a98a8f8f4d24babe966dcc90f006b1bc9e58386ec84aa0
zcbcd6ee9172ac3b838c4128c23fc0a43b49bdb84528ff6d74dc266d8e971f41dcc9fccb802a73e
z663bc8f4082a3909a563aaef6d8bedf2434fa536593f0b65c6d25e41e60e4e6e652611792b3a39
zd90f51825048fb50a04eb7b10aa7eaa2809f7ae8238bcc35f413522f192772b5e501bac3ab4c57
z8c3784f40dbe0057c2d33febf67f142be6b48753611a4b600f1894db0f2bc3b6ce60bd758e1e43
z90879c10f6d24fac0ab06d869b1a9e73da4647b0b3f64721d49b8f8d3d1c37fd8a590ca2e94e70
z98ef458f7e976018385d422d560b48476876baf8396b1abf60a0976a6b8d45d6197ada70b1db79
zcf09b280b171d1e3ed17ee66d66b760d5dba529f25fffd80c3aa5124468f642668b1137e544951
z2c07b5a0c1daea62eda6acb25830a7a789c41365dd4c02363ff2650bb8a026f8fcd0bbc096fed1
z3f256396a262a824e985bb449d01aba059bb4446d88752d4151f0729e7dcda83a10eb8c09f2d00
z036fe050328dccdee70fa59a51037a0f9804ab6c26a75840a8235fcfe426feb597620616d90afd
z81f21a26ac9851b655e558b9cdcb17cb925c524e41bd1749311faf761ce1631571307c658865af
z0fba987eab14ab99e5a29522c76e9468dcb1f24578d9c384d370d1a205ac3fc4804b5e3844836a
z8965a7fa2a0e44ed1af646b29e6d13b3b87dfcb69bb494c49f3013b89258981743c749f4ca7cde
z4711b87e6c6d66fdf05829e754fbaa533616c2f62ef5f8e7ab609e384054d0b83092edfcace483
zf8aff296296790085dc6a94e8bc98e214ee725113298c9daf29999783dd745a5af0d87318474ed
ze758914639689ad0e3104e1cd2c8d040cdd7bae3f73eed50c3b183bca59137422d41dcb44dd2df
zac7b278a812979ef5cc0fc5fe508cbda790751b9a373f0aa732c78393e297357eb6e827e147e77
z6ee86201724daf02615141034be7f69c6a01a847dea6d72b69351b2098725ad4e271f39d351147
zc289c4028097c794ca28a7d0a27e6c66d740a7b0bd8f58c4c854733d6c1a9e235a0366736a7f08
zf3beb978515ea6727e28598c086e7cdc1cd4efd984ee4834288c5b0b08c934b3ba07eda69bbabe
z71c24e45f53618f81104595fc5c67e7b281003fd66b0d78f52338710949de3966d4ecca8a4c567
zfc7a073e4f6c6e908063b1689fe079276069b88c8cd75e24792edd485053832791b1d19087dde9
z9ff1cdaa0843ea7db569a2e79c14bf4edf57a41c622660c64e562d905ed3bf5522cfe51599d319
z04bb00e62dbaba311e6c9781b61cc6e85b250625c3fd0b2507aa555e0b6b6443bbc96e19fd1c6c
zee73ce2b78e381c7633b3902b14e19458bf6f452e9c99cb7c0d74b4d8b37337b6ed5b9b6fef816
zd03815d6ce2b0d01318ce39e42f0e002ffbf4c0a93639a394aa59166d403f2a7ec4b617f119695
z4c5d82b15416da0d2d0386cabd79bf9796e7187a12440b2901d2ea3f4e668fa640eb60c612519d
z99f206c020fa672ef42b03d041055e8a3af7f1058403f839e9c25095cadcaa9aa7070501ffb5fc
zff51e0914c8bde1e7e7c74273cf4526fbae06c9319d6bda3b6a32cc1e2f39720f22b35510e2ec1
z310165bc52589be3b23cee9de0b219d0cd09f4c67334877da6b4f4147ae227db301f9a5a7cf529
z61fff6cbd64b0f4d4ae1e076b25e41aa2c8c538070c9f314598a226e0301f445845c14f403ad26
ze80a6d640291dfdf60a065114cb63d006ca03c5b30f7c3ce8475ff6382e88cf16706b2130eda88
z83c2dbe83a6aff71ab8b7ebe557af4dc2e2424f2e7915f99ee5c6079ae0fec894eefe1417aecf6
z2843eced2834f054a60d37ade7a897df78a62b28f942574312723cdd40534ea759b71b1646cc67
z355bd9d87f8d3cf6277cf83de176c6d49c1200b83b52c5459574bd5f300c4654e51ddaa70aec33
zd640675ce3619c13cfd09292f075d24c0558b85e0b2df9b3ee1abec469b1270333a7e0f09f0659
z7a7031681803fa5860857033bf5f06fba902d30a5a96bc8cc4aa312803ed65952b2814bd39284c
z340c3d30b57f50db1aac0fe05c1a6291824bdb8bbe3de3d263bb9c4d012ca661c2b2275c26cf1e
zd0495318b9ef2b3f9bbe1e83f701098afb1c835f37fc2de0c55eb4536d09f7073884649226263b
zf150be425c0b82068c8d0a629bc7becfff9b15fe0dff7e7f10df837d695867efae13927588a33b
z8ac3acebad5e91c312f3dfca9bb2252bd25bc8feaddced787b5db9be87f3110a5e490dd476b209
ze4e100101cdd378e4c7cf77d371c1499e32ef7cb66942e85ec16865e65b560c8e3de696570cfa7
z84a70fe63af0d541a0463048c07b29666797e080fcb19f7b84373982850d02ea97eda95e66c5e8
zaa4cec55caa79ddbd7be7692c3cbc075bd30b1e11782f3202a283ee9f5d30acf23b454d27683d1
za93194de31a8e6628f484ad0afaeaee84e688cba7d6df0b2c6118d08c76bb800df7475e4c695d0
z0bb1de2a9752d761106b8eae90e9168c316fc9442aceaf62227aab3824618fc571e0f7a1a2a399
z207160d50e0c0b120fc354d70475fbf69ad6dccca41e7768192e7a4b2aafffd30245f1d1e56063
z976dc85f898b8cf7a9b79cec31d6b76b2db7ff8726083c7574f8ca9ba88131f4f8d6506063c457
z6a1afeaad10e4f96e4759bdb7f05cdadf35b0b527f61b414c6e6abf14a22d6a7be71d136cbcad2
z00b4d1012fcb6566c40d6e2612cc30d1b2dffbbd946bf04d22913d812323ac6b89dc26429f881c
zb853ab5b6c4b6069423de5fe375475b28d2b8fc4ac2b34224487c70c371f02306d776b912274ed
z3220f9fef13f8cb775c9abfdf0cc9969195db24d9bf9d0e871eda3e5b44ffb2ad9c21aaa88f759
zd6ddb72fc264c339b03fd1c2dd17800c9e9307be2ba8f6118014f15718cd95236b33c2ea97db77
zf99269ff47b208cf7a69f6a84c81288f097dfa2c053cdbac15246215f8d1dbc9e0696d3240d771
zdc9857667f848783af49c00241eb89b24667f7986d980d217c98d8f275acdb3ff771eb72e82192
z8c085c3607a427e6caca1a0e4e801b375eeb6901ca81a9fdc69660293293dbea18721cdcdd5edd
z6b4dc2c8a2c41309eb257c5707f020eaf98050d1927041658b8b813f6a09ddf4825273497adee3
z6ff6433b88d4039596f973d2ad2037b8c6b7e89c7fcbd15296bcad8257f9e7c3a52f566814b7b8
z226370406db7263d77d26b87530990a9c643d74cd35d8509b5b3c1bb35ab5f1b4c01fb3ad6ca5c
z5680d30f04ff9dde64ba946fc9d034b1cb709fd58122425d93fb7a7a56c25be5bcbbdd4bde15c0
z81f07924a305592c8bcdd1e7b51e6db2cd913b428c53f882a755201a4eca7854f3d88f88dd76f5
z17c7636d1fba8a820f89225953b948e6e8dfaf5f5a810f82d67945b762b9ce2fb72738b4d8975a
z4a6fa890550145b4eed3d77e2a8471a08366f6ff69548b6b3fb2d07d6726c011de04c712dcda98
z0adba788f069b0fd1236ca51ae9598e98067e71ce8c1cd7e93fe55156bd317789283427fc40048
z2f5d2dc8922eb7cddd18d457b062d13ecacbd5635f7b64f2e11b23de34c00029ef19d3e28958d0
z2e59d5df1112d3b8c13887868f76be9a9fdf337900070f614dac2c652f08a4a962eac6d8e13e30
zed27312245671b0a221566ca2f456948d8eae2a42297132e21a9c10d20a7f6c8889463b52b9f51
za6bffa85dc85d8834793a030a91d771e584c6b430e6fd2641cf8a9ccc984488a06e61f7ce6e04e
z88bd0b84366373f129436650910f7748717d28c108157dfe4b396ee78a53c0ec9ce31250502ec8
zc44dae3dce40cb4c8ad6ee69dc312d4e9e9061fab925b3ba1d2fcce6845d19640b0613ec2120e6
z97832f12ec73ca458641a0d3928e81d59f091351dd98e2d8a112a9e0a314391e2ddc9da2a44cea
zb9ecedf0eab2868fccdabb1bcb1054dc7277168ead0b12b55c7563628cd52f0c5fadb1654b2347
za203ea5872da5b9c2942181764eaed77988f7a84693d6305c7624c4d671a70a7460dc47decca09
z72eb90aa27d3689a2d8e01460205db53037717c11f199d432e40e14530515cd6108f186823940c
z68d74dd87a50da38d1698cfdbda8a916c529ad1c2e3a43aac86b1dc6b36d6cd7a0be9312a2e887
z61e1d9fd8209df268126da68e68dc8ee0efccd678e7022fe842c8c9571b2275f36f87052369085
z8640302ae4e683d9dfec3e756d7ed8e451e1cc0344ab0f60911d16e962186cc6a63321429bcc1d
zace072b5be28fcc57dd951557dbc9f8224de7dc3799baf6cf249e75272ab93014bc89539b622cb
z25470306f69034f368492fd5bba24a4176803ee94c0a91e0e85afa21c7b2ab61277d88a9d1e7fb
z24107d7c4e6710b8c8341beb31b0baa4d560a4a6574b0b44d6b6c8cea0fab5a487a2462dbd781e
z46e781dcf406b1bc16a1e362ac26c30cdd5a80420abe2b80eb9a2f725ab94ba0a906b4487b0a96
zf248e40f2b1a2f76a05bfaa19659eb5a712d74fa531b0f3bdf8cfbf89b684c142da3c75789c331
zb5aa8ce81135736cfc24dbd2d0aa3f34db12355a9c302327f913f0cd5ee3e6d000bd189f41eb9d
z23b349a198fd0fc0aad0540c54522a3d3d5590f4561e1a8ecd8b864b728479be0b7e3320773d78
zc183c60edf42cbbc5b2c8b957f0b24360dc281ad5c866f96ab9b4a6504497cc790efa1edb2e275
zd3d82ca6208e24964c2f1761b401a4958b62749c4f249e8706d31248034e52022b2d81cfc8483c
z6df40d36b5397944942c329e6740faf1a53cf19682e07eff2af883a57519f1e07fde25b23d5932
zf3c45b40d424a624f0db1b24864eda237f03cceb6744d9ccf5062e49079680985a1d7311f7cee1
z011ad5259b5e544106bd203491345d98a9b4404fdb11016bf4518f6a2767c1621aa7546e7d2b67
za5f98400931c7785cd2b2936ed5947d62f04e1bcd0083602c412ca9d4d6d6aaeb4db6d463287e8
z2d65c7f166cb35d7b66e097edbdfdf4cc8182b9c6c4f31809305dec5309788aee944f409c11516
za63dda5b02d16cff3dc092ef194102433e6f3471a80d466d08f2a2ea4c0e694d9c5ec3e6ac872f
z5b643591b6b05bc17baac1e0ba4611c1c0019bb5f07e80e962bf44bb7237e9174d55fff67dca4e
z361ecdda6c2765378b7083ece60879c67885ffc2adfcfff969787c9f86e68066fecec6545a7d27
zeea8d1c6c2bb0129fffc072cefe7447c565d0cd7ca2096ca0029fc87889078dc162ea7091fae95
zacc0d83e36088c47f3b6481287b9e3b34f0043e3fd508ce25b45d8d8a6e02a0ea3283e49a819dc
zb05fedf0a5c3176bdaae35bdb7c83bb3aafe51d3af9d78359840ab6a0e95870cec617fdacbcd39
z1d0886eda75fbf0179e75e5ae1368a21c30c98d843c87dff6df54d5d40120371cbed619aef8239
zff4f64771972041edf96e3e2a7139fdffac181accb1abffd947864427f80ac5279dbf2058be336
zd64db3cb77038595e31028a0ae30688d16cd12004faf3240511f162a72806fef9bf529206abb7c
z1fa788f44664e56e70f69a40be6bcf42fd6ac74eac24d018119e9369d35c950c1eeaf4fa7234c5
z5c0b31d7d4b5bf5231870dd29fb187d0b2d877d1f83399f8a33964c5f5e28043e0b82115c3f6e5
z153fd2571b769c0fc1e4a140d212bf48248bc5ce06598236356635fd75931179295995759e68c0
z5e171ce6f8dfa3062879c94e5fa3c4ec53f9aff3c14e612028931ee9e6d61a2942aa55759a06b8
z98609210241346ce0b294597bf3909a799d5454b0617a929565a38c317777bbf659c1c02a9139c
z680368f6f38af7a678534587e663ce18f392af7ca24fc600fd0cf9f3e2b13274bab2a0d2b19bb8
zb0732770c97b2d78f5f24678f30549e22bf2610e4e084feab02df078dcf736bc5ca63fc31d429d
z9a603888b96915177d628222a0bf4cad9334519f2abb8b6e9b9df3adbba4afaf0577727940a7a3
z54c9b287582e093fee7c258dd137fd37a01032390466e4b4c4c207d20bb271cebcd2e40549c82d
z7f204fe731a06eeff2040e4f71e7b0682e0c729ca8429512c871339ec11d971ee6c88122120021
z4830a0b6a893ffee337958f818d48e518cbd0f9f83db40d6fc982363a11f5201f2bc6ce3a5e04d
zc53b2338ac460d8e046890a76f302d77d5f619fb68fe6c568545b791e538dbfd3abfe9c73fd98a
z69ec14281ca0d0e9ad0693db72be37284d7920937eb4bf966c8ecb4f98092ab8628e525af880b1
z2f3442a8cc0395ab36f5ca744333a79d8050f5310d6a39239a957816b54e2107330e9e490dbffc
z95e44c9643288ecabd02c039b7dfa7c8f6c88f6e3cdf843a97c869f3ab751a3791b5df62887b11
z55a46d39ab023a26bdf1da4553ce31761e97ee0954e1ae175d6ab7c0f3974d013a6d220aa1ffa0
z5a158bd9502a482e45f1bd79661eefe78b96a683862f5ea8c556f2bdf1d4ce92c59a2596d2a784
z58c8ef6185d31800bc2f8e2308a20bb63bbae7c964d28153ee941843844375274e09ea5430e04f
z609a7320142572eb186299e292c26836e384a0fd11793a2b527292215e7caf64a5878d57b69b4f
z4bc6cbdf708d1a5d7cde4dc55d3536ab4d3a9a55a63498f455c4496f544259ad2f703e9bbb1aa9
z730ca5576b6721016fd8f7e0d9e9122673c7dbca6ab0c8030f3040c860f7679c18bbf0eda05b6e
z7e4e7fcf67d4c87454299672cbf2c722bdbc7b5e981ebf15632a9f4aad2c5d5558c5deb55f8e85
zfa1d4df06d60a4c106123c14d4f16519d389926e7e00566eb71b2e0ec31e6bdc1318f123cabe3e
zb5d216adbf948ecfd9c37b1c3818d625a23a1f5965a08ecbe64485194340efb733ce2484ff56a3
zc6be51d76bab17c4e097ec2dc9bad1f610db92538451fd5df97abf78cbcde08a88befb54ca6e62
z5f45bbc06fee4419393fa3f7519d3ab549ce680337dcd0b6a6a7da064ada8da576b8675feb40ee
zad1e25afacd19b89fbfbec1626d5e931473a418df1503dc249988de1abc11baca925451dd001f7
z64fc3018909b1076ae45e5e4e3e8238a784ac22298adb680b7c8f3e45400bfdb54134edb727290
z5a91420102428a5966cb10e7a60bcc5a1c0f6eaeec4c0f360145f7fdf313307217fbbd3a250e8e
z1a51425b63bee22f9fafbf14df42cc7cf0404e2e3cd68f37e5adaf0cc4b54a140f464ce30ba36f
ze2c8c8cc93e54aeeda108071bc08b8ae866a1019d06397b7c1058f7abdb3d20de996b7ef7e94ec
zc65faa9ad77ed79513b43dcf570433069e566a624df0e85bb88a20d75da6258c2e0f9ec242000d
zb3c244bc4dd66fa8e880f154a64cb392803252b3d6ef76398ac5ecfa848805f6ecf99b65834ad2
za9afffffaa1df90137dee847c31ea149b3a6d5e00ef3186931254494f5a9e66c90d2e4f2463417
zeef85ec761d431fd4f728e7db545f431d638b539682d9dde3e5ecc93cbfb946ba893358c173516
zfb7ae600774a391b36cb6c78c21bfd5e51cd62fb2d3476a22ba55c3cfaecbc4a6bffffeade2362
zffad22cf9d797f0251ee6817d8d098e3685a9dac9364c569d33c9db1e8e00799c2731d2ede2ea9
zeeb762bdc94245de0f18a571c7bf9b35184a85e5d212af74adcbdc89a07f24a02666206b17de96
z868730bade7ba431ac0d6018a5dd2c6869d88aeaf8b10efda6f6541020b658dbe59eed4326548a
z6529037dd98e0b0e18707a9b68bd224591aefdc12768891703542a3d369bf50844e89d1e5fe0e7
zde8a98a937454974efff8df1b384036d66db562b9d85f90c0cdf45bd55b23d9392a670db464ff0
z8093b8f13ee0421741508f3df068b1762f74072a429407ee273a08f8e8bbaa48156e61c01aca6c
zc5ab25b13fe5eec2b427d502c6949d493e0a12a5811a9084d5d688f3554c0d477bff9a9fd8aa9f
z1923aa87cbf1f5932e89fca59ec9aea59e22ee3df068543e992ec24122ae8c230ace5eb62f1e5f
z53774169106818441b7831a8d6fef22de063f861c6a1f982c1fd9ba906e2268c12d42b25032c44
z797876dfa4dd58f68d707f8ca3975fbdfb963e254bf599e13a8b95476e331abba732b42f8325ad
z7df3e818947616920c0526dc8e5d4790f60ea03c9ef4fc4c0af1bc0cb797f99496186ed96fb6c8
z3d429db973efe36e90e764638671c4e7e0aa7f6a5959005b1415dd6b3459515a2f3796e4a4c51e
z745bccb2aa3c545d4eb3f7c21b879ee45cca9eed04cf7a79e966caa3f3596fe0a6889ebbaef1fe
zdaad59867de028741dd3412e49947bdd1e2b0edc4ea0cf616963c8f408cb6054ec2429a6be7a2a
ze406ac989a59135fa86333f5527afbbc7706ecf75650fd0e39e6e5c72d1e67071899cf2f040125
z6bfb7d703a7926aece8bbaed98007897253358a19121bfe8e85d11c46f76a6726fdb68ecaac75b
zdcd2b50e6f40fb1a188a9e71beb237919674f06c46996c6af1090f3f094ee788faa2d38c031e91
z8cefca846718fcedfc87c5865097ac118d6008e1625731e29fb279f3c48b102cad9c1686764ea8
z27b7cd72a5907d2558fb13991447fd4232d43573ffe60bc6e6d8c08cf2b030b50ebf9a824b48ef
z9e6478ce0dc5825c0d4df5fa83cb8f444a32fd775b909ef65c14d10c72a598c9fadc3d9445a7b2
z798c2d0ac1f594af2e1876c69f1cf3c8330d0ea871c936c1d040c4b3ad2e6100cc628525ec651a
z5f9084f12e75bdd7e5f58863642871f560d873362896ea9b69d6f57303d5be0432750e1bd381c8
ze2834f18f5d592be08998a8e76285e0cd8e8d6f67c96ac407291918db20b130fb4551a2f66cecc
zd2b4fe6755817f9f8e9f17e28c48e4c52c23aafaf4d48f984dd90d19c4560f9319c7b7ef80553d
z8f58494d2df97f8869f9779daf34bedbc01a5c6fa808b1615e7776e9163a8735203790c3354a36
z3a459724ece99569aec81470cffabd15f733caf8ac61af176d9f393502e7003d5a21decb09c145
z8bc85bc6f4ee6269d9a0b24a369dc357463045dfd9eb1e098e9e4d26b96a29f33b78d6fd17d8e3
z209166d52ff08981a3f740e59f5b573082b202ef01e7e4984ef4a8782670556d99f30e9a2411d2
z59781e05c3aeb8db401f8b7cbece785b9043b054b1f610ee064fc18c08378c8231bdb409380d41
za90b480a9e298afe443c5a8917d235355b8db610dfbd1a22714ba7e457d3a7810d00b900a34740
z5a0ea51181f2a0b3a596f99d97373608a2efdbdf12a030e248373b4be5d08e8d1b529ded0b29ee
zc31bb32c5e1d8a6380809265c263c18183791f2814073c9a94f99d4f8ac704e6ee9bf6509478e7
z0718e933e961d2d3b8ecabb24fa22f3eac5af50d765adf810836dda33ec303c7c65bfad9157ecf
z5d108634bdd7335dd2201984129fb8506e3893e22cd6eb3f5cb6aebc12fdba888cd3ec0b402c39
z8e2b457b55abfcbeef2e2c7996fa861693f81de5897dff12f1501afee9a7d51eb04a6fa85e66e9
z0205529f0562d6f4368f570fd7db8a66e6d2cb94a4cf6aa3237f5a8c57cab03511534364e18a79
z0eb3dc374a7c0eb795a514b59cb8ddcbdaf3f06efd3593853b3232b46bf0feeca507e47c6f5bdc
z1d40bc3afc50f8e75767dace926f4aa6f28c719d2ed2ab352778f4e0adee7dd6b521e27089ec20
z279a9a64144ccb1c242d9413b946dbc2562b05d068e5721352688fdd21c20efbbc0325355cd2d4
zce19336f52bf191c636ac9414f0db7132a0232102e3f97f16270d5e2b331d6f5369a382bfaa0c2
zc14db6b7536bb6d29cc5a2c5064c561b9a21e9b6a53da1e8a1e2e70155c97f940de67fa9fb6668
zccbe96c48b268b6b854f3fae6abda595db0f2e5bbf6c209a2905e764552c1da7cef61df369159a
z4384108e41741e437486c28085bd72644e5e0921e688fcb658a45938f5fc3f9ed6cec686096921
z28f68635c7bcdf82fc7f866bad365035fadf165bc0bc7fac7665272b2184c3602491f22b63fe03
z65874e00112480af0d83c8cbe3ff580aeb7608fd36e67f951f9281e5e0fc08ebd07bb639bfe1b8
zdf880d1cb52110c5545765f8f904896fe41984343687dc73e97ac4eafea2589db0583376c6f4d4
z5b483b46d5a1f21e3803bbc604ef41c3ce104eaf5720ea1858dfa85c45c4bc41159eddb7c5d8af
z70750eff7262f97f0cd6c6f1d93905204e4cf3339056dac44461346e440cf522c3eff160f79178
z3a853564f679e170d9ffc2cd072763991a21e223f0837e2856e10b00421d3386389b6e1dede4e3
z5da9a837325be93a34bafb5e249111354d339d7de103b4a011ef4b142c9dbad31298325ae52147
z70fbe29f172e6fa5abdaf04bfb0e904e7e448e670896d3f8e9e6235e0c1a96d71f256f0780817d
z46d426a0dae2e9d632f1631a5f40f6c42fd712b28a72bad0fbd85fa582b661e571e097c7743134
zf1571dbbb29171a2f9b9d03fe5f923271ecb70381e87c00262145af64685cbe00c6f2ad0f1f172
z45258af212901681385a9b71bd318e295676838d45009e2001ca4b70569faf5b829ce04a4396c5
z0a01d615a046d2a96c9b181dda6fcea255ff621eb70d0f165cd846edf195a80bd16f2b276ee059
zc325da84022760653a8eb6f3d2946f38f647f77388c278cb5c474cbd003de371e71bfefdf30b4a
zf792d922014dd50148a3675bf2bc6616895cfb13d3dbda17ac1feff749144aaa9579b55b8e081b
z5f28a55329d1c9afec5a061466488b7a0d77d63bc999cfc9b4925bcf5b628247b40dce2054d23a
za40503f0857942f4c07ec773fbfac0b4b2b393c6a0d5f26168157aa90b1695c58fba1abb058cb4
z0051ea6f3724642021ea2ed51f3fc13779a436c3fcde50f79b2531e211945019a0ee833f0efa60
z23d9553fc6bc990457c438f27ef4c374eed8a259ca85f269d49fd58e083bdbe49c3f0cfd4d6f66
z03dd82dc33ed8dcc2f2200683c4bfb5c6b8ffa56c3e2bbbf57b847fc0ecbefe04d9e8edf529bf4
z2fceddcc913d8f21db0b167eb2d3336d1c8b0310d89ccb7fc2a63f0f636f5e1aaa365eba81b1ab
zf7c7c6654edcc22b59832e3b9974c3d9254413b15db8ac6c04c9e8894a1571091d60dfd876b78a
z6ea756b2d2234cef005fe87c8211f30764f2da73f00642c6b759ea1542ef33c6b87427e3c554df
za61f769a8fa1e4f7c6f077c8e63e694dc9d4db7e82fa91ac9c95f410a3ca336187448e26aa10ac
z279e9f6f1c7614c07b46969dd3f54d5049c1a1f1b51849ecec61248376b0899500f3c30e053cfb
zafc8d7d0486fff82791547b592fa01a972fece2d4d5a8e6a607dec656a7748a43101f0a86883ee
z81006c560ba080a459a4cf6aab74eeaac4b88ffc8fe967b717dc37ba19d8efcc38fbd37daa2ba1
zf7988c836293708b79653ce6b3dcfd705e21dd563cca495ddb08ed6dbc9dcaf0b2116cd6efacba
z697781c44cd4fc08545675d06ba3c371438a183c4ca69588665daa28ebb1476a17163a201d5cd3
z7ac7a599606e47e54e714a13fbb2a1397ede6a541de21553e269707cd989649bec5ddd44c09824
zfb864ff33914c57facac31b032e38ca66fd0bd45446932392a46d3384011246796e522b6b62ea9
zc5444e31cbae62bb65981dc81f7e328f29f51384de93dc1b4638cb33c0cd7c2fc0311b682f9db2
z6163ba824a8635e10380c634d517e4cc1f241c23afcd020920df968891301a5d3b205b78fba43d
zacb1ae4daff7e6909359c8682c1a53a66f1504c9e64e0e28f6e2b3b49ef2292e6c83f8ed8bd671
z05bb957638a01b554ccb0d4460f545aea738bff7baa763b99385be50cf87f1a7718f528d0bdfd6
z6d6260e0db3d535d3d4f9fcca22cfcd992531a958460def00317de1a951f14aa513d6bbb0b3072
z48c3b8724ca9a187d3a38f8603e6c440e43e4de2abfade2947084aff7b74402d67791c709c2eba
z4146760585759a1d74dd863c3fc8d0491714019c766fb87593925043bad21e513ceb836951eb23
zadc853fa109fbc744115de97961d217296fe1846a241bab92aba17f8d70f0ccad382ee2dc9fffa
z66c4b630164d7efa4e2e9a311e81589af90a18ba54838bd11b2f36174c57a1677b9352f339db2b
zfe86e70c43afa58a930e5309d466e355784048a4d43037a36b2f5f6dc5409d6215e557090cb20c
zfee4f68c12b42bbd5f49f22355397810e1a419b633327135934002c3ff376d014796abd3904b67
z77084ca45ef1a43bcc0e88b7b7bcd3c1c5938cca5f8ef16577d12ed345e87d2bed379c6114ed36
zd074b0958a60747c43a0ea9a2fe433b8cb7b1c2432ca88f8291a80a44c3ce721e375a1c407b9a5
zf90be4bada366993f66a21a7dc45aae912131034431102a22a9c99865c928990aac8a658ee5086
z79d84996a746046e4197e2344487911c27b7057793ac961bc0f30d5ec4ed5ab55fd96140e6cfb9
zb601c149894f49fe7a51406a86974fb4804467e772409ab5059a006f1a8c2ffed60b454aaaabc6
ze20a1e7966e123bcdb38addf2805e9bff2f7041ba943775c2aaa73724fcdf9c460c51df881db1e
z746c4dc2aeb706427ee29d69e6468686bdcbb7a5f9618e9e81f51b85de367b4555a1c0b220d240
z7ded1b67b7d9b02516a0f9f59eb3b4fbcab15248a42ef65b113e7d3c272dc4a7783f29fee62c2a
zd1ce46208e9fab4b17a9ead92acb63e7c0b14b8c5adc932e7f308887cb3949a9eff2b3610d5ad4
z878d06438bed85ad73f90ef7b89d3d1d41c73193cca413dfe9271e37c29210ec9a13b2ad27b0c1
z4fd950e74b02a025c11fcd5d6265198e87f765e29663f46454981b5fe4595f6d5055487b431a05
z4aae5102f4f9b13363e1130c327dafac29280b6a8c229164b0d7889d672e15c6bb3d7966ae1872
z026db8b986f373abe585bb87d9b2ca4771b606e45c0edaa44e6f2d557d3092b558ff2424a92543
z57fd7ba8b300bb277f03964485ac6416bfa1e06221a891e27197c288748f45f63d3ba177c97b7e
zd8a31e301ab6b52c1cadfb25365269f5970131bea04811e52bdf71105a6d6f410ca27b43cdb27d
z96bdf25973688fd81d5e586f3d74a884d5916ab77894a4b1563d4d413d67ecd65d5afceb504c7d
z1dab874744218b2bd7f76f9abda37f382c5483fda134fc00a3f284ed3e69c24e07d21606de2d5a
z27c7032fbb201f88c3ad2014e5f50231c61e8108fba5531201be55ec900f3218aed95c9e4a8f8d
z233ec89126f9f5cfe0572e449573b45cc42ced46c1389334147089c6672ab4f887b10f1c984b16
zf71da63eae1452fb465563fdb60ec5e9409cfc6a6ee95c70290458f5779cfa6e96fdb7d3c12eca
zbfec03fd1987913e313e2f857686ccb2cf531aeca2afce9740fbc7b115fb78985bfa389e24a4ec
z2aaef6711e4cdd4f03388a6a3e37d63566ffa2b3e02073b067d08b49bcd8b0cbb7a440db70a19f
zbf3642ccac64f8d0605e2cc418cb8dd3087b5fa7777e6b98b3ffeb38461e7373db6e73f9efcba9
z0d4813fc3739f8f42b287117a504cd94a052c43709fd54aa377b878e86b243a6ecdf860323f4ba
z294804706a5910e968db9c21452f110067b67bbffdc009980d2cb497596d71c01e9387cb743b9c
z45d598b46843447c067d8797ee3d601a4d65684dea5e8dc8bf69cca4111ebe2e9c5d29ac3281a7
z1ec2ef66ceceb2a0089eb224e5b440f5e01845dbdd34adb27b4d72d354a120c2d3dda403a33e37
zfb4fc484bb7f4c65dece4cc8ed861801a3b74ac51a792b3f45e05d1ec4d2f7166cfc66460c1e2d
zce61b99825119369d52d23fb588f40a97130d9a0cc7b1c54f811cbbdc6345f105011c698bcd34c
zba10f02628ac32f3f4a4b773058fdfc1b7f3518dbd22d8360b2a2b3e3c64b16ba17f2244c6d2de
z4abd5552a492c0a5fa4d0e8a7a13c1a21e5e1487f0bc8ea28eca8b16bdb8360310d3d1e3dd4310
z6a672897c00a03af49e5daba18f266120d22cb49f5c85bddd25d13a0bb281c92ab1cc95b4261ef
z957989a76b4e02abf12b7f510ae29bbd2e822a89dfad034061a4c2ac54d9333bb4e7982a07a715
z27a21a32f0e79e46f094d840657d87ce07466990f975ca901bc9358f931952533c19737086dbfa
zb70586b4841008893f3a8e2fa9caac3b30861a7a610279e20559a510e3429a3e691a992225441e
zadc3a21e313a0be5df781331abc88f46d531c192622a3c267f49e6dfbc1abe12973cd73901ee96
zd421e1573fbc8d3a8e786682cc245330d840e1e5378dd4cbc959ce69c3e492b483246f75855b01
zf8fe0946d238c98965011983a0c918b86e83debc02bb6eff15918be21d0f9343f3afadb84e4d32
z58fd6311c36d6f94000bafe122e64b3d5ca72a88658962fc6c62dff26bed3946ebd17df1c93638
z43b2758611c4ca5fdc9771e705c0709f9738848dd24d7a4bacaee9d8846606a840920b850f112b
z228cc2f3dc18107330437e28b0753e2019719c7f8734848266b7b7ed07df5a69d504e9594f669a
z753fec3536d2bc19c7d7b5e61c070b6183358acc8197d7bda7317a60c379a69962895b7563e044
zbb52d3e8fac003e7ed81a52a71c16ed3601f01d115676fe8c42ea9e58074033764de98a18b921c
z86293cdb14a39f98ca0f316356ff1fe41d400b3bed1a3ed7d4d126dece0f74237f00bb161481e6
z073d160382d15d221180751f105418ec9f19c7d06334c0f96ed59b81c9d868a7f073885dee14d9
z60d0052a9e0d9b8a63428c6b3cb45d8b33c423232882a9cc3a6395ec6a39a6391f2e05d7e04e7d
z55cf5e326fc76ff91e8e9bdb7a37d69bf9536dc3fc3946ceace490f4d6b8bf9df6ee78b47ca546
z45ae20c903a1647a83289e319bb64a88401f2b2f7eaf05dc68662fbdb975640630f16df3f5a0d3
zc28cf4cba41e65ba196cb1ffa706233ed2fbc4ba02e5e57a4b42ba49c323d36a507f75081717a4
ze5c028be1de44c84121f3538ad0f0e7b70579c7939e20a839c25d8e155367a2a64f0195851089b
zb9dda958d255a20c46c5203ded2ea13158bff7fe6d6f6bb7e11d7f2de56389cc8cb9481ef4a806
z022a113b038760a2e019878200aed301e9d1a7f4a1c8245b839ab7408945b00ca98371b1103768
z94443e4d3f20a7c865e7facc8d08fcb89cb079180e7080af4fc02cb1c91a2687a75bc12349d56b
z79dc84b38d0870367bc18654cb571d0656ba079690409ff1fba995ff3a2781d8dd40db631ae3db
z4e389a1c9441a1d5f9f036389e4e42903cb5ef6c2c792e2fe4ad62462e3cafb822dd789e329446
zd46da2b9931fcc9e6f847d19da13c42a25517c19309a53836b5a423df714a906dd53775b6361a8
z0d59a4d0fcdfd9e37a0e3fe83284ab4fe290bdcf662fe6c8cbd4f5849050bb89541afde329cf79
z962f3a6062708d05278b83420974c46dd64437992325cf046c66d6ee9f3afacf8866fba6c574ca
z0a646cfb540faf395966dec892282b297e12e74791945674b56fe142e568557d9d0a4a4db178b3
zb2740e97c65ca0c0a1b812e10a4f97349e183618ca7d8570dda4a0bc281985130f444094322fa6
z1d1786d872c918fc7583efa152dec5bfee6249c1545fbba89becd255b403fc024359e6235fe52a
zb8474ea4a0e147465096e8cdc08e8aafb95ef0bf7ae603f20f19fe67195b0d11a3d6a1d32c6d2e
z062539057998155b433cdcaf608b2cc358c1febcf1ed162b272c3083441450265f5b028d205c2d
z82154dbb88b22bf26c851e730a793bff6241859777f27d791ffedc45dff8f3612c4908ee60bd67
za66f9c214d85b36b591e3faf21bfd4f564ee8a7213fd32bd967f59b5ada2cbae72df3c60b5f6fd
ze798b8a04cec178611a921ff584ed1eb5082c017443e60638167a53d5a80f2f615ca794a8f587a
z55bfc92c22c1af35559276316ec546509eee7a592dddfa5b2ea82d3eb380149b0894e05dfd9735
z058125f413b46b42fa735a5c241b77272ec8adb9bccac939de5ab050ae49c8b1d5029ed269fa3b
zc0baf9cbfbe9802f12d5519c4f6a577fbe9bbb3308f56441949892ba119f98d2214c426d63a834
z9f348826ef4069deefe67e6c6398342d5e937eec8af19b15aadbd40562dfdbad04af04b38e7f81
za9920e72a94dc8b52e7d1782df08f7bf278a4409ee16ff7e07553418228dc11e470d8703df95e1
z7ce1d7345eaf43cd1cd2fd3cab8b5d26042949ac6cb0fb255271a77347027899e62df01f1b064c
z72ecc32486846b223d55b2ff96ee88bf23625861275e7bff3e1aaf4abe9ec4645521e4ee4c0383
z3e233c65acea9bf5591f527dcd2a7d8c536ed642352a8ad5ad1f706e1574e87822936d281e7ca9
z44516e6ce840c0ebe1d8fe8af86b1dd937e0f38e95b34bf22e6386a71fe7293c477658bf9f65ff
z39054dce8762f205bec44a5f43d8a0a488a09d8fb7836a4e927a67c09477e3a83b3745955dd259
zcf6d1c680abb14bfda958d01ba1474036fb4604a60db8a91cd80fcd281e4731102ff7ddb5e7bca
z92e36cce46698402f722045ef0122494659150320b4381a890a31ed44fcae4e02f2e3183089213
zb239ac90b5e88d7c633d57a8cf817f85f0db0712e37ab30a278c1ed7097f3ad61ea268649e4b0a
zb149ca215e34cc443ac1902372ed8b2940f0061679ac0d6710bd11771203b553e8a9449f064ad8
ze6d41b80777f4fb9eda6e6b14f3af63fac5ab95b3b63f4ebfd50fec3d291f257d57b585617cd9b
z57adc19467bb95777cefd9288f2a7c7f7b2b131e264d233c65e556121c0dc5884debd8be0fa57c
z4a527bf18e3221166454e8d7b7c60305b4fdb804549d70a9b5f15ef1806b031c54aece60447e79
z970e081e64f569f3079072bb4cc20daf0dea50f503fe77a917e9eaa4cf419127fab0efb5af03e3
zbba6311c06833391109ecc27b2751e0b1000612b56171ff57638a46364d55bb50b697082e92ed0
za2331f50208f1d3b25c534b877f204e4d96cba06910e50b1cf287837499e30f8c82b037b4fb13f
z22f3f6f80a30c4deb500b4274032eeff797558b71126160b23ae28f02ac47868a5347bd04347ca
z88d12aa6b5eecd5ad0ed58f3129d95b70072ee1895a6c2f9cdc2f543def395ac1a828975b7dd76
z65b501960992049f519eb55cc87332398dc5b4f979109989c201a9f5c86ee5dd300265183e4927
z1e3b4f8693a145a43e17502216d99d5c78014b1518cbe7ad5a580991fc0bc98a7a32315e065b13
z2b05a1989fa209de58504ff81239318bb9747e8419c0ed63843193c5e80a5a018559cb5a03b3ed
z1931d58581ce3bf7e54f3c489bb705ec4c206d9017ae062927701c1864ef1e047bef574fcf5582
z9f31aae1d35bbe536149ebb8418686e61f7ea20bb5f0aa96e88840b0fb2832c2a005a14bf7c501
z3092099e29b33b4db78c10e0db0c9ba48c66bb49617d41f24c6399f752169c9bf9d0def10c252f
zc0a4ed38041ed1abb6bdef9fbaf57200d0caeb648fe02463ba5dd784d5353ee238a88cb8245aa0
zf950e1210e958ea96c0bca963fece390e64dc0d1e2aac49bd51724d107b4ab8def5ed8400ce3c7
z4b3af50537d66fcc927bc55b29de44f095648d3663512702fa8d13b2d2a548c7110cc470c8296f
z0e33dd8547568ec55fc55111fdf473e7085d24626a3c1bafd06bfc798ce7c47263abb4fc28282f
zcce883d63da8898cd90de08296e9ec2864f9355b3c437404028d5989f3214e9bfdf79c0e63cb67
z9b3632d1aec1f2de7f232cbc9fbcbb72ea27925b62609cac9ee221eb1522b6831c1b411300a330
za5ceb4ab4168724105165539a607943a52e7f479805d6fb4a7a432c6f0571a677c6cec90e32fed
z014be3764df6fd954079b445e4abb16c2ae39655baeea02c476143feb4f820f07d7671f04a3cbe
zc2265c96a245833d2b688c3db290c588b16482bc129e8963b12a70b56ac10bf2ec1e4180a4168b
zeec8992892bb6b908cd44e3d1f116b9bec5b2a07d96ad60db8d864e2bdafccc18d30e76222ba87
zdc99f32d2c585b608ba4702e4fdb4a755edb5b81facbfe2e764ac3c4c57650a5e2bad64025cb98
z4e9f8017e86aef1741ef2a4335241451a6113fd5fef31e91ea05e4c5fb42ee981fb462564edd10
z375f8a001179b9677a2a0749220a50fa71d88eefdad9014a269eb4b2ab3481bd4acb69f1f493d9
z90a0cbaa3b1039b906f70af1a33c7a8ff1daf67dc29e323dcd1b3774e39db6ad0193fb20099640
zd1fca9fcc4c0de7a67f061920763bfad69270467ee95873eafde2e3f8476d22a2a76de2fe8a62d
z83aa4c1c69d2d9b32c26e1259b215d48a419f8caeef587cce563fb6e2e4223a7034a7a0539d440
z533faa28af066c254c5c05037c6d05246c36a43ad5974f38c4d1a68234f059acb6e497ce744741
zbf5c4623e3aad83b70666efcbdb9bac55c9b33e91a224a145d0aee2bea44d04ab738d6c0674ee2
zfcc3a7be424db63be782597bc3f0724fd617d7a276714e4fdee021d2bea6fb4e60def5a482aebe
zec7cdd0d1fef5f9694995947e1cb9985114bad4cb3dbab5830e676b03565fffb3b19dd8d61c376
z778ae2cfe9164eb9bf56799aea6ef4743ddbbfc382e3e0198283789cab02cc5b30ebc25444504e
zd6728c7bb29b34d895b52b6c0be74cb260c654284bfcacbfdb8b2f10a22d712650c0d14dc380bb
zbccbff98852162a4ffcf394c664c2ae0e27610d8dfbbde92767a448feef0b53a8e048aed1ff6e6
zff5c6df48eaa1bddaa17f258cc8882115d56c5339eb91e788cad00900ad559c6f5646a936f795c
z39925ce6faf523f71b2779e554309e858cc69ecd5cd6a441884b8dd4496140d21af4d2f7abe351
z92b4ccdfea3bf43a0c7be542121339f1c474eeaf87c89c78831a1fd706ba8cdc50fb8a5be7b979
zce75fbb534b2ef7a1db37863468d38e90c641e77f61768df7d7460d64d10cbe04f3e62f4109ebb
z4063fadcef3496f167ea120aeb6348878989568e167d9d523c8d0b996970e94bdd1c92b11624c1
z8d91ff9c875a9e5fc441da36ed6509b3f76e98483517c4378c8936dc308ab9ef519e5bd2db7ff5
z9bf4105653dbb13146bf3aeb29c571d883b181e0d0386205d0693d16a2689fd87b42189c868ad5
z0a7101c69f7ba8a61079a296b4f61371a233c419999565c25cf77444fdd0eb28e23b3b95c386fe
zd1b61df372c3a0bf8ec64fb68ff94a8d2afaef28c9ff2c28e4aeb28c730043f934cc01254dcea1
z525aa722cf339bb95b12f654eef2ff5b82c228ec1980273af756841490eb201b9dee913677751e
z3158a705844503ec5addf409754ea6662354420d60265ca5435d9d689bac8540f24471d7b38100
z2bf88d0c6aa93f77459f579d98194998e30bfe3633cd61a218f32418a57c2fffc48d08bf2361d2
zb1676b987ab7b7cc95bc4de3dd65ec45449b01a7eea42ede362e0b356d82a60bd1f9d9362c990e
ze7e65a60b086260fb5e77b64d009562efa5a81429542a3dff52b786d18d3d3a9afabf988456bab
ze67471aa581a12b2ff393b90beeccfb35053ef863c8923de8294d513a58daf008a5b530b451da5
z62e68c27e8505a7ba44ca5a558f7dae9ef3c9be0cb5564e61a5bdf4bf056efa37c95d0009c5481
zcd415de8701ba559e80e973c5e7394ac875252d4462f4fc6007a11d1443187dad328486a196d34
z429486d1e45d34067cf81fb1adee97db7232c7675c40f6afb4b9fb4358d08d76049fab45a9b416
z29146ef0babf976db22774bc49b505b114fdb8f33f341e0dd61e158afa6b5ded6741f3bcd075b1
zc3b10f5b153262eee6d1e47dc3301eeca444d244f026dd2a023cb20165a107a49261b8d1efd452
z3e8de7b84f6356232e8d20ef5ab1e12d8c9df03e103ceb1173b47a42917b34999cf794d6621705
zdee4a475d26839e1d800452853b99c222deb159a2834b9ae3e8d44e55317493cbd25577de94c73
z3b5efd9f7a7dd90a4acab690817a5127a0943ec9eb5ef2b593158ae2908df26010e536cdc87e47
z255ab2699af64f7e5207f68bc33f4e103dbd073946e87dcd33d6360efabfc3805ac9ad0aec2565
zdb514d6f6d7554384d2796702fb1e38c3556913217ef2a4d036a26fa54f78aa3db1f1b6b32b4e4
z085a2ad78d11ca45827612ed9fdd6e3d086cd686a1e1fcb37d44b719b86d19a73daff9a11031de
zef329d01f841ccf2558717b2d14f5b420348429b31c29abfe3dc22756a879476633e85fdb10d2c
zfc3f2ac6bbfe95427d641213e6caea5276d12cdc79a9ae23edf1915cf17593d224c02db4c545e7
z14df4324ddf5ce79f9e7089a6d5dacf1b5d9cbba0d2c6e115f7ea9110dafcc971b48322768dfc8
zd12a46bbc36beb71bd0589196fd00e84f2066d8bf8660cffec448d60c52a834f0a5c820bcead96
zf682e0b7a7d12ccf2a5109f20468433b326d3b15ddfeec461bb650c7051101488f248933f944fe
z409ace37e0247baaadcf4c00d796a0fee0125b1c84888b9ac6e39102bb094bf87ecdb798f48ea9
z3940ea46d3f725ae8795e051008c165b47addc266598db46ecd38b8c23081ba28598ffba5c5d51
zdb53e9f9944af2a10687d96af29ff54d2c382d2153823f70f6f8a0c9d8ea55649fd250c0db460e
z8c31e4cf7fc02110c33a0613a5f8ecdecc29f1fe10c54e0aa295698c1e025162feb92ae0b0e6c8
z2c3728fcc7da5b3d488fbb32fc7363787ad58054a60e148ab7fdd4cef19018afa29164169587aa
zc645e648ace185d727edd08f13f4f0206a837376959afd416ec40cd42aa635d24f1c8600c02af4
zfef648c897308e05f62a6b5ac209d566de0114601836ac12e4713378623d4edcaa0f446ac7ef08
z3a42d7aec85ecd5aa8c20a0f1816d21e4e69643072c048c669cda5500050529a66b8793340388a
z8136d747927e964926b90b7be361fe9c59bbf0fe770f049d57bedacbf7c240abedb936c3cb85ca
z3ed76476e51e644c2e708d2cfb394bd6acca82c90bdd1a226e423b6d3b15ca0ea1933bdcbadc41
z5200241173f905a4f48a281ddb672cbfda5c21dc484963fe5bc2792591b75d251efcc8a099ec5d
z87dc035082f2caed2254df173f1bac74e27b5fc3ee224460a10e3eb483115db0d90c2439091e5e
zc6e5167b8de0cdc14be74e214adec11404196cb8cd4261bfcd9e28f7e5eecf2cc3681a8b8d3e9b
z4fe754e1867f2efe410e2e58eab8c28426a0003291628e2678280eab56e71f799ffdd340190173
z3bf2e0c52bb574a15b1a9e0e6f18c858cb5f38fe35675a78e359d11fadf03b1fcf6f6770281857
zbe027aa5f66b870f5bfff79817b7f2745a42e8c51ce84588c8c8626682c692cd2e7d33f2125082
za46903756b9f779c358bb810c1216eb2f8fc47a6bddaf1b82697246f82e23efa56d91172c44d77
z5ea6e42ae48d991f8571b8f9a3881d38d955105f167a18a541a0ed9a8609998e1192e27422a056
z9828fe5507f520bf7da6866e9f5e4a846b7a8d6e9041e0e45bc07cacf452611759c5d9fe28eec3
z33ca2f7ecb4d0e064427b157ff4ed4edf5b2284b9a36f4a8e2eef113b68214317fc05ede53941c
z2c5ecb0308133f7ca063c19a0ac1d41e626be9c6becf2d385c5a6752424184c0ea6c5e19aefa0a
z1c35f1027ee5806bc311650baef61027cac9f2700d6a03326bb5901047570dd0f3a5fc01033ad7
z34e26748970a1a35cf1e40d49ffbf1cd586e188ea4180cba3ad593dd5ba66620465de9d86414ae
z082286f86a266d2dbcd92be25bbb3631cbb3770c522ef3dae75c6beba24ab6fdc9ece90a3e8dc1
z36b3b731191ae81650e7576d44d63a03e989bd8c9988d342b373b80a794dc803eb43b15f95cc48
za1794e85ec398b05dbed7c108247363ea021a794129c047348a0cd39f848e042783212f36b9eac
zb89e6fa9eaf37273160ed9be9f0c6ac0471e8ca39f4ab054aea54f97157f21fa70ae7cf893e185
z3063c60f78425f8616b41f9ad9b3dec8d68ad1856e3cf32ae86a9f5fbe2cf957cde3efb6c9d0ef
z4de8654bb599df3b120687d58d91522567e43043f9a10ccd8fb2aac1e51d337b092675c50ea852
z9f117ea80ae4fe9e55b9fefb90f59e8be83591667f62db2f133bc223497e220bd8233612cf69a4
z64e4c8bb94c89739bea3f10fcb640070407b9cd3f1abad35f87c16012ceffce985286dea92d826
z4ff99d4695147497083ccd92bdc075c7eff4341180f60fc66b96f5b5b40bfdc152e976daabc412
z01348765513237b65931148430c5594c80059b7ee28eaf4d36e51b6e177e0b1d07632607183dc7
zc4334c1fc61a29a07c96f7e2aeac3f09033219bbe985c480e418d87bcafcde3b3ffd14df807bc7
z3d1c29e0936daac1047c221908ecb8c991ab2539d826df45e885b62034980bcea1ee60e87aa17b
z9fd17e7c8b5f2456129b99564771c0af6b6b3878acc78fb82d0ba64cf0d2c031473f1c104f7e71
z5fafc279c4aa8c82fb6a71b8ee2c178d6f60f09f406bf34f6e25a383939e127f3d2a0c9804e32b
zd06883d3dc9f17f4bb0e55a079ccd403b2ccb51c9290a4585069368f7e4187de8389475af408ca
z4a68e096a90cdcc515eb0c4832f0bb20705fc94d0e593a0b3a45f85283b5160c3a219aac1e7dca
z9e8cad4ac7c64394134e0568bda56c52eed98ce83a3164db99fb157b90465360bfe4c1bd3bbeb2
zd7d8c9a6d569bb6cab666efea461b8693e349fda26375faab92b7bd2dbc4faa54af479e8dceb34
zaf660375b255f9a5d375d9d4f782588eac0459c1b181c94558e71df724d3ab1c774592283139e7
zb74454e48cf69b7932ce687fcc5a725d7493744adf03d1fa8336ac8befcf410b4e3c3c93dd3c9c
zfeb7aa93c6d80fa0c24562a68ddb767c797eb00f209caca5f644ba4c689a9e463875dee1d1b750
zdab617772cae0b4797d4c51776fcb4c65d5268022b18394abf52007754f124ef2d556a878fe923
z7fb3456c6a72cd6e83c14bf21178942b17d4d9c7c85d28cebee9af4a5cfc0238932f857e792990
z8e2ce62608e118d8d487ec63498682a4bb9de07c1cce3843f228a7cb472f0cbfa9b794f296ed97
zd5b5affd6861ced19ec5edce7a3c82b8462b95939640d52cfec540d9109f7d1e8c20647898988e
zb139abe435e25e79c858ae93ddc17a04568e92305a4a6c10ae0e77ae9522658f80454ee87267ef
z911e89e61af680d0cdde35a7cc0504010d7a3ac3891db049bf4e46ec1b6fb8bf0439e729099669
z9a07dafe1c703a23650e2e561593ddfd6f31c6922fcc04a19ae8cfe6be42e858409f77cfc41257
z4df0619fd0ef7e4af098eaf718e8476add8ec6f09570ba068f0ba8386fe8ab4cdb2869cf662bb4
z4636d25caf178c4eef83f2657ebcbe2f498a3d99b81cd0fdeecb5a399981d59d5976c444b7ef7d
z3074c2cb5e3b7e11c00be81efbbdd9a9de20863bb2eadcc1b78ff57e6ebefbb432cee0259a6064
z54529d70a1122a1d562eff7bab9de86772ef06bf15dba91f353783ca8f70939aa591776a38e5a8
z250d8b25f874701c387b52a44525d13b7f44a4befd9d3cc232587adefcef27bd251f7b47a754ba
z9d83281526d2fedeacaa510238d096b1018aaa03c00a61a4720d8286125950029b4e1ad880186d
zcc5a6f1214920b669237ef2baf37c9d5fdcc057b825fdbc97e8358ab9847ba5713537fe1dc4d74
zafbd0c82a450572a3e0c56f1375930b6c439a15c101a79a7ae0296e1176b77adaedb21817a0623
z5e1efae97814ae26d1dcc78d8de51a2b036a1e21bd1cf350d98d0125774f5a910396378db972fa
z0e9ffb5a7696b9a5242f7d7fcdee234ffe488b454779f3730c1e43e5633ce13a71d65fde7bad93
z5853d747079d4e1d2898f1a017f3effb3961ef88c6469d7957c25c23ff87eda9ffb257e50b4460
za1f3acb80855e55f872e7416589ba175447a3886735f84b0f5a6e08996f8f8c08e60c0c1278beb
za8004de3ad1d8350f4bf68efee9deb95ef3a69122f4fe429e8625027d371499ec74d1dcb66cc11
z9d78df7e12424cf3a52d357bd90e396b0b4b6d1897f34e73852658e4578af0c2aa50a5bfee0e37
zd756843897d2d98e774c48cc2b389da988795ff19382b095c0cc02fa02b03ef6ff8d0ceafa6457
z7bd0bb38d646d55737f9e1bdf92b9b07ee22856548dda96684c9af0ef3ba961ac2db918aeb322d
zcbaef60ddb02fa9c887d1b94366e126a6816750032a4b2b068d278ccde2c57c18d13b625d20b3c
z1bd0009af2520de395e310ea3444d5f653f30b0cf062d1ec1ff75dbe315bb4e0038b7e5492a60d
z02fb366fe371def4d74efc246aa7f47869d541cbf6d75ddaecb7667e153767de871465223119f3
z93578c9f27981facc170008238aea97135e60995f183cf76c88e02717a2dfe1fa1219b35f7cce6
z4b7fb05047f4d48e9747fba6b19af7f23ec38c7bf9c1acfcc89c3238de9954b56c1b5ea0afe6ef
z5789236b783e2ce8074f1d47653db727323b08f1ad9e7601947e5b345c200af5f1e84dd98a20ab
z08a2edb4a4f82e5060c9bc8c0c3a4fdc7c5c8817d66853719bd1aae83abaeee0c486836183fd17
z00d467deee9d0ad585b027b286626ed4b7501a2ba042ab536573e7e795073155ef65a4e8ac2681
z1a8c43ffa30c1de63312f430e1a3fa7a5658018bcc0ca77ebf108495e19b636f9adb08bf6135ad
z63ba5ac945dcd7bcf21efc2c14cbf20a8c8cb96d15d20455a1cf43a09bb15d4b334050797ececb
z4c3746cd9b604fa6458711ee706d4c698b49b4ab54195ff01dfc2fb3bf3bb78a25284440fe046c
z62e91544b5f5f6b11afe14d12e743cab7f8bb5b3e1110d11728e3662c85f148550e24a5f7f58c3
z7ca16a58121771a75fdc27d38ad7294d8debbff52b84c7c25721091fa59abee6d934303a1b1ed7
z5c64747b65401ebe9267ce83331b24f5925fdec56bf9353e948a56a59849583aa7f5714895c856
z437e4ecfa57ab15ee3c68c4dc587315d126933c9813d418041ed80ee302323230ff546d4d3dfa2
z9cb4c1d421537e114927d35ff611f794f799eeb40095efd44794ac57441d4fb706234f2c6cc169
z977df5ed487d3212a744d3939f01396de72f3340e8ae3d953ac068c6ef91dd5e303f4f58632f30
zca624c9f963f38d365bb6e21ec3abf459a1903ddf0cb31ead0b08708ab6719d3ced83c265d178d
z953b4566579f78857625f8fb500149a90da0d3517b6c67d85640cb6a4f5733373164c8bcac7028
ze483aaf2e1c24ecb68507b24998af593c0cd65ffc09f82124bfa4935780c9f50589a8b964113da
z03941f714f51f689a889681a85fbeb75d7346239b2153f90e34fd18251cdee7308c410dfca477e
z474c5eaf8023e0ae5d1f2f53be001756bcaf947f61be42f69de64254fd5d036e6bf2e6fceaaf0d
z3041d9151307fcfe1d1a2f149043780fc441c4184cd9af11d18776b3712a0a6aa75854c2fddd1e
z70172c769b08e392198a8393cfdc1b289d77cdc9ad12e1586706ed9776ee5600b4f67330497788
zdb897c192af1361c8e1c243f62cff8c49676f43a30f6ac5e4f63a4a17bd76d47a55bb7cda36939
zb6b756df51d510bef24bf0f22fc82f0d784706025d73148dfb57408827ff1c81e113ec16032e75
z2bb76dd368351c7dd642268c95fa5c3f3e22a21543f03ceafda060682e416f4694ccfa95e9900b
zbcb80d3c8145b1eababdb8a6186fe2240c50559ec2fc399f6eac949b67d64137cfd58aa2411a68
z03e1468ce0da9a0001778538122dae092af6c379af63a795bad547c74a378fc99380c02b6a4b0d
zd5dc5de91d3c5e1c034a96e948c2988abbc3cf49f32bf0266a579cc99ea3398b30f2cc2f8a8906
zb99a9ca75c767c94017afd4212facef9349a7fdd2732560c2de3fc6154763a28c0e085934b436b
z33d4a86a683a76c0b737238e90d247ee2b544e68ef33da8c1e374a3983a2fd19d824c0ccb73c40
z977c9d116bdd3f7a712125ec14150a2f803981d8e22e78450964fafd8dae178f40e76d92ea4251
z8a4100ea7d336ca77cf21ec78dd79bce516ff75f67d0dc56944dff7a02afb5c9ee62aff52f8ec0
z9c59182e7b80e820d9ba7b51f32d15560fcc54d02f98ab7377520139f678ad044c0269f07cb47c
z99748517a675de3162dd6a2880b9baafbdcbf6a32687d06011fae50a9c92df6d57851bd9e8613d
zfac6c6be7ba49c68f520e90e6f27aa79f9df7caffac3c780a309a3bae2881f62e02f9efb96a74d
z741c0ced1d6d8297f196219f37b0a5c7ca9a4e7f521b1a16d74fed1b64269a90775bb984fc7723
zb1327d95bdb289b98fc803b367f314459c82bfb1cd72b535ccec2c6cdf028a06302bdded92568a
zf4db09eb8dddd660e31aaeb000b2a4fcc903a017ead982011e988f5e48e9dea6ce4b9d8fc120c3
z8e7f2747f8c2634d409c40faed7924c3420b0fa5f262f5285efce650b2e488baa7c54e1655313e
z84d7a88d1d50cab4d2e18451a2ea12e144a2ddf704cd0e91c22011a9b94d312aa0175efb40c958
z3087172afaca67ba1fe16b5ec2bd530762f6edacd97b549fbdbb4d9551d84dbaf0f577654514aa
zc0502d0097059b4a5eee3cb9b430cd6a0bed01a4076b4736b30a02aa2ce276604eaef364818757
z30f21bf29555a82ef9cf63f16ca6ad43b61b5356d830d910333508a627efce110c00ee1a59d7b7
zc2d892216f05a874e7f10d6be7a02684eb8570795a9454c34ac2fd6d058886bd5c351916ba7ce1
z872d4d2839f79aca08cf51601def95e83f90e12f3ba5dbdd190123f33c1258fb797fcfd1a03739
z6a409aba8888348eb9cfb019ea0b94f156dbbf84ef9ec199a50afabd79414a04dd13f651cb505a
z0b57ba72c6068dbf9d158aed3564a51375ada69ff1a24daf6b71816e0695013564023260729afd
zfa62cdfb4629614a6af9c6059e27c12e0fa34f3c4a5a098aeed91001e918c902b22d5bea0a3f01
zb33ba68334c6c565f576379656ded1711b9f19be1bdeb225613a6d1bcdcd05481e21460c132212
zdadacace101e648a462da12b5bf21f6a582576e8bec4e4f96192634cdeef85d10e106abbba7aec
zf20f2453dd5235e1cec1ae98dcd5ef4c82b2a90f61a2d6f2cf41fc093042632704cc18723f7039
zdd927fe56bf4009e8116cd896103b8c53e150ffd9b0b7164eb711523b79d4a8f57a0bd627e9523
z40c4dc00c80cb25f43d3ce557a2166b5f2d1af68d736af15d5d83de439edac153c42214a4e3b3a
za4a5b02273ca0f882c72d717b011b97e31dad09fb4f161f4b9b29f5e6d4dda7265d1d8a0f7397a
z75583d932e57b2e69647464721faae41423aeda319acd68c73c9b4cb8cadfa8759d39fe5c52020
z087de0eb5a4c08910f9608cf04aa70ad2de8cc67498931fa1efa28563cc15f09bec9c66a3ba0f0
z7faff1fb92315e1252b60e37708d6a4f63215ff998a46b328970201568eeebf7fb49ca343544bd
zab6e0b8ebda8349b845fb7162dcfb3ded5a70f4539265ce97aa56394f7afde0f5c21720152f002
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_change_timer_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
