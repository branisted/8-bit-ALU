`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026201628cee5aae21fb892db766c4
zb5b1406e11aebfd6dfacc9da5ec03b70c276807a3eb15e28ec7ab1dddec42388b9424ea285623a
z248195c9f894b36317ca6e59c86f11031163f5f5bfdba36b10b435d36514783bc1c6e60eaff7f9
za2b8eba90f8fd9a9cd7c932ce34efca1757e6b2718aa68644ba032b1bdd74efc688b935cf38d81
zb1f311df3e5b8e4d46dbf459c824f309500192485674c175e61de609f1c94488da73614dd500c3
z680b7fbf510ef6c68927870992ed3376661d943d2a929d90faac51228c485cc4f90c0eee6be4a2
zce41f6565994f8c457ad3f059f0f75d13b595288a756e41a6033f636eea17dcdf0844c8e225d45
z55436586fc78f7c2c04155001676fa3f49b24d3beb3584c63daa43ed80ce015162ba22d33c9763
zba142d3955797e70f433f00a9ae14f9d776b76291d31153dd23eef201b698c8aa3a640b228a83f
z18eedf1d37da4b3680484605b10d0117d140a2fec482eb066a6b3e23701cd7a6c894de53e39ac7
z965f6450c8b1c2aeef13e4dbbd2cfb983fae62219cce167861d4291eb96a217f8c834ac6d8cd97
z3fb107301461c673b573fe10ba27feffb84003be8504678bdeb8fde88ef5ce321f88cb3311d3e4
z3967093b4d555c4434ca75af2749c48959e85d0c3a9fbfbebcebb6494d83e27e01ac4c667ed322
za3b077f2f69273f140dcda394caf8c2a8ce384c08761d34cb8c43346b815742115c69db52129ff
z5844ab9bb4552a6ecfec0617ae18cde60d8143585820e4d584bc0146010ee65c6367bd4ebb9116
zdef9f83ca5f2510db14e3c4c3159d928e5362e7283c09d5d7d951a4de11d8f04b9ed9b2a912a25
z32a274bfce4f54e4cfed937ef40e4a69e595ab44bf66b1acb8a0fa0b91302457e1f4d000e946ac
zda0de85e09fbab1b7f7dccdd45b53c2533a3082f08cc0bafad1d4db319048fcf4c05dc77412102
zda864d6fadb88ed0b50175b782181bfaf3c6501b089c03267dbff78d772e9ad5ec71919ffa3a8b
z0297eea20a6dc97d43737912ddb87addd89af196d58df0ea2eb6596b2d61512b550bdc2d0e25e4
zbd1ed43e87cc5488c07143e89262f655b5ba02a907500c83a8562355b77333d42f2cdaf419cc0f
z052fcdcf2d96ec830cce129dc934b3a9b255ad6245271f167622b385745cb23209dfab390ed023
z6548878399244a4dde01d35bc70f128b2e6766f4a97e2be95d7027c3f59e6df0b6b8e470db447e
z604ed1987145739b28a323859e0ec35945a04ece5dd0836832d2c7173114d1ce61ae7a1b2d4d4e
z135402d9779c00aeace2c84599d517892fd7501d4a53afa9d9f36b658cc40c7d157a0ea4659f77
z93d7870ed99ad90b393d28bca30d85b3e5a2e4638e5b734435c93ae24e41273794207a9bd83d3d
zbb627bc67cfc8c92afe8088c645dc3c729ccac0b64150b5a2ea8ec45be020ea1f60fd92f0c12df
z92a84c7b5889bce16bbdea4f080314a5fae63273d84efc861e3db1e7833b74c9006d3b5fc72c86
z946076df62f85265a2b0b6e89de592293f6539c64bd27b1883742693773dfb4e6ba73ce3f80ede
z00b7696fbe9445902438eec0ec8128bf47230d4b4409d1966fc94454df46a90e7b60681196897e
z61fe55bccaf7672bf403b6911f99e982d14b941421549c47de632e95e5904ebcd1917d2c5a1a78
z4278c6ae7a7a171a0292d393e7abfa1f75b0a63dfaed6c429aadb52e099cceec4bbccf79194aec
zd23cbbd782c50d701ae18fab0767c9ee872fdebbb14ee9282d43215fd1af80b2f3c60f723c6dfc
z971197b408ac21d98cc44c567c6a3724d0a3db9a0f58e1da1d6c87290b19fc4019a2858fd3fa81
zcffcedb323b855fd9937a6dd586cf28f63ddec94e70c1aeb08dd33a6e323976edfa4644211c89e
ze424979b14ab038e2e5295ebc27f7c9eb12f9cf849a35012da657ea66eb23c81c7404db1bb0b88
z98ee0810c88099e0554d7d077fc78cce2411522cc90cfd232a9c67a464f8ada168965909819f9c
za19a72b66c01121640e391717e351c149138ac2dc805bc523eeb65673a051734b218aeeed51ec4
z8f94ad1354636335f16875e7e6a9040a23c9ab8b0a1bbe0234fc936678454984d1efd5e7550731
z7c569b721a77f2a0cc870331fa3a52876335a204c19d6f24044e2698c6303142b1ddb817e9e2a4
z100ba0e26591bc870e95807d27cb736c1c34f421038323a21f2654506feb7fb23d41ca60e1c317
z468c2fc6d0f2df6b5b9df43a89e6802a70da55da9f31bcde5ca28a20f0ca51a1e4999fc966129d
z60d7897e24a541bb37034f8156c40f8cce82a26cbaffc93163ca2db266406f94aa865733e16030
ze149459f92be7690a2e5aafe1b439f6e494889f46838f04b851ea01b4243a9256fdf3ef803399d
z3437adb1b95ae7a698710d15cbbdb6e8a44ed88cd4d7e8e25184193b5cf2a867b68efd17449409
z15487b4c6751e3d452870d5cbea8395fa892d18677059d8de4fad71a8fb09f5c8b2aa0f8c3d7ab
zbfbb5b2090d69110e86b7180a69b3846c879558fe05b139f7392f52a19fd127ff5d499855e4d38
z12fb6374b7b71d78823c56b97e2906e1810b96146a98940e8f60fd75498ffb787dcd45afbb74b3
z3412479ff6f17151d89d1c172f2bce989e15a61315d851edbb53d9a1b8e31c622aba1006d7837c
z9b80756dff81c7794cb14032e8e44fa1c5a9d042742ec7ffedd0418d6b8eea85ed436ed332ff29
ze67c1be075b48c937ec151835b08ceab0b58ffc03fc30e92eb75f78f14228bf071d6dd41ff196b
zbe7d6185517fb1d6a9e93ee0ad15dab1fb31e9148c8531a04f1cc6e1ba7724a3a51c76b13cc9d4
z91993901599cb08b7ebacefff3c8d0589222eb70559ac3d3d15e6f8446bf4deb87e5dc7d09470a
z0f2a403361baf45807c4fdea251d1786a916c63e7707154e5afa726d12150611e3b55ee4b57305
zbaa4f89ab8f976f77c703256dca711d8e03fee6dd1d7c001bd8bee1ca456e0168a3f7f33c44cca
zea56babc9d3046cfff80f4b11677d9f4346593425b2b0e3c08ef60f83fd2574d53b4358cfbeb01
z04b191f73aa1c97cd73d8bdc22e867b09c3796673ffacc9c6a948e6c68fa8f0c9d3a736e22a691
zdb9fa8002f3151f536000991748f331cefe7c2be2176b0a970917c825c0295c731ae309dbb1e26
z4289b117c5857fa18bc213f0738f721fe9b03a7c52a9fa01392e348e13e7957fb78c5aeef630bb
zaa14ec6a9c1c3e30fdcc90bcf760b037625ced920aea5334fb905051034b5f46526ebf9005c1a2
z2cab37ac9a550592c2a8c35470b192a28160b2cc42d6d2def60beb558e5d01d5149d52ac53d663
z185ec4ccdc13ba2ab27cc10453f0d3df47a45dbb57a1815002311c9f5af0344b8dcf42af61b48b
zb0e75929269e8ddb06e23aa9634dd485e0ee02cbc8a5e91f4a250ebe68e20acf826748c2a25f3d
z6cafb85569c89263b7add34217bed12658bfc4c35cb9155b1bc39ddc59be6191d846b7bede9d31
z59117adee5e9a0dfb894cae3861f862d9d65e40b0e56e4b903e07e7ee30888ece8d9ddfbafce2e
z3fb5315e06fae7ffa90d9be58db52ee2232ba4ab70466cb87b5fe7e31e7cb2657a08f584a46a20
z870fb3007fa7bf96057e1ca128acbcbdaf5007b0aa3bbd7e32063190f7f309da55861d792843c1
z2f17b60ba44c9dfdfcc4bd99dcd2cdff966caf7721e891991b30c410282eb51f0b5befa44ae0fe
z44dfa8791fd8416e82aa691d8ad76a510e9a7831c3223d871c1ec3fd0537f529f3eca73b7dd1f1
zd41507f3d9fa9f5f891df1021997b56d4439d965f7539aded61cae241741ae6bf73d3724e845c5
z6810a81ddad475e87246bee39a9e0e4fd7f8e8c1be5e72fa282faec0f1ee21c397307170ee7b36
z276b9691ad80a5d77f12ddfb4e0bc54c2bd8258e8c7f29beca106329e79164e8064a0b068f5ad6
z3aea4423a91acee3041a11436c7710eafa450ca99d155f28413eb774be4d647d95265260fc3476
z8bfda78cbb3631f719e7ae4cb143103691fc1857fe1b9ab7b94bd72ee01684cf57df2a157793ae
z5782afef76eeafbd6a27e2771c67367d64bc7d0b655349aa8a68d98f0bcbce5d31bb008eb776d3
zba532dc6fb1192936985c042053e59bc056a38c9910480a97f201a6834a55011cf2d22942c6089
z94d189e81a95585e1c41b9c1595f6d0dfacddb08399850ae86e91120bf53390bcdc987a417f938
z1f9b34365d73123a76e0b7583465d55e3287e1fe679e34c6687c6f57441d745afecd584536cf74
z1fd7a725920c24d3f618732bf6afaaeb2169b6b93776ffcfadd53675d4ce0fe897311d5f1bf621
z31322c4111a97a02e6bd1f7046c702ff0db612f26f94d0e57cde0cb2eb14c6a42bfc07d9360cf2
zffe0c3037d807a3d4303b7c4c6aa72b7420ead6a5529ddfb44cb57413b5c4e45028042dbb29f6b
z605436daab53ac561a3cbf399401b1046b79180c72961196dd706e52b4660c23226e1f381cd9b0
z6c5ac1889ee3f05c9054d301ffb62348904f4657e2c43f16da9770f781c58cdb2f9ab81faf9694
z1747f6829a2d3160a99e8a3cef4eb30ee14c36a188f2eee6676761bf276dac2bc6108119845adc
z77497ac0c5cb55f50cb103ebcae3f50810906441ef1162bf1160b72d5bff887570865f35ab6fdf
z7282a8be44d962e81559034227672b9530fa197ccbac8cda2586ffa850f3014d2489050e9dd726
z080dc2ed64cd016794d7835d5d187e3c0a4db40a3bd66f1c78b35db8e738c808367a4b16218849
z3b38cb89c5d454870008c97143eb2ffbd751a16b4e4d0fdcf12930813a0b9378408f7209307f2f
zceaa83b6f4f9cca21bc535f4819b91e5b129c29ca57aef6287002563bd8c98b5e6e144a249e87d
z79f1b3bbd56bd46c31c4148b021ffef16438c53cb5475abbd58564b661a9a2d5c22be12a3fce8b
zfee1a47085cbd754715654de2380549bf85e361a319f1a687f73e0eae22899c93feea3c522e42f
zcfc6f447ade89b28ed25367bdb2062850e1319e3deba92f1772dcd2b7522b7a65d97201ca9631f
z5b544bbcd94e365597164cc90dd09ec00c1da4332cd53ba361614c28c6a72090169b3074727047
z1b0593c0375dbcfff56123708519330690de192fefa2af3d9edb38634fc581622807312277df95
z33b40b67e617a9dbc793eeb79124bd266ad89a31d20da62a2a3fcef9208cd5e1ec832bd4b684e4
z59e5d67be7842eacb774c26c986c2c94356e6e2d428261073392e67b6a3d09ef27dbcf8c70ac50
z7fdc630a10fab3b7fc3b51a1bf1dc0193ee7adf47d2cbd1abad30fe04a97db45f4aa34693cb98d
za187341dba65829ee4ccbe8281ba84bd3195d294cdf5a9a731c9f46f8d7fd749000ee02181e03d
z617ce0dd64629e1e70e91536467aca515c53c64c44866cda5e744bd82fab9ca30624916a81dfa8
z2a063d2f70551adbaf91f290f53f9313b774674a969d4d0083e587ae38fa4d559c04115c8fe11f
z39f5cd28532b6622af915327eff41877b215cade64c45e5efdb5f29c11a9309d406f7ab0e3ffee
z4528e5c7e85a14df26eaacdc49732a4c346632d6d5c993bf9c6c81f8479555a3fba42bd37bf5e0
zcac5e8dbc639d22181c04a8de7f52d63e4c98bacd127abadc870bd0fe2cb9b2a3207d85f5504e2
zf2e0dbb2d41db8086623fe083306136d9d7ae742154c5cda8a1fca200172c6d0ec073fd7bab246
z8eb9cb830e02aa6eb92b51a94bc5bec59a8e8c34597075a70fde50c3702371649bf5096431b00b
zb3864e9483feb8e30cd337561a67cbfe2cbc9ab39145200b46177e6dd54eb6a6d6971d32c98657
z5c15d678e61dd4d0693190d819542dad31348eda314b2f78a39377684c01804d52f5f1d56ad07e
z7f352d19854d39248ba91a0535a64eedbe9ec4d68a59aa5212a789c1fb3271582b1b6b785461db
zee7d92523a211919cd9dbb59fb5ecd1349dad5606c293f92590821352d8d7f6db40c44763894ec
z3a6b1dffe99aa40e70b7ee2aaf4cd4abb2917697061401b5b9abc27984b8b7814b60e2491f93cf
z61a594ea9ac92cdefd9952df47bae043f88af4f96219147ee446034022fc216a7766bbc4ac77e8
z226f31eeb2df9010728c3a40cfe3bf9a8803d01deb32b3579f835eb42efe3612be6bc6ba34b184
zab856962e2efeec1bd90087f87475f61dd547271c8c033dfd28ce2ab542538d58ee1f13296188b
zd3c63017cb9e49f45e2660f7d136b9d9d4bf5372aef0665ee58eb8ff76d44ceea6eafe4196efc0
z5ebdc96425cb7d2777b2b4837bb7396c92190c4d7ed43464185f523c719fb8d506743cae3ab4cb
zaca0e7dee02f9811cd50d9a87766bfe209ada31e514c9b85b57e2d2c497e27d7b59ae74a3b4acc
z35ca60ce48bbb1f02d14ce22b59427c287924ffeeead4a0bca24d359a7b41a1a7d2a6a9988a690
zed68c6cc65ea87d77154d4b4dc2e0e1286537c4c261ba889f9621b9385838c94ac1ed994d0e94d
z8b6f37b58966d8ef8f6796449ea21ebc60e12df54ace39d9896405a067d474538d868f08a1be86
z1c4b9905eff81a924fe536e8f4e03350416f58405c2f0d0b7e1d00085504b72d620a8dfc8cb3e0
z5d91c661b5298847e8d33fa8c670d744f0203e1f959b53a5addb2eb0601080227ebaef895cd40c
z0c1395b1fe1d2f9865538aaa23afe730e430f52a9def52d362b731e606fabfcde4cb4465431f1b
zb66fb27ba36bc9309be65c5284d6540bb4e2b3b66c2d9c1afa5c480de1f5087af4d760e1fe2c95
zb91226da7d29e8eba82e28ac49d55e2a4c1856cb97c769527603718d1f2f774375df44732b5b1d
z2429d17bf8655655db8258d4850f5aa8e357b39ed48a5865a1883f2a1fb656c90dbbe6d9f760af
za0b3c3f46a5953ed648ac2a3a966af5550c9d72dac49b2c794bb787b391161dd3188f4b37ef03a
z28eca927f4afaf63b3c9095a5fda89515739514e95baeb9e64605f271726efe1e6acd94959a1b9
z04007625e2a72e078335aad0026b14cebb9b39983b08100e8557291aaa99c89c13705865c21260
z042697831d185c8f9011a93fac4fbcabe42e796fb474b5695048ffc58be283395492a4785ae6fb
z71ca517ee0c0b86a3caced1dd08961bb7651dff83a97566c7fb57431b84a0e4dae79a99579950b
z28e94367c8e6bb7e72eb0847e82839b7380c3f35e93553fa6c24ce18dcdaffa0bfa29be26d7052
z8032cd82faa8aa70a7cec990eafb742ab4fe6033444cb46f9cbdd5e0925ffa0f4a6cf8629c2f8f
z64ae01917ed84cb94bb40e6a50b9356517ed9b3f516e7c7955e10524efc999f539bc6c3eaad093
zb0ec8171091374a0cef044563988891a42ebcd85d7b9acdfb95e585894109f25ffba44a30a25ce
z11d17448f577ee4c8f637f6b48151c043cabfdeb8b8933ccbaebe420affc637652181fa38ca165
z362096358cb288799a8ea9296da13bd7a5993477318e75b3da3fb4afc33b7702f93323b69e1666
za1b7fb89cd2f1e364396eb8fd59a8b70823b9cd1cb799ad69a4bdf2ec8e98db49c181b480c3621
z15546f7a2ca384c88d7b19ebe7de02076c8f5223eff8fe0071f4ad083216ca8c6b2a9a7db3f8a2
z020b464c35ff727dde6c1757f6675109caa8684700bd0d24061b59f85c8d0727dba77e076b4e2a
zdee96645e687f5a9af35c1599f300423298e9b3a8896449b93fb0c0ea035cbc4d994805fdeb7f4
z4abafded7cb0097438ce701684265bc043ce2150a7dffc879539286fed124c3f3b933bad232c64
z97d8443d6fa1dff8bdae20f5450c3b04a26aaa8da6bc4cef2395763e7a9b2971535d47e4656c99
z04c8caecee7d865da8ebed46d42ff49112576ff4795e8c6ab908a01381199073922c765d0e3d8f
z838fd3fa9b11b6c779733ff50849264543779dfca7cad558ffa5f5a3f6656e45f1a0293661b23c
z8bdd702551ffa9fd1ae16d336afa8f3c5efa5ab9b4c222e48b4af483fa16c8be9ac41e960ea415
z3b86004a0dc79ad3cd6404874890fd0c6796d3edbd2e96b02004637a81bab711f42a85ff24de20
zf5b7182b9a75103fc411dcd760527f61698e17f1dce67bcb6790e43d3a6b8e4680a1aa763dde5a
z36f0a3ed52ac9ff248281b047a7f60120b8bae134077ffc2b9a3544ca8c7efa0342afd7bdec6d7
z0a752f117c908f9a8ff3a548451665887f114dfcdfdafb900d1d0bce6a30cc6020d0e9ffea67eb
z6d78e0f20240973e3dd6e33f993cabbdb780972c9aff246f5fc4d676024252a0b2b8eb1f967ed2
z30d2cc94347702703719205fc43f801f704c344b853067f4e3fde97ab642ed4c38bc735a61f55e
z08f76d59b8dc6533b11f27976b02fe3067ac929367a6b68b3dc3feba52f1b6c21e570ca06916ae
z3aaf2ef3d93a0cb8eab3a4bb76ce8f69c3978265955faa69aec29ce85b999a7bf3d94ccd10e37f
zcebb4eecd02673f3f0bd88d4070ad67d6508244bf1ca61ba1249917e0d710646895dfcc3a5c725
zd4ffd4bdd008578c5d455158616242a3a45a8c6a5b34e64b220ccbd1051c4debe36efee4dd253d
z030b5606a1c60773560da7289ba70cd7927ea39faef4a662b8a38fccb536fb461bfd53656ab1f4
za5981b884e105d7eca7e7154cc4ed5bac40ed4b26a86719e2eed91fe200209d493a0af6f221e98
zcd1cee7b84026cfab3a5855c004941167b020dc7de8a1386b03e967528bb70859d677eec2862db
z2cd76ae6c635e8dd8e60f4deafbc7c3ef858e1a0fd384daf79503f0335149167616f27d364583c
z6eff6e099193d343027e0350b984815f1ca23ed1faf736002e5c381f7bab2d96be282c0597de8d
zd39a4da8b33450eee51a168b43424637f87e8b91e860a7c8806d015e8bb1b4d90f3be6da767455
z757a8f62290536875d1e467fa37a3777c359042a679cbba53ae078be0094bd4561bbd213440b24
zbe7a37c5a49089b33b8389807e8110c30bc83f33cb88179416b61344d41e3864efd707ea434888
z7e4deab2051f98c682011dd6ece59d7248d63f010493bf700c677360b5db2734f232203e708de0
z550584502b48efa408a24a865e8b6f12d6600df984ebb0d246dd434e6df5e896eb61859a4fba93
z07ac7d8e6445054fb8e8be154f7b57d808e2743fa38f641b0366a997fa989e56a33bdf7ad91054
zb710c86e3b932711f39dcc264c1606636ba95e2fde8e407c4d9bd6700c499ba487d45d742dbec6
z25f534541c723382edce86cdc3ac287f7fe260a070f0c6daa6e8a834bdd502ef532de7dc13dc1c
zb23ae886c0d700122a7d038cff9cff7d6c88f7e635066f4d1470aad46fe28209520941182592ae
z49386aa10e2dd22b492ed2cf96714a7393f9c600be1335a5e17f7a7131f62ea93adfefd98f9996
zb4682ae88fe4f5858fba05679eba61be16350fed9d0b4216d90a8b766a240b953960c9aabf468e
z0a7e24f955310fa530f887cab6ff18f29e7edc27fe74527df77e0d4abfaea16f5d31a7fa36879d
zb23ed6bd59100c018f2e76aa2416f4f850a6af799247fcdf1f013be6c0523d8f7aee0d65098f10
z35be2adf5d7fefd53ac501071fc5a0b311fddbb9dc1daf820e4cbfc977eff8b684f14ef6291cfc
z3fe47a687f88c7eb921205fc370234e0c4844bf43bd92a9d43cdd2ff6fdaa28dfd188feb0fa48e
z382d468196a95b1a696e99ed36fd7c6e1326c3d963560dac49e59ce09f04c76db660a9a67d3ef9
zbbb8a848391eece45a9cc72cc7bbe78eabe1bda25547d63581e68b09c4fded149c02d22b26803a
zbe795b94853324112a3871360f1c18562cdac5c1ffaf4fab63f310baeec82265e8a0ac98b428c8
z3e96bceae1e3ae1e9c40aedc9d388f28705444d0078ad9dc462fed8845a63752a48c29bb81d1ae
za5e3e614b5c7a1ed21b637898cd5c08c2ee9d0c2202d7d27a585e9756aad2326bacd456b20bb42
z33bd43dd842a9ba72dd8ab33bbb6a559890c89c42c69ba7ad1f84eb73a9124a209d7f9c86b8fd2
z22567681307b5602fc5805815304a438dfbb0bdd7720f6d761905c4a356bcee8af76624994ffc1
zaf97188c05864491e76c423e0f0e0f2a485610843a748c0f29b06eb823872ba98baf686aef06ff
z82605a465ad63984654261ba3b283ec0b925d54b0374f03a615ac70d5e04f2f6e787518578a2f8
z6644f05c461a2bbdffa48863846c63c878971a82409930a54a7d121ec6a21dfd00fdfdfc24f601
ze3c235c927edef1e1f03db96e53cfaf5c18454b0dad8d0ad9c8221afd3fbc697b315a89a9526f2
z58366f970fd974a5853a0aca5c0180eefb7e55824e4bc6d9f284d24ac0eedab6d486d5eb40964d
zc20bb8e419c59df97e1c39aceb106adf8aff9c20436885f85f6c04fbe0c5cd7f8fc4b8c9e6104a
z77dfaa7a8a3e9d530279ed1c5ce2ba546cbe006e8ef4c4e3a19cfd5af4c8d3ef98c27c6ce761c7
z956978066e0d1d9460fde1904c675a73caa52b341b264b8da1ff863b59fcdbfd5028dfcc625d3b
zfc493af0257953d5d4614fa7d82c3babb8cefce9866f4a9f5461631d1ccdea915f947d8ac22b87
z3ff64b1ac28dd851fc09af0ab13dfa4f8a0a75d7e16c7dfa45bb5da275a643456f8975912ee2a0
z34210db06886a74aa369a611b99e360928fa30d3c7c433873ac5427601e176154e60ec330eb92c
za4ae21a32dc6ce2f0adb9f2104a99fd86b2e8ebff1bab0bfa525fc9298470f36afbdece0f51442
z749164413a84291ff18ac3593c08589df7586aab07900e01aac028682861e382b440a8b2e56329
z10a0bba375efad704aeb0abab05a54c7d15f589e0fe8bc6f12a3a01411e28fc57b948f63a2f097
z63c65b5ece4e53c170bfaf272fe0ee57c445da9fd96e286227e7a29e7d93f49f3de453349fcf71
z8ff2a36d4fab8b5513182f1917e705fd1222977a251f1828124d9b57aa67fc3e16fa6da4e04779
zabe7af60c299cd07ff9a4cbe10cd222199427cf3a7f46487571ea482ff10846753d5562ee4efa1
z9aac7eb1c2a39cd461e7e963fecdffb01c38d9f75cc67de6217169c918f0edd5d6294af6c2938e
z61bde4720f6859bab55d01e28d02bdf42bc5ba94b773c610f35ed596276b49b1d7b611fe1b05ee
z8037b65e392a56224a0d93f678b121190f9b4f0a83255b3ad1dd033fbaf55f26ee66290432f9a4
z11ebcb068091d55abc245f05bf80a8ccbe277605f1c7d3e2d378ebe16a82af4fea68da5215e386
zd1a5817bd104b88fb5600f7ebf602b6331126cb4308c797a4cfbd1ccf5c779e0ec965024b6eca8
za5b67f5ebc1d311f792e119aea8a7e0378e2a80ca62df358a64255a502449f8f92493a07e86a03
z4f09d597f4a04f57aee1e96bcfdae8a1f0d4130361ff27422b3d03ccf94b47c63fb3c854242496
zf8899ebb5b41e58fd0525a5ed450cf6e8ff0544660b5d91a710d295cd34ceba8b8a152cb7492a1
z8db4a2f7db4cd5fed19afcc771371256bb43e8e999cfed2d55441b21e4eaa96527c96797cee0e5
z6650baa96b59cce22ac6d2a84ebc5ea1e65f833f68fb98e555dbe7cafd04180e164f16feeb3fa0
zdc4cbf12ef26bc5a1d90ec42b3f22de91f62d88e9beec34f7e4803efebbaddce1198a5c7ff62f4
z27982dccb72709b663925c203ad6658eb61251608424cdf739f2fd30ef5d780618ab54cbe63304
z12788e803a804e453b1c933dae2bc5292e38d1578ca1e0753723639728647a4cfb48f580aea5b7
za673451ed2aa006fe2121e9a8f113c497b953b37897b7f1c6d0811e359ee3df2e3f0dc54fc06a9
zf05579c80a24f422ed8c3b5f5cd6381b4dbb73ef3a2fbe16f76bc2ebe3c37689db328f18b65e09
zaa9935b7f829a895801a465834bc1735b1cdaa928d279fc2451a87bb195ac4f9f98a6958f9fc9f
z3823c068be9cc8073b33cae88d5c8e7ecf0e68b9658d70c35c4e6173ad794e59f76dccd7936e59
z3288ade48afc4ef9793f2803ed1c881cb71d64d1cd2ffc54a7d4f352daae75cffd3c2bc655c8a4
zb14b727c0484ba202f1a63d87881dc0987b7d8d16b020a1003725216c4fc5ccb238f5c83b61363
z2e7a6cd3763f6dc2c915d7d537934167b1066bc0a76225a366093adbbcd81414067615db7ef6c9
zf517381fab003c4c95688a9a0a4de775f899c3d9ef97e227965f9fbdd20ae0702d6cc0f97f0215
zcba66703962046b69aad0334b0b714e06d2de4d3ef685348eeb86b0b7cdf1ad6933b9ba969083e
z3547ebcc14ce2929bcf6f073779f6a0c2f752dd9a159b458fd1224b1b76c987505559a8ac72133
z3a7d6afd2014fdb7541d3de46d2df061ebe4ef88d95e57775dfd84627af69bb760d238cb9ae40c
z51b0b7f6fe33b2cf23efc3c0b8b4bfc5169c5639c80c40d34820478ef65378564424209947e707
z0ca7455142f263a3f28a844d766786efd6a24a18ca4795cd3c4749e204ca7e8086ae1b21143d5b
zfe3cf7618e5fe7885db8d7b67cdc89668626110f7635f293abefd8c64b2a9d7a1b6ef4a848585d
z07caf6256835f5fa414fc0407fdd2c2538aeadd40e740cff68ad4f34232237ce0d1df67bf5ee2b
z418f092f5b40724ff27229ef74ef14b83936e2fe86d6267e0390f32dc8fe29167fd899cf48410e
zfd2c4fed5baf956a864cf28706a559b43b4222e99b4dd7c5248034274ba884677a174c656f2930
z07551d00c3f63903e365eed36a0474a198cf03be2ad69e16c62ecf98597096fc6ab715a192682e
z5b1e1b93a28b9c78d05d6bd59611ca2687019111a1e00a16766b4a11d0688e9676b3a332b21dbc
za13f89d323e02ad167444fb97dc29f3670c53fa02874d0c812667f3e4e7781566d7a7354a90c78
z6a3461f0346f6931f94507c86b41a32838d5f8e48fd358ff33bda39b7d7641c657c3ae9b3b8aaa
z8228729648d4162f8cf99cfab77641a26309ed88c5009bed365f8fe89a5176a8144cc5437eeb86
z9540f7921061962e28be204e43f9253ea045911e3f9ffa6c41e0ae30140840c225d44bea130696
zd387cdefe3c2af5173a2d6f5bafe3a4598bc18b410ac3b42d203addebe0b229266f2ac30e5685f
zbaf72f7460811066f8a84a755fc3f618262e7aa7e5c9032efaa9af92a7b6e4d209a0ed02095859
z3aaba302faadd77213040e7e287bf44bcc4797c495ce47214d3f28551a5b64390bf81dc0892ddf
ze9ac2cb1def3e378abff22d3a7be4f85c4633b4f27946e886494e8be7521a25e105b60cb3002c3
z043b56cbf11f49cb4728883bb61a905f7abef75c084c443a0de2c27ee30c54aeef878d11218f6f
z2ffb8da6c7ce45eec0f34a3be3f6a6cc06cb020969643ba2247fbe3517486f5deec481aee0f455
za7b7a94bd9faa75112e541dccc653cfaab6c7881e4fc42487695f1b19cc08a039001789ab30ee4
z03276313d39b8a018f20b5bea14553c210b8ccd68906a8e674dd90df94bb8cc3f2d4e1755c62e0
z9811b809edb2a05cba6171ccd8d00e644d0e4a4b53df041ef8f854f06ea6c0a84ae26345096915
z5ff0ddc8e74301abe69d5cde0b4deb4699751e3e2e46e4c6fbf920e22be7dc63a053ae701449fe
z4d768cd3a292ce840f797af5ca40d788b45a1818e4e1940638c4cd2a92248f9a764f30ccca6e89
zd8de204d581f3df268799e2db21f321b157a157643aaa63e61a3c810612ac6d13aec1a17c71f8d
zdf549d0589d242684a1fa29dacfb0b5bed012f54dcd4a20401a45869b466c9e3b942c778f47c08
zd5dfe3a4e6c4a4f5a87c703a7a96768c65d234912e7e53709cb732b91d90a576a3dae97edd387c
z1c02c0977a7040ed6f6cb922faad7bbd3df0c929344b5c207a93bd4f2e4f418be1ae93dee414d2
zfca67a5b2410652f7e5df1325469487be7aa5211342f7100044ab090842b397ca83fcdecd0a19c
za6cb94ac23e20ac2846e78431b977d9162415fa27f3a68f74b66ff303baa2244234b27b3e841ef
zd8a9375e0a97e21d33c5720add4d24a77fb404eb52b159baf3dc3f80bd163dae91ba4a162115d7
z4c4eb8f73bc537310fa6365c262a233a4bd9ccfab2319217cf71179d8b915577c4ae27de51a569
z504054fab0f1cf94ad90eefbec734a8de62ad887e6af8a83c8f51c44bcf68642adff7ba1eb9b2b
z27357539273fc5b4c1d6072a6230ea855b28ec4801e0620cfeb932d21e5146c28335ba70c0d7d4
zd0732f7b3b03b950bfdcae8bc05b8e29fad2e26524bf233848b838c9ca6e1a3c6107bf581d0c74
z85d20ba44bd63138e8f55b77fab9635fd0eb1ee9259439e774b3bee53d5e6da5bb4ba5b08e9ef7
zb94c6ea5b10aedd6e6a7019c2c045c71cf624269519dee87e09dcadfe7083065d1ca07c046d49c
z1ee691a018a4b09c1fc13423f982058d18da64a6f227d83ecbc0d2b5c0c153bdf581467014fab8
zdca62e22350458ff39d4f027de8ced1c83877d87169227d0725cbc8c4f8e228377daaf8c80d96c
z32ba96742c4e6a4f2490941b165f3c86fb638c652893969014bd8a63a3871490e4c9faf1bc0f15
z07319c65099c3f4e07f11291dcfd85b0e8f5dc6f42c5ba940bee40e6448c9dfa5f7e9595086bcd
zfbafe618524b974ac14559e0d4fe93fa46a686a8ba67cdd366d953de73d42a9d1fa3337986979f
z8ab8c6dd795ec01f3adcc4d798026cf1f61fc58479e40b9d71e551b42c7312f51671a98c606ee7
z126bdd5645c6f7a917124dc6e0356a9b5764b5832f6dcfa7c567c9ce5c3fe68650cef0bbb2dc21
ze1b1f95241f4df45d3df3cccfe6ba7372032f6f1c6e8b807e3432038228217aeae322ca1ec49bd
zb0cf8340e6e4b6687047c4d4cb8cc2cbc50e24b27e9ec49d19242a40bae1c6f77b923bf10e97cb
zce7fe703970effbeab9ad69b6a2e75deffa04268e607791c6762bf3bd1434ceb76bb2e7ce0f202
z719806598b7d7a8993f7ac6a7a6227506fc276b9903cabe4835875c7451f36f8182067bbc47233
zdc25b8e5a5997993d358c70ead51f1553092814e9a970c05be505a32e2cfefba582ebda6c98518
z89e73b25727c40640cfca84f9e154833598765f4c5104e4de57bc342e174d5c53dab4d017d5738
z157eb4837aa81b9c68bb44c13ef48e7891d570e716875e0e5b4e7e4b6a750e1ee307ba63393426
z193540cd5dbcd0999da35eb84ae52290d076b0d60436f46160806ed1901737ae3828f52149ac72
z6d560735a4d15b2b9d35962730d562ce2684833ff0c5e110f8b8e85719b202418af272feba7487
z643a6d143503c458d29b7f8ea3e43b440af47b022bc3726c90c1decdc8413f3411ebef18fb5682
z7a372b12c0aeab158e987b5e3ef0d8d85cceff155bce9eaf2129afa934bea0ce6e518df129da44
z522707474388f7e75fcc2ec29987af8e0f44e68425081c5cf1b5d26c001542835ab1c023ae0938
zc7b3a73583b0d9c9b9f22217c33da293d5bc0d7f8e1b59f942d508672e443f0192a7141869a69f
zace297013c52959dca33b166bfd841c8e72c19a09f11a7adf4221275d314e38a47384840ce5773
zb9e622e92967f4d466b7d49cec16185dcba2306e123008614257cf326a2d02829933c1c7fcf683
z195afe4b509a26e977dccfe82eb2717cde3ce1d3cc23d54eba2e71fbad171dcf62831f9dfd9be0
z90a008319ca63f825b2d40cdfc627a1a7d734aee1fe20a240bd90f9d0d3f9af0d86edd525c836e
z5050ef0e08d7d02983e78d8bcf34462ddb0b4b4bd7577408a0549bffda60c296fb2ec7b3b8c9a1
z308103c266d30cdefbcd0c068b6ba4ff9ef71037a653c78c03743764b3e22e47be5a2e76a6534a
zfab07e7483ba1a85635d47c4386519dba6960beed2055428a3f0c3f4c472899467e8774d9e95e8
z2b7f7df81677f2647bc626815b98fdd6e171a04c0103d295a9308faec47943177e194f55913751
zff254f259be375efeb8da84e843040d33215a1822e5059738c4164deee34a0928a20462569087b
z60d11c2dfdb6673740030ff953d2d02eff754c3e878703160975045ed15c6ee8cbb6ca0f423cca
z780d16d1fd0a5b999ca4fcff212d962bd2ecf2a0fcdac7d21a6858cf3d6d2dcfbe4fe69a6b4695
z937ef7e1effc89f06b9ccf5fd77254f7c7bb8844668e1ee3140b68c54360655baa1e703d9d333c
zca5daf39a557b18754a480b9e6ad21c4081113d4f9f09cfc54cb5df97daa696bb528f3dcb8c23a
z5fcb293ba1b0f21e541728ec21c0fe9c7739db1b05498ce133cf23a757af44e723dd68dce1c7e9
z38e326cdd13259e513372ee501566384e62efc35e9c04890390e755003a5e68e31115f816d7803
z3e36c57ec12b6a89987c421eb890bfc3420a4186a7e2191413a2ecc4c3709c33ace0aeb8c135de
zc9667e14c56c55be5077470c8260bcf6f0efb8d8d639f9ad527143c368974e4e413f05e4c05366
zd1f6f29177e107a37f6500d088e738af306fe4db41d42f5387cbc761cf2a23836685ba8d8518ea
z5598f272ea972f1f51fff77402bb967f0af886ee6712be5d84c86ee4d102f187d8a3c465b4c1f3
z1cf2cafa4a5dc279bdf1f7e47531cfba9ab2b60ae9dd78a8dccb2d20a72237e66b172278d96287
z9b999d6a95c5593dcbb375b3a138db02a84f615e92eb0808c5d63c61f13e5a43b0474975aad08a
zde3d08fc9f244850fe27cbacc4f0f8d31c56f0aeb2885b18d9bc7f98d83c9f584edff99d7e5fdf
z5cd48e8d40eaf6d1dc993356f158cbd7e46069fb3fc1ba4ea5e98eb937f9b59937404dc001eefc
z75ab3dc852032f732d9f63e414fffd9f0d447536c8a4eb29f66b99cd69c28580928fb59a3a6014
zb8528fe9413c587d1e41bb789be44c593fd197a622622a960d8c9ea9df523af16c9c5db3aa4ecd
z2dc70019f270c5ade4652c02f6c577f23a2900f30a2874966d37cd5095b687db448db37cd7d13e
ze152d525cc9ba857af25c2ec781f5ee46fff2d351fc0332d287748835f5dee7233f055914343ec
z2d296aa4f5999c722f173492d142a93b42918a7c6512caf17fe2ac3e6fe332fbed35503e9fcd2b
z8a7f31b18f9b11eccfffb83eb1fb560433b581e850f359f7c7eeb259804ea91da7d8dd2d83384a
zfb5e8a3c891407328de681a02532113441b04969a9a4d63c42171459eb404e498f879a4204b2cc
ze6638e3ce1415bfab67c8bb843343c77e2118e118cb3ca82dbbec0ab75180f899d8203e5213f4e
z391d3ba19fa9ba6886ea7570e737c2880732c061027a9467e9a6d7ac3d4df64d80d46d9e746f7d
z1522e76f970593e8f54f3ab1f0d91a638183b25a146af3871d1fb72c2ee344b3e94c4e80bbff06
z1f539e4c2af91718082cb39594dee85ab33928283d866aae8e673b70a21fae93c8aefe1b3d8ffe
z3dce324049e5891b803ccbfe25d84d15c61811d08f28e07faacee34a330276edb7b139d4939b95
z0f5979aee997c9fcc35e2de2a00f21a46c8ae290efb8bad62e3b318c31d22d75ebdf8bb4d78f03
z92befd19dd95ac78ac14d9741294017d24ec9840adace34358656da9246a70deaa966365c4aca7
ze92478c77f8d815722b77d11e9d437a6e35b6209a62da430086ba7252ae2e84cb375f86b882acc
z871e63487851edf5ae8b9702a25f9ab47bc29f2fc6c9707c97db1153be60aad78283a6f0464c68
z66c2d1071caa26a41b7246914792c32fa52cfc01ecd43dc785ca3bdda450e69ed377a465c8c11b
zdbb0b2173844d64cd351fd97e77c850ddf966dd888117459b1f730d4c10cb8096d79d4cbba8524
zc40c3361de505760af2668ec7de4bc16ce7b3f15fb1922916ddf1d4bc6bb1e09161e45e10feed8
z3e8c3d92d7a6c6169cc6f231fe8af5b22c6728ada01a4643aff5a531729b03e5e79ecc568cfb43
zd013f3b48f63e781b734a4814ee41ccbd47d421c938d92d90b546d5913fedfe2bf4b11989b0699
za6ff0c97ccfb6fec66e3becfc4a814a0b01acddbb2873e2fb09157120daa61150135a7f3f656ce
zfc46ffe375f1f36b644e7fd641cd6cb4fad1fe56852679b94526018197675e628795e3ca352edc
z322d3f2d8ceb4f381d38366a50f2cf58a00ba6d48c816dd33fbd233ec5f0acf9cda7d819b20e75
zd28379129f512395c6e86f38c7b904e0fa844a6ab2ca9844e46287bba873c330a3689a3e42f7f1
z9e10b35bbb2d8b0071a6a38e06ad6d3102d020b0f6c4109a6c33a9fd96e8722e025bf3cd0d2db3
z547db0aefdc0cbf1abb0db779a1c2cf9a6bba01a953cef611c83c53b1dea2cf24a745e7e392bfc
zf6223bfe01c656275d5f10db487dfa7b1789cb9c111112d48c0ace6425191b67dfb6981d118fa2
z187b05ca2cbc34b1c4a0b47e65462fb9ba518be5e1af326384d7fdcbac81456496bf4327aa4c77
z9b8b3281e505350bf8490250dfa843de8cab9f05fd624dcb75e57f9129bd1675d606c45e1da3e5
z7a647fc7f92dab0d84fe5b9eba85047fe1f81de45d54b2b0d0b34dbaece0c4e80fd237da8360de
z80672ed047c62943d8bb441f6156e62b6e816b08863c4d70f7aab4d37902e88f48ad70fd63fc75
zc63c6f080f45c2dab4ec07eeb6e6162d5c09a4a28284d4f7259528082cdd30c1a9a2a8a50586ed
z3f3ddea587ee072face5b2e725d66beba40b69bff97b9c2f67435652d6a7a3c8b88162d9af8ee3
zee97d3a01b4afdf04f67b6703739f0ad44c1f9ef2627fa4077eca1cf269adc73643be2be59b685
z96a1ae952d0831333a4752c214420333020ecc91a70c7248d223a9f129c9f0ef1f4cc5b4fa87c9
zca9c4b9295e044e24b896f9dabed3ffe38ec06a6aa2ef7e0db7f8909863e98ea9d582ca23d9be6
z84ee460c4677f38041f3c6f998d3ab88effae82f0f8e852787df8475c74c76e2c24017c3946c49
z56dd645debfb0694180dc861030445ec71c2775e499e2eeabdd452c207b9537055446d9c2349af
z1f164f51dbf3df53e03af1bf5aaef651db503abfa7f152857cefde64b45e857837c8d8b4235837
z13af14ea9eb79c86cf2f50b85f58da54e3a2cb7e5dcdd63c8b8197a4015a89bce1f60ab3304afc
z1901a0f3b4c74880a2a69ad792dc922883d6ce9999bc0126083b0fb4a03390a09d81d810f66ec2
z7e4bcd1d3bf38c10385cf088dbe2b89f796075f386e25e082bfa60f4c3cbe125beaa9e0ea5aabf
z0c81dd31b7c2e2ef2d51adbd1ba9f9077b91a84377ef8e880e8533acc96fa560a5b73e6ab5ca8b
z1f481c2df40159aa56c89a3c592ed482585c143c519a37eaf0f581a26d6d50bb3145b384cf814f
z968c60796075058f767269a2342df3d382a65d8c793733933fa4332aee563e3ffb3f42ba8daf1c
zbbf9fa176ecb3ebb2c73a7b697f2573613cb8f36c5d766bb0cd7420ea1acc8efdfbafebd695585
z547560fa633c40343140429f6fc7c86b64fac723967b7e8e83789df7357ed16a7db8e8dd3a3bc2
z7bd20b3d55da76ca55fa913a0bced824ebb9d94fea4a6e670de47d286dae33188089ad41a8619c
za5d3f7f50f75db93ee662515c9acf441c27ac5ec5bf780cd7304065960362e166632e4195b5011
z9fd887731083867afedcb897080980bd6c63e0868e698b46c79fae22e3e8f7c5ffde0240fbb175
z448705ec8d06b9285f1082674ad2fc8df8ff1ac836268626672cfd13552dec7334e25b27a01f5a
z489b3b6d7b3e5852639cff135d9097b74072c33268c94fa4dbe4ebe9155266ea937e18ed3e8ddf
ze651d6a3d0b9e53744ac12277129db4f11d5281ab6fcb47957812ce344b27e273a6686051751cf
z232864ecd87b8469fc0967dd9e746d46db07b3c1ef3824eb5dd53a83b35d6c4d7d107ff233d684
z66171f0b716b5a4dd1775d96ed23499d1079723110d7a534d16f99e891c2a5561ef19e67f5d5d9
ze118e3604f1ebed2e369bf4799d11ae5eae96b22c29d095f0dc2f163b44c42f689ccb020595467
z6f97e227b5486ad788f3633149bf4089949fdb62334802ba78d901a880963d745410bd2e612925
zb34562b7c56ab16be2178b3fa16c1a5fa8bd0019d39ba0cf816e614e057f16e0c5fc66dee288f5
ze31579a535606428f11c9e5f34195d2f75be9d61e6eb376f625ea51eda15e006f26bce677150fb
zf10b840fdd9d751aa9c9e65133ff7ea455a09046ea63b0fd15971cf6ee448c26ff2321cbe3d43d
z8bc51010f4a7cf6c5ad89949f61672f700108ccf5d5ea0e92e4b64c3b348224bdca85de5dcb22a
zb79ad0307a00b52c2d7ca0fba148f8e481ce3d48b87f399da5b8d17d917dc8175054b009e36cb1
z61ce3091cd5ea56ee27e7443b05f9a6c58112cf453fab8eab66021a96b7b66a02afa9a40c82d91
zf9bf98d444a266c82d2f6ac9b469a176ad5bd6a17c5a25a9c575ee1b58c2e0dbfe06ca091f0b18
z83820686c3088fb6fed68c2699903e4e49f54a32522a2f14ca756f60d421e5c4b60b65259d7d5b
z4174167ca3493fd0c7ce99de91f82b8f16bb7e277d99d63708310b7234e8cc822d82bceb3803a6
z4b360262725c11f4b4acf70400e4010269d4f04ab16de5c874ecb51acc883cdfe1f87520b67516
ze8c13768343fef01455b1173a319feb272f3ade6354476dbe74cbe63accbbf6b252a81bb453629
z164a9da261c921e264693e19933eeecbbb671e2b7cd71aeee5cd6a9db7ac54e0986b8772acd82c
za39abc2f11fa54d78700341d8f4b3a68d605bcf1dbe6907394588fbd2fc155a2c50a349c1cdfe8
zfae6d535282b127118fc87327f0d1fbca09b4ce56b173637c27fc2a270ec6aa709959080dcc033
zc94a0423daae44be19c505361902319174530ce034f25ee193343776d60a799a3ae6838ba5cbcb
z86bbccf6feca10542999e8766ba6dc8f5409ebc450ddb62ed0f4c4898275c309ec2bdd107c1585
zbd6141480af7ef128cfaa9b21c282dd9c7c2254d75e264c10dcfe6bfae8cee6d05e4e5332b6547
z485c44a8893fd164f9083233b09438d627871c3972c2c6cde6bd66fa9a72af4ff86052279fe75b
zdf9ca8ca50a7383391608114bcd63edf4799423148c27507eed794cab88a6ff3c851973fa8dcc6
zb38d26db1ac2aac2be697e385a77c550170ac56548fd22afbc7d69e6eafb0555d5798e2e367b89
z7c1cc68879d71dd21ca900df9aaeda527093270edd7ac8d4b99391d0007c7e47d5358c4b3371a7
z90457adac3c601dddeaaedd8c794702dbc3074dc2a3c448822a5b67ca5e951a27c6d7f0e4a6bc1
z66b995cad8dfae042f1beec281ab6c507452eae720fb80c6c9f4eaf71e68520c9fbbd2f0f2b875
z09122cb993d4f2ed53746ac74f1ae867f1444e0d655e44ce678e922b5b8217b0540b248335eac2
z587852dca134578b994c7cbc365e4c1964816bfca83d4f17e2d4e89529c9500dec54290eb8884a
zd045ecc4dc296d35e5f6581845e6eeddbe04f989967a1be795090d5b1c60da69c99e8997faaf1d
z2d40ae2dfea453fe763652b3a5b903d19794be4e2bd01123a59b81515e89346c141871e2a39727
zf8eaa218ff05b5a0776352d6e8946f86f52975e788b299e9624a6fa45b695d907760a4dc28b9fe
ze0cc171048c62fc7dfca4720fc12c9644ab28b2688c2d72648dcba57bee05d51c3152beb4f4b07
z10dbedf18dc1e5e66df990762b4cb9b3ebae419a92ad05b677912057f9e0281521430f29de5034
z1f191c40127f92f2b768a17f11b9b9753d833cf84ffc460079fc0d2a4e7a25418d7f937f95697d
z96654e3e0790c1df01a2254a84c9e7408eaa4ca3a68d12613dda9126370ef2ca6d2cc0810a8e91
zc6448673fe4c5d611ed00c78fc5da1af53081bafd68a168ceacad2da02f661508b160ddd3111a9
z218a2eef50521b7559b41ad54e77f10a74b857b5219e90eeae749f1fb5abb7717a858cc838c8af
zdb13af3cce5c7b844d05eb3d21828b4b92cb1e759e3a60c178e952987b64bbcc0e2185798dc29b
zd188567ba475b6a62f4df917863f40444da647b8ade1d695996cdabefad95fe8985cb4320cb133
z6ae37342a9112cccf7eb655a4fdb5718c55a196f646bad7012d5ee67fc79e84783a46a4ad4ae2a
z7a6835e3283d4a1d38b7beb01da4e4356d956b39042cb841d3c12390207655fba1d2ae56ff663c
zd1653aade4b25e86a74b68e11cbdc98356054ff9f1a6b1827fd587a8e37474730d33daf4bcc0cc
z25581bb6eeb7b6a1faeb97597b0228184d59ff086850d32d35c22bd99b9dbe6b44991b352404c9
z15ad5ab3f95814d8f29e4a79aeefcaa658e7b42054d1dec3e7a685c9a73fc1235dff699b0ff472
z4b6286b6b3cff4a5c52d0477b071bcaaeedc4cc6e069655850e5a9c63f8328557647655c93b2d8
z628c3305c8c2889f10caf795a2f0b0d5ff5b824e4b259c3516701d95020774c3d256e4dca7e1c2
z33b1f9a3b79f97c487920a2345ea4d383173eff56d244637fdb2432ab75c337f7b8a770c737fef
zb5f4e1e745a16d6fb77de4ff942f751bd2366b334cbe80e80d4744e4b1e8c0ea7148eeae2fcefa
zeca37d70b4b7bf0f482c32738c85c8dacc85ea068a41e637564c72b837822713943845b436a305
zbfc65b0bae7c84b0db01a43872acb2cb0e932b5c1d21c6bb3847d3083145a0742cc0158d6719f5
z40136a09783d6114380cfc35fd101ebb70b4e84e12b973e4b82fd003a70cf4e8f3f7934e1cddaa
z1b11d07603370ea68fcbc226b597629f9678f7805b92eb2413b4049acf9074b4ac3a2755e37218
zaabf1a012225b0aa2da2dc0e00c6563a05c5a4e55d5a05488c4a2831e236d35e945b832b8f594b
za5cb6edf599508de60ef88250d1890cec2b82395d72d09162311a68791fe9da9c66a241ac8a1e2
zde53900547e3cf24ea2ce20ba6d7b568180406f5c432a6c59cecd8e222ff1e9e9729bf31d73b4f
z5a2677e22fb234eba7d77d8f8085fe5ef9edd8ecde25b8c32f19d31dfa6f13544dd0ce50d2bf37
zf3c7570646609925c1a05da64bd532157c4af873db66ab3c3701472cf36d41f6a32f609de6dbf3
zc86b6ab63fb7d281f69aad243b0dbd359f73187745a75e09a1b8f3c6273c3f4a5c618f54f96ed3
zb28bb2ab639017f4254b113206de1651fb956a124e9458f01ade7302cd00a38251e4f5e8b69a22
z84a6b212bb5336fb10ccf8d74adfb594db8c1f356700fe626037454c23b37cfb502f673abd7626
ze2d3a49a3f0ab613cb373307aa97faa5710a17d6d070f73a3190485eebc3ce34c56c4c563c709a
z9d8eaac2b7e9d7604ecfa60dd888024f3b14bb11f1b4a8999a4d2929e0fa0f8339d1cf313dd17b
z3c8467f1ad92a6e3553984079fb1adeb044a4560a951cf69559fd88fe4917418a19a167d7dfb3d
zb57c66467b7ca1e474384fd3aab1e6fc1074ffa3cbc32be1ec615e468cf8b0226acc0fcd498684
zefce137d047d19acfbb0340c8c981c09257d5bfa9bda4dba89b61bb09f432c859164abb2a29894
zbff9c33c15d8d8dd0c774cd3c6213b627e941b89c0164a8c813ed64e5be044a77080a81aa8d914
zb315fcdfe4d8bb3a64014b7329ae5062204842a178ffd330b78ae119e22ea2f3ac2c4731a46fdc
za23ef714f9273fef4b351d5b6436e69e137d1e5f5e0ff84f2d3e0f28c70e905e1208c01dba8cfe
z736aa2517272dc31f6ea14bc29c57b3c2f39d3c8b60b080403118ae4d9456ebd3a90e8f672f7da
zd5e395ea77c09d7dea47dad07801cd66cb64d5996d75e7807b7589086dd1806588549ebf994764
zd9066954f3939ccbc2e898213a3d15fa1c4ddc46c834821bb50c8dbd5fbf6943d592f7a8563e20
z528f6503de1ebe60d75659d331f9d0f2d9283494724b74b52334e2dfcca3caf0c130fb153f9a4a
z9c41feefb364a170b94441765cfba0d9f1200848654ea1169f03fb2dd6d6495417f3e4c5ce176b
zf25555d989d03bc04286060608c2f1323a4462e1f6d2ef2cf997bf5b36c2f69dc7c135024cbedf
zf2d5c43baf02facf8b915a6c0a8d5cf324a3cfd9fc019caa5867239aa694baeb2b9a48d05e0f49
z8902d353d936c8a424875d99283040be7ff72de6f259488334f5e65d70cc302ee4cd98832c5114
zc3655fa18bd5b8e6fd2fefbb261efad200ee32e4e64b1fbe228495005f0bb0fbfce4a3ce42ea2f
z9c1170fe1c5cc418423e4a76aa9734f1ac2e93b2a5edebb3a7af2bcbec43a3a257236aae300b84
zdf6732874a7c7b93fb164e2167197bac2b8247e7cb43bc20747a4d1a898cd1d3d2023ff037e5ca
z42d81cfa890644719cc2344ee0fd313e5a1b3399cd6b4d58679edb1fdb53ef09240c0082342235
z281596936d3bcede89f2ae0059ed99798978abddaefeaa71127c1477bf15d08c9941f60e61eadf
zc37b19a51dc206676db480dcc609d03aadf7d53f5ac4d74c87b2a79db2ade943a4dc692861a38f
ze11c4e731f07cc790d476ba18dcf990758e3f8a869adf0183940b6ffab55a83c02060fe90ac432
zd0975575eae3fd14d09ac221975e632e9ebef8cb2c31e34eb6dbee187f548bc3fe465d1c39f24d
z66c6010b0ab74409ff53bab8e3d6978b0a8afeb68f12aec24a5b4ed2d55d058752a4a920fb3db9
z12bdbd995d3ecc94781605d3ff511939bab2cfe927b683ff6d5469ecb7a489fdb4859fdbcd9383
z5a41bc26eb38460707fed2ef92e0b323e7c97a30d23726a47951a383c8123b37347702cb4bf6d8
z9955a160e84606a1164d1d27deed53989c3625c212e092695f3b1e784e05c24b52c74287d5e647
zecc3677b03cfc33d70c3d6a8478425d7242d60b42f667f4ca4cf40b0cf928e65f747ccd5cc18df
z326c71ccb33ccabbe5d412e499952351132c1ca951fa181e042a5cd4f5c1f9ab58c48d60f3c976
zc3e18d248101ce9febbec5b1548e2c62f5dbcbf87d8888ef4e5347a06b2c566ad59a23d93951b6
zc6ef92909c8e855f3aafcc3db4f9dc36bfec4f3d72f6960a4e2f0c6fd4d285802a17e27cea31b0
zad13671889181eb4e2b6b49f34e7f2aeaa4bf14ea2ecfdc8b6074792883430965ef76d4f99a674
z2b6f27ab719a9790a52787e62a0ed41f72e75ab404db06cab09af38468ec5512e22bd3c17a03ed
zbb79a341f3e0e40f38a65936c536dc4724e93f60c49d404a5796809c9a4a379d3e8b18c8f153b2
zdf8dae8622ccc78d413c6c3e1bef7139dac0c222d4f410ab942f29a926420b4b93e74ce09f1619
zddc77fe1aa89d16cd25f6b979a3cf91da7108df38141cbf1465c61241e441d0822074eae06ee6e
zf8225f3328290ed379637efc56493e6dbf30cf0bdcb96c696c28a0f67792e83d3f1ea44c7e687b
z2ceca15274dec405ceab62e5b60e4c307496f007f621e87f407e64908bc682fb20a57e0bdbcad9
zcaff1b13fa74c3305da8bd76bd59f6e0bf1483b7a9d74fa70d1549ca9b06c4a856f11d2eb45a40
z13a09d04ade6b26e826c6cfd0ed801c096552cd8e03436af42737128c0bf88389e7f3b3c027f32
ze2aa1ac33151d32081ee0d2f2e78ea61c95579777619881bfb5877e428eff256a6ba1ddca1beec
zea8aeb5c814016d5b7aa36c49fd9dcd031a6fe40f13a888e6a898e857cafd498ffd98d3b3b32fb
z16a613ec0c0a2cab8f962f5708c234f53cec9a5c49686f293d52a70e5d87bbe6bc5f9ffceb5c74
z89c1427edc7d3a667d000d0294822b3683da655a8ed4d7f96261f41d2d4ea05e7ac43efd7a551e
z5d6bde371aed0420590691471a38058e9d97802bfcecc901de5a999499611def397dc635fc60c6
zb6c3dab9a76f27e80dbaa67eccdb591c4a1a4b9604d798e23e843d8ef67061b67021321797218e
z2cb82e57c661502b404d037deed0d8aa6b90b39c04ddcaf308bd3feb61481bc707c5cccd91b42e
z6da140d81dd124e17a8f25607c781972ac03ab1c2c91a2cf124d35a4c0f3ca544aa6e85fc4150e
z9db785984d8dc5479ade2796f2966bb5e3d057303bbc8dbfcb2b6f8ae441838a2625f95cc378af
z07017d00ed3f22412f6c14c0836153545f7a20df4ad429b3faef7a5f1c8d3b4ff5a31d53e7f0de
ze89b23a3cbf385ea7d7d52e557143ab8310a892d1e50cee2900da9d59a08e7f755a5843b1b8535
z45e806b86a781cfaa5ef1ffd9cb7e61a2d6d716e7be57083f5a7c55cef00ceff298d42e3f2767f
zd214ab0b39859c741811b0aa46b94b6d54e48115d2ead4dadcafb96adf71907753c638cc843f3d
z6ca64a379580ab9e6adeda58e076c265a6f5b38f9a2508f703852b8a70ff87455fa275b9b2244a
z68f70a5867ff687a9ff5b9e0c483cf39e096c9df9ee69a5335aa1cb8f397d0077d95dc9bb1f85c
zd62dcfd91f6cb7340d4398fe703a44e7b410489cf274c79340c5991948006cb71a0c1e31e96067
zd159b8a3277543315aefed8fad480efd1254689b281ef38aec410b48b74fbc5dee78cd46df1048
z302e7e4f637f482840e4a7f9148f133f8722ae95d8b252336327274a57d36a96d8043b8ba64544
z2f8a55ec6c693817911939d7d6b708db2dd85bdcadbb52df015723ab8df89c2058d97c50c4738e
za2b2cc0f015eedf9ddb34e24fd8b4fc87a665de0f66e281202ed8032a3e38104b2a6cece5fa0f9
z8ae97be5f6ceebfd251edf445170eac830f4682157c5ac431464a503151c42a8723565ea6521bd
z7dec51830a6cf650e948767487c32ef47bde0fa91ace524efa7564ae3963cf81905afd1d52ae3e
z0345d350ae514f5f56205593213b1a49b0387c7f763ce63d81b6465ca41175488643673f139336
zce79537c3ec2bed53fd458642a0cffd90ec459a26f220a573ac3125502b44062ddadb6c8f36e5b
ze5ea8a521a5a7126edc6496d6f2a0790001c2b93e3ba6b7dffab1d1a81ae41a4f1f892fd60ca85
zf7e9976aa78e6b62cde0d019eafc3b140dceada24b5768dca90eb58201b6cd004fa99c8b633f27
z729c3cd9d55a35201e052d428026065625067cbaf1e2a45f28f14694608946f5563030607f8905
z27484b0a61c7ab39e0dce210da73c5cb4b7728f4f913e52b2ea57c3aff9f57e76f50217120aa6b
z990483ecca7f3bcca4ddabaf6375cf3632e4c4df70820a36e653f2b76dc3815d7d7d5e49fbd33d
z10b527a55db50d0e1a7baa6c838f2a1d273aa3689cc03b0f67c4eb5f94a20dbb44c2732cc719e9
z3e62894864290ed8ca3a9967c73c2d677fc975ebb364b274dd9a8e72164bcaa596be5f1f8e8b5a
z5b190bcc1cf36d755622fa9ede22b5c4fc48eeb647772cb72d3478390615e95abc6099982836ae
z2e43cd02cadbc5abb501a55f2c301fae685d23437dcef56bfe8dfb28e7ebc3e8cbd2bf50dcc8e1
zf10bad64856a688f6deabe0cc9bdf3ce2f2c95566bc33641f88fc734527f365a37a5b3fb229593
z08bbfcda35a1fee07a384875efb1423e185ba8178c33f9f671c07adb03c753dc8fb0ef0a4f45b4
zb90f86042633c8d2501910f3f67e06c71a652acbe7ce589a1cc91062ee773df9bb74f50651a147
z3ca5ecc735ebfc70eb902b71b9cf376224164b47a1074d204fe88a3b5087e665c44bb4056ccf35
z235a1637eb66f033f49b16f59a028d2393b0a0989b70200ea2d2f640c1bca00eb821835deb2bdc
zb36fd5e095090511f1457cd90021ba4ea3a9a0a15424090a9726965f4288b8e22dbcbe8a11224d
z437028ad644f08ff13b533a283c691bf37285711087c8c3ff565a74e182b6a0d913d0ab501e54f
z64d95408ed0b8fb22f855c67bd34d1a0f448b06e5cf969b32f81947933558e7fd36b6c6182b81c
z01d90f44de8e267645ccb4feaddae7d3a70ef246d7e6ec9b4fdab9039e879de3da3ddde8a506d6
z3d57089326cfd8933d39ac6e8cd44d58da9db00b58e96d72249a6b5eea16eedf921e440a1ca1c4
z7c202a41424284c58129f91bf3df8f96361987cb825f5b9f82402fc377f0f2d9ecdba6b545071b
zab6c35be69c173443ddcf32fd5953dad73ef6be14c976f62b42a880f04b24797c49a6065f119cb
z8d92cb12f112bc0152f414695fa1eb0115d078d11fb22f3bf47a16aef0df6903c5367e609f36a4
za61a0a38569d8acbd0c4efc04596e17164b5e6cb8d121a1fe5801b1705150cbbcf0fc02407f654
z40ed9ff932d8dc4bec5133d7c7b67354e7dc2eebfdc6fe44f38c83f0a15363e2c82eb5ba829aa4
zffd4a4824d24c7e2f774151d9e56d2835fd567ce867986c6dc8a9cd4db4c9418947d6b54d96393
z5fef771155114e4e63ed0791180812d1b99c08c889777e21ec0c4e5ed8eb61f6c4bd945fc779a6
z79ee206490ea489e660f7efe6ab7a7dd30c1f86d08d40d0687743f9a708adf6a6fc0d96b4440ad
zc2aa865d3eaf414561975b289a389ce7d7e3465ae045f16c2ad5c9bf66e71332151a17ca510971
zca8c1d4cbea5b833db198c6f3e105e6030b89ff6f9349501948301f9047dcd006e562bec36a668
z9a09c47aac0c4e2effb05f1cb184a8054089681b98e362c6af3995dc318b84fe02d8db1ac79614
z42f343bd25a958da115a35b1e1ab3ffa81340df478b346c3a814cb77fa2ff0f8c8274b6571c95e
zcb2aeb8be84101897a31cd2d23f3dec8aaf16230fdda4b93b4d2a001e479d47ffe660f0e15581f
z2e72549a493247b1b6d1e5b311b11f7dd1a2269e8c14ce29932a4f479270f0cf7d5a4dde178bc6
zdaf3ffa8f7308dfaf365e360d2580c7a774c39db1990f35e2693bb5751bf82705fae7906bb9d43
z88aed414aadbddf71159c9ae452359c7f39507b4ae4e03a094c58c3b60cbf9d244a8f427f64ac3
z549f91eebdcbe694717808dbbd9f12b1c302da6eef02e01b6aa8c8a217525819ad1efc02bda223
z528be17036e2a648aea746955812ffddacb36576c9c9e932e5321eb94d7948c70c0f720316da69
z52c7233be8a523e99460fa454a4f010e068f258219960cc790ada29e13139710c4954bf4c62f34
za7459538d88eb5a8c545a889d6c302e8403af2a2b2378cc90f9e105cf951a13948a82f89625d69
zbfae44faca4555329d20019d92d4556904932b8b6a8d246be3c7d487bc1229564660a98fe4ea79
z6ae16f680f4531f8a99878740b7ca067dc67a8240a92bb6314003f425f0d429519774dce69cef7
z93a037bc6e469c011d03238d71ae44b7e43bd2c0a8692a7f172fb193d5ac220063787fa4cf3452
zbca83088df49cbfe7fc962800da7a60b65683c87bc2757edb6e26aa385fc550d560abadc098f45
z1e9a79bc31799c4555e0722f5fc06969c6129817a471c99607be1de22a8f13072a7f226158166c
z85a567fef09ab7cbb1144efa5b5f2ee0aee17ca3715d52dbc6722c9ee63f1056e0a3fdf2df2b93
z3a913be582feecac50ddcbd67f216b937546e5f164d1d39f03c228d40d7680f2c8c34343eef4eb
z463420bdf80109c9529db775ec8a5c20cad51ce56f511a1009f9e5c73192214984d6df6871b295
z999329b9478ef87e8cec28feaf33ce4f5c7d10b291f09cd7fa5d7b95ae73b5fd527bb34ae2e9d4
zc8637a6f04a0aff310aa90588aaea2e6034ebe1edb405a3c13a551a3fbc6f7ed004daa68e660e3
z47d17689437503f205d514ef052c0d470de89e87ee63ff7b10c3b7d748ebb0f40e84a9822bd7ba
z756dd451729c2646589359c2022b0f1780f12b622882bfaf34a2296a30d5b3971f5154fe6d2874
z5dfb8712e1f3547eeef4d53d82175793d08753429a7281c624cfde67cfd95aaa6b11f38a7b6570
z554f2dc3fabcd25cef8afb5188610521062935945c5eea9e348d7ee82ca84c4377ae65780025f2
zd0dd061e5378a1afdfbae2578b9f629026b975e29dcc3536025d04a10576d0967017803bdfaff8
z06b4028c0ce5b759bd09a351800cc14085e516ca7151bd8f5b4f804eca1bcd908204560c81d530
zaa7f4eaa9e8eb38a8892da9fda05f998b1cfdc22872eb0badd33db60e2a2aec65967a96cd40466
z1c944fd13123c88362c1b65ba166874746007f9d4baf2032a5f0208852a2a7f27dd06768bd38c7
z2993a1c5bec4c9eefefb37d4ab6f008fad8db3193a219435e79976ed9b6457408dd2014de33950
z0f73db28c79abea2212bdcd4ab6f97e4a304fee0e4d587c045d866a2345b44569481a2e78c5263
z1d32dd58d0f685de45ec850b2f78e8f24b9c49d3d0cc5b2b3b9937a8067501cda72c2a7f3fcf05
z80f7562404973a320c5bb525f2874bd297726d712de239beb357ecf2f845c0135157d9f455bb84
z1766a569cc4f02b0dc0840267c910dd94f2e75cb40ee31fa79d348c1a1a89204e20bd595f55046
zad336ad7391af96f1b19bf58667e8b7d68f5b816feef903557f432c14af744f2aae67909d53464
z5980fea6296dbb8614a798e808987179512f3bb77102b8a6505114a01dbad701372ec624877033
ze875c92449af886e110273d636837e7965a321e12a5e2b48668c4b65813cb2a7310f3aeea72a2c
z2633a49d81b3b7d3bcda463273850bca007cc0470a4ad65c70dc6b571f4488f478b419127f9f8a
z67e549c981565278154dfc766a75eb3b45bffbc4589a09b88fc65322a4579d757dfdea000614fe
z2057a554688b0687754343e89b468586fcb4fac7574d2cc94925364421cbb57d72472328c7e12b
ze7c706a831881d5c4e74365e3fad2d2451b4fc1f520d6514a5fa1e08145267f938e7a74d568e02
z47134e6a67a218197b36fbc58233fa2c19d17b06c834a3e18081c53f8b51143388071912036d6d
z02573696d089fa24f41507778d3b69b65802f7715360b7eba138608683bcaeef98faaf75a231c5
z03321ba426c33c9104948ec9409be568f955c73cd589e0690aebd85b7b61a4e2f51ea304449d7e
zd8136df2fb8af50ec6468732b22d999f57231bc50469cb2bddb15d74bb3ff9af6a06fc64788e84
z591def74f4ba22ddfb3238c70418691ee9453a9c4c01b6adc8539fd93566fee14741ba858eaef4
z4bff61e892d356c003259a5353ff0fb260aec8b262379a8965e5cea5b8ed8e70c12412876a910e
z8275065f6d7bb2be1e81ad30378a6b15cd8342e3ccbe49d5ee7b494ae2834ead96e1f4aa7318be
z4941591c0b2177a62d1467f2dd8a8bf961c8953927647b096046036b3e455391d1cd0fe1c6d3d5
z8f9a0c3a2042b41fde7a725c63d5b64844579b58c218e3ac8a242a7adec02d04dee6935e700c40
zb84addf3a9bdd4c887152d8fe4279bc534fc3fefd4ba215de3877a43162600d79f82c0a8314620
z322cac20fd784bf0eab9283e0170a1938c69f52dea29639385d8ff3ef0f9deac8714f7ffc815ba
zb274fff510d4c14c244915692d0285ce664ac0c7435202cd7eba298af87653ff97f497746b2783
za6c9db5b7dfe8fc74b8a0695ba09a965ab41b50eb269030b818a8543b69484e323274f3c9805b9
z219b49ee5d79bf019b1e0422dddac6194c5dda1f5bf59a0135bbd28f6a3623b699a2bc0c854afc
z43524f0a459059c51f3f9688ba547a716a362ab4249e0143ee868bb00a5a6fcc5d1166d16dfb26
ze604d4a59b411127fc0cf6e07862ae3f43d9fceea1d7eb3f0c226f00994f65c9983f85eb4fc807
z9490173d900d10e027ad61238d12a46121789a2d19d0c9812c09e652b676fba76ac53f53296404
z851b59ee335f212b4ad28bf887c3d7b05f933c75c1f53e25030583220b38b29e4d60bdbb17b2a1
zfc4b5b252fb43574f2deb5d5dda34003c08332c0ce3ee4b97dc6a58effc400c3510f896c590916
z0b4f10aff2d8b117638f28a5527e0601005c7b34c6b35a633d2a2392803321366c1bf7036d1408
z0382692734b04a70364141c6c69eaabdcd9e41da4d67cb9f904bffee523cfa581426b5172fb379
zfa3726f69f5d5ba610efb7f8ad70cca58fe0bc90011843718e28b32f895d577db0c5842e301e38
zc6867f321fe41020c658603cac0dd1ccf16b3504daed0248fa00b4d373e115f228c79f1ddbb207
zc7e8c7dff4ec941b9a2abc129c5e0a4d1ebc616e2d43cfb7c86d5dcbc54d4a6f285f1c1e88eab5
zf75923dddcfecae6468cad63fa33e739a52f7438097a589c41d1812ea60b7a0d162c21c3116656
z12b387a5a4fc34da6610ce9d9670ab60a4dfb302aedeefae993d02a47eb5102c8ee0f016fb5e58
z280133462a64d0b7e14df3d29412ee22a4dbf093450dcdaaf13e532dcbc2de6b340e19ac0f1f20
z727eb3669287ec80a666060935776fb6280c815751ac62b14bc85775ebd64612614443d5588c07
z0400bec50a129e8a4fbf9dcfaf82dcfc1af5d3a019222f569d4d9ca5889b30d297ffa287567c4d
zb153d9a4cd9596c91b30c1463c9d3c923fbf12e90402f6cee59f1c7de83959bac48b772953db0c
z019aa7d42a425a977870ddb348c03b4623da0125a4a9b16e12b018609a9711f180e77389dc2ffc
ze4cadfd0fbf5d09836c631654d2745e9b9fa359cb07ef17e27400dd04d2f45fd99a73cf091b7dc
z1c7a0dacda6c0e94bb074c4590e4b5bb41a6aa820f8c8c6e8a3eba78db404e196314b1d38ce70c
z7d171f53a0d865ddd5d3a9d0646bfa5c2015774bcf1cb7844ac8ab4faea5ae579c1e917b831437
z72824810a2830def94af92857a50a11b6aab449fd76aa2c717af5f03026bd310bb60731ce70369
z2c6c383ece83cd7a064f1481bcbb1ac286f5f94fd6c3e67347b4df37ebe85c79922a93355fc220
z12f1bda91ec78c360324057ca2f2a91e5a117ef1413135a6404ad540ceeb15173a4d788e5bfe8e
z083ac8db5098499b11bc77cf0b404bf5b898306aa5cab8e5be86d100d16a01a0b0de24f7afef38
zb1d2b1af284c9fbca4af0137b274eb0980753ceee1a37f0f7f4c2ae4c2e803844a3eb9771ed91c
z35951245d7a43b51cf55a8328077e98b34a96bda7ad5465a520b337c08af85263cfa77e28e3770
z3497e65e299ac4ba1357560965c88b6688604d2d056e4504e25383b123dac12f04a5f00981cda0
z923dab5ffd170eee1f23708170fe302c26e33f45d7b730424c6b077e92698d7beb605aab159eee
zb0a1b0a6c1015f2a420104d56d7f57e87eb410fdb85671fb3f230a1870254b4acbeef42d87aef3
z6e40326cad3ba714786e61711fb82f03d3e749d4a0574ceb1b30b7a8a75dc62961d322c8d34fad
z3c746af58127928dc5a9367035d6005bb4432be2d92fb67cce8106d9db81fc4b95f390d01305a3
za1d9ec90ffdcb706bdb57a35912551d3cadfe23a7be2ae8f7bc8f13f96872d2b8ce09a6dd1ffa7
zdc11dfc91693359bceba2c515e5c2d
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_sas_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
