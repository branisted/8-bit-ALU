module adder_8bit (...);
// TODO: Implement 8-bit adder
endmodule