`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026201628cee5aae21fb892db766c4
zb5b1406e11aebfd6dfacc9da5ec03b70c276807a3eb15e28ec7ab1dddec42388b9424ea285623a
z248195c9f894b36317ca6e59c86f11031163f5f5e0af432ad71a370b503d5afe29967480e0ac49
zcf7c756f92650aa81b43bb5505acefc12a9333c15090c386c323f8cce4e7934214caea9fd9c42b
zdda79bee782f6c797ee18b17b0c257e45bee7908de093c385d7e8a753e689ff7fc8a8c9e7ce08d
z05cb3d56bf84f1fb3473afaa2d473467ed0a852501771349b43fde42b4344a1328f0b9488ef772
z0ab2e71ab13ec995ee041d04202d900d95c299a1c207aca6e4735d4f3857211f278f025542d047
z1120c7526d7c7aca9b4535ac2a7c89914a071ab6e28ef5a017369bce3e9ab2a40b1045e640a03f
z1eac01f38537c460592b18e6569eeaf3cef2c2394144d0b4682b5a48720ec74e4d0b2c6180f2e3
zb86b55096a5ef9be48293937fffbe514105bba4c72b420bddbaff7c98716faace082ce2b7270d0
z082943369f9adbbf070172be89ab7354b521930c5a900dc87238b1766e67b7a0e1191854639319
zdf1223e075dde8a5cf288060271fb236b0645c68e01c0ec3232b83e1cfa0e95b47ff1652160747
zecde91b28ebaf7a1a398cd45bce9bdfb59d8a39c019333c8c70a92757f3498ba94a1700a22cdc8
z871aa793ad3267f5ff895ad9188610226db47921a6b2373776668a9b2bb5daa92fee02383d142c
z8b55f881e25ed88fb59ba9c730d78bc55a0757a3afda6902bf697868acaaf20ee3ab8a85200ac6
za186225ff0211433acc05f5df1c2b0c330e70a04bdb8ae144ddf093ff61e1e143a2dc7814f5445
zda60f461b3cc96c31c3ffe91af592ab64af298369479c6402812a8f0aef1298bf74b9348aad66d
z7096e30f35ea4205e6181575b95d59b1704055c6530760412ce718eb5b1e106fd6a179f4165d39
z8b30846ff76b49c610f1199062e473940596e20516e2a4d93413f9b79c94cad57b5fab211ed856
z7548faf36b57164d3e598195148001d10a1ee6944d21f69599b7b4002edf2846bfb91c88304bfc
z7c2ef11e4a5d4955d82d2f79e0f61ce32e3e1a32d73c6aed2779ce5d7057401c0b53a1ce86b67a
z14dce24a1141fd5577a376b61629ae692164d11b92077cd1cf211a69967e8e2507bbb7b018c668
zd3a4c8bd78ccd7e3256918367dbf654b6c0c31f9fc3d170253249aace4f7db3b1940d44f44c9e8
z4a1c5b5ca99c3087c8b889dc4e453c650040afa921ec3bc79711a8afad1e6700c6508a487142d6
z1b495436115e5ec58141e54bbb74297e058d57b8bfe505d384b0857689cd22076b5212bd3ea481
zd881d2594bd9829b0183212fdc49fd49b234b87dbaacf31472edcb89d34babfece7ca2050259f7
z9bba58c8d989b4e472092233d94b57dca47dc69c547969363949ac4e45dcb38c20478ad0f76e52
zee812be562af73ed06cbbd1afb19bb37840e41305d5169047d9842b7f850acb1cc71924aa55fca
za56ecd97d5d2fd19bad64f8e43fe3326b6e2ae877a910982d87bd0d607ebc539576f81096838bd
z032f50eea83ce5060df70f577ce5163a92a2bef3b59ffa4aa098c7a00b39ed48748b7c232b4e43
z1fe32df17673251debc24f699efb28168714094231f3a47a9cf70fdccef91cbc3882974cb5a59c
z9e3e019bf96b1dcb63c025425e149b13932511123c2fdc1b697818a84f23c4b899f717dc37633c
z71a63f60774e9a418056c6156492e7fe7f8af18daeb5b3c81a2bb7263f7545eb66317a0b216bdd
z1d7fda29344c9dc228f16f133333a1c4e471f1cc04aef3f90884acefb698424bc6c87b09217bd5
z868120a3b350c3742543ad1b3960b15b3af67bacdadd7fe47bb8fe41e96d14524b97a1e88728ae
z25bd8a4f76309d1ca4ce35f4c4d8d78ae5411bce4f761323b91412ff88ce7b34795f25e9f4d30e
zf4133861f84353669d9a81c7dca7ee2b306a62de23f17632d7792479c2d5acf9a6316e0d5d93e0
z765be2fb1eca748c2a6645205af4c8d9d7c8cc9a840ec8307d02118facaba0388f05df3223d6d2
zf2defa5dd5796e268630731f48d471fd9f16a9ee151b5825bed1562dc5160424ce35fb74015be8
z80db3721076d61e2ed644ac939344ec61a33952e45998f621994ed20760b49849ff1a3deca4abf
zba334e4ae5dd7d794496b458e2e9ddd582a41d0ecbe5e45069072a209a08cbbc5ee4e5e6f5512a
zca68a86293df4bf3881f737a33d8954583ee4fc46fe4e7ba3a8867ed88afe153393cf470ac4d67
zefe5cf87a143e7abff710ac12309084361b46170d540780dff3fbf21312bd3a28048e618cf27de
z9f1807d2815755af6079fce1c2a5531fc98f51e91092bb8dde3f55e9832980b40a0f7c0875fa25
z61be7d40d9b4bc160cb8d3cb144d916d25d3548123059a183d79a9a132af804a02cc548b06452c
z63b3aab32df32f3e74e1c677e54cdfe273eed1856eb8c5b033752423c57ea0c4a22367a539d0fd
zdfe2a4d751a91c0ae87ce35cec2e1c8fd636a3fc922712a799e9ce96485d9dc975d64b1f610c2e
z86aed5cd184133dc9c19c446fb2d293e67a11d04d84fa9cfec363992da7d601a362c43dff8c467
z4e159cf9d05011d57e18051dc44689d8451d40d1c3df36187feb3f77a08643779bb6a11068ad81
z47b4c6ee2d0ebada2ae266464ebba1e4383f6731460493be17493696aeb992ab5b8ca735154a4f
z58a3bacff7fcd22d75970d43a1bb0b1c2af32768c979667ad2445198ff998d16c50494177879e3
z1a7d0e264050fc7395ef8206b590b8ab6cce2ca633c1b2f123d227c33da2761f99ba8b83255075
z4e658ded24e3afde7f8378d2058bdb094dc9e9f8262121fd556e616255ecf65af21a134d41b4e5
za221a31670ea5a00a43772533f91d1e4dd6fd2b007c28c5a53351960febde743ab7c70b47a23c8
z237ec7eb3f584f34abd35a42c8f45bc822ce2e891bb5d9ffd43c6de71a4ec488b06c558ba64593
zedcdb0d596abd40489882279abf38933962072aaf6936640e20714196331915253e92c8b0827cb
z7751a3a4c6563783a7cc669abee44fab4e178ba0e0ec87fffe5f8f36769aa528668bc37aeb2072
z120f0cbf6dde0591b0e334392e6da44df36e7793244017c2b8c7b2585d3a8d3cf9f9ecaacfee1f
z65e0f131f4fa0e943a1543499cbaf5cf4b63749fdffdcd757b154eb9cd147e020583a3717e4e08
zb6ed41f7bf249bb21843904694939075655b0608c63dfd08d8a29ff1cb3b0f46d96cbb350b9872
zbf2dde0c225fa45f242e4becf4476649b54a78cda685c5ad86f5c5d1d9bff7550fb2e508ad8211
z7ab7e53540ef3a15a044672dd652f6d6c8ece1e7ace5cd49e73de7decf4442f9257d459b0085f8
z83bbe6d5f6f3edd894b57e97d44188653972c61df117c1245db4a22a39d25f210590d078ae28f8
z633952c85bc533201dc7e96c4e8b257580c2e6e50141eb926470091530ad0469e8bdc6f6daf9ca
z01218f849e1cdd8632ba031e7a27b80a793672d6a37798548fd79535d518231b6efc99de64e112
zf2325b5ef6a821abbb71d3a4639d677911f4381fbd73660a415120f4935c20e8134af24fd7c723
z3a341669186acbdfa50b066b650e10515edf29445eb172b500f3d2ccb88d323a28477334d5ad25
z0d3e63c306d01df2b67a07182602858736b5d2dae0d2a4c5d463eddf0607c3d52fbf97e15e7b47
z67b07a30ad33105c3e8c0964ef3c3243b7760f251ecaa768cbe4856eb856ddce46d0f43213439c
zacf5d803ae4004f6b04afb777ab5f063f70b80bb6f5e6cf8e8b0536dfd2138366c7c3dccf22be0
z0f147884d0b8def890cbafa609482aff6fbc2ebc40784b56701ca796d1848537af4b87f0dc65f1
zd2d74ea1b3a6e3ee87b92296b9836a1022c7bc196004c96adebfaf0f87ea0fb52af1a56e536ef7
z11f1dd01ea9e1b696c3c6186884697054a2e41208164895e9ffeb47e7e613368d17b74ca396e85
z1c7a095b336b22b097777c1c681f34d0ab22ebddc6b0da7447dd755d7c941e541b979fcbf91544
zef74c354750498fea2a61dad8d39041c91aa57cf30f2f883bb93ade04943eee32f942758678424
z6996c64f043faf459443d2c95d5a628ad37f9846ab230c6bd07c4c21561b71d883ac58c651ff5c
z4c1ef7b6d031da343c3e19e9801a98c98eb836cb807bbaaff743e7c2a6e31b24353b19075793f1
z4b44d53982beeb7882fd6aab888bcd92d7a93469ef9beabd07dda7c6d3bbd0f929f5cf97b88029
z57cb87634f33ceda3485c798b1eeb89294d74b103ef55c716e9a2c3bc05e86bc80086ef39a6233
zbdb0ee3ea839be2e7743c815d6308ec8cd1aca4e7c7f9c4dc567a092bb66a14a6072f7a9e76d3e
z37784a1c07bd06e9d34778de2676821a502057f646e0170e3d9933c963c5f67b4e632426c41b48
z7eac3a33a3593fcd4ed1ac70a060c839e3e7a2e1f5d71d64f7816a434a4e905898cd9e1542e9d4
z3f7cd9970ad77d68dce25381b4f22f649dffe6fced267d2408493b191df8e36d05a9384874c681
z4a4a0a7430d77f0e57fb1d40fb328082985803b27383405cee11e10c32763506434bdd88094711
z5b9a351b652a95d06b9f13737eb7995efe1075b9b06f89a7ae9367759c384a25a91280e439057c
zde5d1e72425f9eb4f967289520d1ad781a4d4058bbf25f74d1ab9640e7b59ef3eab0efa984bade
zefde8dc5cb9c003f79e8a266c8a7f11e5aae3e9e3126c3bd85e6ed92869b07c4ebce25f767581f
z1d9afd87b6f0bc5dff30f3b838abe836bfaa073a8f80d25bc00db4866bf7d6da72cc2aa55d47e4
z612a03a26d491b0f60d07b83616bb3a73701c69060cd3f6dd1da9e13b3c8d04a379038c64a4754
z8e284b1851692d4cdc5fb107d69854ee66d581117933987ee98b6960b56a2291a507e26e4a75d4
z4faa5cf3ad2e764093322999ae56a464f6df306c165df3967635c56a989f7f75308aecb8118536
zd43f0c32e95f88e6469b6add8baa944c496376e9d9ffa682de84d96f9fb98e649f4183d453c03f
zecdbb5b524eb07890c9f82e20fb37ec0fb731592c59cc52ef785f2573ad0dbb3c728a6d1ab9c3c
z48d83a5e48ed1434e13a1808470899f243e7b4f02e0d7a7a1248435f04ed89a2f2115e7dfdd824
z987e25ae525ba6cb45e861bc63e1034567c8f0c39f5f890488d33a48d8c95cf50aaa0f07d9bba2
z67597fb44001123bd73b9a7d4057d5b739d4880667f6a5f62a84d2d973c7ca953c6d4b64b12bb7
z1c6f6c73847fdc5b47a1eaadf009440e219fb3935334a3bf39809aa304474677049cd02748f68c
z2c7d218363eb007ce19181aeceeae874c9f8875154be9d89416fede2e94b74e932bae70f4e8abd
zc3c4789923919270132ac7493b86abb36044e2a512f41825e69de90be8f53c61d425c616e7f63d
z1d2c16ba481692729f9320a8541e7fb1d92303fdf83d8347003f73f1732fa718caed86930a9879
zb225015d124abd1574ec3f817f2f9598f7790ca47cf594ec594050e22f5841a85245aca9aaa058
z4c98577bdb28807ea0dc04ddc5f48953ad317d36747e8ef41127c7218a3723c91be1569f55a49a
z4d90f133a137e3327b2400f354ab54188228cd8e0823830494a345b81392bb94b07e5f0f0302f6
z63af26e8524d6f0476342d57ce9f1c195501f62a66ef576dbc07963ae36b452b90951ffa2c2703
z2ea11c2f31d1f0841d50c5ed00f2af10478af1017add4c13daf665735226ba2d64fe1e9f941b5a
zcd19a457fadfdd8a8e1e95fbe4d3690d2df7b99417e0987a0da4da3042af281698dff9afc9ff53
z485fbc1fd72e11ccba39875f147907a4a2232e55b29745a0ef65ab979ce4e53c9abec0dbd4f599
z2bcdf510e84da3529b6f5c3b953ec4a47589f8751c7700f0c3afc4f769f8dd494cdf953e44cf2e
zb27d80635a3ffc2f73323b8a589b2cd51874d3cf5d6df4b83a7c9a828a37ed631d61ab1aae5343
z6c79186f9f6c02b963c10baa9755325868bf2237dd7072e6321bbf835f3b8f39720ff1710996e1
zdef189d3774c93fc77717aa47f4c5bc3255119ca2fc1fc5a949ee63620baa6cf5652ea1832f131
ze8dd1014c5ed5e9afcb6d36b6aabfec5a5807642c81916554ea970636bb2fe6e865eac0edb5e23
zebb0786eae65d24b256cd7c2ed7111ca02be9a112fb929212adfd87b3b7d3a75ab5cd1b8100d64
z8011375f8e0ba4fa9c4944a1c4f6a93d0fb38bb9bd66a2b5f1fbb75056d89868cbcc19041d056a
z9765aa0f38f6529511d251438b2834fe6050d59280be942e9b7945bcfc71988202b2917f44e7ba
zf01785a0894bc6d1dedb30a71322cf219083ccaa67561e573000198f5a4c5738589d683fb29d9b
z9ee4713b9222a9481c99b5e3d86657582c17bf4b966ee3d94293dab5e8456ef38af468c8abe8b3
z13cdf3c302b2f64111f2b33a552c849f2e0d65a692b1e43537fcad4454190b915aa25f86d65e57
zea167650f7ccb45b79877cf30267da4121492806d383b9c535a8cd80f3b6c3850a7588e6a86c45
z4c35c46f70624d98e8e34ffe19ea8663db619745e0ac0104e2cbf390fe7cf7385609a48f98667e
z84497a20fb3e552893176c117bc8616a8087bdab251683de393737c96fb3e5df0ec71bbd5aa93a
zceec275235207e3ec10fd154234fc9fc71e8f6912eed3f93c240bfbc27d0d4db9f1fd6153d2a24
z2703858d3238f70b4b0b546532bea849686f872a706ebe7abfa8a1a23b0bafc99809164d58890b
zd6f4589afd4217a692e537ccec9caa102c917b4c8a3eb88d7f0c8928ba1aac4188e978fc09d47c
z9765cf24efe8836a90429fba3e3b9e3860596ab7c8c7c4de30f32c41cea8b232ea0e1b7678eab0
zd765740fa2c333b03d84a0f83dec6babf68cb7d8ba6ee364380431bad8171ed4f489c9151080f3
z228f3833c7a8b8bb27dcedb5ef2d157dc8c96bd5bfbf160dd9d9522f4bba70df90f7a6fdc9ecd3
z92566545b5714be3fbf8cc5325a0c9cdd04b5848b1cce91a181ae056242181665c0da1b57e141a
z78601a7cd819a616cae053820406100380007db6071bfbe44adc7ed80e03adc44db188594a6c47
z9f6ff286c3695c46e983484ca8ed93519ed377ce101e36c0373d4aca53b41d457d4e50820625bf
z7e91e2633a0f312cd612b37938028c52cd87b6541296c10db313d85923cf7ec326879d2effbb88
zcfa9b407202011de6accece4a508f1a53e008cb5f525be7970a6cef46f6dbcfbfaca90d7e4534a
z53812a7ace2de08a546c0f468cd3df4c6792105c981d042d96511b1a6893f1a5eace48f119a530
za684e69495ca9ee4f64198cf0462fae2e75f5427e766628d90f1a1a138f336e517ad051a0e5b5a
z6ad2fd81ec7fe1f0f9a047d674af23084d50ff3c370eadad7f2da2befa82baec0b6494446c9d51
zc42f3e79c8395a8c94a319efcc0d56ec286f78c619f75df55df9387cbb0474257c26a17a2fe164
zaae2f98ae10b7399e9bdff31f18a13a89720b05da6089797e5318a24283edb2e5153a6e5b55033
zc4182448f5c3244c69f4ccdb2aa6eebec61c8b108e116fa235bd9bb666535871389d2604e79855
z12321ca14c3f741bdeba03b396ae046d452a7c2a17b5a0cbba8d7d31c7ca04ab0a53a7b56d9b86
zd793dfb18ceba5b8076b1fc9f7b83179dc06f8bc546e874f5de879338e50a42c3a71c224f8475e
zf4c79e3c3db2ecbdbdea6d91427e924d32ab60c2d5018278a1477711521a8eb4696c3e4992f31d
z3bb43ee0c8b0d85ae9e7644fa385802e02c4f1b90be1c081f0e2121d20d5641413f508c40d5d6c
z13bce324c4404c62a9c5f695f782f740cdac7c94a842a1b119074935278ada59d73ae0aa4fa83c
ze8a7058417e63fd03fa3896422b65394bceec3081df8ef63c23ea5d33aeb38238da939f5796f3e
z041b5b467c1b894a9c7885c23d39a2ca8233d1c74ddd28ed7d9a97bbfc1960efd861c219f7e2f9
zddb64ed606cd54052539028a606faeb9de7aaa46f7b158a7e0f626686c7c86e121746e04153464
z377cd0fe485e14adcb282b333161c17fd52263cda7a2ec83b5c600405754dc69dde45102835de0
z3dde0f3b4cc3c7774beaf2b046885839e9c8820addc601c38a13e8d3f5fa8e0396111c0b37ea57
z4bdce705debef826660a3eb838ef79c236b53d07c7e250ad2270df156dffdc4d87a55e1ab45ca5
zbead4181756892e3857017721e1ca347df3bd060551573bed24de0e1201e10dfce42517112c0c7
z540a4b19766246f750db589adc74f3d4ef86a41d465da69994c00ac85a7d226f12d3114b58ec7b
z9945e2f459cdaf3737b92e24dc50eca56c87811017e9c2ac4a68bc1b32d3cc34509b464e7012bb
z299ae7516c37bc55e43cbbe9e10b120c79ba8745ff5ccb2dbfaae795db3d8dcdc242950c1098f2
zf16bfce18d846526bc4a1e4c75bde1bee8add1f5c6470f4b22cc81aa0bfb292fdc34730b79a437
z8674777ac38f89a4a15e9ab3ef097f99ed260e659f4eb5ce153211b4d9c628c7f31c3d8351a449
z0889d03db0ce564528eeac0774e0e3541681ec74440d4a3cf021e635bd786508d7a567614e2bcf
zed1dac1c0768e1f0b4437665df186a1fb33ba6782f8815a358e0672942fb4e186a29354fb03587
z3193c040d5c170b911d9b52b5da1bca7494c6ff6632efb013048991d92eace144867ecb037e2a5
z5ddff81db4ae0c5994a9498f2d04a39878719adc7714f37e213e97086cfa90d44c595c6b21a43d
za168729452949815dae7fa63b2e893ca7fad53622bcbb777cfd5b6c5eb78afda442e2efba8163c
z6ac56a39700725f254972c8fef528191c002f1a852f7d3142976ddd81647c4a5d406946c435edc
zff81adc976aa37fef342bd673dc52b0f0f343a173e8a8ab0249b518516910c7419960f620a6a46
zdb78333f65f2b38d68b3dbe735348d741cd43fd02e34d3c5362a8b3b1ac23427bd00577e38bb1a
z9c38dc1f828ee0b2f51f3f9eff0a509872c1179e46748cfc10f457cd8c0bb615f8577eccbd372b
z7c352a208cdbc262d7b344dfe284225aa0d7f9e01999660663d9c2a66bcca5a74cc8cd8fa90ca4
z23d4ff622cc59e8124697454c598e5cbd38963569f24e3e4bdbcd1a69c1e98f1a6e3fe06df1097
z4646f0970105e7fc2f7c9721f88838ac7af2fef81faaf45e15207e4486abaad752e62d48c56bc6
z545fdff4ede76e32166cbfc68d77faf7f3d41e9be13a8fd34b634406cf35bf0a7ddbdf59dc8756
z3eceb30d720a091c48124e85b4afbd0e75756a2780021d9942d4b24d9281de4fd336df7d114efb
za1ca1506f0b5e926ab8acba4b865c01518e89900dc7f6c25bee308f652c94a0e1f3cdb86a63303
za3d5e05bfc04914957b211f4234923dc8ee8e7c992b6ecc4a13fc2e36e90176f4a8a87b7392440
ze94111b6eebf8b61ca4c6d952d61f64b0da2045e6eb95e6a18798a4f6213f064a98062d5a2cc06
z2d5b95c5fe59c29492f13a640cb0cbe10792120ec410aecfa6ee3210ce6f2ea4cb23afe9729176
z72983aeddbef0f2365c581b7c6d79d358bf044c58199cfcc3bae90f440803e759040d1805c92fd
z5bda454fdd104042490691e4e690c25e08943950dbea044eb483085dbe29e093d7526da5bb75bc
zdec970fc49bd014d730e23918712b8e1f08051ca051f37e3296cbb281034fea81716b1a764b458
z677fdf2b0cea703d9690beeb9c751de4305133dc3eee5aa9159a4d54c6d713cc5b6871e6ba1f60
z2db59ecd4dec0d5b61ea23705507e0f9d768a302518000bc21dd7e8d28d10764af1d8a6dfde1ff
z0ce957c0aea8041a19e8b19a29165471ff77bb748f2bd2904351acb53771a09d17c22c7820bbaa
ze474f9c58fa756d3bfa55073b5aea3442cbd4781e8beeb60c619a10f25e1988e5898db9746fd87
z5d7450c4ffe3257aaefef63e3e12582963bf802fca1de1e06292333a73b24614da20f6530aadf1
zad2646ad5d51aec7fa8033b3d37b7084687d34a6d4e2a784fe18f48b94188736f84435351cc666
zc8637da1e59861e4e767e1b52a79cd22e1addf4dc4cc80869b7fba8b5f99ae5200a2529c59093d
z2cf4e8ad477e5121fcc2fa370efd7872dd5e068267d8e4ba6d185335912b8c907e3562150493f1
z97b760121030c15364937f98ff8aefd69f1efd3757249729951b0236fbe575ba3c16f7425073e7
ze9d16d266769ffa0859b6c48d540811e5a706b75613cc90a1f7075f96345935b51dade9955de8f
z51a6995392adf2bf2b1d7c22d2e540395c5f1e9f62baad7e5ffe056c5f1f4271c644f9dfd183fc
z73a14f1c5a268375d88c26157e44274a791118d749f8c8045727be78d2d8095f1b59db0594a787
z15ed37f1cd824876be9be3ca38fab490c9874cd95bf8d13aa1e09304789701967a16bfddd0bc4f
z105621c62493277e0d50e39e5c8ba5387b2897c5552e9d85865eca66e2aa5392d22401c399b90d
z311515977e2e9ffde435dd055c754ca49163c7212d0957dfa8dba7d529dd3aa6255c72b247e256
zc29a70976195a6b9c4fbd598d5b815a9310656e227fa165e89d892beb315d2df663f75a5957314
z6de56cad864e9143ed66cccbdcca81dd3ffcc4554e1515c3583fd06024fee0254cc48f60cd744d
zd3b4729d8d939f3e99dcae82d00d86f6e329281e790b54efc8400edc460adbb3c0dfac1a51d69d
z303e48a55431045984c91428f5f581c27f0111bb02b94e6cafc8c0a68ea44166391464c80a829d
zc8f0a26909265501259c9522659031ba763782bd7e953135257de5e4cb9200a6c9ea3a6f36a489
z415231dd1a3bcafe84f862030c09d2d48dfc2f026f6f0f0abbfea74b0431d9c7544388ca2a5a11
z09335fa6d7d2cb33c74b103b70627c1defc8eb837c67bc4ba223675fcf7295506451f202a07664
z951ede021a7229221faea75a8f2b4f122092d6f92f9bdfbaa7b5b05cfea46a6789c353c8b6025a
z2c700fb65683552595168fcf61a5cc04700d9469d164adbbb10dbf8048cb147a0dedf9033292b3
z1f55e1c15f09deb5ae400d02dc0959c3743f06e709257f7f2dbdfb234b911f39751ee70b4e0084
z5d466bacf362108608ae8ebd421a00a2a5e1a431e0cb421790efec7230598e51dcfe45051c53b3
z94e55fce6257e8bd13b17823afe10d7fc5d35c8b823d640022fbb5722c954c73bdf12f8c591fed
z8f69b2acfcc365773c6c0f2bcf18e5e590de596c48c66b4753013f4bcc70042ef4175c176873db
z1743213fbef109a82d949c563d158907886c1f98f896e6aef7f5715c53f3066fe5c6ff6ef83fe8
zf169c4f487c2c9d8ba64d78d2064a34649facffb8b5e667a4fa77e2119e9f36bdfb89d6cc66626
za98d00aa35fc02bcaf27af2b8c638b08addeb29a777740ab093d750e151a081e8ced7b7ef7d3ff
z40436d88e9f62127ebcb41aff5b63887a506c9c40d02209ea76165f619f5fbd8c4d9cf718153e7
z9d1c815788d0dc46f2676833232cb222ae673ddafc88b22c1ffbd770e76d0d06c6f50d55ce98c4
z36e8900ba13cc7a7284c2fb11a9d2b9f914ec9e4f8d48264c691ba573ef683555508fdc9f4c98b
z35a8741697b0e2f62c1f6e3fd26e389312c84430ce01a8d06143bebfc958c25eab70a0b49f6238
z3a81fa41b2baddf9b3e94c8862249faf553bfb0403bfa04a5c3ec78887739a29c2884dd64cd374
zd11dbde8873a8c07afb8a0cf0d271ea4575ad49efd29de414a3bff279dad8ee6fd65742d13c694
z8b52bc8a516b9dfa81bccef8b2611dd0cc16199f14f145c0d2545ffea390d128a3bf7c54b130a2
zffa1254b4b62a0c1b310eb0f50c57e9b9ae6518d10c610689cd21ef09ece41403d14ad16bf6ed2
z022f4c0ed71e8638be72b30d144dc09e3b230f40d12792fac13f67eefb1706f8abad4f3b328f64
zba1a637ce42bea0a38092ed4ec95852916ab6a58e59a7c8d0029582018586f2a9b5842ffc9c812
z6320eef9104cf04e20b2fcbc7d038c6a42f5002a0c5c1c315fef96a1abde1e84646decba8847dc
z67817c42c5f51cded8dca05c5b5f9c221c0403d19d5694fcd3ff85fda1271339bc8e0c8bbe7570
z0c6d60bffb7236770035faf75e923ec18ce5fcac4dee16bde144e6e414bfe2be4b1e7e77bb466d
za0cfd0397e005b450880a877ea4da874d40a30727c0e9799d9a44011156c9bc2d04dfae4c2973f
z5cf1fc75f1992d14e35e041d079821f79771d97866c48c85205838cb06fa36c606c37dbe8daf20
z194f8a9629c7104f9688c95e575191671390949cab55a165cbfa683b2ee17f577ec0f768ba52fd
zf10ece2481c14ab850d4688eaa305638603fcc6439bf18d89fb4a1c4ef539508d85d7130a7ffea
z9567425578e1b678dfa5d893b4caeb92db59837cb7960b66adb24c0654dca031e1e191d9819f40
zab4dd2f164f255127ec47bbe777bd73b75d51ead6815fe8d9aacc47eb4cddb36a68359418d323c
za89587aaaf0a4f0dbc25d278f4c26515ba9447a11f991426ddd348b87f0a1ace2ca0e812d3ab0d
z341daf9e26a57a19b4e5f2f445f9656d6712f9af5fbdbbff4057360130cabb61a3b52cb708e01d
z802e3f2407c5f8e5dabfdb27ad4723abc48aaef5eeddd52dcbbb94c423c4568b973fa21dca7e40
zf3a360fbfdee1f5d5081d65050061a2226b24ff5511066b2bd66eb4679c5be6d7d50e9c9d14c2a
z82b19d20b1452495879421a91e6f8e747f030d762909cc908a033d5c0a764567981af890c2d462
zb0afd40433d5d851547c1962567666b1ff72910e303abeb5d1b890009c8bb7fe4e3d50fefcad82
z8cec6b8dc231c0f8c3789441fefa0fe944e542a911ecd835177c0c9d6dffa6175f8fc490c12c52
z0d7a8ba93ca3475103e0dc0e8da66fbde17da4273e203babf0493208282690f89240114bdc186f
z1c51d677c2c07641e5e9e3fe1147e89bbd72e4c72480978633e1ccc71623db97d4df1a8d5eb91a
z202ebd8d9b960fb4e9b6a181d878a1ed932116c05c71012d1a3ab570f9b819dda6e0b02a16c36c
z9549c4ae324df64e1e04c93810c7cde836e70df0f710a5b6d3ccc0e79146b9e22c7e9e460e70bd
zd983f6edda38fb4370feaa177b8905dadea83c9caa50804bdfe199c7ead00071bca26797a89f74
z56f299ce0d94221c015c6750d6b8d40a85d64126ebb14394d356006c3ad86686142a86c8fd6263
z05b8b51c596d7c50c2c5391816c55d43d4e794b780ea7cdccf59b169d12996fd96da41ad52fc70
z964282e6ad340d5e3868b5c002637e36a196a88c31bd5bf7bc5bda93863b590e6937802a5c4d6e
z316a5c709165663bce0194ce7d2c6cf2683f536ba739c88d3d75767eef834b7d4001ee7e924afc
ze0f7741965dcac825c481af502f571d3f5f44b07f60d79980d922eb00c680ebe820d3bf93b1c83
z52ccde76a3e07760a5278ab6299ce5fc3c173248ad0f7492c89dd5bed918acb6a1c8d87fc5bcc1
z71c380fc02415c563719daf553b64efbf5ded1d50e5b3accd6583dd893fc890b525f4b0fa403d0
zde9227dddebf2bb8ea31489a59875b7897f5ea2a46bbaa060618536b95165f4505500d0184cb86
z97e26a7cab32b6c63675da5cfb3355b71f62a1d38e2d9b28259a69390671af554748e0065cab4a
z7407675dd993f3d15023a0a628d7ba636ed63ef896e43006d5331b185bdc227c54d73e2c0d3b42
zd678720200e57988a707edbaa2db5d4fcbe06b32a41dab2defdbdffb216e875e760a65fda22251
z689ef5290fd9c5872b719bb4c25c8e20654efde8c87f2560fd7707fd7571d284ef4e2c6c90fa50
z40940f0e95e54f99ad0917e767a6f93fd74d8c6fd9576cbf8bc5abc18a5491946689772e08a817
zbfb434174af5b3c8e8ef0a6469e6c9173bb00784c2d187d9ebb210148020bd57d8c6c706ae6b4b
zf8d5dbd5faf83ed8005679be904e4511f0591f1289243739c2bb1c304c23404cf4757051526d10
z9facda3ede966383e86b6199f7f1e34f0711fefb6d44ee5f5f94ca291cce4a1fe3e8fba6abb88c
z18f32d637791501d638f82efc0428fd6b695f66a000a12e76be00953f5983d8387727a2d356f19
z49f004fedb5ee0419d82e338005afb9f471581eda16c0fbf3cd830cf11417af4babc8693a7abd1
zfcff838f523f185a31aae218971e6d1d113461b810362ab349bb32eae1b891ad3fdccdc625b95b
zbdf96da6d02ada05389112ffc18e325aa5379c321120897b5479206e0dc949d4d61014b92f6e01
z739a503063921b0804aed491a70ea01abba4a2691c110e9f2fadc83eae1d280bfe5feb6dac3e55
ze2bd25318759283bebfcbd01be74eb9120891b05d6c4a63fe6ff71e86993412ab3c91abe588222
zd4d696ac99feb70fc1ccb84d2ea1ecc4130944341eea1d804ecda07677f98f0e6219d6111dc2b9
z72c4aafb1fb87104fa11ef24ff300f4daa85c68975c4696c56771c1483d94190c89df30cb0abc1
zc339cb33722e3e1a84c25d05db81d06c55908a295f0a886d14362b923fbca393876c8329887f92
z5e92f7963c5b1caa9dbbaee55c417138b386a353d4532f1325c147a66d7b269f05463d8c7aa7c3
zde49e15392670ae774144675986737b9ce72b19a04021ef5c6078a472eca90416bc59eaabd79bc
ze97a866998994113d7b812600ce450dd317c86f4c01fa729c46dd32dc2354d2d535005958ed2b0
z38f004bdf346b0f69e7e6ee7b87a427c0fa856fcca23e30ae1e27b2659ef7474591f4283698440
z3fb9ce93d8461b7f191386480086a4f8866e192b2df2665d19f775b5915578c1dfce4729c365be
z9d6dae5b9f4f0fd91ed64d4a16eac735ba9a443041d6ae92190a7dc5d026ea01dbd7cf3b827a9b
zd68f799b21ac69d38b905cff1b3b728b47613f9eaf1cca715a713ce6588aa1d2c5db06b7350c6a
zce483beba08ecebf290677c0391b4bb673d9f273b8e8d0f7b1ee9427e38906194f11b59f3a5bde
z35981f3f818a6327b836373bfe1fdbb3e545dff4a3f49ad4bf773388cda188a3c023795fbe0742
zb56e9b5dea8dc5a208c83adfdac9c4d9bebf36c6b6fdb5cacbfe1b552a3e22fcac3a969495ea50
z047d97ee5b8168e506e4afcdaf6141025ff87f0710161046ee36147f6f4320a9cefcab1008f12e
z5e608a39c23a65073c19c05247abe2151c855244bd3298f0a26f5bfb29e16c77ac02b65fd289e6
z8e84d0cc10cfcd7557f1acbe51e9c95e3f04c53d08473b7724235bb39f4458f93fe895a0ec76db
zea38b8b734639bb698d6b29863bb2fdf7a4a40be0f0c95a48ca76f36bcfb2d2cbd809b432370b3
zce2e7238de8f5f9f0e12b9056350b744c679f7d109d01ab079d72add414fe8369a60ed5f2e1b18
z5026212df8b2e7ee75178dfdd67179e477ca0d9677091a6c094371c261057bcbcc42f0f228a339
z1a41c5054b693957b684be87d99c33b00503f63daf24384c19a4e11f1f467d3aa1b8bddd9b81f7
z2d8b27fd091ebb478d963a11b2feb1895de25584a23912e71f89a81a4dd439b6c475fe441efa8e
z754e37ff1fc3c00161fa38ccfe67c1fd27c9bff0044310593a9185bfefa8ba7b4e751fc1c414c8
zde0def8ba07f9b59b4c363da4b9164596d917e01e403d122bf7fad5f4407c2c3f997d988104f9b
z2fbd1ab8d0c156ed7ec8ef48ff8e3787b1264a18b0faa2f2364ef66a3fc18e687ccdf561f0e77b
zd1ef0bcfc211137c9215b8e1f0b7fb95ca63b0ff32e2f45802216f7937d4c784cc3874149ec914
zfe545ac6f4aaf9b8a369b2bdd2cf38da1639c6f3f56ceae0cd503d9761e725e88d62594ccedb98
z2e0372c868f11d0f3846df2b2c412c302047ca442091281148ec16090c5a57b4019e129cb3db78
z2407d87230c4d9888ccd40372a8082f4819afa492f952f2deaeccf55300dfea8cddc3df9515531
z09b0ad5917d0f8979d538834b9bc6bc52f11512028ae3124f7ca9311da8f9f07f08643aa9bd364
z01dfeefedb1d1fa6b659cf8bb10bfcb5ee488a94b70b6b4025f578f069dc373a68e6ffa0aa869f
zffc5a72cc8bf32a1a711ad9e31e8c242bb7950348c15cdfec4c22e6733bca62c62e8f200ec8abf
zc5e3a9159febb5149e2db0e78340b3c9d67b388ca39696b84ab7fb57d943d70d656bcd8cb892bb
zb1f8bd99bcac19ac2b9471053a6d5913877861d609bab7243cc1788530cc8475078c1b51c31722
za6d9b1f923d469836f3f442ea8a64a2cfd1e0cafe198fe2f459cbc05dc02f4d81e5ccf2ffdcae8
z762362329e345fa78ca18e8750cc1824e633ed0bf8c0195799cd4239ab11ce77023f22cb523c26
z08cde09d6a0f1219d01f7e8dbd50c1e4857af6e79b9b82091ce6dbaa0f1ad572cd440715fe8f24
z21b227dee7d4de432761f8a56707c5d84c4b736a3a582eb6cd23e28962fe8a796be07993a971b2
zdd35f6380653c2de070756d08dabf3a8d483a6976b22b03408bfc040ab95970c5826002de8f995
z201c4be458e004548f5f87cbd76ecb43787ba28ab2e6a99dc596ce76b9b3625b17200e94159a74
z5e6c2667001cab6e62ecc104ef10794d58ead4f8e5007357a1186a96e13b081729d4f7f47c8030
z4fdeeeb7a1484718515b26452e394e6e568b8965516212607ebc7dc2127f536e71f36e5234484c
z78ba35c21e337ab57cc3543aabc5214ffdf287a9f773e36c7b0b88f2617d1d04cf1e407aac3a1d
z8655efd5c3dd63bd4676686b844bc8a19886fd6e1cb4596e9ef6b6ba5bde504203defa8b5db189
zb18335f09b0bd93a3035e102d9f6c251017d6689a5402da003fcdf935009190ad34fce0d23b8fe
z9d590cca56d50621bf8c365761bdcf0156561ebbae317d1f163ae805bad8d874ffa527a8de0c20
z4cd2c12041657b2ce20aba5024c0bd1a31b0a4359737c2eff25d641d9456070f4c46a2fc1c8a6d
zf9fd44961d8653ee1360258b16cd939c748bd161471c4da3815d86e81123f8f43ad3d454bb2e6c
zbcdc45e460a381f750c0a8074aa8324769f47202b45623516e75d8bfd218b6f368154280079749
z696c5d960c66a2d8d899b111d8643e164cf874a2bcab8af0499899f4e8c31faf112dac0c223ee4
z570b1e2880e5c4e22af71ef1861f221d8ca332c47cde59b9914db29901cf0b6c737fba3286b527
z03c392dd0c2eec274d7668b30963b9136d1b39721304c8d6c34c82b1b730b69f85afa29467d3cf
z9430d4400ec40bccedbdf5a216f6bdc13138a5501dae26d3977c626638a7a0eae7b7ba398df702
zacacc336a67a36211fa41316db0777cb4d7d309799967f42670301d9ca52fc40b93a8f4b34e7b5
z215240212201ab1d2cd0409024e59d5c7fbc38771c2f0e12c9fcdf7f4fbb669c7ae7ff439aa810
z7754708d5c4ea25a2a23740e9b72d686fa03e2c68db883b9133324fba66f19ca3044f3d579ea6e
z1d362db2687559fa85d0b0d7bc20f1996944c4d040a2561e2295b4ab5713103d2f8b7ce1b77828
zd34f89604d31bd8e5de6691bbab2a86dee80186aa9c01a6c78cd55f81c11bbc6906ad496358d4f
z5ed635238f11ad1a4beabaa9ca5a579b378d988d490525eaa4844d47f096de0f94ddc07ea5a785
z6638ef6f505e35c1d1cc89aef97d33351a0a683dffd8394967961e61dec61ac1580a612fa9bdb2
z1aba13c41c72f6d5e47e0a68816517cac874d2ed49c8cf2ab320245ac1c5b9d99eed93a4a98baf
z910f7f470a10d9ec36e6ee0b43e8710821b31a74962fd095881f26860fb28e2afe59d8bf6525ec
za134f2d43bfd73caf503788331f25a01519fb52c98f121195c5f6df3049e94547289f60bd89d6c
z9fdeb3d1ff00208eba29b8c616175b7305d082a07a9555cfe5aa1bca0b95a6fda017504f07fe6d
za79e8b866ddbf1990a39263847cf205132ed8e38bada199afef99da49c966f5eed13bd05dc754c
z67d182336067ecf08ec0d498b4020f07a552d4bd178d8dc449e00c25933d8161f16e95ee2a1a40
z3ae4e8cf2dfe9b859b8926b5a1aea56f09f075b07d1cc9ebcb58f3be93488f09d45a510267f939
zc030189f05455927c7464bec9778e536047e1213300206a6d8ad169bc566212266302c0c2d7909
z2fac9680c66592d0c97728400f171f16bde0e1d780d8ea06d9d288948d8ccc31f3c111f97f2e7b
z6e23c358a9cf3653cae4228c3cf4bd4809864d1d0c348906643514025218455da6129a4ee796d3
z322ede3375e23b01a128f63247fe31d6a04bc7004db5c95f6267736f13b92d8f41830e85568a6b
z8587a4f121c9ef8cbf309b54b859945ef6a85b7db5d9a05af90d058bc59b47785d976074942088
zdf1ddec00e94b4f2c94a54e96cee068cee36450ac61f1bb8697f8692b85d40b3d6ee0b86c75ed5
zcb85e87e09fcdd809956db66ef9d9d20b9aef0810f58e71d42f7d8edbf14e24433182ee0cb8477
z518ebed4effd313d45fb5f182e07b48aa327f8cc0220923518cad8aee25f20b6ee0b2f5e48ff33
zb8a905bca952d1b3abe7043e8e0f47b330a11193871a99f4db64b39bb1de8617581d99e7124ec2
z12b0cce7127c416bda8e548197317d926aa347bf1c553170730be1de6e702eac86328518895709
z2866d26fba8997418b297c4db70ed3dc8dd1900e4577d201aa2149ae0933b5d151560a3fcf4f06
z8eadffe5fb01c743d4e021588eddc8d612a5d07e7dd5d22a6523701f18bfa775cb05ff07e53fe3
z939d21ad5db51d6960054130dd13bf89280cb3ecac20add09fbd1ad95adbb700dc8c4f16c00539
z695b033f16baeb4e4358ee29afcc2f461aa17056e6bc960a840bf71a95b52ff1ff5278a4306e22
z3460902e91f7c8dfaadadd4da40751f894720ebca634206f0d88fd83d0ab6c8d4d64f78b62327d
z1c696019c7d4796027f1cba3954fc0f547b62bdc63aac0c6b0d037f9d6aa2dd1600b69b7e4cb7c
z72e978f321b12064d5fb1711b43a78d0b402f9cab8b19423c3d9d65d5d9699ff4699dbd981c143
ze649f8f3a81c961783ecd12b4968587b3b2234cde864b67e90cdc009eb2ea7ed430a773b85efd9
z9b99bc4b9d3e0cc83d1288466171220e627cca4fa5f421525b249ef9b78e37d8addb0c3289ae96
z01d44159367ca158bd50a045eda5ffad7f26e559a77ec8ba25fe00cc78e277d56240105a176d0e
za5515ab25feac0dd1ecbd875bba89a875fef8d760279e2afee098919ebb27b39bb0b415438e4fb
z33578258f51d38f7678820ddfcdcba2d00837e4d3a67a6a7a502f9873dd3d793155f9282d179d4
z727c91424c523152bb457ccd00cb726901a1f0132f00b21ab8a14a4a127b5abb58d181ede78bbf
z9ca5704b35a3e91fa918a6eb749fdebd420f04f71484f7672505a195f8ed55329a8fac5bf650a7
z41e37772e39024920c19abf522d74aef26ae9cc569ea24bd9bcf8942f7b8ba5c92342220a7e471
z1fc576553a8012c73b4b62ff7ee0760c13adae32b240d4721244bb2b4e1bf29074c5c1a440ed8b
z8c7a70c6772842c1e6c03464eaf714341390e44a7c3c6ec16014add89d9c96cd76bb476711c81d
z632d3223aa9458ce8f2c69c97e271aa08dccf86c5912ad31dfe6f52c33431bb4b805227662a8c7
z6557ecf212c55b7b528b8b9005fb85f25e86cb954e74e21b4ca72f0c515c5e9a1e568deeae7a74
zebda7b0e857768e309b36adfd0057281cde1bb18f2f165aa404d4a0177360187aad344830aded1
z4d41c5f7959de26679cad406790f2ea64f18c62b719e8ebdfce5787d8cf1754c2b5c9b387e304e
z177f6716054743b9c52e493b85151d72124b3ca86725d62370ff14211c3e11573a82d924ac6386
zcd174c363bf3b807401d49c4366cac06046d7e18af9ecfbd01933f58d30cbd7fb0d5be6026bb18
z3cf419fa6c0468d4b36e50b97163f56a3864ed5f5a91f9e77ecea43f8b65b1dedb31c35e280efb
za71a1951cbd1a7bde1ef485fa745c0611af9481b36a3bf5aa05acbeb3322b947c6eb2e3d780938
z1a4d42f1700491d7885967dc03e4a86db4bb63d63bba9fa4f0f5c7790e1f6bfea0e46f3ab6c1ae
z2e3c34dde466d06bd5508472b79104932408b2e36fb28b5c9a20c2a9b088aeb13413308082e3a8
zada61428ce866e4246d45c9c20b4a25b72844f5795e84b47e1966c021242f18e60e48ba2966ed7
z208b3871c895c612b874805867c97dfd325ff1156c72876e0e42fe8491e97119857de058880271
za9e5555f0d6335f4dff7f0303034ff164f6e4beead1d73f013f7a147f071d2e30de2552a46aeca
z3fd814d047fddbe039925ffca740de87e3ab13868c256593b377a4f586ee7fa2c482a28bfc3f5e
zc4fe7ec55dd85020354b2d0b136b9ead4502e8f1cb19848f1d5c2775e5968cc149344ee6962974
zb7279134053eb0da4de183b0f7c08332ca5acac4e8970d1b413e6d4c045a1ef594518a2f6abc07
zece790c67d082b25adce2705d0d411599e3985e2c3d6b72f630dfdfb456b777ef0690e9cc0539b
z04e8aef625fabfeb4c9a5bfa455c73fdefb2c5c2a97db2dbf2d5ca2929065f505a8340db8464e8
z44785168c8e39cce80869b006aa07c30f2fe8afe9501da4cbf448cef95bc648c2ad817860293ba
z4a5eb331008cbe7f769c0342dea5806c25ed062cae6e1b940f1aab9c0c76ebe15040c45f1ace81
z4dfe93811353e8d68c4fe9b41b8cfc039bd4fb878a352068b383efef3483dd8f6cdd5371dabe99
zedfc85a9140af9ad525b16244b5227671f38dc8db5c03f1906b7c89105a208c4e96c0862e6d2a9
z5114ccfbc781370262c995e8656161013a161f52d3f9bccdc13e01cd2a788a255829276bbc434e
z906922c76ba3652e10f5b7bf6f9deb72d4b68e2fcf36b12895e01202b778c3b92ea186512e3cf1
zf51d17aee9eeaaaa9be33b3d58351c257dc380cb8d1a1c7c2910e7e1a1a39ef7c9f6afa590fbd7
z919788d8fed9f7968f5cd4ab747fcd8a7fc610ea5b247a6b2ccaf8c9a75b3716e2931de28ff3d0
z9f60e7da9ca47fce9391c411b3b672b8657135bfdda3c354e98da4fd67f4c84f8c0f7ef983654b
z00d7cc831133632e60b32fad0f60f8e3bc5192da3c34f44d138e57dc024d89db2c8b3bc00987e1
z32b45f3c0d0930081f0e69e6094039f156e41eeec429840b788e214d58744b525c09939b009040
z0d535dd51f2a5ddabb970fb289a5088d5efaf7174b474b3057e9201edc919388cfdc0b7eb45d93
z7fa2cc15d455f18e21618a07171bb6aa8d78aac78101196c4567f6bb96e1fcc44f102e348f148b
z78fadd92b13e9c61802c93cecfad6026505a7114df443de089593d67b96b24415f6381394b7d21
z9af5b645442002606033b017f91e15a76e3b389a79dcb4bf3fe81b5fef9caf614eadfa0e13492c
zc8e991065a9ca02edbc971aca55236d2dd892eb0ef868717f6de3754a45db54d04808926479dc5
zd5265bb384b47d8d002b56e032daf8c53374c5d59fb2ef1fa730a70e42408a286ffe7725c3c66d
zbc5c368538eeaa373a3b3f710f63b503efeedc347c5153355a903f243e35790d5e15ed8000d6f4
za03c5940dbc32acf85098123a4b641e9240c1504e2ef3af96e7294ab9f9ba69d14bcbd1fa94c18
z8816c27eba5198d10c1ddef81c716a98e57564c28d09a23410622cd8b4a643702d21f5577bc47a
zbece81c8639078c936ed4cab3135c74151b93daac8150a8d5835685f2940ae49dc90540dfd9ea3
zef5f262e9ba05775c2ce93acddaca0d3622d25d93fc7a5991a9f338544cacd5c82911e73bc2ce0
zcbd42eb20ebec2dafc7147034bcde2a7f8b7ce746b9de6ea9c095322a17ae1c853d418bc796db4
zfb3432d07b328c3474d3aacf4807a0caaea023e456ef105b8236d6d16a2b106a2e237432962fcb
z70ed834acf650b34306117417a5c8242afddde7d2776f215fa4071b781aed07a054ac39920bf1b
zc53df9dd578c42d3be8e7d744a3aabfff8de605e5ac0557033e8598391e8f6b115559c2280400c
z489f999693cc703e2b61c53a1bb8b885579d8157ee71a3155c02a3f85efdb42151f936129c7de3
z95f64566176296b19cb9ae03962d3a22eec436f3401e07ab582b1a51d78d8e2cea6fca076ae73a
z26e9e6a51f47635cdfde1ce693ca9e3cbcb03c01873e4162a9e8446d942ee3b45fa4764f1903e3
z1c93aad73030a7e1c1224dd623e8d873ac5d996caf016ec43a60a9ac4d005836143a3bd567f17b
z2b18202eb561e93ab0c8369f29bbd724ea576722d8e45863d173c412fe168b732df63c3f16d17f
zfab865953b58365a18843d39cb8b41f5d7593ef3d4f44d73af55296b7e3b5d3ae038e5baeeb755
z302a1e6cbd4e67d80ae2ff49342a8b76f1a112ff33a1c21dc947531d0a9dcbfad2d13b84378bf7
z2fd6c79aa83391b01ea0763ebb5669e0300af6f4d8e1361df9f57df5cb1e2527b3674c256f8eca
z8b96a9fd27450502c699da518863904fe1ca634bfae0547077a7c377e61c6fc2e5590ee1503096
z0bceb34ed5e8d7e5b9616a4c8989dc107d6a4c50d0b0d1abc14bfc4f733cdb6eb5cbc892da0a86
z541300a3c897b3a8aec20a9eb367091e77bf1e116b20c04ae7ad25f766370ba0891491c5efadd4
z7e914a6fed188562851b73c626173a03e805f1c9ec0b33365a51a0fa774d50d880b79e93eef98b
z02d62676f13e988af606515423f5e428111955c65db4f0eb3f2db7e8562cb9a04c9536a52e1cc3
z226179b37bab3aef25f998a651a6d87a45039c0628c7693f85a78a962e483bd582091fefe245ee
z96f58f2b6c0e504c58ef5aa7ba256594e48ef9ed2a5c2938e2197338e3c01ca224296392710477
zf231c1bfbdaba867e6b2c5f651e86a3bddf89984d1e0a5ebfea41567ec86fde5beba41a8995810
z845fc4a9a2480c27e812cd707dad33d1610f6e9f8c4b680801196777e2b6b7de8a7c16b2748cdb
z1eb96a1d0f6ebcd4e379e9a26ce6d5d6b79b2b0a6e972b000c457b8039ecccfa8f37c5848b1b99
zb9a9c9b21faf24c02b53f9d1e8deb03052fe0092b8322fafde7533b696bb6a570fbc7e90fb93c4
zb2e7ac4611b688c17c0f4d36094b7578b1b128aa9d2ce1b245aa7c1c441f6aa343b3d281d786c0
z3e93ff295e3dc2f23e5cb489b934488d65d2fc083a4621be11cbe475fb465df241b21c1096f663
zb2be38dcdd98032d70a3d451bbbb459ed454bca848723641c1ea9eba09f5cfd7f3f557d1b95a52
z5f38e1f46addffc00e80f2f7c4c568e14a8646dca409f245eaa71a3fa3149a5575d183e4eb2088
z678c0c101046011ff5ee2994382d3df2ae0a250901de4b1fac1e5c2bd41ce2c8b55193cb56fc6a
z3ff2edb540c82b78d43b01d7d88c5666b3536fea97a5926515f7547fe6b98b948d67554984763d
z25f870b1fd2e4116f5f1e09da699d52cff199702a0d2bd4b97ebe307eb44e9722c09b840f9ee13
ze06163ec42f12c5745c65ad6ae3bef600148a55b8c228eba406e5378fc14a5d7cf2f3b57bdc509
ze01f5257ba6c208b21069733fd9a2afbd5646817f9aa81b96a4876db48a6c373423f7853528359
z1e8ac392c5d0f6955a97690646a1585559924da593414b608531ba9e0bc1a8ac44936a9a07d511
z6e76a3d5d08ba0219b91e219ac83e32ad760522dde913a0e12ca709bf4562327ea2ec6865be341
z8b1c696901b0f5ab33f5849cb5f6b38fd4278db7a42bd000c3efb5730a0e22c76b284c5d2834ac
zda6e6793fc37d1e2c57765b655c3a22722b63b9675f0e7cad5577c703f40ca756540b17d995bd1
z80dde24fc8a0df92b1f13cea3ca5a2c725858e0c2e09ba64cec486e860d271630269b0a3281b3d
z5c7145c0cda70b613ff5733b328ae3084eaf896db2beb937d132e6f8a8b91603cedbe9b9ca09c1
z31a1790f1132f4d1ed4d94e33a49310c2b3a33b22e6af9ea830b345d17c3c11bb17b69aa0582f5
zaa97496fa826aea806cbe1a90fd811645d854a0661cb90860b8bcfa69665fdfe5048cfe3234872
z544cae8b20b625daee076dc70873d73bfa2b3b0827eb4ba93368b187b9b604c7158d73eb4d57b9
z6f2840e55b7b1c73f8ee16b1ade42432b9f47abfb8ce80e1f7a1f73b4f8bd8836403dae3faf71a
zf38b8df58340320ce027a46687eb7ef0bd7531c72e9852ba5648ac5d435009b0386207e6def777
z0a76831bae8c8324caeba643ad3dc7648df6095bed5953186dc78694da7214d7a5c919b03c794a
zfff066d8e013d7ceee5f74070b6cd2e46439e60871348519fb9fdc43b2e917b7eb4b6849875bf7
zc96f61dafa0bceb785fc3fce909d860150aca017d8e407d6a9f045022977d739ce5055f8aa5039
zd3867858b2015e6aa17437836bd0e9f1e010797332b97ed29782bfafd3b159113184596eb31596
z0ee6274775ea3c6b3eb9c1fd2ee589b7645ab75f300d02b3dedbc834586779f974d515c96fe05b
z17256af6662696a52be0588619402da00df3573d07acf2b548d72b1454ac81e014f56f1428f020
z99f72dde7d4f51de51585f97c4d897fdd8c40d788c82937c4fa66da884ba73058311a4523e0b27
za6f664b6b4ab453b49cac7cc20727a5fc0f9b94d3b61f27b2ef3c435b8595b1c08db6b5064d0be
zdb7ce0b4941b5871a9d489344a39514ff5cd5950b385ed2e9d057ea61a1005904853f7feba9c62
z91232b1b3c4c22cb7832bb507b7a5affa984a78bca8e179e978216fa31f55c0515a9af895d36c8
z6fb0acdb054830f82296c56bbfd730b5defad1e260f93dc712f068a09f9bd67bf969a0f35e26d5
za6896c06305cfbb15538257c1711033e4ac9aa455cc8272adcf79e29a1510f3b20fe100944df70
z6f9493c40ae11803510ce3c83ae024760a9e6fbb406f0ec195f31dee8892a865e635ba782edffe
z88972e9ba7df71327386d3cded8b5357acbf3c302025df29e92dbe727ada591b7fcb77265dac78
zafac3710128359f2d259ff2227dc467b43923ab1b58759c83c4bdbc8d57e6685c55144018ff7d6
z17979b6fc777a860350fa7535d08cbf6c20c0957fc716bcc1d962a30ed94189f305b65f9079ef4
z54cc8c4397c48d1aa92df857bb48cef34a0f6d29bbae76d38609ee50c17488d1808ed259c609de
z71a638125aec320cc6f2537dfa5b76a0ac9017f68d536e642102a072ce50725d9d25fd01f1436a
z0a45a1562b2933893c14caffe3dfe63979d02d59dfa7e09537d28d0a9a3370378c34712df89163
z8e14e6f81cac6b29df296d4ef6d1e23ac5885bf3dcf389421d4ee43453411f13d3cb5b98459017
zcd2bebd47af4ecdd9e1cebddb9f88253c7061a0eaeebb89f847e3ac5851bfd88c7032c79566680
z5000ab61fa8d0aa0d7dbd047352cdfd37cc7e3282d020e1f917878596f85d35794bd05daa8a907
z819b545ca66b40cd5f3adcc8dd5d051d1f1e598aa447c21b2b2b19e623411741f0c2369cd85ec9
z0aafb0d885b6e458e6a5e2568f1b29ea7e42f5d00962c58fcbbf9cbff0c08b837a8917c0d07e98
z52401acfa3208639cbd7d4c21991eed0a1a79ba43c223356277e86009dd5e912635dd8311b9fe5
zc30c1e8c3c88f961d05ce151e65a65f39f6cd88bc0e5acf07032217cefd1e89f03108a3573caa7
z1cfb0f8ac5f0b695126438ecc93868f78e7d5c0fe132347975996ec248dec101b4d1a6329b0b56
zbe51a4a15156906e6c87a3e769f1554b66a8485888339427ac3c15e0ac1ffe18b0190072605107
z3f406d0a07fa13664f82be38e66dcf08dcb293e00571c159f085bbafe48f65e6e66f19809e938b
z1743b6f90a80f26d038725c85f9242995aa9064eb73856502f74d6397f13cc7bb1069411d68e39
zca55a3f452a7cf2e28c9693931d76c6034a11dc9ab2ca6e79751f827a38a353c49e5def190e148
zf2cc5039e17ceeec541cccb61d9db759d9c22ba058c649d2fee4ca9511f457bf06cfc19f619492
z35f296e3c14f7ca832ca843cfb64878d88926fa0b061d8485874366545f665eb54d74a59e3e244
z2cefc28b3a4a1dbc311cfae8ce51878fb62a67e8eed9b1ed2597706b18dfc92c41c3e9194ce45c
zd78a1e371adc51933a3e2d13fd45b98fc3c1786ceea4c4e5d429a0d9bdfd16e013102c75ddad99
zd349d8d0bc2fc6a22204c30d6ed6ed732d97c982f8294a04465ccae1ac88861ba1e14850aaecab
z7534eba27a0611f32fcc6c8d5a5be449bcd7a449f6b3e300c480aeeef25028b803c894f752c53f
z3f0eaaae8ed8bc14ca1efe4817cf4368cfd66ea1e839b2476dcc0184964873516856c91dc6db86
z75cc7412ccde0d107bef0674affd891431e96a92d517704e68d6ce55930c8e53cc2c5ad845c91d
zb6976d30364b07cc8fab1256bbf7f7add78d0dc0933ef81fa1e2fa428d278746ac52c8f2489064
z89fb001e563b7db0a27314c3df220900135faaf2780c61357f2eef0c4529b526b34ac03278a756
z8a0ea16c61fd893277c0cd00ee1a3cb76626366c66498787bcdc799246dd7bd7cb6dfa4ae9325e
z6e7df31f6cf366963127f013afff67f1fd30d8a899c7401c8c347a2d2fb9dee1dd7e562cd71bc6
zea92410c1640694755d42a6b964444b18ab9401c1d23966721cba9801065e715b7058acc3130c8
z77b1ea760faa52ccb3df3cf2302999d24fc8dfc73b408036ea41aef076b29166e82008171edc33
z109f2d4e742a78fbf7c2d33fbe0121e23a9d795221fbb76b97acf1e9eaca84849519f196d45dca
zfb973d0ec3f11114c0d16fc84e741cdbdcb3d25201724ee0f00de70cbddb3c7f5c17919fd7896a
z55f94841f01d0ed18a7a59f4f36d9bb4bfa65b2b9e8f3900e81764b17d6fc58a8f788a859836c9
z058b44a7b3054a7d5b279e5278b3442c1c7172ff963b24ee402ca239f1d9bf85abe790638b52d5
z8c8a4a894fd72f16cb5dd2154ddb350519506a5ba1f21c58c24da6f65a58054fa1e85e9ab8a43d
zcd737d4cbc378fa3b20f1d724384e841374dc3a4132723204d27a02bbb731dd6d0a93b11aa0206
z83f0126ef05a71f88d3bfccea9a424dc232f1eefb4a6778991476e1005b3af01fdaaa079f8aa9b
z8d97d035b2db89b491e5ee5e02696d322392f462932f2f56059d4524a89fc23f05ca93a1f444b2
z973e2f6b71fba8d39e97dfb1fe0afb46cb7158fdd128d8e3a58fc3c0ff9fc5f08c688877b43778
zcd7166e2d4d13f218dc5e02843da16c8d31859cdaa1efce60ac7a8142fbcb1a407dbdf8b90ff55
z36e1679728de298ab6e0826db9a141d6eff850b0fe34e15ced4dfd67da790df98944585d553d4d
zbe8ca620053ed592cedf1b200a053b0bfaa6577b8fd5ca93019c30a130a9c06041d1ce99e1bf4a
z0163c754bf8595ba54f4670cf3f0509e4325ffcedeb955a136055e23d23cb4e46ffac9e3db8cc7
z02da03a6ea6d2aa7c89206422dbdc2f33be39675ea51350887e623154afd9f936bf2735af13361
zf69d4072080687afa6b58acebd0b97e877de46e387ceb4c65a8b34d72ce2627a58bac0399b6b2a
z9dcdedd9012e0ee90c06d2d126c9db8afdf1b2dd0aeab7970889662f31e837408ac246a3538c3b
ze5d6bea99f4b12fac56763ff8809fb4fab0d7939d26ff3c17dc78cac7b327dd4eb082093270714
ze182f32fdddae08627faef6ee9de2e13aaeaf27c6198ed689d11f849cbd91d897decd823dd72a7
zb26ffce330d412347aca1e591bedf68fa6b4e51423e8c947c2ddf4be73868fce48515a810ac687
z7b9dab0a5a60d7dee3e17e653d9e684c1694c325b3b5277a09eb9bd91fcecdb2e617c6b29913ac
zd50af70f6da989e54e59446d5514c4b99c1856d08bf7abc94e4b6ec798171c2eeef3f8d26b67ea
zdd83b9c436ef8ced03293c39ef1e7829d131b4bd26829c28afd4c07aa030eaa3fc18c5fbda0441
ze4b982e16cdc7a34cddb15bd040592fe7373781330afa61395d6f6bfaa72a131aa066bf851f163
z53a33026d6c5301c23179ee620979839f800dcc324aa0073378bdacc55eda4684e4a956f9689bf
zc06a7e8bfab523d559738b9a6b9256d3d73a243ed5eddf82096e72eb5b7c24bfd746ffe2c482c6
z089d1707ed83a904a8d65a0c6036283895c326a4f2ee76470e1a225b22dca54ddbe51b32291689
z350ad0ed3680d7fd59f38a4853f454b506ce5efcd291d22f6db3a2229e8b235268caa3ea68318a
z111487ea2e2fabd48f492f2adaf4b0f7232527619232c27652eb99067dceaa2b7bb3f991ffac27
z9218c6aa3a9810000b608f9975723a37ca0fa1a5573efbe1195e6003db2908028670a52c76bdce
z8e09eca1926492eac6c78f6d290943a3150def2c5a5a399cbeaf0bb7197a8652cadefa5d6dc037
zac30f2f9bda5beab381f3a108dc73ecf1f47ce62b723e0c24eeb648e03ffce355410f2b4449174
z2c9f2158d853fa625a32b9c1db65616f9c6a0f2d1ed3eed930634323c6f85e94648ac65738f8f7
z27772b59185a781d3dc53477c3b39c519b7c686229bbe4a5dd142e6605de0721399942d195a80e
z0acc59c2672312f52eb97672cd630bc7a02ee0f79881969ae59333d9b1901ca4e5d9f9362532e6
zdfbb24101ca5429010038d6c42d82382fc6825adfdcadd693731f9a0be154841950743189dc3e2
z24a35c567618a4e21542bc1be4898cdbecbc6fc0902c86352e695794254803ae3f58dfb5ac1f23
z3e47c96d814695916db2e2e0b9217d70dec381af107427744625e19ae7ee822c253974a1c80341
ze143cc153c0a10715da1bea1e8870526544478b6eaad219ce02fce6a5f753fb48f6b4b97b10d2e
z356a3b1f92f7f81c86c25dbc8ff08f4284be819391d0a279b49f7a318a24f076c4fa3418c93326
z87356eb24d24a0d1d501d61196721f48a1338ca9863697d633410adb68e528209a628c50cb4f72
zafb1feb7dde5a4d174f54642bd0ce46cccaa122b33220fa7bcd2aed96a8edbc77ab7a920136d24
zf06e49bcaa2cb35b7374dc22fd44b3effec615430a8377deb162b74d7b5880bcea3579a0db48ba
zd020015ffd841bf748e255f44e20262b2dcce953814017937d16c7a4e09ca19a2e489ae446d391
z8800e4440a593fbac2cd02568bde283c092f036cbf857a5c6528a98e5f94236a3865dcf5df5674
zcf85e95ce167a5885288501b259ccc7919a258380f5fd72ad5d42055c5916839d6a202b0d653d0
z6ba9e9ace143499a0d25b5b0b85448952b797e4110e918ae534dada96798c7877cb05cc193d5b7
zc5f4354886862959a05090176478c42594c1829c462fab8fdadc63aab24d96bb4fbac6ae276a33
z13cd667b9a21bbf9e3a532085ebc8630d46f097fae88172b536e5b0f8e4fcb630aec35e3862ee8
z1a17c9bc0abd0353cfaf277f8bb924daf0a905d3981a6d01a53be696503182137a18c076d821ef
z9dd91715eeefd3ce74e037f5c97696c775383151337fb2bbf73b567176d8a6f55818af1556fc9c
zb562d6e9803e547688765f15c620ed8e5b7062b68402f2cfcc56e48461454d4c28bea469ef4159
zd994097981d556ea2593d9515cb5684309c1ece3bd70df75f50f4d66cf76939501615f7d9337fa
ze087c157a72f5c2be08e5199b8dc034ee61812591a57a4a9f527a624b21edb206d7d81ee0c60f9
z32c28fa6392039db062d7a68aaa53306f92a08362ef3d612475c1928e7a48010ab9c5a98e4739e
zb8ad3215606574586375dff02f3dba3f39e7b6f730123503de052d6479ecf77d19ce5170f06665
zfbf94e61ed5b3e1aca8130bd3bae8c5a8ea89f41656d720b4021ca54a6d8de78c091438f8b3f90
z257da9f5c8f84198a774a4112f9b97b46d490075acbaf0b4744132453558dcfcb72a6be66dbe0a
zbb5b03ead6b8a849344825279f11b6b205c9bee8a62e663bf9c49bdc1a8fb287ccbccf29119289
z793a383d92690ee45fe195748730b684161ca0dad18679dc902cc8f2d10370e37cdb3cf2a78982
ze97b89284cb4a2c6fab6390595ecd5f2c5f19a27976d0a07508dc4a262a6e3896236313ef023ad
z8cac84c3cb3e12e08272d9a39021fa08140ce29566b574ead1c240b1c697766175bdafa8cbeee5
z69c4e5cd2a8f5b86d7f2add45de82d58632bb4b85c7d769422ff931858a4f387c395b4911630ab
z4a90a5956a1c890e68766a65c222c436a81979855e2083f6f1d762d351f1172b9ba146b438b191
z5a9069bc7ce71eca364becfef60df537756f1e70f41e2319ac4656d93d61252f667af44ec3eed4
zb8aa81145957c27306247373b6fd46bc279c5f62907af8d9a303af7471976b6d46aba7ba7c25ac
zac6472f369d2cffb67ef6852c14b3540340feab6855d25b1a56e8a57e8369c8b747fd2718f44fe
z230b72792ab32b911cc32328166a77118b3c4a309565d2ba3bc1f4d2e384b92a8c37ea2cbf3c97
zdf5866dd27c80ac4b74568c1e445a986c1b8e307ea4d779290f6c43d99448b0296c77fd7303c66
z0afb86f866237a785d1b16fbad4a2e335deac723d74938e74ae2db92b48b2e60a6f45d861afe85
zed0f581db0df4678fdd29f0d4e74bcfd948954f01bf904adcfce8491dfc4340a4a8fe5f6ab1a84
z34e9016b7820cbda4b7b34a224110789b62910c8ad0d6d577534cd51013ea84efca9194d489b0a
zb316569dc16a3e9f6928d8325acc28398cce68893b4ae69d5b7ad42c0b67549c7210b501c24a38
z547d88cb5ed352cc21fcdc78f6181fb18eb6ff51eccee2fc326bc453d7895f1dd4014fd57a9952
z67eaa036ea53f8c20a81719c71abf6942c3f48c6f806853d0da7f4e8850c4f18e8ca9dc9fefb20
z9ff6b92e307482a156fc00d64ff3dddd310706cef1532c4b5aef50e9286ce9d0d71f8e978539a0
z5b9121219b38934450dca43b1d5a883bc2ea525617df4d8e28ea9c053968ba9ca40c8a9b922f04
z0362c85b1f2236c42f6b71ead2ebeaaee9e38048f438873aed8fec95d70712cad4ac46d0fd5279
zaaa66f101b0ee871e8f9bbc6f03e6ee2c529771ef72ace96d6198630b7c5f0cb95ae980bc298e0
zbd8ba08ac22ff9606823f75b90e82f7984ad337d6fea2d952a7a718010d42cde5e12719ae207ca
z49efd32dfb3d45415665b060c14cfe8c4634123f1d76ad037a285628078d2d717734a416dee05e
z765e63156d157ff8484e738f811500aa4a78dd364d28c7ddea05bf6c90df0d5386f463aa2186e4
z8df169f7c31fa492faa4a8d6308635b90e7aa12d70a838e758f51d7512b880a7e1273860873410
z75f657553157f758acac088917b22b8009d9d1dd27f3eef63b8abc2c50cc8ceff776b595c2b9b2
za24aa87c236b747ea2fa55713e6c6b3dfb0fa746c70a78e2ba6415caddd1086c9d72e62b43bb16
z27a3b2ce78a65e74b92ac186e89fd6e2546b5ce6b952319d8b0c4c8775c7799138318f902cd7ff
z503aa8728d45ea4a16a98ccfc3102997b0b03803b3577b52023ab84d1e8270fdde58f5828ca7a5
z374037c6b97868b1bf9578bb1a610c605ecf73dedb2152ef37d0d05a3fd207f3f891a105385768
zaaf9af76da317461c9bb03cafe82e5b74a133e4a234a235654a639ce3e0322c9bf83f9ec16d25f
zc75862f8fe256b2b1790d2a7ddd1031a54441cffaa512542863c2d3ea32c76e19ec56c0d87208f
z0ed8b5fb15792d30e3d4c60a11fe43db62741534909cb0437fbd2f9009dfdaa71bb0bff700b1bf
zbde02ecbff786a685fd1a17a39e31c6fa1b8dfa7ec032642c1a57b8c3652b13c6f850157baac21
ze833371e980f7c8689f049e5f729838e61d3ad1f5bee5337ac8348857abf21ce1074c63c837dd0
zc585fb506947d366417d917c17a0cf3124687b74681817cf7c968a3be746a221aff3564aaa1f77
ze0a422e5f757d2e8579d3431d7bfbdb0d8bbce4d2d8d5a1d1e48b1c996a175cd2895e50d064f63
z4c13bc0e71893fb29e4a928edef5c925d3210ae40bd987a02fec4d859a34317c96537d33542497
z143fed83959e124c37fb587dc17efbc5cea65ca9fad044f670a152f0435c28c01aa13965bbd701
z5e747d335be45b395fb5b62f1e55667539217293954b40958c687ebb65ac89f1e5e3984e23af30
zb38a1ef36039cc2ccca677670a8d6ba696ead51b9f93662cd717dd91b0158985f819fe66e84aa4
z64dd6fb720b237830804478a02aeac87cce8a7dd1d22408504ddcc4e8e1d9f181992c018dcf54c
z8c771a267efde6bc0c476e2bc4da94f9658b455c4f4560a2b4c765ac4c7ddc6a7d147114cb1f71
zfd126427f581aa8aafe9a7ace229229838e3a5c4520a6711a3d7d634717b5831bb27656555b29b
z5758159f6be9b17c65f52917153a385ceda4b5ac51c3773b1e5ca4b841c1d3ac10fe486ca9af1c
z41ceacdd99ddfa602f82fb65e350067e0090a0db28cd57b8706bfb2211536d61691225fc0ac9fb
z89674c7a5b46576946e1740f55a0288b0c61654b1bddf536d9ec23c4ab34bb293f1f51ea16a465
z9c0dd1d548c18106caff3be4a61421a8b61e536ae923f020ab26de0ab3fc0f119f59713f92c692
z8c6e429dae4f0de11077e6590fee05ad251b814a2b35a3da5c87c57c0427b5d2fac7ab3a7438bb
z162e4fbdd238bac6da8bd3e0b064a77730ec41a167bff8b93b2b290017a51e912ea9ad35bd0359
zab0ca13e3878855216e79e14a521603df5bde3a2dafac58f3f57aa879df010d996ddbddfc85763
ze946cc205fa66536789309d890c31e41407d5f04168579fd7ce83410cc30d529903b10503202dd
z40cc603c0d7ce6bb9644391672fb4d6671c6b9356a3226c2a508170965ec1d324d8e6f56a988b0
zdd6b399779a0677896ded9c8d72d72d183d599dce8baebbae96817882fdd3ac177bdc03d451776
z947fb4795f9c6fc19bb356a0593d392c56375d1ae21e6d3a1b0dcc34b6a095e30b6dd6670e2835
z4a8af72e3a41b76824e8b4aae58c3312cfc3953b1828d228c6546df9949bee8746de89fda1a5c2
z8c21e62bd27fd00455da2516cba814869b4d3a0fede93e3e837250ba1969354637b1fdb17d2c68
zb330f114757ea326cd365bf06f7efe1b0e09b47fd3e757189bb444688b869f29b2a20631258c1a
z6d1aed0fbdf35c2aa6f44e8d9c8828671656c9996966ddc4699041e19e0af6fe8c43ea4cbad9ad
z2c29118c80c90b0e290390d0c9c3581becfc17704fbc1aef41ef2141d63c6d4643c529b3212d80
z1f3509a764acd42b549c4f6b18ee3363f37375b477169fcfdfd2eb8c17805b848f855c6ea746fb
z33bbb324ada8ceec77d4deeaf0a77c2b4e28c0f932c0c89688adb7d51cc3cb029f8d2c1a392647
z88e8b0071708bf6b4a1acced175f6c2fe20b29c87279d8f9653d70eb07fe11ddccce89b4f4dd5e
za5b556f4d654ace1cebbdcecf8e828b0916edf2468b72a29356862fa7c60ed0bf98c6b795f78bc
z8441edeff2fea4585e35be21db2c40804629f1ece74a97c62ee1b86f38676d7bf9a1680d7fe3d9
z70093bec7460cf3af7dbb2791a847e5667dd706e3acf5bcb4b6ff79c868acd3ab065032bb8668c
z679b0c47351504bf6ebc63c56247d07cac9f4b6c8373fc8d5f9d897880e47d9701f0b24f0032af
z3246b1dc044f59c3b694eaf3925d71478bb9abdbc2ef46df644e8b475fdf81b7c8cbce8aac2697
z6112b5795a5daefd514981f18faf106a8c8d12bcef3c92155a7ab02fcc0c195024ed4d522a9cd7
z1e876fe71bc636b9c876d5169b254a0ac14a10093a4dcc004166227d6aa7d3994c597ecfcfe8d0
z165b76eb844649b3fd7218960fbb4cfe8a40b320971e1281a00f78a5ec0ec6dbebb9eddd32ea5d
z2ab6e29c8935395eafb8aa7eb43d0a048556224471925decb535e918d2ef8e41aae287464e0e6a
zb2db54dff70bbe55d8638d4cbbbdd901148b630e82b3170b6f82329b254e19dbb9efe3ce30e66f
zb34ca5aea6b768951a2ad208db143b0d3567c65c7aab107c38ab399352aa0dfec098df97f7664f
zb6354634414c4b8ca4e98e914fcfa410a502cf652a430aeed0257247948057619f269ffb4a70cf
z589d54cb3af7c0a04ec02ce44da3af834eb5cf9a8ae37e7b469ba13eb0ae425621e32a03573d2f
zecf1aa0e72f759489665a1a971a62b4c0fc6271c7265ccb8394622830644eb124f1b95e065c66a
z9c37b7782e08fab09f8b6b9810992f955f8ba808eb6d7bb26f1d702638207dc56b790eac221a9b
z7187f16909773e121e58dc1026274b1b04ace07382f8bf6187335824089543af14e4fe7a7b053c
z2bc4936070e72b0f6d0ffb29eb5927537619756a7c745b17eb9b7cfabad9d1d4a25cd1235f4a5f
z83d8ed1d8232080b48104d194623869196ecf7fd2ae0f41a3e8ffd922cde930e5bfb7b7d5c5256
z14118aaf25f166edcdc4d980706c702070059d553e3cd564d8f870b54a2f6948ba23f5f67334d3
zdb5befd88cd65f345f710801ea14eeb9e577a0e3765555a4b52f25bb30e7904cd45700f2c1440d
z6ee87506072e5d6719e0024f4214296c264ea6917fa8978c03298535ce0cb4f499b9c6d93672b7
zd197d8d476dde1f02d4d985757c54445ad1d9611e18ec585c73edc10eaff7652d6e422bb7b0010
ze6129276621be9454eeeb7e6179631bb5c7b06797a02d1ab1e3f33c442e1962c6ed21451b6d7b8
z4e81006581472565b0b01d7c7b10955059ec0e4270b18e4d55e66d0d56eecf10962a146caf6358
z57f08e382b452e4714113aa25a96a29d8b41636e08ab806cd93af9a0f9f41bb44c7d28fa604410
z80984c2901daa3f88705fe5df7cb12d210d6c55c53149efaea5d7ea9cfb7603062b9a24f31d66b
z83772d65b7faa211158fd843a2d4abe63fade36e00ee7456e3513fd6a31c0a2de418affb6f5205
zb109b1719641461a554ec45521c7dd92ef55a519cc316a5e264f86b0e848ab397f4624cf937c12
zca696036bf5bdc19c609ffd000691d1f3f6332a9d65278e71a8faae130f72f5a3978f0037cc0fa
z35bf1cbb1ac805935cc4880f1e55c7d629649c9ca484ce0797eefa1667511482b34c06e14cc259
z77e0344f695a0bf23a33cde0ad8201d9703fee245978b74cad3e18ed5fe520d98f57df98518839
z9349570aecf43db1984ce3b35c899cb486abf685497f8b377736b894f3d57eb48ef90ff3cd7f40
zcf2e3c050a00c0c10a7bd06d17a4894ec99a15c3573fc4140657c0eb17b89d05831436f68d3341
zbea1e552bf97759c991af7db45516329783da094a42555df781e4ac9e48554720b8721a03cb051
z57cbcc3f7bedec878db1d786b9f925333bbf3ebf8a35667bb2c9055207ca8d221f7b6b776c7778
zb3ed6db7ab0ecdcc596919a6e23ea240b508a89390cb48ebff768a6721faf4e3a012be9aa8e5b4
z370714313214c9be1e2da0d91c157bcd1be47e8f67edaa94db34a6adffc53e7f1024c7a3f650a3
z5801c3e2785fa7cdc6d15a04f3560ed2c9e13c497b8935bddfe16670a90058cbc4ed8ea5ebbfd1
z33499f3d2d04291f1352429e558d8e8f8c713ee505227d3f98521843c34615546560e8bb158d48
z537ecb94e4419351c2b0b8d2920c3820594263750128ffa6e90dc667ec04d32d853df7d68d7e60
z79454670cf1cb9fe6de1c31c06cdaa40dfced860c94a7faa0fbd3e3f5fbd477178395aced0e139
z5b81f38ddbf765141a86d02fe3d99bbbdf02bb5b24c503afb38c86673f8bb4edc40bcd59d96583
z05deda72d1de187246fead1b80caf4c4527af5ce59f208c742becc27e11f5e491f2680d26062a3
zd1c472b146c1d6d12b3b742526bc1a2c8ee12298ea64b51356460ef5b5ed85518afd4d1445622b
z09c6435e6530c767be838e37f002d5421734f96a32bde3463ac4842dbecb684a264ed2bd54bfb3
z310c25ec5d131d5a8c044b6b4b1cc933be70b366de4b5f2776f0f5f65c9ea73ceefb121bd37718
z641e2371579932fbfed54c21490e5e78561d6de1437faab3565b2ec8031edf64c5bc2fc450ee0b
zff108bac7dcb6e25211f419691f9b6d364855f517cfa7eb42fdbb5e2ceace089eabec529f92856
z0f8dbf5301f1422abc1f2f9c164f7b33bac39b5d5e3cccbf2d8b90bfba21a23e0b8c5122931fe8
z34ce2343dfff5a7a6d26454ef955a361ba60d4c8a0751b12f4d70a2c01593b8e3c6fc9ad8fed1a
z69b2d9c9eca34d5e838320e9944ffd3f55052571d69589cd696505b55611aa421e53b131f0f040
z4e882313ec5c2957066eaf5b37b78a819b0e3cf6cac5e2638910d7e7d72c2124d64e050ccf5a05
z5d38ae96153c2f4eafadfda95c152acc1af2bf5407c3f435d86711439598d5bd04619d27337dd6
zfdf6fc3530be44805ea488dba50f6ce0c3513a56eab1e9a3fccc47dcc59086ec109c7a49105b36
z101e8af85dd6e18b666c8d2938e74b56d816236d4d3f4540b5f0836d4542e86463e56ab432e696
z7e0a6b29d96fc17304d200972d49d506807d82a2cc2b239d0caeff2e7ecd8645e188e0f400c120
zfa836cade47206dc8c8d6850cbb37bd0e90576b0eba490f310f3ee4968a0b4bb25cba7e1b3cd55
z12adecf503619385c0fcc984a41d16708847c3a8706be88619e881f7e01e5113e0caba7e2bfe6a
za84179929225f24a366b5507e5dffb91e8cbe59660dc96bf4f726dd99638e88f18dd14b531f0f0
zc84709e7b4b3dbfe83140c1d31aadcd20000233868cc6e92d19b83631ad0a0fc88b488f723caff
z89a61ef1d9d7abf7adef04aa83eb9128eb8cb1723a27da40b89cca7acce42cf0dbe16e20525c0b
z3eec04fea068dfcf23221fac5c04115c75fd48f018b79efa300c5951e91f65f289c564f9fc3615
z4b4e657cf2b178e0df6f175b255e9ca4672ba14838f2f707e7dd9d6cee06444f38da590d5cb1b3
z749175938b110e89fda5941469933739a7faccbcf886db6cd2ee1c1f74fd41f08c7e8731926590
z8305d808d64cfb26f10b88317dc4e0b23b1ad38388e63854814fff15a67d866c46e97e50a2eff6
z79ac3640cdd35db3abea91930be94ec05d6bb8d5b531d1e8899aec4ea879f528dfba719706adbd
z585cfa4159e8af736cda22ba86b9efa48d5196e96de8bbef1401fda888384fc2c33fba30459c53
zd4fcb779cf61f98e2343428b5224ff1a92590ccf5291eed521dc61eb72eb15949c75504c721a17
z7299cbadb4aa6e3cd0a4257ca7fdc462ddc9e52d74bfd2dfe0faf42da8f25e4c667e29051e1e57
zaf9322fcdbbc23643a7496a2cdd86ba6c7823dffcbd59b22629ad53586007b4ebc05b5537e92cf
z02d33a12a43f0e4afb07461b026e06813a97cc87bc96cd6952a35cbed23ca9bcc2bb4a3d7d4786
z0fa61427ad395309e30244d4350bb68db9f8e95ed367bfc654abdee0d82dc4cd1eadb6f0bcb811
zcdcdd5f4eafe0b23c1a54a8b614e8af956d40eb9263d5473ba5f2f2053846e9fa2bfd1e9c055ae
zef8c228fbe6fd27791451282e18b8de33d4caac83e2181c8b45f47478c4bcb6a21dd2961eea47e
z8d91ca3a2d6083fef89e15ceac1eab5406aadc8ed3d836ca9b6af1468546bf51a5c2a3883b6147
z9eef658aa88539daf0cf4acdf1c85fee5b2ce456593587f418e334b8b5754c43515b72bcfb40bc
zd163df574bda93d71ed05b5346c9917619ef09409a532d137b2089adc5294f94b4cb3276604d75
z11f5b60277ae371b5adb23c433d91f99bcef48b90c0e69d4b07861f101186550a5e2e8660a800e
zc69ea4c4427b7468a25ee39592e1b7ddfc644ff1c9a4b6ff7af328dbdb148dafd6f4ab41586565
z3c2a73accaa8f86300e191e079b474d99a85f283b4f84948dbd1cde12f25ae5b5fa19cd3651583
zc7c74837d69b54215565e7c9470d324f8395d9464302f66ce340c4ccc320b04468013dc01c1655
z60cf69339310dc4d7a99ff9f78dd3526b589f3b982dd6cfd1ca6c1dd453386fb12ef490a01e678
z7d610619f86d0b788419f9e5c6a6bc811fc7460772895d2c8f6d85846de5bef94755bd759f6da8
z4472a9ff94ddf45527cf1a1d1bdce63743400fba7dc9b19b8151d0cb03673249cfabbbc5816d06
zc2333e5c97be8638540ae478d43d7c90135cc7f1b698fe1bcfb3b0407de6440c9613765436f919
zd24b347e35a341191f0847c9d985184e350b9bfafebd9a64dab1dbc02a4a1052b5791f297e1e12
zc38a86a08d6dd96db40fa087194d84aef198d27d87868ff93a5a8d2c1175b27f708a76376c1526
zf25c056e88a23987c89ce72dbc2433977c77acd2625083bab15c7cce4bf3992348f177ee869336
z5433d98b5d19cd5341531d42a30cc31fdc3a360e0bb04e28ef1b6c52bc55bed84f77538ec1fb18
z8ffab4a438325a3babef3394b7d2845f1a8ac0b9059d00bfd706ca219ecdc1bdd03c640db2eea0
z15a44cce2c9e286ccc97203979dbdb1ff443eef683df1b4642360591627526906aab25404b820d
z77f8de64a39069e169209656945b6d422a9d32136f91785cf76beed4b9c5a1bb2fa0b3892196ac
z0e5dca239074e2a40905f3db2473b3c548a53788cb107bbc4c287af4f2aeb55e29e6647ffd18a6
z351b4a933bd543b336062ab354c33d1a8dc4cfb63d0f3954a14323b99ad1520e0a35ad5b90a7c0
zc45d09bc9777a9d4d168524cf6293fed1745495d103e35fea941808d03e39eb321657933bc3825
z4252def414f0cbbfbee8e63365b1d4ac7da3dde7183986f2725ef5158c7f97c0d17dc0f6b20341
z7d3116b8fb6435cb6483f22f8a9d825b3c73e5c58120b5aab1a6695ee10f563d9b44920e5c7b7a
z8e3852a746507c49d1b9dcfe5cf8ffd0b889b1f042e3aebede8d515d1fb7c2a32588eb6e434914
z0b2160152dd57b42e902bbd9619e8f91fee1724c567253ea932c90d9a3a4d60a36b5cd84e62ce3
zc8289671edf9c8f32c3fa61c29dc8f44f7a25c4718209ae46b089929709e117b058a34a0967c26
zd4102785df3606a6f3b4a1332ff9f7636fd689cf78a7c6b88d339492b7e48a00a5a0ca34d6a5f5
z9f3143d361316df897f9b5964632148b8030d9039c137f7a16292e54f801236b1a87abe3cecd25
zc6f4de3e11527d4413de03648c33a55dc5bd83710f210b57f602c551186c1ebbee80e3e8cc7cb5
z887ab037d5d586ed62d3dbaecfbc1bd4d3e278673dcb03c92e5b3e2639a41d1e2bb1e6db4205d3
z22c6f1b973910eaaba887cf3559e2b34a9c241ceb833cc2b9271ec3734e39a83ac0e47056fa8f8
z0e88884afc4c5f7a9f43ada5001bd5ec57596ffd1989ff3717a40d0cdacedeee5449579fb47362
zf1596bd8a0a1a6d0c18c921d548063350aa7722587da2935982f27c7db33639b6024c5a44938bd
z49612d2696f770e30a1f8467d9bce76dc1cc5ed226482426ef7d49c59ab605a53a3b5778511101
z6bcf1d0693b41820f0ed25a21c4b1bc058c90f92664715862c1b4e21605c4695dba39ac547b48a
zb17cc704e791b15a074d64823e08edf9e2a94e649738b7adf442b8aa007b5e53c4e879007e2c85
zcf661e011f05ffd68a47caee325b8ef6d78a5083e23dd3b455a1131fb99bde3df2820040d282c0
zdab35c2a4dbe001f0c5915111df0933ac80a7d2579d19d95115d7562b27a9ca4e9dfcdc9c3e84d
zb4f40d1f177a28f18b92c34b4b4eab62d7d66d02cfb27d777c435a619cd18ab6b53bd5fcefa866
zc270d3c38711146f3a97259135d804dd78a3d85b0d47ca9602322e87b40ed243168f1788f7312c
za81cb2ade2dd907646e10ac24509bcba33c12eec5539e652fe68b51f19e47335b5e6e65252d772
z4752931d2cce86a32cd387d5ee3df59e5bbf19e329575c11b5349901d6665f3ce561cd70ff2e27
za5b96fae0601f72ebc87414f8625d7449ea479cbfba985e6493423ecbf9ed5882d6ac58e222258
zd7740a42e6f3b2eb61a307f52a8f9d0c43d48b9d4a71330bf8babc052222060ac5bef08d35393a
z066c359d53f6d63367de2e2f151e7472589cccdba4cce352f3f26552d07c3dfa0768ab1a1cf34f
z1908fcd27553158aa27d886793d5b9cf99d9edb7e00cf799aa15deb3a91e9176d34f76868d1cdb
z76a282bf3b2fc40fc3fb2263bc92529f25b1c277c1addc99d2e751068724af10e9d2d1ac559ebb
zd5fe915a036b913b2da719fc1b4c32de32eceea652c70bf69a03ff8134d13a1a232963a3765af8
zbf113effa116879394d225ee370edcb16581244145dc253f2d2d0b052d3afe159d4a2d29803c35
z3ecf40cb7c5fa0b2a7667f7d86eee9e525873c78f689d455d3b594b7e375703bae2f1d8738211b
z147bb9d210a8372735957ab1ff59f7680496f621db3a606184ce9ae1de54aed330aa9186281cca
ze388207f064ffb50f28aae11d057908590a59bfdaa6ca5bcb48c9269b0026bf70ca62fd228c320
zf3a1ff3807b61ed5f879736fe573f515497622ba87b1bbcd95b0d75fb9cb3c7454e14ff062c167
z2b2711c518339670dc17335967b918ae410e6575526f73747012a647393c12b9d8d91d013d7c63
zc35a1809ed4e9706ba694f52dfa0bc4cf9a572d5705caeaff7b44c0176843fd87f47c48910cfd1
z6acdeb079622b203fec03939bbbf1f0611f4b0c2b8bf390bc2e179ea6aa374e64cdfdf7e2f348c
zd9524a237bbdef9582c8cdebbb128db314fea7d4db48079ddebb7fe94000b5af5d62f1aa0c8cd1
z9071be17dfc7310a735494018b1776c89ea3ffe2e023cc52a92435555777d092ddf65beeee36b1
z4b805dbfbe4e34c6c7c0c8a254cae53897fb64e52c91255fbac14a45b11815900d4685601535cf
z92c4b64db00cd43cd8a1e1d78b0d68362eaff04d4afc1b3095ffdb4cf3cb8f1bbc881bc514ae41
z37d8cbd261719cb03e613fb8f0b644721eda3cd2482970eb22930a9d463083aff477996fcef94d
z01d99fc723ce073f427bdf5b6647079a27dc7b7ce28e2583a65b1b124ed431ba48d4833ac690ef
z7f18f7601d3d825fc9e787571c71c4aafd61a233003f2e8c7e953995e398bb666be2e095876922
z03f338aa32ddeefc3e9ff08e3c90179148fa5b07688d9d8ee1a4d5b929c5a86724aff538de26d4
zaeea785defda7dc436dff06dc5125b0edbdf387f330083d4e3fc9f81923bfaa00b05941577696d
z8ed8f2a64c0f157c27230ad613619bc60adbcf7d9a89dc31bcb039adcfb7b83d0a39d0cfd42169
z50b49fd7cd938e48943e89cf287bee8bfe4bdef0f339a776881bf38459ef25c6209d59f8d1d1d5
zb4038740eab3eb16a436e467a3c6cd22040366efaba430e6b0cccbb44707db86fff05a4cedb30a
z96d91d9ac0ec6190caf39b33a6f713a15f7c927bbdf46b8fba004902db406515bba620e758cfa0
zf88006270c6d5c68146fba9722508122d271d2494d8ddca164a0564e3edbb9a95d70c327722924
z67350a825814a1e0253df4cda7795e8238904d94cc359999ad8e1b9c0e133f69246e6676fa51d7
z04a13d053a239328a107498a991249fb8178ee661b4155dbec53e2a8aa7bde8b9b03d901affbb9
zf0af4bd7cd7e1f25f2497a8ea32b150630619e02dc600d19f662538c7a85b42694a0f505c851cf
z372d311884a31998113046e5e5d004d661933e7aea335bacef66b27a190dbc6e712a00c53b6cce
za6cfe3b4f68f348ecf11082c7dbe5601386ba05e532e59583cfd8d5982047a48b03ddd07df719b
z4fc1c814967b6370a5d612210eae1a92e572e77452f319c7f5755af3072c09f3d47a3dc25b7b63
za10fd6debb71662541c6d123066d3cc06f2d90752051a61cc3a4522a068c10864cf71e8c2d3565
z4f3e343ca2ff2b6e25b8a7cd7cfc74c128ede18cbcf0c6dfaa0755f42417941ed62b8d4f0d3a86
zfa2c0545ea16600c4a9f54589ae4827221cb8c1f3530cb11df0c0107bb02fe7a9288985a80d8b8
zdce0c8a004abad3e647e3991d5f609b2092d099deeda8d6c750b142eff343e9583db7ff3be707d
z4db0ba9bfc41becd39b09e88af607ecd578d7a9641eb188b962b75e9f045f612db3ad718187bf4
z1df6c581f5d1494ad96e7c3df844da74ab1193ada2755813ffd6e33bff5ec232a4cf2a221d0e31
z3c2538215e8595bd1e472a5f339e7b95faa2a8d97d8590170ff1a4bbc05505dae61791143fc79f
zee92f121c60910e9e1377c64ae888ae82b04487e05148d316686195b5f7b19d5bdb1373d791210
z5ebf122b62077860dfb01ec0a909ca0bf74d0c5e1550c8bf5b7eb55c7be7934cd418935a40bfec
z14e986f479689bb6225edef76b73abfcb999138e857251255ab17710cc3d45918ba86b621f1c42
z611525f13bd10836837bdaf41e9f07a9682077c96fc9878a802e9df1fc5fab0d836c1f934c807e
zfa8391c8059880de6ed0df0650684ee104fe551e0fad46edbdcdad92061c139ce398c573766ce6
zd8110c78e1973e91bcde2c92ae68098ea4a8109e469d3a62e539810a786f21d008fea2db63256b
z3a47709e8b94ea0e6fbe4887bd5a0e43afb7cc50d5805ba8e65e63a4323d4e544dbeb5192afd6e
zdd3314ebe4b08cc1a129c749844515d137030cc5023df7eaf476f6a97eaed12759b8dcb5c52f74
zabe2f813581c599f385c7279e8747dd2480c6a455559524d7cf43ecfdaca1c1e45c2ce1ced0559
z77f750ea68907bf78525e9349881d678d15f759af460c4e26583ce3d05338e827115e64190ebfc
z6d101bb1ca1e117bdef6f2ac5f2372a8a9e4c32f122c73ad1c76af49868cd38cbfc19e95144c90
z7bad51438904a27d9da7de820bad3341c0630109126787b1cdf30ca4750db4fbba5bfccf678dc3
z75f345bb2241ebdf746c35b4ddca8c10fa041ae2c63e779823a6e458c1bcd7a6c30e5a464bdb39
zaee94a7b103c8776e301499d47e54442ecd3ac036deac0e1b62c3a81b983a3fdafcf01eb59276d
z39aaa5fe4bdb933724640e1a08df31fc68990a90bfcc3dab728f44bf8f5c7399d63371c49dabc4
zf8bd19ac32d6396f11fcd01299f422e219314cbeb59c1c916b56c3e91cbb879bfdf7d3d2caf6d7
ze96fe27a1a69c40dfea1a971925c4b11509f3e100f12eb13091734798b979aa87df0ad5e92c264
z1c98fddb19aa3b538e86b9da0945b34d37c9c1cc636b67c1972fa055c51b8003c61a66c2889ce6
z4c9b6fec4ee1af419ceb08c0bbe8374d4e97f9c735e302a955ecd382d43719c3649d3e46c2d584
z75b9891a277f901ecdc8a685ed599263ac7dcc08f6f9018f5a1fd837292a9fc2cc4518974eb59f
z66b190a60fa37e56d472bec4d9afe63e263f076040164517ddbbb276823583b78d9e575bd8e664
zd569b039cefbedf63fef18c5d8541c5e7271980c9f1a27fc198ef230d286f7f0bd825c2aadc848
z3fd5daaaa725f7dd9e6fecff0df21f59d3c63fd98235c40de02d791abc66a26a60c404dda730e1
z9090a4ef7eaa7e9deba9753a643ccb4c88babbe3a10360569c5f5154b7a5be3ec078d09aa90f33
z4bdd0ce0f50e9912336dd979e8282d5e14f259b6cf6568e8e5e7f5fdf3f82be06238ff816a02af
zea2bf37c2a9ee8e1c2f31d9adeda3e0f739f7251391a470910d255bcea5e4861e9bbc61dfca7c2
zdfde6c0710a6fc4dc345c44f9062f7af422e43fd11426c6a6f0b5f9a05a5bbd39099c13dfd7564
z2101bcf10f5bad03f55be1eef0089ae4f082791d60162cd523eb5fec1bf4fd047ee1414db4b27f
z2bd9ed696b091723952f57cea41c91653fe87eb2bcc344cbfc2643cf96702876dd6673b8e30846
z9248445567ca240a7bc65d612fcecdd5ade1f6b105754620a1c417a6e6c6c0590b90f18303f584
zd12a7a2db7b5e5ebf4731d10c3f08c960051f9076a614594fa548e1522eca4eb3f6b6c830c9d12
z51437b6ab7827ee079007e886ac93cfa5832966346f1ad572bec94e9a33efed22c600ada40cca6
z3e1260d241fe8318fab69cccf0bac27147be477da9b8a282ad9f826502e325687cbe077b653bbc
z679d2c6e7da724494cec183421b68017e517c7fe147987769014118b9cceb368ab2f1f2503fdf5
zfa8218a16935deb99ae6631be273d698c0fcd47bf7873e1d2a355e0c7a2978e654de3fadde2c95
zba70187d6b9f688ea5c5d1e3e9c982d21eea50debbb762f2bd04cbe96698857a80e408bb30da81
zce2a3d80cdf7fad46f0e17d6a1217ea6a617aea8ab5eb3c8a2b162f47626bf1b0371d415a3f30c
z4ff118f176eecee0d869d2eefa9ccd401cfd444905c48e9393799e2a916209401704cd0b07d248
z5efcfded018127d3bccab57268e556136b443255625eb3e91cd9fade8d90a72c913b377c06db97
z560d09522bd97d815d3240f8944d652c80ce38fc87449032e20a2aef34ffbe752b54c0de549783
z4f6745dd6bf6d488730a2b559f232b5921dc8510c22f19cbf2eec069b99af920653cc767f9630a
z07d5a99223e141b1c72dad1971bae7ab87f5ce737180a521afec71ce2190c4a422a22e91685fff
z2720952975038606ddccc250c0a413dd53d3dfb02da9469834a45e9a0e8ddd7f01be4b1c666bba
zf19649fa199b94bb6af892c8eedc74afdcfdec50632e43cf909c35af56a18ac069ea75987febf9
zef582839b56bf44f8f89bc83e1ee12ee5e75d6d463217fd25fd185a8fd51ce1257eca100d8026c
z75677b815e9f337cd5d28dae983e004ffccdfa410a536b409365475f3e2c6eedcc5dbffca92e8a
z58f132a3a12d83a3934d49e2f1dcfe0f7434f15bef6ccef8109d8a15deec28924e09705bad2809
ze8cd376d452e14ed1c0532e7f61ffd9e6c39b8e4d7e7b083a100e5c3379c35c7f3e050e1f5422a
zae0e7038c9211de3e1702a5aa1c97b58b646cf5113f0be5d9ea7907df766daadc972cf8e4f3924
za32a6087aae292d1c8315662b7a8fcddeea5b45ae44f4b1a66ff645d7e87fb289ece4793a37011
z217374d8b6145d2479de2390a2f116230c935e6cc8d46fae3054c1923485de3892117514c192f0
z31cac9f99540d4b3ea95c3d37da50f20d47e33a4cf52535cb2b750fa2ef233d48e6a025d18af06
z7d6486e846734ed6ae1606ddd794cc767a5cde7666b9fad437a3e62fae02325f6b23f4e7a36441
z970576b499f1f5575395c0d652ef73fa036e7f61da05da3ad53b386bd140103ddd623e3f83dcc0
z5b2dcb1fb8a76016dc685e100bde860028c18501c8b68ee93fd8040eee831cea2467975cbfadd5
z43829b04f8ca821803b27998f84d22b05fad0634469dbb851699236eda4db21336f1d9c3104ab9
zaa60227b3ae25e97063053c4a058f3fb2cbea8f4b505a76b246b0c312f39849ea85fae199d576a
zb394d5cc3ebcbe21576c2d5204bed61ecef3d59c0ade4c39edef19908f956b106fda8aaa47a4e0
z2eb9ee1313fb893935e24e2aae7965522989d9ed70c51b498f8f20a42886ea103297968abfa34a
z993ba17ddb5551dfa5b6f1887a7d9281c570c3254ba6e18885049f7567137481e39b6d52322776
zf8b759e29b93f9dbbe01695e8a090b851c0298364e26686b83ad45d045d2a21e4fbe3d6efd423d
z473217e4d096c18101842a3754de55858f5b1845b4ed833432064f16336f8496d184e129c1c6ec
zb7b45ce57b4c3b22e664e48febf2bb09d922eb7a7aca667a4551159baa3515b99a70488cb3a535
zc326d28e937e54a666f12f3648f3403df808e6b8f34c3cd21a51c5676cb8de2d6bb94a194fa8d2
za972fe67d1cf7130a33f3f4641fc400ef76aa5e32f33925361ae7c8d3d364d13c9a84a4404251d
zc4a4297c7d8bb0f6ab8caa72e186239a27043240800b6a4587bc913d03741b941bfba4fa1d0cfa
z08ab02facba46d417d5a761d90c4c6a11c1a8e0497bf7825af1e8bd0db18e7a0e1dbccadb32246
zd069ea7cd9395a566c6de37f0e93e1c8a828e8ccd1d54a706ded38adf61d6f490c30cf74d7861b
z0029fa5d96aa746a6a3bd5d903edc34ce4f9d55979a63709b684a615cdbeeb31833cf24ff30377
z11ffaa54e1fac0bfe5227f5fb367f7e4d6a2ab585e92604557fe7db4f133f425aae334559eafa2
zd1abc60443a98fea9fa4120d0afb5c59b4a6a9f5b03c0809c39f270005c744e3c5ffcbdddc72a8
za73ab58ba6c9c9cdd54f623387e31b6699e1ff3dd8b565b42660f7e121514c624c25dda9c6aa84
z7190d0089eb07bce70c02b70e6ed3dedfa37b7e70532f6659f095738b6e66bea86f3c31d684077
z73b8fb6824944915e72f4f511cf9dfb17f2224536e433f5dc4dcf5035f9e565c84f4c9e6ae5d92
z771e0aa5a4dc922943f28db475bf022d2fc2a53a91a34468b804fc29d4c3c7a2953b421382d5f9
z836874c57b03477888805ea156be5d9765289ca71cc04600c7f890ce7ca1dc52c4eb4ec3aba1ac
z0df611ff08e2ee3a97ffcba88d130f522a958367c2a68ea4e46275d80376d81d31cc5deaee8ab7
ze544bdd6258e98722a26b6645da34589f1fe7f7c1e6eab2d0bd16dd61a21ba05d03e72c1dad677
ze66c34d5634358db3c2fd98c1af4b111911dce501ba757fecc34ff67bcec92b63a13d7084cbdaf
z33375e2d0a5418f0aeaa3633191dcb04a4be9080940b95cd55ba1e9d79170807f1a61a7a214c56
zda6af88528568ada5b52cd80b1992533fb31af93a12f0a512d96b72359f47402899673f412c903
zb708165e4c51955296df21d851fe554234453f02b287a7e9665df189d8e832a06fec929db47e68
z3a79094fa04f0099412005b289fab8addd2ed332eccc1b05873e5b4c426c9c11de7a047b002a4d
z0cfdda40dde7c17145d4d02e26fd748c511e3aa66790c6ecb208652b453a5a7c8452d64c6f3d23
z1f99cf45ef35b7611a261b617e765a8648e53d61cf22fa626ff0efd2ad0a4c5c1ce03735bd7966
z4536306bbd06b2ff712ab9019a81277e8e55d2c99ab0baac6f939391e101acb05f63b77d5d57da
z90fe4a86007bc7d91f550862eada1ed9e42db5073359b7559d8676eb7ea6fafbe8a6528a8c54e0
z0bb43631530ea04bc6543f020a90b1bc40a56c2f2cfed2046a35f7f4fefa24d9a5f8c8d9b4f5f7
zf1e6cb4a8dece3f28e3e32e7402c8138f9c9ec28206067a546674138a77551b1606c938cda16a3
z02983319bfc41bb7409b6c9992df26cbede75d1fb1963903ea8d3164ecbe18d94d7e0abc7ef5af
z642cd4883a0e2f6ac66c74d72527c21fe98f0736eaebe480e6819568c7e852ad7326fbe38aabfe
zeadfc8f7d0a531b6d14d46cd4b2f4e2fa2fa815362e2476882ee9759a08195caa2d1b03da25dd1
z79d7fd66ddbc1f93bed9c5c7ffd5415af5ea171d9f204640184f8f671ac7169957a3d8b428dd73
z3b6e58f3411cfb81c051bc07257485acedb628ed869f8f948b5e07b81319b21b3ef698f40af24f
zbde8c5f61b8b8253a62ec613b658ea524206bf3b1e19a85463d9db682a65d960acf0414031bb52
ze4229f3ccec9faa4497ad60b072ef4ae1a6a6e0f307b3fd99ad3a29a11561b2cd7247d7b73b0ac
z75766c6f162b9c278233c108e319bd27fc91211b6059c60069b1bc9dd43c0e28beeff862bf4078
z246b5af69655884a0851d09e87a2a26f3d7a391cc99ef8fad253b93f9e6c7ceb5c36af59c7d141
z1d2d7129852fd73f7fe1aa4be3fe097c74055fcdc1916ca831ebe4e8f0bdc356370136fe9f46e3
z28e8499c0c9a7b25b23b66c7ac2d14c62458899c9961ef73261c6516b96339d0e2d9781e14c735
z821509c37b272a399a6835ea4ab6dfc9f01627f36f846339d1e928f3018aa3420b250bf0018160
z48930b88c8b19b7bf09f01401ac20ec5025bfc4f180d5cd8d4022e4657045d3e82811b2036c105
z9045c4a4801089d7e6174de0ebcf1e95dd06b1a2dab9655508848de3e301eb6c2b7ed30e28c40b
z09dfb4668cbb8e79e919e385cda0c2031f8637700c2e2f266a9617ae29f18e32f36d2bd4e81372
zc91c6ea858bd1f869364337c7db28fb11988c0318bec2ef38d71c57f9560406469681121b3f8cc
z8b6231b5b01020403a143d1c731b4c963d7fb711661cf8443d03e7d8826ed7d79181f69b6671c6
z6dfd1c267b2ca31cedf9b5aaf758f5c7196b557399987c196f805df3777bbf942d41ce758c84c1
zd090d5fae956d7d0a0c39475d956c95611cfadde9a805588fb4577a75212b0d766c3bc6b932d0e
ze362f008d8df76a90c3ffa2177bbbe70997086f695223211e2272a40939e53d399961e6dacb364
zf70221990b6033f9332ade8a39e9622c8a89d2932a464f9b686b84a4789142ed2410439f0e16b6
za086b5fb093268cb49d57b5aa70247afbca71681f28f47812c9e81db87b02011aac79549813d8a
ze1bd21f3fbb7b090355e742597075f4f7b74035c81f8bb986fdfc61752880916dee8d4d225fae5
zfc88f8ec0c6b761f17e5780484571f863e1b32f05af6ee0d8d742295abdb4e2e383601f5449e9f
z9f874ec4570acea4e8e2523d2841c5d9263944f51bd0046777e0aaa0a79ed71f444349cb70c86e
za462796f7131bf069170ccbcb4b4c8c53f86df5c6a296a785b30430c772cf1df2f462df74244e9
zb883fe309c00b2b2a38b7144340a1d35a5c45d01ae95e9c7368de48d7e3b60052d56e334143a10
z77d2a56259c13462fb42257a80a464344c8d202c5048ec70c7da5b3f616144990c0755517defab
z7a66d16a169c7701bf79395973653511d0069c9eab5a2769f6d46233c48d4049f9d65ba61e79d3
z66553cfb42246c9383836834cf9c0de33feacdf560c22463028b86f956d68c34407c942977e495
z1aa9b30518306289bab7a7335ccc07a3adfb0a9e77af2e035855ddb8a677234be227e658f66a69
za4b0985c34cbd8b702c50b190f61b539d09b7d7a0f57db81600db580900057828188a8aca5e8a5
z959b2f1c2412fbbe396de35505a3e7bab6b08997d6e153a7fbe9edb3e09b818474bab7b8793411
z517f3e1b77115176041b3817e92766ed220abd988b26876b3b749e6f696bf5a0b2e5d72b2f78c4
zdb8e5ca2afc9aa4d1a9010f2d22513d0c7400210908f46275e1b34d5bcd4e97b959692376a7672
z2b9f640f4e04da6a3f7cdb0313e6ca47b3fdfc26e7ebb063f952afeda8f8f746fbb1de6f78e517
z77e23ae099e074866abd8c557ff21e673b3e722b666777483289e6bfe13bbef07eabdbaea94f6e
z90dd8d34b962
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_i2c_state_machine.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
