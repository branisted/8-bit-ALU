`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc5fbb1ff3
zf1830148014fd9394d521ff27ffffb3b94f76e4b080857e93a2352915b210e68807cbfbca4e27b
za195dc4923906c2470609577cc88b90a3d575ddfd816d18827ec2bf0674dbe81d845821e0ad122
z8b1a4759824e7b4e4f5ab8bb7061b336da17bc459143590f1e1a86a1e1978e3fea2f56712e9dff
za7fa8285e8360d90b70c6bf496ffef5bd1b8edc7a1b6119aedc43f059186c637e24fb3fc9ceb91
zd8217f2a431dedb31f8e201346825065a0c68cdbe99dce9470ae6bf90dc1162ff1bf22aaf80988
zefb789c9fc451ec607267d5cb9c97b9b57c172f5fa3d551e6d6e59825082b665b9da20a3949d00
z407f5070eaa33c99559580c066e81268444d137808d713e451220c8d882de7adac1ee5721a05f2
z12b9464d1e981ff3d5aa54accec194392eb408c674207411cbf1b250d60971bb34e1551b8b243e
zcbcda459b543eebc91bce6ed215125decdce9015e1c4bceb75741bfa16a9845fb3b3a686cf29c2
zf8f9f7b04efe27ae187191da9209a3459cc34a23544fe4e1f89b5364a997aff350a99810c76dc5
z96cd7d22d3c1126fc9ea0f41c49e4b6a235408db19aa7e6f2dd4f974b10dc58274e1a11f85b43d
zefbd41144dbdfc792279f7ca742383d21059255d8770ca4adc37a102b4d26f39a0e61176888054
zb7c8a0fd30f404f009526b7bdc6265573da260a4c72e0edeca7b7271968ec6c17c89d971639833
z760839f0b3e985983e25e18d02f837abe061ee490379a84375a86bbe650115e5baaa4f10b59239
z038c7e71ea96992ab48e4160a365da93812a44d6e287a63e7793a4cee601e70251178de316d0ef
zadb7f4cff59ceab0b0dfa25d25c470cf44206b542d41c8c86a122640b719741215be4221ebd35b
zeb0e011a88d75670a7deeb7abd500b52a820477420cf4b1d74ec9972634226d726bf7653abc364
z037825de51480c580f56e6fb7ff4115c13df6d0224f07e07e55a907d4627806474b2a4330fdb26
z4be6abb5b73f49badfaa4467a7719ef49ae8557c0f7c7d9a04462bc78a7f9ef492fcd087b20894
z66bfa4f87466a38e721daa1f28012c0b30686ec66060e31136bc59083a1d5f4a108ae72278ddd9
z77157b8942e97c1caeb52dddedd3fa008762639317c6b56c08d9be349fae8cb962b3b458553c64
z132bd2758fa6fbf596adf0ac8766755cd975b3ac2854d8e1470a99ef2f1645f6c77ab516e13cf1
zd93bac6762b8a6e6c0341f6b642c1645178516b2d3fb301610efa55a5f1d5e998fe981b2815094
za0775ceda7dbab7022ef43505168a86806f4cf92fc2c9afc8167431265af1d4c5624d10b45d2f9
ze6b91d67edb6bc838b798cdb5027c9721477d55f5f10f550749092c9c6036ada97d94874db8851
z1ff98f493d9115d7d40b443afddf78c0c32f6e1624c56a13dc33d6582049983e09e86125be113e
z172a238402e2d5409aa740ba81b4196088eb145248a613da2a31eba561ca6ff0c76ed9ee5954c7
z6b5813488ea75e57ffe276ae3c3ef389667627cc4ae8ae42ad1be2e6987b92eb2fd8496892d432
z73be565b2fc8531317e02ca3faf683e922392ac01b342c5d502c3d5e004c4392a85be91907ce0a
zd074d08e46641712ca44af789f63534c9454136b27c72ec00a55f84976220b9bfb18d921218106
zc95e98d3fa8eb23e90b82842dd6b2495968b7ebe25e868ee45be669eff706ba3c742f0912a6939
z9c41886530c541d24c0e92c07baf765f7088b3698f8b024e30d57cfcde20fb947fea6a53d98a76
zb4d5cea34c3fb5e7d78cb7ffd697f4377150961df5bd8857347cd38b9712f02c60aa8a489852cf
z582aa496d1ec977ade875dcb182e213cb7c02e74e11e7ea4d8a5a8989d197aec69fcb3bb240966
z0a21d10eaf355483ebffd9fa8efe4e3b42b210ae7195e2be9f263020a481e99c235158e970b278
z943e7582a7a6cc44c8594943d2ec703d53b989c32fce8a49f38b9ff85f9538a9ec811b53356a8f
z9cb062e8cf3bf5b9adeb162346fc36ef406b681b072eb15ecb8ede5da9c9e84c69d768ea281cae
zb3522c7127989f71dcdc5198c647f18685514223f4afdd2c180d48ee7c6c59d91ce40f501087be
zb4c650238191a66974cb13d75660de76cee67c2f28464f7e891c4ad8f637764bfdbe63c744f9f8
z47f59c4b0ff653f4e4ebc1376dfb4ceae9c86c6a073b0eaf7acf436c7dea31f1289cf5f7d18212
zd38b491a80979efbb77ef102ebda2d9c78330e8edd0e5d529b7ea8edee52a5b0341a13cf20af4b
z8fd27873712a00b807b59f8413b2fcfba8800283ba5a87851530b29321493d2c4a6039d9448dd1
z96052373213b5002db880d88068ff4917783864f1e50a83186e63d36e1227dfbf9cc90e9bdda17
zbea7cbc78f286568330e9be60a492d33a5090d6863ce733735f80378cf45c23b63f77e92f5bf10
z7f01fbfa97d667b1493fb5597d6a494c14241116db992ca342a47677189957843eda78142ac9da
zdb6356991e5b1fa0a57c4995b6952bae4badfa8753c6c67d47bcb6048d94ba08fa43f176b5cbdd
z87a689b2ab7041d38bb793eac696e6229f5990881e3e3d253e0c9871dbdce456f6dd2ed85cd903
zc3ac945c29c0bf2bba2938c1b6fba0c1c8b24fffd15111d1d2c803e166bcbbf44032874e0c3841
ze20620b855ae7cdf8ca9255903b1f35ea0fe71903627c0674b6d0ed91a17b03a953a8cca43aa75
z38c42873b0a3ebf5689a6e3f254439ef5ba538baf6069a38db42ba8fd527166667b22e4c0c08a9
z47bee5e1a1f6e520244b9600a63ac293b9032bf4dbfea1c6a6df149da9b6ac8edba618f5778d8f
zc883a248e1576c45b863899cfc3675e77d15998a3c2e144d57588cd58be383237bb423e16ab489
za6f0f68d5f4b5d440c91cf762b6fef4176540a17cd02c78d46c93b16b283ce5172dbb8f47033f4
z1dbe02934af1013d7e66a73f3c704316e3ba864273cf910693f86015cbbeba6d58a21573dbb825
z050dfd302aee88d7627117a672d2996078aaa4048fe1ce628ec89815c3ebdf16886355b3a6dd62
zc75c391961edf39751a3632ee019809f4a442e1ef4a6eb81ec50340987bf984f16d325a372a193
z847200bbe578afa64b0a85bcd40d11ebc403961feecded04ff88770ff4daa5d9e9b2dbf2aea5ed
z96908f88102701ce32b9f2d8dd67451231cebd93b393857fa26dbc145b49c41c5ec2b7c89dd9b5
zf5ef278d2354a78c9df3aae4f1f4744e62645210aea7f89febb601a5dca34b278f2b8b4a9902fc
z418e28af2b3641abc7f4cadcba0715de44468a40bc43e9a5414922f137946211fbe6dc562c1329
z32d10897674504efdc9b6264e3f755468f33ad101d4668729564b799a88840ffbe85bf8fc3f417
z7bea069d8ebae7bab49a7cf90884ff9230bb6736dbe0cc1dd07bc9d6c829fdac9b4a30de3f77e0
zae5fff1017b56f2e0b0350cefe8a5de984bf2c400540ed9ff82f74955200686a918cf184c86816
zc4016263001fb2b6b08ca325b615b2e6b4226ef2d4eca24d2b332d47504b9421b0c555265e21b2
z106134175109e968c30e1e7d082cdf35b80374630873cd16a816f7c35f258706586dc0ba189fef
zbb3c6d2f1fb35a765b41e10474b526f127db7aa7b892ce25ec65cba21d30508116ba03dfab6182
z371ac33528c9d71ab696124038792460c67f86fedce2453eea5833ee5fc1dbf4605c7578c89f6f
ze11fa06a11ac7747ac5b39acd875f0d89d31c357efa7b67f9da9d638a169e8e68d59b1707449d3
z8525ab0a440a24cb52bd989af8fb33b35fb033e75979d627a64a772da2ce3705609ab7c1a466a1
z1df04a34688b0e21b677079bc30becd7d18c849a599aa9da7324692e5915401aed68f135862527
z53a8ea36040a0a1efa6540ae524b27a61a1427ad4def92feaf3fb0868748e6abe2f396f329639c
z07d341ab98cd95ceebfb5df64f6c92ece9885242028f8b898cc9be041ab84b054bdb764735f375
za38b5cbd9658a302a392b3bcdcb47fa7c97e5c516b0966c3a4902fa449603f655cfacdcb29d358
z0e4615c2ac5e800cfe14b3abba2443aec5f6276b600c5078c9efba05c2f74bb2ffec9b3af00f48
zb2cec9a41ede48c3bcf6b8031cef5a4ae72259610d62e6fffcdbd57aaabb8b622485bd4d0efc91
zf4255ea2f030156427441df9e3567a21341ddb5cdaafc16dae9c3bae6e72eab7e4e3c82c9dd8f9
zf50f46a8ad061af7d6f4936ab1391caac454a59f12f652be82ed165c41b1a07123f5263c4a686b
zeb796efb72531a95b47433b5b6c56a773f4b324f7861408f3d42027fa5bda67072b2210c8ed835
zdff0699ba2f61310253bcd2ef431deccbd216b9e366db0b77a14e6becbc5f11442a69808b2e57a
z32396ef6055102ee9a1de4da0f9187fcde76eaaa1cc07125853fa282a2a484e9662a036ec8eef2
z69c869dcda826ce33de80c2cefc95e2e69ece2a6375a86dff68108beb2875634abcb29518bd383
z05c050da6e216ca5d640cfce69ca8d2546cc944e352a1f2ad5d951adbf20aaf25c3bbb24f99ce9
z51931da7924b6af3d6f285897ba8e4c8e20d1695123bb7448ba4f7dbfc901b39b249da1b77951b
z709dc926f7b5a1d15bbbb2d31fd0e94961ea3fd347bad040b7963618bfe740e23405bbdfe0b527
z1c5a49d9f4ff4203eccf36671a05a84244a7865270d4b7d6ad1f9db8eede5d5142cd1a19c7680e
z6ad44d8bb3c8bdf07c5c16cf08bb73f944bc3b69fa2f926e3b13e8457a9e8adb58157544281c31
zacff9b3450827177465b2a22366f9f137bde2f054e79ce999117910d8eac4c8cf62cf3ac88e05d
zefbd8391e34300ead542cdc3951cb98a72a466617b0506376808334572d0b46809160210deedb0
zdfd74c04badf7606e257cdf47f9495fe748acd2c8db0bb3ee19c0b217f387427b6359b27f63181
zfa875bec350f88bfc2137b6c5f1e89e76297165332cbf817edc0cbb3fce54b93977fedd323edbd
z53faff41e5774ed0db143186873f0d2cd110cfee0f2674847db924dd4ddcab8fcb314a5e9408b6
z62ff8ad72b1f8a05d06ff6c0c02dbbb2bc4e6d8d63d4e9c27e252f7df307bd7a6f4ec373b1ce36
z027781c9f90e197e02b9ac8625bd82a62a829f312394a5da3ee7ce80af780097bfd9f2880aef8f
z96922f5e769ac39e7aac5510e6a2f34fe475eedbe5626cbbd110434cd806ae17a380fc692a59ae
z70ca1579051469932d3fc1d26f9576730afbbb507ae4b95464ffa4f9942bbe73d092d0dcdcbfae
z1a86070a9c86cfa19c8e8c8b988637f0c15c20a19d5de86b6e2c2036827517fdc20058c7c7677f
zec9ea2bbf23319db8464df08a7e6c42f8008879f192ab29a87636322e73397296e18ccceb7e069
z0e7e3e4cf5d7eed396ff021709c6bc711f9259369ce40eddbb6a47afd9b91b9b2e08f267009763
z0c27a206a9f015a9c6d1b9807d4b228a60aecf404d6305e4698119b3e0c29ed29d289e7ed6f187
z69fb00f4f7e671decc88456354dd974476a1f366154cd017099331949c4278e4e054a211cac2fc
z4f035398cee6e38ace042c04bec22877c860291a71f61964db7c73e74106c7323c369150241eaf
zf68a4229c30f767c9d33492db85fdfb958312fbf3b550220312f1bf17266863371a50b9a30d0cf
z356ecdd92d7e17c7d7648aa1ebf1753ae6ba2d7affbd115df89dcee5372315ee56e0447a2af741
z563eb6c31488046e50b41b77899f9b2b47d2412a5b6fa46188bd905517b4446882647ecca4656f
z166a52c6a76f342baae8b1914adca190ba8afb0417338d02aeb4552c46f7ef4bb9ffac553bc500
z24823611f5d00a6a90560fece596b16d86e9874289bffa7003aa295ad843b2f173323b799230c4
za3e2091394f44602aefdc6324969e85bb0a8d090935275e8fae3ae1d53073d8ee6dddbf5792bff
z3628b7e59fee00b99f9e0e0a9758720c566c60fc2adb1fb5d82d220f60006392ab96ad928fd586
z62e84c37ac8018f8fca757349d1a8ed39242f6d67621a46a0a7453f137f45c9a391e5595579790
z6b81a664cdd1e08391bd86390202a30153c7916273cbe1b5c7f2597321faa0ea97f87d9bbe9b9c
zef38a81e9bb988d0263ce216c538050e1feb316bfd122eeaa48ba13ea4d499a1479c1f63259c88
zbf3cfd5cbea4d9e697af69978c17edade5a7af7937815d1fa599416b0a2bf4be44255bd74d9bc3
z89b0da206c5bb68832d64a7be8f1d9ac0bf163705c39c256de46537a6b53cc1b49bc889507c151
z190df73436344e340d9607b1b83859ab0ac1cf7ab7d135f1c8315ada4519a5ba6a9c9d1e12736d
z261b92414d0336dc88bfc27f6224e1e55ffbae9e3ef0ff544437feae5749b10977d82e47f19d48
z74acb271a3be7289b92ce74c3418385d5a23cac06a931ff47a55c3ec60285f499a2e52a780f7ed
z7860ad217dd6a90ccd04a05b4e96784e1f237833214e3cdb473b7d122d0a4121976aed22f5d802
zcfc830bf2793da663ac86e5bcabaf51abc347539672f6fa1ceedc0ddd24adfb652551145dd4f01
z8c7867e90994263c208f0ca60b186d2718ee29cc193a01270e76c0b14e09466dc75eebdb0cf398
z1fe1f8212523382b1ca171964074c50e91cc43c4b8690400fb201ce3898f5009ebf89531884889
z3ecaca7d1546e0fbde7dedde5870c2c3afe40d8a68e4b2bc1c3ea725a38b59a6328946d288f92b
zb40a07c6d686f0b127d2b181b6efa7739196bd1f9b381fac2b082802e13e0d21ad5ac700ca739e
z2ca2a71f63d42261486c9a9bf23269953843f263d0559ffbaf557530ab8b8d1ec8aee75c64c601
z11a23212fc97de7e3e684c927f376a5bb03c0142d305dc270e1da34d070cf5bb8981537080b7c8
z13bac53480bd6a7ec8895800f2aa7c32881fb426f2a66a88a349d87e454f73c6e0a3248502bf0e
zf5f18b5a423d3f4b4cdbcd35e4f9dc929723a5e4b97e0ff79f5c91f7415de964830530da2ed108
z7991c533ac503b1ec3898ce55c7562b8eba8220961a4e78ce67abbd6d2788ff1ad72183ddbcd8e
z1af36ec21c5204c18504c304184a51e3b5becdf304ef7caa1341c5322ef81ce8204e427bbe7d54
z27484efc69cc972610da8feca8560bf9ff19dc684a65ffb42dee6dd00884d678668f84e5ea544b
z2af15b3a5cd8b177998dfff8bdf418ac872df8ec150fdb2ff678179968101fee2f1dcaf9bf174b
z7bdac0f264b8f1453e95e23820fbb07c5da4f466acdd907568c378321d526070a15497ff1c79bf
zd90b20fd3b7036e446065d4b60c4131e41e1efbc911af5edeb164731af29a69a81d2c07092ec52
z98581fd513049cbc32881a56d3e1eaf5f9afb3fd4b0b8af1a0e3047833ba71582d8d54f17c4375
z017535bc18738b0e9cd22c02948b943b368a15b9efc8ebbb4c40fd122753790c5fd7f0b2e036d9
z8f580f0be079ab65f93555742d4155e457ca3c9870f3c8181c772d2e77123c47d1d40062ab2082
zbd4efe9a725736e00d144dde236eb719509ca0fa592705f0de6ac1aafe7bdfbd0b8435e8c6c89d
z8cb190565ef6b88c8bf2ae68ce60490a3c2ddcc805b01347e1987bdb52284dbfcebde15d4de0fd
z6ec679020370daddb5d5a855b33f6be8ce5ade7caf20b8ff8d4536bb779a4946229daeae4dee65
z6e8a010b86d3c6e64b69259cfb44cfaa42090a5d1bd4483f6bcb04e63dc38708957680bd4da06c
z98e59646b7b62cfc4c0447a0add0399301c9ee2341ddc5f93d0bc0e6a9d7c00c75ad120e136935
zc6b3a5ecef0b9c6b87ae8a0e9ab8f02043fe9e8ed239acf523e271fbd24cb642300424942f2f8a
ze47940918632ad192b6ce382bdb8d6a20441bc7aafc037a5e80c9138390b5676bfd6231c9a096d
zbc42556a80cdd792ddc548aa357810ba84deaf7505ebd51f679397b674c950d44987a0456eb6d2
z067d81164a100bd103d6ac72b4ceda559151255910dfb5632358fd10fd00ed9503697159d421bb
zfe6588a50a4d28dbf95e988b53a82ade66474aca093fffeab0d4c8970d2423d7683cb8574e2ff6
za36f0db9cd087b536305aa7a1fdac65d756a035fe97cd6452c070ab1f35855ea2c2fa734422788
z142812b4f0f6caa0b276c5bb335298db2e08b8a280c9a982a2b4ba049c414fc87e9c226726ba5c
z2e042be06a3ba0b95c1cd7ced3fb96722aa1a74ca3143770f2cfa86136f0bea3b7c92dc2d0bd98
z8567dd5c7a48aab3dad0c1cb675ccf1941b2e20a595008171a92934d37a6659c6ee31db29e2185
zcdaad0ab639e02bc496f8aa79fd1206e87bf4e734b6cd2e328affafdc582a90bba100c2cd36639
zd43234e5bb8a22e7c10e7f1ba70c66a55c9437bb3fe754cb43b255db3ca355a733ee59f7a59975
zacac6b34bee5f73a8c220d9484783833f780e9a2e56403124b4aa8f1dd1b78c2b91d7cc23c1a6a
z58f652fdb06a064c9331093580971aa41c6cd6658d8a49b0bbfa39072eda05067e6fa5cba43299
z34bb4baefd536a4804720b55523e525bc09bbe5c254a852810470abdc64103c4a628d684293ff8
z7266ad98474851a4645ed22b8c3baab08ff82e901d75ec203c3921bc29fa13531388a51003ee52
za1891656ef1e3b103713c2656efcbf8e08203fe0eef06d8213a81265948dd7b0b13717436d9f4f
zea7a02f91083758f4ff3dd23b301247cf301d3e57493331e65e75c26075b7c31ebfa626d8e5f08
zf52c550dbb0c8e4c64d020c0237d68490522a528611954ad5628b262ca7a0b848fb3185f7b8638
zb1e1130738604c04c826236064b89e84d3550b20d6c3457f1dd333a95aad00fc4e4a1878477f8b
z36a255ba26841d548f0b0b62b452631935d437ca7dc92124032a1baf96859dbeb3ee86eb0fef5c
zceeea2d2fba148d3c7b33e0aaba1e4adf248970ecf37112ee0e5e72941994de68750c258f3ece1
zb076dfdd090528217961b7f2b3fc78ec681da570f71755ac42d879c979af2c4ebf639ccbf9c636
z4eb3866e2734337756262179cfffc83349cf043b1c61620570294ff311f2077a267ecd3f438bf3
zaec5dcec8ee102c39922b555479e87d1b300b5588db76cab2b964b305ece7b3cacef3ba2a31da7
z24230eba8d00e3bf5b3e0d41a841741a6f711bba4912c55685d82948bbd9aed09fffe3f54099a7
z44d3d41cbc4dba99b1902eb21a507c67287dc852bfc745f57287a9c7320f95a4b606a5ce62ba38
zc9da98987323d81a59afd225cc604da2d10c33cf35bf50456cc242ccf6e5a05385109173c38b04
z8a65af8b12b2296b4ad4b2edea7e80452d1587f8ded459e52389b2e927771b8a7c471926803e71
z87c958f3007ed749ff9f2ac1c34af0ce1d5ead5a47429f428a0d7623be92a5a8f3b61def0bd3e0
z1d3623aebd0df4ee45fb6767369792a813cc9e5d993d42e532e0c9c767c4916f81343b616113b0
z408496a77992245ad0b87dda4f911eb7cb78d2cadd1376d97c075c64b023f1456100562f395435
za9c7734c540d66d99247dcd6d586a8a128ad4a580b74ad26bfebfba4faf9fc5e6cd447208541f9
z88c1e263d7e937861c8e7f88a80e7e8431c6c904397e812d9e263676ad77383852898c4c2d5fc5
z8eaa6263286f9600dd10ea4b9c1e72acc6105df70f5bbf7c4cf75031d36f2a418146745346bef4
zc9ebb533d89029692d6022e97a7024e8fa2ad728395bf8d4ab2cc3c267d3223c779dd7b103d61f
z4b5d389351cbd8cdf94cb81010f9a6151a708ca7e4256d62a194599b655fdbbf50c08833237313
zd06e398c10475f43582eb96628ce553a308ce76f994eac3782edc98eb6a7faf89a8633bc25c449
z56f0371320b3d4734e5bae35a31a37ef9e77ec9acac6438c71d3e3e763e37c804d89bac9a27819
z9199554b8b718586d9a46db84cfb55ab6fd6cda58faf399f06c4e4eb75c4e47c535df77cfb6263
z3f01eeb2daca08145667113aa92c9b599ab3152511c9897b3d4f6d5410de6d8c1d177babe2d251
z912133eff8f0f8f11927414d7045777be2e87da5f9cc03ffaac268cb97fcefdf79be87ac6753ad
zbfc4d22b9b296cb5d33c77f364e14999acac7f94c216b37c0faeabc8f85faaac8d5200e50a0ba4
z336128d0dece5e7cf9f52a3c9fe65df80dc23598ff65dee0b01ba14b5f4ede10d08d5a9a7730fe
zefa596b1813c3d154384a381f7604fd148611edc400002946bba3aa873ce081a1013cdfaadf0a0
z2e7ce02e30fa1a851b89976cdda5cf8c97df5fb80676d7e952270ea69b63617c796b7423e4181b
z7ded3441b6ae66a182d9b0f20a841694a80d98938cc6bfbed27f6f4ad38683022c05e7eb79d466
z5db2fa46908ea1fb98b31165099b7cb935f165ae0308d3022be9314a3cb3230c150280cb0783de
zf299fe92b4a8aa681105f19b70ac0d74518bbbe21a559fa673dcc766d0137dc5a92d8d52ef3ee9
z60672eacb2ea022e47ac640bd691fb8681a5bce800b1e3cb7d0743b8c4cc2d5e68d0381252628d
z35fa7046257f987a912642a88655013c426e2b2d1a5a163983ef365cbedabc8574bf7f2696ac64
z546037720a30066001b8abbc3e6e2b47a7db2b0601d31d7167c47f5a3b5b02ea70237632a3731d
zfd3039409b5cff26ff7a4726bbd7d771ff16f6dea7b7a417ac9d34dd622bc6c5d667cb3817c0cb
z2232121c02dcdad7429d7eca47c90d0275849b14209c2c8fbee9ce6eff16a397e943f591d060b4
z674a4fa4ab8415295891642ead421af2af9251f9d5f6203bcc0ae09bd5fe18ae98a94557313526
z954291479bcd54f66aafd00ef990cfc007c40af0330bd8ccca2c8631af6e1b1b2f261157ca2069
z75136378a93a9f7403dd8e91426836f3880a91326d47bb78f6dd1efad2db57acc924ee8663abf6
z2f860b8c0fc3bc712fe196321217ceaab9988bc80ac913ef074c0f1e1abc564c784bdb0daba090
zc4a9a7bd454e56d4ad21b4910c0d7322004b28ee819073c84a8be61da3de29afae6672bfbc1439
zc255ff1f831d9868d63ab285658fcf8adca71789380bde9a4aee7d35735f9b169fef16ab7e8a80
z09f8571b83f89baff1975b651d8c24ca42532d1fb737a571d6354520996553ace044b5bac47b89
z2313f8e009ccff85c3fd603d74b7790d0f931cbe4e01008a7c95e9a0736ee5b269a465c6888b8e
zd15781251c492f06f55b57aaf850a19f6008267bf9e5b3a2cd7bb13ba3ae5e14162df5c90a164f
z8192dada5e7603f4144e7fc42ae2bdaace431a1512e9dfa9e4e647c7f0c8f0c64a9fd210590737
z8d284afd616917d7d2e3f8d249366ddbe0f685eb30a7a8c9683591f1488d4daec5628b11362497
z98b746d519acaa40c18ba0b1bbc0d638770e5488ed931205a93768e409fb0affce147d5990d500
zfdbd07721175d8ea479090c6326a2bc3a82fec3c89c501faa34db914b99a100212010d72cc7d72
z3abe2d0e1b60da16b34e51eb21bd806c394837242db951d6129a226507ab498e80f645c0f9aa05
z13762f568115d9404a5590e2f0c12221c8b1c04958b81734b10ae145134d827cd734a8ed8cc05a
zf24b340ac6b98abc085db43ac1e481e6bcb56f2aecbe2490e99a97b803b6ee597cb4d100a64ebd
zb4f387fe96f61e5b737a528773812211c0a9d4492c86385f46f483fbe7227d76666ba20719752f
zc58c07f03a0a795cf88830783e43598ae9b8e3c70c07fb0ad9901630bb973dc509e9c177f107bf
ze6758b76538426d76ee7216591679d19d5beb76e0db0b631478b60abf197e00c305d4b045ac5a1
z27f3905e8e446ccdce4895f2e08b32bb01bac888dee3f4e208584ba95192e17950f852e709a52f
ze85d593ff187676b7c912f00e8d13ba5ae8b3a4cb35e91c17e13260b2f8c31c631caff65a91121
z12fd2aef73c3d5ce0a3e583a2f1099f169a6a049a218c73dc9d36280c9865de71c379542118462
z30b2ac059cf6899aa7ebd5335db66dbe34eea2991f24db562f946239b040a479aa2b7f3c3e6e4e
z3183712fe41e235805bb44d468194684ab87be059af0a0f5f6862b255e39c632b75adbf71d724c
z193018e8fd7ec5f3d502322d685fbb6fbe27a83c940733036f30b1c315265b1d9348c56b47b91d
z53bc570141533af0f2baf73af4f47aaae520250734c14f43fe798aa6110caef864572183b65acb
zcee26d9bb386f6ace6403e7e2dfe51d1389f5a0544c4c8f0bb3924359859c42645519a770766ec
za04ae9c495c717d5002d828bc78184e85e724a0329ae203a2977476e564b3b8f7cd961d77a9b89
z8376f3d71a2680316800a24afcd086c52ffacdad5fbe1f7138c817b66827968f3e1db249e5d7f5
z66b5dab32777dd61d845094acee583d346a220d4b2b905f960d06eafa322bedd2c85a612952125
zf38e11b2144bee970105d2ebbbb84c7a76c645f832a0f434062aa5a2d994c6c0f290a2215eb074
z47f087d6b42122a15abcd9306471286db06c13e05cbb46c3d69ae1bb81130e9d0123481fac2395
z117b5a1a307fe19ab3ecefe4ef76ef2e2fd35937ea26ebe9c71532825ea00ac4df129174bf5b1a
zec3e0b3551f9abb32edc4f1794acd7e171ec92d8fd1de39af3a9fa82bccfe95d9b7752ef3cd3e1
z4a71115b688b00c059feb60784fc02f0bdd9d3dd3a2241a6e98dd1b2493d7f5ad9a6adf1db8f22
z15f0cf7bedbe52b40b3d01893f4b6d179b7fd75d08a75b00b3f69c64e9ac933af4209725c2aefe
ze32517422b786e1c7d8b2cf8d2bcf748f6c058bdc50c4440e7a970de43822eeaab188411db17cc
z7b55f0f38898c39af0eab921b58ab6138610bdb5cf887e1c6dd0ff034542d75a7875802b81a137
z26ef9bfa5e47db07060826934bddee4407bb2c87dd1eb6f835b8bfaaa3c9a4792a9deddd0d5b8f
zea2824b768b663b5f9d1b1d2a46853d103909e19a703c9255ae0e3c5dabcdb7549cef804e63a5d
zb683986f87dd78d8b03c60d9175940312558232f6e6be37d250fd8a818f2b51475d7b4cb182479
zf98d0382bb13257171f64ad8889964256dc9a9447018c8e14c11d331b156946d715a3b62e02c3c
z6f74322c224195657205f6fdcc87f07ac87c56f98df7b89dbc941746e6ebc72fa88f13b7a05c7f
zef6cc03d061725ae547f723a3f5d59fd69df5402a6e7bfb75d0d9f5b3b51b9a8dd2020fc5de24b
z0c3bd3478c6903f34085eaf2649bf9d0ea357233e0d2609a4e9a4270ab2a4440856e691dca79f3
za3f87a2648d191d459443a15badea71ec710dc2ef2a3e87cc9a68ae4905fd3402d4da23e190a86
z67fa2f2939a7e680c2a112ffc57f9b35e49b354ff2fccfd7181bd13940b9b518c9b8ff87208c26
z0d6eb4515d087bc68d44b11485b317043df3928958cb65272d15a1c7fed69317fc30834213e1fa
z83d4778c01f600013e5d9c71ed4d1abb65c507abc91bf9912d6a254ead4f3c419d82d122870b5c
z15bb76c8b0cd3d0db73b60d9dba741e6530c0f6c4d0db66bf54e1b27796dfe99c21c1f9474b230
z57bda5c8c5e121c193a68ea7079c12009fe6a93e721d165104b8daa5e36995068fdf28f9e6a4b8
zad6b25e6e5a4a1139e7351ad5f00cf037438696ce0a8e4b4875327057f6fd1e6da5e31f6c2db50
zf3d7910908d40fa02b0750842fb48ad55d7ce56746b75166c85aa85e2d7a03e5d09fb85f096420
z44ca2aacc824511faf8355ecf9d75a2294ec5de7eafde8bca857801c7b7e2739909fa4b878b1da
z79d568701ec3f52e2cc46dd6eef9140645b8eab6b96f99bc0fa4e86cf6c735e972d9d58546a4f7
z8c5313a45b4ba1e4b1c6f67bf23c52f3b6b299fa3b39ced2cd4a622e91a05e9609704a99de8696
z262df6924f8a8cc17da5d3e06846606550283ab36a9ef4b040754d5786c885fa49b034aea6e567
z67367f43eb45a82cbd43b27c53b80bae42e097df21b4385565a64a01300a24027fd7eafc705115
z5155bf9cc4e64824d3253adf7373b15f1624150c861ea4836c9055a6740f9c7033c30e33f15add
z054cdd50caaa8a3e3b2c2b9dbabe59df469b96b8e3644524e0773d4fa284155b81d9df5bb62fae
z96f377363b19a3ea6c062a993f620ed342a471de03a6904232371de77e46362256a6a4cc768f5d
z011a050d9f8404564746af9e6c3ec729bfe0e09a180bc6513aca95d6605d7133232032775d73de
zf5c8e11a68521d2b7991d609e77706e9178e41384e281cbcbabed397ba83e14409c1ee1a7e63d6
z9df0b9f7dc3547671c9583e0804b274ebec396c1473dc59232e65114731ad5c8fe649c5aec0d72
ze95bf8614df2d738b4ba318856c18e16e0ba50b2f8b181c38eaf94a86d6532c319e50a390bb3a0
z2222244d8b7d177cfcc932f7656152ea02bae7f36a2bcd1b4fe497c69e80c023575775c4cec771
z73459935b395e3984b54419b12a6713fc734c486518f6be8dc3d1a36cec5fa3cb726e35af8dc87
z2d5196948b764737e486c03991092a6e1331fd700f12bb96411c7d1547ee20a184434675bd64ba
zb0589ca699418608bf7318a956832abab256ea5768be789ce74b5c5bf31cffbf3054c6e403160b
z8d1b26d072a64865bd139f5b7f18419a59b5a1df09cf516976194a57f6a13d41fcf160a274ffa6
z9be0fed518f0b89219d7d2b60b8e4a93984b0b41199afc0f92b777b0052e8fbb4e4ea55a16a8e4
z8a1ece0369e8490348a829f68ac3b37faa27a6f6d07c322c185f34c865a353278add3b4276c421
z25e09025e235733282aa0e1883bb9da4bc99fcc860d6fb379e6e06c42dc47ad0f5dd744b3db157
z5f552b914505a6dc53adf9ab38d6fbae80eae4fcf251eb36bd9eec59f0a6db75452408122e620a
z965a66661682b0485fcae801c03f3125206cadc323d574c9d3e610283b012e0c5e8492cdf0a2fc
z4ef9b36eae16279a2a334aa7ee1ad6772ec5a95ce689dd6d58a0087accab1992f72ed388806f96
z31a94af1d7abbf5bf0aebe6f36521d0b101c867e84801fa009142b9583c4d49bb935e32d981834
z3c118b5e20e193226e08c78170d098ff1255c7834b0282be339778334e2c790c3756e25b2b8e04
z21a3c9fb084b28b8ef9d3443ac4c9e288bcff589c61828b537d386efec94b0d921a2551efc2e13
z43fb567e135138432ead1b461e8632ec3c520e66b764e4ad05bf86e1fde00cb47fd04884d1035c
z0471afe16f0efa9bda7137027c8515474531eed037dc3ad802b7ebf723844d0645bbd95323b84c
ze0e424ecf7b44887a176790f10a7763e4b1de23b302338cb5dc4d28eeabbc673a1ca76e33151fd
zd37209f9047495a4f88a8ace9f57958c43b30ba6cb3ffcd1b570f997178cf9d4681c6de5c18c05
zd674304e830861db188a7d682f75c6e13b5d8617a88c4fd69f7ef84dd7dc9c6b4df3071a23f96f
zb3193c36f2cce8b831a2a23a8c6ae65ef109fb718a36cb4f13b159b7b348bbd141d40eb98b7c12
z359c3b39e9c6394422cb4e0554523ff024bd32cd6f242d5cee028a382d62661dd90af36a1c76f9
ze86327699518023111079582420a9e4665a5c0df621525bdcdb12f612f219cd91efc586a67476c
z3b161fcea99bf38118d9e8e83eec4c6847eae4c49032e6fe23c3ab45f309175256f94474e3b242
z5b8ddd0164a9938dd9fd798d9f84ee1ca48bafb9500a7bab3cff164b55d520736633d7575f825c
z70fe2c64f04c2d74ac0f63f79cd71c08414bb6029e6f9a79f392b2660359ca9b3e298ae422aca2
ze20ba24d5fdab37c8d22b6f4c0c5adb1fbcebc2d28b94e5768352813eccb24d12530909c6f17dc
zd1746aa0d9069bfef9d1102fd85ecc2f2646e9501d72c81fafa6db0cadd524c4069438088c0bfb
z5022febe0b08d76debedc8d96531d6d8d07ee935027847280dd12b900fd512ba1656cc732bffb5
z2db5de1ccef523dd0b0462fb23e097bd4fd8d665aef34577a8af91e9d66016b36f4ddd8d0d489f
z49f1aa355cde443551abed9c6a22baaeea8b45229afe03c615b1ebe4778b719c5686b238099e88
z4557ec55da2f142ab82dc11358191ebcd0f17239ce70225f7175db7f83f6fbb6c63ff87afff794
z9167f46493edd1b839990f22cf91fad658c897735d37667e30cb74d690eda1e17f57ef5c9dfce0
zfae1615c31a63c4fdf100e0e4bfcd38e4aaf9333ede81c95204a7c56200b74b08971b56320a900
zcfec0e1719edf6f80fb0800e50e02151360de0d5db736d797bc6f836cd283e71a3d1970afaedbf
z7eeaa6d72eb740d84fc3b6fe3f1966cf97002a9d97342e2a45206be8c3f087ef208563d53d0167
z3e0a52da4eb5f6a8657e04accdf3f8cfda753d84520f45e5cb39504c5e67b9243a46d1f17fb6af
zebefef138ce3251fc92db472af230b352aa8af7034c3aff52e140ad06d4d4f8e0b149f79805be7
zcbf0715a4146459855ecc2cb5008def06063c7087ba96e8430eb58429f8a94f4c1c718bedc553b
zfaae3524ec98de0a6b72349761a346541feaad1f3c24aed775560392f4f1a7e93401c8aa5f8079
z9f9f2c61b884890a22d2da38b989120ca9808aa7f021e65dcfe8c31b552571a7d59a489a07a64c
zc6c6b100b711c7328620a4ce4850916bd514b074a46c86fe8a48bcda3a6ae06e272fb971550e8b
z1d0275ef3eab4da24ce87a81ae01321c1cda336744426a048911dba8ba48a49453fad1aa8e315b
zfeb92ae8a416ca4dab557f575545058301c428e6081a26ba018da8000fd19faa8fee99842f9db3
zd2080b0254a619e04f582672869b2f6ef27b8cb168e6283e7303bdc7696e9c8df0f117e6adc678
z568fb85ffb93cd95e676f5a178c27597107d7d092dae84ca50dabc6ffd6afe7620b38e1481bf54
z1a6ed6374877bce3393f4a5e54a26caac1696e24ab80b706dfefee2af08d4680c7105c2ac3776b
z742e1c8acda64054f69f189206ea42dd50bfd748d13af6d4ba7808f2e76322196562f7b8ec36bd
z6ddc755e62a646403a9abb4ee6a69871537eb2cc15899d3bac226c1c8db0beb991390bfc42368a
z6827ef21725aca1c698060aebf88cc97b15043c61b9aab0192ad981d068dd1d981284baad4620a
zde5670a6eb70e1271ce8a2616d2eb71c8c2ff0368826d7dbe193fbffe7d7e4d56800575effa751
z62e6730b0d500a17354c6f1f2fe71193f908db1c5e9b74957e63b814f22658ef1126dbfd93a527
zb9f059a66c96596658e81f8fb995d836473e59d88f79f078844f227313495f5ec8852d5a18bc3f
z7fa922c9f46a4a75b99ff7feecb7338c551969203989a945f9e295f090ffcef174afd2762fe2cc
z376e3fc20a82fc131c72ed9c08d0e4c51bbcc95db35d1526672bb22523268b8dd5208e4767f893
z29ce1a36c37392c6db0e08b432ec608a739acb60030002b3681c73379cb498ecea1014139d5619
zc159804d9c3dbfbc1e8ef1041bace63527b3183d5a8a6f4a9449c389cd42ca91af10fce06be8ff
z35579f3d2dc459e9156f939cf41b1ff399a35eed76120314b24b3860480a99a4a61e11189dd915
z43891da28a4779738a8afe3e906f7cf472ebe892fdfa21c8dc842fe075ef90440949f0978707dc
zf016ca2e4928d03cd030ea09b99ff7b6619f779f7c85ce78561a35f341677f2b06926ed2a87bd3
z882a587d3e83ae717301287ec5158bb67e489bf5cba7eb5349606a7145666d01b48d538065f4aa
z9eb3b2849ee80d07db1ed30e582768a5b6d6ad9de91f23c228dba9c3903ee63d9a5c1a36849047
z40fa959916b76abf71632f09f5fb40f56b60046657dfe4c00ee64b41be511bed73884beb629ed4
z2989476b38934c9f45c39916573e638f7be2e7f839d064511fa6383fd9ecd0708c403631710d33
zc2aa638750d04f052b8b6bbfc2d9bd40a2e65d7c244a1260e48100be4583288f1f325b4280d1b8
zecaa32197af8feafc460c7d0256be3bb351fa07d82e46c0fa90bd99e60b40f07e0f6df6947e89c
z1e80c6ef25e6cf3269fcc2569f86e206ad13b7c2f51d1955454c85d6ebd7ecc0e8d279acd26615
z797c6c03b6f281a428f63ff131e0dfef8238788efddede75b475c8e3d78b37f400f369ebd15ba7
zc288d59abcddc4518d4bb89d4763c19ab3e51413ba264d222279af36363952dc3083300a5a075b
zf8887e256d10924822e468fbeb0f9304777643a9e1ea51f2456c9f0a428f4c8f40b73962733558
z8e3c6f763619cdb2cde242f9cd4ec0d4f8b0ec738b29f760330fd979e480223dbd054f600186ee
z4f08d56af9f1741836fd7f044c3d69fd0987543d8118aff4e18d350e0feee9c2e315233c72a42c
z3818db0ee65645a3aee3edcb13a2a16e3f5dd2b894dd16118eecc70989c54417ded153a37ce616
z25687300d93c3da9f96a4e1c0d7df644d0778bce1d79fdb3d3cc0c2696c5c114978c20f5c78da1
z10877a3ead453b0562e97d95c18bfd3843ca804e317b91afea9da74287a463af8d9c70d3532269
zd6ba578d8abe5678264472794e108236a44bc883581e3bc004510b3a7d735a93cd299675e5a5de
z647da58f7117030e5bb832755df7cf499c73d7c510612ede65b39be76aa1ddf703a5778a5113ce
z1c81dd08064a4dc5c7e733c77b6c40f700c101d9601f7d2c4b24311050d5868e727ee27689e5a2
zc9d6a0f72c5dad0a3fded6f78a2d3ca237c38960899dec1ed3fa71c97202168c9ef92d487825d9
z2db279c7e8f3789474ad90a1afee36ad977514c6ea619b95f13d7dc44a145afb137c4337743308
z21bf37f6c2d549bfb08d3ffcf67c9e56ce4411d2ff47e04f7efb809a9055fc58250573f0d18b5d
z38252261b247fdbd9778ae107f8a20470284fea47055b942c4806c9d1a47a4a742ca6aa3f8f90d
ze7a12415d28dc4e16da59d83493fd0fb0bdbcd08c8cbf06059b0c1fbb634a2c76e018e7c42d615
z8131d9a85a18be75a5320145e05f88f55cd0bb8d86593a40de53da09aff38e17680c18b52cc136
z607b111028d7c5facab86199b48f3af4fc5202bbf813b379fbeb4b7f676cca6d90543423a24de3
z7ab326e45c82e2af5038475f70c45ab11d22ccf22e63eb645735671075e47f8c97a6349841030b
z925b1954b25dde7aad4fc1d6e2dddbc18e5c3174a2bf9a6dcede627778f0ca1716d7e2af63ca41
z5148c3d08382ee9d471d225d066489a81732d4698fbde92cf5cc32c27dc5f481d7cb72bbad9681
z0e763dc25307bb75e4d4c0272953ae5cf9e53e3f71e61c6401ade65f34ef2d98b3b954ce1dba3a
z5e58fe9bb601e2d241c2a9433583e53add477f3cf0c68916e41a6cd8b918b019f8c8e8cdfae26b
z6cb17b2c9628a672ecf8bb6e310668bada95a8947e90017504ccf3fbf110035eddce6359884a87
za9ecb2166ebf7d94ff1ab41c6e6e1daff9bc4ef8f838a278fc179e0725f2bd780ebe30b76dc413
z36c821171b83c0831dbce780c34f70978cca70776eee76bed0c2d7277744f0b056cc17907e8d82
z9fc93cf57e4b383a0cd03f63fee259a500800bd6ed00cd11c5dd2b796b4ce6e57c34ce7dc574e0
z2aedfc386035daa9d9bf504df2d7e154b021e9377ee1bef76aea26b955d552c769655d6d27844a
za55613a5913e3b1d9d9b66c65a5de80321291362fc94d49b4fe59bb5f4d8db9dc5be45bc73deb0
z987fd146e3ebdf3e8486bf45605ee2d208318780ba9ebbb361fe0e48ce0ec170a631bd04384f46
z47d5a789c5a5d4e457bb137169ceda39da6bad1116d8f74c3041f0acb3d48dbadcb98633ecdc3e
z4092f6de3703527b003c0773398caf77f38514aea8ff147b6c35b545de01d1547fac17cd6db3d5
zb4646dcbb7e59f2128b7f8ff17bb0cbfd4e97a8d1030d34c548b06ef49ca13f0f167f1fda0a6de
zaf7bb5b85587886122c8841fa3bf21ecf1a85f9697684e1e41d65e5e43c35dc6de3f6a266bdfc9
zb8ee76561e5e45f2aacd36f7d55b59baeb3e0b173f77f79a86daf63817d914a8266e41c793254e
z72ce63195d786d8eb4538f635e8bd3125730115c23630aa83356a6bb9564f430252c363d01ef2b
zc8142cb9b97321a54cd560b2d01ee72fbaf2889e14ab057f5d71c4826c20338e1970484a8c167e
z97247451ecd97c9087ed4b68c0bd5ec409ca8166dd37c615152b4fe2673195161aad7c463d4bd6
z28b5c2efc1cb27128c76df2f12c5401e2d61a1a645ac4b92b15f9fb996d722f5be85e28954b9fa
zdf70725ab78df9453ee4a5a77965e879f0ea977e63245e48a305c41978a686b66d036fa20eb14e
z3bcac7d8c630f67978357ebcfdfabc00a6deac31dc144ba0d95c0f4a454aa1e2c4740412096737
z32b4fdb989ac4039284393d0e5552061ae932e38a702976d77b63a0963e6ae491b87c0f6de56bc
zd5a23237f9f427c14e2c0e835825108c74a0af78ab9ad3acad73b1e21a116b7f98f6533ca29b5b
z9e0b9f7d57fdf34d97d12f6f428ec7d7d6b46faa6dc71ab263b16864927b43cf0de90a1b38e223
zd10e2756a4aa9a35627d31895aef813138c583bcab7dca2080f0acd4ccf68b7271744abf19a646
z9a1d6687d633fbfcf074c26e8c8a29554f2a0567c86f52661aa8522dbf7a5eec87693d9c4b0285
z4be9b29e32e49f299a0772d026ea9a0718ec838d817b48d05aa03173c39426483ae080ea5e9ebe
zae6123d013ccd6c57731f773cae4c5759a2c553fe786c16c96c8556452a23ae4b011ff684856f2
z210a65bf2176baf79bdc0ad316f29b4d1dda01b584171ac3a6550493fb5b68156249d01629abb5
zc4c4fcfaad3b4d0e92c1149a8abd43f7ed92d20510e163b36f25a23227286f4052a4d6e9933fbf
zcd72c373f6495675cb3a924c5b7b64a6efd5c3c6a181dfb22e68f5075c6eb80be60e277556794f
z5b77e9ba2a7e2f68e8fc118d049691ec939151e3868aaff8a6ac9133b13515c844ad8b61d7ac0d
zbdc9c988911a2aa1c72c1103bbe7cc6ad0e4e2cab36113c5fda82be320c469df15dd77029fb0f7
z645b36f7b1cffc7a1721890bb319b2830f2a3a9d2c733ebbd0e58a62e36ea69f04c41de2cf0ac2
z9d4193f109c2a73533f4b37de0ea5d24d0c1bb31e0ab5ddc117db1f8046cebdc8305929fb255a7
z2f32ddb67371fcc9a8b2a2b6c1d3b11ba474b85df60d8bd99299d32d9bdb19a5c1a0e373349e4a
zdef3b3d29107a3ab1dd116a0de6142a51cf6e4d011f0b99a7b937d7f7bf8b58fa0e0d89a8c31d8
zf40816642d4c7cb498022f7ac7851342c931caaa5306eead9b21a0b974f7b1f9139e2e575d5198
z351beb50f12a04cf26f1c586a98cba4c37524a60ccdd644201891508ed9ba4d7152a44f2a665ab
zb1b44ebddbebe59891fffe27123b7a9a4a52eb97d92d48a8cab76034e3f3e0b8984400ed383f66
z217879e4968a15f04260cf3d768a638c90c7bf5a3c8142c8d085b1622cce190f78f92c3b5ab40d
zc0f6e14abf4574a19cc2b6ef59a70bd8aa2b7e2dafc4d0d65df117b4b45035068643ccea74467d
zda7f094ca590a075693706a13c50f8f47d85cbfe2bd3bc4bcb90e5bd836f70620d6d2e46e6cd21
zfac08438fae6146d6a0ee83a9cacb0c9919b98881ea2b82851f3dc26776216b3af50afc9c6a117
zb9cda91e8df261e5bb36fe95a247daddeedae11dbd51e4b153da7c4f1f91b933e11fbc2cfe6e82
z23b384bc889f9a73a188e2c1ab218d274fffffb58b8920a52537b0675324f466d424d49395c4e4
z3a6ff66fdb06dc9ca3e579af589aeeda1bc5753f2737d95336a699373cb065abc0916790f69727
z322b5b9fe0ad54226c3d813be2f247f8f868077e7011ee88f7975f4042c6846efab9fd1111c66e
zcf69dc069c091c1123862cb194f0858f7dc1413889b784616204e9df60cea316d0af6bea5809c8
z1184b4083744e8fcf27bc5ec5c4006b646e33dbf2451df3ac47c74d8b9d74c499d7029d2758cda
z4e395be44db03f79e0c83e5dd806b975a02345642472bdc9de3e8f1654b227449b1c90e2923fda
z9a4ab7069157d13d6836f8ea2a7aff444f83a281ef09add2a6a8471a6b0143c9c3e1ce4eeec2bb
zbae2448b5dc5d7b6a8af7da5dd18d574adc794d68fe7eaad8e0f7a6a19d178f7f84198039385d3
z4c1b24cdea1334928eeb9e68520da018dfbd28f0400a3a6a649f168a65d232e5648214e9ce7982
z27f14b8946c99ee4986b107df369754991170ec5f48e0c68d877ac3ca0d42e549a30c86a6725d0
z0dd27cdeffbfd868e9392c15c9f7ad13365e619d9bfe557b1bda32cdfb27bffa2f95a9f45841a7
zb4cc2b0b66809a41c0841edca281a44f4c6a1e0dae6016cac06293eba09c7e99acc0c734c17991
zb855fc1d7236917842e2f5e8b9b1c87b1deddbe249d8272d7582d4111233459112ddbfd9391182
z39539185a2b1d918d12dba7ec9a2607754415fadeb066e0d6bc5d6883314774a8c702d5ce58865
z62bd9e96274405662d63b2c5dfb1b0f36d8ede8c0db46a3e0e40c280d0f005abc785a9b4d3d3c4
z3398f88c9348fb85c1a4f14ed13bb21bf50b4ff3f42de1177645b135c882a31f799c597fd6140c
z729beb44c15b8e3134277d29c805a7c114427078969878efbc6207eda7fabf40f2d5da6662a351
z5effc6a676e5633bb755bed52079a4187cd4d90c4b7fa128f21cbba6133313a34eaa5347a82325
z144a9c2f774eb3948b715f20528210d0c9c38036c9faa19b9ba7dc2b651ba82b4c458e15a69103
z22c0e377bf7ad130882107d6b9d224a9ac509f22c292e3df77d0707132f26a36270631cf586b7d
za834598b607037dff8080d911fd787e4507c01d0c2f5d1a02dcd3cd74d8725a2880e7c2ddb420a
zec4453506a16395fa8ef28972cf8385d06befeb2660c8a2e00d6dd833dc218cdecdbddf8505c04
zff54bb403fd37b690df30502637e66ebba20018584bf434827af2aaee53002ede4c48cdb37e420
z5987b72c25951c3fbaa34da49a3da12702b1bfb27a35eb4514333a965353ba01100607e75ddf2f
z92294210986f1568ecf3ca3a291f3e3ea749f085bdd4f89499e90eaecb2a9fa37bb1bc2ee4dca5
z272510a18b4ef31fbbf2e8c26769e0157ad1ac44845d1523235e9b15c8a08acf1e096c31826a48
z9b640d7ff9082b2847a4a394edc770225b65bc89825291ec19b643472824a9306d7a7d4ccbcb4d
z9e69e2de40081854a648e76a420fe74ec592d95a8cdace850f22c243f976de5c09f9d630d82dfd
zf552a8fabb841536a692677faafcfd67eea5a5535ceda1b70f776c4cd88c3ad4c3bbb2452a22f5
z4e57be3e97eda066050238ba667b9530231e7fb8e7a85de4966c3b422c2b3fff2c41451e1dc9b6
zcfb1c9c99dfa3f78564e96d7fca82f7b219dc9eeff7fd9feb2f078e99446602d78e9a5fa0b52e4
ze8399ba0a614622c7ba2150b609516f6154485bd85d998929ff36a4816528ba778d3b282c2e980
z1f649485f4592365cc659c60f13d1478a20e0adc115347c5ca4eb24168da4a7221adab57e4e910
z180b35fad0a294966490f32fd53d8860752ad2462b01697d952a5d525e0cb955e87a207366bcff
z712ea622f58a17e1dc9f371e8b0ba20b9d90d6b9d4cd74270584af60496dbb0270cccb7bddf5b2
z74cbeaae8832951fe5b5ae87963bf07c5d2dc1be0b79485226298b14bf2085f9871eb0f2bd7a08
zba5684772b481eef458acbbea425b7fe8e07a2e1784709594244f473b3215a529457e786b82718
z993584103c00e2c6073c921fd7c389bcb2bc3165a546c28164fdceae930c2d0dc7b8c956bd88f0
z657477dd9fa5f15fa1af4bbf49cb00dbe088ecf5b9d702dc213225f71afc8372a166b00567aab2
z5f25eca3838e0a6c390970c435dc1d3745f899b88b7a8bbea46d6f75a92a133f674c7dbc046c8d
z8497525469111649d18e7b2987f5af68c466d56ed0e3deb11a96fdeb7ecea90f56c49cd0ff8eb8
z74f3dd5f229ef06da5ee37a2132eb3759597b601e909cea8c958065725b214134ced9da31463a7
zd1c284d5beb2c0b5d1f0b436e94e7ff9ab846ca2ba364e0876c80341c40eaedf74c0a6cbeff0b3
za6d14295e767db7f1ef46d79272e0351e3f4ef471a27aaa71a4e35927c5062631f8bcccab675ba
z66202ea3d971e25c65d15ab473f170c00c4de953bcb8b85bfcbe8d695e454c3c765dc780cd3d9b
z34ef0150c0b90496d6a4e8c7f6cbbea92176985289c4c3655f8a63df1a905a23cf5e77c4aba8c6
z65c3fc2e31712bb8a7b67a348839df91bf07821d6ccad985cf0bd39c7c4820eeeb56851973fdf1
z6401a660002535008ed2bfeb2696e4bc39a8822c5de9af2e010b97ac0438e1efedb7e4c67c372e
z81fe3f532aaa2be4027d35c29b4d450b4aa8f72c5e2790d4904234ca0727dbd1ab32f21fc3f631
z0f33622af352338edc247a44d37da4c0715f97e835dc3d82ba979abd5dc67e451d20348c8727a7
z926f1c22742903d551ab1eba9846bbb089421e21f57613e7f202783defddebded8c4d97e9bdda9
zf3297225ca5d03dc123e580ee422207fa6f5ba6b72fd3a35ebff9d3f5d5809166d2b354f60f5d7
z97a4d553230c4eaf17b185bb0d723f04e89b392e2d78b0852401e46ae2c98cc465e9abc1159222
zc24e20cf98de004511f457aa817026d29aa409410a2668d447d5d234a64cdd00ed1469dddbaeed
zbd1aff872769f0176b7056788ec6bdbcbed409b04875c023ca0bd957c384a5ad8dc914c396a5a1
z3e8185733e5e6812c9eab7a6b0a04ccc335803fb1f9b50867decec8d5a8afc3479b7dcb47a7226
z3190197676260b35a84dc2cd034fc0fc0e407bac2aab10f341b48836b1559f40a78ad09fe12101
z3153a1848906c901ced49d4ab95fadcaaea36e80353c0e1ee866d4c4bcc0a2e549e9960a92a773
z9a676cbdca1254303b5e4ef5af48adf2bc6132cbe27cc4adfa4b946573d3fe223f6583e82a88e6
z3ec2ef467d6ed0622f65b15a11aeee1816261bf6aa10fe3342a4bc83fecddfcf2ede9c2befabb8
z85d27362160f2576965f24bcc12d8d453659471573c928a8bcebdaa522637d699f63816b549453
z534f76fd8531d0d6b08c2888be3062e3f93ee5bfda18ae910836b4ad698a1f7d6fae3adee6a04b
z6c2593e39fd13701d4e335a2df9934afa6b5f924634970cef4892ff57b3bc4f782611e92ba7b9a
z2371d07d113982a25bd26fa3337e59489befad6ca4424a7b2f9825e2def249679d55a4feb94ecb
z4b6185431b95e12ad986a5dfde4cf45c1ed8c6c08a9c914a1bd5740614e66bd1e6313f9b4b6488
z75485a23fb1b294e8098fd259d69985e2c7de19c1b6798570e844785ab5afba13ab20703620df1
z49ae6387e56c2a0c40f96c32c029bd723662ab3626c007393b16519259f37d32c54ce74a7e3441
zc2696ef2da88f4b807ef233970dc71d064bec741a56878f1158d35153bc250ed396c004a62632f
z1f71543fa04773efd0d45aa46c1553c7b15af397197e7fe09cda23d83b0b0564c4007c26cb0250
z5afd652c151aba4880100aa5a98e2a5e8ecd03206984d7a06eb809fbecc4b90d006a6a0095dc39
zce2cd81b27fd2875f4641d143f41359ffc0fedd18f241aff021d75fb7348e6f636e49318d3749c
z9a6dca9042fd4e9a433b2d7038616d14f1fd4f824fa53805b32f6b55f94854ed7765a1dd631c72
z07126e21559accdf11b417767b23febe52baa90033ae64180efca1c49dca2cc2c0227e3c733365
z81968787a1ff4486662703d4cd582488e2c8faa5e8da29e765f54b064b6f875e0b365b3c5f02be
z52d03e8f4b135a01a55ffc3e64efd2fb158d67f125993fe30741677daad1134ec780520a70282b
z9abc3c78fa976f569d61f660a2c845ecbe843262cf73301c476f34ac39e7e63bcc15dbc8314b2c
z53f3cb8a956dae80d078dee198f70ce581e771fff3310853122d27796245178db5f3b93ec1a745
ze5ea7999eb948be1746a04bccb57e19d43ee34eed35f1b3a2abafb134f03158c212d4ca1a2568c
z5eaa3ce88dc9e079d7d218aad7054a9969a5b63ef9d55569a2db233b049f2a76420b98e2c0d2e1
zfec3b0e7ba9b7cb61316e07f1abf82ca4742deba0597845707f9d16e9d232cec572a935b2d7d8f
z768bbea6e401fddbe13a72ec809bd7014c7baf2d79038dc04dafef35dc739e5d25ed92d6f7d1c9
z27e69233754b2fdbd9ff9d200276b35e6bbbfe1fbf5935cd41e1834278b70ffd7e100ebd39ebdd
zcc8f3b9b4da49e998f56773828767af3fbe6a8d0a2d313544c12964714a661cea7f34790227fca
z9ee52cdc2ffc6cb2fd072afca3d390f41e9798c102f4fa9348f4353997f9e20ac91b6fa458e4cb
z78da4bcaab55a031cd3b7fe7d274b34f929ddb3ec729e8ff5924c16b04d8badff072d0ce603a9b
z2345134177346da0aa8daaf7a2b8e9e09dc4616c9e319c55ba8b19c33feafdc66aadfef2252b60
z5c2ca9c5f7d06fbc1523e7421cacdeb825386f683cdc5d4ecf3249176ddfc8dac5549faf47355c
z3036fb9b05e850c7f7a530557d7a3f4d82fc987a396e640a218750ad3d4ca727eec681d1f188f9
zad6711e6c6fdfadfea7e7748b38537d5b0fb462b03d51e745b00fec09e8b1a1df572f0ee70bc63
zb3b589c6dd470a5fcd8f548535a5548ce613d217604e8d77546c9e4c864014110253c4008f4332
z9cc5a144948e9df64f3ce236f666f670e5fab00b6444f1a3f6b09395e0870151c6e6e08fd439a1
z3885519c639e7f5e0bf5a80f0ac2742b3291e2ea58583c71fe82afbc3166bad9299fc954e9f427
z686524c21c3e203f88f5d28a04e93443fa2352c1236f9e44d8e7c34d4808331cc013c7e49891ff
z009026aed57f4b6dd8a7744680d69cb0d7499a7848537d1466a45394daad123964ce2fb5a5a32c
zb279f1779d1ffaeb3a5829380d24f3e6e48f3546551539a66fcd7ebc3386e89de4de2a6abeb953
zbdd9e1e6f7a0bfe971b52dda1c9a702930ab33c5f814c9ae75f6b5e111e5c9e3207fea11b43c3c
zae3e3d7ccd4dad4b10cd5f4f71bd9ffe6f142e3219bb1da0ac6f4f4bc24b0c8d300be4a705d360
z39df0e5c1ae9f2a1fdececb3c2bf097139084ab148856afbbb2b10f6d297c551defe0f7a0f4e84
z4069dbe7b2aa6cf7b2c59b9b1326f0b46cbc3a37125859984113210391fd44f916c04bf0acab09
zbe8d7ac3f55db1b6cd08a6a1d73e9f3bbdb72f55d1a4c85512cdcc9b9e5d0996c8d94bef1f506f
z745743190ffed5b6f4013de4938902101f0c8e121b965e1e44cff3032c289f3195e6495a58bd03
z42d5296f25cd66797348a5cb18d27314f10e54808cc5ef84984b7fbca9bf417501c0594d49c377
z683fb07d05447f3bd8a7357f15bfb6e781914532ff594c9fa2ecdaede04ae51e116bec3efa547e
z9c6c7146bf0b7b75bf21d46dc608c43a775d52c527e62dadcc64f6d28dc8db732aec11459ab8e0
z1ffced400befa975454e9bc756735ae0974a513afedf33e302eacfc0870df29cccd2b892857efa
z3e9fc0d04b23c295f2e3e12992090312264f12d16e28476d1ee0fbb185a1cc333b557d376c6422
zd47d0a9383db97eaea3c101eb4ba4298de460d6c9efab4b36f0c196cd8c6f933a8b5cd40da1e67
za4dc2e187ef739b045c253b80757806c7a0bbf7c47a82e4a74ec06888e8a54d22098228bc8c4a3
z603953b98cb288b1876c5cdb6fc63f1ad3b1632aaae1fbac5983640dc5d16ada0114e4203d5511
ze7eb8f8476e87b6a42d10a44f17c95f45c82f5da50b4a3ee2ce4a9ef4b5383e981e909ff8ec905
z8a75af34708473f56d46d89ac386ae0c6a426488bd62410e39996de65d367e8767a914ecf9f35e
ze3a0e6c123ab368a831cdea608320729c62112d394c94f38a99e4e4085bbbd37ce2b84a9196269
z7a814111fa8b89bc19d6198edbab115398db5a5a0c3de8e1507f2db59c2a6c168b503b665ff108
z68e8f35dad99c2d55eeb95065bfe63f97818f99e8f6f8efc3c1325cc29a4a38e8f392e1078f98e
z2c9ea8b1728f7fb4314dce706e5a3911918f82f91c4be54e16bc3311254fd4df2b1c9c538754b3
z38b011b295c05e705e2c70e5d03b83927593ee2650871294c17f9b29386e09872c06ed5b30b94a
z070cae893075c53352f8d29aa1b43cabc98a178d4b3046c65d91cdc4e0c5424a93a72d20c14ee1
zd60e548f4b09bae5afc7817010ee313b0cdfb8ff2de439f34f8068e3953747bc851d7be627e4
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_resource_share_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
