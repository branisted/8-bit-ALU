`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab30857016fc53a
za25afc8341302f0c829d94450c399b8ff9b0386c187cb854ee330605b7b59da379b1f26f488e1d
z36e675f0b1336408b3a1ad87d0723054f952fbefc8d5a33eaca6ef5be8f42bc59870a29a5cc9dd
z4fec09ce6e44cac279651402e7e1f590df88ce49ec26ab39f12b4a02855703c6f03b1e85c797d7
za357087d98e5b1f45502e45892e5823d6fa4b762932009620038c05d74efcea7c3fdb38901d620
z36515d0824367e48d1bc182335f158c262d396cada6b0ad58add4f945eee634c2dceadbfb5118e
z14969c29a743830a07124bfa78707f3952b96b0db7af7c9ff36f77137d8c490c4f79328328069e
zd7d5280e4f95742c9841340368b9764f0f80413adb175ecfbdf3c40716abca7b8cef6f7fe92ab9
z6bd2453f1aef7f7899c5365c5c83793cacc7795c269413f6cf0dabad14d40e9285afde8c01a47e
zb61893788ec5060288cabde8fb553f21b02eac61ab0b48ad3d54f4d1d76508b22f0c600861b5ce
zcb30ba708be817b1f50f59c0f6fce449203e7355c1be55b662fef3f92ba58243d81537761af8d6
ze27d7864d2dae99372b2b75bacdc0437a4f7e011d68c3487a89759e3625548fcc920ad06471ee7
z2d701aabf726859343208b0a543c73eeff8406febf277e3babff437ec820fb49d6b78e73bc2353
z884917487d35a6cd06d7d73ccff5f05355122888b886d178a03d8eac5505df521c14d1e332b234
z86bc1de9891c0fe4654d9d65be6ba17e0f35eaa0e5fb8d4ffce747c7530d86192c5a60f63648d8
zec2b11ca4783a37281db3c8b2556885556aafa013f24449e0a06d5242cb51399b3e756b814a7f7
z7d2f3363d024adf895ee1f4c57fb3048cf14f737f4f7878d0d0c6b48a3aeecf0d16f61ec999e70
z8673047544b470019ece6d4e6f8a1469b42dc3022d4e7bf3ec62c2af4cfb08f5a5de608628cf8d
zd4665dcc3f4867d0a07a836531edfba94cdad9d90730ba8b6b2364b0eba1514c0246e78124c617
zf6a26bec02cd6601f40650424a431a340361b2120bfaaaee24cdba68de41a962bafca77ee84e80
za2da1ab25b494bec121443cfa771b7300360491417b42658f3967a20c16d3ac0978600bf5db91e
ze42f8327318524a1e54cc36e7ad8520c8c816f80b84c9f01401149c4b5521b29874dcedcb6a724
z7fd67ae188c4951240c65cc56706fe40e0268bd1d996a7edd1a6f87c2cdc6dbc2e615cc516ee36
zac5315a8388a32eb11c9ea78e632f2a835aef1e16a2a705f424dccdf3601eb5f07309e509da0b3
zbbe6cc0aee2849f266708e5861c30c79ecef15362c54a3e708353db6c2b2ef1b24f45a63a43aaf
za90283c32ed5a72bfdce92fc6d189150adf8720a1a7d97e1ddac45b8361b1eddf0e5895b0553d3
z2cfe4cefe1e1a9997fab3a4cdde9ebc6cc5e1bad261c3f438cb0e4b3ac99ddf99c5a72cc0c5c77
z8e596eb486b16b4c6080bd445cd4a251e0079c5e671a0daf28419fb0b7f996c90c507c6b1f922a
zf71b9f59cdeeef8aab6a169d18c5d6972620835ed1834b9e34bd757c1558ac2c7a222ee09bdb27
z54c85265881871f595d15691f2aa22b04de86718328653f1d7e9d7f922a4b9d6ab7f41a385be6e
z201aa0fb774dcdb78679f19502a8057f04e4fe6c77fdd27fcefaae4cf170cece7121c46aa6e6e4
z0e6cf968d7e83dafebbbbe893eef1b3f6555127ab3767f5e6df40b77fea38a2420b84317d8893c
z1b6d1ca3200a3272d949e962e96344dcf53e0d318f5685677438aea318a0576a6a96376c8df389
zd0a3d20a92358e9ad983dfc5724d61325c8ad8f92f7a8369b166e91b4f5d0c5d5ed15067dd8145
z6ec7bc23fc6b2f8ad20ee7542418498406713e9812b09b5c221175e1a0fc4368a36ef39ce4dcd0
zd6d98be3bf9a00ec7a2630f3f79b342cadf5adaf9a3428fbd3c4567f8a9d76fe188b65deba1cdc
zaa3274f33eee21c5f670f78147abcc1f92327dace8b7f56bf10926354c5a5709fb74c67396d147
z0566fe7b4aaa43b897fd2a793fed0cb228b139c3bdbf0104f6d97eaf0b0063374c879301d852d8
zaaa7356b3265d23bccd048520984b6966689b456768bc63fe39dac67887fa130eed2c19f3ce40b
z6a31ebd5b524614c6a025da7c751dbb0c44ceb414d069159135370ed35f9622dda34cb9c348402
z01b77eb06a07fd059c718b172cabe308f578c0ffab681ec25d8b3b8deae69c9f30b97b855267db
z410268a0d09249ecf808a1aef06fe08789947accf8000117e71f73b0d8a33a9d757963c04cae47
z9f19f47b04118250e430f00edfccef8a21d482b0dfaf0662bcad8a7d274c33f1a5b97819820838
z74637844a9ddc2458629d17a7e93f95317aa2bce32797267e9b921dc811b4ce648d6c7bc75b34d
zef145782141d4a331dcddcdcec5aa1397a399cc68ac92056fb2cad099669ecd6a7a7bc0a4d9d31
z3dd28029299e461057fcad11fa8525593adab12b45156e7f92128b864d0c29b5d3746bd76fc80f
zc3c25dced899d07a2c588b706efd9f0542975f7dc6be061aa65ed19c4e47cbc0d2b88fb3dc01df
z589c0c35c40465228ed58234751a3d4c9d569ed666622f09ba81379c68cf33d877641f1bf0afd9
zb5e040cbf7ad2027e155db8f83e4cc7edd960c35b2b04e686a53fea9c347bd8bbedd4f3fc3c73d
z618a94b65084d6fbe031acf78bf77d9f56253705107048b5d988347ad21fb2b1905343a0bf873f
z479a1c3dc7afa86772acdfc2831ace52b57c024bbbe418f55e55be3e2eb9b029f67b48f0a69193
z24e0665041890f7e6980d3902427b0bf3ed43080f88568973d447b86a2cbbe51c7439b38850fba
zbf66587f1c6b36e1dd33d36c792d5abddf1f7a02fa77313909acf62068f2c760d2a988b1b7b629
zf937c51949ddea87ef260c377301302436e153a5da35670897fb401efb02a8911626f41c788e90
zd807c42baf8c119df131d451256af69351b31a80584aab2ab4bb569c5007e0929f2329fac8ca9a
z582fe4bc95d063b8bb92108f7f2ae13c22b00443458ecf7834f281e00886c5d6ca113aaadff16e
zd33e7b8160935eed20ece5645c51ab499c3ca530f235f227a52e90df28c8e56a7ec606d0e25275
zbdf4973fdeaf686b126ca27dd9725fcaf18a8e71b14342858c829efeb79fececd6cb0882191baf
za73f2e269c119aa34081b5d2bcc4bade06b7d18bfb243a288b199fa1a7a0be5431103f091b3aa2
z2f943cecbc1d5eec745d4fb3ffbe528590e5d857c45d1ddcc39954395ae6e7ca19f2f77280cd23
zc1d9d9695b0ba8d560393eb1e21b37eb8331c4aebd2cad19b09c1845cda5d213c37edc1d2809ad
zfba405c74419a841674ea730f5031da5f484b723c459d7199a2ae67ee986b6d4e4ab7a9924b372
zdb8a6c6ed8c9b52ef1968c3352a537e341f624cb71e951ea7b525380a3f60c1ce9b50533aadc80
z17b3200690ca2b8b00136277f9709d882eabf77c1679e01976fd326aa47bc93927f3ea2b01c1cb
ze71862ab77786bb17bffbb9aee62d2e5bc2f6d3edc5cb6bb3dbb5e0e6197859fab68209faa1822
z65b396ac0e9819a2033e7ea1c3ed376a6ef6a048ebde2e91aadf6b53f0b5206170bde7b68b799a
z6bfa3b06922689c49fe123d03f45813c4084101c087d0bb9d35c86fe25316324c710c8a8b44bfd
z65df9b85376c5a825174c1485e02c5d8a1d0959450b02b590cf8efc4a3cdd58aff888f9a3354dd
zd2c815880885da00968490f6e2da0cc61147e2751a6e5c0f4c828f2a996ae4966a1d8a13ad50dc
z00b04bd470030150b84a6dea3ca3a2c248dd8916d590417a2624fcf59743051db75f9f8ac8de1c
z831456911b2621fe30402c2d2791b732f4d215b41657e8e972d06bd9c99f634f7acc0468176db4
z41bced1f052feaf8140bf7f628203da75e3b8c19780da1a81c3d423da0693e47805a392a547a10
za6abcd25267d3eec6232c2097ef3017393510faabcc38dd3fd94b96763d7fe8a6bb71b1bd6eedd
z30ddac7e695936ace769d2077bf5dcd62244575ee55e6bd74907bc4b4129a292d7ff069a05b7f1
ze63727fc94537ed6593caeac48a8d6d84d1516129af0196b4fb8e3fdb79a0a88af4e06be2e1b71
z041a4e652e19f23273ac94a254621d8f4f5c97d2169279df3012a5e47bf2187d8811aa45ed29cf
z74f9fb280e16b21f2a88f15868875d339ca392e5514297ff05df1a5b6cf5022c0dda1a1a4626cd
zdab264ee09479c1fa470d42bf121e2f8e4024162c7c2249672fbfe201bf8f5a47800b7da6fc98e
zaf99841e63433f513c48d2439635195cd5ed20a792c41abced5e19a4b3bd99a5f5ff97749dac82
zc862ab85f22b54a3e06d85b67808dfa4e1168d9f92330d4008c74f0aed2c55429fe9d8169b8541
z76ac07a02c0049f9ea6fd7a113441560cac89f7edddc16930a1d70a448ed95bb63e05ebe7a0f0b
z0bc4ae75588354bf893419bf85b78f59e5f606bf4c651569f09875c133430c5149e3a5d4a88430
z4b37f5ca8f9c3b9011a912ada04dd30b0d0ae29fc31eff572f34d125137cc233693465c143f9d6
zddf1807027811f82fa99af4c4288332f63d8447f4dbab4279af5fd4ff24e7207c97c961874b2d1
z665eb0befa931d0e09ec3840d39852bac0b4644ff8cd3f4eaf381124c0ac46465b971356543660
zc397d39e034ab482d153270f5c7ae1ff9639fff1024313c74e4d7c0d9395c1d23d982da4b4cd8e
z22be0fa798b8838c9d6f0df23cfa3750771eefc563ea38e225b5bc013f6d37607af6125c379938
z1be23f6587041bf3cdeaad17264bc0d4d722023a25c7c21dedfb79b1440a3e08726eb95828f7e6
zfb385e4502fd86ee604f5a73de24cd8e01650b3d621fc4953ea14e129ccb3f6198f3a33d9a0f8d
z7805c93077c6676f4a24109cfb12f6ca60c1c47d95a16fab83887036175cd63ca97b6d8dd61862
z8528be494127a127d755872e9f3154ad0d29a17fff5242d6b856bf6f0e7055e2a14052ef533e31
z09d44f27e31dc4cce0bb4c2ed9a905eb59122222528b92de711284e933d4a836e38ef19338f098
z2438f29d0b73fa53bf507047d2067261443e53ffe41841d3bd7e91c1de90a48266ccb8c50e7319
zc9120c38852fd6c652c8af68fedb9a9706824e485eff3b36635a455cb0c7538a124fec8d4c004c
zc5a1ea7aa7b25fa41cb2537932ceee53af5eb9fa7e331759c441bafb0e05cd39f92f7cae14539e
z1233b6f35d38e0d4547555a6b55fba1eb3315de296093fe28f3962dd75461769db7b068b81466e
z1054afae6b60bfabd314c0171387457f72dfd23d3516744c6c7062af45d86a5c69d18a0f0382f9
z6e7ff29b3df04d2c04778c616677196a7e883f89363b34f27d1b9028318f751b1955f76b5bf210
ze99aed355820eabe93ef67208e81ff408f48d96a4718bc7c3721be0f15b36a6e8b29f94bc9744c
zdfabe36cdcd868599a23666d661b9b4f415b3ac4a1e866d7dd11918eee319f621ec209fc73ca59
ze44b0316209a50f9faf2ed749cadcfb23a0f7c99a6ec424166dbb2d338a9702d0493a57ad0cb8b
zd0b86c53bcaacb6000478cda928c8c6e49be933eb4723f9df39962d3843abd2c464fdff9c1b942
z076c70ae4358ef018a7d432e19882d6d7e9076e7fb804f93892e7c261768b58abadd65f608e29a
z63b5430472fac92ba0220b15c5254cbcbdc3f3b6017784f47d4dff07c64dd0aa9394af007b6a68
z6f87eee3b197d8ef2e1f494c79936dd809312ac819dac92941aff8d3ea2c35291b1752fa503095
z76dc877c684dfbe77b8fc3e743374b189796dd71f47f8d5e7d1bb3a74ae71e0db15f2c20495e02
z6edcd28b1dd7b538aa32100d650bfc28f8981ee2d073ad4a7f4469310b337186686dc0c1c3c068
z4e27df3008d24bbb7e361f487508b7ffd22e016b3abc01c89a9d8f949de7e62991c13044b1d672
z3192af91393376345d72ef413f9f4787ef3a98f4f515cf48e5b047ba97bd6ccb9bec234180c64d
z5f2fcdaa6a9e5c90158d40c4d1ef5dff7a8d0e13bbdc5e2475cf542c1566c92c91893dbca1d3ef
za14aeb8fa6359d89290e6dc41d88e4b866d13c0a46d885af7fdb69d3b7419f8659c39d7fa6d68a
z8d086ab44dcacb6b70c8f60075674556b2fa750519afdb442b510c5ef4ccf851505ce1c792bb55
zc7d5099c4820b2fbc349f911d82f6c6f5089a374779389be3f3097658acaf223b6513fc08e64a9
z7908378dad7469f53dd24d49bb8ba05e0b0ed4dfe3ac06a736d4ed6af28553beeab0a1a16c3b24
z19a4f6cee5a93cc420138ba1e91e3a53ea858e9419ff2a733a28c740887e0ae255cfa79eb69424
zf30c12de9afc85018a61a2e6c745cafc68f3415581407fb34f374a19ecb7ce2ef0d81e66306f84
zc3abb6252642d954be5a8401fee88684269d3e06df33d0e8fe39b535da9bffa1fcd66103db710d
z63754314c26dc84439290fda0ae78654294d46883c44570aa745c1f7abd775e5c5a95f5c7732f1
z2d2445b8bf8bb7f37617fafea8f1068b7d3891ca6cb2dc7d1e0441644e57fd0bf28e8dcb51b878
z51a92f80e98df568853f27b6d6de2fc6b15dc1c7aff364ce77280e8d9e891c0b80332308057baf
z5e37adce44b5b55476c37268f51caaf671dae25b8efc28408c9fceafaa82a0d0d0deb85ba47373
z1e5c5515af50d026e0901bd816118b5250f753ef7a05bc007a2e6f66f07ff4791f43bd14ffb32b
z14e30668ac6aaae501cae47943936d7a6ae7c223b47b73f30720b0eeca1cc2df4b8503713dc86d
z78a63a261ba102c2a7813558acd26cbb1f8e7df00d55eb189b38964841256da77883bed6b1912d
z86af535beb7a145b5172cf07baf7b7d86e46561e39e4c59efcf658964b7f22b79dae8628e0adfa
ze7edfb551dd19e3782e28641625284ded0f7e6297b65a63bd297adeef8466a1b55ad7ecb482330
z16eda1d5e0cb20607678fb7de77679e680742c314bd9f12ac6aa773894c87135d519385acf8f69
z42ce3a8fb27c5aea6977bdcc5f99c02aca2058fe799962b777b664b559f6d1c04c36e42ff7c927
z9a6a4d755be9009173acc853898ab5712d792a5bf725943593e67415fc2ebc83789b117485c862
z99fcd1a50639108a5938bc1eb8a81914f2625e74030cf6436ccd660bc5f6114e82d7ea71c4a573
ze00c2b1ad4aff4618e12962917f37c8b034d11aaddc4561e0efe63c8f602cf6b830cc4d92f4ff5
z1651e9ee955eb0df70a9dac8cb0949ad391a118f9081009eacd883fd46b2a6d77c71f1632e0b4f
zf3e11a3a03ff0526ce87c3b359d5ecedf70b2511b0d71e86afbfd16dc2d5a425d4604becee82e9
z1bb26e5097545fdf11a9c8fd2fe41d4cb4cc4a88ec81cffa97ecf08b45036d03b69e4c33075b3d
zc40d8fcde9b06aee557c702f3d1773fab9d527e02160a713700bc1ab7345c851c944be356a46c8
z143ecf8bc35f2104f408ce4a5fbb274cd4cf770c3e43385cb0862426bb6b69faa2cebf8655f873
z60c9ff19ec735b465c9c9bab18cf36c4be904d417228550ebd47a71e25c5fefa4ecaffd7b1d646
z30da94f38668bff423f47c943eb3eb7d9359f925f37bc3f5ee8455999221ffe5fed3089f5b9475
z4d758bb9200d5b407260ab67447a580c05ffd2a795e5127d822d5fabefe996b644267bf2364aba
z1446576dda1fa0ef56c1288785925c1a02d794b908d273cf35bde8fd010c34bbcbbae571c795dd
zdd3603a7067b3b4b7c3c2e29ecc1367c91fccd0653ad6f7bbf80e8909a5f5ff573e2fff6c0671f
zc82a138ebf7b137b3263800aafee2fd6808d99549be973a6a63cdbecb80e2319196470857830da
zfce39b2ad9eae92ff1b0408aebc2ec194aafb2e05889668f5235b37bc549c2d85f4ec099da7504
zb987f7cac44956f69b2c267a6dc2641dcc7612735629d50d4b2f79a81ebd9da58e2a7b4bd35307
z0fec3380b36240e833322605b4231feaf269536b00f53364a79a356e10274d300c50593d5f8440
z6296be049b53eed49b40c71fc0524a5db66e39c09e16292b0162cad8a1ee46fe5c415f191dd084
z94756e1be8bf63476b3fa63ecb7fc9505ac681054c80159cb15afcda8d7bccf3084d806ce3777c
z59b509bb3e430eae667b3e08b457f109237e76ff5148856fbaedef3fae08b67c8a362c2517baf3
za832bab7a395880af127771f21f08b7f56deab72b5935bd3aec9bee171724ca85646957d773254
z98884cfe76000f2df3167cb60ec898abe7eafbfe7566c789c0efa539210da7b5a7561a87ac4be8
z439b22b0b667093ee80865a1708084029b5e9b7787277149b423521e982d2d397faebfa85db76e
zcda21f7af624600817c3c194581545e5caac593c531ec4503d11d2b140308b0f1dd4a5f1fcf61b
z41a203b421d867e98e3904fdd20b4c729bf088bb5768f4db0edbe129d1ae7eb7c42236b6edda20
zb6b55088c07e805cacced2440e7e27eaae46c107df985006959066d252bcf3dfe25de8cc138cd3
z047bbf75dab6dc51f76c766203ed9b7c2b6479c1d7016a81e23abf9a98e21bc7c421a6bf40b5da
z0db22c76c8fba56bf03bcf795fa947eeaf9da76eb56e0d1f059c5f3dd6e51503f24e2f277a2e6c
z36d8c5288cb34a7a82f872ab29d6f3a45bfe2b4feed3eb4aec9b2f0425942ff9f3c0c3bba7107c
z61f2866e72e2a11894b114d372548ff6a433b70aaf9d581f52aead36b985293f5134216af1303d
zf4119cdaf0e128b42f48f7b212721cb69220096a58bb9e975a9e3904b0ed059dd9e483dd06f274
ze687fcc87161c250d83cdc585051905357a9d4ec08d1065eac048a2b631d936e432279490be63a
zb24f54865ccc4e6b32eec9deca1ab9953d388c03b970a42772532736226431f7ca1ef256057d6c
z6c5fdc88609d561cc980e38fc1e76ef01d0eaed20e68d235549181518605c013564be5a567f7a9
z7bbbc33a3c024d39434f79294adf85b5e7c418498d31e0a9974a2911e9f2309d7f2ec66350fd54
zd4d1a05924fbd07fca95c36ef8ce08c9462c0d51da193e427727667acbefc6134617fecd9243ba
z36e887a95bed484a9c945a403918950ef9aa06398071bf24a818551f819b5d154f39f161de5a37
z2b37dee394c230e821ed08852e62bb49bae3f5c24bcdef4ed7e644b407fe9cb82e260ebf7bf2de
za1676f2469e6e914abd9bb718e2bca4d9bbed33c0b2dbe41e2bd7d8472ff65d1f050fe74dd9fc8
zba34e54ca62aec28690e24ab16c599188e7a511016f23bdd2ff3bcadc3048ccd195f659062611f
zee5c07d18331bcbb19f0d1a9d471b58c75149590d0c0ca75820c4d5b1cd508782bd3be854e48e1
z31b1386b4631a109d037364ef13264035af5a796e457afbdddd1a9922e029f97ab7da3dd8d590e
zae60f62a20cbe33ac77cd1215a9540bc5e08406b644eb2fabb34e0375a2f16df522c42e3fed421
zb1a60411af2e15bdef557ac73226d2f5941f4305085c273d8b442316d5a5ef2aadd293a3a89079
zdd23b22d0c15ecaa57707a4f502669fec707ba04e18765701a78604634a1c40d69fbb1088cf92e
z2ba19af43fd36497dfa49914008f325468f6cbd36a233c6a49d6db1f4253af9b934b9ef7ee2bf1
z37db1ad3137cc70713c9e3ef343d3124261376cd74527c3615fa41f98195d9c8f93ecd551b8c83
zbf0a0f0a8c449beab23ca6be013bbddd30193ea70789a0e0108ed513e6cb8b14216577cfbd5c4b
z9b1639edde131f8d3427429000d783c0fc20021bf5d36f7054042f385bf3f860753df7cd73db5f
z88eb98d14b570f63e46fb02063e70805ebce1d433f018af7d0195469575ea93da85e22fa7edb12
z7a8add71424a26ac62cd20c3eabcbd305a6093fb82ea0d920a1a91c7ffd93a1a69857787272482
z62b0416ee121675e75fc9f7f3a8abed537f6f6577a6fb96c3407df242e3a06ac1033aec57a49d7
z837afcccc83bfbe637d9e2e21da36301b3746d383e674532d8403b051de071ab75d30cef7d8377
z960ab12d99c057a589e0af92e3a0db0d2a93cce3f843457f131b70d99fe8441774e48bec565038
z27d53efb4e36fa26b7f1d7387bf199eba3deb358218a9ffd671bf2b6dc4b994c0b4d4cb0aef219
zbca89888538f0923fd56946a38ff6fa638f50bcfdba601e2106f163b0d17f5966d213669affcbb
zc71f8d0c0885c309ebb55a2d67ca4ac699df42d6b1ebf84ea07f56effa11d900971075c3decd7d
z8ab0aa30dd29cac7273907c19d2a2f865d1d7f37e3da29b48ff5564319f365811a69ee44236528
zc1f2466cb0c138d5d63182c25cc972a3dd9471c9d223fb8496a03b665e7847755a96889f5193a1
z3e2fc608b5f6d0b8f44a80c8679f1ffc379641d98b7ee088d77b85c923ec40af232ba0141a5eab
z7e277e654ad56415b9102689d9ae4444cb7fb2d4384dd2402f2d80c0fea32bd28eec5181a7f750
z40086559fdc5fc98e830c96f2f251f670dfe795f1069f0140dd455e320d4906a79a89bc9d1d306
z5bdec0b596f6b7e0b1f5837248f59d5c451ee451bdbc15c6cc18bc3a3d58a9eb84088246207a2f
z475bf47e1950917ad085145ac2c0928547deb64676c4ef3265bdd80a0a808c6c37e56c94106314
z74205c52091a085598e4990ab29cddba4eeedded6657fe3cfea936374fb26cba0578383778bef4
zc45518175f6307957490b2a73c7ac0a82216ab2a185c31910723d3554474b23e1152a6cf550834
ze3a39c03bf77184c39379c5d54f155ef8eb316dc750ac94914d1dc3dae463d2012b0af52fcaaef
z68b1a7c4858fab5d39fdeacc3f867ac50bfdf532f2af48b64498ef443d05647c3c9c5bac6f343f
z2a7119372c1e827ab25fa19b0f962f87c57e4e87daa425365fc617cd776f4a35034d82dab27b18
z29b1dacbc795b4439377539e14f511f64c11e2e6b2b96859c4273e21c5b754b8c996591eba6696
z86ab28cff95d2ec81626a6aee0c941ae795916fc76ed07071c4bed530afd3aa3452aafac1a1d22
zddb4e8d6ab29e5124647be5e1e2506a0b8d88ce17f5ff42ceedb9a9b3036d12eec079bb61d8714
z9deefc33dcb9350b0cb29f5d6ef6563e2a0196ff1f1981ad0b66928b895c5bfa0cb7372d2a0c59
z3a0ab13aa09842e55d2bedd96dc69e7d6fd8bb5cf919322256d15a0cfb835209f5441db906da54
z469b73d67251e66ee556f4f3597cb6b2e526bc17718f15b903c719c5a04aaa5ca821b44c0baae0
za618b6bb2363903440be224f10a1806c785865150ec28de98992f56d3f15f75255f58ec54571e9
z98b58a837008dd910e40a088e40c44f5f1502bdc258bac66d892d9362bd174de34468c3f15763c
z21c9c9f7583b43b01e8f2425746f5bf0365e4ad112ebfbd41c59f5a4830c553e3391f82836a7bc
z98f3e708c8fc11001bed6441542892d6b160be1dc39a7b5bb07482c88bb864c9bdb9f5de477d9a
z68c601f8373c42b584556030921ef7eb629dd1ea65eb29f7b0b50d8a9086bbdbba902a09130043
zc9358bbdab0fe02a163dfd091088cb3d992ec1f41cd0d3893876844d5c346d4c8ef5e8f6b77998
z192db0b19491cd739f4480a12972e8fa0210e813d4c9a2920bd0627308e41adb14888aa9a53e88
z57094e4da81451250d117f31e7655d9bad51dd2e8a762a736d309ee2f9cf7c5bb30d1b98f39579
z295b2c2842c5aea783ed7431b5a9c10095395aaf1e15d7f26c006ec4bda7a4b68b7f9f1dabc2d0
zea4d822a5341ac965e5ece685709daa9c257547c270b7a1fcab47806b9ba43c16c69341c7155f2
za8c7b70305a4e9640face3780c57f0c8c763fb626ab556523be7a9e5b23067f6cee76ddbe388cc
zf87637c299db43a8fdc4c2534fe83ec066cb24a822968086c1b72988689c3ed04cf3d9b7ffd494
zb7e7aa36a703a4edee51cdad0bbe43e04411a9574ad6ab85bb011c329ed4aa6dc0ce0c4d493684
z9b66a97ace57f7b399211d21bec63034e4f8a055f0c77ee77632d9dbeab8cc155cfb5fe7a1eab8
zb624a2d15f9ddd952bca5d02234567e7923ac51207a4442483652d3ba42a66516560cde522d751
z4a4a9e9bf7f22df2e02a2e69f84ff632ddb3b3bff252eda432ad1c3734f2e25ae498404a75a6d6
z2791db5dcacdedfe43284ca2084162ca6076bbbdf0f4339e208417d9d7b41f4f7921a23fb4a3f3
z56f0b62f99d8275f480e13eccfdd181f9d4f420be1eadf76a800ecc2a6e6c51eb18faaafa8afa3
zbe8a502a4cc67f3b6388d92482f0c35b387911d2d647637720a0a5a42467fee6148db2f8666c61
zef6a86ee1d2da7604cfc03be467a2986923836d01b1b323d27cb0c1cb77e6c98241a19b8e932b0
zf17b8b6847c7ba663e7a857f81082dd1b2514fd76eaa0ec5b1703bb30e538eb9b6e08fa8450b28
z2d67e3e5f650bf3ff162184ce774d411bf3ef1e55e08533d68bc7399672219591f4cc3d73bf75d
z616a97678c290f22c064f0e231bb73890c7b63d473ca785d590637cf691940f8a86aa0db0adccb
z6a75605a72f994e0cbf5aacb01229dde8bfe7b864d7f5ff77637ed5fd6135d01196861759b688c
zd65f0aaea731061e2ba852d0f2474eac1cc39c4e534aba2867518019abb54ec0bf048486c1a71f
z485c5c1068770e1280e86c0967151aca31a8c41894d18d3f03111024a619292f6965f340a4f72e
zd3de7dcd1c23f21da43e901b5f055d38c0dc5051a9b83f67a224c9eb44cb9022493e0e1638c43c
z20e859d70d8ce3bfd269c50bfce980fdc15be09d9dc9bd291bfb7e20271c763a4cef37a602712f
z048e150673c37b26785a94efd36d196f79f76b705d05d14134d8537a8e5a44ce5588ac2d080f0e
z6b1e877c4942db8b487279580e624c14980c9b3e133940186a75b35dff7954649451184a06f2e5
zdf4bd638f7c06b1af01d6700daf1a33aa2783d490bd0b09dc59d5cbcc32051882610bf20ce65b7
za8b9e5995a4f569a4eaa3b196f4e941657ed9930fb62f436c3560d074988d362f1643bd2f0d7dc
zadf9a2d2e09590e580bd2e8febf9beb7ee7d54e1c90df565036b83d64970625d6cc1698ddd5f96
zcf81e8e41595050877fe4af83eba717ad5498c331b9b9a81d4b6a05f7c9e2396982d66c14cdd76
z37b3d4f144e2874fafcce5aea9877ab9b9736df444c3db00fc020a95400f844889d6292850bfbc
zb921e4938b3fdedd76e588a2210005066b004782fad9a4b8283783ec6de9a55974bad5bcf016eb
z8c3ba08c12cf0690d0524686c196ee2d3da698419e9a82bdad2e11c9b3297a9ec66893bd82c38f
za7e7bcd7f1412fa0c62ef3ca72ba98a41a367a994e86e34df8a59574b0764bf458d1937c5a66bc
z62e5a67d3c552a9b195e4308223badf910b476d2d96ce61547fafca47238078e0d7007eb71eb8e
z7319375d5afbc09f51a0eff4208a6480e3db2b81222ff00d7b86ee4c75ee33f74030b5282c25f8
z42314c041945dda6a481930b3b4a50967d99837007cbf12f34d2bd5df1c13166a3ea2f165c820f
za38035d68b035313de277464b247939a79940a70d136997de9f02f9fdda9afc7ff0a3959552a1b
z9570e1149f1c0f8974d78450737a7d22cdeacfaee84dee45d97d730050111ad24d6d84c04f1f86
z8415312a3abd2b497029c6e49e2c4356b83f676fff9e7dd1038b45c9bf6d05be3e5c7614ce023a
ze9c9cdc1299aacd72e0d16e5ec1b4a1244ec54ea53f58d74db2c6a4b16ca805190aa45b7d644d8
z8176e3af46a700cbb759aa7fd864ee7859558a30bf06131d8bd08744f8df63440883197ef5c03c
zc58b6d702a5e8aaeb1bfad0079e331e8edf63f18c7ee1ca51f255fb53b319b8b2217b605739401
zef392ff70c22a98639c82faec8f3032a75a40269c5a3133871255c3d39f07fc785cabe4038e248
z117db0875de1d704fb32ac067c30d0249c74cae4e790c4e76033c8c923fd4ef5f102f1d34a9f81
z33877a906f2db10d8bd35181fbfe5c5b88661a95c63ef17755cdc8105bab770d4240290f7bad59
z8eaab20d1ec62974abc1f54304bf2ed6c53151ec6fb0a62d33c8b3da9e40c45ccf08d9ebed3c51
z1826fbedceaa83c21983f3ea574a49fa7fdf175d4c9952f1bdeca4c566c15fee16cd6e68b037f6
z620609b4916d0ac445b1aab44a9b4e615d716448d3267d038613c4e28840668c195bf1519d1fb0
z5778d42dc20cde0642eca547365e0635163d8fed9e18bb7701be7d02ad088f05c53b0cb5aa10f9
zc41d03ae4cce99718c68e4a0847db448681487d83158842cc70c6902b1e6e090410e7ec304001a
z6cae634dc9bfe4ae8ea903b037872991d7047f2c2cf3c22f159652372614705dd20642c8ee4588
z393826fe87955160aa74f70f4856b5a77fbf19862d0f16f8cc08ac757e3df8b0a61ee9dd8ba64e
z920e54fe89737c18109157b95c5ded71fefd8b3910ee6021ba5d39fdfbaadb2ef81738b1ffc91d
z716c7fd5a234e3ffd779bb3c7735c59641559d166071fa3585a64d5aae83e5e8340cd21512aec0
z1f5a2e0fd82d24fe3d9dd1044017d241c47c2b5d5951e9254961095eb732fc352510832f15c6c5
z749a70661e0a6606a1b96800d69610a9a35aa57bd83115e504f5579dafa1881be5815655f1e103
z15f2d5293dbf10c9b193ff10ef18519891b6756b4d93a94ce6b74250c2c76e7276cf92428040d9
za6a6550a9d8f8899ff0321b9c4253b3220c105a0a68c553c988b200d56dbca1218e8aa39729336
z0bb23f64db8491817afd07bc8f364ff87ccf1090ab3919607d1738a0397c24b0247042b2bbe051
z470825421c374137b668fbc2667264ccdedd0a0492ccb2c575765d2b550285a683de6fc75f93d4
z49f793b640dccca8b6942e6aa62a7bf7c27300122227e8d8b789656069bacb0aebf98ba925f9b3
z4453be4cf23b5b68f714c3c5b25e6d0482761d585b91997e7e8f592bd6eda5087f1cf2b946e6e2
z9026313fb09d9b9b927432682db5329553ec6389b66a176f44ddd465b363731b3f2ae77da5140c
zfeb63110a33a4c7c2aaa551e2a3b2ba8bc9ce8b40a1024c60feb9e444dc77b6fb9c45ae7f5cf83
z9f20962907f9415b4b0602447af496dd975f6b859b7db5d28d5e73b3b60e87ce896b059d485ef7
zdb8553a1f21138972ea9b3532f05edeb271c04d1bb10dc2f7c9bb5bb03592494fda176883f4e32
zf0646cf9bf3dfda79250b0b268b67ed81bd56c001bef50ff7f609fe9f9e4aa90f384f6fff5878b
z23a084dc5a443761fad893df7e43769541b833c87ef369347d16ed3dd5933736a31e8b7bb31574
zf7938e13dd19a22e74e30a0195361e56b394eff9799a49f0d4b329550a77bb72f74b3bd854428a
z46c16791ebc6fe0aaf5bf2156d4955d7f75967c3c2260da3fb65eaa0ba0778c7a9c02378f22a3a
ze80aa80ec1812e7f2188bb96b9288a8fc47170b2a4ec5d9083713182f982a9fee555e18ec8c5c8
z8b65310b5da756c950646b6b9912a408383e2b568f62268d26f7a8c2570a49bbb4dd27a45918f2
z1a1fcf6d0b9dce62c5c85fe718602569566d19c3af20d1af7db45da85a7207a439f5eee7233396
z1d01aac5275b79c7457d0b1e2028172254f87df21051391ded7ff5a8a9762769b27e1f3f2bb974
z6143609fe76caf3e531a848db21a9ef8b4d36ccda0b0c449fb6791eb23e369a8427a5b0ad19adc
zb09b49bf8620a41de54e952961e4ed645b4304f77b0108d67e9d550a5c931755841e8e3cc8fd32
z22abe4bd18f899b1471fa89cbe5b59021d413a531b431764d43ab87c84c05a5b4168512251c625
zd34951e7e5ae130e85b841ee414b8367ab9388251476f5b8c7339c1f8ce346e4fb6461919c32d1
z9aece36fcd12bf1d88324d843fcc02c8c517c8170dcef14f9f055c7a302241ec0658c0318d2862
z8864f99d8ca26e930da9c03ec84fe4c16adc77443504e8cfde1cb02afbd5aa7fea63a4b0044363
z893f47d720467ee71c0cb7fc992627098f332243635e62d027dd9d3236e84d958beacf98e934a3
z5b99a0d147307234ff929a6188ac1bae59b2f214a7208b614669e5e40616f894ca13d41c7c9131
zdae512d7a952861c3bcd7334b281ae307415ede2346cab6d03540e1fe220b411780a2dc1abfe4f
z0715a21f5032a73d352dcf25538095642ce1501ab84384b95f6df6de38babdf04765f452fcb553
zf524d7b7bba9cd28fda3176da6cda6a087ceb937665afed72509a0dc2ff459638dcc1b45f63bf4
z80560172a6297cca982613308a430042699bc95e143beb0b2996637ed1b10cab8634924b6cc723
z41fe1f45e7d0cae775acc477a3cd56b2848f1b4a9c6db7bd9128d2b06631f99f652decfc7a4e9a
z93a9c5db1a9f9b3eba25c9753cc0d4eaa491e01626ed3f275f2ddbdd46ef7c3d69aa4f0143427e
z55e9653763e0a214c43a8a87be9361a8477a969f0fab7f787d354c2bf339db98ea2a79f5592e01
z569a367d4ebf38ac684517707e08ae7b3518d07542e657be00b1096583138004298bef3d2c459a
z2aad6a649d72ed2359f4b02d24725d8a25e9632df852052c6d5f652da70ddb97594efc0b707427
z0d53c2bdae3dacedc4ea2714ca7908ae6c55e8a4bac4274c21487f0fbebf7774d4fe93ddc866aa
ze2753be37a080b14cbdc760cea6abaa4fb87045a3e4600f427efee68472510dfab744659b00896
z83d806ccb3af061dfb9adbb690bb076e96bc4559fdda72aba5a35acec5f4239627b1dfcaec1777
z1f5796eca23ad5024cfd5fd412fb0a59a3e0d1d0969639bd0af566350ef26bcda13ec20682e491
z0729134a228bc9d41ae23ae1aaf4d43f64e3d0b90541444163951b4e2a5b14a3d20bfde9bead0b
zf221378f6cc2d029e5e50d7a8bb95b77b5b4e00c4570164bc971d7f36f4bbd194b456f71d91010
z80330087403869398192c2cbd6e3ec114259d0625c057d9101a10de0c3baadf41b659b52a2d0b4
ze0c212c5150766e934a17d35709458d63a47ac4320ae3c7bc383fca6426dbf9e46275f576bbb8f
z2676bcb7aa3d2638d47c3d4135aa6cc42664d10c7a106c8b6d778b1ddae7b3916d06607b3743c8
z817aee39c137ec5ca6063668b2fdbfcf01b5b21f39043cfbd001ce130d6bd00b47f87726bff84e
zf21977e6769830e85392ce24fe5d256fa53b6cb76cc79de81b78ebaee12bffec1e18203728f5b9
z1115f6a6cd3db6c062cbaeb78ef03151143a40b2d287b7e8c5df623f394b945796fb8a748ecd3a
zb42932783f34f7b786a65a84a5c512f34e2b71b9e403da6f4ae928ecc033cdfedd338e316d2416
z6f7af5d18f03110cbaffc667733387ccd671b9e580f922c806e7bfa60ad5edc95bf41a5f6934ed
z841b2ec03f66d931ab5bc7e451dc8d667305244459da9df171c87986fcce3e1ad9bbbb4b910651
z1d0394b301d4a81ca6743959e04e1c2da06062be70da8c0e72c4182219f6c0a8ff77b6b052a603
zc45601505f8e168df324549a7661269935e6b45f53d8584739228370ac9fc277f4ad742460c5a6
z3b446a0750c71f9ace476baa70fe25713dc7b72da89f208d29c447d61f10c7e53594d203eaf0ed
z843d4a50ce79b2346fdb3478b51b63d5223cad0901096d05e2c183c58f87913ac1ef59aa35d1c9
z0583c04f2cb043a96504d36634a7df95b5742b5548ee26fc3abe0e754a8fb4c8166d69879bb3af
z535bf33f139cd3f1104e23c66affb48bd84832a729884cc01d94b7e6df1d4ddde04b9bb351323e
z2c0371ee0f5c38aa23b8857bec72f80188b9dc84e353cb76eb7353f2fa33c124891485470f08dc
z96c442773b3fadc21b547fade29cef0e01774f1e5db490fbfae3fac565b7d9bf654fe73c269326
z51cc4c7e86488b83a07b15495e0df7edb962831a847c49702d8152206a92caef9378c05f81778e
zdb8b0632c5c97c9281eea2e21c17cdd15bd9ff83ee3f12553875764a2b9b5f627ba93f0ea40204
z690bbd77aed6935a89a4ad72c15c45493ffcee37b35ab40ededcdc5618f98a927818e95ec78bc3
zd025475bfb6fc9cd6abe3404fa66f24bdc983e6b4882f6a3ce868166d11a3c58a157c2221c3af6
zd184332ca18cf6d55ba63872155136a2de446613a78f651e78c531a05eb949ddacd566956b0609
zeec6c3144c29604d01fa2b50daa3574f510ce330c6e29cf329fdcef3d30b443295501308f695de
zbe3e4f5ec5c197816adb3d55dc732caa2434e6642931ce3a771d2bb623108b8341ed0f0945effc
z768ef54c5af34f49df490fb5f27caf44acabc3bb6da514dd14127c560e5d89124e2a0d32751567
z1fe1f0bc65bc27f854d5102312148ac70c8e50b33194a7af5278260c03bb7ee3eb0496a4d67d16
z8a8ac4e1e4e712417e4eb8ad345745b216b59cd5d69dd5b9cef0757cd3f9c34df054d2e27d5d2b
z17bd903995294843a05cf483d299579efd10031ac3691ef95db9db710c013c67401cf6e866fece
z4f42c1009cff4bce058c8fe48396276a61fd48907802ae1043e7689bb5a6918ceaa79886b84bbd
z3b6dfdfc09be38bae1d9c2422e68b574e54c0a170b85694926bc74f44b7a5130b716be9df3e714
z32e368204d8324dc9c5b98f11bd5d7253c75d0db0bb50da9f59358f6a75b2f866d0253ad1c9ca8
z08e82ae9fb91e3ae714bd3829f0b09095ca78fe24d1aaa1e736cf146652387b5dd40291183503c
zd6d2afbf39a785278206afa19a2b83bf60a840950aca82f03f985da25c218679b60d87102fc09e
zb2672d5679423c402adc7e020d2706ad1c733f8097334a5ecc43b5c3b40a62e44a36aaae344fe8
zab0f449cf6d559647d4ed4bea5da9e6c3c1d0227107dcd72958bf2ddf435a1624fd3869438d143
zc19c14785f5d0b2d6f019bb25c551b8225679d226d4f2b48220b5e7b638fa8fe4bdf94173815ba
z4396ea4110aa3473f9ce38d68996e837fc131cdf77b5a4e647c70caff47f6ba4f74276e017ac97
zc192d83adaf60eb87d0043fe8bd516e6f52f70727170ec06ade1cfc34c8a3ea3e6f752c3831e1e
zf2e94319a82cb653a6f3f9f78dc15c8bf0fea6c34934c918ab2cfed52cc270de577bdbc3599bfe
z0bc29c6e1e73b04be6a16e55c1e803d4543eb532512941af6ee39ba601527c7e72f53a6d09100e
z405993dfa0a1e6f66f0550fb81d5233618a5f4d89505baa126336b9cc677012ffdb1807552d448
z291a80785fe94061c578134237c2bf2e054d0502a3a1e58eb389b925dd259dfd15401206790916
z7143291cf8c245e49f16f288c31002fe00c51d011f83b2a7d2fefa8213a28f28c5a462db1620a0
z56ee6a7445106a8104b4c861a19e52fef3300d0f58564aadd7fff830afab382185233ad0aec90a
z1dda2732cd2ca3fc57f415a800ff165612c2b058f4f5e9c6a556ec235fddb924253ff29c435e85
z73bee322dea85d9b441bab8d81e7352d28256dd6dc8ef743b261e9b7d6fc81faa6267c8527e337
z22e58294d0b984fcc1e5187d7f01a56a9ce4bd8e37cc22b61ae9c70e18d97eee2291c193802beb
z54d71b25153e94307d0b79d960d12869d3693f8e420f69be6e3cba9e27e6b01c6de0b703013ff6
ze6a3ce0c2bb5cea8e593e2ad1ed85108d762c6876b45dd937d3f621e9349a2cd68904a6babcf81
zce884ebf2280dfed1c92693217e2b710116a99c335078dcac935dd5c465d26ef453a302698a709
z3945486551420dc394f3065fa5897765a564df18def7bb2ba2e81a9f80802beb917cb972f3b847
z225510ca7c65feee375a740dcf16cef66834e326382231f78eb91020a772158932965a10272643
z58ef9177952952b728e473a3d2eac0e6f6da7bc917ec95fbcee8e52e3cbdb1f181fe09beb46c34
z8f954397526bedbaabf9ff6b58300b7b84bae12f49b21cfd4a0a740cd78b88c4618fc4acc6385d
zd1ad8c8ef960dc2737e8955ce589b9487e65a8f4494fab05a14aca1448051d44d389d277e72718
z9fd975e6e505b19096f9e374845226348e243685af7f7678d0caede5ec07fa5b9de34480607317
z5fecf6ef288f95f208a44015b201c1357a2efbf4a37f4bc6fc05d4cb282ba188c20a1c3b926fa5
zb52e4ae19fe79557e3e3c08f407b18141c78bc3d3469d538ebe3d1a733fd83f253524e4af1d4bb
zc9e889e152047ab1155d969cc0ae8e12368f3a33b8588e034ded5ce3585372c728a9d318d8d3b1
zea38fa36673166fe9c307f0ca7466d6294956656efbde5de25297c3923f7015f7973c8473b0ce5
z5f5e6a7c1b98f57d7bf8b88ccd59b71e8c8e291b557102ed1f4bcd8403791775739ae4dc67dfad
z1bef363a86dbc531b9963864223232f976b15d717a515ae38af6c4bbbb188fb76da90bca38fd40
z3e5ad4edd108cfbc9a554c8f9d9a526c3b5c60dd4715ac4f53534b3b04abd52ff29168273b6ee1
z2d6e407239030f495098df60e049f3de3429ab3d5576f81f1d4ee1fc730e4a3c6249ca3f0f3077
z997786db57c2e436b045419e101d8f125a1187c3b568cce057a59ab8f69402cf87562a6872c4d3
zd86d94eef13034c06e3890ba6dcfca6e20af8f122bd541a9a09c46b8151977362434f8dc77fbf0
z64b336fa92cd4a50749237b7b5de9512310755a5e018eb33965d47507e3309c3341ba68ade0d42
z95a0bc0e1de0fc18ccb50cda04c8fdceaec31eb420e5cbd5933b89a742b8
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gigabit_ethernet_descramble.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
