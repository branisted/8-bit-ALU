`ifdef encrypted_0in
`protected_0in
ze74c34e226135848c7706a11f6cf56d8b49c00783f1d62fe2cc4177e167684213c97c457199d07
z85bce6f4b1df2552721c5fe686568b965d45c530886ff51d724d464f782df52e056f41673256c0
zfdc3d64f035638436788b30bbb008e02ec90a86fafa3aa27ca76b1cea351542dc765fb540e8b57
z9835c62399956dc41713b282cbf51cd3eb799dd44c969360de5949799890dfb617fd4d3e8154a0
z0a0e2afc736c2af5eb14560b32fa244ab357cb5a615b450d312c3c10815811769bc4a7dca77f3a
ze6ee4ed0b1787251f75834c506964ca9fe9b6154f8064f60e6816c22cab6e4874a8226e0393a1c
z104606e5ae362d4beb54c969715a5781ed7bbbf376191a0b807cc97d2a9a40a82c555b4d0b511e
z03930ddd090d1039dab2dc25f8b8db1e5517f4eedaf5e41f7e4ae9a3b176a5a6ea5578a5e349d3
zfb5c3e82c523e5cff087750b886bca029b4501befdb5135e3d426c351f2d93c33a9bea3528ed54
z2780115db5420d53bd81df307d89aa45326a4d90def90574958c6060764bdd9831db72c15a3b4a
z253a0fe1d4070ff20f96ec6e6f59902348258c2faaba53828f3b6fd49f93d700e76d80a4ae15a5
zffd9499ddd2af48afd4a98c5f0924c68d415809163ce8234bbef78baf47abe6382b182d6c28d6c
ze181cd383b786fa1f29e80373bb3830d582a721d8cf27ec70ae5ab4eba672ec30f7a26bc00701b
za3c4332bd8ce8bddced3070a4caabf85cd0c0d84f4a8283e6a6bce15d292edd198f817feb6c97a
z8960d4abbe7eb5b11666082e522bc247b9f9669bd5e0356a73d95487afdf7cfbf4ea5434e4478c
zf20b986143d8b1baf8774398860d11a8fbf28922341c827ba98650ac51822464d22f250123309e
zb70ee516ed1ea9fe50c7f0424c07c9a4d91348ecb50c4f39b7e9aee6a15bef09daf9b8ad03b193
z311c1e9bd045a39dc04347a599f1ca52f5be790c63ab05df7218cd573b57e4a604ab86a81102f3
z4f1475ff686890a6d4a4610a55182d3cf3d476db128f60817c8430643ce4277cba0cdbb71abff6
z6d9a0de90035c3bc245072fc4efdd923004d4e16e0b3beb62d29cf47e1a83f174b4cec06898ab6
z33997cd2ad3f07ea9cbab3975b38ad176af9b078e40dd1113ca2a1a9f167fb1f8cd7887fb92b41
z29c43a69db89969b37fa337cfeaa714399bab4017399162f1e6820468b86d7b855f9546a1a28d5
z05202469d2b73d2b1f357b0103959e7ca3c6a6cc1586414e50935e261027865d89b7e1a968f758
zbe00bca36a95f45237ef6c3470c4ccb8ef39c2ea782dacf13ee8a01e613f446c7d4c41ce833a5e
za756e2c4821070106f8bcba87039fd8ed6836585c0432825eef1acde8144421559e9afd9d5dcef
z44bc17ceffec576458c55661aa51048a5bd68f16e9a6910f1f3452866a63d73f7397cc1b1c1675
z6ca3e2058dddc8d7e9f8ca876d404f29b8e3dc7101c472b9ae7b0b474ccf0b35f1a9e0293ea93d
z8b8e673c4fb614e85a9264905502b01d8126696c8bb3ec65c9dd8e3739f7b277f029b593e1c0a3
z4c1bef43ef3299b3a0711dc8135923a3de8b082ec5ea370f3e1a7cc0252c057ca56569200d3713
z515a7a0b9d2b16c43153ad1cb7e9885ecf628f9155a1ac6e2a16895ab363a67716d8a83beb4722
zb9d19a6ca56379396be66598a37c1cd4ee2a382c764ccff79b886c5e31dbc9f1563a94b19b265f
z6df9b6d5d22563f0c382c3018a280c5da4ac3a3cdb755a6dec22aaaf75b22e68b44dd8d020a4cf
z3157768bffbe94ae672a080933b4bee31d3a79ec037e1879502d46063c08149dfec7b551c07afe
z93c568be47eb6145720af91fa6a7b1396c57983c5af5698e7daba49d73078c431a8d991aa0f7ef
z5ef6ea3af826f5090542063bdd74b41fcbcab877999a1e21dffc2c7d65df0174d1f7ae4ba3b3b5
z38a81cd467d3eb62fd971b8c737e782ff69493e17fca790d8a4131f7d07ccd8b5ab34d26eeeb6e
zb3a89852ec6782b763c8695fff458b5a25331242cd9ba3f7bed4b1998d2c93a5ad9df2b674e58e
zcd453f09f26641783445ff468905c0df450c5992c4c121d85d4c205aa0b0ef5e9e5ee7cc3ec873
zaf0e375e08030249540f313fcf46af5b42de72a6bfe9d52247e19605330df2a6e75beeab96fb50
z37535cddfacfbf1b912bd76cb2eb39bfa99aff981280e9699b93825196c190f01c0b48b38100aa
z9e7d1cfc779014dbb59f3107617e98427660f720e2b0b5a9c822922e632cbdd5da991afec5c5d6
z4ef1db877dd55d10a68b6e2b773b5564eae4650e1b0cbf8bd68d066e69bddb0596f1e0e3296df1
ze7e00a8268b6e8391f2a7c76746f62481745bc8fb68a33d5d9f22573e5f3ca09aab47b4ade04e2
ze33fa64a53fe2e3d165b2e23092f1ded2234842431553a591dd316d228dc84da97e3565079508d
z107d8a970b25f4962be27b563798d089249cdb2f2a7de83d6a34ec6ac907e82f78a124efee50cc
z61bae2e3c9e189b8ad0c3a78b6793a6eb95a6ca725094d6146c842a62123c972c80459d5f45fba
zc04402c6cb2e21082fd58829885586dd04744b1176a2b776a27a76d7fde47657af5c7cd034c47e
ze8d7f2e9604fdd5867f5d981cfafe7a875519e9cf88a19283a523e138fe94ca4533966acd6e507
z0c7d95581666993b4157bdcee38e857912fff32a03366a32aca914ca56b35e79432c70fe02a20c
z72611fc7ebde6f958745a8e36208f9135bc199ef93035aa513e429958a0082a1b38f5ea9bfded0
zc9e372a263a42cf038eaaafbf19c20ef4a740692de6a8f11057262afb1116947507cf400576162
z654a3bee5ded8024e88929927d2150ca739f61ae3bf1f193801c7293658d911ffb373df9e81fe6
zec6bb9f480c8334122072f2c6f0a11a62c326d0116feb3bb3f11d1c0c48c53725117c00447660b
z03e9c3856b33f4e0fb609512a7e5b143ca25cfd2e01e2cb12c39b7139a982fb093c87d14a949b1
z74ceb317b21ae4725b24699fa857663aac8198b3aa60c6098a833ef6dc3833b3ff26269b45524f
ze93a4f8cee5ff89393950d93b13ae93dc26680b1b4a1f20b8049017ce8f562a0b62c9b399d19ce
z06ba4087168ed2644ef814412c461e965ac0f956d638082889509441549e38a45f7ff8ae26a370
z4cd6b28919bf953bbeb3453336c5826892503faa64d4b6aedb0aa9c023249f5df5d1260295994d
zb2e70ad2cefdd6980dd05ae72c67ca06b7d8c5c97f36ed70b7ce7eef505325c6fd634f7a6aea36
z41f07adc733904d3a17bbc28e310b4c4a0287db0cc81a908faa3c8ac60d812005693bd5eb691f8
zb170a58c212f4651bfec73d1f4132dd030d427d47823901c9256190559b8d2d7658135dadd63a8
ze41e7495d4f5ff6c8b3d151078038e51098cfdf5c4e02887e0ea314cfcfea25fc1243385aa9e84
zf69978a69f28514b8003fc4657c0d574964714023f175967c10882f4c966cf435c1adb819b15cb
z1ca375c478d6c4f4886acd3e9d6ead042f8a6d5af8ba3b6935014f1de1411286da796c8554868f
z00bec5da88666135b11bc63c4ddcd91f5e05d132b44b331a3e7923aa6ac3349afd034b1e501595
zff730b055d64306ff61ef6e72580d95ebf51102846eed5a873855e2513e99dda0ef7fd7fa41bbc
z05d835bf0f09529b4ad31f1e2ccaa4c50dcc72b75c6fcc29fd4e2d368fadc9eadaf2279f030f7c
zd07b9620c1e8daea13d0437b39d9671fdcb36c59a1a626099031ca5b43521251cc61404f318aed
z2dab1a6123bf432f1304288d479ebf7d220206f2e82c69f9a6bf067affac70f897e2d66b0f9b42
ze5e765658c917dcc05738f93418ae02d0240b5ca625f8fe538ecaff154a41ccba147ced8403478
z372b2920d93cacf1ec95e851cba598d6d30abfeed69d382e187c965f346df5ca47a052f5fbb010
z51e8ff4669a57aa68908c8748edfa6d9dd688b0cbb7e5c47b467090166955b56dc8037c7b3a64a
z417265219e1c90d1b021fb819d42686572e49b4ef1a329029ee75125416ba16c8fd4e5123bde32
z8cf8a17fe840bf40d221b256b11e3135b88d3e7696e8527ff8ef07d5ab0c945917339f9f163830
z12eefd6725524f73574d8902458df45dc4dcc1f4655e0f666f53f6a4ae7e3d89b66f3e2d5399f9
z781ce3209e0890b35faff6266fafe409cab634e94c2f42f922408343d714b1694c598bd27c9da2
zd096bcc50485511622e871d947e8694cfd36a835fe9a08d241ed8b107b70ff49d88bf5c11adffe
z80d16ea6ad09d1e9f02fc98176de593d8e90d8c24b75f1302a80466790f42085bebe1471febac0
z0a26486c22e08a855501ef421c1d26dbc8bae5ea7c35bc7f4316fa7fb11a000cba347314baeb41
z9e1a7a0d913f951a2f354b0fed25278c44a2e995f040af822e80b99911bef85a0585e58c6e331b
z560469aca01f07dd2d7f292a69d30d72f6cb2377806e592cb452ad042a180f0503fa6b609734df
zfa9b85435240c65a3a1e38099e8fd8dbcef31032988e7bdb389bbb682603e46a1b52a4fc7b1e84
zfefa7bc9d4c849f5ca1320de466b72ecb97e58027deb140d166ab9c1fbd0d902a1a3d0389a0fb9
z865bb5b7940cd192c961e1f776c1e975649ec77b0efa40b29c328c504b26d93e99ae2588fc1ecb
zade558d23e2cd0b98c96253e312b9e76ba3d460772117c21d0ff8d9e06f087134a3cc6feb1c70b
z88e0dd579488e384aa2edb5c714cf61d487106c3449c419e61acb4a167332689aed341928360bc
zb5459c05201efeffe06cfaddfe21bc96a5e2973466d9d6f6dd125105250c85276f9af90d40485a
z5ed0d837ccb9f8d294c41ef3f75d8937009fe5112b616842fb3812caa05756b02b6539b5ec08f7
z381f205079d80b6af88615c4a866f71a57c514af552a27a3c28aa650052d07ce02886c519be355
z390729346a23867290c4008aa2d5a6659cf7eb6f2e15f87eae45bcf54db7d9928b7d5232679a85
z7980924aa4677db3a928001e8d7025472eb7548379da7ad7907b30c5d592d5cdade9e0d82d0d2a
za1ad93dfc8451306155694fb887d92f7990b08a92e3ecfb5368255adcceb5911bfb43ed3857b96
z35ee159e0724d9c64b09e6e35e24545c26af6f892a7f5ea11ba997c99ef53147d04f6e5c54e838
z3cfc6c97ecd85f88c978e5c0ef0bca8ac851c3a77c23b109ed2cb3d13a7bcd0fed05546d8bd220
zdd4f731396b4c062768234f1a686984764c62faeae49783048b76ef154f4d2f582aeb11f8a4dc5
z856bba2087c54c16cead59518d028e8825bc487bcc1f170463bc1b9a1d31033f37b317241be754
z1d37d738b4f8684226421e7a8d9ffdc79dfa2ac50f75e8e15d29ae67c8dea14a60394600409c65
z10d2d60d1925d14b324ef3a6806e752ff05d5598cb73a522bf0fa17943bd7089423118fa886c9e
zdc9862abdf5c589de23c58a43fd708327d197e7d0fa6973a31939090819f17a324a98dc48163ae
z2dd1f69db862e334caa596e228eb79b9cc4fe07a36a6b5f9ee66c446ecc3fd59451d8b4b5bc05e
z61594a331a651be3d32c11ad48df33465443f6557811fa3ce9f7e0f004b10b3c1fe87bd5de80a5
z09b2cfb15d895247e262ea3ba101df9a3fc92ab8d817bc3aba207990698de61c936cdd839ce9ad
z184e4bcbd9aae47b74ac86e449ec3fd33ece15c1f0885e760a78d98254837c269dd30dfc3dedbb
z85fa56a321de4ff60e4de9c5d6e607f4ad65f3bad2f14ebf57b3b3c4673fb1673746af7f226648
z308b91deac7abd8f8cddff16053a89376181771533ab2ce5c14a0fd61b499f81c9ec9e39d03eb6
zb86378df140d8235ba4174bdda004aa85d692e1fdec47f1fa3c98d123774671916c0a011d22239
z419b1a892ba5bec718784a4ed83e77939d5026bbaba5d9a2a2771e089b8c2e872ab7de11a9946a
zfae3b3616f1d8352fe0710dbe3f075c58f2c9f332bb9cafc37193b69562537f965eaa2fdffb7da
z1ca7ab56546aaba8d6f2d8ed07f9ec91ed342e1a41ef29b5886fec9d77376eda70de4608de2098
z3e32bf3f39e5bf4d93feadf770e6f95b641b08353ffea4fbd12645cea9aee745127dd9967a6157
z1609958bc32b46539802b6d457b4aed0c3f5f4a737f96040ba292008ec11f06b354b9d03380ca8
zcdc0954cc4c3758455aa238235d880a02dd31de8f61e8c3f57b8d11d356cc57dbe4785e7c2e490
z6c9fa9a1a9013794d117fe42edced253ad870efde4246672035eb299731493a89b5a3d04eb6c3c
z6510145c07f3a052140c2a551e07cf9b9a5fab7d2c9042f2e1acf4a068250e2326a6dd5d4036c0
z2a0a23dbd0f73ab769dd503585f173577598dd9d2d4f92d28f0e5c282ce60cc43d5ccd374ea0fc
z118b37592ac095ff58b8bf15e238d5e88d5222adb0bb3fc6fc7a4ab5ddbc3b4fd0b5df85f00ff5
z24aac75d5f49b9112a0b97500c11bc7908577ac5034d9455b3f0247c7e241819357cb755b1c659
z87c2c2cfeb63edf63f5f602af66944a5481b2fca465784b669d0d3ec1818f529e0ec4080057306
zf3c3ebbb4b3cf5225d939fbe2d09ba8cf6e788905824d2a95a51e5ce407ef15d5c05600197258c
z98a2cab02151eb838fac20d2825d6fc0e20374e556dd73ddf45c6d18638d62cc283936887c778f
z52db8b795328e65a8fd776bd58b98444c2178caafea26447561186b1b07c95b22d7bd17d71cd25
zce6a4e1f1d1d274de3ff26b51e9c054c23c5cc549ff8aec417dbda44e01ccb8067a08011cb8e08
zf189cda3f5c6238901b357e584466c9db2719a81d42d90f734a3dcad07dce425ed987e4974eff5
ze97ce9b42af277a68ffceba8fc8a45d7b6fbed01721c40e8c3b0126b63da074324dc98cbdf0e39
z08a7397af3c6bf004918233d4edf8c674829f4b1feaec8043358551bf0e2f1ee4990ab425b4064
zb68a68a30901a709d41efaed3d6db0b8e89b6d52453099a5e7ecad6636df6cfb654b46de4cedb4
zcf5b7b446486912a284b2198f96d9ecceb89c19020599590600a8c35f7e8fe5c27a825ac9fe270
z95c066e7e1f4888edc3fda6e0a7748dcc48104f6bb21954473855a0b9baf07a61fd17c6ea90c16
z06ecbfa0ba41ee282a4e649ff7db8ce120f7b4c191e3f56853ae73af0acdbb3c77bb4821251fed
z9e222e09f7b19ea06a81eba63efd03c37a98ff5ad874a573fcc0d908175f5af967f560fb4c1066
ze3a2610954b867e5816cbf11beac9acd42d039d8838c15a76d465e0e27457b91c412956aa87ad8
zcf70b7e3d57800a7125cb5f9c9e7800e1e62cb802631ad747e1d1a9849ff12a971dfe67d2fc26f
zbc0cfc92ed1432c57d1b1f16aef9e4fd97fca4eb662a045e2b2ac9d85152fe16a75549ce8c4390
z1d1677244743bf2f1be7884a2a494478ad15e30c72a8bae0a8bd310f9c712038e1534636316140
z7f891eaa6402fcb1546cd47b283d1847f58bee7ec667905dc7540ed1fe63ffc8614cc0d2bc9339
zc7a9d9d14f222d9cca49f59964a5e536fb8ccac829c013732492c360d84f231687699d1f1fd771
z3d43b20f02d31ffff1979d624b242ea565e8b2e72af1d45d06c1c60ae4acee76bf2f54c668f1a8
z8ec40b072de6ad93c4b7593afef7473c875380c523f913b0b223f0bfda2071ddd26d5b2d793c2d
z76a05040e827772e27b0ed250d9f801dd6fd8f61e9b00b19a523311dca77cc150cf83eee590e88
z70ebdd22d6809dc43a03c6a8444689232a54f2a1a1fd4beefcee0bd57c7f33287a156da6ccb7d8
z5fd48149f97d9a0678beedd4db0ba61163ef438222494b115da87aeda283f21c4ffb09bbcd6d75
zed8fbd2c24210521be89400bfadd6bc76c0daea4b46b27b569fac7fd4c853d19a878d1b1fe4586
zb2a8b1c4093da4fdf3f2279b73e8acfe7bf5a5bbfbab50a262fc6a5da9753ceefb12ec0852252a
z42acfba9b0a3d798c0f9f5c0443881e17b7e9e2343defc74c77470a5ba7919ea31679f333ab638
z2fc24b633b71ad2b3958d9d50e8a8a8cf715df346efa66f0da452448457bc8dc43889a59abc705
zd06f20a1a3057512065b23ab04cbf7573855cc5f2855b0c1c4694e54e9eed1c2000a13177f2fb8
zefaefbcc563b71aab243c888fff3241cc696e429114c7aa22d3a07b972fcce05d86d1114e36992
zd64c44c0e5494f16eb3fb5ac3017870c27aef646d924bd6d8d971b2eef4043d6b3afb7792abca0
zd4fda7e374bb93872b231ed56cb93c32aaf89814855937c37708f467e7e6a07da12c35c25d5142
z72656b78f2d50b738dfc1a88cdedbcaefe87e5d9c87c8741f8039c78a89320909090eb7d884d21
z4ef13345c819f4431863575a57744d026ef45a4b67bcc194602212d73c23789b18bd4e4cc6c226
z17fe750b027d71fbc6144c7fb9e6e539fb7b8900668f4c0632223d730f29acb8b3fa90418fee56
zdb122fc725332bf6cfce44166cddaf11224a648e091b865c26089699eb9b9dfa78402db2b8af7d
zc1e9c334737599842b19783dc083cf830a2ba47209de8117e551cad8134ed52de544495f597e79
z2112092157d2e1451fe29226798bb4c720f2ea5aed5ce5d60fdb78b5b6c2f9ce5ab0f67736683a
ze98cefb0412db4b44e71cf01215ccd57557d5dfa8cf7092b01719604da198da6fdfb9e272ee86a
zd4323cae5892dae46cfd7ab5ed15771c7aac9118a30bd51e228b27dd5b24274dfc83fab3da2abf
zace1c1f1be5fb8301012b43884b4cae52f0869643a022b48d2f388a11355b2473d2fb7045982f4
z2dfd8190dc20c03cf4dbdb49028509b4a6b561f3c2314df5140cc20a32132a86f5a125893a4d64
z27143255a113cc6443fa778ff7ccea590cea50d4449f935e1b10bf9aa1ab767220c0f6253bb576
z0c4c5a6fc815b69312f34fffff51f1357e3d09454c6905df751316eeb0734d7902d1cdd7367976
zf936ef13801505a13416bb4bf8e7075d454d7d3fa73ed9fe0114d7fb066c3dc22dcba0ba7e215b
z48ca30836127685f1fdb643b341463b677c5323a30534057cca4a575aca4daecd15c030585c476
zf8bfc5661281943d859a538bc8119e54cc475641919e7de99a992cc81112227c706ed6db9aa6e7
z15ecb49850b3e458dd144267d6c13b9339536001977cd5f1cfa328dc1ad874ef07688654793048
z04a7efe344b67690ba9a24ce866f9d6d17856ee81630adc90cb4b16209e166dc5cfbeabf115d7c
z2d7322e2e8f6bf44d693fe815d48dd629a98289f5c01e274d9934f9af3ab1e623d6f76b8a1200c
z0baedb179a76c59848d0e66abf852f0c7e0288bc4cda532d9d4f50afa289a305a07a310be689f4
zb2469a89d0543f2d6f1bc971d477dfb6db35598594e6e8d8eaf3a78bc5989f8847392556a0f77d
z79df761fd699ad2f5fdd29cd56a13d741b50cdcbe0162c11734a9f63cdc7fc2c8831aaf11fc15d
z96c273f69aedb5435f79395bfe6ed7bb7036af141081605614b1ab1a2bb7b2af406bc31b1949fc
z3d3f7cc585974d411f575ad334974bc95e106a863acf854cf9e87c9a6a9d6a1449f84933eb6b37
zd562097d439ca5db397d4609313976dc7e83d610f4068e6f31bc3bae40c7cc1a49176e9940b08f
z472bb9a1b7c3b9d42c86207e98c36aa33867cc1ea1b807bf2fa842d9e16af8a8c0e18b6b96c46a
z739f4facd03ba69f0444cb24b74878b60351b9fb6e80d4daa538c23b2c661c129eebb684d425ce
z9d249e6239d793f2891b293a5399f7096dadab148c49b9b76b47cec1944bd014405ba7e0875299
z04384cb18e75fb29f82516cccf247ecc9ae02874ce3a3c77fa594802bd8153e7b164b090c038c5
zc351342e8174f230446fbbc6b6a3f6778d80ea44b4f8a8e520bc1e41d07ec0150e18ce2e36bf7b
z85726063ae3ea3df0c7f549b963a990ab8dfb67a95381fa948dc40475c5f87600f3f9310e676c5
zf8697d15037ee29c4ca14c340990b7f56c4512f5dd2a7ba22c604df686f723b9b6b9aed139ba0f
z38539ce8f355024982419dd93cc1b54f568c877efa0b7cbc50d8d2debc77e41155b330294d8050
z63b971dfdba0a5dec71f2ec9d12642e0b79d2a961685d709f17c7cbd3180ee6b2618cab81a06ab
z7825c8763c0f7aa2bc31455a92f07d5787f1e078afaa9f8641daa4e2c9572185b77be4c113a2d9
z69eaefdb5b46c96683f571e70a84f21a51fd6ca645c300793328cebd3fc3ecbd0d7828b2a61179
z02deed62417f49622aace1ebf81db3b051ecf82c3136241dacc89d24b6e1012d73d4c7cc596e24
zd443f8b3e369c8df0d44e85972956af4b59cd323465d7f6a48e8967acc647735e922a43817454f
z66b6e6045d8876cbabd2b1eeb0339941d14d3ac2f10f867e048c2003214d95b05025f5ff218fe3
zac21f4a5d9affc3049ec4ea317132fcdb229530a8dedd568a7cacfd84aa8f163d3d2486f459ee5
z2de76241b3f0ed652c61f724f004925e0406c30d5c5d89f3d5123ae68e365870f3877212733e19
z835df9eee5f28ecba93ab2f7bac5621c4449258cb50b9b6cd6267f474417b31eef3447245f02f2
zf283a80c1c535db7a9c228de8d0bc51277abb779ecc12c3a4bf15d5879457dbdc4de3d67ee7a7d
zf16d491066242a34927d35b6fa4e1f12922d1526615bf071f9bd3f8b1a96cd533cd6d1255d385e
zc6fa3d696c54b3f41d85c1156ed7372cea0f98dc2dbdade81a6ad7b1817159d564b6e43f88a78c
z6f4c292f15ecfb3af1f71f98dcfae166b4cbab38a8fb704f3aefda6793c1414695fd353f741221
z0919ffda3387669416c31ee90508ffbe287b61a732fdcea06703e3c6583a16dfcb71501175b440
zf1cd880a1c18349d6f97544b2f57d77cf7cef923783c5b52b2d3066b39e2bb70a64cb11577611d
z42408d46917c2dba7d5362032d764ed921b237503b8515185f66abfe84ce57e5dda5e6eee0a6a8
z33a77a5dc49002abd8fa6a4d72726d1348353fba5f73f45d54d5ef82f124c07ad330ebf7593550
zb171c4a648da2ded6f8b08f7909082542648c99f43a7890450bec23fd32bfe60ea92929946d368
z0bc205a4f83a961e5cbb328274425a16ac22b1ac741f833da6fe4711f25af645e59877ea84ad45
z723020953073770905960dbabef27c1018dd18cb3a3c888d41eedf2db53ea250e68deeba8ffb57
zfaee96b25879718e12f8741871b4069d7457e6778420b7043efef0824b9ade7d23b9d697b99b91
z3914a019179fadbe80073e3480cb8867bc24e79481d6993354131785d459060a6be918a8815640
z707a87f8b7cebd3e8269d751d57f24315871313d13c67061e9ceb14736ff1430a3b5f2804f05a7
z1ea595e9d3b6c7c1a0539080759af549866f6d0e0594d94605191768522db16bf6453f9f06091d
z515d998d67e4fc70b2ea6ccecc3e4d3bd83fb250f2b604d380a5a753d88244210fa54243eb983a
z4b66eed3f068bf32b505f7639fd86e4094e3e6df1dfa1322a92bf15381685e439f8e0aa8bc6bc2
z8a82af67adf1c7328034aaa076c5d266b986d1a4bae64d1ad4aac4cd572d0569a5c00f0c500bd7
z8aeb8836081e246e51025b884d3df3a2bc184d938f34d6b4ddebae2a41ee90b6c594ef126a861c
z96c77f9d88fe7f5256390e6e1ed11949b9889b1e5bfbdee213dbd14e4e266060f5dbb9e51eefb4
zfb1f74469b48ae8d7ea4e5b1a4ee0e7ffe6a3e513695182483604ad9ea389657d6c473e90b7bd2
zd082091f03644a7e3cbf80c1d7fe094b20f1aa6dd43d29bd3af706f10a23ff3a28966c599b6aee
z4baac7844b35627b529a2319110eb9c58efe5936b936901bbc63d913dd88a6fa45e8599417dd1e
z64d1f45e31762cad0accb9f4165f8110ef8e01fd2cf4b49fb820c62cd220e40093f73707f27b79
z3112c1ab45c2540f4881162d5f177642a1571f7b42c77199ef6ef1cd1ac9c43613dedf9691e416
z8298565df7d9aae72223613a28556db6e9b0d6c07b66b4bd5a9137bcead2baaa48697415641cc8
z85d619dc60d0758508ed116b42646d6c75fe2fe0ff42c596d937d58cf3312606016a10c2fc0f12
zabf79c77229b7a72451ed0333d9a3c624eb185c070d5e7bd7711dd1bef053d7f739e0f53ea0656
zd3d033aeadadf1e1422de7269fc9651d7a18c2887280ee3a76000360c8b028427643b65bb60025
za2eb40563a6b3925fcb3e96cf42df56e0229bf3c0b901753bc788a09720cad80507d8eb969c799
zccf274c40aa70e126291166f669704ffc305fe5cf10ee8f816f0341850651ea7801d8791b3ca51
zf63ebe032426e555846c5bf30b0f1d4d6d9e710114c89c8f2d549d774e8f2ca3edc2b0f270eb7f
zf57fa9d9f5c41af8c1f779755cb650222b473a722808db147408c7f0f5470bb97f1c1a9ed9c13e
z620bfc534fd0b2ea263093168a621e380dd4152f62436638f8256fcc8c11821fb79ca015b65f8f
za33fe12d7e0d493503d00c65dcd1e79485a4cd4c5dfb988536ccf2459f605b2fb763a049a26b14
z054f3d4cf5be609c296fe46cc43c1097869529cb486746946abbf4a771fb8fc380c30534302b7d
zea1c0eddd0a5a73bf04311735d8609efbf23745574fb1bdf9055932681c3f3626dd4662954b762
z882a278703bc41cf247e5d27d7e15642d430c2d8a4620ca027dc3ee93038ee9f13559734029286
zaad9a38be790d90624cad3652f9e0dce45b15fbcb8cbd9adc3937376313b894a591b87604ee41a
zd45abc9966dc649c1d84af8af304a6d343afff7346455c838b1bc09a70e711024f30eb3574cb0d
zb83e5f89d5a41dc5093714c9ce7fed7d1c5b93396fdc5fac51a1aa97c25b8ca78d5b8053fff204
z8b08c50c726434d8472d1d6e70d0dfafc05d8e22b5291ef20d5c2ff643086d15c34ad52359fbaa
z6e7fca63d46ccce0628ac5490cca2e423bdaa5bf411e37e02a9e59ffdd005bbcb06a80a2aa37da
z9d3393eb063cfcff3611517a434af9f631714e044cd92b4c08d3c16f64817f43e77d07a96ef1bd
z13ed88e4e86833ea683ed0b3e2677f0eb18e293284b450f8defff3cbf3ecb099bd6d87f4f20372
z65d4b2a407eb481919811825a4b1f7c794ec7a3f400021b1914d042e10254eba21bdd36bd5514b
zc4699f23eba790abfa2b34c6736911399f75a8c3847f46fb1b6b35184d359c3f0324d7debca272
z7658d65198dbae0066f06520eeeb4ce850c7d08d87dde912beb3cc21a7477b744fac519e44f5f5
z9a8a96439cdcd2232e88480cb7e3726b06124d98d17ff9cc6200df1a88496040ef1ef5de2ac1f3
z46c726cfd33c071fa568d33336a6bad3bfa4d0a8d333e7ee7dce9262876de2e63680d42a24987b
z581ebd51a53f108d58216d79e5621081b7df357e8d5a1c80ed00936c3c823d09522db657aec400
z1d6993d442f8dbe56ad0f9e8579a42391aead4f02fe00fe578374afe693e24ba862c63cacb10df
z03a87895d9a949312878823e6913546c15bf468c6819dd17bac2bfa0a22e84482bbd8bbaaea3bf
z5a9bba73317ce688ec3dbdf7d1c8f1d572188d0f90cc7d88f6142e4c8223d058b478a50b098a15
z24c21fec6c842ce4b7fb52a03631790713d1c3f380051261d21cc6ab76da86cc5880699508380a
z966112d70f017b7eb92f483439ca4b1d6147e450a92391c27df64cb5af34d4e7d0eda1ed380a47
zef16273dbb8ec892862cbbac702f5b521a91154f61bcb190c6b17958672816bdacbbf919fa7843
z8e6e5914e2f8afce354579356722cd4772e38bc3bc552fbe6a858d248ca83078a68db1c0159f89
zd58993b66cb0f579511484bd04b68c9efe42419507e042b26c3715e6184d3892ed5c82c987147e
z6fece2e86839b8c25076a152e5415600f232c845811b13b5487f65a5289d5809ebed40baabe2ca
zc5cf06bc4b48ba2cdd974619dd0401ede85188026374b52a51f387e0eda649f89d3261c6f74f65
z0006781f3e282d973cb2b1c7ce891bdd4465c465ee579bc5de09ca43c744cf240306f76f5783e7
z0a7abd160016cf65b99028135e51b72a036ab7b97020d8d3c4746a96cd4c17eb05c2ec306b3de1
z0424a54bf1e07115fa007625cc7ab21f10fecee3ace436aba272a9acf9f0ca45bac737f92fd124
zd8f9961f7361f87f23b638b450fe86c2742bea7bedbad1a4553a839dd214da1d14a89e8b2d3197
z5deaa0a54fdc2c37e9122d3fe937af5750f4d78363f425a2cf40c3eb29d233a3a17f393e88b481
z75e1f27c0804adec499e7d11b149b179427b0a61845f09d89a23b3aae09c1ee877644f2d4414f4
z10ebde94e91ef9b8fae68548d9b77807b86fc9a7a46cc942759ab3bbe88f9ec6023ddd362e1532
z2cd61e85bc2336e2bc34b4e3b968b39f77a48b6b60f8fd630ca5f79c4866eb81cbe2380c4c5d98
z1764c10dbeb2eda9ad10eeb0b653735c21f58274e462886bc9f3beaab5b258ebe8b5aec849d798
z4c563e2d1f175fe99312007c37abb4ec3dbbb8731d75c61a1b97b4011f6da6c56b17ec06cee8a9
za4a1f7c3b1face3ac745f3b0aaea3a231b5aa36347c3a6358ac4a62b70bfc88aa6fa8378ae7125
zc9d7357e930459ccf85314b0a4bd6a84cdac034c19912090e4db9eab9c3cd611d05ff62faaf449
zf1b34b4b46e597e84791960e400a8673a6d444cae6ecf7bb49395f8a46793e7e528043e6049500
zc7384b0e9bc0e44606b9279dc4f58a900b5c802bfd3af95dadddf3f1324dd31ee559b0037dc3b4
z4fdcaf85338b156c48acd5ff97a9363693caecdd682fb2d0ba2df3f738b61de38afdccb0528da5
z6d9299c3b1397ee2fbb4c30e661e6d9badccdd3f60c8241b34165a7afb3e320f01ca98a5ff544f
z943adbafe0f1104e838bcb22f7aa03af53fe7b607a88e6da2b826f704cd85fd9f9330f9d201fe0
ze9a1581a6659576673355cf593bd263aef71b0a157ba82349c3164d39399494397def411d1c627
z071c0902da20c77fa82c997412f125cb3589a20af825ecdcfa9a0399708b2b24b7aeca92bff2ff
zc233a0d271a563212d4475322041946a43b7cad3d2ad0f7b4b922ac87647010937884412b48333
z709cf5a51a1e4c4e728f50ea899bd094d2a57ba2226e9d2cef0baaaf9b33de6994120d295f3f7c
z94e1515bc015ecbb0d8f12ef67684e479e5a670e6aac9db861ccf34db35e507797c3dbdde3ca91
zcf9fa1ca6f0223d40ca4101d6e25110a93dfca3b68a979eb0201587c4de3a608e0b97781ba9107
z1ebc90418d4b254dac2f38c893e63cd1a17d107c450cd8d210f64dc5f5f4e9c0787ad4803dc8e7
z350d64beb720199c3a0fb1b6ea4ba5edd14200b489b8179e06f8a8206f9e291d7311d16770e6f1
z22b4170f576552ce829b0570bebfd638f8107078aec4d50c58b508459d58bfc4f8b360290c8e4b
z49ced5e2fb2dbe7d803c878e77e2c018f3cf3538a9e0d914e99a4177b537fd704077000c82a57d
ze8297e00ea332e17393a6194b72ab1a34d3c437cc8ab336440d0f2183539f4f32b4f375b1c657b
zeac7d1a98e0d1e2116acf552dac52e8041bf8eb169e5def28f035c377def31387826f0910af009
ze01ce22fcbbba880dcbb8cf962639f803e02d5b3c7c56cbc6c67d4331b17153f6c1274fe5b5ee7
z7c49633418c2a5839ff93842384df7f7d4130fbdb0a7cca8c76ffaa086ef7be9601b26f6fb8dab
z4ea2c9906ddaf278e60cf6fea73e5c0335fcda49cbf10b511222a7efd3d6875c18b3d10fe623cb
z9710b4695d2149ad5b2d936532fad05f39a32e61c8d5ae662728b5b6243e7f3ff063fba71d64c6
z55682be96c00a9cdb81e7858f7296910f9e5847bcdb9a0fbb1b55041a6b5d6e460a1359421585e
zbe7e48cedba2d07e88ccc1bd845444b8cd456f0cda10ce7258e7cf4ef7d789ba632fde1fec9f02
ze8455e1d99ccd65ea1e0585642a8bca624de67575c491764871fe29c95337dc2aead074af0faa2
z9a35927482ce5a69b0d2b61e8f0facb5d6f398d8c858088ef90bb23d0bcf44dd4ece69691e6c04
z295e78bf7ba9f2441e5d444d0c3d153bb14f4d5400310ab8f33ba35341fb9563753d4dc1e7c956
zccd4678a07b3e6b19b122334b2d966186b346a41a7677af261c95777777b052f84a8f663315579
z386a25dce82e0982c5e5bfba43d1b4369d7297a0b49d3d7d844bef3a7ffbd51d8feade4dc33445
ze110e0eb8775b23015c0f103198ab0bd92b46c15a94af7d4ab6d8a8dfe66fcb4e8f6d93d103201
za77fa776c593fc18e8051338863ce78ea24a1400d3c2d2f877bd473924ceebb07a7e7665af619f
z5788ad6461091d41822d4c1132234aff779f42c6ee308ea0c2dbda62c6e2e3cbd74bd6e45dd924
zab671156c0cb3c5d8d2ca4e9a250a3d9274090112b44ecdc1f091191c3ec38bb326cda7237537b
z0401603639232c8413f4192ce292ef4966066f7cd1e6d20e92d33020ca0555bbdf525d79d55d7a
z94ae637f5dc55e0ca870e744f25adc0fe3c03317a6c94766dcb65c6e2fda91c011b1c3f1e40bba
zc6218e14782ebf94c4db99f35bd20f80f88967ef334f6485233c6bf1cd53328168169830998490
zd56e9ec2bb5448a518b11c43faea20c97fd71d8b72ffd31d4950398b73589329dd378fd1d01fc4
zeb1135bacc1bf435ddec8ea4bc0325ce4c62a5a3f69e5bb0774faac31a9f4d9dc1bbdaa04601e3
z3645dadda52a268eeb7f2539061a151a9aca604fa8bff1eaca42a14d51333ddcb2eadd66ed6d26
zbd53ab431432baab1a02ab47878d58f26dbfa26d62ca0608016acd0829931ef3cd7a8d7449cb82
zf30fc0e94fb0ddce3076a044cf13b7146a4ba7a31133e1827f7928011e53d5514b9dd6756d93f0
z5f61b40b0fa7fb21d405980c17a18f29edfa9d90ee597b92e8cd0e40bbde733592741a87f7d0ea
ze9f3a1277c9c63819220599dc6751bc56517323951dda32c43b72b2545e95f3656edb65800134f
z377c30eecdd98a29f5362cfaa11aa90440e76d01ede1089734f41aad3d02d5a26ca5809fd6bbe0
z5a112bd58389e994336b21cc7b492edc65fc64a48f6da961d0567bc2c69c0df2ca1e9e7eb8905b
zf96a8807c88245e0e7dfd767ace563095534c7a60eaaf98326ef18a69a66a978dee515c26722f8
z4591446338cc10b202eca68804275e2af18cd95229f282c66d3594fd71bc50f70f6aa65e2b48a4
z3eea6a7520593cdbbda7c0b75b696a46303996b35897bd710b2b94490864375b9d9b26353a0845
zbc841782e0ac6a2db5eab63b26654e9c8425595f29437d285c5f6deabf2a532f7287adcc0834ba
z1d57c8c41af80837f52807023fe47647927b135929d32ddb19d3e42691ea1678b48d73820f71a2
zdfe1732f4fc133e09bf1d223aa381917aa1c0b8e9eb3c5c52ea305a2a9346b994a9acd2be60eb2
zfc0ef806090a2853d8f846e94c50894ce898140c53ebfdf7975943e8e87e36415d3fa4a27facbd
zd3719d537df8d9c2f66eea4e184eceae593cf7e532aed59bca6c138ebb551bce8f50fba0bc523e
z937a1cf526816edc7ae2a79f18bfb326300dbde65d627c2508704b4e4d4dacffb4bd04e3acd20e
z1fa036739222b985300740825ec0d3085d60d460f82a1b0bc5aa1f89dc1217abe39d74792cdc26
zb6050e8ab5c177d745761be6f84d1e29fc48ef8de8b7fc874e3e983f3f1e954525058c247b0a4c
z6e7785e3e8a13732c7e828a8011131ea57183c450ebf91244e91df2a47d41a2fe51e0224711d14
z721308eb0b81f42ee7a07faa15ee8053bb9c7bfa0a15d5e161172b9bb1794945e7b281a31c402d
z6eb02667768d88aa6c4de2909d21e0f09f8d28d488205bf1d38ce7ec48ec8bf6a550a490a93c4e
za129110f127ce41e7e16692a5455964afec1e7064784180975134362dc3185a37a33165330b05d
z105afc78a2b8b00f2fb88d2819b50cde0fe2af1f1332f97ec6c2580989d3f0663a65527533cd6c
z0d46c7ad8e6a29d7f8ea0b2ed34753cb288f80745f2e5a94400ecf829ef2998c491566e1073f5c
z327f7eea0f021ce1d3224671c971eff0ba7d2ee127d5657e64f6e018c18c4d5ca46e575e82038b
z0bdf5d0fb0972f1f1ff6e99ded23af80ec8b45144c733451b69dd8d87fec276081238106f670a5
z3e65ffe087383647dd17e79aa8747dbcfa13994a837496398ad2502672d15b5acaf4b1cf57a640
z1e84cf60c05fe96882c538351f42598e6401385d4299c06d535e370c7d96f1349c917b3166399b
ze516f0987c8eb57f7423dfbf5936130530cfb399538becd68144263370dcdea4aa34c2a7bb8095
zf9ef199790eb3c620e143471299154bd079897b41c235e4295a82e19cdfaebbad8d8480227033e
z2123472ef69877c7fc7b5c10bbdc9017c1514b2616cd0181b562d8cac65e078ce538e9aedda41a
z44f44660379fe4a757e12c2197de39229b486f228a9b86ed9a57df93605e4bf7661983d469f9d5
zb2a2637a206f9f01461c7ab9d8fec89fd40780ae5c6cc93430ba8a2f25d18dadd26da926b07107
z20aa80b945bd72bdba3713c318a79e3f00c962e04ad76f02dc717dc5d0ece69b72b12ea9a3ffd7
zfece6d623d0bcdf93983e7e638fb0ca6a1ca45c6a44678dbd28a1d55d04770cb3ddd156d0d7853
z8a961f7e5931ed776269b9cb38e1056412656d9c233344a0f19f99d1d75ed6ab4354c1b3a4332a
z52d50c533b4824311e6b8bb814624d60335d4e62ad7df3292ce817fccf73d9bd59009da5d906cd
z26555d82d0f327f279225cd836412678cdb7c722ebbba8fd3cb1d1d01738aca04ae6c04eb3496a
z42d4efbb521efa3e5934e9e3eb200bb6c15a4169dc457462c4da2ff9f2c4ab2a85093d99336dba
z2116cdbde771c1faeb335fc3aa924b16ba44e5f1bdf10daf7d3d5f5df3dee58d37fe842c3440c9
z63a275058f5484b84f9faea316f8c13cde9d237e5a2f7d3f4f3a8dde02f480b183e0fe1d91a911
z58f26522863eae54b2101030f26f6028f2a2266042baaf8b875168687728422d88762efca934c3
zc9d405b925b5524ce2acd3fd057cee904036441ee80255eb01a88821f305997e06186c3fbc6d2c
z5622d1df7006d21ec27434bc0e7a6af4bd7c40f538a963418136fcfcbf6eee993e00ed3776e8fe
ze147dcc463f404cbfa1daa759e4677a98b8e7550fd4170921f491f72dda919dd171640b964b09e
z078ae3f0acd0a43d1eb6a77f414bf02d442e26edc8ff0db4e9b986da394feb10c18a398fb3f958
z91ec606261acc0ab2a085d4bff0d2e98cd5c9311eb329af5b52dd7115fcde244245b79441129e6
z7daca98b3f419f3988e9436b5e4f621c491dba6014cd2d9458d689366f1abbbf72f50ac763c98a
z45365529cc962ab08a750ae5c74723c4848028f3e40f5c6806f877066792521c44ced5216a880d
zecb1adee34867d7621696226a2593f0558926a9945137ab8dce40756a5a6657e63aebad5451442
z8d83b59cdf5056671df5b29ec559fdd607aa0fef37bfbb023b68c1a0f956534edbf19da07af349
zab70ebbc3f0dd80f42adca5a3e1450ab472bcab660d13b4c7c7d1f98b6b05af4dcffa65bb514aa
z9cf774d3b453356e044e2f01dbba06fb5684d8100cb100e7b237e5caf7e4123624e7e12b01ba1d
za4761c444edcff12832c29079d1d3a1699067b559ae00e893de5613e7a979d387939e5a327a2df
z7f771018c65dd8cf89f9037b0532442ce22d9da0712f8d477c47df62ffc3663506936868afd2a7
z4c8e47246e7b3291bb056793f57fcdae96589ca0f11ef4b4a95331f8f3d8696e8e3aa8a62b4cfc
zd9b58c487161176b453946b4b205f65a6cbb1897fab23a8e7d0a9dfdd60b4a9375d31014653cd2
z929848f8add77258c12c29225985281600ad108ff8072202bf5be976dffb55ce89395d4160326c
z1bd8c6802d2489fbc45e45bd15a7bba39592adbd3497a94105fec584c7c09ae7e218272dd25a13
ze7d24e5dc531487df91ea13b1b2d00972a6e38de2a45c5aa47dafa622a6dae6604ce0d909723ec
zda074ad60030d5f2da8c0aa67fc7061bff23d531afe40a62e0947d6400a7e045cc7b90c340eb4a
z27ae6851748fe5f77698e943f18ff99207426db9026d69ec6369493a3613911e1af0ee750d4f4a
ze83cde9d9c8a21b48bccdd0f39ce01681ccb1295a1a8da131d034cd101a4fd9e84ce43b17e1124
z2b3af90e4071c1411bacb4e343c9a9f11dae659df1ad4f547b16b1852d126379bd14c1dc83ad4e
zeb08a14c9aa297ed426069c6203e03b04a964f4c134fb8ef37e3cc0690f6f63cf414c20070c29c
z6b85149ea4fc6422205cd5f25a97a7aa71aa73e26e56d631713873ad9669791ec08254277c8cf6
z8eb379376c3aa964e200263be43f92d9145a4199cf51dbdcded804ebcda86246852b817adc8122
z5efefbad4b5422f5ce4e6023e699b973e1e4dfb0be69667215c940838634c83952463462f905cd
z89a476dbd3ec257915b65be48064f6022b0e177781055cb56a7845b8bc2edbdcfcde7e3a288002
z2c7dd014623c6367078a74dece08d3ebacda47c2e8ee2b4bda26a5d5492ebf5c9a489d1be3a552
ze279cc0344ea99fd5a5c7e3f3c444ad55e26d09df993d3bedd20741d6dc4efceb6f836e6fceb29
zb8343c1ef202b754bdad26315b8c33be7055607b959c3cc12fd524a11891f039efd4fc0b12a9c4
z4e3beb8969c67231810e8f69c4d04b71952d2f2b97e63e8644a1a67fece0997c69f99ebe6b476c
zcf4e593d337521eca86baca1dca6513d3ec8640a7b725d5c0ede07d4ee675c5ce21c1c1fa22893
z47341a6967959185874429883df16eef0bb6515c79ec34c368ccda1808fe0fa2553fc150f88885
zd538e794e29b24e25b37664bdf71fffed6c13a3076fadcc676a00a838e8e6a8d74a2bcac252faa
z62ffffdd2184484446b3d06bd02455ebd224f4b5da51eab188173d5254784daec47d603b4b7112
zb0772eede2ba17fd9f2fb0cce209cba2437890c98aab7033e8169c8a9babb7b933e08201ade5ab
z2c0c34bcd1e8413deb9848a94dd0370db290408f5da3aff99fe4ad44f326e45204a0f87fde5774
z3d95be6c190939a029f9d80f25d1fb56167af0f74dffff3676c7a1a8f945f2edd75c364f2a9372
zff58a69861c54e8a8dc28ce0e2d8555aa9a1eaceedfde8dce54a0585977f87a7f7ae2749d4ab1d
z2d7088656a471ece75d66a193aed04bb9bc3b3db11df43e484bdcceea8b16a46bd5d69c6d1d139
z6642b7d335149547b559ae40c6ad19565af1c245d304949e6d951d7ce380b3c3a693ac1a2e01ae
z8f45063acde6a186335b284ae69cc520151cfd4ed1a0df3193cf41ebdad5824096f885bb21a556
z17581f462904d2a3c1c439831b7d739f20be2a853c578544020f97621eb7c0326ec0fc8bd29583
z441a685ae3431199dc3ae68eca117fddd69765977ac5771d5389bc6809e81cc4964f3f9436bb3b
z1ce5b03bc31a89a07ed6e13181b343ece133e193ca211f6a78936f9e9a1559508e7a6a112f0afc
zd7a69a9e472119b18e16e2bd262d5e09396dcd5b9641a20b48a47f82b337da2942703628bf33fb
z5bb22bc6bcc0e0d193518ee237aaccf6b9ad11d30309cd211e44c3fd2d7010c1763fd2b5b0c2d1
z05d2ff06643ba93f9a80f25f17db80c9ee736d465161c7782f8d137eb755dc30a8bd2c3429c508
z63b805a2f5919aeeecc83b7a04ebde34730a2de43ab5515197674bcdf07a085a9901ba5f225dcb
z35b8bcf3f1a0a2ff579dfd2ef7298e7614712dadd74dadb3cc3e994c8f12e47aba140686fc818e
zf0437fe6792a951d5f03fdb0f0bf87f66df9f71fa395ff48e3c2b5d36bcfedbb3c684cb1be41fa
z49217f8d7259e44d337bb7ffddf1f074485b40723c5c0279a7ea4171cbe88c08c8db528c023405
z8eb7285cdae2b87b24a414a197ed4b6698b0d1e7b68a8545a3b8c924cbe54847b5cf1f6fab6762
z56973270d4ee3cb75bd399bbf44cbe396931862f2de9d24061b533bea825acc5f79b321c84e455
zbd87fb809bf294fd6227951c6759995450dab555c79e871e409da9172ccb6febbcfba31f7751a8
z0347c9e32bc8b2f3516a9e3370222cc8c1b2fe7ad4bcaaefdc155705daf27edad0d11ef5bf27d2
z9c46c3de10d7575267a46986e2cdada6c6e7e4350267a7f2c5d625b071373fb97e2e718b19fc0b
z0822677c3a4f18f7af694ba3ef1a6be7728dbfd3cb5219e04289a0f64029492cbba0cff0892702
z0cf6027a14b96f1e112f2214bcf619a3e987f3a296ff3b8a1ae390b131ad47a4fa484d25b67ca7
z175b0e5b7051a474a63550b64b94943b97689d60753ae320aa49350091b55b804916ed97a582d4
z33df5d75ecf10db7c9845fdbbeb68d124a77750f58176ff45331febf7dc1bb779a682e04615a2f
zafae7af871f3ac86ede189686cb29791ad51ad19780671cf35e0153938154575aad6eed174141d
z8d1c54730bf26dba0648c26feee181c466ca5a3fa8a4fe1b32021c238a0216162d745774696a5d
za178d9c2aff6ecc83edf9db1af69f7111606e350f65f88a2c7cab00c8bddfe10e98359398af6d3
z8fb8c14d4856502bc12e303a7b9e9b6b66727769acb8bda27fc6ac3c2b69af26dbd5ca3881944e
z5f02abd9ef84985d25d6442ec79f2461a980a3f4e0d4128493b9390f00699443ffb0550efd9275
z6858fc19a942ce15d88a0bf5fd2f71aac56e531f4d5d477da040836fe809d5ca0f5214438000f9
z9c0de25cb83e9d6769b909e8c2b86c353d59ffc327080cba0ac01a78ae106d35197d2cf05b3c59
z265cf7b2ef15fb9e09b58a9e26fc9f6aa977944f383180748a05fe23b99c206a789aa78bdaff61
z20d24d821824874507cdea775d29a42e34a48cef4be53b9e9444e3b666311e00b67bd4c374bc35
z06be31b0c9637740bacf85ef2668424082ea48a353f1ef340f0ad79549ae5b4eaa037f58e699db
z48e34af196ee80ad441057af110b7e3109bba0318b52184d9a92c0e45383ca46487fd2bb2881cc
zbd537b9e3a52c85eecc871546042dd3b053cbe385995deaac9f438b8cf33447bb4367d705d67a5
z65d9a8468e3c23ffa4c9ee9cbadb22b4ce3b54a563221bbce0928fbb3f34d561fb6ea61b48113e
z3106a4b5cbf6fb74e4b04ac79fc77933cd038f5cf3448c2e225182803ef941d371d470ab708b49
z3cd283302da6720040e076d665d0ea8e22a7031181df787b40e090879142446083a6d7a9b785a8
z1887a53eb45ad3b78a8fb2d5d59279b07370b943828889080d28b283a6e0ce452e977f1a5a3c37
z47055426b2c44108fefe06fbf6aa3ea605402a97c6a6982b771eb4da6f318d40e593103fd6d7f4
zd7110a57ea99e6831b298450ecb1d86bc27f8db530017117d7f4b02c32cf4591a77c945702170f
zf0c2d58ba3be2007126f3f8e296784181bf148fa1d167fe79d4feed2d25dab3b52f4f953c96688
za0d1430c94d7b33aaf413d9fb913a6d6c4f27db26a6569c3dae0e06d894ab3d7a6f7f6ab22ae61
zc043524781d2f3f6d6605d8d56d732ad3ef75f4e59cf6383e20f504a7d27111c9217f63565d5bb
z2fe4b27148fc22139161b91098fb056b71a28568fc87a75d28a3244ea8eab9e9d012c950455267
z03330732b9518c112ac45d6e8775d7ed0ea1035ca605e2ea1c27d9c6acce1f7baf11ca9ab30757
ze01065ec02585db977aae2a08c65c8c83f26537f0cd896d428bfeef05fe2c96764cee3a9916133
zc08a862f6f2b2f2a57375554e73f1a670b40e314a43f6dbbbce420c41064a8b38834b0b11f860f
z3128cdfaa8e5f631ef0741efce76c07b80d38ded741bcb5c9de94fca6888f78142d07b818b461f
za16c618098445ce74aaf52422c328d700af39449884adee83fa8aedfe45bc7ac688ab8374c252d
ze53db6ebe9d4cc23196e77bfd8ec9f8b4b745c38049a238e9228824b6d70680c48d57084ed1320
z02e4102d4bec30191362be9d92daa62870f76454f8eccddc136a3e85ff8a17ed969ae9e19f39b3
z06f1f667f5a5beaf0212ed743b5529a315ae7590b21960fc434996c2fbe939147773c644140347
z28b5d604f81e36d4e725d5843874f082c76a31c5c5b8ef68c2983243a99805b7662b8e14e98b6a
z3b7447ab95c10c3dbb3af3bc655e8dc1641e67eea18d72fd9685219f1453fb231d66695d7740d0
ze203ce127a99005c96c1da924c0d2e51e3a74f01bc82e8b4cdbfed898e9a74053021bd08f7e3d7
za7c47474e60a314aff9457c605d3c3ba064cd1878aa4dee3cfddcdb054abc537094e5a6f60f7f0
zc05c8ba52540632f6d94a7375329fc5a2836cd27ddf3860b4edd7109ed52a367a3f2720f8fb5a5
z5ba80172a8907fed63cd50011c426f388f2a22978845c9ed67e99007f34484ed06e98c2bfa0163
z1e49538484083d88cd447aa48be9514fb3fe57362fa25e136e6850bbd1926577d5b7407fda24a3
z07e8bde98319b38a4bf3f5cf7b5084e231f34c647a47b5ae74f13c6b18e5746a580dbf3201233b
z88ce14bf3551141b7e8e916015d641e14eb15995aacf0fa75d49b7c32965fbd91b279f64dc6601
z627fe62398ea1f6e4cd21b6b1a1c6885aa4b7288814ad22e94415fb3a28d04c0f1b70fdd8ed4f9
z8e1f49f69e33a947c960c480b4098b7455d5ebfd3ffb679d4c96ad0a2f7573c1a26d857d448273
z5d59030ff86c249846a025feb2489a68638e180a71f99766c547264ee4438270f15d0c6e3f5c06
z00690f500ace7bf611fd16252a740d745893ae41be19cc457c75a95fcfbab0464934830a851797
ze7221aafabaeb8ef15a382a726ce53549825fa7ba555d3c2d875dad725cea8ba58ae74d5aa9462
zd6c14003937c76c8b13303775b55f76269c0883e3ea05392d02b1124d5102a2cf1ec4fedadbcc2
zca522408b2f64749205d500343092ba5e72b6fc202995fe88f3f604f68f8cf57b8476d92ccb023
z7b21e2c90138dcad3c6d27159cd7cabbb3239cf154fc5b93b9ea4e2e803bb622693e81ee98e684
zb490ad2d50526d40bae21c0ad17235393f4724b2023e9e7664dd178eaaf2cacd659e387e45801d
z34659319a065a0841b27f45f91fcdd2969d1275db9f2a58b851bf14a779b4406f13fe5e6894baf
zd589753c2735beb8c1a5d7607a2e88973dc0040f7c4a3a38b4bfe96bd7c3edaa165c85fd7506f3
zd8658e2d81d5205228c53605a42c8c720709ef7ad6e11910a9e3184d42eb3367ff4eec159b4802
z8cfc28a6d42554cefd1c51e51862d2049f70ee2358e8b9404cc85c26c0fca5e80560a3bc097e7b
z50d276eab3fe4d4898c7cbcfd239a44ba0232dbb335c99e9f68fdfcbe4b822cf70ec8e77900739
z96095ed66a0d5228464b6f2f75b2df78714e293f1a324a1e64ae1490eee04c8ba3e3db87c43f33
zd4a21b8f8d5a467578f4ed9b9a8ed2809d0c207a55a25c7c65a24a9f4e07528061690aac837ce6
z21179191912c967a17a02123304c0c28c5ba2e5543f9323f922d6acce0083a0bdb2cd4edbf1184
z782534bdc733fdbb6f58843641eb4278e53c6badfe2cef811ee3fb1f7761d57917dcd93a395f9e
z5a79547e71f1fdf502620a1a1c7cc94a4ed6ea05d2c05e94652e3903d9a0977c326cf5c6aa6b19
z8584be2296de9751435ef4ef0c9c3a86f8b2ccd799c81dbe258070a7f0a98e40f8ac5641d87dae
zd0ac03c6a222c349e9a99b4a075ea221ef79af9e2d9afdcf5e0633601789b1bb77433a23019fe0
zf2928a27b19bc838c1e94a157cf644e79d80c0eda76c28da1dd1ad04de6622021b0f8f50ffbf87
zc5857d4a978e7e9c1f24e16dc355cd601f47343a44918c69837a80e39fe0050573725360bfd873
z16c1f69fbb06eccb48a65ff2e1be01df06759595d8be544983c15a153cfddc4bdab63f5bed58b8
z268dd641cc964482329e38bd3333a2882559206b3c486a9db143ded74d6de45519089d04a35618
z5e96e801239ebc41ea5e433ee5535a4fd1fcaba1b7b7d9fc14f3bda3d508dc8c943010d8544dc8
z4a82bf117ce665011a8b40df5f77ac1de20980c95ef2e4b43238eff91bff22817e1ec7cce243f3
z19b61a8fae1959294740ba1b102d2dc31c22710a1073aabf09d2e3b6c6c095a05c621b76dbb978
z21a3440f74ad353b8a0e734a2dbba2aea30f243e87f9f61665acd4bbcf64a2bc0ea52aaacad6b2
zf2f5ee3082d9605301ee7f96b0b28aa0c37631280b64ff944acf619bb3d3c3194999f1db8703c3
z912c9af698de3ec496bce153b44651ce76dfa97e8427c5cd3dd0d92089a18d4903f2283bf68d4d
z064adb98af32cd5cad711461bc0ae3da0a0fb99ea32bec88405dbdd4aed0309fdc2de2657492d4
z7650f51326fea7c06ff094a6fb7e48a388b3fa6ee4f81c943302b51ab430c8ca086a0de5a1073e
z901efe29c009558b3c794b30248d2a6171316361b9bfcbc0914e5b2708a07f149b3707f57b5927
z3f9dc5369bf08a5b3ff4bac68d5f822a8ad4009cafb27e4bddbb9bc40ea06203cdfbd6ae12f38b
z7b7cfb557d3ba920dbae878394946cb15791ba096feb9a454dc8b55b2e64d7f40d495ef1dfa36a
z03e7e91730554304cec787b4c8c80e1c0b0c10af6103b045cbf16c2af08da30b819fae50b9fa4c
zb927b306950fa7d2377b3cb7c989292ab3fc5db179c4a7f6a6b3296d7412edbfdf644671364de2
z49afae89c0860c2b908dd1f109359a6b3ee9f6789ff444778f9bfbae2fc5bf64908071d0c7e1b5
zea2cbfd8c93f3accebbf70f0eba47674a8a7c25f511f60f4901321d0066664439ebafb94559b7e
z4acadee10005161c789f4eddcb222bff219f7264631f9307044d6fe3c03a42c20ae9dd0427a1ed
zc38bd18818cd2e06054257ad30c8fca39e421f729bb97daa24973cc56c24392cdc6f0f9b8b0cd3
z21228a36ad98063f36cd124e8375b8cd5e1d1a4d21ff3f93b3ffd80c1b10780b78b4f1ee87d31f
z697bd72a580bc580d5e790624388b19041fa5cb7df84f83b1eeb5952d1a84f700d89aecfd45cba
zdccd421205e9a7e0119869f5f0b8b79c0311a18f1e0aff4164c0cd20799d268800da7b338c70d7
z4e2bd740b22d82a1ad90a3910c398e1dcac0691b0f7e4be7066e676d421d2c50afdc9f8cb0c8b5
z03d31afe9659d78def4d6c74e6339b96dd714b722bf26fd11509991ce4b9c8edf27acdb382b5ea
zce879c56ef1ad0410f261f571b013a64c9840d5efda4ee1d6ddabbb328e528fa03aa91bc005dcd
zff60b37a2af094b25829309dceb04849d4168b322680714804ef9a55015ea0eac8bfe3e4b9087a
z7b17d58c96c85143d70161c71459d55fbd55d36741780410577d32db41c6f8b10b11f61db5aa5f
z5d943ee11b93bc1c2b341550fe82b7ce5b5125dd5c8ef50bb964e7574eeff69953f5dce4572399
zd21c93e82b5537252e4705339d229b52b5c6e7108d114a7c190be9a0e07e3441ed72c6382f814c
zce91433e3b0e45b2892ea24ddad9dedf85c7f4ecd1a8b5a56c1c3a3efa696fa76b6442cbfc2add
zbd8949400277cedb4ed174ceb53d96a282d24fca18d66a0608274d475e5f5056bed13322ef6116
z5dfa16dc63acc714bc96b8315cc86160855314e88e382165ec08d52a59d1b925ecb1b769ceb2bf
z7a3e7c6fb7824298331c1a8a3d087063adc7c308a54eb903edf84fcc37bbacb5c57097563f7800
z918ef9ca32dbadea840a7fe387a0779f7378c1d2e4a8c1341009d0ffae8d1ca371e3df800b1fa2
z564cbfda066520ff1bc346e88c41dbf1284954c90377a7a1243da0daf8dfbd5a79bbc24a08b609
ze3993bf6fca2448de4b6936145acbb677312f69d6148d8937a3a6c644e62c00cd0079e7cc549a6
zac91a1481009757872b0a2dad2d78d81fedb8a4e1c328ca0e15dbe2a4a5590eb735740121d4175
z06c601676f14c3ede8d922c84f9a5c9ab6999fb6c1df56f14d078b2ccfbc334c54c96a76300ebe
z63a10806f3bc2907ac1f39cc718850985d3b9ed8867a4b574610afdfa6d2fff861ba68e9000257
z890736505a08f15f4c1c1be89f10f0375024e9666b8c57be8af08e37c5ffef59a4586095a2f8ca
z5c04c9a3259a049890064a3ffb81a54c9c9e7d079350900dd901ab2b1de7181f22d478ba0322a0
zb71ad1fb77a859ad584c88e247b537a4c99b8d235dfae5735d68270d68c26cf0f0e14a55061756
z546cdceceb25d7d088a7474ce8e1f74b05fc8569039debc983e96fb2888c2def6f57463160ffd0
z44d7a4018d36f3dc02ec7b128623d2afc82c3b13f39b0813d71173348c903b9bc445e532a81449
z82120cfe7621f10c9ce72544a4a953b96ee88ab7e343cfbb864ae72a0b382e032f50440f008e0c
z830db8b5b54144dbbc31d8f2cfb88903d6757adacab35be94020f6f3dcc709d26e92b7921827be
zc9efb913bcfef03418b5b64a213caf2bfd9d19c2566f20ef46b98e4801c4257939a83cff66975d
z074cb3c60b075d816092b083824f067942c43d40b759842967672d022ab8af9eb6a0e2a8e0f013
zdc270a63d0d86536a699d595d4a1783d3a6a428e1a6bc8c6c5d863aacfb8619d1898188e49f627
z07b90918b70d38c1c363d64184d7e71583e959d59fbcfc0934e464b77b7d0966f83d2e17614a33
zc61da062b1f6cef3656d4053ebfdf874214701478e22ec6693a5d24f6c43839ee3ee3351cf0fa0
z157c56116182fd8e931c9702f6b325eed1c82af7f1342e16c09f8ad1b890df79d1b9a91237a0a9
z74dfbc3911cf93986b577473c5e267c0e62a676ad3f221285514f6d161f0e3812d482dffd876de
z16cc9f00c388cbc9242466e023953a01bbcd46d133de750b6b8181cd999e7cd0d16a6899499e25
zabe93d9617de6d6a5c548a62da0ae79bc173e03b4ad9cfde2ed90ec26f84d217a17d8780b947dc
zb4b880ddb4b4d4efd711b17d333c613e58b35a61c073dbfa95da10deb9748b9855e6513a3e388b
zc71468512e14e1f7541446f7ebc24072d24fa5efdcfb380011301743d97c9d97a356a897beeb06
z598a553876836e1ed3a9625d7ff8256488ae836b7d78fa62678bb456561519e560b7a6aec53b2a
z5155948568814d269df5625ba6b394a2e58b1213ca661693176d3e7e5a119eeb1ddb70f8afbe15
z8e074bb45e4affd376613c0ad8817029bb8a6f46e92396613955d0c6ae07794572b0c450513f3c
z67a0a0ec1e0f9c0c2f13ce1b969c01d0ebc49add4da80257770a0e3789e5222caa38324fb61093
zc6a1543596a44b5287eb16283bfbe8e0f74f000a14aa64b88044c5fc8d5a49c64a741e40ccae76
z589cd377807dc0c30ddb4a9a6af8a2e9d21185e10a8c7f9f93362342471193029a686f5de5d3e8
zd4065ef7739968931e64c9a52b220187b3f759840036d04c2f3b4cd4a01eefceab6107d32ff78b
z475b457c873ec8a4ca3fdbdb2647ad77ce2a9e9c5656380e4f1facd6400a56ed833b202e66b3ab
z1c5c3d7c3ca9cf325ca121580fb8caa9a2d798204075a6030e9129e5a95e660baf651fb6649f18
zb3ec2809cbece1691c875429559ed08bf8120ad486ffc6fc410f9957625d3857cc77585bfcc7fd
zc55f36025616fb78e79ae5d1080de12e6fc91251c8af7f747c58fee4898636f93c55bc0856f4f1
z035a2cff1847f3b7f2f95b85e2cf7e1fb3f39313701553c3f7ecad0214111bc6e8a92d4ea109b7
zce7ce8a67f4f2aa3a5c02e4762dc261e899279dccbc0e4b1c6ddae2298ba2ec399986c0189aede
z8e2c1b6b176982b929fee27a239989d243d6f3ee2a01da9f563bccc9f506a168ff8679639a307f
ze4506be0070847bc177c5c6268922ae2383eebcdcea5a0fbc7fc6443a832f5fa5eb5d3dc0ea1e5
ze4e77d2e2a350ed65da40a278d5046492fe40d30c29ab645b93b58dc16435d63e68bf27833c8e4
z3d6cd124a63146b51f9650684aff4e66739bb99384eaeab505016e5902998e848a2a3ef2397de6
z96dc0a50b6eb8fedf877363187122400e704c94bdf1317af61650d454d9e9506fe5dd377f59670
z9457500a5cbf7dbf9dd629126e6a8625593acc92943c919ccd552d9ad7c02d60cc2ddc88a9fcce
zdb3103e90659879bb19ea9b29ed202eaaafae90b876d50aa6c8fa3a529382628c689218b9b36f9
z4167fc6418a1c8bc87554b4f22b7f3c86ee329364b2eed07b527e2958fb0df2ca5d5a181e4a599
z6bfb53e2664e0b26bf6de8e861ee4311c8e230570db97bff2ba44467f9a65c631f96c93c5020a8
zf440d3cb809d2f0863478cc53be2f475f545610841449ffd909bc6e2bf75b5606338239239bf50
zff3c5dffe833cc89c7f5b25758240c2b73afe9f34b7e5a464605fb28377aee08c6dbd3b4a84895
zd105cbc24e2613571379ffac9fd1578a1289dac57f74722f65c3f3647ff2102aa99aa0a5d677a5
z9d57c8eed32dd185c4f435612057b6761956c6bc9f6c91339a3daa6fd40704424a366a5db7d758
z01d300549242478ceb406dda46eb53328025d2912db72084862ee4dcd282728f713138a9b3ad0d
zec8c301905fd1595b9738c0e8a9f05a13cac511903c9280f9cace083d6faf09013a6119ed015a3
z6d890967b3a23d26d34e8aa10a7f6f6c64b464901253205865833c2e6fc7a82e2790315d146c25
z05ac6c59ec8022c7d221670781c6910886ff297852d4824d42766bf819d3c319db527b004d67df
zf8c9e2c946a4a22547dbc26d33cbea7d8805f39ef4133576670f060170de3e98f50aa5beb90930
z4c6deca05ba3489903137f2aa8359f87ba32c75731cd5eb122c9905a6b43f6ade7f11bac49923d
zcf494819427cf9425db79fc84995c61d2142e8eccc544267a530450985a1341942bac83fd39b7e
zb45ebaeccedff56fa1ae3d40681c2e2ee5e17dfa4bba85afff8f38374a36597a12cc70881f23c5
ze168d903d93fbb3be2f224536d948b8a28da540f827b3a3fee9fbbeb3cba1433f75e652a32bf41
z286a87800fccd83d45c86b144b7a7ea667a5bcbc65e911f3fc4a1bc6327aea3464323f01105fe8
z7e5fb908cf534c46fe23f34e03cc645a72d1df0c25e98fe2616605b4fe37888767e59d72371655
zfa52ad2ab1da9208e4302edcd369d38872c9dae1d6d5f95688e9585f19779ba0727ab5354e3c48
z2a39120482b8765d62ad743967a3027005545ed19175eebf65b7ec6f79a97a4d03db61d1237429
zeb562cfd936bffe9e2ff114fb6cfa2424ce1365dde056e6608b2792f59244e6a3044f74f54956f
z37b2ea9537f0c53f3650aace7415acbc63ebccb7c879a664f3356038103881928ff5010bbf621b
ze5fb63dba961024a715d15bebe16a62e721085b55b588204308ba4100ba14e9feaad2570b3fffc
z6f0ab01c5a879f01179cbe231b3b2324c6b2a2ac395a019f7707a3efbfdfe118907dedac467952
z0657db3c757be241f6c619a4ebde642fdc9068c7ad020baa15d7bf9c27771b72b48574bec9e413
zaa090d91ce7c05f5d7506e2bba8c2e3d3758f8262d11a85bf2712e7a144076f2af55c459cfa296
za427cb553cbc8dd4530d8cfcf7952b7807ea0f37d05c03d0ff90eba5e7d43b4c571893c2de21e4
z68994383e149aeacaeb28b798ef33b8ff19c0d649e6f28b5c148254733ea2a2d38452af8723ec9
z7bbae151f030b8955c8c650b959998692607f1c89cc5c35a8f7ae6cc07ca7779f2dc30cf57c1ed
z14fd6741421bb4153b6c927242016a09cbc9b4de7262f1ddb1fe7b3dd1874ae8f870ef2ca8c7da
z7066b07b2882eabe03e11fa138e04897edb6d5f898a44d6d1894ae174a685b895af2e75adc5918
z355418e110b6863728bbd339178b2e6de62a39d10c91c390b16af5c56798dd879e1e6dac4096c4
z63be6f26933953861f87b09ecde945e736353450f71f70db2ae16d016b4dc43b3c731b8b5a92df
z5caab609217dfaf5c57cb8979f8a76a202e1ef4cdd141fb865976b5e21ca868ffc63221a69548b
z443e9bbb2a9ab45ba5270c4e329182e5fee4175b8b98de479af0d639bd20cdf7ab09d1d0384a3c
zf6e8b81050d49e88ca721f0141c2ca357e0cc2abbeb00a9b170dfe9dd76759331ea0d534c42336
z80385f0d95251ed25b1cbf926dd3d183c2cb4414a72cd1929ddce50615b01c1bf01d3d50cbae13
z5f609b1c31d4320347a7516a3cb0e94044c3e518cfa864ad2f6c17d25eadefe2c72d41dca6285e
z2fb8bf6abd7dcdd50128e5560d4d02638ca39d3adf4f793b1f1fd0447ad089010e2d8b0d73bf3f
z2f3d1cf043fc5b56677166f34f640c31e892a52dd5ff2c272f52c8b3c09e1e25fc142333c77c7e
z3392142331001f9eb5fa84be7a6d98a1a49167f78d90f653ca03c1c67802194fd0cf56e95cac0c
z5c4e7f2a1544a08e78635fb1ce67bc605dbe2812382f5a5583c735647af5f88d04b2e525d288ab
z7be6db333c4f7fd5bd8e3d3e5147222daa4cca958bb21aa413ccf5d33f8c2b41b44ebd69fd4472
z6065653d6dfaa31bf99cee16f74364e899b19bdabb34b190e139d314ff458b3b19c936d1dbcfaa
zb9bb53a691be52b58332c0c2befb7435710958e8e6ef3e44c56462dd2b89e6cfdd8eb9d561b2a6
z95ece13ba5cc67dd68cd42441d8f90575dee130acd6538eef53e26a41352de89ca652edf19c70d
zc90dd2281fc09554589385f2a3138dac314f990b591e46df5cb3e12fb2ec0c971ba8005d9f3e1b
ze47ccd55907fee0972b6f7ff9817a54ad9a6e221d102ac0dfd6a20b2e15e49bc88eee2112978f8
zf34685fa05209afa50a97240a3fe71ee91faca84405d120536a0ebe9cb01aef8618a3b923a26ba
zc9f5b278d4bc847d0bfbdd330a32d3f4305df0294e96b281f858a166acd67d6cef649fbf4cffdf
z0b3eecfbc89ec38275306187c83b9a3a6ce9c4190ce3d58ebf1bb923c46195e5024d50611348ac
z8db4aa56238033c568da71e8362302ce67af2d5a7050db878908079c680fa6fbcd53924e9ebe07
zc5fad35ffed1d89d23acccfb793f08457948c6d2159a02c2942d282e4758cce592c2517ee0da0e
zba24cc36f5ee404a45d052162e86beda394a8af473700715ee332ef1a6ecf88d57cbfb0d0bbbb7
z80d26489243bf147b5dda2d978c10c3d3e6a2b5b057054d0169fcb585844d7fb426e9810619805
z816e6c4f97424a03203f21fdfe0ef121155f78258f6ff9590d35b6aca82716aa49202bbae64b70
z2e6c90eb7e92215567fbc54818019680b02eb975c4ed52795fbc3cdd2ab24fa37eb16b8a92a9f1
zcf324c1e220687bec38fd19953b9a0c132acdf9b39db3f3f20cec08b43580a5ec8811115f7a628
ze937818246fda446b16646d6cc450879917081601f83dbbc222e21e0db0c37e354b9cc0c039c9a
z11f27a4627321c357128f162ad1b1659fcf963869f91accb866f07e3d4d9686a6148004dd5ec47
z32beebfe843b2549f4bf4b51b8bf8f84371c02b5fed33079dab8e3151154057d38d57c358d2f70
zbe301972a7e0c08bcbef510cb98f4581b3e5e2e0db621aa7364955097b3b5fc01bbcdfbfc1de2a
z6a62b72dcdd4a941ec218e0597783bc568d77c4f273ec516638e051d1b4ab8ffc3835932bf0d4b
za9e390c8dacb66828bd9dec1e9622d5814c5e8c83f671222999f0184c37cc1387f92c1074be20e
za761b4a5e634609d7490e0f91033ef42b96b8643e5876ea6d4822dd15119fbe913b65bdc4cadbf
z6f52d66b5b7fd52970087afbd560b42d87b0f0f0988353740459c20e2742e06c522af9d2494676
z25ca9cf23acb448242f70fe3e60e025fab6c3d10415743f6e3f96537388e6cf348370708ef1c6f
zf77941c75bac99910d8154bed5a0e0a5b612af05fea023696c15706c8b577132ea14b62ffc8b3a
zb90bbeffa7e24e0e38ab127c2d05dc147466107aa10bf8b72afb87c670b7d51a3d9d38f8e3236a
ze466604b5384de2c7dccab38e257b01c5e9dc236b590c7f89dce4a895bf8e7d5e94028692b51b7
z9eecc18d313bde9aaa05546ce01697d7491c0d366f0688fc8daa28d08be5c534e7b1d037069f8f
z6f3304bd8c4413c2e81c2a1f0c3efd4439b63514b9410000c59259b3db73dde168a75a2e8f9fca
z7e921d82c3db3de7f88e57771fa5716dd74ffc8b8e4f2d983180701027c37885bbb415b5c7a903
zaed7cbe51d21976a9ac446dd56ac741c5a1afb7db4ef07a3a2d2ace5e5a5216b53e284331589cd
z57d3043a4f67f4ce0cccacccfc9c5fcef073c19cd8997260a0f34bf4c714ac8ecc374c6bf385b5
z9170724bcfa90c5409bd013c8c7978cf54b494d36c7f5767f121dcb1a18d6c3da57c9ac980e2bf
zccf832ce0398c415b55b561bf505937e9fc0a2dfa395b0512d8953c51bb3be7110f0e9ab730028
za06f0b2015d5ded430ad174b7753f2d01e279d1c28631e1915660df3073177481742142aba1679
zfdb131fb5631cddae52a28e67b990ee741b1c840626503b1ea118cf3053afbdc015ece91a1c128
zb01f031d93338e1ae468819e98cfcd502926d611627a0865a48fd61d0c82e09f3971feb419c4cb
z025eead3f52d2950282ee160f786b5dcf91c763d9b6109ead9ce865771a18e12b9d594c40d119e
z2952bd06a270022bc8f32df575a51562c7f8eca2e03b54576af641a0e46b78315ae2a251729af1
z2a35ebdde8ff0b21e9bbd9bc3ae9de04736caa36a6b0cf2c8bf340ecd4f3cf86a94fbc2d2d8507
zd9ed679fac32db7f4cfb4c9b981170a62267a10422b9b9b7b32ddbc5329ad69b745b6ba5bcf8ad
zf22d1eea83278bbb21656f5ac6cb4328aaa9794d3650977306a0ca450e6d845b4619e3ec6c0add
z54b3b7cef211fe75177264d6b1f60abb81090e0f31259aa133c497502bef471f078431af5a843d
z2d210a5fdec25cd3435a9fda599a715cb66ffb07008c9b3d08e52d1b3a5400aca90f2bddadbf22
z6d5949d0973dc74576cc53b234a70c4e501365ea3f93e52e799157c323ffab5fa77f35d6e1894f
z3ceae4d5c73ace48f67aefd3c845b50759c768ba0644a85226fb16743f5125590a76d89ca08ed2
z9f73fa6b285e62ca416abed64e613f8a1fc3269bfe30277fee30a0829a48ad82d54d06ef253271
z51910af4ebb2bee0294517c2a88ffce6eea40ea336d8a571ac71d940016d875c6796a5b4ccf247
z4572fde9d22839c40349cd3978899e5ff7f3819ffab2c7cc6e1012c576bcea0f2f3ee5c94989b1
z1839019d806d95de191505be3adb5e600d3aa42ac15b48bb8c3d7b7df56027d63f768bf8de8456
z6e2ac9590a0db50892b20bcd0dd0a91378bf26d434ebd6746ab5ad108999e913bc797884889ce1
z882597ee519fcf7ca2f83bbfaef82c8836143e376c8d2395d0460e8128d0386aa39330d35e554e
z834bbb7554db13c515fbf26b8285d3c9ab51ef1d123176f932f7284559fe5050dbb5cb174e0771
z43ed8225646cd64636fc94936217623a5804b869996ce5ab74e645dc030ee53c48c1aa69fbfec5
zdfc153b3a20c8cc46bcd639aac54a58f11b41bdd783f022c9159a300160a01927059f83a58b77e
zd440f01ddbc0bc17feb9c540cefdeff1e0615bdfdd41b59bf608bb9bfb69415ebefa01b88988cd
zdc2993d600a99732305f0398c2d88e2864df5da2ef0c815e3e6a23332f2a935241721889ed4395
z643b5690c4a9798f78cdf2fadcff194396e0893050ce73a1eb04858d15f44e7ae36517d8e927e8
ze7b197e42270b82d63d1091d8d9fc614f48f050b2e595ba580eb23d0a496f02074320d1f20a3d6
z73b43a8e936a52a3750ac8736f9fb15391b7199baced0c8d4b1caf43990ffbfaf72846e31c599e
zba3bb7efa7bd234f3b556d61d8d7eb233b609be17409a48a2af2d108aa3180a3462eeeca97a588
z417de709e611aa36c0daa4f0ff23169958ce9559ad623a1fe504b78de25dc162c56dae95c37748
z9e93e1c0cfa11904f819d98840021d4540927e6c15fff59ba9b82ce19049f62f47d4f640d46782
z4d0e66c8700c44c4200b28495b09f15f0b8a155bec04a1e822d2fa88070bdaf2328b7ecd39bd24
z2b236303ef9666e43bbc874543cdac3860f6821e1150bb5330daddb470ac84754c1afda62b1b2e
z453c9194122445dd0ddb58b93b5a39341c3afdae025e716bac761986565de7618596a2b2744d27
zb77b9178db71f804717576ea6b72b3e05708ff963458dc23d2602382a9581e0681d74e53ad0587
zeaf25033ad462598f1c73b314421a84f98cba72ba3c7d376c8c0bd49515db634b7d101010ca1a9
z6783dcbc5fa865bc5df8fbf7076e1e1e43c2e127f650d749cd318658f7cdb77a94d092ebdf6b29
z8af4ff6eb5b27aecbb7fd242bc1dab3fb3fbf39dd5377962fe6764809e6cbc09d2b3005845dd80
z6be64918d0d280841037229d373ed731b1f6b92d0a0ad25b993c2a068918495bad08673e9792f3
z55b22850d056c5f7338c6f2a15cdeb025b8a21b0e5a12f094303812bd63d40ae011fc1a48851ba
z28e111466bf987665ad8c0170ba5d5401f39f0c63c62f533cdb3dad3fa4f8599a3c2167302a83a
z8e75f6837ccaed1243287f3301e8d5a7f483045317fe10c75b9e1b4fc3f30951710dae67313f9b
z6e15870644e7cbf343c630888a8bb39d77ede099e6d0686293dca1021e2fcb34a1c7f33c8a800b
z2d066a8e717996e2981f3ceab729499260babb4809d47d80acd75cfca46a381bc71a62a3613858
z23987362ed54fd349cb4ee80ac05046a3e2db17326e4c34397c96eefa05107886f1c4167529a9e
z588b55bb57bae4f6e7477f3703188b91758b203f44c7d0de844c8b9ed288310d4baa594427bad2
zc1bb14552baf6c9ddf3015c9f23c254731b615d162c0d300319b9d6e1eb2b668f8391694ebf188
z87e7d730720dc12cbea747e3eb0fb12dcd4340dd1d821e6c4b0fb525841e829cf7af887e1566a9
za6a7e8f9f1b254b8b003f396b35fea89604af6fcc98ab9326b374a622685d8cd67ed7de996bd57
zbb850321588f4fb2283ce7d4f9921f79120dd940a89ca1935e8b229ccaebce9be96d01acc837c4
ze346aa0b7be6b64386b7d2e69225acfa2a87dc8e1dad2812d7ae9fa69de50f926ad570853c8d00
z71d94f42070abba01699b1a4413324320d3ce3b2c17b52ae3fbc0e6171947c0f1e321e853ea50d
z5e235609a11448a2930f2aa69e030c45650cb74aec7cbe25ca9a0202f040ebc26beb13821db953
zaacfd92835e374f16ba2230f59c54a27e667096deae01193d4c651e96077a2a68a7b4b4d402860
zf20f9deb02b2ae91765d3c462f076d0e69c97f58c922b56e0b6e5580687f285a4d3837ba5ed0f2
zb3b27fd88962822c80e36eb630dca07f22e749afa85f1cde8465dea7d69317550bd1af3c21030e
z4d8edd38b531cebe298b273e8fad577b98ec11268f705f08bd41beb50a04ad4cf0cade0f3817cb
z98eed9401b5866c053c9feb6a9bd73a02de47abaf99d97433a56b631e69a865159798b8169521b
zb159146b9fbe17eec06396fb956241bc009aaad645cbeb534a331fa313a1dab37dd19d52c5fde5
z4bec5552bfb9d86fedd643cc27ccbe536b4a1cfa0b9fa85ef81438e13373963dcd91ffc30bb201
z722172389ddf03d384e955f502bedb53db683c00e7d2764a0dfcd3edc2681e7bc7b410d6770280
z8df04e434aa5fe354a7498e3272273fe196c80203b8f185b890e791a04734d7dd53c0c78c18f3f
zbaf5931b02e791328211b2f07994f93a0a99d7acc4096ea84c73cf264747c74daed163e89f0d55
zb1d64a00118123dc0e538ad7deec587b78cfa5ab83fbbffd436f59387faab475fa4c4ffae1b23e
z824a5073268bf9048d3b483fb5bc53a39982170eccc7bc1c14397aa268eed8d8c8e5086349df65
z33ad374a6e45081f89ee046ef577fcacc23adc2cc3bd7e6d6ae905d60e85866039b243e0cc635f
z0c1e879540f13a57cdae828e7ff091ef181fb01f5614872290b92902365e6a2fc51181e14753b4
zb45ce90f852bc4a313686fa8cf553ed21049a930197219b5710d794e282328a395e7ad2a0d2953
z2a5e29d6e4e647d159c4f024b05e992e76dab0a36845197ade0df39ec51c5250136d0e9938d9ab
ze05336f10b6bdc51af904541a136dd49b05357689572402e6a05770d1010d636e06bf030b8f8d6
zf7af489cd61dbe16be8f4182fd12c4779a9c47c47806dbdb55230a2fe596c694923b98e3553b33
zbbafcf379ea2d1f3ca105f4316e3a72b1e06d1419ef8cc2da1f6b5750332fabff9b9cf1dd7f071
z44ec98102bdf5f1ac3e9d7318c60c357fc01026007671d45fedc8035057afc3b005884e206a5f9
z8fe539a6a8d2f11041121479237d379afbd26a9a4b130b4f66e2865adf45104e30b29ee8add421
z4b92efa40b310e9f8bfe69c4fce75d54c79ade4714d415eae19a10b8c920f159000d149abdbdf5
zb0d4011b101435251c8ffcb81ab0638870494a6c378a451bc0053c7811fbd3709c0a170fc0edf3
z8fe44a979659253b6d7ac7933b05c60e726371ef5b4b32d709d9458b30f7206f0618fefc07511a
z6cc789599bb27b60b70bf26442cb3a8b04c45c350eb1f252284e6711e5f51ff25a4636301416e9
zf312258a18bd03aae409780b3b1d8e0323c7548311ce515262bddb0a54298d566df64e73ffd17f
z6e7b8e48ba505922cf7d396d5d656bc2f7c39ac24996dd1ca2b517076a3b121262ad297492fa59
zc7c254115d6c99c36372df5d9018ee147b8c59eb76006312d56c86d7944677d672c5810b33bf0b
z38684b108051291f0f6675481af29c94edbd44acf4a6c3ae80fa1951fb5a2e89a3de5b950d4512
z74a221f59a7ea47f132900fec7ea0c2e3e79b8ec2d412d06ef6d1e6b4bbd835827279976a44957
zf8821fcae1ffa8036a9448d7758fd0e0f5d4d26f21b480dba28c303c45b2be1fde94347533c024
z29ba1b56e20346f64f335793d1b6c9cb897ac069ebfc35c120ae3ddf8590432d6db33d1f751f25
z038a0c229314941c6d61218813990e5a073a734444c4e219fb960859657bbbe3531822cf9f1f39
zcd8226a6273b2d6be5c1ca74243c70c6738bf300e9bc16a923cbc2aee6bb057622e9fa68bcca1d
z0341364477fccf5e24b0ae646e8f5d649b1643064186b1f736e44d5b6d9fa7fc5029e35b52060e
zd1f4cd27c418f9aafba2c54dd232731e85870abac4de30138de2fc5fc3b5549a6e989d6b7f87fb
za1bef5decd4717ad64231cf2f6dbc4eb5e8f5f673ae7a755a8fe647a7ecf4d6081177d5f06fb09
zd769ab5daa9afcfa1c1f87063fef57d8402dd2a21c5e9ebca319ba1f533a3e6bbda5b36d6087c4
z190cc949bdc530cbfadb85b322b644cfd817df4ba3b95dcc4b822dddeee8a47eaa9c3f3491595a
z05c732f502cb0dcd754477a761bf889cad45d57b5f96612ee44ce30fb14184bb10111ea37d4ba4
z428213b22769a2ca7827017ae3d934e50a0c6cca67c59c1d4c5f9f77e058beedd73d81ab046231
z8c172fbfc073af65cca127991723ed4670397195c1ebb5e8de5f8fa1f3884355193ae2c100d9cf
zd0e5f8f78bfc8fe70a9d3a75c2f541bc20b3a67696d57c563e49c983d9dcb39058eed5c0c3db5b
zc8d810de50e8f4a424ef4edb0ae5380f37fbc585315f6399e16be43515163a9b55ac2dde360402
zb7ff3e657fe8fb4671309866924ffec61696db8983fce420a76c73ceb032919ba052ffd2709106
z8056320fb1284ea2bc33bbdacd9418a804048ced25a67af490fc415093c1257fc6fedef301d741
zc91dc8c2845b46947d4f33fa2f1e31aad5bd6cb47e6af77b2c9271cca3efe50919e9887b738666
z5de1d95230163bf6c567f067970afb1b0bbe59ece8f09e5ed81776175e7bb76ae5abed1a51cdf2
zde748ff50d87c90bda794b169c894444f0fc104f156dcb563e7e243bf3dc12e5025cc5d8a9b885
z12ce6407158f858d946587cc96c4f7cdce24d8632ff28632aac36467d3706198be86cfa1c4a1fd
z4a4505d3234f47ad9a7e84b73cce3a38dc14a1a6530969f68efd98ab8778de6ebfd72407907f8c
z57c75894ac0f7c06ff0ec0ac4b7a3a70a6d7055cdbc88023e7b11bd83cd50e9dd47ec3c88ce596
z89c2f2c985ee2fb74057cde07083e45cbd0b027da8c97a189a35c79a376f2b5ded8bf2a10c5ef4
z019572c2a513ccd9df135676f0bc53103ceaf3d8b247fff8d3785e1844daa09e9c499e1c6b6af0
z5b5ef073f46520b8ff886bd69205a11a469576937867595a63274eaf1c8a0fae1aaaa48f45d2ef
z0fbb6efcb9bb6634cf968056a8ad0e28a6cab438c45c19d5c224c459b0736d838796ab7dbc5398
zfdacaefabf92fe99e18f4adb04f35fca6f9ea89e3363ee45347b1679efa506f8e047243d9fa441
z320c90d7e0fabd02c469c1f46ad11aee6f452c43e9e97235d548359d9accb99cafa46d3af33107
z31f7c72c2a0513eee96294b4a7129376848be21dc3f28263e0f073e7efe14e6bf2ccd9d34517b1
zd6e99d4bfd8e2c07dd62c77b97b48812bc8ca21693fd467beed6d83a3f3ee4a7bcb5e19365ab59
zd2cccd2f197af90adc02f39e63714cda7fe0d02ecd980cd5f1e684cc5d4518e09026883850ebc6
zf905cd773d2fadad252a8437e37cadbcb0ee8da8b3b0cd6efaa21c7f66a5afd825960520fac480
zcbfb9b72006e854874dd0260df473a4eb8cada7ce85185553e8c688150e07976768bba022c4955
ze6ff886f4860ca1f0eeaef44f4e6207f536d86ee1925f6f1809eb68fe0782613c206cb1867c1d5
zecc9654bb8dd1ddffec51a72f01bb746b25de33071534e49f9d3ab6c4707b802a4deb9d375f535
z9eb173855058cf3a5afc5c5f2e6836284ac21bd114a7f85b76719152e0645e9ec13b904f7eea05
z44faf5058e4b960c889ab2b141da61b675facd66b74e1b9d550b8d8a1d8dc67519985a93471bbb
z57202fd1b78c2d123c84fb4b3289019483afc72c08ad93917a844862712c0c31fcb2d843af2991
zbf548174a1d4acccf66ea7c845bfa9958b92b5b82e65f4ea7cb6a0f60ebf272131e3e6973a2a50
z7880b10e77c5411fdefa789fe9e86ed035b0459da0565455464534d25340f7b7c9add11714d262
zc29f7a8a30dce850454bc725114c641e10b67f875178428efc0ec8bcb9e239056e770657642ba6
z4684cf5f1ca8bd57e0ab7d58a979e3ee8465888ae1831b36f99f45d44e91abc615b081136cbebd
zd4c577dcffac1a105d2d23c2643f0ef06b02fad83098f1f0056c9212139aece6d663f724354a7d
zedaa6539be0030308880710d59dc3de4e9c2f401dfdbebcff0e8f953a598a7371942e23e14e7ab
zda06e13a5a224790c52ea7c9849f419384af8cf4e846c1ff10361d5792b4199ab65577be727d02
zf43f882b72ffe3b5083e9c8e8c9fcc296c02ffdf6c2c9a1ac146a241076b8522f7010550abb148
z780365b1202d9c660404fa123fac54cb5ed6e5233bcd83e46c7d76a4a6d768b512c0b9c4ba5549
z40c9c7da1daff0cf3a387f03f7622a1a98ec4047ccf9cf430a7bdf2e548ffaf89bfff1ff99d485
z00d34513eced402b86c6c4700276a2abdbf0f6a7458827ae38a6355e0fd067e59817671f646ee1
zb08c2c846f12bd941c97739c8f551d52686861dfba34e70f0d4c30416e2b0c8f9dbc5b8b378341
z3a4d4d3bda8a3873e1db3f0312572f91d257393bebda48a869450d84c4a988ab9b4c3eb90c51c0
zcfcbdd6759a6a5c12a25b8c3286cc80b34586624571d7b92914b49a659146861405b8e6661b681
z874535f76db9691bbb69b3d5817416fe7a879b3d3ecfb482729a6dd8c879371532ffce74c592e8
z1769754054d7edd9e33a066e55e16737aa0f120910b1a3f7afd59a1e9fbc8feb50c7a08f54a869
z83154bd0182612d57c70be273d011a4da90ec70b9df54d17b4afbf1bd863c2d8b2a6d65a3e343e
z87c0ce112622087217d818fd5c34e926a64252a46f1c3b18cadf2e938d76fa217f5d34d3f89adb
zbd5a71b981f61ed74aa52ef5692ebf2577b1d772d7979c36d89f979a38ce5b8f3a2cf716fb4a0a
z3dcf13ce37a218979ca845d4de95fc19354d59407aa26b6cfac6082344b06c105bec349a6041e8
zf2dc126b10d634a0f6f183931c109cbc4a4c63ae379a9d1dc902a1fb0cc5e5534378977c5418a3
z35f2f7c174de689724c2bbae058b745e2d359908c2166667aff4148e7b6470da1e5dc72e016ba8
ze8409bdd98763abb810bf368454029b0edd0ac87a31c3fba3c58e4f31a505d69b14ede580be367
z2bfc211fdc49c8b3775d916709c4dede1df00a779db19f84b4150db6f32d3d95c0d81ea9bb9681
zc5b9ccf41c948b0019b46f5128747469355ea660c1ede16d16aca3cc67b4e3a2392ce8084ec3a0
zb7a554788f28f3a63d4a070b7362aac4103d1f7c1d15dc5d4c0f1d849cef224e065839b96dd32a
z5fc5e37d0b673699f2383d007550521a3479ec043f8a5b792a58a3a5546f94cab31ce789f6bc1d
z675f95818a8a1efb588cee49410c7f487f0926118b21e79ba786c9f99c2344936ad6352bb27d5e
z2d497975cb3e22adc98b269f09f1a4dfb9aff6c560e9a16262ce0f8c6036b24c0451bd8bf8e62d
z621814e5327e9448fd3afcd5c4dacdf753244649d094b86245197acdd341df921eef4961c28694
zcbfeccce94c61e5dbbf1db938bc75c097e074c72ea62241978b5510a34208046848542d19b8319
z3a0b31c548f472e71a51ba5f5fec4a8282aab5ebaaba25278d36c47d28f829f764e59361d7ac96
z3fe30983baa6e70c4c7d35f2e56ab2eb4bffe9b831a9a756faac94595144b22f05cc9ef1bae5c3
z0aaee72206177e5ac2238c7eabe8b27b2c812b04c73ea1eb12091d3ff0aa8afbbbe9798dc31f09
z71a578b3cade1eb37d7c7934494be097808680a11a19cfaceba53fcc8194118263a30310f715d1
zdf319b4afd786704153255ed056dd9aaaf1e079af2941b89ab9048c46354fe38554c936883c6ab
zdb26e2fbbd8ca3a5d46680b7a3a3f661942f22e018eea95822145b5c35ac5b15e4534215cf989e
ze5af14c81afabea3904ad252b8f7df8988bd67eac078f272c0ce83bc423d3e09af6c6b7f9ef36b
ze01fb97a9f5da5ef34ed7d089f4548dc3ac90d13f5e35c1e9b5d3b7fb2363c6b65e1876ca2503b
z9b7451da0ad373e6ad889fc2a0f6a8ce56e7b0514a51733ef8f4f85f8c7da4fc9a8d5b0c0306c0
zb19f3eaeda5b684e52539f368b433dc276c935dcd550cad9032d9f352c43b276d8300b71342860
z6b068ca383ad0b7097bff12a5fd2ad3cbc8e18865cc9e397c55a333ec13e64b101afd2616dca65
ze96fc5e761c54753ecf3ea4d2be561a66dcfdf2322600c155ba08443061ae0f318bb6ccf027f81
z7ecbc6ad547fc3ed445520708c4639bc30803cdc0be4b5c635ea80d105a5351f84bb75887eadaa
za96a471c33c782b99ab2e37e5c7c2c2ce2f7bfc1b9156cc152c9c916064990e0fc9d967fec7f20
zb9764e08716bc748e4619bb9f94ebcb2135d40342e904dc32872aec648706ab1acfeb29443f3b2
z64f26f83b3dd7452e5cd760c392ddab0ae62297980c1f2dda285069b429803d9aceb3512035a6a
z5aef01ef3294dc932da866a606b32d520b060f6e543c58b68fe4cd5193823aad70ef33bcb3acd4
z8eccabce8d7c51f5d208fbd4ec26ed078aecb40f07dfc4c1a453a19471a16a13127e95389b291c
zacc03794adca43c0e539b921b599d14d1519d99e12dd6709385a7fa48a4f8e72227030ebb2c51c
z97b54525d7bda91954ba845fb4e88fc91cc8f4142b26874530f98472ea378e4c61ff9881bc59b9
zd94a83fb0fc73bc6fa6cb2c1367f0c1041f4aac6b2962d887e98e88fdf3b59cacdd0a28199d878
z8012054b1011f46a64e350ab6f4ba64241ed8ed1c55d14773f5b2e1a08bc6ef49dcb9b32197727
z8c7a34f4a4f55da70da27a17356704eb01006497fb65e8e477f8ef0c1b40288ffa70a89ef25b8d
zd517db7dc0865c2f9e065493a4a10d931275b11d1b376ad0acf02dc2ad8aa273f58f780878a659
z084355616fc105f7df0e6f163b28ebd6e3bc01d1acc888517a7365e1095ab2da1143375579cbf0
z78b08e510ade4da6f79740441469cd49a4fab79a77f9e1d9111a48dab1dda1cf37e44e1542ee04
zd88d601ecbaa09b0b5c304732ab5613e91d9705b0573d744c8149372ba97d1d50e4b677195fbaa
z7125e33197ca6068ad67b0618e7f0af4d3d4354ad507767d895d44ebdd053c754676008db791e7
z4e7e14a04bf418a65c8878ccdb22370e9d221c30530886a5897db94f7d155fdcd905900270b1b0
z0c272f33713e7a75d60ce7ea4c02805e289384f92219defbfef763390c98d06d5caf48da808ae2
zb70858e408f1e92b42e802898ae5976ef6f96b0ba5b3f1b53e0f20eabf3803bed72c70ba226913
z118bd74bf0ed8fa91122579ece703756d87ddba7942fc9209343f863b390ea5ba44a3b2d9ef19e
zeb4e3dfe1647655a26167347993d5d4aafb9a9e2e18ed85f1c3c7461ebb29223f3652b03c9ac50
z7185b01759445619fec022084a7a712e4514867b4822232dc45e7a2b0020f51674f91b1881edb2
zfa9d3dd881f3798515461e502582efb0d8d2d70c89d427ba2ed6d4fe41c73117bbbe8f69cac589
z37449f092de9eb82f865c0ab1c0c325bf9804424cbbb54afdbce158a08da820539cdcb2b28315e
z9543a5299f760acdb4e8453046140b0a194df27d034fa1b811bc56d9a402733397b9b052e4e6b2
z7c6fb8b008065ad0e0f192b90a9f60a1a19720ba6c4712c5e5d93aee9fb63da652e1953a0e97e5
z5ec94091fb22119e4f93b05d5915f8d86815659a199971aaa02bbaf8803577a43979e8b5301a69
z387cfbacd6517589672c0f9778c1e30b68d2bd03e792ebe0a5e0bf2d2fd93bc71ab8eca6791463
z97089f1b2e7aca53c5d1a92d509629143f26b0602f4ceb1305f1aed32061d6530819eb0b748baf
z09099af4b09af9d34cade9955b0cadedacdf67d8f7bd44a657bf96fc15f1c9ba0c39a9792272fa
z5afd5902dd860297a762dcf0dc9da6a66e2b3ca4ba7484431a5bbe493bf8e369ffc51c20b85fce
z96d8ae1bc1fdf5109e6628044d7917dd38992b3617686acc99f09de6e178c61b7dedfce18786f4
ze22db41b0edca6b81a6ab9128b37b019eb9853df54c64d4e80c28b42058db1d72660457c268758
z5d8418a15e30fc7672d6ecb922bffc488ba8f6437dce3385270bb3b0c1ceedbab804bb6759b0a9
z180fcb8d53dbb6249e05266c5b3084f6b3b355d0a40e945907be5865e96b75c964b2f5bf1bdab9
z1a00848bf4a4b2ece2322543ebc355c2ef88ab61d37030d6b454843b5901bf50a0fd31b503cca7
z4a72d1ed8936e6c42aacf6584a927f7da0fc4665a5063d2616aeb7f3f67470a040d97d476d3e92
z8aebf0a6fe7a3eda601f243f3738532320394b76ff9c94c7f2cf4273f6b9fd2e288865e22beecf
zb6b55394eafd9e6731b32d6edccecc3596ed58c0d31f109a51731d05f85fbf65c1ce5266b13520
z9eab35b9320399f3304b94cd50a34ba520a14e98ce33bf789d128ffe049f183fa9338d57fe2f9e
za7c940fea534dc490c018939c71dbd48c3ef46f637fadcbba65988f1ec61f334f0908365a45358
zceb0a7a3659f64ab0b42f0e511773f8d93123f4f607a17c35c556563bd3808d85a2ca24e247f54
z9178ca80e42743d1645eac718141993ae6ef0543544b5de3f4edf04d3dadaa0fe5ca548e71bc71
z8bea3cda6d39e3ce0111cf37c3936b9426732ba382eb7ba5bf2bee8899f980179bf3713b9ed90a
z2fa2cee4b2f39694371c8d8dbadd17b8b228d51dc05fed8cb88209cfcea4ed70e8b578c5310f0c
z65b895fc47e386c74a03c217adb736a0839ab2c3b27071070677c3e1c2568ce5bffe3fc10d6e2a
za31a09c045cdb277069af2c8f3360aba5c0a783b1e15347f5fa96fcab48db0923605b6f6e10e20
za751657075206e7edb3d080e706d73bb1ebdee9e2dacd0df403e5bc7524bc56a2fce5785f316b3
zb42071f6133ee467042cd1b0e6ce935afb31373ef789264e49695c40dc5247e1d2aeb5210398d6
zb61697fe877ed4b91ab97de4ac4e813386c716efb6f8b7525fbbcd912e08267d29100ce0818cef
z2ac5dc76b3f58dfd853a3fa6c80fcbb8fd87f24b9e47261431d8a7dc351994d5091dc29080f1af
z45afa0978735001fbdc67ddd6896e019f4706968105e680fcc1f556cdf89cef58b4078674df096
za290e6735ca41bf8d63609f26a223c6eb423aa3fd17a0ff5b06efe6d88c73f615e00c62f0dd561
z16c56df31a13d2f753b584419702f0e78e15efab18b08d08424d5258a50aa8350722cd116718db
z7e969a100e0bf1e3b7b5ca06bdbc363f7c5cc279c6e02713ddb7f1d27938ce9881d95ee7172577
z52646398a333c62c38f3d5d419e6f41272c2f7fdd1d0e24a92ebe728f7eb91ee1c6af32f7b1860
zec26827cebc62a9e4d847532cbd26eb8180ae1a0612fce4bc1824452daf3fcb95c74ef1e838675
z112499d2a396676b0f1cb1ebce8b273f0ce3fe14bc3798a4856b5521bc220aac8a32f4e8453528
z7b84c6ac30b739c1bf115a242c2271e60a1ffa5c09e10b10752d849b7b9f2447dddca3cf87148c
z9f1c0498c3f06c9b0660629963f8dacf1b9675ebb311474f55a2e4c9b6a511711d85c47888059c
zd892496425de750eaa48a2af71d01fe0e22ee76fce98661b05797cb32b534c2cc6985e54671f09
zdb555d6c76d361a0d3d82d9ef4c273553c6fc086a5044e679111072839fb4c5cd20614d8e0dcf4
z833b9c601e5e51cd4e4bea0689d11e50850273ce74e5fdba9378c02e1ef8d6377d78b98fc2cfa4
z158c14503e2ac6e27ecf6534c06b793b44e6fb54ea24eaa495cbe3f2a8479db06f236071bc9161
z7e9d8496a11b160c82726b5b54272896f0c84ef46e305a145abfeacb0e49d0895caa785863c01b
zc453c454dae914631307d4f82276f2c6809ce1209ebd14075a45b065fb906d936a09562e7867c9
zb92e87ea9d07b73147203f3cc129a3a4763b8b539a8983f4e519e87e39f52e7d4d471b82fe536b
z00ea026f088e83f89501d3a8600c1bcec8abc7e31204628a60def9569493c2ee64d36355d4ba0f
zd33dd5417c7ae052c03a55b02637b747546d7b40004f010b8e399862f1aa8c518fdfba489f5c16
zeca9209c62d4a77a456d7336ffcb5d4041aee1aa084a6e57168a7097d676b8ee0fa5d55b05378c
zb118fa4c845c8d59962f7a28e041eb40d8d1569719a441b757d197cdc80e559c62b27179c6702f
zaadb44a16ea63a420e5cbe306c5e274a40dddcc293e20c8ca0200b74745e0104a4badef0ca21a3
z1862b2add1c409982bd29ead055879d5be165aaef55eaa491461bed5a1552825cc8b1e3e2a346c
zb6325610575ecd2e6ed67f93d273c187457342c70e1cfbf3d828c415fba17d03616014055c9651
ze1fbc51645c96778cff23ae5b69c022fe2f16a1394dd56e362c8e358e53eda0846b5d39a3e5f55
z8c5a5c3283b9de599a798f286c78cd313c564bb09f8b1623b4ec5069f81c65032794b30c8b888f
z88f31a52744fa555d84cdb410632ca75d69941e88c6dc5ff0ff0d708038224b3b8eceb1462e739
za4e23d4ae0ba54e4856ab69238b1165f14ca624223911ff054c80d7d4abc43b98354906e62c2d3
zd89bc0e826f45054e06118c2d17e2644f609662b39822a88a0ced1aec5e244ab94c9ae490addae
zf128948210a2f6aa74ba6fb6f771f26943b8b89c5e8590192de8bde64ca64dfc4cd801ff04a102
z5abfb96e4e53ee38c147495b3a6662735ad57b0c8824b5876c5012bebeb01f204b93cd2a269477
z21fe7f68921d91452da434b65f2238211e25604da935bd83cee256f23152bdfedd7ec95f4bc4ac
z6427569b6659d06c8e6b84b8f9c364efe718f8e1ed7a5691d711d8a32f3217155f54d565585329
z6cadf2e052e0991229da5efefc5b5b36bf2220c18c22e3ec9aac5377aad8cc61de93277a24d01b
za128bc039cd6aa058897149da14b4ab8e1de4d304e1159bffe97216f455ce5504b4700190683dd
z0f24297bf24ebd9d2e7e80747afa3a7eccdc31a6ba8daae633e8281a955257b685c61c46a12031
z90365cd4160342579c3169c04d3f2c2060493acfe0e3499d38366570b0e31473abce21318ad2d3
zda4c5bfc76414d3c7b57ec112e8144059594ad5ae76c252473c2a3ebfeaf5b55f2921bfca4ac91
z9ee191b008c92b6148de8c3c775eec8eef7910c116f35ff69764543a17f2948f86d57b0b2e48db
z203d6c007002a078e4dc3bb8692308ba044f3aa557b4d37350eb68ae39d7eb9aad2374f997933c
zacfc1e727749324f6bfd7ba8523681a8f6c42a9d53ea6f2c3a462fb2013fd5c9e57c0c60beebb3
z8f6acb749647a24c95e8ca32c45443e7eaf71ae10ff20a0bce342e7a08f0ed9ef8b4b5036b8474
z7e6ab1c052fbf608af4416deae4e73174c4290b1579197fa3a8ba64602dbf7b0a9dbd479ec599f
z3df8a6d7b5ea06ead9119131a4d8e67ee6b41467daedd75f81b77e4250b7edec5006385d7b07d8
ze8f277dae40cecb7d62be63ae3c20add93995b8561f43fa955f8b1b3f9c999c13da7a5599f73ac
z00767b21cef9cd874b1ddf73600f348ed5ea96f82bb3264c311e5fd74dd18150b41677a32c94c8
z8ff7af969d32b0ccb539e10d7d00559f25f58be21869eb60118a5f8a18fafab55149709c23ca3e
zf3b0eb260e334a38cb7572bfe9c6464ae7c6eca15b1c289c30a48045a8060f4a7f8f1a42d07a26
z43dac043491d2c1ed347b4a091c05cd749a340b43f05f6ead54a7f8fc7ec0a3611a6a13bff47bf
z26c24b9aee57f39cf4559d7d13eabc90fe66f01cb3998c7f0431a111202d1d8f4cb52bfd0e2d03
z1ebee501e3da8585c3c70cd5bb9379070b36063a48ed0fd760d4747cb3e3222ffc0cdd9a59c5a7
z93c462fda1629109be3743d9f9d8d0de28a28e00942fb9b86a27c062511c74bd55e99c69c26f56
z628c260c9542653037c2d86067aaf854a88a9f291de823dda0af31b6ecbe51a1edc52a32a59b23
zb7a7e084286925e458359f7c2f153d08856d67c62a178435ba71ee18f94d1902980bbdaf1e3178
z872ddf0abb03ef4fb1cd46b249f676781a93395b1a65933d02460d7228b416e0066b90cdec9c89
z5694487442e34f5b2000b21a4b5da227383736330b14555b467967f54c03fe5c8cf329d9208368
z9dec3cbe4666a67eac18be9a56e1601acd36ccf4c5a69e012bc19bc827a414a972edb80acab074
z06860a5cf0524afe0f7cf15d99173a17c526c8c7576c93afdc593640cf4a0f7764cad8e8704b3d
z646f5df14d94f3d5ad0aaea789dc8c9ab935f07a439da2f205f655740992536a6d6377e8484695
ze9c770e2aed101df171586ca0e1e0c6cfb68f2587164af186a5d1f3618ced33ff2b6c4b9e78648
ze114155c2182c267466544d2ea406d1393b405278319df0f4888e8e639b968118b35ae2e8c5aa4
z53751ac45b6291c42a9e9977f785e40c6579008b8a63cc4dbc2ed977aecca683218e6831d4ee93
z1ec44942dab5ad262a27336c8fdaed693bf46046233c859fe5049ebb2203953d37fb884aee8fcb
z747d2b17aa62a21d50bb257b5040c5fd3d6d4214aa2c8a567a20ae93dc46a16dd3ea334fef028d
z8592f076d2719f5d9880a2da70a1cad14b1520442fb664e0d24a1d69f7fa782c82eb46f588c6f5
z07f3d35bd007582a4ffdaa6d3dfd7b5d6259847ea2e2ed3417b691f4463375f2feb00c62c2f9eb
z4029a640f2c28e3ff362275c1ddd073db1fe3161a2d8b26c08de4e0104bf188a0da16cc07afb05
z736970364233d1cb14d9aad052b25d8077394f926a693087183fa8a19fb5963256f9125c23fa7b
z945bc8a48ef6ec052597529a3755eb0a2d321316cca1d83b0c967381a308065c5acd1bdfe12fc6
zd6fd44a538cc1e6bfddb27b98ad7230c8af821aea17ff538edff1c5e7869156dd67b85bf3c37de
zd4103a32a39b940f8c30d1d905cf20ef8e4eed54076940e4e6e9fea2b28967949838f7912b20cb
zbc70e1068583ac602f4fb3df81d7904c7aa7799662a1e06d65e9c86f676ddb85c16be35228aa53
ze364509154e3fb94c88a9e6af2596885269d1dd57393e67f23701a1ec06215e63eaaf4d8380053
zaca91cf728a3f82e283d12119682c479caf82307c42661d80b73a4fec7bb32a525030a138a2c3f
z3e5c06f19341685edc470ce9c6e61e8d4f677c1d68713ee11334e415521e972c8494f6733653ae
z7910c7dc74b6394ea8ab7de884f4157da4a507ce4d71dcdd0b0bf377d24a5558e2dbf713f21904
za3fcbe59d7f50f5c875f2ec5738c404d72aaddd983d77ef764045300f0439c4178a458272b31a2
zef7f9182350857830b19d2228b8fae4f6dd64a39d01656f5decdc58dbf5013ac6a4497a727b99f
z6f25a188b75cd9cdf2ee2cf80728dd932e69d9ab33bfac6b85ad03b75ed5ee90daf36638f73a77
ze416a4fdba9c0708098f15b516895414fc1550e4a086efd7edd97cb7e0d4b32fefdddf0e6e8518
zbca3f7a483d890c780ecf64cbac4bd420c1f6b290fadc303aad1141d54450bda64511de48312c4
z08b485d59862837eff5aca767a0ffe592493c5e7f635c2822d623d1c9bb3330797006bbed95e3b
zc5408c34eebadede908686c31fba8e4c84e5bce05172d60bcf39c22565a066fed92522af5d267b
zc3f9b8e6c91ec85d8a57cf01212c27141ff06941864f3764ff02c581bb814c20a35a43779f9a92
z35fd490f0ed625a31cfef4c72f597310e2f4a1face4d41bec05ccd183706363e1a89b332c8b258
z975c6d1c41b58d8963cf0a961753def1086ba86f7addfc082dd5dba28877ead31c3463b8eb5480
z313f83b4a93d24a37c3a1d4929cf5ca1fbe60dcf1a5fac0124d8afccbf658f1253e07bf210657c
z2ed696f9dc13f069d107ff961a70f92b93fdbcb48e6ca9cb419bc93ed28dfc37b7b8a77468133b
zf6e01d7f0a02dc06d0285436eea0da1163f50467e8ebfe7fb80283acf837b78827f29595e228f6
zf9d92dfb0d588c03739c56254fd72c7251aa6d8e71acc1c6d83eb425bd1c68db4e6bad4e7ae8aa
zc413b85afcdec246cf1f194db1c929e4dea6ef71879d20d6329a7a040b9908a33f940400b737ff
zcc9d61205929cf3e968fb2324520bd351d77153044ceedd63d449dc21656874e07a93a6d1fa920
z044013c3964868f57e7b7f134630024d9c2f8ac9279082e4b9f630fb2ea3160b310928dd162673
z9a3324cb218d785ad1845412e25142e83263fef2a7f46b0e7e64431dad3272bf2a44749d28c7a4
ze8d3a6ac1de2eea67c3b542e596184b855e82a5a7ad9bc792ef56b98b27500d4c1781123b01ebb
z43c45902ea3961a65ed0827b6fef6af6d05730a017ad1c1e0298416b942f8d0658c528ff997d8c
z86c2962c5e9cd6cbb4b3c77d2052a8e2e0a090ce373bc2aa0b32b19ba5636a51c3a05070e78512
z246bccee82e71ca0f94c3ec50bc9c35c0a302ca64a36f62d9aec6df330722090a70f2d0a038dc9
z27f3f1f1414eb74110decfbf7bae8fe64d769db037db764efb1a8a0a087e65026d4d3030d1638e
z843b6931e5c12092fd9d848dad2b4679cabcd479d048f12a69c7836bd01ddc9836cc051e907344
ze27d429b940ce426a76d53fa05fc65911463c3c2e9546c722a5803958075d4604b368bd5b76947
zd4a92e01758aa643bf31a722575b30db9d80e7f0c3389f5b334092b8161fcb0d793aa87ca7298d
z77c5801e7379b1ffe61c4d8e00f14557f19f38e58be0e76565b50a3aa4a9dd858b2daf55e7a943
zd6ad573a5eb98a0ef619f3510abd2202d50f898f6f75a148983ca5e3cdbe15fa9a34e9321c0b18
z1f52daf2dfacae3dcc27057bfb01a8f2be8654e9c9cacf3415a7bd617c78a6a16dc9862aa6f195
zdcb6710c9de8e5498d7c0eaea03e97d229cec82e33375f500b8f8853f59b5d4f09ccc691f6a2c2
zea1fb6655db1d8172d990b51338af7783d667661ff0db7d10a407e535b254e92e6c9c5dae5a4b6
zfb54ee26b1a0e79d7593475e34b350a71382e1bc5be887022330ff1d9b9a6ca6348cdfa9f368d1
z51dcafbaf78dc16164b5dc05c13fcea2dbc128dd4191702462bf66bf7d1bc77376bed183d86d67
zf3b6b52abff856696b0e31aa58cc5be8e30c4d253a91e49ba08a8c5df1f4c3b61eac5fcd29acb6
z82aa798f07ae450baac2bd94a12981785344c6909ffc876ae219c3e43083620cbb084bc30e1254
z17a9fcbb20367a38f61a72e211bc6bc8e7c1151bee9ada48ee3ffc8c583a0b49f25f46c12d55a7
z696540e5a95d1d52c0e0b0f40e5eb907ae46270a639c5f7b6c4e49dcacce24c880724750a3b9c5
z1eb925f19b19684eb7ab2f1bf2d0558cb84a483f01443be3f7ffff3258f866f7ab58bb5faf7689
z1401120b312eabd64a6c74e1d44acd27899620f5bfc3ae240c5b19f41680a5699426637aa6acfc
z848002861c9eadc15f8e02ab24e1526afdd51a35501b7a4ce9e77d19d05432821465daaaa21f47
z269b40fd0ec53c8d0388adff553d7313e0b7c9b07deebdf9c5b851a77c7e99f0c68b8baa849da6
zd014fbcd8c5e1eaf99949404c6764e1aca221721167a35be0c1aa6e80319405c317835b66cb0e3
z6ed1ca979b8a1bdedf371b754fd6ab3c7e4413d3444711f10b1d06133c36732afe6e4d5c7ede76
zbfeda51c05278470f365a23a6887cfa6b4683698bca1ac42d81e5100da7b6f2df35eb83b4e3cf1
z8073c98d5f042242738f11073196fe5affa09c92d860a784032867160aa775f6cf86d51951cff1
z260b8bf16bc6ab5764fad7aa6148ebc35e00df44ba280fb4b83789c33d6d9c07264ec9f09be6e0
zc4f122972ebe7548bcb1adebc808869b6588907eef0e5193b48f8949fb045df7943afe27d3bbb4
z20662d10adaec97b5571f14fc9830330306388a9b334459b0f75b985e8d3ea0d0d6f6b6ebbe96c
zf99446ea2366c29f24bf1676db7d60be7b6dffb2444d889ebe8bc7e3a0c201defb280116a3362f
z9d7a9cf2ceb96e0482eb8719286d5ed7fab7e3504340ad7f1ba4eca538e72ee0b61fe9561b31e0
z0246dde5ba902bedce1e7475f1eec7930990bc9d21ab86be1f0d9339852ca769b0d9f914ae79fe
z22e665a6ee56c85c287dce6a4370ade54e3ff7fec4aadcac84592d7925211751829f593ed869a2
zd7065a36f8ceffd55f1993f3c06585f8905c55d45e6c1298d22b875d31062828fd8ed9bcf4fffc
zfe24310f46f7fab501553b92e84c57201d79c2f9c6f06e7c48d565dad5be7a24843d2cc4552407
z2d08a60a2047aabe2d2e6be6d8f63f6c579f70f6c34c1b5f4665266ae6c8ed58d7b280ca219afd
z5c05372df95e8046a6c7830f350c5f7f8f548b80519c9e1ff44e2220d755a50c552103f0054e04
z4f062b643a99da7c5736f9210a0c259a1dd989f9c3190151446295e73e57320509699179cdb5f8
zee2a8c4d98306fb810d04ba707236d45b60a55faa4ee2d03c1ca1c6751f4044822d3d51fa3a7ec
z926ee4273df1ad34d7cab4c2d93260c4161e643f6cf176329584c3309ae417016f05df1a07ac16
z7e1537934dd12d94a30fe4c3fc08bc987eec4cbb18359caba87d8cae64a290787a08014ab772e4
z5964fc95b9c269dc73d63285de06ec3e2c49478744ff86ba523277596733a28eca222c9d1872a2
ze60a9a66d8862c9b0559323036d6dbf91f4ff9d00198c2f74870230e793eed00b7546141a4f640
z05f295f53f0fde583ce803da622be95b88d6fce3278b5e425f265f986d3f70d24234ae806e050f
zd79dbb2927ad63285f8702c1e7996af85d11c72efe5e3a56ab1d35e116edc23da99485fb2fc333
z01845a7ae076d30fc23c89931ddf6c2886068ba9e57d27a514232582985ff32f6fa1707dd7e56f
za2586e394fc3c3d8639b372e8a27900c08ab138fc7656d15ee7825d1f60c28048751df722f01d4
za1b2c4dcca489b26fdf1aaf1d0eb4733a82b450f68f35dfd0459f7d55ba9840e3b7da33ff4e8ab
z149b436819cf557161ab3b74e555da7496b5f6aaefda20143c4153aee5a73ef6e0cbb2d9327f1b
z75f718d1f690deb8d8c0b715d8a8ec7ed1a02c04bc5c8b8268bbf0582aadd60e84e01efb6ea976
z241920aeb44dd2f9262768c4b980b9faea0e21e9f0be05706e89ab4acbd1b305b027f9c8bf499b
z8e71f54400b423bb85b63ec43fe32d70570fe8cbc46b60c5cbf68c016389774b6d6fee856baa35
zfb2180122e7ae23f6703c1290967276485c06b289c8a8da12036e841ce7fc2b33c6774a8963d1a
ze7d2c729a57129a3670a3145b0b8e1bbb699ad8b7c8c4416376d8281a4ab853e9834b9d789419d
z5d4c25424a41c56619a8161941e19f4b6cc61ae83e7d11005ed1013112086c8764dc607490e76e
zb5ee13c600ed77b88162b6e25fa30dfec64ffbb209e0a0e1f610bd81b86c04e1e5a3333d2982de
z959f6e77e61dba75499b6506153ce7f1a5ad0f115fd608f8743ebe7cad94e1b0f4b5b05f277899
ze91abb11c8d5efe00167a4b2fe047836ec9f2bfded5f3971e00d293462f56ba859a7f09b39bb96
zf80646b37efc48c2ea3e33b627174ba819882cae391ba1f045842755288ecaf09012587dabe532
zc7b054611dc0464283739569d6e41da8fc638f1945509c071926da2e773ee4ccdca761986a40fd
z0f111e63477ac78317c4cfba7101459b1e7632ec3e58085f791bb411e09216dfece4b915650f85
z9759fbea719e8bc325395436372eb1ec3b0b7816a59304a38fb0c1e6827c3a64304d4c851b2ede
z7a3ce0568fa6039a9fb97d608afff568b36a28f1b3e8c916a3379577727f346e924190eb394d97
zd1ee9b1201ff2f1f0f4201b3ec219d700d2b890146421ecc1ee431745d505b4bb73f7927c2a833
z21ebee8b9f9166b4e697552b63b8fbef8a376a31d00f2c0a5231452da0bbf3a7e590d8159a59b3
z97a039aa1c401aa9298a34f3dd8bc5ef9b4741a4b7ae951f717001618e80ce775d31a65874bdf9
z4ed6ef910c3974ed1236663cfe76dc07ad6fd5add3ba36c30b8825bdcc22c3d262e83dc9313198
z19eb56a8d50036fe60e5328827fbe637bf6cce2e37edcf4f70de9a3dc0891e2b32bdd53ecf65da
zec3e28f4586d039bfcb44bc745cf0305f0f37bd54be409c879e50a40bf884e32a36775933cadc6
zf30b61c3be8b68f84b3ce3a3dd64306cd65c6a225b995c03c95cfb56a7152760356d2db750aef5
ze6fa056fbf9020c6e401b30ef983d1f3987eda529df19c659409e68ec9bb85445261ccfeb5ed32
z0bbd17a98e3bc6e17dc1c5dd021cb5cc247144d4adbc04b051ea9263c83ce472423892da97d2e3
z1c21939ea3b984a3d1ed51ef2a719dae372297ab26f45b7acd48a50263314ba3dddc9d38b771ae
z08c3b701e8cd0f89a10122540a0dcb7a490be221458e3278a055ba2bbe144a7fa50d49d1fb7077
z4bf5ee498cb1e83782735acdd2ce622805a70f7ccdd36a3e4acd36122bf72b6a6c3bb46347e880
zff99de175f9277a6ea4b67dd26c2f33fbbbbe9d320668bf67ea883efbb94132f951170aaed6bb6
z33b345d8ec32c371ea41e0644e783e3fd0bd6a14141708baec198874f1ed31767641d2a3810523
z0369eff6a2f7bf0fd4c2f0d15ce85889fad179c05781860311e16debb25259c63f857a9aefa811
z58ce2fd6cabc8b2c93f9557d118cf9881d1e2e8ff95dd7063439eec714d3ede7e1497f2fc58363
z65922b0beff7012df2819f1e493215db3dc56cf40af02b92f6ef0432e974266136e0f65db48443
z79c8eff9ef97419092e838b2a0d4707405f4e791f92909ce4b6e92457b41e0b1ae73070be02348
z1e18ef604914b983567f4fa3b27317e917e2c7f7788320df66bfd6ba21390c2f2688a325316c05
zbce62bd2c1795621b17d73c6355410a79835559b0b1354a960740726c4e5ab75266610a79d85a2
zab3f72ecfe170aeffbd0699e0d14f1a4e5558bba88641fb3a500cea598fc32a40abb59650a1697
z003e1def784700c265b1258c9f80ff4df1528470074a8251d8add5927a36393687e6fef7d69a41
ze0944dc6b9077e7ed182f5c47395a7d065fa8de7f9e1931ce6d6dcf655a47a9a9a049a15063129
z32e5774b6764a2b7a39eb52084b08cb5f88c89dc124db25bdc3d38265a5d7dbc86289c9ff8decc
zd3ef1cbcabf80922f2faa65332a180dc938b66e4d7e8d31733c6a818fd217d2f57aafc3dbc2b1d
z6a0c933d9ad37f004c85f4f8cd3fb29a8aeab7354cb711dd87ba67c970af71920f7c4dc0607d09
z866583bb76997b97da25497a9b00902e2e0b59894f41c114cc3ab6183dcf38d8e9ebf730acfe66
z24bb50203d070dabf670b6abde6e4e56f1dd385512e6b4959975355aada7bd9e12b6e6e72872f7
ze3c2e7a6e9ed6f70ecb3afb72dd5974fb4293be3ef9abdad33d93379a216d5a515b7c972fb22ff
zc0984a03c0df372091ef5099ccdfb62a010bc5370ab6ac6522424b491c32811d2d08191d26eef7
z7f39bffc1c53ff8a4981481511ef0cbf6a075a9759e25b17e72c7a981927f20e160e01cb1fb711
zb6f4d41ec9a7645bdf3b451068587ed992ee2b9380c22c8db169d52d22252757d6b98c7241bfbb
z468d3e47f629cc17105c44d6c20494a0b66ee6f6e0c48c734d36658073ba8a737f08d35091a515
za48f171c782a82b605e00bd4ed45e4bedb62d40f1039c2a1119c19f9a4e53b1d62c2d2e5869899
z931b08c1869b359a203cf4402f32f20546a226ddf8dc5d6b3e31116a806dd0a6367eb3f1d4e8db
z0369c54211ead853a2f97a3081ff95b1e94a9fc82e71c1303d919899d02487dbbcbee83d660678
z66e44819edaa7fc0e191268eef62d244050adaaf50940de0945d492eeb15d87f46119065535797
zd0dee123b920386231a4b0ebcca373f73dc46d4dd60893cf5b57411961cd591b4f04c540945441
z09fd68ee1c6e7618b0d7c11c48d3ee7602bb9142e871b493b42e209ccf735d482b917a24857d2f
zf9828bf89937da3d43f740b1889f9f2966e5da12ddd9b8ca043452995a37dd2c238accc6bc8539
zfa4a2b188b42d48e2198fcefb8dadfae462cd9bb8c47ee3f52bd58b629280eb262dccfd88354f6
zbb5bf115ad275e3a8eab51eb271e61fd09aca62ccc50758ba7b2736943473436d3a5f4d8284f2f
zad4d40d6692d1dc4ff6e59b0f1e9080784de23c22a7f7a030763640f6adfa34f293e8ee3b7fdbd
ze7287d8be901d62d87972f02083feba02dae5155dc4a46d1ab0209879cc01566b8cf9c599eab42
z3c7ff40934559dc4d13641e4af064deaf3fb59e4eed72eb8a0d8bd234c2f37f866c44c608e251b
zb24f5270f376643de3d2c9b58519e1be8967fbe9b54035e82bff1cd3dc519c29e2bcf8105a2803
z004d5421590faefcd14c43302beb86174e891aead5952edfaf47f4750270befedb051b1d8da4f8
z659ee2781708ef5a9aa3fd293d68e394409a26e628b767e17c0941e738b777eb490c63295f2155
zee0d1e6d96316de0c9c3f387b8a3a6d7dc044d33068ee1768b122e8868438fc9081a5e8731307d
z66057c3d7f39155ba4cb12e3067f074011cd70b292cc9891181b09af9384dc224aa54124111135
z4db93fb07d4b5d2a45f2d9f0e03dd305c69c2b3d0823527493d5db37a35e43858444cfdf19b444
ze163ab5f7e4c229155c5430a02c51983fc3f53d217f680fad02fa716f0cd9d055a6401e6d0cb1f
z6b483e8fcace086ff69b94c4f0fcb740d1505caf4d861511c735a66a2720deefa6a4b77056130d
z09603c4cd09f36509bd4fd7960b4463c37b6b29884e6489bf2832b08fb8ff7c4654230c0ed5fa2
z2aad4969cb31f84e345d0b0e292e95b0e75a8294a5ff4c74f937c3a12c0ead085c0b53c3ec23bb
z76f6f697f5fc6230745ebf695ab925b94c209d9873ef0896871a635666651d4b1ed2d9a6fbc369
z8191d633e96331930786af2e8d56bb13f9715854cf7bd9a6e7d24356e28bc1acbd161d3d393bbd
z06d6733172e7aabe3078b40af5651b196d928ce0976d803820d0232aed04a1786851017bde4f44
z55e773bf816a13856046238ba76a303dd6f81b38219ee5ef1367353d529b83cd20392c7a8c5b7d
z8010af02259de4d9463a2cb360b3820897b6ed321d3e5c5234d362673e23d23711e505fbcf55ee
z58bb1d605ab9902a0f887195fbdf6376e6d8a35be40b310411e1cfc867a0499d065c94f69ab7bf
zd38da455adb7438319b811b1142c4e39e6322cf7494264619060770ecf9d4d79531e52f71110c9
zf0a5dfdbf0817fce33bba7b5e78a96fba00dbab58d7cee883145249bd8b82f0856220269defe16
z2cc83bf041c3475436987c84b035c8e9b9e3d9158cf331c31e10caf7e8c5f8d2584031e6e63ee1
zae88de4cc28b1e4a5d41c5c1080c181d04da28d8879cbc80da89fed4345d2181dfc8608a2da7d2
z21645183663020e6bbc17ce7af2a080a35a7e61dbfe4d0c31dd4b69af116fde1e89a25efbcded8
z2687e01a6629d48a53a66c265984a9297f5d90382c3a9b2f3fb07854eb9f467c813ad104cb6e99
z123dd1d7666b078d75de010bb99189235a0a0b4845931a3bb512997920916b6104926b19410e7a
z52b44a81e8b77df03110feee48ee828a7763651bf06523faa77ba2acad9090262d880273c116ee
zfc94e25b3afcfdefb41c3d5d16a231720f8e653a23c368771a2b261dd337fdf864633c336b33ae
z281cb6d6ded589a2e06370412ae675b180f8eb58460645fbfaec7cdfed0483ecf443d6df41fe1a
z99672a6303238f8e35a7cc7e6e16a06c2a22b616d7ea9c26bbb4056f04a905ea1939960a92446d
zeb1bdd562978cef2580cbdbc715a48842c64c122a1f84e2d141517b185faed3d77056117c5e7d0
zb9bc7f85a22c3a15c8f94d09d46626ffc1a31fb4782d96dfc0a27c375b3a7f35162582ed1fd042
zacc70971ce064788062ca463c2fc2e2f3964a90b1f3ffe221ccc1578ff917ab295fc61bf0f8e98
z492938e38ec3f50045ab3243ec8277afb99132a876161472a5b2fca3166af09a1a6271bcfcad6a
z2dbe8f900896745032d4a2f713a053eb9f89b40380a29b0418b2686cda13636ff86880c6e0f303
z3cd9e7d65c9a6492013009ee7a40b7c7eb3f417f55f9cb3f647345a202e20b3b52b4642007dd8c
z28756cbea6f3e01fc0d652f801592607f448f25c71ee462aad6445590ce41e6c31b172bf4d4889
zf0f442bcd64b7430109f89b7bd548fd0775d72d124e0aea432bc1cd8be46f6be4416ac5a63be12
z6e5c68ed716924ee3cdf289c9af371f6009eb8b3d6e4eb765c76fac91ab6b01669e698608e39b0
za0b0c18773ec5f20329e7aabea9644e19b0eada305b8a17e981959c74d74eb249c9a8f89d9b5a0
zca6b90104b3c65e5d1be8cb7c35667fa8b13b1f76d3a19c9e44a5df5dba4191562552101140d17
z282a74d4592634a37bd37ec1e269bad72c48fa2cb8f77bd7a1883537e92999686f1d35bf2909a0
z352ccc7143ef24656ce9e407b2ae57b2fbd5d4082b215cf821174df2cd73aa73814a507b66be2a
z59cb49516658f2a3478725ddf7010cdf5910728900e8649c91d9cf1e0c9f4080fa6b7dc92f31a4
z491c542c8cb5de9d7ca277b681ae757af200c57afd2e8bb41839fb892677b708fbd0e1b9f8d37e
zdf7daafbba12e06b22b41ede6d67e87cf6e566e1cfc6ccdb09506dbcf3d205cb8a7f903bf81d8e
z48e22324e3e69412cdd67fd3880000ff604b01f3e3846753d6bbfad88193c973a607d876cd1b4c
z4a7f3c3698c39c0f41a50281b603e71e8c764e044161cdba8debcd7c5042d2981d02dfc8325627
z684a76997bf10b45b1a6f151798a35565047d0d967df23ad4a88952ddf33e5a9675444eead5cd2
z7d54c4e28538ad565ff9bdbee128ba8c202f2bb17ebce46c4d69ad1b690738758b47e8c446c635
z43108962525adcc5415ec0f638fa20ff61c8caf958df2993360b1c7d6a2a702cffde4bfda23541
zf0e218a3f9bd9a0c6b900a3fc28dd121568119509ae60ba281eb162a557e8eadacee9a610e3ebb
z4e6cebd3e1a84adf16f5c4b8e9a5c439d15334e75690063dda3ccaefb241d94f19bed568fc30f2
z419c8cdd6653f3b79f2e91fa879064ce459d3a19c2d328e419c94503c0bc13c06cd867d02bdee1
za3c211ff41015417f5de541d407013fc0e7d9b24f43476142807a62a5bbd04f7742fa482ef3e66
z8e3bcc596adac812605bf8f14450151e27409d73e054ff81f674165a4bd238746390539a624bc2
z2c7a9719f4b8678ef3b9547ad72db8d92b19e51eac5aa904ef05a43ac7b1c44f4ed06691799ce2
z7565fea6dfb480b9c109cb1a056ca58e0ba6612e8953823027cff159c93a4401f82b9536367ed6
zf6d7ee5ff8208c7775bf2454fc3372b5da84da986dc5266930440dfc9768e109a9298f3cb5d8d2
zdb867db2c63a94f5068f6f88b101db96576990e5e5028b977ffe997de7048bf20860926676a0ee
z557a044c806cc88cd919829304cd9c0650bd9d027aea645add009a180692d791603bc84c88cd89
z4aa64918268630f0bbe0fff27f622866f6e8191de22341fd39accacc542e35b5d1f4cffd0bef8c
zd7083c0ca742cf22385807a78f4ba0eab305f15c539388a6556836ad1ad97c43c3fbc24d79b32e
z4a2bbeee5e1c94abb23cf5f88c9600652483b9cc9ea4d387691b43559927b305ffc80e8f2a6136
zfa6ab61ee2b014aea013e3498cae18d3da170a83502a9c7ec5bca0a946ae0efd237ee39e7b6e4f
z5b7bc5777adff0237cb70958caf40267a592223bfdf45944a77f089e181d6d791b3d94883c5b9e
z28c2ac67bba10401aaa0a3407f1e7b600ab0670ecafd96b39197bc17d30ff3f0350ac09378e680
z2a645a0d6ff9b39e890aae517277571e443f24f39b9a88aaf8aae8a0acfa84e77fea4423422d43
z5b645cd0543a76dcf60430230b7e33eefc5c777db6748441ea2252dfa0db27307ab40b66414055
z3b3089b5bfc2b6d022e68cf23d6e2904040c3a9f7a2c0c33c7244ea451cac6581fc5c82f6f10e2
zd9c084cf44ae4d0d037aafff7d83197dc544bba76d5adacb8fe4f0bf9f0cdc9dcd771df6b06adb
zea57a7d46d5df6f8f730553e8e4ee867d7b9e49fe9df617447b566fc3e27cc5af2e1cffb4428dd
z1c6e87d1a87835991a2ae5b7289ea9b807a074c22966b1e8fe669939bf5f19e4ab2c73bd6b18f4
z7acef066101cc8c9c72619a1e5ba21ca0275093ce8322232e9cfd54c42803c7a31a7534d026386
za48bff2c16b806ce80441a386eab81518ce1452a88a26182809ea49361065df3d3f9e8ccf7e4a5
z858d54f627d8a1585827b9fb13b07c68309d2a3f4451375ca41ee7a8a7e8f2cdf7b25d41bc603b
z6656a7189a28af99d9e154ee721343e52ed0d1e9bbfdb517f47c85666b13748a4316f64370acbf
z08fa5d5c73f24478fd79c4b9e0343bd00366606d05ee55f26522c5d7800d57622369b23783526b
zacce4c2e8fde3dd8f6f1eaa9b6773b61620bcf9750e1d57fd4824d7f4aa296407aefc21690a41d
za216667cba1c5759719988fd553abac0e9c437236d940a5e0ed942f2b090cd3a1ea052cf3bea2f
z3efd0de84914ce961f1243c632ed2df167aa059af3c16cd3eb29cb672bace6ade3c3cc6f700098
z66612645d3119054a9777673d26dbe0af510b0e465b85c60a7ea126d8366352f20b6eefd784294
z4e62905116577563ac3c57c22cf0a1f10500747a47e9da42f1f190a767e413e44e951333842bf5
zf117e664d8058ffef59db0f475af1ff60118f91acfdc993878c85255a457f5d53f20989f0fd2b4
z0dca00619a5c09a48a9adb58786c02eb588a954a3433b168653973a6e7d125a9ba1c51b9df0e4e
z92f47fed79f6ee97b080bf75849e95498f16c91b9cad541367ea658b6fa7d39fbdb9e1e0d63046
z0a0e5f4465f14f61fdc181ef5281fc5c01e4088a1676d87f0742344fa8e55b1d8a0cc1c97b385d
z85a39793c0cd020c199b4f9173d2d7057c710241c45f01bf029402bab6b816385b81b3d5fda902
z8ad9dcfec1b8f929825748d3f146ab4e07bfe7519c3f565a1bf3035a548684ae17f9079cef3598
zfaf3fa29b5fee5135f436955b0315334ab2692b27634fc43f4d2811a63d0b004b2882d68787310
z2e817fe8d692a4eb507881ee5bce432f8e9d396d872a8d56442222d163cf70e462574bec9ec034
z646ef33530c7e688f6fb729c1a2726a750e39461467a9961fba73cc72061c095fef3791f676c64
ze2e0c48801c84484b26ce77168f59222f3eb3fabd54a33888faef2a03f1bcc2324e770e18a0f59
z7a1d5973574aaa4d3859092995f0d48d2885adf7f5d946885cd8e1db82a865ee9845f287f2a274
za94d62ebfdf5098c5c29f2327fc704ff1926469c695955961b99fc651433df6f19f0ea0115a0a8
z36a791feb6a8fae7da818de602ef9af35940f6cb5c1634abdb11580cea2d91a0fd1f998e6cd74c
z20d7ac67b11c59ba0eb0c56841f77ba9341d60f744abd0dace19f25ca33b0220e78656122e951e
z656b6417ba448e3ac28e4c53e639ab4e20fc45f60ce050835b412d73c02fe25f9d2707f975c1f8
z6441ec82cd9db42b1a905fe722f5f5bc2cd22ea4d7e747c00544303800256ae91e50eef2eaa0fe
z69c2898ae664ed6f8e65857e8f91c1a5b203c9fe9e08ba3d6737b0293579094b28d71b9e65aa30
z0c96dc69bb855e62bd1fc68002b831d252573c5367ad3fddee4a496b4e042ce038698bdd130e86
zb1e3953e637be953787c4d7a4a065a4feef0ff507a181cd1720a543a24eb834cc357abfd727680
za2dc711335a51cd9b329d54c53c4747882872cf1363a04552b01464b84a648c2e3890570718c33
z46065a39d385d15b18537e95af2c6dc51edec6046feb396c2d4aa52505647aad1559dfb10a9ef5
z19cf97a33831a5c6631e53d857116d89536c3681d39c90bbf99e6d92db3a696fe935c184f1f872
z784a1ed3868ba5a174be47cf27c842e8fec8b51550a9f1967bb06669e6663c190f92c5d60ff0a6
z17028ccc22a28250ee528f689ec5c93d65ee84721d4cfc84309bc1fca1a6e19e1d22791247410d
z4569a159e56a3287c28da8f4ddd868d89a1750bdc29e4bd8c59c76f43e98a275db9b467cae3530
zca9aef74252b4a4d2afce1d9dabc0b59b7f314f76c04cec2b000e2961c3ac7d8d657d3980adefc
z383962fe52799ac034442b150530a7009ce3c3eadfff9131437f979a3670f768bff3911eace7ce
z11c3586ffd476fe2be7d4587c393df200076abd424f94338315d027c3109b5f93742863a9931af
z51554feb0e3e01f9c1fd8ebb4990ae6b826eeacc780f8fcedeb18d3ee74d70e30e62c87b59c4fc
z8ca7087b7f5d692c958ec1f07685700a9314c0ca2bf8cff951b7836acd5190b9d24429e4dbe1d7
zbf6ada30252b64516f4bc59711ad460161d3640e113fcde0d7368029178e8f88a9d9334c2f0dcb
z23314422323722d145cf4db1311125af40e4953e43f7a8e4fc58515461b77dc5eb93eab5f6d12e
zc55167503b0cc090a8f69b1b2195efd53d8d2926c75ade9f30d341935a43d09c2f3d41ab722fca
z45ba9c9e09c7fd2946a673c0f373c46af40cd453859c1e0118d5ca960071738fb8b653b59ccf37
zc7b3765b793041246c4bc1f3d2f8271ab953208513b31b2ae171fd6feb77a659946acced7d8a5d
z35067870165535d4782b916d07d18b68de2e269fde4c99dda82abb1668d3956425c866a21c4bcf
z8c7fa2e101e79b966d5aff27df0361ec3845ae2da7744d0ba907fee66e71331b19ba932773c443
zccf314d57f89a62f65665200f12c942df839bb6e1d54e8282384a4575a537db6824503f82e76e9
z3277cc5d7727fb489223596f28c4c0181821f970789457cbd6858ef75f8576f56c8b8524a82379
z047bbe66b84d4cc5f24e7ace50b007f99127aedd7881c3563948f2b0399822dee3f3aecf8be0b1
zf09511031cff6822a382c43a79615485b84dd79733e1581ed0e48e4475ae0a19e6b4bbd32a0294
z20b0304f92fbfab1d3d04fe0a6c7820ad59e373319a429b7b290b5227521dc58c04ebf9d532676
zdb1229580c7578a968e15b576511e36ca98e59549771d9a4ace7474767d4081310d87b769fb926
z364b1e7994ef5ec6715b4a0b2ac0783e9d1a42b9977b15bad8dd29c49d63c69428945810f1b5a9
z0a13b2de5709bb55f496855e033b5bdb82b02ae3f74808136624d75638b2d66988ed2e7a60fbd9
z5193458a076ee622cf240aa88d7ae0ec5bee9758bf4b659865e9c16b7abd13deb3adf0ad82b029
z85c0f35d9bb040f95e3399e91c88513a9a4d69aedcd4a8f9fde497bd00754dad06bc36c39d29ef
z53e7c7a42fa3517dd10823b7c2bdc82b53c4353a852bacba42adf7380a21f390df47f3d28ddc21
zbad85b3969efbe07d30a4324ad2c162c6ca377d6b69f25f46cfed604de32432496d91afeaaaad8
zc6331d4a0c0cc8cd854f9a99c6b9347e05389eeb5b346221047ceb0c14a65616c15846472b9a0a
z45f4661d1ccc989b93d9ed4b8f9ea2d7a0573ae44dc28f43a4c92761436826a5c08d5ef8ad386d
zc0ed8f42336a50ea685b3652195bbb88149b59b61c0e5b99da509ca15797bb0df54d1d593cf189
z7020ba168831807392a95df4287f923d69296b12589bbbb475129251b31b8151d56d2f4001d80e
z6780e54363f696197b018b6df3dc8d9cdb2abb850691618af76b2a0226bd03160dd3f81435a2ba
zbc9e49a9da38b4892f54818ac56a6b246e73d44264f97df986fde339a7d00d03cbc8b802dcf603
zf7099df982555f505531f68e85fa85f2773ade6e00a1bf0e8f7ec74027ce60be07431111da22fc
z63c4e18499975d276cffe41bf0ad697129175dcc2943d37cd0a9ee1707b6ccf42f0ff008b3bdcc
zbcb2e629d7574008b1510247e973f4377308eb256e4f75cab11b73b2f1ed58c22230c6a6638cc7
z9a04b9460c1746528607973da59424f9e0ee463e6f1d2bf410986bef0e93a103d08bea23444aa5
zd0553cac086ce39acd69b0d2ccca6429dc23ee4cf16eb8936d929c57d74ba097eac7b51594a0b0
zd25572fec1eb4ae96ba929bfbe95bdcc2dff5577e6f401569b6a67a82eeaa24c612326036dab8a
zb4b24061786081d201c9ebdf983f5e2aaa840c445dcc6cc43a790e3608313973006a2ed0356e7d
z5d9575947c572e1c88a3194101f44cf7cc23dd27156fdf341e0424b0538351623c3e8c0efa571b
z72b33ce68c16ab9273ab79b3d93bf1aaec671bc6d1fba2519ecdc676002ecc59a700e23f021df6
z962c81fa3fcbe2df0c37b783dc3b84319e70bedcc23951ea2dfb87125a658d969d779f207a72ed
z456c00435692edcd6d29c8d2c8f28fccef344de8c22d198ba727036354fa488b39c4dcd7d90495
zdc249e74bc770076d1b9f4630727ebdc85cd3e00a9907be1be92bcdcafc1209da26af1274d5853
z1a6450414903f47357f00133bccdb69f5005148d9ffdc788a0ad96a02bf2086fbf24c6c4591311
zdc1191d23e34b4b5847dd0982f4993ce603549c8cf78b334735f0ae9c478bfe3ee6d2c3ae231f9
z11b9b27088a243089c273d46f6088e692cb18f6f3a25119b9c7f1703dc109b4b82641d0f099331
z9d70b9862cc65badf3c466b5741291f24a66d08ef2f6c6fb9c18d4be73b5c1453a777bc8c7ce67
z109f20200da4f595169445cbc5a44c8215170a1f4e8347f35cb1990487a2f37a377ee0ad7b220c
z5ace6c9d4470bf7aad3507fa06b7c4fe6d33395cb99554b94f8035601ac73f7a7b3ec0522b5c4a
z16e0ad21bf2e855ca2cf335fa35a05c4bbac925540909d6bfd92e6ca4bc0d068e461baef9f8c19
zb08978104e5cfe7ed9efabdd8c27af2deb6566d88d5f8a7533ba639cfa758c4a2070efda659b0a
z9412b71df3ce3de05fda2b0eef0ae52d712890927793422d397b0d04a26d5d70f01ae162a7730f
za71230d2d465fdf28db4ea20e0941ff69ff2ddf15cacbe67dbaaac44de6e0c99cc6208a8576b97
z6041d006dc3855801903127d4ea4287550578dbc1327afe5a3b6f62f1b90f48fa591fb859be64f
z390685d15996720bd396e6c725c336eb3a69dd27517ca624403c764031783c92ce91d844c250a3
z207a7e4e9c5e025631004fe59083277428460619d2ca78a0befa6fe02a888cc7b271358f633ee6
zaabbc34f09bcc703b8971f14a9e0afdbed4625eeb0dab664f90fb83d45eb68b759c3cc743ba8b0
z84909ac3c2bdb28641ea10d4435c2565c93acd1682a7f988d7ff2108dbc3056434235ad3173fc3
z99fbf83414e937b1b4b2cda1e3ed8862f4b18e5d95be117d993de3893a440bdfabcb2d161325f2
zae305831640f91d1bf92cc5bdc6b9e38273ed8ba746272c30de278503fa0a056c738c858843449
zf62137a13eabe770538a3eafbbc5daf1482a4acb8035654eef071927b9535cc6e6ff2281dd8b97
z0de9e40b5dd3c176c13e0b1c6934a4cce064ed99a9fc0bd6409580b6785578f269ceb1a1cac59e
z5a37718fd8f074ddfe8b37e2901426c540a74ddaaf1d2e774adfd7e84679de4f316a2a91cbc49d
zdf990cd8aa26181ef47c37fc00cf559235563153a3c28ee1bbbcbe85410737967499a3528db9ff
zeba49cf263e313ef8c9239e3b07917f8eaed5562f0f95bf60a5d88c2cccbf9c6b0b636ae491b56
zc19dc8b5da1f6650abeb7602472e58a480473fe81ef2df13d8265caa3716535b897fde018a539c
zc77a9279a9c03615f29916bd703728c93096250b889cf5636f9d76484cbbdb7d1b97fce763ff03
zb0e2e9b883474de488cb38813faa516463790d95c96e1014d19370277a04f4aaf2e99233485065
z549537b93ea88528a589a844d2e7fb6a495a3d85411d16b74d7e2797ec10a03375a22e88e583a8
zb0055480c07db47a38ea23ed32b941caad3d9084778531d71614e21ffb5709e57d16b89778d002
z337b4135d21ef8a6061934caabb6e0d7b5ee6f6802032571c863799c59c8642d62a5d47e8fcbbc
zbb19906ba4c2e4923010016c740c00c22e77e1b1362351ebc049c5f0b73863c9fb6fcb68f66f39
z712ae6cb73e3e5dfb5ad4ca1dacd4f3fe57f10863dc2ca6a45038856c65a8e3470989d1a7d6dae
ze211c831d39f71059dd36f1ac11e3829d1abcd91f38197e79740fa15d8994bce70d20c34981d18
z51a44838a224822d3ef150f33e196c78c38445651610cb9f3043a0ac89357a0421f0ea0d0a86fa
z5d8a10454a37131a09bec8c6062af05c81cf990f860d0c8ac14b6652cfbcc321cee67c6eacf763
z907914096c60095f15cc34816bff6444acbd466c91c129397b8875376deebb94727001c009d601
ze49040bc72a5398527e1acaab9b112a8d3af4830a6ea0c3a0010137728a59628de2478c91e4289
z482a1249fa56eda45e38e48a16f669165fc3a543fc8e151f3cfc0cf8c4435961359aa24fb1ce70
z8133a53927edad6b57e035502ec5049f7fe5ffcdde786bf1464d67b09b1899f4daf4836f42b38e
z6c5e0f40d40edf1f9324469d74e0042c6f6683bfb50c334c0790141dc480b1b8dd5e0f1f3be6e4
z191bdf3f9ef080413bbc1f3eaaafb8d604c89853ba456059611e7b9429f37394f98cc8833edae4
z526792cdef87561d24415a24fa546d971a08cd8970f012393c8df54ad4c4ec2fec93a4e554a5b4
zcba373213259815e423cae1a3cfc3d1d61ee9ddc8163eb4c78d306c46cabddf6d6bf008a6c4d64
z859989c66bad918cc701200d1f9ac54a699a3c63c8082515c701cb48cb525fd75b125857cba0f5
zb0daa23c406b9ee80ce3950bfd48c7fb2a74e3e061f57e3234d76efa535776deba227942f906dc
zb707ae61102e82144f9073c0f30aeec6f88f40526af3a16388242f9ab68b9d5155c5d2eff27eb8
z0645949bc56d99d8baea7a4029151d763c4456f65fbcb63969581be22efbb3dc02b2b328f3a410
z841fd94382f3ead19c1932497651114a2639e0df8b2f17bf36164b0d8f0e8d540515a6cce87f60
zae8f854d0372d04ca051a03c6a4d1e00b19337ad215dd83be32b7410cc921bb788d9285e0582c6
z566909d5d6fd9177d117915a28597494d96308ef30d8884b67c5f79b57f97b76b5bf59ba7eb777
z7632ec32a35a861c761383480d9475bd601f6b538169729d68fc0cad765de496c9bf02a3213359
zbbaeb9f982ea5c54e704ba2490395af92e0d8b71f81699cad052b600ac91721e17cbe6a282c515
zf93ee429cd31bb0ce5ae15ae7abc72007af78e29899196f38a2df71346fd951769fad8a0f1c481
z5921165ddf8bbc9dd55b775f5aed3ad5a6942e04ad41ca8ff7d6ba80d9e7bb4a704683704c8fc7
zf7ec9ef1d849c576bcdb770937f87c13d2eb3310f1604cec61eae3b4a0309e5f4a83a1d4eb9f09
z5853b45bc3adce556f7f5947c050685260225919b4922482ee05d4474fc48077619d86010fc106
z08c2034a9aa69fc34764ead519e2ab18aea0fadbd79892b7241ae720fafe7d9b240d96b809dae4
za405fb0fbd678d8c820131f040be3a2d907ca6576ab3ba8edcb46047e0419f45d4d2175f875717
z929b946618a302b0d8df72128ac32172c938913a27aeff90a463050576b450a4bcc54969e26d6b
ze381146795271a41419d8ad63cea194d71616bc95f5cf1b20da9fd2c01f6fdc384ff2b0f757ba5
z2bc38b97a39ee7ea36ce210c88d3dd6998040c6f9c6c2be3e59e9ba947a57fa19f33e55500046a
z919dbdd058332b9f9fc89f8fa415374e3b868a99d3a303096faf962550c31630f149bed78ea83f
za9f333e663118683795bca172c58b837380f3be0be993ca6b98a112fae8de2fe441107a35255c1
zd036a701de8f4171e9c6a1ce01e1a9699670093867675ead3dc4b07681071df3e45c084c2f67b5
z02b1bf1ee6e2c523e61d0e7a820c122215d0aef99fac4247634b3344e6deaa69db1322b2df0c1a
zbf01b2003d881a3d3eb1cdd5c86279932a0137b4e48a57aee9f0a23c2d4e1b3f0b537205bf196d
zc372df01e17c820dcc69b8efd0a33c3cc64c82dacad61a776343804a6aeeb05e1275e8ee214a7a
z810de9f84632c5ea38d60144dc4d0c65518365a704d4298e9c2d767c7a527bf510370bb72b1635
zdd1c6f9b6cdc73dfd7c3ee9324d595927033bf1c28f9281cb7e7bd3059d785c64244fd80cb8f13
z50fceaa7e9916ea50b1a39c7b0a909052a9c5d3e7cc5268972f68e2a95f153e27277407b977dd2
za527452a885b43ede0a66201fc07facf2d123074f923af4f8c4d17a983df0bed7dbabeae9636b3
z61aa78a589296af33807bbd87d2f958191ac146d8165f6277d42dc39875bea326363cb116a6a2e
za2252ca1321847339f029cbb109c3a46f89d876d755dc8ed0c20c40a6f2ba59a3843490889baf5
z0006d480475d9ab4372672733381a9c995579a79a32b07849785c2245f3b1e35e90223130a18f3
z1a8fa97a579cd53ae116e0e5a0eafb9e2323bc41ce72cde495d7620d4b59198b6166ffc49dc8bc
z245c89b2e8b1c317fb8ef7d20694a5a6b68cd74f55947b95eef356eb1f6937bb60054d66730389
z6fd44234e0e49346a0598482a3f717af5652f153fb304741cf01e2c55a5b58a2a89ad9369e153d
zed5417c501f979932406555e816ff9cafb23fa40d02c84ecdde2b1b0dc0a66e4daf2451b6dc43a
ze97c53e50a71de16c06b735e6440aa59769464769ee306b543dc16ce1f0319ff0d4676ad39f090
z480f7716df0da9a44a976dd33b3b54ec4f65bb324a1781a218d24439188d2d428f51bcae718f1a
zc4662cb891774303c7aa705fab6a7443d2f97ea33a6d3ff4d809734bee84223ed19c0acf12fa37
z362ab9a12526b9ce51c46b732f169b62390d33467b1244a118e739e40d90d7c2f7d8d863bdf86d
ze48604d517a4879146a41781b42bde5897ed5a810d5ab18ff85379b0a24bfa4ae851fdc182021e
z83ddd5a7211d6e81ba3e31e7983069beeb98aadbedc0552d464f17c0882812475d41d1c1411f84
zed36a3e718b2736b41bcd09f5ce11e877d98ebc8d1b74d8503192008d07ac8a148b016c4b47135
ze36c597bdc3dd8acd4d03e73f94211a3ff9c7f8cb04f25e717131db0a676451ecfd5da926c42fe
z383b84c4035fabb9e709206b5855b3daaf4b47b9bc47b994ebf1f1ef36406f83bdd0a27338ba08
zfe9af3fafdd699fee8a1675b9edeaf1baf94d8ec288435a5339dc7892fa5a0d81a9b14a027bef5
z4a52c41803a10857a87353d4861b251acbb6e006dec178a48c9868f907b6c7469575f789f41a21
z2d120eb78d929255186ed0026a9677efbbb7199ac2abda7a630139c11ae435378291707aafd969
z09d197f9d18290855a7a9a31bfa3a9ee1dd387fa69d230ca98e673446d168fc9e9c89ad0f9b19a
z1b4b2a564a4b6ac98dc7337274395645d2b8d78d140065a199325df80bf79cd4b3dcc9467f1efe
zbc7719b651e9f825d3590a481c1275b87899d6c74e71c17601c49aebe1e2b2fdb14ef7cbc4aef3
z4305308f256abf71c8d29dd77f5dbd19ecef99918b69f0d34c83dfc6fcc0aaffef8f871f100e95
za00267b53435c8bced6c6e109db4526b5e29d7ec6d32c02e4d2147697aa420fc655e0f4a470d9c
z2de9c9359695f12a9887dcd2e3c270a16e9617720b22ec0a8751f91f198d82a31be8f7c2e9c63b
zdf90ad6fe58e3ab6460a9edd4c668744ba4c7aeabde37a39b564c40350bf5e9c0da724e1c5841e
z4b230c216d9718b3621e256d9bced7eadcfd42c6836ec71d83527500343a672aa4d3116fffee86
za0bc925dc9fa3bd98db8aa97e757d5b927a2c10bdb82cfb4eeb2d5d7bd21b39f29650ab9878db9
zd3ee6e1ace87ca979453a89310ee6af76048ca37eef2c78ec91b41bb86613c93101f7eed130d06
ze4caea4aacb5b205a393cd6def597ca2c98e7adec1e5f7a5c0ba84c5fb718f7ff296a907dd736d
ze5e0a1804fcfba59e82abdb75689b400c3c0bc307ed1a4e6de86f60e97ddf4bba47e9692d7c98d
za4bd2a3b8be2c572bdb92432f05bce35e460a441cfc34aa216fb03d249d8ea6aab2253c61f05c1
zc2d1f31e206b81127067483962e0a259678cb720a71b9a3e464339dcd286c982f33bdea91cf239
z5f7d6c443bc8e4e103d4a5fbe3c8eb97d1b71f7e6a65fb111a4a107ef6df1f4f463705aad23af1
z92f6214f75b902c28860a2b87a9d0a5313503ccab77e2391b664427c1ba56159149d3d46d82dac
zebf1ef5f0f7e229817764021437aebd5cfbd218169a3f8e0c0e88c6d28732e3ef278e3068fae01
z3166c1338f5b9b4619c7eb25af5c762291577fab9ee5f0a75b6f9efa230546c93fd8e0b377dc47
zd8f981a2e5603d1d8744737700dfc0e65d9e5182cd8823a5d045652c21a6fed589ede92586ea20
z73aa149d43ee3df8866d430904bf613eb7372821cd2b59667bfc44cfd545c5094d84e576b3ebb7
zc6b439d560625c0bf63a911d1054cf776d6ed05ecae64219fdd810d75b2ec1b9e1eea7f3ee80fd
z7debba9a716daab2c29017264d2cc61be1b2baccc7e9cbfde4623addc8785ebd5dd47025764f5a
z83711b6cc26909d3d164fec968cb373aa207fea318a6726e8420e58e4260a7fc18894807e0ea2b
zf10615519bb31a11867088e26da2b400a2305d9603e9f0877086da924327cabc2dd65c417cd79a
zf509a56731476777523208aad88566e6108b33a47ce268c7b86d4b1193d99a1d05e9cd6a7e1c68
zb8e236ecb80703f2ff7ca88107ddf9ceba7121b4235a4bb36769cdecad14739c29581c7393ca6a
zd528d0a8ee44bddde9fc50ed30379e419b6d4d5af3ff1e2a440600fffe7b2fcdb447ed530a6a3f
zdd8e3a89a38bbe6b2743295069443767fd8c8c9072685601ca0e922cde8b169261d2095a281584
z869a1adf5ef77ad212a16637ce347a46217f1385b29136c625376cdc6b61a553a965e7688da81a
z03eed5a0e032aad78e2ebbab39f6d12e0df3090c2b492c276554aa07a9ccb5899950846ee9b41a
z784739bd4fd19527d47183c57c646cce8d3a1769f7c8a3b699faa24905c17d771abd645db9b840
zc16639e8c1e679fd54d3edb0d0107a2ee902853897405e48345dc535e2207a47629bfb42bc3685
zd068fb83f073120288a123f3470474c3260f72c7d9cce7aa7917438574822b8eac78eacc7ffffb
ze1a9bc598891a0e2d9370065f1a0903b30b55b1adc9d7e582798614dff05240ee0a3390be2b8d0
z34ff9ca2dc0a801f47eeb2216b61caff6c636f48b24f2089c4f37aa507480deb8f6183cde6d5dd
z5a81be2dcb675b8d2f80dd37b19537ab64453e2608ea3a6be2ccd37e63adc69a4ebfed0741e05a
z7de212581f294c5ce3bb5be466c9fa0c8b24fe278fe80a3eafbea33c16b6b7acf3ddbe210d5b27
z883b35c8603ebaec9a168d8932683a502fb9a5bf973c6232c84c34fec10e95d22195fbeb67dae1
z429bcb780c78538a8f06f3ac209ddb1846329f4d350e14948b81d7849e7d0424fee9bc345da7f3
za70ecf949861ddc73a0b5502f9e6b0d1770112bb5a12f62fbebb521bf3dc7a5fa45f7ddff20be8
z4f425b4a3b92767173fcaa1cf664d83d3e6a72ba063ecd331f923ac3a6e04bb1b27f3e43817875
ze37308b9de7e3de880dd20ddb488d6fc9331fcfcca6837f05aa00ce7ef12a1b049de69d45751cd
zc6dc280c6b7250a5e6cdb8d9eb5dc4fbddbc4ab635c3164a47432c899d7d081f22f187681fa2f7
zdfc5658b12d53ee8cff36e2e3c09b8a9f1baf5d6f16789db03055af14cde039552dad0b0335fdb
ze14ab7c84acc64a76539ecca1d6c42e1ef8ce9f9daf274a4dc9adbf5051b92fd0d536c6bdb9c02
z55bfbade62b75fed9ec2cf3bb6027bacb6f0ceadb7e4e0f0a373fb2e001a71926a290702cb3e95
z9da670709ba439a2dfa2863f8a0864d57554c2c6bc9ce90d05c5462c01e40b01b97bf674fbecea
z5047d0158e21385d60aad922cf50480af86fb9dbe1c67872d93d7c189c372f8b40386b5b4f332b
z69f9e79bec7622aca10958e7ebf7365d3beefb0c7d89b650c2beb4ffd331f1c073c7221a9a7cd7
za67fd6d3242b0a594233a689131bef61886f2f90801e4f933e4d227ebd9d9989dc4960c5e89244
z0c9f4731ff59d7213640bd081ef639f0acbac5dc81b91405efb7bed503811f9fe7e74d7df84dc5
z625b3640de2701754eb99e1500388dd5c19b91ef65ad7ea72fe78684a00b0c19b0dd91dc2323ac
z585ae263e96b085d60db8410df3f306a05db626c936b88da3b8e43242785aa64a40c1b058b8c0b
z3d119481a6748e88e3e6dd205ccf35dd1884331c7148728ef9d74c91552b8d881a1c733050fa8a
zb2010e3acf149c0f9493ce2750da220d99c73f114dabe5735130754e0b2f9af3eadcd2240d7771
ze813a7ad4b05cdc55a0a138efc1df25c6f585119b8dd797f20b91eba64e6701fa60ca4605b0b51
z4fe65752f75c90e31f4a270d135b07b4fd4c08c8d9992f11676fd19dd79d2ee7d8dba05505436d
z26830ab84da9c0f908c1341cdd8663e2fbeeffc8a8edd1a27d4be0d2b4ac22191716b4a01d96a7
ze0af47352d56d8ea6f5771d9e3fe642253cd98e83513761a50be06bd5543f52d1904f83d0ea9e1
z00ea6950ea17b07fb3b2fdaacb6692f77d4d934f769e50ff3a1946063ab7e1a0bb195e3a0fdf83
zf77fbfc964a0427795a4147b0bebdde90d38b20041e1b40576fc1c1dc470bce226e238d5841272
z1b474f42cc64f286ce2a7afba3ecd64565ecc71f4ea84548f845820562db286b3722f1f36a42b4
z1d8c3a324f4d4e84d36ccd774e2e2b2ca675b125e9527e2279652abb882be200f51df6712b87e0
z6d6f7e5429d01ec1d76aa1a4932f6f90ebb1ffe17941e1a4e937866bbb3d4aeb335a17e02f0e68
zf82a7b78e26a72d58d541677a4a9d6b8fbddf2819f0c877455e242c9336c74f7119d8c6458f9c2
z029b5e4a466da1a1c0511492af090d406df0dd13c0c37c2c1617665d82ca57ead299574534fa80
zaa25844cbde3d85f47d92e50f71f2d184a9ed0b13ab414e38ebbb95d4f2c26abea672d433f0e05
z8062e396566cd78e3c50a686902b7ac38894c227bc40c22b4b210289089d8bee255eea7d794f91
z22786044decb793390a5e00fe7782b403f314fe8195b48a0bb83eece0b698265ce61bfdf574b2c
zf0d367698f4f0ca8a71a3d7a5a22f4c180d22182cbc860b567f1b18ccc136e65ea797d5d7f4c8a
ze7800975944356b5169bd6643572407ab113f8f16ee15a7feae87d97a5f75d5ec2f64715f32c88
z7deed315ff48150ffdca804b0002e1f62b8ea11a7262e188b52bf4874aa36c32dc87cf0db71855
zb2f5071932c018cd646b05fb4ff47ab28a6c2ffc8d0ea46e641fa6809cbc25807081c4deac9609
zdf02919af0a6777cfdd35c92b98757be1a4cb178046be4ea47c3930eb7830c1fc8830680f465ff
zb447701ced36110ad92a2b53856be28604699182e71a2dad3bcd475f193b51f4d7c02385347cfc
zc39e2df99bafeec0b159381e4d2e5d6ff411f50d95ca90ac2de81b37de2c62c651c0487c7fecf8
zc51974dc29b342a8491b963cb91f24916b69f4ccd328f975878990d9f5e43903e91d1f16f34785
z8ca46ecf0a362366ae9e6644b5fe2a6d98231e10dfa116f0c98bc5d7460782d93627a0e7a87c79
z912667003c6279f60cb82c625c500bb72dccdf2e05b9c0216dbc466277842dfdec550927d11f24
z9af30e677900273d0e242efe5cea686926cfe2d360c153fb168225326ce629a3cde7bf87e15782
z702190f990a99997eb3706da44cb0cbca812bbf2301f9b7fe20c22af56a75913c3c0b76e991647
za7b8f7206ad527572a6b1a4912495ee6976d0c6288620e3db934d43426df81b8a268a383034703
z66403e23929512ef0e34277625adf4a18bb47cf0f299af61cd5c410ecfe1f4227925f50080afcc
zb299af3e22fde7d6250937a5f8d8346eed2922c1477f26ffef03558e33cc1941419aa5b837d61e
zbe51b022008503096ea353b701076098e1ae0eb782d3aac52fcf8028601cf8fb667b8459b1ace1
z8bb2eee4995e13bae41e95bf9ee5758d536178e8c6e2da5b07128806c7d8540d515e615a3fde1b
zc7f6ff4cfc0743cca5defe9ee4dfde83089166a8b69ce0d96a20aedd3bae551b98d83be9e4a189
z37ff4a547ce4096cf77863da14f83397e8cd826961312e4e2953333aa2f35d6c885e067bb9511c
z746c0f7b688fc1ce70267b6963d0c0571f33672f1209cd0eb65c2e17d315b23bb27a7c627b7a3e
z4484433c0d9586562f2f218da63adbf77eb6521616b2fdcd10d02747ce7d79127b92bbe6855fa5
z5b624d9172588b67f5a0e5ee1bc0f1d3116410b6f6fc6c86d72a7d355cb787e7bbb37e2ae1388b
z1edfc3a872f9ddddbcb42852273a08650acf992db0409f43240cec8d03553b56a56f1f2193be96
zf6034473489bf8aaea7b885ed93a3c40f18c9ce3e53e346fc44dece73c249e7b5b3d9ff3ea5cd1
z0361ad387e55cbbc9e01bc0218c469e25e2c3242fa75d19b0343c1496309e245a59097c570c757
z3789771cc29876f577b068a68b72826f097541a623a6964175d584ef8b78cf8b177a9a6417b819
z087b96cd07bb4d3d5fafb55b025ec20fd1d8afe29d4f67ec6b38e42fee24a3cb8770b2811a3796
z0c63f934de5bc929d020528422fd0791aa727e2037afbd3e44fd6da5dbaa2a4b1e6a233d350aac
z55547bad409390baa9f3f56549073d692bbff95d471a7c2507d9636f8f8298f1418573295e75c3
z271f55761e1ffc14fa02512e16f4e40fea6e5abda17cdfa35a415efd8162368be8fcee2db8b2a5
z9ef74e24a281601fa1bfe9fc0f62a99a29b2c01f052b159389c55a4498259670cb8056be6a5e41
zcfeacc511c06f44098ac65f9c61b0fdff58fe0d26e1ba986eb925ebf3fee5cca37e1217e0748fb
z4677ac31fea15eeebbdfe18e7cb395400e60bc2d49581c095755fc17cd1aa6b9684d3da9abd830
zba9ce97937cd7bb92427fe768c95b0240755a2f371447078ead6383e2db45024b861e9f6dff07c
z0bdb1c78e7eff66f05ac4b80d6ef47884b575d1718db5ce23efe1a8bf66fcd2b6017dbd47e5cd8
z6239d5c0ec98f1920903cf38fa9455765abe67c884314f5cde30af32a3447b3922d5a8bb895457
zb0fc76b555001c6a007db106d7a0ab9d2bffc0d639c60d24a7940a8c6c805a48ae6a794ccf534e
z1c7487cf7bb8e227ff92e71ca48ac2af88ccfb90fa5c35b6cc2ec673ece4f07748dafec79d1556
z35f40d216a98317c1f4c8988c3a73e62b7b51ba10f78bcf086d9a1a7c581fa728b6c36e2f78bb1
z19525acca340dc6acc7e44bf752689dac8d6b620096531d938b396e0f4f1f1652ffcd992f46688
z7347606abe286cfce4d54e035c0af7b6b01a11f362dc28653d0f541a8e119413ce5028c8c2244f
z21d68a3a9539d27a9e7d4fd72b35b9288441c6d87e3033c504208aff2fd3eb684946f150133513
z70b04459da3874f31412c31c9d49e6fd87ea42ab1b952d1fc70bd0001b7d786bc28e3400e43ab6
z88e3f85b3c8187f8a1b8d6aa3bdca125110f0e72734a160fd170a2f4660431af296b8c1972f197
zee3382ea3fa4e75de5bdfaa418e5fc6816997001740e75258a230703b8f76b2680dacee3c91e24
z2ece1d07ef5061429d4008d1622031dc0409c4712fcd908f788ba9267041dbf2f017a34c677704
zb75ad94ed5242b37d844c764e343d0866fb34f9da87244ac6ec26bf02c0caadf1bc9314d36cf77
ze0411eaeebe0bc84819e207d9514c8953f621a68e2bc67a6ad7eadf7bc1a47ad3c7f6ec8bf6883
z80105187017d411735640e3bbdbd3ec95ed174029269b9030557c8779fe5bdb19a232977107ae8
zf6b342574bd1f0e95d7f293a04f3bd63edd421ff0ac86003bbb42f8001dcd48c4992c287db8ecb
z0324f87165d43ad49ac7c5e2c56af76cc3a8d25771acdc5a68a4373d78d7a738cbd0d2771c556e
z9df09de379fc522ab0194a7274ecbd2a6332b212ce8947690eb67b6adf9e0e47c3b77dfe399ba2
z73300288ce53cabe1e4012400c430027a327a09b6764c1cb9d6e4bee32831b4f5f30570dd7cc48
z8613d79d3df5b265c977fcef17fd46b6b7874acde2f40eb2b7aca30cd17ed649e3f3ef1a347f1c
z157591f29e3d7d89dedb76931a99f764123406c0566b212672c1ad95e791c9cd44d995c7cc3f87
zbef59c62fe024ebed945b2f4805fceb4b40a000367ae321657efc3ee81564ffc10c7a0536868c8
zb27ce25f33264137669bb306cb7ffdc16fc1983684ab56a7d7c4278bf765658c8b1458c70251a1
zf4de4ae627cbc3f23d4b271afa621f4c42a4198707365c43bddf4c9e7ffbc174aeff5b1b0cddcc
zd430066c6eeba025084e4a6e4c950c0cd8e7841ee53b94a90ced4103a0ad6209938b5f8a9b4800
z10562dbe5d88d3e66ffb4f8b4ca1b729e1bf8245454edde60cddc146fad5a6cf82805ccd58d866
zb230aab5a89270675c765a9efe59c2ff8a77be76c598cb391631ebf5e5a1546e98776ee3fc9ff0
zdded4d075ea19437b2348a756e875b6eebac2fe7c9830ab38b662341801a7cb920dd68d3bef647
z7e55941a365ba0a1d62a06a4d9111a1aece774e29280838b207a9cc1389ab673d5dfb2f5896cdd
z56073170a6a0239952568749652e16687389c61d65d59ff38ff99acad9ba163ff5142c0499575e
z1eef013cde7cd50b3022acdc862d4950dc4c82942833fb8f2ef9bfdaa2e709e5d02ae8453049e6
z088b9810180d13412ab792cc2a330e1b151ada106a22a6c7fb84ed2deaebaeae0a957468a0802b
ze22292325979f321a876af7db1081cdeb7f29f23d531d1f4540b413fa5f9e03d6d66901ea02258
zd35eaf8be43311323224761c52e43b167509aa723cdf763bf52bc58bee709d9f5796286422be37
z173da4207582a49d8570cf5015bbae1857047a251a983183f47d650b9f9fc8e9aaaf1e4cfaa541
z3072e385cdb08cc6885eec36db84ea14be5fe8c2b192cb398b6ad8220e4ff4d0d712a3bdf89fb4
z2f08acd474a29b6fb46b58990d718b4d9e96006756858a0946877fdb6aa0f2c0e49e362fb73dc0
zfe6b41107b248763e9d483fea965a2da6e40af96b6b6f9c45bf000573abe8fad8254ab527c36dd
z4d421ddead488215f62bc939e9e985a36cac2a990c5d371e01036fd7e85393f80cf74c4b2d3a19
zd874c025e7ce70c42e8ac74caf1d241c73f03fc6010285d1b1f562a22f0706a9b067fff53a6c0e
z2728affcd872768ff67cf33a037929c841898ca34647cbfcaeb31511beba2355eafd76cfa478d0
z0c314926aa7c488da939e344986e1e9ebdf152d3866a3a042fd124d7195259315d9ac2310b6f98
zec01417e913fdf3b50c9bf9db3895d310809aac18860dbda0a285b78d09b1552f03fc4cd749f9e
z2a38cd928a4a9208bd0c6f555c4408c31251f81f07e768b9293e7dde26423bef1d699a6dfab90f
zf1df45368d7d111053aa0ef0ed8c383cc95863a3934d3dc67cdb63417667975b9ce114ba31547a
zf72faf16178fe465a11797fb24f5a33ad0cef6ebd57aa7373c74c5f8fb096f655761983974c0bc
z1b9ef0b018e0a0f764530b4d808982a90079f8ea82237c86488c8a184b52271ccd73a2520945cd
z2a787f3c47fb730043f4421cb33ed1bb8da15f88c06c3d11bcc5f183bb35bed309f2fc0abfc78e
zc8a8232dfc47e6c0ed36c81641ba917f98aa8dabe6ef90f45f783526d71b13b1e5927ac06d1ae6
z73e2e1e96078715de3aed0c52ab6346548363f702c84be590f557209920c7d8be771b96afe652b
zda799caeb8bf34a991c5729ee01cd3f36fd2bed2b8080e6e6e3f62d9f2ce403423522255f06a4c
z61a1ce6d26d1c7b46b2a320a07c98ba130cdf6639c4d3c518bbd3ee4762ee4db8e621a484d4d48
z3464211bf79c8e0357b0baa3e7465ebd07a55c47445587e9906436e0001dd44e5105edef8f88b7
zc290edefb55f7a79e4b88bbb5f2744d88d3a9acbb83e5e8239140822e29daa9850920b28aadec4
z83df59467e7a0ffeb622bce1ec2dc8db0e97f8357ff6c3589adfafcfd80313ffbe88f29f3948e4
zdbf7860acc30b891f54c129afddf98cae9496a953dbd954984b778d90b212b0491bb4336a9a270
z936da71ad9dc29ebe7ad2ec76462bd03c7b165dc7b22a2375a7b18ca92d78e88cd6c5f842f4679
zb07a2cc415e4a8383594661387587847da56ba6d2a94a3d13c3332e5cc9d69c0a796d2aa0cd79b
z18b7519c53b81b183d5910c3c7b29bb3dab6f9f8f3e3006dd73e9f18575881bb5bcf1e20ce2be1
z50fb12d9a88bdceec28d04e99ebe888f072441f1ef2e2905fa8f3f43c638bee802b1e5197bdaae
z8b8d6e86fd5be0591dbcffd7e91b3c2448c9ce2b8b9fc5fd7398a750c90f17c8c17ead18721ca1
z30c1abcbf2fbedb4fd48f97b4ff34b87aa018776d98f447b52b157f5e34a517bd7323136539220
za3a3e6f1ccc7f3359db18b12d3f76ed3d28ab494f5ef97e48bb4958a08eb89d4352fd04b2dcebb
zf46c324effd4d7f9e5c3601b6841bfa2f1dcb80b947ebfc428a4f2bd49d444396c6952fcae76e9
z51c16377bd68cf1fb26e5e90b7949f9dd5f2b88031da3c1d4c9504d9417065d9f333d3e84e17aa
z54a44ec333da46147ccc05893d556ad414dacc02048e649d1d937b4485bfcaa90de8e89a1e8315
z55d88f9dd39fe54dea8a29e08949531289b2c6d5296354ccdebc6d8badb2cf6250e3d647ecbfc4
zba1eda0e8445d25205ef6e9b3948a416ddfd51ba9e0101e83ae9f4cdde602c0991b21f6386f92e
z6c0a4d50ae820b1bd30aa6f035cbf58654edcaa9000c0d3f41495c220aa40951aaa8e9ffd0da89
zf8a99dc73cdede813c07facafb97075ed55e2b99b32b7a9c5b43d7deb25ec249459712e065385f
za623889449c010e30167abc80bf975a090102139bc8781de7547b80fcb0a0a60f215a8a3e9cac9
zf72cc2d45cedfefdca2d44a9a007f4708e521c184544dd935eb507a707b9a2ab03d2a53c345a84
zecfd18658a58bcc1d156c454ded434094cb5255657a6a5f19dbf8cacf95d79c95897459b32864c
za8e5ac6126d2549f7be6117f2433e469488fca8b3a90d25c37173ad04625e37ce25120789e0db6
z33153f922c42e3a2c8ad0abc1b6497adf55fa4715e00db4c9664bb1cd00dc40a7804770394ebd0
zb69f3d9e0241a28cdb64364c99089e563c1e46ca0e2c7e6992b2f5c866a187d4d51632950996d5
zd1eefc91bcad140bc61ea9dad2f3944ea98918f108a1f32626840a9999e0ddc9fc2c7d80f514da
z59d4c95681d2a41980b188f6cefd9ccfe0e48e174098344127a0985c96c082921c9f1b07faad7d
z54980943bfd15494bd5af3e235d3aabf6264b8687ff39f528b7217b8435147f8b2b14fe25ad22e
zcc0120bbe481d29461891dc70d6ae8afa338a56d4195bfd96710d8ab80b60985ae67b5129a3295
zf27d9e9b7a1e50f4e1b80ef5ce2db41756113737297f462bb4c9a1e4856956b82b8170437d2a3b
z55dde800261160463efe8072083bf78077f1e2fb3c3ad4ef7def42b8a72868d48a050609ec37bb
za916332e6f4c2a55ae07d427d407db2bb42ad4579b2c72c19465bb07783b668e6963f3af8b3184
zce3483376c5383054dbbc19890c53ccfb8dbe4f6b186fecec272d129786c01d40d78ea76674ff1
z5146bfc4816e993efc6576858a06338d5f4f513df60b07a3f92cebe7d8f5b220adc191f0492691
ze2a12f55d8eeb2597597e3f3d36f13474c21d08673182d03e030eba14a4fd87f8a852d26d94888
z8ffb9f6856fc75a29debf9889e2a943ac7a2566f880100a75155b4476619d4d8f0899bd94dfa36
zef28d3e08d730cfc2a965d80f13d2b0db919754b0b6f90b682238ba7f85b42199bb9cac3d96e0a
z17e91c77b51c04923957c418a1378d8b1d15538a7cb8ac4b97b27cb87300c206fe88f531f8edcd
z0033fd837d85ce26550c0a52caa09381b11e2e6b8d72b114788d0ff53e8ff5b43ae3112c8748bd
z18ce32d41bb68e28fad1f9bec7c71b4ddef6b56c5dd61a82706c72e382249aba46fd5a077fa9ed
z58a89ff05a25c964f17df9deb39ced5c6b59834e264e588318a399c9553983c8cbfe901f93b35f
zace4c92d8fbfe7681fe150791e0a118a6cc36c3e9205a8e8b11679a66290c24a7c3c3e2c196dda
z4e42cb8fc46f6e9ddabc91caee8c3f8539ecd256bcb425ec3423a0769da73bb14e13845da83098
z8428ae4552740762f294e45956e670076f0ffff7b0529194f1d5f856eae8b3ba1e25de6a200935
zab89643a355b7b2c6f67ac1249f23e813f031f7fea1da2ae75ce147726738acb35d1926d98b930
zc7f51212c82ed64764e2e4d55dff139c0361ce45c8dd2d0c35df6d029c67d9d35a548664206523
zec851ff899638a5f6ff9a0c1857724af01d3d8ebe54f6dfd0a80c4d54249d5b5fcc540f57fb7e3
z307b33db9dc85101dc26cf5b8d19707fa76e968d2e72d5970689af6aa4b3fcb6c8b423ee900839
zaece6a856b311c345f784536dc8c12ee2239a1d01eee0658337002bf0f00030805e38ad11b6350
z4cc5062c6904c697137d220402e94cecfa3549ea5a00271367f915c1a8e0ca699cac059f202ead
z8da0de8179c30295647bd65d61f9ccbd681923b4b860f36292e534cbdb69a6d10f65b3ed0330a7
zbfe02446933ac654a57452b77921414a89362e808e3956794158dae101adfedb4cdc779abae56c
z7ccb029d149e696f5231142c19cc3ef6c51fba18adb4e3483e32b3638dd480bb833ac11523208e
za2c10bbd3ce2880cab2d4367777644513cb9a375c5a60f779df9c2be222290925943e869a7c6b4
z1c92da77f1f9718903b9ed5cb6cc22eb4498482b90ae574e0d071b6c00d661f9f86877f191bf07
zd7594fe21c8b19bba95d414dd8115462730a7e39973dc9223ecf9019485084670be73f378502df
z1b3ba0614a7e4dad94e5ef71fbad3315727f1b2c31407081d6374fc64890ab45c8c15e717f97fc
zc25cde2ba4f9687b0158a885bdc5b2784b54d6f944b3ad42a2f27c883cd3b1082f053e2a0b3bbf
zdeda349a94d28834479f5385c7f37657cbb40a4de533435f17fa471606d9f7369b94d6f546668e
z6f4025e36374724f42f7ab1d01c6af39ce440f8d80323ebc4e672d4b55ca21b6b77f9d18748156
zacffba7acf432330c2d94abc95449ebd1c352bd8afa48334418e7c503d05924dccb7afcfce0835
z62523597cf50065da76d432dcf46df6eecc8fb0fca6d0c9d8d7ba4a4945ea779b67e93543e0011
z3df1384d74237dec6f1c9d0edc93aab9a03941aa5f0fbb503c0beadb57f62425283ed17d46c70f
z25151819a59d95ed770031a9f9a2758e559b61e518db71c4c137f8033fbc0200fb3b0f56524992
z0cf10e4fde3d4134c510fb1eed51dc89a464e35e68a4c246edf82822561466d5289e24acb64123
zc4392d176e6ca464538154c99e0bf5cb71e47782946c3a02372e516f3a7f61e9117824b5915eed
z6259bb8840bca14eb9f92f9dc710b1eebadfaa1660e0e0f8aec1c091b3d4b4afdaab3143635887
za026ad5cc580d9276779b8fc052c4c43ce591254fa054fc3ef75a5d233f04dab375d72d26872e3
z100e390e5b02905509d389cb7d9f804f086e369c7f69d7a51e3126f2f29d02b850114142052209
z8522a64a7ef3f23a767cd2c5c680d3846dad9dea98112492c926a2e467d6cca1a38ff9663237d0
z82f721b1ea66c8b4adc5a2ff9ef223a97266c6c88eb71712d44b6378dc9f81fe98e4b187ca8e20
z09c05b7da85c4362795dea18a41e954dd76fa39db67bae7d315c8d4b530c2b2379f3fa636dc7fb
zfe825f428de8d1af351ce76d0f6ac73321aecd741043c121d25b20f000d54aa9664e712e845aad
z60859eca4f2809e9269572327cf47f6eec4e2da7167e67a55a597f46ac43ba343a7f5f9e1fe81b
zf486b34d8823bcd7b3bb66400e5d1434148b6024c2d92c8417c363b115deba01ead4ac756722e1
z057ecadc7bfcf094b971a3fc5db923fe6a636df1271f235bf59280029b5741b47b07d11fae3d19
zbb693e78073cb5590dca6fdf3bb02ee3686976e9db43cd330d441fe92871a8a3ddfbb8fa5a435f
z26439f8fc015a23c6dbdaf3d7e1a4ca86e9a8108c5c831034f808176d4aa40809efc5116c9c63f
z5f42a8d143d92ccdd902483ace42b3b57b1d2b314c25ba37e505e6a773d813546a8bbd59c63ff9
z25c00c4243ab5022ff5492fd04eb3e377c31a12e06763997abc680498faf5d2b3a315e632c5f8c
z7b243ccadd8607ff721ee0e8af8c8920debf632d37f76dc37dd5f38e0afb9e6830248cb521ebea
z987267631ffb3a47b3766d8f1635e8309e0f657264c8f278845c46f7da69fb930a26f72bb97426
z9fea7b891bdd0672d06afc5d58ed0aa6bb0746523e7970b7d187eaf919b10f13d7cd8a50e7e0cb
z995fcc98b17e541ef6a554477c79f7a2691da826b36ae37efbc0977b818cde74957c7ceed798a1
ze99c6cbbb8cd8e1d3a347b1ef5ccb62566945d5f470c77a5dfaca8d1a1836d18e354a863356334
z6ff104f395e58f8f41eda7dbad69bd75db43ae1c8a63620419997bc3960bee662cfbc6c54cfb35
z84468dfebe0b6f691e8af16fab8c01a4402e34efeaadc4d36e719445a57907a991d4c5aafb385a
z2c287cba096147b58584f1b5393332e9d3a47b387aaef03660e4966d8b0c00bce19203fb7fec4a
z4c809e2c29961763fcf338908959b6f4d8f8c03108c67136a64ceaacfc60c1150a2b7c4a715475
z2a9ac82893039a204f4a67ec2dac37c1f45413ea82765b248197ffe222c998607c922d630187b1
z6423961bdefcce94190b480e963efab97ec63ab0c2c0ba50b405401962fd9ab377d451ce91e888
z5b643a28776361ff075bcbf0f747d1b1581fba57b7933dd59251a2c0e1d4065cf73c0887272bc5
zb7bcf6f327042faa4e968db1b811216b65678f116fc2aaccc0e4fc45dbc99578b1a04d613b4cf7
z77a26e139e2a5b1ea2213c1bd95680f2a65e09f492489b45775a410579353a8dbfadc8d27d6782
zc9ab174a2a7245778cd88cc7903a8d3c5cc7309c6fa104fea7d6b2923383413404932df58739a5
z72cc073f130bb3bd05fd02ae2132fcbf7e1dadde9e474462781cfe2b9b465ac671c9876f0c05eb
zf09c19222eac1e7b689b2464f8e92ef12a052a72e95c2a9923c5cf626ab21e8eaf6c81d9c406d2
z6cf81d090dcac8f9972e1c25fe65eaa2c03e47a0bc77a6fffc102719219538e3c86304cb48cafd
zc9f194bad1b9a785ba118c319fdf60abc044d6e4bf9609cb343cc48e0813b489974ff8a388f27a
z6f16ec8c56396d2092c63121301956ee4a8a8c5ff5ad00b2cb1f7e9bf5a0484068c51835cceaae
z27eb3c9df1ee2358aaf446415b49cbba22854c976a539f46b22558e653551b7184bd3049e566c4
ze8ce9d2d36ab2124177ee7b1b9714c6206e5e9a54232dffe04bfcd317f8554a0ca7107902d8b0f
zb22f849196518cc2085d4838ab8714a8b4a1940a178e4eedde7dba53b9086d90b80d01ac4c266b
z478cdce18e63b3b23c90d65fde1ce281926d7ad4700bef094a3327f73571b0b24d1bffeab207cf
zd1a651ed7bdedfbc3b60f7e3328cfaf610f5ac86d03964f70b3381479b9a1cf9afc78b00adf201
z9ee2025c77453caf3b50e758e2b144aba1e3f102f098272c118579b4380dd07b863b717df91363
zdd23394d93fd531bb42057e0a4ef6d13c8165b6cdd17daffd4648e72e14da3354ddecb954ba53e
zf776dc24122a56372ab26c44fafeeaf9cb9b3defcee1c2f0f4dbdf57acfec955c8f6630a6cb231
za62566e9e8dc080bdc7cba32a6eab541a7b9c9ec8e5146c20c8a00771cc3f4b9298cdd4b23cea3
z30435a1c5406064f60dc1c88b40eeea9c22c916a383a2fffd8da8a0b8d509a6c4c3588221f75d5
z5c85bf44405b83d36bb9f94fd98e54dc48d3799257cbfc87d88fa88664a0c095d3d8da053cf1e9
z432801de471dd4d5674af108711316a6c1e4fade661bffddf032777aa1955b954a8bf94a5b5975
z87218c54feda3ef31383b0634bf4c53b8f6cb9afbea08d4682dcd7b2cf463a379134f4a146a7c4
zf59c2a1bf804a66b1c25aa5eae401dca8741b984a64ed482386b74e802ee27d1b2605abbd31f5a
zab91fd52dcf6e1d67a1d69a4aae4e1d25aa79161bf467ba0dba900377d1251f0b782170cdad91a
z0a410469af020ab27175ae0ec516e289738be0d3ebc73c105f85421227ec549c8bbbe295b769b5
za455ef8529d694cedf40bc21dad15e19c85383a28195c19f4bff3d28c503aeb20413f4e4b56728
z9f504e984a0e24d7e630e4e201a10ae28763ae8b55f22e7e1363bb5363d41437e6c9d9e6ee6cab
zee49c86bba54f0bb2266990345e6f1f2d01a0d17648bb3509415075fd61bb9d98123cc2db0c290
zcc48fb2e1f25213f7b3c1f90e21a8f16bb7fa0d78cdae14542662e397f65a58b3bf72ab87e828d
zff76df6451c24a0558b6d0a6943eca240ecfb0d25290bf10320efa83602be06134a42ddeeb6314
z5bc924d54a6c7075336ab5a2fe22e7714adcfddd14b360b2f7c8864c1b53119a0b22de1898dc48
z27ae509c7b4e04ac53a5df4d82702b3ea2d1eee00c36284db47b8874e848d0b9e304fe6885a360
z90fa32bb7fc8d28422db31c0eabf79849edb405ddb55cb1ac5aed49f7cd281edaa735078b25e72
z433a213f1d1a28592ea8797f13a75414d0e504d9774199ebb67cc9c696353a211700efc8b56694
z5f1e0ef02bd29be1bea06bd7fabf31b21227d9ce0254051c96e0c545c12971cebeb2ad679ae6a1
zab1182bff902d25568874756673a8bb63b863343e005261833d51b60ae45fc88cb8ef6d7ef690c
zb6e616f6bd36b98153cc64225bbac517889975036033727b24dd385ced33cc5b1251437c607760
z92b528e021a5dc226feab9009979973b6b5f316fb0c553394075b0727714767d56ae7a3eb0dd32
z32ca4ff09cae715660b8ad81b7b75260929d952ce80d92b672db8dbf23f11009f6e64bd4ebc548
z0a4a86c4592d66b0c60a2046aea4b0657782624384f8145e7e8de6baa1c892e973e0357a814910
z0e26d8a4de1dddc946ddb1280a7b5135e08c0ba2f5f34eceed11a54bc1c871085a96f0c940055c
z52b1fe89894ece7acea9e5e8f8a4148db86e579f5adc990224bebecad9247e66d5583874dc1ffd
zb7465dd3af6efb1f1e227d330551c1a58c9eb29bd5e8de2d2b9630fab265a2cdfbb92c5eafb932
zeb17cb730a4a6b5cb5bdfc6e3caa002551fe93443004130786048516d52f2ea91c7d8f998ad67d
z85ff122c8fdf649cf4c3915097d29c19a6da8f3bed579505af1e209a8b434eb145695fca899885
z41e72424d49747e3d28fd18330e976a68cdd632af596c3e9a1b5aa59d803f014b242c1c774e02e
z5774b82d604f1874fa94179cccde0abb3cbcdefdb4a1acfeb184d68c3dec4f8068401ebf59b23a
z3d173f89bfac57a676913ee623dc3da881eac16539bfd64aa297b0230922c8f5e170dab6975af4
zced57d9b7e6caededf6756658aad68c4447de39d24115d03738ac8fe54a076a27451506cf4ad77
z4289735503e6d59ffe581839cd8716fbfc5902863caea6a469013575d1997e995e8e9cf6847b4e
zb9a566b2aca7dea547132ca05ea1abcd6b1a89a370c17289a7acf24374d295083b4a14683d2dc4
z895d72c556c988f9f18fb2786dbab722cbfab3bc130c0eee550e4723abc539adee9b98389d5261
z10e33a7d5a041eb240d5f6ebcc429ea4a1b69c304989479a5f5e2eeadcf8607fa541435a973e54
z9f5ff1551aa6cddd733c84f26ceebcfe596e5b3e88ae64351589cf290f55967a511df67916f3c5
z76c7d28f7fed1b7bc6a6445c606b0edd3ccf6d5dd13d758b02c9d00f21aa358f1593dae68a883b
z09c163d86aa9cf3d04aa318f724d6b2a82eb9bd81d98ca15aafece0dad22623900ced9140905eb
z00da3d9d3c189b21a0466a384dd08179ed2d4a522fef2c5a73c32732c194b31641ea66c3417b55
z9ce7a8efa5110a7d515b6b4b0a6b64b41a0667b31957e484dc53ec486ebbc62d00250f2b5f009c
z9de0c85f712ed19349a6d2b13e885a547c29b73952183331d04ddb4db9f9231e6fa245c649da83
zf0dfbc1c07e6bb066aef999688011cde391a7ec1baac7a10847945a110937f347c06baeb26b0ba
ze358389d9e4c6511c7031a58d4e3ab842fd15ddde95475764dafb80425756dbf77ee8fa7e12749
z784792aa47bac60906e3b719dfb54f5f6c9ab88c5aec36b794c006e2a1b83c121649a541f45b9e
zd375c5dee67ef9be75b5ff7ae86de1c2348ec323f2cc2784fc5f63de9bb659ea9ec5937afc3df8
z11433c9050ca5581196b49922d941479b8d3bdf8284920e42adfcd5e1060b1fe9713ddf200bd4e
z1add7f0a1db891dabf9229d0d94ee22060bd7898fc980d2bf74da01137452f939f9659618d4719
zdbd2bbf9826f61a165da2456f8d005219c3906471a18d09c4d40b303d06d4292dc8f22daaa8026
z606aa56ae01e3437533abdf80bb7d3b6d5afab5a1a4f4a8faf5065a7dd47c97eb5281687d7f9a0
z335ea6ac5daa9eb683c8ce94d2c2d50db99b86a7ced25b9595cd067930bdeef015c67d892a00cb
z29797dac41c8a6b4e9f3d659fe0168f0c38ce019623e1948b2a853d50fd367ed3fd8cd6694fdcc
z402a8bfb0f3bfe51c71e291f6109bb679c1f0afa56f07bba587109012a8add2f64aea45a69a228
zed62fa1b4311a5e752cc98b30a4b9ace09dd665934b8b6ec430a277a35f8e58c9eaea0ada0bbb9
zc22af38bf51b291b4946708682e1e11cc4dbec2b34ac1bfe8864f489ee7dd2c2a030dbcd9ce0e7
z1191b79260bb106798dfc0583367cc2c6e20c82bdf69e717df95dec7698eceb8ce701d3dfd7046
z5d2c38f67f435e51b0de57781a110c6e07171647d9dd8c0a396db278cf5374cf59cd92b4b5caa1
z2e4643e28344046743d87bfe14d43ec77b0f18d2204190997348682bc3ec952ba8c1246ba8e41c
z9851bc160172a0b73f51e18456d3b639837e16d41bd7411d21cb01377093f5f13e6cad1fd69d37
zab533cc601117f8bd39f2d04e9fabb1a5dac29223d4918dabb713a658fdca8cb5dbd60b7d73ca2
z98047285f8d0fba63ca11809da4658e37e3e1ba61430aee43bd6c9c140f73faeefd1f2fec19d87
zbc25f060b3f924e78d02c0fab53c364ac60865603627ed2f7f82483741f45b29af43273133e375
z9e81aca55addd1638edcd5d17eb558cf3eaa4d3ccdbc095dcc00f7b66f230efb47b5dfb8296352
za7a24c710313394928de0e39fe270b22e6e6cb63c404a9e14b78bf0966fcc0830421c9820f002c
z83b332460300589b64b4669a1eb8ef99662fab01a231b8a2edd6b21f5b5cadbc51b63e14336fad
z968572fb843c852ddf695579eaf834584ac1a3386ee328eb1348725cba21b5e0da253df5574dba
ze80d5f2737fa9204f6698dd8cb390ebc21efab3e9d636bdce8078f41273863992572368cdf96ef
z7be7ed860a8591b23cdae2122925b96542dce6fabc91f0879be9a7f98a9d2273d8431984488100
zc3a85a5641501962bf2903ad7c7bfc9f6ec0b7f1dbd1e545acd2c80591d9f90023e3e0004cc5ae
z901b1af5e28f46852729d81bcb4a171aeb3078c8b27af27b31dbd0136f227467a6c993c9f986b7
z8c2bc5e8a05e421e81eeeb40135e83db4f32d3a357fcb0b0f6b8edb2af5daca74905e57c061b51
z9f690a524f2bc8a11a523274a95b42b3b850ec8e26253a3a9bd1ce3aaf599ccc35606553c57823
z64f7b2c58265fe0262290bd97e4a27cf7393e86df7956825003c0a2a7da88ab561dc920776e65e
z88db53bc525da861a3382d3cfb758dced685d141ef2f9d15c75c2f230871cd7aac00b38d86ac07
z9032ee2fba9e525caa5ffda74641bde872103fe234aecfa661b3f76589a7af980cb3a58bdcb55e
z9e205d06fba104f9711eb11bb8d5dd6f9826dc1b1129f6f3c6c581ecffb35dee896e73e27f0683
z654976e4c6b7b92b2e0992109b7db1bdc7086014f77a32fd0428b047bec78b0e81e92117f53d99
z7607e8aa86370de182e3a632061f19d393ccd4467e2ec26bcf55783046b2eb3f495442285d34ae
ze364312871159f17edef43ccc28e3b7a972700f290e1ded1673dd3e7c76dbf33bf840a300fb509
zfc10a7770417edd25617783f69840971aa17ea0957c174c59e5bcd76fa42edff5c1dbfbfc9355b
z91a7e726bbc7f243c952e3289b7383d3060254af06cd8244a4da9e6df7460244ebce4e3fa681d2
z5728b6a7480de1b494f7b28a0db378202b6b3ba98185417c0bc279cd602b45d4c54394a41f428f
z282a37e99c587bb03b487e0548d4fbde45d1fab101fa2fbc5e1d3eab28ad0395cdf2e96006c524
z31f7bdf1b9cbab9e7657ef187a5ffde2856b4edf4c84f6f893d713917c65fd5326b35843a98f76
zfb3e42f6c62c15f19662af2949c204b4e58dd85f6cf10e8a64109bc9362eebb16b0109b6bd6d1d
z50cc59c3cfd48f3d8a99b634f85970ec3bf3b39e99cdaea7c74ed733151778d8d21e0cd1f0708a
z5082f688fc6cd579871642e273e1b3eb8775e8fb435f4ecbb0c67e40d58e85d25455cc7cffc7a5
z2395ec6766e2f62673102c29d7cebb84da3b1b72fe666b5bedfb36c694b0cc05856beb22899426
za521b6e4ad3367a7d2daaa93ff62a8de14565652f06ac791e7cb0b93040e70223dd4dd47991f6c
zad372a190dee78209266ec2e2b2291439109ec991e1c1fc63eb38c6d0f7c73b462ef48be3ef34d
z85c3b78ec4a690e0331cf35eab82a3191262ba1e11260d3cc6a5c29ba40e8b3464acd35216a98e
z97a43b10a032e0c544a38d93201757776d1b8745894fcdb72d5174093e48b3dbc5db9830ad14c7
zef3da59556cf384c86a67ec5b560d0f85ba7d92135e2470a5e19a517b0e70c5db9f465ed31c607
z6f451cb94304ed5d3a60a84fa42923f101030ae7b097ea692ff5bd2a1cae96505f5b5d00615cd4
z4919ce4ec1e423de91beb5089e5263df63498728924b744152c79948db9f7c6cf3e492d3d8af8f
zc143cbbe7ce60703b10f72fa85d9833c569ccef4bf6a976b40eabb9706b3f282a2348bae26d0e8
z64e82ee606c38cd93140e2ffa992c8ba052b9c3b9b632f247bf7855aa3d47899211b7e21dcbd2c
z1f90bf4f51e59f0df36efbfb2ed5a12aefd89b2be2562d15eab9935406803c1636b60db1dda93d
zfb89c522ec37ab763155d1cdaf076e65fecb0e0147ec05d417b41dcdc0cda54c56c4344a1bd0cd
z8edccf171aa5b8ea78032df2ef5b690221a224e758112370304ad1507e7009df66b32045376115
z82770199e74eb4d541bd0c3f92c7a4df99abdc33c081fc5dc428df4e8dd414acc661bbbecb665a
z1f50d2d24171f77e76605b1aa436936b754488dfa73e2620d805412e3ecc192fdb70f63323b85e
z41aaf6fc5bbb8f1b9d4126757c83e1ecf7910b2b99e31f41b17b37b810944d6bfcc18675f042ee
zec5ac29401f5fbc2acc004534f11613be6bd2ddd6056c67067c035ee8aa24629668aa5abad600b
z80abdc8d30618490dc33f6b16af5f4a46504091862fa6b44856da612916c7f5e09474fe8546767
z816edf9348e61995a0d3e7d5326eba0b4f2667845875f55c367f9c600292047a6061ed5272f364
z0a04b0411de31395277663372b11a07e404305ffb371f11eaea9289aa49d54f8cb8f4beba81ab3
z2ceebfbd75395cc499ede0a0fba02c4677396439e2a0febfdacb3c4e03872e0c1b9745e3b4e25e
z413f51cc60b1087e996e265d1c5baeb8bf1debedc59fd194e27665cfaa203046fabb7662bfa06b
z61b95ee508cd00c55581e54af21777ad5f539ebe6988434efdcf0b97b70872be80b946149a6b68
z0a8f4b8f65ca448a04b5163ad8026b64a2e8deae38cbb704703d681f7dbca5865adf6ca7cd01c1
zcca26f973590994d86483f4fa6a2cceb7ec28fd2994c1e4466c105c54f22c2ee884f18585bc6cf
z676cd240ee08506ff15b0479a417a28ec9d19024ffa355864e4731aec97ab1d3228325d4379ea7
z6ae018f638d23a10d6dabd82e8c65ef230ef6bf2f0c33817e5d4aaef1c6be2420c99a982ae4ba5
z0210b57b5538be189abc41f2c41932b55d8452c3ed0f99f9fbfb09bee7ac406dd519c7b0dc3eb9
za15ff0fdd7feb22f9ffbe7fe2a7c586d7889f82531cdb431f9d5bbdd349a297349a765ca5048e5
z02dfe2e50007965c9d705769d45c2852909d5e908816432d90e297af0141d3c4485cd356e4f4a6
za77772a9d23b4bd18e346aa81b1cc71a08dca31e77dc6772283ab629de011cb9442c5732fae5f5
zf0fba58f9bf2c4b91b3c3f4515ddfb177b23ca8fe1b0988c79b4e9b95a84cc30ef9e5c5c334180
z2c030a96a0f9f9ec5fd6dc326d6b1df6122ed043c54013630e637f527d19ab2d480b8ef1d63d3b
z88a3c50df516c3d242dce0998a44dcc65b56467a417886d72b5dd44fa1ea460d2e876a347e4e2e
z40e49dd95204ffd5cc3e78892192ae6a6a790070e57a06ace8c73fda9c0046fbd13abdbc7a88e3
z9d297836881af56c5cf765a3dc7e507fac14b45c342df2a6233e5bdfa6b5c2409f64a510f9a63b
z0b835850af0392b0f7e199575f0d7e8c5d92c6b309d25908e061154ce70698af72cfe497263e14
z3ee43cdb27ba907aff804dd6c44867fd407f95a1291d9467151635515043f09fd4ad46eb4f0e6d
z0d28c10f48232db02f782d0e2d465865e164328956a5b146a69c7787a3b7889f62d5b2a6606da3
zdb1543dc417dab672f614dc2b5a821d7d4f2bbae52bda434985ad50143b64cd4cbc4d36b7b193f
z925396ee25449d50c41fb4c72fdfe337548d7d518b3c8384e7a5c01a974f889887817d806a3bf6
z6d4d1eddd39950ca2b9319b6ef2adb845e91515215f60bc5828fd9096bf01f7a591d39cc6053b8
zfdd44fe996f3d5bb471481b8bb872a2c38b97134aa69b951017ee13beab9299a998a7d317ede89
z2f360bd6baa38779c74fb516b689582d30e8318cc337fa1fec3909b21bfcf3b4f01c4175854332
zd435923ef23f433e57be1adb6746a19909dd24135901f8592f077944f7839f83dac1334450fd90
z03fc0d145bd26d846eefdcb399ea69dbc1b04207be96ab81848702b9106c0055908f49c03198ec
zf9fcff9e054291751c4f812ee2354813699f09f11178646d54845528f0acad9cbaac14f14cca43
z9afca069cbf6da0a6918beece1124bdc2da822222f6cc70df97bb09b93a6d2267a326fe8b2e96f
z034cec66a6f8017c1263a2431e575108ba979645dd3917f58a520a1ae5407e8a1b38b25a504d72
z857dd17c0b64c0621a5cdf469773e6725d8a7fd516e830492af3946c66b06deb7ba17a33d622cc
z9b4a6b843f77e5118444872efb71d09990b9380fc61c21e4c16ef28dcc02d17eaaa67ccde22d6f
zdb284e5094e72b52c0e627be7abdd4ad6f78d2938ceb264f4e5122376990abc79f2ee53f08acde
z3ef5b4e634f2972e00e66966f27a530c6a0fad2628de4f04da0171e4594e4da40842aba4891767
za482c2c6fb6baf5515a8657f27ebca3658fc8ae43f3b1171bf9f40debc08d940ba419ec9cfdfe1
z17fc24fde95498523cf3587e308e28083696d01454e4a3ec89812735c679280626e556e00b914f
z2316718cc16b803f838b210e5e360787ef8a7bd4bc2995128eeb627ff470d7f5dbf09110e5549a
z49026c945b64d54d096d67504e433e62299c1036eb7ec526fd9d327c7534a9deba5c12c26167d2
z8b1089e13772c2393ec175e2a95a894c24cb6ef2f71cc310e31d6259b73e64c81a12837270fef4
z47c01246c4ae4f3095589348101e7c3867ed14e0f73c0316304c2f6dc703dec4086a0b7123ffc5
zee725c452f5f6ee93d01ee7289b086a56b86c7bb9db1618a1eb9538300b842702f976e45c793f1
z3b4a971e4e9b46d0a8701f9b0bd194d1f7fc58cd3016cbad429666ec025efefa2651ad925182ab
z88ca3d62b82219c3f42d9e5580798d6db2186a8fed946df40f224ee37cc8ead98500c3becb059a
z812b1157225d4f0c1c778d4dee137f61972bc703c37a1cf989d279a005ebe9806517096ad6078b
z4e43c536e473f12c05d84878931c37ee8b2cfd3181412bab980ff2e0f77b472fee99478cc9afb2
zaccd6267d3a267cf9bf14085417512a8240b8b7dba3c375031074df074cd7b5c8b113923986480
z4de0d8c3dc403aa714a32c5b9dc2fd315a90703627d9d86bbc251f0313c1cf89d8ecc76a8a60ec
z8b7d925ed6554763c8287395fac1f16ca33c00d6e394345b2404abfe2683123a7a82dd4243d6e9
zc9f8b9c5897cf5f00ba252d62746fb9dfc3f3ab11fc77c0bf3fa055f106897dfde0ed8853a0dbf
z9d3e89c2889b4b03a5edf58f325c9b48fcb4a78eb5a726ef6d9a42102cef434cb9b3df43212f5c
ze1e0482629c4c5227643bd6ab752a1d35639cd09dde2f275656dbabc98ea2fbf5088dabb7f88b3
z9acc7b844683b0a5e8dfdc76a9b455c256ecef610e1d216aa5f7605cf5d9509cf883aba887c6cf
zbc92981ddfa7d9d767b0e28c234975611b543a8e42b57d66ac098ffb617ed745e6f837a77398e5
z02a01da48c23977e1233cd1d331b04ff6cf80b042053721cc43604f5a9847d82288aa0c94a2406
z67b300e504701b91c7ccbdca7283fe1cdd64ed668a46a66d77430f6d4c14681c283dcc73dc570e
z0bb838e67987dc601ed5893e33284bea21b08f82f90d6da28c6928af853501cb0882d9106b088e
zf0b81541418b35e4d1b622bd77cfd0865178f20f9393acbad9683431df5cb18d38caec91b3ca1c
za56e041d710c3335da859412ea46d3d38cbba684125c230c9e893b3bcf579e2fb3ff38290ff145
z3993bc5cf7b4e1722ed8ae42be286fa086d85249531e491f047125c2b4600142fcfbc3ff6f59af
ze84a611dda37edb1d863e573fbd9788ea3b1e08e22abb3ef720d154ff7bba9b3ca74abec315913
za10569086cf058391af024c84110e6f4abecc87d2d4af75456c7511bbd9687866e4c5b48b531a1
z89457aa8d64533443402aae07109a1c8d2777f9780059b83de99342963d0efb6832c26c38fe58b
z2ae80c1d47ab65cc0031070a0f86b91212b9479fff9df62cb1741da235e414525221b768cb4cb7
zeb28dc85e47454401248159abd5f1855ba0e3d1fb2a1c1d3cf8bb1ae8f02b3869d4540a27578f8
zf850df8f661b10bc14aa5555b23462079ba88e6e75ece87c6369af05b5f898ac8cfd91f7de2a4a
zaa315f709a5c45a0d2a1c4480378301be46a8cef1b6f9156fd098f6b0b27f82ddbc43082cf0a32
zbd227c52cac01fd9b2ab9f97968205ce22cf7a9d5e014245e878d88462308751ae98dece1cfff2
z6a3cda1bc94e265c847bff48146bbe6ee23b91a43d22a741be1f5db6aff5db2003a199e8a0a786
za19cdc1ed24411024e4eb5bfd9058c061d3219f504c961602d45f8abd36dd31feb7d311bad1c58
z201b0d7046ed214ea724b4021b076644d8abfcc61e9e4d607b1214b88cac3177488c3fb60bb00e
za6d743ed386df9938f60f30ef8da0ea7600d9622e818be95d28a126000c3bdead45d0ebb74874e
z908faee3e9ecb406e758f854e3ab6aed2e5c3923cac0517d9382e40876f98497d667c82deabd0c
z6fb45666fbd2aeb2b4ae0ca87a5c978dcca09a9a9d276f838c5705436c6c22eb75637ad561f26a
z52c8306ddfea554b7e81ccdb703e2b8d50f7b4c44b4ae8bcbe7f0d7dbb282a9657eeaa4e46d715
z16a0c916d5db6441593343b2b38c9be96aa3f5043e53eb5bbc7c0e68247d8a6dd6c11df33fe5d3
zebcc92ff506212db65a306d9bf7d00b73c88c5df88a7a3e58d158b0c41cfd2528156e8b7d3c249
z1418ab8e4ec96ef6eb2b4c7bb03eac83e5746b2c4764177ff17b6ce2a77540253946f7e16e40d0
z276d0ffee4b07be511fbc3ee7253303684b753e5c39496057f2834ebf4281305a282f3e51cb3d2
zf52366a9a69c0806c3bbb84ae75793aeb1dc2678be1e6b574b6853322eaf8c4c206b55e8ff7573
z3f06fac5ec883b62f12333e4d9df33a185022d0353754e2e9c749122347c3b70ade483b1866b8b
z26f75a0ca9157de284d990b590607ae45f8d28568c59c62320ab3862a6d43afb53cd1a24b11f75
z7b4d07b530b52a6f03c6564ac9ca255bcb3030b4dacb9d325a32dfa6e5302838b6edede9f3c95c
zd165efd6fdcf3c93a187f2ed15cad1440915763d4cfa378593da013e6b059baccfb231584f8118
zb6390beb75fed2b402bd1a6c8508abe975e411b5019161664da87701eb811662a23882a415f287
ze5b5c4e7b32e9b8cb2e283eddc13fc25c669ea264d215520dbc46e506c7a81bc950920b62e3ee1
zb87adf0927146d33b031963c494df1f58ee197cb32a5bb57afee4145fae1680afd0e82fab411fb
zc88af3f32677592db5701e866c8e1dc00004643db542677c9058183dcf3422ea5b75ad1b22a435
z68ef8d5dba437f740e75d7bc87a3a3f8a78eb14cb91eeae3d6a5241b880200dd91e610f970cc59
z4ebae1a0b90f7879e153bdf8abf97c7a6c0047303d7b6b516d8366aa508e0cb8abf1b338b4c3a4
zdf4ecd9e6c7dfead90135c98627ab65e8784ff3295ab4221dddc2b9b7647c54c8fd27909817da0
z543183faeeb4c35802755ad91fba48178f067f3c1935ef42a0a525a091ac6391d0574449d2cc69
zeb76199f36d29fd2d3d1d58b0f66f44921562fdc49014f273e130b63dfefb41cce082aa6e3591f
zb25ff37c00e9624e342fc99a33d683306f2114e4780c78abeb583aa8df3de808afa381eaf0c21a
z838069fd02a13dc384088b7371b1e670caffff9e3bd03bd2f5dcc028b0fabd17c419354a237a9c
z8e0425598bda8b61ba1b5e734faf5eb50bcf06721004bbb16daea36f67194ead9472f3ca3be49e
z8a71e9ab8b382ffa3fe54ed6d0b7cb8d13cdbd56110d85977fc87935d0e0891974d1f65b83d35e
z15019802af9cdd114e520ea954fa7f5faddaf40f52998da66256a8ba900b36911d87cabde8c499
z12a45414341ad812f79446bbe544ce4d8a262b349b95f3e54565fce83bed7e58ea6f82614480b3
z0ac3a84bc8169c86913443c44ee5a2b8b319ed5f3193c1b20443039527443e681646248ecd5244
z4ac88023a60cb172c935d1dc07b0c12e3279426d1fa4e7dbdabb1330e203af9320ed997c80db83
z051953610f8575d3fc9336049036065b11ae250975d7d88c267d632006c234e53f5a49e6ad92e9
z71c083dc940d807a7b03849ccc72a5c1677fd4e92f75b9ec532754c0c340b996f86f7c092f0bde
zb82651b9873a56a04e0ae2877db9e310ec490edc44377f7a5a1b888e973a528706c2989c7bf311
z612e6f37cab82d5d039241024b1f9ff24f923f946e8c04e0091972846c3ea484e4435b88146984
za2845c0099d7176dbff6a5e8faeee42ac72863e8f69fd74f7d31b01cd135aa773f52f1fdf7db2e
z98e083ee0d35af51c574cd4574132f95830e8025cdc84b2573a1087c4606ec7b0e0c4bb8a6f376
za5c43fb61a8a6c0d1974250cbef8dd67f48c7d6b0bfc21f0aa72e963052a94e433ee44e6500723
zada3735c5adf056f6f5ad7f4241c17039b5bbbae6a6b6e47a3dc0af1db7a92600dc322ae07b402
z08e55c328b6c0ae5580430c4e2376f755b0d7e4736690379636cfbf8cf6b243d64e57466283335
z95534be3959871536fb32bb68e6c3f3f402deadf5c905c956fbcd3e3309cc140f74a88551a2c80
zee5bd73d683378ac46df61285ef3244375caef2612e3e63b3f62e2125bf8e6d2235a3171ce462d
z3252c9043e9656796e749ba87ee9ea80d08f00c966eff0f21b1598d82aa73dfb5eb78c3f867d25
z847d77ac2502f0afac83c5baf737776484ce7788dcc12f9fdc9437a61a5c344fc101bb005554ea
z8baecc03e6d22f9b67a90e039eeb633d1c32bae979e59da54dfe7637fb3000d749234329cc4be2
zc01ea03082fe6468c7fd63aef16d092e43c35003b042236736b39548594903a9ff80d7f89a720d
z268d2dfbf2a7e95ab9188f6acff3d0ec1aae67813a5c67a6a94355320c5753ccc0a9c5ff88bf96
z730c61e3d717ae818942d45579e9cdb7af71c2588b3b0de465aeb272cc8db8830faf269f0c8d09
z04c53e159312f1360a6528ebf2b9911527537b1cc9ae45b1e23a1fed111837e9ee89a9cd9e5198
z27c49892a4c5ee259e90b36743386469f6a69357701b472f182efab76e1820892e3be82296df9a
zc727180f80c1500e216f7c4180ce34168ae6e2902d5ada4030bf0d492a2e78b81a4367b561069c
z6e4351047049ebf539ecbec4aab6296c3e6e6d942ab6c13ab62e3941244c6423090fe6411f79b0
za216ded8d4ab2df2fe62882d7c8628bf58b6a38479d4388676f54e1c31cbfc72bf9454998f0627
z59d03c4c044f6e2bb35c13d2a832368457f91d3aaf963856a6f8fb2d7c57e112e5c87a1c180caf
zf3e841b4c1790ac40a564aa58af8a27852eb5172c072b2fd6f9efe39142ce32cbf5b6f31f794a5
z7b61b9934dba6af3d356e781e2825f43698c01c8634fe74881341ede87209fa6d5181e5273a84e
z19c8f97fc61198b7e71541b72e38c89a67ff51e93de2fd01e720e61ae42770c9a04cdce19fe491
zdc08a616ffb2ddaeb8b99d59cd754572ce162d35b0d1f73fcad46edcafd4429e15d08f88ce137c
z4cc1ba7a086e4c3f549578ce4011d03efd058cbced61a1f9ab2fc34f374821843e19b5d9e53c5c
z84a7f1bfd1b633ed82af5074b1c60f07bc9c0d6b604199e2958c1d8af2c392147aaee57dd7d568
z952c93bcbcd229e14bcc838ebea1349c0e90ff20f8178d6b7a84585064d4b2182eb8e8186a436b
zb87465676f9d8c89a673c0ac6c951d69409b51e10780e1172088bb4447ee7ae6e2e131b5eca752
z1d6d6b97f132bab351974eaba9e8c787b5e49238ded1c1b087e3b1087a923455ccf61561975257
zc2101e7e03bfb50f0e50e500d81daf1b73a8d2486111e7b4635656639089f843861b48035a7ec7
z48640be1e03a66434154ee8e98ced233a981fc1ebdcf3111260d48309b9cd5e327ac76ec742cc2
z352957a8de6fa5e2540d1b3a44d69539626f2c23408192a7525a5790eb439a48460d77008c7dcc
zf62776b45735ae39fff4a785e9ef72997dc88094abbee9030c31e1b584857ec25e45d77c960734
zdcd7ca533c2fbf666257771b5e1d86ef7d930632a55d1b2550df59a83cdac4f03e66b522bd59dd
z8c9889ba123ef8fd51e4cb62421d8050d2d53f065e7931513fe9e18f97d509a0213161c4fff027
z2c21e924d2102cafd39f19e77429ca31f627c6e24406bb4d853f667c6e442081877c62247f53c1
z0b07afbf577081380b51542a873672529386d0970bb3d8006aeee0552c0924d8df0fd7da105684
z346c67b756737cbe30d217a1f224a17153bc544ed837cb04720b275c1119cf0d9cc539009037de
zfd7a59dd12ae66a3119d154293966023ffd59293b86fa5e31279b8495c3871942fcd9c111d217e
z32b9ab35fe6366fb51897403198358b31d69e1acc6cea0fe09bcce31b4bef5d03c82e0abf9199e
z07474fecc2190747abd7ab6e33d15daaa2e1b443dca059834b3ce3ef236f60af68ed8156ddde42
zb4bc34164c6bb2e618b3a3f5097e87b4eab9aa9a172c712c460cc10390ea1d00126cc7cb4cd394
za4975848f947f6a1c1d125f1b5576c9352d63208346965e6e309d1c0cbda4ad2378ca5f47fb08f
z185a20903568513c2d8d278be293749157cbbc153403a8a406e48ee034dd597d233d0d98ef3c39
z5f890a52b22c69d836dfeb9e89bb636b7e8f3a6febac7481a43236d44c294da720d2edf1f9c137
z9fb6af93b4c40343e7dcdb9700b4d8bc7de82f2cfbe663f6c92d45c27e4cacaf7e869c1c12dff7
z71a8a5638922b575a0e4d673e4baf22c98f166b65f0f210cda665ca21d250b9712e8144acee521
zb4d1d6c66fbf3fa284d7a88b46d45ba05e8ac6f41a09f33aa14bb507af6996f29e46c93ea411f3
z9a51782707931f9a70186fbd5229aebee3fb382b7ef087adf62ea30265d90472ac2760bcdec2f4
zb789c2101e12815b384b6744ddd11b3001996b8c230ecf30f4a2695ef58967f13f1b257c0ac57d
ze7809f2c8e213a40bb4663bca498b87ef3e1990cc4e83b43b116c93701c94bf6c3a766d32413e1
z04429f9d4f6564607452b841590757364dbdadcfe6c6b086799e48893eb6807ab044def2d392a1
zdf0f60c157742e9d02c5862423980d02fd9173358b59a84da13771ab168a35d9bb8942f04506f0
zdfb6fadace58189125c02b5d35b881ca58adc56a993668738d94c9b0417ccd2788a0c481e40c0d
ze1b8f09879a053c55ac1682b9a00d4b1d2ac5876396496b29ab1aa10de2fba6d93f87a5a992b37
zd6c1e4b0b066d7fe2c3b7085270a00c7b39262971ca93cdada3887b78fc47e25e796589887f60a
z042ffb50f393c62d94b878baa85893303ddd1293d45a99ba19c61b99033dd3d6c79e012da40b60
z47f41a531daae2696e409393d68b29b73200b66be41d47c1025a253a7b8c7b9ff1008f574680a8
z24bb1f9e3ee29cb174449d0385c043e35edfeb32cd9b31772c90296a16ed951e0dbefb0b41b2b0
z8aae9eff7049f451ebb5dfee0d8a8be5ebd205ccb8e01711561b1f55b26baec2477d551b3a880a
z94a94665e8dfd94a0fbb3b3b741d555ec937f742b6b2057566700b66f90a7b6df55cbb0e6fa335
ze0fd1930002ff91292f9be844f5cbffa5c65bba793a855a417a8bfa2b899b8c15d8a6051f5c596
zb66fb46513e50630cf68e42114ff87cc6071be62ce8d348c9a1dba03583e79ca3f9043aa62cad4
z3dfff8008314dc29160561941730b6ca8278d981664def759d13962d88791344ca51dac3c0a0e2
ze80413d87edc09b5c1c002fe4e6d320aabb3893c1dda40b498c7e83bea8372b954e98a541b4582
z93c9da60dc08e7ebc721e6fd4d50a7184cb31aa7a8696367542a7a23d65c92fcd76963e72c8b10
z492f569b6d4d7f42c2e7a237bd42cc8e6ba46e2e3b5b24e460fb31ac987256a7369e62b510a97e
z0de062304208866df629cca08d270c58506bb3edccc35f42f5f283d110712ae63cd4268184a8db
z005fc7c2c8eb3ebad669363d156d2592fe04b320f9e195dfb5c5943f2ea43445160ef6a5d020ee
zfbb78a42afac69a26a4365c2c02cc89723d67f3c17c55d5174383a8a9d382afdfe0d6c9d6187e4
zf9ec500757893438272343687b804352806dd83e35c2ca716ce6eb111b75e111a9ebe96b1ed203
z9bc23f7e9bfa30f98b64d3ba2484225ad364f75a721f2aa0472142d9711eefdc9261cb3fe54d23
z33dc776d250d9676efafe5644ab111e3d45be958c20532a5c117c42e2b04407ad4aa86d577687c
z8e620a3945c8b3d708077f0930b7a0063ae2fce231a8f061039b6cf8c83e8d532de472232c6005
zc87cc269460fdf875455809052ea45e86f1b571cfcec51b278ed7ef2dc1691b1c6fcc565418eea
z73d3f3a1b99c0624b7bb6621adea86075e3f13d0d892a2b60ad3758d3226915103e2565d297930
zc69493503e76b2e3534ee2abb5187849d1f2dc5d9e75a4ffd79cb29e191fd3347586d0ca7aacc0
z071b6770cf6a8c06db7a2e3a8a09348cb2d4463debd4a70d73eae867b54a08c4ae6816675714fe
zdab297553a0c197f999456a7e3414b3ad24358bb4a2202064c2ecccc29213028ffae375ef29b9b
z8e52e4234cff03513c012f07933935447c03908b900d7c43992bfd97b18afd53dc728163d02d78
z984ab27966311391b84546a10186b42915a713339a3ef47528831b02abb9701615e37f418d40d0
za3d685b869a58f64441db7611fb2b8dadf3bbbbac69a9c88728a354b015f9ab436f7cab425407d
z67ccf80805743191616f509b6bbcae0abe520345005272b1219764ac656527122457674f00e7b2
z21a29dc5e342e043b79c79f6ebedf821d72105925ff448f02a10a9fa14fede744f3f312650c7e9
z7a08c46b7aab801840c372c824d51d1b5e4f465b84ed379638332644e180c1db9d608a0386adb5
z820df30b78ba369e45a33166b4965121dc36d15fdd12d56c3cf6506ace06d34d7def7387243d56
z6d7f54c4bdad54eee2efd427f99d86679f568a5449b5c62eef614bfa2950b3f908787133e0e7e1
zd0200f31a237eb1e60c61546e2c5fc5a5aa1c668274c2e75e873e0efbe4b77936b032164f783a2
z3e757e92e40769af4749a0c3954471709abbda0b171ef23eac57ca4260b7011f17fdedf2fd2dc0
zd85273e5243c1f8d92295d5cc312adba4844ad0c88964944b869d7abc299fdd40a62f8d945bdaf
z46f7cb2ff0c509528d925410b6ee8adce9873f8707dd93477b0205f4233463358a9c818c85851d
zfcdbc96bc62329509db6aa21f5cbb2b64c4fd3154e39e9ddb0cd2f1257ace024141eb70f091f0e
z39bca00c66e731c8566b385f95fe88a3085140e1187a64114b7c4c35e9a4da226353ba14fdd186
zef39db2f60420ad64fb5e1bd3452d4d56251928a113da63f5164eb38794b653b425086630c17d2
z96d37d877ece556ce4f772bd8964a5e9a2b31a6c7ccf90ed1db676ae20b8255fb48e9e7fdf9be4
z6322818b1b8772dcf4ef4ecfc94a0a3c63f1c67d9b9980cf06228b35c71b70b67e49d452483048
z48499c0ef655aed4afb20eccce22d3d7c0be99496b3e3cac9d486984b7dcdd2f06b8e763dd2e3c
zbc667f20271a84c932518dae8bd097cc85f8b2e46baebfc57425d6ac72cba7b711e265594d08f1
z36a721b68e954be267d8241c99f26736f2118ffdf346f372d472a51a89affc27f7f2a8e2c453d1
z58d3a4537ee8005a2a84026ef9094585eafa2e92f6cdc38a104c923989a62823ad3a5873fb8e7b
zaff763d0c6654287ed76712ab44906c57fa1326eec52408cb5511323aca65e07b5961a20879a08
z3ca1e836b573f06ac169ff60032848997ee40c8ed0d68a7a8e9d17d78424b67fca645418ad9b06
z79a85d6d98b643de8e192228813b6ea5f1b48c480f3fd7f0825aaa1980e7ba55d617028a302ce9
z2b6c3ca767e613cee2b30aa551498e49b72ad9f872084e59db1e06f2db25605e77a4939ea7ed9c
za2fda0f83d87a50b4ccb0547dac362d8944c0fa97e535dc7d80bbccdc73892826d4590de155a81
z77ab6312834fa7bcc2722f41980a1fd471edad3a019925869bff2d766d2a51fba9650bdb8e05c2
zed8882b5f6030675e7d35d002bffd2fc7f36e62c2ddbf3fb34642bf8537b8591a790de9beedd72
z80a696019e7467d16bc40ccb41ccf69d9264aaa0c5c7016c2c23ae3a3646cdfac8d92b15d92180
z5e05b2c2ebf8f455f79f5f75f6c13947aed068519e60b260858c1ca8c8a4c3c01fa755ab10a90a
z23389b84e462150fe8104e14dc5bb9b4cb66400a1c92bd83f0c0835ece871626bb926628ecbb28
z774ae9d1b6c7c50655640c7ef5926bccd0c1fe6fddab6966dcbb8bd266c55570dac16ffd8c7b1d
z524884937e42673667408a5259f51ee76a6ca7203b260f08b079cfd7f8d03d740eccec429b289f
zae1f4bd37b3086c0eeb23f3e14995187053ec905c0d3149f72777d0d24c5c3b029038ecccc70f6
z157045e2e4c1d51cc890310982e630cf430b67a35ce515a7dcd54c51a5f1247b9526c26f45f9e9
z22c4d763d73cba4447c99a83f87b6eff4099b6fa7a96319002a2184c96388f180116ad34fdc48e
z41ec4fe7661f16ba130a2409c72f51c7986aaeddcc15cc8ca88cc0cb01ba1aded1ea17c067571e
z1b842e898947fc0729a64a6866318ed270bf3ceff33748a67e7058643c7994c9faf04a81153099
zd01723deb276522c9400a1b96ae09360082f8c79fbf5fda9fc5872700d71eb9c7c630c43e6763a
za981f502a36b01a235e78b0c53134bbbcc876cbf663552b31c1e1c8ef1e483a1b818309097fc3f
z8c5b7871c066a8ff6a94f3f251392ef2bfe1f903437a68f7641ce0037d310f0eb00fb5c4f595d9
zf0b451821a001ae55aef81405008cbeb4c4a35acc3a98510fbed612f73c210e3c2e16e602eadb8
z3c87705d1082e419729d30c1e8a7f13957748d5b65c42eb3356ccdc1c8cd87f95011a1fe9eff01
z634d0e381fb76dded4316758591a0a48a7871b9731b17652298602c646221be0b3ecbc7c55ff9a
z7ad4bb111f4eb4aaeae80c8dc251eed43de2d92a6a707d2ef21bcc5eb693e2b38380e321788b91
zff125d0b9e7331772897d5da2537ba114ac94c58096d575f5020956c51f907fdc38c8908dd49bd
zb38c025945a6b89d0c59db690408b55e587c37054588085cf2de6b0f7637b5d336e42922310cd1
zbd1fb8c747d556e6bda0c835e254d683ce36fbc4e54e08a4a210d2ba40b069e823fc54b179b7dd
zeab6537250aca97011f70198a1cbaa9cdf51b4ec52be9e58b009b42b2af9e39675a223747cccee
z820517f4d788c0682e1a19b2f9bbad5b793731e6991704376ca843bb469b6fc878fd2f1fbf2420
z868cea9c73055159ad8dd9481a1e45d85def5977e081c7c35f91c949f51d253875a326da385ca6
z80a169ba6c395cbd9d2820cd4e9d02f6ee8c8d04625dcc1ad9df3c5380ac16d65f95b135392703
z331d4afb84985b70c71aa67afaaef643d5232e2e219d44fa2ff0a5f4997986a5b223bbfe031c70
ze8b12087b8dcec946702feb0a21a107bf9e88a702d291faaa06b2c552a120fb11769241355a633
zddf4c82e4740970d3cad7d198c653d085f1073934408583b2303356ea79ad662571bc5a265d6db
z0ea375371f1d2f6e25ae026b0e702e151122c736623c3ce657f217b7890db6f7128278f4d23cfb
z5c71f9487d48baecf1ed83226da33b6069d24d75e40423fb5c5279d6891a71c94da4b66e834710
z76e054518dccaf10aef344f8780f76b835c19bdbabf2dd7bcc4c162bf90fb7dd426c37608c796f
z427762566fee6dd3b60ee2b55b5c6bb522bc19addc82742b7651efe50cf6d8ba5a333777adad6f
z4996d84b959cf10cbd2a96f0348c9114ed2eb20ee667b312fdd7d29f4958b396abf228699b9cb1
zf196dfb3e21f0b8020ceac14d221a0b88d5c38f89229d2356a1d7a8428381ca5b368b7ad4ba29e
zec25b4a975a4b9356b61da7ec62609e6b1d4c946d750b31289c78174158bca842a2b14871682e7
z9b0dfe1d04c2aac2c6a250370c45c6f3962968d86d6ec487c7b13c0782232d75dbf164c0ec5422
ze4ec72f0f951c4b9b01d7f05bd2be416225da51a7d9d79d4a353e9cf44cdd3e2bde9c3da6ef101
z36f5e1b32335e390211f80f006774866de9251186d46fab2dfa2bb3ddb03401ec65d5aadcaca25
z73c0d698b4d642b700f075ee834968e665638c365d984034d3d84ed4cf37de2a3a247109b528f3
z521d6730e102480a3d18fd152562e2cf75a4ab042e97f45476bbe80e6ba72e6a0dbbda5c119d5a
z84b3cb405b5c2a542623b998feb38faf14a19e9b92084db892fc5830e6c55422d75d89dd696db5
z97a5360947a296ce4bae60105ed22669d58d709a19cc1fdad317e774747859cab6ff0b15be32d7
z9a530283486a775713cc1f8d37471e28c03b559e38cc38a5709de90a30ca3ab435f836e6b9864c
zc5503851026991e5a7011a264eb0c2b35989a34b74bc64835ea57d032870e40d2ea7ddf3d5f9c2
za22f50d2d427595aa880b44b76b17e2b627836bdbf0b6a65e7e4d4ba3ccc824578b913f3dba7b8
z29f779132ad3a5675926697fa2baa2eaf94d5e3600dafdd95219ee844b096c1ed6980f29d79484
zd2ce49463bdcedd3f74c449a123140e5f5d67005ae6c8796cb064d17f145aba5106985af96e492
z8c684fd172010252f0dab6421b11dfa058f37cea99d0fd1d618e3e9746115f03c43db7449655df
zc0116a8401ec25e00df5a1776027fec37cb88b7900056715715a6d4a01b03c1d33da0924166db0
z2e20b1ba84afab9e500276008cdc1a0c12a99c916f50de9b4b8195aa512a9b0ffd774ea7e920c9
z406b16e46f4e352228001feeed680c080f3d835f671a6fe7b12aee0594c6b8efa845c653366f9d
z0ba7222d92e2102ecbd86830bccc0d81ebfc98753494e83b83011a6e34b90aee8feaf7746c7eb6
ze04ae399fcbaa50b9fe59d4ac8629061d00aa8289f052b27fae77f38ba80e3c3641e8e6719ef42
z5d7ba640b7b8d2b89027308534a3bc2e186725f2c296d1935b3d91f6eaa12ae08aaf15dfbdaf67
zef4d15c214a8f8059953dd30f597bdffcb2ab3f2ffe0391aa8561522b48e236f7541ab35a63a40
z80e69b6a1132bbb252c1297ce78a03ca3fc1cc15dfe651a5c00dd28c05d487a45392edcd78761e
zdbf53d1f7ffc7066ef76e3670a350e52735d67a2dbc8f24b8651a719599ed4874523e6d8611bb2
zd2439f2f89fb05a8cfffcb34f5ad1d558475b14aba0bf5c6e29cf912193a9518848485c2514047
za433025a9220afe5a8ee1ef1c22fa5c20124fe68bc90868970ceaef8df726ceb1d16cf84c81d49
z7e7757971009bd38644c5a7028551de1ae4f491b5a2c042a26a2db9722405a767d0b44c4596ee2
z3a4657d4f1f47cbdca8034df83afd5f32d8a230397fd51b8ebf3b6efe5643c9be49fb2d5121cd5
zabfa840235466e06960e3e76500536ceeab809c2fc57d37ff2602995a81f2a017743e7fa954b8d
zfe0b8d27e7c9ba7e35a5d48ccc6806205aabea58f002d302ba05f3e6869efcf0251ede5d9e1671
zaf045ec4d767c8a74032e9838b61f294bced56cd393a8d8c6d59e39c5288fc86aaef92153a7d4c
z8fe341dfa7f0782777e19764396fc2ffaa31899bd43eafa67d6e4c0e317d70af80b5679568487e
z4856ab77a0d230e00e8050c43ebec0e82c5733698fe2b8d90073a885a3907320075b11d4a7294d
zefa4c9463a26a76b522a7943435f0985bd20df9056df26ece89257a284885bf4b711813658956e
zaa148a3db40899718a90cdcec7a83c353704a8a443c51a9c3c2e65178d56c2c245616336acfe3a
z5bc5567c3d4fe4b9b9bc5def3cbb10ab8f70fc7042dcd525afa18864f070f6ff7313845b0224b6
zb54599ee3b62e9e5a21a46e4e483c9566ffa8dd033d76cb8250965958bf081031d43ff0fb02859
z8d30a304fe97aea546b5a19a42525b856463de2475afe825bad9379ace28f37c94e8f06800309a
z90f6e4cc20e1b2d0db48ca008d2bb1e56f702bf63e2d9aef10471a181a6ba3b6513926326555f4
z4cd381c508704b882ff396b9a12100ec326e67f5410d2b9f1835472c31dd63fd30636c2fd9d342
zf874d272d452ce6e9438f81235ecf2546d61f6df1822ebe44922054bc783cd910f5109687948d5
zee2c741ff31cf0b000567757be12bf22b46e67865e54c1612125b9fcdafc7e20fbd8a76ef30254
z22912a3ab2be00f6820b4aba9e829f91f5370a8983093f7359b170a3d71a516cb709956bc8d775
z1885705587cc43adf3ff9115dd3750871e2ad5e4d97fc976cec5dab0576141cf2a25dfd20a15d9
zedf7c018b54d13c8a5d33cc977d8d24bcd87333535f8ec4dcd774cf44a2c2561a81e02c6531146
z67e2862dc2d6622e7fe09039107d29e33425d9d005dfa558ea7fdcb0f9cf6313af8afd6e0075f1
z721fa1b8e174e111245de3252c4ff86bd096f6c99fcda982555be186f5ca82857c6083f32c3a34
z853a5d8638fc081d62d69ee0c020c7b42e0d85d69273c9f4158f516483dfb946f7744b3c55f3c0
z9e03bfcfa265a0a4da4c48e283dce1ae355a9907c407158378d929d71496657c2ba2c8c1fcbdaa
zfbeb76a7ec4c889d70ba4779fdb08a7a270578f155b0a7ab9c2b7a57dde5f7e246b31020b58957
zbda8db3a3a988337e1d78292d1314122032874ff2ff23f6c54a398871c1191fc3bace1bda55676
zb41bb934af23348223c3be272043a088a1d0a6c67afe436e160e669465c8148f008877510738cf
zc837175801ac332092e94d9fde52a782a37a4b728192ecad78cbe1c2f8c1f7c91a13a9f8cea055
z874b75fb0470bfcd05226c365e4a857fb3cee3ead15e8018a40944b72dcfbe1cd3c1b03162e5bd
z594a48644441bd1f4a263b281fc216531b13293ad5ef4d72eee00355c2aab554e7ee7782f49ca3
z6d25505afe4ba7e2072cb35808780c118eabafc5bf9067710663db4cdca7f4e06c2dc22c0dd8dd
z2a2061e4ef866c18ed4777d27881e0c727ca5c7c010ab3784d6a19cda5a981ab2eed4fdbc0acf3
z5dc3ad6cbb8e49c1bb19ee54a224a34cb721a5459b386d60cc3c16f4db5f1c314d00d7b064626a
zffe14636b0ba856e2fa7d2dc704afe1d7c6d135f48074d352c2ed5e60914aab2a1eed68677d3f5
z5fe4d5a51afd5c9b98f954c2b87757faaaf0d270539609d7374d26626a7383c9d10efbeb0afccc
z2f738cf3931af09d0e6dbd31671597feb2208a2e719a406c2da42fb1dfe63edad42eade5dee26c
zea54706b2aeb3d88c666b409960e1d7e41f9dd3f37898287fd560ed3789db2c4cbab61d6545bdd
zcbe68e6e175d3efab53726d84cd05c72442a68229d7f462fc5828ed166a427398d44b50ff80d68
z86e488b0e53181ac368850fbd795e79eca8a04da840542958778b6013db170167273f2add4130f
z3cd62a9d379e9977e53852df2d16e3de0585d943488b9a7940bd7ea372239b8de9a8564e5a9a29
zed869f25cef3c8e6fd51c23fbb7be05684a47b9d36e88220c15ae09a1cf77425194b74b3b5f32a
z5f469504f66fb2fbb74e1a8bd3c556241480d9e2896e6ce9ccf0efde48033ec97a5665fb750869
ze015847724ea96a54c98f4bb2ac16f3444ee2b3bee9350195bc27d6bbee7e3e50eeb05572ec45a
zde2af7e4fe806d0f72e9ab3c19f0d0f4a5a6fb8aa6ab7073bfd1c96df8b9d48d9b90663b15ebd2
z62bead2629b7b46293dbe0bc9d1a1bf66207eeae94ba1662dbfc93a45d4742a79eeec8a2565996
z0ca40551f91d69a569dd3bc71c320bae692e766a98425bd897ad1c749989b78fbd05aa20d4a193
z56afb9112b878bfc52983982239875e5c2db394693465b690b806204bd80d49bfc128f8036e71d
z2d2779b64e84ed682a0a4ab1d2bf37eb11e7fdc3b15b19838ee108830e28d12b670c21b4b38e01
zbd53f76da1d04c9b01d2c1b27ef3dce6ac27358927647cfaf23740855310d38162ee0339262561
z06f5b8e69bf9e83cd700b805b19b2534bd757a90076b17ebb23b75e06bf5460d5f765f3442a0d8
zb68b42b0beac6292a16d6286f1358ee78818d6a6e8f932a688678c818725cf0c6adab3daf0245c
z50ba1b7604d7b69965a4edf9023a36f80f29b9619bec2b651c2b1f209b344942c023e4b43274dd
zfa65692069a627d0733a7e7a53b099f24f671c1a88e436b29e7398971e21b6b7011b5d5ff9832f
zd1db099de287d51d6e2343ca2df7a7a82b418138f25f56238a5cf8dd1074bc64f4ab91f5ccf53a
ze7b6def460930008033d94fab4ea828e6c4bc2624a57f17252f660570ebc69ed5b67a40e0a0840
ze0e7b5dcc0d7a9e5b510262e4001003af9899077132ca937ccbce629eb56c1c4874b90aab6aedc
z1db67bf877024a7590cb72a6348e99db0626874ad9330f16fa48d296d045ac1d4c0caf9e2d9cf3
z477b6d47fc501372cb0908320da9ffd154521777c7776fb46f76f016596707d6ac8e5862c2dd35
z740913cfbe0f6d3d3177e6da6a89b0ba2c4a913cb91965e3183fa5a0639c3adb652d8f334babf2
zf1df1655c1cf5cf56c4c937384dfe49926e207475b0eb586ef3512d07f9936edfca3dfc86547aa
za6d387e04d4c07a5ba29f79388de14c26f4aa82f6a6198e682fc65a827cb298b2e80859f3dd40f
z25eef3b4498424f5b7048c16efddf6fa86319403e65721c933674bb90f3a93f4b7d62d5dd2c3df
zfd2cb21ee330130a3bdb6d94bfe2f8dc65c81b22e125556a197e6140107b58b5c65f7a618f7781
z376778d9a9ebbe253b2d7e15fdcce254a11551a29a93a3f1d17da1c61203241f72c83dec0fdd55
z810facfaf47619e0ab8d7f837f0191b874af87e26751de5deacc3fe00e7aba638fefa25154d244
z1dbc70882a990e20089d387be1444f24134806744fe06e1a33865a9c273e057ebe99ca2b57fd90
z08baa5c2fbbebb29b085228d0aee679716408af52062169af5e57b1c470ba03f3cfb7028372421
z1a2c421e8d8874f800851b998e602c3939f5fb56969c7df39c84e251c7abe4e1b1b680fd3d5585
z2192c05c269a3f70fa19283e60b43c9656a74d71f9ed748e55cf2f7063494ccfc9deeabe25f52a
z36944a9607813502dbf806deb4661a01eb67e1065eba3e216604c56f1292bee33f1734c199fefe
z7817d48cbdbe2ee9eb0f81d617ae7473afcf4b34f68aba26600740867589c94ca6de9254d17d5d
zd05725019d60871dba36878199f0efdb13b281d425923e5915577f9d9c2fd493e4efca78487eff
zcdabbbf397db55a016e6c428bcf4dcfa8f04d48fd184d8b431063462964cc174335bb4804f1b67
z17fcba909b507a0ae627533e15051b3358a619addb57d6c65af7a7ed10691b114c559387889c11
za28f36b9d3c0e8ac7114394d5467eaa63fcc85ed1afd6604a4260762554d8afdc71c659a70c81c
ze7cfd71a663ee46ab0d2f81973f60548140dcf176c8a6b064f090dcf113e3b2722fc92fce251d8
z10b4baab017014ce2f7738498d7bc98758180e7651de29aa7101c02f6414de9ca886238da4b4e0
zbf803d7dee8006e12b71dc02856db121ca4d1bff8338c4b89b3f4c473f4026651e9e0b4fecfb21
ze6c8e8100e453b77a2c267bbb4615c29c0b6116ec9dade1c3076df92989a79a7b076a4b306e378
z88979bad855c551b69fa2a259bbe366f4393b1150544524465404112923d2b036bd3b4d4a92406
zbafdabfdefc09bca866abc510aace9b2f637ebc9a42e96f6131b216222ba918456aee5cb254f59
zf9bb1a43fef080fb1dd5e696d249077b444d640c9f962f982c92aa94974fbb4b6b99758cd17830
zff048cb62243476753deadcdfa34c55f847cd839b8b0898dc60b6706ed12fc6eb24c7b01c544cd
z78cc561c7447f76f92cc243d594fc991f0a8d16fbbd73e1066bb497a7d3fa42321547c9542eb35
z1c1b9d2c03920ae1fb59af1c84898f4bfba376f27ea9d442fb7812ce15011b518384580a37bf60
z8ea7cc5bc505f36debb60ef867e1edd38af597802beabfa5ab816236073fe7f8d7b280f20b46ee
z5de61f97c0a299ef6b0cb8bf0dd970475626419ee7630989b0731bdb91a9002c8c1592dfb77069
z248e26a6058246bd3341f110e4617afdfbc4557d0c1503942ff87d3ecaa334ebfb8979c258e14c
z1e2b8424077a5657f19758c66441ae874a4ac0c68743f477463a663804a7fd48fa8a2c0e590466
zbb1b56b5ded2b4ffbcbf791aa649e1f357a17642f4ee9d17bf3ab9ef4b25932f0bd56efbe01932
zcbe45e3231c4466579e644f3c543f7cd4ad0a54cae39a8bb0b479942d5f05aa9ef5108e5e8c58e
z02b788a9fa8e050556cb0d0a043b723d34f6af1e96560462e16563e80c9461f04d105b05905ebe
z4daeb4dcdec4c81ef5a68683db0c5cf32b8c5c76f9a4df21772424a25d82ec91779ccfe11c6b63
ze6229c9fbeada387b99f634af7c6f9cf4890881880e925b04b648775150e321fabbfd04ee759c3
z649b9842355de9bac0947ebbd4c46849083a1fe6d48cf432afb542dbadbf916fd11e27129d1ca9
z64714c334ee603db11fb86fff90fc7e717ec0d1139bc95c808db365c5f5e22c123c336d0d7ee70
zeb48d50f3c7c4a92daa89b18501c21432f4145d313dd6eb84b5989dd5d27d255b6cf82537efd68
z814210d0c689a5bcf74010b6820143ef339adb6ad1b28c642ccbbc68cae7ad67b12cdc042b587b
z62fbb98b43e085c09d2b0e6b2e4e540c3fbca2d719dcbee2b1faec0e05cb65abc20276ffa86466
z21ed9c596b3c46c284834f0ee84e26b5c3951034c0493beaa48e892ac3aea765f55b1d941e08d2
z9dcc4b05d918fa9a3f4c7b639af476d57630922733d55ac46b92d0c4a656f3cb032de61d581ad8
z85602323202bb850a5826e745d5931762c894df734b1c69b2177a6906ff046278b6af4e334d0f4
zb2e719e34dd0b25b75a860e0856cf301b7cb0c919c2a9e9387216170cf983d5bc58ffc41cf3553
z4e1fc5f0cbe74d4f4ba214424ceefdd0c282bc4dfa48262b88698a55aac94bdd11f665b4657392
zf394bf3370841db5f9832f6e123d976b243d195fe5a36d7c0b7024a0a1b583689ab83563d1496b
z27b0e0dacba9ee5fe9c5b5e44d38f1d0fc9b5fe5182899e52e90fe76566386a88ccc0ac52731e1
z0dfff36ee0f581818adf95c5a3a43dc4e3e518290a6636a95f75ba933f92c10c38e7e5f62122be
z61777acdcd82ad55429163ea9ed8b2f3c01dad029a134d566847124281d58e81ebd8d924875582
zb5e04c67548e7105c2398bd6969329ebd9edbb8cb6074910876c6d37b140468abf08dc3945f7ad
z19c18e4fa8a67641b6a94ccf0e21c62971f796417452b0467640a14032bb4e77edff9be3a0b48c
z53a1fc871f377510a431dc77628b96f71671ea4839c278b4373da37f86df69cd77950c3052de94
z595826533bc939182887f544f9b2055b9d5c038b04bbd55be544ee976f8b333dddae8712d6c6c8
z1ea19cafaa1476af75b4b4423bdcc803e97e6d6f431037914c312a4f7ba69e542362830ede911a
zf1352c4626240e79412d08b08a8369d03a2b80825b7b52d00cc25c95392f5b002c36ff3dea4055
z9dd0f54dcada4e2022a4d513ddd9da82f9c86d8998c99162e5b08f0908b00cfbba4c18e6cd03a4
z97446d6573d8d9268a4242a6b730f67fae69bf423c303c90d530fa7e0eede6c5c9cf773aebbdf2
z38c2e6e1209950ff9c3573a5d75a361a4e50c49b5dbf7a314cac4d00586f7433219d43d0e9a9e9
z8aaa8597a010a7d6bd890e2ed3eca23d0091b4b81af228bdd753bf84fec40cb98c95c2638a1ede
zee59cd7af0f34d1dfb56e6c3f1027596a0f178f66539208e44ad0481bc3b38b2cbb61c874912de
zd4ee4090d42e9329372bf557b8a1f1665409b3c17f44ec4fc083853dfbaf780008dd0ad7c86686
zde1e62f330ffa67c698e98b02c8b35a0accf003bcdb6d4d7f428f3806b19d178c871deae7b0eb7
zfc7576d263db97a7e52ece68e09c0150e8a47ea0ef4b814c9d4e43c5c8475f3bed6358608f9462
z1e75529167ec39de432ec279bf63c3008f5a538e31dd4340a4993542e379f7668555b87d46ab8c
z454cd31dcb785eda291019de0d0863cf302463c78d53fd680296de89a604a6c1ab0487bc482def
z48fd2b85c1d01a8f759c161d066d3523a181d56cda5349dbe2fe1c21805df33368085997f93efe
z6cfbfff19e564e77734e7aa7d3d38d65f7c8b0f4fae2cf7b3f8a12dc87755ad69610e8a1a5d677
zff8c67d6f3c3d4765a33ab7ef9415427684fb48b1eba67943c6ead36728e6ad25cdc43aea06816
z0fc8691d5cae6a43553dcc6b5547be7e68f9be8d3b4bea5dc78360ccf95c985fd12b264abc1703
z165566ae4a88bd684ed07cc4ba809487d32ccbf0d639768efbd62f8293d5add8d9d8dcacff301a
z35e4de254e62addffff4b79a33dc3ab981f953096a727af1ca068e8311a6a25f212804c0b50cf3
za5d53290ab0b256c40fedad2d6f9a1b797419a83b64ab738023ed86fe422bbde5c7a906a990c1c
zea590b8c51cf7942bbda982d959f9bde51c9ebc1ada5a8b92938208409e1cf52e92dc7d4e55b27
z8e47c85ad18d25f9a8cc4157c6198d93b3a42538425c2c70352f7cdf3cbf01640da91657a9fcd5
z7643f7a71ca3fb87c9aac2c0b7e814d32e1262978faf28bdf217cfc2eaabe643ca3990746bb643
zbbd7905c76416a19775d7ddd5cb13fc39d8a5b159bdbf15a47f31cfebbfe3ca526e8f40ff15822
ze0945bfb8fcfa83279845a5a334b344939e4b48a275fdb589571d22b6ef8827872493310737d7a
z6dda67b7e636cf824a2d42588d8dd7d5f9ff4bbad97015834fd5856f99f8202dda12327109ec20
z1aeb4912d491f78622051557705a0c407468dddfb1f6f6be1eb23f6a21efb63399ad9b2dd6c69b
z95a3f8e6e33fc6da69951b33328b1372e3b49e53a32139a4060b382826d001634e988a6fac3064
z379e01894acb54db56826dc37011e2b6e7deabc53366ea1e559fc5e80a8d7d3f490976d1f55fc4
zc15f27c65bedc221d9ca01bfc4889470ca564a638a8ee04df3bb2c6814a6339554eb41e007b56d
z751e12c2a0517d6242330e46d2751b4f54f3de8f0c19e2d8eec2f3cc2a2c58be24306678100b89
zfe939a125114ed73de6e8c3e9b0681428ba42314a1c25262939bd69310fe0f6f644d6933ff74cb
zac5bbe228603abf7e07f8668fbe9c7888c1de98b3aad2fd7e56b3bad1f58055f682049844d8157
zc01ed5ac2525e7349424f85cd59a21a07675ae372e0e413ca4c415bf5cb2275fabb28a7ba41f56
zf89699290f3b09a4baa8e8fd628b50b1b7b2e8ea469ad924cab239b03422c81e4791621186f06e
z7df78fd9153cf86543ed808751b721aa5e4d3aa0e49f2f8abbae08ac04f7239469cd7b42eddd9f
z1950820b650e2acceeb778c9e8de705ab224126a0e8876e6d98a6cda2b05dbd12964e666264f45
z882c489fa0dc61a38ab7d05344ec25eafd059e17dce916595e046eedf5189700bc1c9e645ab312
z9fff8ad8e0f5a028c01857bb8a8e7ea5626110e088f2026175a02e13f8e1bd665068cb2b64e23b
z876f82b690d80bc25b6918919712bb53278975456177e3fc37bc8699eb04161c1f9952ffd24ded
za0ee81904fac5f11e1e1fc6e97cfabe62bc649ff8c18555214bff33080cf1fa66ff51f75b5247a
zfb45af1bc3fb7f7a9140ca474c39356001d7bb380d1cf3a9787c06b98050c0e74c37eb158b4e86
z439583cf66def6a626f6cea60375e8a34ee011345d0bb95e9315503733ee3931330fcb7b82a890
z45568d234645e7004b4e124dbadfe51eddf48c26a95b0260e964c67111d1e9ed2d0a0c3399d6ed
z03a65f18469b6c98fa6ecad9cb965362d5265ae09e0339c3aeffd20fe356b69d4333d62e1e2edb
z8eb06e99c12f462ab543e3117c7d1f5e3ab6dc12e924698edc59d1060c4e7c538db707e9af9e53
zcec1246c9e70edeaba54a839335efb441dcb8ccc58d6ac79b1258704c941115017c8d39e010dc2
zdb3bb13757a34aded867f0a04d3e053d061281ddccfcc99748a0d1b3da8aaa2d24b675583255d1
z5e179898661de9c02339634c8ca91895470734a4821823fe0cda931e236e6408cdc36456598198
zdde03cc821b7613b0ff2648562e7a1482031cee24f1f8da90287b60620a2be66afc01cded5ce04
z015fc36ceadd060c6d8c986a7d4d7c399b8094a6dbed1a764ccdd04eadb08c1fe99a50b582b95f
zfa25830ec1298b1cbede44963eaef70339555a0c88b514d1b59f4a664543488ff9032bfa0003b3
z253b20040e916d4837b928be2284d3d3193f3d821a1905df95290583fb7b5b7cb911423d7a5a24
zd7a5e98e755f44b2a58e9c757170f0f5b125ada5b4d66468ed44d879d3ffab8e3a2f5098562bf5
z37a72da7594a9cc774579f7687ec5996bd0454fc428200be6b8ebc076f97262891cd538f5f505c
z52695166505a7959935be09e3ea8d5ba3ed6fe858f2efdc08e3c82005d9b1cab5bf3fbeb13791a
z3e2283912b5a160256fd3bca37dd1774dd720249352725b885ff135fd2ded4cb6562e13671b8b0
z452fd6d81f295b865b568855580c0d33875150fdc8cbc50ac9cf8a9900abcdac538bed468a8fd7
zfb57f31c126e3378b15a8211141d78684e3914ad9e48559287ab9dd0608b4c357012be336ea0c0
z6c3fe728059d14a7f4b7eb4856e2f16ba22daed97969367b6ba9b33da2f7ea7b35cd1e589aea42
z9ab454c3740d1fd3654529846d3a8e4655e8f8bd718955fcac46de537e6834401feb28202c520e
z2e9114cedf9303a97c6c59541db29718cb967fa9953bf68a91c6ffcf2a317b3e9733fa02d15f5c
z3142ec7ae9e3e609f90fe642a232ea986ceb71bf2a4844660bb7b39c4f586afcc3a9bf38af8fdc
z2001f5cb68e8757198aad546691ffcade9e454a89ac7549f1a974fd59e9d07e9791365e041bdee
z116a8b564db5ac8ee4152cc7bf98bfaf9f4e238426ab0de253d26b92fc8278820e04bb98cb97c5
z6baffa597311872aa8b7e57b72920ed6ec5df8bab1e644096d47edb9b63c6d2809aec153152ddd
zaacb81c62d0887fc01d3e7121d1a1bf9492fbf54c070351c5213c5df2ac9f19cd3f57100582349
z0c93428a9eaf954fdbd8a38bdb0d9bc1b9a1702acee4d501e8585d7e341d19c1b7b49c8eda17bd
z1866e618a440ebe9f2eb9d1809c07456adcf33dfa2148594aa734857e5aec550b5b552f5f06d1f
z8cac798c6af081e1d8bf11c686c9a94119aac986e14495c78a493b4b3a47d31a7738805b5d2abf
zfe3494a60f85fc4e1a327faf014e0ea719b0ba6dd413517ee54aad2110c321aa961bb9460cde6d
zc82480771ff99d0d0b71258dbb933399a9ad5a0f3cb283e619f06bb15c10567dbf3a4fdb9c8cf4
z6fbba0f6bac2018712d8f20783397020ac57931789da8115948a2a8948f2cc987a8a635a1ce6a7
z58376b6cda435f2cbe1b110acca1a8c79049e3b0df052500f7b81fc5457bbdb450eed65ad4d517
z155460d7f54530230f7b1b3c203235a34f0e141dd9945dc1169544d835ee2b3602ebee9b506077
z301d716a9b7b98f148b7f93f8ab606a554a557885a007f83812c30b258c304a980220a99eaaa95
z5ca0326fa23e77906a8283026e7dd45a9ccdb962d40898c42f6763ba329cfe48428f7d7b2b3600
z7d815b60be3daa892e13b1b02d4b41839e0343db09a77c2ce8cc41f511f2cb9e23c32cfc6ef662
z96ecf8dca757bb654b79670cc15de5bf32a46352a9326ef9324bcee743592cd73d2af049f7024e
z4cde4fbfb62fa13077442ee1958fc61f34054f532714b644f0aa5c8802febeae4f9a3da3416af9
z6f268534c2cfdb85fd9988a4eadb074e57c3d3d80ce9b9abf9d550dd3f6ea690478525958f5f14
ze3bc57872bff30227355c5a37149ebf002f5722b3846ed4ead089d53b7aac83e8b648377e06385
zc38a619f67d0aec6df895381a6eb67d7cffca73b4409d9a08d774d4d3c1010b8d54592eb8edf68
z280ff6a8747d00c7e82f66c1dff2b2fd4babb78455613cdda88fb074bad1e0320339145dffeb18
z50e3aae4ab979657b1572523ec504ec8e848fc801b06b666b355b57bf4191c9963c49c0ab3e87d
zb27c3fbf5c3efb883e099dee252eb13807f502c170c468ee504d3b31f728831c3ccc0bd179d17e
z7dead1f248f9a0eac904f838edcd05f7c6bcdf7e7cfb92ca660795e18b7907c71a9328af6a29e2
z057545c1864b911b69ab3f7fe93377ba14f1700b6c91b81954cdb51b4bbca9f86081414f6e1456
z23739c89498a0994334e4787ceb2391effa072d74277a8374680bec35610b1012ac04584568fa7
z26db6f18ecbdc5ae3b5ef5214cfc0fcb2801fc11015fd72dd4dfc7101c662c2ba044890e548d7b
z7e4ed4cb3feabd8dce8c461fabbada6326ed91981a8a16da8de3bc7f5ec1b3f1d03f14a0291334
z9baccad9900817f9b1ca14239364f8d27d56c3589750adb5b5e9b35eb53855a3b328a6ccd4dfbc
z213bcf26ce41c9b29056971bcab93b1616df996ec8452a50b3bd05035eeed6f1c2fffec05a1788
z47c30530eb6475683a88091cd3b19a9f17c4597afaaa8fd47b89399bf42db94e2d7238ea42290d
z9a7ade6ea93d87288819a55839e2585e265971a04d00092408f7638505a2f7ba2b4427a831c137
z3b4884ff0845c632171d5f1db53ccbedc7b5994a629bc0fa9b9440900324bd937220c3e9ba3665
z2f1401410b2a9e513a76d439b12a3f12249f69bea83698882663bfaabbdff405016ff2ec5a9be5
z93dd8d1f2e6b41acd11538e0e2ddb046f3f823ee8b7e2228b0e5deef971987b33d6cd1dcd3a5b9
z22751a4e114058e661c5bc46c58cb46ea63ca2f266d64ebf71bafe2d055b09e67789c8c3bc262f
z1fd19f4a768668a3f1d55c1dc10975753be236aa719af968b9e322cee89d2b5d18296d350704f8
z1f33f68d26323e0bd1acba4164203d330231f9d642d3e2bf327452393fb547b7bde0634d03251b
z90326a1e8cd5e68446f368d948f82ebb836ff6217c9df1197b2f3e934aa1776e1a33ad4f16a525
zca752882407ff36690f06d02998939d2711ef45ebf5529f2679f6912a7bde6aab2f4f11ca4d643
zd6cafdf5824bd016323c0b34328dc88e8124f44cf5575107a9f01960e0ee80ef2c1bd1ff3ff36d
zc3258074e4c6f90988e7ff57e08b94f7d6cc956da4dfd6d6cffdc3f7d455eb89aca264c48d8834
z1ff66f0a00774f51bcb670e7eda41d9ee0f588c2c3ac5d3302a0026fdf636c7e6ce819faf3aa73
z909a4c656fec2993b63bd60942cf87b5809f972d3359481a7a61e45e45be2038a3889fe3c8c02b
zdae972c4ce7c081c4d7e8b9d19a7e3d4bac831d5dc9a0fb4464cd50b769be9d28c12b2b48f2b2f
z9ec3f5a48b8d79a72d4b522a34c78d0ba9b3f732218f3cecbb88e098777859ed625cd612441616
z36b6156607c2c95f5ac33f463b172a0faffb46c4965a5d733af523518273138d7c7ef9bd0f7aae
zcf25faf4f51b44c30bbf3537f5be76d2abc72118ce24a2846a2e1539964e4e8881a50ccdb0ac3b
zb6d5b9ab0d424d1b0d70400fcf0db0be3f45eddfc409ae2f4a1689a147fe9b287d5d3e27ffcaff
z85e8021f048d032ae39c6e358a2453c5f27561dc6fc31cecf1c7648be766163a9c077d04ed115d
zafebb289f8d437073293a8ed93e3a1ba54b43b5f4e4c6755ea3f7b14ce4f005926320c9c9f70da
zc03280b5ff8ffb9d42e845d33090f63cd7d082126c4d96432dbd59d0a95828798f59f8a3ab46cd
z1e5978c8ad9fc7251250f7e08feb61a4dd7112fa33fa0dca19b91f787482ba233ae34fba1488fe
z84303a172ae67ea075e81ef1b6dbd57719507195273cc11694744f1b5cf889feebf9c822ff1b02
z69639cc90a45793f21aede5b23a66d18760bc001ee8cb01a74e29f6e8a4b5cff1af8533da64f36
zd72e1110439eef09c318977325d5877d917c7ac1b33990d20197a04711b8e0924aa3426aebbf3d
zf5cfb584580c3bb63e47033b982dc2ef5bb27cda17f8d6bd302c1f160ad192ac17e265e071b7c8
zfd66ca1e0d9f7a8a787c4804545e6248dbdacc6bf89b1ce6cd5837132f726e408208490473f2ad
ze154c6b09d4dd03aa0a870e4a85019435e77ce9407df4b7f404eba195766b214962118916b9103
z1bb18dcc6cd9ee571d5bdad4b5022c46c263a9d72b729e092405174de0193f14455c719ddaf277
zd5334cd34fcf55e632a7c3cc2d9f45b0d55c72edee43ea0c8d00d9b762fbf85bbe5d99fb212257
zfc5b301f29f0fdb27c9b24537aab6805125ce0ac49064d3ac7b7295be8e5e4bf457902f363a34d
zec82c994ed5ace0ce3c6d37bd5b9d7adbc0aec94bc801336132a50e9a2b3ed87899212c1eedec9
z1ab090acae3de5d6667f289408f45cf800fe20af6e08ad81e9ea8ea443b31ddf859bb26e49fff4
z1ff77ad15e9e335611f339a3635a549cdf492cd0c6a97e7e60e1927b22aa1de9f34abeb3ca3fd6
z8c22b8894c4cee50fed8cf446372b9b325780d12d5dea0258023588b3fe941fb85bba7fe5f7ab9
z1f1ed9d1bc2ca4d12c7371dd2b54156a4adb67caab0094d0a325623077d21df1bfae4bbd74422b
zb7db028c0065447c6bcfc0c9c4dabcade3a85b2cbce8b7ecc4ad047786a7faba31b41ee107a39e
zdd1e078452535fcd2f9ff9003f8cb675e1c3280e93817e56ab675e58de1d89618a9c1d8c7c6e2d
zdfc4d3a6b744496d240b061b612575c2d7fd915516822c5ebb8340b5b01ec29f0898c8824b274f
z9ce4fa703c218808015ad529e791f6a1ddb36ee4f2e46e5caf60e7266ab00bcbb870f812ee17d8
zd04b90ed46052f06918438b6d1b9a97f1bc683d26564b65dc6f852a87604cdf387ee5a36ef552b
z24ca799d323bd1b4f025853d015a054781564d889597a68ebebdd67bedbc139328674f03c6b046
zb2dce191c3304e8b0037dd80ee9f56f52440354d645ff25dae24683f32d301fd5e03cb1c4a228f
z3efd205d8a92a3cf377043337b7d8cae580dfc3fbdab4bc5a1726a01e803ce76bf4a9d83ae29e5
z53d90d50a00fe9d2f1c3834e7dcabd63c629f307ee3acd66e618bcd562d806fc22dc94b112650e
z84c9f26c87c1fb56052398ed6fa893ba98087b2896a31ce806d998d7a07d9c0a7cc7fe5128654f
z52031da49c6e84399aa00a9703494a51828079dd7148a6c0e013407b0405e96dc1ff13879cfe6f
z7930238c61011ca34905b44d939284cb8a17a6cbe2f7e6144fd00d4ac5eae3545d595ac8942a54
zb3d6be6ce2e8f249ff278cf597847ab39ab1f4d23cb8d5dc71e1c24e7ffa163b13884d7f6a0f21
z72426c1cb7ab958eb4e0e4aff5a36f549630564415570c2277f6da49c956eb1d512984ca233788
zf545b32217fe7861a7299812b42457756445ffebdbc81485bcac3444c6473d6e186e620d57704b
z8f4c697edc4b19a707c63bb21996bb05a99bde4a10dae463688400207f9f7c0238443ac4e91d88
z4d5d8aeb5938462554612e2fee938069e781664ed835a815a3bed072c192de54435c20ef60c43d
zd724780eff8af6a55eb1bf9d47369dce0fdfccdcac6b12d27db2593ae557fd6f06fc9db814b067
za3bcdc6d464e7fd7b7011581f54321363edfd84f7fa130ae48bd28f252db7f98c93291c647feb9
z253d12ebefd5bd956cc2bad79583ca78fac0e36365958505c4e82bf246af3e5585c3a3d4cfac6d
zb03bcdaa51100433ba3588491492df6f5faa44447cf6d0066b142f43c3d9af5f54c1de0df14800
z62679fa48698760ce379f70f01aadc3a7bbd2bdeb25bc0deb49816601f3fc3998499c10aa812fb
zdc7bc4cc9d25077ed2650295f54aea4563de6b21ebb5041d5d2cd888d5b37488827fe6e477c9f4
z754519424dbd5a93627b613bf1d62d565fcf1ffc6ccb012e942871354f5b6c9875d5835535d2b0
zf32968e1412967deccf1a37402e415d58a5d78421f7086b02fdf0c262dac125401c032f21874ee
zab58606abb6c8195441026fef7c6c445d6b675d56963fd9ec3f5c66cf3234b02134dbf43e7c3c9
z7af9553c9956e98ebfe593bac3ec3eda7b90a3dcc462bba050174a4da7614a35a4d0b8f566c497
z9f94a1112525e275620284e8f72ee620929f8ebeaebe367cd2833b3059e5f0d6d97663205dc08e
z642cc3a2096bbee9575414dcf84a60a137fead6ee506de803bf6efcb4d4c307a36ce93f17fe832
z93a96439c38168ae5dbe7980018a63c1ea061ad1948b82e9890abb73b5a846aca0a3d7c213551f
z29cb9f7127dac3dfd48a0a6df0b9cfd6d0d24d63ac0defa33203b4f8b1f71bd48ea34c2c163f82
zbdde5d083e62f2e8fad9e1f5b291b8dbd20a8bd064899da3d8d2215475214b39ce839429109bb1
z1d91f71f7204a42ef641992acf09077944ade48c5f77f93a33e4868ff3d83070c1e02a29d027e0
z7b0362389173219d7973141283d54b0b208990ca69640242393e0ff1828b230f9093e6150c7f9f
zca95d03019f4a846f0a36014c17359134f852bb8a8d02dba649b62f66467f1fbeb27d021e924c7
z8463b8d05b7578246d614af1ec84ffb6593b312d1a3e6fe53164959244fd872de5c107c6639759
zeec5191589b2ac5225632dfdc3aa7e4bdfca869caa398e44980603d92d77d843578749f5349a59
z4839f903feb8b21b54b558ab1cfe2468a009477e665113413fd25c9ac939630333f898c6362073
z1acca23ad4f6228f39fec82c2f6d7c2c13cf63f1f2156614f806a3a942dc273c87940698efb943
z621c992f3303fd317bcb26e50b6380e5d653947f7c5967a4d4015a87ae3e90f3effb5f923fe563
zcd717ba85c67e75deb2614ddf89ddc6729bfa50cd6d93f84ac8891bc62ef1a17d12f5963c0d14f
z0949c6785aed90ce0e5f9ffcd83e8f2414d02f71f3c9409e82fc6a5efa1439083aea40c394dfd0
zf2e841daaff969b3bae6752bbfb3f5d0810c099d285b1865d4b81199b70f307c4c0072ca2071a0
za63ae9205cf914f6ca08240d739062fbc5788e888f0487c52fa9d2462c374c86a35f42b2dbb108
z2279e93bad10e9bebf360516b8c56900b5a1bd1ebee5f19c73a4db18b08697d064cd74be54014f
z875377bcc57a071ded9e70eb3795fadc538f7fdebcc36ed1e6e5455a000f584a254b54cfd0e2a0
z1ed6e8605d925e703757ce873232c20b046c5381f58a24ba29dce70bbfee5c8a1a5fb2355a8d64
zd0b3a47b07197ced84f7315bded401bdfee06911c4d116b70d34897250640785d98dac8e9d6fc5
zd2a38cd2940e5dccb513e4b0831b4dd22771b4105fef4e9db82a294b2acc5379311ba96c6390d0
za321b382dfc640720912e8edd0a146bb77d495735f87253ca40f27069684c6b42fa6def51ec6bf
z0591ab4b37692460dc4af7358f48d394e78e32b64bbb3711dd735a2e3fd2573f83bb5e4b49642f
z53ae08f2a0b49a2cc0ddb9fb1b591870fcf9369ee4ec5670c04988e5016d365ebb08ac7e3a74c4
z62d94fa4b368c73aaea35528b4a09eabd081c038036b22c0b2c6555ec2c0023ecae28ab9e7de4b
z70a5a627222172607ebf3c7ba4d87cd11a65fa3b90073e2916da6b2b49b3ca26accbbd038569f2
z08486713aeba2a4f714778efc8f760d7862737db42d14ea3a55622779f9b74fd7cce7ea44d377f
z6915ee1348cc210a49413b05b83b9baca7ae5cde7092ad2b97ecbe161dddb0004c3bf1be60cee5
z348a96acc0f19b664c19fddfdec9e78edfc150dfb5e82663b58655937838dd07b40c014bd053e9
zfadc0e4939afd72aab12ef1d4be45e7ac39946a298bcefa9502cb76ff6ab0d19a7fa538c6164d3
z39dad84b61f7b81e891b26408ee44d1ad31d9069796f73e2766eec112a284a2d45622dc1b97b18
z61c8223f31d766f7e184747e13e9e2eba20e0a3bf6dc0e43f2bfb12d9172361871392251382469
z3c245407e3afc2acf5ce7c1501d505ee0fbfdf7027d821864cc9a7d331a79897a004428dca7cb9
z8f024052121659171a31a72a5b581abf0b041a12f0092787dcd7247eea84f80d81e369488d4d5d
zfa59be83f8dc89355a5fb7bfdf455b2fe3fddf8c28bc1d901fa5ce1dcef873981dbd76708e389d
zf64a6f01edf6a724d3f32fdd1ba041d829f2c545562a2c9c4214c382c132452334ab8eaf7244ac
zdd2e00446c5298696d67b5a0a275d923c58b00eeb193d45f59b414bc4a11298b2d4a511538613f
z1f4ad7af4c8b2994a3d1eb8a53949c0efc400401e84aae30d5085d110e6869899bda107d6270c7
z0e0569f96608181bf75d0e89fea3c4b8bf337044bca0d2bac2ee3ab0f2dbd7d86861e2c17fd590
z7d32b6825b25875d7fce915195b8880eb50ed18ec987b54bf09c8bff4ff98e5848cf8d7e753f29
z19c9bc73bfcbe63b35e6238162dbed809806ab4e4b0b5245a22f6c6dbc7bb64cb93298602c445b
za322ab97eb56e6272b60d8bb56103ffeb1eac328264a78ee6e1896a1837851cd7e058f79d541b6
z9e32f991a6746f038674e5fff2e2fc6148880403ea3d41d0f3f5082c8cbeda3ab686d1f5948cab
zf933985ae85f00690166487b3575b3d1cb1b608eabcd40afc3c0bc73ef59982dda392ee1855402
zac1cc92c07b05ee9834404a71b438d69d76032f5e040a46c52883a2fd03e3a9ef0a9e4bf98ab16
z29dd926726b7255721ed93e9a8aa13acbe601abebf4f316c550ca21214ff992328fc44df1b8fd5
z7b0cc3f2ba3f1b8954907e17db45e16fc2fb0b81e828bbadf1d16bf7e08f9dc1bcc46f9ab5d6eb
z5ec8afd7d18f6d142b9e04fdb3dc39515e8b7a0e43242d8a6f72c3586f71fd4bc550ce3eb7abaf
z3428f74c0a31f646b4f1c6581d9979ff5ebc311394046678ed2954242a9b2912800704bef50072
z5f0766e6c7e702dfb946662c87306019539c616dbc2c6917ca243e7ea6d46290b5e408150ea25f
zd1a49f13d5d97dd7295ff2e80db3a5d8f1e9442b9c560c3757a5ae6f6972654506f3b7ee3276c2
z1b894f139ebddbc8d9550ae95828d65f720423f718e91df223b7765ba1831e3e8ac6adf877f150
z80960e026bcd09d26c34d3d43d2ff6b8495c67107f84305b97ef32572c05d0e88e4cc13d12258c
zfaa7575745e21d608f120c448c7664db7cf71758b86ea5181a92c7825dbfd4f418de6c2e30d745
zfb64f45c0b2a010872fce58c544f90ea68b6470225c520b8ba6ea3a061542beb3449439e30c6e2
z0367e5df4faccf134ee6958663794ac28d6b692da003bedc8eb151d577cbe5b05f0ce4fa66703b
z5706f7d85bf47594cbd667e9a346082f16114bc47ff5f9ea86a935fe6153ea33b7d2ef9665889f
zd970a5cd6c43bb614e6ca09cdc676d6af2b6b739c9d906a6aecdcbbe43575d7ac06f36c416b81b
z8e52d6fa0801c1e5dd0cc460b960e2438c99e70f2fd24e2460dd8314794faeada49dbf33936572
z9092dd11d2214d74e4ca18fbb32a3af6141a1b0add38f5c123d20b4a45d9e3411d0e5a956a9619
zf3ebebd2d2d2199d85428277ede6f9cddefb88e55e6df1f238fa90dd52e3285e65bb32ecf0e58d
z9415420d89a7f661c673cd80fb6ca9e50b5738d6516bc2cf348ffcccacbf5528e88f7d7db5e7af
zd0150e6bc110d8b33e3666bc144d0cb833debb09c697e845a122144ff3c58bafaf55c3680f163f
z796ecc6935821a3fc79e004e6f014e2e8266d0d024fbf26aee5de090623d478cb163ac12410b18
z75c938d3d535c91a52ebb5ee5c69a6706abf89c59d4120af02e3a5a66d1bbd1dbdfef92d500ae9
zc1daced4ef01c15ef2a609938ac0292d2b846027eeb98a8c2a10f41b4d96b558dd2f4d6f917189
z170f09eddc9d26c89699d3a1a320aa4ccb47164b1035d9e98001797b8f195c93878e9fb4a6e8fc
z27627037eabaac02177b28d8e86c5198f9808d0d1f990db568f2ee0cd5f4059853c89d85720e48
zb2b0d04291d66349418de83aa5575ed48b2d99eb76af86c466622bfe5808b6d2b991cdc7e0e97e
z751688c36c59ae5bb1180a256537ab16b825bd89d992c4b1e2ae87242378412e6cb86742dd4513
zfceaf9758c6670ecc22ca73dcb7c51a4767427eb41138083b27d8367927f53febf97aefe70e4f4
zb086e9ce6a9bc41fe917d61bf6201420bcc15530cc5c58df0ca4b87d050b22e34d7a214061ca5b
za669d28685e21f3720ca17d2e57e81253f4f94b0a2fa0cab045531e6cfc527e480e5819495de81
z0201cdfb6f45c788936a2acbb62894e9a06100a8693e6e41ca0a5bb5266e852a99f6eb91e7a06a
z5f6fbb9269f80e60aebe242fd392bb6cef7b8956d21479a16943f76dc2f5a54c9f6c911364a71f
z4e8df9f6b915178da6af4abe7bd76f83c06f9a01e2070864ddbb53d610fdccbf2f949c183964a2
z8d44237e3f823d1dd890368d81ef7721c9221175b3bd057e2232666116cd8881c3168759bb477a
z0e3f67600fcf6113e99af46cb63afa7bf32c2ea9838b231e11f17610fe554adf4e1dd4b2e27d40
z8ea57593f43311ff2dc5e64df891aacb2a37e01ae4833842eb508d8dc0455d153429a55f7c7676
zaf54fc51c1c2fcafc4e7475e33793b60c0532d71aa0ebef80a17d067e8258060c339c5579d52f3
z70c263411d25ff98e10db74a69843e5992207d6b17e9bb1832d3b32080f70a19c918ba1da1bd35
z985bdb7796306c2fb139f55ee6c52a6101ecbd1c6539c575797ae8e07db92918120309ac078f80
z5a27b10a5074d610ed05b744fde1ec9486b7ea998f7f8b8473dcd5c9cfe5dd2ec162e0081d69f0
z0c262dc9909bb035acb7ef02608bd98d6c5e7d0b61d0c4550b9d4481cd2b233257a984143e06ab
zc508189b737bb75909d806eed58aa3d5249d46addf40c2773567bd969d8e50b646e3f82c4146ef
z8ca504012f03344b5c48b5390c0039bd86509043cd463389ccd9631656979cec5c2170b05022cd
zd13aca1830e4b5291d0ff3a2f9f38d847feb4fc47b4ec68c5261d26f5b4fe894e274a1067fbcbc
z2e269513262989da9a0d23a35fc3c5096549afbffdfdd3a644ad8d472e4d676c0f5d3dd7430cc8
zf0cb261184b44b2c4221f8b3b31e7d267f2015c6f281183b8dd0d0d733d571187ddb2cc1c3946e
z88f38fc31cbef8eec1e45f5695f6508bfd42cd6a40588228621b1060a54d950228faa5b51ea920
z5321077d0f75edd034cd83b5084a229b670c6815ede371181063105ff3a422d334d3e1019f1aba
zb24ed56c494a0ac276ea2d7f2dc0faf3bfc9c330631faea3c5f3fbe2395728f02db72dcc593323
zba31e73b4a5b7d90faff544bdb58e4fd428bcfc3d86112efa4a3b94a6527dee330e39195079e94
z3ad640ec8dcee1593ff3644495c11b9f09e4757945d35e32ab3c1d83f22c0770adbf91e8be8e5d
z83be23ccfaa6d4441906711eb3f952dff48927cb427231c58de5c3867215ac1d6149f9123aa840
z58f9a79c88ce30b8840b51855ac98443b18a237b926c7499951f40e632569087589f1991d5b18c
zee1fe170acb3d3b47725737cd336554dece02e1bd5bf206cbe65a56ac7cedfbeb7d6a23d37b006
z58a739a0c76c6774ee07889092b194c5cebb49b04a80f04d9964fe56261bbc6555524a432c3970
z2f59a550f91a73dc80e61ad6e23caf87b0b1c9be5ca3b800351c17895d7053b5b1540b7f88b91f
z15304042a8105e2358a8148d5c8a4bf9813e933a2d82255ba88b4a861fc077337a70ca818dd932
z0c7047063f6170da0332757541d5b7d3cc9d334bd7f7f39937fe53550a74f748f4561732af5573
z7bdd97d3827a1c163cc33085b9ccf26b57020d467d3a106e1e3c0add33f832fdd9a07f118b21e4
zb675d0ec41e2372abba55e07667e8c52756bd6366dee4c5bb1c999ca70808c31e7697f48eda92c
z45db63a651b5974ee5a12ec362fd761951eb3036d27858acfb5d40a31cb060c3159911ae690ce9
z1837641d9c5de171c6dbbbf36618bef7738610c707c4964bb577245c2abd68580e2f4b75c22454
zcabcdecedac4f1b574976dc8d46f543a1f2171dc59129cb865932c5bf02fca811c9a994acdfcfa
z78c45aedc2b31f8180ab23efe1baef82c204e678b2bbe897f5f1da064bdfd72dadfb5fae57e88b
z7345774f68e8bc89faabaa8a39b953cbb7dea2a15bbd9ba403e464b9789f4fd70437eed58b90ef
z5fe31586a9f279da24cc55d6ab841ca77b197e6eabcb895a9e38d3f0eb2264dcd56141a573be57
za4259f214901118b5ed9a8ca4cd7f5a705ca90689f2ac7d84f9035adfd8a31a87ae8d0aa8ae980
za1a333286a0ea4e9c02a3aae1300d147983439c6dc77b1d972351a8fd0b6802845f24065e5b5b3
zffb7e8575349b171858ab00ef3ae15014f8af5d66776ee028347823cd220755c26dfcb77f1f0e9
za1f52b7b289292e82a1975a1c7f0c87f12db4e42ceb082f248f10c20c4df305748d464c0308749
z015f3f3c669b14c40df3ddb3ab7523d0a246a996f31667f231ab56203badfbaa42015c551ce4b6
z3c7418feaac45f235fb11fa7bcd8f8d5b563a6326a2619230c10008289e6dd2a91137a138cf67a
z46db0d78ac2740f8c1297bcd174dbb0015b1e0ac43279b4b15f8997f29ca916ca5a08756296d97
z80d77b0d24a4d905caed6b6ef9e5bbf08d828bfc15b69db62b83dba0706d510c1e6965dc8d1ca7
z5dbb471440818d2e4652438a1a4e407d2a763e9ea15edd1a9fa941e880fb9749a5da0c9cfdf4d5
z2908645188f315351373e40b02f941c1c826fbcf2b5bcdad48bfc45cec9c84249e80b923b0ff0a
z02c1b64463deb2945b9abd5cf76e04a4367d278fc752d77270bb6a79d10bdfef4aaeda025f0b48
zc39db6f8d2533b84e9200086319c32a1798756fc6f150ec04d477b86442cbc6c5fd70d6db01173
z3090d6ae937084cea61f148c626c5d797e0f83069af2b3a71a2c617fb32a9362854cf82b200228
zc28e99f8b93048c83fc86175e2a55274fb3d855e0bcfd8446963d7e8fee154ed9ea39a6a272679
z8cb25f5036cb5fe8e260c29804345d9af6f0605581b86e5d7295756a9012b9df00214d8f05c576
z2316b28f0d8dca84aeb7f5a86c970ec697d77fbebdb1d815b7234b96aef0c5ef5cc7e81a59c0bf
z5717009eaf92a95ee544dc6d53df27ccae8d899725d185d11649e745936eff6626934e4c90b5f2
zee66d64327631c3f1eb148aa79d99b5d8824a9a28910b696ec31280c16a8adde6cbcaaf154e6c5
zcf34197bca9a0e759e84988473afd0514eab328631a9eeeeee8915c5ba5b61f3cda2e18f537f9d
zbe9c439a5cae59b974c9dbc59cb493820b182fe5810473cb247bbeb95a21218786371c6be410ea
z44156a31f5226fbce83997174d26bd586aeabe90401f199546b3e0e165837254fe6142f50a5e12
z59f8ad9f52710e5438f0d818b44255629c5044fbe596ce88e01d4966ec34f86042d59a7e54f279
z005152711662c66a2a2bad5bb4dffe3af1af58428f1c843d7a2a257de097acb6a2322b9e88ffbd
zc4f1729b9dcd8b3c732e305ce55af528c1e1b59fbc11db00f91b85fc3a39be76e33317aed5724b
z6c1fb9d2c2679824b4277d8bf93808beebb9b26b51bb113f20c2d87eeee6905b10b3476fe51ad5
z485313566c279fbca32e9ed05b4690c2e38843d5435305b7ee72196ec972436cfd1edea563e717
z02951095c9d971836effe3bdaf63a1a430259640e2dda15f4ec4886a78faab83d93d43a9b6a35f
z07680b55a2426e26dc25f42cf35c08d6a7e8293bc396c1df769f2fd9bad1f67950c6851d77e6f1
zbb1029e7e5700d25a4bc193e792289f6de418cdb001b643b5ac2aebc21d2a82d35c8f4a4b2e7b6
zf0797df1b70d747ad3b4b01a67b8b9fb9637cb17883a9983f9188975a80d35144f83e6357039ac
z56e0983b1085ad7867a4f7126231f611ce60b211af1d3ebd8ab161f83211ac3ba879bab9b1c7b7
zfb6c3f21cb2aac26
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_ddr2_sdram_2_0_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
