`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc7eafbde2
z54611f4ed90e5bddc938938c26736aa53e9689fbf9636fb31847053cd2bbfd5d3d217ab8dc7416
zf8a3ec85dfb34ad227cf64f935216be2a9e692d6fd7940078b873ae6abcc2057bd462565b5c127
zbf19c4447dbcaa08e647cafca73985887dfe942976e77a52d1dc32981585ec480431362c0621ba
z170228dda8222f04c788e3de6c5cb957815f0aacec766dce2e4363879f993680e07d822ce4320d
z5a53a923799c12ed3e609c8147dc3555dfcb353c14032fd72e591b32ef0de2aee4197886b84b3e
zeb6f7b226c0d758d41107b6ca2d2acf6140101fe2b848a54ddb819025d501319a0cbe43aeb0371
zfe755e586eca62eb785ae1505fbe7c3c16216f7dd4f22e55d87c361fdc018881bdcfb3a5c43b05
z980794233bfcf56dc1b7ce9190fadb854a58588a9ea63b761ce9bbf66f1bfef74806d029dd41a1
ze67779207bd6deb6c398c088e1a0c2bffb11e6a77421e6a2ab6255370c41745b28ec54b7194e61
z54c486c7069b85d45dc5f6ebc1a1e44e9f98d81415f29bfa36554c4c24cd1167d7981ff01d8aee
z46bbf43b6ea0a28612c3d3f688cd97ebb1adb12d6474acd4de64ff7a7401dc1c05f034d64c5b8f
zc58714c2cc9ae8c2bcfdce4eabdf1a61a2213458f7554121967dec83585ce6624d498c39cd000c
z2c057c49433309d81415b0b54fa49357e3ed51089e76a1af25b0b86aaba51e404f4bdeb479edd5
z57d52e7b0a8643657d29feb5139557b7d9caf438f6309b36e6afdbd0070905d4c8fe16baaf7842
zdab1d795552624017cb57898520fec98cc04f2febf6c39aca82b3d9acaa9160c3b520519cd8dc6
z6c5bb639ca1db162bf42e50d6cebe5a8f9b7ae75c947f1ef552e0546a904a10e0f1d6c95fd71fc
zd2e27a1893a5ad5c9f593adfd925b90c9cf13aef2246dffbe4b575dccea929d4569a26b655e723
zc36672369f2846a716c543ce4dcb48aa3f988a8acd6bc430402b6647f02ca1401f86f772d75542
ze59ad2ac05286658d88124493f883de7f25731770ddc6a4276809d86e3a9545b3914ed0131e2ad
zcc759bc74527812ae3c0d0e4f0dd1603817c8abf1f9f3de62d864f9ca864dbc067d71faa44bac6
zf0aa658eeb1739531540dca11b003e76a575de9474cdbbdcf1ba81560beaa73aeef37298f26e60
zeccc0f9085a207bacf2d1f72495425bc5ed5d67800272b229684fbb56c8b8a0a247d4c0f12041c
z77e9e1737b3006e3642f4b1728c9ac3da0dcb223c93e0b9cea699db1f911b4b126ba452eb33ac4
zc78d0e2dd17377f7b448ac63fd17f361f2e9115f831c9571134aabdb8d20b0333dd19b41220a4b
z8530022b2762b6b15c088c6bdfb29bc6d147a474e03b1a923f8441c0289a2e0bf9bbb87b38a51f
zae1c7a440044a92cad681f4b19d77bde24627c2dc6a668d63dd00b5c9b6273ccb6210fa06d635e
zf0271a06f314aacf0e209bf9e9a29fab3bfd7c9be0774f99465f333d5071f4c095d08ec963b48f
z37735a9f40a2541c0dea42e75f81d2595e14adb1a3cc9b4dc70e4c0c448e3bcd8c9e1e2be7dfd4
zc24eae2ace926c1fdad78b218b6eed28a932b66fb52b3318e5f1249b90adde7f44c1607a5f803d
zddfa89f2610fece170bef5cf24ee3e2d84d688a1faf64877abd78406955d55cd1dcc8f877c9f4f
z9266cc3c2e757fdf84100cd8026b4a0b1ab5f4a9a9a415afc4011e3b9b33be844dbc63d9241fff
z25576fecde9e8d96f40173294c90ea8ab47dbe984178dc5c50d14abbfe6c08b84a716f45e3a0a5
z463b9d70c71d9110c8aedae582175ea5cee579512f6ed0daef8bd2c060a5cd9f53e0186b741c77
zd6ccdfc206cf33ddf06f6fcbfcd349d597c6444354569d098546fa6c22f1b20749ca740ba03ed9
z873977e1f456e9055fdf99043b650b1d841519c9fb1cdd3c87e80129826db0cd8d786d0c33275c
z9c6902284c059e1df271d633096cf2ef8527ba913af7f67d36ff108869d5e7bf6f09fb543aace9
z2402e20f8d1231058674319312d140b35a5737091649b7a9bb139e27cdc9833c97ecd9a6e0522a
z284135ef45dc76fbbdd93e9ba5f169a0dd38730f5f42ffe723a34c5b77c3de14f9f7729b7d6bf9
z8c1d5261a1dd8d9930ad7f47f5bb5f90965a731c3d9126e989e92bb919843fb4317eb9ff0ddd59
z2c86647a96ae26759ce1a661a19dd917fdc76406eff01beb686d5d07d339dc18b2bd7fd63c873e
zfcdbc8362686389e91fef85402698182e73f916aaf160a08618aa8c1c6b5e92c36d68c7cb0bb02
ze83a7b765ee84ef2f68df41cd7c5ab72775db3014bd89ecaa9ca3afc04a8252e981e170d99720d
z03486b863eb9521ec03fedbd562800fa0b6e1a5bdad910a11f90a885913bd1fdee94e9b4dacbee
z14236c1868729d8f502540a79b3d1c0ffaa1e1f7aad82bdc0c02ce92900d2b0cb576812424af73
z589bdc487519df7f061ec79a3f64fc65d650873b7b6ad24c37e57411381287faf330a6bbd9fb88
z7932b4ec6307b24f3a0d69b05b87ac835733ef6eae4899ba717664a5d52e6d0f4ab5959b8a6adb
ze8605360076074b36c92c2dd882201fcb77a9d14978e871680a752278fc531d7e1e18be5bb14b0
z560bae5307fbefd372187e87b44ddf8d412f6f99ce39d131376332162be7ec2094a44987c52f2b
zc9a8162a175cd5472a4b9235073b39a5659bd551df3435d635daffdc29340426dbe4ba1c076b91
zabcccd2de649c5f838f0a960fadb7139d16186d200803b058bb5b6d267f263416aba62f0948dfc
z91695225fc774cb37f8fc57d3e6eba768660a382a57896bf82d0d629a76a421a309d7e05af96d5
z1e36fdfe85136d7f2e4be9de50b058bada9b2ee0a04aa1d181bf76d44e092be78ad241fc8d530f
z04a92721e21f2477f148c47b1ce99cbd6030d771dfd2630304e93178a55a4e8a63b3e1468187db
z19caaab18c53e89926324be5f5bc99630c3d347149c3db3f9a553249f32f72f725a9b4be088c2d
zb843932c14f8c65597e37a200bdd0cbed08f0309b355fcd749b974f6b8ada071df6252a7b2b1ce
z2f8445f91ed81f5423f857eea8d44aabfc616d7ba253f6f90e67b25e352327c53908ef46346a50
z9ea35e315a02c15e1af4a84a0e8b587b3d3a6351c77c55f70321723100de69d0dee0fe28ca9388
za2cde96ab56f70f505102eb54ea1410e76d672bd7184efb39bc08e1f671ecbae7f164ef3ba9991
zf50130bc6b67e8d115c843ff8964a8df7453a5dda80d29732b6448d32e2648ac9f31d38cda93eb
z2ea7ffa28912f05a79e325f7d89315852ea4b9fdebce07133b187b10ccc24b65086f593d0c493e
z5070bb513ee57ae3b1107f4be7fe2a8d9fefee3a6d58eed5bbf6a5db42eef161ab38e8ea7e7be2
zd4e3b2e4548b9826e846d83821e27bf775bbf2d5f47d40b157c34190535b9ba338879e41058aff
z04a0bf6e9bae40d145b8f0ac7282081d3da13094c124498aff2a97e466db832afc6fb14a396c96
z0d38f72579c38805ebd47d0321473376b6f41c2035c58c0688d0b314c4423a36e24cce39adf939
z42dc9a60f82308f2f567ecbfe1fb37f7e27abb6ff7f9624c5a5a1e263b153e380e76d46f73ba29
z340908c3a338e4bebc3627230ee09530b42eadafc7e58f9add03503bf820335af3bcbdbafdd3bd
z784cec7e855473f6fbca0dfc8d3c957ca02820f83dba09be125c6ce1266828e47a55fa1bf476d3
z9d5c64325ba0f192c60014546b7b284a852ca56a76ffe1fc40c6412610c6ef4603a29a81a065bd
zec62bdc545a9560321314605de47c572f7d4a2aca5d32e8f4599cabc2075c15a8365671f6fc2cc
z74484223b91188c28e85a215cdcd9c819ddb335272a1760c0142bb9215ed3ad2926451721fd69f
z37bf5c4723e3c346c58b5cec46be9a63889e0db6d7877e29a505b822efeaf601125022da1b0d36
z07cda2206bb536724c099f11ef12fe124a41d57e7dfb368f7b36090b500a4bfb87b09788252501
zc8cc74b79b1264e7cd5a91105fa92064b93281278d775a2c46aeab859de2f358618e0eb5a276ce
zc6a41df8d7e2c9ad5e58f8dfddeaa4c67e2edd3ee4cde8e3748105096702af68669597b96e4c42
z0fda13351199b1e353ffec5bede77b9ed7a66d6a7fb28f5b0debb419142a621ff3b6de91324165
za66fc4f1796a92caa584c5f25ce606d480ea78cd2001d2aef36e96c39b07fea49ca12d59430cf6
zc48b2c9444f8f0478ea0fdd974b87d28940a3d726710bdcc6a184446da21e9f54c6654f9cb5f08
z8b0f84381123e53536cb4d0c6bf2e93ff71bb1d020569147e5200fc6253fac0bc086d2d375919c
z13843d3d98e759db8cd3b095e942546e3811bf027f3c68f2835e57bb01adb7f52d3eea65387b18
z0bde95da0c2cd2bf6e2b8f07120b5aa2a1de7602c12ba9a99cc6f9c5a3394812e6099295317842
z8e4a977e15d77e1857edc68ec6ff2d1d923898c7df8f45cb2f05e2cf1db4e4669ef814a8205f2b
z718d388af347988501da603377f3f5733562cfe3708fd123b1deac96799bd8ccf8468c6f9ffc9f
z7ce849de782be9a99321b4afdf486f70c26362571c32d4841a270931d9326b3743d3b9bc44cc68
z31ac510b299bc70df18911580c709546043ce2206b959bb4eacaebfbbe8684dc1aac5506559d3b
zbbddd4dac44204d0a058eade3a9e15d6d5533c9df86868b7318ee31d41460c9a5af42e07d01cc5
z62b8a174648bda2be8846138ce6a688c04848a0d54768007d81e539023f3527fd84eb1ab4fa6de
ze20752341039401298085d2af567b557864dd797c8c13052a672423c4598d5ac8c5d2a5cc76987
zb8cdbda23c406cfad75c43e7c67918c3dd18152dd7675b62ad71439e24bfd8d940511796f5c9cc
zc72d02451efd683c14d7d6c8a21fc83720558a3804ecf62798d0db63d68ea453ceb1ff2f0e6d55
zca467b4dccc5a798499c83a030fbdd249b7d243f777f45f6e82aeeb86550f8c593556adb16eb89
z19289a82f8ca5ad50656d2b260ff38b763ce989bf47230ad7edb699545c08905d14f0ec74ba932
zd13751802213a61209f7e6cc2e20ff4bf692b1ddc38dc615f6204c483b68ab70fef564e7d90217
z4897c43c71fbcd6cfeedf535530d4f544ed73a25f3dbf28c53d22db2f0e9d5af8c03be88c9b2d8
z90c66614384c21fe8a71c8d994c618955b3d9d59012ceba8cc3d5426217c51f73fc358815e24b9
z5abddc15e72690edf7ecd94f144d9d7aa998e547b33e4070e92ae3f2f67491b9b77624f5ac349e
z99730c2810f90b5bbe2dce37c5b1704090d618f6121ccf40aaead18d5a2bf6beefdca3349f943f
z6c34f3fc91d580df99e25715dda6c1e7b11c46a4cbd28ea1cd4128496686c0ff144d1a32f19b8d
z89fc1a4bec03093371c4680007234f5baa92a07c9c8e1563f5d1fb4e8aae0476ea41869668f805
z70076ae00b9809704c5336f8042b1aa446daaf5f981392851ec087dfdff40aa94212c53c689c9a
z022a5e98643d9e92a9b4ecd308a87152ec8b3739120aae97ef78aabf2f32f16cca81ead65cf7a3
z538d0fe9264a55fb448c37604fc46b86059f706a1e255388692011f3b0fc3e5ccacf5d18a9f737
z460150af0dfed60dedc2af6146f2b86eee91511a2c3b7f6bb264e69f2fc1cd3aa5508b67e40644
z5213e058e7ed882db62c8f797af22685da2eea04c95d5242c04d6013a8f7dde72d08ceb6ddcabd
zc82dd0b17f84a19b879e5534e93fb2d7ac7c3f48c6e96597e3dd758f986bb84c6d5a31e892bf40
z5d18ee096e23df5e4d6fe2b30a39342538bf4bcae7923fa0896586d41676dbb48c08cdaf123d11
z7976492cbeef4416e03272eb4711556939557c86d16123ba19a8ed4bd2c9e7d41b161553d8c93f
z093c0d9399023b02e9f77289585623db17e5320e5040d8991b5ad2559262ac29d0a5e1ebf79a1a
z1829215bb3b454cfc25daa7f102af207c67a9607c083417442fb55f109cc2a622dc9bcfb116d7b
z0089f860cebd4d18960dd4f00bd1fcdda7fda485e17f82c11e56a183c109e71e4e1e3f158bff2f
zc954602945d691c99ca4752bf5cf2b05de0e95ab975a819a0b6e03f5a18a6517a1b35c89dd90b4
z4124c932057d5103505ef54eb408ac58ba578acabe499cd2811ff78e59f2b05f0c275f9fea3378
ze5047b04ba1dd6a5c94b267e1dc5581cf237948934a5c03fa875f674d1632e76a1810a58325225
z5a121599a5e392a653a1a4105c5f87c6ed380f8f4b3691f83de44e07cb68867ddf8dd711ca7522
zf9b0384baf0e14ae2d1fdf8298ce5d33a0c5750b6614cdc2cc7c8bc3de0576c72b5a6cca7db8f8
z492306086a717539db1d5161c585456d1a544546f4b86ad3b290a6b1987f1a655a0809496e9b3c
zcc3279826618d922cb088a8368fc5eae52505cecfb0651f3812b8d10fa87d84e127e3e31d4c40c
z630c32f693fdcf6b3e88079560c045b4773fb8b988ad397aeb87ae7a9547f41d965ddf41d5f781
z7897ad3a88d62cd39eef327621a9289df1dfb52ebe952dba63ce45978fb4a4464ff1b9f71db475
z8b9157ff25be2542d075445c3dcecb4a8db51b22f2733527967dc26e072974e5b59312e2a808af
z1b92cefc187e4ee4570536fbc1b59ef3a4a2d5b2312d169e83a74cb5e39c18b9ff3866f214ab52
zdd8c62574ab4713c07fbca2a6531fdedcfabb9245adb04f3ccc44878d4493438c01967cd60b345
zbb59d6087a134a70b17e8b958a1cc265162fbf0a848bb596e12cb8bc53f81d96dbc94d84ed2728
z245f577e00c8eee55aaf5aabc8426d3dcfa3a8bc19bc12c8f1c6c879c9c2c0f182b732c07ff3ac
z6286bbea4212b0d0942415b2ad87e49cecb2c98e84f8193b8f78d9c1398bbc423d7386e177549b
z31d7afb55757e6a1d5bf1dd14cf60a15cfb7e9aedd7d39a16528a86cac19aa564f3fc16be7eca8
z43f3d97fd36ceb47b11251345ab15806d50259c5434ae60b6e45c44bc802993ecd9f7aa48e783c
z6aa835eaaef24429460ddedfb512ef5708044ef75339ca6a7dd4dbc400d9ff294ad71eb98bd8b6
z771a0f34dfdfc7f794d7bb843bda69fef442d7ae685719182afb92393ccdcdd8acef9e45686ef6
zbd18ce14803a88e04dab8b6bb8f67ac29dc80e1a57725d37029bfc5f0b1bbe1944f98db27d887b
z21da9247a12f46976f42dce5915f12ccd773203d308229d9c59f098ba0366a067376289d465b8f
z93522dff7ed50ee6c5f6e1fe8f4a13c3862b7c448c47f408388236c9b24c3bbb3149199948fdc7
z2696d3c72b7350ef575de059ed3cfb06caba05db67426e415b1cf617305060753984dbdf461ca9
z05419d284a0d7b6300fcf4fd37d24beae4e600dd6772ff1d5b363b260f5d135c2b5ea6ee79b79e
z467086460665d5fbcbf8ebd4f4d3a6feffcfaad6a68f183ba659fe6aee586c4c9d11be5bd115ce
z585df0c07251573e748ebfb1ee332b9a5fbc1da5cf94463730a9ed07044c62df9cc66c0c7c9b31
zc4a0d2541971793b0b2b18c55679c664cdd39de28b6c42e5bb4694c50c2265b31d59f963bf17d9
z2cb69a69407d132a39a608512c5a01713219f3e8fb7fe897fc63f3accfec7281f06b3d5e01c180
z3c2d500cac842d1eaa6cad1bfbb850beba393b2c6c6f1b129b663246baa762156ee2285217540c
zfe5e56294e173e44d70a38d995eccfd6e790438c339036b16ce8a9bb60a749db332bb359a53d15
z0e11bbdf5dcfefc07f08b94794ae78e54a5dfa40e076b6b20665669914817354a00d82121e209e
zf874003b8d05fbf6107daa1856646a4358e4070dc725fa48d2cb9c5ca0234e5b3bdd81d9fb6112
zad3a7a8367187c6f83bf804a66bb81e2bc65ff558bc9327d391522f3fd923f08a7955333a45038
z3a3b27f788125054fba43e3cf7bd91ab985dd3a772949196f2791ec638d17841f8fc8b2ae56a75
zc415aa8dd825b3ea86eb02c1dc4d82de65fc7d5df78bd87eec88e1a10b58c451618d7e680c93c7
zffc8f8d92c69843150312dccfa7e40ce0f3c8ec473ccefa0444a8620d90874ca008596e55731b0
z6fc804ad20adf4d45df5324959b364251edf3d696e968e66a0218bf24cc2e6b2be0bf7b86e32d0
z8aec8cc8d22fc1198ef4320b90a220a2d18d86d14f1ec5a5f6ede79ff469f9b665df84aa5a2d13
zaab2a39e0815a3f7f29879be38165ee447cbbb65e651cd3c2b4920daf6b6d561f490090547e503
z35602e98d994df35a21236afd12ba5769bce4ccd25368565b0fcf2285301d576d0458c4631ffd0
z1f608f4fdb5cb4128cd006195a7a691325b65998afaf1352f1607704b7c490db8b0adbe2ea4a90
zd462a37b43caf8e6ce8ce06bf1269acca15d05e0355eb7ad90317f5f3e074c5e2a0e37b842d71b
z69ffb093564d85e1eda6eb2d652d4e1d522ba1a7cd3690604e6be3b5246a447d163f044eb0a568
zf20847aa36dbdcda81e66d725fef2fffe6d670ea00533874b523dda43d58dceb2e014b632c179b
ze2733a4a4828e61126a48b5f3c162a50b3e810af53e6f2cf20b9d33cadda1eb40aca47c8cb0333
z0b3cd28344cb2c85b554300403bdadcb99a47d19924f216729c835871b76a0ae3230b1a22b6ca2
z39a03977352cbe3c15f41644a9c2d67cfd35e6716dc1b99a3d45fc84d83b78156c7ed5e69637ef
z51993107394a947cfade09dabd4ece01a0ce6622e47fa760043705ec9db4f9503e0575eb45ee48
z2a5840b4ab3a4c0260570c7ae51e654d2c80837be1bbe36df2449aedb477184dfe21ff1f54478f
zc335e61ff546c8e1d77f3323a7d1e3a15e36d5631aaf34dd0233192d320aa0312fdd74beab1ffa
zfe2d20a0c3bffb9223b36cb8c5cc8ae7fec2ae338fd50ddffd70fe40dca7a4e0500d0739ea4199
z898a51f5fcb0888a31ff62fa0ce80fa79a4d480b38e16a1e0b227ce4953c320c25d1f5a571be66
zdefbfbcddac1196dfdf8ecd8916d948aaeab73ccaa5f243c6676477a68af998d3edb7f2fe839f2
ze0c2bcc040a812e3e38d5dccc4d1b63c85aaeab7087f6c82d61b8d50d27b3d9d2ad3d350eb8896
zdb52751ed1e5873ec4a25f3523cc454a39dae301e8fbbbeb0fdc25a7622ba578debd652b7899ff
z3f4e085ddf8784f6bbdad50a4a0380853cff3a8de08eb05e96beff270bad946b2e4f329dce2601
z3b583636f5e24a4ff69d358e83166a28a6ca15052192b4e807c65f286aae833b6eb78c3f213f9a
z6ef4d697a1d05e76990c2c0b439f880e17429e2b8aa3f475606e406adb92f7d735e4f9c5311941
z8003de45096cfac1b5b3417e9cbaa3e33f33a595d0bed9d05daa29bcbb891b429431021bab9f04
z0e4c9a4de49a677ac50da4dcf574cebec9ff1a334ce33752e962fdb9797d078b6f62a8b481cc17
zda260c57c52dabbc0eff30a77a45577bf2a17a4bc04a922f0d4e33087adc567a186a6a4f76d558
z19ec6dfadeab9beda5f89bd647defd2358cfc7a5e9daea29e80fe898a3993746e3cb3c60013eb7
z562d03c60650562e154de933a2ea218da4059f54d44b1a480994a4ae017a66e292e0fca62a1736
zbe5397712c2e7c9fa30e689de7093c2b327f39a630e0e1e2ae9f5219f00ac20799dc4d0e22029c
z7ef3eeb52aec3100b952dc6dd4471436a42a051184f2abcc71a149be8f536a6817dd48f12e7778
z44499bd23caf788f16cbf6440938b7efd15e4f7e3fc63a5f2b08577329c80eadf156a0f60e9462
z7c9793740685168555d0f0752fd0902838d04b221fa4ed567d0ea09a46d153146ba3dd674f9d9e
zc87d540832203739d3f0b96f20a4a92e8cb744cff4bdc9ed4398f3e8407b7a2a6fd59ccbf1e96a
z0705eca9c513f41e6c1f713a2a090f52a3f702c54aece4b0eddcab2bdb1999962172fcf209cd8c
zb7b00a6f36c6ab4f34c14a9d371d3791b2b113f9a78e0e4244bc8ed5c7712393347d52dc17b86e
z26cd9cee8d3218d2faf24e4a49c03bf3c644dfc6565978d242ea9f6bfc2fee77c87534a1824154
z25a389da4fd065a25480f5598c999e846031274c25b65e51f14f62ca66f5d3daf8436210cea09d
z1a010a9194bb2d06285e467701f49e8eabde1d63b322c40afa52d7aaf11095b68eaf2e983a418c
z90d5d77543d4f5e358243ae2e707a60a45c41f2ecf21ebc7bcb5e3d0eeededd634d4ea295f17fe
za3caca36f05aed0eb04e3d6c104a02c00f0ec121952e314b1326380f3922c5c0f76356d8de019e
z2aabd373848bbae8672490f5a045c72cbc05b2daf21ba5c06dbac3c4754dacf0a503aed735dc59
z42c4c12782ebe4a228aa8d557e7acd97778f9f6c528f67c389f62cee4b8716d187385805b2dd44
z24f50332caf2f61ded9656e5c2ed9f878a79f38ee7da51c925eebb3517dd804974f73a3dc2d507
za0005435a5cdb8b6d611a1c611e37d984d81677f1e9344fc3c9efe3c6f8912f47db0644bad7a0d
zc81628535c979707814097b134511077cda3cf54bed4b521e7a841b25b4df9c7493c6c018cd696
z8cbaccd43438b7b56a7049e72747d7eb5c648112d4addee86fbb057cdd2281333ab9d96ba098d8
z342a3683969826ed1a373024b47469a5e29dbd1d2475ea7d39d87fa44fc961e175577c7738a599
z07b8b25ba3df40d4da9a59e5283b0e1e1ae07a539b78860117f09645a2e2324d3d86a553ed3ede
za04e36fd07a7b25c84f298a614bb060abaf87d514440b5c6caa07363ad5dd36d0000c0be334f03
zd58e4b67f2d0b7e57938d908335083125240887419431a5c2d84badd376c6ccdd5aa06435e96a4
z09cbb0dabe2c62fb0f6e2e96dd407895b654d9d0ecf09bf58d0864427493f80733dd316876aa03
zd633eac3584fb1d59cab9c8f08e2838a879eb07e0e0974553af4304e2093dce6ee91b7e211ed3c
za9bc3f37ff3ede3d307b6200aa0345d29e9859b48dfa981fb82a60cb691d333b0269472646d616
z917aa0f6e814ebfc5e77a4aa4da5856fcc83f167586e20b8e8534cab09cb2c2b2346d81e20304b
z128ddb20bd8727287331216e4d4c1280068a65628d0debae0ca17a5889a49989be28be2dc967d8
z128e3522664c910b79852bb9fe08f3e333b46c3aec06bc684b2ed0b9f0bf26223aef763ca504bb
za2d58da56721195ed422340659a4236ab5ebfb0b92fd500a5c2c6684504f79642de58f1cb04e4a
z6bcce67b2cc42727ec2afd80d662e9d6dfa2ab9366fbca1821c8d65b28ff8f297c272c67369d7b
z0a03c06f4e84b4e456dfbeaceb6102c3c21c7f6b9f863f1b3378c5360851c3ec8aa3d076a4171b
z751ca72ff807b9ba3313237f01b010665358db5c2b5d09290f991db463a4e0f4269188c402a1e4
z83342b2bbd95250881f074a2e201f4aed9b944affebfc85a6b3eb23dcc73ae26eb7bbb37e67c7f
zc5278f725e78e7ea02ad74ee0160a24242c268f269d8c96e6b61ebdac850d2eecfbc8e864afb1f
zd34b1f67ce1a02d41a9a3cc4dc62c9386954a58c91b441ff0f5b96779e2449fc3f199e1b851440
z3a412734c8251f879d5f1c7bde34ca16d7db49ce15df6f7ed03cd11fa383a9e63942f01454e695
z73b67cca1e89cddf99dd252599c3b3edf2911c18445de5408941e8092560e75e6facd15961a048
z8803bbd2491113a572acf9278dda26eb2d8402c5c32174e4559c16e447e61490e784716a136a15
zf09e4d0cfbf3ec135890c0e8b41f250d1773e99a2ea492a4abd270978a9feed033dcd10d1652b1
z427e254fde82d323ac0c906328eb71afee66088814ca97b5b583011503ba642c5484b87147b241
z9df0449f919dafe5ae7547b8eb4fe4d39e8a8536f229b83f3c8503862334cbaefe6e79813bb514
z3e4e7482cd465703cf61c4e4ff7c71f9eb98450b6fc114b200b1a16ebfa1b25a0d15bb3126f47b
z2e97786c73da0692ed73799213b5720f7172669a1ddf513ea12ee74a959a9fda3568c8caaaa97c
z33f0c81d6e7ff74aba1859533361b5f6b8c6c7dc1d4d2e49416903e1bc930cef0954b28340c46e
zbd12702423a7dff8985924d76f8e9c393377617f5d3a98b2614e75603c856e1526f779300be713
z7c818f4971caec4ded0b6ecf8791b1129faa7ef8548a64c797e35b5ab3f49a3d0a46394bfc3994
z65a584935a32bfac78e903cfcbffa45c96b94ea492d754e21c712cb9c05c213f5e0ab2440bf86e
z0ae9aa9083a0c371828e46b68eb341b63af301fc9366e7277aab35679592dfc3e7146d46934586
z184fc8a8ed3cc7c3dc337a5ab73a02ef18c90c60307261763835fe4dac8cab4ec1bfeec416df8f
zcff756e9ef86f636584710a10a13603f811dd1c59c68704a76c42ea65ccebd512d597471550b50
z9720c579356138bbd6b1577ac047a9e5a57b9736504a567f5d276a5f62f437fd81ae6ad12b4544
z46d28fa20d12c49d2a5062011d121686c9bbce055900fa3fd81930c6808fd6f9203acd99cf90a4
za48f63ea0154ca2bbcb39d2ccf436731835fdc40b4e913edd83d1bbaba5b611cfaa2a6cb597faa
zd83f862b8c10dda193dc9097337dafc0c877ceb62e5dc735a7af5ab7b28148ca6b738d7946af30
z63b07260d426d6accaccdf6a37bac0fb99ec46092e1fe0d690edb63057225331e3075c47fccc89
ze503cc4e601300b71859971b6dbbd5bf6c6d5c37ced699a84f8467a34c61b86be8f23cf5d0bebe
zd9f987941e138694c10463ae97da26c6e7f1238c040fc0a1d1b92e451c888198e7429b69461ae1
zc63739dd81b895b2c51b156d0d332d9868c0fff4dd3140485d005ab2c55cd48c520744c6cd92a3
zd4f2b9cc6293c8fb5f4d3647a8cf032e59f2e352fabcd0f77708a7c76417e9fc5bc926705515d1
z2a6a0f58a9aedb85cd52f0b22d208181ebb650349632ce00f1e60cab83d89adbed7e8e720f4878
zcb0b595e7245d32a1a2ca33afc38dee507b83f6b85489bd678d663fdeac7a3f217b179bfbdcda4
z4bd406859ca09236fd9e01daf006d2b501d494c3fc991dac5f34d2d414c7f5e2a5c6afffacda5e
z93149731fd61586c26c611877c0bf57c9232a3d3beae44bccf979f4071a919719e4ec4c5ee8423
z82f3a28cb7149d40ba643c1a25e29c7c88ef4d96f95450a5808277a23aead0f3386a3a5db70f2a
ze7611bd48d903a13008f14a990ada01821309494cbd3fdae395695d430123ea3f054c432f9e685
zb5544bdbdcff3f1fbc98771fe97a69b010347f3b703916dbe885282ebe27f6e6cb9b4214b87e7c
ze9d8a80aa2895c629c363726cd5b1bde68f528c70680472154166b31a82c40d662fe546ccd0410
z7e6f937bef0a85939c3bfab54029507fea98bacc82379d4331fccfe9e75a7e7c5ad39b07d494be
z53ac834261606e2e81429d68d50d79497d69b7b5bdc544db33aa2a6e3585f69bb71dc8590baa51
zd08f5846bc5b050c9f024ded46808f1f0415956416547ffd3b1fc9153c0154b281e9d1e1a610c8
z2c8b42cd276496097ca4d37367112ac0ff4e42f584e2701f75c340eac1e4cce47e51cb23ca69f3
z8dcaa817ad0413423465e663f61aa1dd653fcf8e8b01e1daaa2074d1c25d3868a3144caa25e93c
z3b076df98ef75746be0bf37cb91305bee6dffa406b6c30eeb8d6d5918261ba6f1b294f3c692240
z5fa1dacfaa6dd9c6d73e229afafa138faa0f96241f128c56b76ddfca39b1e9e21a34ee94267879
zb8766104793b6c9c67b532d316d82e9b8d23f27fbf5f04936708a3e17565e2519536c2e2917264
z55704d6a8d12a3f1c07378633f7edf98d3af3ce33bd0b3a798ca9346cdf306533f784fdd45aeaa
z1d762032cb99120cb7c8fd13d85487de6be480f1024a77e77ed81db4cd956509b9495ffff00401
z7658eb997a57a8a6b100380b3eae394246ccfc3d0bf31bc2820601c996bd61af113f84e48055a5
z5afe912d9f0b65128698ca33a260e5a1563484bb4b1cf26a085db38a309a9a0af2f848ba6e5731
z6804cc162fa0af29567573319a21840f464437c1c6e52feaf4f9855f91d02ac41f89a3f51d96ab
zeccafd4d8e1f235d41f87a7f9552ec345f80ca8887fa6bf99fe385e459b6dac4cc794597436212
z8e637e42a65422995391ae6e3d044c3b1d3599ae0493c2221a2349723912fd8301e1743d6e4fe5
ze3969cb03f866194a194d0baa116485bf681035b0aa14f9ba5bdadf61a644b5847f6421fd8ce53
z9854d69af5073484e02b984d694ba57c653270dd99ed1f8a2ede7be64491c9c0b713685f55c349
z6565b2622066cdeff3fd0401f936018384061ba200c29332dfa65e37e594d47e5b30c0a90132b1
z6cad24a98680041dddff80b9492db998dc8a35f47939f78dc2764718a1c8d8d47b467a836d520e
zac92b127b11405ce52311d5c55374ee0d4201e8e92d6ccfb7fdd7a5f2dd51eefeddeaaa4b1fa32
z6070bc15d6dab43ad6dca832585d599173e47fc1a4a8e97b2d5ad364e8a490b7228975b072ccb9
z2d7f632635715a28e400f5e01ee55cd00819b84c21ca53b4f1181c884f8ae8c9db7b8a353a6141
z9fed77da085f2165588beff682792563e253f4467824888a3756770ef4d2138dfc3bf3d110cf41
z8cc3766cfe90a7d740711a7fceb19099a8d4b09aa88fc9cc0c593926a795b432d286400bbcbedf
z7bc6a3a99d6fd3b750bd29f423928e1a31309e2e3d44fdbdf21244e820331b9636679571797926
z33f32d80a4b16f6e41a05d445220039c45edcb558d2870da0f7b0fcb8271ea33ffffa44698c02d
zce49e3da4eefb9fc6704c56a4ca6b239b9d7bbf36013db6e73552d02d0f03e577e23994ef7d683
z39d83ca315c0de3f69a779fcdbd0142433556a42887e966c95154b2374b29917216fe3baf9aae2
zc304b4b5eccb428d19de53f6369508762f8b0d20ffe2ce9cd3ce0590c7a1a89323fce739d724fc
z73b4c2140a6b03ce5e90c3fffede86fa60f7e9a0d1415b21140eb9f59393385fbdc37ecf9beecd
z578ae193749c95a4e17fcb81951672dc09489571fda603f4b3b12235f0db78922f117a4af69728
zaee3fccd5e2dc5f93b18d20557b24c6d1ac19b3050733b71ae580b3d54996f469961f710924cc0
z6d2eac0b522e0a49e995ae2b4cf05c1fd38f4b8f0c0f81bd2ba0b71581679163677c238694d20e
zfc566c40dab31c3a59ec10f2624744e080d958bf8b19a72b753489e91c166bce6bc17198c81c8a
zeac785fab83eb023aeda72d6d9050989c2e1c486835e7fe8d340a35dc401ea876bd4004950214d
z99d7474d10d21a8a67fc3e2b4f14cd17234a95d51727e01cc9cf8b54266b8c893464bebccfa947
z9988e90fbe88082c33e3d96bd00aba39777a5a4e55cdbbc3f18f5c8735c6734d96900c42858141
z7465bdf0450a7a491262ccd6c3a521a592f2b071d0972bd02093ee034011394c7f0f4eafa25e74
z0bf7d961b46d01009767295d1bc97dc714dd4aeabb0240e11a5fb137f1549e1fbefa77ce91b599
z923063fd227c9e8361c2fa2d2c580a3a98012472f08f053005d51540e5051206200f19a5a55cca
z267a822f1d33ac06889be57e9ffe8546d40b52850c7cfe35f841d69d1599c8d9f13b7fa902d0e0
zb4331353478958eec2a91550f461312d5c3318ddd084481ba44e1358ff3c329da1b2886c5b78fd
z052dc826cbc71bc732396ed0aaf62273582c9b04fc00e190d7de847a17d936269aed101ba6b879
z849a4767db137c8b2f7604f78e66fbebf9b342c25fa618351883f28a63a653e1ffa3c99e7e360c
z59fc317d84447b4d2aaa85fe53394dc0d3a50909f63533612a8b5d79920d6c92f7b983f19f0ae7
z829843f0d2a25d745c8e589bb3ebd193f0d1dd621034d16d8fbd68496f3429fbcf41282b933064
z65bc3a14d4dfb64c52e8d93da705357f4fc6fc2708739405eb8e31fe1455b5b53d65f2e2e3f424
z86f0e34967600968f82518fbc52c41a48fc50ecb49e6995ba5f53af42115367382ed20b820fd18
zad2ec1a550c87a38ce4e93b6099f79bd082220bbdc9d7961868f230a6226ca76ced3c6caca003d
z0fd74cad98874f278a011ff7926b6baf3dec89c32ca6bc2e52ac922f918592e8ff1c26696e206b
ze022362d1bbcde29e67c715ae3e04eab51a00841e3a6f6a1182258d2168dbc0c9afa3a78d357d5
zaac19eb6a76b1eecb1dc605135580a79cb29499000f6827c4ed9fde150492135f556740b355b8f
z4f164929105f75ac00d3aaa6b6f89bd779421d72079be47ac3c0cd81eed8a00c6b1f125e696460
z22c8c5587902905970be0535bb329100689299fb6c45078d6a9ca10326b3fdced0987a0562e15e
zb26bcc0d0aec9d4f55172d98679c1cc6a34927a65a7b97783c5549b895ba63f842cf6c4640cf7b
za58d658d1eb635151e09196638545f639c51141f841eeb138bc2cf6750296798368abb8267f28b
zcc386fc9b5371f714117bca04fa093f7b1443500e52452cf452aad4d31bcd439d74d8036405de8
zb1364f7f14ddd5cc220bceaa1ebc59434aa962dccd621968185769498572ff93449ffc8b457532
zefea4dfac29a20d9a2d57a0600f3e3255485670f30dc4de08a99895cee5697257aca191f306001
z08efe5ebc944656e4cd2528957d96f71750ee568fded04c97e1fb17120ef89b54e6897fe103202
z0648ac00834663bc234a015a124f69cc905028cee511fc37278ac41d210792ec5fc99c5f5175dc
z132cd04b5daf07a7ff765dd297211f48949df64bb7e5b6099703d9a93368e6c3b2f9178681356a
z013983f5247b1e0fa0f1b48b05d9524a05df82d6ee5963a42f2dbee1aa0c8d05f0a65c96f5ed9e
z9273cc3b3ce5ec4546ceba1a29c435765f16f4f462c0fe3d2f251da06758c9e7b2f1c64d0f4cca
zf07b2c606f0d69a8a8b6a2d0af547393915a960d09fdebceabbbbe1915bb59b85605bbeae8bc1d
z060826e155f35fde8bd7b8406bb31bb1be7b0cde13b310c984011c3c3d48d247ea985ad7f5a4c0
z93fced1557fed6a03ad252976f4e144d5c1d8b45644669ff5e67257bab1563bdb517aa244b9da8
zf07c69be5e5743d5303adb5800f4f588cccfd8d4151633634aff128c5e2b3b5fd813025f476e51
zacb91a0e18704c193a045803423adb57f7c91fdb86ce5e5d8ddf810cfa3b0d94013e2b9ab0b7d2
zfaa9c52dc20ff16686527ee1a28d08720be507aabcb94d7f3d64731ca197658a5018a3647deac9
zc1d2233414f7d26cccfa5249a74fca69b6b18866cd18d4291b063da1346581d9a01d281d595d7f
z0408fd3c1620e2ac8dad74f5f0a61174f4be5cbde789095b88df90efe71fd31b9e11a801f4ac79
z36546de093b9e9b808984c44148ca2af34dc19592b6991fd4fe2a724d64291b2e6faf9e26c690e
z446ff6044d7d98001a9b16f6c5b7e73fd62291a9cb8ffe92e66fd318ac5e596164d7950fe31f29
z12a22f9fa26e0333fc902790babe874e221746cfdc7bab209f149d6043d17798a085cc6e2ecba0
zaa82fcb9f0a6255df1292f32a50c7eaa0438a8d2e2555461a6ed54317c0bf3ad91494b3d47c26f
z3087ec6fbe4529a7016625722aeb3cddaffe5ef8f46bb9308931017ed1b417516db94dfc6dfc89
z3b6a22baaffffa3418699add8181f9cb52a349d023f84df233355d9a7c574d7915959ead7835c3
zfa16980606f95b68e6c59b24483a702f59ad88e2ea45c3593540b5dc528afa294eb66b14ece2fa
ze959ca04da430dd12a0417a269332f58c3ef6227e7e292ab0719bf60db48d034d4cfbbf2b36a1e
zfa89c08465116f35d796b110d98ed5ec30ca7aa6c797fe4b072cbb36eb1734cafce3d3bf08b2ad
z6f8d3e7c828bc976cd1db0ea81be435e2d42c4a11bc44381750255f10b227ddf97f33dcc54da35
zcc320999c6d0c39da47739055fa5e595c2fcf83ef2f32c99239e26495ffb08a51b016ed2e77305
zfa33f51db1a032ee6bba5a9a6d28ec8b3b02f28f09c8f81e9cd3c58d2eb8c76ebeb0d882a26a72
zdbbe3ba3de9c38466e91fbe215f153d64f454b003503780dad7a6836693f2275ef36a06a468aa1
z3666b72f3dc6062437d09808db4e2e7393e6c108a20cdc06305181e97cf8912a311a9607354087
z43b59310a64f7b6bed8b7e3e295b9d64b7e9b184d180917d70dcd7bb535b4ee89de8583300ea8d
zea5c328687b9ac053fd70bc1073a2ebcf47adc6d36ecdfea7e7b20448d8c7a2dad80ac53840127
z6066e1e2230ece6f815b2f3eb13f8d3294a57aea0b216e1f62ce40177f03603fd5074488971803
zc9e274476e6d149c7b1999ad775d08c5a6334a944962149d5d99b0a2d19ab19883d7e522e06fae
z03cc5081bd32f987b39664884d4f495396719c42a6b999b17113479996dcd419fbc56d752e0087
z47b1eb825dee44c6301c545b2a70443e7409854b879b4219a5097b519588d2406a31e82e445d8f
zf3591e2e43a0f94c28d003276be0f69d8e73209cedb83e2b015895491370affed81d0d67767c16
zc5eaa4a6b1d58ceae33c75614485f4e86506d480dd75c1833032bfb983ae3c07520fe3fc47f23a
zbc6f6927d9a53163f9cf3e0d1037ca9683149fdbc566a1605b3f51d1d079c9c96e1bc0a10d1559
z92de620c35d2be38022b2dd9d6238ba36c4003a402332528008b66ce08c0f937d0974dba665736
z81cc559ce55e02e4f556980ebc9df1ea00efafa2aecbba73a232e4a52870ae6194c31135046337
z23513acadc52f157307ffa8ef9959e6b12af6dc50affcad31d87d84a687fd1ef64c5cb7844008f
zd8981860ef34fcd271c6c59b81e5aa567f73ff9a9d56332683394ca16ed0f501e97b26854313b7
z6dd8fa36a46b37b8afeac8ad6b935aded481097e5ae3e27c571b450f207814d7cda1d237b05e3e
z88d85ba79e4c0e4098db51035ee5c7319651199f19aa75a7c1470589f22a4e42835141a1f1458b
ze6f516784b48eecd17794abc5d63d8360d3aee062b20c1dea48e30b3e0e76d82368eec5eacab5f
z541f216732bbb0d816495c36b2faeb639b2b4b6fb82574714a400612571756fcd9ec1c7f742e24
z1605185f61c1de7863139b27632aa68ac690b461c20f0bad4be6d8a6128e318de86911753cfab5
z150cc36ff4181a4610fd59f1bcef851541b3362ca63df95c39d956f141b780556ebb8e0c1e0766
z86d5bed4b330feb38d6503c11859e2d63d6004f204f7f8f2b29f3a5ff250fbd0bb23c804de0f2a
zea696d407b21aacb3e767bc07121142ef9ccbb6194ae68938b4b352b5882eab94ac386f05595dc
zc57f680e644a9f06def1ec8bf14aa20bd8994d85dedaf3635b6349afc7383e410f578a9f24fa59
zd387722038946f495e5ff08f801c12e691fd6c7dc5f3bc9720aa3b7d34da9e963d32b8dbc553c1
z58b8c684ae4eae2215af13afb73d6b720f3ddc13fffbb3b2e1162ba9ec5a4605155892078bf931
z585eef428ae9d576cd26981b111b94950624b11eb9ab91b51fc0f0fc53fb227bd8244bac6eba51
z0dcbbcf8ca2fac2dfce6fd9238b11685516aeaa3adff2a576893a24a1040dc3a3ec67633873c24
z87d00c241fc7d7c08ee3a2b810ca06dc77569adce321576b7f16790e265f21fb124130395da3af
z65f678cb73a1641f4153a4b45700985188f06004bb161a3cdfd27c688d0c9dda8f542fc742f295
z75c78fd843d567ecb91987e1f6b31dfcb1a53fbb88a123bfae840d7b79073c6a7e2b63c865e4f1
z487c2224cb64fab49d736b24425957b77ec68f4648910901a32dca59e9db31aa1788546a6125ef
zcdc45c3fc46f87b8b2347fecd60fc98eaf03018f739900d8c86cbe536f4709caa301565b0f231d
z98f261506776828c3bd0825266cf01fdc4ef782888b0aeb9131bb043f56c4d3409d0e17d49f359
z7f4c52e3c9161e99c8b419ca6b8a168166cf0e7a0772e263d4de582143536a8acf54cf53110474
z07a82b9e758395d9193422572be35192c971535b8a24454d0a80fb70a7ddac938ce0b3eea8a108
z74c5b7c368ac0ae1bee9fbfd198d813aba396b012a5842f30477788306216f9e6ba28978bf54ba
z938e3fa07eb8c432641ad97022b8cfc2652bcbd9ab8228f3e19b21d9680ee64f18b7c3c5181f8c
za335d24875dae4ac7972eec085be3e688cdd283e5dc1d6b5117d1c018dea8414ee93d7a52dc943
z094b38944d4a499382507bdc11f8f0deef9a24795d12d5f211eb7fcabd76d0e639b99f9de741f0
zc993c2855f1f1381c6146f207b092bc2b3fca0f8f0a4711ea6644923a89ef191c04d52c59485c8
zf64fec86ccdf91d99e27ccd8ae892230f69ca98ddf886faaa230e15a7821f7e1463a701b145524
zbf3806511c81e5782adc9c07c1f46573a5c5b57ff030fddc68846850b18225c2eefd8ade61446d
z1a9765f34eb8397eeea4fc7a178465d79ba839266c4e848ed470c8e4725911d39a842d7dc7c9a8
z674c3352f56ed1aed3273b0b916565a96e47a7965af758ced2a656fcec3393c218bb4c377876d7
z35623d9a2bf5b7c76d85330ee77b77304cb0454ffc896a58f8fce07e5a4a9b98a26d499c8a7833
z91f614f17d1c590d8b0b47c6ac8cd56c2cd23167dcc71b6b644e9b74b45a1837881b92e6d2c71f
z9c1505c0991a2aaf51d461f77645d91ff86e4b0a72f2c55612b3be3e3b36bdc1bd163fd7cb41dd
zef42fd34115c5ec7a42a5dffeb6e9fd9a08212816bcabe53052935a7ebb1ba73f18e8e92f4f337
z7be54203194e394175e38f7f8432685e84819c0cf94cfff8d3fc7b58715efd3eaf27dc1d1d3353
z01a42213e373a69562283d177e479d2bdc436c522edc85e22bf02265f3e3da9e57c2941ea1c99c
z316300faae19a87fc1cc2683857c839abfe79030dda6c33ee7854b743d04ab931d176a2334359c
zffa462e2d766e545421a836ca39d2f28bdfb253db9fb74b0645f3816003caa8242133bd17dac69
z2e152ff5c2cf066b488bf1622cea0390c6cbe8943a425af7c4fc5c4409a2730086f93063f8db56
z02b19e117d53906d64002f407701be23c9bfd1daab553195e412407740878d0307ff4820e2f580
z11c4e00c34675667df827a8cf6c31e6116ac1e4d879fbcc083ffe88d219b99f85e178b31c9717e
zf18de9c6b3b3b228d504ac1ada20dfa21fb9dc72de57939c7dccda0114098dc8305d3889f798e3
za57bd9fada8cf1115e54814451b3d2f249b0894b5d7880edd790003450b283548cf97cb3bf0a70
z9685b3cce1c04e9be858599ad844d00f3b855cc7a850c1263553d0f55a8197738525d2ca8dfb40
zc9327bf4e81ebd2574e508e672af4abb212594c5a838438cfe72bbd74e6ee59f5d740be54d1a5d
zf66d320057297f36b8ccc0e8ff4031046dbc9d18bfaa231d4a833d9b47a39a8aef1cf77a79cdbd
z3845acce01c109a2a32adad83f4bb75a15e2205a0667b3168f1dc49e0332060124fcb535e90821
z0a7a25bfaf5f65d9da9a8df0a13134474632290ef95393fc28d95b4774abd8c954a85680aa0119
z9fb6866faeef72f13c4b5f472b83acfdb399fbccfae58aa6406aee325120f2a98c11b311f5e0bb
zfd6d1d645002b1ede4e7aba214221d3dee4066599235a6793b86f9dd59089b27e6cd1b7170205b
z00c3d9a2481b0d8ad03960871d47416bba7119c64ef98935c369d9256ba3a40b6df12762e94165
z8201321c00a0fce76589184c19b9568962e547d26e34b4e04a7d3911cacaff70b841206486c401
ze85063527beed8182ee0aa9c83b4e9a96fbd2183281b296789843970acb4eee37f943eaf6b5447
z036bb3dfdb7996ebc1678af06f2abd3c4e5eb1687bb30bda929de33e7905c486b80758915e217d
zae7a8074493bd47630aba6171d41406cde87394820216d6e5cf7704556416e15f08cb12436ed92
zdae6604ab896e8327d8a36f23dd161d2845a6d99a2952bb2cb97091840aa66b7f8e61cd1022202
zd2c43c6573737a1a92727352a9ef05bab9fd0e2b5c6fa78d3179b0e7c2c81e3fc035e07d421f4e
z67b76f2054a9b233136b5654c5eaeb34b0072f77b1da7f0160a4f2f96d8ebb364fb16e0662e55b
z307a86bd2505ff68354a96c1ecf85bdba87b7cc4bd9595e109e7ac93ff5c594d6490bc2070d62d
zd239a272426aae025360ae601023667ffc6c7d3e4128bd478e35eefc82b09e8c9b5c401e05b7c9
z35d3a31bb403f43f6ca4eb52cb21878fd8f3355afa26b6f2118cae554952df9e5e4f9547e55c1d
zb6cb2314999757c78c1bf5a1c3af1a52dc0b0802a3f8c9b5b8d8b0783a5f1c36b05e30ea111675
z74359cdaf58f0dae06fbe53ffa1ec1d6db85fa5c999293120e7b2633f0c01e4d085ab3218d0733
z258b8e4a0b75f74470155d641d4a31ee0fba6671c3646486b39ba4c0efe50cc13c1fa009bf072c
z8680167ac397fdcc3cc41c1a24bb499553d23f362d59b86b96799ad1ce4bd93f9048056eaee155
zcc857de31ca188714d30cd85ed5c30b2a4018fb642f0499b4d0875ee1aa68d50803b865f1a9034
z12ba142f9c396b962d5579b3dc3e4196fb6101a25de126bb7b04b46675ac2a4d311b85d833b842
zb0b35924ec3cd3f1546b12ae53f2d1b27913436614fc139e5d6a38f54c3846287734f0b5759a93
z3ce8034584d3a5d9d37d7cf98f69281a7599910a07b73c3fca570c34e90054f8f50a7096f62e50
z33f616c8e81c51fca4ad7683373338c63ccaff4febd6fe8b32e5780e7cbd7e2d4be0ea5bd5f10e
z357d5934d652318c3eddde0a5dd19f5064d1bed7df73786272d95f7501f70492c7be499ec7a39a
z7eaa5d1bfb2dd61e525b35611bd18789763e8b2269b08f8c52d25a17a0f13e65daf744a19228c8
z288e798668de1912117968e04f763b253270b052ffc037742fcdb9bf2cc7d14e2e10b7a55ad17b
z8df1ed0b4ae38edbd429bc4fff1c106e5411293ec5bf154823dd4fee04fbf662fe9d42708bd486
z4c470680e15996a6135c66917aa4441971c9faf5592522f373760fc7b6f8954949053c8f80c92a
zead731087456a14442d1444ce549aeb4bed97670ae52d239dd822ec2be8fd6eeaf9e74fee17804
z18431c921d0b279e5dc6585e5079ca1d038c4ead15c2170ea993a20cceb4268e41cb54cb54064c
z31bc7f3d97579f9222d9bd3c3fe54eaa5e08365b457b63d92771165de71307df841f5b2dca0ced
z5acac4b6e66a67b9e2a1ec2c9ae74659911edc48a956e9f83767f5fb64e2df72e904b41f1cf09c
zcba568f16d02602083500a7209d34dfbebaec378f1809dc67cbc8bc0ae037274aa1350252e3165
z5f5a706e797f9b595dc58534400df34b8d86468d29c293fc0ab058641534b2a215f3bbcba74cf4
z24b0897753347378cccda22c384ce692b8a288f9d27a5451bf6c71a4ff16736ea7200209a558ee
z7ca0cfa73c9ea6a12fc224b022c0e6a4867111caac165c482fdf9429f4afb7ab1d11d37fabb6f6
z5150b43fb5dfbe7b700e947ba0cdb8126962e33afd53ca78e51fd0626c0e93ddc7311a68808651
zba0d378c5ac1647bfbdfd2dfa3b3be168b7f909081bf9014f418dea7f0ffc653665a94f7a2a34a
zafd74d10bb88694022eea10ccf2e9a5c4855b819d73b757c3db3af3d4109afe4ac6341e0ac2e9e
z4dcdc23030647c50b013418696b6bcfe2062dc884b7018418b3f088c6f51c651129bb1cf1520ee
z876489d088634585d01f92166f58870136939b257dbe2bfc4967797fa8c34ab180a1a35fe3d3fc
z068828b2f0c03e3484b48d9e8c1948eb00c3e927a16b7e3fec8201960200f87ae601bcaabfd49d
z5fb6e5b91563f58e49f78715d29cb98fab3ab1ecba9757d8fc7f93a05565026f79e459e0ac19aa
z0bca672d9de753c70b7e986eb054a6c9c6b42bc1430ecc6be99e9822cc071668dc37605070acc7
zb5780a44c56acaf3e24e4ed247ac5ecaa2e40994f6e926951109ba97a43434aa5c3d46a492aa2d
zc41ed7d2eca2dbc88560f17dff8b2ec332762947305d3b27d52d349ea48ad61196f8e5182396a3
z3d65c83592e6eb511066377c2127fc50dd0b57cf62b8991231e235308f4fe4dde09fd66165e525
z68220b9126955cc1afc1a7f5797604d7eeb62422391963a69b16c398ef8ccb0ed4b64befa58aec
z606d869dcfc3f2182d1f07c6d78b87bcaacb7a61a7aa8dfa40d7779f2d5ae23cfa1a28d366070d
z450f48695c169510aa965dd1ec14bd154f7a88cd7c9618f3ed9644e4439825b0760d78f8344eb8
z5714524984b8f78c404e39f5d5ee2212c502c00a28f02f21d3d081fe4b2af266a0a64ea07858e5
z71e12c64858acc3996f59c15e66deaf1cf1fb3747a9f7562bf8b47723ffe2066cb918ab61a42b8
z5235603856a614b9b107b0e4ac978c4c2aeb370d3821d038330d0ef0b42360ae28ee61a7b89ac2
z9ad2067818d66678a849b0b0c934c08de25fe70958bc458bd53a8884561bf97cf0a67e2a452cb5
zc88c06eb65c5db47f057073f22a1947cc2147c5be5da73f92ef57aea4bc41361b37b6d64dd3a95
zbdd9721a42fa753ac6a2b1e2e6bf50b4469c741289ec787f920c786f5cc655c156923fcb82c363
ze374b7d8bbb576f4d9d158f462fafb63b70882d9dbb3af65120a04a56e2a19b8ac3790aea66027
z0108c1876b1eed6217dc915dbd14ea332f3b84dd3fc857fc6eb5d446f78ea42dd4bee652c6194c
zcad98b7fad22143b0048f417d4f9dcb02de09e333f26702855b1782ec048a32835e3ba00b15970
z99e07f3e71c8f27e41d1afa776d60e5389ef252bf3e7b25fdfd6b7d1f1b9aaa94f7161e412f5ab
zfa804df2b9770ed8866fdc586a5676ed18966fcdd58736f4f11a129732ad93a3c590c930a130d2
zcd3e3c526868e44c53b8349139f94de3d9303de897f592342d7d351d13f39ba1f072c65d911102
zf79d32c300765567f5ccd52ed3d883926a5a935413afa26d6313760d50cd237677da9d087c0f4a
z91308c46540e312a50dfb0688940a31024afc8fcd5d414b094316adee418dbdca7f814022c53ee
zf54c08aafb4a72dee539f04e68241dbbd4bd921dea3706690b16d79d482e1dd51b561582fb5e5e
z6ae093b1102a1e186cb39352bfa6b4a2a01c17a2aec9643bbcc2f9c68fea4dacddcad18f4f1c29
zdad768ec5dd0fc8d418aceaf86db86ee43e318bd4a56451e07ea796b20fd76fe4fc003d5fbc813
z4a0ec45b6d0478732deea1f26ad59a7e98ce06b53834863ac28a6b26f16bf3d28b314db17acbe3
z06e327e259f41d79323498eda7376104c261491138ec901da2634f51b450f499e98532923619bf
z774fa3458df2885b8ff4154f07984a7d8c71d4a23c4a992df853259f6b2f0f55001946a1b13496
zdf09d9f17f05e64e9e71ca4efa520ad5a6d02128fe1df79804fe04cc0d8cc21bb667bd1c9f7a53
zcfaeb77c0541ce06df01b6aca109f2bc50c3f8180c528a63d2cd09734807036541e88fa2
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_bus_driver_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
