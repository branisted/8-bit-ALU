`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1bf3f153bd631387c118a296ca10cbf0349426
zcf2ea5eb241fa84c8ecbbf7180f10eb9ddd4966d421e6ca571b198ed195474578ea51160ffbd6b
z0f73216703aef2bba31d04f6d0877540c760cd2535de4136d5bd4771107747c34c07fab3aaf6bd
z67c5eab3938266c996e67839bfd448cabe88dac2c17438997a3ee0a0543dc656070eb3dfe7c0a1
z57e24e01799b1ae1652a0133882b63649084f8bfaa3118d2448218b5c4119ef2134dee0d7a292d
z80c07e69250e6cb0856a07c01efe3f869b070b26474ff619f1ee9676ce10b0179ed9855d8e02bd
z3e17bd42a654e974019a7ca7de85bfb3ac5c169726f832c6b918eae789fa38ca70f5115a2ee7c1
zfb52b503ce6ce35b7dc5989bd64a1623ecf327040db427ea1518177d9f8bd73c5a5f9a85144832
zce11043d3366841a1a219f20d08af9d4197a26c0742e77ce0e439132af699837b50c44ec0ca068
z87a83cc53f69c7354f63d64d6e082face2034ff5b7851fcbf0f4d3ffcfc3e3b3a209b142a948a3
z370b68ae858a75f8dd7971759e66525859f09b792ba0fbf728431c52587e7d8523ef44fa720f3c
z0436c86f8a131a2bf23d43391fbc8309086056651b273906326242a4ba4b0212ef6509b93f9530
z362d388b4193b89b1430fb4aa1ee4a65c7ec1fbc29393a43db0346f983d1b801da8d2132271e35
zd25e665581429d363a0aaf17f5b8728471d97a6b84fd98774368cf0c8f8f5e78bdf184134f2109
za762a2ede8afd7dac92d479943ce6895372a5bccecf803d7041c4202fa52cba1f9330cd1702fdc
zd4dbe9a23a563e6de07d97dd27786a27e3d9bfcb75ffad89c47a7aa08eb6293fda57b218c8fc07
z35354e1aba6a99c0b170dc7c8e29c04a487f19e037a3777427fafd568284f349d65a3acf96c2fe
zd5bf44aa2a8dce3c66e1dcdad13950f906360f2afff66f7e76733b9c740ad5352161a3822623d2
zb42de3f3a0e0f519f7d9a1946ad7af175b8d3b1626f772092fff9c66841046ae222316a91a38ba
zb0161f17852ccac92a87240f7a5c67abd2fe6f0c2883fb84b46f1b1c7050e21c60e85135f398bb
zdd2969b70756ee4564c58cce85b02812c2772c4e724c3f265b67e47716a97b81b2159ac4d5635b
z44203371c8bbc11f413476b470887f5baccb86813c1192ac3702bf0421975a343e079faf0e7557
z0afcd0b46ec141b54bad47d8d24e21d9a1a0fe7c734fa13b3e0307226831881525a65d05541467
z0a4086d2ddbf2534d8d116ddc008a0cff79e4a1233156c5b119a987b9ae9e124e7462a0cd7d88a
zb28a073d6b42f2061bb240a1d38efc4676f748f0e304fd1c4ec6f30cfc86fdd38fb636b7cf712b
zd328e152f2813fa5ff08c92262e518429edfb305c7d09f3194431be8e8623f783d2c7f1e15a4b6
z106b40d839aba7475620662ee643ca11b41e286f38cd1328a0cd113b15491b53aeaa69664fbaa6
z40539a8122eafc237ac0eea9b4096bd21583e5b5f5f581e7b822d90356a6f2efd7bdc547f1fef0
z7964bcf5b46e20532a19ff1ae263fbf177cebfa4e4b0f49451f06d282a3691015738aaa8da5d94
z0405948f00c819fbda7ad627818e968191c67f2df04d8aab038d804fc3bdc4c82cd871b7df31c5
ze58d8a7f01395bf608f7cbf8ced58349a769d507daca0e54ef8ce5312fcb74c1ce90d1bff27950
z6bdae233fdb4eb109868b5e518bb26845c29086689aa3195e5cc5212cbc6160dac997f1adf8a92
z19f31865d005c1caf9b7a883865709a70b0d647062214f7d9585d1e96dcf1bce47674d35adbadb
za0bae81801f1274ab25bd3a602769ce43cea07f11f5ce540b02155083097c7bf1b9c827c479bd2
z2e574a624bd77a996e2a15c1aebb61f3394297a6ec3e6665564aa6174d43f123427d1c99c88320
z8c95b3a03eed988c7990fb321724a9aceb1572469d6b75f4d932831f75b36d26a34d11f91f9888
z38f850da9ed34fb4d26ffcf13050972250e60f351161c8394b1d95df25d4989cf016484bb9a126
z2f7ad323694068f478ebcd245b210ffeee3dff2adee3a13fd8d433c2681a35816293ea164bf4e4
z2d4b0076bf1e3cbc23eb9db5fd96d51bf28938e679f1092c08d97e34c8b26bd5a365c47c027220
z9e9a1055ca1c648fb1658ac31d5163fa212047abb34c4fd22b73912b78dbd552dc02939d16d145
z22278f52ef8c3f0ee39d52e6ef782c10095398aaff197950986d3274ad08ef65738eda4bb337f5
z91210db101499f20137cd86664e09b52e6fb589667278a5f83fe3ae7049846d8e3ea62469e1dc7
z28e94c8c1f25053a512ff72f0653542fbd5f6c917b2aedbab33c5b4a439b6d7fa5b26d2cfd437b
z0a2376c27c7522fd3e9f38769ce242fdf0c3b296a64966fa242c57fdd2388bbc42bf07a9c021e1
zed53ffd5eb75c75649c1c6d6954123322b2dcd3e50e6d4d32dd60fc5f4b0d41a62de58bc131a44
z10a0f8859153a4598a53184e8e3f1fb3f51f7886e50bc1cc1be0c7804b060b7b09f2e0527582e0
z7d8884481ec5a7d22e3d54dfa2381d62a6f67c0265cdde6d7646fa7d2347543a68f7473139be8c
z97520d719bed77fcc11f21c79f3c47d464d8bb64a5b2a011a19335680491344d4dd9b5609324bf
z33f95d0db93efa11a25e08bb6bd631ffd464f8cec97e739e6a70b90e08c70721c72c38822d0831
z3229930e37d5006ad6eed71e88243a16f0e1e69eebbe6227a911707a02010581a752260ab6dd9c
z045255dcc0b3c24ef6ffb18580d8b29382bdd7250a8ca9214b7a72f2754cdf6fcf04910bc64090
z1234ea00a100a86d216d51074bbda093708faf358c4619db2c9d9a3304287fba66ea86e1a6fd37
z83e2dc40181d3caa6c0f446c1808089f25f9000ecf8974231a54dd3a3173baedb36c63edf0a995
z39023f842ff7440575aace5b0be6dd0d159a22ab8806972a558ff379085421c681bf7fe1b93adf
za4ceb1ee8d424125752306e1b9a49611c8cc0f5f5804b069b6bf25d01fa9c6693e98440708a6e3
z6596b8b2a33b687b518260d8ea15946182c5ab4f95c18581604786a499b1b29529f820a07e4944
ze4e77fee829dd7c2e2981da2e2ef899c31cf17ee67953a4fb98eed6d11d80a0da10df0f78381a3
zac7adb9913222dae458a8e483f1ef1a0cf9b1d200c7a3322eca1f3daa5870bec8d9e76dea0da8b
z9475969655a62f0e86bb4f41c54ac4c783187b4cf70fd3bfb41aa73bbcd9d3482d6627f8fbe095
z488e34281c3caf1a4cab5c4e2d6c713a7630ab7fe64fd93aff4089d395c97e1d538b07ebeca2c3
z3602ff853f2f9dc75573f77f27559ff6640e7e8b632d18e845131edec7bc198cf5a2c9d4987eeb
zaa6e2d647daf930d84ac99d9024f13598ff63e3b2f96bea482fbe2270dab1185bd0d2e2ecd2fb0
z4484ecfa4e233e8406e729afb1eab8b81e6e90781bf2c77802fd74e7fc20296cd985526270c8e1
z177e2470861592b515795f7f0895921ff5b321eb55bae4068614ed7abd9d162865ba65608d4d6f
ze67eaf5aafb171ff5858ca737d5d907469da9caba896ee24fae163bb0ac4d29a257cf439c18f04
z32dc54f2ab773a59efecfae17a522ab6dd8890c4187593a65fea4fe4e516c5c3b2001d58fd463c
z46b5a94361e8f8b9ce7367a7e054d73265b2893e1be60f8b531f72f98284ab08784edf589edf69
z1e3f4c2162624ad0881b0e967079ec3a03cbc88d5f1654db71db8041ca8404db11bafc2208c02f
z43d0bae1dac5de5d9381367e2324e8400ecf7ca84d2be2741cf67bf585a0508d5775d80fc14a67
z6e1e4e13b9baa990e0adb8ca4c8ee8256784f0f71e919f150e94a62f2e80bc1e2e05c152c001cd
z5cb9574e12dfe8c962eb7d8db76982101c045dfdc4cb19bcad9fed9ad553e5883153d0860226d0
z9bc4440d0c400248b5c26c8b4e0d655331a370d2c12f39f72a36d583f6bf136d908ab7dc093cdd
z84939f06dfcb7acc167dfb257a7b9f0a76cd5ef97368ad09ff4d8254439abdc63f9ced411c2984
z3d6dcd56bfb76f54f557ea4ac79534aba465ed98bd4611c85e6ae5f682b7c744201633851aa045
z25bd8f4daa241b930e538070eaa24167b08f0273781fc206b7429ab415b27482708309f743c959
z36da3d4a42f2e5fac90fbcff214a337042e79ba772e1bc3098db4d0646e83bfb7dcde93c08d30a
zda42ec98801e50f6737c8bb665b11397473f18b7298b4e8e8b1ec74c65e45a2bb8ad571898c5bf
z230fa8fafab2ad1d90bf5ae4f0fb4fd739478b221dfe400548fd903660a5b4e46ff98776576b22
z8c267cdca3345c1b005ed3016ff1ac5def16c456a75a1fb74ae4a9aaa977cd5c1402de3ae14aff
zc809a8cea80a5afce3987584b30f9e82d21f430dfcf0b546aa5279260daa4fd65e91919afd546a
z61290108f5434a94ad3fc2e1c11b897fd7a21af95d5eea1687d5d6e575d7c7b7dddb7376c2ce49
z468ea7aa13f462a059ef7b9f69fe41c450be477ead4d17b21cb9b058609b380a895ae75cd5a9c9
z5957902ae0cca45372987bd0c1d729ef1a738cc872f5a0d1f0995b3ced4e19509c5ee9e8258472
zd895d43784843590f3982410cb55b12fc830c26a1f31e62c6a7a1263b40e1e75d66ee9283efcaa
z03e9d44c98e57b390a0f34bd2cb887c0ef73f58f49a6e0cf136b41ae8f58144395fffcdb1081b2
z4a7a5bc9a970d6c48b8510a9c650d3e5970220acc5bdc843c0aff52a342b40b00682748634bcea
zfdb2d35792be732ee43bc5832346fa385eac8ca5251e69e53879d8ebcda92a3d8d4c3e3b25d5b4
z1db0a5f28c2550299ba35558c32a78787a36b9189b76844b449fa9d99a7096444cf13b610f9b73
z2c7c340cff94c77fce8b81828d1c96838f0878b85b148dd4e96b82879b59e31680ace39ac50318
z28c5eba5b7e6f554bc6f71c84244206ab1c82015a250ccb98176a1575ad1d9c59168e234c01792
zb31d2a54240c08de3d0e49d13d850ec0dc626aba44a09efb4528e19074e6c922b9fa8fe4fb0039
zc87343a61127bbc00fbf2f6288168db8b4f4f993cf08d840f8e749edb359986326f7389d071de7
zeefd6e077bf6f9cff6fb64208f63ca8b8a711a23b1d6d50310350ea0cdc53367439dc19c9e7be9
zda0726d81280942c3b7cedda73e374116ee6f49a4780fdbdcfa5230e803a5b1ae55b130d6018e3
z17ef6c3ccf90ddc3d7c49c4189342f86213fae70e4da3b6e4e14cdd88c93fa47a92859e9232051
z47286ca98120a111864c25259026e68551d77bc93f9ac84f94fbda5adeeb125cf4dad9983b1873
zbd1bfb12a936043a27d8991d9b2f94e688c683a557ef85a71f7ce50d6ba1d4d361d844cc75dcb9
z107b90d1d87c82be90ce617e3cb75c5c7fb0b6f52971fb82bd0a9456c25869a445bcab2660a8df
z8577befa8aa8eea21afaae227c980a04c0e8e8491eec2a4e8f0213f0961218f2949f148a16df48
z82685d33b51cc554db5db6a4e52ef6d396d31e5cb2e26cb65045c6917a6f569a60314203b64b25
zd315dfb22e2394d336070475014bb067f7b898bc38a1d6b4dbdfd48a1f3e3d028b7bb0c0c63242
z4b2b0f5b527a6b2db27b3071bad39a3b2645a5b8d490a0f113d29a501531d199953e8916de473d
zd553c7502a69dd831aaa9178bc0727da58a650d2241d1ff5def893ef7098e8071ece19bacca600
z61c5bf5caf4395fe8a1dc2e497c57d7482101e1dbb444a6e5cabab597ae131d081c59eba8c6deb
z852f61d00ff59c51bdb42bf73753a512262f33eeb7cdb540129663a786333b641c3f67d2d62bd7
ze6234d2dd042d5bdf806194e8449a7dfb45b7eb7714842bd6c65bc6bb6c2b294b0941c16cf59a5
z3a8c94fe254a40602dc5762a0b73bf343cb78947cf52b01e822c2973b62d7088ab97ebf5f26dcb
z718081693c88fa6c86c2a47ff022436259be7d0d41ecaf54f621a1d76043875583c0e444a456fb
z9802b754d1db0770194a85f91beb9f1ed3ac85232d75691ab8f92d1012f0a8bd863d7b646353bc
zd878334b1111c2576f55bb45c437ed90ed1421dfc54699be155a8e749f23de81e07693ba1a93b2
z59569708475a6b6e1983cf0f397dbe6521149f74c5dadee74642c91242f7e9ee4c155fd2802bec
z0dfbc24418debba44617e6754e314771e173f66ee055e0ce8d99a15bf6b976f90839901b531d6b
zaff91204459e1a4bd7e22d75e0f6fb391784cf5965b21ce84e9fe88096c0a5e866abb56265d22c
z46ff43927e6551d27b74a8cc9b72ae30cdfdeaa4c18fe29bcf2acf6eb8245faa0ff8cc6d7ebc92
z9af5146f670d83de71e4ed7b00a874700b50cd0525e66aaced0f64d1d7133c2ec303a9b0287ff4
z737b9386f65457aa626c647de62693f7b0e11288e57dd7274b87573333725c97839e10c856d415
za88636b041b9dead2ac609518f756c4dd5e3708146c0969f97d69e92b968906819f1a298aac8ca
z3e1d4d4e7360fe2bcd733394ce55f1c94f11f7e19d9a1a009eb8eae65359adda08b5c8676a255e
zf3baf6c4a4860f729f95af0a3bdc169b4c6f9e0b4cd6fe4378e257d1467ee872842be45bea8bd3
z9456cb32806d15e5f964c1d048d26467360bcd439b878697aac9fc5ab6142759a5ea3bb9878acf
z0d2a3128d9931ead8ed3e7920aee9a53e9e3700ef70960ecce7fca51d9d6756b051f4c3e8e037e
zaf4800d7238ffe4563d499aa2dafaf2ee14e0b2b5c59ef5b069ace5d9774d52c1db2482836ca06
z6bc28d492f77f29875c5225ac141e4ca046c2958a4b3c7a72e72fdeda5f8cc0df38a6282540900
z71428860878e17724b40362bbe11e169b2205a726655fdc760387284377823eaa45b2950c1db5b
zd93e57c3feb9ba36aadc851d8fe3573eedf5ba63846251639c2c44654001eda5ca9c7750fb0c0d
zfaad49c1c1c615c1b7f4894666e97dccf1325dbc589fe5e6400030d626e196314e0c9b784e5094
zefca5c3f7a3e93c413f4b41b2a44d8ac031ec5d5b43d80e3d1936e2fc433491d10a8df6802c00e
z8cbc0633f86febc302193ef2bc2fb18361de2e36eecdb928c00f7f64e8b89c03b52ec2beba7a9a
zddfff3ce7ef6a27743d74d9aa5eba780f6b0773b6dd938f9f01e3a40db154040aab4423b34cceb
z27f458eed48611e32715062408efc3fdd144eec679e303f33e347cb0c48e65ca26b9edc4d2340e
z9157431f37b09d98717b932cbada44c86fe37adf10e1ac28721ef129fb9d602ef9e16fb1c585e9
zdf8a71655b0396b53107c9e413e91dba18df8a69c61e5c6721a51b3d024d313a966973916ccefa
z519a17e74c29de9e7ceffaa1d55e9de910325b0710d8fb427b8dcad4f791167cf3baeaf255a645
z5ddc64a55e234f77988e704a75f0f92daaf1c4bf456528cdc125972deb97928873fffd14ecd305
z5eee7dcce62b49408e27c6f215e8eee711dbcaf4f8dc77850991b70e5a513803243e00b03bd22d
zc7ae4777c6e0486bfbbfa2abb3ab76c2a4498cb88b48670aad54be626e1b638e69b1b1027bb6a4
z7eeeaaf3e5a72674a03cfeaf71a73a79a022c28e8c9372ae573fd4e8afeec9543fb1b85504f5a3
z426689ee17ca6fcc54936863c33fa1d0097be69dc0d6b077b131239545d371e56a33353e238a21
zd58eaff91d0dae51dcc99e2667f76d3055a7f3255a9418383878f6a0827c7976fa452cc1de364d
za2a9c886a4957c7d25f87cf7443ea0eba56a996c64382b92c681db55391e059e59a631dbc79eed
z934ea0141f85da04088b13dd199e9b59ade85ded6782ab518d9e25db843a532c557f697c3e2f9b
ze6774d1af80048571b9af668b237e6d37ae96b712933d949524884cecb029fe4220417994ece1f
z75fdda383ed328fb108ad91a24b8a38287f1d7c71e077587b90fe860290828aa4553fbfd0422a2
zcf1c5a3ea2b6f46601648bcbde3d8dddbc785f8675efc7724f8e58c64313f8832757a40c02d935
zbc9b23ab620cbb62e586607ee44cea0c771e617baacc2c031f659d1d89ca056d577a0ace67b801
z257e801274ff0a75ee644813b34f2f7b4cdcf96c0a9f85694cb47b4dbee9b2da67943ce14f60be
z0f86bf173790dccfc5359feaf345eb4447dcea7094d0596d617c55b917f6ba731034775f98907a
z26d558883ce367a0f7cacb43e45fc98fb76fa1adce0299623058d9dcf9fe602f80c8f5bf5e3584
z92b51cc56791dc1646c6c0680bb6560cc326e1832569ba089e7b77e35e68fc1cfcbde5c14351c7
zf45617e9f174c6a04caef3b38dea1805772d08f5f1528f5bf62f04fa35a14a98a9274f1f8cfcd5
zfa624636f8eced55b72c3e537ea16cfabf17e755d3b3093dcb6bf0e252d40c4c937810ed091e48
zc9cc81aba7aa99fac147443862e7c6befa75a786c67e0c811f3d5201657ceb787f5b7392502316
z0c6076001f35428fdd37c5658c5312de00fd1bc6df94f0a3b8602e00ce11dd335ffea8a5b249d1
z9323f185e0d433224b20019d1768711f2160252075636ee9d9aae06d38534bac03d87608b19613
zeb71c0dc656ecae84d515efda7850f91439af52011893f001e4d176d2a05d495e43b3880124155
z5c7f2084e15e8ae684839c69af66bd504b4aa38975cc21eeb3a78fc9e8a6e643f91d2a06eeab7f
z5d9c2e0fb98ec41b7382de60e3a56bc440f136f3dcb73829f68380561ea2e7144fddb3e82975a7
za2ca713ab9da1d93821ea737cf54d0ce99abec11400403532e64234464d52634a329a4705c163f
z57ca62a90674a28bd0966e4824a36b12cf4e6b8d68ac85d1bbed04ccf94fdb304f3ff413fe6ce9
z0e7a9b9a4cb4e8ac1112570c9a002d7b68c7d16246368c9a02e22c6326c518878a37a9a934b4c1
z2726a5dcd5937bf50259996f2d01030e2d3bdd0b369cfebfdc8679fd3e59ef1d5e458359605a7e
zac16fa56d45366eaa1fa9b6e4db637359a7189ba87379a63c448fcff3cc9d4ace9bce11a6bd70b
z2f662a8aa42bfff7e2f31b29c2567e0a07b1a16e3ac4ef725699cbee041ab79c3434776ca72c1b
z3f927d0aca681690f1cb9d53c1ef8774065e5cab1372c0a3c38ebcb13593dd32c856e5cc6af301
z1a092614ce8d73c94690d999285d7370ff33f55be0a70e193fff448ae6dae5b372719c6b3aa0dc
zf9ce75db1589e3805715cd062d3c8f5a024bd98ed6104672850d295c19d773928e3ef7b23d37e6
zce3797f6ab9d4d835549e0f8250fc8db339dd52fb8a2cb593b70ff959d52ac1bc60951e37e4789
z0a5ddf2ff1dbac0d1aca9b1968d08e1ec99b87fcd66bf06559eed063ae725948795f1f427c8c6c
z85f105e7e78eadb76c6dd9611c213c0a4573811b1af7c2ba6595d56937ccc1f1338695dd6db0f6
z8dd154ec17419cd674720b4eb14666df41d9898a3e939fdbf67c5351e1e1cda86248dd58ae4daf
zf7178dfadb447a9ed2fe013c7fc2e1374c09ee445c12487fc28142f3a7e9e3cfc7122b0e1fd033
z9902e057e14bfcce18dc680a9b4a5d19a33014ad90b0b2a2b41bf4735467af8cdb5d82625773c3
z221470e5ee78045cfdcaa58a3f45a0ae7321b17a1070fb3df7f35cc698e33d0ed6ca8bacf870a5
z1118c5ce57f81867af96b80b7f6b55f4cb7bbd9f72e6779ec458b9e8e3c6c9479b93d2764e0d6e
zffe5113cc8ced73cde546bb0777ee652bc2d5f7d4603a8df435bcca2de06802bbdc7b88674ed9a
z23eefd8cc4d1153c66387d1bd30ef7f1242645bfdbf5e23f1d0198d163354f4ccb288237111091
z9662231eb6f1521553a912dfb22f7566e3c018675a6c831f1c2f1ad303f6ee569250dada88a671
z6cb5c25d793c4a51bdda5de93fe1e5e2a4176416568b999a40688dd4b145384a56dff91c385e1c
zf63723f2438d1f3a0418910247fbd99b0de8e0048aecae1c808f072712505ad7351a7a4bc764a1
z7d80a5bee9079e73c8d1b4be9fcf2733ea3615ff7848a9b0abd41270c2f25aa1d424db7d42eebc
zcdd7bc0f5756f9b9679895fed7f5049138359b225f213431e35a8762f39ca6d5db714415d3bcfa
zccaf3e01a04d1b7698bd4136a97f99724d1b4495a819e07587964e28b167e755677d9c1c5a8464
zdd1b1cf4f9d6544c9c7871151bf805f6b771b19c89af6055d357bd6701501b2f05f0bbdd6e17bd
z3271a0757c9141ce3c72ba21a782726fa1012d455cc7b75a5880b8711e3739baac08f3440c42de
z86664ff8fa8a0ccdfa3f4937ed68b388e7d1dda4d279761f161b1eb19d27acf22c7f50363b5553
z94a46bab6c033afe466345bd740802264f7f0a7334731d4ed9c3d3a2a2f101f49666631c3c1296
z0b87b51270a20f202abb8ba51954940d498f1fcaaa6a977d83a269a8b05d21ac560a58e541c6e3
zb36307c89bcdb0f89e761071b98bd1ec6ed36d69c8176ef43aecf1be6f8871372278d444a5a7e9
z2eb6300dc18b32e7e194a1355100767578838464d37360696164fd0ee97e67ab47b37b5c7ab3bb
z5063ca4558752af1ba7781ef42ac8b86ad7e201fb3e7b4113461db45d19bbaa70ee521831526e9
z1d916099406b102484e9222025cc9cb87b897825c4a6421a00c2c343eaa96e61bb269fb4d7c08c
zbf515fe78e377ba57fa623b4b53c26d5e8e91b37094fa7937a715672b1a538bcf568f46ec20bf5
z898594a019151cbfc33fd7c9702b3e446753caabeb92852e3fd3fa848cc3cea53e2a83e8157954
z7a662c866307147bee9f333fbb631f54a7d6595ac77826e2a13be295970549ae0dee27b6d273b2
z3b7b6e31e481126e84cc17e35f319a955bf2c894f76669c3e8ada07ebe95d393691a717fa04f64
z28b362f5efef095c53a300dc0cd970efeb2aef2354dfa066161f179bb797bf5d6ad08e5fc245f3
z96fb83e322f5ea37be08dd30e10ebdd090c2152b2ef791187de08acb05c2e0b0d2eeb55ac8786a
zd2f9dac0102cb8e81b13d23bb6f698337c95915752f3ef4ccd40ef6c39496ee192238e9fc6da68
z03fa7cdeb5ce8f08dede4c681abfb6e926ed11e133fdf14b3cf1298dcf8155664c87daadebb1ce
z949aaa39aba1ee19a4df488171ce13b78e01525fac98a7f99046aecbaccce8087ee1c3d82f0acf
zeb7a1bff0296f0a11a364dd4355aaaffb390952eeff03457ce941a14efb0b0421ebdb22a7a0296
z1e748c839a8052f959b62546326db7f0507aa957561db96eeacf975d1b2e79833c00f5ee8838a3
z819ba4df2983f218e122d11469f523c2bbbcaae638a9f2d81a546ce0e5bd1b3ba52e408304e295
z65388cb52729b1d944fc30cc4169e4126212137f37daf144c3e309826572bde6848d1a372764eb
zce77a695c79acafda92bfe09b3527a12d3d3e2ea8b3bdf414bceabd3b720867deaed8ea5d0ab7d
zdc8722fdf9effcd1bc5a9b4153f0709254ac2a05727939d8c4d59c0d351d4df14a44b9068311c1
z37c5c8aae3399728501a781d7e2af847c8ed7f0218223301a9b415871ad0bb34867f6750dcface
zeba037ad3c81bc6d26dee6473f2d50e48bff041b14d4fbee376bc302fe0d5180980b2a7aa4da37
z7aacc72f0393c0a0b7f5083be8fe089c54bdece3a69de4fe9b49bd3e585f68fbf88e242e93710f
z366acfdd756b570a0f59af1b1da2cb7cfea9cc2fd9ecd516f017a8ef47efc32ac4bdded0c1436e
z882cd4585a289d0bf3bb9bacddb1e8663c31afac7a561776f6686c82ae2cc564919ca73d93d039
z1736638d26c80664a8e9bdda9f5e7880c98b90df6f45a7fac7f791079e1dd600626b0eef948ac9
z40b279d9e36887ffbf1e0b78bbef6846749ac411aa82d57dfc441b46622ea98b6dc9975690ad18
z34bb95f2aae376a733ca14d2218bab5f55190e6faba84af2a8f39b6100b06781d63d31f1dd6654
zff8ce071f33b58f79c47b0685efed91ce06ee583d68afd1c4308e7d669fd6e1228f45481371cfd
z4d39bc6b13164a86002d1b58e0b850c77d45882d60030c504a8e132ea82814ab0017fa5ce6ecbf
z654f8e7fd26fd3b378e84fb7ae97fcc6a0deb6fa8911c9dc179a51f53badf74c3b676bc7879b06
z57ff330d5e1462c9f2b4b84a08c469cca7a03053d7f6bfeeef26b6eab45831d536a376ae6c83bb
z8e6410b434feac4834cc4145ec4be7670f5c7c5be55ab042df24e20ee201bb76d5eb8be5508c38
z4f5b7b7f98c8fcaadce0b14a1824e92eb51761cbbf1b4c5fbb535e026d1fec798662e8fdf634b7
z6a81f66234acef5b92d154022e0b360a6b45bdf084369aaceb7a99084a7bf0fa9644c13769843c
zdb5ccf5f6f81e318fe6be587b8af5ec21c5eaaa8e06f3015c82e963d69054493ba558280e7b641
z3096f2a11fdd31542b110b96a133efbb381ef66a4afc169caebf6c21a7713a837001823620a64e
zeea4f6642f7ab9338dc37902264bcce1ba8d54f4a13164f0343dd28cbc8d172fcdedc41dd75260
zef4c7be87a655da4897dfdba17e85ac05097485ec0330aa4e2c7ffbd8ef35a4d1d47de90f8556f
z09818e400591d63d62072465cb7e3e229af186105bf451688835f019569eda775c6530940c9ded
z378f02ea37360a0a05449484aac3bd8045aced176346ac8d3d42f2ad55abf150fde45afb120ad9
z57154d1aa675e8053ff5a7beeab9dd69b16bd918d1a8eb21279a084a2d934580e2211778723f68
z7002bf896c5adbf6dc03950502d0e9add8271fc1be34ed0f48598c32d169db2c6d6560e806b85d
z4bdb7046db6bdc3fb110ce2d7174882b7764049e8637fb179bb4d4157b40b19f1efd83620f61e6
z774588856edc68af7f0cd94d6f81b993ba24e69a305ddb9e064521dcc2b6c490c6afb63ecc7e91
zc744d77e191ffe9ec8c4e300ae4279fe118f6a9ae5578e17155cd110a30d717c4ad5ab64db892c
z3bc547f66524c1dc861ee7df07d12d02f38bd81b9f93b8f7f788204187f083396b24b076e2cb8a
zceb8e67ea038b690479e247ca54a4e9fea897df1e46bf714e4f8eafe5d9e822eeaf0e51f9a92c7
zebb958e26c59f164aa9f73cf29a245e8ceb0fce5ff7f9bebcbca97de7c7d0a0401f03f794603d9
z310a35af1c6adbc31c86f879fb6ee122659c5656faf153faf7a42af5854bd670e8b2b8f109a9e0
z253f9f2ace67a4fec8316b73d25b30a91fcf9ad91c128941eab23fe34c8e49ba96471565505b42
zc3445fab331f07ca9bc036847dfd6610f3a10f0adc48a7c27674bf949876d0b1fbf8f0748a013f
za72e99193e23eefcc9e31ebf417bc6dfbf9a55a51dbfd56c6809aef8e8ccf04f04bee449466b4a
z561ef8c045bfefd58ffa3b7a5f0fb6e404395581064faa1d7b0fcd8f1911b502035738a463a8f5
zf4cfa8992d7ab453013f056768cf07ce93ba69f9b49eda914c691f578c9015438face13c909d6b
zbd6c21b62b5261ccfb816244a4b8937413d81273cb0e4c8cd68c5c2f7332cc61feff05d24145bc
z2e701fe5c3c7580633a4754ecbf1edf629c997ea2f1c2b7d2dceb8bb2081b86663b9a875df4776
z2ed72ee89256a1d2293ed33eaa03d33c65078bc77a39846c99943be3bcc2d299056ce576f1a4a2
z1f1434b997583a84e900dde2b98a2dba2f277522920ff37a39cc88e397aea374afc98d850b03b6
z160b71da8de75e43434f9d39a2ee9e66251136656e35f2ae1973a6fc12431b03e6f59b20132aa3
za1d22e467f6667a3fd7254a81dc6d98c708b54478483f74988965f278270d22ee86ac41d4f0c36
zd69525739f31a141c197032ebe52268a68b06d5ee6c9b57f7db57fa9ceaf3b4a76b59d710c768b
zce3b333014cdc484ec25f2c09433370bf6018f95beb6f19bc537936da6e0cc6db22797c6c6fe69
z9442d4180e8e99f8b459dae7e3bc3b3c2466e6e5d9b86be9cb72ac8ab8d13da65fbe1a6587c277
z248954eeb750a167f1a72143ad3bfb9399c9409634428ff1ec656f7a632b1d96edc3c2fd9ecff2
zfc4d58764097008bd634b523eeead9192f26d241b582045d921bad1493c10da373ccad92ade975
z1d16b90701863c260b6116e2c1a582666555666c6d6cf274e66d1d6c4192e2bf3c4344a72b2e84
z59f9c662a0179a624b9848e7928a8a54c378a237825bbb73a56d70315dd7e62552cb45f47a36f9
z5644feab9ebb47fc594d5e066c4a8dd117085d90fa859249ceba8b6e96f36600a8209bf0e66878
z1cd977fbb045f766254bf782b777df82348d218284ae8e3801d9a1cce6af03c2b5ef72c867a116
z1751fabdab6e206bba37a5d01209ab90673c64bd9d0bc29ab2f0bb2551a3e153041b4d5afb6528
zad8b9858019a4fce71eee89af63f2031790348ccdeb24fa21f4776d503b557150cfbb2becd9ee5
z7199b312061e2d0c166e7e7f8a23d5251a4ce72d970709cf2f0b3aa46c2a11897a14789d2fe1bf
z74b7894d3bcccaa38befd500f5b16313d822d678227fe6211c45ea40849ff0d9ecc94823280788
zeb32e1e56c2fdcc251789fe32c256a4d0d2f32873296bc4de69337c7568f8db7b91025b8d17105
z2304da1bbcec9ca7bf92b4e6ff92cb83909db7452e994751fdfb1eb11fa5b99fa5e1f071f90236
z9b1fe89e00ec8768132572a3b5d11976d7076e5e1b46f32a19fbafa5fbdf4d1936a9b273564b0d
z15282e230fe04b3dac99b29903e913d2083470407b9fba436243fd7ef18358554a9dcd0d88e40a
ze94ab369f8cabadb365d6e4ba40bf3a6d14609d6b99a19d4fc98c0985a3d4a83f5a45d28b24369
ze3e1598a27d7e4ac0ec7cfc360d334848c0cd58b4fe35cb69a74bc57291ba3c783be9d143c5355
ze2d0bb064e715ce478615b30796667727dd4ca1b370970d994fb301625277443baa7ed8befd676
zd09511d47b19acb7c1fc572b4ef9f8c97185e19ace0280eed71760af738eff0a190284a3e60fcd
z272b5a5267e1f37522d246aedc361f54a3c23489fe7224aa444bd237d349df7abac433ee1bb11d
z2541f49730bea6fe4a99daaa8d59f4dd1692a44ddb64ea5f1fbdd5c8518244771f4121bd52137b
z2c9abb6090e5ac256b1685621a170ac8edbe51236d6fc0c85f4e07140dffb09f5232a2f9c64a0c
z5ecea1a0f64159fbfbbd876004eb74755985e85c46c263ec5835041db93a1a8eab50132fab8120
ze79ff0ddc16d808ed62b7ea855fbab6c028a1a32d59cf8acca36025e13b13ef9a602030825a9c1
z7882d18c41a9185a1b2b990fe24ea9b7410dd4a579169ba283b59f41f4e7841f59f4d637cc6d4c
z76c19ef567f5427b5b3081f78225c236ca374b55d170d430e9c55182f1b7f6373194ba1f0f4028
z01c4cb300cc965e8f7c751d318a18c5dbabcf0621d3b836b1fa8733303f2e74777a1b955ebadbf
zbdda7211c47fc6f8b4b35fdfeb36a0f5b764ac90e7fac3d088c455f6b448e981f877d38c295709
z72010dea0a8356a6c18edc4b8ba53a29fd8c92774b9ac97271fad305a9a2a105fc8c173c082da8
zf7891a8331e96e3300c3e8e5a2a28a39c081daa4ab80c012a5e93050422006ad8a1eed667c1dc7
z6c98a0c37cdf6a68052686eced28ed944cef7fa5668e5faa8a4d01b9aa23f04a24ef860d5e99d8
z11ec97b2e5bd4142aaa48abb215cfd463b1f759d1cca18ddc746ba7cd7fbaeea83cc67fe5966aa
z0a73d73121bbbd5912117c33584e94f9aeb86c527c2555fe011f285abef76d0805718d46e97093
zbf62610bbd28381ff9af249bf837c5de98dda28adfb1df2842ef52c31e49820e33c1b2aee774b1
z0b78a011d2d7596336f9b13250518bfac572dcd7640f00fca510b2db621449df1cb9ca4162463e
z7c94c40f7fa0fb4047f2be86c2cbeeecebad4548d19f9e2888a9819c2c473fd35a1933ec488935
z56da5117b5ef1544375b51d3da33f0ac4ef921f6033c3da8ab242c65ea043b161466fe4510af0f
z66897df5b6477fcecd2828040b61f3177baf1169f333a544ae5f41c3adff6e35d5ae04e579e814
zcd18d941fc914061314a6fe30320806b3c45c4534f440fdfb36528f230f77adc2ab19718db662e
zd1347e36322d6749b970b7ad4784ed7749a375d514b6f2a7a5813298c6b0d12ddbb59c3ea0cdc9
z2f9a68ebf19e23d68048a85fd705fc230cec8e90b7055d2fc9f5162cc1ed238ef741718a0dc133
z1545d322a125c3b5f94c38065d72defe4d61e41632d43a6aeb2cb446cb52b8746f815e24555c05
z3dc8d3f0497890abffa7a25498c5929bc903f0ad64cf145ee05daad005e0e88b6836a224acbfca
z63cafe7f1abac01431bf10ffcc6bb28cde1715c2c7a94738ae3712db946fec2cec5bc9f291f18e
zf32043124d7bfa140c467d0742dcca34fd1ba7c15b0fb600ea0db66ea6f0ffce841a1e5d3d847d
zf097ad1c08d14d01ce8f5fd99f6ac8c0decf955162bef7577f5010c9c7255a208a1dccc9cdbc26
zcf2d065b1ac9a6487c6f4608a443181f7bcdc4790bea58126972d32c3481dc287cacac7e5bc6c6
z1a07bc78a0849e33420e32d8b63c74719e4c65883ec4bf807e558ac8257150ed9016c1cd2734c5
z6a4e754776dda58a67c1ee2ee2c79e9bb4456a7f1c1023f3ac25e662d350a9ae65065b696dba21
z61e3bf0b80ad6d265be265d9afa0cd1f70ea04e2deda7b175c7909f5643aa2d634dd9807832e8e
z84fde72610e356afd9551de42f194b7ba274bd040a53474a69f8f1cab7c17e7bb7a48cb70111b1
z4f2321979508f56a86f1f261f56e138ef96d1a9914dd5cca7bccd35264fb116d5ed026268fc58a
za351fae01f00802234413d6b19128754f1a645abbb9483a4d8abbf9e1399ac7e6f6cd5ccea7cfe
zaac43d35e6177eb76548a2f9518a68b2c1cbd502dc9476c44c45c79bac707ce9e931ed81ddbdfe
zdf57c679348399ba88425d7e641c66010db08bee202a82d94089458cc38e22d0343bbf4245e554
z59671ae6b08133e49209cffd1f83b138a1e06a5e95c113811961c0f3438e641d9e9b121f48cd4f
zf80f0a306208b5009cc7611fadc9e07a1ed5156d22674c3d75e3da02707d9565cae4a03eb0d516
z0271fc574b596f4375ca44f4ac61f97b26d6ac71c41384615a6e5784fa1408456b0afd6387ec94
z15ff5eed1970e14ebb7a32a3e477f802ae7fa0defaf2ab1100a4a41b491c976abdda7faa92bb3a
zc76c8966fc487375bd2107a7479bd60311dfc51196843140e8f342a8e2e7f0979c86860520cfe2
zfa7ae2f73977fbcff5f33267cb7b454d2fa5bc2e3f01b967f2fcc62bdbb8928d3dfffe555c72a1
z0d66c230173cbcb5d4918c91f40e66c1b4750113429fac97fae206d2f631a8018dd73522a68696
z1f72f9c1a6e6200bb334cb2ed4badd79ba7fa166252db1c264e3d6a5d56aad85a27f9427ab0545
z52071f29d40d194413fcc11b4729d9bd77d6d34932d728735ee375055a988ba9983bc1af5f27ed
zae5e007d4bb3efbd899fc6a6499635bd0de8b3a0f5b1c2a11ba2cd5371ef5665e9754bb77bcc7d
z33a41aa597d551c3a5125cd01b2b488906ad3bafab5324aa740a561f55c5335e8c188e1dac8280
zf104da80f83f389f824d99be8dba1e7b729b048fe0b6a66918f2d450552779820072e23c6df868
z086815b759b5e1c6cc942db959d427c817c51592fd5f68ffdf00a259106ddbcbff4fc06cbeacd9
zde9f24ff9feb32ec21e596924257f690b5f33955be167eaf3e0a97d2568a1190571a56031c4fa5
z0594cce4fad311ed0324a1b9a7e858fcaae73ed8d183fe29331800c859dce20953b0e75f5a73b3
zdc4faf90461a4a7b3b65f69c9125e71c14d96ecaa6a5bbedf99edf09d2f35f63c67862a259a942
z59316be49c67266a11a8fcfdf222c081884e2b26cee996aea7a41cd3b262cf79f8cadc7ab04228
zc3cadccfd20e8e933edd1595f663af4394c45211b68d5dce72a8953c5289ecbfd6941e67141fc5
z37a1f2a77487619c169db77a53a0f2f84939a7c656d7addf3fad5cdc957019f4fe6d4bbe4f8896
z9dd6fc1c13c60be927b732d7b7b0f0134270cc6e22ff46aa35d5dec75de1f3344da93673c70388
z0aa995d28707e5b4c8195e4ea46b7cb2c33482884f3a75f3fda5fcdc341647fdb5f15b3ba863a6
z87b267fe033ab64cee04469476fc8947d2b26d7218c8046e226ea262e7c1b161fe59118a007def
z0d2b0f2928960237ee456fe30a6b5d58f2b1c7d1736d81772ed57e1ccea5ead480b68dd43bd9b8
z1e649295c5bdaf0081f4d0440a29a1daf7009772bd21ce13c3114582ad4f3cb5a05264ec48bd5c
z37df2d1ea7d49018392e9171ad59272c150bedf2a30ef530e05efe78f0c0b77748a6978a74f82d
z8e1cd85bda7b3e5c8d309075637f5929fdd2b3f718ca5741c3516183eaf76bd7f2a25306b68585
z5338d05460504aaf941658bfd68b14271399d1f40272246dd3e1d2eb58764440326a4dd21a31df
z0de3617a866be93b9e53f48f3fa629fc03ef2cfd84bfa4330e17d5080acb755afec75f1aa5a96e
z35a3c380b5aee3033932c14c451f31ce4a97e893bf05a11e50a8fd2a7da545869007895cd59c1b
z064db76969556f9f932c0ce2b72c98d65d057c86bb4ea02ef11089f792836eeabee54562794387
zf49be3fab2afee84c5ea8f08c4f23e466daf0c175485144220abe2cb0d186f0771f789943fac30
za483704a75ad30d0d015938f26534c99f6149352ea8c5f2f7b1589fb1ad6a6e2a1040607d39916
z7b42e0339341a2ad25dc6558d46928524ba63d02bd299abe2d5a198b3fae4dd4d80a58c74dff73
z6f82cb6bf697ac6b3d82506e763c7bc050663e61b3a4b6eaf9a5c4ded6474b0a738cf2895fd3e2
zddb0dbba94ecde4aa53a2db22378feb16ede9aa1337e579a3a617001be36053aefe388fd928e05
z6d23a539514c3a6c4ed5ff831b8627bbc5a9f6c665f795a00d1149187d5043252de9167208b629
z11e08c219abe6930a4e5a1ea4ca035b8eeffd3977b8240a6db4db2bade2d9ff395e4dda4edea67
z8e5b7066031ef351dd8ca01b65c3b7acbae4c2b1699d1e8bd8da132454707461b8ef0aac13a641
ze18e810324fdd78d969653a156fdf0fff73c3fdbb13051110a61ff176ec5fcf0263993b72ffbe8
z91332d84469d66739cad9f6f906de00d89aec0adea884b2c1ead9c0e3e64b1bfbb83caf7a5fbaa
ze3bf468ebbf28d9685a884388c4684050c67e10bf549b657e2f6b9dde9f3ecc916cc37adfff9b9
zaf425a6bdb2ad77ffc4ef8eaa09090fe64ebba703027830c4c7907229a7650e15931c34d21a4a8
zeb53ebd6467cd6cbc8852e6ceecbdac7cb2543ec3b72d49067b319b8af272dc4727857e6ee3547
z6230ada0dff7e78c81cebd72281fc4399c979d2badd46f0f4464461576770e5dec9e32feef4d85
ze3c1cc233923fc0d273f72159297f66cf74148ad69210586a94666502af2a7f5d45bb766130d2c
z5f761e5dcd8645a80203e99b2312b6d7479ff1424dfe4b6fb1cbe80ea38d4e3cd8821f20331962
za1cef5719e738f6c61c1a34ab649f5168a63ed09718a3fae91b51c51904d68875aa0ec328e9a73
zda1521efa0ec28bf8f3e61d6c24c9a6c544e1342a37c496fc51caa65c30440d839d9d9a5c48273
zb4a7112d041d7562ad01637aa03ec700374b91744e3bd4b7405eb77e185743775938d224dd58d4
z0946c241aab2d88f79618cc2925f952069117a0e21f3b3cf1abe891f145e1ffc6d77c598709d97
zee65ee9416b459cd0fff9f0194acf8c36c815dd0bc1fe8fa9b4efe220fc609051d66bdf90a914a
ze51f38dadc14db752606fa5900868381ab434a8ee7238eaee7c2fcaa7c3bdd785a464431aeedd2
z9f573937dbaed1d4c3d12ad285545169a9735bc01437383d74278b516fc66783c358c0b190dceb
z3bc80f146b8461b896d0916d62e056579888c5f0cb5a83ae2ec2fa6955a6badc209801e35db531
ze47b72785b9db8ea6a0166b8db8549130d9d069d9257ef5b83f559b4c5dfe825c8006dfd9bd1b0
z4fab72637caf91ffc622337feb4270470a8efdc081a7203e601c8b90a33416c4e60fcf3c7b1ce9
z1d2862e6124695a683a7ba01ae0364e59913162c86aabd08a9e49c379dc4706765edfcee87fb85
zd7d5a388d9ba93e88df3ed0d1f003bde1b5d3b8b93c2933a8f3f24fce1483142238c2aa7f525cd
z812a4f5edd9af7b7b76c6f7d87c3f5ff547c590706aa61b6e67cc2b38fcbcad544a919994bf74d
zf72f441c941c7978d119eb96743d3d6872b83978f80fbf481403e14f60fa3aea400613a145f38a
z6f3bec24933b432241fac75d968b4eb88e8bb438d5287edecc64aa6412f91e540d10fdbeada6c5
z31a0a2e71fba575a2151f02fbe221d2edb11336a465b3a6f73974a4457892de0c14bf366a3dae9
z0a435121d100c8dd13434cdcbdc3e135d9ed07311f5c71784732f372a41727b7443fb75b2259fb
z96b429ae60d3844d5df0e8b9327fc381a3b9e28b5f10d4a7ea0757b54f9ef040a04ee89b2d924a
zb731d761e0898f27d0edcdb57b81affbcc58c988863ccdf21c7e00744d1e4ed6eb56b473fc00b8
z8ecbb6a6f70f668f84e1ba47361e5c902dad6810146549b13ef5b254a38dd97e99dcbd32371a05
z04f6fbd7b1ead530ff92b66b3bff3e076819fe644ee682f497e1eea8d476216c7ad88ed3d4cfaf
z17f950db2b0a65b75f4addb41b6e1124719b5fa6d106600d59f1db4da24a0a32771e8ce8a37d27
z4b41108c63aef173af96171d7e28ec2b995dc639b2572980d4c76979dbb48657beeb1245b1f38d
z6aea0514991b0f630ca2e35ba990e485deab7384d0a941eef2193afd8349bce95940ee23146595
z9cfa464f2b1cc641b902cd0828d5c490cc967b3308797e47a80781b76abe9aadfb3fee31c80b99
z5c82a65fa17a611105e7c82e18d663d06115937c262e0d5403f517bae925b8e1c4f3caad0bc8ea
z218b613a0d8d3cf39a0dbbc9933a205fae160414c2bb9d003e13e341c2896988ea11feedaaf4f3
z8225484134e6ebc7bc8255d6437a23e74371448d816ef14ab9a5a93b1888adb902afa71c64f545
zd822b0fca913bdbcf8a01724caafdef7d07596352220cb58c75f04a37edc583e4b11a74df2d558
zebd646c2ababec1bb98715eacc9ddf00ad71c620429b6179444c01f203111c74081110022bb02e
z1dbbebb139756e00b1d7a392abf908604336f12784a85d391de30fb3bbf7044306a7b7c1f4da66
z8388952fda84a89558de3fcab9a665667098227c5863635dfc55be9f99d2eb662924f0567cd284
za1e66ec5e66cf369d757c2e770fbfb36212298e9eea9ff054128f957c9fe28f1188440bcec2ad3
z1f1364f5ccfbb73984b979e4f559ad8620e33f4f911baefa28c87f504a44c36a07fed33ebf4ed7
z761c026e09c97e969fdfe0d3d55751905257f218ae46542c5acb57a4bdb1219f1cac11f7306a76
ze17f90b7300304520ee06ff928c9674cae099dda640f12d31e24347b6abe404c7b0ecd5bfc7999
zd34dbce0b68c9aa58e03da97fd932658c57df883620c0d0ca928bcae2f6ac36c4cc1e834d9e3c0
z40600598d6489d84114ecb103ccdac349d3e8c95ac790eb5448fe0b7de3640ccfdf89b1307354a
z3db77e0f024668621b85080ccc0ccb2141e3f0499093081b18f641aaba03578b6140c3d1da4f0f
z0050511ffb9501cf078db0ffe0bf78d6d82027a7ce2375cd854c7ba95517356cd8e81159d1fb86
z6848e811cbdfe2a84aefd7403d4de2d0d66d1f3861f32e39a01008331ee271a6166964255d84eb
zf27ad7ae917dee30650bfbd31c1b8e72ee2e554c009340af20cce65d0f3bbaacb97e4e3e4a9dfa
z388edc7fcd19108b9e0f703283ef8ca036f716f3133cb7517eeaf2e6e69124b324f3f412289ff4
z9da06b91c805aa375483573828383c2e7c5da99ed47eb9a4f3d83ee101786e97e3bca752e91cc6
zfb19ad134cd32cda960897104d06d6bb726acdb21d9b1983be76cb48047dd5425adafb144e5efe
z345d46ad17c13ecd2730621b99ca48539c537ed432aff676520d3206543af1af2551b7189362cb
z97ff492e66563eab83f16f7ae16b5344d400353651a0c4c9918e6acd51876cd89fec26347ec3ad
zafb3d41e592b2a43d99f0dd22dbb9e216c91c9c18f8500746d4db5ad9308854589ce8bdc722452
z51b7e2ff3fd1bc3e7f0fd5ce01130bfde699ac96501c6880e60d8a50c7d9fecf8ca0b181ff59c3
z22fb265d9cff2e27cdd171f450940c69f152e303a076b5cb0700e522f48c9860b65160e5a6de26
zc6a815bd998481c7e1be3195ddc10912a110c87ebeee30b1cc7ef7231b0e5febf5dc3926b0203b
z9aabea2fee90e722aaa2008e9b1ae2a57498a2dc88427455bef5c87a6cf9aa96317e0aced8c8be
z30622ed75d3ed9de02aa4ab59e87ed4c0e1a0b25954b96fad98217f55fdd6cbe11f3cbf6dbe7b1
z1a248a3b1163c0f9a5c6912faea9bc530a70503a43bb930c7c17ddb11771e4bc7ba7132934a2fb
z3fdf38985c8ec2d5200d5147bdb6b197e09fe5706b024cf9c9d033ce8485fa0c2261cc9fa4888c
z22ebde935fec5747e943ecc4914d7704d62e54ef8c476821ce5fe240e88c91b4d4b40cf6bb632b
z0d91aabc10661f23c5a81bcfb80d9ae15de5113714f97711a6c09b1d58aed5ae028182fddd2a77
z043bbdd352bc897046f1a260fda386ba32c5e898bb1d7fd787cfc0a4ba495a380c951071cb530f
ze426bcae9591dc843d38eb64aef14451bc356f3d11b013fc344d7aa9efa31166c828e17577b105
z3d9be9217b539697636a6c23c5036e4549f2427c7bfa1468ec84164f0fdc75cf5ea8d1b66c7c24
z654336d8198308d417f9bea8e594cea499b490f5001e1680db2371c43f6036e9466b6aa01762d8
zb7136d2b2543f107a6a581be22a0d28f729695a1c60d228c4e80e194631d8c57ce183cd3aeb90c
zbfd7406d0d400fc62f18ce5f9f0d39f09045ffeb07d0afb09a6467069efa66b9c43c72465386eb
zccb9e9e2205550ffe66d0d294cc0044bb5d4c844b94b5282a998946ed551f5751d35ba27d975d5
z0fc64ebf2016c69a8b90ba78d88d623d70718b57cb9513058862fa0f007d6ed57c07a7d747d21b
z5ad209452004d1d4f0b06b3685561a757271a804652e11365754585491f396a80a1c4a06bba217
z1ffab01db1c391d7113a4c13f444970074ff815bcc134236969c8ece20aeef6103dca9e1be0781
z35fe8011c88069e6fb067df48deebd0dedef6e578e46f81c6b7c7dbecfc47d65a354756e4455a4
za9a914ef8e07a1aef0f227812f73e7853218c4d98940b30e230d54f01978bb8be646fb050b973e
ze5f0a40f4d02362229c75f23e9aa028a02a8591628ccca68fbf897af3fef7eddb1ef834011089e
zbc54cfd7e9d47db53c26746372c6c59273d7b31efc72316e0e50a29772b3fa0151fb46ecf7ebee
z5b1fbd6bb0c71c8b226d3745ad5deb935003171ddfab928341db76dafe54f03208b6fbe5fd9aab
zca67f5e7555834138ec2a74c47f76249c9fdf9295523b3b636dba573c12e02f5fe7041c75027bf
zc85a41f03214cfac621555de756dc16b5d0287b008f2124c01f3913d28cf3e3e3e76b7f8c7050a
zee6ffcabf88d1acd93bb45de6ae5d15aef6610a76adee0c197d39f73a855d6b7d62bee983ae7f4
z773cbe658b720652f0ddd43021a24eec2119f0ff2d573b792d92340c58702f4762273daa53bba6
z19c55e0b1ed835fb712d0c978d818be3eb6924a86c9c2e63e2078fc5023b46e497b1bd11c66410
z73636720bcf30d51d21da5382612d9a3d52b6fe22e56c189f94735b285ac2c5c9ee15e80686512
z6ae24325fbff79a6ced48c2dc5bf5683037f45ef3aec03c08c9e20814706a88c008bab6f00b44e
z2f4f0b8be30b4f97e5e69a02e91b9a9e1ce42d7d0fa1715f5dc3cac4ca1ba4a8431293d8ab1c54
z35ab8f91ac258ed523555b87cf79dabb0ee2421226a164bbc180d66b094db84eb85d077caecb3a
ze14f03dd5581cfdc33f5bf65d50dea740ea8223741381f8a2ec400322a55e7b8a63edd77304c56
z7bc4ce199f184e03152388d5698ad67adf6cf6e1bb5f61ace60a5e5cbef40d1f812d035247fedf
z2463704ccaecae290df10f47fe4980e97b312bcaaa27d3ff517d93f7d0d2ff8e4bf65f61c7700c
z2e373fc5a22363042269a2d1e265c25d5b3efe621795e91dd90813ab7d1d2fd31d13c6671a70b7
z5ec18bef30bc559b67c3dfabd4f9a5a0bfe591b08de49fcbbc07f0c55991fee6732442119bcba7
z3101fc529dc22648bfb510c40a751417c8fa04e8bc2db631782bf0e84d91da3953f297c9daad1f
z9207b092d16be6d60bd9589ad9fa2cc319e6f1f04e09a342ffe9c9f80804c7e393a602daa4e01b
zfbf365a5bcb0478447bee94f2f8924ca6fff801b28f157d4e5e4fccda19bc49d58747fb9c3d62a
zfda994bbca7d57617901ad2eecb2eea76508f07428f8ef3135c546f5b542d045a876b846c986c9
zc63e8d5cf86874fe458f96ee0aac03c00325e322d224519fa5c06e0fba8c1f2919ff03c0150fc0
z6b9698019197efaac0168192d8e9471bc33da5b3929eeb94b8b368a9461ba6ce962acf2767097e
z5b8b65ffeafe2169f86b5376a4222be44cef32a55cd2d5f603fdd9d288793b070f72eb46027096
ze822cb633e16f076a37ae206d56c1e7649f614bc323558dddd34367ba71d713eb4760ed28957ad
z7a6504d050fcb4f20d1e81842fe90e2f2c7c225dba9b750f26fecb65bf50c2dc6d142dac38fca1
z8710a82c1be7f64ab84e073a1ebc6ed1a7a12f7c73524945dc18161296809aa0e60cbb0d4735fd
z49fb411cfa79d9faaf8ace06742750a80fbeba409caf2fe32b45847618af1d7f631d64e504b494
ze7b2716908a490210db94a2af07f7f4f27af8628c34714e77c8ca5f221aa6f2a8281378118db1e
zec07d24b6c3ec1d9feba8165c9a1925e34e7acba194aa7abfe74b688aa92f12406fb998210c8b2
z1914d0c84989dfb9c8e61957061c66bad0dbe82687d56626592eb100534e7522a0e3962d08626f
z6c90258e424e09c86fc137a2a2f74f21e4143bd3b855ae34701773b2e1a980421c0271098ef0cc
ze8a931b25d4ab02d676537e2f524fbc763f453aae19041e6c225348e3be76c18bc126a522ead3a
z349cfec064bd768d28c1096040dee5ab1c1a39cde9ff23969047168adab452a71c8a3aa7232d33
zc1055e3f3bd334bb989aa359b61a90aae74023200467f1767f2136371e8d23450b95e937f0b0bf
z0dd6890cedef1cc7514298a68414e44ab107cf606cc44978a004c996a31f69795d0b42af4da931
zef7311efa7f147e39ab57dd4d384790269e0b6534f8f05d6fa6147fc3dbd19ca60abe13ccd0af7
zb6edfbace35561515ebe2922ee98d58de28b8f8b51c6d9f39eb3b41b8fd68957ace86043f5aac7
zc595cda09db1606cc3c24397e4c0d91fbc05253c816ac4c84a712e4081395095a69d38c9e04343
zbc4c25c44a3870e74e8f970da580611c926791ab291412779a82bb900d7ede87dafcc75d8d8bb1
z1f193aa9304caa8ca1f34faeff167eb7552ce84efc53bd3eef7d4da1d573776c1f09e8d2821e17
z5334924621df63fa314de599a83a5d84baac60b5fd1c2c6cd5920f07da0202629a4d047444b3e2
z1a080dacbc63dd440932cc0e742ca8ee367131a6d0e535af5cbdfbbb65cb952d94a0f0f6604cfa
za95cf9790c3ce1a086dc3355a2c71b0f18604861cff597731c518a6aeaf0063b0e93c8fb71c534
z4f97ce6ada4385c0b08391c3fb57bbcb92ccda7b20d74baecb5674477f26e8babd2fa45308cb4c
z341492d8644958f2dd73eeffe28a0fd55b4f9a94e9951a77a4edca56a3e128284a7d57181aabdf
z638a637588073ac2bd9792fc1c4de6f70dab8e4763da1b7945d92aaca5cbb8b6b7ac4e2ac6ea5c
zdb1b51754973d213162ffb9f650865f7bc8c2dcfd87dcc3783f3e6e8d973077af14770b80111e3
z206192671f740b03cc31ee0c5fd45c55a5584d8783d3542448a0328ca5b5e46235dc860cf10cfc
z81738920af6c475d75d35425a5d100a0f22e9320b28a9bf414dfc853d31c2e860ddbfa3192971e
z90faa1c0f3ac1d7793cc3c21b1236ef4116522288dbe8e8f6259d1faeb63025e8166a2306d4dc9
z508e467d13b2a0a1f3a5f634adef12c2afbcd34b7f2e5cffbb6306b326e31979c3060c69567cc0
za79f9261037ae513339ffdf4201a929feb02f5c87f42f6b4c3609e1167c8fa86604026c19f8c55
z0128a115b96d0b944a7f344abb4d6d4996cb7df204be480502c2eb09ed4e4c077bfd0ae8d377cc
z6ab09349c3f4b5e4fe504af9e71ef42c1cfbe8bd50de634f09d946441d9e8d41534943d67d80b0
zdb5421354d4b10bb28de28834e1fd7df97041997b33198b4830882a385b5e8bb00e9e0e0ff4971
z6481cbd73cad5b85f2b75bce64e3b414e96ab14e552fdc199af45271ec361168a596119abe17c0
ze4678b4a3b7fb68a81d4b300b36116aa7a1fbfe3f0f60d486e27f1df353fc3a239b041189b8028
z2ad1fe5281b75ff206d8b8b769aefee748a15785e446635f2b9d420bc31c8e3a1c1d5047fc3832
za13803efcc108c3219fcb94ead6d85a64a5415ffcc361e2cbe16edc07b45fdf12d0076f587398c
z66cdf1bfdc5a618d6abd38be6a702ef529aaa9b6a7b59d3ca05a5c9d0e3f7507a7647b20a61c15
zb12afe55e08224b54448eb79e9bfdf19252c7a939c31f3ba13ad825625382da1eeb2731df4f8fc
z7fe8c33ef9dd0e94e096a2729b0dfe47bc72f57b0a0f3898b18d26313c31c71ab2c003729aae4f
zd34b2f09da355a71e793db75fce36d520afab2f1145ef9ea886dc2bc88c62cf153fbd2213b6633
z3f373aabc67c032b3e2288d7b826f9e87e16c75f00a10290c3d6be3ff9a516882a68e072e961de
zb998a541bf8a0c4d55741a7aec4693087836b684a3d7c5cf1551d148b2067b3d45d004d734b825
z33b5185ff7f1f8b381fbee474d77ee0d62d0b1003c2fd119656cf83a70640d19a7fa563e9d548b
zcdc96ed206c5bc328b9374fe938cbf9e258b9769e3ed11cabf26faf48408551a46abeb69249ebd
z04b782534af144027fc49bc048476b34d99b7ef9c780bb6d938f2a1de354497b820bb05847c268
z1ca9ed14fbe0d8dd8854128a6ad711b10e9572cdced3bc6105f217dd6679577a64de8f7374c220
z8ee9361be4e89d957e1f96ef5548f9a26c6dbba6eb61cd1c7664ca86c5fe13d5088a67a4d16865
z4f74eb443b08ed894c72e815346135f74d37f42649bb57eb7dabc08e0089722bf865cb092219f8
z8d1870347fbd35ba1cf153cc5dc489c06417b9a7516688aaf1e49355e90a634633508819808f66
z29bde1e0e0ef67d1b7237e0c66bbe8fc0b183fef1844aeb25e5d86ba65d98b28f44b75fae58367
z3db0ce057890f5f2a5fe15556082489a714a7ba1579abc93ec0c46d82e8c29c2f05faa296ee9e3
z2c33ab29a89e981aeefcbce5a83f98d774aab5cdadeeb7620d9ad4d61a568bad55ed26ba9445d6
z6a4578e850d5bf39dfa2d60e0a6e204095f7f62cf06477e54b7efa47b7cc0795cdf017c56773f4
z8921adf3ba4511ca57429ad5ee04e2607b38c3bd54dfd0bdf6a854af10346de7de99fd9ec8ff67
zef9ed1c904b1ffa90aced54d64494e89e685e7ef16b15c07bbb35b45a4c0dc80c8078311178d27
z8e7a41c62a9c7a3698df1bda0d2fc85c0cb243b6144e4ed0e197e8b1b2ecf87dbc5e7943ed0213
z9098ea0dbf04540c7dc2dde207633dd47e4ebea9549b233f2e89a1051ae0c0fb79408e363a417f
z8f84039e63b6d4c8613a5257f11630e7728a0779845256ef9e1ec9d0410e18122641cf1e2b572b
zb8f13bb94d46a6d8521736ec0afaf7cdd36a3923cc75c34f34da913448486722f4d7adf979880d
z3949db42c33a695484d7763ef04bce8423b10c48ee200c3bb24f4fd65880db7088ece1b884cf48
z23b8fb364dfac8fbe0a19a8f8f43fce423aa2574c7112da4ca7409ca09ee518b993e848dff2f2d
z78cbdc80fb2f154c811bf6116d4de0d7c64310759b3dfc0f476fcec031aac8b734b2451f5ca8ee
z480b2a0c7cff252fe84b3d5743208d3ec68b11bf6e54d094f046dfb9ece3afd5116d804e2e1199
z036a3d2990eeb7ec496cfcdd6b5bcf1315487322b0e487cfaae4707e1a1cc40bf914cd2ccdd3f7
zc6ef83a6eedc94161f0c6971f865a361685fc8269223cfff0cb9d7a3e16171399636d3870e3eb4
zfa7bb5b5f87a54dbf2ec8635ab3340992ad16492c394c57a1be0e12a3933ed04b239deb0e3812b
z309571c4c90b53bf8028ce98b1d6721a1d7c6e209d268dfcdce74a4a332e461306de65e9f4959c
z793992fa8e869b3f73c7670423a578a0087475d1b3d93840626ae31e3dcc79b4e84273061e4a3c
zc0373a7cf7120a92b56f348a8b3614c9fd9ff6a6dc9f86429951b9a3fc800054429ec6e06acc62
z578ed4489296de1811806f621dfb4b0e5e95ab46e95b9878faabde7662604e5e18a1d1e2da9194
z634105b0e1eb2ce7fec7431f72c04271b8bf6ea2fbecfcaac5619a72ffa08477596081d183b163
z944ca59dd563eecb0d05d01d23c6c89253ba0161eab7b5dab00786fd66141d9e61ce5aaa79e746
zd8e17ef4dbc9c82e68d5a6fb63678bc327543329cbb9bd13962635017ba2540cad79abf1173ffa
z78052062596ddb6cf67c8d64ad1801a991d4a41a22e174e2b35e6b537d65f9c6a10849654ed431
zed383b557d60e52b3e059db75fc7c4aaf06783ac687172ac2a669eafdcb1f359cda7a44f68decf
z22ace0ea904aad3949c6952d96960b6e4a19d99c2ccd265866aae4a87994da2ab0c5a5283b0415
z9c25413acf9c58adebc04abab0cff53c66fbb5bccfa4bc4fea3fb6e637c56db5d0e415eb638ed2
zf37e62db607395cc4e065aa06db8d7f24b374d44d67da591a89e6ec6d0609b0ae8ad8a15d945d4
z1e0c788c0ccff353e66a4b3dd531ec5f12707172cd8281c59d41e9ca60337bd26b2003887af58a
z007e12fc130f3c3faaa0de7b563ae791d6ba416499f525d8ecca782f93079ab9ac710464782ea9
z53700e2e334d941263c9736f50c2a9c317079881b80b91f45ecc5f50d704c4d2fd239445a0c89e
z90edc2fc54e0ff8ec441372e08d57e22f614e30df2ec0044154a25f0f79c1a7b25f7336afd2fe7
z6dc97d3949fefd416c4162a90b98bc96a665bb7cd896450cf4eee926363309f76044ed49e6bcaa
zdc1e85131ec5571e8d6c6bba2f781ebe903e29048a1710aac1baddaac54a1c4e16df5ed63c67f6
z5e974581a9c78eda33dc50254585a83500599f9c92d862a7c27bd6f879ebdbe2f58517dd2ca28b
zd06a16e465fc3d1a525f3ba62cb1dfff43b8cbf4ca75289b4816f7f17861af4e5785c8d9b2b555
z564f736691b49c27fee8b9b2f075b66386181896e7afae3402ea7ae7cf989f244a312723471e44
z6329283fef621b7c15c8e8d9981aa90526e6e2d0357be6b519a1ab0541e0eab7a607d6ffb227af
z33cb9a51b4ce8428ee93f1d6dfde8765c18a2453a293fc54e4ce79c58c608ed55490af4e0f8adc
z4dcfec867386cbf60e0e5b84c732705888119fd7373a5b08fb67f8aaea9879583e839a7d7cb2bc
zcbcfffe52fdd22b8d30c39d34e27dd6e47635d6c3f3d8dde300329777e4057707cdc5d17357c91
z2d0f49e8837e2544afc5198d244f7715b24c45df579f030955c816ab6132d02ef58ac86304afae
z3b64f796f19de8710295d58d78898e2097f573556ce8677090bfb3d7d1b3c0afe60f6303f8a30a
z8211f97c0ccf910c71b2b42de0ad22f7d2b94272da98185854d354007a331cab119d7434718f04
za10772d090d81aac19d29eb949449f55d97858841473c7ee65109c81b210a59347d0c252883b6a
z2c1e36c6cc94208657be5ba5a64e31878b1b5293c1c8cf6307ad152a83d36f5f0dd4ee2c6afe59
zca1fdc2dd46d76357f5a719ba7f443cccc64999d5a07719e2bbbc9d4e41a6747abb14b7a0aad42
z3b29fb0d4cda267016a109b6e2ba6973ec05e1d11801dd14757c9d48267ef555b38198fe67371a
z75124816770d3d0d38f2ca3452b40b7589649ef8182ea8d4a64c7a82c35caae9207dbb5542f553
z7ee4a6cd3d378107ca589c023b35d7f5f66fdca28e7328b5ab50d39343463602d8dee921cd872c
ze87751fa4b895627ac808a4bee5e56f4f849fdfd3196ca6fc64865f0f8f8db01dd6e19d83c2a8b
ze21b834d9669dea30b31ef372cbafcd29dad120a87c3a8c91f5ec38e6bdd71145396e50227ad39
z64ee6f606999c4d5d94dfc3e640d35c83de6d9f148d074bb1487247bbf810828aac93c9b1fc97f
z88e3319b690799b66bd848250f8fe83bd9dc57640517cb12296b96e81c2ac4bb9edd9ac212093a
z4921e342d335b5031091c891b2e73fa9a69b643332edde8b35a26f80283a4f541ff1b60332db7c
z0c6c2260ac40fda694a8e3863c64933f273ff63e7f4bc8537aa456de64b527a3a86fe0ec85290e
z4341855d56984bc9972bd58e25b9efab903e97aa96224368e561ea897e4b2c1b55479234bbd772
z8269073e76a0266ed9ba581d1d0873ac7b8c5c7d0f87e6030d214bf6e5a9c635bf95b477cd7076
z19f8673edd3864e4cd7cc44b2304dbaceb381452f4cebd6b5127c59800588be7d4d2c1c41e35d1
zdf301897b791e3fc5ec4108cb33b558674b4b7163414112bf08696c4058cfc4cfa69b41a35a25a
z3e4c06deb5532faaa907cb724026d137d1367913210eed92f2783c438cd64cad40e144660552ed
z04247e29b50161f7be4a0defd160beab9933ad588553ff127bdadbf8dfa22be0848b45300b2745
zc498526003897aed5939a68229c84f2cb0b96e67f325db537356efe201cd117e5e859193cb01fa
z28a04288e3c6cc77d54bc071d6e66aaebe90088ecc5de528fdce7fc7bdc1d82fc964eece91b9f6
zeda54a936adf53d9057d6e91941e841c705b4c3b43b8be59382f61277d69fd017567067fd935bc
z2cd61a52d56280d197f4d818b0219c523fb6bc2f7da349900ba19982c39af2ad740ec42955e2de
z0290f1db3ee00123ba21876609b0168e290d95f5639fd228d66a518477d1874dd58efcfae327dd
z196495e56f3e79af7741678f669366bef0a04163ef31a212822fa9653f242f1ae73cf3e3e61a04
zd5415fa85f877c1bb55e5d7860b6d7a9fc2bd0fb95c473f8a8f0eb79980527ad83131075a7df54
z651319eb3790a885b8a7a5c4fc10867d4b1cd76a408b7ce3619bb622b5c2f98e7a70c722a7dc68
zfcba80e0604a910c0eee443962645b8d2aed491019f155eb5108ee504a3efe329e737da1538cca
z8eccc8f4ea49ec109326a36afa5ad7594e5bf69f285201a6a97660ca63a3f957e81fd72c876dfb
z81571692a243917f2c05e7775457522d9b6cbf4aa56cd56d155f4dc81e2c7cb65b83e06241b34b
z335bbba0d2b832e146ffb86e4fc4a40f1966ac6d2b0c26b215cd08453cc3258783b77fd3854ad1
z689a7bdbd99fd5ea4135e5693b2a4b877c6bdea18de02972434700983cf996483c7a1b4a745a10
z1ff3a4a710d427dd95b02304f398a9e2d0bb11b76f5845a8daa860174a86b2fd24885831c987f6
zc06dc13befcb523dd7487b88a80535d39a9f2bf1c1374022044d84a284c4b08361950caa49658a
z37c30657eeb506f05171a5e16a5f56b65f06af53c4eb91f37f2fda31cb254b54443d3a7dd5a3c6
z88cac887262b13c2727d59675ff894ad882d788c0f63d6e338483efd72fd54e7bb9aa643addc01
z8c43934a20033c1375a13300df487f839cbd914794952ad0f0c5c75eea58a5ed5e536cfc832bbf
z1c0614d3310105b3c13edee98529489f94f27aa19dce7ebae3cf55dda18be0d0a2238e31a0abf5
z880aa548e8b181c37561660c3f292f31732ce00cef31a9d27d3090e5cadaee39970704f51d8531
zc17ff88b0d91f6bb00082e15c856b66d54e93c6f8b02ac65ace08c5fb4f679f7ab3a755f40f6d2
z070a42471c2e6b3ef02d3edffb720a8fdede40e7da4fdc9f8a048ff212e738799c0cf2d437a38b
z6e32b0edc95c5b3d4a0192d82f8fd964d00784c4e7a6d4ce530e1bb46c9d368611153f39f2f36a
zd017d124c1797577ab3607dd585904fbb5799b4c63b9319e0abd1b732aae62c197684a625895c3
z48d1143d1ee3b699a6922f4ae901a695bd230c6d1d52078a47484848198748938cd776a147fe2e
z4a03fae4979593ee96cce3be2d3b83a4d53f4630407d799179352e970988c4c60815dac65bc671
z1d1237005412d8c9d0ee52575b709f23e03ffd6bd510e6986f0813027b0a483eb1a77c604579dd
z2987e0b31a7ea1a85d60e7cdd747a06f754d4cb1bfa9f7a6537d480062ed57c37dd16cdde77a6e
z03c965622ba9cdf53b2cba73fcbd564c762da105c18813c59522a8274667cc79af8435f623b1f7
zac3adf88bc8bae52b12b34877d410cc7b3922aa0d04fbd1b626f084cf53c2a407116acc7f4c265
z72f2a75e7cf5bb8d473fe96fcc682b094fb7ab799a992226774dc1822a7c5c841b23b91f9fc26e
z3684bc64f751e282e6722a547201d6462ac66fb869273a611b4cbe2e76aea4585cfbd62f97289d
z5040ae0c968c16640937cb20fedc4a08a76d6d41778387748d0b6d33d3d3809266a7bd0a0e5890
zf6c132c67490ed0c15295256f7e72a4939130da26f6bb5be77085d0e4a4391f245a2f31d7c8db4
zf7f55335e7a52c8f14f4e47d9825ac6bf4f9e87d341bed9c194a1fcd45e4a8cccb38d66c98028d
zcacfd333af10abdd128cf5731b4a496a99623803a2cf86a4fa564b0e33a9f3674786c05676c310
z82556408dfdd36dd27fb14554ee96f2c93a8afa272c504cdf7ed7b93d4a7de409d1d5610327fb7
z4a9ad7ab1819d45ab5ec80e269377862d1b8f2c35811cb50bdb07eec5c2d6fad6d43e052d4c528
zf3a3b77af21659ab7b746d0a8ff7d0506001929b656e82dea3b2440cf340809a1afc68bc38917b
z778d8efb3c047a07b390b43cc3a30d599b3550f687d634fbb344e8508db3249bc425633ef0a7ce
z191c3e4bccbcfcb836f6c8f579083a04e05a7af7067e28f9a335fa5d8c2a77d31300afeb32a81e
z921fa9aaadc0b0a29e2833f8b53ee3d4df3973bd28e48e0d40d90ca07e0f193d23f7abc010fa19
z683f6bdeccfcbed5dc68584a7e4c23d5d36d0fd911c51816c725de9df59a48359b4909aed996de
zad6f455c36b1b2fa3b728daa603f7c034038b85acc8954470605e11dadffedf1858ebcb585f6c9
za5198118b489cb312171bdf94354324324d114ede07241e967e58f3c9e12df8c22544d88b72796
z0faabc9330d198ef4fdf1bdc5201b01ece54ed2da4ac8d63a376587a777d4d007d1908e61b846a
zbb1a9bffe9b0c205401d423c5357d5e9f1e624266fc0dfabb6ecf3a7cede54d53d5f4aac637ffa
z91a5285cea6aa21470bf66722abdbf02e7d09cb7452e54ea77c22c715e689178c1fa85aa596ca9
zfaf771d256be5388b3c35571529ba6926d5648b3eb87391fa36985da5bd20ef0ef2c4f80826eb8
z1c3ca11bc4228e66f5b79443390ad01bad0f7f887193723cdfa1f069ad347788039b32d60f8294
zda0b1bdb951500902401ee4b6dba5969db97c089281c8399ecf796cc9a794fc1da1b31aaf204df
z96a1f3ece6482dc0256b62a88587f16e2234fe08afd68ebf6725b3fe4648c13bbb22f71a018a64
zc3565dc318061dc37cdf27f50ac62b38fb60f4163eb75a31d16e7fc0cb58e9579bbd60c54b94bc
z2a1c8bc26ccd3ad7f183445f88cc89095569da9ca1c10d95b3c675eeeba94d1cf026534cac0da9
zd2df6af6bb96d864a1b728b47f7629059db37a7e548c059e99c3fe06992df6e35c5824689ca430
z4c54a1d1f1dab24162a5f119edbdef961572ec1f72629a54240099671c4a0bd35b387354bad404
z619ec3344d0678620dfb9410bead2c44d214d136ff4f2bd69805af96219b35cd7eacb5656c17bc
z82b94c07565431688d83dd0258ac92703fbef0d19ca083502db9dc4f3834209d8051fb376a7c1c
zbfbe1382b4e962dccfc116849f5e977e30cf9ba92b64724e0b3ec1d9dff31f5c68fc81c5509289
zea553be0f5ac97a5a8cbef0dad9ceaf41c889d048663d28ea14f6ba3d0b7a29427b5613cfff0db
z087c3c010c4f154d199e7759c4183a7c9b4cb0c738c751118df9dedd06e621351884adc9890355
z93248ad449964f3709307107ed3f05874b7d2007310610334f89995f2d4e02857b060c0613ce21
z00368cb74a1ee93db0e1ee9fa1b0cf0ee2584a583e5ab36ca31ae3a75065fe0f2425d237c2b1cc
z65e1154946fbae67ccebff0c43d205a091e916652c818a860c8e51ac4d38983e4b58fa5466ba3f
zf96f015107b035e41a70ac5ad0d0eafc40f5a333ec4852ba4ec7f106854c55aff3656e3b7860a9
zf431277c63df988fff05039b0f4546b0d3f9f964f6b0bec04bd0f8b33398122172b7a719a74eca
ze2b4fc3c160f921e998e88ca47fe499e6e27c8cf99c7aea07888a910c07b3f4aa24581c114a2a0
zd57e9d4f4deb20a989b9cd464ba139d148ab4dfbe3c7185ca42e4966edbc2bcdaeace4ed0e6fbd
zde3e33cc93eb331026f9a6ae42f4bad6c1c696bf9f1771c20ca8d282b60be7d6f1650239efab38
z0f2874f577dc17973de9d934d76edd01673849d610d2da02eaeca7466c16ebaf35781234f5c9c9
z2fff1bcedc2e8dfa502938fb664ca6aa1ba3997ba7056ba3843594fe58f00a3bee37657bcdcda1
zc5437b872da978a8f4cecb6367405fd69df0d62c8cc77fa364e3727bd046c92e85ca838c50268f
z17a8bd110a30f08fdb8b68363e197ae281989e7f70cc93adba764047fe5cc68cb7e5f3f02b8f5f
z88c0d4216a5a6649da71e7bc73295dac5e5790f2ec24692f4ac61b9e720d9154a32736943ada1d
z18b65f2f7e83ae044416c8b289e6ffeaa1c1d82c4d3eb464e96666fa6648bdcabce968b2cc391d
z3dcea2571d31cc2a1f2f1b55e5741e76074637b51c255564561f9d5a4147a794e273b1ece4fd87
z42de57fe813bec15d3d729a89e04243687839526fafc2485844edad679de1542379dbd3a6cee21
za8cdd39256564bff4abd77b31c8885e18a14333386b9a23891f6e317428e451dbc58e82ea7c906
zc7d8b967d0f6e507712428fabc6fbf1af61160cd66ebb6dcb2ed9f4892f6ba81f103af7264508c
z716596f00212219f8b92f6a2f43b551bd1d337c4ca1669c95ca99775ddd8d7e62aec218f4234b6
zc02b7c365f2aff0fd9812f6a58e3597fb19f0fa7ffe1e4586476941219783fe87a7a331ab07a45
z44bb06b9782d17ff4936ba596656413fafadeabe77b243f3f309b55b58ab0f8bd3f1694f455897
zffa7ef3249863288f8ce3fd2670a529625e7de63b667423906b30a2b95b17e7d87019c7764a542
z6d84db4a6c5d0967a0c47a074272e8c78a9b2c0da083f0a89993979676841e44d954fb245afa1f
z13a61791fad9614150e3d8f063e60aa8cfd4e8b3184dfeaccedeea4ce0fc1986dfe057e2b920e5
z02ab33fcd9d69648c92c5b60abea332d3fea76d4c196d9095305bf88cb5a83faebbe9fe276d36e
zc2668d3a12c9682487aaa1cf24b5bb80ef7e39b3c56ddff55a0562ae65c0058c860f1ec5ddbea2
z791af328b1696dc318bdef80099fe7295ca28d3792fd3891c6c13fe11a628b2bbd555b8d7e0e4c
z3ea366057790eb1a62b35febc2b1d946575f0bd432e22e4eb901d793fe2e05008593df82b09791
z40fc614904bc1fc05d081ee56fd43d5056c6331797a1a312fa49a771ba9f68b6c807a2a2500cf1
zf08406063a3662a887a04f62daa4535093ad93dab3564602aa9c27b42c922e7b409b48eb1a97de
ze5af60928534b27eac4188b6bb891dd2a6ae6aafa5e4d6edbd6eecab4a96924fb30116382ede4f
zb46acedf2bd47ea51e9f2d8c2980b1f95fa79d71a09d31479db40d2fb6094173cc7eacc6094dc9
z38cffb272fcbaeb063d09727db2067427fff31a8dde98c3d221a37b6cbc3767b01c4e777cc21fd
z712b83470042f92eca07b27ffa35219862c7d421284cdae5381add4e2e1f42e3ad6dc487812ffd
zf80b39a573a78085cd68e25d2dd6b36ea4e6ef054d3d84e5e53ad9b49a568bad6b28522f419a2c
zb76b4b9bade624aadb3c287513d5a2f53a4446afffe1478b4e4fc0a9c12a779a674030ab09d167
z9c68d61d58b5026324c18051f78cdb98614a295798a5b06934fe2adaadd093c9a318b1413d05c9
zf311b080ff2e82ff2796180e21ad0f681af87721442ee7362f3e7478f3ca8b70cef6ecee6e4c6d
z78136643accaba75bd0eaf2108c28cd3072447c3182d1260e1325233b48c82ccf9c087c55b043d
z6e87b6a43329257cf80467c9baf05c60ab4ffb9eedf010bbd5753cb511506a65c40980741a1434
zdb91061ff42d6ce0db2b19d835efd72121934309d819036dece851680b00c3cc347b893bf700ae
zd5f6afa6bfc23ddd0e8ba7c19fe667f5fc6ea4c47e3a3930f6a3b02ec47a2dc3a5367f4991452f
z8bc4cc8a7e7bac1494c961876b641154206363a42ecb7918292cc1b9c8c19ed266f48505bddf75
z7e1ea7632c078a6816a0144a79a637693cf804b4455789f556f02a1ba6c45c490888da1f9f2209
z5a8284616517e2262d7874b02db2ebf001b8fdca1d317951d8a760ee4f2bf86c4a463b25696994
z85761f2e3dc69fa8bf7e35bff4b28be44681da0f556ffa890b1a8caeabc582f5367f57ab25bcf5
z6d2f37667454e37adc9d6c16637f6e45699a9151fe6c57a7b3c48bb3b997537fc6a1392284aa74
z8955051e2d2a42482dd8b71e693143eca053b6f3e7dc25f10e611131457326aab0f5fe7118ef7d
z67746ea57d0ac8e49c609b15e427c0b07b8f6027ae70e5e3e3dab9319723d1b0802264d114b640
z06a21ed5c2727765fd638584262a62db2c9a8a997471386942fa779ccea8b62d0582f87aeaab08
z31c425d41f22f04777d6a467474af36784f274e12c18319f3977371cf47a33001e9cead554c49d
z4b934ab3f3aafb2bb9a8b8da23b0100057b832af76c1a39c2b5db66395146b1524828ca2546ea5
zce6e02606eadf7bf69af077c86a418bde9940a189fb586e61f9141766b60f179f5d48dd54eeca1
z98a2b916b6034501011fa4f0709248a31167b5b3d8fd10284bc7893914e471de32912c8b07fdf9
z10b8b1a39c57871f521e2596e2edcf286fed99619355f33fdca57796b41467161247d1665844c9
z40961291ad00d7dd383f7f094d8249d98284341db1e59eeb346a688230ba0a2274eb26b7edd7d7
za1d5a5c11aa6f5dfc28a395216084a8e386a1b8d3e86469a42226df5697e16d78c06b2d2acad09
zb3f7319b134fc67462092dee6b84c7bfae0e276ff590ca3cc11be96b7797cd9ad6faef22ada9ff
z18a688168e597d5ca19dc260352c610446c4184faf3280a99be727a11a896c57b13d1dcfe3e804
z4fa856ce3a8837d2fd4927ca60039016d23649b1bcd20b4094ae1ac40fb223a046da068fb6279b
z86a81e6b062c16875e7210481d1c9f367f376639d20751e1ecea9831629ba4f052a533ff9e24f2
z95731a6ebc98c2b8168ea8ed6c07ad0b76970abda3a2660e66448aafcecdf3d46f265f70164925
zd204c7a988b01ad6c8009749ae2eb0a0df35ef620d5797830ab351f1f53acc8c1dfeb4e2032066
zdfa519e3aeff5dbacab2ecdedf9d130ceb758aefc1800099c00052bc50f6d62367efe43f9489c8
z4603e2b3ea01f70f2686d2f3c0c802d9837999f4df6e145fc0dad074fe21967b49a16e5803e4f6
zd9dc393f0a420690910cf0be78b28b58d3631a4931363d00b40d7de5d6ad41fc004285966ff3c0
zcd33bb56176d5de3359cac93307c9e28235b6a432bf847ec27adddcaea9538bc26d142d8fb1fa2
z7fb6f703c49940f0264334f51fd292bf8f74d7429defddd32c5edfc7d518c3104e5dec6d74b8fe
z779b93185294d0c3d7850a5119bf99451ad9ba5a3a6a31a4941932dcec9224286587d48f81ea90
z7135ab84b677baa4978f04540125e9016a5c7b5ed39078a7b01cee52d6641674411c99b3cedb94
z75c0e4988a137dea68910553a9a4cda128176f0c53fe0ea232e4d9dc8201fd7adcb174b07bb06f
z45a4b38bc77a71304f53e90c5802d9af95269cce52e0ba09ada612addf119be9713e1c72ac223a
z8eb2f748f99aacbf813d425f79fc6d5f8f97ae43a4e1662370c3c969dec0ef10facd55b7aa0ccf
z9526797eb60c83e9fc40e3927de1c76c7ae4382982d6ebd5e15cbdc8f003a76a092e8d69fe5911
z5d25beefc2280d0ebb12487d4ecb0ee8b75a12dcd8ceb977975d674563c8cd773892b7cadfa676
z69c748daed0e4a04357286f949bd1ab5cb4c39a6bb0996674e794f252cd749bb97cb344215a7e7
z61fe10af8dbc05637794dc18b8cc2ef3a7776b8806293497f82ed75920cdf889e982c4448efcbf
z148853e7de99ca3f2963a706bc36b877c085a6cba3a899b816d47d70eb8bfb019b0a2b7e4e9c61
z26d610b23c5b0d4ace8e1be073a94ff226710a5925f0ca532c39041eb64402496689eb8989ab4e
z1e7bdd7a1d074592585226d7a8a7f54e890c16e6c4d8afc713fea5da6dec6cbc087da397c43f14
ze9f66695503726af595faa89754f4848e5863544ece1d1128efed42d6f5b9ece2081d7e4a21b9b
zda1306d937000d954e5f506ab92e569f721eb508042e3d772918d906eca6bed7163fc285ac5e2e
zb2d4cd0ffe2895e7f36aae8cf20e57a74d03920c4e1bb35c8da8f22264540e934797ecc7a86f48
z3b944604117029bdfbb330c6f2339fbb6e421a25bfd7ad8c1aafd13aae55f1a4943255217b0477
zb58442f65704deef8341ca0743255844037b0df606b7d15dc3bd3320c3480d6ae4cf74ef6aaf76
z97fb19b0866b7c3d58ad20980109826dafb812ac4c99a87f37233b63153b957ca0e1f67060b9ee
z5d0e3e40586a67c7da7c07f8baf0f3ba7b56688c756c05720f95acde155f470dc66b755ca0e3b5
z3f9ce175052c9002ca9f98d38124bfefbbfb7e7124b9393c1f51c5d36181e65f55d11f6e80e3f8
zdfc020952a18a1f571ed24e2a29f3a5cac3f6397bd70b98ba38965facff71bb37913812d307f33
z330b164d160d6027dc7caf02fc2a2ab2ffff1607ab604bd458636b42a6cbc5f4bac12c5b4cb5c1
z49c8dbea7b754fb6a74c839e3a824f9a2380643cd5c7703db3645825762bffcebc80cf7aec6174
za7f7c317bfe58c8d1732b3e1b35b68154e3058e0572b691164c5ec2e5c1a1a2077a4295f8123d0
z1fff418980e1673705fecf0c2297e6665b3e5179b6a18acba06da96f7899afe71831892bc37325
z2a3c9ea050437948e1fad79500c0d470793620986a9d3951193b87d260fe3c161c545dbbf273d4
zccafd18a021ce90e3fa783a5135d5cfd20f2839262268b8e000166216e1bc4e5be7b9016ee5517
z8a1021129284f1ac2653def18d0237dc4bafe0c66d126583cf34309af52467a5417a68432068a1
z662b0ad854f3c1afbe34711624396da6e9395dcbd4ca26985d57325d675d6970b4cdd36b081ce6
zdd03a323e3366b2aca788bbe0ec17223efb83f0a7cfdddafe671f1ef7e033bd75204ffd528e2f7
z4b08b9dc19966a62e759b58a4643fa440399f46717e253fd390965e1cfa299cd30fe56309a5043
z6164de5789baa546d6cfe0272fedf7d8dcf9aabc2a287f36fbdc86787812aee6108135bbe25f70
zc73dacc7c549c5cf2e7f326341292b19149380929e9c7830e8de9d9a7d6338d515355084b3f226
z2fa507b48e4ff6dd507cef277cd8cc91dbff607e8a6a88ecd014e4c8db3d7fb907779b02023799
zed8e67d722c7753dc6d07cd92289f89edf7b20dcfe45d9f8851729e3dd6c8e984d95a64a7024d1
z16d7c8d42dd44fbe1ed9f1e6208c7ac1c070f49d05e3063a948711e68734564663842a48d3bf1b
z3fd375a0a7e78fae7e007fd4ca79fbddac3efb60ecf791563c72daf90bf12229c0426b0fe97736
z938dbc0c7e2600326829609e5166fc2527c965f8eafa26b85642a6b334232ab7883b5133e70312
zf281c9c003c343e2f44da6f83371d83b80f6ea6b11fe7d15cc197b19f41d3bd1c39f84a6ab216b
z1540629bcf81dadc422eec5cdcfc5a2ab170147a03b5ab27c9edd3b3ab6d779fb793ff1e259131
z60871e8f0e1bfa7c72dc77aa80701c0546b3661c31d875bc9d3316104ef50780404554f647f155
z43aa5e1b37fb2ddc54dd32127f310aaadebddcbdf407dd4e0447d0e2234ecd5070fde8b903033d
z2afd9dfdb9c0a8ea3ec819f74e6aa83c7cbbc42c092a70f30dade006d7579e2c04ee07b8654752
z1f45943b171bc57a87f272438ffe61b7e352ed0e983c1139e9e9f22ff5ef7cab5d536228ff96ac
z924880be698873beb9d2ee6de6bef6c0aab4fcc334a042fcd31c6f2f14fbfebb88893cd14b5212
zafd16e75ead4111a38278bbc2bb0969de9b1ca57475030cda97a2ed92caea78458a3b214a35441
z5531c245c7c3415c6511fd4300702b17315d6df45a012c2a4b47d77a884aab2dd9e988f6ecb69b
zfdd199a0ec8758205dbe2d3b8c93f5cde0981ad0c8273ead46e99998b335d137ba2799f3007a0c
z70df0b04da2785edbbdfdc5027ecab4b3089fedf2e84aa46f56522c2105eb20ed7957c1e7ce933
z2ec3f7c6eaf18ddf6aa109ce7dc812b66d8ab62d2a5afda21a4a3511c5044aadeca73d13a53fdd
zd4fd1321dde1660acd453e878a9c55366383194894620bb34f9ea4a35c6af63209a68c5f99d45d
z090f187ac59f4ff22ea291e3e98cad01dd0894092be1a6040e58174c56ee810df285ade002f33d
zd76104e7637a286cf62ec1e48539049ac14c2a58f0836d8557b9f6dfbe0c2deb6ea7890ced77a1
z77ab9cfb9404f4bfbacad3a77e0a6659e9f3670e7b51e26ab57a1138022161f90a6ea067bd330d
zcff0fdefda70af0010dce1a5643297002e56f2af515b570a2a6faae711e0b09500f519817b73a9
z2c86fa071c31a7b59f7dacfce78315ef1e789a01f82f564d61328bce2f41f7f5a5a5a12194e284
z40c59d8cb0d14f8c4e468cc4ac9d8675c0e94780444a5466dea45e75e39203ae2c97b11dc24470
z32011829ed601244ff9526e6bf8b11229c5e2e532a6d7fe5cdab1a3df2cdb59121313d7e177beb
z9b162e935d9e951fa6d6f45457f2babec133453098a44dd4332dafb400fe3502ef541e4f39351d
z6c71f38687120d211f986b98d47158b987669da4497433d7f5843b528c81c0ff28a5ac596876a6
z60071f546b8df351b4036852f498757728ce00390849e0fb3421e8ea53d472337c17fbbf3027f7
ze5e45b7878d8720fb6c5cd7b13c30a7a84be9fd827583bc40f0a8ec75a7c3f2b6a8b3f7ae0bc68
z1fda14d5a6d698181b83f18ed1b80d24d9b1eddd6601b5c8a44e2349318a0f8c26e7098bd18cb6
z7796eca5ef729f6d11c0ec1b769d3ba767f06caabe3443f953c3f08f7845e5bb61b88ece41c23f
z21b36612399825ba3f39daa32475c83546be31984ebfd7b5fa97083922b4c25a5b5da40d00da63
z5f0bdd720c055391ee4ed7e4afc2303c69b85ffad9b46eb54e21ed816891cff7b32e1a2f627909
z9eb87857a84a43c2ff01485f9b2559f560ed8765ddc0a66862fba2770cf8328459e7fbc66fc1e0
z48c962d68306d9d56718f9ef145e744f428614426ae4281fb76973246149151cb94abf169b6000
z87a9b79f1248323252bafadd93c8640c6170324d89456e263b6d6c7838c3a970684aac6b3de724
z950c368970ffe3c50cfdd82018ddcb02b3715a6bd1093fb8cec4c0f99573bb9e288349e0d884e1
z2532e51bab6225f7a9766aa49d8d7fed4c5bfdd98aba2ae62d19f74ac521313d758eefbcf6d1bf
z53209cea0b684c71adf55693cde51eeb27cce31cd56058f4e7478001f405965e2cf4a7e9d7caba
zefe43a5f409ccb97f50e3fbdc8537975bd493c9e0210ae12204da08d523df2aa22e306c1c8bcea
z41e880d214bf9a5c118a5ff66eb95ad6a29759ee6685b127edd913fd393762f60e5b874f36927d
zdfc84238c98fec7912871ec9d7f9f567352d6f0768ed4bc09faf78fd5389902a90a0919950a17c
z7391d4b039b109e1390ef01f363b0dc768418389319478eddea090a0a9a68fb0f96ebbbf997fa0
zba280168f08670cd1727496b8e2a975e56fadda775a928a3bdd48fee10814b08cde5cc040d3fc2
z7092ef21e40b9c8f6a34d52f5c259b122293486904e31e23a47051adac7e9276be53104b7a49df
z4e996faac1fa2cc098d4f48e6375ca2ebd282cef0916fd6ae1ae8752f4dd6916cb49b0b30a6d4a
z869f9b3421e40e9f5f9602cf19d08bd73350a3f2c373fae138d0d88410eac82be141ab3036d752
zff07ab296c51b4e400b16ca66b27493979ff349f4e59357236d08e2c4af72d7f86e30cc4d6dc12
zd3de512bb07f0ebe123815bbf83ee3ab608ec149d80f0604239f22de67ee5d0e90e51d5d7d8a32
z610723134eac85fbe325463e72c66b71949f2c06b542f3ce1f425977fdc52a9c7110a9bd015d07
z3e5d41edd0fc154df4584889b3f839fe3d47f054e6e3b42cc8b838939ac8517afaa0c832143d34
z620eeab87ebe7ddeb919b094fe84d67f79370c4cb3095d157b8be6b8d59fcbbd3d904e5f9ab692
zd92ac68b69232971427c0302cdbcca5a5e35f5e75d7ec2017baa7f78dba02e150f84b28a6d825f
z1e9c768edc3d15de79df91522718db4922cb920d0189f1978646d63c057d52f159601aa1e2d37c
z14c538b3474ab3bccd54761737495317fce78aa46c079800a1dcf41b9ead159f5cbb8a43a630f9
z72dd17de2320dbe4f9b0004f69eadd587eb5d74e6cd0cc81de97f386d354660391dcca73aa0a06
z7e5deea3448eeb4cbe38358f0445499e5fd23ed7d3ca99fcbce828bee68fe66ec4a9f178522a39
ze1108d08683a36df802091757686f4b7bb27c0c3e6f22de0b56aa757f03c2dba03cce6495b60ef
zcc02fdfe4b758ca1c78689dbf1ae8b4cf8b671defd5c1b2eedce689d9754e1362085db615cab81
z512e697c9b8529984d7a4d906ea2a5cf9c4e132a57b896f15c1760c9fad93afab09faec52c3fa3
zcf1934270dd02c12ca9953fa97e791f66205eb9c143ed7256b3b5347e1c3a1aa0d38e32db05889
zf6051ac18d997af0d19e3205e917a909f307962dec4eb0e97ac756d0f894fa85876cff89b54a9f
zc0a8b680219234cbe2f6d11941b12773fc736d0336dd49a7acaa44fb2d250b5736cd6266a43dea
zbd03e28811b16ef43eaf29e7e0a20219b5d3aa0eaf39c0da0434d12287d93294ac799ebbdf71da
z26c4be3bbabb7efd49e3e70c78d12f4f135f2374fccc1428263580963f56cc1d403f3c74f360c6
zf738f42492e0b4de8da7527c1869e9d00ef0f123400cd6c90639d6718b8339f365c87df0fd7dde
za2a66d15e79cf2fedfb0b465f26be2f6153cd81c8926a1ba0ca2a0b2191606948a77c2c03a117b
zea83c343e98d11b7f544cf139f87fec0b08486b31d04806b21ead7829d0de06a29c6525dc188cf
z7a37b2353e4c4147567ace842b7b0691f645fc9456ba299e51d29d59fdaefd58c1114a737818b7
zbbce49f22b97f93d1dd5babcc46b44c4d096c9134ec873a1ee0c855049b82bbb289c5483cab81b
z2db4cca24cfb367c523f4d7f150cc5c977618e2b0ed72d91546e31bde9d52102c57c92f7902ffd
z615fb7fd7d8b039a93594f3e14d8822a8f9f4ea4024cdfaf956aa204faca034f10952527cd94cb
z8033fe7e37d2585408a1f56cb5103b0f0d403811e03c490c29f1a1cd686ccb98dec9bf2c94e993
z3b7ec83accc08fe29acc36002dc98baf914c778447cbeb64efaafa4b48f7d170b33bc15a88e2e7
z712c61b895055addbc9bebd711b35f873d5771b825e26241653d3569ff60d3a283b1f027150224
zfa0c15b6a52f2be747f97e83f7f5ddcc73f455b441bf9edd21c40135d54f8827a81338a682dc32
z0818b8f3d6e8d53f8c32845ce91b0b4c05f76070eb50c5773d184684949b7a3125b6912308291b
z7c5203aacd341621fb89b1568b1f3fb8db7cb7d4919f8e55e6986e683a92c88f44c32c2f591345
z66e47f1e5b047c420e4815455b5360be2f6a7f812d1068a0a35c21b65c997d077c3d6361812284
z9605ca7e6ad1db8c37c36b6860525aad5537e9591eac35fb71c07015261372c598310a6a73e371
zd181ea56bafebe9d297f2411319cdc4680caba7c625b1abd61ff4cfa74a43eb210c84adbed695b
zce901ba4ebe27162804bc633765d434f87f0e247bbbd526942f0af53dac2573aaf395067367415
z53f04535daac171373095dcd646a6a947471e83ada6537f3564056523479bfba795d3830af7f46
z316f850d09754cba39f603525a3f5d22b8dae53816ed3e23ca1713e3b9839b0b08dd76d5c2c60f
zda88552a0484c6628dc31035d7fbf6767c40a0d22866cee9fa19d3024d32ae04b070c21d880c28
zb259f227b3c53a7a36c8aeadd3d11b2c5986c72e778bb468e6991871b029f8056c25ac2593ad9d
zcdb15edfad6992f72952b39435f9922c1d436314f6e2c20e702ca938610230c1a1aab35ed19603
z6033695526ec51330706b229aa216258f6be21f9cac1b8debbf71bbecf02cabb0e75b9fc0f32ad
zd4185924d74b2bd9bd794b1b183bdf56b1e2a247874264e2a1e100983ca60cbad0b43c54bca9b2
zd9e7c992b25eb31886be0d9785d72a82bd4d8a69b0a477f653fc4c765646eaa1122e377d220a82
ze9e72e7d186aaa76c7d5b318553e58bf3ddff6e3cb781372a36856e0cbe62da8f391e6dff0261e
z0d5608a704577733a996b0ac687da9f4f4c799cbb0fb794d513492cbf164c1cf023fd22fe4d09b
z3dd7e4eedfd076129ce0229037a0d0def343bf3b86341948b94564fc7952aa35bb17ae76108b3f
z6287b97d901a874881b7717b9f9b64b1ebc775c74a9b4fd9c3b9b5dac6448a0f1a3590e8a7e282
za67a3edd4f71e74af537ea7ab15d870f5d09758a5970f017ab8cdb1dfae91774e2c6cb3cc2aa3e
z42bc1b877d6162801ce3dfbca848f538093ac7653501326a9663a42c5731f0e3d3579ff1a4a239
zccc183d96591268803bb4ddddf373fcfba994a063192dbfb2dac1c6f940bfad9871061e6438c65
zbe1eb4041ae9969bce4e3620f2dc1eac71b6848f10763aa74b81fd48775427341848d7757aa5d6
zb7c4d0e145ae21370cd8ea63f95f9724f64f116cf1f527ebdcbe2bc69d5d85a10e0ca3c0839e48
z7be72fd0c437f20b9ddc3ad52e23a1e7177bc51f4eba0d63486b97a824b21db1aad0c204c1c9ca
z86a86fb4da43d99545a8809da0c4341c68024f621292536ad47ebd8627b1be1ba3ae784294fc97
zbf311d305bbf84baad1fb8e9c6a264b19be1af40538c74bc9548011a03362e5f9d1aa74867d9c3
z7bab0fb215d648a413b5d9b4fec04258ae55e1ae9dd790c9d403171bcc33a8a8b9db64dbe0dfa3
zad493c659d166da59bf9047a3ac6fd05f36f9f28099e15ea58cca5d265777d56e4ca004b57cb22
z041713984a182550e016bc170ccfbfa9f24b326f414c4330202762b59294fbdba6b461a098f78a
zd2698ac7762d42e0c892c4a29b1bc4a0a87ffd9490d07bccfcc9ce3c303abe634671aab126a7a6
zef8e3fc9892a886491f9a3f61765ace08f1325437b67be2e66ceace56b7e80e1193041005c537c
z1e9053aaf2fb0c9656bb8333fc93d8627885cabe991a314ddfad871bb9e0a336320688c0972915
zdc6daa72fa8e25e3926a6656467d14e867594f391c4588e7543ed8f226d975fba4a112148362c4
z581c6fbdf6f012e2d301fb59d8d178941e593a98d188362e4539ed7bb0188be953247caf43d778
z7b347882ffa4414f2768d5a4418b6e47dc38aa17ec0057e31bf8830af4e4c7e728cc74994f7f84
z658eb78569bc935ed6854405c15c4c632217e5708b2277d8a963b574c55dbc21b45da2551b01e2
zcd1387a711cca1cd2eb0aac8aa5e30c6f32f65ee50b634926c84900384e16c1ba42832813ef29f
z78ce174e63bbc88b633123deb652ff61acfdcffdbffdab0f4f7da9fc7603dfeb9e9a9f892019b5
ze606e459298e8b4c7714792c450ec0904799dd149f9a1593d8d37a06d2d144d434ed13035ef7e4
z1334b51a7076eec31ea418315e98f2cc12ff0f2cffdefca8797d39579cafb1a00e9c58b3bfb024
ze01844494bba1732996ac240b7d131e5b17d6659f48fccdba08c5a49550946a2a8d69f3bdba3d5
z3b16d9c4389cebd94f2378b981b519d301ee97628b271c119556a6313c9da019501672b24594e9
ze32e5763a9eca4fb61c9dd7ad0a0c52c2134874c6a15d1e59cd4590d251052f25e14fc4db38cec
z1600f7e6e806d9d7daa913dd73076dca98b1ed9b05954a0d1e32304664cd518adfbd1e11dcceea
zeef0155fc02aac7965fd5d0f834fde86c74bfeaed3a3fd2d5576ded959bf7ece77e6e0d0c2158a
za0ba7240a411b1ebfb5e99d056cd545b2aa29678aabd6f5836137abacb44010f7d2d0c87c05071
zc26bad93d436919b5f9c214a3928c76e6f870577fe18cfc9fb1d86b843c99b8929daa385064d24
zc0ad79959acc56b6403825797168f7897564b36a020aea85b149fc59bd3f373e1d2d17c29c60c7
zb32cfbdf6320d98be2680425c5ba7e2cde3cb8fb60a19a81587edfffafbb68728c3dee15e18f78
zb7b5d25bba6146fdf36bb95e56012e3bcd31fa380ddba7ffbde6af17c5f9657cb59d6ed6b1e53f
z34ee2c6af3d90730be670976471f44ace44a2260bd88b4680dacaedfce5f579e9265ddcf62f97f
z3d1e7d9d29704b1433dc4372fe1f0778d3d1e1bbf7ccb6c40de146f463179a93a572201e76ff2c
z46092232def0beea21262516367c1abe7c91cb4c231ac4833bc97ed2e0091c0548fdc827e181d1
zdd6edb8ccff3c99ba38c7ccb6a2471a70ced1ad2ec12ca34febabedd75992107ae46169400df83
z2e8baba1a833edaac52efd0af89f2396d46add6be056142f20e4f830c0f581c24a273d70be0259
zbd77142772577f58fd16f83f25c16ff8178119426b0fe1db9fa740482640cd774af2ed04e3f925
z9ef6a907e5dd0a1f96fed20645600679cba55aeab0b080e81c89158f324af0d1a56c05e459f3f5
zf2da2c8452cd13f2fbd74ffac47284ea25005a9f5124b138345c5dd32472a088202c4c0e6e25d8
z41fe6d047b6eefc928db2db8f832329c9a3e9fed84d165cdc182a64d624c5e856da535b43289c0
ze11a7a8751d1edd972ea1e2d2e7bd7e44097109c6e4d4dbef1c1683fd4087afdef1c90ff2953ed
z57d761271b1cd3b254dc992c04b57a939e39d3dcad8f090f0dd638767b4c45c39ba7ef150d22aa
zbbf4bd0ba23f08f41fc3c952f72124147697ff1ee92ac6d932de055c073e10db4c8629e8575fe8
z482e1fb61cf33cdc0ffc380114f018e8c93b0c38ea75be3b32bc26186e0715aca79481ffe8a0e2
z36deb9ae3cb9330f2cec23fa15932b4d2b2cde1852622c6398f157f24663223fad84a9178aab43
zde4ded8ce0115df3fb05e0babedb3d2c1fa31849149cc3389424f4df368eab8c0762eb563e6a5d
z54888fe6bdbc7dcc765544973fe2f21c6fb552a6ea2237f3dc0c5914c2d71cb0ea358cf55923fc
zbf9dcac55084a95ec5f260925d799e1b4b6d2c80c21fe46a9a3a825bc55699c26cb8d965311c25
z97bb6c8dc41544a319a1b0c720e98d743a057590f1153e12865921587649ec4d18f38969efbfb5
z8a3e72fd57575fc8987d38fe4a386c60643213a7035e4b946609303c1747c7214a9bab473cecbf
z99c84546eeb9b46a218555ac010b43b630d5906c6e290745a4baaf4646741b412be4a11fc6ce48
z64f90e2ac7f41242539c882e598be90e8a8d3969cc6049da65b6b33b22f266689f11d0de6434f6
z9ba0002e6a45d82f441d409561192e594b69ae8b8dee521448badf99b192778180b1df3a08ad11
z8cde043ae24690ff447abb240be6a7b8ac9af2d40e08cc514a07e2ec893d9610d66608c0109e27
z8966b6a951915df9b1c7727db7762b02ac93028fc13116361e96e48a51daf12c9e3ab0f0c21183
z1a8b501501a6de6deca5d8a53a3643c547e44028aa4d595b01b1f4b0e398df7fe8ff94a89379d4
za4f62375fec55146a698b9169dbb21a993a07e8ae82d1284b10b062b0f5c2a74d90a39328e4881
zad2cb0a8cea42367cc4b9e989dcc8e2f231de8b629ed857e21b31b6c21679105c6aa86b24ee5eb
zef8c514596596995de87174ecb13f923c7e391819eed3ac3c30e9dbddaaeb51187b6a0e76e7505
z63e09484d649f954a4dff827f57c600da6b29300f129957a0c24e480879d764bdc937a5af9d588
ze89d74479adc8b21b3e78a33c3d02ceac5eb381beed26f53ebeb2e48acd914c5e5acc19753cab9
zdaf5bf73541a4293913267817d0dfb4f2a109df32339dbc0bc246bb431a1be2287187c225b8e5b
zc61fbd673b37d80338563c49491ef8a0fc03c02e3969e627ef702a867554ebe9f0c5f13911a408
z7628584717eaaf0c7e0e4abb485f99d7f75de295b840f4a108e854bb84a41bf4b42a36dba59b69
z89a73625b7f087a8218904ad5ef1b1b7ac48eb6d78228271c34a050a2af7ba5cac5a3fdb989aa4
z529fc0803387d8f02f3c997833f5923d4ab419e6509f1d13382b7d17f74064c9a43c6bf0166c70
z195a324035c147dc54d51336eaff5615679b437f44e3e671f9f3ed078385cd0e3187daf95d9724
z257f66afcd0a0df4517b890746cebf74935273beb7a11d08d9a0fd86e1790887f19227a21482d7
z3ed92e2d0757a4331d6b6590f29be92b2a62e340aef6f942e255cf161b04ce0e7ba4102acaa2a5
z801a815e410cc1cab758fa7f23a752294de7db5e52dc8d43726a3992a4a4787da240a6a1923f18
z65706bb2b9b93c05a0eea35d3478609a7b1289540272c85dbf3a7126e8ada6dd4ab5a9b65a1bde
z70eed77d2dee448acb47d2059a76fc3eb33c9eabe346e9a25d8e3fc3cbebabd47d12a3b467bc39
z4107476e4b6439b6b37400dde8a24ecf5930a8cd7cdfbd65bce6ceee2fcb12117729507a652ff1
zaf8500e76b6977e1c6effe3d82ba31d24ea2c1e261d557e1d9b2a50ac49e55be0acb98cf2a191b
z72d26f0fec5aa68089e7b8c249d85bdfbd5864cf8b89e514e4435d6f42395fe5575fe54a485044
z0540c24c97fa2ddc03ff6e981e53def460a3a70a35f6d25a7d518b3904434e0b426d7c59c27b6a
zbe330fc11422c519424845ffb975de0b7a4c1cfcdbfa6434cee796c70f2981b3561c48238b6db2
zb60aac564b7b9c2aa416cbd911f3e60e4031b3c5b8401e54be2f762a1b7db5d0a7c7a589f736f6
z8e567e82ee159e353b0159d60e87f1d6faafe6f37d4b57e86f0f3c6bfcaa2625dd5cce13fea8b0
z10d1a0061d2bd668534549fe8ed2d3204dc7822b5a2e4a68ac04d207cdab818e51ecd4bf53d8d2
z3ef2518259ab380217970742c86b65fde3a28210e49d6beeb17c93f870f75214fb89fb5d083af3
z198d55c7315a0432f13d529e28cd4ab05791883f29e2b46ed191ba18b82635dc63b9e1a0516664
zcbfd365c2177dc06f48b028e9fed138d1e1e3b39c0a63f416450c9d7123c36a7271e23137a85b8
zb0116e64688a2ce01ef6cb93cc1a75d5c80c557942fa3345c5eee335c5313ab52c1530861cdd29
zac1eaac6142c5ab633ccb32c5e412e10f7acf2754bea99ca82827d011f74134a59db93505a0d00
z043b90555d8cba88946f8462360a8a3460cc91f6ceb812829af1d1361b9ee7530de6ad10eb1537
z3fcb8d6245418d372fd3e67989bb4eb32ea1711748db0ae784ad720a8f52d2e8dfa80dae4fb5b8
z1213a46f3cd49b43cd82eb65013b3be7482f244442151861d21c85a876b2b5c0c065d50d7d0776
z819af511750ce690c4965d9f1ec6da66bec86c33dcf0bec8fc096a3b11cbb0253625a648596dfb
z4334e2303e0352503407f539b457ceda16c17605bb7e73db384ebe437fa6bfcb25f31c3996d2ea
z0700e3c4a26deaa60ad076e91e29a65196e65fbacebe523ff82c033551f2fce3481e46475eb548
z1a7479889ff56f9961e79a2d0142fa13991cad59be0981fd7fa288bece2b0921e7b74f3290e662
z25210eef1c89011c02bd6b747045416aedb912161de5e2849e2af7403c49d56e77ec6cf2c69ea8
z7fa2385a6d12a7d76222150196ac5a2a82d783690c18d8b7f75691ca8697fb05ec50c70ac350ef
z504f0120f2b4a819ea96ac45f07511b0f2411834f1d190cf8659d6d9b83bc7cb2bc086c372db94
z2a99538a1b91317cf598490af329e3b0e28f082f9138fb6ab79932e5a820c19a495fc492c74696
z263e17a80d195c78a6070e26bd62afca3bfb9891baf716bddb194bd893d3657131f8b73368d4b6
z1eb9d6516c8291c4c6351308c60c4dd2112359e208d180e1a274466aac7a0141a0621edc47fb39
zfae672145eeb04954fe12128443abbda578af38db7abcd67f91da80f23eaaff70671aeb6aab262
zf7aa5fd32f58b6321d03e9b3ea9e5a1d7322e1b7a71d1b68c44b93a09ab5e7b4513bc538b22d69
z58eeb3f2df89dc6de81adfed8840a8186395b6865f0eb2be4a7ffb8afcd6153ff908bbdd094dc2
zd4c680a290bbfc538e0ebe04f46c5f2423d28a6f9f6ea23c9bf5a4fc026f7095fc3a657d9f6499
z6b0bab1858ac7aa572ca6688a4ec2a1a922586d91ab15679097e61b3edd833ebaf7f05366de5c4
zf081ca495043d0a94f94597195b3496e32b22e1aac143e33928e5a22f170533f7568c939b4ed7d
z5108cf7192e93df42f6d68147f8d6ea1f874f41ca01ac1695b29e53e48c0a1ceba61047c483b85
zd761516956d835451b1685ceaa654e0e9814467921cf8e62fdd97a8560794f70d699117a5839d0
zf483a518755a6593956c1bfbc5f9fbf2f4b3ca51175da01903a5b777c15cd8c5aee06baa65c20f
ze473f2017e1913451d65cc3706e3a6fc8d20d319d651760e17f11687e906c7f7de40acc838bd42
zc01bb49b07ff4e2fcc01cea0e3f54a320740b7fc3431ab009654ef731de766791757288daad0d9
zbcf6b5342920d69e37355002e0a76b1e6a04eb7ebd242724faa00388a7b08645e041634b57a0e3
z4050c239387959545089e6680b0483be53ac23e14698bd61ed93e4080564c4940febc2d90a94de
zc7a7981cafd95ef2a7af775d0debfe1f7215d11299dce855d1a49268f400f594413de5ae0d79fc
zcc0b1c934a3535a202eb68aa681460e3bb6b2e1eff59bdcd77f7f15c8b6c55fbbffb2b150b8179
z07107502130f30d7d249680d229e0445082c3b433ed1001480a33e518b14a91e880f6061f458a2
zadd29ac3b96b71fb252a99bd4fadf5fed8939af3507b22787bbd88612a2baeb19529694006ff1b
zb9c3859c65b5204a58b9908021a41684689f231e6f415e343487e643731d5ff2420295103aff27
z2f781269b22f991ef3f17a75049658b200337dab183833c4558f53bb28fd572bd8b463b4dc3f77
zf450e72b22fa74b5dc4b49e1c690a824090c1aa85a7c9526597257de9cfc3b227aa3d60e5c2094
z19a6173f48406c20eed48cc2a4fe2494200d4e20c9fe669f3e38d5a26006f9f2df85627a380498
z0c06b809a20a75862918460244a7db11d92ec9222ddb4d95486cb400d901418b2031ac1287c8e7
zac214dd36f93e2ba560d3590c7c77f90ddb439b868e4d46804552771ed36a9a72770e7b81779c4
zd6fb36959e8a855a47c972cf6210f65fd872cf6311aeb1ec4274aba7d6b379ec0a89ab2e55633c
z64882c8e05d7769a3a10735e556a71520bc3929bf4e0e553cf586c2d326e9fdadc73a00d2fc458
z40cd3c56988139287463696f9a56b7bc0495dc5822d1b854b49e07bdbfc0a6433066c145d344f8
zff35743dbc932800949d9fde8dbcea3eb2636c93d4549968b2156c7b3da1d3b07537880c7eb69f
z66fc86a65f8214af5ac5032b4d33677a8cb959fe4753b055211bd5c9ee14a4d25fe925f645aec2
z8695e9b66ac5ba7289bf29e1e2cb0d04e70963b451602983029aec1cd0c65f711ba43757f9a7be
z2ebd613664705ff03f8552888de0f5b90ba46be0a49844f103b4139c0fa3391ba1b5281a854003
zc7f742008b6f2b0d714acb14d85d87489258f18cdd383f164949915e15abf8933457bcd9649668
zca83f89e6d9abfb307827c3cc920f43277dcb2a825454cd1078be894ff6f9b9751f89be77167a3
zab25efd4c816e355a24904f637c1e3eec0b0a734e4b6467aabc30fcda0906981424dc7347ccf89
z27b2c4617775e787b07b17c890dbeb233c1a3c5f42d5e078f8c3df93ab7cf6236a846a49b5e76b
ze4a3a2eaeaa048f790441e2139f439291146dc651fc3c3474186c196eaaf5901b066f3f6000870
z1ecc1c9428fa620fe7e821934d873d09a600c4f83d3e32fa4dee535e5d9e9dd19b9ed6c892239f
ze348ff5f73d0ea3c0d3bf322b297d25b651f605f79f9c227c5c58e2b73e16bc07247bb46954542
zff8b81cff65fa5c71ddafe6bf032f2a2103b4a40e50d543eebf4e7cb28fa967cea31338c6cc191
z88c555ccc2d1deea08eb9699dfa88588d776be28746632e8d2b61023ef137dc65593d5464a6590
zdcf3be0524d60284d3a3acfb8cc1148d83c07dce7d9a83833379a58c02ab1300386603bbd80085
zac95aefe026bc9d446309c1b74ebd49c1c4911082cfe213665174130dc339bff48eb0e855577ae
z847de82944409681a5f8649bcd42de00fff8eb4c0b015f31d377a0f692d5191a038f3b99505867
zb5ccfff6a45817cf0fa3b54414b97584c7928cb9f2050b45011d01143a6082680479afc86834e6
z8f890800ca64eb63c5a35ee884fd84321a5611eab0a4e1e7ea16e4c1964e5141e8f35f7d33009a
z6666e3a5a3f4cb5cb6e1157bc21f3b76394bdbc5594bcc4be087032f188813096b3c4f3999f8bb
z0809c782859d4f71b82ccd2cc74080757ab11ea4e020fa62fff0b1477319af2174d4861c55077e
z341dca55e3e6b35b062c23fb28c19961b5c33f214e92253c06dff71bf19548840f34e30bcd765d
zc667e9711ef142bd3b0b87f7b3bc643c464d35c1f73d99cd1e21c834166a5076d981e6c5a7cfc5
z1463e706d0fde24a0f2f733c5a9ed04d39c421ee40895d106d737bc1ffecfa81fd87b0998fd3cc
zf9d0ac408c200c858d3a85ec7efd72dc8fccc0e3eaf7527d38f0ce6d5481c24d54b7e04ce8bb0f
z25ab03118cf972974e042c1a992a0da909671d5b9b72d75726f13954a71379f96fc34e5c1d8339
z76e0b6b3a84fc19b6ba875a4014b79ec91e43d522a23c6172c868a2ab5c381fd6464cf677fc8d1
z7ee94b7c9ca7ed1e5e17447b5d81434c371406b54c73078e288e5745619ea12e8d1c330a5cc1ea
z11e3082690b66dda176dc8cdcb825e10b4a2954677e11e63238134c233131321d18e18c42e08b4
z9c2ffa2793267580df52e1e4c1b94186389c70d045a118d5f159464944bd9b85403eb1174d9ee1
zdb4c9ab143cb697331038afbe251b44c9f323621f0a2a6014f0797e65638537389946f168d1e92
z9cb0feb81df5ec41c71e037c5024bcaf8ea5f5c8f9686c3df64622054a54653b168fc8e5454e81
z5b14b7b5457a372db671b4f480f07cebe23dd3a390e070f0686b8558224ed62491d4242ef9983a
z5da6f4131f4908a1cd568af8613277bfd0523769ed21e3c245b47306c00d89f58d8c4e2c4819c0
zb19ba7d81c20f906b45c33743763b463b0418927551f6d559856b806f8b374dec134e6c9812cd9
za066d96c7b28ee779453e322e535a94709e980d9c61bec9464fa96968bb2610187c7cd4df35767
zdff8beb8e5a24a05e6eb9983250b8dfbe7547463690957c8be5a01f69cdc3eafe15553b3ab4944
z047277bae742925f64c82c1b2ff8286944f724096b1db5bd3f6c5881f7a1eaaf1df9eb6763182a
zbb5a150f12dae917454d19f9e75d3f998b07122fb30b33c344199105cf65e5b4486485041f382b
z92805c1579b68b408095101103f12b389b745846076f9f05bccae4bf4e044011cf1bc7a7b5f337
z94e7295b84821a1912a22ac38267befe94dd78cb8d432e72f97a288e785ae7e5c12275cd4f6654
zb60420dca7f2f7e9b73fec896bb2287963cd4deebf355940c558157157a317e09fbe8a4f461ccc
zf254b4a957ccd4e63f1ed1285ab5c394c755e54b9e2968756a8d76f5105dfadd1855b6d66ec38d
z245e29f88de0de4c9161a5896c9c0387ad7480d48e8835845de53c8fd2de61255d93bd8e06b338
z04f35f4f81184c32d95b64a65a14c2f744bf2571103c09c756ca6a7875761fac5be8e0ea2ebfed
z816e5e9510c87c879c2bcd8231b80f3c247ecea9bab2cab51a6891acfb67c29becc7de730976aa
zcda67255af7d23adeab4925ba0ad4ff30c2607daba8624f0a429588aeb2558bd1c99b96b513955
za9286fb7bc434865757ec54e5ea5c735ce42a3cb7d20d9f4b9acdcc9ead3f08cbcde4cd37dc873
zf7e47eba5b401134c934e6b7ed6519a5be1553ef67037616c9fef9ed5099ad1e76ae97f85c61d3
zf9fd2481d7ac2c5dd7118a4ec6f55e248d517ea8b99baa2824b8e7be7521ec550dd19181593c35
z1b7f384a8852406e4ac2cdf3305ce8d1daaaa9190a3a3afd048b1d8f83976310cf121931b9017f
z490be54029825fc4afec14f19e6cd3704ebcb5c2e893d35491d8fe54d76e2e92b6c4a9e9ae2aef
za3a19aebab65f7e381f08f79a15cd948b0c45f80b85279a2b96652b4ceff44fe65c5711b4c49ab
z278d0c2ff152aa3a3c74c12cfb76f4685e3c4e987eb85e4ba69f944891f990fff02357e472bc91
z1a8db8b2d3d94e282d6367a77ee7218177f2aa88643e2a01a11016ecfdbe58e7697ebfedeff858
zd462644d379693c213def72118d58c342aa2cff511a428b7731aec38a2b04de6bc523d56a5d5dd
z6a5449163ab1943c8140cfdb15438e320e7d993d4390979d0cde278f1e2221b4d6bbb0238064bd
za1092d337d0d9f659bda52bea7bd7dfdef253bf23ed04b1c27f51ddf67d065cf08bbef6bfa1418
z89b97381f8dba403a846368ee7615cc7381bc5e74b74f744f5e13c712865aa7d8cdc74d2dde844
z205a44b6f92bfad1633e3381f161548c07b15325e220653a235168f832118871f4da5a3e6eccff
z9aa7502a59bafcaf71451945667f6d0c0d9fa03d6a44bc476840ad1a8ec48ff44b7d31a4337158
z5dbb376a18aa11c5703b24e9241db82176a4851ee3c0091fdf83fc8fb6ba60a3deba6f0317c761
z2ab54034f722691f8a01799219c1141c87fdc016aeb4f3322760e2c68c0b26bdd3ae8135fd989f
zfbafd0cec62479b460063486ef4cea1a0b5251a13afe0cc8936fe255587ed5e08e7bed3060543b
zd9c7d8b3d6e979ed5b1e8cffc0277201dcfba3413ee0b6281a78c6ba60282db4f635d3cdf6661e
z9267db7f8a09228e51c77dcdc41f195132c1b538ea4f929509eaf120dea830e728ede5e8e3ef91
za276550d4bdbeb438ce77d694a25ee43836446e8f54c7d313b9d25a007cea6ab29a2a05f1f9925
z472cd9705e12b7a013c08ad813b165402a7933be9907813870036b624beb31c4dfd655d71d8086
z0db421081b88a8eb217d07a522c8683a3d12c945208a9c07f3a95573a8c8c9d66c6b07b2ca778e
z5ad7a6602f7adfda420fd0983788e3c895158c3dbcbcf9c4a4fd670f6d5e471d56821b9cdb042e
z1ca14800d80681beea4136caec563d4fd7ee08524e9411bb7f7c96dfd3f643b0e44f17cbe992aa
z726b65996deb2f5f6bb5f44406fc127dab383ce475685502040de186518b8c78a056d73f9e7c56
z7804c78daf520f63291092cd2b03a4708928f9caf46548a56bb1cc2cf7e289f6856ade6b55daf9
z0c45b6d5beae55b55aff13117ac59c793fe6635de179b3ad1220686fc0ba52bafff709a5cd8d02
zc6e80c6914e28b517d5c0c7bea6382a53aba22d44513ab40e86c48b69275feb0d75d8d43c9d906
z30f82580d5fcf94ed0ac7150ad842f03b528ec17fa04b26157342950b32201b04b0dfbbf1d3aa7
z5b8a0ff0e5c54d3d78d9db9e9ff5e99d45a16b497bab8abf54ff8fb36f8bf9afce36a9265598c5
z53bd8330606b95f5772cbb9782731ff9f5a98e50b91061cd4f145ace530ff23f9870d398be9f79
z82383eac95f8502fac6470b4d094c61024166962451202f276d93594c8283245ce2735c84e7f4c
z1186b4526f9c6072e3c6d84a9fb2eaa46b28136f60052061472bda47339c4c44f98ca0b20a3e39
zd22367287158dbdec3a54136ca00250265a77ea991fd3acd7de19b81ef1ffe4ee85796d3bc5093
z958bd80f961ee6fc13a21dc322fbe1858a6914601039c6919d39ebfde28a2160b7f1f72e7e2392
z1b22d105a3a446cb87d62242c45ad98f39edfb2a3decaa0559a6e36d5cf419a8adcdecee4949e1
z4c58f6050911b6f493a164f44f9030ae747553b0db98bbc0393e2944f3fec13a04f47a44fa0904
z48c77c492ab0fc39d6ccfb2e3a40fe4585f2f23826d8a0b63dc6f04e44348afe535b3c49792194
ze46f18d085539ef1fdc725d8975bcfc4f16273148b71bc13d38d862f0878a85a2418cc64ab830c
zce4ce9e8f43cbae9bb482209db82d598b1b4f7d3936bbd4de1d022d2421fdc00f8365e66338633
z6bf76844b6fc09eda26741e3164c7e654b4c6ccc13201b921d95c8946f3a9d0776d32c308be8aa
z2f62599ad501e041c9a6447512c3e45b207d625dc2990700968d064904743c6821257c86f8e0f7
z8b6134f2069870b5a0572288250db62e5b63fa0de19ac50c41d48e62ae53aa769c898857f64cdd
zb36b10e16b87a1b8652dc311806f66e2b371b1c051db34989956c47cb0e8983f00625aebb2f411
z95f5fc809aedd1fca6755a5fae29b4cfed48fb55918902d922ed7e155466c1efd9dc4a30c12ce2
z9e1286736e5492595e7d17daecc003d4513e5452aef12327c2b0daf801fe2c85da24e3a40a437f
zc24922f935595b7244020d60a550dbe987251ad2058e4077d521314d423fdc0b5e1d65105cddf8
za7879744ab08fb972ae2a5847ef7729d3bc337ea67bca12c83b65f541d08ecd16d55ddee7fc13b
z47bb2efb129b3b16fe6f38a808bb22686570fcaa75b178e1bcbb36d90181adb11cef5d2c662de2
z7e74ea0d0520279f03a8c0877342a9d738418eb31018ce67f699f287514b668e69c2a4ecffa944
z72c43647905cca61759410341459409a666eff541ffeb064565fcc43481d9352bd158ee2eaed5e
zc1c4f5236f537d7e552f9281c34b65109b5fa807ffb973a84414231a36a78a026eeaaaa445a7ab
z966dca06987e29741dcd4e56cda376f0360e9c9541352b722fd36d6717ca15effb9d01ea2ae0fa
z8c01a4ef233067ba6ba5ccd6b6f1f13b1733b09edc54ebc0
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_express_phy_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
