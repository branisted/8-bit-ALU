`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026201628cee5aae21fb892db766c4
zb5b1406e11aebfd6dfacc9da5ec03b70c276807a3eb15e28ec7ab1dddec42388b9424ea285623a
z248195c9f894b36317ca6e59c86f11031163f5f52d70922c037057ec3eba50b955600900b32628
zb2250f2b4fb3ed6db7d81b8ca05e994209e236669db511df2c321dadeee74880d12dbd5092819e
z312f2e640fed00f965c7b0e1d2007d987dd08e1042332719768f689f95a8ecae54578598cd4014
zf52c9aa29e5602a0a7c0b59ee67317c72101e7d1c45c07570c0683c158486b6e3157427e0a2514
za97901c629a01f6fd65b5a7f6f7538b7ab683549194b5767ec9f9eb38f388669f93633863ba210
zd15b4f9d05bd96c35341c02c93752c2344db76edf8c697562b3a09dd9e6ea71115a107694a03bd
z48c4beb95a5fdace643d8acd8693678fb3c10dbc716d343185d0f8c8b090128427948cc61f654b
zd79e08af23d1f841dbaa5dc1936e4660e1f04efc36d203629f18a16a4829e3b3126751fa196d42
zfab93a2769d0d4af5366799eff9987e0ad2be0898f05a8a7fe7be72a09e6e962114c35e028f985
zb4f3db4d71c39b999c96003b9bf32fb342a15fac3c4446676fc11b463a9620113254265646ecae
z71d7cf3381b7e84b560f223855b0b20038eec96c1ac4f1af8cb0110cfe327c79fcdd2413920852
z093eec9cf19ae3cd8a67022d07fcd7bc14320c1ce4d9db0e528514c98a62b5d3ec31605cf03599
z4d6eb850c37fec85cf69e6b474e171d53ee2bef5d245d9cea5c101e34ebfcfa73468705933e98b
z1a22aa5b32d9f8d3412392ed7416ae93ef2762a663e61a210309cb52001dcd4a952d8799718756
z65c1db60a4531864be9bdeff4cefb56beffe2bf29fc5f3345b63d7f8ab90e88a20287661fd01eb
z5e716c090119d5d4c08ccdcf8d33e906a8990d677657f34d4716cdbd43f372c20c4a03b754b7fc
zd09a688dec478294aa8052d341050720e84add185bba28dced0c27c13f7c8c7cf2b793b02369da
z080bf6eff0124e7ffd1e395669b8e0fab00d0bfbdb7b4de8907980f17ccc6a990eab828e203546
zc08cabef41d95483de759263a68379bc58694349f4d092ce1c8cbc4d8b1cf9a2a993a7ff3c5dcc
z09f2675b286e7c0bdacfc3510345f25f7fb48b7e6c7f9ce1da3d69c5c34d4db08c56127a25342d
z438ebc9b0fc4b41f387865b25eca0c1c664f5ee46d631b1a7b4d9f584843a2492f0e6a4375f36a
zd408f01e8d60caa0c7ece9914b89550d320296303dddb38ebdcb4c0e7f0efc8acda6e6b587210e
z71b5deece77038173722b7fc945257e2139de2f2dcbf3aadc1d4275bbdb85bcb926eb21d7915d3
zb4505e7608d3cacfd452b687a6788d931c6fee286ac5d74f5c9f498cc7bf8e2d6a6fa197c9f1be
zd7a9bd147265b94b25997659e046511eff70d0206dd77b5e79fb7e3597be5514c639de1d19ad0c
z05f2c3f18ba55f3e7c2c8f092141ffb4ee0f913cca02e0bb1f8f8095244c00ebe259e435dc1712
zdc483bff00a38f281dcf7256310edd6ad95ddbb1c63d82d04456f834dfce146c520a936516a50f
z29a39addeb72adaf9354cedd5aee8b848376fcf1e0930ff8e2955d5b97eac946abef96dfc634c0
z6d65c11e15339bff5a665cced0fff422a2050eb221291d0a204f573861634a82d46ebb13a2e7cd
z54a1d8766affe05b30f533b4430aa6b644138bada310d7e9324ed7ef40e05343d0133ff335b54f
zd0d1c9cf7af527f1fbc9ab345761975776946876b9996acf2b0a5dc1c7ef3a01b979d3c8335fd4
zcf1e2afa4711a10ea38eb5070315628df9f656a8facdea3cc8fd85bf05f0efba585907a683e2fb
z271f5adac55b7d0cbf1f923dc6d77da4ac065b2384eeb11fcbe4e9c4e286b3e0c8397c9338f4f0
zca5cb05d0221de519ac2cdbdf7c08e1a0d16dad14ae8e380d9909c159557fb377b8fce383efad4
z45ffde49c2a441c977ad7fa3d21d5968c4f3a81a3e92e97006f07e017bf15a9ce2ea866c3a1266
z726f8bb7dc1de780ca7405debe14b37ee80aba4e7b76374f984cadaaed3580ce6baa3b3cb72960
zbe04c1b7c04cff28aff46f7e3f9b9bcf091f352d657f97c0a6ebbaa0a3a3001ac19742a265e178
zaceed05f28ee4a98d5b7ca9524c364f47bf2ee066fa1c7b24bd3f92a37fc7bf54d05e1135d49b8
z5ae86802077f20b120dee2b5f8b0ebcfc182c8e312ccfeb7c5565e05e0d92e9b004e270557636c
z0eaa4af7fdf69fdd97f4e917e9286879d6a905abc5d3189863e716f36baee1e21373197d14934f
z200239586e40591852f3643e60624677f80b662e95948a9a41e900d5f6c23f565dfe90df61c04a
z0f7d290023a9543e70690da44322df955e5018cd25caedc3f54092054eeafeec2cc984c8520e86
z6145286c957ce85aa0acd996cf7e5d5af3357059038ffaf73fbca44d913ea5f60761be04bab3c9
z2478e767e0241bda4cee164052e43967c4534469f54063e9bca3b2811d694dc45ca7dbd9937e6a
z773c817a1b807133773e5db0d2f32e689321d06d57ed5a963dc83e3a30211b3cc8f052fc82629f
z119b3a5c9feea68b4363f0f5bfe3725d9c528b2e9ad558a81a9e43ba75ba67931311ed351921ae
z38cb0fda266ca34c98305f40d92421b393f8fe7658cc3684827c0197d88a62e7aea055ecba909d
z93f23d1cd6513ad88c54c83fe93b13bf48352a644055b0115da01c5ba6a14c482bf8d8fcd7b35b
zae4ca8396c69ebe6e229164108d506e0632556aedebc0256e06b028bf00dd9a70dce66c48acf25
zb5451026d6249962f13a15f4a1c215a4f24bd044fc1924dd04f5fc5a7a86b8fc01103fba9e9f17
z5a4b7d916bb85b5bcf91fe3f255906acdac8cb1860eb79ff5032983a578f89a934027ad5e4a03c
za0d64470b622084a0de73abe83adfb0d2e4b41cb5d929de63cf88e7175bc14aaf7bb3abcd35935
z92d1ff6e72e6a77c13b3b2934202d1dc5a371c42c2426645f2c5920af881ff7ca22c0e95d135de
z70c0a78b99b03829ea8edf2e441514347de79056a1b64d02529d6bb1119b515d321b58e739eb1c
z79e74828cf8e2a5379ed097e60e4259b854c2bf84f5af00eb38b920c2623885a57ae81182a602e
z78467b72725a4a106a09a53bd6cf4b69d7b3cea9406d35103b52319b1a26e2cf21b2c2b4321302
zf845a8dd882acc1edc800f7e3e8eb094e9ee738e95fd8fefdf7e58e0509aa6b95c4058c5056748
zc2d1d30f7defff1e4c88aea9dbf058bd92a8d2784050cb4bcb54b881566dfeef527d45154810f0
zcb6498ef5eb60dadd09047339b2bcf92f1b319cb663b708ce0229f187bdcf988c166ec3c72d3e2
ze7eba3d158c68f7fb02ed169d75bd2620e3ccaec149b03f6ed11d192671affcc6b40511bd2ffd3
zf2ee0900091e62d9cf1592b830f40ddbde28a928b1c483f6f9a52b9c3dab361e30aa7311606c36
z808e436d7e7a968e5756ee057eb22c8e2c00c96323a67e8a8e8a2204d5ee369edba6e62286add1
z3f485bfa08d555f9a0f19ae9ed796847f76ac09181af9bdc18835c13c5cad793bda219832ad956
zc64c22d20cf88fd9bb905083011610b8d2b97910ba9eb2c37a73f546e04cd872d3092e4b301bd9
z2b659e124e6144acb1d75c1f8c9a06b5254ecfd9ca898681b502ad6c28c3f39dad1e6afb8afded
z76bf60679879d0519fd3074134254c59eab676eafb0c7fae1713d07996eb58a73058ede0181190
z124b68b7adbaed52348dd24e48e74cf6441ff004f50abcb25b17ca3af2a45d6cf9e84bc3081e0e
za4112a64b02b2fc67026f7843271a401be3663a045f57f151cb528fb20be9986e68c771edf09bf
z1022ed17cef9197b82ec780f87eb2bd677db2efce79a61a6c8515fd25167cea226541494c26567
zad1b87cd50c89fe35f95db2fec6749426580ebc054ca76a8951a8d35339aa4038a1c7c45abe63d
z6dcd95286b0d8b597c2fe08020f10963a518110af9b3c553aed3e16fd6a04b3493ac25b4dc2870
zee37c992953bdc7a72aa3e164622f4f0b4e0398efbb7109010e02330d0b1a60ba5c32e8b6b29ac
zf148bf37d2b7bf29c7ad7a39bb3589f9adcc41b55080ecc05af85172e61abecc619cb7c2b04fba
zc4bbbe5e6eacb2452a3af7c9ac24c1a21b049b9a68cfc54282777f152a15a0b5a5e66a3272ae59
ze5f5af9af996426238d1e07ef601310d1cd94d3baf7985b5f4843ac075234eee28e5da50e880d4
z1110dc18be5e6393d83ea0fe5858db2deb4bb0022ecf4f56aaf0da9bde7a3762c29d27c4d5a78c
z123b51d2ba5ef358fc46c99a28426bd2d31b19ce236c8eb822a4ec0888440a259b70a0fb16213b
z16dafbbdaabdd02aa7aad0b44498772e72562b453dd7656da6a96a9012d4f82739fdca30c68ca6
zd41f02ed0df11ad470316fb34f8b347824293fc3d9c091152cc02d7153b3dc45cd35000917a18c
z2ee48018df46aa59ec64005a343f3c7258f4c22f49b07321dea4d966a6def7147212c2be0f192d
z9cbb75e1392e4ff063adde20aa3f8787b5ef9fa5cffb2b03e55b6929530a37936841ef7a2e2b9f
za9aee566c5eda2b48073d63c3411f0b958b53a8a1f8cecd1bede7c415bfeb4082e2e4464d9c7e9
z71091921b90309d175f21c2a3bbd6dc8b1fee922493ef8f80de2f2888ebc25fdef6deec7b7c349
z210568912611aed3f7aecb456cb0ed5ac4a91e37e5fda1b7dbfed3bc0b40f3d6f06c887a390154
z97eb62f77f6d61b54d7ae41b7778d7f204853fe8e089b83ea420f8d8186f1f5dddb4561b1ec303
zd34f256ac3e67ca9b76bddb7353decd2d13980997a3610e41e2343d52e10ab1866e7243a87057a
z6067dc75f1ce66680f746b930bf448c9b067bf8b915d47f4f9d3915a49b13c42df0fb142eaa64c
zd5eb26f2b05161a938241224413315425a11a1e90000379cefc46eeb83811860e6c26b8e7215bd
zb3c153f9abf9fbbeb7b4e3a64f3238c1e4c480a6b382d8f535190a65db1bb227114f4ec2acc78f
zbbb2f26c63950ff43a491374f1e50aa138c12a5ba0de4e79e8c9cea452e0a6ff8fdac33653b5e0
z9a61890192b0a1d79be66b34eeeed898ecee8ae09c53558c7615814ad05e07463102b0ddc9c600
z8e6b87154259c0402e5873c54c650d861d59ecb86c2220b66064f4f4d6b250120b0e8903e421bb
zfae2d1b3a5f1b055d4bb218a4955628b627f54713d64cf19ea2c553cba16db820e3e6b30d2aef7
z8e8d5f5368e7da22101fac44fb6a170d5c86eaaeff5e06f26d8d4d90a5221a66064c4331774b33
ze59fdda88ec8eafd63cb5c23f80d19625aa90d91a12873371056bf5df0d2dbd703616c01f10771
zeed764482ce852c9920be2e2a410b7fd88a142166a807a010d1cffebc48efab4a35ea58b79cdbb
z8b04129ce927ad10e85c45533ad828230ad1a32b378e728d4096e0a85b4cfd2b2947213aa1c533
za82f610df46c4b4bcc0e3c188a5de4130f6e0280df65df414a213436e34ff264f85aebeb8eb50f
zfd71f3976e21cbadde2fa4dae405521e094e4d450aae27ab666f563f3cb6bb06c77718055e52ae
z0599f2374ddd5246ca55f6c469ada63cf4a16f43d8ccfe03dfe94c9564c36fae4a738852728f6b
zcda3113d98e1ca988fc0bb0b738f5936088cd966f3a9d186053624cab7b879d912f9090925f0a2
z3f9a6600039d473f3b23c033fa577945be5977e350349605c18589ca7c15a9f298871cacc66b60
z3c5199e32e4157b553589357b462852b8b49e0e2e6e10c00d68a24d522c55ae14f3e8c98458b2c
zfd56ddf399776f9e24c69eb5aec32c7281e802264aacf6424aa53bc363628d10392391bea1cf62
z5df6bb2f539c0124da9c8db5c655f9b7c172138df51cda90a576a397d3cf5630612d4ea697298b
z9604e1972f8415eeb665718d6605f8e0ae1d5a77fa5443562d446fbaca0fbeafda014821cd2ae7
z958b035d7ac9dd96a128b1980c8322cddab3446276ff9751e5743ca6c5e0cbf1494d94a640b7a9
z07412b2087e05894163e06e5f7feb500aafa16156442f58a5e1c8a63e498694d216afe81885d92
z0765dbbd964a1c18c781b1007db2ac28fb3e35ab2805ffffc9b0a27ce598d239b9942946d58abe
zf8cc321730b6daae724842a7e48c17e184fad430334c9bcf33cae032f99e5aa847a23b853b6523
z485daff3c29f66a01c82d2d61f03bf16c42d19fad6701feb8613c8029bb88ce806c0a78de29170
z9d7bff9eb5c8f7c7531ba888912d90c668a7d187c336570d15cff0ac4f34b680c4bf3bb6e3e79c
z6c0803b42b5ab8b224f07674015f87405b1687dd07ac733d80a771b2a11ed156a3b4a58e01aaa1
z4741802ec01d248e125a5ec6dff56de828bfdb9760628f731602dc0ada14d80ab26120e4fc8eb9
z9c8a084d029fec90ff1b06c711fb776ffad10112829c8bc60b427663f913b837cf84f3c030abaf
z353c042eaba43de94fcd339444dfcd79a7f885e392a58f519edd7436586ab82de87386b0d04724
z8e22364e0e254c3dc42fb86b61937ef46bfef730623f6c19d5d2833106bc732ef15e794ca41099
z6b781201dc2caf549c5843ad9d982cf01c701750a68c6ff5266f0c6368da92fbb96f0bef62a086
z6af595039a71137db0a95f9780f15c3d24d7e349b95dadd461957019d18eed16dddc7214c0f056
z08b56770f4211533367ece892670fff38c2f2b57814594925992430dcf9d1f8c0aa07f624137a9
ze4d5038659e4359cd4110972755f3d4c32563a8975e9455a5e0beb7da51f16ee08134baf2efc7a
z8fdbf3bad306486f1d55bf6d8ee7d289fe70a4cce7411642ca1f636be4f5c474fa57a99af424f3
z0a0c2b58e0db881498b0fd2a282fe80557407365170fb2c3aee5e53fda12ae8240fb637e98b821
z55c4ea07597e6f67defed3b36de35165a3549f5375b586240378ad5bb1bf13b968ce542d4c922a
zeef838e2646c40c0d3111418d3730087c78a05a37522a8bab61042973dbac563826d2cd84053d2
z7b0408b5b8749ea79616261a27be2c62ee18e6efcc68eac2584a4183e6d7960be575d1ec1cb734
z192176aa701ecc8a3e7efeba1ac620a359c76ef194b391502aee580f01472e8bcc8a93505acb96
zc82a75f58aec53262c231e20d674690a3fd3a1ade7cf40644c1cde28ce0bbdc1df887d4fded3d4
z472f183cfe525ce5f21b435b2b37a14045c4785a5111e0b74db970dfb6750c97ac517e70f4d1de
z416fcafde37a1e3ffae185a53c858ef1ce9884d9447c4be7600bd187d8e769db7521e0038ec5b6
z9358ec5c917d7bb3497298401e05bc8edf7da4044483811c518d7d1298de8fad460a6c131011d9
zde899b0366ee8f7616477b92ba0c6133f7ced3f0f843446e7b44f67e056442cc3cb6285754825c
z10d648551f40a93bb7185cd316cc71ef83812fc49463a50cc344d1bc070ce2860bbf27f9ab0561
zeda9afe8374a76362e96b60cb4c1fac8263d785fe1b8d7903ccafffeb23c90d74dc74c177eeb86
zf4755c4dd0c7fc6d0b495168e492933bd856ecf341208696b2af6da61b4e66575777127f327a0c
z4facaf7f2f098e6d4c0e85cc5f2fd7c89c108d1085f6283680c6fe8a0b5d765cfee5ac497ca7cb
zc84d692916d071dfe93e5901d108c53c02b50ffce7cea1465a1b0cf4bf91d62dbb70093fc9999e
z721a66ea725514cfc1ea1243dc66b66492621be6aa7716d830464170e631270c37378dfbf7520f
z2bf6a8b131e40d99041f90589f9a46101e6d94754df779274141bbc8bf74233b8c7ee422611414
z2449a06974d623f132de4fbd35d68a5ab91f816d08715b97ec7842ef4593dfb86180e2ddeed546
z380775e06a2960bb630345f4161149fd92bef7871912f8a291707a81dcf83312edb41c348a9e9e
zb5d03c04966b893143b5530977e4c125cba9bd4b845c1029bda3e72564c30034ef7c58849ddc32
z209eeaca689907632d68915f2a0ef43b058d013ed660905393ff3739cddea0d5a778647140a959
zbbfcdc43871f910af5ac19f4ca2392e01582ebb04d303ca037258cbb7777646beb81a3e8ab5a94
ze41bd70b7f099308bdb41b02194f4d74fcf93161a59b01833426323de5291280d9e5e21ba205ff
z886a2e117df99dd2f3e71f831c61c4c895bb8fd7a9a4250012dae7c867d529f3cf277a5dc596ba
z93c316ca7857158ede6ba553115fbb2b26f98f502156d13eb419f79b05d5d504ebc328d1b1ecc6
zd226e2867968532d69eb6f15cb83401975f62930a2bc70062f86342c9d030a9fee801d240460c5
zb24f8b7337085633e332bc84fc041ab425e10008077ad3bc88b5ccbd62417b192dab77a3dd065e
z5c07e94e8988827ca5c282cacf8983c5b9be6edfe4bafc4ae71a0ce84c4d4e21acb8d1e1d3fd2a
z2a5d3757ee1473b9e1663d82e0bdb6d1f6e8d59abc9171f32edd0d635e67f9e3a60e8e2611ba30
z0346e531ec7cadd01ae258eb084997f72d6efcecff1ecf1210837c3c605fabe07dd25d30f648da
zc18d14a91e500f4becbfff02f8c399eb4a8a58ceee92a7d8f4d707e0f9a50200aecbabe3873dae
z5ca3a52fd28c521c91a800c020b9914e6e933468034b23b20563fda3abd337516a0e093e3816ef
zbf47ce50519f0ffe8f4eb01175df05400a2718002ddf7300794bcf50a36722555f3ee69202971a
z915e29460281cbd59dece929ac23187f8ed89958da73c3a260eb4df2e7943011bf4281f0f6b4da
zf561f83223fbcfab501c80361bc142413cc822058151823b2aee8bdaf7578014275a40ba8052ec
z8f9456884382e26fc123f706d8ffe9730259d0f5c3f3af3de56c7068fff217d8b4dda4eaa61f36
z92ed57d33d1f680e3fc1b281c84570b7e08d4959c35141ed76a7704156a0c29119911ab722c5c4
z75690bc89321cab8adc772d0a4e9d4944615eb21484eae929949725fb124b193bf7fa8e0b5e3a2
zdeb49a0b91d1fc93c646446ea7d6cdd0b0f4b238284eec27be37181e956365bbf2342c8c71cdd1
z637cad3cbf480d9267a7be9bb34291d515fa6117c35b585b5e148828d7b1bc00bfa6818aafcffc
zfff97c8fcb5657ee12c274a591ccc10962cf09643c05404e6971747856239a542812bdd54d5e66
za8d7bb0894c5eb15805d1765d1363653c9ad6a81b337093d0bb0570c8c6b764d95fa29acac07be
z79a657023343e6ff69c5b393770c5153266f32da3ce00e7782db98d95d61073447a77d622129e8
zea241e583080a2d56a3ad889260c5c9025e11cff952b438e783f3b305f45d11be51d4c3938dc30
z32237fbb5196b13887d6e847a14dbc00f49f3e967a76e78e0a1de33f3128b0173821a017964900
z55dfa4e710b5d35d273c8839e04001ac269cf3547a8eafdfa4beaeb48b43b03473d942ba984d6f
z76d01e544c623a6a2fb9c1b2da395bfcc8e044474c6a289e513de0581a693d5c405e9cb1ada49e
z667e543c17ba100d586ae3f42f2d5b07f4885382213ffa40c66ef3365f4213b606876603af1f32
z667b5f10a98057eed30e461fcfbecedb3e150879906d3b61736ba9f4f954e167f8d619c1494052
z47e7b61908217b555a3c8ba5cb2ae83ffcaa2aca4688cd99758e7fb6ee092bbb842102c86bc4cd
z9da56d62cb10ee3335c604c96dbd1515c9a1f0d67c96f01860c6c85df8c75045e74d9e087664ad
z4a577884ae21cf7d16c70bb5fe4af095b7740c2387a871f7582b5e35627dc2a1ab1e00ba34e21f
z3ab0cf1913a76193fc46c5117c3fca1fe784b77929162fc8681931817437c4125615fb734112a7
z6757373404372c48ff4dbdb203f23c9aa10e6f433c79da597540f3c3a145152450875d0bb6f1ad
zc443e1feb027afca25d4085fde816ee62d9b6a73b16f10e1d1df4c89ebb4d70282def987591e1a
z200af7fed08befb44b234544c801674b794417959f683c23dfda4932a7bf9db677d9bdd9085a24
z877c0d508e8e9a71b32fa4a3ed976e66ea7206767c54d9c61c15943e1d91882dbd7dd2841059a3
zf9ba008cdf1c46ea608c9e7e4efa9ced6086fbfe6b1b547aacaf1fdb07b7c4a024a36e97c01b5e
z71873467f2c6bda6b3d02911a6e572eb6fa13cfa7a40d668a57cc3d77fe3387c865d318eca1064
zface2c548c983fd3ffe8294a8e69b3c39376864c68e7586042da870cd677b0834a507af10b4900
z1ade20ad2965550d0b8230d73942576d779776ecf36565c5c940d901ad324ccfeb012da6e58529
z4e85dd68135404795e6ab54422e7644f291550dee7d916ca961185db2551a67b3aeecf9121d0d4
z1cd416dfb29dd55062743df5b8db57fc0ccd6058750aeb9c11148a0dc8f3b7863f2fe1eb7ed372
z6d2a58847fdc190a3c5dda3805b12c2e615b103ec4c7bc7759a0ddd7223c4c9726d9e9871dfe41
zff4918e75df377a4e241da16ade72515fb8e687071e2a6377123dc5e652d0ac08b19cc6fb779b4
z91a1e6268fe5aff4aa7718b5ec28cd3b4830708d8544dba086b007a7d1f253e0c043030d44a86e
zbbf0a0007f828c0da376a796d29c668dcfbe08f67e5916f3f5e82d6ab182638db58c1338b07abc
z1f1d38c651655c377fa7cbffed34d6246b35a7842481744b8974de83c54593b7e7dcaaa8238487
z6b1372370ca2d63ee1f649c458c667723c5ee2b249ec3a7f93260ebaa4b687f3ef2dbe63d3816d
zd62faf5656dcfa086deb212eaa6f186c15bbda4786cd1880d793bf161dca9a862e20044b71156f
z99f9779ebac424ea0bf3018561220a12e5c75bd461438a344404c32eac85127a2d303da1efe994
z515e69a87c8c9ac966ce3b4269cd0e28e1f31743a45882fe1c152c4ce05383a1a7224a04245685
zb0ec0cdc9714104f2cf86870e94d581e4accf977d5fdd396f729320c4dd4bc03a3720188736e7d
zb82c0ab6d4d75e908713eb61b5777da1367f5d800b0dc82e2c43bd44fe5de19570f0225cc85552
zee4ca96b044ee6804c5857d0523ad4028f33d7278ee6c7cc619e314023a92e4e0ff773f45e3029
z093aaeb07189116427355fe4076a7e4cd66253a1a92138a6a40918f9412d998cb0f59520dc11f2
z29e23bdec85dd269a4e1c65fccdcbf210ca230b2d72059015a30252d8c2cdcb01027cf9b5595f5
z1128506d1ae245f49b603eae7b61a6cacc5a5364ea38a665f7d9c1e4a93de95afd59b7f7658e56
z27b8e191dc4ae35fe376e2bc2bf48e46918b134a72c35de1cb50740b6a6b81539065545e55fb9f
z7c318b5173cc7d54a35b66b4752f79c701155b20614c63302f8da8a12e9d1bf999434f68c883e6
zf7163a7843754f8935af1e49e03cfd497e8d5f1c433b670919edc89a06e070bb7624a8b8e4443a
zec5f4086abb8574d94bb2d702feab12b0365ebe6630c4e98eaf7d7dbaf11d41f579c51bd9c6f1c
z6b26022ebe984d6a4f1b1ab2886db70b9f80606eb770eef23b5cf3e9ee6504f5ed73214461ab0d
z58838ae91d6cbbb2e581fee1f34c75b98890b82c5fa94d1a07028a0d09c656a5683097c42bfeaf
zeb1ec798b16855a5be366846d0ff01062a15f819abdb02eaebf46859332e10864e5d305b436ca5
z0345431abf97a2706c54013c8596da34517cf2b5ae9af9ffb02881ceb1045ce0c0ade28999234c
z16e3e15e018a6637bb66029b6d28d9b5a4bf44482bf5937f393eab9fab0b5adc2686051ed8aa00
zfd2b20e90e6f32239e43acdbb40d1772d01ee9256de94972f7d744abc9a3c28a4ad3108b81d2f2
zc826c01ee4279bf4cf8c0673ee421d19f038745cf139e00dfbec8b4e78ee10ac03835476b4bbeb
zb8a98cbee81b9a29d37e127f06c8174bc2c14840304e915204a6b99506e57d4e4a67882a6239f9
z2ea6e5a92bed349f7ab549b1d0afdd2a577e5eb1108cbafa6ce2a0ae82f2e527f3ca1780cd507c
z723ee28254ada2e552216f4cfaeae29d65605d5f1c5151f75af5db358085a34eff68b5ba46a4d8
zc2fbd89b7278f43d749457e34c574c68912deb24a20c8b25e0ade6b7d9120ce64df612090691de
z1085522fac5bab7c0394d7eacda121f7e701c30cc715c0fe45969f7734bae4cf1e99fb3d2b799c
z793e4da73fcfe0b538761d53774ca0b4f62f9e74e9777b484da399c79b8f26977d884b4f20b1b1
z4c2dacce57d1b530e7a0841158b876a149d20d9b24c6cbd1f9e8188fdaeea7869fa2fd30a58214
z0c5de64ff46d81f0d004b8f53e3c857747ac0683eb8ca9e92fdd481b865c824b4ed6e98cdfa7a2
z9f76721fbc9f713563579c62d1b6e832f7a50510b14c321ef44da81e1370f8dc6273145c039bd0
z201bb262ac155b8ff743cd3d3c2344c570835d960fc808d55c204d86b04c0ac9bd9335519d7e58
z2a67b62c978a7dc1c55b59b3d3203b82dfded9164b6e1c9964b5f0d890f9ee0ef2104f3bd18484
za0f429746720dc90a20466b088d33cfa013ebcdfac08745446986639ce8385be09e2d81a17425a
zcbf4d2743f1b3baa1514230c86a138bdcdac4e73bc9d7681295f834aa39f21c2d03ed9ac82ce48
zb9fde38a3f493f1a76ca84dfa5a82c4760c681904cae448edc547174c766265e3ef46e3d5004c3
z160d43a5a766c3b27d4c091cc2d3a9ab4864149072c12d6fd4fda18575a4d71500d2db38f99d3c
z474a2177779118c44e0fa16b7ae3c0a4e631192f87532744193dd75f6059ce0f7220baedde3172
zf89f997fbaa3256b011a3f030ba29679695edabba5f66d03c939c65bf57a85bf18d382b0bb3ca1
z9d896a86645fc7999307bf191b7bb846297b6b578f1c8519c5c3efc86e7799e67cd878ef6bc12f
za0cf6535b876d7db009686d641b5a43573a072532de861a3914b96dcfccc1a27eefebe79c89154
z93dc84f7ab20bbdd1d86d246b639427675ff4e027a909fb784708640c9c7a05a94fa1dbc91c490
z5123ed124b81f94f670882a686d2d9c4fc348e34b33c24720675b297f19171a8283e61ac1faf68
zae606185f68bfb43a6b2653ba09c5181fb97c4b2620a7d772d15b524811b168b141e8b15a4bae4
zd5a6123c7646ae1d1314b3b9aa654e86b1efda441e873a5a36dce17a7b0f692cb618395176ac5c
zd9d125a9c96ae9450ae810a9bae0315b430a62a17c01491724218271fe84580e930fc03de11d07
z82175e201cb3ea1b98b1bd0b14e97dcbc175041ee787a754c5ea0e86240f5f4c115c354740c5fe
z1d71ac208aef9fd8bd2332077ae7ea0c2c9872762c08509e628fedaba5c00afe2ff4c71d6a22c8
z0e8987957e1fcf90faa90fe30fa814307376a1555afe1a8cf125ab50c373fbe9e86a7669fa595d
zabc58c80d276a1caf3627bbc8b65d8d9e9011fd47794bf58cfa8998df66d67daea2920b8de4ec6
zddd82b87deae8300d190e40aff11cec81f66a67da782f2b0db3a7ecd08abaa67daf8df55e88b92
zf0a3a9f7d8ff1241d1a9a12535dd570c921f1618ec17ca5b4f03db733c663cfd529b797db13b79
z58aaa73fb4bfbc13babd28efbadd0c0d8dd7a5a104018cf7091da5f022c8b78ad9739567962b48
z08b41ca261d45e9060dca78fa340856e9dc652f5268d6bee6b7acc9173830995cae88700d452e8
ze93cd681946ad34ebb796c6d2a8054d41dc453e0720b6e7d04dfdcd733103260135220fb45fd81
ze82b5ef9343f61281e894dc6f3baa037d3b71bb0fdb2a853587f8ff6f6be87bdf82a6f46711f24
z02c4728594e826dfe4ef298f3b5ed5ef7c9266be99c258ecac73ef6ea765808d187e8845910cf4
z69b3f8888edc97ea431e3cffab0035fc8ba968757f53a1205b7d3a3e2d22bc0da14243e9ddea5b
z3e8c3b17fe9dd7b0e1fbff114242c6539c5e39e1138467cf62e88fad272915694f945305739fdf
z0ae774571295c5e4a33121d5dfa08c6593558bd53e2a6fe99c551ddfd665d5e1bc44d505708fd5
z63e0a55720e11a4c534bf0dd53b00221d9e12fe3ca84171dd54b58ecb6d5078ac9cf298ecfbe61
z140523217dcc54e2cf5186ed068cacc4102d1d3d8107311b200019ca2e559304df636724333f0e
z5d8d3d1916d1a7874484eaa12903ef25cbf9b6684313a38ad58818ebce931563d62014f31c4d7c
zc33563720053d80c251b46c2f81d50ea48bf5a7e16c45eaeeff689e05ec74bff9b6a524258c8ec
zd633bb5cf76b1d8d16042daee7b463d8149fa3d32c73d8c5207ac001f526a9fbba8ce9bae63678
ze3f5cfa72e15e94dc97c35eb63ee291e8bb78b5ca21749b8e5100b540d820264c19c2dc1842c39
za24527615191b5adb098626953086c27479fe3f591a4c045bc36017b89bf4b874dd00e09b97949
z054e498a7203c52b608365802f9879a19ba7b87b7c1a7f0e3539b4e17ce23e9a68443f0fef34ac
ze27ed1f2076666bc1f83881d0e8855ff2f0d69d0f5a9a7f553fb522e160d8461fe6922230528e9
z2e310cd87c341ac18fc7c8c6240cff996576bda195ee84b84f480be75d03fee87e4337be0d06cf
zc19059701dac37799f4a2167ba56a59600b4acfbaaf7a06c7fbdd6cbfec4ba947f4689f79fee27
z27c0c39e5cda613d7d204603c437fe6ae10b1de156f1367fc27980d2056e29318e9ee689074f01
z520a28c6b1fb5971f80424bcee96e70d4ff19554a6d19d0002e7bae03ebe69b32d50da8565b81b
z6afaae713c3e00d5bcad584b35f57bba7a1432506d700394d78febaa1940a57acb6c219269d28b
z9e613b2464d59c122cb8cb63f8aadbdf563c9b3906f7b8672b73b635539f05972a304680a67dfa
z16831ab2e479254435da0ef280dd2ba32aa9f603a811059e359321047606f240551b97b4e2612b
zcd8ce359b9e5d215443f158648f5d73d8799d391d4500c64410423a5d12cad60980590bedada8f
zb3490c576b77c8d7b344cefadfe834e5caf41e3bca35659ff7d22c61fae86c4c6fc7865e42b59c
zd2d5c84f99a19d51a8b7f204c1cb0463e7eefa9682d2e35472e51b613e8568dda28c53bf23e39c
z719338b9a63a71befda21ff51779fdf72f88d5f949e1f6f3e2e5f4f4dd7ccd551d99af63d6cc65
z1fd56eedfba71879a6fec23970a1f7134559665bc22dd2192f74fcf717b5bacb5510c74879227e
z0be443eeddd259c7ae7da7330e10c850f03063e056844961046e330b2a12f46bf8a5db1a347cfc
z87e132ce872333243766a27e5cc7d74dfc5b633702ba6af3a080950288edf6caf1e573a751adf3
z7654845cb8c17400c6e277b884a4d5da8f758abe46ee00732953372482a07408c15ed4bf7f6f32
zad2a3d3c0575ea391832e5f18a8894c98df383ca10ecf0bd7212be9125fc56c2a1408f1d1be1a2
z76c7d03a58ab0d1a9af8f7ce7cb369083d5d190fd3589ace31a1718508635968a5217b07578e90
ze036d5831007541e1b1503076535e4ac2566d2ab3c030650843eb38e1eb4321c3c674902c423fe
zcb67f63bde423106d50b680b0c063bad59245d743b0835ef6dd4057ec8aaeed31296d1052c4e98
zfc3b87b1be3a57e0285cfcb8886f6378ef23226d0c8ec37a5dff0969673f7e788862d1bdcc95e2
zcb8bec0245ffa90d1d1ec44d594466c667b6e5d785c27f6e6de874a280b39c7c9b868017d622fc
zdecbfad026862ca3da05ecb76d42957c3d79f82924f010f33c85d0a5d599df76d5dfddafce9940
z82c1201a737986e492970dc45d38e0520118d3e8e257df455bf2e73755421fc40d30eff88ef3bf
z78b2b5c777b5dfc1c7a5f520e25e80766c87494f02a88469fe32c0040101049bdabd8bcfa0e9a3
z7f528bfd7c8a49a1a27e58672d1f6f658688dfcd0bde2e69e6278ad8fd0717e5f93c927986cf51
zceaf3508d96cf21dee227c72e48273e057cd7da063f2ffbf93fc5a024826df2c83c0c4fe4cb2c8
z10b5bd7967266957026297b41f5036e4cc4755cf474fc8cf3d8049e24ecbba50061b4cd8adc481
zd29a2b678e986c47bc3439e41ba4e55c77cb81451e409757c337b37e823c20e6bdb5b7047d5779
zd5413d9b01e47b16b2b9e77d05227329f9b15b0883670797508a25a5693bcf155d68f2d516e764
z7579738783f87db4fb517681ca912c9688901b47ecfc992c29306206259797a4f2d7349771ab78
z98db758d1f1bf3b8499d8b0c10c12a8d15f9e412d48d474a2a6fb3eefa6fe2295553c2aead98c4
z464170cc33571da7c155b06a2af041bf453f277abe6009e6782f5eb134e599afac946d1000829b
zfb412a3292e0e37a73518afdb1362436592cb9dfcf147dc470a831e30875bf2e170468856f4fc8
ze2be5f1073e10f23b8ddbde4a09a70a18f80b73d9e3095d68bb56d896325b56bdb03dfe86e8909
z47daedcca5a6bc9719c89caf6e4bb13a6c4893b818910589180f1f925d80115ab9d1cca0d7ee65
z15732a2a6cadc6e608cffd855f109ef55ee3e0362a9800d763253f1f536d9277aac140f92a2208
z48e69ca77ee437aa25926e7f072caa00e85ed6ba76dda4db2efedf77309fc4171b9a084f74fa89
zac59c6546e4298b5c55c17058c7b26c7cc3e6b6a38625cfdb8c8aae495070fea05600c4dfd2127
zc022311f5cb8bdf016d5ab6f49843d7eba0902c72dfa27b3579a2e5bd7c91ced4bb59cf4edc765
ze87936bed9e099bd89f9a4b00c61f826c79bba432d8a2793216de927809af7af2333577f1585ba
zec7e37b649af0d9ffb9062f05b5502e85dd148808b28ae57450f6f2254feebf75a490fcb404a4b
z4738afe267b7c44196d9ef37ac6959dd8a43a91ad9f5bc49bf6cd7854b414b24e0a525dedd0688
z9ed07aa9650990f546682bdcfca6ecad878354a061ce69f5b6d37b44fc8b707ccd088ee8c59dfe
z2cedc47353bc148311eb594e2f40ad5f04332220f9dc5845a08976571bfad4fc71e39329fdd60a
z82a89fdd37f7c8fee51460ad2a0b7a082a919295c18ce76e302e8ae7f53906738483acbb56c7db
zdde465ed23bb683f95e7912e7aaf976f7839546f963ef9904fb1cd385b28a325a2ef3f8e7732f9
z9308a338c72a437da30834647a6a442f81df865f3700785bc86328471f147f134b71f4b8f9d95b
z406472e8a0d453f8320e6ad863137d266c7bbb82e02a9656a4d803236c01db8a98cdda1aed6832
zcb37f9be57a7a5b6a898c4ebe30f3f0fe58d845a7189ad8a4be67106fdc57738664e8ec446e693
z3d35eea1356d211fcededc92df61d457ab836e2e91559045a315ff4f5a80900f333cc079a825f3
z11b1ed13c2c50e9566cfc5386bad4b5e603adc3ded771bfba3e153c1fcc94058326213a1ded152
z982c6c1db5444985ff6ece79c188d869d070e8433f767a3e3834bb5309b16252ee74e221f40086
z49d7c045ebeff3fca35d0110dd079e4f28f4d4c032f1ce905cec1f4752b57a9783ae2554ab0875
zb2fa3863fe5ff0239313cae29f3bc957ddc7700fd3b850d0a7f167dd0c154c68e7bdfbf5453bff
ze999c534627b57e8bfd00db748b991bef0228af80fa39f0d2c54c086662014d436feb4ee57c6b8
zf47b8d2744f7a1d484068adca14b06aa4276a414605a516c07b4aad5a111d950e3f03eb90245d6
z60e2f90af59ae3687cc357e89026bac784adbfa1bf5b2d09733bef04abef05cd131693df4900af
zcfb96933186671644aa7b9ea0455298830c7ede222f12e9a8127fae441ea55e0a4a0fe72ede168
zb4aaafa7adcd32ed7471d494189c575d7807688be8d5d4fcc7ddf722161b78cbc1013c328703c2
zad8610b4fc6f36b21790b3f5739e54671afbf63204faa428ae777283b69ceebf6335f1ed88e493
z004a59e1ec4e19528af357d5ac502ddd89a133ae06464f1d6ac2e58b3804d769df0ca5bdcc8f76
z81e09f966c32a9350c88e940118fc808c311bb6c2d310d67247095705ce414087803d13a9f82be
zbbacb69c89c7ffddd9a60b83585519f5bf6ed2dab353b3d4605fbb6ee049a3d8dad51df2b12939
ze0a55a0f009bdb1bfaaea249fd069da6f02e3d34c439b9282a4b320a3a9e734eeb4256d3fb300b
z2f67b4fe424570e4b17b3d3b8cdf6d369ef6d45532962987a664b264da50a36af3d5fdf650f109
z077f050034b32ebe9cd63f0d942d53cdfa322e6729f7111f2e7a15e30b20b284693e12a9212207
z94e60df616ee239e25855b329525983c92328c3358bf5b2eee7ca31b7754630959ca34884be3f8
z70cefac5a7eba7e139d48442864f89c67798b8daf38059126b6d6c765a421ac965776cd5eb0702
z43f813881ed517737cc6dbdd20fbb27da78c65b48a8a65a83cddab2ac91c94aa9e2cd491f62261
z45fa9789642bee7dc2e063020d2d98af186fb3618bdbb4ff61d33a61245f67471a561f8999836e
z5d5faca1d5717bcdeec2ab56da22d49a6f019c6b6b7a984ad8affd384984bd3b3a24486c909e3d
z27bf5ec31de15ac213313309e28524e000d03bdee4dded560c2168141702f4a39c56e29eb797e4
z95139c4d8abad7c83073ea6ec91729a5b1cb4439e16e2cb34bf4435f243519a518f718425fa13a
z7c41ed9a4eec141dfd0533aad9403005a712e9b1a2bb5b8ccd8bef669190ce93e6bbacdb25088d
z7e36d6824a8771e8aa219aaefe70c12df58b63be59823c4fa7397d7d0de0aea9099dd93922b84c
zb81202e0b72d84606eb77c3443a9ed248ca50e653aefbc3024f6cbae52f8b2b94c24061f2f0435
z14f7abb14795e03e5083acec4a92543ca5d758f021b38a9bf48a35e88201953c12632b5f965bb4
z68da742e89136de2783456896b3142e57216d5f12dbcd047dc8c3a74166cb1ad15871f0bf0871d
z1e50c67056a426dac134a44258e72e8cc6e70526fcb65f2dc453036d95c252875b185f3ff315c2
z67c6ea4e80297ceaf95ba801d591d40d662727f1ffd311e92e53b7f258e2f4294a46e63ae3249c
z78f759d2fa79572d017cecfab678db60d2c0d624aeeb595a7e76fdb7bf33daba58c5e58e1a7698
z302e967a6a62b8d40c63c42029788ea8dac456b87e53c0bf9fed51a03e772c89b7bbcf6555718a
z6459be4e3f1ea5d8c081cbfce2408948ed7dda5ab23bf2892057001162e834936676cd3964a5d3
z5e35872f732dfc2da438529828e57be41cb9d0b18afa84dd6aeb0f190bb3444dcfb5743e291270
z34eb3bd54cf30147c93afdd0133d90dd5b8456ae9e596b1b94e1567c6c1057db35314dd1ef6a5b
z05085eff15ce3928a0ef28aa0cac987955a3992ff712a081967901798914251fad7ef4440a3a7d
z6b05513d6b49c463ca5efcc6add7931392004c43a24756ee0332f7f7f882fef1fc8402b0e87dce
z7740dc76451d93785f0456cbd03b60e7fa0a18029393bbe21f192fbcfeb5c306fcd528f05fbd69
z9c4761db41e20dc1645272b65edf23c2e53c23ba0945f7775053ca196e12f5620afde1302953f9
zc75362f93c012551b80855754965c5edb87ca344685aca1a4cf8e40960c87e7193fd8f9bef2278
z68b08675e8bafef25eb3fd4b8f6da679a9b5adac05bcbaa625b0b87e16968f85141b32e459eefc
z03236df0d82d8013e3bc706c3fb874d9305a33cca255e6e0100a09cb7c8ec75f9900c0399849be
z480188f778247722e6a86fa998d0471a4025e7136b5a5478a83852def6c66f04d28eb75d8ccb26
zaa99e0464f7f19ade3e1ad4a5f7f739633135022f2e02aea645fd48be1d44e91c2f6e6f22fb7c0
z1ef9f3927a38838361f6cad6621eba4246fc7792ca60eb30d1fa21d400dd44860ceff21b146394
z0cd7a3d5b409d6816ae1ca8c488c9f248b584749843574ba3a9a770487cae5e31dc56c9d3ee293
zdd840677b503bf2816d5939c0e263268a067a0dd39c50542da9f63d38e5d274cce5335dce3743e
zaae2b5f2c77786a648613b23fe5f4160fea24d245b87e7e6feded0753ebaf0d4d7eea29254fff6
ze5ae21b48719c46774a5b44829d399a0b485649afc8eff3a76bf6262056b9517a59718b50a0aa9
zd9e1818502b46d0b3999c6ee7ce53a0d1949f78abd7394bc3136c672ddade7bcb8af9d9c78feff
z845623a7ea2e3fdb36b33a91c6c95f90826ff833a328abd2bfbd1d8774983baa853279d4e76b96
z3fef434525406aa3cf08423c3f738e1b66148f01f2e482fa30c222b409211b8adabe187f0d91ce
zca1f7d30b937f33d9eb09508f5022132b8a2b7319afcc2a9c4c1c1a3643a27b639606981f486d2
zff68bcf9b8896c4472e026dbfcf4c19a41f1920f8686ea58c590f439d945200bb0200f3a2c2fa4
z8a97c218d119bb15839d1237107300f977d4776022fef0c4904679ad438d6f9c630352dd5dd2d4
z602356d28ca01b9644c4bac76728d54d7200f6fb388235b09afb833b9605b82d94e3aa61bac818
z27acefa68f53179dbcc99e3bd1ffba94f4591ad6fe48f7256e4dbf525939e1660a3b0f79a2b89e
z1aa717c8a17455b523e3d4609617007cc4f9d0ddb207b84b0d807f00568629814e39aed50460ab
zb6b0cb9686e28399fb498714c4c1d2d1d8956389fd2756a0e331d19397c1e2b4ad93cfd883d401
z465665941406a62267b71fa8ac467a5d646083d5ee375a070f10ef9583fc0286bf879ce89e10d2
zc169e853775287e799fb1e08665a216d66701cd0c8711e7f20270142923b7d32cada2b90df2095
z5517696dd9034a8e38649d54b676aa59045012395e4f47995bd64b46ad2e720a65f2cdfa5ef78e
z003d14b8de2c86af5fd7eb41102220d859891f7833b91a64436be3174de66a92297ec6622415d8
z07de82aa43fba6e3fd9343184ef20ea05b3c83f95f244d284d0baa77331a010693572e6dae0264
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_i2c_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
