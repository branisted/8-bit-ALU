`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262e96b75598c81b19220790e3a0d
zac0e9cec59fa3a7263133e4e4c54ed27d6f010cd2be3fb7767eeb444f708ca477cf85da9e49072
zecad6036a0395642e2b7cf96577620ab5d97fa265f262bc31917a660e40f512c01144e41bcf570
z93328ca57ab128f2468b562581edb4b6fc48d738d2ef42032d2ee4d32de1225c9eee5132642703
z815d6d52c9de6848a675662d1e3a839e490eb95e7c589e603dcf7f3cf55a57ed46c2087081b6e8
z4a5b235c4d7ae5c0e87920b4ee54de87eacb2915463b37ad1971b45e768650f016271758ab6322
z5076d5659ef437c746302172c55ee35882e861b2ec7367720bdad325906cc89294ecab9cc5460f
z89708c2a516488318d197cf92cf986677868b105bdbfc178fcc175b9749de5161ace23a9d25bad
zf3047c74f552f8f0e8f9f048cb8780ddd312151b47893438f1c54088fd657a5294f1d0a4fd1307
z711e0269e63f44033a834d3832c41a66f775f333d7871489ee355f5d4df6a95579dd8731bec839
zf20da1a0a220d5c0d06d3c5cc356a3f339973208ea4c55ed0cdb956a766623a486f8e21c1ce8c0
z9eb3ac3a10f1380f338a19dff906fb0147afac33da863e282b2c094622efa20074849fac7620af
zc7e576f18fbaee41a11972e7acd581273c1edcdbe9fd9f8ee23281f86bc24e4ab438d7be05ec29
z7f7f730764cec476a130d30689224639ca1fe6f4e9e26ea0f6dd497208e911b7e1546a90ab1a61
z0780d9e7f1c795546c0cacaffa81cb3fb7749c04f008a9bdcbf24ea0c07a50278f2c7534418924
za3a48335f7ea39bce45a70a92e2f3830421aea76896ca9de37c8020c9ca04fc166a58b4b26fcf0
zac02117fbe7b8d24b50435ce53aa4699206742bcc83910a541228039c067793d26b881043aac07
z3c1f3664153b8b24fc2b6af7e8b1c165c11cc52748646dda83e0c14048ea2d10907b093f7f23e9
zd77ccb342d9a124251a289516d2e6a0781665d36c7575c4624c65e71c02e2365ceeb8f8f522456
z2db2bc436890754cf24a1b6b5f72db5e2e5e5cde2b0c721aa26d87f7236de27c3a219867fcee95
zf5a0fef72d8bfdc9b2f4c511e8ac80d14596d67bb687ea5e4466e34d9e09c4c4e959de04201145
z0c6c472c6bb3dbb09d4df70f59d99cdbed790f2730e69811205bcfed5b85ab97e78c1cb04dacd4
zbf0fe84a36ec3fb7e2f516aa1b895add14dbe9af990983a24ec57346fb52f25f842fdb2186ff54
zf06e9e033fd33e32b5ed7f0337b290bdb9bd882b062ad74ccd7b7a75b24b8787dcf57a7ea2832a
zb206fedb09d7041007ff69f6b4945d7ba018196456cdcdf9d9ecf7a82a78659d493d45a2ec2ce6
zae1b92851881e612807608d7d6b3e11a583a28bdb5fa68819875a4329eb8d37230c3b8c9951b57
z56f64ab80a282fb1556e633d46ed0045c5ea9328013bf8314842417ad39f4fc3173bdc384c6b97
z5ce53d8930175774c652c52e9ac9988d7d04cc4599086940f9e85ae13834cb0e9c874ee7f24548
z8f02c215e6190ea3ceee97e5af83b4dd98ae8c4fe93f000af383a63929b6c40c8af6a1c6248b89
zfed6db3f680997c992ce43c1a3f658543923eced6cb059d666d66b02a0f645e9687375352c8117
za0e5b0808ad511c5c8d637c5b2d54a7a0a4c9b670df6790a5048bcd91ceca91850cedde570b502
z185b76f66a6589252dd901bf609f4d5ce855249cfb99e78d69ea6dbefd15c9cd9ede65080ac81b
z33ea1084d72849051f80715d65e5878fe7271844c6ae2385b922b616121be4000951b4a12e6aa8
z16e3193694feadcb297664b1de5fa656ac3a74251bcdc27536f6cf2157bd55f772a87117b58c1f
z86022c7ac057e128bc3aff3a44c08257521938582bf8ee16b4b1046a2fce920d579dda71e2b035
z62e83e71368b08dafa39cc7267c3f2209b66480589152f99484259b5c6627254ab48326f2504d3
z1fd1c014f64702af061b2c4a2cbb8fa7d3f22c3715e3b811798a2a776d5381cf347a4a0752f1fc
z2d173341a71d3e6e2a39193114483fcfdc8e87ef70bcc77d8296b391dd515eccb2c739e09f6acc
zdc7b07a8daa63869716dc7d120639de9fd71be6a65bd04f16c5aac71a15a0a880313601c9c469a
za11afd149a71651658f0556e4e15108426f09751b77434c1688b98552fb0422391ac7ca22cc4b7
z9ae67b8f94f110ec5ac7ea4868264483584d5c151ba42ffe03804d4a1e277c1e3f732941783fd1
zb9c179072988cac81e6fcdfef115ab2b4e77f9a42331d93d2ad8c5cf5724a40b33886819d8cb78
z823332b39d7d3015ac928621385bf6b58b198a948e8c7cc3d2f2ee9c04ed33b612bd7a201d6ae9
z3005af8a0c43a9d27758e3d91fd070cf4407f5590755d5b408a9839f5c39e0e743d922112e1f95
z4503f5f0cb45798863b061ac22fc23218d78ccd08ff9a5afae9f88e7ade160d36b7fd784382b3d
z7ff7647df197526ec6a15791d75b0c2136ad5666a2e34d7eea5aea2209a24d46522895193018aa
zd97d384a522a820f0f84779d5683a5080e94f0179cd02c0850dcad9d3eb4919d705f4e850061e4
zd695f80ca3570b680f63fe844b3e9590f339a85e7bbc747ae1f94f67b0df009f900e81e7db894e
z46f695481e58fc7ee566f7dd0aafc74f9c0fd321044bde99b84c6386ee1b28f1de7b313b068172
z27ddd7e514206cf298b38afc2563180409a0c70dcf987fbf3fdea870bd1bb5e927c2b844fdb4ae
z68519ebd979c5061581c7ce63255a739d9337e6d7644bbb6072ef5b6a44f4e21c8396c13b669ce
zb5599b5f4b8595a82f381028d914c0fe2855eab87bb33084f4fa40ee340f214b77dd254d50ab3b
zf00ff01bcf2370d7c726eaf5381f8415ac6e403e43582764cc9351ea4dfa349fb62466f7482900
zb41ca24a8aa454ad923acd81c6ed7ed6ec12d6e72f455559089bc48bee1c95486e37415c85659e
z1da907d3777137cc18e7b08d40ba0df9f2bfb840d6c57818b56b5140c70f187c7f76df3bc0eaf9
zcb7f16eb020dbc6a692a663615203ce72fd8e1f3f27ab0cf3e6df4e70dafe4010614a3d4c39dc1
z17144359dbcd47cfe22752a57237342687b9b35ef652053bddc932e73e4ecfca8b44b7cf9eead8
z893a6a84a945af2f70ba5f1199e8f28272d176c074e2fa75c3e7bf038e63c1f4962b0c7234660f
za5b45f43dbfb483e7bdf0602e431e04af4635e5d1acc7f7de76b402babee9d071e297ac87497ac
z4fd4bada55bd5733b1e08eb022886d8b162eea1ca47248e6eb7434066af85e033d8ecf0f8b4470
z9f9eaba334eaf32614cb1645c4ff21d242ca7a3d154d5da1db1b92ce184026bcdb3263c9d951c1
z8ffa009dcee9ed5df51e348dff16ab8a3aafa6c75cc804af89b37362203abe033f5959b704c0b8
z7edc5af264701fb5a9c231a6b7bf6cbf04dd73ae32ee0951c5faa545d00364ae5969a5b51f8c7f
zbcb60542c4fd7505c6161a0f2abe58c96e17e83bdd9784753d98c0698686991f627c670876484f
zaf1e8f2209a9c8bd8d53c00ec3bd79b66054d75aa9a8a480356f5f6a04ad6f6a057499f127d5c1
z5ea763aba17a8770be3a1bde6801b32948c72bfdf6ab40df0ecd13a2c6a7b39f1d89df7bb75c48
z84c987df6723f440cd1919623d1621fb0ff475698502d7662cce0a27e60d5ca23db02de5cfa506
z9dffddec139fa8f82b9a943527c862a49a530a4dcf2aa5bf89a5768dc749c21ca94b686bf17599
zbb9a2d8f16bfac6f261303eaa33ed9f2217fb75bd7176b74915440ddcc132c98dac94ae79f13f2
zdf8be372f46a7d09d22781b7bc85b6eb065789519314231752f37bccc141686f791a128ea87e7f
ze52e9dd8a277efe869074af1fd5f41917fa4c5090a361746b76bd54ed363eb839d8a02fd1543cf
z0f5bacbeb75a3a5c97c2c3608e72bd8bd178fc126546898a65d6e04db6a8d24af8634d9b4ce1a3
z2cf945aceacd22cea2d71618f14dd5da8fac3d7e1a7d31172b3024d9294a2156254b1de7053d89
z6b6857255c107dd832861628d535a14d95b02db762fa899de14cebc16a4deb002aafde49c809e8
z8e947d026c391139a469a8d95db788f277896ad098692d9ac501b99fad93aacc349637aa1d71f7
z67be8d9a2e5dbf4993c0971d2e286547f03cb749d1d8e9c9a79e2bb25d8a5137a5e6389b1afca8
z726b0547c1ebe85b80fe2730347a91b1e06738ac4609884306a9eaf512ee11da26d267ed5c288c
zec656fb182029363e147841403c81f6e3d044741aebd37763435f4ad64003b99eee3aeb9ae5561
zfd2eff5f4fcbd99b37edc19f4290b07644a819ec21a21a2d38528de7a758ef4c0ddf658d746bfe
z3d9e17d864757e61bda79f0c676c1c231fd2496b2459e998eee72ef961dad573dde5c5fb59a245
z9aaf2fa5fe55551904203af7abd0d6ac65448698093139058fcb201ce2f6dc95c40165bf58c2f8
z9016b29613fc11f9fae14da369eb7103c0e1a1125f835f606325cf2f87bce51dfb5775afc2ce8f
zf70148e7df80d0247bed530b701f8b024a17239347e331eaf9bac9bbc8266f18807dd5f8da01aa
z5be350d029fded77db1ef6e86385f0bd0c370e7da4ece0c663fcb1f2670496fe9720b92061a7c3
z2fd02d9093fb31667677fa3ef002b6661cbcae2251b2ce30c4c639633c4b57760fb61a0697aa4a
z89aa0d894fd5a877f943d039e433260ed3c581b57caa12480fe1352de7b134904c9646ef50741a
z1cf962142ce700a1387929e47608c42296427b8e7cf1e5902576b946ffbefa5d7a7d5eb98d50a8
z0affcbec064412d179bb7c1995dd3fb882509b261848e37bfb54c8cb16aebae26cd0b619cdac93
z4f697b1af390b2882bfe21fd8f445bb0b998b0b818510b04692a0326227258c3bce77d44527681
zbe8732664e05d65b0558aec08ccf31266822782b447b394a63dd48d3744395236cebf0f6c38ec8
ze8705ccf884a1b0e4605e6db56d6a92a55dfb7209f9a98157d6fa4a67f185822696756d43338e9
z22df3483ffd434bae089d656c7e5349010e20e1cde8652779757bfe7312cf0b6b7af3f634e2b7c
z96ddddf1a2762a6a79e19bfeddef4ae797aa3f5c9158ede1861b27f88d7096db95f60125ec38f6
zb1ff818d73547145dbb0d49553b57bd45c7fff3821f60aee9bf4494c4a6cea3530e29639818f22
z9aca01a95975c7f126effaaf12b47519eecb5b73ce86dc3d8e5c1c2881fd2f37788921dfd0c771
z55e6e1874268e6aa19c85fbee252af860753816b2183c1d424515d850f8f177de84e037e490228
z7d72366feb7149884079b315957dc00cb3f69d5de4fc37bad001fd4d824980a491063fcb3516f5
z47ddd9880ae96a27dbe7aae08c4f4e3e76be457b41e999a92dd3d38363a75e864d146d484a790d
z97557cb6358588cc19b24be6d45ad28d39bb27a9772e33e0cad95e87ecc8fa9e74876aac62be6d
z49a7a64c9cfbb6801a6f372be37bb3475b916af8141d9704d045a3eccca4dd8609f33bfa2d181e
zb4a6bca173a9bcf48f20978aff049a4acf10dc80d69d65f6bccb0b9d72da4b2072d7c64b084569
z288ee6e9d3025fbe0dadf4ce7e32b8e03df245d74f859f1e00082606ef3e5025e580278d936a8e
zd0bced56e04fcdaba85bdd9a8a408947362d124a2fc0ecb996371c30e438854ee932d0d97589a5
zd6a0b820e5cbd76a2c455d0011407e1ee03614c3b748e89e9f5ef6441dde299e73776828733d70
z4d7b8f14adbdd549758af3d0d291eb80ae5a4f62236e0afe94dba855488ed7f3b932693dc5e7a7
zb73ded28f86c0e57ad0ab84ad179488cc494c64468dab09b3746ff1a03c82bac3e8cb9ccf3803e
za61e43f613b8f93d596622ef01a2dd497c081107784c4addba5b6be018d7d8d27ea928d01a68a3
z51e6d45b2de800c2aa92af860ab01b503cade98798295fa671a9fc3e862ffab2069be938248ad6
z055a014c952d17e9210dedf6ea4cf0a64841e3466323d8bbb4d792ee34eac4982b62869b066a59
z9e83b8134bcdda994a6ada027a72a7e98070a465f815bdcf96b85adf9a28106363873d70e3c8f0
z99b68c2e356b1a00032cb7705e043f3d54f0dce194fb68e858a29ea2aef705b8692f08540a8d20
z38af61b03c702e03916ad3e139700c5f9f24ec0994b1482069b9cdac682d9ae6c884f3317e73aa
z499ebbe8a7a9304c33cbf18bfff2985e6674a7f88c03ba62d40766389472c0f00d81fed0abfafa
z9fc75f79c57d63b037ac4026b2e592ffb6fbd1037999fc0f48e1fba74bc8c37462a80396983cb3
z8f9007a1e8446bf764b3eb2999900c005f2f99bd83382857f6105eb61214a665bceb5777417450
z9bf09d14e26508d6a278c0d35b9277bdf08a7bb553a60a9d77082e69f8cb446e9b020afb6141ac
zc65c1d956dcb7898709c2839c31c5eb6aa77270f776db56db140280b0a31c7ce132fdc9187c226
z5bc60e340261bf0bd597e0ec8663cd76a35ee5e5a31c1a70354776d681409850eaf60ed2e8f946
ze9bd060bd0123033a00297ed3b6be3ae18ec6fa58c63d596d6f8620b0e1547d0d776e08648c484
zf8b3dd5c8466a9fa209c5dcf06329356b0238c37073c2dbf3859c846dd92928daf6b31ed957668
z6d7fe0639cb3b977e3385b95bb5f30265e8266725271bbac7b8d8192c964597ee0a47b0b4e6cab
zefb7b455cba024dc385e6b81683b5e70e0a71be3348fc6d1ca35fed2760e0067ec6b578d4ef68f
z61524f413f10214d7a087ca865ed97b396923b33d834eeb701587d79704f6a950e2e4bb3b8e157
ze119b01ff38d3fc555593f78e65baa48712c14566b29ccb65493fb07c2a309541e4a206433ced1
z01b15914951b9c0582636b544b10a59ca6c9619633a700f1b2d42f9d2c0bbd6da92b08f6439542
z74546e9ee8462a679eee4456c1484530f551019dc4255dc5ec48849a314704aac5af5847ffed41
zdf8c0e465e6d4b77837ebb6a9c37d2dc065f840d37c65950adabb91704db27302c40a4d5357b6b
z6ac61d4249e03ef3788ab769f79746b8a868b4ddb7375597d9664d40953d46000834dd390b0ab6
z47656f7ed2af384bb3613d9de7c1872566258bd89412f3f2b0d3c38ff79e300375b4f10ae6ccc5
z7eb283e7ea59ce78ced750aa60d316a7509c3396937f863efdf2c4dfdd29e635ce110e59ba8e38
zcdc6264c101a53d09bdaaad18797d1a5c6471491ebe1e5f021fd7a2643f6e3320ad0c7e4fe6137
zd1235ca384a60f9d8fb41d8c974ca6e55e511a4f979c9e72ee8f832c147184f56524fe68aaee59
z6c3021daaff45ddb0679f264f0b498fbe45673fbb9d2673976499241cac2668b1e2e8a09ba0e14
z1af0e52ff009e7a520c2449f56f9589132a9c04f6f1b888f89995cd84fd213c899f862b8b18943
z9af71e081fbcf71d0e90e53a67eb0a716e1dade0beb4f792d272a2b8784b01877445034396c8bb
zc49ac13f1a082fe043c0ee40406c4dfb4b28df5f7f179bed3c21b2843f245d5d221297e6591c36
z8c6453d62224c457f9c563ba8e8a7e0983a6be4c8343bec037d743bc9448408b71d04718f264b2
z430d0908f2ea0ff3c47adc1927f6a6b2ee93339455a736f65821c1a4682b97cce1f2bf9979f962
zd9052f30f22c7f09d457c0d8044d129be59de1aeceaa5d7664c375e7404d37b6c3b92bf6b50c57
z0597b3f1c235564991867ab226024bffee63500e301a5506ce73548b475ee7feb71035807811a2
z73eb5b56c5aa2dc9bd06b826e1bd6b420d2a7f51ac3fb9274f57a039aabc92eb379fc652f75e19
z0fadcb0f1e5a127fdb588f0e7aded1442e1e7b20a84ff6cbb6d443118689fac0c7571dd0a819af
z6c38b450630a43b89161d03e74f71ff6e0a852d034ad3fb9b1c90c21d7aabf6615fccaf41ca717
zda8df85bf0a44611f278731ab8e8c42f9e725cd71e9e57c48c6eae3f512235d311e3d884948bf3
z7cd3127f62122f4be8d35c2ce64166400e429bcaeb9780834f91cbe8deb0a3baf4835fbd2c3297
z45d82c333a1344ac59d3b289ed7715a709cc7f1e6a6da824abb73c25a80c93aad5a96a83eff0b2
z902ed7f1ce213851b7eba59c77f41eb9101cdf9ccf5c46aa9dc1321e98f8e3b509deba25f62672
z922398af07237ea2c5570010a42cd5fa95288af58e1f28b493164dacc0f0af7145c7a66b20e4dc
z0b97dfbafeed80426aad7a4ebce3d4826e4203ffebaf22be627abbba6ad4778e535cdf877163ee
zbfa403c802acc311a387a0ac203f5a1ee9ea1bc0e871e1d621d562abcb57bf6e452a4e76a282a6
zdf9600eed3294d689e75986abd642d488009570468c6993fed4cd54ac9ac3be3de1edc5918b3eb
z677cf7d2a582a98614d37f083498132617d2da9fa3573fe5543ebc1fb3ce8ce688ce1dbefb22b6
z314fead21390eeeb2356123610adcc1ea3237189f6374dd7264044a86802bba229ec05bf7ab51a
z969848a0631dc81a6fd20a2a841cab6eb6a7fe7c3164dc6b7de25b02410ad10eed4606200b0883
zcbe5b7266062bee908f9c33387f29e6c3d376f79eac732a845af9dabb4fedd91b7611c764cc94f
z9cf927db8fa7bd36b6794a00ae70d374cf0cc30ca0076621b1797284b40788cfa11b43b7576abe
z94d50897f13f7aaf488ef9d904eb0b4d07a7d1e31fa7284fc685e5b2956eb8bea9ac1110ae9639
z4031b4a7fbd0093586d70e51715ba6b150e6bab769c5bf739209d2844dc23c6c5f74f507442650
zbdc0a4de5c58fca3d196f4ea1984bdda0e9f1b6a4bc313dee13a1e92b7b17983c2bbb9050c235a
za37579dac4d6d36a92bb1acefb4ec4fd34007c7d5ee67f519abd43b87a35125e6baa5e8e3e6248
z0a03c3c028ee3537d3cf19e243111ba11a9fb31333250aa8d94a92417061cb92412a94bcb0f799
zc6dedc128fde5a9c1dd10d97a7b2581261f07bb7464b57baf8a9e9abaf9806ccf4e389dd89cbb7
z0da99970919d9a4b6c6f4d35a211f594fb030330351c0fc514889fb1ddc91fe72174d671b2cb69
zee0c811ea3031ab02ea5e1c7fc65a75f0caf407265267fded3ffb9f9de0665e4d01eaf694d33af
z371e8944b31caf5b14a28195c6fdd1efaa56bc093682874aaaedb8778089f5ed3b9ebc19a05dcd
zce6a7a0c8842cf28a10ef999431918cb3e4dd81e308995ad766aec85eb528ed0490efa3698f3f4
z868463a7e20cf43421bb4338e3e9a6bea5413e40c87e96fe3cf1421c96b5f3fa848181a20fdc14
zcebdf0fc2d3b15c0924a528a0beae862196e9455de6a9b45771cf619d39ea8b09868354478d356
z60419e600b79c02604bfa0e36442d00939c66a4e685cad2147317de5d0afbf38c8e5be0b8ea287
zc0f57c7265b894ee876df8992a494cf55e229c8c37ff3b99efab4b9080c29dc1ec02425ab3e950
z5f3c16524cdab10a6b7dbde0b62edde5cf6c17584bce13a42639abad71519a46eeaa196565bf2d
z77469b9b899a198d63b3c1d91cc9105a9af708f26582098f6127b0ecca3d50e256406f3661d247
z46c3ae0aea403aed8170005ced6d5bf1d524df2576c93f8485525897bc038b4701a4320669ebc8
zc5a7ded38b751e7a01068d12c83e0843770fe0681252f1c29eb60d6b2306a0a37f13b3ff0267a7
z7f779df077f16ed79fd0ac20e2a6efe35b5c4272e4aa658cb3a5e0516a34b63b574b888a79a270
z13cd2415f8f1ff2c9731fb0546a89bc9321b2796ab186d69be6c6c3cb617765f0df935bd8499f0
z7a8262ea4eebda559aba28430e63f1c2c9ffdefb85dd394538b963a4767142233aa5f32a076a8e
z270ce3f7079765ae5d0efc4313a0cd7b508c06b24e54c2333fb59049bde73addafac217fcd30c7
z688b801f2367c1ee0798358a4dad96ea8db0d6ea0688925ff3592ef0fede54d4ebe1dae1aa0492
z5045f55a3f776a5fdcd7fde550495803fbf26ef4c0aabd1a87790805877f1edcaa25b475e1b7f7
z532686e7fce2189559192d210c1abf62e3e28023bb8b38919ddf75e5b997988ced854f4d9d1f81
z96bd90f7a018de21d224d4e7c0e00d56827a5675af6858e21a226dabd29db166d57a53cad13132
z3a6bcbae8b3d22dc03de255550f0073230afae40e9e644a8157793dce1590a1f6ea091dd7f0a56
z3af89bee32242b35f8e0f9bc4a999334f88cf1188f680630cc4d6d03459f3c55a8abf3afc21951
z2a2241fb685df9fe553dc67e73242b12264bf17c828171d266ad66fce8d9d1e54f028a9131a6ae
zdb0a88f9a128395a4091c261031f2348872a270c02b2dfd8371e91a56ff2d7d4884166117569ee
zadbb1cb38df51ee8cb9ee09d1c34b8f7e2adf47ddf63979424bf538a3a1c2e457c05b3d41fe9b0
zc14a5c331d1118a36212c14b114471008b3928fefdacf7037bde49947f24d81c7fd52f503db747
z16ac66b5560918438f1f30e3fe7405a8478037bd43653e4c5416a795dca7803611ab02ae7b7fe0
z5a80ec3fdd800217b4188c2ad8bd1a92c0d570213a925b8372df90e6bc57331d47f65cbc6cffb1
z76ed1faab82905cfb2eb619988837285e2445449af415f0774d5384a5c7bc0b2dedfb498e0534f
zba2bbb66e0e1486e3708f93d6cbcd0df74366378ad805ae93b63bfea42622f414ea296c6ab2622
z39d212f9a13f45eec205262dcb7c25de86709b3045f3defa3aef170a091f66cc6fb111b68ce044
z39d2d0214c85f88d614def5fb4e12187ef054c65878e2b7481114bdad8e595d22f51641b9f957d
z2044613bca4d14db38c60226abfc8a76e52763f7dba9a7718ac08b760fb369458ac52574558f2e
z5f9401fb22120b7bec832813c71c1cf54e60f29e3257c29adceb6d1e2131a14d92a94338ea2539
z9fefd77478a89be14a443032bd7c31ffe797e7e74116a47b90daa561c1b6d20d9f38bdc045fcb9
z024aa78104f508a3753235b28f11a19ca3362f9fd6380dc78c274aca2ea8e0b55072d075f5d3fa
za3c52ae99a52a2131fd90e9aae1a2a91b853ce1bb8adf1a3bb24ddee99ea9067efaa43a3629ca5
z6b29ff47660dc79407730d878cbdf1f10c7bf835f7d9f9783a362c8f25a8de9348d5f5e9a0c112
z021ed7211a6a25d874f644dc360e757471288c0036a099702c2a05b8504362d811d6834c18cd38
zd0ad28878604e8f7562757ce8373fee7fc51381238a14e253a2e4b49e070231df70880ba39561a
zb77919f8206091f1b5af582e246bbaf100c16ef13cce3370f41869a52a71f569e708b758295528
z90299daef97d8109058687359530df650def81db614ccc23919c0456e65d6dccc8ec6439748f09
z5f3cc4f2f75ba60d6a695302e57df96ff609948dc646ebe42b315149074b0c66aa97cd4af73012
z2644603c97b1644f12601be93e9cc3bbb57499d5dcd8ca11a358efeaff19cfab43f26e4eed6d8c
ze8e19d5b9b56e41a7892d4609498dc850615d73d3dd495e8dc6ce98da8a6c9ca9887833855e424
z9df489201216ee30a0a66a11a82fec4f030c841295c76518ae9eac38c08b71f749b8451448a458
zc2a4449c47c51658472396757d4a8cc8f81af798e14c8c30f44371f1a58e851d01dedf0a8309b0
z9ac11d63c9d4d2b98653de8a874df43a09e4d371d06bcefcea4cf958d34d2cc17cd8c1925fc94a
z62a9ef4eac577b47c3f686abb06cdfdc3227d1ee81fe08dd36a8ad3147148e104ef2edc292d10b
zdd7d106bfa7a396f3911bf65e55003ff5d5fe4299eb28765e633fc84a53595f8d86cf2dac50a26
z13d08f0fba4e15882a3a13ed44c578c2ce033c32f10fe7e9492702df2babb0f419a39e71a15e09
z8e818ad58a1db342ba974410eb46a18ffc4dd40c4eb473eabed450b148da32c6a5a590fd79bf7b
zd2d4b40c3c0735ac77fb5591f5cb603bbd132d7028d4222d3c0587116b2b978bca570106ea03ce
z34105d0f9e07a91be2e0a5e5bd912b8c11b1ae3d61c5f3d75705b909a570b6c3a4d515d3d2865d
z8d0b779c965e9d98abcf885c9f8edcc88bbce519d85e9a1df6f0c392dc12de9de4ccb78450ca92
zd374c6fcf2ec15e72445286b3be3d8ed0084bde54899987e73922c1005042998bc795d5920aa65
z3feccd8626aa8baac72cc5e6bf6c333d178ef5e30f0f91510f06a620285ce5c3618acd746ca40f
za733e200907f01444a230f698051bfdee6fc970953c7e43acf5e5c5a830419dfc4156790659ffc
zfc555d1bfb31b2820798bcb093af7e5b736260b846f82547ca4cb3c048a16ee592da350b3599a5
z04cd8f0603024aeed88a8277a9dbb59ede4d61a76beef96c2a5146bad6a66cba1324e640690983
z044b475fbd528f62d510bd01ff50c5631bba277453b5eeaab4f95e90b56b011cd6287682897f9a
zff578c1b0295d80b8c41f96832a1ed71f461d68da0bfd2d8870cd6ec4a506aa013aeb62562a29f
z91041a9b908586f7e9f7dbe0233f097bd9e317f85700de9bece16886107b2b5c5fdd5f6bd1041c
z08fb2f11958a5d0706f2a4f53d8527c38f63fff3abf1cc20e49fa4bb38eba0fac2df69cb2f0f22
z8cee4dc97bcd6a4e9d74799373b4708fd73638536e0b9095f08bf372dec8885c467292ee60ef1f
zdde987f5e4964244765b3daa4ad393930747f808d57f88c3c9c68004bbbe7fe1ee9cdaf82ffea6
za54d81422666f0f29b583c5282b22b43b0ab0d96135165418ee2e521d4f2cedfb0423c061986c1
z0e020ea573f40b951062d5fdc19c170cbeeedba04b6d177265200ec6a69b7c36ff263c08577469
zc3539548681d07b6a327e2fd9b0c9d5dac61d84684ea6f7013d0ea5037c5b1eea2ca1d3df99b40
zfafcf7dcaa1e45c2a281a4adc25e691a3962731a13ec6115f74d0f42f5a205b0cc30876bf153f4
zac575959ba13b8883fcaf7d17df08fa17a196d208e4a7f7954e5f20b491e40aef79191d5ee0d07
zbfb26218853b41daf2cdac4967a0936d73204d6be285cbcb995195919dee47e83d5ff2e5b47fa4
z42399890e3d32c59171653fee470fb1b9758d597927cc4578844b6a1463255fd12390dfc1f06a8
zcdc81c2a452683989f2daa1f9143ff8e68aa37180d30ac63f4b6d5cf1ec39f08266f81f2c56418
zebd17e116e6a7ef8db729f130bd0a8b4016aff0e1688e11e1f735ec3e7d003cd9ea6e40affff7b
zc047dc1518af5bfd828fd36561bed23a2c7dc033c57f5bfac80da38be3e29168b7aa575c71dc4d
z65ad4c39e09706579ab00ae6d6fc98ba79687fcd448b079ac1b0e383b248e493a632229bb0178e
zfd3535d6163971ed0cc724400f1d971543b947fffcaefb949d4b90bdfea2a7d05a6032b084c28b
z0c74453eb63c3f569d82db99ab3bbec328eb36583d9ad6ce96ee0cb9351d65b38b1feaed39addd
zd3eecfa4f5ef5b9e35c0375ea949b01445593c1bee2d9d5fa62fddba67de1f2b4b60bb439c9d3c
z7d04c16e73268d24db038206bd12b786c7455ed73406f31bf10db92ac6113d81f3616f89c38aeb
zf9eb175a6104c02742b5885b1eb53e8695d8d4f939511ac2335689019f99804142d5f497262b5a
z5643146cdf9c5809ac80ed4925a6c9b63fa482865fdaa4ab3e997b73ff5e7ee7224e44db5d29de
z3bdd9b8a0b85127852d521c4e8e56a36d2bff93ff40befd69d93c4df7ea163911bcea6e0fd8442
z3ff15ed7d09e2f47545885bbd1961ae0a1bc040b27418b1165395807fc2157f7f50c6f2774da05
zf4fec6e9b4ecd7ff6518c82358daf4dbb655490bdb502aae2683d317f2c4bf5fab8805f128b2c7
zabeedbe24163d1239b1ba4e7dfc0bcb3298af70ff9fc8b6cc2dfa82499bbded00e5b1a810d19df
z274425f89ef3eee1d3b58508f885f617d4055eca732707d86a56be19812f56c3c7590d8e18026c
zf9b09a18ad454c39f5b1a9d6125da29d51abbc44889fdd99944b300a280a8532cf18db16b3f4bc
z592bd4c9a682afcdb3e854e36f9a2c53bba73be82c3e10dd06d3f00212bc71cad829a29cb77ab1
ze1f426a4dd10395667d14eb2e843c96dfebe26402d1a0a2b188a761c68c2ed21bd0e8e185e8db3
zb5d22f85d664ae60ee86320ecaeb9f9dbc80163e797fc27cb39c20c6e01bef69b7e0cd8b76dbb3
z6b196da26b40544ac63c8ae016c4575277c12b73e385497afee30b60acc5e43ff81823b0f2278b
z9dc2946589cac404ea9403d7714610ebbffd1381fbc4c9858f77624023afa5189be0e4ab4f63da
zf009667b959224c600488a408d0643835662b9b56b621c3c4dce0bae5d64f57a0d77255cc6fb62
zb4d53b95c97fe4b7fc9d1cb75622ada15fc719dc7bf06bce562350450cbfba07cfdd0464620376
zd469c628e582b259213e5a448b91919882b9eecf22de16b3074048d88c447faf1bd0558a8a5969
z95ec54cc952b2c99319e2ab0565517c03f9c20bcdec3641691f7363f750ba6f795f14e8b625fb2
z36f11449c34a4365f4ab40dee236ced89157f93f4e73df4060d5c562184a18d0c591b8ea95aa1c
z0323e08272e8236f4f0de00a9ffc910f17414361fda7e6194aeda8d4b091b9ebb1f21502feb7c0
z23f321622a402f550d9ded2c8f1dc2ee86e12b004a4fbe68bee93a0e23dddd500a1c914b72d7fb
z141b2351fb1f8cad2c01ee71df586f231a3b5f4eff1febfd2a5405e5385e83bc2ec1276108f52b
zbab483afcd690312cea522e8ba91adc1df483ea22ffabb4cd0cab9fc4f1edf10e7703b7bbafcd9
zace7cbb1dee9f0f4eed9c23371cfb3b1e97a0f22d6cbc7c2b14ba648aa42ff414946bd5e224e1b
z1a3c5060d9cff4ebc392f4b922da9c4341e7c80e704964549dfab878b357591c71bba070a9a803
z328c590a0cdbd0bec951708440ccb9cfc8492625155921d6976e382493966d5488ed37127081d9
z4060463a75a00a40f9f1f2062c2aeb182b94d797020f56e1c2dc48d9497362e4b855c59f9c77b5
z8bf7bb88435ada7f15f798c362ba056b34b9046907cb388cc9e9df9329ba8a448cde1849477e1d
zfb7a089b010516b15927ff2146a7e190213dc721cee0161f94754c47306028733b3a7384c620e9
zea4f763f1ad1ddca2cf380cc77295142922f0d02c25d08893afc610222157a0b3d7c2ff6e19c8c
z79af6b274696eec2b77e2c4f0a15190c19998faf302d2538838bb078d52566e257d9ddc0d84db4
z82fc1b2e781fb567d1cb05cf23bd6f55b313f912d254bb200a2b3ef422cdac964fad4156c2026b
zccede20be9338d18b97449cd66ccbf2847026bbd000014af92a359c3e1accb66a2ca6a43078613
z13884d36825ff29b1658b2f80f0bc352cd5aae83b6142b3a3a2ad5a91dc6aa79f7dd702654e64f
zbb1cb41132bde350cb11fd58160e1eaa7ad0e1757053492581a87e1d3b87acc3c4e726fbdf3d81
z6c125e3a2443c31468d32ca842672ab62cf62f6e7c351da63aa7d889319a9c8db73e9db47f9229
z88b55404d21ca4a8bf224af546838b8e166d25ad966e8695e7a359eb39e923f22657d629798730
z2c0184252616dc80b6a574c6f7366dc40eacfa0bb08a8d986a21837390867ba17baa332671255b
z0eaef15ec3a3626c7ad89563f9132a0c6f6ee76fd565dc91ed69710c9f37992e9a3f822c53e450
z433883b3e87d8501a3a8ef3f6d59881b4af51f39853931769099e913f3acca03ad767116f368ce
z6694a6d0e629a9a0d016293db430da8802d5fe9e4fe0e1edd6b3e6ef27371beb12b6049435ddbb
zbbc54da5e01e05a74ecc1b8a3532eb7e9bdb202004577e2ab7bed5a43aa506d2b36c3bed475093
zcad1aab43eb36f32d069a3ff4c08e34331a168ec95e3225f18b9663c867c910281e3236db0ab5f
z93a98e2e42cc82fdd81276bc39b3746ede6d3ee282f8ed472b5a9237333af6f3bc701f165354f1
z1034e883aa7fcf879d68e19864e0579f93feab81d076cbd05782bde4bd13ec438d0b04a982eb33
z76de6b09299ccc28a57f3630c4dd36638209acb2cc441bf09c62db12caeb07cdadf2820659bc04
z78d3bb3d592de45c1995e46e267b780dc9e77040ebb00e59870cea5d0bff0b22a2de4399894e29
z131828277bbc0a42ff7faec1e62f7a822ca2a50c13b6e7d2cc50fde780c07a573e6e37ae97b8b4
z02bf482fbda345ccde88fb9173f362898e7958a805f9165301609e04e83b661fb5d2c595320450
zcd2a8027675d7ec06e509371c7d86858de51ea23fe8b86288dd3118b855de8fa75db4eacacfb4e
zea8bcf6128616663e1c3507c773b7be0c476301eeec68f12df0d627248121d48dea7ead8b44a69
z912d78143afde1d2b27a588864906420519ed82350daeda1ffc1d2a08f19a144f4826245a403f5
z538d9fddf58d1c988116a5c5cce31cc587243f8a7f10715093a589dcea64098f66a97b6351de06
z2fdcd72948ffa23e6c79feb942f6926fb30389d669c6105de54230fe5ad04955f4d0245d6e40ef
z296c3ffed97b56e744b6ec8b99631acd1bddf41e889ee6ff4c6d12066393817e96dda3f5802d55
z75a778a0cb71066fe651a5d2b011d6d84cb4c681ed8a50a335f7c29607462f575e59333630c9dd
zd524d7ffdc8ab40478927406c953ee1a24908fe20c978f4c74e9cb9c61c2b538d8bbed1468a691
zd9a68390a9adaeff617e3fb8770947e26a2e95159690ffa5c6588eb9d8fc061d0d315f605bba3f
zcbb45e4d8e700166a02ee60d4eafac6d057cbae4721205fc8663e24d6aaf6eb33f7d59ccc9f0eb
z5e686634cf4b6543fcbfc6d726f7a7348a46f3d21101eeb8596d9cd961fcbb3acd0725d016f56d
z1fcc33b1636b8cfd25e549423726191613a74758aba0a504ed6a1e1e83a6d4c0ede7ab46845d55
z8bc0e26d374d8a690d215179c860b04035ed6c0a4732b21db27efd1d0db9165455a031d458bb96
z33bbbaa39328409a38a25f9c5903e01343f0db57fccad1c8676ab469df5bff46ce097df39d91eb
za4b6bbe96c435f1aae0d4fc0bdad47afede8b3f9a1e3a6cb612392b04aeb8b8946ce924d6460d5
zd4bf5437d89f977bcc2f115a45cac0e30ad5cf2e4e1e580536d6ecb01fdd904d937a0e2d8e66f4
z198dca1ffb7301c635c7fdd5881ca440ae158a545b52d38e6534af50fe915fdc26c2f092f815db
zdb6f9094772a7a3668f20c3a5671f05918cc62f61aed8341fff5ce535d4dfe9bdc18fbb86e9d34
zbff2e87d41e7ec815e5a959bfef780aff5f25d6ee8ae0a28ddbb18f37010d3e3e96a628feceb86
z31975823c6b312073d1d1bd5e7afd8a312c7ca807fa9b2b2617c65b7393dc3efaefdc982a45acb
z2803928e0f66d684fa5b4441c3a23b7c2aca6ea95d127688600e0089750037360b2bfead663709
z4348b774668adb27cfa3ef2c06f123b7e66ec0761b5a6fb3e86a46d28215ae44ded9bb2bc3854e
zbf1a042033aec26c032bedf208f83ebef50d6dba8d990c5eaf62c2d19f81805503af22c4547678
zacbec23fbe43b7354f3f285e6a94d8fb5ab55ffbd2bb5782a0482cdc58265e4d06c0d4b0570e72
z164f3d0e8a739c929f8d30a6913f69ab20c8fa5c97ab8e5edcd2459afd73e49e10ed8e4fbbeb81
z5f31c58a2f293d476bed6e0a93bf52088716316b8fdd99b157b6b9a361fc6e34cc79fad0a5a8fd
z7e8d3c604a5056120e10823557ab166e3cdf8db0bb6b45d3710174ddf01c5a9255c38aac8e5f33
z199ff064b801a292cf7afd2dea0a86adc689ab6460c848945a41479795fc3cdeed3c57bae1b748
z73e684dd7130ce057c67045cf55a7f3f85e9de2ea958a00d56132de0efed3671e936db229717b8
z371588462c6e2e8f2c0f76dd423086c21843c1ef7999b22f0233632de8da858f832e7b37616b32
zc891b1c58d28ea1dcbe503ec14be6d17f48fddded7df6be01a27e6044aeba78ecfa6bd577be47f
z116a2e8168071de41d264bd6064ef46cf377479263eb6365dd76da278809278f7ac2e000ceb6e0
z9c2ffdafc97871b92495173d7bb7180c2945e64bad6d959d179c15eb5792b36b7025722edfbb9d
zc07e23369030e839cdfba5e974448e6c70b82065d192e689695923c4db0bcac9b7e2e81326b1df
z41ac3266a6870149ff9dea0abe3b726de17cf7baa5723da77e64896f05d8a75a3ec131f41da69c
zdf5a16e63f6ffcc40607e07ec6b21fe9bd78f24715b02a84e3161618fda13007f8a337e5608890
z3c2937b849ed9756e71568e2660931edb3046dcc1296111366a040f4ae73f0b93f9930c11b2ad0
z86e4ce2fc0ab0784c7329170318657cbdc02ac14440413d4d5294f29a0752efde8f43cfbd015a4
z0e3921d8dfe520fead9d9d672d71bb759162810baad3990b35401114b0a9fe9a6d12c99b138cab
zab10fe359b8c9703b15b0eacb93d5c1ae9882def8ffd01e0c29dbdd208cb233289bb9c6d0f1e8f
zcb1161e98e28c48b239463d338be4f16adbe304f0072c02df5a2161c50a462348474637dbb51a1
zbbda51a46bb3dce5516da2dbc99fa61ebd6d538797bea0d7294947e126e2d56e6bfea74e430d67
zba9ea87d4391222279ce41f8f16f788b58459b15fc216edc6b6803f242899bdb8b556a9c1b38ad
z6d6b30ebb08889f3f2757cce2cf4e498278d219e68af08d9ef1fa1104962d564eee82877682237
za9b2dadb292dfd3c7ee152f29ca61205e9c10e0f4f7f83567ea525ba203ba4858a1548dd7c139b
z2e5102347dfbfa9cf04c4e9dfcf07caf4d02e8d7c122dd0b6be311ecd34607f0cf5adb588fd6fb
zac59151ea20bdad8d9c2ce7d0a6f17af541d01f8b960348d7dfafb952869d7221f4c8643f1d5ee
ze35588ac7b0502f4ce82d20a6da5fcc072ed91dde783ab9bc4e268dbff23728650e9c7298933b6
zc8351a0d05a0c68bfc68559f2cfc401487e73558c1a320e317f4408dd73b884b7f0200b576db8c
z3edeb95e68fc731337021018b55938d68fa3f4055dea809add63dada5d77f4f0b5b190e73abf4c
zbb3e6ff00fa4805f4627e004e340d03387513bc1f80fbdc83ae844f21b3c93b28db116d7280d63
z954044751d89b924306a3cb3fb6fd0c5499f08ebb7d4f120599526ef49d902a5dc1820d6fd9406
zf705c8f5d2c71f524478bac5a403d659d3c08cc8e9c502be79679c9c2e030181190090da0e9008
zc6ace6dc2eb567f52ea06a2671d17d72fc13e1173f2d98e4b52708cb10dc00557c10d2b274d0b1
z6aa0be05b76fc00bb1d26c20f9d98a8420321edde579e7dfc95074af58018f98470253b65a4789
z0c371311abca6bd775d15c546251d0113d7eff17f5923b91f7b5429f0dd9b9cabb21d91c7eafee
zf90cbf5f5257cf7211855bee5f10b9c6472afdfd69e1dc0e27ba79f04af2f655566d7077c69b08
zb5b34e16595203f02dce429c292084b7286d6929ff8ca928a0cf9a74ab18a2737f7d896a6290ca
za3fb6b4b81e0899470e3e068984909a90916e57e65e36b6d6be58dc53c4de7c66eb5b1a8265d45
zaaef03449847304ea333c67efa07385b833419836fb864fe9a1605cd3faf15b766019f4a11cb14
zb89a61835b92e0f4e285443b5ee539113e6fadcb8cd8b2c1c99661d951ec2c16538575dbfefe7a
zb8af377e074d948bf3f9a3679b5c9ef3ebe4c5811450e9089dc28f20187208dfd5d90ab52a5f76
zae942c6df5fa79a67abf4840ad421e1bbb8b0dbc3bd11c233c76bc6f194007b074357dbe92baa8
zaa94cc4ca268a9730b2127d94aeaf4032c453f83c41c1a742b422b53c0bdc6eccf1b2d6456e946
zca6d4d713cd04135282b99351dff6a6618c19053c30ab3a3876bcdb8c20ec68eaf67e5cdf44993
z62747fd85df353b4c517a6698ae3a61d8ee415e4a38a04292a3b52d6e254d6c0099c253cd9cd1a
z796198cec6d1621b949c64e18f8f29126561a47451bc9d1518f56bffc1e4241e3582fcb3e19b7d
zb24b2a36353b7461de9e0e47ee9a7449efae4e7c443cd9c422fa27344c7308f3aacd564fb2cbe7
z016c6445984c907c33fb590eb9387439085ce8b2fb7aff0cfb618cf90a761ad4929ce6a716416b
z4f6e24c95ade00258b22e5fce8b527f8746772d42cda9bb89abee400561dc403a688fb1e1d0403
z6d27723c0bc0fbf271ce1ead3a167a87c122021211617ab41b2105ba327d107ff9933f4e8bc484
z94f928ac2df87160a8cfaac321bc0e74036660f97a8b995d01034abebe6238acc7d20d3cabf67f
z0625d646fdeeb597a5a40fef8ca0ff7baed1cf59f41f4c3a81f4bd1d779b3fd88a3bbcb9a1dacb
z78c09e40c2247f56e46e1187518bce55ec7a8166112d1a0322d1c1dfe190d792db403648db6951
z0fb257f96b98eb0b6fbc4a55a9772b511409f1edcb6e674fae387353880315b5efdfc8b9205309
zbd12813412010f5eb836356c41c010110f8b322ebeee45bb1c030a7387e37d9939501d62a5ea6b
ze5c7be5f204974891e131857a7464a8a07e1b2c688df12d36a35db4c315ee95ddeb47b1e31bb1f
z260f7c3a4ecc58bf128510b32cb8c3b51613d474c1b8da8ae57b1146d91cd3b809cc56ea83d003
z6a8df31b7bb291c3a39ab0db78e483b97d3f290252ac65c556e5aae763c8bf531e4afb912baac1
z34cdd6ba0a18532706c76014a2e0c4ccae118c554f4b7086dc6a146e4dcbdedd9722d749e4493d
z5359f236a4fc7e1a5a68c167e4cdaa310b414ed4041cedc5f9aa346fb22c58947b60f6ab53b1d9
z5cc5eda6418bd1ac13ac5301d967942033102f8b15cbdc183b0cb95203c06b3f3046ed90e4104f
zf544f0c076930d7f3d01510ee7a1382563fd6dcbcb49334fe2cdc21ca99ac09707f1e3abdfd6ef
z2ccc48d35a1307abc75f033c9e9b7add7fbe565dd2dd0846a5842df804c9ab33c45964139c74bb
z53e1c0fc94caec0a12ddc66faaf8168ed48f142f7789e5d06f6cf008962ab1db202d1c839af411
z3d8d9887efccda10add45b12426e35ed238ba50c9eb47b920f6aadbe0731d75d8911cd2eef6d1e
zd84ebc872e1ebf042850476412e4d56009b257f05735764945db49556398ab7599fa578796664a
z1827e9f392a8b58602b8f252e9469eea699d44e754d427101af4437e5f97210f1d210fc12abfbf
z234a19dfe030577968a0889a0b151aede5db99bd36bf33a6548bb3cc7fac75aa6000e049fa3fb3
zc7491bf51eb5e564a24fd46b31d8d7c0f41301033cf3a41195db5329ca110a2779021fc06e2da6
zcfee68ab0e2752d65808478e2733348d830742efb583968c3bba38d43915109e71741879e8c775
zc83438c30f5c1a03ca2152715a7c4600ffa60c680a6513022163eb9290c731d12a44bdde39af7e
zbe6b35393d5b018ae139a906f678471c3f0653d412dfdbad08c470d0c6e6b47fe69a00c4d31fbb
z4bc541130633ef96500d9aa9f77c8382523e868c71b80126e2c2139e2b9f82330177945f7da6c5
za2e1b6a3f559f48a4ff953889ff53bcee3738bef820245686a597aea1b7422f6ae75a61409bde1
z3b790ef5ad21f208cef63ec1014c8da5c749ef3bdb2e1af8bec0d185435bc342d5e266a60bd0f5
zfe1eb9da57ffa0289d9746c6f1876c97f3df2555163978081a375caf87a0f7b3c61e027e5b43c9
z3db72c551b3afbbe3484695b24643eb126b35d3669414ba61fb2fe578165781542d110856d67e8
z0e9680892cf934d948e900e3e125fbde414b0f2bc6ae9aecfb58f1eeef3503ddb58d27278afc87
ze29e0a417cfee34f6629e205526b299589214309ca2f22a9ac67b77aa16acb588a3619c8ababad
z1f52c450f9c6d0ab757df535bb01a29e36b158ed5dc8a6146f6fc38c451a6dbc540f5626654af2
zc4380897e49ad848a0e3f8a57e364178b1f6fa9b0de8d5af096818b36795fb5ae69cd91a5a6306
z4a6f1cbe97bf24135a80938c9b77e650a107d9a067642d7f4f1f364cfb3a3367ea0761b634c25f
zb9baaf8f82bc6efdc6ce484da2d61e21c8edc802a5c9f787f2b50ddb7df36292109729abb03c32
z711f59c734c0c5d431d0a4f0a22b1f3d1a43d43012dea256f8701bb4374c8dca0a377786c44fa7
zad60e769c7bcff8f012349b3d27e00cb913f686a9662d56f335173b1a64158569ff0044a85823a
z5d9660314e9605790ac45f8b5cfe69ab06821fd74fa1f75d31efe28a0d874c96347bdfe5cbbd77
zbe54ee718c879ebe30631f405e03d429ac8d33656d4c5a9ecede9ac472147fdd04176e278266b7
z9f566404d2ecd9d351b4fa0382470c3bf46060b656e9f9563cfd68667ddd5574f37d04a75ff10a
z468ce3f321ceb800a11c4c441094e28f42f4d21daf7dca1457fa1e1b2a7563ca1db9a0ca0f4d25
z9c8e9ee663636505608134b298bf5075d0cb195a40114f80d54b20e78036983ea70ae38d63b8a1
z6cc51a09826b98520f9e4d70c82b0d9a13ad57a0872d7b81bd1034b2f51e7fa7d3c638baf9dce8
z19371165465e75f537bc2d87c3e9b8826374e1d1efe8cb941b736da3fb926564b042b6f77056ca
z0f97f04e135afd91ff02fc4f47ee5c90760f19d74a5bdb10e330f494062637b19d407ed8f161dc
z08a27b198072b8c93e34c346b3e4dee27d01d95d3cdb6bd71fa67166e87349ce12e4c4f52e8eca
za2210c6cafe29bbb5150fa0bccd764a85e21ef7d700645b9182fa0cf45aafb1e23cc2d3c26022e
z704caafd154d3e74ad534ef36559c04895e10e21602bd739ef9bfa7180d64b00f6241bc8d4e65d
z27fea884d7fc006fc633b0272f36e49b749165fcf12c831941ab2458aceb56947de4d65f4916f1
zcfdde1c9b59d7daa0668bafa7ec18e96f893a5461a7d93a69c6f386089b68f8d6496cb309fd020
z0b653eac26fe5732039a94913159c22d5dd710b76592d140fbc0c9e5bb64bcfac9711477c4e2be
ze6ea4de3f313d17c2c4bf6653a94a1729736be0ae6746804df556588ec87029d66e70749d787b3
z85cf0600edd420a13e98bbac3cb4fdccbfa65cbe69dcb78dc2676fd71f0063b74c288e2ba2ff09
z0c789bb5c9d520ef59b6bdfff2dd7a4c04f145af9d98366304d0a9b981a15c15fdd8f4dfa16011
ze83d7cc72d10ff03c33dfae9b6829c2c80954ccee57107b3c217e2b7f87ca72ee7d5a0f05e379e
ze2cce8342e73487f284ba90c0d4bf80e2cc537e411b2fa2e8c840ab63339bbfef7f97de31c69b5
zfecc7e17a3c44f056a338f2fe551be75a29a1c2d8543288517054f479d31b72926b3e1510047d8
z22272075b903f22f7ece74c47cdf089f8c19a9f3a60812685a7ca3a81d96d335564d495c7574a1
z1a59239f435a18fe86c28677f27ea05a5ae522576746b4906665e9dfb14fd17eaa49a26584741b
z38ba832a5fdb5bbb18005b1c5e8fe8fd7f6ac95d50f062a512692041ee72027106c6a1e0328a0e
z7d0d1737776bb33c9ce27367d75dcf10763a84a5895f3c5788ebc8f858b15e8cb1a5ec29c354f2
zf61e29c1fdecdf9448d37e3bb7e40b1628c5f42f2d0301b1e2ebf44fdd5f84580c6795abfa594b
z4a47b9440c125b746be83a96179c28278200941abf01492e08f75adb991222723e670554a37c3e
za5b7d342cb83699e4f2916bd0528073bb5f14ea90f229eee6b48d7f15a6ba0fe5cd5a8baa15b2c
z48efbd747730d5f032d71a7a0c6d0f6df1e103720d664dc08581841b077983f93ad6b318dab17a
zed40024ebdb706516455ab50d9acf88f23662adc092e1b27df1fdbca34ca7fa9d067db66900954
zc484b9e4675d44e627b8f0a05dc922bc720f5bf3183fabd9072081b844af6c8f6d3a6dd337c2d4
z96cc298edf1ebfd0ae65949e0f751b9db9ffb7edc4ffa0090599a37ee9668f26541b14b8403fb8
z8b9150ca1710ca7eaacf58de68231b6dc30593c3b131706504c0639a9038601db3f7c80ea52dae
zada8813e8fb3bddcfcb4c0b9b8a82683e27228d68d71bc3d6b75d0747e58e77f224c4eab9ae250
z0d15ce013590273058f81e7380ad315dfb8ec89ed089fdb45e9d8e379dacf3ba6fb96aed7fdceb
z7c49400495e56fc66a16ec1f694e115bee06246842ec5b888b5466af384dab79b66c53a7270491
z213118d4ff20b61e56c7d0413d543fa9551e
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_bits_off_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
