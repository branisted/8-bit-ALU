library verilog;
use verilog.vl_types.all;
entity mti_scdpi is
end mti_scdpi;
