`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1bc235c2ceff4f6e3b1ebe72fceb7af9adc96a
z694b4bad7241bfbe775016041d7caaa74d9c0e7b507ce89e8b01980415bfa35a8e346f54c548f9
zda8767c02ea87d27eb7a843f4cada7dc3b575fb5cede69da7a4701b2d725c73f1f7375e85a74e2
zdeae70c30f1127407402c955b283d7b9512dbb3cc85aff97f613d57a4efe57b3c092e5ccc5b6dc
zd01018bef01fcb6b6afd138be37349905063433d6fc88423f78d0a5cd8c325dc906237be6d3673
zb87d9fada90e2c892651aecfcd04caae277f299df76d77ce870132e5e40888bd3b3b1b6bc6e799
z48a23782b89d176bd848937c64ea2b6938c5a6c2c52409c3721f00cb676ae49dbce756d647186a
z2d5ecb2321a08bb462a97b513b2f2f7e1913c836666420a662f742f4dd090636a3381f28becec1
z1708d87f1f0a00e76b7fab8e82c4b58a7479b0d3618edbc64d306b42be8b9498e21a252a9f7760
z4ddccf620c22105b64d3442eeae29848475b6321275c60da85fcc15cdfce58c0be67611b4ad217
z85faa32f1a391d7896ecd2d6a476653f33c744e342ca0bee6222cd817d247928bb48ab87008585
zf4c934887ffb02320d1f5e9901371c546d07491c6dc0560188ddf7660969a0521bcf06899960a2
z846b97706440dae0671d4d93134b115147c7d3bfbfec814d2c532f2bc7b5a866f7796e878f79fb
z6352953b57e9db9e47653b1e11547331dc0137729d159986fd727762f733f71a51abb4c40cde6b
z54c31bc6f8d22c1e7a4b1496d59e544c58c7ac5b5c2afc9f78545153e5723168b76fd133b724e8
z3403b93744942c53afb201e1406fc7e4fe912f4918f0a983ddc083038f980472dbdf3900fd6334
z69ce561392f33f021ff6ab00c4f53c57329859658e8309b2ff322d785bf61240a5f851012cc7d1
z8afec9d8591fb118ec963c3fc41104dddb3d49da54baaa2055a485bcb958723a588d00f7b48f8e
zbef4b52b53cdaa25201dc441b400e15b450affdae195606877ef954d4bb29bba7ad092353b7a64
ze5503fd79281cfc72d3d8a3ee6ec684ab92121a9c7805b30f46e6ea2c43acc01b5ff3f160848b5
z5fbede0d09022b87b348d1f6e1acf47a160208a23b68c990fb377020a462872b70d15ffcb240f5
za78e430e9b871f9a17274391bdd635e8f86d34c1ee0f698211b460f8a6840c79dcce551d97a78d
zc7b58fbe08290665d04108768f2cf2bf5c3bc6e99a48704ab47fb53b068ad52c1843972620c4cb
z33daee1fc20cf34cab86ae881c6b84c93b5991296ae91ef9e375e5221aab981cc5de17d35532d9
ze3a41038258c5fa0c8d376f4db6c18936deaf16f14e17d594b1c09f09d708b6de50dc41f699941
z85aee06b6af43beaae31b79f046b04e57bcd2d85ad910ebba795b3aff7c62a2cb3bf7c5b811653
z7db84730f63e4511d2020d2afb54d02244527fcb7c686d8694a72ca2332b6f01704aa3f1f59960
ze088b00201620f1bc676d8d95c8dae99934d8c1f24a1916298f6863f1a551cd1df8c6ba28ba1a9
zbd65b0cd95cffbbf524676f9ff6d0cd234a5742807f3ec9a4359925ce462918ae1b0272768966a
z3314cb46f7d520f17b04c6a845d9782186d990eb399a8b4cf0e76165fa06fed6187ab16b8afbbe
z3bac93042029ababea86e2be90a65c9ccb1b6d0e153ec1ffb70cc0f01890fc3dd2e9f032ba0073
zad5660c9d3e90f77720ca66df61ce9ffe98f0f13cc4716f2b244eb333a1a672c7085a8c50e7c83
ze86e81b58ef32b3e7939d99288c4aa311b399cf05b2b437bf14eda36cf041c1010dd86510b6c94
z8da1d6e86a114bb6d6202c83be0e5672c8eae6e5f170094c14a69a6cae0bda706389bcc4c6cac6
z776517feb444c969e84a3746673d40c7a05aee80ec79612ea541edb8ae765811e685abd6bb8f18
z31f87b34871c6abe98ed51e344399c48099126bf7c862c7929d50e67b97a603e522281a1fd5443
ze4d3e55c51108b084d55c3cd29b1cc8b4fa89226438a83462f390c3381aa9860780b37992a47eb
ze673c3e2a48d786253938787ef7e05884f7a83f0dc524d4bf0f9fac24798101671ef26cf497ea8
z251591990310132ee04e5e9ac9cef8f20c0a7a354f95789bbfb0c34cc6bf10f9b93607e0c270d0
zf717e9e669dd4c1d93db0219c1efdb3266032330f0d96c35586381012cba3ae7078c7d560d7104
zd546e29dc3ccbef0f03a41c4a871369312634a2abc94c1e7e5a72c62dd7ba2bfdc7022b81efdad
zf9fa290a9b27109d6266027a683acb65b30cf777b5929aa10812619131281f41a92877c1f3c998
zf23320b1011c7f75e8583ce6fcb3ef3e545d4bd97e5bf1178991eab0ec1aee756dbccb3b714f3c
zd22d01b9c1bf5018e86bfdb4cca25a817ac12a96dc2199aaefbafc1525acbaaeb38c7cc82f3382
z42b1d3a17ce593888e4212007c512b4db4353acbcaceac252945c510bc9453fd4789bf1e759f0f
z7cfbbe21759fe406692a24d6f3947ad0a2567754d4b66cdb79b5a876a7d0d0b27acc9d5630cb5f
z33d21b79341f486629164cd04ff2c0b65cc8c7c873c023cbaa9221d6e851b91e0751f9a51f6fe4
zdd2e4a1627486833d54e37fefcd55db57f1d3e51d2b8e3c69caaf3d16142211be8d732625fd36f
z974045efd8f8eaea8c54b0f7a9ba69687ebafc74827a9ac20bfd97e014ae78074e09d5adcf43b1
z9133600700160b81eaf8e28a45cdb0bf6219f0fb56d20dcf86e7edaef89378f76e181925339519
z3e289015bb06f156f18edc0535aae903b8135861f8b5f7454bb0d994dc1c394181e3054ea6937f
z71a2536e7162149fd13a6b9bf6e51c3f43f873d48e3ca9b65baa5c4b35c42501a9f966dfe1c1f8
z1365265e4d04e7daeb357f466532031038004eac07aabc16ee0176e78f6c3b7ab98501d8e8c55e
z50a7ac4a994714842f7066bba7e04db077c37bd29fc995479d439498d56176308b181b6a55e27e
z3254499be87417ec210b2ac17a651d6125ef12f816a70cfba3a94d922d1e2f04889001fc1890b2
z99f9d304687059269bf8ce8e0b8fb1b643192f604474b7929047e68c30272e1d547b0597de4de5
z364a485eef516d3a65454c9a97902ebf6bb9207745ff94d5eaf285ec9a6c7f652513ad6237e4cb
zb0c03d11e0e413602dad47314557733787fa2d23bb1e4f4886af705d87a55195819ba98592ff5b
z52629bd6b7645a6cdfa6b1a20728c4b2af7fa6c912b6347a526b2576f6d3e2942f8284e64c3197
z56ce697cb4331ae2ac5d6a4b06beed6008128cbf1c3392ffbab85e1cc74d609c537b43ea29db04
zc95ac612d4d7f741edd5dfa5a5e9303078280bcdccc2eb5ad86579c4e9d8b99e6e078dce990a76
z88429fc65f03b5700276bbe7c6a21959318e430461950b03e4b64df2a894ef4dbd9a3cdbd386a2
zf1387698ae9f33969674ad8d425d200bf25dccca46711cb771a23503e1571ad9b2c629ce89c092
z9d19ec2e4b8a4e128cd1f181be75c27769646607549bde9f5ca34acca85e74d9c4f48c5e71ac1d
z2614dd5e1006feaf9f4f30687db0c0d6910ce20a87baa9f91f9153b8552c07b27f8ef0dbb17d57
z73be9f7486529cdcfba6423ab16d4f47cb6c9de375f78b9654ecb02fa271e0cd58bbbed7494dfe
zc2bf47f84514d9d7afd91b715bf7df350d61f6a1591fde752342b1ba9e40bc586337f462ac3eea
z8a8430c27d8bee4b8dd2ace22fb47e993320f5eb6f69291411f90f07f0e11a10ce6e8f77888d7c
z10394fbe20acbdf25041edb03ef6d7860359147a31d9669013faa47d9557ec1ac7a5c176e44607
z31e25094ac63a5b076a1e772209ec1747145b80ee2feaa65fd70a72a37b23cbcd7675cc8151c4e
z01b108e041e6de032bf2f4a5cbc28d52dad64ea7cacc10a99652b8de488894d1f320614a322597
z0ccc8aa82fbe2b222e3efa625cb9a458bb96d1e8cecb676e6506fd65b09db0c453c228b5ae629b
z88161a720598311ea75feca8054ca867180b0dbe47897a731b08230e5d1de9df5206a06f40d8be
zf60bb80fdabbfe1f8bbaf7a7a01dfee93eaaabe62b57f4c9f6fdd219d85ae596d398549262b0ed
za55507f8323fd4c4480d27f003bb83145b008b70c834aeab42c39c1b5ddf7751728a352d39f52f
zfac053f3e0853a53e01b49ab70f6a9e2eedadc404a6bfef4a2b474a8735cdfd5d1bf9878ceb4a8
z97aa63dc5264c39a4547e9df46eacec7167bdc8ce5e523bd01bde2647500b983a2903b5165f307
z7ff9108db0feb30f50f24040c7c92dcd067cc951ced9d8474f9b342543846e1a70b6214ae23c48
z7702eb20e11ccd8b9488514b8d81b977fdd000537805d93c6bd2439c47b735ac9e4a1c745b10bb
zfd774df1b19dfdb8d7a9d561d4e54a8842582b80475086ab36e0c172293b76d8076705763ee1a1
z6e940a7cd030b752d187b2d2d23480dc0d2a7f0f1cbc4048d85225c471248a20185444b6e37dd2
z1445aed9d5e331eab47bff8b052bcd312e9fc4d0d8f685720ac12bf69abe46eb160003513be767
z29389304d3dd8fc331dd875a4b7be8454a90f4ea54c0a376bc6f02a75b63aaf0aa57f5e887c597
zbde69fc74c68a5a8dc2264a830f4627c81da0bf600599c8b336be55db4caaf2052b0bb74beee74
z5ec22f9a41c9a8b3918f48ad52ed09a795193737455b40c307c0aa7a95c28ee345e4f0c707f0b0
z15328fa3589f2c2f22640fe0285b55f29a9a13ad53b52f89065a4526a3ac4318a4c1e15b1de380
zad63a3d3637e00aa18bd2cd8725eb12dc0b0d7553fda2ad5dc74a597eb7ab39eae507c9e9f2804
zf0df8a67b0c80c5461465e875aa67a3dfbbeede089847a613a4e99651f03e448ec4eabfa94f3bb
zb5fd691763719b043bafcaa18f7caad31e19976f40823e1d979bf29ab4d486e2c04ccc2d84cf81
z5a664d54aca548b090258a9bf752b4ef57a0c62aa052d0a84835376b585e17d673b13ad9b2f591
z729c5089449242eb30c432738226486f871eb40cbd17f9a06cf37440071c96d37940dfe3743a1c
z6d784b76da154e3b0a2b2f1e215ee49c27fb3260ea720dcddb77993eb81016f72fd317eb882d5a
za81db32998dae3418ae855ad9afe9f5875904e3271792b13fdf38d05b3307561ff5a73b4c713a6
zaaa6058f77935f310fbf8009f8411cc8c159f825170f48be2d53a5cdee65484302a0731ea34258
zf32df1c0ec6dbfe8ae7eb21087df051facd5e7e90a9ac0fedface5bd6f0cb60e972b6544f5f211
z6941dac57ccefca397ced092ec7809e1a618e3013feb0f0c99f93b60d60600ced1a5db54d5d118
za76deaf86ec8e69803506d4d082dc2ee8ba464f25238e3b57d863eff261ab72c292febb2eabb8b
z6ceb5596a26895501568f1565588f0328d7e9f10653a9c50b681fab7162d1b9e52b8e9ac5c02a2
zd00663cad9f3151a54d49aeea5521f6efcee916bb958add028c42e1c1443ae94f524156c2109e5
zfd0d1c773bb6bfd50e0166a37bf716a10afe24be40d1bb35cf5898097b04994d6c730406a6ea53
ze059ed847191b308c7c6dbb107f5a85ff5817db1af724369e27babd86c8722d380e43d0bc09681
z11276553b655bab12e80a1cc3c72b80c0eb3d39d2219dc5d0d2e661ce4fbda3089d249d85a948f
zc119d2efc392806a55dd82dbaaf0dd770f5f53cd0139cbf60ba2a81f0114e6fc961ebc1c0dfc61
ze321a1a83cc808a49ba3caef14b3aa765e0cb5b0e51862d0d748dd435e65b23134e5d8ca3a288a
zae6ff6e46b355d07fec7fa28fca43f3d5be3d653ca01bdcf6de6ebcf286c4e2e907b3290a13d34
z2481235ae8b2302ee2d9165f9d8140159b32847a53afce76b9694cd43fcb2c26c0cdb3c4a23bed
z63520982db8f7a74afec72c825b353adedc410a5c8be4767ae25da00fa335d28f4f5b45b5c9fdf
z69086bb715d787aec0f0d7c6ebaa1f2e8274f03297d74b0dcf756fe89f06d0e4a1c7e6df643b3b
z9c7e8e7b43e23c74b6adcf9d924bc725cdc451a01b978511185c0d3d06e274fc224f69853bfe9f
z09e3a707f14fb3465f90b81c920c428e7b06cf24b84cd9eda69869b23111a83334bfb1f9554177
z2144cff84f74e236130228f0695b814ba06c60d4b09f90f9e94053d97d98d5125ac693a2349af6
z41812ce66c914d2c45b53bb795e6dcd11ab232a657921958541dfe9b24847200a14d7e65bf2018
z9571637893b075179fd0b088e6925fa8ff3a0b649e03bcf0b5ae1eb7b1d8ac216288cec868356c
z1955e5c591a625b1b456164c1587182f1717d0e4aa69840847cee9c8083fc4ec86c539f320fce7
z41d4e4296a5e208ba7f6fc5edb8722ba8fd4e48376ece6fe6e146c9c892e499e8afc18594142ae
z07db1e9bfb7af9704d9314f89e7bb919048c48efb75a79a927a5d0ca71ad312aed90bfb4fedbd6
ze33cea8bef794342c69af1311504d9826fdc439eb7e26b77ece857d04f1ca62b00a5657f101f6f
z5bd4d49943b4ce4fdcb5fac1bc723f99e49e5dc0f89d7f966d0110cef62b246592cc189ea158cd
z02520fb36db8dc57c6cd0f003a650be24e3964ec5138826156e55eb0dd9b890efa5ac6a06fa533
z1f769a853c2f977b464fb0bad9134eb8f8e4ba3ca5ea1fce676235fe80b457306e62ab419ff6f1
zd3dc22c66340121fff4f28c1d10b856ebc2c5e29afc996bb35b0c7e81d6ae2e28187a181ae8783
z8800156e8e23c261493b17bd1fdf405534c489c91f6e013bcabb5b1bc5e1518fc5ffcec563478d
zaa7574f980dd3630db747a11e115746c4aa694642673455c6491511378de8cc9de90b895c9e9f4
z3f1eb63401bc2140ad577e614a5c56689223339b359251deef423f9178d180cce04c27a83da376
ze4bc71caafa6a724b0513388ad2d1c2cb93e60764736dc861db0720d50b0ec7d78f73d9a3e30ec
z7dac39bd42be1276c5a8a38f4ef7347c8ad608db31df8cade3a8c701f2c8dfcebd3bb1ff8ce2c4
ze9c379bcb069c109232b1b9a6a1f6d48f3e35d66e43b53dffab39cd1ed4655098c5102eeeb22fc
zc8008e8bce28ead56fc99209c7f8e954cfa159442a74a5c4d5ed46d7880bfc7d03dfa8d7c02eb7
z3b73341e6ff078c5a18ced7b06861435cf37265ddcb9436c06633cfb449835d22f93790b03a9f9
z7830f7a2cdad1aaa0a7b054dddee8d6c09b6820baf35a268d84dc86e6c156e763ce13075ba6e9b
za163a458e55d59685d67541e4cad17429c5ccea57f9ba8d1393bdf23b6b1babbdc9196a5947198
zd77f6170deefe3e247823b7ea3d8b08047a0d30637772a5b61506008de821525e1426cfb3327a2
z626093c1fd20f8c57116d261113022af6d16577b3271f29fcc79248cd8e33fa214ab9b93eebc8b
z03ce6ee762590f5fb1523dcdaecaadb5a4dc97910e66e4fb61d0129c108a192f57c832cc02dfb2
z65b2270b5a9211dc7536913309dd409c0871dfecdbe6bd439267f34c525549519884f6c541c9dc
ze1e502a7de7a79e52bf9e5f1e660d452b862ab77ff836aa6d9c910a77103ae782d20331b1f9421
ze0c5fa1433687a4f361256e5dc978efb49ec8565ab0902ea7328438f28da64d72d6d3b44a296c3
z15f7c9e0cdc36e89771998f609db43af4fe9671494c042a6ffd773a5dbac2754c8cb3201eff67f
zb072650985c31593c45b34c77b98261477af2aaf8af17cde3840e86e1f8e80ad4aeb5a3ad3d2b6
zdd7bb2f9735df0825972668a6f6cff70389b293fb24694af2979dfc0b0695d86ebaa1aa390debd
z29e26be7e2411bdf909dc3402e1577d7969fc9db5d49c9019f1a76c20aba4145cc907609d3ede3
z5b7b518f222ed5340441ae17f3470a94a3c4155505db985e2aac1977d97784cf081faf3705981b
z9d1409ca1781594ce67bec32ac26cfaf57df7b2e13cf680e68495528056eec62bf4b34a94382c6
zfaf2cfbec8dd829d0bfb58723fd7d87afa62f3e53b172e7e29cf96b4275b7282cdbf70fec6865d
z3d0bd5805b5b63c8084fae7c6e20d67fe9c0e8808e9f4389b5b9cbf862109bbcf45e768325a816
z742e283c9005ebba0d1ac63a06ce06abfbc8910e3ea5cb4a850521feb37f8612189821c2c885fd
zf8032530b73103fff19094e5412d12316b1747db70159943f66833fa0e565ddf0690348eb2dbb6
zac7960306027b257d7f4e198dec161f5691a77c567cfcd884c137c694df98af838debfe5a56d24
z7a51343ff077b2debadecde326b0f633d875a69626ea5b49c20795b47821c1e5849f24cb4a8e28
z8ec1945bd57235e8208eb40d28eb976e27e0ef4437cc1162b9e3fc19300fcb9f2207fd17db54ad
zcba447ad515922fee08e5433a58d4f930a22c989c5c8cef463b2728bd33fce26f436496f9226e2
zcce255c67fda5acc90e7616a2b9caa59b34c899a78eea6af1f2e082c5e8221bd53a757f3d9eecf
z95ab5d8ebe3e84a1ccd56d6567731db6d8423be7e23c64623cde83988c3c7ebe961f8bdfdf4f67
z380fd29a4df72294e8de90c2d461acf8884ad916f5be291c92001d1ff43a6883a521947cb2e82d
z1e9bef1432b96f3351f8500a896f55897e57b0dbaef1c95546719ee76b6a5ef3d5eebe50ee5fb4
zd973652272cf3c56a6411288e92508d165a379abab483eccc7a4866a433d5d47336fbe30f744c9
z2ecc4ab31bf99970c42dad597035da1cbcb764bc95001fd949280cdcb3d949192f2f1d2026e260
z4b078797c3a9d5f54d7ceca499bee03b1cb3988616c45eb06860fea205c6d60593500276df09c7
z6d8378d5d523e6fcadbc1ac5d577b250de967bb760cb1dbe457b761a2f24c59a5790e3b2018a12
z80952c8bfb9e2ec5acd155f0e13c60d9d587aaac9a6debf0e2df00231d4b7ddb4bd742ba527b7e
z8bc1a9413034d2c8e487bbbb38c3f2118f30cfdaa0d5a62119d106ac8c87d7d9866d6ef693ce81
z0be688b3b5425bc4f612ed25d4178c8cd75c305e81949c925245809f7ff3a7202813a4f9e55b8b
z4e10d47930d9041b485e3be78bc7489b90e1e2e862eec62f771c235a70e641201708646ed16546
ze0c3dbc230aea02289b79b590d177d33a18ff5d962da3b8c11793b42fbea505e2c64e63c0d50b3
z9bcdcbccb55e6e9dfa8e47260a06a627d402373562b78c057ec3b61679ba0d5997fd82dfb0e453
z83c5028dd9693f283e3dc4f9376c37c13fca6ac44c49757060c1204e99b657679588d33d5dd6f4
z12bdb059921e1d8823ad855026b66a327c210980cc2ae32a3bb11f4a29263f89ee42bcab6dec0e
zec49b54f42aa987c7c3301ad0bd4944f94b369bf035563398a595b98e939c4aed0351bee120005
z76a45e51af7c9ce38fb050e3ed049fdae8c77c6ab87afde6c91e6da6dc19473bbf095cebf35ffd
z3ea2edc81a731e74c63895ae4241f7952a4f4329af404d71a73503711bf8fb518f4a89c331287d
zce8ee9f4ac0e11a58e06667ef2063ac1c29cac6111d3834054a2ad33fa8766726c31699bdf9a5d
za1ee3e4d138f0f1ef656a6c87f19e43d749127daf14a265ccb2d4fc6670b407ed8d3545b367d6a
z4c02f2b12e2663a83a403db6c40b8a57c814ea73d08ee1c8d615bb95b56b208e197817f7168c7e
zfa5dc225297138f2f11024cf031754ce0684f67d1eda5f11301361b1c9f35aeb957ed2dc9410f5
zb57d3ffa9a1db0f472947192c82d27dd6adff5ccf4979312f2afe4c432953ddb8ae1501e2f8de3
zbe8f82fc9e5beb28ebd8b46f0a56d83d5e40a3c73be603d79433a49dab4c8bf0172323d9b10074
zca4b9601ef8b7644426f4cf78cc9dfdbfb169caba96fcdd264e5f52f4a212cd4ea783a3b406ddc
za157272525a6ceb8045a00b530175e76b0ff4caf18bb435c2c7e8bb6801d129806577ecdccf858
za6d219850dfb803fcfac2196908a19a5af61abfdb33f3ca9d60639d90970bd6aef80a9fd3e9dcc
zc739bc723879133e36cd3bb2c238278737da4365e17158a1af39ad37929894e041f8dab478ce08
z15061ad3964bbf3bcd1c4f6b5146044bbdae8ec6867132a52358a91dfb5a25d1baf881b284a3e9
z1497bb26e267287de3ceba403419c992244a79eb5e1c5630655c197937ac3b5ff045efb2021b8c
zd0b3f47156a7107c7cef59e187cdf88777f763ba1b0bce1a9697808a8a83332c48a253200bf995
z526cdb659c4acae23f92805220399ec124d744f2cf231127193e62fc7e8a9d94a63693bce7aad6
zdb5f2b270cc4083bd17382167c581e29172109ed288b3a9c35186777c82d3ba05baef9e28c91bb
z6c379b11a980c3eef71f2feeb3ecc707bd8c7f6b4a21e73874ebeb5e5308ccb12dc9fe40ccdb1b
zd70b56acc6c1138aff6703a7bf861a9655f71db634be8129a6f0da223a0fbc53d16f1247901b4f
z884676b8c5e223b2dc5dfc6754f5c286569bc61415fc46409eab8895ef3ae7256a37d427351bad
z97db65bf3a690fff9c3c14c8c00f37e5703c173a13cf8776f638fda2879363f1545ec60807bed0
z77eda04a1997b093c0cff61f5ea8c4a89882b58fdb444ff710be58f82f01c5e373d9c6530e21cb
z63aac7d59b79a8792ce1dbb459d3f7b77d9371fafa7c7537d1a5aedea65ef03f97b8983d372ecc
zb36e830764ff1018c224816e193e273aa42338c4b2b2822559ab07c853102df9ae8b081c8425e7
z3ef1a083e58ea560c604bad8d36635bd90fe69d574574cc7608c80e126d067b879d7a2bb7a1e99
z6be907e2d8ebf90412a8c00cffeab0c7e4928487a2f05e4836d4656d513f96c9e033019a3c5f34
z154ea84419e20cfe4b7827a7a853e8560daedbddebd75cedd04906fefe97d3f34df65a682cfa83
z4b7867d8b408f589e09d3d67e51da89dcf69907ef3c2d3603a991086d611388c4e8002ee0f23d7
za18cd41e9004e97f5291a7b088d821917e6b5edc97c6a560c4d497f3e38fbd1ea3287004056c30
zb04725db5939c5afcaf01003b43c520ff3046c66fe9dce73bc6a322383bc0895a422189bbe8bfd
z859d69b325360c95262f1eab7611f6f1a019cc0967d04838d2e47dfb1eee1cbfb8a7e7e9eef6e6
z0adfe6976add66a2f502a8e39789971d9f05719cac2cd7d0605f42fc71b4fbe7bc57aa1143c771
zb59b02da59034eaeee7ffa3c6b6343dd6234f3dd3806275fa7a764e2b6f85b1e8b0c4b3821ea7f
z79084a9f16e24a117eaa5537b0d0b3e4e4b457085ae236218a0022b2c578741d56e4a41e8b0131
z65584e6d85416251b8d793467fee3c5af1b3004173fe2ce8200ccc0a5d82f3d18c692eabd3c594
zad5a83e1c3bd63e9ad8fc7babfb6304a3acb8080ff9d8b500a23a105ec71c9a9ac408814c42d00
zbb931de8765f707136d332715a451a25d0d4566f98ef24aa0e5d4a5b649c53bf43b00f778854ed
z794101e3e485c9524541c2ce17dba662fb2ef5f06e3c6c482e1734e7e57f335073ac93aee62f77
z69a2ab2e3c471728a77e9df20acda10dc24f87845b56c492f736a2e88c3bffcbd91b3ab81aa9a5
z75c042d45d483e76915bd1fd02cb3768d36a39e1f823ca1f56a69ed7af319ef72731ca2f42d44a
ze8efef197e6eb4fabe9c8b11616602d636e717f75ba217044d8b39b83ca58da58877c6f6851a77
zaa6622e27bde07105ea87e4e8a08c0fd52e602cf4f691fbfeacd65ff5ca972e5966c3cd6d28cdb
z274bd753ac65163dd5ae679d0bc8de37b77be897135c425d3f769942cb3382403f1125a0b308f9
zbace4e8f4218bf464f21e2c4e93ae8200172170b84e46deac0df696ef69961b4294c2c93a8418a
zcda12943e73de8fc029dd8bef18236504ed18d53311adbf00210d112e24622e617eef07ef3444f
z8f54856b3ddfaabe476295abc2829a9d6fa4bfccc12ca3cc24ad5869f19f279c941c10e36cc460
zb46a876594133750fea81c87c69e1bdf0bb491631a8d923e9c12c75f1dadda8807c1b8a53c8aad
z117c98d57f3892044b6f6dbf897ad1e13a2b90e97c72ea871922c5f4c701d56465aea66c4c518b
z7f553083b483c62aeb3adc462970978456cf659eee0d2100911714faf34f552645615c5ae6e8a4
z31aa4872ef390973e4747e372efe5f2eb6011f289652abafe00e88eb32e52db9c4f1596696be7b
zdc0355cc348f801c20652f3fe46e84f63d56033138c23db58294bbfc889a8403eb39a507fd1a38
z52b11310a19c8a9827cdadc1fc2b0543406f9597f50524eed5572894410dd5c67c878e7ce18b3d
z2f72d364451c88abbb90e707982caaee6762f25767ac97e5ce4f629b1288b446f4b6a474ace250
z3169f63eaac75dd6dfb5a3fdfba7eff82343bd45d8e761aeb2491bced7bfca50dab159eb257570
z5cd8fccc6d0e02c20e7e5b26209f7047f6880e8a02a1c8deab37b5a63e43d6daf7febb4ed7aa1c
z0c38d77b9b397826427dfa3214cab8560ff1c03f83247f0afc034561bfefde1d58c9b375e9f083
z44cbabd0603f049e0b9532dcd0e5e4636288d3a4d87991757fed4ff4329fd5096026281d91b55a
z78e634d251ac2589dae357481127b44a10dd2d7098468ebd832ed7e74c31e9db9db35a8fadbfe9
z23683053cbdb9a7e9ab97f6211253e1334e602e49ba61b3f184483e40d96b64cf62acb8a30a252
zb95edc1e0c74ce1bd1724520b4ef1c22f4c648f42bc63d1ad802fdaf65928be6eb8512f488a1c2
zfba34b3da7ea02e1fe073d72cc70fd902f4c9890a641c64fa3fde749495c5bb2bdf1321b742ab4
zb72c4be7741bff2bd96219a5a52aa2e4d64fd9125164066c03f46a137dc2df3a3bd51af613d501
z6fa219a1d93b7284a3d9a24f756fa9a172f70209145f6c7071e35df1d035ca634ff15a0f260def
ze2ccc46270432fad994a0fed1f51c95472fff72f062225b143445b85d34ca50ab06097c25ec2c7
zaa71ad73589defc7f17c0e82ca51e4b1ba1791baf8b2cdc604e51adfa911ad7e862457c2aa45e6
z3ccd14efc73e183951d0453cc01a42647b197ea8e3ea6c64101051bbf50bca9c9c8bcbab598809
z1b7699cd5a40ab0f32ddcdb6bc77fde3d3425b91b1c5453541586f597db5b42ca8182bb62899c0
z960efdd1e02b37a46c3bc5892131c94058b92a1bcd17efcd394e13d56f00b66890e0ee79165cb7
zb6a95b8a28d3736db8323270081247678e86553fdaac230b29a3f83eab8272091f9e9c3a4ce739
zed88b37f01baa378d4c2347adf0eb137c704c21af6a817478f731ce5a3f3ce1b921ae470ef6c95
z0c6cfcfee427988f026f8316f3699db54d17e13009e89428c47a33a7a5dd4b9b147b4e84d5dbbd
z4edb3474eac8c36b8719b873aacceb573ff71c4d8a5f92099ed66a39501120f8513bfa7c61dd27
z0bde96c041b72f6acd1936ddda51fbb184e077d775293de1c3206b2b58a5e62698d4b8eda2ee5a
zb584e388af0441d0c5d538b0dad10510631e82dd9cac5d861dadc6ac69a8551a9f118a84f15ab3
z2a65cfaa9626ee1e74727fb0695d09382efc04f2fe40769f47fe061f186b923773b95eec4cca28
z20cf9b2e35bac3e09a1d3f3866ae265a029df7c848b61bd8f44a30e791bb7b15bc8941d68f8044
z685efcd6316da9d50cb69b4994a36678393c3fac9d6608e88ab991fa07120e61ffd9c521678bef
z2769e61eb9633ea5eac9f2ef7c770d3a1929192ca997a99e748d784eaa921e1a1108a60c64ba55
z972f9350756571cdb68c636571421d6051e83ac277d8b9a9225b224b5525ead271a30ddb31a8c8
z0e65eedd5d14637908d84b046f35fec1c7f6036d8bd64ef3fd7b2f5f32c140b165028a0b5bc00f
zec3fcac12d49a4918cf23714084b476c8597c9be7054ed8506b8abe37d72780cf1083d92e326ef
z0c0cd60b21ad7ae876ebda0a0f202334e7bf5b4fa5bfcc30da440edc2098d14d9a53f7db66c46b
z3f78b6b343b19d58c106b3e6acae945d57f9747a54eef392f0d21af6fdb9dd7c8f611dcd0bf831
z10ab60e7424e29c3c4e1cf65b7c51200c630e30e5ef8e4b5d07f70086b6e73cfa42d9180eb0e5b
ze59246eaa9f6c050e13ef46cd5239f494ad780c1a834c2c7840696ca76ee284b87250a4c03b814
zec701aebb6a8a87d15ab5c03db4fbd2e2e989f58ff5d73fe7c3a45d8474457bc9cc521f7d1c812
z68d338a9d63b7b6338f3b8016b026365541c85e391c988413393f171233d7d3e842960bd5a9f5f
z9faba0747d30f9029c20726b781441de968995c2d08406da3d51b78d0d7a0a206afa5ded53cc86
z4bb006d68a499502dba53833e8872b116abe73fd64286cfc20a386656c82475f28f74a6ffd7150
z9195bdf5e67e429e395905a171a2ab8da064d2e7217b4d1e7ae013e482517aee0fca8e90ef7042
zf189d4ec2f106efff95f094ca98af914ee1c6c9a7ad897f8d9b6a12875a55b980b8e2529a01f95
z81361e5d04e76805288ba51b5559533873d5f3f62e7ff8c802e78c6c9db85a09bcba3346184859
z1aeac838b3987e575a0bfa993c3c73c4b58ee932bf319049606c65908b7093c2eb4887aa7b368e
z5ca4c1d8b3420081fc4196a6e4a4529f4fa1f6edbd02f3fe07ec549e70d35aa03dfc67e6a0353e
za5e22a3d2fec39587444d16fe7f0f9bfc2a2e3f1dd5f2cb2b7b95322cc695797746f5be7a3616d
z3b0c43dc3a1111f3b27bfd12d50e012b2d216b8a2466187f804665926a7a31a52465499f4f7396
zf0ee158a8c08ea8de37612793e3750bca999e8cd37f789d014a6518db3aa6cc990681af7daa341
za1357b9d2131f7b297c1638b509291f70fa254a740bf3a175c57aff3912e71023c193be959ed0b
z32194407d62e5755bba5cf6a658a4d36affe037289476c96618639a6991c7d94b3d8cc169c7725
zb99716badf520d99fbdb127b931a1c9032a67da774fba308e4f4f86aecb230e2052e92cb5c1073
z806816c9df8f4d67c79892ca4494e5449094c293eb870028f0089a389c46e69a30e7c40528d3cd
z4a384e9402e6eb38c188898176be72539c41e499de03eba2a75569edd06e1bd85a08812a62817c
z5880913f7101b4faa8d87d59b7f43bed2e92b0c1744ccf0ac05548b5a974b894f823c373f1bb40
z513d2664c89c255ca6210c9de7fc63011afbcf64e15058daebcc66f80d15d7e3e9061850d2e20d
z50b55d3d27a794c77d97fb5ce050c8edd762c1f51b261cb6d1c62fa8d72e24febb78d7d7dc5c7f
zf3e210f3b9f0f7801ecf33d192936ffd04cfa3a87927c87231d7cfa5e9949591bf3030ae9ff1ea
z61d961dcbe0755246c8bea7acc38cb12fca3bbcc4e5a477b739a7dad3f37266874adccbe577d9f
z398f7993ed4c71cb5ad3fda35191b8d3e2164bc0a4352ad8fb51831055fffadf006a89b0d43f3a
z6261d1eea338808c00fe1d55f60a36c338dfe2ef98613597561434824db9e53c8f0740e18e7d98
z3883050ac858b23a7c67d011412162d2cd00dcf19bfa9456998686883c2472056ee2aa1e4e4e50
za1f2e506410cfd665ad43026adcabb9132e20e6ef09e942df8ad9cc0dd8b22e8da198e21452d57
z23bd0f863fde1726484630da7a58dfe036be7cef3582012b99027dcf7feb3a754b4474e0cdb05c
zb7de40f5d477be40e99ffbc6c1655f13692786e7534a62569300debe71af09604aff041cd6aee6
z4b0bcaad4f59dc1b33b8b3aef3b7ff98facf9faa17feba670130125e364151aee8e8b091304ca0
zf16cd68196d9346f36ad671ab8bf870f20a1db9689d8428183f317c42e44430c3019d34eae6f9f
zb5f1ba93d47e995a1bd278f42cfc6c1139d402cd6889f1ace012d12d5c7c9a7dd0b7703dab675f
z99094eb8ee7524ac5203b1578b0e1b9f0b57f116f25e80a77c78d8ec71c8a3eb8b729a0b4fd54d
z923ca3c242caa7f5255e60b6c44d868f075a694f065fb5401eaf77c3012cdd00627f892f33894a
z74591d4b31b2b4ab53f3000185787378af2087dc00e86e5e1abaff7d4ec16d67459a3a6b9400c4
zbedd20d07e17bce1e4cb62a932c68aebd6e206f2305860f5cee12f81e18640fc4adcfc75c9b35c
zff50071421937ebdbaef4191715f4fa61fea4d209abb6c956a7eee3d438f12e3f3233428a18b70
za337c93b86d0dca07114fa9128d5858e188f71fa82be4ff906b4dee74ebc1f08e569ef52daf20e
z615e225e20a635cd8cc8ec16d8fc1e33c4e6b2a1e079766c8e904e55a953feb51c294ab2495f9e
z19cf91284157ffce68ceb72647b1197e8d4992869876c9ba3f13de1c3761ed7b8c3a718080e7d6
z571846422939d80d22fae28a65fad02edb1c34ca0d77fe67781d03370f248cdb16420a00ce6d6e
zed2377e355f8a9a19a5f5ad82f318158fd86a5b918112c0ba261a1693e536de872ef292428d997
z352402137bd765e4f4fa98b5cad1701c67841151534654d4f35412449c933faca69e97d1a58bae
z5bd20c77b8ffa9f784fac556eab3feb753dde8c5eb5f3bd9c6807ff07c03f0eabf4864439999e0
z15c3b80af7d8281c2f88c8e0d0bf4d4e546b2de70d7ac1e3fa2fc2cf2edbe9fe31789c4a42cd76
z75f9bb1a1beaf983055706a6a60f241a3fd027e14f445f672e83c2d7c5d9af7cd7ecbc86858799
z55a577f468777668b827065cb7055533cca633303cefa2b17d16057df23ed355f3a3d10a77f234
z0760c12a4c3a28ff8d452cd2d09d5017f105d2c9cce3285f845417a2a00960473ac94af6d52cac
z28a270e4e518d2136acf818c6d557dd889afdb5e78d9dd075c1fa897a692ea36c08ffefca3572a
zbd6b976e10300cf622a8721c23b53b5adab281f5055455ea97f06ea8ac66a3acd3a686895dd141
z7daff93557bfebf40367485f17bd374ee5309348554369eb7dff774682d397470e6107e24dbc78
zf069fc52ac00e74c26cfaf0b27ce3f5e3e755e84b4ca34a82d2ab14bb0a76554cd7131f9359023
z02224f8e051fde7025dac1abde94b2a96ca31bc60aa4df9818cc76448a8ea31a54069844726533
z098220633bb6c50824fd85a0f63adcc55d98ce485e86f0faa0d67f17a2f5310f6001ef358131b2
z99c06735ec7b0bb4297b83cdd20191d07d4a440b06cc31b3defa454eee1e56b52b8e348dc95392
z321cb8e33db4bba5328984f202d9f7cfdf05f8b2f8a6e11a40522f841027e874cb8ee60f720b8e
za72d156a4a04235ab617cafb2b1d915c904f64aca1bcad815d05bad7e9f60c5e66d1ef3278dcc1
z773f7814ca1a0ad48a32ad37c0b232c89de1727019ee842c1af61322cfa5f849aa1875ce504cf9
zf00cacc8a3faeeff55daa0bbe2427800e64a0a7a10f75324cbb95aa254ce651d937b966dad5163
z6506525682d9342fe1127b3347d6a5e021b8d6cc45c7c9876c3ed88b864ea0247486f500393f20
zc1a98be719bf3a01c4479d00869df1467b9a9d6e25e5f3cb3d3ec3cb8a9def80f9a497d5a4d64f
z4a139b8a061bfbd36d74f40279aef759b0264e08a47c0f9314dc2b862a28d9266fb221d00a3ec0
z971125d1cf855d847cc4bb2f52cd2e7d86a844c4b4e88413af9d904a3933dd0c9c629965889db8
ze400c65ebc6347106bb91c0255c4abb24391a6a78f2ab6ee7c49aaf9593859ad78215367b3a257
z8f560f338a7854f3227333b18de84e71ecc8a297144d3235b49df63188b89843ffa9964116bb7a
zc3d85ebd2f62ef1c9f031590fed50d2b317df93b12ead5dfcbe8e74e27dabab9d97b106e4a5f8c
zc571de4eb523818b292f1191c949cabc28c04bdf0f3114c4504f1618eb95fe339e531bd4f83fb3
z87398971573e4991084d01335c8521809bdfc1106f974256665b6dbc39e96d12e5232d021fdcc0
z7871b2c031464402bf43e05a031e70bffbfead0c0f04c23b459030ac8bf33fb6e7a2269aa779b8
zfb2a6b98ad83af7d61ed12bc8bbc5085287529347be73780f3c89870b11bb6df9d1c981c10e0cf
z57dbb5122de226946e932429f41a5627dcc02230b318f597f53b3836a7ffaa8d7b24e92a1d7a9c
zcfcd346928e7659fb8e0c00cea072b8497f371cba4d03226c1986293e8f4d102b085dd61d0cd7d
za504797593638fe90b869d87910acd7daebc9d0223ffd3c453f121797bdb9ae9d1758de87bb586
z05a98e2745470877e516c45b69bf88a62d01701d71132ca8a52a5ef7fa4a0ab1fda2b704418ccf
z85c8ba5116c6af45c8c3902eaf733f106997499bc74bf7b44d7db2a3d2694994eed45371707b99
za0fbe7d575b3b31a574e2ba8ab65494f4f5a01cb3586faa5b2a17acd8e049e8566213aeefcac64
zd33211942cc93f52290297052025e65d77e1c328402dd4c060dae7a9fa073218e46ee8b57e7fdd
za8b40ae86478dd8b240eb94d2eec82d47e03eafc0e9ef1ea066173c2825bfd563fa43901146063
z7df1aa2fdfc4c21db87de6630bb9e22ffdaf17fd4c5f3a58e4cc3b4b8229d357debc5948f90869
z631d69eb2d5cc9e98225e6e965191fb294634dcb159f7be155c7725d9f82ac196d74b0da96e46d
z52b10fc5da74eb3a1bbeba14e3e863af537aa7667ab996bade5c8775679ab748d39fb9ca77bba5
z46f238ad775ab68a0e97c74d70a0bb6d4d6c13e8d311d4500d103416f3ac8e1d59b1990f9ad7a2
z07795eadc2000bc2a412c9206f6c7638024280b1d45f11b97df3be26a372e55c74e9f8f7c5e607
z962c83cff34a9fbc3957bdbc31c0db4eadb2feaa817a6d1a3dc2cf68b5bf07d1ff6b1ee419a053
z5fe72e4b7a1df7838feccc44140ff78d952d54ebec2f9365f364bd442128c8d545bf5be9d09400
zaca2a464a69e2be270f4ca22e310ed9b9347ea20da9dd61a33b7d7569cf799cadc579dca0e1e66
zdfedcd051e7fac06ac15a2645016ef3b13c49c8ba95a43d06f814ae82e9212372582c9bc2e40d8
z1dc6490e61f06e4c04e88c43cfd97dc84a74afb178958667fa59d1426a5372c1f7cf1dde087fb3
z269fd4da7419ad1a2797e7157f8fdcfcf2e65a764bf29bf0568d1c7185c212eeabf59cbb0cc46c
z49e0b361006d759836bbc5b947d94ce882b488eb5f696c6eac742d3ac30ae382b1916df3ce4c59
z1b0bd8759a513f83dfdc03007cc634998e6d3f8e1447b1a6ffc12cc9773e455a9ffbd842737e7d
z03fd91c852c4a0ad338e556419199241d314ca6a224d973c2e0357dbde2b22ae1c0fa294f30314
zc7914aae8ede9ce39749befb695cf55d288f94bf2ee37000b7a071c018f646a2423199b4e0c726
zcf3b6181a7761604c4195678ad39e7ed3500f0fd0c0838c1f09c26f9ccfb9b50947f774d1e302b
z738f169471e3cfa975a90fa4a5c966d7780ac87ca049ec0f3c09fae1567e4b15e7edf256d3956d
z5978dfb5e1575d5d42aed0d8d6a2f434ce8ff683e288eb554d80841b3fae01bacbe56d45ef88b2
z7c14502bba37118f7d6f1f34dd881d4d2aa06d7eb1dccee9fa94ad8207831624725f357bcfb790
z566cdab95c4f0cffd54785476188efce47a7ee4c9859b7a31d91f947e4479cdcc1b97564863e1f
z3bfe2d29318bf80cbf26b634b3e8d7a6a9d37f7fd7ce5d8081b2f828e73bdd5914aa3c4854000e
z67699f20011a4528a7d6905f89e0d815745cee87d6b66d6cff1f2793f9f6dd5a9eb816545af93e
zef3a04b35dbd4a8c29211878efe944ebc62c73362671f8b924bc3a04cf0ae37074e8ee9409a0f1
zb32f59aed663ebe59aa9b0feb78804c927507a8f79a1282ee396570820b3a6fea4a0c3954a23bd
z45451624a7d7093b6f52920fc0421cbe07b4f9d2c7480e41a5ea9ebe242beea17b3dc3b7084645
z130300e823ceed0775a98d9acae08454f16498adf566a2d3f9c73230e6ab8f086e40dafd7a0c5f
zaa4da58b802732f2fdbdde45803403a3116c9cdea818e3fc0f7afa2a8337bbdfd001fbd02ef77b
z160347dac82d06e44aa263a05a68bc2a67787615cd8425c7b45ce7a505d2f149c1664de6d0211d
z4e0ec2cf1028c6aeaa6932a85cb8f00b9b5e6aedc66a6ed63aa146ed300203e269423d22f8ab67
z1a60aca082008981a5d56d1555d6f11893de060afd65b662aa6c58ee27ebfa752f64e76aa37e6e
z1c83fb057bdb70f92952e97f9f5c0aafb56b97003d2fa3d1cf34024c654e50064c03c7189fe930
zc9827055b61d3f914de2735ee4b0250a0c732d690e1704686b14c65f696ef8484c4a73fe6d0d42
z811764e64799e37f7aeb0532e47bb393fd7eda2dadd40eeb994a049087953e463f61ccec41bbf7
z7847f18da467c02974b0931c666186b1160a7072b0334b47755cfffd5e25dad501788b6f790414
zc7be9d47db9f9181da42fc092c406d0d6dd27544b545d3030b51ef2a7b9bdfd0d287ab1f4ef260
z9ced95adc70a05fff81d82f19714696ed44a4f1cf74c367ef5279fa44489ce031ab69c765adcb1
z905a3379b1a53c69aca15716d146580bb01605f9a9e99152e4f88ea6429de3ef6da733371d8e3e
z4f30dcc23dc94526d2951712e44a01cd041f7820d741c0a2a01990bbd3ae5f7346e5e851bd0ee4
zde4bd66a59167cdfd18a901098193a899acc3ffc31487d5f53e9c61b977b8dfd83cc25fb3217fa
zc495934592f11787cc64154f55341fc6280373d67c5ced459ea4b5b7086c9b0701a757ef3edcf8
zae26eb0852ee3ce1b723cb3ebf05e9c0f30ace43ce96cf5a1df6c3743c47798ee90cd25f9aed7f
z4279a8eeef6ece72db65f35b05ed9d57a73071472695f8ed8a37f9c53661fe415265ad4a9f1c01
z717689d5c363070e539c2b3409c90446bb5b4a2ea961a1c88a5b88811ea1ada34e26af78324c72
z8f156954c9f87247e1a78269f3c8106130ce7d829e939bcf08350f0502bddda7ce3fef694c8ca0
zff2f72e3f93a754c3a4b08e54afc9ad66b50703c4824fc697d3cf4b5dd503e725df24c2e68caca
z52c28a0b9235fc1fa6d05eb7425b6d6aa9595e5568b24f37f3cf8ebbc20873e2b9debf3add5606
za3b68c8c9c588738356ec56de1f58fa04327d67e446aa85118fa7bff5e0992def114aba9db3abe
zec7a9ac1b5605fd9a1f98a2d84810ae959763a3d4a78531f7ae120499f7535afad95163a54d818
z924fbb4a49d5df48be65706cf442333289fbfbddfde5b115fdf804190463461421ada3da1e28fd
z0fa9e8bfc2e305531c7ca01c107ed07950f99c6370c7c09b96607ae3c22bfb14525e1993a30487
ze210036a4a7499721a739f185f6bb0012dd189b484fe24ba59c82136b8fd235b2d453d80ee997e
zb32633c91cb5e91c208c9e85065df269325ece22ee55b4f6704d0d7099747436b0b8a63b47f27d
zb6101207b4461bce6c509ee4ea1850908d6981b831d130d8093cfda2a5ebb9794464371f5f088d
z904b96216c8dad7596bd508f417535642abacb01d42603a35213ae683d324cbfcd7080b5e39191
z8480ae9d90dff9d3fe3f400e7c080292c680391918feb99ef9c21f6082572f0d67768fc23c6845
z0c300216a3cae760c20e4df32ec67e2e81e3ec4260b7ed8168542a257d51835e409b2b0939e62e
zde91cfb7be098ae701ee1b184a944da0056578960b5beb9bcb55ace67f88d8e988b52a4e0510bc
z289c43cff66acd8d84e48c42a8c84137fd9ce7781d47199356d03a4751e5b3beb9581f5d63cf4a
zef2d64dbe8b9fc3a975ab8a480f22d8778fb6dd693a8dd86139aa50c165909eaf54b7c6516bfcc
za50b3ae2786bf7967a9853ae9dc68cc90b660101cb604936c8ae86ef770ff5b40862046a583cc2
z0157cc99ab814a7335575059f4f839802769a5899cf920e28685b600a5c56e725752ccc82e917d
ze3d73f2840077c47f08664d126e73882491a1cec13166df9404708f9d510af9a18007b12b31aa0
zab578beba0ec166d906207161e96abb6c6d30a4d56a30f3eca64beace1799a857f236489008902
zbfea238cb1a75c97f0e2d1b2453de55cdc1f69c81eb4b8cb50fd59db0ebfd60dac2ade8da01f46
za411ccc68465764d09fb87479bfbcab32956c8b9fa65ba9c6432d286c0c6e44b7b99ff975e875e
ze1b299a44edaa01d4a3f50aafe451bccc50cae4fabd8d711caf2a99e8ee0958aaa0f3ed6ca2bbf
zba215211dc598ca9332ee57116e542c6d67223f938968003469535f23290184673038691f7ffd1
z0e538b22301d3bd848ccc97b6e776abf295be0885fbf6755d91a44cca00262bf1a8d07fcff2605
zaefa27ea72249291b501306bd1742d4d53a889e366bd00a28c0ee46f8f08e707e311ca823c821b
z2c6a8921e3de83f1fa45fb7f91af86bd4d7d549651bf78318dc64665530a3963af45eac7b3e555
zddf714d54990b197a89c02308ee53361a2099f3f3f1d89c4814c7f2b7c76dc8703859374b5cbb1
zab744576d48e9f4254557a94ffe7a065f4152456f86483a68a1e56d4f59698fa372595976de38b
z0ea6f9189889d6ff27b5abccd340a2716ae4f6ce0fef836f48b5f7339be817402ea02d7bdd4582
zaa784e9cf4764acde57408cf15b5bdb77d4ccf857d71563394bb0436ed6a0f29598dd0b5f4c40f
z269f0e64a21054aed827a82153bb7c0d29b8c687055195ec15a64d2756908d20a386a77dffbba8
zf8fdee62e2fd8544e0ad3df9dc8e1748ec745d0004a73a7847615d735e48f516e357a848f5a94d
z0cbfd3538302db405b97c15bb2c6f2608f174fbab1fdf92ce17906c8550d5b3652a6dc8fe953ae
z718f17d45ce5b89b64f2b2a31c80e6e992e27b5ec5e8d7b8ff41f033b139e96d84722b4e474818
z3848783b6a87fa58361b395523a0b9c365e62a447d00ddd8e31d7b01ba6ad838ddaa95dba23d8c
zcd223f11128878dda2dc1a5c2d43a93519e73cf13fca918daf0315c980c856594232eb1dff3fb1
zd896e8bcd84ad1ca200a38b9d3c8e60aae63ac0616278e6a7539a5b15f47fdd2b6b1b3cb7a6b1a
z802ad0bb2be462e7e36585e6d97986fdfb2ac9a901e591762f85fd4943f07020320529d380cd74
zbc955580bd3b1d44e7501484573f7e0e20a990b1b086e6a151e7d9db45b53188d85110f2e08232
z1264808e16a782ba645cc467c086ba1af08aecd8d843bcb9c0a68fffd0db8ef05b130a2486d92b
z9974a60538868e153ed7e4a5854bf0f8c7a4b6749138a145bcca341f8984fc495dd4ad90904e0f
z8276a2db872538dfc3a48d08727d0e7748042475ea5e4078745e810671f1ff4c4b2f119e9c0d3c
zb273433e52ecd6b7a505beab2f4b4c57d16f00744b0c678d3684cf49255adeee872d0702015d56
zb1be505c99f59a320bd911da46c8737543cebd45fd530000145eff7a76fbd5fc06f24118dbad02
z22b0691f09dde6b1ca71ad9bf2ea8cb5bb02b18978af18be946804886831e9a1de9052b3592e87
z7ca8a73523ec5cef384703f112d8ed871934633cc6fa614f53899f7aad6f82d01f4b46e6051cd1
ze1b9edc04dfe63c80f3064827a8e70e1e9c7882fce8c7fba586d03b5726ff2669d20a0417415c4
zbf92b4993b5a200dab8bcaea4fa808ca463cee0eaf4d285967ecbecf7e541540efb42dbd3fb712
z90dbf49bb78154e4bf50246aebe5095606e2d1e58742e178a920683cb4337f658cb19aa4f0a353
zdc68c7cfbf62537a4a37a11978a3471cd5c3726b9a99100ad4d9848c94f92aa9ca9575a88d338e
z688046ef88950e2c96ffa3e3f81a3e5d402e1ca45e31d10759dd7ecac10ffcbee53c9685494698
z2cebfd516e4dd4c21f84f23c93719e58c33bbf592c87ba884c6c0f107a7c6bec0126cd7a751ad6
zbd90d00e9ad094f3fa51307ca27d45f169861e3a95dd281312b40ca7d2d960caf3075573f61d19
z9435421c56a549f0ffab2877a9b9732d458da5de1c7e3ed20ee279913f6651853e7fcacd6d731e
z6511446df6e55fce47ea039613a5ddd39ede80cf3d420e21ca76a77d5b2dc9f6a767709c7c6524
z67716ac46a345eb6938d293a360e18014d888fb149076db94f6c3027dfbe9e32be14312eb70dde
z7e5ae648ed4a76777287cb991ad7363e99bb7cdba125e6a1191c1f621477e191df7322cf5adf18
z31e36728e9b3346ff3c1909e2e7a97c4544fa9de8d2812e3f89f31f2f827d1e55f885f2357c562
zcb3a28ed493d2131b11baccd4dde89bfb87d056338e378f04926602c3006d6ec63252b8d2af2a6
z78946a53f2701a1ba3a0d01ce8f20c16aa2bca103a829cffd1463087b0a2dd3802eafe06f53dec
zb9a0dc4f92eae3bd30918195359c4026a534264c7fb2079b1c3dd5a7c98b4080d67592d89103d2
zed5df96765c06b5c47f5ae03063305e23e49606be46d1e550fa34ac01fb62bb1f7d24513137efc
z3f982f547a9b9a5ae5e9bc164418b731a82195cb0c1b64b564535342291ff5b43a1f6cb6f248c2
zebd1a65f0c780843aadd6f6392b0b0b330ea4d1e66bd0b0dd093902cf462221caac013fb3f1c57
z07543398fd48892b1dbd674df95096f7c84800cf21f86ef1cadc0e280b0170e5dc346ee6a5b928
z232d9fb5e9d5566498a2489f491e291e77a7913fcb6aef401ef95a031cb09cb52c8d5919973f1c
z347614b466f42c29b25506e2ec1075d2a56dc4b5eda1642c477529ac8a86d7dcc7f33cdc3e411c
z9fd9ce02322d69a248330b0a48578bfe3564fe56d8c29280e14556df2640e0b454293b7f726353
z287d410409c9097b0cdde1e40f02b66a45085bbdd6b1d7949e5d455ab90af176a2c37068ee3701
z41838878fad1467aa5ba62524fb4ded12d7d108aa5799d3ad01054b0dc276f857c03c97bbd3e9a
z7fbce49e5588e21fe2e26af9be0f440e81d9f2250583ff516362c0ba42046a65451d33849fc8b9
z1abfb390e26d670a520acc831d1f60fed68bf2ed7ab884d942dd5b0f76ff171e518acb06c6c754
z3e3a5f31fba7ca3e2f262dd501310f0284a0fd95ceff9f024a3ac023565cf804817e25940eb67f
z68e36333ea24a3bc9ba6f321c9eae68f41370a2cc33d575e1ac9ee4cedfd4d502328d00e37cbcb
zef2c89010468ef75aa1460f2c0d67d6be8c0ad3959c7725e4c2e27281a5b39dbac3cbffca8bddf
zb328293e0991af0d563f82a2c308d1b2d2f9e11edd16e90966866714d90f493b852ea577cdc181
z934014c6e2222a59323f266230c7927b8a8f615c199e24037b9262d729d6da56d8ffbebd51e2a3
z1325d1a30be17a8110658e1ceaeb924d61db554dc75c976af812d00f519c3f847f44e56aaa254f
zaf67a57348e0cd77030c77ad5c948c29b3f2a2835594657c8c71448ff7a7e20a0f21856a2aad45
zf021986a49494c373e1aefb19b47b38fc22ed9608baecc5260baa3b54396d55571efa8a1887fd8
za210eee39c60b345d75280ebe4cab4cad8bd9a9c8686c9df9e81e412457da8fa16eb2242dc3ca4
za628d19853baefccd70413e9954f218c3723b7ddbe7ff8c7add9c2900759303e21432c5a32f848
z1c2b1ddc1e6e1ac54ac843211083bbed57db99412ca8463d1b37e57b1353931c4e902e2db7c8cb
zc0c9403d459b1b1b2d26c1c4f273db22e054f410fb0093b79569fc44192d412ce584e7d617e129
z69de071adf524d98bf8c75933a8891a699c8c55c09d152260b8d9e01da984849137bc7e2414fa9
z9adee068c5b0de2104c89e55e3be31288533ff45936385531aafa307b20d5e36bbd5d7c0f4bfb7
z38b3dfc2948afa99f8ee85a9fc7e01318c610d9fb0f4096c192aef6a221329a59be001ab150f74
zffb1309234638b714df13e601de664cd0e689d6e214f6ed3cc23183fccb84815f4082364b14b13
z93c20aec055e8118d8426e5d9a4ead34ee2fb2b56b84252f06352e28331c8ace76e626c367b0c6
zed38a36e566f1daeec5e8e85f72a1c41df031186cfff1b6c214ac335af4db62c03c34a9eb8570d
z6e27c50db87703aad1242aca4af993258df1dcf63dcc1681ffcc37cd87e4e4cb933dc395b087d4
z0f537b8aa29fc06dfe9037108ca6dcef548d39f041038381514a3acf4d58b07d9ad116ca0b0121
z10d64c72009123a95ce9cdf9b809bf035a7c035246002551ab85b109f43447f547aa94b0ce1c6f
z814f78abe77b9b20d674bdae3a5e5498a9ebf4cb306b30a4e9a58dd193368268edc0a1eacc391c
z85ff4d13d837b24f6382fdd18d5f5490f1c0c34dfa565bb577916232678e456014205f8faed0cd
zb0d3a413b7776375545cf5e4af4b54d173eeefc83fc9920278d1f8a2b04ad201dd98ec27f7a06f
z4e72f6eb194ea1f0c83ab4f2da678d455d0cee060dc12cc7d2b86b43bdadfcc15192b7f43c370c
zcb272723ecb04cb86fa9edfe927a10ec7fd8a6397c863fb6e913da1f42b625b98efd293c42e728
zce2eee9c381158573153c17fc277519c3eb3588258b35615daca000817c93a057cf904bb148e6d
z2645021f275e1a70f7a6b16fc3d8eba0f37a8330af935ac1bca9271cfa2045497730e45aeb6fbb
z20048423d2a4ed1b6ad19e16502c6d9ba1aa24d3b3e642b5db18c41e914e91e76cddf4e45d4071
z31cdff9c0db059d15774e4734e2cb6a9627f9829ad99aa678c36a3caf68688c2d367154d276801
z8fc0ab6875e5121a6e0f9dbc2eea3b1ad493ff90b766183cee4d1470a751a368bfff911f88665a
zfe0d2edc869aafce7fb224fb8140a8e6aa1ebcbe3f6b7672d71bfb3cbb3c60969aee78f01039f3
z9f951e764f795e2b78835c99fedbf6aec5d284efdc367d8f8a939423cbedd7454e96e5653e215c
z7c010fac4f4c4f103e0a676947943d38b93b9965779c2df06587a39ae825be06326856c34918a6
z62e165d0d1b638c43d47f1141203e5259d7f16a60d8008932a7f56ea5e16186e5dc266221b31ab
z323f81fb06f0707b31dcff47e926e00912c26047b8a8dde96c3eb7c05d5506e35faa267fb0c851
z23493f1357cb0520fe8b4d9d5b37294e84ad2425c2394250c67470571c3f88b93816324a45fe01
zf39a40e7a7612854e4631dfdc67b9548faf3eb60c903a7e9930f827e6c73bc2ebe261b57df0fb2
ze26242239a06a4f9515d356441d6f9ad8aba959aa95c23a9f2fcae7cc5ec245e8ebe35351e5c14
zdbeb58b8a731005b225e29f88a334f2b49fee6dfd7b3be1aa97a77521bc79d15fd988daaa39c64
z0695f5975d5688e0679b9a08be6fabb312ebe5352f2a5b30f969ce1082c73b51441ae67d4809cd
zb793b31e8ba7a01539c24a42aa9ea675063b3bef30c69d5d82ee6232f0b1bc647b2bcfa979ec87
z2bd0abb596af24139c98ea80473e5aece061d113dac7eb027133c94ad9a9238c09780e7c23bb73
z4573c42ab0e2b4f7837b32152bfff42355361e8b340cedbc146a1c44a2a86d9a88616ea2ba7a96
zeb7dc164f945146e83dbd91d6d5c2a6e0b5aea6d666acff47e9b6caf2f4ce574cb046aedb37aca
z7e0dd019adfd85a84137470fd2c4a8ba86967f6dbcd06a9f8838f104e76b43b35c85042ad619cc
z596e8f7e8e970a6e17ac372c3467975d440d1a44c854eb14526a3df8ca57205b17352370a01416
zfead6f16a6a1090321b6e8696cc2f0352df1350e28fe63000f24079c171f35c6064787a505bcb9
zc6629b26883f4e4f39296d6d6efd9515971884e0b734d273ed3eb421bffb82e8f976ac4698db6a
z37e0bd9d60a375d76ba441364e781349b478791501151e5724eff0d48f7f361fd18640970b5ba6
z26d1c1e1220a841d39cde6413beaba6cf575b0e4e08227a4ea139404b9630001018de3ad3d354d
z0299209e863a8eb03c6634814da057797717b47e50ad8587ee980e91661aa786353351c182f460
zda860290ee6313af3c9a2bb3f7fda854a920b4e014f05aabf367e2dd2e70b9ebab65a34589f1bc
z43d9da0b92eabe6bdd0555b5a0280705b1017e7a4f2adfd5dddc6d981b67a6d137d6d2f114d20f
zd3ff734c4c4a568d3fd60aeb202999fcb33d4e0b8ddba0f2a925c07feefa96f1116fac5bdeead4
zc3c3e0d6bf53c2a27c907ed42a34352b9e54147211bcd0034e38fc3477e83a92deae6fd0a46e67
z6432fb94ab0463a7c6a24511874492e872983419b20b7b8cd5ee31fa50b791b70f846c103258ed
z195a4811193b2b68a4a6e11f89e064aa46e1dd0862f15a1e02bf505835fb7cd5b8bc19aab8adb0
z4b5e0975e6bd70f8a4f97c337d5a73719a3688a6371035245edc9609b97d2ca34dd04f2b022b10
z4536dc34e11ab046d086f8513432fcc74c1b24a2a08ada1a86be224d456bdf3034e583cda3e28c
z10f3b76331ae3b8fe43add3115ca4f8ea1ecc7f585fb0ea150fbe13b270248156fa61995444d92
z6bb72c95097e42317cb5eeda92973a6eb9e0ef5161efa30f88ffb1630957bca86458901227767d
z2e615ec9247102b385a0026fd8b47a29d834cff8c2456fae756b505004c2ac082dbc73c64739ba
zb577c7b88bfb53eab1582a8338e3a77f5f6089f62445d60d18a3f960a95a219b2ad41f2698bd69
z817182dd6fa20fa886b8db3406ad4aa9c379fe883445b6173e796ee1fc43e3f3d8f0ca76465285
z438f185f99a92499dbaee41ff1e2b0bfed69f8a34d79ceb79366104e78fd414ddf827be2017d62
za7c62b9c92060287a8f2bc1980beb51578a0e57e844748f8bcc2b7fa90c964dd5fc47bd7b1316e
z7e565969f9b8cb6d0c2b4d0ac844b2190ee61fd6ee56fb03aced3d029218c3c1b8f3c4fe0d36ad
zeb24671d7ab73655ed5abeafacd9c6fe97cb697c9ef9c5b5046da85e5360ceda682430c322d22f
z81be10a2b95e46e06142fce6ec9db849db88b95f53fff3b6b408ed3143e250d76ad0b388af9c84
zfcb7e56e79d09e147f1d619fd0adc53d4fac058fbf32ddeff965a8037ef89538846605028fd10f
z85dbc160641911c4be287b73f2d6b51523c5b5accd04ce0833b74bdadbe3af8013a2908ef32ebe
zda09543afcfaea460b8b8e975357fa3181c6041e51e82c5e720221765fc535bd0b23fd770dc7c6
z18a9975e69988c02fefd9943672c8ec85f5085f3b794c0bd5a36716d8e94d758fd305253c48933
z552a96cdaa7a7c8fd0715ece7b20e88a8d781a7476d29af504b6c4077f56a9902721cca0ae0578
z4323c0151d2a4d96b9ef3fc119226d83ebb864e25dd4b2cf2cf29e9ebb438725226504947ca4ac
z9653d4ad9b464114792be079ea632bc355030b0ffc4e62f17f928724a1551c566397a7d114f4d6
z7acc2d6a1e1e454f84bed5b48388d0d7a740059dae2312b1d84c69137f73ecc7c68c6dae127b66
z4b98f689008d280e0f037b8f513f6e27c9385913d166a9baf18b66080b1459b529031f0e431e51
z960d3744d40faf79862a5e846801f6e7cdb3865ec4b67e375143f4a8ded79446105a78ce2af9f5
zc5dc50d5f410eb1cf808fb050514be35c7ac86cbb4720befd80ccf69773c314592104805555dbe
z21fadf0a4ab3ecba2b261f903160589ef6b933dcf0f099bb2fae2fe4d852e32b5d5b30eeb754b2
z500c958e1cbe65e1ad84d1b4b97896ec6486abaeb47d560fd2f63def6694ecb69b3e0a5195b32a
z502d3d6888b6d21433482c99f8013221b4e954cca313b780f00898d5e535fa396309b6d84a149c
z577455d67a0d9d1a573172ec2460ef10f966ac20ff9d14a0030b141e39335159c841e3e753b45d
z2feb804b2b6d155432aa2bb4b658cafb359be12c9bb9426585bbd573366754cd6ba577ca9e6dff
z9b4fc9fceddf88af0652a39d8187f7f94ecb0790857b5382ba764dfabb1eab375aa3269d53cf51
z39d077e632729e73cdc1d648ae2032be00b69947f6e4739fa30804f8865152b448f9aa1625ca65
zc8c40e0afe091eb4f14097d71432d3e9994af6c15b241c939abd59d31e2f23eaa10fd7a1eba6d6
zc84870550b8ed0bf6965f44c4fa01f7da37e4db9e17d8dfe5006e4861d6e5baba4d7701167684a
zf51907bc50608076dd1bf9adc311b802534e502e6ee9c2b0f98b10c895df8f52d2bd98f866601d
zb2304903411035b17fe7731e0fe3168892a191d7004af8c61cc5ecaf3972e0d72890b614a072dd
zbb2f07132fffaa442703e7c0641987040d118af69d8594640b5913c32618e284652a52d19ddf8b
z0ae24db6e80742f3630843d951f316628b90212caed266860b1c3373f0fd30995b1c14b7744ca4
z92a2d75fbbf78533a889c8ce154b44c5399e480226bc4d859e85ec00137bc0e98b4b509888fd18
zbd5d7d7c6f857589466904c2d80a37932c04a786f674132c70628218292109619258da78d7069d
zd7a289f99d42c5bade0a27f57d18a579a52b3fbe01996d9c72adb0d43c5fe85fb2138baf062bfe
z96598545847192f3f97c2898804e7642462a2b7a6f8dcbdbb722cb6f63343fd3176a8fcddfbdae
z74823b35b8e03fe6986614f06ffb3d43a794e0d9f8c7b41fa110952fe2a50d915e1ab0c2b004e3
zcea83de168a10fa16f85465bba9dc4cfb54495132560f665142e6eaf89a621e3ba304d86fd1652
zbe546271a243bf6e06eec01821a37ca9ecf400bc1fa8712766b82fce3bca65bf728f456869ac43
z1594a7289aae6a5b4eaa384d38a6cd3a2ed8b94b4e034586cda0167a675183a8c585ece25c0c6a
z02bc8ca29650386272eefded7b8b7b2018ed6c1b9b8727524a51c65ed754e644a17dc49f213ad6
zbcd870f5295e056c4c1715688c50a0ed9bbcadc694ada231a4e0dcf49ec7cbc942f72d77564379
zc4788b8af25ade6d4fdc2a3b90832aa7872295d3b6d23ff91a4d303951bd22f3d1a63883d70001
z7aeaba829249898c276fedc70017b9105fe24ba6a6cf0764c5a5a4e642aaee26565a8c9f18b8fe
zdc2cd0e24c2553e0548126ee0c6822a2eeecbc99152d1a86b207cfe5e09630719abd44911ec529
z1bb1387ac0eb619e5b5e238eb0962a40d5d3c3deabb0d381d8f5e2133d9bb183fa9c75e12043e0
zb18a3b0aee928243fa96ad8ea8dbb8f0e5aa9adfcaa3581f8d95edcebfb07e7f08b3be92e0fb35
za8ea2136d0bc5718ce07c31c6f6d5c2a64feade4de26bbc4ac17ce47a7502dbabbee64b7782f1b
z2f4e9b466df31916b9d5c48ecfd63ea7e885c6fff87cb881e59d856269bbea0eb774df5c23fe1e
z02ec27e88b8330bd4a85c0a31906ae05fdc19dacc740c014828a56c1ac752e896e3661e554f98c
z8b97d07e7b3bc670f904be918c669153005038889e8cc442effb676b13c974314645d8855d8f78
zb8b545f2415a021adff6a7a623f343d4571034cc2cf7ff799b54f0795ddae79a61d8a8a5bb4092
z6ba89c67ab152a1088737c694bdbd230c9ea128ab05c5d1a3b5bb4906f2ed7906ad642e62a5e88
zd2224e2d41d303ebc07e149b775abd66f03f770d5bca86bc6216853a8476d4671ac3144b0201bd
z4c0966fd141816890f9fa26571d67d8b81829bf5f0efb354d1845bc850e6c91b2acdd2ac835a37
zd67a5077fc3d5a21222f7ec41074bbc7a45c2b7c4bd1b09f3e835a9a486fae81dc4fee14d83b86
zd922ec317dfba8b96e1fe0819a9f689aa86072fc7c1361f471661b8351a5d2ab467ceffaace5aa
zd830dbefa1bd1190d8a35ecbc64f67ef3aa0a18956a53e2c3c2bfdc92d105110fd800bc721d869
zdc4482be0a6bff1774ca9faf4a3d222f0ae26f905afdcd9b8b350697a0573a6bc13fe09d04f3be
zd58e631532246bea82093ea86abde1f715154617b1a615724db6cf63d3fdbe159c494c76133957
z35ffffc153fac6a78f156d5242d0a2391ff25f0901b4b652d5961226c0d215c628e84260ec7eb8
z28bf6b5bdf4ca3bd7904155820f9999887e6f4935b97c5ac016f7ac3dd2cf0cda5eccfa0bddb
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_sata_stats.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
