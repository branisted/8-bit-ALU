`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1b396e1048595951af798d8de75c23e123dcba
z74156e068eb331e95842c597f3ccd341bf87af84cccb15a44d811686c10b5caab6338f8bd390f9
z35e3850857fe16a4bd09a1f73b16fb4d985cb91a2a6e022108c6d66aed9c9b28b7bfcecdeb30c4
z21adcfcfd1d3a705ecb82a7cb228b602c508facae7d7277529f388f1ae749d3922daf9cba774a9
z7a2cdbe51bafb7233b5a04f9bb9c3d371ea04be74069b3a4dd10e4f6c35c82f6cb174014a35e2d
z402e001c822d16b1aa1074708a615899420d065a95dc28756fd5bbe26801945392ceec1550bc0e
z515f0fdcc539c420f798c16eb9b9a870afd7c2d087012d56c6f5d61f91202b9ec8e4e23c2f42e0
zcca954964eccf2c9a8fcbdb189ecbc1414ef7760444dd7b8da02d1eb9890fec73370650b4ebf34
z957ede5930c6977e92eedb14f0b7a339dc32f20f994d01dd3c5317c1c2082975bfc237a581d64d
zc8074e2c08f317cbe7f1667e3171ab757132d8b950b61bc2d35a431f66572bbd8eb14674623c29
zcb53df71e13cb1e1644ba85189af6e0b860a88e897e0a058efd779c076f821aa87c8804a441b2c
zc9a100d69e12be91b37bc1beca2ec7348e6cbd8c1e4bc31620d31f377592be45577bacebfdd441
z4e20fdf353524730f177690bccde50943390b2a7789fdf9526400d7411e69ea6a085eb65e4ad2f
z0d7d638e936b6a102c456673765021abd616e05824f91968d5d698d7be75a3dd7a676936ec1258
zfe9c853362a5a5f82171645717933cd9c90978214aafd2ff4f1b842a635b702e48288c4798821d
zc1c5d7916e30904630e78b0bd97519ad7b612d2fd860632a173486fa0fe020dbf44776b462792e
z08331229e3d0206a89fa000179d9c1fb2f774fc5abf6c2dc1cd64204cdec7e446ffb2cbaf7c792
za578ae38b3c87850423cab5073d30f7f472f21aef3ea3c627dbce0a15e4bf7b5cfcb2aa5806953
z3f4f5ab25c63b8ebe1e8b13a27d0cb8e79a313d9662c532699322645e7f0a37bbf6ac4c55654b0
zcfa851fb81e28bb150006698ff64a946a8528c881f626049e58795f6db749d367fe361d7490dc9
z31566f440041fe86947e3cd23a1b17d2a127a2993bbe75b248066ded6bc32f3b350ac30ab35829
z2dc2502bb4ae34afbdf245319ff5b70c7537754a7c22f70a225134b9f93900c1bb4f57a920aaa4
z4aa637c64687afa9cb07f5a28658e4bb0e6a0cf3cbd6020a024cbd3b916433d8f95abe535bbef9
z3b95855fa3d52b2b79235ba10ccc72472841303cf14dcc01e1a130f32891b39214453767e30a28
zd33e5e33accd99b2f94ea2971851db78ddbed303f7fc9f091578d8d9fcd4a475806abca16a015d
z2e41978e141d24f3122bb553390dd56733307543a9fceddc7688076033960dca6a734a49ae7ba5
z7f21b9b7a0c0bc55beebc6a07c7003fcb142a3d163aca0453cc0d6383b6af3123be3ce775b735e
z1df1f522b14a73d8922db7dd24f05b1c8c2a777add88223f118174495dcc4f32361dae8a6e02fc
z1b061ab77f1c53d0012e991d54a6f577ac4454dda052346568807f192330ebd235326f089d6b1d
z69dc7ab7fef2d4359832ac5824735e38196d30f5f37af34a2d1c7ca493b87b2bca5c4b814145bd
z4166d506e99901bfbe96445986daa62013feb7b20c2f63e2ba72c8bc9696687d98febd781f0b34
zfb7172ee4227cdfe414bd493ab84d4d9e29f66db3379d70db9d3673d3832c39b84876e53eddfdb
z72150a9454897b6e2202b62831722a3a482d4e300c234ccb7e03e2ecaacf36f7a8733e658b99bf
z66e286f8eb64f89772f84d1b4c339817d91e2cad9b5b78002277e5cdbc2990ed8add19a59ab809
zf0c3c3b0847d4949e23a2ca97a5e6d77319663cd0b7baf2b6c62716790f6108b30f1bb48ca3d75
za90ad563967088d2872fbc4d50bcac4f029c867ef5647f7bb1c6aafe2b6af6a63451d72155ce94
z351d56cf719a8509fc6eac12f5d467f8abf500710b223cb7edc7b48c872a989dd56342e25eb577
z25da318a82f9d8876f5c58f497d6dbc6a90554984bf27bb386d06a1ee0665cdd9c4006259efa72
z2efba71d638dae79fabc5960ce6f54be5291bf878eab1f87320f0e3cd1e7ac12e78d644f2433d4
z9f71d2c33a45d937d47df8f9fac0bba0a57b855230507c71cadd1cb09c5332686f6a3ba7ae7c6c
z5f327c146b96113e834ae58435d0f99ec5c6682f6827bb44b05290e8a793435779badbb11ba9c9
zff8f69be9393fcd94eeca44c14b35a143022a133d5100c97a52412e3bcd1e40c18816e09c3282b
z2f3032b7a4201dd08c63e6e396b839c59cc74a7b84eadb7d54d06c48b7fc7f2663250a53c4b6f8
z371d3435ad1e353d33de72ce0b4e631842482264a471f29e51f43273c54d545e24c0c7cc384068
z9a5714795e1aa4890a3d2c0a98595988ec06365c61b397b8cfbd38808804e4514f57f192bbd4f1
zeba7c9d1348177580f4c586d20e6fc2c5d8422a5c3308313d45c292ae00fdc20f73d0addb039b9
ze3de59e2563122abc365b9f774b80e6eda5430f0af0e6659f7b0e76d687272891fc0772a5e55f4
z1dc6f8412469c77cbe5bae2435faad0e99b1c6a14e416a83ba5a741c691e643fe805450f355617
z575840b322978334d6d73eea1cff132afeefb75c85c6a933093657a7d1af8e9232d473a07a7183
zc396173debd030fcb477b547c5e32085f9e4e8addb15b6fa7ea69f3158764b55f893344c674980
z042bb8f7474c7a6d65fc02de251462859263cb923170f99783f977617733580e29a882dfd66a2b
z3d4a32eaffb9607d0a4b345522e120916590a4fa009356f1dc3776f7ac354b165c8caf71af0634
ze5f33509aafb0ae44cca68b6b47d10485082957ca38d6a74cb2599a8bd905674345279775ba7d8
z2dec1293ce427090f5834e692d2974fa8422f7e0e02b92fb1dfba0c8153ee49cab9a05a5ee6613
z09a568168fe3b4f0a406cafbc1dfb2bb51d19beaa3cdd917fc7be5d7270a13a9025eee7bbb260e
zc059db3fcc4a5654913222a06fd09b936be571eb5df192d93452e5688db91b3a6a222746a86ca9
z9410179134838b16ebcb60314eee08dfbea91ebe40ab688e57e42113db713bc112595d802b5f89
z99ba44cf2741e8b15abd03ae287863683b5a7cdb8557726ddf20128cd3e0bdce75870e26912bb5
z3c3672ae3e2cbbd494d8360b6379d5fe0b1e71639a188ab92dff1e4463b44652b762f7b86051ba
zedea546cab2fa8685b764fad87008e6a716959acc266b552c386e20c7ef0a4b8b9c4a7f0892f92
zb35a539d4e037c622a5dacf79d55f925404bfa93f0076f52ec0ac2354ed0a7db1cce7724b37fc0
za5e06ed7ad300fc1e25d1b60b6d0dfb0b600319b464bee72c491b7f05fe60eb19d7911ffd9240a
z86ed0c95ce12421f3d220e35ba455158d2c89c5c615f0eb1d193b3c8a27341628409a1cfad1437
z1336adc0c47af3877f600fd74907c73deb4eed58689dca9373483eb46d8f6e9c2a30e524ae201a
z79da584b2aba4c27891352686ae399b0a33d8664c1a6dc4c628c49aebb59c0bee7ff48a41f0f71
zbb85db2256da12a2a39343a01dc89ee50acdbb7157d4c7d5444eadedf8af0217cf4502a2b4102b
z93c2c6f83a40d57ed2b28edd3a4e0f3952280071ffa6ec238acbeea05d48def102a1d48c8b30c7
z5eb04385a9a83dd70ab69df6f79b6616f9c2e4a900fe7eb05fa29e3efdb69648cf1d01f682c79f
z40e6087884efe20eb2a1162edc00e84cf0334f75917b9174330c8c44a796b09d2d12723e6ce0a7
zfcf35e3d18abc95711495a362a2f4168301673c0075794075676eb70349fd06fe2c53770fdc299
z61dc1430475a5c37c2c2cfb30f3301aaa5423eab0b9d3112052b88128afafba74ef7d20a80576f
zf2393b23b5f515d7330c6d59304cf8ad1169315a2903debbddb77402f317c40c02f063ab5d4d2d
zc7f8664aae0f0bc06e61c0641302bfee838734676e1c1a2a90c483a7a4c029d7d8e314435c425f
z0d6b9ba934bb31d385eac7b075007c34c2e443837faae1b73ed3d78b94b2e7ba3a0c2b746eeb38
zff9455b0d841f5b1e2354ec01d17dda6e21d44827ddf44d2aeb56abffdbdea0cb9f308e337b7b6
z4a596187d430fc6a9201671a45f90bb3def1c14d7a9ab3bc36f2072693dbef09171260b33c1776
z95731f221f12df14f8309c796b4cb7ccecaa26b6b60d3b8bce09ecaaab06adac75c80baeb2772a
zb2be6d0edb1d7e37111515d9e5567397fb63edc709b40de768fbc8eb40d648d7918a06b1ca7efd
z1f2d5ca53e302564fc3dd36d08f71b6f4b5c43fa71589044326c0c278b766f4ecc89cdce2c1082
z6bc2ffbbd28e2d1aa55231f6232e724e761fedc636359c0f9bd0f5b3f1d08e4150c18cad20944f
z61037521e2de5cc5ac664c2927aea4e1cc9e5f1e35f4a7f1bbdae5a2539419587fd8b58cea40aa
z08393ddf1f56a262d0a7c2ee461fb0a0d19fc9de906b4630424cd571707a2add254b611467b62e
za0c6d38dd1efb637b642a0d2ee0997f8579f9e141ad0855071312f668d1218f4d74c1f89f1ba42
z4b4afbc208102c501c5199dac27496c8d8325582dfb24de0cf68203502f161a4e98c5fa27b0995
zbcc435b6d5b0a9779f90526f16537a7fd90a58607be3a4412ff6ad63007ed3792efd9df76d2fd6
z173cebbe208db53e65fc724a22154ce49bcd499c323ffb739cc7d67007f11d345a1ad2758ec491
z1ec8343fb492715c80a6bf5b2c335da62649b8f2c02f72f28d145c101b0a6a05c26f08c0889418
z671dbfcd3f0cfe2d7da69131f87cd08db45e9188bd367390716ce45b20cbeaa31d84708ed4c0be
z90355a968af4458530cefcdcd78328db4a5c68bbdd56e869660f8c93d37a1b01a4cb6519cb16f3
z91ea79a5bdeb7e20a6c7f9448f223f95915e7b547f20f9b30080e2ebb3f291397941c836842266
z5c55c71a5cd60898461dd501f43a893851636d7e7a48b1acd14e437b1538e1811cd3ab5113ce9c
z3e291737cdaf08ca4dd24724f98a6811c90d5bae06b95f77132489121d25c08d9e77c1ac6d0cda
z9715e89bc130f52b80548773e8d1243c345944cbe273a4c8e7f8644310ae20fc09215f977043c9
z7a98b15ce0fd62802b921876c732292c6ec48373ca2a41fbeefae30ea6ec6bb963fafe498daa9c
z78233c98a4393253715bb0410f127bfacff1a131557751fb90f79c1ca407f4ec47f7c9b6c3b1f7
zec735feecda42d5847936dd6c0cea9aafd8d22cb02a95888755f73521a4d4a3056531cbeb30071
z49ac8da351944199ef9a1bb8701614a0da229b695271420f44d0b2fb0ed8dcc8eff1f41b618a9b
zafdeb513c8dd74d8d15163dc15a0541c38adabd2233ae86e4ffa00df5f5eefc70823ded0923d49
zdc4c70bc0d3732f0fe72250d48f1ad4d8c6126a49b6177fa5c71c67b46e8df128ae9d1b085195e
zf1f86f4f7a1d8ceaf587ee5d76a1a9b6b6c2d36e4d0c0fb94617066c6e7b2385a3a0880e39c83c
zff6c3bc1b044b482f1be0460b951950cf6466cad87dde3fdb0bd25b58057286437e57e87d0b12f
z6ad8da8d117103b99a07239c2b15dff497337697dd92b97650efea0ad392e92544a4339f7b8252
zcbfaa97c93fe8f69458406a550ceb86861fd18a99dfe65d8a0f2e5fd96ed57a2ca41160fa23afb
za29d8fb5da32fc70200b8ad123d0df2371f9b2a6b2d80ba2c3868e2a2465e7dc2b44addce944cb
z20afe02e4b02d192db7fd88b06fd04691fb3c035d75825b58dab40ec2958a582b9e58b35f8c582
z94f75bc38a386fa4595c5bb4f73b7c3a514a430d348ca29b3ef6532641a71941335cd1f5e191b7
z49529191751f3d8d9feea88ee00e4a3ae63f30e4ebc7b6c5b0bfc540792ac3e2e97f5d69a07979
z108fde4326abee5607aea1e3c900196c85b7b5a2b83806681b3032c70c6766ce30d93d31124b58
zb35b6b976db82f47e774101913618f8924a32d27ab4d7bc5fa1800d1f7497e766a0da07b7c2652
z94f20380231f749cdb3ddf467b72a6936c1cc06a6e15f6ce8d54bdab93fcb1323d178de2f5faf0
zee0135142fc6aa0c8d19b9ba88ad922200059cac591a83d187965920980c84f5713f57fbd38af9
zd01a6b6dd8b9718d382b560edd849a21d6955633a4595c524f24abe55a5343c9dd7836ec25f5b5
z596741027aa3f8ce91b19b9f5568ec94a7f6ffbefecbf75fd447cd7c6c10c53a44bf6010964640
z2190be911aa7d707bf87b07eeaa951109e368922a4aa447be1c84c10dd95f138c4cc7e9200b0bb
z5c4c0640f95ed6f01802a9aadb5cba21ee153d4082b198e68557def1fe16589b33657c3460f2d4
za03f9fc9cbc021206b84acaed23554792c5c7373def4de7f80f5416955deb3c783c840586e9482
zc8c90d7ed5d52f92ab4542efdbc5fffccbc34bd7bea2c39150f82ec706b339ae45df0d32940560
zc27556062c9955a9a6ef0767df3e346eb0ab794db42c468fcbad6a2627ee26182014220a1e380e
z0a1083179fda1c93a8578ac5deffb95706e75555411f3286981941aebf5daf6ca2a1adcd944118
z293fa0bf94af450320cb3caef1b59856cbfc526a0c11f3bf0272cfc9c12a3b0542922605c99493
z11c10b182407ab98760403729c85130a2cf59575a0965199866b94558ec26d4bd0a272f7eb9e50
z15bfccb570a47acea3cbfdd187919cff6b929b58872541743e18f8319c802decd0e0062497d516
z025021c22bfa7501002beb365bf514b6c6c674af077e6ee535b820249c3d3e33efe38dc68ad340
zc2e517827e317933f407be0fef86e7ecda34baebe847d590748f7d5e9a282d344eaf2ba53711ac
zc3c5624bba62edf7403d6fb116ffcda82c9841fd2b65fd7ef9e20a88592363f2c196fa4a12a29c
z99795de33231bdbad543c75d4695a8887fb29de025f405da160420b12ff598204188f83ee652e6
z9b4e64b8c99872644a7fcb5c345055a7f6ca096e707066c6293bd2d4ac5d6a6769855524de88a0
zc00c4542e79163e09fe39360f593c81bce30aecacccf2a8e0565ac1f2a13b28ac67ec9ca3b1775
zee2f9637ad32f0c3b0637d6e4eeda939e311cba7a135b00eee488adcc7e874bfd54c675ed759df
zdb25e34bccd63aac00e8d38be278c9b88eba30d47b3a2842395eaf3b41de28c403f57b72d1eed2
z2887b265eef506862758224100c3375e49574bab2de117e46bd3372a819b331d934a3accb6160c
ze01f56c5920b303d9b54619ab2c3967475b63179dd7c9b500295358f0d9a91d78916b48c1e2901
z98f0b334bbcbf63f6d8b678789ca20bf501e4ab9f21827b7f07a1f7746e9f739fbee3cd1c50b47
z09bb888847c1a6f22a35c55b6adf1e832784cd259dd0211dc5deb7a4f03a46de101816a416aab0
z412120f4ad21af90ad410237ea98354b62437130f3a91e25d8f586c10f75decdc70afb5a4c12a1
z6f6f5ee8212ebeabb663b42d6dbfde5395b66ee706090f6cd877af85347ad904a70ce3409e76b9
z15c68e7e7ccdc6c00424720eff4202e572a838e3f8bc2b69be607627cb2b87b836c262c607936c
z623bab53ac614483afec31aca7669fed472e32772db50ddd9986c73faf9fc46c10a2dafbfc71ac
za069af3c8fce4b80cf5925f24c882b1bf652c86a78d877652952221a6df70562344f8efdcb4f65
z224b9c0e6570e03342657625377d04e070da52f1f335607dd24670920d7d1f765e07df19b8f787
z3b9e35d56b6c44cb20a8f73ebf81f2efeb896e78cafa1ec1ae409166058bae08a1fc9759924c38
z40641e73e4b696da056684be7f23b91dfe86e0c8dcaf8e1e253c0ee4564be95b39890be6664e2d
ze7b2512e0062383164a372feabe0be4210b416a80079b0399c9cbc8645337912e49a733e0558ea
z5181e21eb2fb6ddd9569dc7becdc44cea11e9c0dd87e53df2d341ba21fae8906608050b84addd8
zc3b9696d68c6f4f60ef2cb05aab876664f49e9665f3ba71f316c0a311f158b391363f6048992e1
zac87d094539f8690819195b25e585d3417d53b6716ee0db2a1912ca9c082ab1788c180605d961b
z691f4f2b46b4842090bdf93ffe23b0f8f5c5c280ef36c81b6837d8062c4a967c943acb3ea0d822
zd64e6174f5fba995165ff5a7e83ffc85f50a1f2ea36b69562736928fb0a7cde67fd887aa4a46f3
z99e3639f35f57b44be6620e6338a1b7725f639400884c9c20f31f18e52495852586218d21697d7
z601c46fb020f972277c360d3e0e274e09e927f4215b335be63842487784e42867caf94c39ddc3b
z37e6e3047312afe73575e80cd5a5d106017a738d9b150d8e5c5b932dd7d74b48b85984e1d09c44
z144e4f73e6024095dbc5950978b6f54583705251b40cce3a144a45fe935525730b661244c0c634
z449768459028d8fee09fa108d9c82d7c11c5e3ab3038f16b5d7c8070a99e4f4376a545e7e66b08
z5abcf0d60c1c9461a8c63ad3dcc78bcd834a0e3f486e5d0bd299ce1ba134531d011ab63ebca4bb
z55f5bb386d28f08eeadbbe0bd2be933d2bac4fe634255a48dda3e8598f177e9936675c0d35b6bc
z48551100bbaea267a1b86a937a5703b5bd94cbde4f7b3ef50dcc915d32d63e8368098d393b06b9
z4e56fd2339a44188309a416b847e2b686129042ba5a09392515e0039923bb1964eab9b839564c7
ze3d03dbf1f91ad2938512b6f1cb02fcc3d11e709dc254f48bdb552067a71294b7d23a115f2417d
z4e36a2d2c40d67d74a05f60e7c63cd0c14d8267165643931081034bc9094cedaf339f7515a4c73
z74cf208b19e2af1ce2276fd09adfd6f4947b33b7bad5653ae9a1494f31e0b994df7222930541c0
z61e6af86faf60bc9711258f2fffc55f08581a180a97efa59d06926bf20a1175f1d5e33be81fddf
z02bb9da83fa10b2c79dd88f386d492fb99b63531d16f51d21beccb43aa260619e727ea946aad14
z0ab8a3c9013fd19b98319e3f83ce1a185032db6bfdd83cdd0bd206d155c4bcff115d3b27681c54
zae298f4f433dc7dd17af1c147aa4493f63a039bef57ab766508af5aea4b2107b8dd13627f50b22
z904ffaeeea9f07f375036434308753c6958b376f5ccd5a37001a2b57d6777d64c7c763e3bbec86
z01f2288007b6f96ddedf6404a2aab4eb20f88100debd2b944771a54e9853393d5c9adb379e433b
z6f60cd694000ef5300fce860509fe9646ea4a5cdf5d8f00d2e413d991a87d7ef046cc1c9d00ae8
zc320c640f349ff40c586dfc7efd5f4d1593b90f1e788ebc93eaed1951f95dc3afee038a96147a3
zb6c26f92be0561b4906b83105c926ea12a25f0cf89af1ef26f7bbf96ab214864c3060dd9edef72
z7bc915b5a96e53fcbe779bdf64fe0e41b9e275b9e8c063b0add51f13256357060b468f894ead4c
z48de613f4874f641e7060fe80c1d7361c13cc20d4cd6c44a51d76221d6990d07e9ff2459323867
z0361972f95fa8a190338ac09cb37b96918d2fb5c36a9fcfbd6a05a2421ad42cc067ea542194bf3
z0e0b6156bb0753c2948f6aca84d9038497537e0bbf3e68e75dad37ab7300dbf09d2b30941e0879
z997f336c9f9511b3fdbdbd6a5c0e2f312e2671a5a19a459d0d685dfe155d7f24881e08079c6036
z13a6526198daba7a1f66dbdd3ab5eb16d4e87ba119ca046d4b34b41bf4fdb6beeaf8e9330ad0e4
za5c525221a4ca0e7fb11913947e2b9afc08d7c42da6e847dde29100ada1f343fc1bfd37949e923
z3b5c88f1ba6e7da151301033676f522850d8ca07f96e2f2292ca9b6cd315996c09aaf3a184b68c
z2b62cd0dabc580e775cf24e630108c19c6a1ffea8002e3e9b6680c2d49c0e1b265987b4e7a0bbc
z3037959aef174724479361e699c9cb36e847d616d2426dc6902ff3503683acf998cde7feff6fb5
za76758bde54aeffd542c78069946055d2f4b62ca8529a23fb8b04a91afafbb6c26edfc8900e278
z4f2eaaf5644a5dfa7a1bbb5f7d6c26c893d4f4a9f3a8cde1e768967bcb1cd0ba38c97b561ced97
zf06a1a248ee9aa7427f525dcbfb395dabf449c5ee8d63e3a2eb854e6f3584d662d333a5db5d652
zac7f013f5bc737e27192e789fa7d6d71a0ac4aa8817a7fe45197807c494e417a969631f9ff9507
z8b7d29acb17647cb4c653b1414f2bc44491a1f6317b3a998462cef85dc4fb9ab4a652f5156cb42
z4062cc1049a42caa774e4590520449867f26d4460e50cf0fa79d974cb94b9188f00c30953533ae
z4d9aea2155fad0b88d35eac597ce364129639bc539fee27ec21a2c7f791e31a39956fc06cf8d19
z52c13c4801ee9484c7c3ff62e671d12d50dd44f323762078664895414e0c66625b230a4bf7af54
z39d38cd42f3e1a5b1129be28a7a0212f682b9ae7d853ac84271f398bf873d064a7a9a3cdc5d563
z9ce920288bf877d0566c8c4f8152c934a84323b3a5d47eafd4f27b3c59a0f5d9060aacd21099d4
zc00987af9af83b5f7bfcde3ecb89b52371536da66b84eeb564289a5d94d6ee49bfdda9cf9ab70b
z75855fefc63364d0feff593bce688bb396eacbc7f822dee078fcd77ff5d9290aaab56de091a894
z1f2103d35179ead5b25ce94159ac48bd510ecbd04b30969a6574820fa868bdc7921c080a6fedac
z6901fe4361f02e6d6bcfd9ee85006643151d9843a7a58547bdbc2489da760c5372e0525ed32785
z3fd77331a55064916019d55c69344744874278772a6d2ffacf63c04b9b5c4915254163eda6d397
ze37fc3cf28390f5c6941b182f9c0a69b2861b6965c27c074f294ae4a7843d1e160551b1a87e351
z786ccbf86300eafe2302264e6805e0ac9e7d569e75671f9e03659690b1753cb943cf6f155bf6ba
zf005257d6170c6a0cef3699c47209768aa1e6d1b751b9c66f99753c9b66451a3511419e71b6eef
z0dc63699744d34710db06631112ec64d61c234ffbc35f787e0b533ab2264d471903deef4172b03
z3f3d00e08d7f884c39bf8c46cbdd13767d000affe67dd9e4cdb27c59fa113cb64343552ef8fb82
zaf3d025582f23b80a6609669822af6f7e61771ca6610f8ccde456951aa1ec8a3a492a3ca126f4e
zf751423d151a29d2233a242f2dbbbe3001c5ca8768bb65f0f73f58972a1a2770166bdb1bdbeb9c
z2ec426ce0fee7b86a6ddf1c6f2af274e802aad5bc2667f1604fae2818d47c0d099bdab97029511
z0c508cc1be3d6e0becca8e0ea5c21866e650d4545622126f18679af343d0b94e232a36ed457530
z7d86bb9f2319f2bc2a1e0f0033cf9007e8c32401087c9e1ad8cbace617b358b54a387526edd30c
zbcb6d7706736808acaaf880ba7deecf51e39c9e9d1535b3e5f1e7b68f55d9cb5666e0638889bfe
z6544170fd8ee09d7b3289889996216d8113aeda8e3ce8a25cb1cb6873141f5160e781a0c18829e
z05b5a0c87465d650c602055fed2ce18e58f11239d0e48d7e70d8f0a80f91343f64bf541b248925
z08edb40a72ae07b3fd19a200cf6e38a90503255a31cb59fe241cdb94cd396f2f645dbe3fb76318
zafa9fe53805042845beeb380a32f73cc5b2dc4defcd2960fa7e625015e5c709141fd0d3c0fa3e6
z06df7884a51a376e3a9120bde5e3a6009cdd717a6e66a3b2d3277a96c4da00088b0fbca8a71a2c
ze5cb7bc8bb0dc49239e12c0d8a58a31eef73bb35926076d6f86ba2546dfc5deeb74c2b4acd4261
za449d6b17f6248522dc453b29b61bb1d4673c3c011e1a648ccddc584e7aac383cdcabf0b117545
z5624d77ba688d8a17b2bb74a759b3081cdbb126e9a53e99a4724d70348fe3bec45a7918b2812fd
z2ebb5770f186fbcc241325a2825890687901738745fa5a18bde05d871c5e41b71336be79be8f52
zffe59d71b1278c39e965c8fd83ff3b0e9f9f22a9cec513ba445c3bf8a6c82890fa300e7e939113
zbc3930e9cd8ded466812f277338dbf9239cff64af9d3e9680c94ca4a2ab781b21d110cfc15535f
zb87333e7e60a87730144ee0207019883777c9d3d82c41f1f7de92d7552ab47ceae9d3f98c6b08d
z2a814f357276f32457c83b6ed6fdd1e7b1ea448802db4df9ba1ca004a3a179a5e7cdada2241016
z900f9aa829a4e4bcb0a5afd8cae5b23bd50f3bacf394f193817b1daf6be52cf1c09324491f3a78
zd2356a2335060c9b6be5e3bf60cd0e8e716a38f7d94be664d083f51873e80d2227df87e83544cc
zbee5207d4e6ca3832684c1ae83bd627db255d86d87f24e52ef4ce7449101fbd4c75b55b3f4ec9d
z9be03b939ab7ca41358f643c8199b54e3ab556bd89ddf16d678515f03c05daa908482003251976
z670e38f2e581a880be3ea9281179cd4890dd54ee728d12fb860788e7dda1dc01c36b5a553a2ee4
z445c400213a8b155247c32586236cebc40f80e31acd82a306f8c29f0fb4e82476c23a6b60cea46
zfd34fc16e786371d31521b0d89ba8f0c2479b40f5c370bc5d21437ab92f2d4351684cabee0b162
z045412c87e5953917593527641ba3bd33f1d8d3adc7ea3707bc72d1f50477bffc358d58eba156c
z6ca80edc83f78598bf239f68770b0d309770fed4f374d66f98f45af6563449076bfd2f0095a856
z6edfda20488f4ed29f3633c69ed22e8a9f5629e00032bb7915b0253416d42641bde19e5bfa8308
zf091d49096cd61706dcd5fc559af733a33bb4e525284365b9bc7c779da81a160c07988400337e5
zb45bb263130497f4affd3fd7d2d859c90abf7e1ece4b3f120e3a12bfbe7c12f5c16189ebb442d1
z073e81624bcff5a541fc7d5955574ff4383c85e7f4f57370bacc3eae17f010f07f12b57bcce855
z5cb68815e5144aa774164725938dbfc603b5102b334c05a49a5bcdfa5ae062eca6a75778a5c670
z88fdc5db21ca872c87e48ff746ef0ff28e08d71032123265d88a1b8fb4513c169d5b79a0bc2462
z4c12be50be76908d6f0566edc466d315d9b374855024e62cd74ed64cdeef345987bce2e81cbc24
zc8b5ae662340702b972facf40c0495b9d4910b7bbd0572d20b0daf25a82fecb73e55e18e3a91cc
z7089969120298c7f1b57c706269aea5b4283c5518b23c5e497d02d9a733f691d309c0e73221ea6
z82be96af6e30b389a0049ce3aead7a0a47e7bdfaf35a8724f1f53162cdf2e4bf98c87f0a8166f7
za22c5755cb13e8c1358b2bfdd30fa3e1100a2bef233ff8186eaf73fdb839f8e1b73658862be306
zd720e28d609099317e78d47b3f9e201de5d5856a020ec30f60829ec0d8d4f92d5ee1a3ce1d1aa5
z7904317bdb2f57645582806c0cf67cf9ff58a268d672a2ff6a21e5420a40632df82d3c822ffb54
z53bd91a4e051abd03dcf309edf23cd4ad8d2fb6ff7efda3eeed7e6799558cd399dc7260a9290ae
zad6d031a8733fe89aea43ce0ec3e97f004f73096c9cee379e70863445b82bbddd9d2ac623720df
z9a91aba2734b1cbc6aca80ca102604f7f8b83768f6771cbe860023c97e5531798b8de696ea07be
za535972929f3b2a0f434c2fd1a3e2b64c6b5cadb7530d265eaf3fa992a57d06161a54b6b053c2a
z9eb90e5e35bea053b8f72f849a3444c7def144c41a994446e62bdf10e7cf4b5db195374f212d6c
ze17ffd9ed2818c3ea857d54a6764424035a126c49084b8d73aa1679a19c21af406ea4152097a2d
z2b60edfd818fec4fa60e390480d9e769e232f4b189168917b151db766374325631c7651431c8a9
z2ce89cbe6d89b1877781873303856d3299f56f9aba91638d8a533afa886c92771b5325fe6870d4
z9ec094df336f3203aef94952b7fb74a91192d5bfe563632b2321bff38baee139077390d75fea6a
z42e68869f55c05e4498e7d54aec33c3781dc457040e0e9650c8baa419ffddf2ee42eaf9911503d
z2ab3a2172b0f4ba9eadee8448b24bc4388350243ab489b519c6c0540886a4da75b854915038be2
z22720d2042dd9566c132f9c2633779f0861fed20efb1e2ca88e12226e7ad374e31bedb97e07678
ze0dad5ff70384f157b2c55157dab7f74042bbb18cb6599ef71f19f20673dbb92b5768ad030f3bf
z5f3dec1406326c97bc79c92c8a6946bc5e6093f2ee2a6836a839a3a31c535b2b663ac66d828c03
z9674cfe4cbc5575cac34f83345fe868edd4015f11362149215c5aba9a7ceecf1bbf91d969caaf0
zc29ce0f43d9ad49dc7b7112e45cffce0724499d5b3b151fc62b90f6df382270ea9c525f118da60
z20928b9768e4a6ed00f8582c74086e7ed0cea12c26b75a9e591b05d174dde48f58aa7a96e74001
z3e6aa300b563f09eb0036b15cd7af75cbed0b1186ccfb8f47b6050977fc96849870b787c4e215b
zb08ddb45b3c6c296ac4a1e88730a0b9912fd7e6c427389a3ec29c965ef2f6748fcb9d6e463dbf1
z0cec5a7e7523ba50f6ba0cdb63e2bc6dbaf4c6c03a5dd38eaa7a762f92a95c9fd17267c87bf23f
z67a1ea6e468e8d300daeaf7f90133a6fd836e332ae35d8eb6067fe824c43514c776e34e0041715
zf65c4fb08993032a43d632f1b077dec553c34f54ffaa33a1592dc6f7a4444999e72223b56182d1
z0c13a496894d1433da665b329dcf4cb54886330fa7c9431adfb134b4683906594261131918537d
z02b123bc5a2f4939e6bed345f4ad305f7b295e9eb99be935cb293375fd391d074ee7f3dd58cf10
zbb901116d8e6a2d55f5f9576268006a533f1f39ce5c1a6b2e200216094ad70520d0dbc2f1fb694
zf05b7c46f85f2691c564f106f51d222b0c276935a364346bad72e010b7f04f07f3452f663a6f8f
zc64fc99c5516ef0c0bf51cc96adf29c7906139f5a87519ed974ae2e92e811c27c66410bca66b47
z6a1babe9daa9da2aa7bfb73fccafb3fd0d4d0ac253746fea3285b087f0e0922abb29f55084d6e5
z31978789ed75c775ffffb1c042f506767137d56335c196359de8dd7613ef75b836bbe38d8c52cc
z230bf32226a289c288c5c8048cf7c9e4a45f4204008e5b65e4ba5b35463f5775d8e66e1f5a4d65
zfc4f1085ed493a6e4f02ed7a3d2cf529ee2b825a016fee59ab07d560488f8ea868522815671c37
zea8fdadf44c4b554ad3d03efd614d2cb61741fac1ddf6555a8c10bf38402b3e747f202db8c0d9e
z336fc56827d73fe1b424f009aa9679ea4666a1f40e816c0a994fbd3d70fb508ac99749ea0d685c
zac13e79fc0df9f1ce76c859121a87a49cc4841a9984573d27052670d0040248510801620335502
z28478f90c6ef7cab2764bf745512c7876dc9a1ca1592480332a4c47d7b5de6ed96e4fb29cef767
z4a3575a0d568ae7721745218649443f5f24836b625be1afa6e0f3ebdcd29b82c117c16c862e943
z93a2c9c1bd5919eccda4bf86065514bf21ff9c079a0abc85d351707ebb5172de8c099a390075d1
ze56e6db89e91217dd4099700925fcb8af45eef5a463aed12c0dbeff2e33661c8b3ff5ad110db4e
z753417926a72eddec478f3be8806a25ac0ef045d2f99ee06e879bed87e1eaade6bf1d6822c73fb
z954a8e24aa9fb7aca6d95f82d7dedb60fbec8d057097614cfe2a7e5d60bb506b8d0b796b1c7de7
z34a6537d472977fd115b694aed7a70f2a9e80f7980d31ff1124717bb41a4fbbd27176e30212aca
z7ba8b04e8153745ed946b7bd22706e87fee29d4aca5deb68866a40e6441aefb0acbbc8841cd7f3
z8ead54a8e303f61f711cedeabfa3631abca86c5b1860570d864559724d41af8ce9b3b98d1e2c1c
z37d6cdc2f0b0d3adeb8ed8492ee83b8b3f8c3c5b1f23425914c634f5a93271b1e499ecca167886
zf3196bb2fcf996c891cac293c08602824a7dc9a67ba4606cc7919aeb29d8761122556f41f03165
zcc26e417fab93024b3871da51c0d7640f7ea6485f7a7e50e1d3a211a73908937d2e73d02ed340e
zba454683d73bd6dbebd0aa2717cc1a457da8f0eb043fc1c4df6bed67465a680595ee9c27fad843
z8bd905b32f9239b3ba84aa53802d95184ccb9f165a4cc1ba83bb6ac44fc2d15ab0411d72bc0f4a
zefdffce290d01fa7f815d9178ab88022e8a40095fac80651e3a10b5bec294f364a996614bb86e1
zc104379a06ab5afdfc2325cd2c7eaac7e6d72c8e21cdc2f2513dfb71720896e1e12654620317a8
z6b67e3a8dd52fc0c5d789a18b19332e7d3af295979587c11ff991d80c43965d478527ff24afdc2
z497fd1df6884a6e44feb1974ebd7c50e5859f5f6fbb4d6ce03bb56d33cae3eb9c506f5bfcb79a1
z716a78efa7ba6f3ee58b85eb13d0cd1c47c40c2848331ca8fa93f779c9f2c7bd3b4527cc8ed60d
zb71b2cecea3dbe44a73e5574bcfd6cfa11208669b689f307562e9aa4b3d4ebdc465c65da2a1619
zaf3ca3c60dbd7e825d50def7276eb025142b8ec4eca420fba28aaa9f3386d9bfe4e099f5c91098
z34c5d4b8707fc8047c5a37e841c2ddd05e27f77191acd61fb0fadd6ba241901f7fb4470a1a55ef
z1bc717f8747fc5298c21663c3cf5f3ee36d05d1fc5c6974edcd43072cb4931399f832a36af65ad
z544e4f498d9aaad34691e3f39684eae030bea9a3a3eef344362ecb5e8fa416512e9552f7373938
z5748ff7ebe1851f879f6288286b2dc0bbc0abbb476ca9c4d1aefcb99d468708e107f6b1cac5b23
ze662317ea1ac595a039a09738626d8aba10e997e41aed6bbe9a9013b649d6609b87aafd2728083
z039ebdfd324437c6233b50a3b36d1d98e29fab8c55e46c993e158de1b40d4bdc11eeaa0366cd43
z17f0eb50d2a51954561a59eeb63b640a8f9410ed902772183d0b6eaccb330c9300f83f64f6bc72
z671a094798b6df9461af68c458d0ce836e81a6caeea6cf8325251edd8f1387d0ac7a90226402ff
z6d418d78b10ab86d097cabc557d8745d5e3abbfbc7b62a9435e9577883b46dc5be1942f584f895
zebecd477c87e2e8e229e844d5feb611a729f210281d85f86b81eb14fb3eb83965cc1511d9d093a
z3247d737ebae6e963ed49c6f6e6e68779429c7370722960581e586adcfd55b3aeb3d926e9b5138
zda4e7c5faa6daba8b0b44e0124a238a383c51f59dbd18934d5c97be5c497d23f5d127d62530a47
z6e16bfc246b473e1676247e071bbe357b49ae5def919f08d1df952350aab4cc3f9574334076fcc
zd5778d294bcc12e5d83204aa8beab48956aca4ec9dbcd4fe318199cacddcedb8c64b90618df2a9
z7cf175aa19f0b590178a7f54614ecbfa01f04af40254c8422566fa31338549b818dfdf8a6363a6
z59be7efd5ce5761c24c5ec48f1c972114f293adf09d57f982ca9d4454536a4fc650204ece83fd5
z28a34517f03c865a3347db8c163721104d055910b2d6ae8ac8214bf24561f9e2e65e041ee78eac
z2d70a86584500bea082c1860c6fbc8935fc0372688e9ea137f114402aaa8d5c8ffc6609f8fa705
zb159529686115c18f6cc32d9c588fffead9d10e7e90be912f21dd786c49786b1c071fa38205ae2
z503f11407d5a986761daec3f3b72a4ae2429ecc9770b6d595c0da8018d963f6934d6b3d3217bf3
z8108a98895df664cf35ba28ae704b0ca4f98a4ab1b0bc33ce1af34a0f3b5a32f84889107dcd6dd
z194588cdcfd4aa80205d2310b7dc8ed902416bf3e6f61daa31a45fd9ebbe8788095798f7105087
z254d33b0ab9f0ce65c9ac79593bf28dca026614f60a40c31e725c51aad5fcd6c0cb8b0d78b61de
z1bfd4fb0d42a99aa62237ae04d7ce398c8c629a8536ec1cea6fea5df2e84533f34b2ad52891fb3
z4a33109c58fd8ae855aea2422e0867515f10cba30b89c655063f78daf039ddefdd9c8ab01dabea
z5c77386890b479d23388ba17ed26bd410db927dfc0e0b97b9df53286b8c53b9823bcc05a8ee399
zcb453b30b4064993f3d08e02e8e5d7cbdf3f2f66ea6da239f428142931a04b3be831c1f05778cd
z15d1460bd3e033e1c85873b80167e0ecd9ef250c0d6c15873be379966aa478f510422b413e5afb
z419447f33607b0ad5325ce8b4ef4b8302928eef185191767977b00fc71f90b0b66d172f2943db2
z4eeeec622227b8c027f2ef125e4f25a84b33971c3d9d4671ea5b219e55323ec00a0b5a96b601d4
zf6b6f638981176d800441e05e8ecd828a6d8827217e87de11974b30837444adc445f42fcf4d5d4
z0943675acab864ac6f045afec394c8efdd2326c3eb3bd56beb21d20743cd63801bdbd99310675f
z5c8fe6d6dc92ae1fbb06ab5d936078129bbbe6aea25c2bfc1c5eaf012ffbbfea03d638d5f277f3
z63407eda19cceb7ec8e78f7d4ce9c9c3b016322e6122551254b52c343551cb3099a699ac612974
z9a18bf23463e61ba6c416dce8e708a2dcdc69d4ad39d68e6b900b3e59da529d0917e9d84fd35b5
z012fc4e14d2c76be769a9e5e9ea286c5fb2a6987fc4895c9132fc6301c3b51266a8550cd5c0c62
zd333f2d5e717ff4a077b88a0b92667b30b111d66ff325e2b692e2c64148d9da7d7814d48ecd88d
z746c27c13ba940207c3a76521796dd761695808e101cc6bd9f159ef82aa75cff1e2df28832bdde
zca62a4d840b40118b88f575c1ea0fe490260f80b64ae9a130082fc5e91d3f965b9b04711007605
z483e6506f4addee19c3796eab7935ba713bb72432655bc728b04582f6711f6de25646d9cb28099
z628fab1d29dcf7504399bd7af39a37b28627e74454fcef912e177c24a493163f9a844ceef9c684
z58142c7896a8b46b8e2cd9cdd814517b65ebf22008c6998f156593879cbcfed88fe3f2a5010a23
zf1a379237afc84b6939d9757e266f0ef6f02897b06a3a64aa898d2ae108d5db9e343784b9a0f58
z93e8283d3666577153df5b6973aada6d695f5fe5bd311d1670f8d3a5268f9f30e15a4d58f0d372
z382858e36b5de04ab886613020f5f483259bfabbbeb567301ef68c54f114c15ebf3dc9404463e6
z81a064aef6b084e530a0366ba962bd59058691dbaeeadfef2d206ed58cb99d3a5ddcd857c44244
z44617d42557442256f2b1afceccfc9ee3e9a763690268f9c76f34a2411c32180ab40ece4f9b3ba
z418e1017c041233e6d6cc0b56e1e99dc4752fcf228039ad3993b55a4d6e5dc5ad4f4ecb24af8a2
z088ad6e372112d53ca3b807a4c250e4577ac8f78369e004a61d0ba5395c87233feb0b31f3f9341
z310e6e64d5e42dd6704828ac82ff840b9ebfdce0bfcd34125a53d1d2263c4a02e239b2264ec0cf
z56797cff927d8dc28e68cddaed64907ce5fccd8d12adf95b9681efeb038e379654ffde7e50e79a
zdb6d3a78e66672b44e6f86058008eacb08cddb729cf5021bc399cabfd62f6d739290264519277d
z4bb8c73a41ea6d7f65705872baf0f7bdee7fa5f97b7f35b820f0b876dd5fa1bd1bbc2059d6e4ec
z116f25d0491831e59410a107574219e4d94a1a6a66e975eeb3a2765b96ba2aff9570752ff25529
zb12744ea476512fd3f1a916157a8982f457a26c7c0d9c4cb72de894dc02fe4bb8d5aaf212b2170
z0de9fd9d494379f4127507571138292dc9ecc1d76685ec1b23eafd2ff624ae36ec177acbf028a2
zfc4656dddf40921c2559d84bfa5d8c344977b0502dd6ae3adca740c192dfc08bd2ffb8f38edf4b
z4bde366d3e7c7b2b4913c3fc49295c3f6ebebc1ab6ca5a503acd40cab83d5aa27dd59e7bdb3274
zc1f560e1e47ddd367506e99caf982459961f43076f0cebdafa774a02e960de455939fe8c0c6ee8
z59102bd5029c104855202408972606e503b671b4b4d498d79d0172d56b181b08ff61be6c523743
zd5528b43d005bb64a92479886b96b822292e8b1e2c1e5c66ed0149b9fb07fcc8a935f726de00cf
z3768f8ad3c6a34348628f50431e3715c11e85ee0b6ea582afcb893f2545eab0480f187b89d8aad
z441fb5fcbe6cbff98c37d27b85d06a7506913bd892848702b991a762f694df3791ac003b104eb6
zb9b804c4cb90c1e9e9762d44f1f306ce15e3342a7c0fa25bab3dcefa079757da3ded5dc7ae210a
z29e1f84dce8c8548be0815dad621da6e7a2da0ffc8488bb44a3ead9d4721fbb0ac99db27d047ac
z33d6d1eb3908ac2a82f2913e8f3a1ea2a6f06f4a6a95dad6ae206c93b0d629bcc19b9d286d8714
z81652d82475617ed09bbce3ab1de0a62457e6ec932009aabe0b4e7ab6a2ec630049fa1e4d0e1c2
z9bbe5815f77064624110c36f632dde91323e12658b0e1ca21f836304a67dac707e852acdd5183e
z7860d797adce71b37d76266ab34c14509ae0dfdf02798daab413e3cabc24f047a816746e538721
z0b7c5d1a25d7f38609622773e4b302da2dafd427261c58127f7673d181445b656e3cd6e72f1f79
zbe7b2085c5f85aa21c77ef10838ad48f2d0ccb739049dadc060d450cca954136ff2226f27822f8
z29692c4b9f92eb7348b021fb4ba43533e7cb26fa82190e1de323e6ac10b703c742ba78ee7ed833
zef209f4ebba5da506124d156d444ba339b05cd276b7a821c8c6fec4453aa412f5bf01c57fd18c7
z9433557647f838f2d884bc966e78ceebe1901be08abf2eed57babf96064732b3f3c0e869d746b4
zdb72571a5bca6f747c850837a86580efcfb2aae2e49862efeaebca320de508a5dadabf5d4bfbe7
zaf0e78930b8775f0534f0c0e521178ed5b59b4c0cbb8c5b04b14dea92fe89b7b83adb1856b1d5a
zd12bb837331134fa0bfcb5e8249e5e977aab869c22307ad3cbb11fe6f8618430bb5b5bd4b56d7c
zcb083eacff52e7798a504c537b07e1f600465c8ad9eea36566d2f74aa5e14da2102a038d33ec04
z22d2e238435e55fc3b3b5cee5d40fc4463dc8febd58c8d62476c5bb61a83d1ffadbc978e375a1b
ze2c59c73045a7dc025146910ee186df61913a1594709868d2f0d726dbf8993f32daa63b4b02bce
zf21055b4f298d2bd5ec14ff9f9e48c85b1744ff8772034765429fe8961c128e7f8e78cc8f28dd0
zae6e03ac3049f52637c9c5970ededba300359dd6af330617936b6eaf8c1825ff71fe62ac26c558
z2923104163071830c44e5746e06d374f47667c1ce8145ab3e01d3b4c90d96693e0ed60194e8186
zd76db021a3f784fa01f81e4a6b71c24fa61d47040bd1aba1a4b38cf38c59e1a75c8ca797c2903c
z9e927c7ad27ff9e2395d94b3399a8a8771dcaee8850ff7ebf079f2caf2f2fea2c20cddb7dc9439
zaea9825ab8914803d0ca289d9b8f86a4203fc6df356f0f762e05a305aa04ebc4b5e93f0e52f0f6
z8d61cbb8b104acd17bbc3631790bfdec4f62e07917bb0f6462ffd65c84e5dd150a11963fa487b5
z401cbf559fc16a3b90c75d65c7fa4eeaaff7c3c0821ed1982b1a5d31740acd11ac23fbdc0d0e6d
z6f13a4b5f17b43448dc0a001a5dacec20955f8af26fcd9177be3ed88ab69a2128ab7e7379d9c1b
zace6159f4c14a825e5a1ee593902c8617b2c81e4e2e45618c62ddf64ad6290c0e22b7c1160dfa0
z1a643543a47ee13b25aa3a9c66321f5ebf487bf0a757eb4941ede1d3cc935898b90e0b5849ff9c
z1d3d991e12db180e02427951ca8eac570b0ec5be119c7fb63b1f495689abed05eb756abdd32aa5
z1e3631cc26c2e68a9beb6eed72b0d3b22721300152102b29a5758d8f051e1326ebc192caf9cb2f
zc34f597dc99fa0cb8aa4fcb190f78ef06d2e9343f02db56da8fb1c0b90357f6320fa545088b8d5
z1952705bec7c2475272a560a8d3575323b3fe9646391408fdba590115a73947c20d581edf3d59d
z4ac020b9d36b8a49c076cc8ac24f3ee48bedbca040bbe34e88939d3db2baa3b8b0938633df89b5
z9def59b22b1a5abdcf6319ddd668460f7339e5fdba32989fe0417f400b1ee0a70bc0b599f1c74f
zd5628fdfbce0511a56857c40b0cbc153bbfb94ed55312d0e50f3345a773504b8c9444be034b94d
zc3381549aec71374763d3ada7ba310e51be4dad09b12bdf7020da545be7fd3de0c268528b51866
z64f07c0147febfa722614da861b96f2d772f914dd790063b87799a6472298e3337fc22ef90f736
zed4c6255194ed174df241cae94531a7daba201866c9bb2f9660564ee4f29c713b79476a1d32347
z1c420792d6655f281934671488434356ba0dde76c6fd7892a66991e49121a040fc1c584f86ca7e
zc47843913cf0cd6f5cdbfd778c50f95d7633e95ca41cd9a95727d0772496ece0f23f3d69686e6a
z13af102af82753da239cdcdc1b9d2374d6ab8d24eabe665bbccb34f54d621bf42b369e23fcc209
zfe69919672c46b0dcbabf8cd525b1e80e98455cdc27613026fff6a23368b030266fc9c19906146
zfce80274f18f3d5e1d8488084202b2af7e0046ba54068ac3fc325f2a758b8c5f3894130a0e4a76
z5891fb97817dcc02755f355c17f721fe0b1fd5efe0dfd44ca5ada77f3617b6c2b5a9a55bec691f
zd5091b62dcef66c33e8c373586f37faefb4d017cb8683ec9081dbbec92074a0c827caae2f20686
z99672e66117e53160ef6c2f6cef7caadd03d007de47682dcc40db5227d3a8aea96ed516de7a598
zf967e3359936c14ac50ae3e1041737b0b8dcc888af5d1593ea0eadeaf791707d7fe34adb5e635f
zf963338b59119e239c9fd24dd6ac1adb24febc4e6245a9219454fa1631394988886248a092f06f
z18cd4e7ffc91b0f59309c6aee74dc84146cbed75844beec99eba71bcf67e4f9bccb31ab001e81c
zecd592b92645d6cbb1f72e07e1ce82498c9be63383a3e4c5570026489e64d86a620acbeca93deb
z625c4dcef409a9da4c9d5a7bf0c5556a2de1fd9ee99d18c2ec4a395318c6105cfe2da143211ead
zb33d16f8c6c0c94b10c9e236c01e3d233d76c21950751a9494ca6befc0aa447a55baa951f99ced
z8d781e076cceb2192278f02800d57aa3f55dd8e9d3f03d4878a5e84555f59310ce54324a5e6f0a
za5a3d7fcab966d9f895838369dba7bf9f7d74d1ad01660b218ab3ef9d2ec96697edaea84f6882c
ze8ca7524b29e9bb0dd89226c781dcd75bc895b63239e24c9123a322d0a629554a67d9672ac2243
z4a2932f7b80d52a3c947a853d86f2920a2dc25705c1d7ef81b93a396f2d3fe62d95fb9add5046e
zb6e81f8103b50adc9175577e7349dbec34def04252ef8f294e1f22695431bf86199329caee3483
z15e2799e5e5ab174b3acdd6fdba0c98f0b63d40a4df9b288f133f5139755e07183f9aa1e151aa9
z930a7039661c32e51d1b893c9d967011e3f0e91dd9d4ab8d11f69385f93cb0b0bd7b6a11eceb9b
z04ecce6c27c6ebcd5967b686f046ebc37adb1f93d0644080c95466d5282ec06cf0324b3a14771e
z3e84f1d9764b8c0db654f668389ac23715ba6557176ff665f50fc0970aea54d2fcd94f3c7efa1b
zf5ca683aa5496287a2b602e506df293c107b57834b09ee9554efa377a84ee4a3f8511df27ddc0e
z06850e0eb7754b99885e9dbedd6e1b35fbcb73f122cd758d4cbcefc5e1974fb27cc6596cacc676
za7d32e5c4d35f71d6a76354091e5229d5bf1bed1bfaf0d6da40812b7b245943322d626bc8e9d4b
z1472db4ae5037d0fd49bb9680c0cdfb60decf764b05b4aaf18ab09c01650d6e344bdf2b6828cb2
z1545d11c03626f537153070f8def981f291839bcc1909fe4e67172661a6b82c378355d0056adfd
z9b220fa748f55c36102f6c0e7f24215e55dbff380a37fda669113cba739af93ebaf0ed154d25ef
z63ef8efea975a6f13822b5cf66ba3d11c8e53dcf8635e08eeefa24e1805608e1778dcf2c61dd0e
z9aef1f34a6b399796c050da438eae808e0e86cd16d24e48e1837731438b7cab6ca2365ace4084d
z1443bf7b22fda5e0771110b4e7b37a21896db5475ed58928323c613fd65122bb43e8cf3de56b28
z02ba21669546bf67a51eb320705517391444952d1730b1a9f94698d489ad1e5e584d1b150d8ae6
zda99339b1fce5e209da652badde1cf647df24fdf1e6ba900c252e3fe66d775b2b221aee7cf63f4
z7fb2a4af658293e4c974aad9620e404bc481e845c4db785d7970282daae6b3f832703461440406
zdb30c56423dd92e3503a3090d7c505cd12004d5023e319e1603fa23252c8e69db769c4b79552f4
z3e108ffd94bab44ccaee80237a9b7ba4f63f2b74f55187e1cb959f72c7bfe9b7d755bc3b58f10e
z36239c21ebb09e835213757ea9b5d1c04f8c204ba50eb68a48d6329b1daf0d1593bde47eef6170
z95d54163ce9ed6e91904c5fb1d1a37bb7dbedcccafa188552901f9d3fd3132f6ff0fbfde900aee
za083bae621a62c16bb47c1e0d83106468358b2995ca6197c71597a66b4035436c7663a2433fe5e
z1c323d61fbc89942a3d2130e6fdd40e4176ef8252a5897a29b463d697b0ea9365693192cc605cd
z55aed31c52748c29876b9a64fcf5ef6c2936fdd65737d12312582cdb2185986f5588d9758a5200
zefcb56871d010a249a5066250a831c2daaa04c72eb2fdc04aa12834553295aa5767945ff4a114d
zba3261c2decaaf768cfcc41db8a03da85078a09726eadb576e2c2ef40c943df2b9f659041755f6
z1922ae0c7136b4d79061b8950f5f613f3a443f1da92508000df08914605b60d0c8b560322e9041
z29cda0f25db9c19077292e50d692954fc2512572028fdb7c66cbcf6a222ceacd2ee0da7cfe6f70
z32d5202a91b4fe1b53e9e2b5cfb8a35967b669fe85759f1928e2fd470e8d36c41bb6a7d13d3c6c
z8b53626616795a83f6a5a9bcd616f9b1cbb96843f1c32e3ed94ac6524ba334f15fd4f88a06c38c
z0cb6452dca2e3c1bd43e40e7db8ea0353937a46109801fa3e1661ae7870dfd256e8e5ec8ff66fe
z3071e0d41fc7941a9e6d3009720bf7d104cf7b53bc582f973311f688d0dbe49ae2ad5ca35b76f8
za4dc93029c6a609bfad86a70c6a261aa0e30c79b2450f3734c090df78e7ec4711c87a1b4e3120e
zb69a64c1333735a14ea5d5cf55fea6a34fcb0272562fe3809c4a48e77a960d77084881b78a54f5
zc8b18a82dcf5f899b51e95e493c648ae9bc0ae74c1e58fd626de6a48ada2ce3a1dbe7516dc4c28
za5ec13fbd2fa2bbeea8b62cad29f1b45da5104b306a32cd59b38c89422ccc11a080aec338e06bc
za8bd3d6d84493227fb3dece296e61bb78813468f3e90b49d66c843b5e077c81f1f726f0aeb7023
za8d210ccff9420461b07d589026f8274adf9b27476b86df3be093a2e1b301f6cba3d4de7e0614e
zdecf0d49809f47311d0b2958d451cd0d650b2951380bc04b32f24e942ac97fd661b01b537021cf
zb5d1f9b3be21c0f88c57a493bf958e3e4e71cea81d5df2baae9642b50115e5867c2e650c7cf0ed
ze67c1ed994d745c58d71030c872b59d51dd782233bb12c240336fe279f4ba5c7bce355429e0d45
zf8bceecc852b70465b67b5239a94de74d3b3c47a0c878129a4ca86227c92286d4beefdaf9a8767
zecfc1ad58abffc6e142593388f32735b2dc51c88fddf2aeefd7fe9971207c4189cab8d43063807
z2b5b137d13de2d96e1a5c1f4326feb80f5d0738d31e6e90689cf7335d5a5b9c09bd5fc97c0b2c5
zc47baceb084366514dbd9ac261516117326cb33285f545eb84f29a27cfe621b67b83c633f25654
z1c71f08f12061ddb1efd35cc80f3a7ddf228826706e287ff9931cf21438c430a037eb8d411270b
z9f76d49b88b34089fba5cc4b5e40bcb689ebb1237bcaa03a694d0191ec50eb284db77fd6bc569b
z2877dc04301a6af642eed31ba6b5ebea8f677bc49a9c0e340430de6d7be1fd10ac6b60b1e8ae3f
zc141d94e462e402b8f2f65a2206a925a79afeef876bd193102796a73f3d497c0fd4876520a7449
z5d9504427a72ad66a24793777abf2505b2ef2fcbf15a70711f3b136ab988764cfe37cadc8ae24e
zd671a6d96b48d0fefabf12cd815d0be10808f8ab4c0fcbef493ea9070f5bad3f4010f540e279fd
zba8a1413d8e0bc983f680af8e7b1dcd8ee4da7df4174ed59780f67ed9920b9892c76929e9dc4e9
zd54b8117c0b7ff4b72f5142c411d4b9311cd73045f8694fe4f9e5557c32f0dd3488cd9d5b8903a
za7baeb29a59bff45f587a466db715273b1fa119d77923d80b577f6fef54895fda9de1bb503d380
zba02d55feca661df8726b56c0489669975f83b4db666f130c64dff39255a5e933d28cb55c676a2
z864f05c182ab53f4aaae1bf7e00ce1592486d9951dd3072064f079dbe8bac1e7e6e5e34ced80fa
zfda27e5a33539b3fd32b0c6e62159c182063b4201432eb7c3979edbb35c8b8d168768c514fa58b
z847903d90d95669eb640131930fe4ba524150ed1eadcd96f392f82379b02f97117bb822807a11d
z72ce3df205f6df717b09ef77953b3867fe2234b8d414b0a421364666d333521e3880e3e2718c75
zdab2e7cbc83fcdb5ba9a31763dfef8a7b266b66b661ba5814f965902a02267f96bc92e71283f44
ze5a624725f02325520f5511d04835789252a6b7be9f6069e1e5c53e4d4fc943d4068ed25978320
z06bca6a9bf9ed1331ac9ac9f5c90790b6382b94a747348beb288de95928418b6a80efbb73eac2d
zac91c7ba901357fbf394a67d32f34d43562bb3b6a6f0443a64d1e66cdaf6da852825ab30bc8022
za2ce48737ae4fa41a0b4c9fce7596964d205fd93b97b484bc5c7d7b563b99b088e0b312a07322f
z74381c44fd3a9d7a5d3105d4411feb6fbbcc3d3cd5d59c03861fd95fbae8aa6dcdb3f5b075d160
z054340ea49de6ca6874578541bdc235d90a88f1bf98e1477b2009ea4751bf495348747806d58bb
zc3a8a18122f999def93a8603c591bb6a801cf995a62294dd71e30b10efc3b4e218dee90f67582d
z4eb8d86e14183d2d77dad63476c381e2a3e9eb47f1ae1c35db57a1efebb2ac174116f93f9416c3
z8aeee2db5f0192f9476c5a0949f10ca7c616724048b8c89098739382e5ed31899bbd70860d3889
z57996eb5274d5cbeb00b4e5568028962bb0c9763c08568bc9fd9878f07ecd67a0c490a28d247e4
zed34ec4b531a3d70ea25edc2aa3cc87440ca59782d2413e355c6ae8db2f4ac3d5308cc435ca8b2
z6b386fb851b99453894581e98e1a7cfe6e2d08efd672a59c579dc70b1d2cb7bccd74cdeb22e71f
zc114cf8cd3ac6ee6534c3c342b2668bd101ded71b473e76b50b7aafa5b1ffe1552f8179228084a
z867b9ab690795d84fde1c48ffa54c4e2e40c53f10a7e251f3e335dc528906c6ebb26cfbbaa3d39
zff18d527b67c5f0ecdd52460c804c17cce7f59fff45d48db8994da7846585e1717b6aac7add613
zb3bc258de0f2dab6d32cb1413d88b1f74a86c6f7173f52608d207f4d11e343ef0fc87e709148bf
z9b95de10cb67036e9d1b1bc85772989ef54feaabd6ff6c7704c97b736900f18cb33e99648b6169
zd3963a35da8d7f630c21a085cb77335f990c91ecff1642e6fa4ab1175389ec42bbba3a39029a67
zac8b1f1219cd8b4b2b7233e836ce11e4f4970efb8de2ec348ed6856b8aa18ca65caa942d7b62fd
zdfe168db77051f6fa7fdf977880336e373ee16eed4d5f2e8de9b41ec34cdcc8c3d436499afb00b
z5e11b69258e1bb64cc0caaa68117b99fb707ba9fa6173532e9c09a889ea828daf5199102e22072
za6bccc28210b11064801204cdd27627ff41b77a3c4a165503d216d4e801c3237e2f98c72a2e3ca
zc3f8024480c80963c45adfefad2be59c7678effa50f980f3b4419ae79ee3dbf126682618011ced
z2dfcd03697a5a5a6b97426654484144c98068a835272281874c8314a5b5a2b4be532d28a400905
zcdf5bdb62710a1148781bdde662eca061591d7d5dc9aacbaa1e1328557e95c4a94de1ce1d6e09f
z5845110a45491d7de495a8a576bb8f144e714dc23e540f4a1e92d23750eecf0b305cf3a02bd1d7
z5b0093ae586ac4bd129d107b9f8f2c523ce6510c9194ef8fada1359679c1857dc56e1b0b955373
z540bae28ead0733c5e05de795247bcfb3a58e05ec05e866bd16eaf2ad9ee1b002306eabdaa5521
z3bb62465a65865eab0b23b306a24a6ccacbcb6c5f075b2e1d8fd9dd96f0c26d5879b6e1d8264c7
z1f76b87af3652fc94f71abed1c7dea69f2f922b9d8362283fdfeaf2421c250c1d8ba7d4de43d5a
zfa27ea763fa25ee1d17c1ad34cee341b4bf6b90e4010fb2f65a3fc786c85de58a19743a84076c3
z1be6e2febf7b6cfd0b0041461cf967b3a1ff35a9549ba8dd55836fd898aa7545acbbf376759839
zb91a179f649166ee16957c686c8f71a6ad510a8135f166000b456c5a74ffdc5dd848be1d19c1ef
z18a0277dab062e62c322f0f12eb646b2090d6b3dc199a27243723039818f87b3e2d3cfa6aeddfb
zf9deb7c72c259dff73c46266d0a4cc11b6d81d028f52ea516f184887b0ff2a2e74ff9585c23081
za705c6f0adca52519bf7a27f3042e187cac40cfdd6ebffd47db2a4e54e877ebb8c3c5d537f07ea
z0d5e684ed6cec54fa9284e089916d6c830547fb8f6207de437c6d23745ea593f1e355d6a855419
z26dda3285767695d44398851f30494bed806ea1edd31975d1e4c5fcf71df31c23c66e7d167298b
zb4bb9b9fae771f05023e7aaf9f527710e5681825d67798425a4a0ec7bfac869a96dbf3f1f8d0a3
z4688d3c5d4a0d3e9c97d9f134bf6c7407d667c71b09455c9bfb1ba797fc698222d47d6582ae4d5
z099e7935ba0040dc3076c8d41f833ae5e12cb3dea80b1f90b1f2ff9d63a19d85be884b7b9f22e5
z853c05d79f5a197bd3d5ef9d66bc1def5facae7225aa1cb24f9da031cb8918d320f60db5710366
z64e15f6771a85e369869a96b7b1ec4522534427adc9a4743155b0d29666f87838aaac530729969
zbf839ef165c3709224ad8932d755ac3bb9a4b60ed806df65a680b8edc6ad8b9675dcaab0580a55
zcb17b5afde72711ad03c2acd1cdf40c137934f1fab9e47af819f9a607bd7497a5472a4362135d6
zb29908a7ce70cd95cde1c7e8024434a7e4839fbafe0a6e612428e8f92b438ce5d90d2d1df4610b
z2059f9f78a7d37995192e979e753fbcee8910e3f7fb9d5c8396c38be1b04243146c561fc9123e1
ze7132683e19399fc20f9d867740d109f6ed4808876a0023c2916fec8b3a7a5a430ce44ff7e4d95
z680e8e888984754a60ef3d16c9fe0fda4ba6c5b23212431e01327f52afad9bc62685b41658a8d6
z02b777ceba099ba63f84d8c60087da81c31d25cce60abb1f96bfff6ae737dff470ee42dd525df5
z000109ba44405494e0aafebd9014f3f9c0a271092a0394b7425c0867a9cd18fa3a1c2323678c59
zc8a9fae6d0892be6464cdb127cad31ad75a66db020a35660929fbad24bdc9f8c969220ef1f4cc9
zeb395b2c8271872ee98ed169918b2f14f04cd53bd79d4980f31f5931557f7da509766a2b0018ca
z7d92b828dcd91dd25e3506e9468bcf81cceecc5b64caa6bce5be9e04d99f3bef120c9125f6a51a
z1a42da490017cbef64102079cd378a4b75b14c4910403bd8cc43154af2afc8a8703b1d1a10d29e
z0c4c05d0d9338e817e401ac459899479f0cab7da44c7f31044e648be75d29b9af45673104a0f6c
z175acf74aaed18d13626810a353bbe525a3c895a204f8ee3db926b2e550fcd980209d1c087f2a4
zcf8cb2381f7c1327c245e2f389710c90cd7f1a7e089047359295963b19780dc5c48532cc977623
z7fc6953f244dfdf92de3d1f8598240a214f5e2d23f614d0271681bbf9834984579357face148d2
zd573e4406ac791408f9ccdf4ba0ee59829b366d30225a4e9d67a71b7c8263e96792d64bf817495
z3e54b216dc2e86b8529dd5f08ed5bdb22e2752f19aca05d8bcc2553ef2847b7ee39b08336bf1a2
zfe16e3b4d4ea13992c50fcc47b8e4d5e316f2732bc954d46e01f9ba027172dfd06f44e87727617
z91d9cd32e7c7370524ef4417058ebde948a8108e3efa8d76af666c06d23f8f345ba3a10bae8fef
zd55d101951575850af349b27710bd498cb4af180f90435dac349e65085a4a734d24e24a26e32e4
zcd5d16037efdb9132397d5804b5ddc6dc1cd76549e32cdbe4b29d0a20e88bcca838667e8c74fad
z9f010a918535e4bb104e213dece1d597c5afde864abc2be96ed6b9639f33ab43a525bab4b95db3
z64bfe5b9914cb0c26c29fd23fb982017cee6a894c6d1f5694319ee3406fd0ddc9952e85a9f7683
zbaf2a8ef26809ae32339be4787df3377541d24c188e8683b71cae4e9608b8f2805ac35051037f5
z191588e2370add9d0b2bbe9b578238e6ee6a4e7339366f762b0825cdba5ba7f1c99df62d12e5dd
z178e0f22514eef73a6316792d87d9538aac334355d71677b126fcc6b125c60526ad26a3b1be699
z7bebbac92ab63441b473fff98f1a8089d250e4c0497317fa8ee4d215579f7822e34ff7e82fb856
z01347c3e5aa68c734db5afbd3abf51f379c74385b5d7a6118acbc845e5fcbeb69c03a17f7f32cd
z998c709532e74c8a6da988924fd3e8bf9e394731552479908fc2fb342c75ebaaab4fda9b37b74a
z7e345ab8e2b7238ff3d74fb27f5c28b5f832818d083f07ae08e2907d579ba1838266ce7775eec7
z717f4029f75e63a4fc77e965c4b530cb52d7cfcbd54c5a10452124f660f291b29fed1888306ea2
z7f3aab518fd84701a9d6cea6fc7a37fc5abfe45370a08b0048864942f025f4ca65104adc724e59
z1acd1766dbe11be08b6a72acd997e427dc5ab58a77b2ce36d08caa59ac27a6c8ef0058f35bc375
z43ff14a0ec5efe13c6082cafb67bacd00ea4dc75172ff9aca99a6e8e41acf6cff0640dea2b6657
z7c91935e00adf42c22c5491240e66301f39cfb973e8efc5bf3db2f15cb6bd87712d55f9e3165ba
ze8a96dd09cb5deb362967860b880a2bccfba9fc9889d7ee92f6b3d6b00c488caa07e54e9f8454a
z04a02640d07971bfac7a15c74196d7a51de718c8c1e6ea14558f3a4023adc37fdf3cca01d0ed8e
zd0c07fe073b51fe03bc759628c124fdda80f92c568d3090777419aa664c77ae4981de0c14882ab
z1f11a00023a174490d59cf7181be4874c933de66d0b7de0796d8f7a42e549437b6c6ca96b57d73
z332bbab4f33f9b46bc88100c8926f071a20a5e353d7be7aaf941f47ccbe3226037ea66881b6e47
z1dcd1cb1ee90436db7df0a33a5b748b6789099ad2268127c9fad1a22e7dec09b4b337e01012734
z5ef4d1c277ec54cd98cfa014824fb874a5d9ba1ea91572388610373066bcb29f9650d17bd21d16
zf2d9fee661c20a5a0850e60429ae965afad47110c7a1dd15f2da09cd4470525fc9c1fea41eab45
z574103033860b8239f69cccf34126c7637c010024bb72d0cd8c905a4b5d1501c8f8e4e2c17d6b8
z32ba2031f2764a065bd679db216bd43dbac84e5efb5536696c8ea7644869767c67c01c9fc99ac8
z7ab4ffcbfa318be79c333bda0a6e5a72f09bcf9dc8be2cf1095c47c029ddd92e2c7033a270a801
z1bee742e5196f8cca237ff5bf549028d0915e55a2ca552634372e6af285db76d0357f6d25a3ad3
z4d293b491d89c92eb3405bc0b0ad29ca729e053c706453e77443360bd1bab294a5f7c8b62958ae
zeb1d36f7ab9b79bca017f8172debedbb9020d909d2aa37877c5054ab00e1b2e41d0221f10157c1
z156e00cad3befeee8766f5f7056f37048a34ee87a75f5c97ae41b3711530c6cacf813e2d22b21c
z5bb04b13eef8d3c35db1a59e61b3167156fbe886ac316815406881b51fa3b28cfcb0959ba6715c
zf263bb787d893091f253332f3aa0de44e9ee85fcd623d687bd53b3e01b4ef2c3862410fdba837a
z82fbafeeea7cd56a491cd303acdbfabfea9d5029ca2316e9dd08c367b45105b69fc093a7d7a5c2
zd9cb3fb8ab4fa77dd000320803420dcf8a605b5d7e81452d3054d85149c0b0a682d008ecbce7a7
ze18b9f1b5138b5c440ca962c7e29141fadf9effcc8ee551c47a8e703b87a5f6704b9158cad2617
zd8b6973a3cd3d68002b657106292d52b4c5dc98b9936b7d5357b6d0fe257e8e9d1d2438d37cf00
z0c62baba4146b247f7b4328b33e23c13f16ffa8fa231c7c0eec5b34b14a8a47b3b39665c815c71
z20f224de14795097646f1a716c1cdc540af20903d91e16e3e83c2e7f3d87e5ff0b4730eae31968
z94f6712d8438dfd78b08e3a165bf6fbe1d3c6ac010681956231f48d95bf16805ed04ed0f3c45ff
z88cfc0cd15985540c855537b43e04dc778c7714a6fee849ee7254e95b84490af8025780bce3daa
z238b1202ee8cd4fa2e221b6b2151a00ac22da81b8649d9009d4fca151eb26ee46fe63efd901c07
z64ba10f84da2fd452ccc56a17c44c6d3b789ef61b208f140c73ab20a794bfc158064251b2375e1
zf0d6552e4e2fa5c5e6295d3b829cff5208f5a526bcc7aac73a94f4e243ccbb4ac8e7571d175bd0
z9548ba8b58c4757d76e29ea5725587e8f65c9ff151ebccd0cdaa5e9f1c17fc6cde71d9fbb33a22
z58be9f142286e925add1f220041be37a5ad7233dd5256aef5f9cf2f6caca52e7f3e5c33c97a7e2
z74d8ab3b5e4251eadcb533a8d80e1f71d2231ce5d6e43a08b770b5b7cd9a293e00000895786009
zfa03ecd00d0c248655adf69720d1041506ba5c3c746a7f585b2fda1a28b68b59d70e5b17631152
zd575de4eeb8405ce2ed13ab0464418fdbfd7054ae1ee4e0f1b88d4d71fd63f5966a992b52179cd
zfabd10fdd93cc29a3c096b7920f38a8bf89ee3943e76ec4e722bf8336ded305223823f4f891f4c
zbbda0ba9152027849b5edbd7c5efd9775a6dc07f561f58c5be2ce7a3088754455c16691d8fa0db
zb612e079b193622bbc6dc511e1b2c85a95b0c346a2c0dc3493c49a3a7bbdb4597ec92ea5f5d902
zc07d3d3e4292816eb1570aeb9c47f9ae8feb56f84f4ead5721e62585b8915a8e1d08798c12086a
zdb10f06ab720357c35389ec010842bc57a1f4755f9b9c923dc3b4fc7488509b16d62c4c86f2dcc
zb5dfa044293bb70f857fe6a7a74a11ea9235806756b9447043161b79849480a9d8c5383590e27e
zfa36b54df78a092efce4d49a08bd09ccfd61efe70db52ecaa366c94bcb8b2778be4e436ac068a4
z7b256e5df7df81ffa601b96daf353bcbacfc8a1b6abc2952ac7d4cd0956e4e2d638c5a8f085c59
z9b10b81566bf58a58479f5d54429ddbba93325c20028ebe5746b42e1cb1953888f36fa5f68ad6e
z8bb91334f85dcc27ee1c4c4d672b853803e9e81d6a254155e389015569ec2c8769ed712263aaeb
zf27f6a3f96a133995359c19c738d7266a2ec6621a2716422240ee44b024d70fc133d332be04f5d
z114ef763ecd30cfd3d194633c6f45dc5f70e749c432e03ccf234bdfde58ada803098f10a2299db
z5cc90dd0e14d732d21ec2b4777f1d38db7d0b7295df5d3b104f83ab3b092ea6d314409840ff144
z34056e6d664bc0963fe3e3592457d49461c86471e9cfd2f70ce666c7426cbca0f13b37accd1422
z683acb7b319e060bd606f9bf78513b5b344617f53bc81b7f233aed1cc32640375a38411d2f727d
z17489a1184d54279850fa9e72e74316394ce7d6a933dd2802a7912976927bdf7c3ca69340d5471
z476911e62e55108840231c76586a6305f7e52df010e0e0cf0e38f78382d6efa71d4b11c92bb289
z2cc174e5594f6e7549be3436b7a661c5af2bc335485ac8341871475623a58c00860bc46a6d1c2f
zbb90f872d43599ee07f0285cfa79911df458e5549df2619576bd4939e35d1be1ba0f012c4467a2
ze944444b0aa8d3a73a5d44cdb64161e3505de72ccf1aa45b1e55fa37754ca451393af3908bdf8e
z7338e8626cf4d16632345b9e6164ecbe55c0375410f750d5cd4540aa8694841f7b02a2d238c5d8
z3f5c9d9a40994feeef997470577b79b4f27891986b5e5eff905b55c7f5db9d1064d95fc915731e
z26580dc1ec3dc056b483ee2b2d28d1c3c8b444e90e8afe7108bc3bb8056d6a7195f2c8f37cef45
z90f25b1be8db0511b0e2f85b96511e806555e55b36c90af885d5ab54794199c5cb73738da5db7f
z3b7362d7853da14d760c93a1063077662f6a8e45752dfb00a5268c87a7f66603b2fe437001e78d
zca4968551c3c574dd30662385856b1b225bb8788c848e64694df2f73ec245818e10308abe5157e
zb243734e0ce4214288904d64cf35f55e85a1113320a504cae084bdb4e8ce12987da39443ff3fef
z7f810f1c466a94df052f7905373f957d3da706743cb9283c312e362e4d5a5382de0f4a46f3a46d
z8dd2e763021db8343bc806fbd45fb657022453bc8845c30eec1b200c87917efd070be9605b30a9
z4a247f31cb6af871a25cbd53ea35542f1a18cddb7bb2d79112e914dae89aaad573db943d4bcb88
z56affadc42f6407e7fbdb0eecdd0370143d24eb59560540452779a330811f16ac43b12b15b6782
z89f8cb69b7c2ae3d57d10fd99dfb74b3b3561817266fc67baeb1a33f15a9d6fc986b7c057bd525
z0653d6b37c566f3efc2ce33bbef3eebacae769ae5f5db2dacb424abd24d2668333d1c9f46b991b
zacd8d58fce5ca1324b0a8da3559a6f7f59175a69e2b14beb67df785a93338a677c9fef6c68a7d6
z67ff43602323f2f7f0d61c35a9d4d979df41bc78593574ae7e89f8c092c03e42980f803da8db9c
ze3dc046e68a21eadca6c4df4b6fd0be7a9fda966fe35f56ff70591d97eee8d2ead4706ffd62344
z5a7923fbbfa74d2d685a47870dfd693aa8f3a40b34fc26ee9c12a3f938b91f429e679062aa4569
za6b32a39590f015748ff6cb22a4ba8804c1341decf45e6555fb4032297aca0fd95e1f5f0a4e495
za938e26f2b8a2823c24a01b7531a6ffdb9d4c1e65b7a3a1dfb383343adfb908ff69739ec87fd30
zad6b064097d48ce0408180ddda35f863181ffbd897967e045aa9ebc8723bf66501d1f9d88355bf
z3fd8142751b17b66447f0fef4d1a4cd6e16a5547f10bf0dcc51e6aadf1456b22694141db0fcc30
z860e8873dbea99cc98ea3bf37d2bec36c5dd72b8b6a6d9bf3607c6bd0dcc24ea3638ff86b08e91
z8467b5fe74495b988a0f228ab869b6b20316df435d9565d76ee1065f9b5f36e85e87ee9d9f9584
z6d09d724a6d80bb11b698c962bd97903c96a57f07ed08395bddae2690c256b4a48988e26e21475
z318ef5e0d45194902488fc91211aabcb2b1e951d31485b2c4e2ac4be1a3a9cb2190e9abec090c5
zce6c29d9580613e93f8d7edb71baee3ae0ce77b90eb1237fe2161480444efb85625b9610927eb8
z9d3ce1542852c42a3356d075d65024a0473c7e2f8b788ddd5b8fdbf140e0d5913f3de7f108a410
za10f8654a82015e73c04bb09ac7035356eb93d06b829e595f7570c6407b6c35f84d66ab9057fd3
zb8f176479048de54712c66835d382839f10fd4fd0ee316e0f7d61af29f5f9f7a4dc57dd262d15b
z59c55faf4bb30c22d8b00710946e3c4e5196f57df61701b4ddf2959af86e47898e70fa993cf484
z5365c4eadeff92dc7d4d785d0f4967b92b613d9379385fc9ed2a7dac1c4ecd550cfc539602c2b4
zb03767e93caf4f6db0251819c17b8b77afbd88bc5857a39ce99b23aeb72f20245d56417c29550d
z161cb1158cbc9815b208ead501960da0648a8d9e7a30b83783d2b2974250d13edd9827cc8be031
z86fc91de0fca81efb4f6bf863077d462fbdec0400a52b6dce9c9e3e98afbc17bb225185f482009
z98c62f8ecbc0668556f97c7fb33f6759e2e1e7a8c8e10ae362d074bd35be363cfaaf81e9b57d95
z26ee07c300103f658a1fee2d7435da1e54d10ef5be1dcbd903c1edcc980f69972562b596a21f26
ze394ba3f13c6ddda852c7e75ed85e36669f729ea94c31a34db9dc15697e18c3c07c95fbc7fa9c0
z3d35a69474d682205686389d7b79ea8a39bb630590b59bf232e869c67718a1133bdfd66761caa8
z24d0d844fa52e80725eca9f4932e3420fd5abf94d40a53e5a9055cf1630134f30a8671e9eecc6c
zb87ccc291fafe873c1d37c4211672b6f44a17b7da9567e23be275aa7965b3dae8504183c22c20d
z77bdfd0456f4fb1d05191f007f82f94962fa664638f17a707fe92e08517b73cbcfb2c55e07194f
z2ebec4eaacbf55a6124498c3161833ff4268d9fd30e51175a3cf9de4c6e323c8404b3f0dfa9700
z421df22a88a98824a48f648d7e4382461ea08056174e11384e42f7b364bef7d75ac04402a15449
z7f9a5c2b2499945b87d77bc879de25cbcda548d92e1d438279045256828746f02fd3bbf0db33a3
z908b899c8b3be558fa6919e92b5f7b5d948ac5e6645e207319061aebc56368e6d76d2989978b46
za3597714108aeb74b2ccf3e5cbf10b08009a94bbb64a2aa5b436c7c6d27dcacbc5cc18e67f12b2
z641eb18d179a641c2c7085a1ec33838aa534c583122257f4d110497ce8e40785be261335982c62
zfede53a166ade71ef3c2551a7c8e5b70fd54b4b52f77e92a944af9751fdd667de6ffa812dc03c1
z1747b5cb33357a283f92d663b1cf14f458d0d37a56e9a83ba736371031837aaa087c8aaa0c2925
zb48c37a8605785a29332909d5b5eaa8a783568720e38177b4417675129d37980de5ce1073362a6
z6f78e8d4a7f00c6ea824dd0832c82ababa0224ef7d3376873f488d395ff8796b026ddfd0e6d1cf
z1ca069ec53c3e6c00f989f1679fe7e6dae1982e0e31d3321b392a3f8d893da9a769568e056e48a
z277633bce40eaa30a8e1a93f15bfeaefff5ca8dc56dea5f15de86f6a8aa684942f97e03476aafd
zb26282c5186b49c8aa7e6d054e7dbc40d40da3ecb14beeb2aeeff9b74283636af0ded84360367b
z77e998e20e4ff4275e7dc97a14845c857a39035479a6a257682e0598535fb65443727da14e4b5b
z5799a7d11085e6dfaa66a96d5dc257010b2045637a369e8f9fb6faca93a59865c33103b74d5c57
z16bdc82bb581b265334785e37081fab6404f7ab52f6ae2713d64323bfa02e1a4fcc07d8e7c7ea7
z7ce642f2669b67fb21d0713e57271ee72c819f420ef808993845ffe4fd9c582a14acbc34aa9f03
z86e9fe7e40a484495268b8e2bd5f71c9bf24742b0dc9b47e15acc034ca63c471c67721f9bac954
za8647139abf71c2563a7cf07351d58f99974c2554a9d97c991159107881e36515e1a13b58fbcde
z46f1e2decf51e4e15f361d13e4723b8f9931b0d7b8d7be334bf042b7bd75422d6e4972eb2129f1
z6d45ca01ad9d49081d3434e92280af6c4b07d5f8dd10006c54ba33a203c8f045f947a4e532027c
z6a0267361056715791958d443d01d5f614895b5aee06d95ea5f1a5fe55ebcf4df824ea6bdee796
z5d4534d0b4384fb9142e66d60f9853eb039ea5baa2d466fa78aaa9e495857a0dd9e550f128c969
z40e8c32b3861479230596933197100e4051e26503bf88689439c2a1b8ed64b7e89b7628c6723ff
zd92fa3bb7d3ac958e38a68919de9ad10fb42ec68de30db755444fec2d6e84da0244fc10b574ca6
za04d5b8126f62212e84dd900a43cfd7bd85a955de46e7c3cfd81c5aab3aa57d66ddb39fdd2b39e
z086ea331c5b5e01f264b7dbeb1edf60caaf41cd87df3aa093857c8bdc5d5fb080a48329343e5ea
z9b51086ba6af1e83c9a167f9469847d549eae422a5ab476a5b7eddeabea3f2143349aa1184a55d
zce2e791cd4f7a74248894b19b3c8f5faaa70575c4e676df2b3628ca13b91794f96f1a142490e21
z5a996598f841210f683a9a5d68135b43c49e7ec70dd5c78cc270b5699ca3a93222948097608bf2
z2f8a9f7c43cf90b0caad3284af2b4d27a478ab2c34c34b23ee2d40af5fd972be90db370ea1684e
z774074c5f7818cab36c27a48fe11bedccd9af90c44451f5d3af5e9e3d9d05279f210e6cace63b1
za25afa79c6115b7926f079e8f85dc89d26f89e32ee084b2bf231073911645c88e3f9775a5c579b
zd7060e9ec05e3f0640e91ac2384fd7ead7e8dc858ecff00b6506db2883185e67a791367bdc7327
z1a0cf951fa8319a7cb9c4e19600634007a3163d067ae11a422d0c98156c5e7dc37cb6e6f65bbfa
z123a2724213134fe7a62e951fde6f1700ac118f988d95d382472316d449c07a3f83b0da411ca3d
z88637cab18f1f180f0379e569a8024be12236a7a88f1b9c82f6c400d109d9e8af785bfb4520363
za1e10cc66e8dabe52458abc0cad0e5d1ba88bc2794ba0d521e7ae99b665cf1f89638d5e54c4dbd
zd66de8b20f9e9ee49af00a16ec61b9373dc99464504fb31e22ff13ff8cb086e669d5b7a2f58850
z638e60b782e7b40d2b3f53fc71c5f4b0812470d5551fe898e2c0387dd1f422a83b792baec661eb
z0939a0740667549b892e4494c32a970a695e0b45bc73171b7686c5049cb16fa6a3c07df6728f95
z78bbc01707cf441d602f25c9a8d176c65f094ac4855d7de124522715ccd07de2e12e99d2d1c8bc
z5699af38070f900f69405e809a3ca677a422afdf1f90382ea839a7a7909cccb12658ccfb49a434
z60f8f87b64218bd68f9c6a7b97238da06a69902ebb1d78d39a13a78755c8c9a9bfa3536a69926f
z16732692febc16d504b3badb449d78a2fb30d2d47acc75d84411894af597e07daddf3c63865cef
z117942218d312fa375c6e0be373567808dcc89204cca29a57f01a5fa4f591c578ba129e3b94b45
zd68468c0d8b365a94b9f8d1b04cd875cb7937ca515b0ec9d857ad98303cd1cb28301c03bc2e740
z230d7f25b52fdd5c6ddc87c22e467d9f0ad1bc30172cf4a0907f587bc9c0aa41eb5e9597377c42
z031e49da2994acb5c2908cc0131bfbe547d2702eb830a0f77366c84e944b43c5a269429f90de42
z5be666e29a88149c0fffbfd8bea0cd6dd7c6a564d2b5711fc11e36036dcbda1e9018571903b7f6
z1a6995c00361cc58a50e4e421324c41e4aeab284d05d4d5bb639192122543126a4e9e27f3e7361
zbde76e352316f6e2c39bf5de39742369c5adee682615039ac8b2285693c7c580449244b4478b30
z8cf304e560da6d015ade731354787f1cdf540c3b76daabf7f7eb2ec44ac70423e88fddd1e270d3
zfc3a8b7bdb3f201e72d2a6c9fb16f21851c0c8711417c69a7729b81f73fca81672827922fc4bc5
zf63575a88ddbd6395081db2a97cb152f0541f7b4d1236f16f28b9295870b3b910159601dadbf39
zcedde4cfa96b193b26017e116a8cf7cefa6b0f510a6d6b636c8ad2d821775ba10495ae82834464
z4d3f9e0a32da9b140f49adc0a4b8bc6d1ca21fadac1efff4acc6c39f816c231e8e01dcf0bef66f
z74fca112cc5d9f9192884d1eb7fbf7692c6ccd219e858c41bfcda1580f76cd9cbaa3945176a33b
zdde78aa392981c45e8fd8b07d79bdb207f6c00c08e820e851b6149957c8cf16b5646e2317072f9
zd20417f2cfd390b97ad4ffb5614c5e6c86068301be7028576b88c1425a125d30f63482dffcf8b5
z5af211e3f0a291ba1a08d48a071d1448030468d8b0ed8e5b15a834dd38577d03c76390a36db997
z0cab0067e5a0b048eee1e132304b4d12903fa7454308614735df43e7fc895399db4c68fcb5c88f
z286088bfec74532c8867b6f14a477991247708bc8e141bf92942017e0861834090c6f0d9030212
zb6a299c89998d2764c356f0cd2a82d583f14f46414f9f8f7c3ccf904bb5f2472dfa3e8b3a48efb
z5e146f56d5c443820da8dea7afab1dfc2f36e09aa95bfa4c9752035abee250d0e4217cad74d6a9
z584f4700a79b46933c9be35d05412bd4c82126446f9e3f49c34b38fff4dd4ef5484670607f2f89
z4a0199e8e74aa11d6099b4598fb0a11a9d75b25ad4097e56c81d167ce85d811cb46927685444b8
z42c45eef2a5c6311a78de51698ff339c37ad593e15091c857ebb0e796c7c5a63c9184d977bb6f6
z17202f22ad4354fb5b686646d3c8137ca69cf0d28e46e9cc92e73ad83f3bebfc44b76bd629f901
zb7441a1f61be3594b0b08dc24ce7d20e2359e533317cdbf86e7782c8009ce72bbd95e3e558ba91
zb415f9ccf2aff29280b1f1ae29bd36f16ef13a7b655738e0259053519a27a73f89f751759c8b4f
z5067f4d841ef222e7c7cbfc861204cdba08efbc14952cc05ce800f41d09aaffe62f022194d44af
z7f5d75cc47aae2d2abd69a6478d6500ab805b5be49b6b2f46d0e6f2eb38c40b56aee593bf38c81
z519bd352de21d44fcff2b4f4617331858f11027bd6cf9ad3f705a276acedb093e6143ed0f5d921
zf58f7ad7bf986861936b411f7d5faac3902825d586bced09a2ed914c8f1265bdae06624f68e12e
z6b1c30344a6a78871943f35b33c14cf2fd4ab54bbbc264322318ec2cc5a13070b6a2e65f8eea59
z033b1c45c9d6c9dbbe9a4acb812c4a3ded2286ea910c0e886e6a7fbd5a3f6247d746a7ae9c2ea8
z568b39b4ec07a9ce0a99d4bd4de83628a1a86508d9a1e236106691138e46285db278c1c3804148
z642cfcfe0c1ba64bba070143fb59dc3e6c681b911fcf7b3b632cf22eec6f81c7d299170e7e16f0
z5c8aeaa55e492152a2a359f194b603096d4f0809c81bd1e2be53d1a23fdec666927cb027aac881
zdc32b291b36f5a999fdf3a536e573b5b0baee1e3b8e52cf5ec357df5e532ec5b122e80a96f301b
z3ae6d71ab0b3f8b4b24f532b6e95d70f41cd24dfb1571179cdf77c78124c40a24bee176b619165
za5cc46dfd798cdde497bb97155624a47e7bc99effe4276d2441dfefe6779100c4c66209838021c
zed5678ab8728e90e0d41ab97ab974b208ec01e0fe5008e2245b31d1f7fa05d1d00efb7336b7c4f
z21ffea0a5a1abdda9034858b79eacc158d2ae52b18aadbb52e878cb322b399c04036af67b23533
z2393ded4e6ed7e3c42f557543820e89e9c85163d3e56f7a223f984738b620de0ee3034e555f5db
z1b3b60c29f5382f473f8b769ba3da6f9c6eb989d0a0674c317859cec066cc8b56c9f4128733aff
zf50830c81c815bc6c629cc7f27ed0ae0661f7a7a7ec4b54959caf35c0f1754e9d84abd4d2b9490
z6281e2dcfa28e59e6b6f976e91468fb2cb8a3b6b7602e40e1a4da4d3fa9f2151a4c4d4fc24ef36
zbb717317c14900353f3ba544c5bd683bbbc9ad54560d9132843465073f6b2c43088ee94f388118
zef48bbf733737e57bc19774382fafbe92e00101ed9a9fa90036d5edc0e71a89c2b0cd254d25698
z9b4069716404059619efde709f5dc8393e3d6d42aa53167ed94ff40a5c49c5cafdc6d667da3dfe
z9cfaff6c0adb4c223709e070d6a6445fbaf96c3ca28d86df780b2bb82a9de2ead93a33b0cc2f2d
z2dd169bb7861044b74b4024ad7057899e65bc71728211793c76b4f7697340da4f956e2eeacb871
zceb3b8fb4d32dc5f873fced70125de9211b0bdbbd0cd3adbb4f5a3bd5f9981c4930171522fc1da
zf06652ec7f0d80c956f7c2740d1ea6bafb6f74f08b5a13586cc7bae1f2b645936de7be720aca05
zeb521304994a6ff68e5807326298c0f529ede5646433412a040031d6c7cd24f5eb52a648181c73
z5fc0a377d5daef01cce04cc08e1e0150125c7158468b7cf0b220a77dd0f147ecd662e4db5537ef
z55b7141611b4a3bbbc5eb8cf58c8e0223f755924dc3aabe454bcc5b04ae3ebae9f59b5bbe4af36
zcdf0820b613764ebe4442eed458bba0b29f63a828dcdab00fb629661e3250c9f972cdbf4fe1526
z67709cb5fbdd8207eca9e062b2fdb9ee934b876aebabc32228cda4908860db8aa3adb742b84ae4
zd278406c27d85534b5fc454242845f6ed1255c6613f97f6726afc333760777c4555f7ffce84b00
zd5405f8bd3c42258f8f9495af656c59a571be6ff83bc20a4260a141e1b7f7b1d03cb4728205bf5
z98c61aa08647d4ad6d933b0d8c09bdb6dae9b5fd5e9df9e069cafa278fabb83e612ba8590b4fe8
z1fe1cdc8d92b213f43588f75999ad57b6161efc7a539807a2dc7c634be46487c181fd8262199ae
z650e321c12b7a7b04695429c946d6dea5a7ee2a5416afa0146afae9a12ac0f4fe251cfe3fdf870
z54b54876f589b5961fc972866153d21a366699e4e774e3b1b901772ea0561d4a533ac32322f770
z44685a5a977af6ad71fa97b18783c3c735507a37c91fbf5a148352e282dea59f780f571fa79e7a
za2b7acf3c1b1048a2ce534269bdc8a9b900268b5da51b98ba668768f2b2318ea703018cbf4a1a8
z6d2a7f792e3e31e143d2cffbd934332f81872e3ba6ac298c7b5e5bf8e6c92b64a44bfa26d07350
z33b000ac55312ae3c408a37a461806bc62c28401051e528ed5c5ccf023c26ecb5e6083bdcdbf00
z18205622815df71985b769532a0ba7ab0443d93e10a17bd7ff1a27d68c95ab740f9a4065e88691
zc76fd5d8f410e7aab1352f8bc1a001cdfead6b6d8afa654bf2dfa4bf3624976fd8b17364d807ec
z49673d929d99247e0af9856f72958856e0b84462d6d266904b373cc71c98dcb893d1f8d315167c
z0bf60a85f221f7fb7c0ccebfb85aa7595ae265fd3f8dd867c749bf47aa0fb6844671be0bca6175
z61db9659a6d31fe69d85f65fc048b7b09058dfa181a262d0d2a6ef733017badf0c0e42d528aca2
zf9460468e11b04c3b5d42e7b246dc2bd12c4c853fc1569c344d89af952623ec89584808e1fe99a
ze869a00c71a20ca7e7315885b940c63be705b4fbfa94c6ffbd9fc8962ee48b752979028766c6f5
z3a6bacc54353d9e14985dbaf08c3988b9775fde3687a80502a70b5b003feda0730a3b6d41693aa
za2170ecc249d1e2eb423a1da9bf44db31b7800987a9c826457e45a451916eb8119d568cda604d7
z968477fd51a98f0463f02a7031aeef56cefc4272acaea7bb02e9483a96b27c42415aaf5d238ae4
zaf93afbcd942d58be4cd467b08e02010cc6bfa94befa444704a7a6b45bb58a3a90a3e30f128a30
zfecbc919042bc387b1de4af5cab3d176d337375b75a5b05a29a07c8b866860326afce4f4f67885
zed865a16d9e31e04e0af53a980e571e9602e43e94ff42d0e1f3ed211871696f5b710229264eb89
z726232d21a52812531f80cd9e749b30e061400b5d734b9b878788b25ca8498e6823f23258c3920
z08c996b4e3e734312875e462d30a4996ea1d1cbb63bbf9fb924a5ed233ecae00e0080a2e25a931
zde880d32d1b1d860477287e1f9dc32f38fa4c158bd46ca3c98672c580eb0c0cac86cd569792132
z0f26967ddb575ea7252b54a9d51a0d024b06fc543f6f1e040fc84bffbb0d78c8f98fbebb7450bf
zd042daf67d675b55d19362d16150da3f19ba2fc7f09cbd7d54dc1a10a62bab9ea068b59d0dedb2
z394becf852aa04ae6842ca2579b18ac55575b330db9bb32a9ead2f26e1c8718467e0e0496a6d8b
z43e3ee537c7be5cbe0a6b7766b378d8891bf3c9bd1d0b9d6dd5737bc6d8667944176a8db83368c
z553c35e789c4c4e5d7ff6a1700576ccdd68bce0188d1f26ba3eb59c08e827c9c9e20228480e32d
z044eef9290751127fdd09fd8954ca833e892992bbbdd7364f26a4a1df85aaeaea8bc8b6746de92
z42313a749e0cc971e11a8ff55c110f6c1023e36bd35c4bbf54d11c86ae8548a31b3ca8f26a26c9
z950230b19e1949686b946a2c41b3c685bda13ea96c1336e1130a54e6ad05e1d02917916cf8adc3
z7292648bfb007cfbd63d8ba7f03da0cdf29b96587008f6c74c15d281dbb46b07f7ef361061afbb
z1431554a99941e81ef061a45068177afb9127d84cc06d1d0d87656edab660885bd057629f7d9fc
z20178bb9179a43ef8c87643799704e0f3ac9584c35ff732cc5c3d606edffc683ab5a6c5d10d44a
z11e67bbab1f906a58a0775451c9bb2749c902aa4fed693ce7a667f22a77c17d2b16e0bbfa94690
z3e9db62b0a6247915fe4eda8fc7ebc542792c5845ad937118557686078c51bf2f32980d1eb2496
z9ec1a2175004e2be10036893c92ec76b6cb335e736ddd87ce482791872e4732edf1cb93fc74a45
zfba56ce286e00c3645be3fba6a3d9db198e8bd2bbad9edb2477603a4e27166ed98ff877340a098
z8f3f409b32750af73b07716a6757457c626175ade93722bfde852482b27f5be36113c9f92260dd
z64c26bbda6e4f5a5082cf9926951027d13d213a4d166fa7bf0c7c6b74040ebee1d015ff5ba0213
z4121df5c7edd7787394d078a318477a68479581cfabab34a4b0d56f5872372e9a737b1343ebcaf
z82ece7a4418ac34858e0c64cc11492f384406e80f1718a0042227fc14322e965ae713ee2e3e7ff
z1e7cda429faa1ada7fb44f7e698a857283bda48f7e144c10f3ea1ebe3b3faf9d3fe1ab81af83b1
z04dc049ca6af202ee074013cb00c14cbc4b36a892578812791c7701016f842462e35523b07ff65
z20d87890e1ead7cf89c7160da8a2ffaa480b585c4ffbfd4e12e9ce80a92192e869bab412ee67ab
z9b2918993c4534f6f001bb994e41b8cf25ec9e98173a568cfec457d53905df2850c960f04aa3cd
z02a4f82a33b627ee6753f1f5b510413d28b973480061342b779d18c51e84da9d4a06ea7a834f4a
z65d60cc42e54c350abb0a4a81607795f7305753fda29cbe5cfdd200e2b26a49068878a5c1003fa
zffe928935d6becf11b5e03912e14a5df6ede4a51ea37ad6e326f8ca760798f3bb0879a4a3914e4
z6e525b7bd09598d0fb6492ec09f5f907fe95204b81633e331e7295712f6547f8779f79e7e5a1bd
zdd5f7bd0e999bc50cd28e24ea2d7856856c32adcfe925710df442bfc310bfa1702b31b99390e2c
z78c1de00775cf435e093fcf6e3a1f27bc7ee399f4a2df0ef7c9e18866a9269e04821a791941d62
zba2e698988fd827bffe88032ba59b4bb1a4b26f9d223f671497bc8c637c698beec435f036c2c51
za90034c38f343bd42de4ee5e4f0216107f1454eb1e8fa8987048e6fb1233e1337879d2ebb1806d
z14f81b4e6f223b143703f26b80087db1bfdab4243c60538957f1298055716f37d084b6ce5e324f
z8744eba006be9f85135d92abc2c09d4c06cfc580bcc85e1a363d5d0a3bf64497ed385f186f79df
z1067a5439bc1b7692b4aaa389a75cd271dde7c6e91e8c23fcdad198914c5b48074281826ca6f54
zd6257f82f36be51b5ea5c93ccb334472e88f8fec8ba595c911d2d9f4a7e70539ac00d79edf83d4
ze2d8359faec0f31a5bdfa36f69484dbbc8ab8c36e6f0864f3cf45f0dab7a7e16fd4cf51994afcf
z4a988e6874eb9e0fac659fcec3c620f333d9cdf22116a8687bd4cc88171b678315c681519d9f8d
z48c32d9ea7bff2c4da9547c37ac2b5fee97a87ab3718a331ce717a27cdefe3baba6119cd70f45d
z19b66e02c348b6f582b087baec014db2030692da25019e44b8b75fc09d675b217c117daea287cc
z1a568de7fd4457134ba791ff0c9f8c830741792ff7f6c39174497ee6aaedc1b2cc2a2c4ae53973
zfcabdc2209013c6acd97db1f8f44a4739f0b12fe8414dfec21c2c081ca6b361d76874aa025577d
z874159895f65e3b2c9e762904911702849309e8b498c4137305a44a53ab58a9379519c6d638063
zcc8eba1d41a827c834b4107f3d1010e8f4dc221ca17a2fcf12d08e55f7585d175c0dd7694000fe
z655eed279d752434e5306415a791aac70c0d3b5ba4526f7189ebc53ef82fd56b4f398292a0b582
zae6373ac1790c5e36029915ea0506b2252a665f00a491ccf14c713409ab25e8a5c457552a2d3fa
ze0d3d852a794d0bf2a4b164c66cbce17b2102fa71a1ab076887033737694d5e652d4f32a691596
z3f2d82d777dc99f0d218ce71df5acbc26dffb30ac7beb0a22270568c5f233d989f075776aa5048
za6adbe0cf14c3bd9093156acab1e8702a2667b4287f509517c9e2a18f3da5604d0f4d5e6ff4789
z0dc796952473bace6e2024c336e05aaad587983cc26d620fc4cb2fc9af757c96de90b75d0923c8
z88c0764912c9670965f2b89fe619c2486d27d37f216995a76bca44d498476871e237034d04ecb8
z841e519e8f444531f5bacbeb3e20f0a5e6abd81a5182a2c86fc31ac4b77d2d6d873ed852796420
z6fcabafc36cedf16b8a896cd378cb621b68f71f49b81125af5125be53bfd1b0f8611b1a99d7241
z249630eb8869dc23ca512172596dcde1076c260c704302351ac92b0639d9e3471626514cb866c2
zfd3c97fa99fe183c3c9f19d11807fd12c8fc991ca848480a325d0d3ac6a4888db85b2f016299a4
z1f1773b6b50913ef63aa761d225124e15fac94a25d8397233004cd7b3f736a9d4ce9ce337e4526
ze7d75cdae70b27fcb6ca730cbbc09c21543b0579d7cdbfdaac674985b6a09b569ba4752622e3ad
z292148cbeb7b4e2761f44292cc3fce77c92bfda59e0f04a3b551db6a2a49cb2b4b8d9e81a7ce93
zc3cbec95b624f603e5a218bdf9a180768608795c2d908a66ae07bd9ade003b5e79d30fc3f2dea4
zdf644abf60d6d476b6d568eaa9acad9497836cd9757147baa999616925229db029784a3ec5fc42
z48eeb4c53c68b90cc8fc49244ed37afe5ec4f1b1d87d6255552707832f906146446cb3e8808abf
zd062b2dd1981590a0f5b579ba9efeca145c7a765ec45fc6ca82e313b6a0418d95a9f9ead597713
zc7ff87f878d25cbc26beec5ebdca344df989c6f1b9db4c9af88ec1666b1fccfbaf9db6fba65fcc
za245e1410e75614ae0894f432ac953a3dbf403e424f174793ec80e4bccfe64612f251eb905eee7
zba8eb1bfd828ec10d4256dc0d196d1cbe0917735acfeddb5c607ca50770518a6ad282e4d13f8cc
z974455edde77d2edf4c23f71f0f430a8f345dd0ddf258a5b147a3f4422c281870e0d9e1770119c
z0687de493510db3dfa5be8b9bca2bedcac378d9d5da28498bb76279bef290a366a57d0087594f8
z8a29571577c7e9770de53c964853363569b287f759b21bf9dac3ebddebb57b10878a392d0fe56e
z801e60ec9f50a97c66ea1ad729a294f929c3bb723ae3a15ffaee11cb2003891a27cae4a87657d0
z263309fa8401d155d447e36937ef8f5dbaff7cebc49711249edc5386bc515461f48b655de7b5af
z64501dd115c2b69b274979eec030bcd33b44571015361df4cc22ce32096a1286bfa5f622f168be
z1b31b65513d1138cdb22b257b5b3cee05b371505d83a7f7cbfd11cfcb36d5d16d9f7cb3bbaae5d
z5681ea1cf8a9869059e0780d26ccbbbf3e02c2b36acda04c8c6e7cea34de7e5e4b3a387495e2bc
z6b73dc44bf795c0bdcff5835d80ed1cdec23196ceaf1d38f3a8bbc94d3d5b131b26b5b4ccf0d1e
za649031a080cca346b1adf9712d99cab1e747616b3ff00ca8b1d405b5c927db9a36b3e3a579fe3
zc3379ea12a980149b2587b6606a7bd8f3dccaa556e1f981d2719160ee4830f3209756ec9957a6b
z27d9b93c18759b0ce6d132dd716378939a472c85b392b7d416cc93a00dfcf1acceacbde2770662
zefe65650989847e449f598858e17e07e52f7a2dad20bdba40e07bd34b78686f401b1c92d3b44b3
z41d01d854d3f67b229175bf7a1c047459fb4ce1ace8c5b1f11da29d049fc8bcdddcc8e4aba470a
z946199f966b397079508bdb46cb1f03d97f8afd044b810399a8cb5951f801981ceaa00fcd13fe3
zecabbda1d948d2d93859e247ef55e5113f179d0481129a899615c4ae9ed5b8b1d7d28be515c343
z8322a8cc3d5f9e9d15aec4c98f9a8d1a47867e7fe96ef9735cc920ea6822fdad952d16351a2c19
z5589cd3714c93835e97cce795c1d049234a926439f928abfe24b5d9369c5349f8914bf3056c6e6
zafb2ad44a009f24b6466341c3b316f8769201a51dfd559d8c0e7e6772acab5ae854f543eb45ac1
z53e4e8dbbfe7b8c60e4f2950d26b0bc3d6c0ef7587acf6696853ddcc99745cd1439ec7f9db7c85
z8bf14f2a17a2f88ff097b25984ef2dbf041a65c913c34145b5ec28761710b7484f9326e9200e76
zb41ead13d25919e851a7935d064a92d13c718098f1104f4749f344413c8d50edf549303c561e2c
z6fe1ff3d83be93474b2ef9a1309994692da709183cd7f6242b47f863903aa33c9d6cfeebaa19f0
z5a0d8b5fa12d19fc25a64ad3172ed3600a73b03f2cbe3dfd50d670f8074e521ba929978132b8ef
zf2963c783ffb3ad5876e6c41a46a5dbf450a3395f9aebf68ee1200c50bfd537fda292386416638
z511995b53aa4e06b4a6291712cc91be7f0dd16d7488fcae6676587fab4637a03dfccae56b97553
zde625c1366fc50636b1465a4e3b80885beb24c23846b61801c97da03228e39d19f4572e5b3d747
ze08c8b2625a3575efa8278208e1d8eac85235c552b433a3f5f4ee1f88c3e09b5f95be436d402dc
z50a037741c62579661f79d94324c17ff8c791eea0aa94afbbc84c584f5182dc324ad26c5bc84e5
zc84d91dafbcc331c88d02c84f396dcddd951eb58af3aa8091056e4b95dfb1f9a16f3bc87ba0863
z3205ca84043e32a92ccecd4bf88a6e1a7ecdacfca7d445069aeaeae9dc7ef4bcdd73acd0ff2dd1
za57cd3ad1dc8c7d5aabd88405180d5fdfdb2efa1e20599e11dcf78970344a54c0a8908089110e9
zcad0c1baa0c3a7b26a2c8c39bdce59810de20d9c037b98434ec86cc0c8ec40939d71fc59ee76f0
zb6198aa6c0ea2b9e197544bb187c8bcbcb88acba1ad2cf26f1c83b5715a29ec17233997bb09598
zb800ff996bf2d3a9a83e47c79de10ba26be2c88a7cc75d4d4decaccb018fb0425eea662ac399c2
z2786b99715b88dea6ef4c221ef97372d980a6e3d131b9925664ca06f88c3ee550378e5094b2e91
z00e830ed003dc4f3f87b31b11a7f3381c279c0f8ed5fb6d789372bfc64db85dc7d649e0b7e23fb
zd2db7ee4a8798f7421d15bdb3c03962b95c8a763c8fb83073a49af535cae3ee960cd3fe9dfc1f5
z011a5b56aad58ac8f604939ba07a60bc6b10718f17e1a5fdc825b1790f61483a507fc0bb84c8f2
ze6c230b6b77b52d04ff61ea09c4125fb5f41620599e71309d0d270c50e60d1c539ce6105117caa
z65c68384c0539bcca9588a055f1b6e40cd9de8eb220438b5a5f380f09e350a10ea5357a86b8250
za426b7dafd84bf77d96187cc34d47796e2d5d72db84f66f21b4e8898e07695103f3195c0b6a7b5
zdaa01566f4dac5f4ec1506ed4c3a1995b17debdd49070ce2f535ba598e0847206ec53dda52d151
zc7de5d8e32663e15bb8448387e7a495162b353fde5c5d14eddf7d42553acd8449e436ae1dc407a
zfc3513d2b388a0898aae76c8ece88e74bb56c3c9be01bbd6e9aa3eedcb022ecfa8aa0f94c0bf2c
z56bec4366723a9bc0484c0c87a5ccf9fdbb185b6a885a5a00ea3b4d5a2cb56cbfec90802197f9c
z8154f2147512b6720d81bd3144727c16ad94bc547ea7f5ff8280d43e868fe59f8f1971dd84e011
za7eaf46b70dc870428c458903369560e99810885568898475f31db05a572e1146550c31bc86964
zacd3d4ee5aa3a70fadc5491922fbf17b43efe7b52e9991218137e6fddb69b678c6ecf67f2fcc10
za168525ff443ece42407ea1613d02414a7d28a2df58c92dee022bf97fedfd71a7ef0bf2df04ce8
z2d6d9d7ecc4cfb91cdd2918da535e623b4eb963e92406650f1ff7535250fcb78cb6a3350730e98
z774ba4c8abff3e79915f5ed828a30f0ed2afba7ef9717aeea1bc8f81b577bb49b163824219b7b0
z47a72b2b75147e80522301dca061bbd0d2d131ac51cfc420300ccfec0a1f7aa5cc2e906f80311e
z1e7f585ae295ea7a12404a132c9e8749be24ffcf2137b7d8c38a18a8c032c9eea1c3ea0450b51a
zc22063d23e1886b00b8bee20720ececfd43636642872e43b4d2fb67b9d08f76814f93859839e46
z8fd7b4e5097d9c55805b0456f9507a0c14a567da750dfe341683a652e7f6e53b4976880dae1a04
zf618610ffc18dc295752118fcc8bbee8bfb758e87215d7cf387f5d4f37aace717456d0db9c74dc
z3dc667cd262a71bb37152d48ce05d666a0b445db9272b40034c078f05f8e3518ebbd3071d59f92
z02215c1f0f664a42105df749c68191a47bf36481b5aed4d086d428e7daa67e7147bc6ac661eb2e
zf445f760cf0dc0a196ffcbcec874e982640731c0d0a565b1601cc0ffc2ec5f83fd10a7f486a3cd
z3ab8b21967a399f057238e184cbe92fa0bd07628027d31dc03385295cf5c0b6dfda191e2c25c6a
z130bdd80107a741075dee214f36d69aee8c7b7b51fba325a8f45574b78dcc7f555d700e9988127
zc014e1fc50498e35ce47362d8fb948c90b232cac3ac90091842b00f011f6c21958a9d7e55f6def
zc597ffadca771761f488cf4cc99b2bf060bba712ecf581f21d4bb63957272e03cd9b6e9087b8db
z3eaa57945ce3a30051cf2efca74356999f5eb2e987f9299b0508b6863132568313ba3677c1519f
z453b9a7f8f8117faac0b5904c8d4c6c7d7482234aeea38b9997d98fa550522e606993b25077a40
z5d952fccacca966a1ea04746b22524c9933aae82f98d294cbcb12c4167dc8685d1a1ef1a9deebd
z9a9eee9fa89dd654eff80f25c18c99e38513f0dfd4cc81723646739122d5cbae850c6f841169b7
zc8669954670c7dca979d82cce1a9dd4d662b4269fca0f5c4223f6b51c3fa69e7bee4fae0534ecf
z2dbe331c48e53919f165e57da5d7713beb7ff10fece3667fca6df06aec18769ac00d4505364379
z7dc3e3d501ac2d4271f1c6c0bb8e6ebb2869cd684befdc6ae632d6453e7c0217558a68b8cb6c32
z0ea6c949f47807371f7b5dd6e4c9d788ecd87ca893edc7e0ee69336318ad08afd9fd3fd6d05aac
z6a78bf87d8d9a5232f8110e60ee7917a1b28b534e09c96daa8370c69b25c4e6b93bb79c9d71077
ze7f54a9a6663c5f3f9ba76de037ac163cab63f4ee40f0685e1850f509ae445d2d0ad9fc8652521
z491af44123016fe0f29e459008172b9f658dc00abcd1d0ec0dc57dd450f3fac465a5812128e727
z59e1f20608018343b84c83c74f9074c877479fd166f201ab1463e5cc7e20e412ae131bfd8cd367
z88932959f773461417ec501402072f634ffe591f9d0101c46c8cba94d91391e43f6374668438e0
z65a25c2e1cbe53ae47ff6cc5e0d24827cc0f698eebd888fae256fc06216ae5267e1b9e55c4307a
zd6ddf503bb8a791af4f14aa3e0ebb7d9b29fb9a7b8ce2b683505d6dd1532f2dcfc67e7f3f1445a
z3d762f9fe2b1fa79a290b292d33cb35fc7771c1006107468bf8d3111017cc4b569f16df3699b02
zdaa94fcaf950edff6724a9a034532390db864270e28bc97ff60ab95666cfeba39186710fc1c943
z0a6c86140e6658b1b33cc49b96528aaf854138b82cbeeab8d59d753b1411fd3b914a4cd19fedeb
z73c8637056e3815b3123c523a4cc70cf4bb01daa062ea671cabcf74c818959810fc8b18930bc15
z69a1deb3663e3bd308691d9cc0abced0ec9e748f49803326199cf263b7d2df698628412df9aefc
zca229be6ed12a1614911b5c815b6e7b0afc6f882808f788e9c58d1afd3481cfd72ffd72f7ebeac
zf5e4252c8ff32dbdc4e83cdb91ab7c184edf0ea5bdbd84254bcc93451428e281db2ab41f399c6e
zd48813a9a8464067809d8ecf9acf0fc90b082137eae9f1477c6a4b739b64d9cd646c36b4f57d7e
z8cbe19edbce42f5efecf1347da48ac67a911077b84268621e6a45fa173d49d399716c1753be316
zf2783ad837d5a1617be2398d2953fd63bb9900d1e4bd13c10952ead64a140ce13fb0fb5395e8f1
zcc682f475dde35d0ea30eb83aa22673c0e346a93762bbe9aa6ed96091a687b84be1a091e248a20
za9411c9e4e61793e5ff90065643f91c4f3f5ae0e03b347c7f349068a064c4ce501b860a30d57e4
z004cb4ff454cf0f03e56b1370997bd04b678fe7d74dffc72a0a01d8b6544c7feb9ec9eb0d5f482
z24364f0874763533c425633c6445332ea1fa559f85c6d6818a6668382b648a3cc306a7fec6e930
z107d622ba14caf84c25ae5a209493bd68fe412ac119ef449cd9301fd0654ea6f34252607440a51
z938bf4099b3ecd26ba3fa8e583c2501ba1510d54a21f6481114857438b7d4d8822d8b6a0ad97bb
z040aa96e283ccf61c2cef01443600d54d6e2edbdce49ee3386cf3a71389d6476da0bb32086354c
zc020b5e840318186d04d6587d10894707635ff49a3181378b21f0af11fe8ea01c8451189e0afe6
ze656c901e31b2375af7e958754bf83dc7a104a45183d8540d67a36cd9640479c6690ab93e1ee5b
z9f69acd46f49322a796e9cef3e2f958b7edb2ecad579a71facf73f4d0b4c0d3754dbbbdd36a495
zdd5ab0bc1ea33e7c25f0327c4be9e52330161fcdc5b031ee2d50360a3f025010cb1fabb9d974ca
z0b7d608a0d0503ae9673f5732b058dba02cde6d32e45bdf36e9607cea2596f3c00986e82935b0e
zd0c3699b200ce94e50f21ac0a3a8abe56c37044c408749f32f5c624e135a079c8f921a3bb849a5
z63a42775b94e28023716f629199ac0c0db7f0598c11398746988df1a4d15933bc2646f62e5975c
zee4dd7f204989fe98679fc7703925da10601e4c6871f0fe9db7873428a8a78ce794cc02dcede28
z9cc94d7cdf2287715b86de5bac3b15ff8264e6f3738215e564327b52963af0d49da48a70566f5f
zef2c99dd7cfa0de4a573353b62d1bd03f405dffda273ef44828b2d91f259a7f8db6a82aa10e2d8
z687a9086ef1a5bc300df2ba9e17cdeb3de4088f264a0d66d5a40f236c4b7d5a09bc9ed0d933c04
zfeddda0a4bf45a254d1f443c86ea5ffe3c5f3ee58921053eeb2bd0019c477104223b745f94c0c0
z14d1c182e48906309238b93442a98b535ddcabc20e58a005007e5e86685caf1deb7138cb24e27c
z7d1875f76466656a823c99097d4647f4cb3218b500407a07a82323c2938d33da54d132d6c2a77f
z2244b569da662653a5b65530ef67c49b42c67e08c299cdaa8f2d4abb73b229d45408372e0b7375
zf32e2d9b7f0f27fc86a11c2c56a65c636ca2970fab7339fba039461db0460e75e5b7f55e55f895
zd7ac22b94a61d202991fdea44113a53bbaab2a28967ecc31093867589996353663542edd5460a7
za7ee646c976fe81bf32959e4e0b804c367525059442448265dd352d21cb53f17f70dcd8847e574
z554919663bce60ba277f900a3f4e95ce1070292b43f6255f0943d4fa6afda564f6d89b98901707
z4abd6dd3444b731edc956af74a5bbfcc8a7459afa0505232749fe69935bef10948319e66338355
z96fdced383e1d4a3e5212e2532dc1e6053a21a571dc1680d39628a1bc878026aac6b28cb141e28
zb89fb68eccc0f9f48cf153e8cbefdd3d95f50139e57273ef369576c7f707a74ff9e844f89432dd
z19a4d1fa5e91ff2606ee6ad47823f37b937f61169b9295b51b1c8d3dff97e208c235329ab918f3
z1de682229a290cc88e2d96799f7d831604ac0368ce58d05af62b7875fdf6ef5fedd1b443868015
zef433326d4e0943543794d4b2ec13b8b30bc1e8e0856fd844e7b16ed7a5f4f2fd62f881a7e03e8
zf4c737a6eee2bc6b1e0e0acc65bf1a51d7e0206c6420b8dbdbcf24d08bdfe1a42008d358cc3fb7
z94f87a6c324932a8e3dae7a09cb52d532a29bbd755d2888a12d88fb4690443caa15bf0a7a8662a
z08d8eb16a03f9cd3642dedb59dba2ed0c3160c430d365c9380be256296263a6098cbee1b36c0dc
z813ce910432e1611a094f50f2850c4267329dcb5887e32d8f43841009b34ca6a519b7469129eae
z717120e3ed2e9b477f1f789b6bf6ca722ea12e34726ad266751acbe985f54985d873b497a166e3
z3fb39f392882c0b520f9733737e66e33202cdb8a141c86fb233f7f26433f3630350b87b71fc7cb
zcb6403eb18c558e0d13488743a122243e7808656ad58f3d3917c51880cbf03daa93060139b55b9
z00bded9d22c5708148cf30e0d99cd3809ccf22bf1849066d765b94c9eccd811a17cb87584f02c3
zf65e2285103c2b8f4ea2e9560a26dc52727d166fc16d863039abfeeed39fa4b3aa336a98880513
z0c22f211f6cb7faaf676f2494359b0f09c914afdb867c5bb002a2d6b288b2fe81b9e9ddbca2c1a
zc47976e8b2bcd4f070b152cbab2f93f2f0236f371a6287db9105ca3358286fd4b4ea6da78b400f
z13e8656dcb157e6cb9d995bd720c9b93994ca02d1d49cdbb85e423caf4432f77a83abc6b506a34
za24fa35e312b1501b22390521dea469203a393e2ca052581eafe07a3a4ae81096a306836463abc
z3f54e8a66958f1e1be0fe8fa53d49b343170ab693d22457f580008de161708c4687362f73a2697
zbbd7cb800011752f1cc8bbbca949651950dfb46d5b64910a7986555e2295255f3966183b18ef11
z7a8641f4d05c0167733e5791d26f1bca46aa833c78e5854010a51d24838aab48376b9c6afa81da
z121a5f81b7eb5e1facb2240aab9473586bb05cb2ecf098ac65664b119616143c631228a4c05cf1
z3b04bf35c52208377fc57ff135e0f549122fb75caaa95d7ab2b515be528223d45b45cfc8a67822
zeb8028ef319a6d3155dec28aaf9185aa3387036f06bb947f121408e5353f0b63fd2c1853a97de8
z452a2ae8aa65a7e4e10586e8a1c0405315f815952f5535b7462b4dd8192452ea2b38b08382b789
z08694b640a6ca1d6ea7d03bad59e364451eec0f40958fbf9df8e1896aa1465db9d8680d128e540
za39fa48dd81b275f09eee5959d36a2e3289cfe75a670fe86e7a51bcbeb69261cf03586032c6c1e
z20f25bd0c3d962beeb2080db5339366eac7c3ba7c68f1b26da0c7411df96c8bcb45ddc34807ca9
za67d5ad5a872281c2a36af5faf638410e93ef0f6cc977b386d8150c3e2b77501d703d58d5f0682
z38fa1812210e12ea5bcf0dc5a03ca2e493b085622898c1fed78d6d8f293c0b69519e4cd74d30f9
za404ea91643eb37f38b0c25750b1303f395517a116f5d36e4a7c2f78c5314a44bb66c81958e633
z4b1f40328f219b3fc67d792cbfad25d0ed387605ae0fe4ae82f44363c928aa8dde80d227a99ea3
z8c7f240f635b2a8a7c7cdecaf17d4ba62e1c358d6ad0cd11b9029082d4cb9e5662d36a2d0ad0eb
z6185608631153c5f34f6340fa97bb803af291e3d1272eba57e13ef5f272262dcdb16d5c8fec90f
z10fd44f9a21d5d8a72796852cb442207d11fc8f561358bfeea54c857c391f7f1b0724b50891d89
z93b124dc5a332a3d80aa515aab2654dd3b62bb48bd70281095b3fab6975f4fbced6be6061a63fe
z0821e169c91a416a7b4b29b08309a16129026638150abc4eb18a4824aa6ebb349a76840fefd802
zbc2e4cd7b8fa60bfe81d7fd4754ac26367b5262b23081009b1ffac1c26837330ac5c22209afd78
zb0c8eca86ca6e8228768e982aa40a120a0cdc85510ee28282ad28ce12146e29874ef13688e6e86
z381864001ed01a0537766716e2af56d2fc21037cc54a46a9a390785bcf3870f04b0609825c366f
z8198133fb49afe612d23d807e530d23835c19f31d16410c735f84f615982fb51e86ff0eb44fc57
zcacd4b740a38fbccce382033d0aeee378b2f7b556a3805f39a52320a193082725ca4383e9f6e18
z32bfc50a40618aa0ef9db0d0297d7c9c46197f124b077111589c4747ae250517062a4caefdaa08
zaeeb88f9e8a39acac3d4674ac840a23ad5edbe2509729d1548f393beccd1d407c70b562899c9ae
z53c45934ae6599c563770dae67c070658eadeff19b155999340ce33be56cfcf94c119575a53d51
z65250a42846964b5229e35f2a79887d785e2c5e73bcfbf26ab1b8e6496cf4becc039d71abf15b0
z4cafd20e452b200f1220ab92abb152eacc22f58772f281730bc9d5164a7ae939cf054cf7dfb42b
z303c93cd0cb0a76ba068b7764a703eda13c455b199d9827f1eda07edad3c44679fd2700caf1219
zc34fa190fda7fb26c46093e9aea8a7b49ef54c7f07a4c6cba20117243ad5cd93d61e0a1b659f7c
zcc712f2189632b706bc0031015f4853f25699792d8972954c659d9e05f3c8dbe0072aca351f7f4
z0226f105b66b3b3b70235868945ff3fcda7afdb7e0acac0e8b208b07e917b312aeade4979789dd
zd5a3784f51cbe014bb5ca196c655e8749f1987f0b5aa33d9259f705f991b7337149dd3a11d5943
z50328f5406378f0d4c73a3e64c58187f620bafa990e32841e6a12809c0ef7c6c5e301f790aa847
z2d53e1c1e050a73ca58134c0f9d20fe5ff983c8c980e7d4652547d330e9a13b29b57dcbf7e73dd
z061b4edfedc1cc2328e98df45667977740947a5c3d67b7e50db1829643c2b003a0d6bdadccade0
z7a02a5bdfa0ab2b80e7a7dec06f5b004afa1db1e9477707f3d8ab608ae4cf76ff290d80cf38804
zcb3c11a9eb36bca4136d0e98d6ed0fe0e1d7b3fa93d36e59b1381f580364404321475ed2414e16
zc85fc11eb4806034ef25be83c28ce4d0a7c79ceeaccd46c23054073ebac6a81bffa448f23203cb
z38539a81886661adca3ae7232da4007d14a926c114d10b02b58b6f67d125aa60539a16c1a9a34d
zea04094964c8a9555f7143a258ffeea28de5008d2b53141209a211238d5e5902764f8a59538755
zd429258cc7501aea07534d25c51b5df1548493b9b7806b6b876eefb2119d2a5f894ff72627eccd
z5f642d491d5ec6f97b1987cf9e317502ce84018cfc81f6607db459962dbf79b1a7b0f397a9fe29
z85b510d9f325dda271f368239e024b1c532076613675447a0d8371e22f91117c220b19ef991491
z98e27e2a9e008b17152637abcdf089717d63655a5b002da09d241469086462f23e4c2499bc83f0
z8a6f0299b71203e3854f17e85557e89d9032208a64a6c48611b6447925cadb205eb1e9d847f61c
z419a73b127b83612bf5cd8d8aa88a661d1fc9dcb5bbe03edca54fb12d4f7074bf4baabea1f9f89
z0dada66b0b21f09d1411550790a6c78134399763090f31b7cbd7585eebfc23c894872706b508b0
z39a827bb35690f6e00c2d5138439d6fe3734e53715e965207f53efc8c31ed4693ee4d1c71e47e8
z051dac48ebf757ebfe3abb439f2978ed28ea88da9c63f8c470ec02dcf5096d7e82c5c18da4ea03
z81ad6f4406f59342d7b610fa89fd23c1f46dc428129ebc9611c13d5d9387529ae9a56abc7c4b44
z88ec13979bf79393a2278b541bd51df1045a3a267f2726502dbea9c534e7ed9147a7f53419fb4e
z7a11876019a33a650000821e29d3536c6522bc495237748efd55c46b34ec2f2ca343535415a8c9
z92f567f16bff1f051dbe46be45d80f972f1508f6d9dc1e22eabae927fea4ecf4408c0e98f4aeac
zd997a54109ba83989bb901c4626300e7adb24e579772b2afcbfe0b3148c8ae5ec80ae158e0847e
z4d7a527897b12d86051230d1c410401138774ab15d04af309d2c2abc614d064ef30ae309af7a62
zc35190963385ae311f081fb2850253d8b63bcfb99c72f8b7e8ab00fa3f7d6412e931b009e3de77
z3edee08c7ad78c25098b54d525a15cde6509051a4af91f74ac3d7546932463c46fadaa823e4d69
zc127de14ead392e81407ec2ef0cabb27504d81e6284192a48c692a8a287ce5eb9c0242d1aa073a
zb2c1063102d2700ae5d3734b184da742a5a5ce4ee33ca3d86faf80139c82c9ee625a9aea08ee36
z070233ccef796472bba5013fbb76f6c35b1474674f2d4dcd9e61065ad8470c83d86ad42f643809
zba43ae61499c87b3672fe8aba212400927f06ca295261530a57cc0afcf703257e86ba1230a1725
zc8255f022d52fd6bf63f1fcd4dc76112af512507dfa08f487e84a9f4cccb747151a3e76152a4d0
z45b0d772943141cf9694206b87c9a02e8281bc2207108efff9525f8cf18aacccfa4111d9053fe7
z57851210c23b049f84a2903608a5141345869405e09d8c5f52fe36f3c0d06295c61a984953fcdf
z1c3d0eb97908796e15c86c3eea9b7442ee1cdb6e88cd874c4648d5e0e0511868b1d6eceacf8db4
z5da8f0822eeeac7521b0027e1054bf66d319047888351ee11bb6e0c0e2526ab88d5dd286eaccd6
ze7ab05c9db2547adf3d9eabef83b55de7b1d96fbc37ac969046f57c51bc4b858873f9d8a96f08a
z49c327a0a6f887c8bd8b38bfcc6312cbb7e74353ae7aafc4a5d0ce7a558a794056de79e01ddd71
zd85bce103a28926e6ea52bba950a602fec895c7565a49739f5810ce5fe16772945915ab59fe7de
z7f9d881374e9b019f1ed0833e0d3f231219aa638f21852f9517822f2f67c450eef658b9e933b00
z109ad996f9cdf94b30d0d2ace5b706a9a8415bbf15eb735e43e5a7321d09a81137439fafbafbe6
z4fff4cbbc0c97240c98a49453598d66d831c7a3e18bf50eb930a9b42eeff1aea2fcf4d8208513c
z68f6ca1f3b260859234202276cc424f5c868f4204efdb931e18bcf8454e4bcc0bb3a6b23e90e74
z5cf15248878118d99508bf059cc12c27529a3f76df759c906ce3930663390f26d31127fc18f3be
za75c897f126bd21e20be2caa6922de435b31281eff96d93f4000ce8041e85637bca516f43bddfe
z1e463f8c3a58825b05f1d85b36ca9b5bf1ca8bc929cd89e61954c586d9dcf885e9907714a4db8a
zfda15d2def0b8fb5642b02ad556ecf9ea9a2d820965d9b1a4061cf095e3fa6571d0acc4dcfde1e
z819a500e4e3cf51f03077adcfd7b3a88de1165e1bd36223b21fee91d61343f4ca9eea1401fcd7f
z0b66cdf6e23fe43414cbaab4ac16258afdb0dc0b3cf7d78c869c91eeeaa6fab47dae46ea3da56d
z76d6dd67ac2a4a69c1c96c4f2a6c1bc4882163bfda28ea92e178febd9cdcbb76dcf1929c1b8592
z236af1c52915f07898d28b48f9bf7179d18dd723b69a49b06e6b1cad6810302f05be849ec6960f
z9e880cb14aeddf6891b5c05b8308cf20491f9e877e60c995ef9f5d323d7e560a0f525eef692c4e
z8c6859f13635757b59173c1db0a1d650d8e582b4a350a44a7d440dc0f79359d7d445a0d159583e
z1878c01344eca25c1ff20c68889dd2e66a3813375d382dae3378040f7c41148560f58bfee252ed
zd751fdfe6a6b57c0b869b696ecf0da5772e424d4d40723c9dcb74a113071857b7e96e63ccbdc8b
zf12f61f1f26d1823f30607b4a08912b75c92ff73f97fc57c5f2dcc8a66f4c139e2fbd103083de7
z7061ddfca40fae8ba7c46f18ee62c6a0c8712ed284600480c71cdc265738d70f59171d06082f91
z79458c350f949ced9ffc3e326bd2f69f98cfe99e50ac845e40382da5d24c65b8b32e9aa9b79bf9
z9979fd0f504a06130cd4dca78ef6ff4b696407232057721ce9a057d789cea78cd6e78820ae81ce
z5d8e5bf232b2fda7d12201b37d84fc7613fcd60b9f4bf41b8c93e48e574adac3e6a883bb412f5d
zea6bd4a72c904c60ae5f137343c58391cfaf66538e040ab46a467a32c4a27b92d893a887b9dc06
zd806d990b7b2a2270617a65d7388e2043c6a4988104f93ea654e0eb00daf22763d4945331cc478
ze7ca45a8bc5404aa6460306d18e5cb1e5221a1589593842f276732f7ee4df5c8f70340d44ee49d
z02d73309b764ad58d561e0d4e58748a75dccde6a78b56958c10450c29311e610f5bac9d0150c7a
z45a7dd01b86e61e7111da5b6d094f145ee9d445836cb31051f02a0b3f569ea58016fafea69f8de
z9fb8e0a7372ed365e745c66de16e6f7177f555e2fcb5a15363b0e5a8e0de3ac9d3f9e0bcb03b3d
zcad42167300ee041863cc5858b727bb185a3be316228a748adb486ab711fc7104759e24880e44b
z8d2047747de7beada876725169ad8e9af8e01260628406e888fe1a1cd57c56c59dd49dc1d57479
zfb3e2a3d85d7c4282d91b2610fcccddc2d697db365bbfe9259be3723392716078b2738636b5582
ze20ca392962a60c63e153cdcd152c887b00f19ea9a6db0b8e13ee6f1115c6b200a4ef749090ede
z7fde536b8c1bd89dfdcb8de2c8a8907c72158c56342c0c4e0bb3835b6ff52bd9835b476bf336f1
z2552892482d203f2d1b86abc61568649b3b9008b23416f47c1d843b07a130c8107552a4b8d3205
zf2e10a3441dd53e5d2d4573d9fcdbb104961463ac853c0c11126f7ab4b94f64e16a1ffbca832e7
z6b539b1c60de733976bd216a89e4b8b73ad21ec4a6caaf98ec979e0dc6343537ecfd79e4126d75
z2c5aea64c5f2f92610ea46dcad0368eaf873f11caede786085a048895f4373c89d569a4daf261f
z46150aac04c8935d53eb35a4e13fa26569fba96d7aa9349985dea120b99ebd97212f2823f13410
z5f762dc76c914c786f66c428304d5f0fbdb6b5bb83c7b0a0b48a43c42253f7c778732084af41fd
z0512ab5b6049d1e8fc574428178a2c2ea80009e87c0a7fc88366901ed83134c3d0c0ccd49cfcab
z904f4146786b0727fcc2b780df36e2fd641a811eb8126a1949225afc3faa5cbbc6b8270399321e
z618f8505c64127bdc39f59bfbc204fc551e6bd0c05059d8c97eeb5728e45b01783526cd7fb646b
zedb9d5db5fffd7611c808ffec12768f5474c8fbbfca993b165db17b908618d7ef68ec2a7baf2b9
z369e9b473163752e8e1522a9b15f4d4bcf74f51528cb1f00341bc592f0bfa36a88ba076128475d
zbf642d66857147b630c47e18bf86c00d482a93ea5e2d5d486bcafe739c051e432ccae4316e3d94
zc016c848853c4e7807eba1dfcba50c0e238344ad7430055af346ab9e8f34f97658300d95400cc1
zced459dc8f840c4c3a93974e26a41839d806d6661402e8888e489aaec69d1b687d2200321a751c
z40f70e040a56692d97505f0ddf0b2e57eeaede94ac9be3349273a39efde886e49322f385294a88
za922f08f0f0df6e6aacdaa3159f6a6dee3418702bd6640389dc7692d6ae89d1ba3524945b22546
zcee8bd594c5f11d50035bf2d774aee97bddf8c266827f2788bf6a53d9e879e0517fa1f3a5db70e
z78673b264242600d82f07451f3cd3a3a0e203bc401964ebaa40c6c184177a1721e4d712a1fc3ec
zbf8a832c03bfda58da7f537fefc6870d06af2b7978ceedddb864e2d2382d7986f81cc4d41adbd1
z7cb7214c2a23d482b8cafc850f8d26e3db740a79d6d1c8f1c5bb061adefc9e81d5b1d09049fd99
z0675c2a73e0ac80552d8e9a01ef6532ff438a6a913bf8c2910caa8f5d3028f44900c1a954d62cb
z17c0a6c205a4ba4a0cd7bd64d2a61962bb52855f96dd5723a2a7703d42a6195c0059d4dbf678a1
ze11ca43fc706e136a463c57a8eab85ff845343ce4dece97aeccfd8762a13822633adf7f1679e21
zd79169c5ec03cc286060aaa9bf4582ad2f231726c96f38ac9634253b9b175e8b9a4823e2b32cd8
zdafb5ba77d061f5694d8158a661fa1b8ba543833d23fcff2a49b8cd06d3db9991a54957415cc6f
zbe91672822c4b7d7608e0285fcaad7c8746c29300fa54dc6c941abd9105118705aa9dab7e5a1c6
z5cf34dca8c2473e41fdf3f0775932a0d5da8ca46f36639ea9e808a90be2c51725a56ff4a184f52
z28db7e1c0e4bcd73bfd197a4f748358ec4928fc47589315109e3479b53979398f4b0208a2d4364
z1b3fe8c8f76c5931bcad2f058339c29bf354756646d2ecc607b472f30f38f4461508a8fd8b846c
zf70dae22cc8e2cc76cea187d98fbf65ebac91277a565862fa0c9a30839e58b99af30b50dd631e6
z4b63e6d2871c3f12e0fcb937ed267147fbeb5a2775975e14c8be25e1749dc0f14d135856a260ad
zad6ca4aa5ac2e88e7ad85d0850cb0c09622db85ccd8407d4bd3d7d677fd1f77a9187d7a2405c38
z6501e5fb26df5bcf89014e6e487eae15e2bc2ad18dd31d30b869defe0d03b677878f81ea22059d
z18cf3a4f217bf921c7d562512e709215cba9941a9d2a60da60e6aa95c7c38a86686bce8d6329a1
z1b879bfa9d8c53e1e683bf3c7f65b0f6e3b99473fa0aef5ebc99d9c23b72d63153eee246290be4
zea1a5bfeddedacfd6cd8b03b5ecb35e9cb8d0cc424c73166cf13dc012293af559d3de31c4eeff9
z57840da8e8164c14e014dea77c71c470219fb117f3296588ce3800645a2eb5637daffc4a22b788
z52d9b4cc80f8bc48c23d0aee0ff5b1dfdc069bf510e8b4c7ea445a1c508fd2dfee928b27e43dd4
zee7ff6ed82929834aac396d8049ba93735f091673ffc91a34c7e1b4b4b35337a7342560aab1f62
z40e731301585ffbcaeba5af46eba55b4432b95368749611c0edc1bf6a0f49e99592c4347c6b824
zb8aa800ba9e7f4473440214705892d43a29aa01adef2110f63d101a7b45f23151a8b437dd93fa5
z3f252f1184977a092b02d80c95287324417156ca90c1f42686de1a023a7226744337d9bc2c5bf0
zc851a149f66462f068bfe2e19112aef24e5ae3d95cda2edeaa2702c58b721738818eb312d6fae0
zf51969504c081bc22bde24547d40ad3765c68c218581df697653d76fb7cbbaf8758147f09e38f5
zb478c1e3443aad2f102b1e03eca3615b14782db76e018c9ea335e44eda9c3e90c73b90f9b6a2d3
zbd8d364952f9d6fd9b02410e32d3d23868119b147df5ca7e7e1b1d2a6d2d3af7553a5c7e7d8179
z714541e8bb0971d16a560e585df619988d2b0dc09c544b3d00e2633326ceef9eacb3fa84a441c5
z39090f54c9cd24ee3f568972b0022dab8a91dec7b939c6f9cc6f4aa60e3613e44542c7954a2f44
z6c633d263332095f1aeb4bffb8c60326e07ad3ccf58ea62e182f26378a8602145af20edfaf2da6
z8c75b08a71b7390ce64b258c8058b2a91b4e3be9fdebc2182b0b432bc2e96abd111e1174d50427
zbcc8639efefbd94cf1be1c30e16d3141ca1e6f6ad2522e75bbf4737d732243ca549230624355c5
z1b3528781fd4cf9347f6001773dde9a985a0e413af8b60a9d3fa56e3f3560ecd5fc914ba5cd7b2
z863d5fa35c9e86498204b56d9ab4c886eabbbe842695bd4f65dd653450c0b4274be0c86eba0b04
z663fd58aea0e5a5435c327b91a022da09578a10159e63909388cb62e201c7f21822f5e8c667ec6
z3b9a6aa768bb411237e6bcfe23ae61893f4f595b05f3147d3d191e5509e01c6b8c01f70bc22c63
z45f74b2e838fa7a5dfad3211dbaa2776c1d95b64cad63ac8948a625007b3d8eaa28913ed8aee96
zfc59c88c03b0988137ae7791ca8eb18382e35b81a10b500ab5da3465f81d191778d6b370221476
zaddd3719fbdee4e744cedefb46904c92a79807bdaddf7dae6e7cf285312f25c868cc058f5653a1
z231fc6ed5bf32ed8e2deb62d2175d1b966b19080ccfe47db21d12258eb652d1ab1f290209f9d1d
z1648f20b85044a8df207f3727ecffbd0260737c6afb68c445d265a540bd93de660aa6f5644afa0
z13dbe20baef05a18bb3e8724b16fc98f7709827bb9f4b580d2682cc287df389bdb9cf6a7fd64fd
zf791c9f11d51f0001b97a32b287401e2abb249b6e25ee387cd93d458ef9548e20f8f8782f7d3b0
z09f4e68608a5e5dd636c0a453a1f5ea9144f8f0824e8fcf060b1e02cb175e3e69da95cb02e5e30
z86e1bf22f91aad45b0522b98e9437429d1897847a4d87c5434fb20a5dcb3a7cf42d10f3693c863
z1470d882599d08a856c36784e3f97dcc9511339c32be70b1a97bcb10c0faf5cb46934265927e90
zfd6cca6ffb10a2c6c7029b25d7015b4dd36cffcfea873158e11b03ce42d25483356f22d5b2cf50
zbcfb74dbcba7639fe2947740a161f286ec5f6e70b4d7fc7e3cd43768633638e25d861a858ef7e6
z4d6b18e7b69ade9d830ed261fb3d8f0bd3508cd6fb76e9dbc4a38fce369565ac3c4a249d57b00c
z73e9f0e7e478678ed0f1805f2db7d9f4d9410c37db04818592ec3f2fe7efc0ec23110304723caf
zb4e13de2bc7b41be5812b167d6340f64c99b41720210c4b559da0c9d4e52e866e1a92f8898c126
zf6b2bc195307e3d1f102a07e6df44714d48412db0606273f16059f6cd6d2e02f9b3c6ebe7b8e8a
zf44e809394fb1c2b3a0bf5dce31d24cf35b72ce95fbe51424078793ab9e2fcac66653ede01b46e
z6bcbb8adc657a6ff5e75fec2f81665d74ebe094cf13d2cda283f228a45fd6e04c2198437a6353a
z5fa6dfd7c60e302eda819397d61017a61b5d9eff4461ab99aaa72f8b9459dddb911ce876f99050
zcfa8a4d92fd19bdc1f6a27e1c63efc9683b7841c70356ccce83c6e87feae8c392d0b0170cecf21
zb5046e399f74d2ec772bad4f213d2afb48e2f90c83b257dfebab143f788b16fa055f42df53991a
zb5945c07c292a3d323dc83e0d1f12a28e17ce742e113b6f9c5c7035fb4e19eaef017a1fb540eb3
z385061c5b0af38aaa84e629dbee3f12134735e6d96177a0849888cd80c56f1d63fbe460269ceae
za6f0aacc94e6dd4f37a461243f10635f129d9e714451998f9b199131b7d3f89de547bcc4e97c6b
zb13d366acd4fef8a722dcf96e3082e7035ab77e74ac10644c02978a1e0ad0e7e50482ee84b8eb0
za07584cd3587628c078ca0f144f054bc88b8d49dd9ab64f3b8d8a2d11fc18e03112c9f921e13f3
z8f54bde3cfb43354537af54df4281ff71c43bd1a12f4685d9ff4eb51efc802dbdca1295b160fc8
zbc6640fbb198e135628f64fb23d9f60653f0adfa79ffa56718ee8b51b5db34ba4e68c3050bd881
z495ff5168d45001f676177bf3a02a6345233db85489a53fe1084eb307f5e4e1d702b0ff8b80284
z26498715cb9179312bb049a2483eb3a5095525ad4da5c01da7427fdfc68d6714a3f98fe777a5d1
z8f02287be785e3a99903672a4d53f64e5d5a26b47ff13e8bf6436e84eeb6ae14b313d708db1645
z3f939fb2841e1075230580c496d1da2203a84ad878b9dbb3ac3a2eaf42df5b83a37d2777c95d46
z0f9da91dc4b59a54ec84d8388590ec4762677b89736167fc67a88a4802153178876029a5c9613c
z7d6c91678eb4e938347df6d3ce5da356e51ce761637a860510a9e376c031968f6a7b6ee9a7b866
zc77957496b6459cb1fc77fb581d973e2235e728d7b690e38c8c9f034f2a1ae0c768498c60f969a
zab213d9dbee63278315c2f60b87274375854ed8414f1c49b4ed956a78e721a76f3407ad7c156f5
ze115889114e38fc5428a25204e8f769166d3b7e2bff1cca473f1c28813d2c78b5caa5eb5524c3a
z23ee5dbbe400ce1721e33c6dc7e66cc084fd0f93491c46721cf1ce282598fe4b061a768d3ee423
zc0a4d0159a8afdd254d1e3461622e9552cd854e1b626c85e78ab42bf3d82e1f4fe9fa32489b8fa
z31249248c4349e38689398b15b7faa2801c68631e02600247cf49a010a7233fcdf7fb285f7e7a8
z764f42dc80a18b0fb950a582d0be2cbb491423f487571824262070da50b696fce3d938e34563c4
z632c38e40be4ad3833015ffad63cabbc249c26fb96d77a4a73ccb74f616474d0f1ba296dae37be
z815bf7a04fa21a1b03756d71aaf78f91c19d5420b72c5a35d955cce0e065d5beedc6aafc09b872
z416eb90985589c2723d9d1eb68e9c225cfe3e7a9f1eee3195d643e950061d3ff762972172dc729
z84fcc56925ed4c62315db2e00155de6473a6fbb1a5fd940d9b955ada5077b5b0d187ed7fcdd493
za7a040fd221767f1f219cc9b077704f2fae1534a3fe12f073c57bd22ecaf2751b397ec392325fb
zddb35ba66ff8004337efc75cc6f03779b50b62c8bce7cf1ba5f2de6cefed1359ba6af0694af742
z6be26a1ba0d9290397c80a00726b010b27b3b9ef627ad997c49624d16573239ed042fcecc344d8
z8d5e12efe993e8e6f3b703409c465fbe90d981a663dd1ad684b4e794f2ddbb5395b595b4c1e6aa
z6272f327735ea4ffd77d198fbe1b6a09f14a7611099fa3784d325681ed1739261ebd9d13e156af
zfb7ed773538d87d422e93ed80357f40a30d3dfcbb132300eb6d3f2ee471eeab6119913c43022ad
z53f125b1b6892d3ed0ba4931a999cb9a44009c79a0f2b5e503a9cd1129bd0e3a2f2e8dd80181ac
zb78a017c1f65591e4eb463e578ada5630e646c0f37c59852830f4409844f3f1723d17a6b9b6a95
zba997172239e1a36b6bb9bf16e14fa4d3d7cc66e0dcd8a24cf817a6479cbd055b533201c41aae6
z08bfb2c1af5606e5234c3b9e71c5a44d892e30cd07d9751b8259709926078a2f08e856ebeedc02
zca3bbf702bf86c1c672e8721fd4b175fc9b362f0ef1c0509f38975276a8333b2a40a1411b00ae2
z499d9e8bd4c6750ddd9df7ed22da0572e258f45b5c46c6283e4e03d90f347bcd4ad9b2518fdd40
zd958369d8ab3c2524773b21c2ed76cb6c00b6f6c8e73bde46a6cf4409486f0f9d944d830559ed4
z89fb2f8f1d9050c26187dab4ef411cb0d635a5d8f1c1f10ba51258053f74c6633f8f9cf92fe66d
z4e162bb70c24f6681f75748c28027c6b60c6e6c00750eca711006d7d6ea8dd5479a3bff18b7a85
za0ff7a1f904e9f0abfbcbad0eccda995eebea319b7ecce8d0b98b02624073c042d0ce60e12650a
z3b5cda806556209740112fbe92612b11d4b01d41476acbd741eb72ee511b79963b0944e0d156e9
zde97bbd7d8cdf6f000a346ec7ea352d4ea4b196833cd24217d7aba29487df2d2986ad909e83879
z17c5bec4866a0698661e96aeb1c2f52662a19c52131590343f4a3f5d28526f170c8c9f36a716e3
z4c6fa560dada3bb5aa62277ca41dc09ee6a5064dee0ff1e9ec28e4cd848c16b4dafc7f5cc0d172
z13ccdcc6c74b66fe046e9a97a5522ae33555dde71625955abae964b4a4092939a34022ffe1f067
z94ae84366370cbb85b1c9aef8de38bf3b70afbbb555dd72b821136dacd7ca4f1035db4c90ca00e
z9337515514d2e00e595b3a442d776d2fc6b520018981b213de013806b19bbac7368618de6ee97e
z0da7750b1d5a4e132f61371c98df9093233f100528265ebb20bfec91aff33c6ad085a2f2d1411d
z97c4ba50cb56cc6d3f20b4c915e0304d549291de3273ff760e23bc73a9c53ad4edd2378648a19f
z51375d0ec231dc40e99b0eee55ee2f3d349432b6de11179359613fd95de5db9b60c0815bdc8e47
z6ec0c940ba52b64d5cba1eb246a87d8f28b31170fbaebb4cb11250bbd6513b3ed180577a277eb2
zd7a9eb004a91ce48469772da0acedca850b0584d795882a24cebb34115b5a187f96018650f500a
z11f2616f795ec0f6f0c736a902cd7adf094d9ace46299d61dbf0832c2bc4623222ceafa53fbee8
z2a475ca030f1356c1a4a70a79ce1cddfdb9b0a2edd34624ae34f424f4d7da0b416b624beab6158
z8e89ef083bcd3ea57d5cc1ff7157411529d8f25ca13f7c489d68b6c90811656aba90b51bc1a817
zdff1de9d6da624bad500104b853b20c4585a4f9187081b18950bcf4a2f7bcfe2986d2f44089fd2
z13f20a67236b0169119e21e84a15ec546732af5584904485646912ab5535b0903dc63612f8d9e6
z706812bce1d412d6f6153b3903af92c0cbff603162ed4898231fc6bce8a61e46d9cc251aa23249
z8dcbcb43d9971d0dd1b38cfa850b9ad8385460641d6f71f0cbce2e57199b2ccbee983ca04446ba
z997179674c0204dc76c8cbc45b19aac4b797ba49f54292b0bf23021306d448878dfaf8d4ffaff8
zafde274d173488e5181080904b964d4df3d509cbf9824a13f8f149942d8af9f54b7057e44e4726
zd35cf645080a70da4a494b5263d2ca114ceb9390ed82185b88de2b512ed8471e5a75997652f8d5
zba9926a50e1c60921de4978e1a6ecd6415742c733fe2fd64a95e7d7b49ce9bddca353d2e8c27f2
z4522ea39f75c02a6cdc23b21cb68ca4514b9141a53e2e90d9c47da4f4dd8c75af1393ed7e81db2
z6ee70830377ee413491b6a238d62341b12c161c002dea7957aba748b740bf0bf05fb82bcc50b96
z8cbd45b52c07fabcdd6a8245d0ebb5f19b31ae36b8cfca8bc9bf5473521c524e9567e273c52030
z51be56e0766026a362dde12f2257dfebee8f61203d65d1f509fa801fbc7756460bd34dd985edc4
zf2251b9660c3a79060d16f3e5fb1fef96cf063a4ff5158de049601bd1bc92485f1c789bcda73eb
zbe24d497bd0d14b9d0c0322d7dfb503464df9cffc6bee8eb79d40e20221f73e07a1292d210caa6
z45205deb59807c21272c9a7fb05b6d153fb753126ccd2f18587dd2b8a3008fd850f55ca29ac00d
z53ad693185f789f15216057be70d567e0c63138033ef87e5f4c6e28fa843b7ef53b51dc7288fe2
zeccba1ed324ad7eaa2bd33280dd71c918145d7492aeb22dd2115a0b3b37fb1378b564c3cf58ae5
z7140b972ac3f9e5044d4b7b929b227f6f07e76d45f19003e0630ec9ad1dd06005c66a5896ed82b
z47dd9a57a91cb4af3fa10f8664cd1e0650ce650ce45e0ead3d093c72429b4be5b3b41e85d1eb34
zefec74a3cbd872ade64e0894735a615f3f2525d6268db3f0d68aca573132d6c65c3d72b535cb0d
zcd2bdd289db956787a3dd94b8f5588ab95250982c8a515d6f84e7cbaf8f7dc16ddab8ca4a7bcfe
z2b989072a3ed3cace663c2460de0c83842709f7d78cdab13b3ec47838e9de18da1ed05859b832f
zfe9e4d9944b6ac2ddcb8ff35e1cfb9400740c24329fabbbddfd41bb22bdb752874c0923d1d798a
z3dd9cd73b963107bcf194ddf586c03a20d0b0355bba7f868562d8ea44bfdcd0951e4de27e917bc
zfb61eeb5bab33e98524cc9ce8fa189da9c6ca9dacf9b57c8047cc6821aa76ad473fe4badd0ef8e
z35588571c42f94dffc416ef5561cae167ee898ca4db45cf6943b8303007d13f87ca7db97a43093
zb00609410b5fd5f90bbe6e58c41676f9e23df709045b0fa05d409fc91ba6f559cf78a508c27597
zd67f980a4099d92be9952239e5c242d7299718eda723ab6091ad19345c5704504294025fd605d7
zb5ef3a8aed97e5f2de8b7da0d9dd63b9ecd30d6c0f7479727d3d909b6174084d672aad3a850946
zfbdcad3ec6695d343803baed69f98d8a19aaf3e5bc6ec76ed280e1faf28b04be43230eaac75317
zfaf3a3c24318e7f2f8425b05c0a0bc1f7c16a2ab1c2c96fb4d08ad5ee288b96783428d9acff97f
zb9ba56d13902c79c274338fa86984eb80d2ed841be1aa850711fd4eb61be453bdc0a9e8f8865e8
z6f8224352016f6b8c4efc12df55c56e8e4f0fd5085f275d015ef423d1de472aff9313792cf103e
zcced12b861b74d46ce1a59e14ae54fdaa96176396389ff0de98e2cc46c8db8ee5b8c049e6f84f5
z61abbf328a415de0bd700b20873d526c8db2602c1210eaab1b707be94cca10dee2c0181f5698c8
z1ecaaa33510e1a8d2b83ccd4e21dbadcb61becf98d8159ea5debba574bf3a3249d48bf59dc4b4e
z9288a475a4bd2d44f03da435a34c7df34b946c0955c238018575e4611d95ee7f3afa09bc474956
z011457433bf9e4da2e6fc9a145be5c7cdd840f047ce0c7d2bb2e59440714e51310495943378f9a
zf37a1aaed159abf9950e1d4014ef2e7f6714c8bf3f3a636d42a895ab236a7f1c30259343b67920
z4c7fb3966944e0e8f5422bd4b77289e18bb48866c9f8e2a9797fe1a0a60b57bd86082942e09a01
z83f5c85bfe800e71c8f24076b4a3c6f8d79b0d14f1d69720e383d65e3d236b997ddde8b4a4d2a4
ze7fa5ca2fc8cddc2db891b77baff2f7e59f3300708ee622ac22043e95831b267d07381d157c6f2
z5c3c2f082f716f370b3a4589e5486d48a187341cf5e4d72e959857b85f798ba67cba14cc09035c
z918ee1fadd300e63e80a5a1c026db439bb16f4cfd99a7429133b0a2cfd82c00f2e049a6f63914c
z877263b8c751fc0fafe5931726742cea22475314443ae8a0016a999da5340f5c36eb66e1d5e4e9
z54a58cbf188566c31525e1eef1956e14d8e09c4abe0653e2bd3bc6c16a5a7bdb9e4fef7337da7c
z0187c5a04fe8c419caa28e70fb2bacba1b4fc0933556af436b7b2fe69d1254f09b88eeb6097e73
z0e0eb3eed501113b6237f5232aeae12e09ac2359704e133beb96abb500ee8314f757ea551da674
z8066c4098069aa8180e9ee72e020075b2702d10c3bbd0c819937422b35a7671cc2b0a2246e72bd
z0127d1f3abfb16fc474e86200983c216c5fbb4f5751e31590a87b8c918872496c45288b169db55
z022f5671a9fb7e9c35e9af44f7ea40c6580406d751424791e5922b1f941c1b0ec551719bf60b09
z0ac0f29c2ae74e0166dc233a2957ac02136ab536c272fd02ed75807a93d48502cb681ad2978c98
z01c231014780392cf66cfeb80f34fe3061ae8444852cc45eb5c232ac83bcb95b22439c46f0ecde
za13c87c014065443c941d500747451d2171d36a457093de0792873d71828989bf8956bee715b75
z7a1f14d3cb3416bc204087103574e45dc0446c15a454c4b526d4fb302cb872e665c41b4dc2baff
za2b34911384eb1554717b0e0808a6fafc8faed0b9b9bbf8d1c4e324e2e726aefe9acdc472f258c
z1133cb0fdc6ef525e5da5946d1a81ca51ee7533e0b2d25644228674c7f7c0659bc31ebb3657ddd
z71c9d88be1313648b16e1edfed17e1f95f3d17e72a5a290a45300f88fdf2c2f902a5014db675fe
zdcd462ec6546d6135bc2b0fc6e31d67ddd6699647040108c0a2d6db3412d41b5cbbe81576bc5f5
z7bacf1729ed612756414ec331178d25c4c1aa1c09eda3f9ee08a3169c09340768a6f71e28822ff
zf64a0ac58619677bed3e09f18fff6982902e092178155fe3e45dbf2b9be1e5dcc0152b8de8aaf4
z97754d8d4dfebecff41170580a4bbbb2dbf32dd57431f4896d9e66a81c056997ee58175016f69c
z866db82a1306b9e369c1e4e0527d92f659c278413ebc12026da9429b9032986851625aa7383f79
z68e9b2f5ace54303b5cc2df05b118d876aed0b90cadbe5884a7dfd5415d151c7e5470a0ab313e8
zfed8a5a12d68259805848999577c907eda848cef79db5ffeb3af8004ff47828aa64895d5af61b8
z649b05706f862eab9628fc25acab12dd259a473942bffec942eed8a44fb3e793a285bd14824ae9
z345b348c17af645128121bf680258ea735eea312c3673c6f741ca0b19dfbaa616038cb0add989c
z366eb876f8ee00880773470311aecee691096ad4f173150ad541467868836cd4595ccfed8a78ba
z2faca072c2f36c6f2ffc9a11f3c7397ab5150ee5dab9c00a076767d4883cfcb53cc303e8ab6580
z7a258b5d5ae39e8b6c8e7af9c626a28468de8315513ead218de5b2afee266fcdf3980ab114f48f
z84680512b2444e8af18ce08121fe6740a366f2cb1667adaef0f6233b6c4034c80604ad0faabbd6
za1d70cd0479dcbb25aca7554a0de7c5039b941be67787c355d923e4b9219b08610c6b85a05d724
zee5760be25d30865101098914dfce82cc3feb345a277aeb85074c32037978fcc48f2a80b6814af
z7dfaa4ee7a1761c7c8d7942ec67bf3951446452c616eca92a164ee01300f6f8fd52b2b86e34bd3
z080b809be27f63f8177a0111cad0326250bde65c1c5234000ef7c017928bf887730ba2e297e9c3
zd48f5a9a0c4fa0897712e722d080248280e5ff56e26eb1d15d448b33b6066f51ba81ba413b04f4
z50250dc527dd2bce5af885c00756884b445b967395023445a01c9f3b32bc44cf3840b77fc42c79
z03ed842c34e7065aa1d7a03238c54bed5b16625c0d5cfd43f2f38cd89bea44cccbc624a8881334
z9cc5a7eb8e57536c5326afaf6b583a7116d56111b7242745b43db4e4ab65e49e26e39cc867928e
z016ba54d6d6bac85bb03d4a6e16cc23c0eabce07778f0828744d8f48b11a13ae2dd7c8c8c472c1
z884430d813554af6386ea510768a0c6d12663e8434daedaca85064c3c10a9b2015c12ba817bc97
z1905052b1bb735cd2e9bfa0584653bb0dc841a32cb6a2b8462a31bcc05fe49ca019a0041410e05
z839ee85d1f9f1241a2fa16cada34808937d5535a8d0d7ff6eaf1c1eba17f4aa3cc4fbdec64f0f7
z5e9dabe86453ff6be3ff31482edc165c6149ca14d4ebeba235d17a702e8385536e7b49f3aeff66
z9ff421bd4c0c663661bed1711e90250b370de1cec8d82edf29faa57cbb5bc2cd1f251e3ff3148a
z9ee89c6d0998abb4f1023ccd002463b4ee8193890736bee1fd0a8a759aa7925beaab2adf7d6edd
z8f063e80d506f125a0d1b0b5a71972ef171c1cbf5c468d16bcd2edd92d365f639cb22021e976b9
z1a0da4c064438b09d3739bdae666e6c01c397f6e7c23fa6e2d4f53fc02b49f20fec91170bd050f
zd806b6ef1e000293892df51d73d3c324cb3034c0c78ca97a82004a4246bbee5f4da60c9869fc2e
z80b464746eaa8f4220398c1cdf24999265236452d3582c85eff3a8e80cb8c027c14588e0be2707
z05a52a9a77c12526510e703f7bb6eb4eb5c933a533ad50ddb7550db4e64675e323e460173f69b6
z3506ba090d78eee5cd2758d84a912de68b61903882eb90908d215443f6e8e3c5bbab6875d338a5
zb76759497aec16d512b4fd9d33b0afc4fe2bb7ce76a802f85fe4e95769ba6883e651f5c040eb50
zb55c6e796a312532c033cef22ea88a9384b69b9c6484c94ffc87bf3fddc9335adc5e93ec55db82
z4a156973cfd2b646a42e1d18c73d0d4e288b153e53a2abef0a8d3e0ccfe8059df423d6cafd2c95
zc1dba5a70ed8cdafa385a849ed6318f0b8c629f21cc2e07a1dc4a8661744ea1ba36224373f2e86
z52d0959bcb14495197138cd8f5367921298445ef541db8c6b0c50d23788f34d85ec69667f1cfea
z9c27c970571e2ac2ac0584882997d27d49876aa2c80495e97e9850f94df797411f5c3c0f2bacb3
ze9367e8197a1a3e603e1fdf74361e934d92032c4a8d4e08e48fcb260c460329e0f3b54b1d7769b
z5de3e19fc7495772929b48d6ce873269a98eb7f46842aa20c2ea7ac94ea79c2c5cc22a0f156207
z7719c9780cb64a13ee275b7e1f0b6e549871ebd9e44e4f21078ac1b443ebeac9fca5d674310338
zb89a1747d781bd281b54f8815eaa179470388fb47aeee274ede5f5a300ba9f81cb0e2c7a5b2b20
z65efd8f9c3200571be6ffaa0bf128bd1b7566d12baec7c3f865d8abcabcf8af873fb71d3a0a833
z14d5a9ac926b82167ea66bc7a36574a507ac19d0b3ef01d50cb92234f1de1622d8048abfe98ecc
z8917dbe4af32cf5d507e466e16e9038aadd3cf18d02f829df4000207571ef1c643632301ac9010
zad1abd747fa89f90d536f244180b6c91410a3148bfc207b282c58e1bcb45911661f99efec1b796
z8707f6d1859cabdde9d82e02f60e7d5cd49216f30b1d2d3754dbc6b97e3de986f8b887bb5bb62a
ze11bec005dfbdd588eeacac2c7e38308fc45286dd06742fa673a09769c9a798d67da4fea2deb9f
z92d52bc722ec1194cca7ee28684d285fed41358009a1007de8c53e1124fe0f38dbf53c1957494d
zdd05a77fb0d616f266cdb0cc6e3141d97b068a2785dfc4bd2c4c7d341a538f1af62f5b8958d8d2
zd5be4289295840d39d0dd9ebc2b9fa2b2ca997495c01ea275bd6e9dfc9d67084403697b1700785
za913fa47b67fea5bba81853b1e936b2ae463f418b59eb850ba00144f123014adabde0245e53b06
zf15bb5bd72c23c3931fe296fc9876cdbabe6836ce0e2d4da736a8d296a6195e3638384a430b5fb
z1421d88c8201e9f05903142b281d7b07cd811702d934c7411e2523a6fec0e85bfd490b3342d11f
z87e9212da7a90ad5681eb6bb0ca2199f8a080cee7b56b10db06553353d1dc312d4f10edfa1c6cb
z391d375d4b8243cadfa0658ca905b76c0320ed0af5fdf1314c4cf5449e57020f1a1e548e364a73
z4c468826aa1d26668397b2318cfb8b671fe3c378845abf0156a94d391246d90b391004c5a18c25
z19f045810d86ba59e38a4d6e33cb6ae05fac77031bea673c92d2f5374350e996549fbdfda1ce9f
za8c5a554f62da125ab0c96a8080b1643ed477802294163f09f4b6b0aba402dcfea4d27e0229b3b
z28a780a3e5c15bf08f382d59dee80367e3d54ee53109a17a932b231b475290c6beb6fc09ce2915
z0693e09128ac17c0e352696d54b3c34ab9d2a168f8a88413a44740c2be47c51209f8565a9c8783
z2c7173195d4b0dc16fae7fe6d87fe413030972ec0e224b9dbf459965d7c1eb8669bc611dfbe647
z36ac16d44cf364a99f30ce7448807e40bd8888a3c21edccd065ec8d8f6d9caf213637362c51327
zf1a0fdc6fa2f1cb9bf45f95bbc3885cd1da2ba328f4bf06ba8c2b92cb433a1070c8ae963d29aa8
z57da7ded94449d866f41fd669b4457e545d004132d4574acee741f9570c558057a1e4d8dc79e9d
z088e7e1fba05fbbf0de9180589fba1e9b0525f2545573ce6da40d379b7b9b6ca34bd852cd05bfb
z7d03c60a3c32d77fe670bbfa337a39cb69a1007ed7f404d01776d8a6d10b9731f3f1a0b024e36a
z3960d19e4fd8d69a287f870188c61f90f6af2589962e4eb1ec1cb94e33264397058ba804a37fbb
z1ef8fb43b595741115e9d6f00a9244eb1273fa45a3b06211c8a43e3a08f516c86e2d4614651705
z037a2c851e167df244e8bde151d880b4926d0573654f675bb788fb046c7dcf9f21bdc180b30781
zaa03255b95672c418d7868d8ed6c8f76907c9b71025e5d5b13ea98365dc44d0e7e5d769effe07f
z46a1bf9329c6fe23e8b410e93aee40a3ecc282bd4b441f876d42e6375dfae025e7395764e1247f
zbd7a7ef7135f1d919667559770a9ec24f74bfe683345cb28a09b6d08050a8a53b54bb3526e2d10
z882ce1da80d03b1edc265d1477e6ac143682aace67d2d113317d48f68214e121ef311a0689cceb
zafb646ba3c9531a17e1ec772a79397f1ff3ecc505bd2217b7fbd92ee18f0ac0fef4109874f4b87
z67c4256056fc8ec3a7cc46ca5d5334e743a91501e26ceda20ad870c6bc1faa4dbc520309eadac0
za6a23f6d09cb6f7c83590e5dc68883541f3935655a3f6a629874208389f8c595eaf5018e064acc
zd25e2436b8606bc0a4df04b485f16ada0e9689c7a6c029fae7aa213a0279374b6be3afe5847b10
z32e28ed0d7ee6be6aa0a91643b42c9cc121069d74ce8ef2b0ed95cdc414374ad71d6675878fbc6
z2ecd60d8148c3f1697c09d5dec0caf8d4cbb68c60451c86b6ea1f64a155f8389adfb2a19f2c861
z12b2ee388a1870cc3ef55181934310b8c2f9e48ea7068732acab8e4a0975de9ae3769669a92778
z548734fbdf0608f32863bf98b4648c2f443618d13ad54d3a461d1f48ec7335a1c8ff22706f5d16
z988e56a11cc7797f2b53e2560f1f552150c30a3d18f3673cdd73a79cb420de259647cabf76385a
z132834c6b607a58d1f37af211e6971f902db7648cd73ee83de50dc90dd84368c45763c9f099d0d
za1ef43cac233a64a4f0a3c4f773c98f81b6f60b6d710ccaffaeac39325f0fedc3302e18e77f29c
z7acfe1d543cd8d32f08c4cb7a497c8b139f126c7aaee7f007841f1371e074ba845b1e10fc41ce2
z0baafcaa21d962b693812cb964e4771514c7e373bbb2707ab372c52b546cba9aa3956a2854dd8c
z0dbb2559d176b7f00c4020c880f8b24c8e967502e8c6d4a28f4c6498f48b7570731df970bffaff
z2fa969b14703de37794d4176c23f9eed0ad0b50866debce2a5e92bdfa9d686630c4d9bbe935ebd
z644af6974a3bbf7eaa94ed1edb1ac2ab12f4592b5a91820f9ecb3bf9d43846e5441b3f9890e211
z45467efd2f68c23f4abcbf9f5ef1df882f7738e918ff279a3f3bd977450f580b480d16b3c03bf3
zc761d1a70cee61b46ca83e66bbbb7fa0e8427df0de70d17bbc50969fc520fd23058f09c516e039
z2ace6b714a681a807c0bb2fa28b97cd623dd871930c857e706eac6a8d9cc4791c2ab7bb8540976
z394c9284f7429c03802bf6005c5ad6a4cf39f16b6c96232071e65a383f6175b91bb16c4357df89
zfe21e5ea27215c3ceef5f316694813e3565b3c0c1365911f3263e0c4a02b9e6dd8dd875f9ef0cd
z4ef9a2c45264898da085a635944708dc7c3da562f8076d713064b8ae778fbc2a3db0b07e5aa2f8
z36926ff7562b435fdbf99dec96138d00c51cba9cb8d91c59b0f283c6887fd291b1694c7de5ba8d
z35393bd352939d2783071cfea64debf25fadc012d0b39610609ab2cf5526b83f7635cdb5e51945
zeb8c882850e51b670c7895ecd1e75d74f28ce8c2327810fa514c3b435f1e2df9bffd84bacdc6d7
zbd782ac41710ba1228bd7c1161de4077c812f70d84e413e619b8d97cda9df7afd0115a467b5ab9
z788bc5bb474c2c37bc53c8232d9a4457ffae083abb1361a0f2f6bbaf0af722c09683235e896bf8
z40f6c8c6ad390a86f1ce73199fc8bd582940bd202c20d3e1fdf706c0da5bfd97d230d9e0c48a7f
z7537e420dd7a88dba11748e7c6bd8a40ee32d13e952fdb1bc563199f327271b943f1d012091f31
zd8786da9fcc90b7d4e9072e3733e2362f1bba1a8eb150ec689aa3b5d012e918152089589fc9346
z7789f25889225ea7cb25073819771916b37f6d89afad2567ea9b424250140adeb2813f7bfd870a
z37ed9d2e3f68099cea3b22a35bdc465338481bc4e198d9dca829c4f0591cf10fa3ef8bee375331
zd53774b2bf5914b314d6434e939205b673f13285a20c3fe9c5ff38f6a1632abcdfecbdfb7a7292
z735de77acfb6fefafc41a94feb8dcb3af86d1848443718d2ec4a673b6461513d9352f19f41d7cd
z718da8b8053cc5f08c3bbaeee00ba320c5f90f76b997e192aed55d3043305de7541ac7b383144d
z721c69523ff012692580c6cc2357ca5545c94e0ef2674ef9bc23d1dd23bd2271cf49ac3f24c557
zf5fb7a97fd73e0a5b95d305f5c932b1ae521c2a4e3d20e593153c1ac4e12af94683ab5d3fbd49a
z228703ac3e817560394d3a7359be429738e2ad8daeb259cff13b68b108e4b0e55f96f9751d9f9c
z4b880ececbbcc0a94cb6597d44d4b46a654d5da37cb337a8693262540832aaf1c70a2ee45370ec
za5a29d1a13e5645834dd60c364e5d61f1202a90fb8954ae4df4c0399181021e0f69c698c7a93d9
ze916773a553549769919360c94eedd7754655b78866d5a721263beaaebaeb91382196c89bbd2e6
z83e61fa0a0af772559ad11f121ef18d5a7aa45047d9735778c9eeb04e84bae29ceee2234352bc4
z96886cb9c114e63393a5ba705ec3e6668c4a2d46317ba71ccb1d7eb5ae0af5f1844de4d5c80617
zdb08cafb74b8ece4090a43efa6934f5e32819ecc476b5e20a988b6644d15a3226e6e08e2cc5d59
zfdd75273895f5ceca0e0ad78f8a9dcf9a5b743fcf73abf982e0517f64c6dda59fcd2762f275a2e
z07116f34b340b8478b7aeb55ef7a78f4e93f7f7ec2a4a9e4262b4145fc45f48d59a7e8bdf0fe60
zc4a335a49283e919fcb4e451c8b28e374d2f801dad421c04409f688e5ce333a91c6641eed9b232
z402f314736ce5518a503d52576c206f8c7ab15efab3eedc34df2ad997908077b263e70d30d14d7
z902b915dd84cba0f32df4ac82b24a01e61e986e49e3e63a2a5fa2c2ea8060dd20a079ea48c804e
zaa0cb2e8b3bca239ddb48379afc72a95c300bb57302b68528fd5db01d0888e9860df9a96df10a8
z3f817fa29c77712899e4693862aada0f2bf62377ee74a9049a4f141478bf61d6c3f1abfc7a2319
z58b0cfa719594ff588626a96297d5d05ad05dd3aa4204604f4ceac322035373aa60c7fa69e1de3
zf2122e54ae7583fb7e9d8fd277498dad134576b405a192063d6235409b846e82e104d12ef995a0
z98edcf2f276101bbb63fefcb054ecce6033a80e24f8692b41e4da54426231a837fa81076fdc0c7
z3159c5a7326d2af6736274bdd8826b884e376174ab00e2bbf3a7046756358299dd32697aef1714
zc2f5f69c094ca4f3d40e169313fbdc9f68982f17dfd5b6924b6428c9bf907e391e261705f7ca7d
z8c73f72abf283bd44394c00c5304084b32abae28cc6037292a9019e566264fe470bef0b5096ce4
ze1d9a8f4fbdda7af7070e0b46f80d4d87b499d30a11285002ff3b091b9afac3b812ba10130cfc6
z7b4ef45369e55c6c94b25456c722d5236370b3ce6ea87f9b18421b503bf979dfe82507661b37a4
zdc685a96a5fb7ddf9c2ac4513ab2cd164a568bcde2952ba6a015411dcdae5567fde2b8b5f77cef
z5d6c9f2e0f04743b7fe93d751212383ade1b54f1bcf9c91b71e3ecf7c389f5fea6189f6e6d3daf
za7bc26df74f1580adcbdb35146cec514617098cb093853e440e05e9ccb74b7564aba74d848d180
ze8cd5ad8984fe6873fc4bdcde0de0262f2603aaffc08d812c1cbe8e0fdd0ab58a8d71a9332f512
z5d5e19276a23d4fc200804e51f64cced875ccf37afe35ccaa66823b939b13c68638060a229b9b2
z1589aec01db416e3100f5f9bcebca0c85d331e2495da74ec0e24e16fc7193b78225617bb0f6ae2
z46684e8e5d5f956668d8eb3aaae989b33c795d8a422f669c37e7d2b63098106a27df2913fc1b2f
ze7c1bf1fb8f288c4823c2f26e0df9bb5d977cc96a88f51f741f8ef428b024e2e097c5e80cd591b
z56eb3bf3b8019baef5347a790e9b70f5bb65cbcf605382b0304a73da26341d01a9bf45292440be
z67cfd31b9d1712edc8ec38370f8fa2ca1082f45b4d511955ae79de579813353a52fd6ae200b3c0
z9af18cee861e71a38b9939e31c582761db77d856fbc0633ddd11c0851573923cc40c6c9ba13f4a
z91da3dfc305ee293b315d7f6dd251552dd688f18e0efe0a0b3c13600f14a6d7768abe452970184
z65b497beea6299067e4123d6b3d7b3449607cc5769f371c1fdec9616e21f26f8626b7320ee3087
zdea23ae20f14037f7582351549ba1e9c95073d187239c1e39e31e84230808923ed4966a0892dd3
z1ad35983b2ad16080ec2a9cbb2f1036efd8c3e4b89aaa3ffe8dcccf98f333c4616d00cc60b544f
z6ba98d7127639ab1e1b6281ebdaed78a78451513c84776638f18b86f863637714ccff9102b2e10
zd855441daf1aa98b9d735e0f4552f2b55e1fedf6e2c5c444fc1ed72d36e04758349bba1fdd3f13
z4f3e6dde9268fb598a6cce0b72bf04896764d2d70e7aa0cc62a37756f4c711f0d5f77e37697dcf
z220bcdc24c4b2f9aa0b8e8fabbe7782e1cda5cc3346b269ac777c126b1fd4b4cf8913895a800f6
z4f8d2ef4f0f9c4fe4fb9d872ed89193855bd39ad4d66f6d4f7bb19304a4aaf7efd4407c8374da9
zd5013f9859651ada65e59b1b45d6556ec4f4d62b09797658fa96846e12c8098ae55f0ab2dfc826
zc03d3046e2c7f360a02ff1f4595d44f471b8fdc9d441760efa787f49af562c112dce7f7ae23fcf
z4f2cd41676de2796ead8514be231ae98f162f56375ed2cef9712d68e08c9925a74713fdcd8f24d
z7314ee0c8c6c968f51f10fa9deae1bd6c4e477bfe8c7de403243d880d3a4760b0daae926ef574c
z7d2379d45c9e8d161c619f06b3f493d1c4c6fcb27bdf8698b54be39dcb482a3d358df7385bb845
z0288c7c3134446576321a7bee606f5cd2eff9d580542854f326cbd185cbc8769ff6e51ae49da8a
z64adaa393c71f17b228912b68f7b4797f775b5b17bdda2b61e496eab927ff5b2576b3bb73c979b
zcbbe6b47b0eddbbd09cc7abb5dd00c970a0b8f3f1e31b85fce08a4eb719f7189b1bdb401ae7fa9
z2b3a5ee7f74534d7b4ed4ff1cc20e219030d94979e46b2ca2d942d2cf85dc7259d84d20ccab49a
z2c79fd32986091d93e7b18ab0381900707cb51c82d6dc3e9ac99dffd29d00b474561220cb502d8
z783469c467998be0ddc727e55188f2dec4bb5a8a0a23ef542910b351002d7f0fb5e49a20405f2f
zeb4cc34e51b2a617de11cc489a61b454b2f4a1ff2df2a163718676e983151ff30428edad41f6df
zb49dff9278f5e887e65fc8fedaddf3aa2727508ecb9a2084582d2f117cfe72a8d1210a51a0a70b
z82032b4aed44c3cc0e78072ea7a5205ff5b41bebc0367f9b0a1fe7e831d5255027ec5e5860c50b
z62a673cb18b833ed371170f8b4d66d8553e99792db645d429fa73e43ed15c486e5fe0829425cde
z63a26267f6f1eb5b8eb1cc3ee213ac6dd848d172c20237a068f178ff9610193c387580fd254b36
z870abdeceed415d6ecb40c2c64676a6baa2c62d7ee3a2a8ef92fbd1b861ba6cdc076be1c97f2ac
z9ae51d378b1f2d64d8236139828b0ba0410fed628206d51d2fde11f5b50033b011a3cc7577741b
zaf2b11ce7b9756a6565be90331e492df27e6db5c8244ebc89a8d61e221d16c27c84746c65d4f65
z588a462b5fdfb53f5d9a884489e9d4a7dcfc5e95a5a9dc0a772f3eb78c3d742a417e233ecfe23a
zfe5e5bce541a4490db8c8f0e3715e74e4385f349c4d994f47a72b276f921b25bbfd0a88d314949
z2548d05ebd20c3e7e1d3538ed156e179a18042f04812e94784c5cbc0bc5f5633f7bb5c464363f3
ze9ded936f11af5f26054e55c7749fda2f6a8b035b7d6f05e97d8e5888108d752d1d43391c5a88e
z8cf06a0e47af9f3317e77342dfc34f441fb1a14cbc37e86a8757091dbcf83ea4db28a794ff2dbc
zf522d08c896e2f00e59eb7438dd9c49dc03667ddca500dc00a3002111a896dfbd96c15ad94ad85
z21ff0bdaa1c8c6468f1e6b11234f6cb2bb69183875e0729ed8e3831697c762afe76d3fd5d15332
z27699cd9abc1694611c168c5487f072b535d1743f4164a2e0d89b2a084f0a1f4224a1ff2f54e92
z616a9a0fc20028f5a3740a8556f53156a65e24e6e2120ff238f239b4790ba099f3553f53b1fbbd
z61112187e9a7b2a5a1f90c7da97c04150ae12c2d3a84356c7d5d9661b1b4531c28b3f97ff6ceb9
z4e32d96aa7d3f5111259d19f8244fbba194db3f909fbf38bcd073ef141206893691d2267cf4a89
z2eb629a933ba71801e4c6b01081a024ad28311bf2b865d68effbb4abe454635194718c86463512
z4cf5509117ef2852257cae14af4452de221698c38563933fe615a9a9aa5c38be4661fa00b8d2b5
z378d2fd7cdc4e2c82f746d43862ef71b5111f022d30157cdd499bf512da4267cc96b4875bef148
z652ec0d4fbf42cdb8c75d2e328193365061ac7f42d80fbcc031878fac3d448215c358ddc678458
z5930f2c1335dc81eba4dd756b348b73beb225112cc7bd0e1e9a00f44bb15fedf5dfbdaa06955b9
z4d98dc87c8f10ef23ef3a9b5d27eaa81ddc6fe5df3f58f221381102ac1d6ed167ea6cb0f514e44
z846ecefdc75653108804f66fde8d2610e37ae1beb37968693495613220d1dd6023048c619937a7
zf65674897189fefb93e8a11d8a7e34315e6bb0a43e01636124c3fc03e032fa6c110ce67057cd8c
z048f0a02b8b3edd5afc1a2188140fc44e00af2ae3f683ba908f50f331c8204810eff8c80b48bf1
z550bd727506cd7d86bd8434d25dc8d9ad3833151b9bab6d7c0870a4fb9c10198d51d4ed869af68
z840fe2a764e4ce1d11702ca000a6aeb071192b4e7306b7d560038f9d76e6b14598ce4a1fe96bd6
zdd95b151d555e15b0f373d2453c7946e1e580255e92c603eedafbd942baf81ef192199b8b4826c
zbcc130de43920797530272bb0dd6c2a6ca7d16aa554f3ad53ada0b959c0e05a1039fbdb4042919
z82c36ec4ea1862e7dcd1496706c06ab1e00d41cc734810641920d6bf5ebbf2f9274f3c95d5092d
ze04225e3d8ad96826b31bdc8dc267c75a9e1bf00ee5908582784dd5edc5bfb5005ea45cde433ba
z4d9567642272955cc433ac8ce9c1221e0027add8b4151254f96568c12c348705552f78a2e05c6a
za8807a916e21e18c5d9105e72609fbce6185a660f0d0533eca73489c5367121a7fa09c2b384b65
z98d6ce5235bcf7bce45a162e73d57a846ad4f0afe494caa491947ca5d508ff3d282c17e70fdba9
z2e090ed5b1a1f06521cf5d1cce43abb575195f441c1f12e1be9966ba076d8a9b059cef57dd3db1
z02336907e00c30172d5e8a65c0aa45d06e5356bc433c6c3126015569da95cd7a4c3ef81ec8986a
z8448340aa3567f4db624c6863f36486513200b4f560fe7326410606ae695cd809229dc8c9afb6e
zdcad3a55f227a6f2b0833dacfd70ba5a47628e6057b5f558ceaa132f99deda13d8ec33ddc2bbcb
z8627ad7707bef1b0fb6d4099ffbded8601028a165bff99bcf738a8b384951ea2249d8e149e122f
z99a98712128633af580f6a2fefcf5309c6998c69011c8f0787c4b93833f9c454a0ef2843a01eea
z96409b3d6fc79a647822bc6bbaf70dc9efb92ba536917de7f4dab2955f240328331f67304d177d
z2a7cdacbccaf2839b336f4cfdef8c83811561b3f184be4f2a595cafaf0d52491dd6ee832fe41eb
z0f27e4fd64d6fcb153b1eabd6eb6fb14eeffcd08b1a5a53559a5d40755e0a62f6e2f4bf90468c6
z0d78d1a7ccfab4c251e82da5701d790223e76b568ee762808e027fe723de25b732324d966ee929
z01cc836cd9799a503c760f4e7b17b51aa10760a8987ea65b7a40e8442034c5f700f60ab49b5f0e
za445fd5c54c1aa9bd6633dbc106d4532fa33d8a686284a0daba8cf53ddb3143b2b3d3b126e630d
zd1b53dbfe219a4b09959ab2ff4d8b3fe786727842c234d029589a5939dc64ecb25d92c8a7c7a44
z56c23242def47af12a84c5f1ec59c470c4ee560af1b9ef5835eea6839e4a9c3d6aea92e8abf89c
zc320ffe5e6c04cd212034bf7bde69002e113cb2ef3f651f3a20b3c13ab0920164a17ee666de892
z0c74c3ab1b9beaee4930fd84ff49dc679399bd6ab7c69d5f6c63d1cc1b5f2fe18eef629751f564
z8c7705864556ef3aa85b45d0669cccc9b1fcf476b75dafd0844c6fe661e3aa3b6b88e9a0718b65
zd894fadce31110a7ed6448df479903959bc76d714721f15f7857e5444b38c6a516209b0fba1adc
z125141d7f6d5030997113b383a3414a69eee319d4826fc6b0786d203309c196270e52cb3d8a798
z7131dff70ff1117326ecb3773e2bbfc2fb2683bfed4fb6dd41dabba3513b7a52eee61dbf5d6a1b
z18bf60ffac7d71a12c2434f37081ae5854c29f58e6a1be82df5989e42bf3440d5bd47f9763ec55
z5383de4cf486fa6882ffab3f1f806c34a586d99fbeb9710d8f1922eeceac0f753d7cc6b0b12576
z8e4941ac08d03804dc666e0afd54af2cfc786e5514b0addbad644239bcbdc2560ca1be46fa655c
zd7106bbe1151465adfb62acb84e5a0e7542581bc4caddf0b34b43446eab5a21cc1fd1aef32880e
z302167904f645af8803fd6d9678a82102c249dad8dd9116a0005d425ff38baaf956c323f85054a
za1116af576e1d8600375478e34ffa28bd04fb241c6a3082aefb7f335da7553960845ebf34c9666
zab7e4522b1f1c1718e7b610278803cfa03e80ec5fccc5bdcbfd22ea91bff533c216e9d782f32b0
z932e161a1cc1ca47c93d40d2aa174bfed13db029630ae0a9bdc9afa389c54cdd06ccdfa07b83ba
z2c70cb58d6569fe8dd14f9556f55ff64a411a9f58e9725876c9f781216d6c8e29ae9041b4067bd
z91f65cad409290a6eb32fe78ae5d7b88ce29d8c1085287a4705b33994d0f0d621f5ebb5248b726
za79a4fbe97b01f875e8ba59aa918a518ea4473bf4ebd1794a23ec7c8aba2ae0a0e0f5f27799a1f
zb6283c9cf4600f4d0fb456c61c75c29464ae86c0abdc1184f824681c1a7e8743f9db9e7794c448
z6817731a6decd1cdded9a9e3f60657e3b386c3bf23cf852a6e1096e7a498cb264ff458b8dfd791
z85e01a7c2334669f59d40c3c93185a7ebe0b2bc80e015739803e9c0a03257f69047c33aa0f0f1f
z60d9ed89cdf314a693f1c7b2703a7f3ea03975e7f86d960ec552151ccec1c298c2a0f6a78051ca
zd9e5c11c5f8607401728cc2c5eb155382bf8c8d38d579189b0c4cf0c9b030cd0521e0908fa52fd
z19e804721b7e650cc2b2aca7f52c58edc484f9b775b5d5a2a6277a537fad68309fc30892738a7e
z70617f1633e72d5737edc5518a4f8455ea6c20160b43317036c7083d9d79356d3333830fb494e0
zd1e430aec580666f90c03f3a9fab3362cbf0f770de6fad0185c08fa9226ed54f7a08cdcfbfdabc
zc7e721465996c15d3b97c4749329f0cf9522550246b70580cfbe02cd56df53b8d82535c48a941a
za02e928532f84c5db9ffdeb5881a62b27ec0040d8a5bb0f1de9e919043d6ca7c120dacefaef873
z2e752337484667e4a82c5f1b1cd8468481e2b9d7e411510f2e67d6bb25edee7b1f13b6937884b5
z80a01f07eab7bedb09107cfc41583ada3917325ae52d4cf2b51437278a81439bacd7f476ee5448
z2da685547c187f31b91a1ff491899a02358422781abeda861e1a9463e6a475c62b763d805bb98f
z3bf6eb26cf7f9e6da6fe6e2187c79917711e32bd24abc885f9671f76b4be0f5d7e74ba75b67d87
zf1887993e5486dec1686ebc54a6a72f2d5da8e069b48310af241c5758ad6f829473fc9fc197efd
zf0ef7d7342a5a58d0cd0db11c64ae6b6daba3bf9883eefe71d601a8d85f2eccbe5522d7a8e11c0
z906df095bd5eb4730bd1175da169955504841eaf60f856c037a9a87ae4e43037b32f83b0fb29b0
z284226a8d1499898af1089d8275640450806530163e60b07834c56417e03087f1f034954953e14
z0eec8453f826be3b929f6aff91d8dfb674478c707d54ec9c0294abafd1d3b9706fdf663a242b17
zd4a7d684d019406ac1e5fab860f70ec796fe76e984b95e3484674b3265301c29dc4f7bc1c17d5b
z6af8c2ca4f3cc031be19f0092e070da4a3959619710228a25f786828f5bf25a94f7fd88f60fde8
zad2820711a96b74c521557b4ec181ea4d50b1b2107b4b0f3d9f536276869fa7f47b55e36b4936a
zadbe09b1191b9557dcc15dafa523f1f5e4fddfa20d593107238ddc8b3133257df7b60a1bb80dae
z10b2a80fd0bd90246702c3365b8384aee85db9cf8d94790da4a406064275997540b3f5179accc9
zdf170b613c2da2e1551a8bcfc059c38f2b93f50334ca86fefaae645f6b5c5ab8e2c87022a41a58
z4360b73064ff939bee454539796b7922390791317c419c55c65567ca85b542b83f50aaba06ae47
z75c39a8d3a1b2fe3b4a29f2cb614ad258fd05840afdde0a773b4c670e2f00201df233051909092
zc19ff001f1ea17d9a22f78d7985d68492cddc37ce85d6ddb2c0ea817a32309d2b1d22fbda83d02
zb15d3f9fcea7f18430488787cd65a9e19d36dc21e1e5338e956cc591394975b06a76e33ea27c0a
z19ced100c2b0db511afe143bf512b48921135b23fbe8dcd7357f49faf4c2c2aa1c45cfa779c4f4
z8655243e162e2da996d9bdab8aee1bee654887c6ef05cbcd4ba8e43679bdf26f7e58de7a7f8703
zab84dbc828b8477b0a5b966866139aa21d6cf7b0534d0f65292cb9db09dc831ec0070c594c07f6
z9eda80bb8c307e00518a753e3778fcf28a1bd46b29c6756ddb10091e7bc6e1f4941bc979a2e572
z265503434ba15bfe888a6d9e873330940e412e8a6942437bad03a41527a14e7fcdcb2a21852228
z9b3a4793665dc971de941d4ab733fe8a175212b34b6e58ed1011d8be3efda4b833841de44f402b
zd8e3a67b149f8953f109318ccb38a9b427223c05c3d5cbdc3f06e4fdfaa011918ca3f1ef4ef1c4
z4457f9a7e7ba01b211b0a6e327ff4acfad9dd153b50623e5b94d41577a6ca1f6db1ec9dff35850
z1b6458d5cb1207b55efaf94eef1a6ca38956598d45225396997a467af4614315f8b731197d7a7f
za02dd654e4775aaa4b64181747a61fb00f1fc6b38ad99f20265243be7ba11f5d67f488ce71da69
z16e0ca4f188dd1575cfa9d1c267353b10f00a2d379cb8a564f6d7cb34584a76944f926b9d6dc9c
z0c21953de724b292ca15b2319c02245c62e0964e1c345bb493536a934aeca5634b8fbea57cded0
za60179281fcb225f743e37eec00cfd8a0f6e36a17d8c426f8e66f71bc48036927fbabc04532989
za208489fdd62eee5a2ed0c86ca3173186a6d9e9c018d32ef7193d74f8a4ea0faceffc752e972b4
zd66238ab61088a466a42172edf5de4f03b3c56214e5da66622f95dbb7ba940fdb390673f559639
zd59c13ea8e54a8eee5ace6816afb94b346ce448d749f29de9e93a6d42f192fbc9ca98fadd43a88
z908c0908f223229afa5ec2070a3310b5ca5e176972233b467c99d0c80f0a99ef5e37489c3a31b6
z76a512e9a3c2415eeb905fbe5cda3c27012f07d14478b420278151a8fda8225974bf42a6ba74a9
z60fd534f562c03530127fefef16222a5eb375ecb43b6202e466a813da5a79b4562f397d8a0b880
za46d9e763c15cc173afbdb7a9065b6672cbe5b1fa8ba3d1ddf5649eda53891e077d570acd61ae2
z1689742bab3f35f6da501312729c6938d63d372074fab13f4e007c7eb2afe343e06ec1c7277e1c
z12bf083b308c82a946ebcc3af866b2900166165fefc4590df8cb5a785d201d82b377ab5380fae6
z4dd15b893a723c995ec36166dcde4c510209291f633f2d7a61fd68712c8d75465ae96af72a6cf7
z0520d12d5318054d8a8dcd9a924089c55d6ca639853c084a962b39b089d0fa1e0d3b7b85d9ccdf
z585665feb647c3a2de601dc81104af24b1f7eb0984f0dd5192037d0da3e49cf0ccf5a9159ebf52
z4bab71ae542d978c8313e09ae347d9c5a67c6e7dc5db0563f0d25fa06e48a8f7eaab596918760a
zfe7d311894c2754f741a04f0f7fd172ea045e324c09090ca80b893252aa2ede4ef78467c1bbb33
z3e432331c30b790b6d35c97b7e803399e8555234671efee0a67bd817398c4b717d583fb883d7e9
zfa22b6a98904b067a7276c2ad05d7b3d3a66efba340fde22bf177ea8deeee16beeec3f6ada735e
zaea89da92c78fcf7bb379ca79f3cc3935820620b651e3ff719363d196506b80f60f211a34bf982
z2ff7238ca74bb2192f29c3f97ccf55a1c665ef1deff5b569165a905be42c997dea8f1e631e389a
z535863e30842db757f5faed8fe7dffb9dbfb95b1bc0dd04f96798fe5b2c07c2b0ea00d5a7380f4
zd4379dc1a681719f116ba143ec5f866ddca635af6227683eb74402a7762fe1ab3765d320fb1a59
zfdbb610b7a79fd65e6fe2046618c6cc45077d8ca3bdfbf9de2949376f3d65f004b430da3b89171
z4a98ef905e4f9c3f1a49e9ed0af0bea73f3a389d1a0773bb92e2bfd1a6af6e0387b3de3a914cc5
z6969f5e86eb5bb69fb4b733f32f6483325b769aa80949cd4978d267b5997deafac70d317974ea6
z379aaf7b3fad8ada48533c0fd3c34e781db1c83a02558b5b2c0b7a7ff23220845476563e0b6e8a
zacae27d60fde15de76718d901d18d9c5bf3c04b2480e2c8b3956beb94756f41a29e07d4e468783
zfc7f7f1f8a51cfd9be2e85d8b24c04d00f4bcd0118b751eeb96dccf952be505f5276c968004296
z7a464fd37a629a36c8d6c577f09cbee6c2ae22f2d38d3366635fba681a635047da4138e3a492d3
z36b8cdcc1d8778625e721133b88ed12fed1d6ef5ba76f272471c34d45f9213f1354b17a1992275
z7a8b6c5609d6c53a08b9d93381e4585bbaf1f2bd508a26bfa544376277240f30881c9ca3d0857c
z20d5f6f6fed3b8edd61df46004f3e831f7805581ef08e2c9f6b4d0b03b3037d3f73e948b6938cf
z214cd7c5b7a939d786e37f77b48811a750dc04b2c554bd8ae9fde5176b38db62fe0f7d72a16c56
z8a6fd827b37b3c5fe7a25f9193a0b4e0f382fa84d33f873560740d33501fb40337aa9ea521dbf4
zc6b9da58584f6bf1f187f5a5dec1dfa61527261da73a1b9a6c7aa888c94ee11b5040e76e5abd4e
zfdf71461eb1766bafc0348725c8b61a24d8e3411760abecd0d65ad345b784ac2ecc3c399ab98c6
z06565e06965d284a2f80eedfd2875b41763e4f847ebd1faab83eff4d3b2518032a3160822cb95f
z16260e35a10d61cdddc8af2b1cbf719acf3408799bd9ade05f8cc8c7d82a02b8619f75c2740ef4
zc195d61e2205275b6b554a9a4c9a2e43dbc3b3c42996b7f273ef19d011efc93dc3f1b18b597d63
z2e11437d3154d4ab4d5538c6ba71b86024fc20fab2fad90a92a0335e07c1e6b80fb9645c1c71c3
z18898db09671c91693794f09dfec7a5fd2cf2e5a4cfb98e53568455c96ec40f018963b091656d9
zdad3053f7517c08c7d4a20af3c67dffaf84e429f55ef82904bef2170ce0fb9400b12606baf8933
z2cc9cf92b2a57cb4c2b1378402d8ba72e8bcabe0a9a20236f956609093fa599d77f2f0c870e4bb
z8def3ff29167e42881230f0d27ef42269abfa3b2518c8b9e3def972ce1c533c7b5107de2f15dad
z2e1a4e3afa0fbb5b356bcfbba81621084871ebe4f8afdc5fa256698f6102a91433ec09a2c54c2e
z0dfdf48b749d84d095c75abf0ddfe5a48c0474b495239624d413591e2fad23cb5a65cce20bfb18
z2123ab3b7e86843d352b71d901cfbdbc4ef4e62602b482219c25042bc7c712bc4bc673519371f1
z011ac8614532c584ad2a1e995b20374e35390dba3d7f7c14a9e64a1e91561827ea5a4a5e706d17
zb84030c81e158089e2e6ea391ea7373089184711b8f6c2eb749ec9ba944568ca7ce82036ffc902
z317b1107c24925ad1509edf625c01686ced36f89a291c9fbdfaf0d7a5b7b56ab45e1119732b7b8
zde3904926c21ba5ab97648bae7052baab8a045aa08cb37d157d6f1893276ed062033bb7edae167
z4bfebc6ff2add145199343c1c63168f75883cf8ed8b7a4ee1b0b9eb8a81e6aba39b783317a27f0
z7fb04f82dde13bafb4ffaf9c5c1cc20b409c5e83d8f6a8fe7a93630041096002dec1592ca6f974
z345ae1bd33e5bb994e2c30f4f9b4fe9f0edd1bbff4cd5de099277953cd927bd8d1db4218c61f9e
z0c0e9101885f79b549f84c73ce3ae06a994e200315e9940b0b9e42805e8d62cb1707a40c7a2833
zd362e7236d3979997673a80a2e2d48149992941d98d295ca358a31a2938b2ef15a957098fefb07
z338022da9e577b3832880ab6dca5446f701a34996b7f2ccbf1ffc969b9ed8555df0f99173cf15e
ze953182a6c0ce610ff34e756056416be9e69d81d3e531d77e62ef3dace6295e0413d2775dc84d3
z1714cae96ff3c8c88736fa7dd8a5bd85bce09924f04789df66a6b19d2f6a7df7ae47a53cc03525
z387de8e64e9842d20b83be36cc4d7afccbd6c8fdcef06ffc5f762e12bd2f11bd8a9c464fa8f479
z7b9e0b9498909a0e10e630556694bd32e263c74649f21180564e8a85341ed7fd265978d2f61b5e
z74db41c5d4b6f152d0ebf3f7e90c1925cb1bbe64aa831a88fa972df4888c1244589c321d8932a1
zb95ac5a3d1a86e7068b7428a9c7b1aa1738da6968eae7597ee6ab6064e26b79a40bd84400aba7d
z29a90e8ef6af71b13137232e8b218b73839a2d326594c6f2c33b93ec123c1512db96421c4007cd
z4a16bfa4f6c9d895d5d937ac24134f88a53c964f1ca8e1583b081851f5233b02a9fbd96cfc8418
zcb066bd6afee59155a16e1a65da24fac681f0f426fb504716dfb391149e2fb4b50cc5467d493ea
z2e536c98d77c128fa311a099386277b07c5da640f0482acd1e1e9af882138f061a7e864715d240
z38577dd3776ea005183653a9e885f4c2a08baaf8002c3df6482b40fba92229420850792fbba2fe
z94a29494da08326622506cb4810f4a83dd559109167b5a472cab63a4753041119940d8bb971d5f
z4e28a1c88290b390b4b017fc95e0be9959029cc3ff06cf154a158f1f622655b0e344e7ba70d1e3
z52bd784cae2dcba1e999867428a2512967857ebd290b60bb14258b607cad471b9483d17cd97288
z11a0c606f262a235177b896cf8e79b651b8c25d83fedabb4642895014314de6bf1ce8c16d60026
zc003077684fa5cb9f04560999915ae25b2f0eba289559d6a048843a30e45514afab3cb436eecde
z6d8f176e2c6043e3ce9c4a146cda7137114da7c9179a434f747eba90addda3d1121eb3874e36c2
z0f5eec6cf6bba022f01249fb4cbf368cfff54ab467358a3cc85736f6cd941f14a9b510c59081fe
zfc1165de4fbc195cf31c72073d458f0d62b788fe6302cea5389a15cc852b0f8acc1d86680be254
z3d33a1bafe50c101feb3abc97ad4d72eafb80886c17f44428556115718ff20cc946c32f51853d5
z2db9d31dec3147c942cd0d05a48e20858ab263b193a40cad23c6159c1a582f61673fa806e3eeda
zf8ee88f3075d017e38a17ca78c1ea598ff1cca0c76eb72641de0b3d0590ab539896798f82baeff
z820c37673c2ac1f99df46adeb159f1e6650b50850719e83dd1d99d4cd691187d5648cb74684ad3
z88ab9c1334ba9bb1ff6b41e9d69270bd0cf5bbd13b232b570d8a903a6ea14acc5531d83762e3ec
z27946a3b6f35bfccdf2730fbb4b8ae1f48de30f7315bc3590812bca0b885e07dfd278d1fab15af
z0c66dbbe41345074eca3ec84afc0bc3ead56e70a1640607f5fb7fba896ee4dae31523891d11a6a
zf9e4bded396d70f1e80bafaed32551824ec6cd97e06fb8c228f71cb53141f5ab6da6bc0318f64e
z80123d181502549110364ea7508c4064804955628f8fb5e2c665bbf4d9711a046172a68b4f9c08
z7b95b2c81617a51b1580410bc61eb3b12d64fa68c7143f64776467117388b7a37ff40898a5b1c4
zf8c08838c67d82eb8f97c129f8ad1155a2629b11f3caa7c8213c1ba7b5f3ab27697cb2bd0d000c
z44dfe77c081dad3a120a78fa82d12a91aa4b7c5aeaaa567d87f0491d9a649301c1f9eb427c0686
z8fafc14b2c8abdd8dab77cce95c39f057e977bbc2386decae45c9fd8a21fa7b88022b1906275a6
z5ba38534785f429ae008da6aa7657c5782954250afdd07727babca7316b8cc3ad43d6f1b47c3ec
zeedfae0664dc7fd9495b0ce152157e20f7182b7a99cb322f2b54e18dbf3edb6e8f46a0dc312910
z75a9025f975965b9e7b9681a818216a128ed43e71144441d8ed91df68bff39f2d1fcdd5f769545
z89af6ef5b9a0b5614ee5491614b5033890202840c1b76134492c69f0973b0b6abb66390944911c
ze8641dba317ef4658e27a188d842f4c1b0fa55f3a337daf3edf4685a1146451640433a41151655
zc26c78d25e820bdea10f677991cf426779936451c1c4f610e09d6fbdb9a7dcc854d74b67da6675
z1bfaf3251059c98d1026bd461725046703f9bbd899e51d70609383b4b306d5c898753c3643ef68
zbb0e0afee76ab3f77da53cee00d5aaa6c74f0ced20b380cc723f6f8a096db321e7dd424953bd57
z49a21488ab9e8e834b83f6aeaa3e0d4c7e3294a241f68c1bc07be3e9454c425b61e2779fcc0a93
z5d3f3454be0b33c18a59ed49bd996a5710976d42222851733f91fb760d644ee823daacefbf2976
z3ab3fc1c17b171f9cd7196aed3457eb8e35234aa450e38f905c96813828372eaf3f540f22b9a3e
zba80faac3696e0062a6decc1569248bb5af54546acd46145f252347ed7c24dd0f4797d74332a2f
z25fa4c7fe30c6af941fc5e7ddea76acb66ed698ecb8f42c5cadc9f7eed8d0b75a16b1b7ea14b35
z433a906bb1d3372350b35945108bf506d27077f5d3788ea0010f82a90aeacb64e41d3f265a63ab
z79450e393cdaf232c2ffa76caf63db0a9bcad1d7f7a101e162978d69d2600feb3282c32b773a0b
z802adf80a778f205827aa69ab04c3899717d149c7a1ee3766de7ddf947f8e047a777f7ed881066
zfa883bc122f2b42708e146d88c0aa9970c46535aa796100b1a3bbe36ac50319bc51e490e2be55e
z351b43472b1e4c48c7a93cb9d9fe2b73149c2b5099a01fb5d30e19b35dafe896fc38d3e350cc59
za9789d8a5ff4d8c705f39c2b1b109d1dd8f61e0b91dce4d6f60c3f6e26b35ff146dfc12cbb6f1f
z59c063cb0d36653115b76ea576d31a19b66a70b02e1e4bb60e7fb59b21dba6e37a4c12ea552180
zb6282ec8e02970aa370b4bbb079f3d94db4fbe0aca437bca60c705c6ccb416a898e372356f31de
z094dd74cd3c4b79de24bfc3207c43c3b6e91d9166bb47019e3a26e777726eefbfcfa27176a8c9a
z51d79a8f8175aa634b3a3dbb3ad14dcc54280e27048e667c5af21774f2f0f73f7bd743798d3ae2
z3d8d34bb9e3bb5e0c32f96967ba6f0262e454a77c3ac799e4f45942ece0363e405840d47b4d5de
za88beb9d6b9a4af62f6384713eefe6c0d95705da8d7e6f921600ee5bca49de11f71ab16ea945c6
z6b6a45b1a7ac8ae5796380416d92ae0d6abca48d6f17e7a34d3be884b146c463316a1229bc2bfc
z827f04d34a3cab074c7cbc9983e27c32e06845a653f881a95fb5c7a6a7d0b0d73aeb85f7f51164
z9341e1a685d5fb968b731b6e902e2bbda1bb8e81038d87c3f9067ba19d6d202b2790dbf817c4ca
z7185676a6fd7c6d67d037db48c078e749dd9e893e5b53a95fb6416935c612ae2c42c354272e556
zfa2959aa137a5cf43fda025241480305be78bcbac74338a2913ecb116b7e2b4a6374325c024e19
z655ddca2267be0da37d18b21fdc94d56bc970838c74ded22fc2eaa69d730e92434560524ffcd87
zeaa0a0a648e0f76b7524b3b37e5d9eeeeb1a27549c62873a7f8e2a54e89b85d0bfc803db698832
z221bb3ca9bb744ca3c9aa667c7e579ae8110ce9870660c5acac15ea55de534560c8d6c8bd11d1c
ze47df7911b2a5459536389770cbb24d71e93bf82deee312bf481e330ec75401d0839f175e13c45
z466306f7896f82ede01614734fc0961ce9a105cc32226fab3a39b15ae2cdecb342190a8e19d192
z4ede608f0b5b4a84bc9fbf39f38867afc3832a626ac705cfac64f4db33dd92f2ab0d571a13cb69
z69ec2c688ae930dd928cc8e96a9a81e43c9e15869212ca4d9ea1ec32e7e310108d76cc39ef8216
zb15ba368f21cc222b1fbefdde7dae16175a7ba0a52a8c738515a8f9c19049fe6d84774312c936d
zd042f2e75b4e7d3f38d9a0a1825aa1d6e541f479664f05654a53dea6225ca90136f798421db390
z60ef0b72ab2c5e1d011f117602edccfdc914d3b5f67901d3952af3aa765c643ed71c946b00e9d3
z40ff8fc885eea44636f8dc05270bc332dfe4b7eaaf11952210022e7f1bb08be932d5fe4f2e6e2b
z0142ef15215dca9a119def5c926f795aee8683b9fe3de5b3e1d09d141020b4ca1d696fee6e51a2
zdf82eaf62c200939710e054c0e45e4f1d5a2512815539de8656dbca6226c1140175b77f240752f
za86e979ee0cc94ede17ff968f88a415565928c33d1eb52f2a6372963516f6380efe271241a8013
zb5c29e568ee248c4f0afd077164db5e89449b52512c89c5fffcda707bb16bd07ca5228a9b83204
zbb56b92685e452829bc2fc320e9078a28d94e2c020b07fa6329b8500ae338a04817f3f3cca1eff
z1fffb207fd739ba2bf97e4e0521407302d3f1d913f7de20810802682db90f8b93b7374fe2087db
z310827b740f13b930b4ef75ecf508db808751135cbcd91757853f817f2835f661488f3042adbc3
zf50a4a7771c2a98a8dd589b607dd5489173638b10f3b6b4a2d427d2fbbecb30c774293a81c3504
zb7d2189bff2c11b9a813046ceee4761c5bc2147a66a8842ab73a51542b1ae07c90202b67566d90
zfc501f540f303ac2e92511bd3c1dc39877b5c2237675e64860e8740032feeffea5ebdf99bf799e
z7391086a6a61a431ae526c8671b38a3d54ef3713a56d19aff195632db8ff150374ac877bcafdf4
z59f1fce33c2f1753d4ea57b87da2cecbe5dfd2b88164a017e9832a01307544e5c26854d8321c2a
z29fa6102f345742f9d385f3a1ac0fffd3f73c96c9f1eb187a181fa0878fe569876842ae63237b8
zcbc791ace9a4d24bb5682b3c9a27e4491d5cdaefc210e7313a8cfa0d1cd192c211bf7a8f674387
ze46af0555cd7c25496142b3cf3be13ba34b1c437ce3e9f73e1fe297766fbf1b53d3d6bdf24fe24
z895308a0496c10466ce09b2f9a23f0e5eac08bfcc9214008d8391312287e71bc6a70c747fb43fd
z7aae665860fa1f95f403bc08ea57a1417772653edba0747c0eb27ab02d30653d771b1d44df2675
zea3bb68808c72a74de9155f7e2069b6bc1c58e074bd385e2e893eae3f0b90bd308bea65483bf4f
zd59d7ebc6448f74d966b950426efa7700354b9c498fad68223c2ae6e1661cb24dd03d7df97496d
z373696b19a7ba7a10ce4cd8cc5dab54a66f456dc542c70e92a41c36bf11a3e8192f0c012989201
z8bdffa244aad7ea612833ce635c1aa0269f3f07d580fe767961baefaf50ef71bf69191f04c7d81
zdc71c5ef5a5ceda50144fd732f3ef36fd4bdda6297ddb0f57fb5d4a16e82ee8afcf5c37e7ce412
z0574c426fa41dcde0c4f1129bab3e633825810b345889143783844a2046929b3f92dee8ee7c2ab
z973a890194575bc48eaa6df601d0e52c3c33ef3ff119d64965f073494b1fd46ec446a0f95143d2
zf012cf2f4a64e616ae27ea94e46461a47598e5cc30755d44e6ae5ea5831dafddd6ea9441bb4574
z0a92497dc511e884088059f2b2f4668056237e0a1eed6f599b91db715eceddda59d79bb5d97174
z9f035784a5da866d4e6c7ce24f5e1f300807088a4d5ddccfd491eb4abc50cc5116dfaca6695560
zff6e3cf3e72611a3a19a7dc6818599b6c038bd1e298f3f92ff5b82acb221cf85120698d15222ab
z14c047afe39a7ebdb6bce66a1d032026d4744e0dc3ca5b765f1e663ee64dbcdda934f64f7e88f4
z8a47d3180cc146cf9d669a2fb793ee626f3f3b0f9cd99a1f49fd9bbac968f43cb2231249130104
zf29b4441e7738f617b6cd42bc5cb151865757263536645975554ad8842784bad298a33e4b0a1db
z28ca1e80e44c156e7c331f93e603b10e7e0de17f70daf01fd23d7411849d580f9b8d2b78210b83
zc51142dc932b2902a2e4285253e4e1566646ff46f7cf51fd05e7dbb561ac90932f41adb5534880
zfe29d648d8f16454ec088caf54ba659be5555dce9b625d9b3f4fe1394ff653f7d4ff95f8ab7720
z35388caaf566a6415068c9a0b332f8dc7f98612f8aa06746de510e2ed4172eea2e527a56facc8f
zdebf66dba51162985cb340913223ab48e27219eb24283ae55d450bf470a3ac73197ec4f474d406
z90a89dd4f7e6312afc0d0b04c360bd0e446e4373092a2b7a764b3b42a30ccd04e84084557bc781
zbb9e5f54c8e0445e31264c141e40c051a720da1f2c015ada349f61c6cee3ff64074e7f45b2c942
za86360fba2f4291e3d53c326833b272e868f8f50906847bd3aed070b4e22a8d746c0c633dc1345
z3ec3dbd0eea1682527eeebaaef9d9d4c44d90bffcf1579ab1a93b0f3c9e3008e7354493f2181c2
zb35d9af21eed797c4a61846a9518dd2d84d798dead2c8e0740f3bf109f62246b6e71d46208e2a4
zeaf69f13dfc1f75f5fb9c9f881c258e282ba33718c6b3b4bef394b3dfc434b5fec87432317a0c6
z15867526cd75907dff66e1e0b0b860851d03b322d53a351e80d35d7074c4abc0676560b99d0ec1
zb296fc4932546557fc3836d208a557a1693659181c64702fb3fd277f8ad800ed3837d6c21bf83a
zf37c7b2f8b9fdd638b42500226b7b7e8b21a2a2d5d4586dce477cc257a77b0027e89abedc20422
z42ff03bd9de07a221ef862f7b826d5046e116bcb38c6895aa72ed2a873eafa6c4551ef21f22438
z52ccb52cec9683870373321a29170f7807d422e47ded0686d1f11c8b21c28442f8cf38686fc789
z302c8d4167f66a7407075963cbfd76bd7117b64530c173958691766e920ae4f71a11bfe5167600
z21657306236f9062785800e9ff7fc18ec445be06a40fec31de1743bb3392669d2e30cd8646a7f6
zb47f16b382c70faafc57563a381653c659ab52a4e778a97e9f0dba791b92f78019486cfe914ca7
z35cc56f0b2d1319afb9a7749487489d0ff722902c5f2d54b5c5c76ecc42b7fc77c9c47cf94bdf8
z74672803f1be084b117919b5cdd6b7aad0ffee7dc7fadbd1c1a9a4a3fba49b859e2fe845049f1a
z8b0e5d0eda9388038760f10d525602e7451360789b8dedf0e82a1a6fe68d31c7f246c76b36eac0
zb1c653d3df6d760f457f2bdfd1fdf6ad1892815fb3416d1a49c4a1e9cc01ea3dcd87669abd56d2
z5aa5c2c03f2affc44616f687358544f2af25c5ad2017b897a102ed20f34fcb0dcbc89e8eabbeb5
z80ac6777e09e64217845e4d989048fb7df416ff59e1a1e88af8ca472bfb2c8b7847984288db114
z15b804774c8eee8d8331778e1bf13e98f9087f9cf4ea9d33635c639e743fab8ef7c8d4e25ecf2f
ze96d001a8895c012d56663e684698d8b504b009d5f0c0b4bcdd8ea483384537cce9027efb6b8e2
z9f37378c158f8f91700b814545c666fbf7759512d4a9fb6ae0cf642f9d5be0ed0f6bb337d7845b
z5c7a683ad17048d855e08100e2df1a9e377d6ff1a56e793a2ac68bab0de2c56b6a3e9dcd8fe51b
z9ee7e2a4845b59440aff7edea306ce5c1c019a13e72cfc843413764f80fb891427aade977a9425
z92f4a1a19f102737dbd42a8c816715c1089f247077a7adf5a1c2afe95231e92be09837dd141b55
zf3d194b5efff831b691520250d56822763c4000bde19b1dce80d8101697600834367f9b09cfbc3
ze651e711fc5ca833db13d293e82c53e48f4b126a1ab6d12559ffb4fbecff8ae46978b947e7bedd
z98bd847afc2e94e9420b1883a3e2269e69d6083f43db6883aaa01290f3dcd125c1df8c4fd27b8f
z566008059281a0c2c7ff2c98106f0722d12fbbefb88ac8c914084e1011f26ad8b2c5ac107c2fcf
zb61144d934bd528b0ffae151e59ebd9c2718333a3cfb795d23b2006a2808b728015479b8ac8abe
z9fef4fc64100fb2b151759b447945f4f1d7299e15fbb2a960abf8d08726cf9cc6acc3dc7638737
z6f966a6e04134c79fe31bec1c21aae9cca89c34d43bd997cb4e0c7dfb8ea1e329e65fe3167c665
z0b85dcbb0d90c868484390aa32adf366bc4ec2d7c042126fc0bb16ce9e9c031d0bce0cc8595399
zb9f260d0f3b0115af57d620af1a2cbbc73becf57b0711d7c9811a4284732cc27a4823873c2f2c6
z86cbd97f1732492515096aba3729003c95328ec44024100f65937bd77b7d026f72995cbc50dd42
z366acc1e0ae1734badfb171c1e1c087df38b797779f376808a0820390956f5d688be8cc373c386
zac79ffcaa9299c83d3591620cd985c6f229be4f9d234bd6c844219769ae47cf0a1cdd148558d5e
z6c9f10d6e01cb6d6765bf4fd5333a88539f8f4b189c22aca95cec506b60139b8aba72bc1113ff4
z66db3a43e4d5b3497cf5e7c3fdb0e1e3622d52a6a9558be0f337e3686a12f17a8c308df8fef09f
z06266458d226ac7d26e72e3ccf397a8466e312a7dda851a82f282270cd8b8f8c38d48d427eed19
z7d299d6508547184ce533120bb93f4e3fe5c16232dc2192bd15007c82e4495b1ff11f436563c9f
z7a1c3b749d8da3d5e01b391fdeb1b1d9ccd26c5d8586ae8b714a6bb3c521d296f6bee8d245da89
zf1356cdb598906a4f0e7109858646492593ae2c17da082f1caf233843bc13a16de0274d37c84e9
z7c7314b6be4551630918fc2d427a390914ebc5205334f10a0cde6cdae0a6ab01b813ebdd378bd0
zc1ea47ef7aa2ec5284f415293f353db987220ea5ada77f39ac56e6d83e8504ef031cbf674e48f5
z22836b544aa33c2c06e112715962ac442a8363f66f640e0d2a7c6aaba68715d8f68672adbfa6ad
zb848209d629ff12ba0417fa797a4c7afa5a190ceae0f252321ab984688b718a650a854aefe2f98
z89d5005c3f134703385be2cf7ff14f715aa6e56deebcea0157ba422c85eb0e23c6b4bf067efd29
zbcc07e8fe0bbb3d5568b25f671c0f06005e7ba068c7e9fb5f83cad10fd6f3f079d31ca59a52588
z661193be43a8f3ae5e501cb914be100f2a7148524e28976740bb3e7a4c7eaeb38777a7afa99ac9
z4f066b32044c9e4b12a8adea40724d36fbe31015e27d73cd95ea2a70f9ab50089d3f96c88ba11b
z7a7764bbafdf453c4d38e3e2e03ddaa22017ea938535e2ea4ecbbc2c6698032eb4ef2db45c145c
z9b49f08792f44445fb1da55ed8db5eded7380048061cbad49ca88245ae34477cdd1bab6e3d209a
z2993b696e10e5e68758f9fa0619af2b1d4777b05b63aa77f86591044764b95b3fab6e8fdf0f8ec
zb2c9c67171d30ab8c19973d17210d6bed8e50f495c80002d21d53903d8da1f06df4020a7e58688
z934ea5fc7f35c6c13068ceea41e0b027dd06a2e7284db6d5894db55745850d4f1bf35ccce95bb9
za1c0584e3cf96e24fc4dfe70be55b936a93038806752cfa718777c4f415a6d869f679265d1189d
z6b4c157969cd0631774c3c6d4cbf1808dc6986c602164b28a1aba0002ee1e2630859deb057fef3
zb66b51f5b5c20e1ef08f0ce3fe47aa3cbaa65b6697d91034417783bdb7198389a09c5a1502faef
zbdd622496868048b60b04c00b93fc346ca90bfc702091e9b4909bd08cc1f4d0db395f5fbc58868
z1373c48275ae4765528140376bd29690c98c6b5781d9893b159ab075214c82c85fd81c968b8ead
zf278c4739d89ee1184747d001162d2b6a07db8fedb952d4ff77bc2d6190210b70900a92966a7e1
zd638e8d667f13470469e65963751c4f2e2062f5a20740a60c6f4d6b244a2d92c086db12b93b170
z440f71df05a7c8f6619b6a4a1cbc7fd382d9fceb28c8ee8907c3e25c1d3dee7a370abdb52960ae
z96014186d78e241204b2b735e86f41d04e14480b7f4403d46314c85bb6e9ed8a266d0a46f97bfd
z8b3af092b6205a3fbb613b2678afc398431de09f3c89565a1bb354803c1f34e2d3ad2878211180
z0f312d4c7b3cd53aa2cf97a5015314386c9c81cb04dc56308cbed7c4d4a690a940a12b78912023
z098337a7e45f6c9ed1be88f33cb1b3032748536875e4308dd5cec1e8c2679345935fecb1d14728
z8818cd1ec159506a04113a3164701452d5c22eb9c477312cbf4574bc54a1f41f4d1f4247b30e8a
z9d4cb2d1ff921cf4a29c104e4fef7134b017d9ebb1bc91c7fbd8a0ddf5b72ece063453d6157d2b
zaa72e2613e9295375b3590c2fa1045d019b220899e7c6ff384daf704777f0c77a0a8dd84319a68
z10b7898ab6a0a62a0e647f9c583a856fd96e223eaf2207f8e114d81364131762c6c3e6353a8fcb
ze74597ef628fbe2aae24a288d53c06b02f20375ee4ce03734688a6c7d61e3b89dcc3351c036ec2
zc5a0115c7d6ce62abc024a6c382efa39ece91b47cf0fc40606fc13302f3486deffdb847dded817
z0b3ad802a6d897ecde3a03b4da02d7809937f22821373a031bc51ae776df15e980fa33ce17468e
z5691e1495f688bdb3677c80d93fb556157bbee71981b7ed79ec824022ad30c48f493738246ae40
ze3c7f7211f11f0549cfeb097dc413cde22a6a3205ea1649b7efae5d901281a0f2a7f20e352eeaa
z031b714dba4f92cd2da8154bb92aaa17b32798383fb18a3f09d3f2659cc02dc0f76e8e61934c99
z0e7c50bcf11c55b39588c479cc1d657d21e7cf573f8760bb9b4c163eef3e000cecb0976535265f
z489334815dc12eef1fdc3b90cf77dbac1c160d5510ae63951d5aae79c155c68ead26048626deda
zbb37e80cc66d14df84c588eba7db0eab656febc242767eda2a11dea83b6f39c01503b6bacca331
za47f227912d70ef080f4014649fcbeb1a77ad6854337f5d9b66b8269681b19e3ec3994e4d95250
z4eb854864f621ee05b1e2ac40a792ab88a81b882e18bdacb3a42c3a228a7d09cf32c8ae076373b
z7c9b4dd2aeda8d3b058839dcb0e541319e1917e07a11d6787ca8617b87f50a72bab5a04a0ffee2
z5a8940a48832b638c14d14c5bfa810b8f0a4775437a4ef4518231106bab132926e5fab45ad5bd8
zefcdcff22b1a12f2f55083f90b9ae3cec13bdeaf5f9ed0b5f7e473a69e6de4632dbed5a0583da6
z1c87e9c61d923866da475d23f45157e275859a48a5a5e57ebaeaad6f74574fc7c93dd1d43dd1af
z4a4d8f64a2eec781471d1980245a2fea525e82ac06cce16fa6b154b069f88233f575f0bbdc32d0
z7f04765f386e933346f298db37b2a3e423a7b179e8177ac2c55b38560545e4a02f5b57fefe6ace
za95b2b804fb40f69407b5b16c71bf99fbf32c3205483193b60901d47ac169ec84fb1cabf588076
zc987973f12f6cb3ac9cc839d3d8b46211ab5b7035baa4c60e682f4a86341ab2e68b23f52e71f56
z183b0a831fc7f8fe90b8462027e2862bf19a082cc3e71994ece714be74f3b774f56959f6b67ed3
z5246c33c30666ce5bc44fdd105fc3f5b1e13f9af5b69cfa9290951ff424d4eb79595e5e0272cb0
z6615d2ed500fc8b998259283b04f55b68635866458accbebb5f6a485f9987b5d05e039657be0c7
z69cf9e1b5e80076ca339c63e38370ddd76de8d67ef218b354be6ceee4c51a1a3ef72562abb5b08
z4709b3711636b089588ee3b07c151689c2237c45938ea4b707fe46d3d07981303cee65bd7c6fd3
z42c067184186fb51d3f59e133d5855332379c054ef377b98404333e96bc09e0c6f0f1d0827d471
z83ad60a5a4e32a31162cda25233500d858a16a0a632edbf0bddfce5eb2627644e3ee7882a48235
z2b65fab0962f355cc167006e1b372de1723807ce4db90bd8dd3d3ab74523f04df31e9c52285339
zbfc28547f99d903b07747928d3a64636e9941c751aa687649211debb97457ebb4c5402d9c3e41b
z07e47b2a783c4bef84356f4f77751baea8b607f4551f47d1140c38174f66f9d788cda5148e5634
zc2b78121ecc5351edc9fb395ba558937655a06986ac775cca17b76c3dfa193cad93d472a8eae09
z775145acec908f6fbbd0e24a5e054bc8eb6c3de5da78e1ebd962dc6c8c2750472893c0d84e3fa6
zdc4e42d6517298d692ff87fad9db9b9946033e0144eb69a74c42ff80e89416c3877cb2bc7ad2cc
zc3257bdc8ae598a1dc15d5998557c512d6b587c4c7d49c11bd8236dc83d81cdf236c3753d560f2
z1bdd8df26ccb50358f89b75c624544adab313dc7fad1fd27bece1be3fccf6c222f491680f0bee4
zffba2dc03c10ea7c64c57fa548254168ae1080b548c45e41d1ab9e8ae7d6468b6bdaf30a73207b
z294985c1ca79c572eda4f31faa3d0fd13b7423e0d029354a0b294d915b765ce11ebc276aacf742
z9ce909a1736112a6ea7785b12c821b0454f864ef5a8d60a75e3cc270176c583a30fa35e9411c54
zd894abf1cf3e2fc02edc39809fc80f83d7182b9ab9aeac23fb219e206f6934296292c2166ab804
ze8da786c9fb7adcd73f38b33ab1f8e294f91162225dee5feddab131bf8216c482161e2d7338ce8
zddfe3c7fe7f23ba4645f2f1050af3e73816763c108a7f8d97b8b18bc8b9a2adb3df652c3b6a014
z60ce2cc0bebef12fc4cb0e535fee02b22ec6465f1ba1c89d8c54985897a8f66749ec6035aa116a
za83eca03ef59732a3ac1a488bfa20eb9172d27f2a8e1f13654e953d44d358a7c1b3f156833f605
zd0d95cffa48a6cd99e0cb0f1902ea60ab7f6ae1859ff83d173a9b31f1b2953a6f3ea592d8df81d
z9e7d3b741931726c8e15cd52ebd3a2cc10fa8351d8227465a051fb3042627a849f99b533f8960b
z10372a6b35c681a7f60147957b3e8e5706f0c77b712290730d5acdedf12ce1c9a2bf5622a0535f
zf3601392f052e4f53608a8c694a78150876b88ea1035a0b90e7c95ea1d3303c317b86787e49fa0
z2a518aeffd6a2ec9fd4ae60fcc725f16bebca5d6afa724b19e4d17603d0b29ac7c20d88163a7b3
z3c359bd6f9c47d077f8770f2adc1202db430a6ec50dc7711b9d4b80d94ba2b1fd3d1f71654963d
z3a6289b65e7e9e731acb2a0df265441cc487bf36e5696f35d8b538f9692514182ae648f2c73530
zde74f5ac3fcdc87455ee2240e07198a961a209d1ae6a3dfacd72acace9add8950c2406594f162b
z0fc8a9a0792699ec4298e68133f91623e8ae0bf211472353378d64779a539a726756811b4743af
z2604ffa82a7ca4261d06d992fe5b2a04b6ec15c351b69d77f07c91000d15f897892cf21252e240
ze60c9aedd5c74e8278f1a3bb88d95e694dc793194061b7ec871712fa8653247f60f54d62617ab9
ze32bea4200428f30ff6dc52d370499e88969ec8c8df1768d971ba22ddb046b7b05624778634762
zf5bfaf53e069b6783c9c9f3fc7d544c75d515169649887cbb32b2b2a4ec621baebaa8241c3084f
z9584db661896700252eb968900f5067efb78603484598787aec233aab8aaaac2f0d3d79ffc4720
zefedbc818401c263e74b7b6eeb75b04f510543c6bd20d3964d58246ce66d86145ffb5025d03c64
zdc9383b0e7b99039d56971aa1faffcbdca3f5add9f1eb894ae7da197b18b9d1d01320c553b2081
z4ce1fbebe4df2de31ffb350fcd29aa1593304628c297c6d9b8b333fc34275f45664fb2505ff0db
zf5ab6924835eed83244bab8e80a47557213906b066e12a15f3d8693bc011a03ad3ae1eea2f41e3
z9fdc9615a713f4a85adcd563732f38a0915555e54c185e1b33e39c8cbff1f3e3c9c92f8d26d3be
z94308a1c341ce66b6a893e2a2b9d179154d2b922f7af76c00bed64e17ed88f49033d2dcdf997fa
z322468dac92aec8eeca6d51a31711adc84941ac66e5da9da707f5158d11eede5e69a8576e238ba
zaa8251030d746bb6a24f017aab297fd9116f3aa8a4a5ea78dc400af4b4e5fe81bb9fb0b150d882
z47f03fac337c575a61ad07d380fb18b9ad4bd1fc4edf02b66c8812460952f63ad74c2c6d62bf9c
z6ad3d390b90b50923e9021e35450cc1b274387370e7a23e17e12af5c063d65bdea754f760ad078
zd0962ba66b742a6d6344ca6dffc33cdb6714c972a4bc9a617dda53d768d173ee4a7ac750b01896
zf9f9fba7f85f638e8a0ba8ce84b66fe7424aae1b850d9c861ef173ae7231a3246cacb065cfca9f
z6161fadddea4c80d7460f68101e7c9933f2d0290a3c662aad4fe302e779c0dc85190f564776604
z6b2deb52a707183bf7c08b91e779e84b6e0a8a67c8a0b96a93279363b5b11fb9daaad1823b5d68
z56c422b535c34b901bc2ee07a4562a7a19c4f3d8aca67f64ff9f5363fc87aa4079f8e65e39468b
zbcad88892793bb844dab8b02ff540e2140509da44a79bcf6eaa1a2d496c610070af87703897239
z1ca418bc1069cc850655eb6c803fca26ab06816ac93194fb346a50e5f0f9e2dce7354c37bbefb2
zc101ead71dd752face8706f7f896ea8006e0bc0f017a48cd1041a0c2d2ce2ee58e1cda61c77d17
z7aa5e1afe7040b0f379cd8c83a7b6628ca9f53bbdf35b8194712682b5aa41e56ec256ad4c76158
zd897bb87854c1d1e9264e02cec89661c38bbdc43b83de16985f67868cf3dcf54bc24cc3fe411a1
zb7a199b5da1ada7d475dc8c00cac57a94a94825e7f87a533f3e564d1571774417ffbecd8952846
ze4f8cf227b119606ff8d9e7feb139d1552cdf3cfece26ab5f66eb29b0e7657d6f93b81d911ff62
za159127fca1dd340a9ae61a59f2370666bfefe653f6a99a326d8514b9a8a1dc50136f3a378ce53
z2df6ac147a888b7185520910cd71428ae4693aef261e6e587bceeeba6601b61cad5a5d99679b1f
z212b788f0777fbed3a9ff0904d6a017ffe733ff4ed40be252cdfc4cee66811f88f32c5f9787df2
z900989403ef10b927f77a566d9e7b8d665132e08d8165b9c933d0d1815e7eedd27db22cbebed86
zef04b812d6bc1fd940e1887249c65f8ea4c9dc8cc01c477dd920a2ba00473093202867e7f770d1
zefb1d0719d9fc5e2a572b4c088027632615c56db04aa30f57fccde2534ff7b46cf73ae17daf5cb
z71da015cdfcd913047305121dd3b882a043799c0ff885715efae6af0c42ab730abd0fba3eaf7b8
z4702e9dc6e726c50cab77db1c63c8680973cca32b8d5dc0e0bc22938dc4f51a94de2412be36256
z931dc9641d1f975a320bcf0716e177258ef5e5e5b4fe7f8257b39fc2fd5634f25e57360e0016ba
z5b72809f1bd4f3cbf6ad0069768cdf033f7de6a07e902d69b709227a2e176caab88040a0ce7f06
z3ea068a0e7eb50b07fa53f9fac18357ff3e9682021cc65343c0038d2a2951f2a0268c656a98b08
ze981b5fea7fe6725e92ec2ce8710c75a21dc47b03d678b4506d004c20ba3a2d22ee33677188c04
z1081ee073f01e8d20f1d818d4d8eb37701f12a67126eec007742dea4813265c074b436a4ab8829
z3363f274e201587ebf6881dd44675fd56d275c052bb8d7e01a56d81dedd4e9d5a95cbfd817c584
z5548a2f2110526de1b8f9123ee0c0a25233af9895993d11c095c45bb479cc8a8e61c70d6f6953a
zd2d085dc640208227a6cfe6a70aad96e027c5fd2e7b94a832e5019ecfa87351344fff89bb03154
z5d7153631f688be5f7dda1a8d9ef79e9447adcc3cc2d65ce1ed36a6cfc9e155e4bb7642e1b004d
z0b09198ee194b06ffa13d2d6f82ea7aaf3a798e32dcb50e542f18fca9c12449e658547bd4726aa
z930627e866fd8f62209661cb3a9274135bd7925be22c4cbead901a8faf017b15b78d4e0f690703
z1ad906eecb4271cb68ac0f09b2e90bac8b755ea047d541525aff866d4a15c1a48117881e4fa626
z9b42385f36f7ae23c2ffff1a63ee9b419e9e97693aa7e8266d5b8fb835318f95abdebbbc052d69
z79e6621221042f0f235cdee306e33162f9eec438751004486dcad649cc77655556b364b9bbc946
zb7cac715d574b225f95627e82d53a0c7add1e815e4b702d99c8e0cbffdf231c84655d96f942ed0
z334be488c6acaec39a49156a87f7fe6530d430d52c9bfc7733309e2b788eedc6cf7cf888727820
z82c5d8edc2912c59e0568fd256fec4586ac390a5c271a16f86a0a15465734005d33960571e557c
z2bd88cb0a5aa96f511dc55ebaed09e39c8baf58604126dc7fb196c92693d6e3d9b33b4f46227ef
zb4f0ccd1bdff5203ab5e456ac0cfbca5e4fc15514fe2cff6eecd10ce5930a27fff02d52e09b601
z54a33e7c4b36e5c0346ec7f217aa090d35033b6e9760dbf8d0f9903d81224d62b535f4b451ae12
z49ba825b2719af9c7c3864d75e98e6ff003fdff0097184751337cf273d2af9c8bff44b1069757e
za85f5d76a248d7c636b33cd2d1e5b607b31bd2b88cbf0c0cb565210173ac766aafe423d04cb506
z6e8d7ca0782aad50b3b8a0567787dd509db9a7781c6ec6b65afde1f2794e7d6f3203952b228a3c
z2fb76cd11b4fa7d3db5325e16b1949b7204ed74c3fca6d96396cd43a0741f58814e6d25cd130a9
z2331008f40a6336d85514c7f549f7bb421be83426082af68020bb0e67d1d64cb6db72b4ef371da
z691fd530abd4134bc1d3396466c479f7656db4e99f23edd49281ae76d51e7a7975d8623152ce4e
z56c843e10b34cf36b9bd3d66fcda416694c2c0d4bb26bd7d0637d7b1e5bcedffe10f6d9da18bdc
z761bd5f47bc2a98578a63ffc6b50fa4b532077c41f1fe37a0decee6ef6ee8ecfebda2b2d528404
zd5a0da90e71a4e269dafd5bd2f6bfbe73ce030512f2c0d414e3a8de3bbd3dddfe7e68c2b3b5f83
zba61fa6a0d212d81ec160a0fb9ee7d577ebe1efdd23af69a101164cf1a61c9c019c555ccb64318
z7cba685a46555aa7abf0f73c37479846a6b17459e6c96dd87e9037351bbd6544d92eb42b16236c
z0b6a189bc6591c6745f34b613c1542ed14adddb9f1a536efa3f0b5ace204e5c655ad61864a5d19
zf250e295ec3e3066b3c3fc1efab801b47d3666d0c697224d110de5dee85a576bc060fcd742c178
zd48f139bf5e593c3f553dc868e368326f319ab4fc38ba589709afde30d8497587b4dea5e38f693
z2438033db94f426aec45907c6962e5c333d55af44772a3cef6eb38e7cc4d5c1fcad008ad8914d1
z81d45341126fdc9fcbc26f120c2db987f32bef1bbd82cd386fe3e0dbb7f7d6c917c6eb61f649fd
z1448bab4a6a43b0230cd007210e834e710a73d1705fd3860d202b01aeccec626626540524c36ea
z3b1b5f7650fac0c8a6b146d6dc8ca68bd5030aea815a6ee378869c05702555518d872c06719570
z44c9412e1a968ef33960d2adc9d1f293c06a1ae29566acf71e425a9b336e7c31676e1790bb2fb7
z06b7f6066f01bc598fac51d3b3b6752c23c70ba4105b79d5c4627e0fbbcab07b23eb3ff33a5a4a
zb8013918832c05357d2e1b5f38120a787becc20386b6d4f2bad2b3a6973f37f468d8d628770b3c
z2a71d347ce09b4bd028bcdd4f79b6029fbf0b9d8d01283a464f9754c22756f723cc5cb7273ca7d
z8533378acea60c2961037fcc940629e7926e14ee48c1c87a048d0cdad2c800338b9ad37e35b9cd
z704e49de42ba8c0f0ab07bb072d0b47070a77f613e236965729a0aec55c7ddc1c6962671dea824
zfa7e5d510db861695290878b7940b4ccd87ba0dc3bd64df3257c998e4c577161b42c3e8675c3b6
z77d2a5d6094f7acad111a6bb49809b6c9c8b15763c0f03743f5c28a3f7e904d0b41220e2ea4d01
zaf33a8cf4662ea9843543c255f75110aff52c8ee23ea66ec20631bc72ab01abddf2b35eb910a49
zf0b3646c70e5aacdc1f739a7bbe764a525004a50c75ea4efe0a55766eeabc52019925f00d3e7b4
za64944728cc71c96ed0972fda6a99e658d087d177e5a94bb8a72540c133a36e67da0adcab99fd4
za7c5c2ed4df70ecae68bf76fd06a4f439eca63bd682c3f74ca4ec9eb63c2f007aca0a66ab7322b
zce7114b265a0ba2af079faef7ea1ffaf04d7ca2dc7cc1f43180a3e031f0398c34fcab3f4435307
z165ed44cb72ba148cc07d8ea84891ddb2e05278d8ec0bceee6c9f7f30feeb6a69a9843879c7788
z4389463a572d6993204e7acc321c60879024781624d39806032cfd4dd0009724d0fba8470bbae3
z4e1b452caca744cfbcac55954804d8b268d284357337c4bad0e1b4129a56a0501af2f5d5856be8
z6709ef772b4720023c058b7ddc42cfed81f13eee292a81c0510eaa3a00e677ae3467865315c5af
za6406af61f2c5c785f879ea1fcd55c0c18cb0c372a0b5e6f9363fe6439feee4a160f16e2ac1fe3
z97114533abbb9ea339553fd9b72d080f90dbecce323141e452607d9e958670a13f3583014b859e
ze8dc581fa9c1086d5b56d723730c32cfd666476843cd797b6b516bb618f9661c0c95535f65b6a5
zed307111cb8a62dd14c92da74ec241e916183ebedac7c952b7b4e23eb7a972c4a4596ce3a1b896
z7041a3d3501a092b3a485a27ca51f46fd7f205e6964bacb3475a86fbc26f6c771dc7f1ac79223c
zbcae1396c51787abc8b3ed46eb97a8175b1e323fedd080752cbe0f730d21185f144b51a50a7639
zfb36e56d1da9e44398a33e7be8447e6d352167d34b25332c05ee9ab8f3f739182037128581301f
ze18f3c576174c0cf3d69696a63f5d2543b21d2e2957ce3081a18ee8e7d83f944cb1ffc64348425
z2288d1041ac381b444d91e08dbaaad89e976b566085628e4e6c3b1de11a2c8890b694cc9a014d5
ze645c5f7bc746e4d6ce2ebf49c82de51807e5e600801b0e8f615f535ab9057c9a1d9e779efc3d4
ze8c181f61525696e300eef8e670eac38da54982b5dfb80793fd46e584e1c0dbe7b2aa28ef80116
z7283bdde290663d7c23ff8080bd0839623c7b450a7c24694d9d4c186572673937aa56c106f2be7
z9b26070b1fcaffa1f528313c87988f5fb11868c68296af0639526ad987dd5e28b55f88ae12f0a2
z3f594ca6270164b965cf1f3fce9e9767b526f9532780a403709c27bb487d20af740503ed87ae55
z627187e5b3ee7156989b92e6fd66c39a85e8c9ab1d3589b3fae6fab7e26de5e48a40aa3cd3e4a9
z54983c3666af316a2d76bd09d2248b54a47d8d41f2e9939105f57ea6ead3bd07efba67188d86a3
z9e5660dfdb993173a4c9f56258789e8703d9a31a4e915f12e51c1903c2afe9df004300bc8e4d99
zaf22156eca866278b430b7ee352f5d346600128c2ae78b637422d5fdfe5bce5f284443122c3eb9
z2b787a6196bf8851e012fc2e587f46f8721a3205c0ea404586c6479f0b40740438b8417baf8933
z291d6690e7089c369f660b0f34594e830473721d7d9a8cb10b60450c7227d16e8133d5dd7aa6c8
z9d45ac83fd2bcd2afac626537b497c166ea8d5a48389b14d8e64a2a24ceebab867af6155517ce7
z30e8d2cf1b36bd149e3f430c1eca26a74f4d2c4cce410dcc59769a9763181aab6769d754fb980a
z0d8104202cc1ef9e5bb2ee3701a9ac42770a39766b415dd55df24301d902442d3d8a0ba393d46f
zd68c503815bf123a152896e1891c4492460ee0e02f70b88b015b22f5cb7767b2b1c04c736d27a7
z6bc982c0d1563ccd81679fee898681f347b492cf82cb994d66020fa5ca92f8fa4ca980bd915a41
zf40fc68f8e77bb7d28ba4bbb495903d5282b1868d863592773a69690bc504b592c2d08c5f2c0b2
z5338d1fe751736647dc14ae6dd5617b0396415a337b7c9b118bfe194903791152c0f2e2a511d99
z419cd27fff19d922392c6b503edfb95dd044f706e3611d3725a728d35c68804db74ae2df415a50
z79632badd0085b183f22dcf1f41c173b8ff06bdfc55ea062d9ef5c150216272229563a8cd353a9
z0b0f69b3f74e41c3cdcfb01e2ec814611b6e304a419ea3905d24c11d80c6ee38179651ece25364
z5c7f14b9c4adfdd3fac86a2a52ad54c99d96f29e6ca824c0c561633b2f27b3598d3f1b60673d07
z8951e6305139bb23554685b18ef8f53461d43a3ff7fcd794fd866933656bfef1558d48a558a7bd
z4ddd9f78f6a7d13703f19bbf28dfceea4095f86cc45f45b5931919fc56d7b3dbec5b4072ba6f3e
za32e4f96a19423dc511db98a0627d859c627ebff8546b0241631d5a416756d5d41f1e79f7efb0f
zde6acc798629fd219ff9a3f9f6658138c7c690aaaaf8c83af3357e71a37768872427d5660d7f44
z8df0ce0d9f714c81e3dff437b5e151fc79544724bb4ae4759afc6adc085b8175c4ce5853b11e3d
z95c0df9204c7e25291e767d690404141546c93549d3448fc284601e46f11a669827937c5cf2d8b
za7018de26e7b85d68d36ff387fb863a9270d486750ad6599e87c2ceea7a44cc5f5b1ab15e61508
zcf05b0c0396b595c66fea800bc96daf3e051693c8314673722427ad40ef479b73faaf160ea316b
za439f9a4e36d7eefa1d42ab744b597ca161321c9df114f3b06b32eb733b10ae2d5428c5af2866a
z9b3c8d5a840ec80b20cea8df53576b2ffa0a2454941ebb6be91e2cfcb54bb0d2282ced53319cd6
z0cf1f3602dbb7d6c7ddd52d11afa1c02ebbce559dfa42f41e0445ac543db0f16003486962347b7
z4ecf32e006353a2f9e53d688d050e6545c85f24cf4a34891e89dd11e346bc9b3378cd2b8ed2781
zb5e8d1f1859e04fca470e3a39f4de117a87e1703e92ab120c896ef11a7ab55d8a9cec871e1ec4b
z27b9fb8dcbaac1f3aeb54cf1f9ce6a5abd318f80d05fdf56b82771d844a5c27a0d852173a56d48
z8741f9226f55ad48827a6cee619691700bfc3acfc0af892b4614bb788597d1343b3ce9d927a655
z041a0e3a9dc803c796e3b7a55e0c02cd51438ddd271ff5bee220febcebabc31cb9acfe22757931
z6174e8db5a2bed3614d83110ad84b72154cdf6a012e608ffc848bec675b9adf7cc08d5369bb897
z70d54b3992e96572df9efd6c505d13892bf29ec8c178905d5bd5f16e9d61d025dc6c3f457c87f8
z4d46a9fe3183a99fbb2690ac179aa40a5b4c9a67e6422d9eaa6de2511f36dc874eb790d944779d
zf12a3964fec82e3f0b236afc661bc3f0ffb72f882ca9d967d923a1b881e1170240652ccb23fab9
zb2d10c75bde223956a3906a9f11ddcd522ba0aa2f1c530c7ff33623103e204f5bdd08c7e72be60
zc02a50200b60589997ea4f35c5e6472a8e6627f1591153cf9b8d3c2fa74b9b495f8bfd06c25db2
z2e09e5c279519dce32db29d15775dfef19261d7e8dbf82a9c3507be8c2906a7cddebad6d968311
z7f4f82c2256978baafc025042cd8f3d9395042ecb853accd4d62bd454a6eaf4e8d0df90f94fbc7
z27acd1514bfdbc8be351cd74599979d7b3acdf3ca1f9cd7d9e00efd9f57530cf37efd0966c69de
z5bdfa4c08af87f68dc61a24a58fd5611d9c9eec42df93c5bfbb937b40867dbc4ed1435fb2282d5
z04cfa060f35ee54eedff95b4fbc48a46ed1d671d9e2551824ad1f4a682e26fcaf2415ecebfe48a
z096421bfb5b7f1be4fac6d6c1c55decd00e372672b4bfb174ff23a13303df5931f1d128bfe26c8
z134dadd58491bc0e71519fb03a5c761b041822eb6b98574a3713fe3230d5ec7295fc86aae96173
z65b80a252f477238a795d29dc39b14e94758fdae779d781783106c19d0c074307d23a2d49965d6
z68a4db46028abfed10c882413b48ecf45ef52d99efb36a7ac522a61d40bd7e2024056990310452
za0ad1a28ed9ba7e0c44688bb463ed992802afb4d9de38adad3aeeafbaabe3ad859b9227143bbb9
z5aefae65c4e67bb376988df910f0c7cde806da0e573d90e905ff5e08ae643bb445f63b9d9b1fc2
z45eb325cb732525d01d22fe24e7c9038caba7f7eac3bb9d3b835fe22646be2385d2f0e070cd3c7
z8ee5831141f26c43da759c781edebfcc96197b7f440091a1299e36b084561e5084e01f17e061e5
zce271425e9e1c80cc58efd431ae2f49c88019ab9ddfd1699021998b1e66e4d50b14d3a1ae3de4e
zf9071406f0ae3007a8b54b1ce8d00e79f658f829426a3271653c08201ad3141cba8e393efd67f2
z9476bb8ec2cf396667d770a875da832319bc1a21d945dd6d28105151d19394d5522fe8feb2cb1e
z2fd263e991c644e965dca6bb53b1028344bb03739759fb67ba12118b5b9b92bb4af444ccd0a7fb
z46dea29da2be83ba91d77b3176b9cd2fb2e1701fe59b36efbabac3280aa066bcb39b4b9efb05e5
z4c1e9a16f2a70192aa006acae2946599e67fcbc2c98a3e91a0dcdd71639bf5c26314157ad2edab
z2ed7f8cba3e7dec04b4420c40d2a5371728775f33d0a6655649472c18a4bb0958f57cb5af69087
z8706c58c39e2211e1d3551524210bc14db2fe6f74d90bbe9a55383883be910a2060998544faeae
zae130c2539d823a14ccc1b2de423f9551457f46fcb428885116f87d8e689e252ad1b12b81055e7
zf6339fbd159630e4b0431bcceba788f55fce5107e48ec17bf3ba052dec6a5e1f2e92a794a3e54c
z61cfd8f3be79af906c255fe04ae435dfa7bd1aa962fbc735d9c600e7528f95e47f77dccfcefed3
z5c1464e4f601c0c0c909d229546dfbe3f84e856b33e59dd9941d47a9c4fae36ad177ac227f61a0
z54509724ca6cc83af0f7fc1046e9a4bb7aeaad1691541fe90ded1787fe6db11b192bf4eb5297d9
zdf828c388d26656a76ca3f492b871b65c62f3c25ec01b318c680fe1aa457f903d8b290d582d824
z4df197ad1d82bca8e83899d17df66cb8cdbdfba9e3c780ea4e5e9191ce240157af2066ccd7eb01
z45781d3d0db85f7b1e22263067a8f46494a5310fb8bf36bd61576a2b17083f273ae1c53cc88b75
zd0ab967afb9978e8814a800b587d833685e7a34a750845b689e7397bc82a51de67bbec6837705b
z2f5b69b8a72ec69ddbee885d06e0e81b191dfac5e96c98a15edbb34ec790d778ab190e1005444c
z01f5b8cc0bb6aa6caa98e5c4b72ec8ba430f09ebe77d126c91630ca73efbc3ae7de1cb5880a6ef
z5d86f47ff8eb9403eb8927c9fe7b6b9270baca6c019150bce70c399d8085e99f676540c352b6fd
z87936526f28821a5d4319efb63e3172478720405f8061c384f22162a7514ebab9d11b400513651
z4a60f973e633f6f13eec3e5a7cc91a3452bf19efabe65fe7bf7f222f976dca20956d8fcc10a965
zb75a97426a93f88fd38496028e434e606748a90cacb955d8a5ac08d394affbbcfde0c5dd4aab20
z4adbc2949c7208bf0bcf28a09b9f479b1057a5635d06749166c5435cf2d8193210173379e1d64b
z2e5a439919b7f026ce153824ff55d261cc8aeaea6450d8c96605c7113108e5ca84c3e5fee79429
z060b5b79cb95a96f6f42f3e6873fa210360bb2902ff67d3d92961d5a39ea331ec0a0b336d09d5f
z05a89777cdb01d2e39883a42fbb3047047bd74e0d2c414a4370e7d235ef13cf8f3336276ed4a96
z6c771acea8964b1e7dd5e481b53552b6ecbce5e1932f181bfe12786b07ebdf595e3253aca6c53c
z668d228baac2616670729cd924ab262f37fd214947fd91f8c986a49f8619cc35297d0ba08298aa
z63a9bf82794678fb15c634f2b987b450fa55abac52b1b9eb82917f362ba9c2662373b848ba8ef7
z70eb07627f82a98cb7d52d812778095d44d12a604d69d85ac314c1ed42b12fe8c4cef9940a5135
z5df59b41d59de43bec8de7469754509a328d927625ea6368582fef5cfa55a3879a571e76966d2d
z7f69c50ef296ca64fa1745168a24580139a7633b3a31e30b8182acb795402a8c896e047369e62d
z5537e0d61b0a66871589550490ad0633072fe153076f40c8ec28ca30dc19f7e2fb4d2a18d354b8
z49ed355659e0560c4d2e83130c79ad5a7346f0a6ffb1848ab822c02cee1800a13011ae01ac29a7
zf0586553f83b3c1f67d2b468d71bee1af89f85994c4a437d8f580f66ddb809c1ae38b247052c66
z4edb8bbd3055720af690cdf8ecbac5f6ef18397a2654ed586a3fa919a248167541d7e6fbfbbc91
z3e5f54c344ed3344732db8cc5dd78c33a82d6631147323f053797bb380a358169491286a40752c
zcf3856f166d6c55cc71bd74b534378f47182379cd5dfb676ec8a8cb56db39016d826341d938b26
z24166d6c73181d49e8ae6305ecf7cf21956bb4fea50c02332f8bbf8fe5cf8eda90b224130c0840
zbd1eb701dcc243be404140081de3e717207ab86630a9e0642887041950a34aee5bcd17f372e016
z65a8e3d4da5aaa27a8c056cc98ec6a947c968c92a7ebb8bd4342bb38ba22b83872fd4401a4b2ee
zb3111c59f77360d718fc0379cabc73098bb77da5abc571cffea1fe7ef27536cc62c92bbb43e046
z6192712075a932789c16b1cb90c7c6448fb73b34bc3d571662211a68c60df8815cce28fc9e44d3
z3ac86c611f5b4827074bc32acfd2f8c85844b70938b8e52f8d92bd83da1f69652f79dfae0caa71
z47c293cb875cea029a703a86d28106a60894f39448420225cf151ce47861fb354ca340b1e42e89
zcffc3cda78fd5a8272cc6d05f744dc809bd34bc6d2844777db83d3045b7e1480a8d75a278f8250
zd0d280e9025dcbab054d07cd5172c810329c401961da3bd919881b1c8109f9cfdcc101adc071c2
z10c18060ea1c99969f532edf646d44ab72432aca174c2b68096a14b91e2f81173c99c6d2751b1b
z06e3ddeac838b0f412597136faa5617a081dc0f8e2ef5f6d0f3339b40ee7f4a050cf434ba85ddb
z90286e59ff48b4723553246f42966e4a2c44a66b2a4401b84ca1ce82975b70b80ef033726a77a8
z181c9ae9409a6e2162273a704143ecf003397e995b5de89a32fa0c760cf4fcb97d88f266f8b1b9
za9886bfa3ed0a359e20112f11be435e58cc9eb2b8ccb2500ebfa9267dc7c8fc6c62674e738ef6a
za3b6b0348ffcb8926a369fff39c2cd5338ab382de2ebccfcd64f12c1d05bf6207440ab3811a7c9
zf058f1f0e37eb5013eab9cd396db4e26c9e0129a42fb00f568ebcfe1863a67b144b50fc623c9e3
z6b6186aaa97649dafbbbc097da81ee524a2216cff34d7447b2dc4220cc59887d1a92f15da6ccc9
z5492eeb0ae340ac396247030dfe2cbe33f9e230e12729e6388739c488a1d94dfca13738ec1ac98
z0ad08f31476b6bb3303d87683b1aea82bf41e6aa4c699349d6b74fe22b2331c98fa8ecc3fb8be3
ze49ae96c0ac9e15ca460aacca4b61150b208a106105f608e6352bae14ec301a862daa919e6dc4c
zee5e95431ae0d9aca78c61fc95b2562f40e5268a96a1bbd9fc5bdbf493b96cbce7a9301277b103
zb23251f4e327b2c9694e20ca4883d6ba0fc0dd1b8086229c8847df61169449239ea85587252776
z46184efa4d2f144c745931da1166aff78027be93e0fd6b1b3b90bcc21d9c7870f6029ab418cf77
z1c6301e08353c3f23e5fadfa70f96ebe5374f84eaec1d7b8b9daa6da84a59fb082897f28b4eb5a
z0e256dac5c36c8618cbcb683a4ec6ec7ddabbf584fe6fa0090c58a3d59207e467ab18142abe32b
z680201a5e462bd54c261f10e9e94b183b159cff3950b50e41edb12715e5f3b99e82b4b1f7c810c
z2ec28d2ffb1b5558e49351ec36674a0797538cbc3712fd472734550e2fa319b1e43d2e3d5813cf
z22ce2a61081b7805703693cd7d0c397266cc4bfb9f67a1f5135bfc87718c15db455d7fbbe76ebc
z70faf4692ec85f22a5ed56625c504400bf582da6c6d9aa247179ffc277da2d1a147811324bb8f1
ze06160dd61e5867fef037bc0067a77c33e9c1cf3fa619f7ea2a5ec4ea9792556c2d7f1ead41f19
zbc425c3823ddcc82c1df10e748a17fb7e93a8eef85f993d76d56d30af2dda70eb56feef5f8e3a4
z9ae57a2066f66f459de16c8b595bdabad0190f18cee15ba30f44e755294d38791c10b4c613482d
z591c4c9ed8f5fe44fb784fcf5444adbf7139da4bee1a729e450ddff3b681a7a1d3526d83830906
zf41c5b86d732933135b21b446731bea6ac64d1250df47350886a2dd0cb5db2d5a8fac452c25724
z6f51262b27081f41762c203ae10e9236a0ad371bbdacd2c6d192794a01596046aedec19dcdc331
zd274b151873faa0d47b15f89115b06ac0ab2eb68e88eba998ffd1e466a38d1eac2c6cf9d219eea
z9a02f672b91d8d4342d1e64aad8d9fba2e56249e650b1046e4447728ca487e25212171ea9e4847
zc68b1948b46d09ab76e4b4549596c402fbbdc057b631f4e45c92c40ae282d459ca85bc6598bc23
z045ca1b17482f792a9bac1d84bd29a95ec4db9c25221f29a08d7d25453a09955c723ad34c4fcb7
za2fd7437a9577e690d1b9db2ad480a8c804872221e7267d1dcc634a7443abbb4f5982ba04bf3ea
zc7bacaad8017c8aae5d0fca59bb1d0dae7b856e3dd40caac6fce5a0a55ffdd68ca815642df11b6
zefd91d7671a7d1e7c2167f779d3303882aa3523346e056f69828859361991941adeb4e3ab947f2
z92c17c3aca5f2fe835ee550d37dab3808c62cbcd7a76eb259cb92f6cac533f9b98942767ce6b02
ze8e94570faebd298d1c1541b373d107bd5c4a2665aa071af5da4866b7a555870ef1ad3f8221c08
z205374dc8d722d44be83b380bbd375c4c27c0374d30f11cc2d71b018d622cdc0b5ad86bca471ce
zd9b78edf878741a335b6ed54d5c51c78d2718fe6b71781e73f52d5cc6535a12415a4eb71b1d841
za9b7d6c3585cb84c495f2334d5479e81a65122f0977d2cee798f2318956a675346547cd15ae9fd
z47a3d90def1d0dede6ca6baaacf319a62955ad6604d4bd33008948e13ec5c119847afb34ed8e8a
z6dabd917ebbe7b5c05268fadb3c9237cbb7e1d7735ad71ae5f32f7a166eb05cbe83f2ec3075fe1
zc2b7f625137ef7177b3965334c346007100324831b9075cfa2637ccab5ac85cc74ee490284164e
za5975b5155a75e7c476d4fea8704407befe63a7465774810a14051bb846ef2c7fa945b94c72b9d
z77326f82920bd80c1b84c9db2ccbd685ea6c4e2037925c33e33ff864c21066c21f3a155112a0ad
z3260d899b80099b0fec2043e5d32a90a3110c9aca93e07e9b89accdc668134cf08b854bfd1fc14
zbcfa0fe6cd10c08344391b5ea7c8e3032489acdea95c7af581d0dc87ece6b9b53e07de2140a3b5
z0ecc3a48af861d5c5cf62c162ebd25623f1326139c099a84c09ef2b47ecb4bc7d4cb6e0f9cccee
z3df34b48015784a8eff747b3e7291645871b92006071d068c6f26e6a5b518d5144baa83e9fcbba
zd4214818b42773ec1ac01b7162868803a4c0960d68c6770870d8a4f504192ee772e75c89bff3b8
za3170aa0f0b55747831b90984f6d4c3b571909e19e56b2556a32643ed1bee80a2f8ec48058f4c2
z27bfe70b05fc6e9c2afd6d2d49ff1a1ed43c7a951ba589e5b060e4e1082dd8b1c7c11150ca67d3
z9df7a4ae31bd396a32a204b3834e9106c9ee7af328b27913f794f0cc6266b457fe0ad9d930822f
z5c5e9ce646952bbbaf7ebe10f4f45173299b6af845924cd82a1f3980d11c387b3f31504a5d2075
z53f61ef714d9e393de66f8e3ae2d3d230a961f644e18454d4109c3d516bed87d684a5777c8824e
z02604ffa6e5474cbb83d7eda73c53d5701df917107d28a5b11faccaa7a8c41124caaa836e5e531
zafbd9659959c79e13493d4f410dfa18d313fa17858cd00d176ce2cb23cfc080e669fa33ded800b
z5f6d532abc1dfb569955b4d10efce059b1090604a593f315afadc1e0434ca6af91f8135f69a2a1
z18cabf0de0f6d27aeb5757dfecc6f59507d9cda87919429be7f215984fe6d434e2c31a06f40a13
zb7dca044eabfd3da2ca894afe57fd9facfd91e50a90147389e79392745fa68fb7bf44ef72863bf
zacf61a81f0da909c9183c2b747aac8427cb3b92277308b1f9bd996ddc482978afbd605f5086b0e
z417c65e3a3c0462bd768e6ebe67887d2d2d1a7e53cd195622027126e396754c88a8cd131955c42
z77e6a517c8f89ec162c475258810a7ab33b6bb96f31267b9c5cf46b7c337569a2db8e21e034308
z9d09a29fe89b3ff6b04230888180d891d453837e10941cf1c26384e31f420dd847a1cfa53545fc
z8f2ffe23e8ef336d912acd1fb89e67c3d6a45058b53514f033699627a613f7f4cf6b4e2218970d
z68f4866266dcbf35bbff02a3e9dafe745f1439bfd45caa31f46817b3ed6df403e504a4f6806a74
zdfb0eb5da608e5191758ae246b335e76f70c81897aba89b1616b7ab8d1e84dbe1af13080968737
z794e4d5ac522b12794429eb69dcfa688e4e1f8e2a9392874b1685b33d0a58e0fd4751c32a8db9f
zdbfff24c59ef2e8013e892c30029a4ed94d9c7d2a4c7eef6ad9b31a739532ed0027316cf078d9c
z085aa2106ea0b47903622131fc28f3ea9a0d093573bc99ab875ffd5b36183719369db1fb30142c
z69178b17883e12cceabe9ed58dbbb81b9cdd18fbe26dbea4977b057ccc6dbf63dbbe864a7731f7
z7f3ce732917183d4d9dc187589911b8ccf972039ff5088d83fb4089d13a0686374234f1e7e573e
z993c834a8c453edb6d4608405f0c6b239382de125f255738e199a3e0efefd957cd38d9c74777e8
zc33b944be53d7e8bd5c9a01985cdc13d52a39b46de506eb1751a8cf80782282be7040c26a566f8
z5c1ec2216b5c3c45313a3b6cf057a7914bd70b52245eaaf37d5430d7e8614e4d4bb6dba9e86a4d
zf37357ab12e190f4e42d90cd1f5d85c5d91cb178136103ce17c55ecc13d92d3d3eb33687a1610e
z8c01657ff2f411e31cb679614da911a056e530a12b0190ed9012405215eddcf60bdf99e5d05d32
z64e94ed6a60e0486f95b86ec7f5a5f275e1798567ef236b4b413fcaf53489cf17098bb90753ded
z1000b099cdbe4fe5ee80543097cd8afb7ff8d62150b37c0b635851a27842c3287af25a6c344417
zc5c5aa04dedc0f3b50dee5f18701e1634e59e966eb4a5088b40b3a6c45518bc8b8b20a912fd5c1
z55dcffa42ffff0ea07c5208f2f242339f837a1169adead64f9df98ce845ea3baa862d862c9a048
zc559314370c6c4811691412bf4381d163e94b9d8a7a9c07e262e7cbdbf2db9ce382a8bcd10a193
ze717e76c27d4c6bcdcf335de157394c8c91dee3e3cdc9faa759e95f5a77a26d970b2a0bd9d5a59
z75be003b33697302627850e3807e87877cd2e868319b3747dcfa3b15cad5cfdf86ccbadb9c623f
z61db3e4ed91ae390de865c03fb677b8e4ebf5aa678ab1bafd79aaa1084a872d13aa39969a80cf5
z78be49e7128e7d87d8d0fd6a6332de0c44b7ed165f5fe83abec3cc67793db7fd7b717f17c8251e
zc8d72763ca3d21f6e103a9c481e03ec984df0e05e5b4e202973a31afd123b04fa0a5189744d2c5
zce26093abb7a57e51babd58611483c7f24c1439375c5e166b4bb18a4f615fda142c1e998de63ce
zfb231b6894af341d7421202958c416e11af1d683a45d76dfb03b3401fd9931a12339770ec7be85
z95627923ea3e0fe5d9fbd010b0eaf0a8091aae0e4571c640145cb1f9450e2b29ca432e318dc0be
z96bc3e7dc5144cdd96173ee6ef4f2e3eccf95b137eae4d46351bf3d1206ff715f70f34e2edced7
z6f91af2ac8c4dacd94669a3a2a65477db6a4126651ca16d656451c42ded6e1d6e8541b84dd4626
ze850e4bb6e7aca1b1045872ef38f7c6126e53b580c208a917980e09ffab1d34526226eab84d94d
z16398bcd2b36da5bbcc9211af06b849f45fb5cd29c98113f14beb021c41add089024f589b16162
z07a8f423f0567307cb2542d5cfbde9aa818813229b6c3a8728c91fca61e6c0b5d88bb08b21ab2c
z74401172c73ed31a26659f8859f8125961803ae7d7d1dea65e33a4a201a134b9c8602d318286eb
z93242cd043f278f0edf922e2ed5d01d4a75231695f68207cf729ad2c3bd75c85ccc1472ff20218
z01c019e222e95b45e5a17443a753349b356904ca7e89e8ce29bfd3e8674e5c73a5a61876496a32
zc8181a0a61e0423de03dd1916fe6a41f22290c985ed79f2471f463ba9bb70884c3237605ad79f0
z4412bcce9877a9c27f3cedd55f6a12f1b6efd4c6f03d0e08b6a6d62b55ba0a8d09977f2adda42f
zcb1d9db97877712e5dcfc3181312c77fd30f08bddcb9b538fee9b4be7f39cdec693f5a8413d541
z6bc5d328670cbefe18f250a2bc2f414525b7a01fb99f5b9695606fa04f029f2828d1c37a1b6ced
zb0d95f2a4149299744d444b743266755c5d790b847d5e0b87520fc8cbafc2bca54d1f1ca04d897
z0b398b8e21498a07c92d0b13f3d6a86ef4826da9feeb90ac758a22182d3dd3566d492724eaa4df
zcaf6bac1a3280f292faf5efef899b3b0aac3d562ccf2be3b5c6f820ff28faaf7e22bba47f5cd7f
zaabf8be8024c88eb3494ad3913ae6bf223b0e347ab1809ad26f24e4b12ad77a69e094d5f07f3b7
z83ecf48ff5951db7827d41b31d601d68a836f2e62c2c875bda575ccf8f946a039681d38583721a
z5f148da86f9da7c64a76c2d6db5f575827948f9d6c8296c6955a12b2d2e0e6f069f418343e6c69
z67d9bd32fad716a9fe1fd92fd1ebe803826cb747c7191ef51ba7c196aa1a37c5ae2089db21273d
z0f97d84029058a7a753901608363c1ea766a99b4af18aa0ed6a6806e53306e78d839c1aa13ba49
z4eb7356409d97cebd648d86ba14337a091aed1599524ac344471d14517fb6ee25143f0a3f53807
zf71016fe4bcefc3ccce3db9b3d0fc7fe9c61789f34598a2a361d288920918d27402e4c844cf68a
ze360ae871c7677858174da8185a4f4323fb85a3be1cd6bac75bd646f813c8ce89e7ee6d53a9fbb
za82bc1a25eae050f8941bd0d8a0e8928943b1446ecc99528d5576a7027f373ffa21f5650140f03
zc0b91511b313726470d3686f00c3714ace338087b9331586f6e70fbb0c7dceeaa8580fb3d3fdb2
z87eece9c631eef81ba4619b0c86ffea2af824a8f70af8f3f7a163efd146369dafad10b4e3627c3
z53a49e779874a878632ee2eed4066f2b767dff1f4c6b2fa80ac9f7f45f77aba47754495ce1b69e
z9f6a95933f7f3172a9afee445831d4ad24e320ae24b98b330f4abf4463be84af1f89732ad71358
za49121c98a525114c0166ca7b2667f0ac055cc25fe3c8bbf73b7031fdcfeb6cf61efd68f9cb236
z3d9aca73fbbfce647b42325caf3678a0f7e8f613c3adcd6e111d5bed80306954d08fd1c5d241c3
z1d61e59a5b5553476d6ba6691e59f862116864f2cc2919bef053ce9cec97fbba0403aefbbb3363
z1ea4ca081e960f1b04a6574f3ff3bcb1b6f6a4fdec3aede417a5fcbe1695e0f3649d803e447f4e
z43e20e98542bf50e3de84ac9eec4b3bce4b8eeebf26539f57250e3959bd798ef0f2daa48d313d1
z7ed6a8e1c31ea3b13e0a569ec9b1e9d5a1c69acdf0fed6925a8f3d7a19ebccd2e7b064a302b931
z5a4af99380c19f97cb42b70b6ce35546a840fa81ee06bc9440bd055148e661932ab8c0e302212c
zcea4f941db660dca590dcac1c4df6de63c02abe72a58e434c2ae24473980a499841207762357b5
z6d60a17f3ce7b93802debd2ed060091e976ba2fd11e1f1805b59e2fc689a2b151d13460b2ce669
zeceb252c4330a9a0a1f79514543aeead77f8c8580016ff2971bc461dbd4b1377dce8215dc91cbc
z36e3ec9b81e9433140017a7877efd9be4f59a8206e8a37103ff500b975584c3737c742a2257394
z7596d3448de61e12e46e45ea698fb88204201783a62b5d6c71b826e3737eda00089957c95c9136
z2664a05f4eb9ee175eab6bc0544611f9b9df121ebc8bfaab8b814b528b166118c3cb453b5498cc
za89c6839239a07e679a87bfe842ae930300c0614f1d5c173cd90d478327a595c7c15d02157db9a
z18f9eb7ffa494c105c312f6adba8724387ad15b24483e46b4525c023d2db3783ee98abc3ff44a9
z0a8d72a9a73d06229520f9291a03383448fa9697d783ae0f7ef479ceb8853013e1692578992100
ze6c1fa6ccf43d6f1271bc4213c8b91603cf12903f3883cd31e4a14602c25338d8e7fbf725eb44c
z7e78519114f127f14d030eb4ea750f3a315138022ee56fd25165e997f4433d02eb44af9f99becf
zf298e6b8daf879741d5b6f7a2b7af5adc14114d8d29144ab860f1442a117e687f3fdf67fdee052
zb43aa74700adb393a16378b66e06f480970c913d21318e031d75098226a068c8bb7d3a6d24a9cc
z0b3580723cce35f017bafcc354d31ed15cbd76f0fe221167bc646a6c8d87d3fd6c612923cd3251
ze18acf03a82df2fa1a2440e816dff7f7215e06cb8589efe5539e8dcae107585894a5e49d09dcfd
z64ccde7d62db56d2111d4ad56956c65877df341108b83cff342838d5fc98b5375d947acb224335
z5d62c858bc7421756e669028e3761ff1c9505ac816d13391a65cb77995ff705dbe6536f379f6fa
z1c3655c5a68ef453fe9bcb119f3ef9194b98ffb72fc35a988bb98f13393b5113c08309f5cb35ee
zb33081d7c77ced5618e8d4277643bf7ef0b6daf3cb69f9befcf3ad078e8dd5598799ecb33a367c
z9ec10aa62a505c565273e85bfbada357cbcd5bf3055c4c728905f65c2d07ee3b6f1759252635af
z46e7d3d001b37d67182f9aaf54e7da496e412846e49bc17e5eec9a3aa418f46777e49390b07e26
zc781c70706da4fcecedc8386727b32d94e20c18141be443c70403266108fbfb61d7a5dea767a5e
z89c8eebaaa73811485a646f8bbd1dd9eeeea5eb41d03b3746195ed760fe39ad8196eeb9d0dcee3
z2fd092629033f349a38bc54f07a3a0dcdc6b1acaee69ae4a158d2273ce709882fff7a141eb914b
z56255de0f797c0f782c89fc1dde3ad03e1c8b1ba80ab16342bf16cf9e0fd080509b151707dd229
zf7368a94c388d5424fb11eda5d794fdecb3030675c5aabf662c76ff3f8dc1430322a26407f1760
z3513a531fbe946565e827ca327d4a736d0c6662f0360915c57a80210182af63ffe757c0f381e0e
z6c9470a70109a8ad70bc4993dd9f506fb105eb5ef582793542a3c099e2131716562ccd8ed394c9
z21022e39b81e5008b964a80f02c815573ba4a3f0cefb95c3694aa16193aea78d164391017c0867
z5557a75770522671037d8ad963ca0c05c7be7a4715d0daece8a43bd3897473e02fe32b2032452b
zc51e5c931137965b906b2c29bccc380e14f50e61bf9f25d4716a30acfa571aac4620c2cf5fbd3d
z9babf49a20fb1190f32dd9bdd3f1e0a0c1171ebdccd4ab66367c59d49386e0a8ecaff7b2e8d346
zf8264bb502c1acc7f07a065a262afda7736fc9dc4011d4b412f402ca3528858b73d5db575bb1fb
z6c2b437d1acc8c4a93cfce18128ed5fdec4c18ce64a95107543c5aa6e5d05e3a18752406834168
z4f544943c403a308546eb7f4907a05e3bc7b934b82ff10fb1dea202bc75a32b7c8bfe3a173cee9
z84c22f9a9cda412467016b65b05f1c2020ac67ce846af4d1937fe4f7bfdfebb41dacff6843690a
z782b6f50ba9726dce10af9bcee08eb1ab5e0caf8bfd7785206d90a34d700172c1a17f6594172e1
z16b2229e3cc393e96e2d34c94ee086f517934888631734848716ff0166df83d4c60999b826cda1
z151b00757115e86bdb419c8d11addd68888b52c40ee8ea84af0fd6ace2ebf24ceb32d38a7b7e1b
ze3151ab2a0b39f95baa09ce85d8b3464797c189be09987b38d402ff9a7286bde955f28c255b154
z67daf48dc5c1560ac0aff5185e6c0c06cec22690b10e08613718eceb133eda3accfe92923ea13b
zdabc8b911f28d0736fa98417ca0aa4fee328b9e624abcdaf16c0ff9e865d964ecc81b39129e8f2
z1072b6f5d0604a6d52b0f68e0b27758b31e1343e79634a1d9634be3504f97058d96749f83e27c5
z375ac034e1da3f93d7213a8112bdc4636577fdf5e9f0330d2de52141d4d30cac92fc224f782f82
zf99efbb348efc14e8482ecd7333568f301718c8ff784c79a0993294e70313a23e02c018c4a9ff9
ze47a51e090708bb782e963e53bcd7c56377c8eda6bc4daadf216741ee1e311970db421c6fabd7e
z95dcb2cef21ee0e5085f930f86711b0dc8bcf8e5e71f9a302a97417dd99b998a0bc635d504d413
zce6d4f98fccb68e841cb6a26aec08e2d6403fa3fce3acef944b64c828fb0fd26b99477929ca7db
zab8e64ac0adc2288d5b1bc0f3fd62386bacf053b5aa21c3f9d7e478c42fb68c8688e2abb362e4e
zd6838922e8c1f10057654e52d2b4b65118ee0a71a887c4b715c933988759e5f48f22311cae9a16
z97c1e258f6c3ee69551d76da06b4211d2f4db2707d2b02e1c52b8c29b550a943ac76b61977bc1f
z8f015fef773e92b989f3b50dc920dedd40d83a94d9bcfff82187bb8aef5eeebfae7fa0f69cb77e
z8549575b8f047d50b1cf6b56455017fd0a0c109ba4759d34f6c34992c56344d52f73a9c6d62fea
zdf5ee0fa924a4d9a47ecb915f08d710960e63f3ac0e6cd0dab0fbd4f675b9c3e6e14b5af6ccaee
z7669adad2435439a6ba4ebacc4c60ba4848b49be76dbec6a455c8b66d7f9e597931b53bdfafca5
zf1a81d4b7336dec61282e5ecad069c9f9aa70eaa7f5b61b4a6f7ea0b0440ed231517b4089e34ae
z449d4956111c5e22a331054f26d04fcf2baf2acdd00f818f8f474748d77c0c822218bd0704baab
z4eecbd8514376db8d06313128c0d8e9eac60b66289a917ebc4d73c65dc524c3cbfd3b79fbdfc04
ze482f58655f57751b8316ae0439b166be8a3353c0dae83f9b4029adc8650ef20d9affce88c3a01
ze55beefc730096f6e4921e7b3583cde126533172e80e63f62c502adaec5ad7db07997cff8b0557
z056e61d70fa5e030ddbec0f2b1b46585b7e1ed614f1545e79bc1e79dfedfbed0fb99e92671a49c
za81d54addfed86f6094e197a402c4ce229f3e59717f792812f0b4e86c603220374e3354f84c4e8
z9634bae1dd953e9dea2f5ff8a3aaa0e0a1d85750b0f9a7bd21407e85d55cdc06b15b3442ce0f6e
z1683b1ea5fccd222447a37025d9395e116c3432c3d9aba733d4198f321b29a0155b757251cbbdc
zb0529b036f4c23e13f9ac41bec57f2ab9592f8cb128f3ef60f9333e44a400a21d3433ab5f70f09
zef51edb72243e919145733fb8eef57b0049b762d23c8960a8c124b6f5b9897dd6d61e8dc5ac0d3
zf955892de24ae473cf9980cd2274961eb521cc7d4570ed5b66dfb3bde75b3dcc7e7266e1f1fb22
z373897a03e10fc4c2aee6a28b2a39839443ea62e6c470934ed3b1e95d4fd09d53129e9c169e396
z2883fe4095e47c4d7c3ded4d37c5c4645ff2e6f37b9e8799b155f98b7601ff2df9ddd5d08e1bec
zf26738641ca83c275ca9d718f8b2ffb9736d7c7f7dbb2fb9e56fb114dc149d3cd35a8265c20f73
zc588837c4472ed8fa8c5f2a28d09312bca48de2479ea2793b978b627b67ed2cde68277ed724c1a
zd77e9ebc1293f0dd5f4a15a976a26a4863064ed4b0955406a26a0ba8450eacce9dd551b40b237c
zc46d9168f5de7541cf39e62be0428c1e8047eca1fa2796dc0bfa3b85a12239f03be478fa9fe8ea
za47bf464e67483ab0127a92fd5b921dad03b248679029b448048e6da816ad924cf9539fde251ac
zc031d7e3eb8099834e82ff4318c906b08bea9316e52bbbe6a155e424b5ac2d9d125935f6cc2c83
z2b43a75d827d3976c9d76c754fadf8ab1108298a1a325cfe052cf30a00bbc2c35f2d91621ff6f6
zc1e4ba5cee5515dcda90c2aea93f1de782dd90c5cc2a54383b4e2f06d5013ac07948f44f5de4fd
zc35e7344bc22b9a4c6d6d52252d18bdeba5dd53b1e3bcea0c136ba2148bf47b58937477c5f9eec
zec57971d1441a72f125c6a52bce81eae3ee1d2ee33f51001fa355762c4d220ca88d8cd3417f056
zee519f2eaeb2eddad8e72059c59207a75497396c9e4cb979a933bf4ad1d57872d2993318be42ef
z139502abd9431547fa667081550b20d485151c3c11e6f265b5924a6976efa227d6d03fb28e1fed
zd55ecd9d2e8d987d8ef47a84f67457ab727eb34a00adee15465b66e6f572066b918e7a9724ed69
z0a631edd95e93cd68f2afb37d31fd2f8a3aaff32a06618ff329641f24b3b27f4a27873913866ed
zae0123f9919a64c62d450f08aeef9db4f1525dd8d08212c091f10c2a77a7f044f39dab002c24e7
zf250927324218711610ac29a81be5a8f7b24e50e1c174f450c4b999a02de8c9b78f20870d610c1
z8a8e07cb90abdba971ca930065f347b036adb1bd3d2695f783fd8ce782fde154ae10eec601fc62
z524542b213e667ae6d8d29ddcc0bcaacaab1081c574dd3de0c257506c543057fdaaddc5f50ce34
z6b18aa207369f2cecc5b83f05bb1d7a549a8ddae17543d85e0b62ad51227bc337a8e80d956b480
z5c8397b71a3de76d6dca7ac47f231a111a66e27d6e7878177ebf157500e6fd123641a381b1742f
z0307f764e0461f5752ec1cba01a0561d12d2b7f53adc2ade39fe6b9d1623d71b0a3a8b071d9aa6
z924df3690c687e79c449ababe26d4b44e7dbcbcd1c370854a4db015fcf79fbf5f02da2d8ce4348
z73079f655536a9e69d075057196799559113054d5202c67f098a0ce6876f5cfda960ca0cfdb966
ze6579ff9aefeb1b736618c16bcc31dfd160f5b00aa7960073b808431aad3b0a63c537423466000
z6ebc0fe35fac77c1fafebfcf747db933ceba0f49ba78157b5e915c6793189237fd8bce8262a8bd
z9d7cbf3dbc60a303607f09e0f901310c2a4f86d2b1381e3c2657c99ccdfb4823c1669d0028cfc3
z0a9065894a37a02a5c1ddaab3616975e6591bcea1f5ae8c391f98a5b892a26afd9fcebc52c2f6e
z8693a948c68b2e7517c46ee034866f7aec71654251c31ea9c8e87274e1362f50190f554bce209f
z6e04930916e434fc3607ac01ef0b5a0d9459f5f5ad913db0ca9c951b1d8c00efdae890fac7df21
zcf1f75324a1badc21521ba8b1e078d3d1b6ed848883a193f3b1275d29ee53b4eb7a298a14e2fc9
z5de5494b8a5c215ac2a33ae83acf4adeab61d0b474d4edd291c150e7fc547333ff1773f395d381
zfcbdadc63aff8fbddcd5cbe3f88da25279c60b48cda159500a8fc43ae60aaaeb2ecfc5862de992
z40f578bca6cee1a3bfa5c7a5805477585a8f4d8cb6c29a20bba3d598dc472799ec029b4b3aabfe
zac8a83f50cffb8ec1fe29a15ffe53a25666326417db1d03b7bb629edf831cc7ad219fa45f6c978
z4a370f0fe6324940046cb40430ddd2071e497fa26ae4ff8ba0314112535169ef0530200f0f46de
ze3e5514e40d2c4f3504938ac140d76b5fef6e1753d8b744b60be75bd603c38ec129bfa92a370d2
zbc972fe94703dd51506a6a8ecdd12a7979e9b3571caf6766817cb5730f2edc31ad018c9ef8a567
z0e6b3a12890f12713d966209ea043f27fe9e10958d445ea6149cbfd2bf93ca17229a2533aaebbb
z8fe301f2b3ed71470589743fa4ef975a8bee53ae0b124c5682aa17621dccb8502cb9fab56295f2
zdc12234c61e5119f243a53f667330237cea2196bca92c53c4ddedd649ddda0d92eeada970502b9
z3b44c8c09e27dfb496b2c0b7cbaca9a41ed40a522597c4d15ad205dd11925de16f316611af5fe8
z55a53f8fb0782dc424b96016f1e7db4b6db835d0651fef01b10927558c465f12bf6f9600e3d29e
z3856b4d729e73e7c258d3c45546e38de853b87d6d30f87d7191223eee5ad10bd419ee119c895a3
z1bd22864fdc685dd521662354beb1f84939c603b2ae0ce7b0daa12608bdcf586a18db97c3b57af
za70aed44dd9efa909648c060fee0cb0b82d8fcac03ad2d3eedf6721e40b91fbb904f6eca2a9cb1
ze5ee5641e931072337e344b9b598c62171e3e37fa9f1a10d9ae5199d201a3f60a0ce3ee07fd420
zae40dfdbf2ed3ab8bd9a04e0d4140ae16319f7db435ed6d32356df006234822ce81c0b56755c35
zd94a00e4bd07405c62af117c944560ec11c107208cf2eeadc850b16b951652d4a385ebd7f4634d
z6c9f106e50104bed9bd1e7ab05a670bf652ed095acc64a9eb0767149cfe0fad937ed86ba6f412a
z15808a4c4753bf26cfd22d0c142e8e47462463bb28a9e69f00c8edaa0d03be3ddf973df713711f
z40f47b932c2e4a1fd5ec4bb9d7a1ff2ad3bb5ae00ccb0aed0b1612b856a806b4566d6a162ab895
z2cf5cbb0271cb33dca973e9336807d64cc4626dbc5d701d6b07374b987e4de9fcae4de76708a66
za21e84b7c9f1d3ce9a8b30a46b3bfcbec47513631ac0e5813eca5adf40c3f53c9d406023b07b6f
z624148a86d888ab4bb37e4f4971bbd07e150dc006e9404c691c3fc8f5d486bef57a7042424adcd
z65205585ccc2c167269b1faf886cfd373ddaf7d82dd66ea75b52cb34c171b9a120109fb67683a2
z8f31abd05b770c751d43155683e583acffc0af9e3917540d89149c403fc3e21e71d2b501ca0ea4
z12465cc9f9fed89ab9c7daf6dd6e6ed64db15b5d4009b4ce60b40f2db6fb3f339cf3fe1cbc341a
z27bace1c6dd9ebc4a27d4b60ad6549bc81cd664664b94d57b1b63f10830814d7dda1c517710691
za355159f0b11cdf9c866e1a5d1e6dd8c91a126f14d05aabecb10c52b4a6eeb39ff1d38e8690ea6
z11aba8e2eff16cbbe707b8a2f593423d24db2cc34d3320b9014ad7a4e00a082cb247333cdbe8d3
z96ac3a627cc484d0e2fa4d5cbdd31311c8aea352ea9897adda6927a2f8d85915e7d3c465bc7cbd
z19620b8dcb4c63d02e77ae3f6af06b89b177959243aeda5b5cf210316c88722d3655c890f25c0d
z8e2bc5608a7833130256b9f9e3b4a086d0fa42fd9eb15ef4b077a973c73f42622b90d4b25343ab
zf7eb598b10642bce3bcde1ad64331507d6b354739068bbc3d454fdddf7641f76aaac252c11cdd6
z22dce3b33ef0d197cdc6282d96ce2ed896864fa69d862b20340409af5b62b4a101b7ec192e0871
z2877193754e5fdc24428075f6f31d865add99f5d9377ca65c7680336837b96fd1f42d6b9ca691f
zb6e5af31b6f3bfddaba2a9b995b196bf4cda607696578829a1bafb4b57f7a045f178c309a49b91
zd5e6c0aaee0b822ce55345edb0b819aa3f2ca20cbc39eb81370a332782093a3b4b991c8ac791ca
zd6f435477c14c3ef6ecf565627317510c1196646daadccf71513a6842c43e801cf1d0b718bbd5e
z24f6e17de9602944e2b2847adde5ebb520bf1bdefca8b16eed7868a8b1b09c4f68942306adf671
z1b385ea9429895caa0b76dd90f11e6886d734a9950bac79dc39a88ad232078419363ab52e7f038
zd15de89858e44625b0c24de72c98702282110bf1392273195d955499cabfb644a4159236875719
z5d7843a3400c05ec6de8f859e0075a8658a37cb1fe31715e476f1696d161e35911c71f007b9d61
z8a637bab69a0da6f6818f3429f0fb1f1f1d6002e043b009ae7cc3dfd402098ab7cc2435ecf03fb
z43d51057ebf6446fd0452a376ff1831b67ce051ab17f1bcc71d8ec68b1d0aba7607c55c09cd5d8
zfdb15dcf99a31d9148658389fead113af351d3e2c95ee0b4e3244e569bd8e2d64ef1ad20c8f9c4
zbc9e1deb53790881276f5540c1cbfb53833de4dbd6427103a45708da1f020c6c5a385aad1f8aa7
z3ebbe6abdf27ae5e47a5045fa869824ef1ce9c43061f39bd78dc3efaef84d830767d60b4215e6b
z90c612592a0052d16a843245df5c81aafe496ef7ec6ca007fe3064f011c9ba210f99e7971674d6
za415219c67f79948343609a7460a55e0e52c49f609db84afbad1fc30abae7c082169b84e7aa2b1
z3ee14dccd8c39189f5b2ac4f21c708fbf497c5b78551a7dde9ec1eddb48312dd9b31fcb3f69ec9
z9b92f085adb17e9174f86c1dc5f9fe85452dd49b0916d789c3683d80c050932e160da0c4cc8df1
z60aa41cfde18af41bfe7bb2cbb7a2e017ee1ae0d5d18f6523123bcb40208fd6d38ec16f0c6f5a8
z59fc0648681b68b5f3f8cb6e1aac33b14a12c596cb08da8af02f331d09d7a8d7fd5a86341b0ffb
ze4a6ff0631794a0f780aa675ab3fcd61d68d0a7ffc59f69fff6e04c481774c25b1c254f1f8df6c
zf94f38ee5f0ba8d292fb40b767ddd9bea6c8462d7d514e5da5a1dd88e3bb8f295e947e1c7a0447
z4611b46bc6b30b099a3d8809a71cd9965d6b0e640fb57f8a295b7748a7c55dc90524b503285743
z2c8c8057faf7b019545113c7b735f156618ffae0ca6497b04f693a38adde57311829653e4e1d2a
z6cf81493ae19fcd706adee392334bc2629d63e831c8cac935b6cfbf2a83bcfc1cfeaf3ac3c99cd
z3ac68a5bd06e144a09ed7c5b965e1a4fc8f6ed68334f31fd1ce3f97ed7efb32303e687e63f5bac
z638a27fba2fbb4ac0422be26b4e5dec2e48369e50028e4045ac7d15ca56c106580e77eda43742e
ze3da56c539445794d25f229c8101f59e48873bd384f54bab9276463319528c9767048f2c7ce7d4
z72e41b8e2a575021432a38ad944af1407156c2b783385fdbeab9b3bd5c47395b1d9778753999c8
za83edc736f17ced0ef2784a5900f6d1ed4470a57e93f8cda4615a6fd1d276c4524c3fbc38ad73a
z5059741e6fe8ae531022262f88aacd6db227bb7121415dc389ceee553c34654b4aa89026b18aa9
z20fad86abce300086e900a21ccda7babd707287b0c24301c55d0fdb331559184b7b35b2f1c37f8
z14c26b57651845c60ece9073449aa342a10e98d6cced3fa714f64c9f1ffc99022a3bd26d0bfb14
zc9a8dcef432b6f7cf7ed03f3997cfc827b982322a76e106ec49829bc400276c3b19ea649839179
z5f877c4caec1f25022b9da0181c7e54b7cc96a1c02847b62f93e15f4ee988dfea9162d27da880c
z60bc6f187af92c53ecccf7680f59bd15086a1544b7bc8f19f44b9c1c5d46247e1beb7c2e902234
zfbc73ff409e1af785f5bfd796109b373ea5b8d821efbf1d778ba497f67ea64f2c460f798db0acf
zb101236d2f1b10f2e4ab3cc79c9d64ec6db285e3eeb71f21cba823d8ca30b37f1bc745fc4764f0
z899e7246d9fa02828a79a664aedac1c15b940a21b56690791ef400683e0734484a53726bbd675b
z82ca137040e84f602e614851a6d1056128539abf9e5c541cdaa9cd693f71c44fea120b0a76f63c
z38c65c402b41c69c381b97b821eb0a1fb7e3769bbfa2c9a66a0173d06bf6c4bb14b258a5d4254e
z2b0d2cd9d79142d79fe29bd89b72eab9e017b290f15bd9175f8460b32faf2de6bef0dc8cb0ea4c
z6dc3571b3e1963a139005ea1d311cc948c71a731a8e7d3b4b02462f3180b9162625b406603e37f
z1e1f66898c720e9a84599f737abedc20ad6372ce9640e49f6936ed53cf530bfec7fce96a6cbabd
ze3afb65fcb693852efa37ca786e330ccca44b04cc493b4d88c712d00abe8d0eab4b7af470ae615
z981c582d1b5b3d1cfd20333e14af13a2e8929ea8f6bf34f622fee9a7f6cdfa778834130a963c50
zccbe1379f317bafa7248574f8623aac3f41c7ee6805cb6abaf6750110dcff1051befbdf818e283
z2a87a7fcbeca19ce01f8207c69bc4bf42c377c6d15869f3074b4c039e9bbf2d93a25d5e708a4bc
z2cf27896b0bdad380129a03a6ab23785eac4a65debf7fd8904bd014513b9d337599c399b0f2fb8
z82feefb3e38b398d601e6c6b0b314082f696d9089dc77817162180f13fa5b4ec0a85705de31cb4
ze9de563c3ef16871f9327b28397dbe3cdbce432d2975bd95a7734b53efdbac9cc703f2fe6bdd75
zabe71d502b8039d3618e64178cf5bdf5e22bde03e6174382f51062206aaf675bf02cbaf9d6d215
zdb9af8809280bef0a61e1ab8eb5e0d4d61a345af3a3369f79cb13fb039a80fcae6c4689334ec66
zf92e5ddd5da9161aea87841098c806ca23711bc7d956e9429c6e23f58ab8de3ab6dfcd4c4db022
z27accb9a3f4303f060eedebf13bd12448295ae49bd73b14bd370838553c2b7d5c857dee27f28ca
zea9544c83ecfb6d9fc86ba56c1fb3cabb22713b270daae5447b367cd1b4ff0966bf68862adfaa5
z3be1a4c6639522250741fc7eede7ffdeb0d2d54b54a66489d40888a184f6d34523c99961b18c69
z87552289b5a13ee7a66ed275fb6d811225d4ca9cafb772311f9aacc9447cf6f9c99b597ec8f9b0
za77d90e2fb829c50ea1743d889fad82b482e44c13c0ffd25fffc713599484971aeaeb87600842a
zfbfd2bae8e95156775904efade98a753f1dd1eb3926b3b99ed70b9ade7f3d1ebbbb442b475c11d
zfa0b18e6f25ce1d419fc91cc68d5ab574f677055fb1ee018277ac282433b5ce8cc92e3f1e79b7f
z1c29160419de586b17edd0ca5f5f0a45dae228245fec146f0639f63e0a6f120c60063ec286f973
zf4f38405ec8bf7ae2a7db95817f740c381150fbbc5f0fcde97a3a55282b5b7098edfb84d95cac1
ze56927820c8cdadadc93ce278117739177e7aadfbb247e04c93c204277f3a16500624b96c232f3
z136b85a50c7f9ed5f596a354d572d5db27872f230d381388a7c10d9f4b8669895d538a53ef2f73
zcc41aa7d1d52458d5445a6b9e339b5e5e6571893aeb04380686f7ac8ec308d636b1ed8f1d8a50a
z356272f2791aa94083339e4eefa81cec04610ef04578293654d704af39601ef20f518938ccd5b3
z5ec6700ad6ee6e4b8f46a95f62fe0a25977bc4c7c97641da18b2dcc77615ae31ae8d5b57566d5c
z4eccd74ae7b0be664819eb8addea4a4cbafa381ecc87c83e976b51bf93aa37d57e2523a5efb401
z5af02ef8a3e93987842aaf5fc28b040d6c16a5709fd05f9419c800d4d26233df4e3c7ef5652733
ze8ee8f57fa6a40f9227c3f88cb1c6421d96b844f0f084a31e81036a09081b61d3df4107ac8b91d
z7ded928e62988fea139710eae839d49cb03484348741a7ebc75e3dadc553e402b8cfa585027ca1
z497fb22c9b73abbc365f5223969b1af5f70fd998f36f8c745ba4df18612589e264f971074ca953
z5d6bbd48f408f94d544fcef338683f3486d20b1c13431d252f8ce1ae24857a18ae6802bf1b309d
z306f0ec87608f0afa5dbeb36cd54205f7189cc97492ea7ab7cf3a0f3ff78dd9a0c5b5aedbeee49
zf4058811beb478f0f478bf6de0acfa262a521229f46c11042255f0ae9f327d843e8f92a1502ea2
ze5034801399d564cec69e19d8dcf5a24de7f452721d36dd77619f7f4c57facf7109e616babedd0
zd6a927cf783fb5ee7ab8481017016efe1a7c9a2cd1474037e80b0b4a6c5a54b126979724e6125a
zfe97289051ef850a450f3d619d06c909a0de38b3e52bd475ee2569c361feb9f07605338e4fd32d
zc8a91dc9678fb315fece6fe88b3bb0e80d4f83acec1a6120ae8afbf53138150179d34d09d187e9
ze0463982f5be4dd53c89c621e3c9ea499fe6c61e0d934f6a641dad322ac2e628676ccb10a06dcf
za2714e8ec6df3f2ea7dfd369ab82e444425d8d449da8390fa086f97488db32415257e83dce7ac8
z80489bc55d3e658c00a3c4fb95560a68d73301eecbafd6d2953c1f05e1512ff9de3c57b4c0f8fb
zf0488b4034bb32a73ee219371bca05449068d98d42ebcea8e831e7947e5d5968097887bc74e2ae
z4922d25fbf5abe3452aad29f323e2eee088638726c2d47faf33f46886402c579af6f4d1473366f
z1f2ff3ecda40cf0fcb985e564afd463855fd20defe82a82e12b228caa0de52a39fd369863c2048
z45cafaf7b3d0bcf1e085ef3c5af7d1e866336130d731cda7fc11238c7a91670a4f054b9f6cecea
z16adddbb60556024fcd18195fc30831267e50d2da1365877c78e4ac9f4f71c9fc24bb9b61665f9
z464bd3a8dcab888706593dbbe735a13c8584f6aa1c6dc80e49b31e3e52c246c3792f6812c08c69
z75684772b8bf1ccd2502468c12f6e82461070da0b4e8d14f9faefd16685e178d53425579e5d66a
zf7873d88c1a69c140c4002a0be90c88acec22f702db4ffeb6ec101e86b97b3d51220b5fb77f161
z7abf9bde2d9c6d813a180dbb69c07f9388f940a0b6a6cfd7b724f603eb28c853b904809cd689a3
z535a9c88bbe19925f09bfe794ca17934d2f6e7c9a1db4dafceca2db7e754965be56c51d4f281c9
z2b909fb15823582e97cd052121b68dec5c07136b01d29eb36a4b839afaf93f34e1a60fed5a39c9
z03d2ad808faa88e3c13370058023677e413f1b3c55f27a7f441e02e8bea9791bf47f8a0c65f76f
zb95f66b91abef0eae8db991d9be82b6092b9921dba59f9dd7746bff80ec9f446d42368e8d48381
z9c99b583160e88d3bf9372fa32aa09fc8085d94a9033efcc191d933f00f8d739183c82d31003f5
z2dd65afc7e34c2fea7a2455676b795bb4e2ab6487bf93d50b8ffab6d7b3e24ce6f97f789a25b8c
zc0c530b028aaaf71387f729a30b1eff158189b246cb1b71aac260828731c24dffad507ba5fb87c
zb833b8784312667fdbc9dae40b926d8f7d019e20935f3712806cc199d937f19879826babff788e
za6ddad4fd8be5bdd14dc86267d7032cf81d03648b343ace741d729627dfef4e8b6f9a3415e563a
zcba30f4a091201860224c101ded9830b22a419aa2ac0c326a9f401f57d072fc6dcbc233f1cba18
z83be5061d501c44c194753aa8b50c4311f6d72c740c6b162d56dca74d95491c9a7f441783d48e0
z209c47f695bf6432b893567245485b4e1bcddff15f1e93b6442383ec89e88c35eb3fbc6405635e
z42837c5587e0d90889a13a6a63fd704353f1d27579d2d31152eb540a5c53e704abab07d8c41fc2
zbad627772f57eb96ae5772a1b21d48e4571d72642849aee2a4313fbaeecf41b889678499683ce7
z742980fa714bcb49e505fb14254d9a151a33c678d4be9f608bf42bd823704ea3199405229843c9
zffe511d1e6a68a697bc75fbce8440417ca35082703fcf37311b7bae0275f5a2e454b485dd86eab
z83af4284f7d1e59fcf00bb9e3e5b1ed685c76113cb20ee74c3a0ff54c6ed2ba666deb53e7fdc62
zae80ffb062570597871d6cc5b600bc56746c67c8512e48442d1811bd1764300dc3cf6901eb5984
zee21b9ffaae3cccb2cc978707c30b36384101af765288abb41fda49b1a176f47f6a7d2c13547c1
zeb0f3df0eda2b6aa4b1e2868860a0a1429efae57fc4dc397eca003b2bb21f13e784d5f9e193726
z6982e94f68c4ca39d38fb10ec3aed9408a9313898ae0c5c461abf16b2bb23d93b34bca4be6bd95
zab39bac6de23dcd2a32cd500ddaaaefb892ec6efead624097ecef433f96bf464b804fce735bf9d
z60a0c0688916a6fa4ae00d1699f30805592a300f1aac313893b1229c79e871b68b59d5558ee429
zf3c0355e8b62e2f4921d8c7079222befb3ddcf87595b6907ea47fcb77ecb0fe6ced6bc39c263d8
z2b8790c5ce747ad6f991ec7a635c68956aa348eb57aa352f5bf415593c2d6a9ef205c0741f6ead
z68ec11520bb5f6bb785c2f341de478ae941648f98a3b585f9acdbaa4b50743c76a99968d41607e
z3f76b4a58bdb90ad762e909bfc3860fd417dd8c74a3fff6885dfe8e7add6d15476df654df051f2
zac504401ed7dbb5a055ac32668bbc681d05cdbae954f4bedbafffc542eff882b978f240affc66d
z97797a6eab3b0b3caa3c6529b141861b2490bbe8de7991fbd7e5455348ffd2dd6128cc6396627b
z96b086efa9560055311bcb5d2ec0cf7644dda634df1f0ccf8737419eac8ac15c2b8b0a79d7df59
zc319be5d228b3dfa7f6ecda7506ab9a352bb2686327f88567a0fc25ae457a6e58f55a244420e03
z8ebfb67f6560e7b9f96d508f8e04d86397ef36b34de13a92178014e653749eb0d73dce3f3b8942
za6ceaba5600784e2c95c9dd393167c9321abd3bded21d9645bd94f3b5dfe523aff683bbb35af51
z90ccc23c9a4f0e4b9b81a3991f0acd3a847f007c1d93d8082207f17a831d3274806ab859a85da4
zdbc460d22bbfbaf5a161ba291121dd417d4de1681e03668631294900dfd38fd10ca7f3ebc8baaa
zd19dc817caab8a14acfba90dbe8c3e120dd82b8fce10033a51d529c92e6edaa829f9a956d50fac
z395ede56f544a5139db7a5d8db07c0469d32236673df20c235486cdc8fe7932e31e48791968976
z3882161f35328a4b482bd1e91439a1d52716023c5cb99dc5ad81a57dc32c8800b753f355e94f9c
z5e816900ab1b482a6d2dfcd9e6a44ef9f550c6edd423bfd0f94f241bda8f87f3580654632458cf
z73941e4ad518de4220881dff26b92e6a4be1e507447e88cd806488bb61e6074a943bfb52506a30
ze233809be0fb973ca845b32ce7276e0dcfc50bfb2f8a25de9dc7cc9c84f2d83032d33e19e1ac98
zf191f2f0d4f3ac7c65cef0c5fd4df81a65ec59ba34f65901f50d8a116da57411fbfd2a097a96ce
z1f8617e8c2a09a233a34c6e2b85e699ec7d860688b5301ab98196c85d4c53106dcd2fea1b811e2
z124719eefce77296c9092ae7b2421b07a9759c8812f35771ed1ac76085d968185782e224415488
z5dea3a3649136a580b79ca1ce673ac9fc303e16056b018e6ca10ce54124336c9c50fc58fe35427
z1abd0ce7dd22f3e672da288d48376a454396c24eb04b0dd5cf75b91b20aac6a0d3e44d2a7f3fc9
za8c20c6d25481465ffb484be2574885ef9643641ef76c58d75fd414fe0bc2e49b36c13b86b536a
z7eb878e397499954a3aec42eea684b03c1ea23fb9525efb1cfe687b56cbae9c0925c159a9d5bc2
z761d491861c64d5e9b2825fa3f0081b9c4b4c46ec8b9cf2e82c1a318e523ba05436289c5b960a7
z7b669d1e1136d3079ddd2c1bc2e2389b77f1cd01ce3f3a625a4f673c6b2497da8eb466a3e15931
z28911c67860252844d5fdc4f5abcf0c1ab68139c640096e789fe74fdf3fb4b6baba4db518f2c31
z55fa9d5ea2df22d46cd11ed588da281ca039d37f7fc0b1e5757e7af3a5517b78c2347781369c31
z887031273f245ffd31600d6d2488f13b0de8e9d0823d29ef7eca92b1f890cac8bf5954cc518331
z96be748905cb96aedf44bd763e07c7e409d4ddf0255085cbc855f03e29c3c67b9b1a3f5bdcaaa0
za01c7c5aaf658021306ed0d6b22490dcfaf1f381532e21b29389690bf59f913eb9f49204ba2d82
z444570353c605d39d6a5867c26d7264d3445a3e1f63df76da78de37b671c390db18fe95e502ef1
z6e96b11cb99bc9779f166f419f4bc7fd480641a5b2fa35e9eea5b7a2241327e76415585354ae71
zfb8e4d53ac6d9945b4a5dfe0a6c7e528a05db0aa847b58f501bc6390e4ad7fa9db74b4e2c10093
z5d4920a2e634b3f6ad6929c6762d01f8d28dfffa239262168cfbd290bfe6d4b0b423fb5fb575e0
zd3c53a89074dff7518381b1752eb68fe94c0012d7595b19228b3ee65fdd5f99ed8f0aba44cc008
z5302610f2025cce3a4a675eb716aac8f21e2c788e73acfa018d4b00f06a986ac86f6fc45845810
z2a87f431b09d8d0473be10ff87109c82a803d62c9f48c04bc2f4728c5f9dbacc76dc68dc5fa745
z1e8f16578da142b8b53fb640051e5410e06c72db8a7452e52e095cfbb41a020fc684bae117138d
z09b58dc05e98f595f99c3d6fa6b78f10e65186a90158d9e05c6fd85748fc6c2e6a385ff6493c61
z7c2f116f520bdf7794c7fa9263fc365adacc602e4ead9f42fc48f697a248ddd02f6983f79fb570
z1b75db83082dc5678e737603b9d5d8d4c7ad9789d20d2cd76b832093825990d4a39e7f45b4950d
z61e6c6a7218109587750e2733115da80dc281db97cad469ba0c14fa314ad92bfae6fb8c4da670a
z0fea15058f6b765fdd88c84a580bbff4c22b89ed0160a5b7fac1989fae6f752414ddb86f640e5b
ze807835d9057442d7a62c3adb365fb7972a239536390383e4b8ec047a1152c8a1ef71cf43b45c3
z1f54746f5d483eea5cab7e8301b41d83cd23e6bd849f7883e1722ea01d9479a8701333c9a096db
zff6ed6dce56fc2d95b02e99052bced1df5b0e5a1dd46eff73490e7815b2f570309ec7062ba34fe
zb96f7c077f7230525a1bf87ded40202f921c3afd3ff672e33127266f60a1db1f5f8a4d8bbd8c7c
z385a49597c85af2dcfc0f101ee24e61b19c13d48dd1623ac07b99449e31faabcbb7351422c28d1
z5db47407e0bf1412a09e4b3e39a20afed5b3f68b35fec3f6fd09af84ce1a4623d160d2f4fba188
z6561d16175b4681b0843254e5c6c3ac7f2a0be4e61ab6617cea5d98920e5f199628127b29ff44f
z70b3e4b37df715eb29e9dbbda58f5f1f29aad6a5a5fc2b1d31be5999df177752a8fdd95511f823
z5690b3fd5f407a1d10c501b26627195308854c647e5c9019424cf059d1eadbcd4ff080211f69c2
za1ea979ae4cd445bdcad41de67f2caec2ab21d2aa2eb0eb4c99504d24767ab4ddc6db41f378bf7
zd72f1dfd47ba1d40e4754bfd0809966b232ec0d3b38ef93340aefbb9ba9cfbac70c17ef95d8a9a
zecce4249479d106e3f8907eac4ec6fc2b11eb11641e95748588c8f3487064d2a188b2c3ed2bb69
z4cc180f93aa6c7a29c21c3c50d5f51a5a5f59fb427ea8f94e440fddeb60d105cc34d965bc0ddc7
z9a3f050a5b5ba250400073d2bdaa7de78a4db31a985992de364bdfd17dd6766239e6bfe27c9263
ze552aedd7b6b774d61e28b323f4ff890310c5d3aa033fecf979fba0acea79d50895780ab649895
z9e8dfc64116677c7380c88e02ab2a285195f062a0951fe00bc95f2a2848b2b5dae49f12ba54307
zf756e7c8397bc90cd977472491c0fc6a50a7c726bea257844615d7ff8e0f3662f818272d593030
z337e5fe35b8de6b0550c99d03bf9cb3b6a1f4f3ed9f2f85eac0430eef53e215e7650cc043eba70
z54d0e05a6e42d73fbbb534a7ed8ac046d94e5d3cd282cabe14d9430d3881ef853305f3df6c421c
zcbe5aa465c1c061e36c771e9cda9099773094075321d54ec66ca81365ade6cc0671acb150f762b
z5895790d222e4850d94bf3d34c41b9c4278e57bbf41bec417f74d4c8afdbc51c21e4858ec0c81c
ze356011711f51885acd73e9964b4bae2c933ddaf9b3d27623f194bcb56b6b6ec02071e2561a6ed
zd69a61312c516f841a728ba9784cc2d85de1fc00f3993df504dc17dc16961d3e074e00a8e6c4a0
z83c799741afbd3501dbe75f2ba07701488f2b40a73aa9e96d8e9554d510b0c7961a965303b5958
z7e38d6ed4a4acba81c4ad45fcc1553a63ff98ac20937cf5b5635c3bff07e324823cc66a900ad6c
z5bbb002b499dbc66f781f0d000c2bea0248c7f6e1f9b7e30457971c9229480bd9d8ab4ff2badb1
z63a2031fa054c3091428458db0d4326cfbf38ca3f698672980df805a96dceaf28cbc69f7e953f1
z96da6bc8337c69593b42408a18406d1d18bc65a5fd555d09bd400aa6d61e2b94146c83fc1c01b3
za41a16a2b6334a67dc7c1acbc275824942ce341dfa0b2c3b29672b27bd16f0d2e7f3bafe017e8d
z648154ee2ee2b007d19430e535e84a14f14e3a6e686e4c1da3b3ffd4d8a9566aba4c0acae799d5
zedd2d0d872bc2a8268c876666b3074c3ed0f87a2c2bf084d527654d596d7f0a0608fb11373e84b
zdc8c541cebe25902fcc3d9ffb39651121ab1f01a7cd01d8773c6d038353f15eda2ad60ae030026
zfde502209655b55a3f40e0f3aa43d9fcd35fd7d8422e2ae15427abae7e088ba8064789dd57224c
z455e70fff1babb72a6b3577dc00773245c9fc7b6f9d53c11aa4dea6cb63c0788866771175f025d
z85cf03d115f691546fcddd02b3e6406145883937642f9fc78437291fb7db474d141df7a11ce7c8
z017bc19329cf53d7f4469c789f1fb2afa0a253e564b0c39c401abc6788240fa00bd0a5b2710be9
zdb2d87acdf8b147c89a1fdb558a24c586b3e5a94a1e239d127a34a6c3f3cd7b4acf75c83ceff0b
z5c7b3b7e49a7929eaf9faeb0a1f74ed1110c103514a0f684183a14775e09b66f6eda4d88c80646
z5164651589a28bddf6b47e8794f229f40e3df3671ee7ab034844cffaf66b1c152fbde4fa019710
zdb094b126bf603e16634f25ca20f8a5add4bc43bcc95ca1ec825725e525aa07e05b90fb48a56b9
zf6975cacec86a76b44b1e6b51f01f538f963e1959093cde42f4da1cc9a5f3e16907e8cebfd94f6
zb2091bde9e4330fbb1eb1df89c25891d65b551260b64e4d4017d73a103d160fae9e73f8ed47d9a
z8dc9472ed1e67fe45ddb2a32bc4f279a9ee7c3c64636bccdf98bd8370793fa6c98ab717161b374
zd0416f6a6de6602a3213e8f83f69b4c1a25d2a7b661245761812d37344a59917d5e5ef446bae08
ze9f9f205d0043c97530278ad685c530da577e9578c8d773e54c29981005961a1da8f175ee801c7
z7bbeef2f5f792df0b549f4ab1e59767d18803d177d1b330d1b67ad6ee307c0ec10c7a281802e3f
zf7859f7e42a5a73c28199cc3185cf77e39e66ec4a1f1e6c0bf137ad31f29e11afa9287136a5dd1
zb0e5510618d7324841eed7cd6f3aa04b4936d63d0f2fe4bf161dd19a0d466623ce37e51a1ddd7d
zfb4fc863b31316102fa0c7b1c4709551710e93ae13d5934006ccccac90b1d1dfe43fb9956ef353
z09ba039e7403ea906ee73ae76e8386b6e36aded82f770ff7e72f8f338997a92b6586beb5a056c4
z9643abe49ef678ccf305c3e3f2474b36db7f265a8742b7c5c28e85b77272a679b59ba606d47aad
z29b8780beb5415417231ebb0cfc457c639c76d1d2e0bde2f91a3a3ce54f4c6dd0a740e5009fdb3
z41b1b88bdda32b639f770250b4d30a2a9654bb65ebedd89a55246f1e0d220a9968d2acc5c16b4f
zb4958da3e52a3e75c48ac9e9ad691c56db2397d11608ca2d5b06ec0cd26321146d6d393c5a75a5
z4c6087df12a4068cf13a4ca0f9f4034aa4891edaa9a08432875ae8ee61c8ddbef2adf19405fe51
z0c41fe1914d5128df7d52a95205165920f5b491788e9ff75daabb7307cb69d5c09db5b3f50798b
z1a2f988a2a51739fec7d626dd22b5c7e0eeef0ff348a08d15fd85611f4a6666400363b7dad9fad
z2c6ef98ada2901df44156a031da023a5348422564d4b8cd0cd815a18b657140c9157c197b8b7ca
z53daa07754daf4b34849e532750bc5e30463f5412c4d3fe9db7750cf2dd51c77b821d7070e67dc
z93daeee39a48f920548da0738ef755bcc9bc7f9e0b651c1b2d32b990e30d37a4aa4a341179547f
z096b2e22cf4ca052fe3a6385142cff49c3ca34c09b20a3840c
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_express_transaction_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
