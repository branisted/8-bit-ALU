`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9e91dabe8e7975bd7e1fce653bb8d6c5ce39703a3dafdf810acbfa88a75a85155eb269dadbd
z9cab6e518f61194d972240b3b06db552addf599795da8e88ba3c212233d8455fb159cae2ee1ff1
zd9ac02aec24cdb1aba7c7168dfd44d844950772c402d8fc60adba297c33414f85885094385de52
zac58a4bb9892d28420996d3efe9a9f9f7947fdfc55a06ff1e0e41013a4f48153e6446eb2563dec
z6747a0c750768a1adf162c9120a1b3f3018ead5181dae5c28eab4fe19ccc291e4d98e0f664c33e
z169de7b377511ddff4d0a4b56352f8008860a70c74d0e5a974af65a72f662cde619786138fa84f
zc69467645db6e0266c5f7b634898f1d765ff9f843002a9872bed6f0e1347b2ff4812e74bb7517e
z29cdc154ed3443ab30b8053a054281d2f1be5c2a3c7dd8008f56f82a56c92d4c5e0adc4a3aca80
z174b6293910ac23a5f640e4a89efbb1639b70ce0f954adf865250185ee48871425355c0629f2b4
z4a1422f023785ee32c9f8655a5a8a608ac00c951afbe48ee94e65f03b455299a93790e14d2ceb8
z774723f40fd186afb5f11fa5df9493b604e0d231c3e6eae4191bf9d5e242fcab6ae0d142434573
z3aa21f4ef85e9f263a31ce705cf8620feb9c679984dd12e07243c29430ae51cda44cddaa4b2c32
zced667af65d0438e0bfff477d187e060f852557f6daf8a9c839b4137ddec566105f87347544271
z2176af33913577000ca1c185e05a1355265e2db39e8e8bab844f211778887a8417fa0a51acee16
zca8082d90de215e78ffc2fbfe33582776ee4f897ef779681633c2605970b540047f907854acc47
z6b9b8c00efbdd216ca22432401ada83d158e0b303e031816e22bfcb777107e1a604a56fb4fa734
zf9c95c71a519f56f65323d8c7b16d7964b933edad6fab63ce0cd2283d4d03bb4b16daf3124a26b
z037d39d1d405095c052618181a632ac7a56ae6ee162294da7af640cba42c4a830750a488386653
z0cd29b32ce6c13f73c641103876bb4392e414a42741446653880e4edb5c4a69ffc6be26352aa60
za2a1fee3d84f4bee3c126e16a2d15d828ad3464296ebda2248ddfa373a2b4e00b87760433a8507
z681291e561438c7424ead0816078a75588f20711ad1f8ba7e4576448059927bf4a99f0a251ffdc
zf7d9354ca83336c88f20b95e2bb4953dfca23f979389f6c03f0a46d423e506f8e935c8df53db25
z6780277ce37308608dce51dc63123542dfba347e244438f7548184961a4d3368882c2e6ac37a4c
ze6a5a99b2b523745d13ef4dd5657549914a6d7fd9ea4b00e90759df0ce832f0aed446e94a5442a
zf2d82c8a8085662e8847583c76aee9904effdbbd6fee83b63239812c14307e9551494e1d6f2880
za6af3f0b5df8e1f00a99fb5f2078edb82cb50895500d6afafb8f1d780d22530fb019f790db9cf6
z0907e5c2c14d0bec2b433d9e1ab319efa989c511ff78e227255bffd2cbcc27d104603c99359622
z51f8cdc079a668766b22b1902d085da0a00133637cbebd2867a8debdec2eee1c4a9c940f5c2c58
z7517c8f8636b5bd44fbb413b1b74f8f963499139b7cce0199a3ae613b8aa65a4e86c160cf42334
za87c99e0b655ca64cb2e35357a596f02f20d4f566c2ae3d5a9bfa252f520d5e5493439b825e5dd
z3b700b1f0778fb857522c3ee13291ba49448ead74bb420746f83ed57f541d258f3700822bbc947
z1476eadfb0e5f2e72ed7060560f1b7fd03ffb10e0eda7f38d3958dee9933f486df13e3edd9656b
ze8064380e47121c46754a26ec380025f0cd4e8c60763e5f82dfbe455ac71f64f46f5d3d71ba208
z28f3d177875d8a24c6a54d3e1f5f7a4ab271eb41dd7b189ae24dc1a2accbbfbdecad9a89c261c5
z548ba9ea84e77b162644827ac5c3c780e762e1ac51be6ee85805e987149ba5f768cfdfb47818ae
z2c28b678d0732fbdfeb6f7cb15c1e5f73e524b82b5cc74aa08448070f3002721b02d4c4246bb68
z0c319450426f36b95bdb583e970991b5c93addb7368c804f8f559757d7b7686a539e90a5dfd7c7
zb0b883338dcd85a66248280ce76aca6294131b3fa6151a9d044ebc32ad6dae20d95c0b0d840efd
za5539c92ae0d1353f1af1543d2c7ffbe73b8a5ec1d0f9cb4f638e7b024ac8cee97e04f1f9b0970
z0f6f6982f5ea20c61ea39ec3ee4b734c126586514cfba3001a66686a8a5631f85c7a2e3a5b8ccc
z05e2876d809ba6b1a16c53e273ae84bc61faf7e086419d88df984a3e75822d21357ee5b661e1d2
z3495ae97a38d0b6477092f7df6775f91f7dda9d8002c8661d6515a1b7328c916eac623cbeecad4
z10f38f465368f566d39347fb7fa01d7500e612bb304ee2594b0e8f1a7f6eb76bbd6cc616373ff0
z1cc03fb7520de2d2f4ffcd094888fd65e69b19f768f7f0844728afb9a0de8add4fd09218ec78cd
z1ae8a1982773ddb6cb7d592705362302d4cc22fc5bdfaa3ec7565ee52b4dcec850f5fb0424c971
z3d635504c75b11c73bf31629ee576de0a7499cb01f97a210fa1734a939066c2d845ea873c68ccd
zc56b7ede31fbd68c28968fe66b9deb2c1633ebe29d5acfb22a32b9e6639320ff2d8e97628ab929
z8d1f0204fdbc1aa42401bc73a18df1e8528ce821f8794a96f8c2e12df56eddbbf0e6bd5c504ee8
z051e45d21767171b330e78e04b6eeaeec15084da506b18c7f189504f0db97dd1b48853220b5d58
zb4b479eeb49bba0b0c345356380de623355eae0cab09966ed8747ecaccbdb58544f1f309720763
z524ed76fa43967c322ffcabe0ab2c0269a6544447628613ced65ffd2a55462fe187e6e2e052f17
zbb3496157554876675c3887d978bb8521541533ba49aa5ee132b78ef8b9e7214f099a5b9e9956e
z0f3c64e35d628ca655e31428c9d2ed627608522cf32d6584d6b74bfaedcb9f6189da7b3aa992d6
z013a12a10d12afc37fe67647fa7714a98d3a1f37e8052fed473eb2c39f3ef01512bb57a9d0d5ea
zb62fd6db481fa58a6f3ad2655dad10f3483c7089d25409f4e11953d4bd1523b7c2bf14907e42e9
z5e8be9e7dccc1f7c339c20dc4be33dd368ceb6daf4ace62d74aada5f3f86a20daa592aaeadbe69
zf8a458f0d09e87f7251479849c6761aaa4bba4c6cf0154457c4ff0f5d002aec02d50aec7c25efe
z4bcf50f4f980c8f6ba822dd3f251d0ce251c3a5b8d8992c6d1f0c43a0f0367398318a981b0a486
z7ff200a11d1b5b6f251a20e48ff0e47f293ad22c473a3a37f80a6756a2f9faf6542aa095a4f245
zbbb7f54d55dbdf0f05fec760aeed0c8a7540f7488c8fc52f0064a91ea9e7a03a61726c5650f525
z00f2d0a6d47a5fdb0f0da5c9433b342aa0b88e1991c68934938d395806bfb6f03255f807ad702d
zd278bc724213a42841d3c59f042cd9a7b6828a48be1fa7b272bbafff1422f414d6ba6c426e532e
z07ea9b9e7eb9727296bfb50f321a846cccd8349ff2f9e07cb481b3995e3e911e2b5b891c0ffd98
z30e5e27dc056da252bb16462bec2c429000cfd8f6bb418ce8e0129d6741675756b6e48e98d4987
z674f369c41ee6acacd7f0092568080c8edc3aeecb44f6c53323c1a72c82fa2bf7c9ad42a1cc9d3
zbedb5df318fb6cd4d27054f5865fc45a0d321176b9b73834e45d12ce4832799756803535b4a558
z8b440eb7e0f12e37a07e9ff3de627cacb4c9ba8439a286c400d59a401079dd9a4a1b6280180a11
ze79acadc4302b56f02e94f8fdc17b9aec50b64b1f31125d7e808fa55db5f4b6bab7abfe793b450
z4b7460a12fff89e9eb03a7611c1d26b8d81b19867df3ccf902318881925226b2628d6158fea0e8
z3716f91e155bd75bc58db424aa0da0ad07fe21711f26602d349fcd7ed94be804c13cbb8bd2f100
zb971ac3170193980cb0b9a3207bb1a083c3ea75e1657cd516e90ec319450ab2597fe4f4cfc3626
z26377316ab9dafb6fb33e58484a6c6c4591d08b1dc54bce84fe415cd1148e3429eaea8f4ff345f
zadfee650f84d359a9a25e59504bd5980ffd8ba23355c9dbaf22ddf4647e623bed7290f710eb113
z1a77ce81c0f7ed1413bcdda3f134d116e6399b5d8234e476d07b0433c69e843ba1026087ff5e74
z3f93a84f0c0e548fc254091b46b03387bd7d2220fc4a80a6e2abfb1c67128f41337a8cc7029dbb
z0eec30234c494b36646746746b0848c9a7c4850477c448375e2856196f2e9e21cff54f213d46d2
z2bb66d8eb4033e2c0714e186ce77010bbd7481fda29b2a6f805623bc6ea69278b9c3618fa0a4c9
z9eeeb3d6ab7e8c54c89bc372b31165f612552d3cbdb8c0689654b32106e62d76dfc7e2edfd0320
zc5574a747d1267a736ac35ba0f1aa59f2a2a2fd315c7de0ca4874bc1fdf8517d8fff5de1de8958
z41c5f04413f9647805036d405f6ccae110ab24a554fe678de3325c2adef57852d32d39f8c1a230
zf32770c419d89b1fd388967695911916fa9230c6fe1099ea81758736b15ea74bf8aa2be060fca3
z1d4997f7c97572795134d8436bad238bb8a5a1d5cc0b985787c6b57cf4871d47a5b7e4eb464067
zf2c81221c8a7767ff15007d27661db9a4a3c311fca94fa9fec9e9a794d91f0dc8d952819441c0a
z33f638fc75a34a9e0b1464cb9694e51474c2f3c749c8ab195b0884fc58f77005cd4f203338b58e
zf279eb714eaa8149ab9da6615cfdbc4d8ef89c3a63cf613e3d58381b0cf2ce9f999313947eb459
zed58632eb998196d0fcca3c4799d07bd8abf69cc72ff21612eb19c75c065bd0c435ebafe85569a
z17c813ad0d263a0dfc4dc1258e515636e506aaafda3ff45a059279c5c842b034731c9d5564734f
z2e534e53ff05e84c2dbcc51b851c968d5beb178991775c5a131c4ee1bce2b62047aed89a826f6e
z796ddd52ee31b91958303cea62380614061d06fd63837e95c2cb8286b150103cb45adade62cd74
z16d333d659ee7d073d4cc7a5324d6724a0dae29473b47945e1277513715493cbe493183a2b1800
z773bde262cd2f65f39d8170b048b2ecff770fdae9294020f67bb623ca936f26f1aeb5c10184a0b
z4cd3eb2afca1224625536741577739b89c5527175097345f3834c34e6bb7ac8f0e2607d7846da9
z91958aab8a3035de33a43d46e635072e58f0de3e3f8a6192f54239210f21bd2f330738cb5bb1e0
ze04c522158cb3381221a9e30b455bbb6b28cb292d0bb8cdb79e00e4fc675e61d23dba3738d4788
zb1ae5823ef488ba5724bd480d3058b825f679251910b1153ad6f6b9a69b83f2c527540758bd2a5
zf24700a0328200c05203a0c09cedbd1e9893671c0c22be0d1145b25750a2cc48708c265605f6cb
z72ae99954c78718553d49147ced84bab53645fccfd30915aefe19eb450d8ad61439b149b61622a
zfab857a9b5e5c0459df781e65614c2939a4b214376ba6aaae3460b025c4ac39192e1907ae2c360
za107714cdc3e80bfa6747fd8ffbe9585a4b4f0bec1c20d13c2dbce3c09160e0fdcc811fb7af703
zb9984435a46da6f8ca8c5928416db34d374a73e3f5f82871899aa24547e14f28f0d7068a5245f3
z4368239159dab3722a890565ab18d13bdfdb01317544024870ff8c32583b981f66423b1eff75d0
zb0c7446858df5a5f208ec041c7d2beb5bcbabff31f42ef6b32b3bb95da55c16e7f5e97bcd877cf
z84fab1697c0ce005b4096739d38b3ec7b0e5fdebd514144d09a5aceab24b8ceb0fd9ea0ec5b649
z1bbbd74df44fc6de11f8ac928d568204b44ce175733b01d901b251bc238c99fcccc3cdc965df50
z5f70321db9c478b4239547213e77d4313ec610b04120e5673ff1eff349c9afbd3a89b1c471265c
z194fffb748675fd55a034df8908f4821a60cd97b9262bd92d82fa3bad4acfd302124119813ee7e
z612a92dd80de4db920297e6160dee0ab55c484be88ccea9d05ba2a507f8317b133aafb61afaf3e
z50b3749551122e2c4dad07c27a847caa730a3de0ce30e8d85f9dd45278f16f9240cdc80f2ac8c2
z1d202e200a1072c31b8282e007f7d24c1ae72d496fc2500f682cb51e3e584cf4fa1d3de5467409
zafce21a2d4189396a0784210a90fa969991bb7b880b924a4b608706698c828e50bbac4b922e125
z6eac644a514303ab1ea0d0e962a9a2d0438478c1e7d133d9377f8764e8bdb71160340e6fe0bfc7
z8c46b5e13d89dfbca7096c6a4f92411ef23b19a162a527fddee00caba9df87398404c9ef9878ac
z02fda893eb8581dc21e540767b9ff219a1db400ed3cdb5c1020fce3f6abad5a9f4a00a7690c74b
zffa1c72a96dd00e245857c2486b51a07fb262a9aa9f650f18cabd86133238a816d3981b449b2ab
z61ca6881435fb995843489ffa8a271ea21a98906a5ec07c5ed9e7e2b6cedbad4e8d79e01096b21
z3e87375bb221110407df4549f42869663213e0405589da73be9cc82fa6500cb140a37aff262b72
zd337b3e947c5167ca850889d3622e13706ffba8fc65ef70e62a4002703f70a06f64fe6060e47cb
ze5deccf05b1231be8aa22620ee44a1589d50b66273f7fde154d465f77d0a20de471b98b9997281
zd4d89bc43f118cd932ebfa649a51e1516654ab6632a7455c5507b64ff9004a71aced282342241b
z2bd839edcebd5c3c04747bcc09c9aa4a9522cef4d2fcc94e3bd84860c5c05b56d0740ff1ad9e0e
z9f8ed1be4336c0f529ea34900dd8ba4e2f4d80d040cf905d162d96a9c0562e21e035c968ab349a
zed0cb22c0fd3a397c68b842745967320936b372fc8a507bf5e12dd5b58b68d28dec27ab55b5803
z970ca963d72edb3cedba4268fcbb27b06d76d4fbfe4c64f34206e5b80e7410b13ec1ec27fc4841
z86ea284c5ac290a991bbeb264ef4bc468043c6c5ecf448f3997a416edc782ec04f6e0278ba42f4
zc0de2686ea1bb5cf31b3d1945ad1098bc0a65f242d55dcf462f5100099e9c486572ff02aacd2df
z9971210e2b1fa27e77b832df4e2b9e652500ede592416d896d098ea9bcdf006a954d99b7d66433
za829872eacc2d3222f06e43e98493b034f8ac4b013205ff6494d16ded9d010b40e21dc96b028e5
z9dab493825a07420af1d6c10730fe445f1b16dd3706bdbe0ca452a6abef615d00fbbd013819686
zf59d252602cf12b1bd75fafde1840657f9dfc4c5739aa7f8071e5a3e7704c61f484c1531fa9863
z4a715328407ea4decf55d8439aabdc17a1e55efa92b95078ab35e518b89f624f172f2db497afb1
z921e871cfcc59d81533663981b503fa89a02530f2020a6250356c16ec37a49f73b410c81703985
z0203d8f6203e6033ac0272b20cdab342ef461c6b1b8928947b72f610bf51e31f9dcee42bf1c39a
zf8af5ccfb71eed2711f5951c7b8d33f384f351562a56cde87eb19c8cec7a514ae024433cec3393
z24081050a04e49dc4f5df6deafb630dba8fa00df6313d42f74df171741393a0e973c3fd9fbd549
z5be77838e5c48d60d11bb49e7409c98cb76672be40d5e4f6cc0c548be79066dbb6730cc0fced78
ze07cf602efcfbf58a60831e1e46e7ae88d69bf3eab976feeef5c5b6d7868f338fc463cc17678ef
z2e8708863b3e65b6db4e893deb7f26ba0404df771ae099ba8c3d75b3b37d313431ea671f32f020
ze2f373276ad6391140140a670ccb954b672b7c560949a5f69346c0277f43e8ce259607edb78c79
zc356c40c537e78991227af6f03d8e98c1d2a29725b0f1e9687877fc795d29437b689c75bcf9900
z028a3b16ba92bdc06da1ab7f0b1de2adabb92f639ef87c0c33212342c35c249791836f9e806d3b
z21b4bee4758444ac74ae571e796fbe6a9ee60d98f8de9ca3093d39eb368dfd91776b48c239720f
zb1b40ff0139d891a666cbad446ecd90e98410ece2e9cf34c594137dff1b79f7ceb2a877566140e
z7e9af6cb48eee6518ffeee8a8c01401834e259a5a3bdd9f5c068d5ce95094a395aebc5ba605c86
z65e36b40b0c5edd7b8f3260f69d1d8d4e44d364ce5cd8d106597d932cc5192aa2c84d2a83a72c9
z6bcf7dbde9726413b0cc0a08f2a4afe3e4e960152508d64bf5090bd82ee44cb57469f14c79daf2
zae188abd2c7160c9efba47b081fe34e1510a03c92c9d9d6c76666ce3c30fba4f10f9e4df9c5089
z28bfbb15c9b1addaac65e7b939ab417d1a72f3f89def3a8511ed1dfbaba9dd690b4bdef9e5bcc9
z315292a929d3368d4f7f19d8055c75264b1e2b60f2df8bdc080065ab63f3512e67447ac9a371b9
z2bf7ad47fe8f89292f984d23f5d755313889bb64a9ab00eda67ab66d505fa02f95adc0ed4a10e1
z45098ca55a71840dc85de4f4d313d1f830661c87fb50e8453a7465911e4b8ffe729027344b5d76
za4eb8e9a038f26fa9e49c70ec18ed386d477f0dc0451255e4ec39ab1a626c5dcaa986da5308365
z9c38f57e721efee5bff27f1ca605e822713b50a58d18400721ff9216a73818cbda3d0b1cb856f2
z9adb480f75db36743d90cf2a7af67be4fc0ef4b95001a751e502e50a51d211341659a6fe7d5246
z0490ba25d428d60d8ad2c5ad6fb7258d219b55790500d23bb80b7a4ff7ac63476686c2a7528c37
z129c694f796c5993fd9fa2cad1fc5191e23d645f46bb069bdb790964f6aff1001475072f6d688d
z1fb0d7c99819864959ea8f4128e87449d9822ed729b91ac463a0af039f9d3cb3fe7bd07414b168
ze3a750d9811496d7fe990787e5d5acc07e2c55afc651c7a12dbbaddd5ec589d7d0e78e2a39eded
z57cc20b7fd1715ca34e30e51d913be1a540c9c0521f7021857959a94b221b9ffcaacad52319297
zec122dfab48589566d4be55556b7bfe65e0b1d6cdd925f6edbf412419cfc228a8236524df42716
z99bccb47c625d952c0e53f58e78b84e96c2b151fddd218ab2a68004c4c7355c0bb4b9230d782c2
z49ef199bd3dc010149c4fa1ab7eb3d25d976f1fdf3884b2a0bdd2f8a4fc1153044189388d6d40d
zd57d7334c9629abb1cfe828fa1304e5a252b57e0159de1851d6bbe89c4b3cfc5256e8df76a4d2f
z3254e2d607de504b164a5bb23921068053eb27724f66053f5214d818a9f30bc62f54ad0231eaef
ze4d664b1e1aad926b73c9ce7304339b56238d3f1d4495723ef571a3717be025acf0cbc1b4d5495
z80d84709967ed50084105c9d32ba97ab7ee4b476b87a92778c5c51d439ae144a6937b26f1e5d37
z28522cb331f26c31844390f95b34e8d56ad13d6d43dc043e80beea2080cb5904e61737bac8dc7f
z3425cf76cb3fe94961537fdc97681682f7eed50f06e644925d8a510a172b8838a514dff97db1df
zb16c5950bba83e4228a24ad8cfc8fe3f2451eff841f3f820ffd1ff60407e304309a2f1dfb329ec
z5d53e9bd3a4ea96caac8f6a243a8ebd81b4d8e95444825796a7491486166220e8633bab1f20157
z974c2e2b22e5e1e31c847fe9900d7bc321ad75550e1b5b76dfe4d6bfb7fe45f0338452c7490d12
z63ed5a8965f09cb80f25cb4e9f2f2069a70308b0d8382f377c4eda60542ed9167bcded6fa25862
z224bd95e7d2eed65152d44df0e73e859a946773f83375e6606f655fb49bb89198838622496d7a4
z062e466595da
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_three_state_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
