`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bcd350d8b9
zc71703b3d6e1b18f9ab7b0b63d0d3cd99e08859fbcdbd2c3a70031369ba06de2aa52613af46a9d
zef0351bdd4f344e3e1fd770390f1782a301b2d4a41e5b0728024e583fd840b734fbfbc2539f723
z470c09d9e1b587cd379db4726a33fc581b18676fac14f107324abd517b7c6787930a3b628f4a18
z0cafb36d5f96e9087cf62f7575f95635b6e174b18a545bbfffe03667abbf543b6d1f6ef0e4a343
z6b8165bc876c5dd1d5ea659cde1dcbe304e2d324c20a0ff27ad3ad85b724ed25fea4e4d23eaada
z239c6b59af032b8788085248f6144bb594a2079fc8c2c31b1e3bc58305807a49f1725a9cb26c49
zc4a949f2b7c00d9787e2461d7baa48a21b69c56caae6efa436ca9182b382c5428303fa7c5a7510
zfcf5a4e1c5bbcf3cda526b8103915964e801e2b1c5daee37113fff79dc54bad17e82970b003687
zd0e4647eb4e9924a8d57722398b91a58afd7033964212770beb282eca9638e02224a9ecec4d6c8
z8eca9983cc3f0c8be24e1d983fbd9989ba5251c1434d3c8d5bd056c970e5ac49b9739ccc983ff8
z986d58a615fcad5cdb74f0d8c56e3e3e7b42653ed82b2dfe9992593c75f0d217e707537f601731
zd75aac013fa113359e7e53bfcf4d1301b07aa0260e5fb5a71072ee13eec061b314621a2f2441d6
z187b7fb7cbd3669b4101a8f1de06ba6b7c4aba8cafe5643008d856f08c07bc8a461b4a9f8fb41f
z602d82b644829c2278944d0b34d020b12190631c138ce7d571bd484e440aaf8f519664086f5cc7
z41ad5c25464d3920199be3af1709f3234eaf183d0a5974d50b9154f33f2c1457da5cce7fb0b734
z3c480da224b5296a973bb386b829385cf3191ef80b7424e63c34762e6400b6418ef7e88f375918
z7772650948d3327776b28986c99f509cf43f031985363b1454631f161616bdb9b4d35e28f6245f
z06b4f5c7627645515ad95d47cbef0743696838301d18cf66c3f9a9406fd7f53e74c4227795370e
za095217ec50b6f081849f562369a8de96057ee89a1809b94d88e6810b18e2f5bc68454c26d7e77
za1607ff7b3c9b36d0008b1a374074240f8990db4d0002cf0dd79cd26da0c132aaf25b666c59d83
z5f84593f811470b352383dc2eae4a74b8240130d829843853f580f8c6bd8cd5ffebf3b533ea8ec
z711fbf11b1a5584e3415ee3eb8ffaacec7bd98a342b78e6fcb8a1e631572a64371cc0a7ab3db31
z24475d7fcf58a4c7b76a9b7b14383dcc265bf176d65f2b57f6b55af5417c0f1cfcdd3961dace74
z896c428c1779a71f74025df7de4b6288af5888e560773fe7a166cc2a6a4eb8f7f8bc2f9396e37b
z935e177ef7155a0d49d7baa5ee4a769d59bd815bb63db7fe7ae381cc37861717ff8aa5bd9185e2
zd3f231bdee691b8ebb2c49b601ef303bef648d076c0f64d987a897a410f031854be115ffed19e3
ze9deec8d9e529eab32cd48a2cc46352f7faf17ef5aa5c1d5d061a41b5df5b74fc8c35a8b26d8c5
z632e0cad9f28d20800045da4c8e29c31916835f0c81829b878f2bdeb4aef441466d02dfa60103a
z49465b4d24cb56eaf3cf0eecf51054265c83aa8144923223d49fa8ada0f8cea46694b1752f3cd6
z367d7868027b5ffa512a09629818f06a46742eb0e871853022fe4767531e213bec1b20357932c3
zc0359333feb946ca37666221afeb3aa196c1eb39889c7f0d41e5475b027993f6e404e6a7e4c909
z4336c7ec31c14baaf7255578fb25260ef011e691a4b0e065ef9a1d43efc56cdb019e7d17ea0f89
zdf38ac5c0d29610b850be13f98bb950917ebd24a9a5e885ea9078bdb739d28117b7fe7d8773cf6
zc8dc7321312163c2368b2b0ffd99cc47d289bd6cba74d89dcd249494849bdd167ee07322c50a4e
zc689c423ff64cb95c5d128a980a9529848617140875341b74fbb24d5f2ea5988bef13a02b3e5e4
z0bc1cd03ed380f05bacc552cca49d29ed4fcea5ba01a10718fece13d0a72ce9ce2f1e61f2620ee
ze3a3c87824ec96ab8e2316403d56559f4a051904bc235db8eff9626fedb59f5bcbc49d0f7f2b98
z565ded58a1635aded59cbd363c25aa29a7ee44c3c6c5b0764842678bcef6ff7b31c5deafb23995
zeb0576342094ddc684e022bd62e50f5c99badbbdc5dd2ea1d744f6151515bba07f97bc3e1eec0f
zb8771ff7ce3c04978bd6bf004921a1c81199d3c64882f9d6e0f9a956ecbe9933416b6beb084689
zccd23ac0f6fa756f0b1cfb08c94a623f5beb17ff18ff92a24b8b9ae6c3c1d04cfa66756e7229ff
zec10b8f6a6a08a366db7b42a5af62ee6f5f5d5688a9dd9befa834fe12ea463c630438a78ce0360
zb58306f53339b4c538edcbb42bd934d98aae1814e128b9e0432b1d67215296e7ff129e8be4a472
zd63929a5f49c0744c12ad376a155c802b71453b59cd1b63d70bd5c9292fb1df2c42c345e7528c0
z73239c57fd65c1567d7827202e9a983e527fd23a049383997ec8ad3fc3535933711d1b693c547f
zaf49fce7b33df549fef1362642130c23ca4354a8e47f81342ae072287e01715396ef349acac57b
z5f2a7f9d56203a5c8a99ef2ae223780ff5bb325abf5eaa91ee98862f025f2304403c621e8cf03c
z9e64444f25a1adf458cd67ce68181530f377719b5bb11da98eed6ead5f2855c014c18e760a9f2d
zdf8c8974b5a4022143d599c76d429cdaa26369aff32171f4ed637f42cf12cbe75dfc0481f88e8d
z6a6663ed24b58b5d0e6982ddc29c9c7fab84613337b9ee18720c8cdbf32bcfb920a0cb6ba6b931
z18f7824c5d6b1b3ecb0e05c5012b1eca0d610a1e85b558ebce75f8aa276bc587f4b6c87aae3bdc
z3c4fb960e81e541efac8fd399be84e0d3efd8b1ef759fa81b2b5ac461133cf5307542026322798
z2f030642a9c244342219721df49afb873647ae956d8e2e14b496b10ba2d950bf1c62fec74675b5
z5f68dee2cf3a6241eb95d302d9937768408e2a5b39ebe2333aeb48ea1efc4caf71cd0bb9880929
z7eeb133a1e0c36b4d1267e08fbd4aadda288cd6230c9ae18953ea343897f60e3bb7caa4929234b
zd00dc47ff4a7062db0d8f08bd8c89feeed07fdeff257681ebbfa41aeaab8ac2d46b52189799871
zb1bbb870b5aa5aa34d8ac14754d8d3e3a0aa2919d534945dbc34b8aa1f85503e38502a7b7b2674
z1eb3104a135819152e836640e5dc2ad8d713987601622684253fa086a59767e3f96ae3bd1eccc2
zbac5d3d25ca1a5066090dd789a4f95ca0eeaa1957e211ce3ad079dbcf96f1a645ddfad6c399ac7
z747a3778b03de1792f649343186ba910b7bc0fffe4f40c60ccd8f99246435ca62a9ee210b2453d
z19836008ece0b60766d15f0a9c221de30177ffb0d9981efb82da867c1fec29680fe7e1ff475dd3
z930096d5911d52105f3d9c59eb70c29df9df28b0b97a2f9c045bd69ef091c515e657576690ece3
z12ad4994769f8e7d1bfaf025433ac527645bca35d068f9105c56ef6d2da8a08253d1b6cc47f4a3
z941f0c781aaf3d6d9669152cf7554bef4f8b43fc2516960e3382dcc043f1b367a681e3d8f0b353
z5d1d5d8b8dda372840fef830ae50f826804ee20cdddc682d684ffe7ad1729205fb2b60b4439a25
z76c431c05ee0e413a2748096517f42a4b304afec772ceca57129535260a1cdd09f921c79d1a965
z51f302a73e323b48011656f3036ea3c638627096b957568b386d4f3de16d8e67c3d85c3ab11223
z20ae92e8e6c277ead7dc50b2ab88b44a9d465ceefb74fadf1fc79f868b831a1dbaa34f37afbfb8
zc106f61c68911e8bcfdb400594ebe7e40e80313dd438d3be299613b98113da797449ab8d961d9d
z84351fdafeba3d16fa5810df859af416723293349553d2a1614176f297a270b85baedc429a34a3
zf493a9bf854365fff4665ba123b64c3e27ab2155823862a493dbc04f14f66f0f03a0651ab3db69
zc53ee334783b97b3f87a0ad4a99c57d8157ed9ae8c4fd3062912e65631dee3d8e6de9b5f202eb2
zf1a151168f6414e0775472b6703f41169f2449bc0a8a3374d501af1ac29202b72b35049ede9d80
zd8f256b5976f612ce41a37ec42dfb69dbb0ca1a505df1b16e77186b9a2ae3b1ea5e19ca135e939
z08d49dfead827a20d2366c496628853119ce8141266a63528301ace0a906b01f4b4c57027dc1ac
zbb6ce7685bfdd7ae728b8940f538d75ae0ba6fcfc79aeb747a0b8ee3158af3fd02c24e4c072dbe
z33227a52904479034670599240e834b657b3cc71afefda45415db4c3d6764573249262da2cbfff
z1a8c1805b7b5c9f7edf1d10a774b1320fa264bb3e1ca9ed1a689dd99ecc95fe7a375e8e001fd86
zf771f499805295477993f9904a98e6a351532652a88304ed161021ddf90490f64faff103bfdca7
zbcf69e0c9a69c193369d323e151eb5fa011d91650adc3e3b022650c60bd2d5e588039d341ef86b
z50b9cbf13bde34ed8d6eb9d0cd6ba801d47ccca6e4858828199a2088a63d81f1430339f6d2fc50
z7607838f12b0ee25812cdeb2803dbea8b419cc6374af69c4d6bd46177b0d6f01b2fef24e039604
z32f4c1c393c5fb70a02ca5313b4b9ac25eb94acb487d5bef1a01e7cc39ba91dc35453124ca2bd5
zeec6558e7fee2ba08acb8ff7c728c3353e97d3119cf5768d1c8967898e3f4d8df2dcd62dc98ac9
ze2b63f95f5d8221b64c4051b182fb79e41876ee7da9d898d56ecff2f71cf927ed65cf346846c81
za78f3bb3e02d99b0f61c27ed518a46cc11bd71c3710fc37fcc269d6f0cf7527a4d49ad7c75f97f
z26cc2565a8ebdb8f2d8629f09a9a426a2ad6d1a683fd9a259d1de92a848bda4b00d1a4cc447863
z6d1c3203c5ddb475874551558f8b5ddda76877210f695421094cc5baf7ec3b5b732b7c2b28136b
zd45e75fca337334fe20b36c8667ce6988447fcd7e736ddd8b534185da73ca8e8549f083a6a7082
zca09ded680a75337d4d76e7da2879300cae790eb95616f88242b6b7767b816b056bb1813597a8a
zaf8d03237741165c9f2517acbe3be4488900313861b6373bd51c627b16c926e427b2fbeebdd602
zb99f79a69c1afe0597ad3fe3bb9178e4fab7b1b4f4dce5c083e63bb52313f4583386855174a8e2
zba3874c5d2007543f034ac5ba4480ca5b0cf67fffa9087c79400e639ad142ef9fe5b3d4f9a85c2
zca1ced9bf92dd145973eca1e24f952a3a8c8bce620d43857d6338ac3ae60f4396175571d945c82
z1e44bb805ea35e1724afe21c8bcd905be771433580071cd7a3a5317ad6d9e5515f7cbdbf01b10f
zc0021f1573805d16b173a347bc6df285ebc89542347f668b8ff41c25068ed24ee773d3fc091208
z466dc38f3a6b504b8daf6602f4929b40b44688a4cc28ea2a6b933ab2d0c3ac9f2329b14518a037
zfc11cf4c0c6a21255fd1af0fccecb786202ed57bbc0e27fc4721474bcba833127ffd85fff467f9
zd38d1c37046cbf973221ef1192928bc6b1e5c1b3025d20c94e9788e0b612199a48543106129f24
z4ce4c79c1fe8bcd2cf4e6bb369126add5a5cac34cef239e540a7e04864f6389654bbe34c29e137
za756d3930f32cea64b25dae425690aaf9b297b3c415b1aef26e3f5bbbffff4934d45077cc8ca4b
z702c218cf95d1f99cdd3685a4956fa67e9941b61f73d1fcf6fdf119d0860cad2cb2922be3fb57d
z7fe55e9bcf38cfb75df2534845c405a2beaa7d2d7516761266739b3e5019344a6a92046cd7d486
z60c2b7e939508c89dd62dff2b40f5845597474fe7e2c6d26bc018604ab562a3a383ae4e4d915a6
zb0d3677515261b250e67817811156fe9b2c45dab610b179f6a1a4bca04d59db685365c603ef8f5
z2cc64b252f304d073c92645f6dbde9b08df4ea1bbd66643e5650ea4d77e0f7912d073dbc95eb9a
z9878baf8c63549bb514c8026e84450f70b6ca2795fa476ded5f282104d6630cc7da35dab6b17ea
z215c79bb044ea188c0931bebe9a3921e61a7e02ddf34e909ee3e6b05aaee4da9f6bf86e4d8c375
zd6c55bfc8b7419e65394da87d247f96f0425be04ee0d8afdd302d7712d4cd49a1d0a997e832912
z050876e2d30acde8bb839557de8172117207cd248164df0d981af112fbb6b984b47661b7f4761a
z43c5624fde24df1eb4bcd9ab2906b8a16cfeb611efdf809e1c772c7a6c5e4aa9ae0f4375469fd4
z6f0fa45ce34a9601ee2e1a93e7bc8e0b7a3ee15b7787c6d866809d50116707b609b94c92c37503
z3b6320235cd61ffb9059dab8691f10f0a3e5cae6a505a51585df62c45088026b14ddeac88fb447
z5abd55de747d9e6c20bfc0bd0bf2b488e3a9a331f9b33b350ae44e1ed19ed9979ae3967b4188b1
z025355c500ccc393c3ef91d4da4142e92b413efa5e1701f09a0838f622ecab723d9af8fb1e3665
z4895519f3cf6e974902f02d80cb416bf0b138f01c6b0bf408220cff7b99bc83cf58744f7eb7fdf
z3a9be7a7a82a4a3a66ad6bd8c280d1d44f5e7ff390af64bc9e9d04b7dfa11fc0ee429c49da357d
z353ea2dba300b7f4736915a9ba9396e1a8a79de79873ac89235dd1bf06db1654905e0321464e45
z49c88eaa565e1566a165eb57a5d92057790db07b058dae28199efbf8725c12627c48bf1d316736
zf15e99fb002c003bc8d103380759f0e11ccb67a88de55a0e1ab7fac1fb66e3abb2f7b49754ce4a
z59d80636f3fb54a588161eaa4ac9d73af15e2b032f223eb921df52cd2b6bfec83eeb529d214437
z4b8ed4c785ed356bc094fc2caa6f3f6b61af89483763f8116f9374ecc2da24faa72d8057d3bee1
z699cc12e7bbda428aadd14191dc6d72239d90f9648699f815da47e751a9e225e498803956baf2e
z0d248f00af437c34b0e622e944a189e97b9aefa2b81e2f5201474b74e39d83377cd6df88467b2e
z369781846024aaedf5b1dd1f25ce1069d92400ed32b6626548a3448309994caffeaaceeac9303f
z8b7376f43753c1076c633ecb28309ba9bb11df5d1f7e700689a13379bac75b3235c8ffd5f76c44
z841aef5b933ccea1deed7b149a112b6c398044ca9d35f63d091c7a4a0f44f1d8ccb061976b42a1
z313bf183233ac4adf67813407510b5e04d546604cfbf64fa3bddc4197450199f62c96c1942854b
z40af56fea7ac1c37b4b279fa5335c8818bc25dc18fdf6b39615db9705811c7cb28f6ac0ecd77b8
z0aed2025abf761eb686649c095c56a647798d2bbf38ba71fec71205252c81fb533d9ad015225a4
za91e12d466135d4599e938ef8a7f7d1028b505ddc8d15af5a7189b75cc7c08f1448fdc86fe7de6
z69166f5a54cb1d0d1fa6b5d4528aab4ba54ad9375794076a16e30d344abab279c158a0057e0172
zeac75b59a412f8f91284e299df122b90e7873926cbd1e517b1327c70df09383555f1fe85354519
zda11542143bea5092316c5d7af2bd7a22102fffcb7a3d5a6ab996d8c0c7119fbf32770a008365c
z9391bac788642c8ae09a3bb4acd91f60afba2ce0a361742f2131e05b47e6eca9565bbf8d5c7f0a
z36d980f718f68f0e9907c269a6d197b4efb070393fd446c7944c5dbb7ed9af8cff5ba670f4bae0
zbe475540e296503360aed882a89a50bd6f751aa014652ce3409f0ec772d75d073c2ffba02459e8
zc8df9cd937088ecca4bafc74071a7fa48070dcdd831e5104b743de2eee4bcef359626d36771461
zd4d6dca4b525a45cbba26e13feea8206fef93446fd9a0ae25cf3f3515987b445198d8a31ae1ea6
z78a05675b15e48039e0d336e894364e03d543aee7d134713e94d5fc72548e32c003f2a586b0a27
z40fd58e68f90b8b9669ba031b90725910f3526d783c13557d0a737ab5c688645af0870a5dc64b0
za25694d77c033f9fd7f976baba6ac2cc044627de49e33facdd2bf8ab5f088537b9e40eb8c47f3b
z37d62d66f88f2b543d908f7fd38593203fbebecff2a7f85676e1813ded7b4a7091497de5e659a9
z3497a7eddbc8b9fc7a3fb6321927cf0992b371af6ae1d10746a861dc865a0ab33d948528371e66
zdc6addfb1b6f9c91d279dde2dd04c468d41e6ad3275647dfa8f30cb949f59022639e3b80c58ff3
z42bfd35eb19a5d3d6aad42b5f32219092d31c8b0069e340e9c4368df9aac54c762abcafd85316b
zec268a7008f7f71dca7d884571b787fef7abd2470ad957503c59b974aa8a2125b7472ac0dc7c5d
z073152600559b29421283716a38997612fa116c358a5ce0f04cbd79ca5001dcd5820e52b31076b
z77e2304dc118ed26bcca90839a99d7732e7b3e0213dd53760de46890bb4022c500c4e25a9823f1
z90c339fd2c715ae6497a10e8e5b56856846ce75a7b53a9c129bbfc530790b7eba87efa49f6602a
z134602dfcb7ef865cf15d68d8d894b56de49a7a649a7e839d4571158e654450a711f6a96569952
z504e54719a333e6c8344945cc9fb561994ce9c6e18a2e36c57f525b32f6e9886dc94e88d26d104
z4011286d311674b1ab89cd15826ed535888b0897046eb23f431356907ad447ae7b6d4e9c8f603d
z187e3bb414c9fcf190ce59a00dfb8d28664b7f644f7506c3f4f8f27884178edec2e9a4b60ae65b
za5b7f06dcf28138ab0b11b22f030eb79e3d3fbd4a903daa8a6ec681634cd714a692f6f29d027fc
zac5979d850f1418b0cd976571c30098f5bf7b025139d5c21ada3187c27547b57960dc5ee66f0de
zd3b086be34cb5b1931aa584a47f88b644ccc01e83e49d71938b3add53457b0bc2cf89ef47b7558
z36b0c7a77537b49084decfa5131bab507061dcdc10740c7ac9cdfce06381d7d264ceff2b80e482
za9058a7a1a7b1885a9c8e1e3bc4872ee10878a3da1976c0a587bc9f72986133cd9f938891682a7
z112ca4a2be2d4063cf818304a65c574e9f4c7f77bfd14117b22ed39984d48bfd42594259c2c763
z970575363c1a57fc5b100176f1aac6b6300dc03bd49327c48fcec3ccdacbde398fba44ea0a9436
zbd5c067c1a38e7263abbf555f50fb71a8fc7815bb05ad5c8d624ced09f1e2d56cf54886f8dcb82
z3a9a7e25dd60760d5caf886c9f9d06a4a4487c7d704ee9eb0303ff6325fb589236a1b6ef9a14c6
z3d538a80fd026197de052a08af58377ad95f56df73cffb40a85f296ce11c89d9769b29595fdae4
zac31b2fdc1c1f886a134e87ce49c691cbc8c3c60cedb11a2f6eede3a4cedefad165e48089bc718
zdc15042810b28e04f9b7c43e1b53580489fc76d89b027b1b314bcf4400ef85d99deca88e7a71d2
z4f4d16000bf08049db80faf790d64d54362e949bdd705ce17b6ac54ac6e3652f60550c7a7a1db7
z920e1681acbfe352d1e319e1fac2dd41aa2bf15a17f1d5a1769bf70b1fd993a164e8ac0ac76a75
z26a3617926572458b61a56d234c9b627c9c4da492233128ebd114af1c84e1a4a09a89c6288b00b
zedc0fc91f074ba63e9d45d7110535bbd24164e62a9ebffe75b6e969560843d6a800ecc70036509
zb6e46b36a8bf1033526589c859cbb1d1f970ae15858502f4a53c23c0e6b97106c88ac11406c224
zf1ca465eb8b263d84073ea502f3dd7e175ba3cac04acfbe8cb5d14f8a43190ccd8fa41998d73c0
za3a4de56710e54bf2077d2ac5bbc844ce0f93dbacf064f444b7f1074640e3d118699c5850c76ad
z05b954cfe35bf1905f8d3efbf7d2ac478c5ecee23ebdaafae52e8ab41aef0451269f3069894457
z61eacd6556f38fbe81b674a2f388472d07d8fd85c6d6cd5b41362112d5969017e1ba098ab85637
z0f41de47e7fffb5d4a3d9091814b70580a515e71139d2b2818f29739a7b9807578be9091bfa350
z969d2578208240bb446281e8b5803d2a99686bfedc1b14556b3cf212da804299914a67a4acdb82
zd053a9e94bed67ff41ecba77fa316ca21d2422c59a6772a86b4126848cebde21e2b16c2e344b3a
za43634bfc68f7577c6ede55c613b6fef1837610471d478121244cf927e5c13fe9991c17e5d8b13
z2b5d03d0cc524a0c54a2df5653d5634313932381838a3edda5195cc3654790740e53f2792ceff0
zfcd25c33dccdd38ab6ebb57ac0be10a25b230284cfc631b5fdb4b3cd35a402a44aff58d0209f05
z39f82f87af8a8c127e96e0838539c6dc810292f0e1610b825737fe8cd66ea4493c06ea47b08fd9
z8fcb71748971b591853d3a91556b9a0f4dab892aaaa2e7932952bf6a7a52cee9824e4d23e11a69
za5bb66dda4cc271ce0f9c8fcf0263342537321716643081f6d40bc10e305b6a819017c02a902fe
z279e570ed6edc5641846c0a4e53e45b429bd041407a892e6586630e8fbfad5fcb849f0399c25cc
zab875cc83b83bfd9d999705d2956c1423aa005b1c81d7ff5e26b9af8b3eea3cda2a5577e9f6c98
z50d2a3f3f1c5891f8c39cdb019c5a2dbfd359f17e18959c7c7e9d625d33caa2c7f07c1c5ff2306
zf979c9f075088e03046ba63a169000f936d5fc00ebd42f77d1d92adf7e5581281e3dc35639db82
z5c334bb4277b96e615eb7eccea20d620f3d5c9bc73e6117190d263ada66b09c401bce7882bf208
zfc26deb6e9da309b1405d065ef81ab3536f5b3184155090a74f68b8d59f85c5410a70806395014
z06a3f712097963e9465a2eab56a5da9d40ba60f55d4ae377c6d690b4befc0e1e573f10dfdadd24
zbdf2f8baa3cc0832c30194d9bbaae6c31df8df6a3ce3f90da0fe89853857c10df6b4f80947b08f
z9df5253caa08bc82ad1d7f96110f84472ea0d6424c550771de96daee4bde52044c9e6744d19c65
zc57de932a3c11e6c980cf250447eeae992480b637fcd69220c717b64ea95dee89ff6e73ed16e6a
zcac804aca3e55061e2424739cc8fe13aee63fb828397db2c192edc23d3290ac16d9021e4154e29
z720503db775bd8181da759bbf11ef0ba20249a8ac2abfdb99b80bf27387e1d9a7b774f52be089b
z95ba7d926abe8a3f3373fb0ff81d3c3105179c7bc575ed2680fd2b5e11ea9096bd68782fd5081c
za43cb339ac6962aaf07d04f645ff474a249b2522d6c1ac1960633fd4de6b95e8b48c9f3708a68b
z7a4135d01ee084cfed3b5d79ae95fd8473900eb24066863542d72b542e613668b4480eb7563b69
z1cd5c99694635f4591bd7f1dd5d67ab209f566ef841debcffde73969e34b907a9b2548bcf16730
zc17e1839b947f95743ac4cd989371c7887c597ef64b72469119998c4636c669e5aefaa8b5726c8
z12f8e0006372befc3008d43b86f967b9811ea2fc4a4fc727ce557ab9ee19364948728c9bd9e434
zf99e8ad32881ca027b5ce507b4262dddfa91f4fd463c80f2a4afe9f11f4ba9d7e6bc7a5b8ad10e
zf737165a0ef03c8c289154d6e12b6ae6aa02586da4c96838c5310392496517f874d566d7d35a23
z42eabaa98b71e2abb6b6d56bb9c5b240cab284ec314438539a2b5c2a92e0c1b48cd277002e5ffa
zf83aeb8127c0f0f05663832c320ba2cecd39f3e8e78c11030203e430f3b7c99abed900db2faa8a
z1a875b03e1bc973da752fbce293715377ab6936378128e0accdb1040392e6dddd3f658a7d8048d
z1da7d7da0f819bfc8e4feb1f38d06cc78c4a431bae72b42d88e70631e935657ce1b275c48dde88
zf3ad6b9565f93687a88195c73e435a85e90435ae1d3b9ae0e1e5cb40691ee470976bef1e9e50b1
zb267a5e647e755ef263d7b25853929b86237637f78a269190d0e83c76ac4a7c28554fdff92ac5e
zc3c5caf184b2793f2bae30d3b21a1ebd88fc99336b3c9016c8bda8f531315a00ee2cdf7ff0ce70
z5ff7b6d8d698e3cce94a6f4020b6f8ee11f4ffdf8658e2f3877d462f8c43fbb0da4884001ae54a
zb38548a8d2bb89580e2e2374dfda86aba02ac0acc0ddf096435b35bc226cdf3afc085c431465a6
zc71824aed09efe495eca841c82da29a898448d3ded10b403778f5afeb3bc61c2b8b9dee96c75eb
z870ce3787dc7669838c7c8c244bf1e5cc6c26c8885a2cf47f94d992cafca56becb711f2e8a42a3
z0ce0a91a2dd3f3d5ec58b17d7437a1bcf30d1789c595ec8b211f3e853bcf0630d78d4c335d6ade
z2bc31770bc3624ebdefb472803646e2467e38ecc9a78abcdf16e12077fd29b366f994775f4516c
zb805e690130bb897068ee3bc22aa63dbb570ae06e28f5485b3d98ca27fec6131a716097d63f6ca
zc779789d4d40947d64773427a9871b90a00f06064b73877c89bc752bd4ce3d9aa2ffb480b724bb
z4e6e9757d541f0e53fc7b0e744b269b43274b109950dd1ec7256b9559c81c452823418fa50133b
z1ede52cf3f587b9c5428dd4c654f98551427fc6dfd542f01096a79bc85436db56b5ce6d5f2b39d
z63b0ff1a046d8e0451bfd8c09165b81293712516bb43c6d21825b0db783a090937831c20467064
z56e5d7bd13b865829510b74b4525f852ca91ba75ad5920075427ce8947a81cfdf8d2f0daa56a9e
z45ed3891d3bd93d50b2a9108b831e69589ba826bf708016337a36dda7cfd502c5b48bd5c770cc6
zbbbf19ea47475ace4784ae74bd0d2810fa2923b1131337f8a1dd52ce2036b1cad12a2881cef300
z816db5a1f68c83b38b50fdb660cf71293fcb026c4cac0ce2559b3007d43442d67f884868947c20
zb46666a5d09de2fec20161354bea9a2acb28b82eb3e70293a397884095cc2cc2e9428a03c7f7a3
z979cd4b57026017e5e9fbd8b6901d965e88350f1752d075a8cee1c7228eae5242e3a7f4178773e
z3b9795db2a8b63eea0a7658ac67a06c12198cb6646f7ad93e4cc7e873e377e01ef995773a05a3b
zbc6670f0368f45ae9daeb54e6401145c5b19916d08ebc84f8302a039c526f408dd843dd34c98b3
z03a65d76e8dc9d7530672f8659a162eee9a748d989e879e421fef10ad872f7819be8488e931f92
z6ebe2bcd55149976aaf5f8b13c9da0aceb882ff64d7f3248f09f615e6366a00ff3c7fc21f9a324
z04c150951261f5eeb0dc4a08fd557ddfc847bd6389201ee67ec86a7abff502872a4efa7b3f6bd3
zc393510188d192534a1d5b2f5070ca0f5ce4f0e6748963fefd7f2b32a19bcba3b383238c346f45
zde901b78226c4b1f4230531162832fe9bd334d655ed852f2da45245714f2e61752e4d7714e3c8f
z971e9392c3dc2cfe3ac2722606a43c05d9c6e6a0d94ad0cfa6635165ad9ac50199649501152c42
zc0ecfe1d4bdfd1b7d920dfe0288b937f65a5c3353559a42c755a7f8fbd2f11a480e72a1070714f
z271338d40b4ff8e16ca6ecab25d782b2c8a2760f7ef98d4a9e9a188d4393dc3636f182c808c35c
z906106a57c463216017143fca572f89fd27928dfef40e8cbf9ec3afba86e5c751507f2303bacba
ze90a05533360a110986a1f284eb0fc6f24075d024b685866410c6259a03a4f001cc48a09003402
z326e973f8707b8bdf7e2d7f5675f4ed142e49ed1d4863422c8683dce09c5c1f61b6e0ce037bdd4
z62d321a93dba562d81d1d64dcd9c82ec0248a0192694966e1c9092be38730bac16c85a9877f71e
z0fe5917be022e971e3f61d67a941366b1e2724ca4b5163bfc46a652bb52d4d0551abd56f070e61
z9b0fd8792e5c5659a85f78b103ac1ca4e478ac081086a9c3d3a235d347541544c21ae12b067201
zf22c72160082a6ed053aa0d4a9bc432265eed39466bae68ec724a5086e5fd6201cee8b634aa6ad
z451d89825b547ba87dbe095149e0d6f225780cdd6cda151458ebb8df7cd4790eb60bd2f92029d9
z02e97610906e0239bc3c46e476bb5f46e6d623444ba3cb2d8847fc18784fdd644b4d47f8f71cb5
zf22e02970dabd33791f89decd6e147d0f03d902f8fa60a1e30cc9e918a8c67319a8e2d0006f94b
z631bf7e3865af21605ff9e98392a03e3c2e258ef20d157debd84c17c154c6da910b73268abbfd0
z78f85b29de5fffad4bbf1ed33af84c1658516c30287b760aca5726e11bea22cc74345cc4319f30
za382aaa4d288d1b97ceafb5e2e600554fc27cc1b1feb6f5f5bc2b6334dbaa0ac76a603597339ee
z962b041f6c7016ed1ed778beb84d6cc47184c30da79793cf1bfba76a37c1a5625877ba2711844b
z7039e51eca857fb33c07fbcbb05790ee09baac09fc173d9a7eba0b69103e7178c0bb54a7f5065c
zdf093fd5bcbfca935a19743016a760089142f4ac63850c20fc874377a653d6931d452b9e7ac354
zbca7026c6c516a3f3fa8e79453c46bf1bf5d46fe0b29d286bac43615a850f4aca12c237ff2ee32
zb210d418ef2b62bce85e04c8d42b9baef051c3d625072bbc8a5664b7f31b658140398d8c52a7dd
z69dde80419dc9f3e80d1711664db5a759c34ee2662bdd6163d29fa7bff9f848dcac3ecdd77e577
zc7c21bf50401c4fb8cb64bcfde935bacb3242ef1d77472a6fdea7c786db4febba4f2e3c0f7b990
z04d2c698d3cb1b76ef12fccc136c807e3ebdce109dcfeef62e217be17936d0d5bcc15fc9b93fdf
z2611f7ed5b83b808d39d1696fb262a2bc955717d226d1bdd3c04454de460bbc180187aa0473cf5
z68374668860698216739fd498bc8663e43f73cd832ca1b0157e360d0ffb2076cc280e9d82cd94f
z8951ee6da63cc72abc10fa94308bd4b1c0232fa1eb31d9732a8c1bbfde5d456108aba5da89423c
z17ca61e241c964d2a0e84181ccf7a467e7d01d0bfcad9b53f200430bc2e42786a8a571e6307ae9
za661f38ef2ae8a360ad2533d93df50b5969380d021d61c4ce3adce22ae78efb42218c2a09e9889
z6d4568415edc487ee9208e7c18aac153aa873791922de15fa05d1f6aeb99d7c1beb26b44629a60
zd2f190ae216faab48a68af13eaf4a5226871dc3207e10b7b906649eb27bf70751c73bf44464786
ze40a95b4d157180211406b94707a19bd9b3e67f4eddf88d0c757c96a93ee652285489a72d02c38
z87efc7cfd15e281399ee075cfcd0e1b75758e755e0159f1edb90ec8955c0b22911d199b4fd28b9
zf94dd87f54f5823a70acab58a41054a0d2af9f2640ff6635b32afd2af76b67a043b540807b89b2
z8e9a2cb7914b19b31db3aec7a4bf2421aab5020d26ca356dbbb16984e2bf74a5a37d97eb4d2255
z732deee5dd3bacca9d5108c02e6ded4411731d904f839e2563a08e6cf3808ce27e69ef13d83034
ze36982921992e0e6c580d47ebb17af8b82acc02336f210a1e847d400f32fdd2328dd85c29bff00
z5262d0d5473dac976b9c95ab0831a5089929b18afa888dbd2be789d9c35835dcea6033bb5ba98e
z5d512272f31f9f426335409fd3c0fc9635fd54de4c73740c3bda3d3dc4efea71b89947dd56e5d5
zb1d7bbb96ea15bd52757503c5e56cd034d15ef29b1a050143c4017694bf78fde106a5993580192
z52964c571e0f4a5c30740c8a3c214f2f9cbac3c27cf3cd0f9abb98c9b1c44d209f822f2a3dc2e1
zbd0d1e7457ca480ecdf0cd78d66232c5e4ea03baef61c08d509cb26aa3486e40c3cca17b4d28f8
z274c11fbfb9561b149cad3ccb480e0e91005fbae8a2e9a1d9a9dc490ff86dc70003731bd2c7959
z0a6ed9dfe7783707049e09591cf9d397bca843ec09823b43467511ca75482718e2aa280b95e138
z505bdedf6e99da985d87f189494d5680f03f8336d1bb6feee66d52d56362713715f1edde39a02f
zb01ebeeec72630670eab248a02599626792b8c6342ffba16dc96f0d5f3dc7f4cb449436e2f48c7
z404a6216d01bc0e5f337ef0b85e12ae23f9a35f2f6871d74f2f2c25061f4155816e48d9b82b667
zb77892f1884c34cee898ca1ea146c7c5fee481faa97af8cc4c39b284f27a9fd61761385b770043
zf0000e08389a34d2f000736d6b67c3042e82c551c8ee236ea80fa778a49b742ac3fb0e7d02c742
z2c5232e53df689fb93b437c889b7746e3df897b91dfedd307ef5ab83beb465406fe82698db3bf7
z6e95dff5456e49a36d6ea196036383b348e14f575b77146873867aa8d2e2d9e6f727f60b5768de
z08b0f222608af9b9ff1d930190e7e9ce17e509e62ddade7c04e3ff05060c11bcc448b556f08ac7
z9d48a90b4144be69e78b62af563c7866407f357490ff4c4fde8b898281b9fe6dc6603b52f56cbe
zc438382891bcab2b1b38d4cac07af4b6089ae49409143c0978ce574fba14f2b532ca2299f2bc80
z9350a5ed5b8b6342ce9037bc41c10aaf38d3fae9342c6e88cb633ec8932bd68c07df551b6e395c
zfd630c646c9b35593d1d62f63628ae9b0b2203223cf9f821f4bc84e9fbc265f6bedbc3eff71a24
z91ac444bc55ca33f2ebb1d5e63cefa7c2eaf560f268c48f95ebd579d1c7c7996e7c67ce7ba9970
z1f76f2629e0670e59603da382d7e591166cd9481b2b5ee282bebf860ae0f52957a6fdf3c3a6f3c
z0c5e74b23175289e53563e51d0e682ddee2832da4039ce8bf13a4521c2026f5b079c223b2b8162
z23165e63183e8c47d86068f258ff45bf6c5821b09fbd9b0e179b72b71efadbcac061965e251127
z0c82997fd011d18388fb1477b5738529fe7276e4d5a0e126af472b2a5270f158c6210671ebcc60
za232c985e36e4f10d6c2a38491851505f1d1d692cce9ba26235ebfecb17f220536e4988a03de84
zd97261a4bbae90408d5070660c35940233aace1a35705834f2b15982e8c053cff80d56c8d219bc
ze3ac3bccbe5e1875e3edafc8376860e35d9a1e90abfa1c6d010d9b513e69b48746bfed79bf7072
z115736e4745b3a05854aace571509b7b756fe6ed7e36809e5c3fa55c7af676ce1bcc9abb63a9c2
zb0f0cd3abd44a24d34cca2ec6c93e4cff7e88aa05b4710c8184d9781a3bf7d6ed1169e23f73295
z09447880d4cd77e4a0ed286a3985e8071dc57307f70c6779b8ea8595125b218d0eaae4781082fc
zb5dc10ae678df0742bf41606f396e274dbb783fb6681ea9cf27fc8c04748f1e4d057c001069cc5
z8947948a0edcc159e2bcdedfa3a4433617029556b9b9b70db83c5d915b0af02594ea80ed6cbbed
z9a8f3f7687bb76ed4efde17d4e7a780372e9238ced0cd72ed146543c4334c13133ef465d1c5afc
zb0bc25abc565f17e421135d6fbc66e8f06d99f802c00f0602910c1f50454e8a4719e2b11b26473
zd2370decd3d80b7d56652958130d397734e9f8651cac7d66141a835ffaaa2f5febea77262696e2
zbdad0edc80246e04fe5551e5f53d65a4c8490d6ac1a8349948e5011ed1b721b4a7cdfbb956e00e
za1a5ee8806ba4c9dff2504944775f752bd2ebc471d7718b9e1f6b42e891fb4b8029c54a71f2400
z19d7751015e160baf3f71d5a7bf8dbab162097da56b6e3ebd17f93af983e2cc456a7c5457ddbe6
z3af08c6cec0ad879bd5dda024e295a55c3861c31a71f751c7bba1da355badf4cef69ad43595b72
z679940a0504e913df658160ddc956fe22b92dfa60073834eca58923bd399ad53b9d6cbb6f0ea6a
z81ee54b8fe586a4ce93d6b88ad2b70d5b75d052c9a66154d8ac276c9a7decfbac563492ab69161
z21351e438be31f0e09832ac842b461ffc348e2e72bb4d404bf052910efb356a00cb0aa93859628
z6b946094b2e5ea557d5df8bdca637785a557900dc06b1d2e26c35ede8893f9144620ae95498ef5
z02427549e022bdc50318cd54b81e4e5c0528d52a277c1d622d17ff5e408a1d38f2ca350270dbac
z62ea3034b32000aa8bebcfb900b9d6adc736dbb70b0c07685354d6f6f8364c8b43867674d6c8a6
z7a158247b3a8a9d51e7befa53de029ce0febcae8968b97d30a4dbd309d9f7fb29f45867cd8914e
ze9c206873acf0914e00a22b7a49724313976c1a8c20d5390c206922f25f92515aa8c51e7f9c102
z943b7cd332d05cf84cb13ef7c50f7585c254866fbbbc225c9f21abd60acc6b3427c02cba0ebfa5
z69b82febc65c1a5ac5f63daabc83b49a04ae8529b1146e82a8f0b876687f4a7fe912bbe8e7cafc
z0dde95b87c73f4fd6e639fbfa7a869570766ceccf82f2fafdd183346c4bbf2eb5a351f7f14a291
z9a043514c638edf7b9546862c8f4f081928bb20b09f1dafee82c05d827f6998c28b768ce03ff82
zc0d5ebb2c7700f362161afb0464f1ac15375953a41f329045a631054ffdd6ca776e9b8f8fb64d9
zf0ad21729e5bd73c9234a246c998887500ab9726554f59ca53abcb844f236bd3568cd5f5552ae5
z429835e04d4f32638ce483372e92aac9801ce80380846e10dfde4bbc7551be4b1d32ddd40b4a9e
za74eff7e159437ae6b0b4f232fc8f02417cc68c9f347d31b2807dba0b8d4eabbb6f93de95b8afa
zd0388c5bfbb4dbf1b8c3353add15da8974da303287e5cbaec63eaa7f919b079016c71d078d18fb
ze62219bbfc3cdc62d67497433e7b34b02c05b982a566242d0245031d04f711072446ac19f875a6
z4ec97449497298b656a6a7d20e2820694bd237db8a0f730012637ad4173209e887d7479b0721f8
z651ce291ec01176b3c542112e306889c75747935de07b6501f64e8f1de44a0c7701d536ec4017d
za7eee457e140dbfb23db20b80529d3cb1d4cc4b1c9d15b2c4c1f82041bd021fa245ddef234f281
zc51019d54b78703358077e9bc94b172203fb6ff4c0dde15bd4949e645a5f2c0968e570e3d62874
z4b392289cfe7d89a4fd0f7546a7c75c99b1e7d13cc097b688ccf57684bc0b2fbcff08d05ffcfcb
z8e4296c7a1c9cb56c46f5e36c2c7887a2690aec679509a3b881278bd8d8f02f437b2a7ca027144
z0e6fa39615d3ef9e5f9d6dfe2a4bcdf3dd79511ce87cf59084a734837a4335d30257049a170f63
z2a42cb1f350a8d89f23bd57e6e8a082632f502a6535ef0a1c8545d6055401a9decef1295828f8e
z0a68d79642cfd743987714d51ea3faf4e22ccf9e7d9eb8ecf4cd255e304c7d493be3e8f8e54127
z141b7e06ceed1f046c46feafdf0ee72655f346ffd24fbb0f7841687e02fca37c654827d644f1fd
zaa44f1bf8985361b09198c1508e7852203c60fa9cca6ae96b49fa1cef528a055631d96dc03da33
zd3fe7af76ea3dae3527162355f3e82ad63c42b11fa45add96797a4973d20c08e97307b57ff6791
z896d4f8047cc36f134ee0b726f04a18a41d088605c2638a4103ed04c7642651b8d2a6349b89e68
zc5b20d6ab90777b80c55bb6f0598986b5d2988ffed0a81e16d79a67b6610b0746ce24cc0b389a8
zd6694e203be4616082e515c4fedb141bc00ff66b3450d9ad5c1bbe88b26bcfd48559ef7d12896a
za21089c6ba2b2e3bde8b2cfdc131d0aa7254fa7f671c2a9f1df328d84072fa363eadd60208d331
zb102aefc771b2eaa0025ee4dd8b08fe056b07a897c424344c298ead8d07d1c23635a4f47548504
zbc371442b12e96501bf542d00ea239efdd5fe7305ab62041095a72aa8c000d5c6b8df5f2b337f4
z7d125d67e5523a8ec4712ca76e1742c9a653065569eeb990e5fe2fb6f10a97feb7ba99942f172c
zc0ade8166d80ef062cddc3e6bf9da16c07e429b5134dca3788d1c571928fb3ac4ccc5b1089be4e
z930c9580cefc8d60cec571f851a5d8ac1587bff5dc1e021f4e2dd2ac066aaff34faa5ffd84f774
z2c4bf75ea9f242edab7d81da91e042eba8da0b422fc000b54c76eb3bc0ed2a4cebda327be3a608
z620c822a4e16b4f4aedca050f4e9d183727d9280f936118a81c963042d4f187095da69ef6c0bf4
zcf27970c1e7ab40a1902c712e64e831f0e5678ff4cbefa65d0de5ac695ae8cfadd8d82ba7cc868
z0096f7c280c7b984a9c86d713542f667dd2a32f5b5a0e59b0114f092cdd4d9d1415804878c0201
z4bd1132e931eee1bf58f79a9c6740d9390f47c198f8e312226791c2a138da750cab22694ad4033
z078e36a6c66f8495b6322e8175e2da64a663203e97ff6035e23e507d8b401d9d57817e6864a630
zb42d4214f07d9fad512097c16ec7b7f2fbde17bf05ddab90b1704bb8a284ef1ea81117421992bf
z3ed72486afdf6b17735ceaafa474732a64914a17172dd30f35a5db39a7acd2cc662d0f637d5fee
zdba916935eeffe1048a473624aa657b4fff4798c83e7694352872c3578a6315f490ed7d90d25e0
zb6688aec0d1c5247dd967a227f1d1a8cf5b73f4a27fd590e762419a5fa2258155c4404a457152a
z7bb5ae32aab47b789bf48fef66ece3ef4bf2c9f7989218b4a21d507ae10bdd236410403f64f026
z1ea536955b6e62751462e8ded6a67e574c0ce3c3c73c4c0d23e1ad21e5797ccc70d3eb2e4ab4b1
zadb675525c0791db2a641f7584d1302a84859302b5592be241668c065656bcfe504e5d412af331
z75db2b7f1949f5da930a43c1b32bc4cdc8cdb21ba9d162cc7c883231f814c57f79d66ec85b5af1
zdc1a32c3462b0c817fc37aa7cda7381fcff8efa9ee87ba03a606d4d7da56bee1e6a5260ce83d53
z6b07df1baa4978309fbe3a048d767381a36b98f9d000cc5b02d00c2fec798e3df40f92a8686911
z04fa4a337f661252a40a8d28163b645df7fcd6a24aab9a66e4e7884ab841012f4fbe9291b53703
z975ae9edc338c421db58ab1c47e68842e8f956deb66e554854d59f240ebf1ddf2a6d26520a4120
zb54a866b2676bb132c68e008fee3fedd945af1cc41c200df88e362f6a2ea97b6e47d28d5ab4606
z80cc52acb60cbc6939fe017ac74c8f3dc13ecf358385aff4679b5a18c13b42fb13702ce9d50b16
zf3fc3bfc64fdb972fedca436edee57dd1a7721834d05a16f6c4a00d81e522523c2f3a36ab7b6c0
ze2d6f863109599fd188a7ba91c876dbf0b10e85a16f08d508e181e005debcb4cf49b43f3ec412c
z4f1142d26ae631b2f63e93532198a316c04f56b554cbcc85e65623e92e8c084b399cca0919ca06
z2f81c6758d054f3549ffaadbaa0c91b4b5aa752cf7b3f31b7e81c4b2f493d6d57aa22751f1bbfb
z8a17474aaee3289e1c6fc2026078fa514af7bcf171938ae4fbc373ae4b286fb66a32a189f4c7af
z3d8a4c6ade41f02d3f4c8f8c37134597eb25b2a3697029bab30599af9767532dada849be2c5cc4
z996772e9191320923ee8ad9cca66b23629d9525b89faa22dcd4fb1c34f554a86605fb0d2f01e48
z994d1c80c5e331210db7d2537d4f1636f03305f3c7ca663e4a555ea9ba4f9925ae0ac874d7b393
z3492745cb429945719141a469ed19a8cb2b2707f514d3cbe5da28244f7d576e63db6c7e12eb5e3
z9050c464a6e3aa38f0304af32a7b7b775f58a257f61bba944c7feeef3fda6dc96cf7c50e4ad81a
zc886a9f371ead348a54ef006e5b836134447f55da044500b217de77f728bb0a5cbcded1978b52c
z4cdbc586f967a47197a4216e6782a89fe6a9b1b516a685ac445ac416b289aefacbd8fb2a505fb1
z23b6ad743139a118ea64549c5be90e59371e99ceb794f940d1e0d76507104887b2f42b6205848d
zdc117b111966ff7e1a453302f1fde623f1a77dfc6eaf1393c8e9e2f83d27bd91cf60cd2fb3f499
zf62948860138181bdd95f49cbb755bea9b1587f32d5dff7a56d6c456fb20908d8d5a2b958708fb
z6aeec67da3de4d787b952667c2f79a78ed2ca4d52438127aca092bc0729b524632d3e4e9f587da
z6487f559a4b18877da82c65786c53316d53807362ccc607de0cafaa6eee87a232002451d22153d
zb45ed1903243a9ac7c1d4b880097db159351d9c55e173c182b6fcdb6eadd2e08ed23e2bf18e739
z38a8c52454716fe9add894c8fb43b5636dfe9d7397ef6954bde24394dee4585bff3c440f98dca3
zd49fb026729f103aa51036729d59bf52d8b604b8d10447911f1bc1d8b3e1bf70898c17ae4fb0af
zd6eeb15176c9232fbb58b60e1ee77a3ddef41a1eb4e62e5e8bf0ee2b5a4b6fe3a7b81ab739a0e4
z69a6d593082479c10866a8f8d7215507ff56764c21b8a7043dde71e3d94e1e4cbbb6efb6338503
z521e97b9cee9631c2e17013483e9470e5ea51b286a1e5231813cb40d940a4267e46c9d117ad84d
z8ec61e7bfad21083436da41488db3ddb7104ba6613b5f8d21638f6eea23e89acba7d0d1a410424
zb1ee443adcbecd93000828d721affc733a0c3a69636b78aa53a10f980e6de2882a3d0a97ad7ef6
zd7a5ca84473cc99a193161bfebec4d78301d9dc786802e150e446daa030421b0cda17807f41360
ze5e2ebf77138549cf9e063bee929ff8484e6ff3d9802cb67a963d5dc9425bb8c1286577d7036ab
z3ac35651b5fb1ccbd68635b2f7d87d6854d5f9c28ac12f2ca602f7a760d459c9b5f4e2f57efcc1
z63ac285a333e76b93dd4e2ef7022aeb145abde408f92e58d9d5725ccc8b9feec3cd418577143bf
z63f3efeb268503bfed31cda19911ebe65286295fc9ec780f7e2ed5306bab352e017eebc431a1a5
z505189feb80ccdf1d7e45853a64d6f6ae3444676f1aefdaed167f700817c2fd99cfdbcd6c851dd
z552870aa630a319f12e9f9d421f655b7168db07ca0db80a22afb776537ce1430beb0c9d54eb244
zcec03b9bc9965dc4e84d364dd54df1c79de3dcf648f90fb3f06ce511a833406b123e5ea57b04ad
z516b55a75fa22dd19ea52e40d3bb727ab9b4a2e3643320aa6155661d0d9399bb9ce48d8377b603
z713f5f9c70910d7450d3efe7ad011c356709866dfba22d7739debb4afe460e775e165641e0c8fe
z1be51d9fe8af96521e4ad1e60e3eee9bc7e57f18659bbe0883da87c8663f779f5e1e938eb1a670
zbe786b662a378f262e62549c2ca6b27a1c91d01c92550522599f7a82a7424460e063f12c7f4f78
z58ab3ea6dc1f1b1b179e785f8610eaeb23bf41bf1a2de29833f7d23fc802b02df3fe45107beea7
zd8e560a4e5c8ab3f37fb49d254bb5c335a8b9c9471aee3b71b49f6086db116a53659c96a8acab3
ze9a820cb464c1c18ea8ecd62a687eaf4847423738e6559fd8ee1dd2d9d32637e1aaa2302d1bd7d
z562eef27ba4c5160b4ca7e6c1c8656663a8ac9486f936d1ca198a85297b94853044b30c249f6bd
z0923d720728e43fb26cbd48f01aca34896174a130619ba6c2a5f8b28b62f4b7b8bee1e1f017777
z02ad6447d381fc6e29619e76eebfda48934ce5ff9ed3afdb9e9b915662d7120ca485611bbe024a
z8c7361f81ef179beeda54adfe1039cf39a685a67db27dc24e0586a935f400f1f1b6c433925319b
z136d22382fdbdf0553e41721efa834c10af9b6b8a9e0aa532787267f7a101ae83963160e5889f5
z91e2b67ee445a8caafe2ad4cda3629d1247bf53a33ec7f5f752ed7464bb413afb75f0e17ec2d92
z11a960a2e0882523436d24b48de0433e47ad2c4a5465f3289c83f2a7208cb3231c113988b10aab
z56383bc75df4418d08e302d601f4187b7f0af272843bb5bfb5303ab6a688d411a4872d08abb84f
z5a676e4283fcdf5923a5043e381b9585a7d20af111852aec7f732418a919be49822dbf3bdd02a8
zeede2bd0a74a07c5535782aa5a34a561ee86b0a6bcca8ace3b49376edf1cd64ff6487c2378a630
z02f497b9edf6b62fc6bfe8e5a2c8ec7f898002f93b47c237f4486e0f70d8d6803b31789cdf8b49
z573f5303cea8bb60da4ec55573b9d02cc82b4767e5505f84940f6ddedb9db5eebd6686dd33ddca
z813b0bc192e150c51df5b38eb386c81dd695bacaef08c1a3cc1e30e752c0d9608430f19e226e3b
zb1cd023bfd4b3c75366b5b6a324fa59959e8a8248196121f8711c82ddfff15f0888ddad1a8000d
zf7afecaed4bc480ed6e2643be991d15fe8d896afc9f0880075d537f8865859595391f6132a5bb5
z22023db7fa0e4e923141e9d1d79bb535398b30dab04111cd0be853cb4ba31c36a224f8681f2f9b
z25483e67234c5f22ad71eb144806079ec8f1eaf8ec4cda8269db2d5bdb3c3acff1f01bf6ff7211
z36b5a55230fc5093732ede5eaadc7337748e6f4dd77550b8b96c8df6fbf77b9f517a87643ad565
z8410bd6a6c39496ff96766b73e1c8a59a5e74abe20f0061ba6a156ba80f2809bc76b979200f7f4
z4c0bd48effea9c44752a60a791c600dfaefd3cff3117129c324cd003abfc00b2ee09e2e70d5b53
z8acf29a18d2d017e87f9e532fc0f0f4d144231bf55fdc007f8eb6cde4c42196f454890c7636518
z46312838c901e4bb1ca0d8d51eb1a1d9b0cf5b7464c0045cc016f86f82fc61756c05e5cb4a5e16
z3da1f6643d3dd3a92befd7ec8ec51a973a89701fe5972cedf710d476ceb7122b42858ac68b64e5
ze821f221cd18dc0cd15559a4a4463d96008ffc0e6f594688355358c9fe486f25fb64d36f60bd40
zd2439fd09fc403bde1393442e6f079d12a1d950ee3bbeaf81592899b971771269d97a7175d05ea
z35887f081b872d7dd4b877e48a95a1e4f0e9656f8a4055207c208aea0ec303ba35cfb856ce4b95
z2c7263c7ae26040bcfe57eddb0852e90fd420387f9b0b549b57ddabb3e5eed7aa044078c0ae43e
z3941461c7d57944d270aa12bed1b8dabd8e950c4301cb23c4a7b2a6d88ad659c343ca7e11ea49f
z1f534879791c50995384c168f4278884c0e150402a99bc71017f7bad02948ffe364dde25d64dde
z5328dfd65db434a7a75f034445aa34777afb56554982a041faa276792773f2fd45ab44f3a7d9ab
zf7b60ae74145f419176ceaa6b89e5dffd78b0d9618781e2415c19f16717fa98c9288e04bbb678c
zfa5a51697d3b9b9d3e10e2b00bbc8036790f0f74fc2c0e4593e19ca833d772e51fdcf7394106eb
z5c4eaca515d6e004849831df109732b5b530fce13135d736a9e180b470176b886726556f03f7b4
zbb2b82d9cb320f8eae725d4e6b04ba0e86943b87d37c9852f49a9b2a0ad023e77d3218478760da
z7eb6ddf81c5044176bd9065a84966d1c7d257a7bc505cafda9679f620b14bf97a3181866f86aa1
zd42aa30aab66423fad5cd64c8aa8c1740a248a9da1a2e79899223ead94bf1cdbcf8f0a7cbdb0e3
z78a0027ff96eff447b5a4fd55a920caaf1860cd894347609c087ef317135f2c3cafa487b8c0e89
z8d130c3a60e5d02ac613425738cc5b6a5871bdf6820b5f9125c92c7745e2b3d986db654ea80d74
za2445db6b5077ea3cb21357c79335f5f5436d3e480f398f7aae2d999d2e60f6adad4020499b3ff
z51e55b0b13460878423969b9b58b1fef0189df4c26150134b85829eabe089e4ac81a0b91633988
ze5a1cb5dbc55ccc8e8e873a20778e411e5036b20a98c7957ff0916328fdb5d1eafcb14b8621227
zf2d84dfdc55d7076f7276fa97b2f5d3b5505159103724000470c3471cec03f886d77b79fe86c14
z5c8623bfbcd300071d7dde3e3c9623338e424cc62228304cc6b05bf10d70cda6670edb75d72e00
za62dea8dec23cc8ce8030bd02c5a53fb5a860ea781ef8514baf39ffbac3260761dc22b2c1a261e
z0c9dff41ae7947e409b998edb9edbc6659340e03f4dae005a2692ffe74605a0d307a8bfdb89ddc
z0f9d194977113b2045b09d83c576651e272df0ad4d0f04f4b6a427657fe0b6316f4f469fd6055b
z73485ef2ef861c85639fd00c6d5db7ebfcfb76157c199cef66fc57e9939188d6bde0549ca49cc9
zc45ea105fa177f56041e9bc0340ab34664bbb131361e68b9caa5f1c9969f7ac0bfe2a99a04ab18
z17807fd313a30004eca2ec95c14569fb9b4764bc743adcc118a996cdd8405d67921763b057d14a
z067e972f08bc4601702736dfb7aaa1d11768a080da497ac6e92c5966652fd6b8dbf90bb048bc02
ze8f6646c312fc2c44d42ec9678fa2efc7511c2f16866f5299cb35cc9b9cb7d6c756506ef50f361
z19266ec59c41096d3fb63f24594a0b6d733703ddcfebba5293a9601caf09c774eedcfa9104537b
zaaeccc57f4e2aad0290f3c0dcce6fbd41ec26f2b8be939993a0aae3f47f7101047824962876eca
z52c8a402fc4ae2ef1027a24f0140412be62a27feeb849d38b3bd1b6195023bff905f574943d9e1
z39623f7a2ffdebee20a3a2b988b1564866da8b11f7eb897881ce25d1cd07ca17fc6d6deb5c4323
ze7e96ff0ba1ef026f5590898f0a7dd19cc1c2b795ef0acc120ca369a493deb6ac96fa0254cd9b8
z028e3a71cf48bc302660e2322e288db6a7d64635069ee91d0041796222511b7a1fdc4240e4da3a
ze494ddda6261e01da44fd03ab8e22e0840e7cdaa39bb12de449ac821a6e92c3b92c3a769de7a65
z572ed3c2ed27ee348244506c9ae32d0197e49cc6a1bf6a7e23e7a49db43aa1b7a1975421bf14d0
zc6f7122e0248d42af945cd25003caa57736bf38c43939447a31d753a59cb8fd3cc145dc2895492
zf718543b2b49b93da485dc4f485a640d84d026dc0c950f74a3d7e61dcf3bd8df5e9fa372ef18f5
z16f456e7e4d30402001312ea8b4abcc7f1ff1ec0d25a1e04fe450b68ad66044b4cd9d4f1eb9061
z2cb3c9232a706bfa130f185533c06385ba7c4893a47c0d148c7d1ec88f428e519bc17458827a6d
z3f124700137c0c1434238c6e28692b3929f5d0b4a5fa112fb529d28e5d739908b39c4af2933f87
z5ec9f910aa0716b0a6f07a4c3d984939bdaeba6ee8846d136e713e4d4f3b60c4114f995cd0dd58
z215e9789f7d84058af2c2774137b73763ba85961e93df4b00b074e91c0f2b47e9d1f2ba41617bd
ze2aa902ed891ac0f2ad6b35518b8a218b7436bfbca4b515f4357b7887079f2115c3a29c66f03c5
zdf6645afb5936c56d7c92d932498f5a7f522a5e1f91b0c2de46f65aa5d7ce472ec2967de76240e
z7325627aae971e266232497d59a2cf63b8629aaa78022437eaa9b95401b33e14ab08848a2f2343
zcd1603c1c9780fbabb6911e47886d7843629afd11bd7da3d4a6f13ea7954fdc42869873c30d8bd
z326e24968dccd762b31e5a81208d3796811426b1b4fd5411b36a96b76a37e328695b218332be9a
zf3db822cee429c827e78dbe3e76c12093f73cfd9e1cf2f521dcbbdf59dcee7b9b9d9450ad8afa4
z3897cb65de6aca754f6e49631b569643fbb70bb1d972596723b79b83d12f28f5fb44d37a7b6d1e
z1207bdb01a0f8f231964726982c30d00c7de4922417d8f5a9ec3675963bb1f3e06945f959f0b3d
z2f5eff3a5718023e3714b7654d51ea713abc19f9a3254b5ec13c1192b01f827a3cd1249b1fc706
zc31fe174e414716578fa2a672773bebedafb4033b75f931810511820157b0a1ff8131816165a6d
zb0b46469075b47b691363f3d73874c3b80964a1e4210e026b387ed76f2426a67c082b117230ebb
z44ac41307c88d24f375f977cc16ecc3a44aa73f7a7f1f65deea6a77cf75cd346fd74ed2cfc5763
z9d67d5201e4be4ef9ca5e4536849b12f219f951cfd4d03060a7c53954eab90f08bd1a4c5280698
z0c112f418e0ed3c108eec334f9bc522c202a68e8e1a2df5c66b2d8a6032f9a4d53f8d942d5f7e3
z94aa9cb4301eb749cc04e351cf572c867ac6385370f3cc2d5f34b904d6d6dd37e70361421f1b67
zb0e938da2419cbbd10f6ab3af118088287249bff46ee699a9fa7bbc28ce26b5d81ea9d7c493223
zfc690bf0c14dd4cd043cf04209a75cbf39a11d311fa1f3184569cc224d4686b6863465646a9e19
ze54c8c5ec767b6400d9a7a1eeb34609394188e0c2d431acf3ebeae4fc5e6051894040d091ae31a
z1b4641b649f070c64142789b618d6a8f8266cad01e4760a7671d8cd9b375ad1fa8be985800ef94
zd223b3a54f74582208a801f95ec0f3203dc8361d88aec02192ddabb66215bd54ddfc4eef518674
z80a4631b1d9a767b2ea86d3db00a1cb94a58acebe11260356341c67bdc952d962e9c33f373233b
zbcb1798e96731a97a2afa508886732af3fda8e1642038a40965cf795937a6eda802bcefb717229
z782ade367cca4067253c8da866c08308e7b494f2f9423ef31fee8d59b3fc3cd28fa9ed42c48a2d
z5c1b119872a74a89a97adc6474f29a1f3c48a8d844f369a758ba829cf270f1d1d84f215700cd20
z7d593e240f443793a1c8489e61a836a70dd61366a1c9acb185afd85acd8410ee2cea3f4b544dbc
z2ea694dee9c76231d3ccb81f1024928fe2fd322f047afdce510bca306d3193d959708e001b3f15
z098be37e4aabef86305e24967692ffbf889f30ae048316ff39322fbef2807460cf4560e54e0e25
z7db9934badd819e6c70de0a1e51ed03a45a17bb772da8331b3b41f627a8db6911f219b4b543375
z20bd8b98a1de0c1587d242d45eb72119805cfb307b751bd8a9ce0e0fcccd951304d7edc19b9492
zcb84d975f3f6dd1de2e1a2f472beb01b253f7402121fb6189f92f72eebec3823eb65d8d1cdd96a
z363bbde973c4b8270186a497366c44dae465b49e43c288a75601038064b1ec818f553c6d741006
z9000fe5c6b35e770b33a1fe1dc6b47ef1131fe2d6c87d46d4c9ced67aa18d1c041d08a6c7dcf30
zfbf7df007a6cc2c4e97f0db8baf700e3084696e935e2898170c37d4bc2a14ac39f3ab2dcaf9c51
z235de8c0ce5664e2aa9007aae4ffcddf4267b182d3e6db35ff29861170a52a0d66ab9573801455
ze37b46aa79fe360246acf2912e1497ebd33b85c9f59f1b48c9dabbd4c607bb927143b54cf6e1be
za05d5058d9f7ada2f4e97b44646f65d89259aef354c75be4f6bc5ad0bb9053729255af7cc88798
z008d240b4f95e86da3bf73e3d932769d1177e1780b17f9a9b1224231e5885eb12754fa17921463
zfafd3667107aafc6d2f77276faf71c0b8ebffb65f6098817cd9ac3a49d182dea7f22a031262165
zd2a31eb446c068c97df4e6d5e7cd427cbd1199893ab243d008726cb50272b20342db1875baf18c
z56dd7d00817be3128d8bbd81fc9d93212a4f9f681faeae6753e3ec8d83d16279cdc23b832d5934
zb4dd0f69a40010c664ca4aed5a1a1431039dcef956a8fad5525080cceb60024663186969f59a51
za745a17dc547e91331733959fdd20c0f4637b7086355db6d90647d74d301701b0d782d266868f0
z5185a915b6cee6e80abe975d259727d85a94bae75cd7746bead5201a914f9398d1395166fcd95a
z3b334b26c26eddd4de8819d1931f85f747269316d81c0ffd557d20f6f0f585a40bd0b82a782479
z0eeff46f00d101ac9caaade2f4ad16c73c215fa14c60a3b8726f8e56f3a8428ce32f01149d9a40
z9ad5997897cbf0d326a0bbc1e8f295c649dca55c5e692171d6a30047edf720d994ac49807a5ae7
z5c5374eb312a8fd91cb893c69568ba2fc5b403569ac5376214f9df70561895da8b5aa830ddd07b
zed2d954dc855cb70211974cefd596405dd9640bc2157380a598b893f2a11d7642d2195f0bb2782
za102df7af45cbdce9f96a09d47117609f2639480644959abbe1f575025bc4dd0ed1e65c429e763
z2d5d60e1364d4d667249d29ccf241345bc3b769a8eb54fb1471e5ef1d2ed2c831ef123cc30bd7d
zb0b4b6116f30a0c75ff044302ae613a4a192ea302c4475d99de673f216481a872ab906c1cd8844
zc614692ed077f3753213a236aeff9ba086210ee6ae7d27a47f07443395c4d1b93ad39390289131
zd7037ea58ebdde56cdbfcaab88440645655c9b8a701aa3b747f48176c17da466df0889b98bf149
za8036229db5c347fcd16f12aaf7e3acab0d4c597e43916544e9bd76ff8cfaab52d7e35f7ec3467
z449b8ae5d2125818a3517e9a0e1375489b0189a2fa71650a39acfdacc1047f904d76252234d0a2
z1e223af9863e21194dc3dc19f69cd39bb6d797e2b6202701f5af41594e1a2440978ad50a625707
z8a59c6601ea5db3684b671c17c098781d7500dfe23543c589e99d01647b2a13f16173c94a6f873
zc54433355a09ee786ee812da7c62a1915ac6e1eafc179e910faf338bb99ee8a7d7ad3796fb588a
z9eb9a95dba1ae20a9e9fd08c08d72f773bc3f86cb0a61d7e2783c45707505c76fc4245d07efa64
z27bfa9d49722716e36ade885c820ae6d780b7c07f5f8cfda2ef239f00ec46696de0745e169ed5f
z003d3914eddf9fa2a6ac42761258dd21eaf3e25602a4d9ea1773dcdcb9ffafd247f32d53119016
zadcc6efb0b406695a0ca9e6d10759aa9e02ed43c3fa33c3d979105a0bfd0522867cf8dcc5ad2c7
z7d4a929c135d2443a942e569b75ff2bdda620545e0d608bb0801292cb3adaf548ad0125df968ec
zb149d48a24877406bccf624f4ceda458571525b23631d7a64440f7d9971bf4e03e97f3879344b9
z1bddf757cf45b5bcc9798160d4cd2651bf920742a7e2f8123f4d88029ed320a22b945e76e3fd93
zc815b78e71be96376dd50b37fb6135ff6eabbaaabe19b3859f9885fe6051b4243181741f5390c5
z44092035075bf29bfe9f72c42e66de50656b17b3b1dd622f5379e7f62231402bd79664dcd048c6
z2d50c41e1737286a736bd6520565ef3960fad38b33b24018caa402292a181b9c1d69b3408366fa
zee05ba4866d414db8e9265e4c458d1bee7c24ebe771e2023e18e917dd0d58d8496a97fd69f971d
z1cc8caf21165e1681ae3dc834fa554b07f325f404b401b4ae0e5b77657518dc4a7a71f515fe6ca
z5606d1d3bbd6148399dc5399d21d898526b88a4fea3f292f88467b85ec11ca0ec72bdf4b955a46
z350c62ddefe8670eba8faba4a0642eee6be6646947d996e9cd1e62e3f453c4143f03c45fdd26e0
zd77c80407436b628145e88f311092373
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_data_used_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
