`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699166942afea5fb71013544a379d857e146892234d38e3a5
z4d7ba7c62fa3a65f2f4d7424646d44b510488254a74265698a7d7061e59dbec7c6ba2d153ffa62
z9bbdb6b0d94277ca46d0799fbbbfd05e5840c76a44c76bb8827cc70fd94aeade2e109c923d1800
zfabc4556bdcc931c4d75a1f77e2bdb07e4b5791f120f631958203c05da9a77d6b8e1bf6b79359a
z3867a84688be35edcfca5755f9e68eb0fd78d231d23c41965723f0fc86a46cc0ff42cfa62494d1
z800bfbea9764ab39642a354d0afb1e579af2e5c001982f2b3e975e5ba318f3a2f581ed37f38a80
zc76af5372f18fb93935913bd7c8d9c9bf519a32f6bf92658356c3f478657d5584c5e80b7684085
z74f8f041a1934a4b483461bc98df97e0e67587f1df5140642299954a9ff9286bbaccca2303e1bd
zb9a41b701250f7c71a330e5c2348325991513a035d23151d5be51498c4bbb70c0bc659dec2f66f
zf3d0679b2478484e3adfe5c5920e8823d0f93906e4991d2aee2b266fb4594e543bcac71f972650
z3bc9b677abd4e007e7e5ef3e86b183228ecf4d23a9cb90650922949608a704f2673b1efb9e289b
ze60f10cd03a5d19536c0d3f2b78249e2d85c9b7edb06bbbf0a4bb72ea6af69e181bc534e3a7c96
z545c7a3faff1e5582096bf20684132d5406f906be4fbe2d602e885f14806003956053e4f7f4676
zef9cabe44cda41d12acbd88b04b83d78c1f7deac7f9eca38fd758de0e91c9e00a89324907288af
z3cc303d9f263462ce94dee2f7868ef7a9b381a8479a4216003071bde43eb349cd2a0fbb2ca5573
z0e622674fe8ef3fcd4b8ff4caa9c5c4899ab6d4d312c7c6228dfe09527494dcc4700a689e39ef2
z0dcb2b7fd7d11ed2d4e9ff0573f496f7633186513b4384d18a1dcfe0676276af02d4d4a72dfbe9
z2e2e96c0abd728fe9f5c1608f9d4cc4fb73d3816c8a993dd712ff89a3e20b1a150d78bb7494c0f
z5ef9ce037de29eb7015ba41202ae5a5b39482d3d57bf971c9ba76d8e13f47675de0b5d627ae081
zf600ac9e83b51377dee54415edbdf6cf56a2338e952f8a6220d8a2f4dc2b5f5e8d5202efed85dd
zfaa63da36b29644e36cfa6a199f80f733dd7b0c199856eb5432ea6b200dc15aa79e4be3e1be932
zd524321c620ca6172e4719b47dd1729a9f2d837cbef1ced48b2e7cd4ede9eec829668da1f77406
zb3e9cbd8448a44cb9ed29625788659936ea47cbadf15ee77b5c09b42452893e98d10620002cf2c
zf857134d939563ab622e5a2d85add5a2dce40cc83fbdbbda88c49a04ad7467e069de1cac85f7c0
zbc8a16d1deacd50716e8c8369e74a1d2537d3b3fb0fe8bb31c47a16b98958087f28230b1f5b164
zf6d67ca60a64fdd531bac1494deb8a46079b0a8293305293a8e2ccab14d648bd5cbb7c0a7e7ffc
z9fc964485020c07073d33814e03fd67f91455bf2c0121ce0cf3d5516e0365a804ca790de687ec6
z8b6473ff7a8fd53bcdb04cfc1dee13977c1e3581b8c1c6d4aa30ae664e83d53e76e2fe1c4c6677
zb7adddb060e81562200a53eb2583123e8294c2a687a6b04d7d8ca4320e981cc3521d5a538d5662
zc00376284072b4de71b2cbc6be8066b27a4b46389eaf49cfa53debf1f606a28560e595795fee24
zfc5c0514c7d1a414ac990bebef67b119a786069123dd1d22a20c1eaa69ba530958566fdf1ce3c9
zc97a8f5c78e007a7984145cf02cf3845af349a334756d5735772bee145f2044d1b2fc4a0100b96
zcbde57522e7fc26de2c7d8e6fc7867cd84ee965cd6259c3fc365118a6a9c618d626edda0ffaef7
z6bf8a59f1e4c4c668ee7ee539efa4d3cba0563bd5517d76b83bd2a4f6fe72d0dbb00d9f641e004
z9c86f848c0cb97a8d944c5551f76aa0a9d243d4b1eff256fa1d2773fba7e382d0b3ff12673e940
z13d62639f291b3ac2126e55c0754da8093d0e2385751149ec7d67cebe6879f2c006b9aecddc3cd
z74c95879469d42f485c9000dccf5d1c454ddfda0e1c1960f35a1363cfaa962657581bd8af45ce8
z92226322a95e23d7e58a4a99332ddb7d414b27193a691273b15ed8c9c490bac983459a9973e45b
z11e3a12973a86e549a7806efc1adf7ae280c5b070b0d9468cf9942ca3a00676e8273e542da462d
za7e726efdb7c1aca9e3be67f4d8ce749b520246fc64f6f21a673a5fa7d045db68f316c90afb23f
z2fdcf210e2af6c3284dc52d9af2d8af2e16d54162ad7829d1d20e41f0e8ca95611fd7dca8db38d
z62a2832ba63712f517dca21c309a652e79ab485359ca43f0ad491fc569cc37512d49ecae21dd2d
z55d5f17f482c1f9c933a09ed969e78934f3db3b640db8e0d2110dd30f917de57f0e2a914bf60bf
z8bca398c973a63cbdeaf3b8fb1589c09e6288888e188106b7ccfb3a90ea2b5af32a84fdcf3fa7a
zc736eeadac3281131eefa23290f85fe0fe1aca3923a223703552fb4b80ce8ee7046813622b2637
z634dea8a09339941f63347a6943fa372628db13619baff2a47b840e8af6f4296c90363518f85e6
za9eef9841924bf10103345fc620e144d4f70e977ed79b0f7f604953c78ba1fa34b8cf04979b31e
z95a82c6108af449965f81ca0d1be8a43195effdbe2e6cf3bde43a0404eb4b7d345a23d51ae85bf
z653f9ac655dd0bb8accbe40a1092e4e23ae67e84da4eacee3b67f6d334c7433a182de83a9b0564
zd729412e9255fd26fa4c353517a148d2374d25c7b3cc4a964818f1480847a1cebdf357c700e767
z88d483833b95465dc9ba6830a04991d673d4cf1a645439de02f4ddd4761d71dbb67b9f7ca5d7a8
z5e31bf9db9396f0c8a45fdbb6aaa84347c3261c30791cd2d19b805641609ce2b787c4e1dd8e868
z479da3963a337cc4ab9fcc2098d9fbae5fe779fe3e3bf3cf61a164783e243eb13a9d0f5d5d84ca
z2cbfaaf994d8347b9294014f605c11d3ce0311101d54b5ff2ac925be074cd4b102e5cfc26e774a
z5bd9e6350eec51b414c3a0fe864aee301db6f3378ca1d82a46025dc09bdbbfb69cd044d13471dd
z5e6ac5aa9c08852d5e8c69e81b0ed2064f96073959d6bf7e71b599c8d4a84d503c4bfdc2013836
zc6b415704bf63a8c9525611c78d8c0e9021070375f38babfed0c4f45bc01089af7d511f826f229
z3a995ef0befdaa66f24c6bea5207040d5cd4596de0bb388b7c7e1148b37e74d4711e3764604186
z0f72bd7c37abb10a01aa0c7b961371393414db900643cf12a919e910e5452e5b5776eb789eb7f9
z69b0acb33011c31cc3b19de6d1de15a64a41911a7b9fd12e7e4778ac35e8240c1eba587579e602
z57081debac0d26f126d3ad79f3c497581a3eacdc9290098723c4479fd611e3fd182e865442243c
zb346599bdb312d3897093205fe97801492bac29271d7d5264d738ef2f94e9d7581b9ae828321f2
zda8c719b823e9ebafd3ef4c13bfb47d6bc57e9d2d0457875236e80b0826811ce1d78d6a9969f68
zc96b64c2080746b0e5110d825aef5e646193e9b4ff42adfa0772a3ceccef98a95dd850a7f91abf
z930ecaf0205ebf230f78438358290dcbee568bdbef2a8fbdf5e0ad42af28af12b0ecebb44c34fd
z02f20425227263311307ef892f21c9346d4c363a93d4ae9728eacc86d6e286824b83e1a275f29a
z7bc63fe46f51c31836245b3346344ff2ae4582dd6e2535bfb527f46f462dc7badcd0dc04769582
za27c4d8d1f08b7a9e783f07486bee5f62d4f16d767dd31e18c7c135b6710cd0349714f726b172c
zf1e35e5f98937ca48a27ec6efe84a485ab046cda2d3ce4cec55b2de4f2473c10a5dbac3b33333a
zee78ee810262dba2e6a2767d0f797ceb296dee0ac37ea069096c132b4828404821da45982dae5c
z2ad3c286ed8bd9d7ab0c72e4f202a48c501b3140bea0e8290bb1ddcd8292cde1512ff58ac2f934
zbb9729dcb34b197c41c9ae6c444b7f849361fd0b13ca149cc83ed5c0ac57a2e2c9df517b7b7ffe
zc2842ca03bc7250d3533b60070c419815748d8e5c49a0d67e3678c406d508b7cd9d2ebc0100128
z81e0cfabe0070af3a188dfee9b8c429a27552d1f9a96be15b64021e5322b316d13d5061869792b
z4454706f7aeff6d1ebf50aa34e7cd7d72eface869ba144dd996ae5dda2781f9ab4851c97bac7c1
z1cb2d4d92c7697eadca58830587e8e081ffaf68a2fd591d3b9d9d57088bb8b951f502d2b0f4b76
z83accac76c64cfaa5cb44dc35db2c9f5e400b7c7f24cbc5eefe79eab107429d2eb431c5fc89b9a
zf5f3715b3e0764d65f1a2ffe3c8cd5e296af1cc65432c25aabe6aa4d15aea44a05806ed1ad2bf9
ze46cc4be595f4ce35c8e6430ad45a4a89f08812388722607fca508c3685dc135b31efcb6392772
z88d1d82a0f7c9ecf44dbed78bffe2269f04ac80e1161a9a0dc59504fe233320579d72e51f894e8
z22899b99d560249ad3596a531bea1f13620d7e74657a124b1a2b5f17f0c7488649e467234f8ab5
zbf12ca9235af1d13288806d87b97f87a4408cd49db521dd58dcc3841219b9b301e5870180b3b81
zd131e8de4f79a3ad8de23603e5320656d2d8ac1b9c87e351c94c719e7bf6880515a747f6afaa0f
zc7e0ebfc22ab571f20fd6e424bd18a794fa8c78a78da82136681c90a324c8be25dc301534ae591
z53e8fbcb1c2db191a51efe3082f850cad4814c4e9ca958036fad677e13d70676dea503525270be
z9376bea147f16d486dc091eb4a27cf91d2d0db516cc725a66b0497b19de665222cb16e01fbce9c
zd3d4df6cb193906566bcf37bcaa2aff63fe43d4ec7497e94c96ebdbcdc3ea1424191e2bd0200ee
zc3b665ad6bb8db48ba9b5903f6eedd598e0c684c7f549378ef94342acba99a98a6a2ff92773c3c
z335ddd842c9fd9d20012919540ee593e5963b8bbd105f56d96fe66c84360864aee55a338441b9c
zb8a2fad93e8115be0b28e801eae0f05c84d7d70047ca55a87f22b5fdabeb79f85e4db9cd5dba76
z752f1f6ae9fdac6063ac5217afc873a6c79e1826e9bb8c00e79fb859f920150025c5e752bf28e7
zc28b4d5df4930b4dbee77d6830e449c97ab480538cc0535342851c75ee8e9487d885183e2188cd
z713e23e31baa3dc8e3c10a7c74ee8ed54b619e1233b9a39f05a8fbd833488c0996331fcbbd199e
z79cb3ae09369bf2e2c8da5166aab53717530a77757905b81acf7c62647525870783db6c090e36c
z64608a10845c8ceb767f2a8e1acae6833c8727666557369679a2e235a88f8321ea554ea6dcc379
z662631f8bfc60924c483a83a1501ef4920c9c2ea32da1ee455484620874f7e285892aeb72a7887
z515ac5df3156d7f0c8527a7b84d17ffd07575eb3f5bcd9e699fc5dc655ac056868d8b611d28aea
zaf10e09e76ac7f7aa30f183da7ab582318e0fbdea7344e582570bf263f31fbc6c1d398924ac00a
z2057b28b843edcf6ff5bff943f2dd321896f3423da66e19260b2423b83aef2fb1798fada102238
z6c30553093e984e9ad8c4560764c7fb7bfca782317a59f519379aa2e3e2ae62e9369d05f1c65fe
zebfaa59d0b944bfa8cc5aee4236bd6d1d613ee5a8f384c700d42831a1d1dd0b28dc9767c927f97
z30d43ccfb3078fbb54100f858780ec75db60dab2aa93a3df4de86a916c83fa45bdb36d1cf23a4c
za652b8952a4eda9da9f9bbeec22a78b4b3b0fa34263eb2bf160f5d6c340d36f3283a94bc5e1c33
z056853b526465db519d355547eb875f5ccc7b283237a2e5830c1813b0276d140eb06b19c54d5e7
zb4692b818e1a1a4d5dc9ff94fb136fda6357d31625af877a58aaa0c364f7a1aaf9e41e5d7b10e8
z4425628398c6012209edff192e6ef8bd390688ae4ac417fce88f0ac3bcd27b90764e4677bef0c9
z94017bf328692c7d408d8001af51a1be6d221fa3e4b2ff099679900ba8d6eb80b767a001722e23
zc2ac85a34c13e8164ba9680e4dda9796876433b0fc7aeaa384cfab2a9d1222797c8d800dec324c
z035a711ae06366552f2a108dddd386b17a597b6ea91926d8f52515d938b6fdbf9798baa4fc104d
z3de232434c3bde65e53467278d85a23a7f3ffb86fa7a4f53092730658508fae879985274b624dd
zafc53de3e3f4582e4135a99aefcd04e66813a00644a189a80baadc5254fb91e6a8d2c716bfc96e
z9340ceb1463273bee5e1787092f144dd17f36c0c18c3b767524701b8d47163da046d4b14f05ca4
zcd1ef8e26bd20a486a3d0a80ae172e98183d8a16c2fd6e2a29bc7221ceff48616c9d6de4017ccc
z63a83d9f5c38eb6cc588af70957a82225edab27c3a6a1fa7ac90bdb8b282d6105affdb70099dd2
z9f8fffc02996f6f914b4077290471ebca8cdbf10f0d43002057894b07ad7046ddabfc86c31d370
z704566d66b12fd52eca0f482ce5a47fe52c619d601f2482c970ce8ec823449582b619eaa4396ee
z749ca3d01e7b6f10cbc830bf05d52e67918c3b56d9bd532565a5b62b038b7b256dc9293a1ab582
zaeb179d3da0bed8c5c1d7c9953786c6b02bbfe965fc8be30eea47322e9ce2101c89b9d49cc7a9d
z28f6ec48e3018123c3b66f32cd2ef32c31fdf0d6428236f2067f17fc4f963530d4426255452a21
z26cf18fcdfad905d0334c55c2e79337a503482ddb6783d3831d7ca810f4dad953910d908bd6348
z8e37b99b8d0a7f023ab91830e6cc3ba1f9ffcd0e49bf02cc4f66e5dca2cf2f3c957160e39a9ee4
z8583fac03473ee96ff34cd8a72c6f950984d5264ad0095f119af37aa96fcf285431caddea36c1b
za31b8fff977dadf8b7396049fa00c9d59c423de517c7b998b2c10da6a7df892430a9502cd0485c
z448f655f649198eac58dbd0d6f0309ae4d95acf87158dbccf7296ca61d4c8b66f06d8431bb93de
z7b74457483ae20192eba162509ab6847cf6d2006bd16a694a9b2f216ed1f4c64312cf9caaf87da
z5ced0da39259c04d8eaed3f1c62f9175deb8178eb1056cdad8863b11f882c311da272ba1fc753f
z15906f5311f21677bf374c136fd4743e14270e4cdabada23ca853583a40688e2e3067a702b94a2
z4348a9fb4a14bc2b0fc7d3b9d10e337dbf6aefda55384a569a79dd64b034fe5e66d44e4fc7c213
z6d4a6bdc1a84d548b0c7e82e8b5742f8dfa2d6b70b27e62285a251cf374fb0a03f75847e476fb5
z97d1a1f13f9561fd85ff2c3f63810f33e9b2aa89eec1a60e0f65a736aeff4a5f8cd003aac588e1
z9904734a416528e6b7fe1d85807be7a53badbf1199a93d3998b3a1cab6263cffb017f8d06c841c
z9a3976072bf243dc61d70c925a54d76e4d6c0a815121f3b4ad41f5dca53288a6c34b8adddd5f6e
z844bf0fd361de2fbaee5cca9b83759b5ed83ec8fda36fc5cb76bab0da5b03e3e7366b11a8753b9
zefd1989bc4d4e902d91e9e3649e3793c984f76584f1baee2636492950c688c37fe9b08e371c16e
z0da92eb0643891173e3496e03c4e3c1a2f35a96cb164c99ece71d6a2aa93e573e939bd249cd6f3
zfae1aa7e036df354d19aaea59ac0cd57a7640d8ccbc08f9c790af6da736286ee419a5461d94548
zf1d3046b49cc28003c0353070775ca4dce9c99aaf99cff994a31312a7151686b8c6ecb9635a2e2
zcd196237a71be1665ee365f897a455ef2b5b05ed50439d552b77cfa6390e44af9c7893a676080c
zcb0b3b2123850b29f9a1a6abbd0399583c89e1732409e2270933cce570373914ddd9464ea3023d
z4bfb0f84fffcdd38750efe3012d11b81ef90d6e4af8d5792fb65fee3ad7d39a6850c902802c318
z6a199683fb80edd03f0c898b4b66de6f1e48e7948cd6901d9ca9e2a0c04d0abd8a6ab9ae8b396a
zc589c74f4d0ab7cc55573bf533c721ef60b0ee5d0aa87137cbcbfca9aedcfa3efb112310396625
z5cbbab8de36a62aad3fd4926ef536d28f6b29bfee875e6cca8a11f51fc3450a9e26125d91f5fa0
z8d95d431b820644facbb53acc0abdb11382c1a2b079678a34db2a776a77ad024dff76a35b27b79
z6106321a397ea6bff5b243871c78850e3c28f2b85f0625c2dfb07758101a0a8e3b62a64f8db0be
z33318d126f6391470c2a80d376fc1f4cae3a195f3dd8ae427203bdd4a110ecd02458575c3b1ee5
z02433a2f9d4707aff94fa9135dbb2eeddd2660a7c7cc969a1ae24f5024ef2cae23add03c56d1ab
z497d309ec5c981aecc156b200405e34a3fbb326ca31ba65fa0d9634592a8b87a6613f7a0b380a5
zac4196d01b2110ee79861f2aa7264ec985bb0cac849094c7d998c5b9423b8e0ce0aac80ed7eb8c
z271dae396a36115e24e607dd83a77ab0005bbfdc3f0b8d25d5c1374bb5c0d234654acc49f1f47b
ze31e70ccc565e7f0ac2e190ce74b9ecc279de6513564289f11c3411e7d3f31d4055988654ff322
zdcdc36c098ec6162d827edf1c77e26e20359a1a23331ca511befdea4de22001c75d2053325ac55
z26f1a9f3d42613addaa69fe026303a9fe7092b47c929435e73f8227d58a97c3d92e3e397a0ee91
z7c059fd3a456f78fb92da9b7053da5d8e7579ffae2158078ceef0d33f9be9097595362540b9575
z6768cf648692ac7a3deda648c5780ca9b68444f8a1de33404a17ad876bee7742f8c44a8f9fc207
zefaf68c2594532d39c20995f819248d84cb1463342044a1ce83b1028957b945fcac63a09bbd3f2
zc5801541e2b0cbfc6eabe70206149097c8b9c0fa6c9b7385969c2763d2ca3cd84edc87b6417642
ze01a8cce4a20be959c619aab5e33afb41eec74fc6729b947a3cf3be462acc58e463f865021f260
z2913e8bf30cf9dd6205208bc7cdd4017ba8d66c3533dbdf8a0d9e1c3b62f552339b0ef53895885
zd9927ff27341ffa55adb255deb8ff53fcc892cb8ca13f309aed73d84870f2ceba97a04cc92f30c
z056a5f98fbcb32e92a440bc5fc1917cf86552a8e8ce5c0cd652aef7544c5511f7305345e07f4c8
z72a1ee19ed428f16da38c0be8107423c09c4a425466f1803d394f73bf5c765936037babc8aa5ae
z27b80cf29f2ada6d5557bec4ddee19051b11958eecf7097a486349b6ae5783e60da7d4c8775e13
za497d9655a60f46d17640faeaba5ea65e0182f3aac05f2a0cc480d7a41f8b710f1403f612352b7
z3d5adbf2b1edc6eae1868fb524d9fcb42987538767fb0b19166b4b47b30da4b7413272c96fca18
z53e224b75175c54ed0b39fa674b275ea125adb37d7cdce945360adf84a221e78c75f2a85e6b205
z76962242263bd95d84e2ae11886c41712ec31c9ff8933672de5200489fbccde15879cfabb32d59
z305236633106d253fc9a616155ae962c17d4fe0fcdb670a4688373641d2e8eea1257a9a97239bd
zda790a795a003cac8e12082c9384ac9e4fdc79cb2ee42b4cdd6854a184b114a8c690a397edeb06
z54dedd18a1bd2ce49027076351a1c8f94710ff60ebc222926ad9135d4a493fd822b1776bf76abd
z7ba6b258c1e663b34ddde4abd38b7d28c3b3ca6e7969ca4834fb739ee1b3228cdb9c208a91eb70
zb4eb796428079191350ab260713233594207b31079258268b20db014ba7655fd74e4b1d554048f
z95e0307c06955ed972af7de9b60da8adf8f62410b22f39bb9fa0cd32e254d1003b0c902162676e
z55be1a1ec166afeb1f2870cc5ada6bb21a8fdc54262c316a620bc963be0cda74bd65fa821776b1
zbfe03aba0cf9c37f90017adcd9a182461117777d3d7a0847bb590326902b5cc58e638f046f95da
z7a0f5d4f5b606bd452876cb47878cd6dc21aae3a20292203c0f8068f700bf1992bb16771207f0e
z426796f1a27786826068155ed35c8d41b7f06e8ab1be1cb1da26447e273cace4c4605e81fa7e94
z481c5107e18fc515a39f6ca181e15b0fa5d4a43a70c8d4ce05e28126fcf494aa8b6c21fe7da8b4
z7d5e647bbe743b41b3e97f778f55a39522909ee90d4b701dad41bdaedebc24e987a2ea6bdf6874
za0c412568c05560dbac527a0017e589eabcb02bec8081080a6537507b349d5ba9d7e521da287c7
z779a9784b906efa9fd0a5262b2372fb4a75488b7860bddb64d4dc697b50f2d20ce571e6e78012c
z8bb9b1f46eda08e185add5f3abd9afd5b20634b02c6ac9231cf0392f42bdd3a4aa73fc981695bb
z52544851b86a66df52cee0704a50a5947af6a1c6560c7d51a3819cbed345b766b660994c77f432
z42b91e8b71233e9d89eefdd7855f3c054ae576a34b11f8eff05925d86605b0b3f87eb6851a7736
zfd183ee41095f0973bd44c20e99008754dcc0cbef2698a08988e3ae8f4f9759d2150b253f00fb5
zd21e931079a236bd33bf34b94828a62596f2f97fa05a9e589e6c6ec8dbb76ab1d701792f149d94
z761cd991137fe6837d9a69474729707979a256e2311b0c7e0a14b0b4c57ca96539f545c68edc2b
zcda7b8c24087a58286f03d6ace8e35b3f008d1ba087946dd654e7e07e037671a8a37428a911695
z8b53a3532a6e7750b3ee1f7065b45f3e0d6def4d557878b0cf5f8388d5b27966cd2c49430220a9
z113a864b37ac498f729e2b3454e08eb1ad0f3af6fce024c89c5d8f7d694c8db88cd672f82aaf23
z1ed8d5e5675ef388316b95a687959caef5502d9e25b2e9b46506d169794cd3572a2549ace5b398
z0ecba6a91ab8d7d3daa94346bffad6ee0a0cdd0a42ce4110ac42d18f30c1c68d12897bccd6e31c
z8fd2ac1ade97a6b54da0c4fd9da686c9f317f6400a575ccc7bbe50bbe4d3e2e443897490958700
z7aefa03ed62d5df3f4ee4bb0415ad746ef6a3e32bbabc94c3b87c32b3f77b260f974e624e5f022
z821b6a7b7a90463f7209047db5c1f17d1e67fb9df6120d00a9ab11578512f9e0db60447824f3d4
z8c27b9fac62d021b729b753a82fa56f4a96ad355857cb42d2f7e7ef6cfeeef0da8351ef404ae05
z233a093b2d6630781206f5a60c714472f3ee8a30c5678d371bbbf3f835d658bfb66212d27e8118
zd654fb26500638e9bf572c093ded1ba82a1b0333682078a2f7d819674666d47dc3dd28ae30e144
z776254a1299c900a03897286b0119a199c151e5b83f68702b2ab13e6b4323edd9f7cb9e6d413e3
z9b31b928a60939afece2984cc480ec7ef94389c466a9e394902aca5a70b8fd8e6f2bf403dcf17e
z26aa5680cc79f47f24a8b873ba65eb9eb04671fcd3bc5c321dded7605cd58a657ca9696563018f
zcb1d20b286a60c66d28a08673afb8559bfb42f7419291d64d7ef4ccd09403422687954f042d303
z80ce6bae01f23eeee8c577259e93d51054533db7bc47ee86bb3b5ee19b6b896438ef00874858bd
z94adbc22713a46b59070a5e009f774160bac6678e2983a35f832d696f9f2c204b3fd7b5340dc4b
z0f91099a6f8569fbd9a1b3a530c0d5d5e8d03a9241844e26f354ceae85086f248b2fdfe77a0a79
z9f2e6b0fc920f826c455c59b8f0bb64502105e7539840da4fc14a10d7618988e6779d986f216e4
zec5bda6f6f2138d0d753a19fba68198cd383862cd9f0755b3a46867eb53bb841a28cdb9c599d03
za0e71c1a550c4ccdba4acddf9ff78af120f2b34b56f17349250fbc80e528e66bdd6bca79b5d5be
zae54d04b548ac0ac2df6414d62b8a920840c8b9fa733bf074e94fd123f63b7d8b5c85c9b9a2c59
z9346ce7b9de534546b8ba11e965cf76dfc68734149bfcf474e1a0979940528df83f6079785d45e
za8a544b9a29b919ec9b651c8a3ba90fc20374e908c93cf0f4149d2893f76cd9f82a29f64dd8d42
za070c226a5ce0c520e9941c3646a1e3af482e0c73bfe4660ac764de96fd7d434070612cfb34611
zc9cde0ae6b35b5cfaf2e91dea0fc7d2dcb5a8fe1b59882b512ec8b3b72653007bdc6ad647dfaa3
z18f73e93bcf637238bf9d5a4a1f663595b30267f3d80777aa43e83fa9e6d1dbd044a29305ad5e1
z0babbfb7a7b32cfcb1c47d18ab5f660bb7a84aed36c32cf5c29e0c8d56041508e03107bfdc9317
zb2165a37a6aa411e143054a724fdaab9c69caad591fa7a95196ad591942a1e8c3d16b77cde57d7
zbcb9c26a58b8c5b7811eb095d1179af01554e0cc1d4ec4e352dba27e0ccacfbabcea441ddae90d
z9b206e5e20c06fb401cbbfd05dd374ab75b229e30491d8c3ad5be9cab5144db80f1b7474cff111
z219c03bfe6dc48e32006f1d4643586f173e45d493befd060abddd391b2aa6057304533b09edfa2
zc71b3652d0829c109680f5792cae102aecb1adcbc79120eaea834d9ae2fe8cd75f595e4d378e10
z20aab9641e58fa981cf4be7f2ee78f4cad7128cc0d1db751c36a37d95e256b45214f0fe80c0e46
zda006c7d84aeb72a6754b181f53c733dd54ea48d110c9f8c5806970328534f06571044e493a992
zeabca6edffbb6f93b0f3a8372552b7789715dae431b984693b4c9b20fdb5d5ad8d0ee29cefccac
z52e78b435e554a8359e6d00fc40f6dac2db30b69a6ce15cfb6039231b3fd3d77bf33bafc48a75f
zf8d8d1c742e74af486793da0468b8115ab0796dcbdae84b56416a2e088e7ac736f865f074a8f56
z411cbffa207be5f79725a0b02e9a2735f74f538af0ed71f7332857531b747b5b1937ee665ab750
z2c266d0837a63ed118c40deff418226ea4d08da55377e64da1efb989c67aa5eae9a5318cb5a027
z667286605176d24ea89245cfa99b7df758a9f274e5343d1faf18b707ea301abc1b28cfe41c3b49
zb156c900cd86629b07b9ffede6aac6f565cda90109bbb55241e710e98238558d8d9788ea6c8511
zabd5dbc9b5eb5e3d9ea2130ab32bb9151e91dade0ba1bbb1299a598b75c38215756cae7b8e256a
zb7702435b95155d6350164720d35bef48ae0c80dc08cb4f2240369c60be7ddf6cd716e3a61759f
z66dc2bc9190e1d069e95e1c532d95b11f7d9873c5620f07cce0d283153027273c05563181b88cf
z1a70c661cdaacbf38237c0a72ab03be48cac90c29a0ab88ed77669eae3ac030666edfe3b33272d
z507e62ca6055b724353bed49c954ba4655b21a1eb58994ced6cc70f463266acf323a12805eac10
z6dad2cf79d7d1af88f860b326ed82f4b395f793826751ee62e809e5e6b530a3594d160c9a33e85
z13b452e27db932ca7c7bc9f0b22303dc3120ed64378057cea3672e6f366ccf0dd63a418f4ee557
zea768d5412b30fe9dd1802417cd6337dbf3300581c3f4ad25a87721e2fbd566ba1d000fc40b287
zfe66586ef1a3a429165c6693850d77b2d282de146798dd4062c1381580d7619ae97d8be40744eb
z3b7519b5e269c074ff09a63d1cc0fb65303bb52ce84762cf415c4c07319a7a9c8be00283b7db1c
z17b59f9cacca546d1ff19034b7977d74080a1ea3cb08a3109cc1c6273e37a18cc6cafa01d60f32
z3f5db34eb30c209c3ba2839fc5ed45b58239ceaa525e4403e45f9683b0797bd2526137da08ece0
z124cb23bdaf84782f7dfedac35a7b1c8cf74e456c020f7e61a293c0d32cef0248994a0e4a684f2
zc93f2459537874cf2a93452f262557c584b23a0159ce4e5a368bda1e5cf077a3bb3c06384c6fe4
z17c48103702ec3c95309473b22d2f9c4772fb1e88138c653bb49e38ab5afa6d63b8e58c2cd8a12
ze409c48e9856db837c4fee57f60d335a4cb3575ed3a03f9f0c2e24aa31738c5e04ca5e6845fd8a
z3cbfee192607ced304c83bb5f67347fd37262b678bbe486a8740dd873a336d17cbbc023299af5b
z9409b11571612d5ffc984631ee8c1b64ea1cd204c577cda974a5e128cb5289d115fffeb2e084b4
z3b0db22f1a9736a48c1933976264b41aca3197c802e2853ee7b9a3cd1321dda49e32922017db6a
z0758b0b41f5f2e0bcc83ce7c8299f32fc3caa03ef7e2b2c3db9ba457e517c098258b62713266c8
zf4a4da3369bcbd7e2ed5c0d8396cbd7d99bd7b6371989f96cb45c44e0cd4ed5da38ba0a4c57cdc
z00db6233e7909369ea0aae7dea6e4b70200837d625fa8dd5a9e6d99c3aabeb04353b04ddba6b85
z0332010fc72e09451eefadd53901be69c33b7e8bbd39327a2dc4c7f9a9a10df33b5b754c6c56d8
z685ad89d01ec89294420964254420113ebbbe2f5755dabea66c84afbe6703efdc9b62314cab9a2
zda0a12beb45354575f7ab31c5a789b849e1826d1696e148f19dd328df64ce2717b0d579eb46415
z14db8874bbeca8517e97c79d701d3682506dec568f82d34993c1f908f53d53fbb5531f01cffbe7
zd7e3cff8d34dc5802becc578eb8098bc656d31948f5f0cfde9ecb7ca761b2ef5496a572e4efd68
zbd1628ceeba45b8b2b34d411329f76d5e34277344845cdff6df73df5142d6ad950952896d87200
zcbe79fa8dd7e57f4dde0db40350cda5b77993cf7e7a095f0954a880753381bcfe57b4aa791e768
z61ed664a60345b322cce8e1fcc56b2d6cc81fc3cd1e4ed4b71dc3a7aa5887a0961253a7cdfa8a5
z975d7ea1dbdc1f0569fd5541c73f8250620636e26cc61491bdcc9a652b5c664dbdb2edca12c75f
z4424c32c6faf97c080ac806147fe2ab74e9884166f4e2961265661ee0ce0f725a970f8ec9729cf
z9a88d73cff8955ac8140563dae784991d38b3b8a081328aed984c0ef32dda25c9b3c4c2a280925
ze0e7b208ec24877b7c7f15e17ad15ab2bccab2c6b3ac311b015548c6b0692ee95693a40c9d238e
zda386c35eea67bd4a024591e09b1efd28c0edc8c132fe3f115e9ef66f95cfb9ebab51e505222b7
za97285c8e255d590cf869964549cda114ceecdc78b80bb747868de7723f934f61ced38b0979d68
za9bc2c9d1e618f234163711391d43099bd2246e801968834109d1368baae5e6899eb5ac248b150
z55caf6bb69b798c6fd8aff9872ba85d9f34cbf0af6f35aa540dd8ffaade24eef4c22a1412ae407
zab5b5ec21252ea4d293bb55a3984a63b514fd554f17eb2a6d49f049988dbe2a017b355e56c0ef1
zd581e9a216fe552d432fd9d0bb0509f8b256a1daf81ffacd308c16307dfbda176371e6fc233748
zeccb16764f50569de3cff4709622a731b49cb7f25fda8f222bdc01775ce3a4b439c71fd494bc86
z88947d4783cd5e34ce14e051ac145d5aa86d93d501ecb943b3414fb427285899393033952b0eff
z43ee016dbc733cfe048463223f2e54d4c640b2e0da2f42bda7d614a54c46e454bd8ab7f70c6401
zefd7fe0e2580f407294855674bf9b995c06715c6e1abcfbb7a87b3f55be670a1f4696e4377a7bc
z6d1d0c6219a2184d1e016fd4c86fa0f067a32995bbbbc47d0706a1856528bd85106f45ca84766c
zf7383a2cd7ec5e76b633320db2487d3b3ab84d99938c4d9bb541299f1599f4fa75b535f2aee001
z327c09d19afe4c97901e1c9080a01890c3fe77dbe51db1d083327eec9311e0ca53f0667c182b3b
z3b01db508ee51ea02434ee8f75013689596aac93247ead89ba00bf7deab1ee7890c519954e015f
z8b6c361692c9340a98d1a417e6b20db349960decf6f9da6dcbc35cdf332f7c40929831ae0945c3
z2c8d6e3afdb5316331078abfd516f97f1348030d51d3bcea5c03c9d70f625381d1d69abfe60c84
zef50ad5c37c358f17f2a71d773a449e123b9b1a9e3d8cd90725b1a827f24ff55b54d5ef50dfe9e
ze23d32b0ce170e29ccca85f10f54755d26c96d22061b3e075fab9d287fa663f2e9b9c85e5bbfd7
z2f332510fc12d5618dcfd45707675db8dea5995e447078fa0021fdb270bed8ce59edd6d96c8f9f
z6fe3b44caaf4bbffe104e80f18f2200b59624c584ef4982ab03bf473b94dff0f3a94b511b28b0f
z92d2584d0003fa13c436578ab3c4ff3aaa8542cbaac5185f0542d8254bd43eff714b2bea430a42
z379bd97ff6031e417e4ea12d853fa03c333b0b39f2e4647d984528be5461bdf1b1b4a59a7b0845
z8e2b61682fc9ba128d454963aee440d7010d1b8bf21d9a7869fb8718286fe1fba30641a5641ac9
z56b743e504c2ab5b422fa8769bd022b9f262d9ee7b095753bbefaa51e9c078444193f1640788c1
ze4f81e4fb565b5e0ae72a45a2f196ce0a3be6b5dacf198282ca6b1ea3e7e0dd05288844bcdf8a4
z4e8099e677b8b0bedcbc90e30deb940fa7cb3d82406602d29f532a06eff4879173ee0c299ffb27
zcf470a42c3afdb48c0f67ae2700b9d41d061518238051b12382627ca68d28d04674827102b3939
ze6b84865046033363d81ba5607fc9333c2a7ee3dffe8b2b68129b6c1c714be0c63377d81f925ca
zd1f6fd1155a35bcf7cc4b67c7b41971455f0d042f38efe372a6671eca3ddb69a92b953619d50e1
z3241e76a6460fe7e54d0a7b5f30f74bbb80923f4796a3b27072900178d04b4831ef71dccf7f69a
z430cf1a023ed2f5158cb8ecec9d99fa6beca6eb1438f9e9957d56c10235ff016749acf47b4106a
zb75fff9155e185427c13d06baa6293c8f1c4d109018339b0e2b06b91d84eb04e16ec491c38f47e
ze4c4e9bafeb701d4b2cb2485cc882d37c9374f92b2c9db93abdbef4cfe7a1fc8111f9d709fe285
z8c338b3654732bde02f0b19a22df412914c658b06da3681ae58e3c69683142debf37e6a4b08e4c
z3b31a786053edf069f95f1bda77086dfd9e677c01a7a00f879d7255c2b77c19e4129f67da3f01a
z0871f57ce2394032d85d0606944b341514a9e049e02fbc133576a070cf0821d3d818655eefd29b
z96d5993790a9061b66be253b19d87ece1c4461c9438521795eda55c8cd0c0c5631443e9a0e1b4e
ze7391420e2effd45641f72aa3abb752456d21b42ef07b44cb7e62c95faec4ca9234aa85973d915
zf163f228e019ea0b745045951b330a39ac4869b99e1e88a257d96bb8888d51aa0a41fc03c6bf64
z954ae6eed8b72943e1bee7afb8f22275feec95f30ab5f12261db364b522f24e67bc38b80999a9e
z35ba2f2dfe4b1c4306507541479c9c4b57541e0111c758c952cbf9e121c62b6b2e9003b401b36b
z0d918de5ca17485f4534d38683d251365124b91731ec3cc2fbaac088a702ba9447a979e09b898c
z5ed3a46c37edbb2db5a7400395282f6846a49b5e3d05a0f075cf1d1885db810308ff8a1f5682a3
zcf7f800acef5563267ac656efd1ad7ccad623ed8220c4fa1426cef9d1c26a27e4e8fcaee867f80
z7277bb7fc3b860f6124ca9ea229633c36c374d1fb2112ea8517c1f5ff5946279ea06ad61437f72
zde969b8874c326e163116e0ba25280d46af98152c442cee6d61b34d29bdb463ae499fdf7bb61e9
ze6f0b68897e5968a9f6cc8b041329a73f27766004647ff21cb50a7eeb46aba7e0bf725a79d4e17
z822d35604a965e0eabdbbf1c686210ec3ddd56543d7e903cec097ad9d54961c773f43d54a27423
z86700837cfee167f59e696584c354194e2eef961fad6971f9da1d0eb5c5f11e359be75f573fd08
zf606b16ba156f648defad7f6dc47b024754468b2a190271b16221b43275ffd10b9eebac7b16dcc
z1dcb6bd094b317ffc118c8cbd3ddbb966af95c4a2be7ff0bd3a47a5546d4231ef6ec79b2d2aca8
z093a1f4df057cb6076a36fe3a5457567b4ab77cd1b2ab8779b8c57aed8812968110f05d7e9af2f
z1f08eb4ccbac42cdc7b6e68b2d09f820c98cedc04edf78ef30eb40f15fc1f3403c23aaaa8cd577
z4e2a64853a932c75f91989da6ff1888e22d99818b28c0695ae64e8fb816768bd5b390e75024301
zda117e5e4335d8061b3b2016ae5fa19ad436fbd38d978b4515b6bd8b84409e0ebd015a8ca7feb9
z65fc700d9c5d7e89a9eb8de02f215a3afe1e53d68d5bdf873cea9bc175396508e0893fb1321612
z02d33e9dda3fdc77b029fa5c93a235aeb1919c461d4a13faa1f9ec35984af4b95fc7afabadcb0f
z93efa3d13aaa8dca9c3fcf87501748cfc31fd70229814542e62868071944b0d410f8ee42a520be
zc78e425dc4fc8eddf6249b7914d922d4af90d3df65610d03ae62a29565e125169f61e510ad1189
zb7c50355ff6e36155dd796a60dc3ad8fdc30abdf20a3ec7bc664a6126f1de5e43d15d62be448d6
z1358dc4e7b11a355c43aca725f401d05c2aeabae9bea10bd44744467cc53f6a969860abcaf3b7e
z2b4d97efa9c51000c7fd8c2354985bf341e665b22b8f95a92b9d7eab55124bbf25e35916843ce9
zecbc9e43bf6c7c6ac838b1710c61a20f3141f129b9982c0d30323f480728ea8fc559a9bcb0fa33
z4f7173e52eb1589f1118f2ac06349e36a2ce1535c5b752e4fc85bb5aa760346c079d7b608582bd
z23985e98c692fcc456341535b4e202ce1b3134637bcac75ae8f33521b2ff03793c764dd7db4852
z3d1de56a36a63e21561430b2cc37c16fd34d8b6c27aa4e5f034e9ff7acc3b7a23b40e7aca01853
ze6b7cc63e049e3cdc4da74bfb04cf164e8e8556cddf074994718906b6fef0832f1fec81b14dc4b
z28372ca5569dbde5a7b6c0fd7607a6f6fdb5da543eba88b9bc6ae19dc57c530365d54abef66736
z0355ccae939be169b36f7db1a9f702a3efd8925253e9694d3d4a6be6843ccee51300abdaafac4f
z22c7106716b72ce51a9d12db1da489946d24f460087bfb1f2895c65290f550f8724555c320602c
z6607b9aed65df93130b2a9c8eb49ccbfd3c3e00a95ae8a0b3ddf95eb05f31a25d38c9c68d4277d
zb7766ce767bc63973ef5a3ddfcc406faef72c7c9455ce50c4c3e0c139140e8f49184d6c9102263
zaab9f7e891d9de690e5e3ad6890424a18b264dbd792efef4727b5fb1efdb21832ffb89145f41d8
z8b1960668a66fc9cf82f6ca26ae012d18c784304c9e3448dec10ebc4aa7b75bc2d984ba826c28d
zaed2ba571108480ff71dfb2d148c86a1a9d72ea4ae74599abf9a5828931f6bd2a18d6a01337710
z7905c8f4c6fcc71a0a46cbe16a546f84e28a3f922f35c93896b67d26cc58274de0e4108c546dd9
zcadd98dfae9790c788ca455734dd6dc9500d9bd91d0409febba7889da715db1957e5a8b664a1dd
z80df6c3f471bb341e550cf19c5026009ba4ff0da822f73e90dec288acf07f9a9b83001e74341aa
zf13ce2084aab41938d0e08d439b4e998dff0943b37c1b477ffcf066a3a7819f3c8c3a08358810b
za5aced50cfb1085683481fb46de5395a7ea61b68eec575a072ac336e944d2b96f3b2c041684fbb
zda3571270bf2b0201fcdab7868ea521a1cd9c6b1d2a08e7394bb7de75fc93d7773072c49550058
z64ffe084100932876a798ab36cd7bd5fa2826b3c6dd7f3bac25f9ce06cfec238516c698f18f481
zbeb0363b25cf05d350940b56b23f324490d93061bc0c6822a7e216e96d280bcf84e9636fcb0f18
z9f8e63f498015cdad3494a89a687b944305464e47f91eeef2bae3289b0b86c86ad0523d0c28978
z7eaa674a04f0e41ee6357209040ac7ce67fc4dec1a764fe22b2b0aa06408a05289a6eb298a68a4
z5030cce791c118872b1098f7a4249e1f03fe564747dac665b5d48e9c1435bf37ceee90d4a0b1c7
zd35bf801859e53fa47a816c928b64c14d6102eee2b2d4267a11eac018d630e2c1b2b2d681db25e
zd74502252d7197a68dbe0a3235d3bb45ba6b06ec70a87b2930eeff07dc8d474465599a72b73634
ze7faba59f34c97c5e821f62b73540d449cf2889ae845825f3d1596d130fa7f4df83ba24e2e20bf
z67d079938c0aa9099a3eae3a196d7a65285dd9b9441b8f91493148729f7ffdd8e594a87bd8389c
z4439318caaa2608372c38fb60b4ac56552f969af4c1b5fefd7b3f7a030c163790e9cf01be60981
z1e6b139e412646ddd369bd35b99c7f82a535e9650208d814521912a1b15a29ac37354fbdf7bc23
zede31a9a5716c26e8c22dd80e977c0e8f606dd36e4254a4da08b3882db14caad330bd62324f768
zc52a16c5b87325c9f247815cd0f40049ac1cca58d54aaf24de56b7de6c5311874f0043c2ceec9d
z65f15c278e2b001d350ee44787e64a26aec38b17981cb79097c72ff78e36a4c8a0d099d7615c35
z32d02d737a0d24a85e7a24b75941c501241cca212ae2c1ffff61e249145d42c503ab982b6db5c0
zb1ae6c8502e45c48d446fe7bb02a9dd891425f2201d4466731ebfe9e083ab76fb90689e5d67894
z58753de6987c0ac113b70ff22d226dbe840f8b3802cd8eb9020ee958105961281e89207ddd1186
zf724190d94a8215bc88dc9fe4b25c84f14c06a7c5bc44e50be172a9c29b76caef3bc2b6d2e469b
z6568d10361cf42aa691435ff5bdc1afc67888bc17c177c02eea27c82192574f05acb3ea1585494
zcd47f756fb7618c0eaf8a83c10781b663b7a11dbc0b2017a748845051672edf3424dd9b243b9e8
z461761fc91133f0c166ad8727ac20c8ae882f1e2028ac35176fb30244b4dffadfcca63e7a70f5c
z2c92e739ee866bf683486df0700bd72f67a41514549940249c570cba67f70376e84ab55ed7934f
z587e4938e8c1bef59d2040f18f74b0307b4ae86bee6b05ea1cc0e420d2087ce49b68d44bea1e48
z07d53bac48c644d6fe9adcee569a3c26f3d2bee1f770cffe7ccdb189b78aae44fe731acf6070c9
z25688719211e733ea69e53f115eab671a8ec495d9c8d2d2662b8948bd8a8d295d0bfe75c6fd468
z7aaf76af90aab761dcef2c97aa1483013db635d712ef7b1b9b1c547baa88c110dae2c63106e2d4
z63ddb505512c0493a8ab93fff8edb2e822df4a5a592e6fc086c51c33d8d2291aa00fef71b7f6de
z7462f3e5dc90f30b75b0e9488447c3960584127f1a76e794a34f7939adcc95fcc51e644e9c2109
z4980f6a311b1bac1511bc8cf1c1b7b6f8eb26841789cd5865db1d80bb8fdd4a3aa8339d2467508
z5efa7c1126362d5310c44914d2764b066613516eba0fc157f508aef91235daeacbe515e7c45f09
zc76e68221662b703d6bdb71956472d077466a6979299999c8d33e426fd625ea3612405bbb3cbde
zd202d428cfd3b79da18b4f68c8a33afc4bbd57c7c1a23172b8aa253013554d489e9f746e8d4c22
z18f1623bc5a651a35676db7c5f795722a1db558261b9e01679cd95e5d0a229764fd685865ad532
z03772c2e586a8270305004f60851a0ec28ac3e43dd7f4077a748c3cb377bdab355a42a78b28a78
z9a07d45e96a517fb7323c9236dc779ff7c91c6624ab1ee75e5820016310d62fa2a948941a405b2
z8a8a6dc02905794eb9ba7ac428653aacc743e2582feb8bcd0da18b7a5dfe8c6e085217a004ed2c
zfabd65b603d246963404f89cb398ca167640896d04dcb286c7699abb58df97caa0f2b3386dc3d7
zc21e921fac4e698919ea265ce040dc66f4476e1d2187d7add829ed998a793f80aba18ef0737d4e
z2d53c93200e74070286154e452354f7487b278dd2308fe85698fbd396504ac0bf911285a763f18
z2936b8df9729e2fbe443fc49851539cb1587981d48ee8e46bc14b532edd7e5f2eb2067967768ce
zd99b924189cb936e5f1cc6cf0e8178687bedf2950ff039329cb7d81e507f62348ad30f1d372fa0
z3e4e7330e4da750a60a89d62dd711f641ccb6694c0a21a88c2c54816995422b176a15364aec02f
z4f5ce6427b8f9e223d4cb73670f3111c5e1b493499652ba63ef442e27306ccff89045ee8fb38c2
z1b42e43a44228fd0f596d430fe2318e882bf0e7d9eeb7e76cef9bc2b686668a3007595ac81b19a
zab3a1949c428607749f3846786885f71eb72a729f36d293b12c7aa4647803f8ea69d338a200f84
z16d72727c4738929a4a062a35ff9d0336a3776f2db4be9b7bdd846d10132c997d3a18218ec5cb0
z80187e74089d7fbca2d582c1b21a061d994fb3b5009cf3db06f392e2e1144a8c00890958d1fe2f
zd7cde098430e76e73ff5a80fe428853834a07c2543b4026706bbb8c0cb6031b63d1ffe900a0767
z5372bb9be4b9c9765a0b98f31d69fe7f5f0736c07c7796de9f73f6d35b41bca4a856c1e9bf4d8a
z163b499c2845e720683ec082b5afe6566cca6cdddbbf73a62747d7ac477dacbea872cbb54c0782
z9eb0dea8eca28f4ef56bd339c47ef1b383453e498a697723d89a7186ac52b8e36cf3cc318379db
z1f591002939f5efb164aa09fd1a6bb365bfd4443d575814abd11bbf50080a5c1782ea8507d0582
z0a7a08d295365313f83568f34d3ffb55da343a26b9a002c710a140ca1516510ec9845b7fad342d
z8e9ef1ade068609851ead2c0261c48abf398e9aeb7769f4be5dba30e9224eb8c65cb564ff46342
zbe89f95e152304bea781a4e34c32d75f4b6a42fac42f3a473b4449049174002ef6bac30cfe0c3f
z367cb264f8ce211fcaf8fd2fbcd527bdd7919066bd211c410142c2747b361ae085609fc3ce55e6
z1dc6ff3db128c69956bde12219329c9da0d463318dd339ecac23e3f8b99e3596708110a193943b
zbba564fd3ea321ad5177deb4b8b356509d8a1d46a9b8ecf0cc58f64f2614740a764f7d8dd84f9e
z15b5518ca3b5951af2ab2a32721881b422a5310617144f966da651ea1b0dc968cdc5643ec38979
z488419b1cdfa648d29731917c23fb84e7cf5d661a59cb9678539cb269863ad8219a9c3fc8b3c9f
zb2b5d0e28c907e0a1456a55001b2c9d0aca7381ad685e7ca87e4338519bbb4146911a0c66a26a7
z3288995cc0595ea6f299ba68942d26d8b120eefdf457149b38d6a3f009de27ab835cd755b8ae6c
zb84e1a961184ac007ba6975b3ee40180b1e2dbf097a707279d8f4db4267c0db9e940a6c324db89
z44146f6eb704ff75baedf3ad81e9169462080fca777d05ea26f365124621f75549aee585f0c5d0
z91f074910cd170715174651b723da7cda7d007e84cda82c7c97dc81a9be7c3ad5bbf2e856bec53
z5e4a0b130ec7177b460eb55cd3f0b197538f9ed685902e39fd22df96505c3313b3ba14813c6851
zc2f9970d66c6682d51f93ee2188c36799892619e78710b27b2003c26a586c4016bd0f6f8877304
zb9de363e751562e7aebb43e597322166f37c3439541dca7e369d10ac666554a2e04c257d80c636
z7f7931b47aa281e0e4b9323d121b968715e55f3f3f7128ed20f6edeb86fc02daa5231e515cc931
z6e796fb94a369dd6b87d5b9a0c4dd5bd31d1d867f0824f7c34dad9cff1a5ce21d715e242d00f4f
z5b903126203d1af0a4de17185919e6339a8e1cef7e90241e733b991d141dd681b4a11ed7ff39e5
z6f6786b3aad366c3f4ab5226bfb003f6b699b9336122393acf54473b6c91f86c483b526bdadb4d
z8a04cc9d158e912813442802dadd88b770e6bb59e81ce16ccc02b4f93ce1a00aebdb8fda532bcf
z03f674b98c5d3acc3f0b600908a098f18c4318b43b6a169f5639862a5b4e832663d504191b9411
z7e2da1993ec84891dbbcbf29e49c578a918bc6add7bb442bc543880152214b6896377cc12cf6a9
zedf0f8fa1bae1fbad3b53a34251e7d2f13ae52e0155afeadb2113b5b2100b23db207fde654d7fd
z97208a9309010329bb1b6218917f774453a1c87d83680462a4a222546310405cc76efd1a340335
z6a0eb1c7bde382d4dac7721a7c2cc69bb8ce87bed0acca70e7bbef57e14c4cbe2261427f365071
z966714f533b2910ce79d0228342f681b53b1f71be017efeb8cb06c9dcba7373f71462841c2b53b
zdce6c494cc8132718f35ab2b3276e6497987c8f9f25fdcc3f198dcba97152ed924067f958b1c2d
zebfa6764b1cb10ca5ed4b3ae306c6cf661ff729d136ad854a9f2556ffbf47085ee114fc39b589c
z303da2bc5125aac356d24cca173925745924cb7ba67d42b39e978b762125b6ec9ab6cebe6f0cf3
z8a0ab304b5610e427fcaa4f74e9b07cb1c75de8a348672e005bf914b4a5fc060bcebee3b032efd
zb74be83f16a1d125b86629068541a499f94fb5ed30244cebfc59e8a3645874ea19a6c2857e405f
z8fdf02c26e9303dcf97fa742b9e3ac30aa162a9d80a753b7608c7f5264b9bec4ad6fc8a6bd46cd
z726aaac8076287d44b04c9a30c86e3d98a6fba6fdf689d148f31a3501a3cef6d786f1c981d9cf5
z15c70a529dd1ed5cd9161292a19f0c77d3f74b77589f3d4f68fafd2ba1746fcc2c7d1919d54dad
z83ce80c3bb1516f9677340b79dee6e1652daf24cdf710c425e38b47d494a2e2b71d04cd51fcf15
z6f70efad063d78ecdab77095dd928b1f9bd586a863545d92c01beb1dcbef1b1544964a1ede2b00
zc7fd11c6db2df238a4ea3d9113b7e12c4d8f124c921ec4fcd37a60dac2b87895cca0d8534f3d4e
z73278338f1ae689158b7b084ca25e204864e5b8b3d9ac2f359d36d28799919bedcf288f308622e
z56d26e67a1a8d06bdf802834ab4d6c939905e5b91f84811c497272e11bbcde474b4355201a0fe9
z8b3a792ae4f5aa30d7b2dbf8fc2bc27bf1e3b501445eb9419e9bfddc7e86186f70d32fa9adb3ec
z3d6e332da5b96b4673475cbbf5c4099db80ee1d5684eaa3240aca496f23b5f405f6eebd677172e
z5db354b0a2be8242cb4e6d78f53d0cf0772b5c948349f44def5da36e2d1ca37c832126c44a7cbe
zb356c988d62ea77b7d9051d0d73bd1995c2afe1d92a7c72fce389c70ddd3ff491a4204c0c57070
ze5bfcf766a64617d6177f4eb48a97be128df1a7534493f6a55458fd75558b7af515c8881e0279f
z466bdd8e4e612ed8a56fd0b392c21fcf6811d5e99fd17354860bf44b19355302395c1ee8072779
z36828f0aaccde913c35f2d14ceee9ab7952bbaa9a69e660c1a0ef8758c7492db5582f7324b11ca
z50641cb00a614b07d22a3922419f4e766adf928e61f62d1d61e57aa0c3375cc2181f04afdf4d2c
zc554ac114d68952af2b00fb3f4f33d873310320ff1373592c794acc2ee58363d6aa427bea60c21
zb0ca98dbe5a4dcaad85c15d4c23d6365d4e1fb9e3ce8ddd5fdd8c966f3291841c6ded21a820aee
zc8ae0ce69d09c388cee06dc8c02b21bdebc683b09f27c1b228357dc28dff7dc77587c70aedb803
z4b5eca9dffc72a3444ac75d9fe2e1b9940c9213718e0b717d71fdb5b1543003c193fa459240aaf
ze0fef0047fa44ab9c26ebc60a97ac888c6164bfc8a4f4072d6ae941ec7df0e577e210960b65c0e
z6ab863e506bbe543656efa4897aa0a396ae04e484fd001d0608ff356cd11843e92a327f56c71a3
zda9b810e42ea02c148d59e23620960e24ba77e7f16b269808c93b5a0fe7568843796e5ee12644a
z210d1527f731b7c3ff80a7caa611264622f9a580bbba039c7036c320856a86c9991fd00cadeb31
z4abcfd2f5c2398b9f9ba506815a33deebb94a567fdb3f7c20492e80af4cbbd5d862c7682d0af22
z5469a59c1928aaf0280a6a3947bae396fd27e88410de485684940fe6bb9719ab36d7c97c5cde4f
z93d3e662e4679e49993b57d3c2296ae562c02270a30cf383e690a05a778fd620f773b809d02548
z7098a30c436b2f3f264c1b88f24adfaa556c046d8a87c7e936404f96ed8573a4eac757986e2c4e
z3a89ad52d4bf3625f4f314955546ffb5f382270b1d0c176ade087f024f42f3ede60a7cc2268ebb
z92b9cfa81245f413204b4871e90bd738f6b5bda83bb08079d1ac97219d395444d22749436e413b
z4eaa8e4b86a1924d4b069f9be5943b77c7246092448699537e6b7949ae19441e3f1fe786f9ab4e
z86d30d1201b36de86b91a55fd4360e9ba958756a5d52c035f4bd34e2e182d89e6e8bafc4b77c69
zbd88485b403451b74924bcc5e731eceef9e2057c74c08da5e9e8d5fc024a6396817a341eb6a4cd
z4a5c2f99ff19ce6804a61931acc5d44ab57c5df5d7aaa5029c7936f433a4460f9b748d45ad5cc9
zf578a7b0a53a1b538905cab0405b5e08ddeafd2e5b74f242d593f93efb1b97db0f429cd3f48cb4
zc38d3e11ee259da2f457a40159194e66d82daf2a37ac59b9e2b818359bbe8ed82aecc964cf1b4d
zca5caf2b29143b0fc0
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gigabit_ethernet_gmii_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
