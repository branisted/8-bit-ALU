`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1b93f3c788f25d5318c12e50bdced91c303c4d
zaa95dd5240eacb0832aee7cc442fee02c4af069d6317ae36e1befdeda8feb65e1b4762b1aa3dd6
z76acaf9268a261e49b1552ff575c951a2d29c0fff477e3a5f0d27c921a25fe5f1ac5a422ce443e
z2cebbdf7d67d5697211cd7a00c094c1175290ea4f1103e129171ca1111bb6ca801da60f30baf38
zb63695e2266b28ea6d640bf6d312bf0e308065c880181889f24ab035d38a79de2da61c1fdbf5bb
z088475952407c829bc82a5e6b6714597629b62dcfc085381eec18302bfb57d74d2cf982d6c55c6
z8593b61c44083cb6bf940baa1ee288bca40f4422209a23cb04530a45fe7a180d990e0857d04e1b
z2f4af06d071755ce79cf4712dec9ebc126336abc65b167f80b86ffe8e10b27b505b1247c55f03f
z85449754bf0cc53979fcefba941a037b77c55b65457fafaef987b9a913efdcd9eba2c83b4e58e6
z45ba60299c1b1ba2fc0487a6b9b2589a09e03a1365ca8904ccff544a3f38d68f3e7178709a63ea
zd17d19811d579bebce938c9bd7854e5f639378010181bce3c8de28d38ed647302a5c09bf7e2fc5
zbb0d7b84202227b92330b9d0f9117844db5f37896f2b31261e5957969b7536174c858c17feec9f
z0ae6effc2acd973f812c6228c013f87393310b9395c6b85345c1f5c719b2b6bae9269daca6cff6
zf2935f17fac1c7b30b17df87a401d4ebe2c2f6187f57b3560f622d2c7b5273f7dd364bbf8eee29
zdda47293f5e66f18f565129c21eea7715a6a0b676f523ef191a6c7c6694ee1a82a812a22a9cbdf
z4cd80af898dae46e27c2cc36f2ac0c35c03b6a6c9f0672a7b94008768a1f89ec7e9e06ddf8c8bf
zdb75f6dd6e7be7ea16fdbc1561bfc4b27747c6e4f31e39abb17c1fb65f8c31d5f73c5c67b23c43
z7442d8f9767f057652b1f632b22db0d10f1a808f0a1a5c35fd3d96cd271be1e8e7f97b3fd9afa2
z22fcbbb234b9e3253fc9846cef98308260d7ea40181a66ae241d1a7889bbb84765171a830bfc81
z06a896bf98d7820082ebc91360adf31f80228c9d4b32458321977f8e08ac9d3491efdc2fae40a1
zef104423dbbc7c55346291e1b28542ff37c80c27922c0b083a06243db13b0603e7f82afd5d0f00
z11509e2ab259dd027466bc7bf59f1fe0f59abb0f43e4af57dddb8e407173c77c1b475c5775577c
z9997b5e0a6238b61fb372b054cf272a3d576bc0d79e0e29214ed722e1a257f619465be9b8b617b
zfd63ae5d54128893837c347cb58433c41519b4fcdd5f2fe314d675d3dd906e92969133c4204346
z6fb11a75dcfecc3dcae6a6e887f185c424118510e9a396d744ef4319620b92dd702509bfe883b6
z4c1bc7ce4baf04d7073bf47abe19259d8f21240480dee68f99405aeb559ca607a24ea456009465
z801d465ad631712b30eeed31ccb0732c48bd0c72eb73e65e21bc6d434e10024d86f3daa4cbec1c
z665da4d7d32b262c2c409aaa4411eccc57a9158199ac0d03e3c206aca829f9ffbf63670169e314
z8747b152afe3f8459768ddc72da2fcd2f0ba36404452ed230583c3170474f2c8c152de3fe4f2d4
z2e13a7f8a73787c31e3bed48c180cc603cf8061e06739bc42423781190b6d7dfeb46e08586c860
zc200947b122e99dabc4e83613d8c6cd810b9a868b41c8bc837f132b09620525b3a3e1530a2e76d
zd35d98d8240deae2fde0ce3ec4275f776f57cc38391d249cb64c8f8671297dd49cc9b39cc7545a
zc8fe23edb8ad8821fadbf8d1afbabf4bcb347acb3234e906b5a42739406a7ebe08b98fd44f35ee
z9afeb742fceb73e0604c17667e17b4b56fcf46d53a342c3242421980c13ac67e5b86599c2d9a14
z697f19f76bc498e63f103d7285ac157921ad489cfad086abcfff18ad420fb664a69639910dcb64
zf9b8e1b5c4bbc0ed811493b13fe60eb2637d13ae78c821b44703ee7ed577ca74703ed38db8645b
z9abf347b8e83603b99f8477544265658d573e80793022459527d5eead45ed500d8655b3a63956a
z00d51e60e375ec9b798ca10967a478af2fc64bd9b0d326d18aad851817103f393d4f0f1fe81931
z3e782f5b7be9c96cb16a706bc9ce59849d19e80eaa91e227b3301c0ab3c223447f4345cb1977fd
ze4ec7f63b2c013ff625a1bf073b09c79ad607accee03f47571a956b1fe29149e0812886ec7e9ab
z627e6f7e3e096d3d628cc2c78fb2cf741e9970fd6532f5fa348d7357dfab29e96dd1872694b781
zafd1f32ef6a04d26687a4ec1e9fcf55ae41a4b8d79a3c086acd7e2254c0b35014cddc9be8475b4
zbd7dc3ce38dbe39143f60dc07c055b7d709a4f35d50ecda1824cd5c0f9825b5d8c1a8d291a3245
z5237c4eedd2433b26266399919870048618df59294f7f1d9c07d3ef85d9e8bb82889e6e2f56b12
z6b242ff9d1776a5b505fd5224212163b695a0eb24c86910c1bf095d523f4d0e2624cab78c0971a
z7aaea4097097b0523cc3e5d6a0cd3536eb3849e0f7115c1939b76bdad7715722905e9f1af8ec1d
zed647a6697d00cf7b8dd75abd2d1ab9618c2f6ffd2b0ba451c3fa2b7b0a11d35f3abe7239af7d2
z425e70732cb6e2935affa7942259936c305168affb48eb09f22fcbaedaf03b25daffb969ada7c6
zc91852851343bce70e722f0765f7cd6c0f5bfc972929732861d8fcb0990f94f9e9b877597d0c13
z178b7817f1d2e4c35bf67f6e6155d13d2b9a517a29561c166905c4961ff958a40417e286431f99
z5c53504555dbb6b58f5c4520df16269348e7d6aab0ecc5c28800b71de358322b7832c0a98eaea9
z637053e411b63bc79adba72169b0e17ab822c91119df95eaf669303997ec188c7be63c7fcd3470
zff57c9d390c53b6f0e0cbba5b5b7c3fec37b303643e87583c3c273d028f6fd885ecf30b114603a
zb156db2fe2e7b025df16a163c5872e5fb391bf0fda936761c1d2c8c8759697a2de144cb1a2b744
z2900d202dd1569294b5ec616f5a2874d3e0d1b51607480fc3ec77e1b7148b32f73153f59e4866e
za60f5bdd4855eabba4f79243828211d9b0761158699d8564781b81fd859975d45d87f14aa790a2
zfbe50452604bdf3889aa068e107aa3113acd3234988f3d00ee231b0e184613cda23ab03d62452a
zc30f6c2947c06232da43e436082ba8fa3c270a9d7434a665849b18549fee5b87a49eba50e4a84a
zec58b69fb63a532e203f0fa5b5dcfa9c1f039339ac66f08b94da8cea4938d73ab1ec329e29c291
ze7810ed7c2c12e13a00b2cf11d044496f6b16a00e8d0813b4d45b0a197d1d01fe08153fab8c27e
z10fdedcdfdf02ad191a2701a9aa9c0c5cb3d6e5401fb65984454feffcbe32ac436fce3986583c3
zf0d47e72ab011b9da48eb734655182dad1056fbab5b710c0083f746644f81226cd3ad8f12b49c7
z164a12533326dc463137f6a54241b0543528a74d3340d6238d31d57b9d39d13f7f37551f6a720e
z9d70a8b292e171632af6c791eb126bed68b19f4558634564322f5d0dbcd0a89b3e13844407aad6
z2271f9ceeb6d146f91031c932c36a8e3eafa5b19f532ca52f3c57c039e7d0625778abc3c3f0444
z04c26482760497867c4e840075224a56ec79d99e10218305584fc5458025048946eab972648036
z43a74281ca5f4dbc87343e6c7e029c0d3870c46d3f9a52ee5aefde40817ddf8345cf1b4985b187
zfbab81ffdfdb144371cf1ae6853c2934f71155a4d12981c5251a9b2fd44cfff7823bcca3bf0369
zd372a2c1eba7cc81daf890bf7bcda7eacbfc40bf056e901b08d05b96fe4760db0739bbe832d0ee
zdb1fe9ab018d4d80ce002c4037ee1babff0dd1d330c3e2de027f97fd75c3824c1c36db88835998
z9f4cf7997ae01721e92e52932052b15765d92039e1870c548772590379b557d309ff5f34efc2f5
z0a0798697887522985d9693a337827b87166ab2b24e177626486202f08fdff1c0b0f5fe94244ea
zb92d749aaf8e40130f81e074dcd9bd604d871e05f6f89172c14d5281aa0bc3d74bd0d4ca9188a3
z4bf4515c1e0363bf94bfa4fb5ca504e36c86cffd0118a193dd2a4f7809c9f3e2c51d680aec25ec
zc413e3e800a0ca2789a1f9ad312d29b40ac90176ff575ef8aa473ebe7e152e5d3ae5be33d86f3d
za242794758e69729a5840570757dcda84a6cc5ce26653286a7b4f3cd73b6be79297320a791aeaf
z01dd87e8231eed52e6d296a65c762c995fa9a0de5d5f6eee2854b810305337556c7e0a3f5d2dc1
za5df6de9d949904d55583c5e6597eeaf1d632b6a86710cb010599bfc3d8816a1dae46e6a419e83
z85c9d31882c90adce3c32fd1d44f8b56f92a9f84026d590692803ffd861dd5b245bcb31e67c222
z1ab5ad31fc25d63760edf9896274cd265ecdf3584e8ce238b2c339e19fba7eff5ab0cbce0475a5
ze1f72d21e83d26749c4c68e3656316c4535c3422c83cc7adde6e3ea27fd4d4869caf55175b9443
zf2cd2ca0cc4418921e4622d5bde26aaa98eb2f203ca297f73f2a779fd261e700f9e2af6c3f7a6b
za775e7b5e49238494d3c4bc7f54a41da23a60e79af9729e9ae390e4444a333fe31f1b9b7f2ab73
z9520f3718feefedd01ebc4d76cad2d9db9d85a8bfde809cf3f2bf152bc848069021711da7f16c6
z0d71fb5d0c5461ffd48f09532870fbdcdcea28c145cabc90063b4de59bca76eb056c5be178490b
z05492e47f811b3d9d57fafb1a2f089769a762983049429bfd6be74235b9b726414bffdab10fb11
z4d12daa516713df237dc16e064d5c43348b76b3e39c7d7deca0680bcfde43c1ff6edc0d834b659
z7c22334b4d60aeaaa65fa4362d4762fcf66ae16b5c2fddbde2dcdc3c38fd0ddcede8139e6afc5f
zed849a07f1a3acdc0e63e1767351880163e50ee844d525e68a5198222bb1662cb1ca1810828d0b
z7dc40afa90ce77c951822d0d5fb3921a075ddf5d5fa219f70a1637094592c6c867e134e8fccab3
z07e75298f998f8845d867a160a613f836866ac35a2ade38ee924c1a032f3f9fa9a00f5a8fb63e2
z4735ad0a7048508f585f7759cc038985020f7d41c27a19928e94107e48ed4e14e2d90a3776106a
zf275b50500f1c74070e17074aa1ef768eb6652db6a30e9832b8e6b00f8dbbb5465fa365f3dc602
z8c925cfa321d71c55d4e705ae3623d7af3512169bf6126c8026d422f9b8159b7425b7902420e06
z3e696ad40848bdd7c54d331ad6648ee3957f8dc8b9be61e8d8de3bc6d468535192fc98b08ec93d
zb2509eb13a1711d565b5c9baf8ea73e90a92f1e86d13e84db9c6ebbbb56f706ba25ee87026ea09
zd28721ee3cc8f757229de1093583df2a14377783a3061c89952db45e1ed066d77b51069e36bef8
z9d7ac489298573b885e8331bec08fea6a209977dbcd2996ff385f05e74c2b697f1d6192dd92944
z319252c699845575aae0e48e400a1faf5ccd65c965add675bbd3ed97d9b3d3beab5772ef0373c7
zb0930ae61ee1651f4cb7052c02b9e8f825f70b10bbcfd15cf1e07df5f9a419b2e532f59525c769
z4e66d849c1b1b15de6060167bd755dd9fb35806d66877568e0c8ab2f386cc1713ef1ce4e67c153
z1996b20b5821c726e02b75e050b6b027a1f0f8e5b4498ade8da896c0d646223cafd6b1427a2b1b
z1f2d08d9669a86ee88f709809e04730a38d248c6e0832360722936bfc84cc8d4defa7a4ef03b3e
z7667470d543097e61cf9b96d46bf1dded682b684a8ba4b1ad078392734791ed8e71a72615e0f7b
z6cc509d18e03c43fffbd2696ffadd2e9f64cdfbd1618dba4290bbf014c4423c66d9e1c70a70fc8
zfd64818e49791514393f24e061698ab04f95ae39b52c3868d7d6d0ee074cf429ba76e486934a99
z6153bf7929ff0de8251482a593c45b8183780ce117bfd93b3cf5dba2f42c642d86a9fc3c7a0e98
z6132c403e41b058e2b4ca41875de82675dd5ca2eabce18414f4340de5fed876be90c47cbabb497
ze7a6f5eeead075d39ad722859cc19a28af40c1c5b664615c846f5f19dbabb435e3978e25c087ad
z3380ff0d5159fedb146363300ceb85bba6ddc585d88e510142e5fca0e80c822052dac614560301
zac9b59d842fc475ec22ce87e81e464358635411d686c39a25c61463ded7105c966d2b85f9d4421
z0df417f004849bbe57491f5e658b711805388d227afa6b76b07e18cacf00bd69e31ad5a2304f94
zb32fd0d3395186d59664581f91b4a4355d15d32dad500490543f7ff8ac7d4ede69f807237fcb6f
z822f51c5b64ed01839afefd5d29d9cb891d0821ab1c8055e366a9162e9c027c41100f2b3db8473
zd985ebab706ddff6ea68c4601a020add058849273dc542ab188fecbcf0fe1d059ac0aafcce2954
z356e46b0489b873a768c7ff7c49161d88a9dec47d225316043e4ebd94f25d41d4ce3d8cd403141
z7fff1a24feeae63eeaa83b1938951feae9c15dcabe2b034153544abe3963b8a8470c03d3f431aa
zbd1c57eacde45850223ab59741490b1bf5de08800e7213eb042bd3de9dbc78b7f6d6bb6a287d79
zdfa087a391f8afcec53dab5745d9b12ebba7c8e9f57aa4988f700b7176ca8096e2c4faabf9b1a6
zc55ca0f0741e9228e810b72bb3f716714deade9e47c4af7ddd1a9bb74a9f121ac58f5eb5a8a657
z2c2bd7bf17894aab076d31e6bb67126f80e5bab6d2adf709015648fb4e634938522ba3726f18d1
z303fadbf36525c45f8a0126cf37190d5135be2b4e4dcf46cbd32512bd9a864ce9471e102d0af6f
zf3a7f849c28072cec8a5577377084df3d6585933c6ba973b7ae221d1bc4f83fb3542bd1ff33221
ze5e1f353fcee9fa14491c2be846a9695b37e22e413b61c918ca6835e66e87b7fcc7688ce8329d5
zbae194e4b804d8922eae25e6cf7737b412439cae467f791eee656d631e732b893c74539f70b82c
z234f1eadd44c1ac69be9a2f1d3343132e6d4106797f3f6c78d0e607990b9e746967cffd6047b27
zfc9a2aced04b1d062054aa4a937fbf4557353b1527d309a60cbad15c116d3952d4e6c10feb3352
zd610eb77fa4876f1243fe0bd7721c18c1e3d2c8c458042dd6ca8c33de7ecd69c7d5c0a8e94ebb3
zd7b5b3a1d2644992cc713931444be6a4eb6c6ee4fa0280b49e8f693fe623c44bf3dbd33a13f24b
z6097fbecf8e729128e1ca694d09091e3580234b73c56b2f5a5f55ab3a86c0339ed7861f8fac243
zcb50da95e5e8d09b1d12bcca873b5054f050edc815939a469e25cb53ea5e308b933a0eef36be03
z5673428edc728101cb728f8846bb80f877abef3c4c8b474c0fb0c0b75819c9810a62365431e477
ze0b876be80bc873ac404c8a35c96568f061792f14bec6a9bb18f56393c44a0537772366b95b50e
z3a5f889970e553bc93093d61b2baa3e2018d57c5fb55fbf19fcaa949d2595060d4356802b3553e
z06085f20cfed7f65983c0178350bdb4cb3c171ce04ec5b20a199bc7c2250398f7f59abab71b176
zfb77973e91862415cef6b3daa43a5ff24c8e9bdaf26a0f57ef2f6164e40884eae2c8b61dbd38f7
z13a459fbf207ff8aa358cfd3427ce0f5ae0701c47b6f789361617485ef02a944eff164e209aaa4
z5cc583b796c83ca14d53b55527f785062a09fc9650b26cc495bfef7c7e6187c28f145cb5851645
z89b7677523f8d06ef885de1409084fa11da3041e6b5bff6a98188ff2ba43a94c0361b13560698d
zac4789e3d7704bf0b93ac67932c125e894d42a117cf2323cf640e89e3b7335b10eca2270cae3d5
za69a322b16b7e8fb919831510a425781446d2ffca16a9d0cb2a1a32c5af623e8f0efaf857c68a1
zaf8c56325442de0af1da3dd171604e04680c6db2abc2cc5459e7ecb648ca344bc4a379dcc91e24
z2685da58ea37365874de424e2aeba888ba75d8008f78bb572c3462e1d0790212e27c9a67ef15b5
za4eba84cc9f9122c0bfaaf8ac601a71484c2af8f9589c4fbf533774e644b0d4f7a7b802d7a2285
zaa8d67cba0db86f6c6ed92367deab024ea4db53869d9a9ea43c466b46d421a4f46cf58f3f1c7f4
zb8770bcc9b7b0166c310274ffae1b672625c6ceb4d47b912e8a78c45c06de5f25e5c5689b60753
z1fb7a5e7916257e0cacb4d3cb2ec039716805c6923138c10fa11c3da532f82a2bf1c2baf27ce9f
z92b6b2cb1b03b228e3d03a37a6ed44b642874713a7d57a16e527c2ab0ac84b2ec1526f3c196fc3
z9f29414e897eb237005b82347b5e81b02b521c0f1eda5e43a83701ac3c74b897622a4893037a02
z43852f85c21a4004340df70ee182ec3d4721aa714467b62888b5ed70ac8b53793bababfce39a7d
z5b3748af32a46e7fe53271130a158f6be428a93120933a081257a9f07e8b8b8eab81c79e598bdf
z913bc4db18ae3060bc047cc2c97f6b8a7c7558524ea4c9972c5a02060e9b937fa3e81107a65e32
zbf93bc6a9b2d26f58f736870560750ffa3baef116f7ac83b5910ed4785b5212c8ff8b2153ff7d8
z6aab574f7e51eb9a653595604c6cc78caad424f684b3c7418fc88a381c217a7e5bbd3a8321ec2e
z94deee526898bd021089ec766d1f2ff2e5a48362bf7f04bb4906ebee988c583757a3acdcbb8d5e
zbca6b8b95016d8d98abf810d63495fddc71edcef7882acaddbeb050a79092bde0318c309606365
zb0beebac746ecb38d95a16034737139c0a709375a60b04ed49738c719ee6e95bcb504f4df027b3
z71d4f85848b5655eddf08958024bcc4c9fd1bda345c3acf83af9a7d819d4ca22d8cb11b04a9869
z023ded38eba2ad89ffa94e58b69dc8faf0cc241fff9b322b492472ddc807a36ffa5143b094d5a7
z853786b2867345bddd039cc00a1cf9de7d454940823d417a8c94e42ecdf88a0c6137306acf2c11
za635e637d258066b620d1bf4df58a1bf341f171fc24b8ddaca6f06a67b346ed45bd963d282423b
zd92778cde0420782e126b1aeba5858a68953bd74a22d2b226a133144f7519bc0d15d0d12dabf97
zf5d976c57e663d9f05ac1f454bcc8b98b850092176ec25bd993fa66f9441cade3f26d422f04503
z07737816a388ef81b750ce7b5d8ee1cb2696723ee59ca7465545fe215dac8f647bddc4d7c73b65
z9b3251631789c3fc5929ddb1ab800810f4d46305c492ecf286c5b15303cb6a5aef3d24c8e3e68d
zde47b04b30819661a084d63d2c9e8e0a570c1c3d7d2fcb9570ab9d2a155e995369515d64f806d6
z0854cfbcb51a80a86d0fa03a1242d63d797300264bad8c3c0b6ecb6122e63eb0fc30b70255e771
z615461a6a0f1812cd0fb785cddedeeab1bafe86e59d755313de4de228e6e09ae9e45879df1f06c
z143b8dd95d21fbb5dc9becfb8b1a76fe8632135c6ebe1c40f80d8cc49a1a385f033320c73f33db
z50a41269ceb6dad53135057376e22de160ee98cea909c609a9bb2efcb1609759879e1b3e7f99df
z83406bc2e291f573372ef0692b50783e43c9879acee3b3239b7e9bfcaa1715fa2db45af7432d4e
zeff17296dbcc07fe3569a3d7e2815e36ba94705347e33cee5dbf58f442ad49731bc5d72aa78020
zc277c97e0f2472384bcacb0af0e45ce39b98007f35d5f7a42c28090052c6c4fd4c68308d5c43e9
z7f3c707074f4cc8ac85d195369ed09091d0b1cfac3e5e5fc9dbed2d98643161a28991fb76f0c09
zbb9eb7ec85ca56cd2a5aec97b19fae51278989ab171f36d544061bc1af05d326f41728e717be3a
z6ae5232ba4f394135774b87a268d4ecbe7ac245c24e112a4b2156477b393cb9e4305469a425a85
zd63342123c80d00534251d37145a9d5eb6066dc0807be9eff38f5177e4c123131d6ae7a9d4b873
zb765ae8df1cda10b42bc1fe56969e60f4db46f8bb935da8695d213b6ba7ad6a58343c2ffd92c61
zd4bfcc3088c4e34f282a5bd3322bf20a35b1f81b9ce710a83031d7bf84ffd058a79aa3f957bd22
zf07bc5cfe9e82831eb1df451c062302778fb618ebc8c04d2af9219969779a15f8068cc220ccd20
z83f50e28a0c0b08374491ba921d47f8692009c4cb78935564c0b4d3247806d4939e4e19be236bf
zb657b3d310ea6a5324c4d52d524bdeb9123a2e6248eead928447ea837eb010a5a1d4896da61fee
z55184e32394b801c2352c07084d124532e2655164582adf4d013e77cb12de77efcc46700e35c98
z7da73faa2fb485bcdcded876d8ddaae9c6e48da944cc14aaec141ca95e2a27933100ea7bcaa98d
z6d42aeaf998c96fe643fdcffebe4f5a7ae799a06ffdbac156c8886b400a3f648ed4458c4d914b1
zc77f868ae812e79f42ee959d123d66b57dbd106947e82562742ba0b2cdab227170f645b7fdf841
z0df00093bf051eb716eb4aa96f515832f14831132ccd9d3cfd632b5ecb8af850940f0a15f9fa5d
z9c5033493f9f31405d003107a1ff384c304a248a2e3fe203e263c6365b1b65350456cd3cf8f2dd
z182a45e483406027971e35e38ee5d0ebb8b5d43e005169cb0f5d37b05941c84c297384c90f47b2
zc95e8eaca055985949c1b2d1df25bf6b96c3a83a0f3c38c784fb92b730c3113d84abd52a8d15f6
z07e911fcb34e1882699918fd0e1a46eb9622c22e309e92df9b0fd6fb228d35f4df9a3d2c2f4322
z2672b386d56823eb1a7fc81ba80a8c8e653a49e413346378d889c48f6f5af06deadc58267e318a
zb007d292b70e5f85015aa7b315aa4b42d998e0ffda033f57b1d5c19a1705844773cc6dbabc60d7
z6c534ace0de0c0dee62b1e0ce3b33d47cc7a28e6661b2a3021867ac1f626d941d48b1a02129a41
z7fac1f533336faa95f91282ad923ca1b634df4fc0d2d25eb6a7ec4f752f7eea799375227350584
zf8d05db764a43567771199e465d9522fc07df46c90bab1a8f5c3385c99eb2a5dfc6a7ad635895b
zef6039abf136f8ec17938f5705fa702729feaec37810fca3fa7b2ccc2a7bc3e69bcae4862b07c6
zb5d455296870f2ef67fee4571803ae8cbfce2fb9f7b472da7616be56abbc99d4f66450813a7fe3
z7f4a928219c3c289de30656acf29bcbba2e17c5e90166d750b9f152144758f3be98bfd50133438
z0106a575710127e52dc44325d8135da0d4b180fc60361be335c220db91b4d43f194f86b8394513
z5b95cea1bf0c876bc005502fe9f4e3067542dac87220067572ed8cf21c6a71de1e1bd96cb7c126
z7f282ec451adfebcf6195ed004fcff112a8c53af196bcf3673121b2287e8e5fbd60fd791e95b0c
z836ab3811f2060420cfb6b0d78e4fbad5ca78152d27bfe7ea7b2ec9016a99a8244c6f0ec699cc0
z891f62c888aa7f77e3d01e3b957e2efe7f8d415fb7070267859236a33f9f8cb6a45af06cec0501
z823f764f4fb4f54c4bb58c789b415e2098ad7b5981bb7000d9e54b307a1f99e04663fe8459edd2
zbd28331a975a9acb3d753b328d42825ed1f6f42557beee6653cc3cfebb728170d188d9060c5b29
zddc2710ae6b7ef1e30b5617d5a8778d535eedb242d0531adc5c5fce4f9458eabd1ac83fdd0769a
za30acbc01e26c9107970d9e8dfd78b90234ad0bcc86bc99c73f0e341ca6159cb8d62272a0d8ec4
zf1ebf9aeb1662569a658fafbf3064504c8b9d5156191bc186a36538f2f014b82b3dce74cdb0df4
zbc568f85f5b82b61d99d1c061d827a14ea21cbc23272371f37eb26e309b2f24043c69a6613c4d1
z94061e81a30535b36b3e9ea4dda471417b4020d188a1bb77172d97c24ea3521a4c56056714cca3
z18f88d4110a73ab04aa3ddb3cdab05a691fd6fe189dfb93b4ce1798cd8993a18f83bb141273d30
z8bd466890a210c818ec756379e98abf54d70acd0b19b9068ae5d0702f06da88ccf36e1a8bd53ef
z99a731ffcb2b4102a3ecad7c041e2cf310e6f4638b4d96f18e2f2f373ad9d1afd6ea6e4f39de45
z0b9993f2f856f4e47d419886dacf26cc7982d4690f67ce8a887921dc0539952a6fc6ad583af53c
zfda5e5cb50dc1360fe460091adc6ec67a8fd49deb029ae38b30c403e37c3b71bc873e784f72b52
z6e95aa1a36b2b9ad23130e00230d224ced677e343f70edb77865508c2e6e0a64774e545f29c1d0
z8f484a358a179e1e9d8e1617343b2b3512f3367e70ac8ef21410ef644dbdeb6b3963b6bf826f00
zcfa49cce8018e283222e92f495239f7cdb3e14550df9d8ad0b2222b027749ac02a87cca90d18c5
zea9821779bd5b5d3ada4b4d35f6744f96f5a2a25477f6d8de4bbf63c40a51f0becb9cabe4b4e49
z235706eb0cadbd8053b281e54829ef45d5a1042ab6dd34c132ad2f140bcacb7a6550b489aebae1
zc626be85f57b19fa5064e88d2768eb76ae55ae30c8a602b0908466dd1675cf7dbdeb348d5e581e
zedae6ab9f9c2e40bf1af1604bf7a7149bf996df7331b953a40edccf167af5512d3f521202cdf1f
z0efd75e19356548ee5204537c55257e72ad3ce6130432c2948feac36928af687735941f9d897fc
z417d70cf707af15b529a9a9a9e626f73f5d0147db256e0f5f8f7b8e8664bd6b846b8e4e93b7e30
z144d45dada19724ca13f20d7efa6417910f630164d94fc571edcb039fb2bd77788de57751dfc86
z7b99d75c7bd50bde8aae8b11d6c56624f609f2a1f4aa39a4da77045d6ee367ebef7407ba240717
z7fe74040a54ee548aa941550f6ff9b36e192b68e4582bec7f324828b99be1b74e5246346785736
z48ca51bf961ae4f56fc3efa8c2c1de6f6d8c429dea7cab06a0812336424071213388a5166f388c
z5e1120b7f0b75bf8dc5130fc003af504710ce100ed87d57d2d7c83f63ffc0c52ac34465b557f90
z661a6bc485e4c684c6645e5e679ef5859e321e79ad41509b21f35cb067e7b9ca867bfe643267a4
z8d3857ebe89f277a21fc8249c945020546ecccadaaca2940a9d3e6781dad974f150ece6e369a2a
z885fe454fd65bf11b50427553c5b2de758a9f9805fd0668ee72ee3f5434c0740c1e6fe6561d5fc
z919fca99a201b4d4835b7c8a18816cd6daedab6e2c97b6e602eb4a3736e56097ae060fbafeb66d
z9a85c8d145f2dbd7292dbfdc5e42d52c3c54b538cd527c28754f3966e2866053cd1fe3ba140da4
z5e45774c4526b33446f92d6407459d4a23209f727467d857eea0316ddcf714dc2e84b0f3624def
z6531d754e993e00574110f4b1a5daf5630b65ce0093921edd07e00e378c315ed9d99d7c8818cac
z117011a6e45deecf2b2ca7deeb6e3ebbfda17a821ce9ae5c675cbece5f96d4fea53e167b1c9103
zff7f2fdff382535761a73af0c27f0c6d6c7d90cca56e45b3d6e85e1474b59010dc234eee46fb8d
z9e30f50905c42810d3514f79478f5002ad70788b5934df491e8ea72e81ebe985ba82afc7804fb5
z178e889087fa4a3156970fd6ed749c0ab33cd3e924b9d1c9cbe0fd03861ed02ed9dd70a37eb608
z86549cc8018a861aec8f3faf688818be07f50721f9d76faaa332c53a353013e9aa9d63df3c918d
z4fa5a9bf4ee0c81e87a18a67602871c4f3cce8c77db3e8d97cec9f0f70e183ad7cfb3b8fdd768f
z494b1a9443b54f999c1f192d807d26d4805800ceb40e65d08eebae9410f234e0ac1bf46c26daef
z569051a481b81e2058abd567f7941a843805262bae7533fdac6bd3423047c3e9de6049b4be6a5c
z9cf746a1acc822a75d35b964d1edfa186b3957440179f254a419aa2ccf35bfe5450d39c745ec26
z79098eb764bb5ecfb7808c84d729d38e1a1b51ba754f44beb67180377088ae403b7dc875798da5
z09ee7046f162e0e70dd73005bb1493b6f4d04986bd3242bb9b9fb417ee04af80ce532997f5301b
z135aa75b6338b367c5bcae0fd2e9c2fb80e81c7ac962fe3c63f145794a4c43d9a5780d30f20772
z85f7e4d88fc7c10fe8f4d13eee404e8fecbd0e2654df6bc364e09807aa80efe1d902b276b4df06
z69bcb3a2c1f6ea649529f33c26583af8ccdbb090735afee695c62f0fee26eaa858fa75a284d98f
z7d76cdee1084767c2434c39eaa8c1828d3ddd57945dbbac5e022ee46c5b205e01f7d509cc83982
ze976d9832e7d949515aa5f990f90592c5f82cf7dd90f18a76b241a28a2842f8bab964b0ca1b489
z6222ca38eaf3284ffd2beff74ea62c511b0caba19c13f8b18444bbc7ee234c98c4586478d473d0
z671ee485314266f1d1750ec9280658fbf004bf5ef1c1120e324479424165623928ee66e726c849
z455d13b2148ed5e56494b6e699b6a88016a67014cccc5872c5096b798fae6ae280d8ec278db824
z33cc6b6f2a7c66fdb44284538e2aa0801e5e7a1cc91bc6cc503fe42def375fbed128b23e09fae1
z229e6cc6384e8dfaf55e038fecd9d8e9efae2c598b3bf1a645158bb9a67664718af46dadfbb4db
z50b9d8a03531a96e95c61fb1c128d8872fa62499626ea85a72b528bef05e3b9a11bc77ce2ca61c
z22fa5c4d6d4fee70a2086d19b217a0a400958669b15b1b547734238c551c5c46ac9a2d53f3af6c
zf030d4aab9513c34f6fb758794d0f27b66aa0d2d72b689a002777b2b04438a51e3aa33c85bb4f4
zbdfe2afb059a9b1a3b9c59248d2d34768f62c54a9c504a2ba5f89e8f38f6c8a19690c19699381a
zd544935d14760bde14b366f6ad8301ca754415a1570e0d1c3a0dcae5053a52f9c9dd0e8755dfd8
zea667626691e0b2dd84f012e10c4e1de1d408649bdcd97da33ae962a5e9aba9a99fdf1e178acf1
z1ef33915d29a55c8c5a08ae168ee956fbf9e6104ce32f38c3043df6bc782502f9c02b886d558a9
z8b65e3a5986920f0a39e8b98666e58a5b67b17f10731a677e94ada2757a8dc3c0a65389a7b2876
z53b9d47242964c46325fac2125291d5c5ce77267e4c56bd4b5ddfe6d29ea473a57abe0d31f549f
zf2b9f38a2ea27b50bcdb78e156637903c2dfba1d8d3b5fdc9654560972b6d934096b0ebf3e037b
zdea3ded282b913621a04d6b1092dbd9b88767690237088f56d1c3a1088d1dc89a9c7b3d9821f89
z3247dd7150130def95859990a07f7cbd999c48d8325c360a988f011781bfa35388fb398da53f81
zc71566e7fd05e1098e5b13bea57220151772d825b1b1cf27e0a8ddd6770779bd9d3c298d1b4d50
z5a60bdfbb227fe9212f0e0e77766c52043a10332becd2b6f134169adfa708c90c122c51596b995
z97e52a91a612c1db2050a2f776a5659b0f7e46bb6e13955b52924242433aab255c501f8e803f45
z2f16b090185dc6aad918a4f9dcc1804eb8d046dd7f0068abdea41783143decf01c453d04c2510b
z602c91deea32373d9b9421c885543b8d3b5b398b46052e62f28a70c5aa3fbe7f00f9cf11411b91
zde42c5a8a5856fbe9996a2dd6d460f8916f39d9fce357727ed293c490b7560a879c151595a5185
zb3691ed9916d6874a59637d9b84119ed3f91dc6c42076e392e0e60ba1b0573a15b1182b12ccbe4
zb4a82c51040f805ae473bdf076cd3d88ff768cf3f8eb93c7dc61b535d62e32bd38a2492a9fab2b
zecdea2659f3e6d55840f0c2a85c52787c724ba61a07a3b09e697a4da5468c84da76f918271f7b0
zf12baade6bdb9aae2c728b72166fc8a2657f2657bc8e51428d35a29d7d475fe677945dd0a7daae
zbc132d88a9e1a174eba8096cf83fb340d1477fd7cb23f938d9424c32c50463fbf263bcccfb6f5a
zfb9f6819e99a597d99d334f2ca8d4e36f90bc07e09e95d0e1338108ce57a1d0ad875e5497d3d8b
z62270087975dbde3d8ad38918253f4caaced97eae4d8d17de4eb174f5f676bb0dd79dcafe362c5
zb43c4011885fbde82268742f6ed72f9666d6c3b186ac7e06f61e7ccd08435f03d06a640f29b969
z1c489f169f1c73d4ffec3cc73ad71866fff2830a241ba6b2717d968c74660c6c5fdb7f37a795aa
zd5be1e2737fdfe6e1e3744315e333a83758b244f9d4b7c89a76db1ff98517f7d79934d3ab099b5
ze2925b19db181a69f195effc7bb43095f1101050f3c2c01c6b3915b8e396a2ba2a24dd7902c01a
z9fc7cd4a4352c5ce2fae20eb3b5596d70864b5d3d043dc48cdd0860284d6994aefe5093869bd04
za9aef9def56f114ec1ea599b011657fa92f2257c170bcc68f7e107401edc77fa6183ca33cc621e
z1e572e5fb7d5ab064e3eee50db2a73dc1405adae25e560e6e891e3dfa5ab15d2f56d6948fe0d46
z03800ca4b86d45a1471183812edab43868371f03eab83b5d45bd78e0eb7c96fcf71cc984055d20
z533c81191336c123a547e4ac62bc007a12603317203a59ba89aba67a1a2eca535e4fc7347fc3b8
z949bf767b819ad4ba70cea6f507e7e2088aab36c1796c5076ca4d4127eb4edf3f59c1da1235a3b
z3c26cd65b72ed57ca3027eb3f687814922de76dd3049aa9fb8d2c2ebe44b5fa4d2cdf9b690e40f
zcdddbf6b4eb6cdba2936e077c2012d4028c67ba31a9841e16e201ec9c62304145fb40064af5baf
zc77c721a582e1fbac2cf8097f32c027949e7d45f12322a06d4b13a36eb32c87514ff71f6da4518
z55a88615bb4a49f9c13ca81d6ddcf3888396283e035792366609be778a118a934da05f5245216a
z9c63e95efe98ea630f9f9280f8464e476b154c52c4b6736c531a16290ba2f3e44400c43c67230d
zda4f3965ec744b2a7734ed7423c27d58211c1e09c71da9e247b6cee96ab9d556cf724fdee8f1b0
z0376cc91ca44494826fc6aef53a19118472ad1e72e0bf175c39cf18ce4755dd3cb596ecb4956d6
zcf04cf31620f41e60e0445fe4811dfad2af2292a8b829746e11b52e56016bd337da5e61cff5bef
z8f4c77571f22da55834d860329f867667f4301ec2bd8fb69062ca4c936631f51848329e38aedde
zf059043439caf982cba3cb779e89d2250c4de024c15ce85418e4f4926de41da3e3a7bbd420c047
z53006c58fb3557967f50efaacc269d9225e54c900f636635e407e6c3ecf47fdac947a98dd9b205
z29714938fa2f4f09e7a9abd61445e7ed0ddbe95a208ff21e8d3b66afba90f2c993a2257b14d5cb
z062df7c8df323943ceafc4b6f1520b53140f82dc36d60c21189cde9a57fb2e590c79389b25f960
z4a9f84b2da0e84247f0e156dbda2c130f49195d8015a40d5d8cfa06dbc729ae25c70ac6f82f135
z068bf5f293864d7d5d23168050e1e4d3ce27e6afad11070eae811ad987d91412453b935874da91
zbe47497293f5462fdacf75dcbf51aeac6476d1edd5b9f3432dc668d488d4085fd99b8cddf32bc5
zdca684cbb6fe88249d6e4f4051951c98ba83cb9a3eccb5fc274b5119172814ee6ac8913b32de0f
zb624a7245708a461641afd42c7e96226d46d3c4700b90911da2ecb774d69374edfdef8570eecec
zd5a94f344364dee219520c6fe0a3179374e5cce0da572470f92509654077d125393ac07983d815
zdd8d3a738ffdbf1c86fb762d3c55b6017e54ed98f684ec9a6c263120bea98b2659661c520c5097
zf3087c031f4da99d0ec1bbe37bf762b0afb3f68ac732565c5b3ff51aaf8e596ea5a553d95fb812
z8abafe04c015872b56c19bb779b31dcd77641513ab84dccf5680ee107270fd31976b8238015338
z73072c5d7547cfcce2cfcd5a00cce7270573ad88c7c0eadf87290153b6d5b35330af67ec74d6d4
za9f42fc9e62953928f85bd02ebc0d6882080e6feca9c2e33e6425dc55c55f4fa542d54b030673b
z873f49f98725052d7d2715cda082bba9891870c8a0b99c6d574776fb5786d56bf47b3f96c0c5e1
z4c74b425764f9abcef8efc76bad1bed8ae8a14f51436a9aa29b053c0e51448b9d23920f62b65ae
zd855fe11b5fa8d5714ba0ca0e1903b486bd96864abd6088cc79cf90622d33acc86fadd26577662
z0d7ccdfbc1f5aa9f6a77459943b52ad16c97113c90313c705daf91b23d08aa29a90abfa04221b1
z38f714edd8063a2d7bde293f68baac2e91b247d6d52ed6d0b1eaf8d785e7b6fce5bcb936a00f80
zc79912eda615b377d698acbded3e23a8943006a76dbc2cdf4fde74a3159ab860e36b8017ad4a38
z9115008cc3764d89bc93e017bd430da8934e38b0e358e9ba3fd445a60304afd95f22517177ca95
zb7fa75e4f0aa2f999fb6f3eda3d1ec8c55c13e98998dcd5c2265982f7c4906b14bba7040f82690
z011fd286723c2e6ce92a085ea851be5a89fe07020eedeecbf9436593a7b448a0b86d6d79ffc66d
zf7291e2c5925ecc4404815a47fd4fac7f332243e7eed510d20c6437dd5cfb283eda459b4fe99fb
za00b1cdbc3f011bb02bf211ba007f60f5a26f7ccbd0e6541f97871fbb3e9a0d8b671a65a2d92ad
zd5da53bf7285fb7bbc4cf3c46f6ab90356fd3f31c2bc5d12248775ebdd4387c1b6706d4bd951a3
zcb7103422f3312b77ee70029a5277f8ee47d437b5bc0662f8ed95603cfd73046ec3198b14a482f
z91175e9daf3632de21076ea7e1439af7f9c484a0498cf5c8b997ae34ca7c7dfd44a871937395b7
z79f5aadb90bea6e38a9635d6200ea759535eb09e2dd561b502277662535628633a4874ed3fe808
zea13dad68a3266222e9f38aeb027b3f1937ca0f575fd3e6b2d1fbbd57e7c68705b7fea24156a6c
z639703980e60d31159c6bef12127f5824ac1486b56fa4f6e98b39e5f69352cc57a437e16e9cbf8
zb7ad308c112d54d29c5a24747d9518184ebebb89bd002f08255d71e9da939cb41c5a19f6806143
z940794695f8056fcd34b5b4b31b37729adbece7bf1923b448ac1ce838dc641060e2637043100c6
zcde76848db4d136adba658fd9db3102cf882fd679fbcecc2d7947542aedf5b3b31217d6a0be2f1
z4b3592725ea318463753eaf1a876b4692563f8c002634bbefdf98a708c55e63331fd46a25319db
z8baf952ba002dbe6429374b36b57409fc873ee73f89afb9dad5ffc2eb7b3f836fc421259873c7a
za5c2acef4e010878ffc74d16a2a5da23c238c8ff52bfe83f042cb4f12ed820f696058dc8b48643
z25c434c0b06bcb1e8aa409009711003286765a4f8a9dfdedfd9e033e0d5bc12a03795fc2f307b9
zf8d3c2d378da7cf26c2d3751d2eb6acffe6f1aeb92de3e27ab3a5c7fda75eceeec490bd8d7c053
z16aa150a5dda50475a5d792c73c9d6a85a9be42197823f8cceef119eb4f0a49718e24b0f95fe31
zeb926f15b1c059420ef4c901b2d4d04536e778b95f4a89408915f115fdb11671f2d4c7229d91f0
z106700a1469f8c69e33ee9dd56169376cc92b6c0306b84675b0ecced0003ee906ac7d028f9e221
z610a0651becdcc6bacd3634998e2759ec99cda8554477275eac989e9c75350f7031c5c7ac21283
z73eee32d7242d5ff311fb774045a582e66c071eb9964116b83f3aaee6dec3bb96712f442dadb82
z1dda62be8641b97446b5fc165b65ff1f6d78a72bb18d0d1a5e640ae7bbe128f0f7332fe6c1130b
z8a8bef01f3991469703195f49e7f6c688af4dd44691c4e2ff6866dac30d74a53e1f1bfcae886c0
za388ee2dbb4675e87931464c72993a88509e1cb3fdf4eee92f66b0455c0a61a331015677ecedd8
zd32d153ec4eb431fa87fe146b04cebd94bbe7624e49493eabcbe7c225f6b1f8122573195cdd31b
z40ec2fd8404b6c28bf5256552dc4a53360672ab2cf823f56c44af29ac65c722a2449eb744a236e
za6fddca403e9d166d136038bdd6c5e4c668c69de1368c2ac49a7c4373468c83b548032f5ae748d
z802df87483273547199e640c10167046f6300f7aeac73e7af40bdd4969eb5d5faae6da6aa91292
z657ff4644d320da77068a961e98f086fad3155f83cfe22172269a02cbfac9c853a10d1e8c5c704
zfeec145fc0f8aa6937dcfccd6c3fb063b63241cf9a151fc82f439b7c302a55fc137d5fc836d9d4
z2a14e1f16edf5a2fb8edd2e89a60e68414523e2552f7a7b5faec591235878849a365310a331829
z30b0d19422e45b2a17c100099736813352b36995bfc3c659a0c950b672b4f299274ad1d224b446
ze6517399de0b20f84df9fc397431c9b04ab8a882a92d8584d8a9753ea7ae2827956dc869d3c62e
z4e90f1ae6028eeb26878ec34f2baf44a0909f1c0c06e5201190c2ad520796fdad88895851e1803
z7c55a54d9ddc5fd6d966d5a27ed13a81dc0421f7d8686349bcccbf13d1c1d8b2b22733579b632e
zef3a99974906ee55b9f102c8354f4b3b65af551ae3af332bbc12166c3974b8fc702b9c95c61d45
z48e63f6d26b1812ff11f1341418d101c83e0e27732265c3421c771da1b047800ad1494e6e25f52
z6081ced808722c1358f65407001a31bf9046fcb042ac6adaf0128dbfac21fc700f48a8e2a978c8
zc961076280a981f1553303b232e259b64594d3501e6b8750e84c8c5a086f8a125ce69f5559d862
z4cd6c98e181efd60ecf0e005b750441a6fbaf7ab95989ffc07422209d8d9d69357c16c7146fb2d
z61a4d3aed98be65b46c7297a79a67359f240ad656d74f4204a0fc8745833d1e3329ca5802a49a7
z765f106cd32f0de0d0b8e31df594c7893de452c1432ec2445eba4dcf02700439cd6a2e808919a1
za3d5716206ae147c7dde5f9013f4fdf29ba84a267424133f2fd94640650ae3d84724b266e0cdbb
z2bcb554c9254f584c067a6a09de2dacc77dc34d78cccd470165dc3317995aaaf4fad3a908f4152
za10073d91cac032f0ff741b94d92a798f71d5eaac7fddace4c5d47695e9bc53c16b967fad05f88
z4c5b90e49278204bd4e32958a8579e9ab660b8d7404e3f48d8d728204fdb117a2560cea3946353
zd57788f002572984d262c6755a23a339194c1dfb00060d6e7277004894f07e8a64d7976415a639
z02fd0e559bbe8d93a9071b5feaadb72388ab626a17e46b9de057f6eda69bad8f67551a699f090e
zd6e83e42c927cdb0b25403f52fda17c1c75d2ddc22303f9ce228a09d06144ec7de80e1bc457e25
z340b58dddd301497f95544d254e293b10972d160fe80cb675065efe64b5394b7b267378e18a98b
z1c11284886fb889807213c32b566f21eb7f4f4708bb2848c32497ea6dce498249506642053360e
z73fb1c53c171f353a6af8d06211f302ec652fb3e94677bdced017c6dea786453f0066c3d9c0d5c
zfa2752712463cdd21e30aa6d9f032ed1b93d2be1074b892493a26697043d90948848b063d312c0
z30b7965fe1d4c4ecc5f80ffbd4f510ac1bd45284d42078437a520b026a4bcfdc4b5aff1dbb3691
z1ce577c21f5d1145a136a1e4ed20948f4bb518fae06a772c2213c201518b0ef55e969766c6156c
zf5ed2fb6cb1482eb2dd01773f64a5fe550e68ddcf4fc4158840448ff05bc285a086389afe8cbfa
zec9c887332bdf3f1b38da51b58c4f737f43d55512c2bd4061742ec5330e52dd2f1d2cfbdadcfc7
zb83cad1977fbe80e405760152ef1c6b38c2909904af40dd1842dd59f52304cb7d56521851bf11c
z1dd6070993413edc5fa4e8539a52f02420be16d333a7f461ed546944991c117ea4c12347e2e505
z8f62c6491446c8d82edb90768dc76d8c7aa21a73f3672f333a82b02a9b92a215fcb8fa1c12db06
zb9e2138f25714e6691d471a46d23c901814f626bb52a630f346035b64c322b1e993696ce7d52cc
z5498595905166f7cb470a3a4529e6b8e0bd771b46311694d1d2ad5f0175c6fb254900ccfc3a4d4
za7fbea2d009ae14708577443f3b082fa2be710ef33ee76593cc22bb6f9d18cacd2508d2b94ca6d
za4cd9d62373115d57a3ae8b1d741eb0fa30f8ac3fb5ab3c0fd3cc895635835758a81e757d3264b
zd7b5125cf5eb3fa0895e4f8b98e21885e6612c841f7bb666a06804b99a0b45e1a8f351b6c7df59
z25a885219907ce3b9e95dfeddca4914730a3230f05b314d320211aa6dcec0404f4422243848f16
z21f704f8ebfc42503c7cc402e9277b7da93103f28b696c6888f3d83193600f479a1ec503b85f0b
z3c48f83e76b28b0e6da972070bab7ba908c989cdd0a0d85666e993e67b5a8d422934015f968f64
zabda3583168a2ff702baf6c9233a63527e7849c1ddf9f5cd9e7cdf998d7acab62a12268e4c4400
z1d04f16fe37b60bbd6b77418a22a22509a3adf89bf7a5d19eb589ac5677c2a2c195ac7d010a6c8
z584c4ca23b2313adbe2a92ebf6e51409300c23e49d64f56889c41d2bbad5e206733367f8148125
z7e86c2d81f0789efd3d5cae9051755fe52e62ae786baf7d7dde8bb7deb7767573314a8e2e97dc3
z9d7d8315dccad8aeb7f4b6c00e8d31dd8d130f1a6661684f6a0f8aec74d01cbffe2c9b92ef0147
zd887e9023dc582b1a3aa266b5fe840b0d4d41128e71e06853dcced532efef8150ec1b1f707d945
za9f25ff7333f37aee9782687d2456b7c98d664670cd87c70503fbe4e74ba359115c85e89314d29
z0c8434eff1f53fcb0a18124871cfd9e186726da4bdcf4b0a27b5f4e0b4949ec90c29a43009d0e2
z0561f04f927574e1ef5f888c8d18a7242fc85bce9a69ee8299ea6e1f294b1b7f0aefc1d66d5ce0
z7fcca19f8c2b2b285afafac38b0f96fe5ea6504a3f4931e29b5ba86635756de462516accbd228e
zcf92509ddf7897026c753a8029fb6c96332219d4345208ab7524b04adfdf5782f224cc9a685551
zf7962262cc7a6a916a8880a75e723ae1a4bbcaaacb69cccba8abd8c6417b28867fffbaefb318ec
zd64b5d452673e5b925d48cb7b35d3d33788c1a0fa2b25170b612fb13f813f8ab83c9c2206e1af7
z6d83b51d829e938a38ee28536a925b22ade1f07cccfdf53f45458143e2839b2492e3549a07dabe
zcc8c76ac7ac16c3a70b0109ba9a22cce5600e05685eee0109b3e70eb30601c89024260fd9dd760
zc67a0483981d59870ee41b80fe402bf7378ff1a86ba6b93a5d5a7f3bed9a1619b8d187bb622ffb
z2ea97cf46805b3bd00ca949402ece37aab1cfa8834a2130033f298b60254d92c7818820a737184
z39d3ecf4262cad8786b166531707b3dd261d2337d647ba2ce3cf6f8d230c076d1d830abc01999e
zd99f4455726c631b8d6302660a0c50fd2762d34dbe39ee896a969d02dd25261adcc4034a9f470e
z75c65cd82a57098a65c883bd90ed6e0672e1455766726e63b5526b947ccfff983e4dea037a1a72
zead77c50eca5b41186669fde664f7bac6c914ac82628bcb56c597fe8955f57298bcb84b5ceac96
zd8ecc86faa346c6e59f5f8e9fe23917c5fb66f84ecd2b357ce5b5a089703840f432880c462909b
za25d0fc392caead2b70efdf452a9eb0bff0694de362b397650da81db83da1903935565db01b991
z332bb5c76a0eaa28e76e5c997c80d1cb91c1e058de64e256dd391dfcadcc9429a4165145976200
ze685a0de0c68461af6d54568fd69eccd6bba8ee90ec662c2b3e0fa1b7a33947b18b7230a8cea9c
zd7e1e37a76793d32556462213ef0349ac3632fb7d99e3aa572072d1c3018f3ec07375641b5c9a8
z0347406e3bfb4723ff1a808dae887c293d43d83430a369514a803aa38efca28c4e8e11acf44df1
z6d7086f68fb67382adc15472cd05bffe91b718c11c2d22f54dd8dc478235a136d5a77e5e32da2e
z9aac708956262c9ff351814932a8f74c1fbcd22b1c1f20ca50368f229a5c3f181dcdca41bd2f53
z9c42dfd1c032fecc3791cb781c21b27e65d3fb8f48b0fed9aea1a8352848c57287336f4e33c038
zbe54dbb36ab4d9e5aa10937f86e00d6bc25c29fd23398a1116c3fd23e4d19d68c07ad2cc3e4854
ze6c38ae1cb133fa241eba38bd25ed5a4c7f4acf00c6be0712f154aaf0a9fc0c3d015ac2a866467
z4b713864465cb487a827c76e871fa7df3d94b94eddb30eb24efd0defe2275bb222538358d9b96d
zd2dc71fe998672f1fcc28334da3c689d3fcf9531334a0ad18904419f287df9b648d2e2796d5923
z59cb4ef21d8e0b75b7d951ceb99f5cfbe8505cdfc35b08e383d2fce6f71e7875a38ffb3cb2d3a1
zb976537d865a7a10437ed71ff5719e52d64b49d469b9727317a2c5e645544375f8a3c69ce283fd
zfd58347d1a48253f3507e9dd7c7e2f964e5465570599f0c20abe14bd57898fed2547394eba60ee
z09e230acce3fa85f59e9c5d1a6af94c136a5f37f2caeb0ddccb47e6a23939158120f3fd157eb3c
z58034bb1bd8f7525ade6c35dc05e691ca54c27be7f0cf6691fee3d83296539c80313dd56c545e7
z829d82fc832adea7bd106ea6b5c867e96cdd807085f326ea56f0f274ee47d63df52682a4c27ba4
ze4cd691b25cac081835d59bd0cf5b69e9b60960caaa7e2fdb8da34228811852b7dcfc128e99978
z423fb6b803f7d044e7d2c9e437944efcf2923cebd2a1510fbaa72b83bb768dd984d45dd95d1b6f
z2b05844f0b38b44eb88fcf22283bcebfd2f80eeb3fd2bd31594e248c622a509d760fe9108d6bc8
z81e479b50631d258b1ba3688d4787d50aee341a5c4a00f9da5ec712810a007f3e4bf3338817c76
zf98f0b469daedca496062139fae8107ab4858901c0c65176b7455ecebb186b93d822e8ffa2ad56
zc662c2dd8689b816fbce10598bfb793fa46343037022ebd2d06b44cd44f17f1cbceff409ca86d7
z8738e940691aeda9716b53ae421aa88fdf90f935f879590611c0c2728ecf148491c2d4bac51676
zc68ba440593813821f136c2c402220767882febb696ff9692cdec8a831de6ce1d82381be56c2ec
z612ac6b9c7c96a38a166dfa48da48bf4e3235e31cb319f539d70d9385d89b62f76dab6fbdcb30a
z139b1d6585b657a30977c2f9cd42a63890212b8b6e8c4d0a1bb31375f394a866b7c4bdd5c3698f
z36e64747ff2599341b31caeeea5bce5a90988129c8986c257a9f2513c78a358236826d993fe7e7
zfd290b5d9d7a41bc2061e19215482d9cb896aac66f1f811c1c0feea722e9b566ea5a02bcf008b4
z376106dca854c6df0e996e0b479f7e512a70ee867e83219580380f5c8e6b2c62106a510949ca3b
z38ad68e05915958e48eb3b45bcc6c1d6e4cbc795bb6826b503c7c69f77322357f35e655605ebb2
z6e50876523bbdd48a0cd5be128d884858bc3f6503ea4c5b4300c89f3925cef44187be63dc6d2bf
z5a6bedb6ae14d878c8b91c905e82f52e6280d7d76883a7529e8d4bdf10deec02fceea6c3d0bfe1
zcc60b05847ad538a8fe34113e1d70985ed9635cd958f6a4c295a451a1b8b5770c91513261e633f
z3a6787ac05591576755d01263d83a42b12a6cbeb9e1579daecfe49c7f2ba000d739c2652788f10
z681dfd518cb756ad412680b6973ffc6dad233100ac0be9d09f5ba23162ef311b806b14d34aa33e
z63963883f5636c2cf2c90077c68a05258966a21308d001072cdbc553ea61bca93b7e12bb946af8
zb258ee0d1db21ed8a22820a867d940d68fb0c27bb2ab5c57b0a242979b0456afa0b2bb1a790658
z4c363898c585aca0c15532ffb14df7f8f6e09a9c404d3f6b7a487be68649095819f79dd7f05ebe
zec75157924bf5e2b0269c7c0760c299169108845296cd6203067e52d5b5c137f31cc1904bc3f96
z7bc1e015b96c5439772fe839a0d227c067190d94def5a67d5f8a8aad68268857565fb450752c83
z9b46f8d010785f5088b6a83d314706dfa582aba769463f899720f9dad5f55af4db8376659efe00
zfaf7eaaf2a6a8283a6a98e69d71e4b3df2ff4d113a44b3bd502c93c21237546f4bf3388f50e7b6
z5fa9d6ba2e255050caac85445fac81e7f2a5b3ed1949d59522d40672b069074e676fd7ead931f6
zf8b0682292d3dec09ed42e0cd4bae37bbd51f0c641051c5d1cadac43ddce66b74f93273e1205c4
z30e35c997224f110da77717243bf7768c2f69af88a2b3495174e0037bfc2c1389a502b4c5e0980
z0156e96d0cc1f832ff0a3254ba880cc8ef74087adc31ca55613ffdd36fbefb383d3877d30c276d
zd2642e78016f9c71abd5c59e5b3056a189b5aa5a829f6bb85e90448a34a6d053a474fe1aa414bb
z3b656ec60f1458b61fc7be03badece64afdee5a68b1b3587c8ae3637b0124146fb025dd2f1aa42
z254202a3004102f571f831a2684c2268eb0ff88d0b59db43e279b13a3c4d3db97448069d8b48b8
z1d4de27695a9628e83ae05e1711e7dde490951484bc199db2a6d3f4f456c82f5d1686f7f309e8e
zd3e5def5f8196c1b94729bc291a2a2f2e467d788db098b5e270eebfebe2dc36b27b9686081295f
z79738e8e6c61190f2f60463ef85a4794785d850ffc3809b47a4c242290b31d790879fd4adb7310
z69cdc70437977a94cf803be72e6445f0267b4a7c8d4d840b9e6f7ffcc275d51377ee444859084e
z45eafdf921848029dfce1c6d0933c78a54bc25372ed6359a2d6c30f9280bd837665a5f9ab489ca
zecf54f7e19273bac7267ef222f39450b60ce5b473f6b4f4fb4826df1d21f9bf6f126d5078f2201
z860b0ed54040d534ccb3ca5a5c8636505c74a410f09968f3f437c2da60687977f1ec408c453d39
z926f77729ce542b578abc9ef16bdf8ce6827da5618c4ae0bba03cd873d2ebddf4cfec10722925c
zea02d3f27302c95db8366395ed08407927f5486f1f4134020b160aa5c87fcb0da4ef06961f1877
z169dd39ac5dc94dab8939e78b8421706e4f1058831511c025ab816bc930af8f150708433573093
zf523ec35ae50496e9c5deed39dcd124400058ccf3d0f1e142ed5c601c5fb34a584a277fea8145a
ze3f399b3d789220315e0ea08cf354b5861d21d5a14b0a497fed569d5aa6cb1caf9df6aa8208018
za00b739ab5f9f45bed7595881d85c8b02a683d58e451316ce416bc25a0e157c394e315f3d9e44f
zf34d80fdf4fcbbcba63b5a2229c9191e7c4cd50026a1e63877b939e28cf5dea288aba1b97c9951
z0a462284d8d0655e831b02fe7d5de384162da9ad929e21d253ccc2eb2f80a5db617ed72fd692b2
z491bd73d4e8e067be09926018c4b04683dcd855cf86780d94839308ebc4e0c4f708d52b0b1c4b2
z834de3923aefe46f1e913ce507a6d7e37c6dc0ec4ce452ad2d80eac929a1469466453d432015c0
zc54d82f31877f538255f23064e7f69e0213aca2a8f448a3370c4f827da8302c7a58f59ba28a625
z51bf83d7c4b2f5fc215e15326da79667d0e928a9acd60e60f09b1b9214b4b7473c6d450f9fd1cf
zdf33fb7bb3fb4e4a6d6253ab232d6b5ea645c92e5352012ee71a545fd00a9c503eb545905fae98
za00a865c6432c4b8591b654fb4a60dca4cc3f04b8c3f593b72bd9cf52eb927a70564587f1e9d7f
z26ee271fd26a0c0c0da49613da66f201468f97e72b3b94963fd1334a3b41cb37c5af6dfced8485
zc8a47b22e7becc9111500508f5e9fa93f6e52a584f9e3d7988be8d04ea27df12aaf053bcf7ff28
z64acb0616197fe02ee959d017fe53297f2c0d2236d28ada316ee0cde6057c140bcf0dfff43deb3
ze69683a8e2b061ffb2d835698c330808d2ed55f94ae4203e27c5320bab26037bf531ef07ee724b
z77890d66c9bdcbd5a771aa0ad43562ab016188df307c1c55aa5eff2833eecf9fe8489fcbb44a20
z23f2bafed0caa570a45145102b3a178bd2b6d3d5150a2ec750b5669261a67c4ee9257c465d2d67
z7856478ab554cf790abccd303db18646aee67a4a2348ffefca2df99267a91117f0f686f76e157b
z75c4439f42e76788b382f29c147419239cd141b4e1384fa94b4f880cfef876a88f3626976d392b
z7e57018deb9de64a7a75742f4c0d0a426dc1f67a288620087779905e299ad8c13f22135132c6ef
z2aef45600cad2d649b8876df17678ce6e3129fd5c049e76264ac337a06a548d50285dfdedcf251
z0c933e93d178025fad9391562fabfdba748131e451f7d6db4753bfd8423304e510b3bb4b122e4f
zcd44b9f2acde12148a26cab86e5a8210523b54166c3d43b401a41514da613e3999dbf701171f4c
z1e7fd438b3c5098bc5c063e1822c6fba5ae2af96b6f034880fa2b4a21bb303ce425b02dd32fc6e
z04ef44e01f7ff4f66ea3a1031d2a0c826be251db4b43558437e6c31a8a839494451823ade2221e
z25449fb8775126bba841ec3ab842724626724060bdc9488006c88fbbdab51fd8daa9543923ccd9
zac46ffd8de8778a2cf132eda15cafd46b78f61e9ea4d8ebacbb5d4610e9351ed4274d242774bab
zcc38a7b35794c9dcc822d25c7628fa46057d095b610aa91a43df99c091926541388431b2b54282
zbc9f3a6a5fb36eafc757bd98bcf0f2f8bee3932266d92469cea6fe1d83ddf479e26a7c9288118a
zf4eefaa03b2b0b57aee001b8e5f223b3b11707990916eb25de72896476550761f5714e7d0572ba
zeaf6844ec40bb2dd61daa3443000b0ad1d84f7fecf88532ac14c329249d03afdd004b5ab95280c
z474cc0f706094f2315a815981cede32db977e9024930989b099fa5c9668df24f7e2afe095219a9
z935cffcb9a4e2f5734902d133b3205d4df751c7f5e323bb1516486894705ef1b8c96a32d1390d5
za080d1e0a821b592be6e832febeb7d368b52904741c5f4efcaf3802989b160eb270cffbfc1423f
z204a429d5dc92cd70a45f54ef7f3a427a7e16fed6d07e84c9d3ddebe7a176c7d8d81a1083e1b74
zcad6205c2153fd062cd3f2095707b6c0625a47326dda8c6613433580054299e3d60e7245bb48d8
z4ba9027d12d54c57391a5db07e45888f50a4cf6af4faa2658a8de77928405b3e3b639b439b8996
z07e704dbc985dd1d7d6ed339833938cb9a94d6005889fd2ec02812461c335e21d4c7d32b2614eb
z4a11c521fb96b79c35782069a2b73667fe93816e3e35eac1dd5fe01dabb478820158dc1f09b37e
zbdfc5295f6facbfc9b03ee73aa1588e0c34890cf6a9b904a9872eb604c8fadd4e834bf7593fef1
z8eaf401bad6f9207aedc14613278281233f8288536985f2213eb8985b17454d8cbc478d38b09de
z99b3a22dafdae57adaa43af0c2778b46f2c0ef6b1b2cd3c0d730e12fab6fed5470a71844c5b7b1
zb461605244afd08435d3bc66b8f8c511593036e609b08599c0468a5e9968925a82d4f8fa11d3d8
z21177e4b7e41252effea1f35cf840d8d81ffedf45bb5fb3794c11d434bbbc7f979c23694d108e2
za496d2b7ec4bc8df5aa8b400ec12cc156a415356cb00d283bcf0c5dc442b66b65e32ae9252cc2e
z7447e28c0cd60e8630d46e3c02d1cb0b8135b464c3b47a2002cbf6285512e0f0b099e73f05f5e9
z8f6d3498b0d54dbf9242d22c8fb4646fbdda0a9d35c5355baef4716b8f03afee136b613684c22a
z422fe7a0eb16d70e8eebfac06a965370987f4f94c85f1bd6fbd62b43bfc182b297aab9597cc128
z085d8b889767f88f948ec52609e1e0d1d67862378970a18ec4309f0cc741a9207f4692d021ba7d
za62ffbe8ae339671788dcf462809a393d4689fe7c416a5ac7825e5a487757f0b4459683e516cc3
z6bb4282e6634867e298f4617d82384ae28c54c1d92a54a1f36b6ae7e524251fe7b2afef9c5281c
zdb4a74b9c9975c45cb836a4fba7b7ca77181213fbf953f84fdc80f36ce50b899c9457c13f74a0e
zaeba690bf56c5e7f74a825116fec31f112d06afaaaebf856df179c7c7155e24aed0f4cff127e56
zb140115b4d2669472cc4f17b50b9577a36948e71b09f4bac683dad237d208c048175d552b5d283
zb5bbc183f0a164777d4fc44c34d9268895dbd792941e72c4743122b64b09de5a40a84fb28a40ed
z4b629858236cc414eea433ec2dc53dc4dce4a566eeec3e1aadc1c5850068b0abb6b7bf0ed9649c
z63353963841dfb070808bd4ab79c921b2aceac4d91494cf4fc4a074f071cfeac64abe8afd1144a
zb2f0974fe8551e42465ac574c118880ffb5e0ad56263868546ceeff90f6ac20a91341acdd3c9c8
z108a89fda0f29aa77be4ba69f177e8e6d36b9ea8fd5633db6fd7f2d555c7227e608cdeed8c4cb6
z0dd40781ee29bda79738b66a7a50a9202f97b1df7fefffe97de308d8234fbe97ffdf252e71fbca
z8d3a128e4773d4d6f722704326f895bb5aac1cf08b9cf48d78223ed39a269e77c3886ea796738f
za4758b2503a690e9cc82e6bf715e3ef5030811a60c35189ae5dff06b7ade022f3fcf9193e68ad3
z197457d18af8207f1bf803876295996c17c275dae7c35dc94fb8d2a955afe37e5beacc9acf2d4f
ze52d730aadf1c483e98eab8f74b6ae19a071a0dcd192aeea323d6cd47e3e9d4bdbcb22209b1931
z968c0cfd4c0232ea4b574f0267c9865e8cd8bc533bef8f32447d34bd8e3eb1bbf71fd090fd13c0
z1c9134f1f452cfcdf287051b3561afe4aa6ad678d39660ea3324748160401dbc88982b700a18a0
zfb3b61a881faf9522058a62d7014f9ecf5104e354952baf790db2d739b811ba8f9f49731622b65
z597f54fc94d4b194e74b1ade5f12fec1d0498626ad8ed2dcd94a66940e5a7e682b8cb7a6dfd5c9
za6a746b971d9fde7ae455bd139deb887d364062e1819afc81d6e95766863dd8acc515d026b6934
z67bcc2ee2ab69597382d0eec2302766dd18ad4cd26d4178263923c33fbbb833656b29f59d33ed7
zcae4806f68d9d5084999346eb88400e989aafb4f3d751341c0746ee479d3dcca7b9b566516b966
z50e0226aee15649df94b61c578311bb7591ee70809af1f70299df9ed5e4da9371f0319cfcec276
z5b901bd13d1f2aa83e4d1a58198c7ea58e469d051f1ffda40055a593796648afb7dab6941fa1ad
z6e50edc0590ab91edc1c88cc10e50bb888d065611d0b9cc0d0fbf0d533bed8efcce7120d453d60
z0e6f4c492447d96729e05848775801b0837470c14eb2557ce1db3fd5a12b1c5cbb72e46777dd10
zc312364b64f90f9c697494bda20910a890869a03a97bf311b9e44bfa0d06e39b360644c5e4c13e
z5eab00e49af320194cb171655339489b535e8c02ee9a702d55729585bd1bbd11fa4e344dd253cf
z003476a8b8d7b297fa2abf077d6bbcca3c7924b7c5c472ca0c816f3ba48ef8bdc758ec54bbc48d
z5f258f44825ce538829f7739bbd59f1ba453dc6a41bd6b90614f4108b68eab52ceae81ef258a93
z001fadcf844402743037bf7f7b66c7e06a434ab306bcdecd8482e15f2b63af22529eec0c46c023
z56276eb2795ab8cd7b7e8a174d144096e20037697b19fd4dcf254d6853ef4179f82feb8b888d26
z5788c8eb2c43911d85c572c2e72fede7b41751385d6779aaa0ab61cfb0a0f443c13fcd0cf0aa6d
zc8c995ed44519eda5a4722182a8553867a35b9d83a496135c5a9cd453daa4eca1ccb9598163e28
z5b21d513dca4885b94285de374ba5a4c10d8d27e710160a4546138b3741c4472b86be54bc5fc9b
z9ac03b5713a7b6135e90c1f09e49edd0aeff47f63d0d770d969612431b3b5fe1ee367f719b1b99
z212e1d4e5d6ca72e08b7815f0289e0d34d4efa6ae3fff139856d7794e97e45dba080c2347b2111
z78bdec839acd4047bb805ba9f897c09fdf3ad5c5a3dbd7ca42782a3810b2fef9c5c4305c82dc20
z62a9df12d7fefe3a2db97db57c7ad5b6e46e1ed6ebba2ede21bf5794c9e17290073c54496208a5
z8c994676ba62ce8782d76efca7f58ceb6235599eb456c8323fd67f18422a9cebcd48d2b06b1eee
zb62d8c50eedbbde04dde896187101a091f5cfe528a1989387b6cf2a4ee34d320ec2fa5976d538d
zfbb6d975339af72f04b0372a939158630cc86b0617cd5769aba14260442bde81f72446c7b6e0f5
z5d089addda758d6e7fa967cd614433c57f2bf50ad442e96da69e2e5085aaed45854897dda5bfc8
zeb3a86ac91aaef3c17349a102e66318822c56be829f94f9b42faff1cfdddbd912fb3a9b863a2c1
z56d9743b1a84aad7f0a70434068fde69a946c90b399b591fe91a3e8f703f00ded448d64587cd44
ze1987756a42c1166ff947ed1857b1d2e9ebb503ddf7df5bddcf75eb0c8fe867196c8a0d3298fae
z30cc1cbb1b78ea974d86d541ce014d0fcda15796c4663fb6fd46cede1978128e792f83b03f3e5e
zc53dcf54a28f5921caad4f8cdd27cd56f07058ddd8fecdb3ca68b86042addaf213d916d4c584a7
z176219ab6a434561d7fec168f4cabc616ac3964b8d56fe7eeb8ac3138167c10afb76ba455a8d8e
z20afbc4485a75c5ab8e9b12b6f6a1ad7fd19f6af07d4bf9fb2fd75ce75bbc3569f993df67b3f2b
zb31e1f936a7759601b4ec349cea580ddf3d0aecf4341697e721fc9f24359e7511648fb862dad8a
z5908ec1d29264f29e9fdcc5b990892c633958cb4a77eab8c0ca29995c4a45c9e84cffe37eb4996
zcaacf97ae11abd609d3f2896da1e9d60f413a64f7c58a140455430aacd3de4f471b32dc54ffbd8
zea28d597eae78de5b50c7a6158dfdea8f4f15858b2151fe2bce661e7fc6bc1bfbf915d3242d4b6
za9c5dfb705291be48d0fbf851f89217da4cb111810c281024b80cd26deea3225975077f59f4e73
ze3fd28e33dd7b60046ef74199a17f1662492b80d29e070f8039733f6a0cef9917d5eaa7f4c2a79
zef6bee59d194e338bed0e42a5aa40cc8042871bd4bda528333143c588377e1717e6dbf1e7900e2
z5aa4223c40a8a060caf0406b77c99651eb9cdc1b1a56c7243a408bc69cfc16b2b4a87309f0f61a
z519aed0cdb12d223514310dd08d670fb6e60e2266e7d729854d92d7382d8f6ae3fceb4dce01c21
z6891d0f639532d7830fd161a4e2d4591b99434326a9deeab5e4f26017977f1674d074a41327c5a
z85be79a7436f1d60585fa40dd3afe404cb03ad38597cf6d22b35fb3e8d05874aa8e9e41cd06b9c
z397b4118c647b1ff9cc2cbfe1c9213ed11a6b5f65ca501635ae907feb149459586814e17dfabb5
z48fa6084880373148751b2c389b8e9ec52bba6554b99604c653a28dec1c7a3fd76b7e191a782ad
zfba3ad8789c754470a59014c15e43e0e98702ef0da40134a88d864e1dce616282611728756687e
zd128a4d3771124646106e1f4941c70d7792a888e037a348c49a26be6737d66b4af296349f538e2
z077994ae26a40a4f6c81ea6fbdf8c2a0714c5ffd617c8c1dffe7edb361b839f815127248b1a6d7
zb1a951d06c3581e7af4a2472dfa93d3575f5ada61e1c4c1e8ff5786ac69ab261e3cd7b9bd4cb31
zddcf1bda6354345c4f4b076fea02445f3f68897c4d8cd01cb41997e60f020b330489bc8f6f362f
z4f8fd18e506c3864c4c4da0e83e58759649f03af40916bcef66f508cdfac4c57f58bfbcaa2e47f
z61208a69cfd8b133d70820ea9e3a3422145ad4cf33a8f554e254a536cbd55bc6016eec0bc30d7e
z7d7b761ec4aff9af11fd956ecfa51f5c68c85707b59465ea323c589e1ed4448783e2fed006afce
z3713ceca180d9344628526335883a0a1120d5b32ca7a32accf1884e13b5ff97c2d273d72cf7932
zf5cae3354994798ba0d9128340df5b0bce66d35979c2f621067c0619feaf4906905e41040d9a49
z79c1a3d2bbbd99c2e9e9dd828348e8688099f3facac6b2eb7119cf9ee2b77120b4e64dffaeb2ef
ze4c9010fc0bc5bc56126a1b553e327c980e5fa74b10457de4c089dea0cc9c2250d0c2311a26347
z1c14bc88bace002602878543354403e5b5f8f3c68dd4ad3acad5b8628915a59c8c09e548bce70e
z77e734b2efb8e2259069576db58250d4699c57f90d567c07c23caef71381fa298dc4770536831a
zf2d128b21d919a363938393aa455350e4fbe8131a28661b9b4b219f55070f659139ce532b0e85d
z5aa7a52a47539addaa578edc67845b6f6572fbe3037617f4b49648745b997e96602ae8993deec3
z02dd9819c6f092fe6db8ba32ddefd4c74fd59b4bcd1932bc1afaf6b82f755c1ed8679a8ad8f391
z33becc01a656bcd302ed0ad2fc647eb5827d13945e934fe048a4a067e8adcb6118e92d481f43b6
z0775f3ad76b4f1a826d47de6e72b69fc188733de7b2f70f6dbbbe54459a0c9d243322b48868cfe
z15d94d8479a4a103cded3ec1cdaf59c24a4ba17a39aee22d69c38b519fdf6cf03983ddb18386d3
zb927755d13076ea339e742344be3ec5ac052c6b129f474438e3d21c655e911544dc56d44d1cc97
za734ad3f23529e066afc2d3779f206f356d9ec689ca7af8ff8023c4f09adb2687b6de455f8d644
z7d12da51e1997b27e8be5e7ec39699770e2a19addadb68548151484ed1abeb1bef966c7996db4a
zb821d4f2da73cd1bb9a425137772886ba5d9edfbdb48977f344ba961daf4d358c443503cd15058
z2dadce1982258737480004a486934edcea7f0d0574fdc4a14b25ec9b9c4fb6124542c5fbd5252d
z8517e7e5608db058c9bf677d03f026341c55b3035ba0b3bfa5d398956744a8f74055cc06adba92
z25dc567aaa1a23d47ab9d64a5d8df0cda98876015e281811973d07c1fd9687e70cdfce6b4e1c3f
z884f6c0925ecafad0c9323f9185bea5973ea3a4054c723e98cc26bd39a32704cec97e2c19f5e87
zaa1f38c6619f2b1bea3356e69673625c01a419ef7c253dd41c39160fe5ae576cd0e038092baddd
zb7a969a56d36b1329587f62114464e06c8e88cf1fbd0bde9617ad8f43aeb9be87f89c50dd7d2fd
ze794aaedd5de4f2b2046a041046141ed2d7f68c4d3d1c53c542a997091526e6de8c89f9fa9682f
zab35e3bd7869bc43a75e91fa2e5cc5a57f6de356fab6b58089bf6cdf8f6a2acd07aa0d738e517e
z57c1d1b1ec19c44fca743c06d236d1bfc64fca8c02581820d4c56fad460903437f6510e1eefeaf
z91ed9415a8fc68aa10335c88e657d9b1f3c19de39fef487996798b0238f615d490b6ee789ebdd8
z2292ec29fbc98fe0acb26db425fc276793bf7efd9f59641e4c7de1f53b8fe4e041ea91306855cf
zf35a05b4dfb848505f93db79cd8648aaaedb597caef47cf4708e66fb667bbd510bb3a04746515c
zbbe994fcd67339cbf5a7c45467cf894138417e8647327454f0e478d3307da8a4193c85ea1dc924
z1ae1219ff3eaa37f6bff687e6724a80f326972cac1f3464b8b82889e0384e42a9145728f574cd8
ze8bc3534a4ff749016d4ee295693c23306dee830b3621b789ea4755f54a388a8feff2db32fc1c1
z33d0456a52529426c20c1cc7518ebf63116768854b3c87224aabeb8aba03c3738147e046c9469f
zbcd3e653d74579ca964af0019a17338553ac74c4bdee627bfa9671a3085b650519fb30e6ce6f76
ze6e515b72ee02f9eb1f57eaf9f1a90eb0b14914bddce21cb6b29942d90bfc543c480d0652decc8
z9f0fc228b082a153dbbec3c33c1de1584c285f1186d0d6e3541ed94fa34ef655c3f9b1868b285a
z69cafb3aadae7563269cf9348d151197019904d5d1526d4deb3a89bea02fb025ad0de16f036a6c
z258ae17b56f191eb9c375e365700f60bbc3981cdf98aa5edb22f3e88e79b8f4ac4ee2af548cab9
zb18fe98a7d6f27db774e429f1e464b31cd8dd9e37697be6ce699bff7552d61cfccbb4e01d981be
z20e26184654729f48816ad697d881cdf2f32da7ff14dbb1c1abeaadf16f9c129e83b42e0e8e2a0
zcf152f94c1db1b51fed7dde62f46455363f92bfd686578f8b29d26ab90a8116d7df4044daf377f
z70c7af38f5ce6e885db97c57b1fea9550778c2d7010fcbda36b66f10676b26e253b616553e4168
z5cb397c51d8595cbbfaf2d257ebfa9030d0d9c298bb125ca611cca6b47e6492897d99a2e5b6941
ze209e038de05adf9e99331805570cf087119da0740362eea8afe0338e53be93a2331e8c81ee7bd
z7db72476a6dd9368e5dcf3f8f26dbfa6547e0e3321afd25b5ee287f50f2309451654bbab04f6d6
z001a7178ba5a22faac693fd6f0fbe2e24f4d7b4db7e83356c44b8175d5b74c12d5f3cbf34459a0
z6f6837e33127f1595ecdf4a96fc0cbcaaf8696ae60aef8eaf20e8fe95fe74e56c7e0c9f0249aa0
z97cf16c3ae3bef9fe621c47bf735600696e40bb21a47ab69bed061071a304eed5bab07b85bef1b
zc075cbb3a3b1600de37075ac693b5d9bee545b8955745fdce76c92e4d4bb74089fc4eb4f1e4fa8
zd3b8365a2e108a930aba4d102a0a0da7b8f6b7b131b5409b15dea335709d39cd9e1906f4d83b7a
zbfccd5751c82a4bc6666dff7d9740dc36d30ad854e95a477ae6e617fcdd382333a236c70864e58
z685f1b2cd9d5a1569e630e482a1300cb45ff6dfecb389b5b7b5e3784b809be7269a2e384c97eae
zb753cf7394e9bbcf0ebecde2da0b3e045176c140ad0b6012e54ea4bc8c96ceb215f857dba12bc8
z2e3d631c47521484c2cb22db548a4bf0b96cf03fe0de109bdebff4a01560cd2a7cd48046a9aed3
zdc6f628ec6c08e2099d2c335b719e6a7b906c0a43366a76f27d1a4fcb4acae687cab27a00e1cac
z271a1505dc0f4216f3b5700da16898f88302fd1d6a14edb3d3bfc47cc3e74bb3355acd94f3488c
z41f2ad709e40f04774b7f13511de8f99d4bba85cb0c3a226dc1ddee6a9a8a23c1e1eba5010b6d6
z263505d045237b9b25c733256eb3484be631cf982df8c3f16712de2aa8a0bcaf08ae60cb71c7d9
ze393d08dc8fd658c3c32221e07abe3e27349e5e181c5bba2d211bd16dea0249c541802a17894c3
z09c2de3319d4061fb938809bb7a596bd1dd0b649d326616e379fb8e4c0a6eba320a3b61ecc45df
z8bdffbd6aa3372be546efea278fbb5be624b322ef0d2417fe0a4657a7d4e709e5b190e0429552e
zdfed8ba67a99d5a431c17803aad65363187efc3adf50209e6b362d0cc9e717b9d0a14fd9f356a2
z51c06b1506e3a348834b38bd16a685dd8114279cc060b0d139a74129515c46e83f75d208641284
z389577c8f1f3b0ee4f3ec6a0fbe031b70acf226b1806df34de757a66fc063a7783acdc944bd691
zf20b840fcc3f4158d520b7fff2389a83bcff091ac9265fac707ac8aa3aaa48587bef48fa921ed8
z98c61180fe5da63930d8e9029bc17401cb05c801b233e2bd1e6f6c3b8eaed364b095f5df7fe9e1
zc19c70face455fea58c79f01d4600854a0514f15b7917cc3c4f73208da77a787bd69d290c29599
zfbe0d5d2c8185b64f9d314509362f55691cd8d842b439315f8455405dd1f58030fb18b8d6f8447
zbff50cbad741b14c0cef98d64c6e741ba8c7e69335da184c5828d8f48dbf7ab62dd7420f5f4779
z93237ea787f23f62b85caaf805c5d5f66bc3d5aa97884f5b568a06afd2d50b02549473c1d36b61
za8f22554c6a95a4d7961fc63ce2cd6d76a33985ad38e0c80a5e53cda4acdcd2bb3fba82ea30f81
ze4bbb3a64c29174aa0de272f94a336947e44abe1bcad18724d8923fa98370e3967de8692ff6408
za625470c080f8b124386aeddf87bbde0d8c25b86921d02eebe01a917779f4c2dfef0892d15c78a
z7b1b969699df57f4fc24bdafb91226f27ded53f0f8244fec5c0ea89f32219b70af741251ccf70e
za3453449cddb3ad367c80550b7f6e3226fcdc26e7c526304c30d2a7ddf93baf8ae22b2630ac148
z691dd4202bc5b14aa2a8a4366fbddc5af1a9b2581a86f1d58743c4b655666cfd126360113672ea
za9264e873f8084141b53eeaae62e715b89770d084b28848a1d6779a42fcf4a549ac2c6e882dd62
z55357e706b92e2d5b86c0875747cd8b4ed063870a01a5cd021f6ec842d113f8b5f4ff1cead4e24
z759dfc5cff40796a2d7a99aba49b5dfc35a794d8b789fc5a52b2060a30a25f3b2fd7e0e4d71629
z51cfee9af40a8cd8fff9b5cb7da984565718085523628599b4b8deaa4bb51016db132b6b023d16
ze4dbb325c417f9250fec69ec9029a809069dd70b21f6fb65a9bb95d4433b71b3c8b08f5a04286b
z3f8bd90f2eb3c59f59fddb7ae2f10d42e14a7b482ad06955d056a4470bb431d23115bfd06e8600
z56cfaecca5001c72550b16140015edd029430fc7fe325e97ca3bb59f126fc32c1898ce8d793f75
zc53b24547cfb7067cb6c4b7d0b33461ac647b44e2241bfd70cb20a185ab1cb7677ba5f6fb43f1f
zb8915d7172c0ef327733548e29a28ff2e4decc1436e1306b605587b1dac799492b19a28c950aaf
z0c403827f9055b2982ae961b33301a5e2e11f89325dc970dd3df55d571d80b0f3c4b085cece257
zcdd77b53da7ba7e826020690b9811b6b9c08ebba647b2a6d922d82269f3286d98a7bdc6af4c6ec
z47e33e10e03362a439cf41ac14996de8f8d3281c13e30ee62d8e11dd69f0f98a369e5fa159cbe5
zb5c39db2c670edc67e66dc8c1dff79bb530e23205143398c0210a8a08c530a6893b336b698f7b5
zf9dbe5734b24853c65cb7ab34db992fe77e01d5845f5d45d298d8ba2d57abd625bb5d86c553061
z672c58c8526e6a0011edeb27f4b48ac0c5ca668a26810481a9ac15f5241ba9d86a6feb19945f30
zab4d781f74cb52c8c1c2c6eac202121f0bd6830662cb4df7752f763d3850c169e3a32099191b5e
zed9cd9806d7c52fe7c47850fa3d33da3d9bd5417eb717a28b39b131064e2d984a5f36b8c85d619
za18439cb687867d1ff6269411d6589d0db6e0692d1f4f1fb8bb9b22a273d3a5628bf6d8103179a
z0d412f23c6f69c7b68b0c80e1cc3173b1d5c1aec530993ef900a63b09f09273db75ab9352d35ee
z55a76ec061715072de4b846b583c26ccf47d5a1f94d2b2a47b7d669991a16e5a5148a2f4d25e6a
z71562a4cebd306b51933a4662eedaf0f5a3bd9cc8df61c353b6d758ff6b7e4529a4f954d9579e7
zc907ee68a3dd80f111a3acd1cbfc548dc0bc2353b4bacfb0bf85a4b934fab4fc2dda5648e2a63c
zb436c09c9f3c733f0c848b020a5c93f959b40b35f7f6fa806aedd5b0808ebcb04eb2b78c74eef4
zf340f2f24ceb314e97595cb6458c4ade14e2948810068170d68acc30f21d4b4c0c39bc714be728
z9bd48aa905017730173ab71e3df726d8c3a8e03b555c74a6303b9d33149977c9ed828f033f2633
z06efb19f75ad9ca6eb89c79d0098395557c588230ce5798e1656bc04b9e82578c336192960e70c
z478d2198abe081d9933195ee4af2802a8446df69b3450b7341adf2253d88a56bd451280d6ac02e
zdc8088bfb1504bbc705b7163325b91d5daa4c20bd56d8aaa43cbcec5a6c31f425798e24fa5a401
za52395bfe0b2b1fc7fecd0d8373f2ea22004e328354548d09befb59c5796313bd6fc9b961465ac
z5a7a2de88ca9efe807a89bedf7a5b31f5ad223838492097650383c1df43aec72512628623e9609
z4ef97074eeb1f9b64030c763407d9d4c6ad14869fcc0c9094a130d54c4983d1591041f14a76fda
z6ba122dd7466ff1e272e8c921d0317f27fff361675c16a2d19829b05f858606f5cbe22c846db91
z2691699370ecdbf5befce672c55b01bd6f6259d9507ea5356bb23ef342c49212d1e6f98afbd360
z473806b5708f197eeb3fbe75738c00d558147ce2ace8eb0d1de813b93ecb1c091baf298244609e
z88a1f5e2f3d7b0b297032807ccf74e99c1ff44dbff4e87b6e8c734246be3c64865e7b638a1034c
z97328dea1373a3072c140c7ac037b633e280b418f28adcaed20d5bd5ebf7e49e21a79fe74f606e
zce90afcd0c1c01582fc9d2a2300a27572dab6650e697fd41df3ed9fdde70ba7923a9e4596592e7
zd573572dd2a6e9ce4da0775e86dbaa97e01991640cd4d1b76d3826348a0027af0b33f632c52497
z9575f1079784b253837a55f3bfb691939404c0629d5d1117c9b26708f81e68def88ae98ba45683
ze63b0e95479c3bad58103082382960291c67a5327b07fcc491e444864c0ea936b69f7206ec9850
z878f8aaa4b6903a5a9d93aa8bb22e7bdbab45c726ffa88221bff9f930f48409d7c6ee89f123e76
zb5ea048e6c12abf1a63b700f20b2e902a85f686f087adaeccab4d77785f97de8c21cc0e09a228d
ze7379ba2cebfdb989b9f61d0e0be6aaa12d8a681adfb0766b3f69754275ad9ea2d45e3183cda86
zb3e1a6e76587ecf3205516f32bada698384463b8273f0678ee99acba10f23f8ca35a39148aa0df
zb79ee79fc615c5126b8df7c678195f2f96b25f5e52f7fe774ea49b03836ed94c12164ab92f95f7
zd0ed0964ceee456c7b386d49d10ab6c879a3d09d24d8d403bf56e5bac8a1130dd1c08e3fa680e6
z6f4e252a9ab76ae9a936b3fcad9de22ce094cf7704412f5c3684077f170e60de040435133c3b6d
z9568533184adf47e1dcf648d8fa71d2264e3e3be876681fdef63bfb3ecd1b2636c2e85cac5202b
zd810cc2ac1e0dbd94a1a290567b56380e1111bbe2e231f67083368565144483d25382ef113cafb
z81a87de81593d1557dcc856f74ced74e51ef8c3defd86a17359aeb4099ecffe50161a1be14a5b2
z9bce602d699cb5b0367c74a4d35268d3afc9984014a760221e2407fd173e626c69167b84dfb168
ze63f57b47f4dde1a73dac2b91535364937e38ae07b90898157c60c342002be42e7ef4da9c317d5
zea42c551105033d6f0fb8125cdc31c0191f42f242acfa856c6dfb94b16100702ebc3efc96ee640
z5705a5d63271c24c3b2126ea285b520df4c6adf52e9063f64a6cdf859c940b5ae123d18279650f
zcd65a9644f890a9782f07b6da8611b1938b2dd6667f68657fe7e9925f5365e5481c02656832794
z36a176f459da32c70610e994d82a44fbeb2efef09d2d57783b59f7d15d88f51bb7b3396bf6133b
zf7bdab0048102278d8e90b0d02a5291c5693ccb156251b40a0ebc57f0cc6927a3742648d2b861a
z0dbfad957d04dae39cf30b04339303c98f95d70478b65cc3b12f511788a0c1ac6309e77d149b55
zb72b1e7e0272b4d2951cd9649f8d0914f3a4fc53d1fd47f0bd0d3b88214548323c28be2ef80595
zfae4cb91e33c509f26fbdee4c3873378fea4a65cd82f45ae8474af8e08783b844b77fdcf769776
z0b27a738639a6c49d31f2ff96451d123f08fa2582f17c1dec3f85676248741d87af1e2af5c521f
z3933901518305b5ff269fab7c9b097c07d54f465fc8396a01cac4041fec42510c6ea87976a3076
z85927e68a0af8f1d24448d2fbe72ff239c76eb3cee1881a94632444a38b75c2c444fa503e4a023
z0fb026595f81e9be5d939f1d27da88fea8d2cd7165c79a948c9cb6c9ca62dc23ef23ead001be76
zf523024664765465b1b42afc18abd30f13c9db7d1d59a62554ff4f1071177cb8d2b8c4ca33521c
zd4defbacf152df8000cfd478e00116b5c22d1fdf8bb8fac95c316bd593081bfea085500c011dd5
z78ea03e263ac7b3624a8854a055d414fc9b82a9f84e9fb2c7993ef6b59aa8c81a53cab088d0c73
za413d13790784695787f7032092f7e756f661b9be3d8aa3082bc21016a67c8a4e6f9a385d9063c
z649db646d74fdf92f61f3b1462e6861b1250a49ab72d386ac575f68c6c439e9029f964aba1cd25
zb28e8f234361ccb9913a5066a66e10b085255c4104dee41f3a4ea0a4455602404af52511cae319
z923390785efabcb5d0aa1044045a2545becd788de445ca7325e8b92f25a2cccec752a90f829318
z2acd0deb435fb0f81553bcb591e396d0d2213a2b00915e902ebc9663430a45e09352988998d683
zc524a0cc780a7fdbdc082c9b3d23cca6645d899d961d5c67f970e712908e2ee12bbe854031694c
ze59635cd93d25193de5926535334ea944deaae532099bb0875a31dd8174bfb8589803ff9c5f672
zb3fa140cc2c4c536c2b6b5bd1ecd534f65704088d46abd3e495bd975f590247a551e45dda49434
z9bc41d1ffa8bf8aa4065928adc0baf913f3bbb8a4b84347069394c19ed19d29961f2e4f903b3e6
ze3468cf5de1837b264a7cf6a69bb6adfcf1fa5008d53ea57b2528f0317e48d4491ae82e62af4c0
z838821daed7278d9da685875cd8d6e1b0c2ba0d0da02baca4dd258560400c6ce3cd6fecf80b6fc
zced48816f933d73389860e01325545bd2bc0e876400efff4825f81b42b642763c961dde0272197
za1e2365e955e35049c59b3bb79f79213ffe3cb52b842ffd1686868c54ad82960c77f5ead70ed96
z27199daaf2117c248553edc7fa877c66f13d8f555020492aa86b8a5767dbcf346b2e6e9e79860b
z01e4c57120b52842c7b173bb7894dde33b207d078f0536a393ca5ca748eba989d3eb7b9842bc90
za48be50720a083155ff63623a098dc3819db170bdca6613f60c5ba01f38f55e23c1ea3aa406f76
z2b7f08f7a240942f7cef3a72c47bb0307a3496aceed7f1f99b1d73f0db03f872dc0bb867127da2
zaa026304fe8f2611e7e6e2372f431154d222ca161d287a739ae3c449c434ded6e0b88a5652f134
z23881c24e09949fb35813c0476e2fc12a91def15c8bec32774100de7d4c69deafc53ac57f3a44e
zc15a7d75807cc18bb5d50e8110be4147d59449984702f89f15982886f129e4953863e121df5232
zdb9272f5a267f22db9167a237db7db87fa294e32046d68e0f4f489773a60bb694ad85c8dc6f77f
zee06a4c4674f5476334550471c2a15e0fc78ec11fec716903b1f78d922820d2d9266b5d9549916
zf37b6903f4c94a431563e67cabff3296a5f9d6415749198fe2b1beb91de8f57afe80070134822d
za15613eb8c9520fadfafb8ffad37a6a80bf2167ac006a6d5ef061fcebe83fd757d33ab41cb3f63
z4ad004295beee663b331715ff12eb523d8b182e963448abd29521be80e52569204b523c8e76b9e
z3c4a8489453ec2b1215fb08f2fb4c1389be9b6e3f8b2cc2083996a54da0ef2f75588a120877c06
zf29b591c0dd0d1619479a62136fbf5330e35a0510dc2d74e3c37d7ee8abbbf7604910665ba0501
z0d9a2264aad684fca049a08c58d7c3c7bb8324ef3c8701b605c9cdee2c5c419cdadf49fc359e0a
zca9b864007832d6a1c70062a9298b2fca82c6166ee31c24def9b9c8308c2b078f2c0119f56f4fc
z5c1d4f41f6019bb3c8ec0bebe65918137eaed56099ff4ef9a650d6c262544c5d75615b88c80524
zfc2549b7b16dd9f4cd2994d4cd742b1aa4023d8835ef814de7677ba1af0e273427caefc0a5c070
ze185547d33f61333a1447e7b417f52d5f0f42d2d94d34341ccb974f8a166ab3c9f4d7642fd340b
z6d2f54386d0ce69bc0ba57554d2cd4c66230ff266df25aae341d6a7a8179e2efae592ff1758731
z5576ef60914ae884269b86c6d263552526fd4eddcd03c8eff8353bd358ab31d82e4f978ae02ce1
zdb10bf7d70a7e6dfd3fdbc6dd417eab65278d3d542d218de371fe9df9ee6a94846cd7afc95aa62
z29bca3f07c8ee7931cd4f27fa00e9ef3430d58850207c141a6736b2e6510fedc51ad7dd89ec429
zbcdcf502368b7f58c7cf21586c71eed6858fdc8f03ee6deaeb1c84bc80fc590da53a5caa9d35ef
zafec9c4ddfcae9386fee5b8d1ea871be6981912f4f6e9bc4dfcc9f9dedab53fe88d0c891b7ef90
zc86906b70cb91b6e08ceb4c6b0191cc814e49de1772879726f59f1041905a5e9213ee01d7d3ea9
z5f4af0017abe942d634342296fe61c9c1f7edbc8acbf352c2df64b68928ebc44b5f607c66a4593
z77d96c7ebfc44948ab103db34cc44831262850cd8b55e92648644f988859d11c6e5d8bf6c7b7c1
za0c386d0e822b4cbb077aa13eb51bdc4b5f3c63786a49ce456172d072c03e1eee466dd131bc0aa
z431a54ffe47eadeb6afb0a0b3ebebb1b1739dfa1b480acc530392e2a2f1b26e0e46c7b63e69539
z994720f2b6d9fb42b8063e61500161e6a48e5b4c4529350b0f1331aec9b4baf86143b68a2a375d
z33d4120bda9e46e84eae0277d458d808343fa65079c8716d0017c1fd8e0ab24930db81b3307a9d
z334979c26dfe09c2f59f2a4559a1443d618171c068b590cf117d5ccda322739a1b7d143ab442bf
zca8be782b619ecfa92e43a7cde94b94824ff7ee6a675aad64d69eeaca46e2d36bd06a925bf7c18
z5b000757ef947560bb7f861b8d9a1c2a4482107dfd9764f6226983dfb374a0245c617b2c235121
zfc055ea5efafa1c976fdd25ed0122a10898a309332f73d304a647af5e7da5f4a50ec5ae87ee0f4
ze1578aa5bc5c5d17d7eeb02b19b02942279dc4a9bc7f8e55fd6f0dfdcdd9fd96e2e2112b58fb57
z9b7cc29cd41c50a8cb97d45903d0b5ebdb71f76cf718c1174e9344913141959c57f596f6770b39
z016fa55f894935ca750e0c919a9d6e01b2aa79ff7d205de9a180cabfb4245cce290220383c79df
z27b40304e63556d665332d104da674333ae1bb2f7f4c92aa171cab216387ac2c2c37a7f4dbf329
z5ef46aadfab3da1597db4eb86e364116977e451fd27adad2a14456ae8bbe7563cbac27d0e82114
z4347129b551bd3f3d1896b9fc22e297740c636221d08033f041e93ead144cf4cf2c6e2cb0af9b2
za3fc49ef5526a6258c54e0a7af6a29ada5327b3884e02bda45770c22b0a9fe412e65ed5d1a0c28
zdde91570919bab80ef2029222685997621746a29bfcc144424a35d66719ed3315c9bbd31c1f351
z7d1f87eade52073a210ee2552b7884838956fe01956c42c882ca7205e4f0c7c650df0277c10955
z277208e1f09bb34688af43dd78ad5220ed695072092702d430ee0d3b72d8e50a5f58b7d146e22c
zd61af0dfe2efe2651237bcfb61c6e6d82c5648723f5755148820e023b4ef874922a8ee2fdb9faa
zeb88a3aaaf7970d44fb2cf1ef8a8c2ee9c29c10bd709024e3c2b8e65b3bc5e1e681fb6c500677b
zd78c511a0f0660f0a9dc139095fded5f14d3aa789e20946e74e6d12b712f647d8e70c0d40d74ca
z5e2ade5fca8d87e7b8f63e972f2952f4055460edb97e12617affdf44613790c1e62e07fac2bdb1
z8213b5846ade0693bfbde310416cca3d848a1e2a53a0bc739fa4a58bd95d2579a7f87ab5302298
z47211adeb435e4630a399523596f115b075be69637bf0e47dedc5690f44d4494dfaa0d0378b5a8
z6932191eae31faae476c80cb3144c9b68e63ca82185ab1771a7e273294aa69437e121fb4ff30fa
ze775bee76d7eb184c1349593b6a0a26c89f1c3caab72fc035a46244ab1b669d388dc9f4748aa26
z8019b8e3facdc120b9885ee07582f1050a52f5dad422a6619d777621837c757ed4d5a32eeec50a
z681af1f989a4cd1ffbe68c99d72cf62cd6aca5c7c90b5c007f0828088d8164c01ef619ac72c4d5
z582cfc1185d63b2225780495aff456a9ad1cc72a6af04309186ddbfbd3a23550f59143e432c15d
z6fbf5f2fdf862e32f567d19f477ac3bae525660a3ed27c1b65a4211ba1a9688ea5f7c5f785e6ab
z532aeb7acad086860879a1099090ba559ddb4979743162db6f867df053b64efe7cdaf030b1ab88
z6c512fb761232e0c013c13d18109a1b02884340644a6a3b381c84fb6394644d3c96518649064f9
ze7864e2f9bac03e9618c174e5ea321c475e3e5938c98bbd405d88446880e223bb844057d6cfe6f
z8e8a65bf4b925fa5d3e8c2916fa1fb555da265cb0ad7d4029e88941c01af3ec81c1ebff2099913
z9c31d946304b4aa40955b43731a374da08aec64a9a0607b2329603386d7ea4d0677bf8e305ffcd
z3ed847af2330e0e4481fa9018d7d559387bab9ced545a57f1fb152c03a8e1412b0065d306bbe8b
z39c3ee063c63ee7597794f4d84f25d2fc2b3aca29a7feaf2d326708dbb0775931da06cfab377d9
zbc913aea6f527945f2804d3ab932217a333615a61cadee262d32d1c4a4af3b54bd60460195688f
z63b4c851b257036ac85ab77fffac03c7ad5a63cd597bb04d44af9a437dbcacde7cae6718d23306
zb93bcd4e9be9b304ba9c29b8cdfcc80edbb846624f3b707876079854aa62691ba4260660a409a8
zc3a695e67b815cb7f67790cc94c931a269cec064a972f61a06156767201302a51df1e638fa475f
za6cfa7d53203181c93edabd89b87a0faa45821c9b8b3526914a18991ef724a9e199416727f61ed
zd4968c6cc1ada3db1fca8121da91cf8d379337c9c4e0ccb8fa87743c289609f5c217d74d7420a6
za56cea6beff476fa7e0d8e4248a0c52e78212095fdd9206c390e6d7a26d519f6046fca41e37323
z5816d0fbd1dfb60b50d30c3ac295a35c15976d590192434893b08f4edae779e9b4e338ce996631
z2f97dd45f2402d76fee703129eeeda34ee9441951d73823eb9210327853bcd68d1725c1241238d
z97cc74b8788f502b8f60020757b9a49a77be07455dfacd273765b797486b8c4dfbc4a1a05f2b9f
z2626f47f571dc6c13c24ea436ea0708f90f4b791dfcc59c217de9418998648a270c2264a6cd19e
za17850824b51f5f260fba8ae605c108fb1728e9246013e1eefbc995c417c6d6a662c5db1f8ad75
z4bbb65dd5a01b06502243c4a52c3a53b717a43d0e4a1cb2a10f9175f110e5c90164ec2282ea13f
z4972fe44b38aa52f534dca40274c19ad7cf4aa7c5ea5d1ec4095457e34537126f9c7046d141e50
z78cbaedf3058b84eab925ad2398ee65f4f8474e1ca78a7f64ca8e21ec4e28a7d55efa94fa0322f
z5a074bda069fad825efb67e6288e78e2fe7b1b65823d173b87eb212ed9df5e9dfa10e8b74253aa
zd7958b6d6b0160c5b89b815624df2714f4387bfe719bd86133f990e2a5973384eca7ff8d1f6ccb
zf722e7d79fc7c230e49016a30ccfe6a78f20aa448873d33cf63c6b9f357cca70acbc86e7388be2
z9c0481d88d9e059ff49171aa56c83a6310cbf9244c2c62b2e6cfac2792bd1900ba59eddf78f8ab
zc8fb66b3aac2050d34077a6dc7454320e7cb63ac778256e0c1e853f7ec7df13a8799244f12e221
zee6e0a2df70b8f59e4a6d9e052d899765d91a577fd6cee7f181b2bdeea18d5b47cf244c0be9b42
z5ddd28f787c88b2c161ac80f12a7fa668277dbf5aee7c89623422c4513f1d6ff9d48335de0d6ae
zbdfa7498c9bcd8489904278efb35150223d99dd8902a2faf597a4a7fb9b716fc0a8f32cc45735d
ze1f8355f57269cdef7c2368ae3a9729428cf023fe8c8f90b54de0546fcc165c08ba15aa71d3c7a
z73eabebef2afd092d2d92207a98fe0ee006c13c0f5a4d37b2e7ad61842534be57905c87053f898
z5e80a7a86603b6226865ce567eaf8fb505dc10b670b35516756b1949360c6ebdf43ed87afe3cb0
zcd5b29e7dccf096a2c99006e4a46779334d19043ebc7a19093658835509e3f79366aac8c2f9587
z75ffb5af6b3c69ed283f01267084b59f8a78867dbab1874f7a2b702365020eb8076216f1791ca6
zaae086036df12d7935ed495ecd12a51253080a6af72822b627d0157a7cec25fcf29fbddc1f2d69
zad38168f22770211f184a58d0c2b1f58bd1ff30fc48848cd91b0f2cfb5b2caca3606ac3814fc4b
z80b38548390d650cb530d023b864fd61be95ce8abd4cb1fb2cc7324faae2348f96b2fec6fd2808
zee8832ed3931ac97e28aa0412573eb5a352c05d16dedae9748058b77e705b6f3eb244c301cfcb5
z6edd2905e260a9df1250d7acc658778bc3efc584349fe9313c6776a8f85c4ef31bad64149e3df9
z499fd1d8bddc3ec05e0bf0b9c80546a490cdfac64eb16fd3777681dc8984018e74b239325173ff
z0a871e945e5acaae15b202f1cddc37a95322d1f4b45fe0c25339dcfe0ed07a3641b597faeb9ec8
z003b3d663949de12f03b79778f63ebff78cee8b572b69fe78b5233bec0ccd0e22f8c9cb0ddac50
z378a2b0c393487f95a8fd942be2b4b5a60ee7b7f55439ec869e77cb691bad739dbd778cda0fb33
z0195109b24d197ad8c0682c455c562673721597ab3711b6e41c84ea7389ce7c9dd88d15852023f
zcb3b03db8fae5e71ae79e0ad18e87b8d028271d67cc0f18bfb154557e4a78a2cb0febb309ef06d
z6c3a974c5473b80c2deb35e67d1251fc9a673109e5a3a7478376384fad60111e62fddaf3674f74
zc14b39dbae0fe6798f76e9ddfeb9f41801670a9e89c1fa5572e01662564488284670f0db522f94
z78310b5d07cef6f9f07af4b027739708d265301d11d3a31af058699f25c491306abc2358d0d588
z437bc9fd1fb00506d32bdaad40fe02fd43ab443573b83c1e3d59ef022be9993581d810d30cb74f
z34cab3054b731eeed08e18e54e6e058a8a73095b8213245c1db0e728ca9588dce0fa8950045bee
za2eeb119ff0040e7297ee8b8dd603ce2583454e885e7cffc9b22053926278065ad69c092e5b96a
z1d1555fd13243e069e793a01c488e17330c34820487bb1d10569066668f4d2b30e6b8f1c1df5d6
zf4667d06aa982a770597ba3c7045afee9b1a90988872bff42cae64b92636f91dc0fe491f83c675
ze355a6cecfb964d0d4f59a698e94902933d74e470ec51253748107516e74ccf81605a167bc0eee
z495c49051f2b5caf84ab2ad018a1f7327c1a2ca5c814cc7ee6d22cabe907da1d8fe38ec871c5bd
z6d8bcf9777d3bc91f94c23cfe6538937cf1187d2962ef31430b19718d4ee0dba5c7c96005d74c2
z9c8fa5329b05a673b8dd0724f610d8e2d5bbac04e69fb62581d589331c0e7a8fb4ff2182614b61
z93310fe5e09f0dbb48d537c1cdb8a13b22824ad479a284928b33428248c6f5dd6cd2e6674c5d48
z51e5f1faae7035c319e0563114491173468d16819f21efe10f9444e577f9a51120a9b5037a451a
z518b5406bf8c611341abf251db62720d59d43a5e88dbb7d0e6e05d01c81d62d0ce0d9ae45b7870
z86cf4e543f126e2273b2f5c23bb37b0466d817455eeb8b8d5c5f00b5f171d831bb0c8296763dbf
zce065b1dd52cd56874f4c0cc7ed39b55e0fb8a6a0c7334f7ce3c6b4a9e8c67b060c89e32a043af
z117be691d9a1d19d0b1d41d3da501b004d9c48591385a307bc236d919318a5e2c6c6037c3359c0
z6c7dc40ec151459162722cb0dd94665808ff712bd0f5c9efc156596fa3ff402c69f2e467783a69
z1d543ee9834fbe62fd69579bf75a8a301d75f1aa2f886d006704542403ab3b8fe31ca2b06c33cb
z8a170c8d4b63cb3cfd62600a746b55ace81d9f773fa3986e789b9218c64e2fd372f8248d426d1f
zfe3cabdb5f666b3a4451b1e63a33416b972accd60d8483ec48eafbcc3533ab6b71aba5bf419e1c
z63cf083f279f3701cb2a6498dbd71fb8808c6828892bc9dfcdbeaa1db53891f408bc92712b2d6f
z57e61b7765ed6b4dace2c9cc8eb96f7cb621b1e5e3248cdb2c25566cc3e823164da6ad9e0f4406
z4a9f2cb3e26c14d43cd28b267528eec3bb9c970590ce6dace01d78eadcc2fe072045be43dbdb2f
z5d3d23c5bec6e650bd5723709325b89c13cdc80e38f5df607b78cdb308ba08b34842b362e72113
z8a63220fb7631ea121fd00965d1d8237439b80106a17f80ecc5a7d032820d4875fdff33c879f74
zfc09d4b65524de2005761fbabbd23029c6e9a3cf319cfaa39e035e1300b1ade13a61b17e48ea12
zec6e898ed44a6a0775f0c771d8e2eed8bcad8f42762021a8258815809a8f5c159612c61a795300
z820c8bd20d55e1c8892947ae5cf79ccfb411a02c5670c9b419d580008f903c90f4884a8c0a115a
z10e22200908fc0b25f165e54d8e3626564df48254758ac0a474d7b1e0640073ac859983e7849b1
zdddf5082da814eef80c137ded8808e1a03b3f439cc4a72e6a513f7dbf9f3b015de08012fd0e4e6
z84549077fe89920154843e9a566efa644e161bd4d6423ac057006194af314b193982b05f6040f7
z907dc11854343991c1d73470a94bfd79d1e562fa394618ae0b5c8e28075c42c140157a6601efd9
zef0ff43f3fa834929dca9010ec3c4642e58daf3e98bef611c210d957812e664ebabcc75b3f1425
z55007611a287cb3706abf9ef2d815afaa3505c94dc920ca2eb076d9147510ab82b449f5c05f36c
zcf578a51148ec917ed6baa0902b9c96f4265e5c9bc657bce81152530c224f04fe60fe934deba37
z6a9075af1e8e3dfac683c22df12d10c227e0a11a723a3fdeb27243ba955fb83a65737c34e3667b
z7807dcade8890d491565a006cc06f21df75ccb398b41a65aa532409214f6b1fb8ba3700808c2e2
zf915b1d5519c850ce7471fe7379fa16ed71529e06e5c5f615569ba594e9596185d5f5985cd46a1
z944f35b738755cc73e856c3396fe1fbdee0f83c82fc9f9ee99431e70c4dbd64b16e34c8cd75b16
z26aa99c07ab60a64868d87f62aecc5d99fbd872c88ab51c80c0c55df3b5c5f19ac196b6d5dcdfd
zf5c4022c955aaf027c0363c4aa80c3e377f86781ffcf3177acec1f682dc7b5d7b618d2a7f9e150
z5f23005d65d4bb987a318fcb9cc8c3ac09fe7f2ff65576fc1e080bf5559963d93c5c84aa9aa3da
zd1d6f76b4972128e20a600ca522900b8f77cd147844634e908bfaa768f8249f53b26ab2b0fb786
zd0cbffc16402cd2461991a15b80307d6e3e3a430eedd9833cd94a2b60b692dc5c3bab48bb02c6f
zfa09251d36ea0a7bbaf497a53634a0108c7a301013200b0b2a6efe6a6c983dc1fb2f793a944c51
z29e10606ab3dcfcf5470512a61d90e6337c5a5223702973b7495baf6cdcee289b475b390a7773f
z28e30e2e5f6c6faf365c200908babd067410124b621ed5ab164c61d4363bbc8f4f757d7ae5ac53
ze155208c3b389086395f20d84c26fbf393a536db7773031ef560b117843157ac990e226743010c
z3a19c197ca0d576075f8b5ac03eaac7b41a8d8bf881f811ad81dd25877c3833592296c37a05525
zb15526cd3544edd79cacdda1c4cbd788051e3c53351fab99044fbd43362eff9e8905d944ee4734
za38bf2a8fbfdd1b3913a7dec02f4c3fd524381d3d56f3f915a172524d718fe27813ae615a9e678
zbbb5b40eb54e3dc48449ca139f156204b4c0738f55a7aa4bc26151e3b603580944bc4c878cfddd
z4412ad064aa4df64f03ae406455e105a22d336da56998b9430aae1d0401c83e23067a220057076
za7c795e13a6d095d3b45e21b7faf5e83b7b2cca245bdb46174724f1f0cd5b159f1e34cfda302fa
z4a9f119404886773a3cac414721b02605fbda615378e14eed7ea6a7d6f14c67137ce71fbd7eaff
za7c111161fa6f64a17655ce404acb213dd373fafddcc30958d51da21f44fec367ad7dc7e3db0c1
zf4b4ebc7cb7b016f7f80fe34c7cac20a5ace6f233a23304bd5a5b2ad67c9a1a9a5a9548b77d085
z0cd70f14e0208c291657eee0c6242f6416325af467f208369c8992f5ff87238ac17b555ae35be4
z13cd7318d32b396f62bf2532fa7cac03a5592d78c54710d9e5760c4475cc15126a7d75f619a21d
ze89ca70a2c18c04ed8e23ba10c95285f63bb20159695281023fc4413acb8f9164840aac4725bd0
z2f4b4f7708c6eb12e478f42f038f4943924231174f3af48899e0f03ab9a6d02d1de917345c6aee
z38d5a44dd505f16f16de7763a5ad19eb6d09abce524d1b9abc7d2cef8db7197951b6d8c645e0cd
z91c4fe8bcd79ce5101e54e614c6941d0606e41ae3d72a67e26639608f7da9e015436e88d9e4bde
z801c11376e22fc1806fc344cade7664945f8392187c5e4fdc9f37429c60ab8b0fdd453ba2bf4b6
z266528116f8852ac33fc3c770d9563bcf961d1cfec274dd020124d1d7ea9dd1610a16db4394cd7
z55bd4345178a00f96d657e30d373dbae85a845bad9f14c824670e2eb1a534b73f13a2c1b3ce6a9
z26a25d1bffdf5eb9555e94da4a1b030537728055197d8d50c56c9f84403de22f02128e11c228cc
zcca2a186f906121093177402c000423410f497490b5113484521709ac6b19febb43dee26732cdf
z7324e371d66b697088518108621926605e57fa3d18f08d9b42e65c5961e2740b001bd845d6727e
z56fdb5f78535ceb3e1aa087b34f11f14a534b802419e149e333f6146b690ffbe48a3b3c814086d
zd867ac4594088f2075a9bb10fe45f7fac5ef1e6409c5754c69a40ce800410fe8b8f5ea1a3dd203
z5c371590f73e09b387b09b02906b86e54afad9f84c87f96edaf627dc868076f255aa46a0ea833e
z3b6e9411172f39629fae484f5d48c0a189cf91329d9682867ea21e0a9f20758907096e07ac86e8
z0c78ff7e4c979e22060a6042883854aab93a3a0ddb381b2e01529e22c07b6f0ac753ecf83082b1
z9d8f8484d901034d516792969dd3a3597b9d9a9924b8d3a37efb2a71e4201be5f838fdc1c326d4
zf24ee93c94eacac884dc6f00aeab1dd2be8b303e6d54494957c969cfb63b387f41a6f0cb6b2554
z0176ceecd929588273251931efa24d4e887b2792ef4091a2369b97e78acd3738971a160ed1ae91
z5ccb7037540bfda9388c088d4bbc01ec88d0508812def92e46678c24f2671f661a787ee269ff67
ze181069555f53db0cc405c25a72b68422fc127680d486c8c1857792a71346a9470824203bd816d
z179ac38a77dd2584c9579ba4b10070630cf597b74ef97a8108d9bba0417c5707e6446d55082fed
ze730875a1648d22dc70e34909dced5ab658f63eee7d62a0aa7a33c9521628f5b6f08b40c497a3b
zb323262ff66d3af638a27ca7e0cf854f00752270d553f8e95dcabe22d6390f730bfdff4286697c
z782b6b03332aaa1f98774931e021c8c7ef297d02c2ce5c50db84af4a83db8646de5272fee5de99
zf816ba1cc5e283504d46771f22a6af8915437dd2d1215b6761f886257627d8f98b5c11cb17036f
z7cfa9f14624582c44b994e993bb774725b9cb6a8ea5ef86e954bb5766bdedf93172fbdcd95c6c4
zaa98bcea215fa926ba7f677cfef2f22e52208e2b327bac81831ffe59462afad5b11f5c93ae10c3
z52f0b2aaa3e890d66bee3db5103e7e74e08933bb0363b24503df46b983d3518790019ef20842de
z9cb599683757423a9cafbe9150915feb4401191290289b0704f8055b207ff4e039228aa2980bb0
z067c369486dae5137393d9603b52d1a23782ba47763e2f99f413904a751e79925aad3ecb656148
z1cf6853353c95ef758e63a048f988fc4ea0c1e3ea2da0431e2b300d0d91a2b4901ff65ceaad8d6
z7b421177b1aad489cda77a1d9d0f017093e0231cac74a05e29362d2d455de877b0082ac3c4e5b7
z1ee86bfa77143e576ace18bcbb44827fec738fdc07980d26920ba042e8f70ebe3ec8c86dd01d93
zaf40075d8b69383feaee7ff1623025de613ac61915b35364934a4bbb3424839a61671e81cbd4c1
zde177520e8b581099188b6094120a1ff6f17613fa8d01053508f3ace74c3b9307cc4481e3624b7
z7d2b3bbf647f7f2f5628a8372160d03ca1d6dbd4cbf638ee59db60e4d588d80bf1fa987b4aa4d6
z9a89a207537296534a398ff396db5afa29bd2cad2ebc9bc2a40e32223bf168e9aa0f34747ed3ac
z4b97a22ff3986ccf75481751df7f434ed105554484fa94ab141fc8091fea9a8d749fcbc520bc69
z00f9b3af4907966df017f35cfafad657c305a3b39fd4961dd0791402c52cd51f8b2e5445a1d62f
z577d20b021a8b055753ace5f5dd7c434a7d47babe9eeaf2eeee2fa4646185b06fc5c3917a63f30
z435b1b46dc79043e59c0f50e7d019cc3488985afcdc2738515802f73f8f71e7004dc2100563e8b
zae528143e611f6b7461e42456f848f2287ae7b3362c3a3f91fcbfc2606b2ad4ff23d85d14d9fa1
z9f7465a45ebb37d089e876a4b45a2c37126efe7886a3600b4dd014b6abcb49a8bd491e419b07cc
za176c88a62c43f4927ce3103dd664a94999cd00ec2f41b67112ce100764bdd018dd6b7b4a656ae
z72f22a74bdc619b9a36256b8110214871f58d898e00927ba562ea286650ea81c968c592dd9655c
z882fb88974c7cd23eaec48be4422ccd5c45ed1b691d84804113c0365261d95c4ff6df1f2365193
z1300180090a31dc9f19001f12c55e87c7219814f61b539c3b051e5d96fee2abc1df886a523ddab
zed281c5e139e0f7899a04c615bdd9f136a6780ff3c8910a9d6301e366184e03eb7e9ddb23eec65
z51b1683d5fa5f7385bb144a71d94fbefdf07b5b25e367c0edfc81c880839092e53d20b5a3b645f
zafda34a3517d17834f64d12ecc3460f3f784f19fc0cb8dfbd0fcc6be2d04e8c6ac21e0ce126fac
zbd335a5eeb70acf03162a951a672efbc9e543f9bbe1016e12e2dcffa4504f86616dd1e3daa01f6
za5a0b14989916812b0899aae35df6555f4a8ce8b3003ac22a00a8d1c7e8060040df3fd06960b71
z3bd8b709664cc4fb45a54e46be32c1e064c6675600d28b909072a50a2b9da2dc2b7dd06f85b39c
z1993be668ae4b32685732c3bcca697a69081482a52cd7d4dbad658aa58a027bb75717047baa1d2
z3ecb40afb8a5e3b116d3082c7a1cafdc39bb012fcbac9b40056900aa05332d430e600248cbc524
z0e4a67ca3c17c58684ce47380e4a62eb443afe454590ed851008160e458996078a01fd13c84fd5
z68063e664895838c389053db9be6643fa498566a9d9d4461732b77e477b96c3711e09d684d4bb0
z9cbccdc9631166f6f90184290d142d704cb62c3b78e40baceeaa7299aaa7ef8e2361b00e9fbae8
z8261505fbed428341f6449d605eec66685cf45c934589ce6f598e9b24ec79d2edf92a4f87515f1
z98ed70b97910ba61cb49b3bfd5fdd6100364d83a8de1477213b23691f21d9d8affbe40967a154e
z03dd994a34fb5173b58f5b9fa7408eb8651aa0b03d805f715e223e2e6dfb8f6a717c9039f0342c
z78464a74201f1d639c000f42b5ff341c8f096785c2be12499285ab226a5e2222aa59443a62996e
z4c70b19cbd56eb038ce457e874987e266826e2187761d4656a3718e5b60bddbd3e016bcbbe53e0
z34bffdbc1046710a3c16958944b0fa16b76a5a747c315a5a9f8589f01a470af49f1e757c93fddd
zc928e3de4140d374117085886e88a511b7e62a1991fb9aaaa9c16090e11dfb76d1a27c78ca3528
zc647d56b52394323676dad39ef7a9123f6e278bc8bb2cdb187b6bd80a64b2fc3ea6315c096a764
z34d2bca42798729ee1448075a66d7ffcef75437b2ef844047c0f32e74dc7866457860bc2d054b5
z711f0b4a9afde14777d4d4876f494fd9cadb802116d6138590d07a798934be0ea59a0e6843c51f
zf307f4a2b27f8a86877780dbf730aa409251821f387190292104db0e5c71f28d47a09c0040b423
zcc16848e4f59bad98ba04b093c873498c7c5aef6e7418ccfa49c16eb8fb3ce18965cdcd63cebff
zb5f4b8a0415b2c161ceccd1bbb77e0b876ed9fb5a3fecc20ce9e96134082393e50916470184fce
z0b65c4a0d0e20dbfb22c1fceb134834272b85ca5b66e1b1373723ac4ceeaf1d91493fc6b8c8b34
zc704167db39fd087646dd7da4afacdc5533170a2b9cf997dc47a6ed582af01e9e1fca0408b09ba
z0c9abe20742a58c3250cf08ef5d45cd20d9031e0b33c6fff90c05a957d7abb67de19adf6bc1d13
z699e83d52f953e97003179e8b4a1c053b9423c7047ed982c95c34f83158165478fea941cdbffce
z160c8be8f3d3b090dd99bc843320691e7d30711623fa50a5d6f193cf7710c3a869ee5f4a59ad0d
z94aaec423f16de3e7cb6b8dbf015f86225be97a285d8ab4036e3bb64ff9d1305ebebfe88b78ad0
z25c4a00eae34f21294a28307c7f8df42ea53fbe69c9b3e856eb3dfb8cf9752a9b0571c0daa73ae
zf986c9744856f4e07a51606a359657df89ae825b47d856497d128e665b58263b6bc818f3d25b33
z98b3ceb5fb4a86c7698e78bc66a82ee3f2e1ed28b88a85747f5c5003c76b030cee14a3de94adc0
ze54b687ba1dad3a3021713501f936273816018c1ddba9925ef155c35d701fe427694dfe7477c0a
z219410b7c32d225d2bd244d8b9e61232f8d4f2e525ad9860f77fb59828aae825b0f3d905569373
zb1f8ef245b323e11b188b13ff3460d14974fbcacb205522be597726ecc37b1441b2c8b0ef7a3a9
z4c98835ebd2a72a5a5a2193c066f23b14e44ca6d07051e5edf0dd6cad24afcb58f91235f3ec58b
zbf65521473a1d6880962afab3f69511955913e147977d447a147b3cf8796d58defef469de3ef90
z7fe48a5e0e28eab014fd4b884967e3e9f050b6251fac1b63cb47b115861fa327893d6ca6bc62fe
z4e884b48baaa6c6e965421973f4a60d390cb39579a38de8638552c104f4ed5373056fc809eddec
zce34f7a19e87c890b5b30442a68bd1023beb4fa687240aaf51fad93d0a29bc1b9c21d39cea2e80
z69092f4a24649c427607a24812f0a604b0c5904ad1c41d9a5ef3e3241fdb15edaa24068eeaf3af
zb9a59da15c91b518bdc2a03c8846a3c7a705775cff7ee4802463c42f0c4ec55e56aba22309a08e
z28b1aa7219241f89fb73a2b0bf482caa4deec75ff363c63dead935bc191af097b2a8bca124008f
z1f736452b0c3a3bf2d068246eef722d452f9abfd35736b4c7c0272326afb6c9483d02a0f6c156e
z87eb189760f18de07409ee925ef33e9e3d8e416975b252882a10fc5652c9d6b2bc44a155ee10c7
z33e07b1adcce8a337b4b702b550864f1e3265875cbb35f3d0b5163e28202cb0dbb8d07bf9fdb07
z1f273c7ac7ef431cbe01fd71cdbc2a42a73d14d341a4bcce24fa9c0bf58cebcfe9fcc98303bb59
zcd6b893635ce689b1c20041781de6a65853be2f8cc89dc5413e0de3aaa70eef9c1e12213ac3dc3
ze1c637bed280b409f8b228c57e6465d75d0af30e48e77cf043ba7ef27b0f837d45c84575738015
zdca31afe21b230447cf31fbf0262dcd7037e6a71bac00cc656e01773f2ce41fad48b9056ec1139
z77ebc7ab2923381d850131223c6baaa60d02ba6983e124d42e8f24886b211317c840fc482cb8ee
za1fee963d8f9c1daa1933cd0b9031e8d74607cb69e424fafce02eb41a0e5399203430a82c9e50f
zf312286bcc662f1d247a78f2242ecd32f83adab8c18729f0d3a5987cc724b915da5a6e561e641b
z616d61318f1247e1084827e28207b8f639b8a8b875e648f0983d4e8ffa981973506b9ce080b071
z33d426b39048d30764e2d703511c163d94fc90cedef0ce7f9d4ac99068207cb67d646023339863
z1681cbc7c299979c445d08b473573ecba140278a15d54823ea6d809976c8c1c90027cba3be3efd
zef3550211d0581a0db04e97b350c79de8d6f6bfe0e72daa465cef99e1f14d99f15ce46c6bbdb0e
z3011e3b74b05ef591c3ac8ce054b06adecfc445d23e5fd71498a50818d6080b04707d4a37ff3bb
z75937548139625aba4a99886e87f9ecc39565de07e7370f3e7a4b7d752f987551905bdd5964e70
za64a55b0448204a2457c40bcd40d5f7f101d4b5fcd61fbe9a94d9773b0f084fd25d516056f2b98
z1780d8c50ba2390f231cb7002ea2d26062a2732e48801914e67e1da08fb27e27b174aaad634e0e
z811ef4c3bf662c597efaa28622a5d33b409c856cc19815943a144a84b63712401ca4db66a4a4f6
zac0758956b9145be66cb30fbed83a70d45b8db55bb40589489fe17472aa7822230d673a5921d73
z92cdf4cd6a2cc1c4881f38c7be0b390645b9b1a857a7d86a5f1655958a71b2c741416e26aec861
z6b6bf930d40ab9c3ec812fb5af26dc6c3fb4a6d4881a0bd7ecaa1264740cbdb8b263592e486752
z465a02b58229c84bada4be391e9fc34a3e512844b3d51dee2b9bb837c56ca6f824a21ee8258dfa
zd05f35954dd78e84115bbb481d37e63a8b358c870ec22ec2b50bb2669ef562b35a69bc6a902ba6
zb2bf9418aec0badf415d39e2bd8f0b3c5dae3c4432db88607e37c633575363c4d00d0a9b7c17f5
zdc79899172c818e9850c5bfd6695fa7af9d4590eae7d8441e30d1ef8a3905ac500bdf6d0cb9059
zc4c8fa00ea30e7a5287c655c3c16ce62307ef479ce359f7bdb63f54cd70f902aa74edd7a66bdab
z6d21f567d67fc2d127e36cfd2ccb5b8de89956174c5149829ba8e16fa6c5cdd3851eaf237c22ee
z3cb0b053573997c7d4175cafadd60f0c02adc42c5e97627391c825c8af8afd25953fdb88d930fb
z6d81b6937672f8e9862079c9090ee28f09b940cf70ebec97cc8baf20cd732e57b6a816f3fb856d
zbcea0e02e57ba1a1371d2f923fcb97dacc66358ef401a381c9246d229ffe73faeedca0fe528b09
zd6494ba3a85fbf6844c9657db6f9c272bdeee30f30e5c514af40d4b1e208b51fc03ff4ced269fa
z936867480002901dfcdee4a7082fd091fca1abafcb380968e2af77706ebab57f27da89c7f94962
za7292123d6f44be9b4b6c502a45a68cc9711138fa0f26ca8dc132e05b207da67eb9221cd1dca75
za48b327c1185b49f4d322d3f9ad8052e433c67f2097d95523fb20425cf10b70b69e5eff6cc4202
z70f1a74cf7f14b4483f119771ebc5a95db8ad5df02994d9432b358b3c661a36604f8531f615a23
zae7bd1f23ea6fec05518326fd071eff3a8fbca7ea756623ab7545ba4ab953d0e9e7bea7579e584
z58fda8c5c44f0b5789e2f4f499a0f648235eb47aeacdc3b33fdf390b7387539169c1b4aef49e02
zd56729bc821404065c8b8dade25ed0edda5477263b1292078479bf27a7bc9d2bd16fdf37e649f8
z8b2c2598b59f07d8dbe928cd8d87e2d668699fc94575c01c5accccc7a8dfda50dd50b2284d0140
z4f5923fb6d5cbccedfe68e83db2a090014b2941640fb54ae0d5e9cf309d930f344f8a8c2082014
z552d046390441faa2854a4a5aadc87bc15055d8e90fab22dabcd55ffde442269979451845846dd
z314f19cb4941ccdb6294bd6b9dde3df2dc6f0802a81e16ca14b22fc8c5ba3d0577de000b086b9a
zafc3e2746c58d0f5f6f123cc141ebee3fec45a3a53f36d3732b9cdb1edde8fb1bd219e610b89d6
z30a8a39833cbe85ab05a4556bf36fabb24b9746d14e4577ea4bbfffdd0a983311a19098a188986
zc1040e455a5b6ce9786574768cf6dcebcf0695ba6a91514254c2f8ad037751ab1dd773e4881979
z8557154b2895dcdc37201dc7ec833331514fb84a3b62637032f8daac7ca3c78e8182930a972336
z1195b22010cdb30d4e522c1b804af7220f75a4f6e478f30f9936ca8db7ff684c3bf7613fbd8cf0
z369d1c5396a541aca658ebba4d5be3ea08f99df0e4a687f236c183b792660374b5bd3c6773b85b
z6d022319e5d015b2e832032feca4df8a1256328ce7034b1f16911fceb21ebccea9682bed7a234f
z6f4747d8c739577d2db08ac67f54d2f577cd0a785e1c2ac8a288126e7a4a49a5e71b1fe5b30d12
zfa6f3605ce062de98c182570e2cbe581cf0476d199266d3f7ace31b65beb24c1947e68a7c669dc
z6b0a351f33ac67e50b184e6b06a6a6947640f0ffb77401940c0ba4ffc5b0ae05b04ccf8981625f
z79fdb239800e5ae5dd99d93b1e7723e2c9fc0f575a2481ad0b630bf39ebeb574831f166a092066
z4ca06078b32f30ad60e5041f197a6f4abbe9e265f5f60b42a41066e995734484c92886a6cf7afd
z6c5a994aebdaf72bf1b32aa597fc32892bbd031e13abff9418bc734df5fa9ef843c131235e8918
z88afb071b4b1eea5d68c1ae374fb3c12aaa6a31d4a667c1823e5ff4cdeae35380220d5e746b61b
zb6cde49966870a7ae84d373439ca0457c525a1aa44a087aa88b2b5e4e4177ac62aa830d54efbb5
ze2984dc5ef24ec4bf24456dc58b3aa05561154f5c247298fa947e192e585c62eade9fe66e667a5
zf13bcc4a7cb0beb934b942636fdbfa904d9dfbe4c2e103eafb365f1df8897d70bf9cd104e0356f
ze2478e9faaef9e0f86df96a5165e6182621a9b7f55a32321670ed07a5af4d8b375f31e1384c22b
zac521c03f345bab4f7911ebe7795c70edcdb911c33118ffd135ccd751cc9a5f550f2ba2ea32f6d
zcecfd8237a117b8714e08c2fcaa1a302761d73a32b480991f0c6160d1a8ff245885c74957e05ee
z2335f40f8ee2da5ac7f1be77c00bb1643acf9a606cf54a352b8d967c98db5b91dbfa21582ae36f
z8180815ca765cc959136261f43a5dc89ae5c5189340817fd4de320e92b6c20c87857c8320424f5
z87b1a12f244375ef6c33d35e15c6d723bc8f57871405ca7d5ccf19396677720b39c1e3870636d2
z322990c0dd779ea8ba10f0ed5995373218bf53e13e2b96967c3af3ab2681e68f37abb4c294b5c4
z141fe1fc5bd700c1e48270062d883c1efe17444e914d986eb14acaa5339cf112dd9e38c6291585
z439ef451c980b3e26922328b6d3801eee10f5da5d84ead5714a74aad01012c07dcd475dab5c5ed
zc55a06e6a11b922cc4b97544ab79d519168a47c6e1dfb432f7c374a4ad5d06e3e2e8f2539243d1
z384fff0078e11e1e4f220e6a7bba4632578f54649ed78b5d5dc1d0a021e43844a990018326968f
z6eca4c6df8c77e505cea07c38d2a41befcdf2445c9b41fd93693f9178f6b7aa03a461e32487003
z312ae4a57ffb7e66e5846ba99802b36948eb00820e18ceba585d03c0bc3121931ed3a7627f1977
ze1b30f40c6c687bace5cacf9a05a85f7d42c2bf6347595b2c7508b6fc31b95ed7b9152663834fa
zf322b304d41faefc0acb371bba4a4c2e7693183ba32b94e8078eaaf4cbc91fb64f24e67fc1ff64
z36a5be6fd106a852b931edfc93c8302334839c09fa8c88cd2e580c4d7fab6791e01e367e372d06
z1df08e3f53818210205539fb21900dec95eb3b904394c91e1c18ff81e52479dea828355473f080
z8ba3e06d51e7f5982ba6b21f07a616feb26f3e7acc2b886d1894373cad433aa2bee10b0c9d050b
z37e4858d5cd65ff86928d1aefd483236428ebd896e4918b25f9eba3b13d9c7c637a0be54f7903b
z6820f5a9a71a5bbb088d4b813b2c41d68365ad2aabbf7f3b3e3f66041b690140d1fb7586dc7913
z5df0f65bd591d3558e29beab788c7bccb76812b12eb2855d98076bf2d9e6ad4cf226b6b245148a
z2121e3e1ee528041a7a08ad6331c44917366cf7bc888c05f79805f24a8213beda2479c4796ef60
z13694096617ee4fd5594a9eb2bb86daebb7e2f91b58f932fe23e2744ee27cd109ee7d49bfeff6f
z325fc0ae44b9ec21e91987fee5e7aea1ffe7a3199f560e9c7550101b311b626d896c948e7e2d60
z0aa8bafaf91bd9e66157c1531f10712c03ae49cbeed6115e12093db53127f6013f7b027fa2072b
ze857c24d0f22b7d2a0899814ddcb4c72953efe256518b4ac98fbee01056b6712816d5d1da61501
z84680ce590800d50e94931212d6d5eb855ae69df5d1895d92c742918fa621b204bb06a2545bc6b
z81965787356d01ab404cf7c5d9bd5cc7ff59295995c01c69ab2d82951c295f70ceee755b5249bd
z586871d5d7bd3c712ac3388e4295ad778d7011e119f406362d7db793f8335f10af3e1fa4d30fdd
ze4790a74531e9ea25990295dfe55b98bde51dc6e27e5cff1abbfe4edff7019d4f94dc5f4aa716d
zf5f2b0162e5839e5574b5ec517f1e565660504016da19169293cd7dfd46b4602c9aea78a55faca
z7d9975e5c29275cd195971846dd990de4ee89661f90ff92d93979a1fb07897950f8c70746d2a04
z454dbb441393e1ad96231f9458441eb2168787e08e4326684e03ae7f0ac83c0340cb3f138f3cd6
zb1bca67929d173517fbbdb33a566ebdd087e66524449debd51a9e3c49e9331584039785b5bd03b
z1e16c344fe1063c2259c8138966bdb4dd3802fff632e16d4437ec20eef39bc6032e3a18d2824fd
z1ef8c2565cd6b457545cf714e2ab1c162c181a2498fe0d9500d2e5b4c6a058e7f3a64a7a64bccc
zb53d9c9d403c17874c18b12f89f1f12e34501dbc7453ba1f8dccaed91a1c224d6cffc3b6f54d5d
z0b38123575be9e431ab89d302272177ad2a1aa57d1832118977330dca138dab1b316a76cf5b6b0
z534bd47128943825daa565e14056836746c5bbc42f9258d00b657587c2c042c17602bca6b90269
z6ad4553a09efc61d54b01c6617c8f4d58ad97b0a5e2c043ed530a21bdfa92a51c1067d8642b361
z89a31e6749568b5251face3661166230f308836be665e0c8accfcc453b3e41f4c8abcf46ada994
z8458e468d11e1e236b375dd93c114d808126f6ee80855ea27e1bb53630e001d3dd16c8255193f7
z58dd679870292f5564405290d0533683f4f0bf298dcee585c7016fa5166820a49ea4c5f05f2551
z54029bf1681aea0567d71fc4db632bc6660b0419b105507ffcdbc8e0c7b7941b866a181f6b1625
z4fa77ef2f028f3e2b57841e8b19c9cf08d156d594c290d5e1c08be17464f5d9faa325ff0f51d46
z02dc918380b904805d97b6d377d6b46a3aeecc9e8e05dcb67d1ce0528a197d19ccc53666f5e130
z8e336aa00817f71b24d5c27d05a883b1a794aa1faeef83882544d753849fa56b98006e0c59b315
z28ccf1814b5d4b6a4661d5f599b5248419244718909b03e46d44bf599d5370fb2beaae98c73df4
z83e00398b0abaa124cc6f7cf071a5ed8699b504909e826b86cdbaa7847bb4814361e5506f4bdee
zb92ed7b02e13daa66c64ba7dc3dfa50f10747fb786f2859dd5195f8ac6038f0e2da516f6658f95
z581150054b1187d0dbb332682e9af4f9f8e92194a030ea0e0dee069885fcdd07504c404a7d8417
zbb3be69671e4d75ffc6cfc4885fcdc99155b564276cce10fc33aafb3dbb1345997427b0033d634
z0db858401ad690c4fe88e8db69a48144158fcea750c764442b5d0f72d419a62b1a4817918c3924
zd97d54d05ebe4fa1af677697e1e45b57adc5d04acbf09d6804e2ac8303caa8e792a005201af2f7
z74a497e3c95de8f65cadd59e6e2b23683c1ee4cc666e974538d9fbdc797aaaa31cb8fa8b05fbb2
z2171e3efb2ac6330f2e1adfc9477961a710525517f9eaf178bc6158d6a7e8ab5ff2a42596ab934
za59761dcb25792cc3a1a8c345145e744e6f62d9422c85ad8741fc8ad3ccf70078dd6e97e96be42
z6c137a4c029dfadc5df3d86b5a293fd5aa0d60494b2d8869fa6d4bf7504ee9094b9a7bb79876ff
zd7e68879f26d85df046967d41aa54e8fefd25ccc6914cc7ac863c78d7489ba9e093fa15627679f
z8f8bc4680074d5cfdf64157982788c324188a1d1a3fc68ff573e970dffb88fe6689694a72f35bd
z19437a38a7404b7ab78f51332cc46748d769ed5ceda2698f50786f9981f8d9681e2f1c3878538e
z4fefcfc4285f61c22a35ddcb7413291a77fc72e70ab5056df9933ffef1c656dd57996af79e0e9f
z7fb43301bed987a6df2166ad640202483fe6ec40e1a599bbaeb89c2c17334609ef68632fba90fc
z4db35b4f84ec6ca0d7a2fb483dd66e534c849de0594098039843a02d0640d206f6d77de526a1a5
z6b76f005efdaa209bc578f92c7569c10f7d928490e8e0ca3b70391a9c10d3e8e3b38dd3dbaf556
z1db4c29ae3f37aacfb677e6c3ac80263716a6d2e53edc6209bc778039d100d2f404a731a88f7a8
z0a6e852e23b17c3f0ef91a2a2d242a9fccc646942451791222f1c970e78f18d3703d075cfe561a
zd5c6023c06a92a506222980b22c541997457a08ca64bd62c3e2d9e3a896f81eba73b7ec5587baf
zae52a8899dfd66600bb99c3c8e7043aa9ba38958cd6845459711c0f5bf39c76d919a598e65b4ce
zfbb843c519553d889951dbb8564b98b85d4388c45a5df87403db6c5ad19b6988645f19f975722a
z9b2154d62ee9f2adf4790ad04618676afe80849abbdfe03c26a5c18eb47485ad3915a083b9837e
z65767ef99594b07606fff196aca92ba0dc96c6362ac8a3beb098ab97d2c2c49443286bb71a7b4a
z0de2d02b596ad3037ebdb98a5817a057368b03a0e7a1f7790e4b3bd6c233fb4da9deb2720253a5
z7ba58d511c19c37e225da9a9ea1a046aab84397eed565e2996b7b6d7ff1c9d31042efc7eba0e4c
zc3ba38433fddaa0721f8087a1b46a8e94ca1359842578b7408016b59b402b1d343ea665fbf17c3
z431f9e9b8ed3eb16e06b74a275f54f4e251a0d095f1149475db31980661f1f8c0e2ddcc5d216aa
zce889b55fed5fd4e1b211289495899bc7503c07b82df64646fb6208cc31c553501fb37bdab3f31
z6bfc2c251d9445ce2f7730cdfff5f27f7f0e332c706c1d2f0d647d35869dbe1cbc9cab08a94e59
z8d860f1654d275f606cd0ac0ad196a48d0804c0de7eac3e149aec935bcffbac7f928725b7d84b8
z63cec6b3c19e1f631270dec7b65fb3b61508f14e8944d152c6ea031194d55a54889a7e4e0a2b45
z928ffd64485cc0be2d79ace70ccdf876e7ca58c64cb39319d0d7e35a05c1a5936ee9afec856640
z9e2066c93418e8c835aee6abb30929b9b67d9854cf71c2c02b9a5e3c6d0fc9d8b1a9b5ed3885bd
z2453d25db424a2c3d51d08cc86f47f13a54cce07cf1a22347f505d6372591eab4685e1beed572e
zd85454a4bc9bb5c67b7c1d709c895978b81710233bcbaabf62587c8ad011007025333870557960
zc86c13fc8bd2f03cf2fb0d1a7181bc84a663a1abcce8afbb22a65c35344355da30010a02874457
z64c647b5bdc1d259b459f1669c12a3b274b5503ebc28ebfba7b769fe6474fb90445187d0c3308c
z33d340624bf7228b0bb6710e8492ba7ff7bfb6781821a2e15d279a17c09be1345c5097c530da1a
zf941060c6ca89ff1404513b892097783d4d53d8b11d9388d08d6297678af3b354f5a4c1a3eefda
z621c06b7ea7d70429ea4a2cc55885dc8026baee5a97076054c06cd34b5b5a5e5940a45c85118db
z04cbfa7ab7960feeb565ed158646fa17ecd9288a9353b41f086a1b19768eec568f04298709cea7
zc490b5942d882bd71d112c085dc4547d6f6d47cc490b96adeecad97a97471ce160de8eae4b4026
z649f18610753321f85b8707fbb63f8f83c078d133abb53517b6a57e145f6a394d0b797c4073d4a
zfd0e1d260f2173077b44acb6fac8b31d2c1d093ba225a37f91d6e9cffd74e1d70e7e3f75cc19ff
zd3a1ff68beec8a0fc6ba7b3063ef4a8a81fb2385eb8e3335c9a794cdf0165370f901d730442006
z5e369fccc60df98efca136942c8658f442e67dd479e166276373e3359ae0b62659ab8a36049614
z079d3991a88fdaac26fb089c6d8cc834ce26e1bb67748393669ea8e6a0efde0df6d727c16e96c4
zd3716d20f7444611f2bfeb0f731cf0335aeb647ac6ee715c617448cdf4e97a9407e53c3a960e29
z51beb666ab0a25de7dc8e14adb02dd8b7a196d79ce921ef8c9e8d1b9ae77e8e6529973c306d63a
z67800b04cb3011eb9e12edfb0d649f030da69bbbbaebc80bad5a57d6e13c04d95748e7c9ab94ca
z6f6cd9e58f1d0c06bde13ad03b9785df32a646ac38817c15c0f021d6485476e7d191b0403198e7
z4f8292899fcf0de74ce9bb982e989281e1dc9b07122e46d8fdeb51d09a766f4af5ebd44bf6fb4a
zf240ba7b26759acdd1a1f25e3b7749fe34518ef27d2927b0debd4ecb71be5b030163d7b63ec28e
z472db0990060a471a5104ab94cd9d918bae740d77b810052ce2c3bb9c19970b4acbdeb070cfc53
zea7e1add38df3a2a0311064b310973a98ac8796886e740d6c1c3ae7bb2ef1c395880ebd78f8a16
ze14d976ee29e6a92f38c86e211281db6e0ece4ed72256c29004bb8e4c8da81dc281422d10d4b0b
z3b534bfbd2ace7db1ce1a3b30d68d3163ed42798e1123bbdbc9d209ae28fb78516c9ac4a85b968
zb94cb682ac7156033e033e2406c2994d96b0ef57f44520c061c29ac9387741c15f9123f0eae6c4
z1a9837a4035a8171df90449b2bd5445eaf0c93aa7021a97e0a932f395526c2df2df35042ce773a
zd7af3cb9b42cf619bdaefbaaa56079b723e8bd2e585060afdef34f02cd8b96346c9eea25a2648e
z5c5c23744f16f852f9b8a6b3b81e9e64b0216f49ee554e3465b1e30e5c8d9927e9cdb69c33d603
ze1dc96518fd0cea4c491e254c15a9c0284eb662ed02b167b5758308afb0ec2141e2777a0c2711e
za55944e4d0e58c4ebcf4604151aeee4e225a53a100afd69ac2a7acba5007187d76d8f55e1c5467
z3811ecded00a74ba01904b8c6015039fcddf768e181fbdf6544d59d9a91dda1dec72ae369073fb
z42d9e709912e0a36f987a399097b929fb678187a434de39ffbc32cbd04a8aab17c414672aec474
z0d979c794227d3b0b91c624fa917140b00142ec8689429d58e10a642ae476d5878495c73d5d867
ze859962448093c2a0f5fe2f6b995ca5354bbfab08ac7dfe2c1ae8a6236b3d054a1075a6770240e
z5c7b8adca27214f5c9e5242641fc34aa8aa5912b4f12b9066b1eaf8a2278f65d8775e45a0f0320
z453822ab8e64fb1dc1b6ce455e681343e4864db6bea494de5de246f59534358e9408789e2c9356
z1a1d05871d9e2fe1b03aabd39d55bf212b1d2219bad20a9cb8031ea3eb7dcc1576c711f01b3ac3
z9062fe43aacdf380131b59bf8a0e4b80e831e05eede2cce1ffb9e08bccb04db2f0ce31742ea8e7
z9333a790771773d23bff1460c3cee58671fce85813ffa8e5726aefd6952582f61ffccda0c2d535
z2afbf2e4b1dfc6ccc9bf9fca1dc2147bdc73173fc8d61303b6f75a5cf4781b1fb3fafe45d3755a
z18e418c5f99b56f3470910f249a9ac83de32b82e7e43072060d7e895fa98c0e61b66786878461f
zc524a0d0a167152626251246a7490718bc83e08a0d2f4d601a490d9e0b010d02ab5db98cc1143c
z3ec0fe4bd01d89319bb2853bd89534448cc5a2ae9c90844b03ac86695221a0b485b301e4e1b1bd
z4277679bd3b968a3fa0f915432f3453503220821f8a868d293368c0d59a3765f92c9da1bb629b5
z30c52128de29f8a52ecc78b84a29a345cd53f2f2dc2de42e8c57cb02d76160397bd08818cc18a9
zacab5fed6232843354e037aa80f6c8923683eb07f5b081a31127c84a678b623d1ee2f8137eec19
zb1ffd3738ef5f5f886691f35c46dd83a0d71b1aa413053a4a10f4a53ee17cbd63fa2506bc2569a
zb6b22f1048b4274fd45701f0585523c76b307bb4e244a2562d4c393bd012af9e08df534828dd84
z77a955f0f619f88b749911b0e583b4877bb951db512e61426d02cbf7a9ac41fbc0f83c508469f9
z54aa19615ae30b6c9f546b71d814afc66069fb86dc8af227f7a2574ba2634f3c6dcc3b8d51ce6e
zae0ce397e96bb44503a480fcc358a6b7c589a1c73c7a0c8b393fbaa3302367982629fc9d46ddaf
z33554c36b757be94d99863f9246d569fa56576e19c8a0a36a498d23460acad827f6ecb69ffe789
z16bcfdf0f7dac7d2e090839e75fd43ad985dea4d96c439ed0978ae7128d4bc65cc7f7f941fc009
zc84f4e26d4b51626ca1d4ccd5af79ab78d3c2f1a2a1a0ff236d7d2b270090b6f6e6142d2f959e6
zae5a2bcbe7446ec91c069641c48afc9286c71a5468eb85cb804166920c101faa52f4700f848583
zeb63336411dee6a2eced52041bb57ab2db3c83d2e4702c6d720ef9c2c04735509ec255be0f5c22
zedf7a66254d17b11ce87aaaabca8f5a4b755a1a3b4c1f0245eb6e3450880fcc0a1cb8327091347
z44223ec0d313ae2b6db654bc52c3d4acdd9e76c1ebd1b214dccbc3e59582e84eb79bfa4b8e9f10
z6b56c433ebfd7b9ccf523c3044bfd3bacc97107501cfec1f0ee01f50e7eb479d67f00bfebcc1e4
zd16a1a567e30c8e767f2c29fa15fe41dcb44e0a6557a2cb9f6ef9ef13f60243502bb0867062131
z0ffe9d54d57de8d206afdae87ce1d373f34352bcb2ac3bc7de1679208818d222e9606f237d1ecd
z4854f6ba0ecb36cfa92e43335263df60e62a095a55cfebcc2df3fff73d9dc79ab9479a2a36e1b6
zbed0ef309e0e2099f5bbf6d8fafbc423c7b313d2a511ff927166b568c746b9ff21f1bdf24f10a5
zb730e6aaba238a0d545a9fc4d413042e7b7e48c0486fe8e95a608324c5c7969bae3941aa0f5168
z3231e2f4545c2043e51a31005bbbe692bec6102bd341d6bb767127bc1a9a6f0547ce041b8c4568
za579f15eb16933f4c555149124b5c43921de2fda067fe5b18aa1ffa2c1edb8de6bcd7d51e689b0
z54a74c5c8f5819b8672be7affe323cb850ec36666a4150e500e326825c6095f1829f227bd42714
z6d235e2022d1e56b91836594efb1457674c76080322de300aa30ae04a958d31a5e62d754923c04
zc3b3f7d8eedbb7dd1f32f8b447bba86afe0c80bcf886ac313175fadf1fe7a8d085624563435a4d
zc69e3efc0f5c9f527214d5b9717834154dfeade76dbf085448d1eaf50a49bd91db6cd17f81d74a
z452f2247cea2caad754b676e9335817fcc357590eb2fab6a625b009d6fb753edcc70c363dfe810
z546c33096957cee6512dfa09b605a3b342658291e5415b9fb755241d315f509ee8f07911ba1697
z2e3eb423916d4db9fbba7c0cef000915c7938bb55609a3e4d8b3e0248f1e6daa39f48f1348688a
zd9e039c9f7f6c040db3a92404713121d2d2c1b9f10b7addd60664d142cf3bcd420079ba43a7a05
z54c3523c766447f122a45b2e3098b0d010c45bf2e7125dbc5ff383987994d9494899ba2a8b7e60
z2600290918853bbc53e87519326804a6ea82298232a8eb8a92e0c4053032d7896e02d0fc459278
zb47d4ffd941d0a077cb099df24e0dfe77849e1f970510d8d955a4ace80914dc80f096d8ce94827
z425e66b89e643d091fb193918eb43f3cf9f74a6ad2ae3f23c3817e6a6fb93abb79cd8f5ed2dce9
zbee2d4084a2a05861716ece56b605a96183e88f81dacbe486dc7a181ca5692e6fdf301d3698c57
z2336a882de8224b9e9177a93f25736fbaa488e4cd5358133cc34add5400dc1bc1b2a22b502039f
ze6490fe99a4acbef80c51d44392177dba5f0fde724ef31d7c6f8812f39f48cc021ce018bdcbf62
z59b6df2937aed31da5154db762ea94142d98822137244d94c8e3c172b67d203ea4a332b43ad985
z8fbaffe979e02dca7f573fa94e0b6cdc0c195f9ffe880ed8eb668db2c74e281d6fcb4535d2b839
zb26d02e29a347510e96b404242582b208ad86543af7f9e988bd0a440e010c308d23d52a0b8b08e
z94825b279cc962fd08864548a3b1a905c00c72cc0ab810893e4ab27121ba9a641e8b9d1c9b3fd9
zb430e4e752291f12abf640909cb944ff786404ae04dfb300278b738399278757e273393e2af8f6
z59a7961399d1eaf41a15e276458faa68dbb3daba3f62f672b3c4d6e58ac492f0813ca5b2b43118
zdcd6708079ed2ace90a469b483fa4dd37f9cfde2130a4d3698244f68e988c879c558816bc9b4cd
zb6f4f1dc672606a55ee72d68d50b33b9829d747be7fefaa69ce2129d3ea9351330c1cb408ffac2
zf8f69bb03c232fe5277796032237bc3b1b2656262e8b8070e3a71bc0f9eca55fb20014266ea57b
z596c61b21110742418de02589394387e206501e251c2058397985553e72560efe1c1a18f8bfaa5
zfdfab170a9c2f603f34a40dd767db97503bf15610d4ba4c978c58909dded1b9392613ec1273eb8
z55659be4fdace48b7ddc1880b0f31e5eb5c08f52224e9d09d3e41920ebbc2f77670c85f12afd48
z5f4f55f66ce23947900e8e228edbba97ab16ae910af339d30ba6269aae13b5e0327b3cffda7514
z475b0db83deeccfd30aed04f861e792c0ed7d29d2035d8cf33bbf3a01b1dde24112a7cd140b457
zcf69e34c3f2766525413065d7876ce3706e079343f72bcc65f32ad22e76282bb27835717c48fab
z7bf4828620233dcbe4496ff39e80b42d24edb65794762d51f3d2bcf34f4aac466e9c4562584ebd
zf07ebf0bd6edc4c0c0db1bf603ce0c63f754aa61be8caa94f7de52f9df9f243fbd2850ced28931
zebb05be97bb96ad690413f163b854d1302a7e7516ff01579eaa8b28ab02b8d5eee1afafc150298
zabab05fafa1ab236d6fe24aed3e03d71f5b093fe56284223dbf60d028faedc8054d8e89fa76a9c
z590c5e41d2d385d7299f2f0f6dcac56b7799d00883083c94e1fd20ce2570193f140a13fdc3f2f3
zb2473f4e4fe53fb483eaa165b58fcab2108837d640fdaeff5916e4f69d8886343a66de868d0d15
z9e2b3a77b601bf96f50e12e99078a8aa822f4427fcb0812758b3c7973fac691f75912891f3247b
zeefdfef1afa6c711e7470f2fa2fa1a1e27766dcd5bc41c5008c9c552aef1ddcc6e8fe2c4bc3af7
zbf0ba8f6732a598f1f8d1592aace08cb571292009507970f5afdc92fa3a5166be5862da66ee845
zaa009aa2a984cc62672eb3aa4fd074bc21b228303cb53b811be40bcd132032dc95157b75fa5b7b
z8b312e8148762ccae92539a2f04d850ae3955e7232a77f9a9a4d3b21f687b4b32efd03dec36b8b
zfe10c8fc30054d025f24607b4fde948631a4a0632a76d9f30c08e05593eb0163efd0ca97a05cd9
z9b74296e9a63967fc7d0536d31e1249827a0cbcd0bb58b317397f2fac94ce94cc6be4cb265853e
zf1891c1cf84d4fbf4916ce067cd38ba43258d77cc85eb7f9bbf680707f2bd82f1eede481a5e77b
z164850d4a338d4215a4b1e6652bfbba83340615d9cebaaf32e6e838b5a76380a0b408df1364736
zee30498bae081f3504899cad39b370e046db16356c60300f1ec93a814e77b68af6fe0d8aacab82
zf253782ed06463c82d9dcc8a7c21cce6f50565d48f1c23d2c22d6cd87a39d78cedfeab82f629fd
zad802ef847bcb1753caacabb588cbd17f133c964d729fa73b87bf0d0c23b7fcecfb4060e72bad1
z5d2832d3c9a49b7abd3a920b32841172ce936e190c6d2159003e315b4fd4a27efe30117c8a90f5
z16c2c2225cc170abec443d79ff3e8d0d96481b9fa0d481865519b46789b0c742d8d6666ad037d4
z354d93964408c0d808343df316ed424fe9b2bc58360a6e83b7b4dc45ebba3c4bfa1679eb56aa37
zac2163ac0e99ae6cd1099e915b492471e9e5796f644b111cd913788d9aeddcd29fd0b47683fc9b
z84a475c4c881547efa146c4a05f47448d357cd6f77d2aaf68b7298a62de7e2c9690a99d3b39d58
zae1303b9a3d105858fc4670445e18e7d070d9b853437b2bf388959a3034c745574d071de8e34ef
z6e26751c4cfc0b76030e70ab0e4ef21a1f0e8a89c1976287f4b2dbb52fd9bed80d312b6d4f4e07
z1760a5e810da784a56984bbabfc9d531bc3eadffe80743c5aa61a476e2b60cac738c69f64f3154
z2a829cc9eb4661fc94375537a536bea6610253df9b16a0650cc965d4a32f6308dbbd2c80201bf4
z531830afdcaba420a3f7d2cf56ead14419f06878219835c4cc8091fee4f007b96fa4849650f7bc
z74190441239287c45a30e099015f77134730ac0e208ebc0b8238046b6b856a5712e17f4eb292e0
zbf8d7914f9dc73490ae130c6706f9a15643b27873a7c3f1b5290b82c118d5851412ff07b6af87b
z531c2c6cf1059822553d79fd4f7c2817517726d6fbb896aa173e6fdf9ec5698fbe8d45b6ad17f8
zc2319f7417b0c7fe2e08328e512886aaae40977ce938fe4ee44d8a3f6426d9cc73dfe87edaab9a
z0150728ff3de7caaa5bb6525c9f5ac1ea3f224eaac5a12ac1e0858d906d2d7cfdc524e71cb0bdb
z14f3b8123190d87417b6a701fb26453cac3baec7b3df8aa4a81968598a7f62b42c2a1a1f3ed29d
zc9be48f39d7cf240863bff6db9b6795d219a91f9462d70cb5f5d63c8466cb289edbda1205b8ea6
z481c9bfa5b2a78066dfea22f6a50cdae2d20f822fde74c2d19e5c464a5d21be06cb7b97de83d27
z3929df37934bc44825b74192e1a9d01614b5d297b40c90887c7b97ab982f9e483c9aa2be748d5d
z047a53a5665a229090aa89c766597319cf384e0c6b44937cd5511e45f49f83defdebfb4ad42ad9
z2adfc83e1885498e31a72642151a88ded82825f7988b2b79c90cd54e2ac90fb90b54765106b8d4
zf9cb516b54926e0e7250d8a6b6515a2af3451511ff0adbf62540d7048dcc85b204f4e10d0e772b
zcafadf0a6f3776393f24d17494b0b0a5c19251f00ffd6069c22789d0ea4ae3f70c780bb3631763
zfc57552f16dbf4020591967fc475e6783e8aba68c19186363d14cfe695a7d41394b7b7c124d5cc
z40f1aea34f754972de255d633f1f4d382c197c817b27331aac2bf2a8e1ba86698cf27e3d790209
z77edcc529032ff4abda40a7021376ba70bb4dba732776bd252b39ad04e417bea0509dff23177f3
zefdc61105ba50bb11b5070349a66011e1958295146890efc2967769260ac00eb383d0cc0f869de
z5dcd27a5888f619a24046aaeae1aa26cb6f6ced53228350a3b6e79f527c2f086d285c184b9e448
zc0f34990c545e92529318ccf9a5943325cdf529cdedbcc2eac46ff695edafa988af5214dc1aed9
z05400ad303ce69ad3184f40cb5d62dd27397d8118d48f5521171f79ac433593acb29e661f54f9d
ze69babe497df523ab4133fd404c45bf0d46ffb6ba5dec45547905fb85f3e96958f75654f4c8e4e
z473d533746ad6c433d2b26f665edebc0fdc55cd47ae4457354b875861046498abdac99cb303850
ze0b094a50f96c2f5e00dd06ad1e438f8c87df09c69cc72a512ac88bfda7bf2668e23830b8ca2c4
za729fda5fd28e72a9e0f40bd2e448a54f6b5bedd4f6d0a7371c95afc44fe1bc7c7612da2591032
zc341a57f8b59b653bf1c01dac8d14a42edd5bb15844c4b9598552f3342f69f5303b8ee84a648d3
z3d12abd3e0586f974c7e05a00c2671603dfc7f9a2a39ed7d50fc42987c0039d437cffc29b4d426
z8d8eb8ebe5f6d3506d0444c29fad1f1bcd2d4648081012b981c4ba03af5b21dd2371d59b951680
z2cc0f62fb31ba35b0bc4184d2cb65f4db20a3fb54010cd9f9321d612ee6d31361c3e8db496602e
z0d9af2541ca1a2e929694212a7dedd3a68b420f26e0ca6702365e9cebbe26edc27035687e8603a
z4d131cec4176c0cbba1efa4d27ce85c44b17ef848b068ed4dd43f7e90e32e403173c33b8162207
z83b131d2c94cb4edf8a0f2b8df5a60653ed8813b3f09b6b502c2449e6c4b005f5c41fe5028b6b4
z97cc93778fd38dd54fd16cb53e980cfb70e5005db3b8aaf7b2c5d0f67c0370ed2b5397a1cb39fd
z1e60dd4b2d991538270df619e77e969fa0ef8c850ed0521e32b05b9935264bc43eb7725279ba45
zbcb34343c4d7252be216b355b3f0941037d06196386248c4e2d0e2b0b277ee4bf3d8beef24497d
zfc88568322a534bd5efcb0e231a850d38fe2cef2c7cb902876d30f1b47935fba4f9cb2b45b9c7a
zc4964856d514f8838ba7e8a4ba6e0cd2d91607f1d65b708cc46dba56658aa2397aeb37bc888e33
z8903cfa27e5e2d4c7659b61561491eadc6f196c1e490ed4c4740fd9fa1fd32e01a67d21495a800
z9cca11073371597ead1ecb6114687d40de222e0f0991476a1545bb53ab1e082efe3f4b6cdf3630
z490e45e9d243ddca0c170ca3625699426d3ae864db105752d057f48b9ba6acdc0c585462803129
z7a52c2e4594824ca79b3c63fb1b3ba29656e6fcac679c89a7d42e201f0f83e3b517326a2ab2b99
z63028a15fe5c6718258ccbae2d2d24937665727aeab62f8e5958ad44730756f81b54820a86cecb
z839d879b033d214769220dbd40092336de13682e2c740b8f2a11f143f59a0676df94b050323da8
zea1f2e135fdf6c4cfb214cba49a3e866b5376352e01b6106198ebd3fc96d0e51811c67d6e59f78
zff701e5a9c37f65a6ba4b78697e796f7a4734be6921ddfa65625404998de17988a0c9736611983
za926aa8e128d9d9c2d24d1c040d0f9fe98559a089dc6cf75820955ca53a333b7e12fdc719d81e5
z670a784dcaff3a1b0db0cdfef6e1d6e196cf6f212328f510fa1d38d361e0c17c66e954d3cfe973
z611b292df53d5badb4cf97fd6c050687c2f373dffc919ff1bdbb95ef163294d1b34a57cdf9be18
z217c52f181e316173e2326ebc1c51b0ce0bc2ed8bef15eac30c206411d1124f09524c09ac67fe0
z6f9a70071dd3cf1f68c8fab98f4b95e36db23741b9668f207e02c242e756ed21b4ad54c0fdd283
z749e830623bb67c78f9fb076e251414dae737e6ba7dbf448744165ff2e59c6798c71310c46723e
z96e97b250226f41497206f4f7bdf8380a73d63af430ac7829f8d65609eced79512823305ba0a44
zd00db0396e72288736e0ae04492dc87b5a0aff22d94f89fe1ef6c6ddaf3f5a0513a6a7f2cb9233
zbc94555f900041455b51631e88af07596e096b9f9790e9663e76774f822e3018885d305d8565e5
z2c5e3f815faf1ca2ae0ca49613677dc309a8b376f74c34f67d20f9e0c943a34bdc37ccb1f22e2b
z538f076fcfb860ff9c4d2792822472fb37762a93a0d263160e6dafd0c53d2508ec6fba14dee22f
zd3b14071f78929aeccec8ca3ca130efb2eac05981f1d7620f567a68b1f3ddda664807f2c6d6c59
z8e7ad48e1458e9ee7d7bfc635a0c61d605e29752fea60584de34763b12c057c1f33a0534758a12
zff37fd7e8a50063206c181e89c4905fd098d7692ba98bdf731525cde457c4145423984adada6d6
z3ba6c0d4c9ab5b05295cf49c9aab2b02645924583ca4614a6c76591c569a11082787e0ef0b69c5
z3a4143534be32590cf21f6fba5f13ba09de1d89a64c28f8cca5b702c74c488c0c1f7c2e5f97678
z0d7e94ed27b6b5ae5a9c83d4fa1eb5ce656fe66b7d684c25e0cc8892dfada61bf03048f7eba993
zd22cb2b8b3a926d0e10dbeeeb800407ba2ddb86802900730f9173e716aa85e1ceb1e921b5cf5c7
zcc3c96bc17fecaff3c12eaa7156b693a7c559d953e3236503314bffb0b900e99f91433ff57f355
z8bb96aaf2dec6383b209a48eabf43ef6b937d9f159b69a4528a647ea4121cec148d1ecbd1a5d0f
z83ff32e915bd0a2250f16550783f0a4cfdec4fb22643465fa9a2ff09791c534b5ddb67b92f7530
z54b8a69b817b649d190cac167d4e430f3635afc2abc81bcaaf3caa64fdd74831400af1ff2fd454
zc4d66153c9079bff5ed2b870706df6c1a13328df872e0d0c0429b7910b428c8b5cd5220f317b0a
ze40c938a2faa1a30f4b9e6768ebf1f87729af5093a56f864c517b6f63ddc2c24f7f0297a285a76
z7e6e86cacafacbd9c4cd6278ec40932919040c4017f12c10869faac8e4340219bc577a5bb8103e
z5c737aa9ad6711c0252daafefb2b03217bd8e9fca9188fdc6a955b5d487c7f2915d0a3de618d9d
zfc1f86499bdf72e7c23b4411e37460ef821783347bf5bc227f4b63a57960aa5dec3374b90689f3
z03a73022373edfe2a54b2ecfe403808bdb517f8bf9a98ddf2874b007dbc4a4146f7dc96b657bd0
zde74a549ef3f724dd961aa08df7ab41a24fd1a064ab0749f6d00cc68fbb95cd1dd20a1cc500ab3
z46d6775d499ab122331ef11458561b684b31fec5123db644fad0e7a90b12a78f4bfe3913f1a603
z6ca6d2a50e29dbf24820fbf3c0fac7f983f590b3cca846d3290758b97e04b37d7900586f84128b
zc6918310e456078926867d78bf3f1262a193a1bb5514901919976b627a76665b8d5ff5ad86145d
zabe55b4504574363fead6a8efdb2f9844a6414baaa5628ea338ae5556dcab11234b063f8941071
z45c5bd609b333692f4bcddd9ba1735a2f676b14c1a3c628f86692bd696006c1d8815b18212ca87
z7520df47e4ace521d6a63d9092ef7cf1efbe85d7395e06c37f425fbb0610c08e653e4c6e70980f
z14ea612ce5e048e707e7d7f6fae8e7a4c0bdd2b93186d8563d3edda5dff5472f384763def94140
z57a9d128b11ae35edcb29c637f20f8d061fdd6670685aee13fa67ec4c43c2953831e955094c2f5
z5eb0779e2df7960fa60a23d8687e3504732b7fe4e8259ca25e1f0cf707d7385be1f17749b5fcbe
zac0929373023100bfa2ff13d4de04fc249653ed4c1b1896a2a05dc2d63c0b041f208ada10b5ebc
z6b0ba4842e91f725ba4328654a870417835c0fa9b9fa4bd0cf7a5296497026ab4a7c88251149ec
ze63b54c41cf9b0bf0954bcdd41d8cbc21378567cf7a9b963096d7e9d531c21a13ae8343073f1fb
z21d78f97181c01d25ca35b55a3a0ebb5e26174eb2751a4801238eac3155dfb5f5e38f1441d1b3d
zc7430366817644a265beaf0f568776d0929562b7a5331d7bd040baa1043bf9c596cfcf9888f297
z236d864ebae0202ce40cec9ed28a798d6bbac4003135f63515c819a5d7329a108d89b769101c87
z1091bca4ce81d40c36767eccf9ae654175616056352d1f25d4b37b9e276f61298aa25be3d6dddc
z15830ff6500cceb44d7d63ef48c8c2480124acfbb3f2dfc86e536fa5375560c353190004fe1923
zbd342f7b179da5d68ead2e2df99f33e0763723683b48aca66549c24e3151b42e94c7deb41c974d
zaf0e1cf7adcd6156fbacdebb8c104edae0050a578838734ed083679fb27722e024cebd45da1de7
z300b2fdfcb37dc0a781f6a6deb3c667aca2f27cdd778afe28b2b86775811a33c16752dc13b60bf
z7b20d2a8d0226f3ef6948ada615f04c192c7eb122712c581163a199715ac9f199201b4b1baab74
z1b425e90d95488394dfa27e87e3df783eed3737d1933689e8eb3e31f290ba9d25e6a4e198a2b0a
z07a410e725cce777b4839e076255db0f26aee95dcd02df29a3c16da2e110c6de90fec262eff3b1
zd72007c45ed3b4bb7910aa918fdc1de0e24382bcdaa872a8074baa2c68612e3bd60296ba412ec8
z63d3160058d7bfb2db10258d37757c6d3be15e34682eca88fd02421e60e4181ecc2322741cccef
zf806ec2dd2f97896ca0152aa3136fbd774762fa7fc977550af3da04e472419aaa140ff293fd75e
z2d385ce6c5201941e77ec6af803d9d8919b24509dc1c5c8ccc3ef5f6c109cbe502bd4038172a0c
ze014360443a733d08dcdb29704d80188bf7b50730282d62871aaa07dd9bc10503646aad3a2229f
ze0f7071e01b7701e00f4b3862bac5fbe8e5ae45fed5bce21c9541dd1179b0fdec99c5f3d91210c
zee6d4354c33ec304a0cd5b13e053822ab0008b5533686e2ae46aa84b8fb3255f58c6d25cc6a185
z5ac18ae78cea325404f54d07da64740556b167efedb50e19cc66ed30798ad1a011154e5f53799b
z91dabd15e9311d0180ec370b77a3318631b532feb95c1e97423fec93cf88140763840f3b2f499e
z9376b2ea322a6671f77d0af4d397ace2f1b51969144a13fd91b401b9076517929498200254df39
z13b7716d5aaf3d72125f8411f29db90182bd5b24a7e8ed3355f6b2cb5bffc1d77d02596e4e1d59
ze37a2719a829cfd8a38e282c924bef325c08364c2d2b2660bcab14bd3620fc500ac93bf041d1aa
zaf6e8590d75830f2c0700854025c93e81282c3e0c1e065f54933f4d3ebacd510d95bba0d8c9482
zd1823329da5f97792f6033523ca74f7b9bc0f6ff0f6842d89269125fddf13d23d7c2488e89d329
zb4ca559d7c8a7d0cc443352525c5d5d5f76a7f06bf5a515933d1c6b0fe1aee9e9144408ab005e7
zfbd0265a6eb8c393ea61f1093c2da552df924f738d22967d89de9e09b8ee73dfaaf6e4bc527e2c
za9a9effb62bc7eb4e8814322f5812ba185e6fce5197c3b714c1acbbc2635a26fc89292b796b41c
z26b9294a2b4aa88413082c65391ba121f6e04f8ec63b1cd3b44e50f8b6002bd67622447e08026a
zc3c10ca8f891fb5129c57bef9157c037b536bfd174cdb476ae91d51134c667ad9f36cbde1b4eb6
z76564bc5547f0da239799684d70587ed03358392114030322b128b956fe20b4b0ce6d4519f2ebd
z1a6e43afacbf3af7b2b00c1a37c07d07ecbbc1347a8e84fb14d807b71f69955219b66a6d0c8bb4
z2ea6eeff6536ce05272a7b303a3d1a4268e68bbe136b7697275aaeb54476dda4eaed8bcf8556e3
z31a7bb61cfc91b3f179617059e5159f163c55cf0db8f1cd367818f7b3b1676f94e12b31f734cae
z1249854c75138eb7b1b751756ad97eafe29177b99537a4ce5107e47c62683646236285350ea7a6
zee22d1c84f951ae4ab731c254660d263db5326e6417d17562797eeab0cd4b16a0b893d2a8257b0
zcc5b6a61bddecfb18bd3ef551fee86ebc4ea036801de1d77f45af90b746a953090264c224791f1
zdd1a58fdb9f6720268d74c9b2c71194037bc2bae09a96d98f0b6cdd1fa54b852a614fa3049dfe6
za10bafa9a8cd3a911f133fba544946c0833ab9932dfe3a802f1164f3f23842ceccf686959b3bcb
zcad9571b10f7e581d52b658acc2a9545724a0d0d0999231f7febe6013d3bd197512414d2c7819f
zb24d20c90cf0d4e7458ea7dc5a4ab451eade42ba14e755cd165548676906d51e2440f94b6add06
z9d3bb0748e84571bf161e6a5fc7d4bcdc3d38e7cf09f723bff20fedc7f963bebb3a16b91d2b9c6
z97f30bb61beaffc4b2ae290a1ff2f3541c8f2028cf785f68044267d2ea96b0cbc51c1ef46775cf
z024453c7765c351695291b791fa24dc47d237c104bcb1471a0dfab9d2440ddb9bbe7a15a2a6725
zc72b0f48ed2a91f29a80c528ee457fc665502ec33f1bc9bd6d702db819cedb1326921062321236
zb014d95dc077899a35f4f6b8be23b464cc4aff3ad472dfe0fe91e2fd64e242f7785e23583cf4ef
z5f0cd29385d5c50cd481f88fe5da8b787a6ec3e99f637b7e151cbc7a092455d887875ba93f6e85
zc84875945b3a5617a8a340c258fefe29765c53b162c50c6ad2a2b9992eb54ffe45a88bb664d6db
z582e109e3b93eb52da638a86846eb75079813c9528d5e9263bb0c0ccc1f3650a12cde4dca1026f
z73c3a8a76bf79ab89068bed4682f8aab0b5eccc4a18ed92fa85cf577cab0ab974170e9ebe5e998
z5549c6ac304b7ab6a257968bdb800321f4abcee103d505ed7617da23ddaa2752910d88e848f7b8
za94f182ae4cae7282ceaba16eeb1955c65a6ccb4ba09e13625b11728ffe5e599fe988cb44c5a6e
zd18a53dd00d804f87c80704e901aec1aecd7dddf33c21d4190780832e39d182013a28a20933c65
zb3b01e83ecfd4e2ded3a1217d223a4df342c189ea32eab1207485a8c2601925c192ad1d4e6e27e
z4348a7ee19379356f0410256f0f253ff41fc97630707bd6911778658f28b6952f4ba3ca0984f1f
z715a42e5da7721b2e33e08ace6156ca589f199587163db41107f7c66f7fb979b740e2eaab6daf3
z7af9d87d026dbfd7160d639209613b43329576aa071cfe641e18ff69e3c9b26e830625a92e12bc
z03943fd322ec2614c4c92462f354e1c08e5c05d8457e5cbebc51b64dc9012763db7ee1d5cb39c2
zd8b58403a872bc9d5f9c103f493d3e6301596f72520710f979f56c5b3cefd4ba1c24b30022a785
za4e9c4b4710b2afccfcafa1e13df540491c0c6423146fe039b5ce80e8840422cd12ea0303999d0
z8d84f3c18ea672b3db9b9f7c164278fd8fb4015bbd2cb3f1381bb6560141cd09c0175f7171f61b
zffb2671845f0801e9088d4b17ccd85d3f32c472b8deeafd7a310dbfe9eb2b62e87ef7e09fe59df
za511ad352ee6ddcbb2a5e7736d10438f5101a5a3a9a2f158300d9a4f4c14bb449d75792de525d8
zf44a7d048290435040f0a4459e418985d2fc72a2a641274a831c3d5420c7ddc2a4c132d8132827
z79e6ea892fa0ae2b41cb10f37090846192384dc7f3191d30c479a7f4a23706e3154540dab23ce4
z102a612949ec630817854de1e797a886342d8e62aea079f7db0fa207f13e2b95039476fc8ab09c
z58180c3c746d8fd2a3634926f50c7a92b9484e3619ae83e03815c9a22c49150716789b0f9e792e
z302ce18ccffcdd66f99bb46baa2cf7213e500f8d431f16f4d97a3f6e4b67e76f753daf40921a74
z44052d7d703679151c256705a7ad9152bd4d37c134003a5af083fa403cca47e5ad423366060ad1
z56f1e28ae40a2376fd70701cdd12c68f9877abafd3ea86afb3cad3aacd187b7801d57be7b77a87
za26ee6e0a8599f677b4dd9fa1de702016dba6aa1a00ab0b836ab1e2cede27d01015192a41dada3
zd5dc72dbc18bef6fb5bf6dc8f60b66f0cb32e41092427b7c117a6039c74c894c63bf6b21b1bb01
zaf0519573da8cfa87f8cc03a0bd526393dae7314564237b1e5b5dc33ac2297da650f89eae321d1
z633e41a6f15579a43314eb0bdfdb9e501814a13e507ffbc426a032b6ac4d5b0e91f4e4bdf3d486
z406465d97506080b3af1c94354bd4e40c47421b71d6613cd63130a8a5640fe89c23504b21b0169
z58c6d9d67a3dde5e3d503d0ec3e63595052ff3c2dd21f414cb952f870d760e1bc07da1838e756e
z1d374c1edd7e1bb26b7398cbe479ee5d071bb3ee5cd6d54a5da6eb3f7326e3f9903363a85ea3ab
zd333baf32a5c6b84749a1b1497eec3915b98b4b0de9e732ee1064b00d182f7e99b85e528f1effd
z2278e0afc7143784e1ac5106b24eb3d2aa515fcadc4d7e1696259f219deb78b87ef758cfd670b2
z6ef070105c5a654fa2f066140558d49d5d84d52eb42e1ef823df42af33e4e466898c127bf8eed8
z93e09562f4e78b960aa0c6086cc837498bf5d963d86a198a8490d7d3ed399405d8da485f8e5970
z37f6f7db40b587cd2570d09f3cebd7db97e47da037410cf0b83561cb827100a69f4c93068b34bf
z7170bae4906356fcbdb63184403ac884c0ca85c4dd4afe26250f4a206ec06828cdc536dc0f3722
z6ed238c57c0c3c75b1ce6cf95b933a6fe716ad379d5fc563421e75731605ee80b6475938ca9c0b
zba99232a26ba0e66b3850caa91d164375b8b780b32f91d63145a14cc612d9de1120bdd12f49ea0
z778a278ead5f92b08551f6ae8df211e4e2fa214a681bb221bf00bb415f19f201f70300a3bc3951
za008630261c3c5daf453bc5fee8994e3d58b3a88678bf39180319b7ab0d6f9b13d6a8e414d40cf
z0122903a06703187840b45718d186a00bd67babfcf0e514ab1c21e8e6f10e89ee06134ec3e9bd2
z422734a66ce19f4d7c0afc6030eeaff6bcc5793eb77687132569b99ba01be1d19b101d55862e3d
z88f21515bb0642d371a9f64b6750647e11eea8778322d7751dc8df9445e9d18305eb18dde61340
z4e5f8f6b97cf684f65d8b6b3cff266d20df8296e6bbe07bf207c09b9fa47280efe473e0067f219
zb26aa67e990d4ca4345251f1ea73b3d93f0f1fcd53bb46db2e5e94260c3afbd0c1c0f693049e68
z780bd21b69bd821f6e6245fdad0ba03bdd9f6ac7659d4cfe81d88bb7beaf7ac525192d5b786e77
z3e9d568608369ca8064951971dc8fb734973275b3788503e9dc2fbf7140d8d250ed5658fb8e180
z0abe864c42cbca13754f99d5cf5b98024c4842c301a03d0c2822938e9116fc7e7fe440ceff8d17
z13a3d964761303b8ebabfd24af0933133d16fdd839e40a964a9148418e36d6ff5c4ad8b1f2446e
z55c79044f1896a739ba709c6818b1d6d369b3b2b9bd2e7c13290f7f8f56d8a0bd2fa89b4037f09
z56f277ac5ea26a88c39e1f1527d9a36a052e2ff81bcf2380509cd6fec2a4ef7b5625b36c19d718
z1feb4a895facb197ab189b5bc25c3e0ffe10b841c7d653a17bd5427731f407e6d97e3381e982be
z42ce036ead63265bc88feaa9bf6a1757bf1da7b2c973ee5ca79ab6d3cfd4ddc50de96f49dec065
z7f922fdff96a3a0afcc17cb52ee6d95b4fb9d0b1467963919e47b83ce7ad7e83cbbef54ca72259
z05dd1279169dc19435922b849c7439eb5dbba1983d15d85e4074d0d86c930f45dfe6adf310f3ef
z81bed84cf36bc7c6df788b9f5ce965ebb024f62bef874fa6a82dcacee941e56fe1957651bb2618
zf966ef1b2a74dc76b01209b9652754cc854fd5602a20f0961de7dcb9ebefe437854b7c5b2e4154
zea55677363d54056da36c63dc0774c358cd9893a0c854c6054a7069f8d46449283cc734eec353f
zc0efc57b81580243726399d1dc706d61174151ba19164fdcb6ee635b7ef98d4c025090ebbf8c21
z5b63175d41d1c39ea7cc13731ac092f2630c28c5d16c0e97f612d1b7b6e6f6f2ac121fe8c0c288
z4ddb03939b00a64c2177cc50bf4a906f5050f01d9b40665791c344784f35770c624e2339405fd8
z8d1f4197359f0ee31ac8deaf49bdf2900a7d343a04b7ab48d6cfe6942e041d8005fe37f6a8eb38
ze5c219fd45290ee7f60f5fdc28d0cf6025fa139acc9de0281d13ccb5ee48be37b9e526727bfb48
ze29d89948850217db95a33f5f5278077cf567bc1e38981233ac661933e2e1144faa0d5d7b8061b
zc5edbba41a17515227d6e94f375a511f90b1d654791bb698297749d43514dd043cb9304e551021
z19b3752da133b2a4e2ea472a94491d8661fecb148e2a9693f6b22b7a307957ef5186f40e8f9777
z8b1396b8d130248661335149758ac09ea928bb4910d864fad7d8474018f0df7d20aa16f4017311
z123b290b1d1ed5740e19642d8893b3c32732802f63945452c7e38181ef965a7fc3582ac7346720
zc93897aa90680cf59c457dcaa102f1bbed65ed1726d7c5ebf117f933f13059a9b542c548a24482
zdbceb6318407701120cecfbeac7fb3043ee1b2c545af6f13c4bbe2f362c8f51ba754074717afd5
za2ab39afed6a53f20bc867a22f155c84ddfeb659546d2335c7a49ac67e347848b3e2fb1e381c9c
zc5bc8447bf1a180500137b5e586a02f705482087fbf85abcb14a6b6b0f28cce03f4d1e3d130e1c
za2a7c23f4826367f09012414d96be08df02a512d824d595650e210e0990a2cb310c89658ebfd4e
z88512d6272af2f3b9b25d1cf53ebe0347ba6aa3f9b1f458bfc70f584e97f274cef348546d29214
z4f0a0bdaa7ff0b82801dbec47ee1388e2b63e1744540a6c104f87d3f04751dd1ee3289eef9208d
z2512eb69ac0ffe3e10ad141581f56927010d2b79dafff70293c41d278be63f8994a6d9d613da69
zf1c4573c5b98ba4c18ee8828ce24bdb2501f550a470c1c281432eee1e68853c740e911ff564651
z02fde9c1db071a6696e8d94c0ee3640835a80c98492ff6a239af7af7e066f2667a1c37cd3282e5
z487edd0246f7d17fd285ec6a7eb0a61894854ec053386318377ebd643e5eb43fb7a22dd0efa533
zac0fdb9d20cac73a2167824557250281f32ff99b67565b5f06cad9aa87a5181efb7c73389bfeaf
zbf475e8b6e6a23f7c908ba2be9b1f03a7eabf31cd8301189e7f3970bdace39301e4b27ef310ba6
z169ca6e9705b8d0325b31e21dec3534590fb0d01812514a82cdacc8ec4a79a2deee9026325e013
z6b7aea67f75ab1a819bbc7e1bad91a4aacbca203a2fecce07c5ea8405d8169b2fc427d8792307b
z24144bd3a20b4522122648438a631da672129f435d644c3f8f9db6a4e0df486da663a06e42528b
z2346a7bc4817666a360e4878619bc6b81b57305c28246b4185ab5a41abe827266a903e6fbe8e51
zb92859818c22c02d5505ebc596fbc1fb79bcbd1c1b614fe57592dcf9949d30693bba8b030aa383
z02a760051232727f4ec2c2f4b91b57db16dde3fb49b58b34605ce0075723d3eb9c7686ac643912
z49d6fcd95173cbbf4e75343615a2c81428509d03ca5e5cd05f2fc00f76fd1aaa8c9a8e25c13823
zc01b6724a4f337cb2145c28d855daf77dac929c607dc1a09c3fd94838bf0d86d133a4f785c4ca8
zabac1dfa2c3ebb8368211272dfec4dff09914e03dec78cae49a907c97e0de6252daad3b22aa5f6
z5f627847c9906805bc3ab3f435e2cd8f75c4a484377ed21f0e0c153b7dc1cf51542360009a2fc8
z55a415b1b810b5e074275fac1f014b049c1865e4bee5d65baf0995c18b85a66d9dcb15f0e89107
za7492493c51d4153a8f0630de841b8441699e2dfc868c0973976064dfc0d33e174e2210e6ad015
z481a2944d573867fd647280da3bdf219f083fbee50218083b1ea29fe53d4993ffb0877f8e0d5c9
z70920bba140243b4ec3552e7a4302e5081698f62114e7c4384234201ec8012ad2d20af068bef8e
z00b6eeb4d8d6f63ac38e5c7470a433ffb6954cce19688c7b14c209c82a818b1504ff4bc7c43f52
z7ec06ce940b326338b2d662aa2ec16cb44eb62f7420cc1b79d56d2e39a5f0f1e8b8d75d3106728
z821e230267bcc531978cb78b3438670d7669dae61bb4098471318fb1d0b092a5bedb33b9a1e06a
zcb492e8c85df3afb502a2e83964f923030711b83146da60132e1718d3d84da2d033c77528eb0f3
z506b418856e52b06afd547a2e83bb2c7f666c1b865157c9c6899eaab1805434d0b67a09826181e
z5652ed28665cb7a1fd46a991b84e40bd360033482f1cb094cac70dd23047336aa945a120df0921
zf1da5b679cf277f09e36da64e77fa66983d778ea93ed3ef491863e29dd65b5a2a7ca4662ce124c
z0dc822516d483e44c1157c5047b1960da1f94c417abfbaeca852323b1cca3cb90373614cffe388
z6a28e9186668a1bbfce0a9376d93315f97a069fb76554913cd5ca7f258a926bccc708f9d80aed6
z02d0a4db9aa13dc30cd5b043e4a124a82374dd13ddc4678faef08b62f5d0ae3d1df00abcc0b5ad
z40a24dabc40ec810495b3394b71fb1fa951c4b3494f31a9f97b21b4ee44ade772eaf83a26baaa7
ze334e52b53ba0bd7f54dfacf872a55d9b664e010203d01e610e2143259801a7ac824ab7c1d298b
z3def8da8f9efece260eb43aeb808a2bdf1c43dcf4cbd00cf8bd9bdbfe7ac5fdfcc6ca653d9b389
zbc5b9c97c7bd7a06fa84f8b8ead56661ff4debd76a3727418fbbe2ba589dad33bb8fbd0b2e5676
z06f51f4ae4c9f025be9326f08e61fb40aaab91a5bdef37407e6f0308b994237f374ea96e19dfef
z748991ada6f378c8bad099c4ec7e05d5fd55f4004c6d1f02bedb960f77f786307dfe3d8ee4c20d
z1bc1c3f1f3b29b54c1a89fe86691cc43c7468bf68554bf62634e4747eadf508ae67649b5c35e83
zab02d251ba522c7fc8694a8b16c0a0aea1271421fb08158b471cfc8890054cb720e99918b90c37
z5bb6a8856c80dcdf6d289138558874f118d3d5dd8c8ec8ccea4e2fff56939fd19f9f225ef8be70
z1b5b4e139095074af70d5bee7843b93c3f4a5510ec43e75be33530bb3f497ee819a21c69ec1f0c
zf5b87eb304c590d2b0203270d5369e765e6ccd600ae6d2eae874f5f4b8112963936fcaaa093059
z80110a6f892b9593334268e19bbbb0935e34b55564fef060c26bd73e5dbec3be4a0664a72150dd
z699411561bfb0aee3d45b8ca3c240001218479ce33f62d707926428f7e283e6fef5f787d4f9b24
zfc1b5999728c80608f34be970122aef3395844a253baa840699465cc58c9b1ba9fd8649fa97a92
zd657070fc1d6de62f555245d4aec2694849f16ef6a134e07b32422176eb87ad3c36653f2bec1be
z3855c2bd0f9b1e9254a83e39275f88a72a0eb0bf56a096fc90f64c122fabc41cfab1795e3712ff
z71bf79c963752fee7a2ea12a767c44d7692a8ff2a4108edaceaafebe077a1d0f41733f5aee70f6
z20b337df763b3114a673b5126320c9222f72782007eb244fe1df749eddb42d3aa5512580ba9f2a
z92518da4f3c3786ddcb01c53a24e9c5c6e1297d7d9e93974290d4d3b240983330e211d5055e8a0
zd3e8e20c80789135f8f6c2b14c60d862a6b499836026bc8544f6628dc13357e5be5a23e59abdf6
z569f93b1743d279fbf1e0a86abed72f68491954836310440609732a7d3aca864f2ecb6b18680f9
zfd8280fff58b9c0f8ad89884a382c3bbf745dd6ff8b56c31370c037f0e354e2a465d52e9aac4f3
z321671d0284330406bdcde0a443cac837a0d0e492248adeb7af21ed6edce5955ed5a832f81f87a
zb37df37bc47df13801a62bcef400b5d74c8ad0eca1eff3677fca977a1959c7dd959ce92a5ce9c9
z32543daa59d1397d1f27abf94cd90fee8ed2b7a168d1953947f88a2b2ed22ae53b4fcfccd210c8
z89096e16cf92e70253fbc5bcb63eb44a2f9e859cf05eabde0ba684f254423bc7e44a748b9b3753
z342a086e2c681659150ed46fa1d8cbd9a5f0215ae26a5c69e2bde418b2254cb640c5630baca999
zaa92e98ad33b1868d9824b325c0427f2a8e0a1102aa1af7ac8fcaecaa1bc002de221934abca1d8
zc0eae549538206023fb719ad9d54cebecb1191ab1a949e54b407085380723efaeb3ad4e0dc77af
z335353aa097f82e05207bac970a1c703f84c39755e8bee177babd4462acf50190cec963ba5e4c5
z674d3a5c05614381791fba312df0925bec9b0279760d4cbab6d28b9f0595bebccbe882200b65ca
zdebd479de236ac3e5ef83a83019d260473a8d8652cab739b9b6c64d12df2bc790ae61a5492bf43
z1ed4fd11752877a3adb4079e14588f7b466f5c6788119ea14f2ec87fcb96c30c2d4c392ff22a0a
z7e43ef4069694a63d37220441a0081b98594eec7b875fca65f3849f9d74d055861a8d6381afa76
zffd81de23c047fbb76d1fccdb4d5f6255b899c788eba9341efff43d2c70fccfe927946d4b47587
zf98cf130531a06d88e6c8d32bc9217f5aef5fa0f916d32633456531d432a397b7fbb7bcfc0d255
z57e28aece8c5f7e6c672810ddf1870270cdc8ff06d13ed0fe2b4434f07a16c706be68a0a1a0259
zdc48de412c3b76412be33e201f3ed3bee6eafb4e20063ea58027ce9e6a8ee7d7e0b9b561f2dffd
z4cbe396a9cbc8ea107dfa8cf8c55d57d89b42b0e36fd1f4b9899fc329600b3c2618d7a08d6e384
z47fe712f5d3e6cbb1a286339c39ebf3fe7f2ba429c66bf78c858d037df666f08bce6e93df91758
z27183cbde45f7a0d073ba4ef0482e6d9b1d58d5814aa7d9fa092f686108d8720d236491f71f84a
z8b63f75bf468abb929926e3c919d397a1b428457beb5613d217342b78636dfffa3fe4d0f37994f
z551202a720a65e1214823f653124ed682514f082808bf931f4ccf0f172a5a85ca2942d854dc891
z1bf56b9404b4b5938b3f179e4c1da29812ec08379b72c58d04efdab44e7110a357e49e8cfee558
zc587755428db60df23d1d59ea32b7a39615292814853bab944f5c559e326bbc8d88a5d243c8c7f
z7e16a5a646e17ff24a8b60ec4d0d30acb1a402afc729b91e2d09cc06c6396dfcc4ceace61dc68f
zcd34aed94078bc354ce44da422d02450ba775459c1d1a5c9763e19dd49600bcf035101470e91c4
z3d6a7c71fda40ba5f0e9ae4fe43c41c05817402a984a605ef918cd0e79f87bb62164e8e442111d
zfa182849a813eb2c20e08e6357fa458ff1d70c1fbfdf2bbbfa3c16fb2f077f484f25e701fc95ad
z971e4b1140af4d87896b934c670eea1df269b1c720a7323b41b510ef4eb068456e7fda0f8a34be
z6a137042e1990dc5d523753dc8de5e27601f956bef538dbfb1dfdb4ecab9897abd7b0570134a3b
zd89abafe6617941a5d69d8abc5bf340585bdbfb76d0b9ee486522ee7cc97cb9b0d781be24dd1c4
z701d9d58e15b09b57a1696fe430bdfda04858edb5e1617b704bcd18545043bc76dc21b1e3339f6
zfbb8df9cbf4bb7896ac90e5582e9eee3b249b6335e63b8d98e793ae17620e9d2749ebb9ae86390
z8b10ba3d09acdf4f90e846c6ac3379c2affacb61c49a9be450b73ee0da38c8aaf856b671a22122
z94f51787b72d9859d78a040c830b95d63a4dae92992dad594434117e0d51f6caf2e7777dedb9d9
z63c54f3d0ee93f4f1a72002cae3a81e436af623ca57fc1059e87a63ab46ecb201ca3d9940caeef
z84616b154c874f9308945bb727d12ee889fd596396861ac4df61c894e96f65c0c3468e5a1d9e5b
z0e19891cd2c9b75b61b2aa7e5c6db387c3fccb7d572e04ca09d7dd78c30ef7bc0ef63a184a6dd5
z1cff5c8b3d34d65e9dd5979c3a4aa3c073f1d322130d9176b3da500ab1d9acfc6ca22e919b7811
z45a4440fa2f4c6b0e48f344d58f2106ea401abf6329cb1b48a45dc2905f921b081497990559d75
ze2db3b4ef914ab342b4932a51abe6721da55daab249b9c2d56b8e76a35f94ddbfa782827eed8cc
za5728ddb9ed64945f33f251ee4c88d8fb713a52eddd978c36b8be8bf4380c83824d37681243abb
z37c73142c3dc96ce9e176c281c67ec059d4365239eaa7d84cf91ba5f037a2a43df99e623d06658
zab556ae5b599bb42bd2cbc1d751ed00579435ca804508c45c5b91a21f4445dfceb300bcf27a402
z805e62edc8781e45e037b6067585a003885bfcbf05645e73fcc58f979d30cf6f542d148f7b02dd
z64da34c08c9c15076c22f1f47f79fd43d427842bd17614cf9c76c13f810dee07650df270d1497d
z8dfbe5e5b4dc4300415205604096c37b1cc8a8b09d746bf8144bad34f47c19023a45072dd3b36b
zd1f1b94f610b4cecdd6efc891a3f390f88858cd7be6a077df57a497030ef77c1d6e1d6178c33f0
z979417497632ae6aec1a64c74ca517edade76f637e6b7d851eee07c77d87019e5914c7b8b8707a
ze069b680e30374745863d3d79f483cd5a2a90c5083cab2b5e3fa825d6062c8ebab36c64ed431d5
z5ab561343f1891dcc1792e3fa2969778def229b842ff2849ecc4d5333270c02ee7db100f87ecb9
za0432d826e30fa3aab1160e2c0ce820fc4cecd9bc12e4de8f7478480be550ce7862958eee9ff6e
z890a9ad00c7f4ed18123cb718f13f0db140e6a554029c62f59f55e01256152fc3d24d96793a081
zf9432f5610513f8167f787ae7a17d709fd9b63fb20536554e11690fc5192112edb0c70a9b4a449
z03ce3e2e57849faf1b3db219946ea04a01b18056708165edcea8f37e136b9715177f91c8b506aa
z0ebb7fae1b17ad72b86445e7f39065dcdc01c427a96c551c937f3c3577e6fad7a068901e020899
z5893d46ea53f1374ab405d7ef045203a4a256205d2b79f3b61b48e7ffcbd09d7f2e5e82968a7fb
zfb8f9f21c0d051af22725a0c431898279fb6e9f19c21c6906db9c0511aa3312019e5a2f232a232
zb5d35a6536a042997a2f2c8f177dd000d002f3ee8b4ef2d80510edc42e5cce326f40e327ded13d
z105a629c49e341d3a54ed4a9bc89d51b9a142e9322e40172b157a4d001c19fb4050c88aa4138cd
z22dba2ddc50ed792cdad5973c6a78226d6d04fe3776759fa7d6a7ae445e9a8541a7c83c1d1c0ff
z74ccbe2825442c2a52afd0739d9a7d3898ebad1b37c6f7577b8015725b9e4969b125856856518f
z7164fcde09e2e69c32e02651c7f5aa7ec8a58b03c640f8dd03709e25b7725fadbbd5b886e9ebc7
z4371cfd6365435e267baffc25c96c1a3203c681fd243b5fae560c2e2dca5d39587625b2877bbfd
zad74c00ea1d67cf3d06f9987a50c7789782fdce8390dee16891f829409fb2d9f295b2f63615dec
zd1b871e98e18326e217f237b5bea90ee1a03d9a5face9b1637a3401e8d0366cb3c5ca7d8db15f7
z1747e95c2b8cb9f63b0c9739155468ffa728cbccd8088b754b78387c82a67b88eeb543625b2e2d
z132cf8afc758ef83f005501cb7f57d8cf142dab374d73ae86e6944c0a2e6b7e7a3b69e43d4b64c
zdc2ff2fa39268f32d2f3e8cd6c5d1669152cdcc9fc33a14ffdf71f340631ad8933c8b9aace40da
zc996be01db829ba9f481eaa756f67e01b414421826b25bdc000b26c16fdd5fd2c36ce1eefeca45
z14a80067fad78a16a226fd152388a3400286a68909d4bdd7075c578465dc3b565940fa4d980032
z3c2fa993538b095334186da6372ed0ee0803ece500bbc22b3650123336cf0c15a3ee40cf5f0512
z0b6647a58899f9b560103688242883e06aa572d3e8ae39b71c490f9da06a3dfe36f5022f6b6c6a
z5715ed7e500ca2d0bc8797049e1a22cc9bc39ce67aceec0451ef6b5aa5f4fd0837d2d51d7b1a14
z265057f8b7e4d68ed6626ffcfe063d918d4120ec000c785d40268a9beaf0d30fa7ba842f4d2a39
z59cc244d903c3eb290d7ab592ad1f6cece6ab946cac90548d8b15a61c50d105a4dbc97cde688d3
zd53554522ea5043a8c44a9a390dc0c9301bfa1411b4049fa8eb8f52474c02a3f55893523c78ab3
za033cd16234db184eae28d307b49b05a097a29c299238fc4d3bc95b3e2788d0556f56cb43b690f
za9f4e34da768ca4341f519a0ca507e7eb086ebc471df5819a8c24a353662501898efdf0b2ce437
zab64b0bc59fa60a557e8cf7a6e1e5427de7c7703da6d00dc7672b989ee020439693e0d9aa28ede
z895ce4454611300e82411782cc2a36c901be80420d647726bb93f47bebf9db8c44d79dbe65d82a
z5c66301dab10ffa18e34ac211671f44916cba85e610c3e6a69db05b13412ca72383f73a657e1b3
zae32ba6d7d8a461e3991b16aca7a9623d53c8237ae81ee7bd37a807f074294adb71a50c1b74f84
z006855e8b4415436d2142a1c9355435c51e488dbe37b6b07e7922db7f585b2ff7727942643e411
z411411d61b983a2fed9d9d4cf807dccfcb9149a20bcc062f7a7a4bf1220a42ccaf5009df354670
z4646fb46e90a5f34872b0a265ca852c9d2521bdf20e82aa234829963fdac7bf2dab0722758de26
ze01963dfaf29c66b98123b5cacbe62294ab891e0631e79c6037571911d80a11931acaa09511cab
z4dac261823eb533d98ff3fdf248cad7dab4faff1b4a580c1cd87c831abd64de728debce5fa7f08
z5ad66966950136b60ebbbafe010f3322199fcb92f12281a9b0334ad698c5ac0ea7dcbdd6791d66
z1cff297e0b7ef86b72600f45a9d0bee46cfba482463355aa28c7fddd494a26ed15f6657c68a294
z2c02c90bbf54d6d2a4525ffeebfdecc4fd586fa1a275fe7fa0b3c38c95684bb5160b06542e2eec
z862b6066ab3f8f8354bde77c2f32d310e56e075029cbb688e14197dbc3143d4996ee60a497a46a
z73706c6314a6b6b4594a70cba781689c3dc8d545bacbe0c604787faebfad1c3cdd6cc2e345e0fb
z9c283b6641d92b0a358e7470ceeffe14291d068403eaba9df376e547528c191989de88bacaa493
zd4972de6ac463f126892fb1abad471703f73b310880edd26ee8069757cb0d66cd61fafb995f9e6
z2aab7309fb3183c1512f41fb2e50221c1feb694d491f9bdbc92fb967bc2753a785826f903315f4
zdc560d10355559ee49fe34ff0521563b2c1e411d147cc6f98defca31b426d99a489264d24b7358
z096ac9a2c02c8882b74962a9e0141a0aebcc45256b933777e85ff0ae175c10f58e97480cc95ebb
z54dfb4c00151f0962df217816cae640912be3410708b550dbc0c1b4e0f4896684b9778730e45ac
zd525fe4658e211068ec84951717ba10a21f464345ba7b11d2b6dbc8abcbd753b64d68fc89600f8
zc8c40b1be1c3ebd35302980bf50deb64dc2f2846b5a2413face6b6690d83238671ab95906bbd66
zaf6365d1e322f70da11a74ae80538f92656e432abc97aef75084a20c1e9f9f86a2c4002de7b47e
zba9e9e6002bfbc43a2748d94328a62b505d643e72f0effef4f23243b224f6a9db3211c6e5be360
z2b0cf506557e232ebfba575701d94fa87ccef80ea5cb1edee8ca9b63ced89dea5ed713b10a2e6e
za67f71c0ce58801b983f4264307a9000a6651ddae56997b08098a40a61d1165566b1909f8eebde
ze926997a2918b045852c113d5a4c157121fba1920114a6b8a740e4fbf9bac8181de14486eddccc
z31b4dd4783fc4f97982863683788175509086cf4e3b4edf46a54483e5983af80e1f146ac31e10b
zecb9a6ddfab4ab56687b24e3ae0c8bd5ad10ea4c7fd18e0a0364a23a2e6ca8439a3c168ae2dfbf
zc18ef344f0a301b8269a937d3d27c79d8470393956940d464948aa42bd28278cb265d33e10e297
z7365ea9a69119c1892ecfc60f9d660d953d15bc646428ce44042a64dcf6256619b5493b9e5ef05
z6c2258b1f4e96f7ede0ccf2ed9d6476291eec3cb01fa9c6731bcba345f20ba0121031c55da5f1c
z0b2197012e266e163fda7677b28016b133ac38f2bba0adc8c0b89f43927f8194834fa19a325eb6
zdb00e579da3c4915bb27f2f87dc58cc15635883ec7bb6e7b8bae3b63faae0f5bbf27a9cfd950b2
zccf9e64ab501b8c16ecf7f446e382c836823e51a5c439a4285e3e05c98721b6ca3a8d0d3c56189
z834d6110bdc4dbc09659467b21456700db2f42f8e1f230dbf30336685ff5e82795808f2a708706
z4d4bd1eb49be227c2567f8e43d5d70d5d6053216af8e694af8a065f0d939082b9e48e683e63ac9
zb764ebf5090b2e686e465d11c035206d3e161f897f71177c9fbdcd3c637fb6869a4486fdb6df14
z42d9f6945602fcfe305e81374e91c225c553a9ddce89d212e212f5ee1b3593eced1805e45d4945
zc731186e81a922a36fd0100da98a8fe8e1e1baf5141310328d81a6d3567abe45464d79f35211e5
z242a952669a8d514d815fbadc48d418ec7c71d84c41211d3dd688340dc27a04c62e911b114380a
z79519789d857d11563bd8d5f3deeb5aa606fd1074be4fb0d9ef72b154c256e198a9deb380fc285
zfe918920876c737808bbcb836b80827506e94c01c5be1908d1f6c51f8326043272edcf88c5b179
zaa23c7fd27d3de66a5cbeb67e9df6e87c9878f4d5733d7915250274d2650fe521ce4a7d3421d0d
zf830e7da594ea6b14b1dcad5ce5734b36802061374efd8388ef3662c837dfc1cdddb7882df119d
z14b2d4c0964bd495e1f653a1bc21aece4e4170c52cff7db96f49f591336b0dd3b11e2dfd4c243b
zded1266693da6a5f7548a27f9399d400f9c13d13548b9f0032389fd4a92aa1f005f841e65c4f9a
zdb0c5f5148644179163316dc2eacb9c3466709a47a07b7954190185baa69a05a3f79623ca252bf
z7aa93a146ecfce9a1c6ba895c1ef9c238621e465332f8ab200f52ed95de95156f0cac9f5454306
zc94ce9dd21dc13520779a13aace2126e48594eba0935a3aa2a979d011a9fb2678c0230f5621d6c
zf0dc9e52330c2058ccc697725611b2767cbce13c5f86e1cd0837e448b545497ade6c32bfbab6e0
zdff40a225942c12d1f97d8081b3843bc11608b7446ee63e0103f798a3e948107d87a5c66079a56
zb6b232f71ced87abe430489983d75f13ef2be81903acbb062622c90c5b0c5a651f628c464ef9ab
zd61c5e4c1849b5ad6d1eedc08e2d09eb0e439373fd50205cece5033654fc93ca8cc01ffed108b8
z9b376ee0cd5b3fc2f5b7b06bbd8ef9bf3b3f708c8fd7e70215911b9ac565a5cc023ed3dcfcd097
zdcd0738ac412ae5498e59a33c06bb7a1f6391ab560d5a6b67799beaead36331afd282abdf9147b
zafb0a806197d5c6ce406278813351d6a1df59d64157535b2199690a11e30bd10b152f2c6c5293f
zf932578138686baa92250792906db849a52e388e6ff366358ebf4e26ce0113d0d5b2193d6ff5e5
z59aecc87afa2012d5bd6fd89b76ff6209aa0ed6acdef4b4805674f24f92f038b79832e95ee209c
z64c42747a55564ff75404307a6ee38ce46e09c6609c7a4c09ff159bb3446b47eadd1ee9d6c9eb8
za8e7d0ebd5507d9d9e6b3bf67842adbf24e929f0f5c288a0ecaa19eaf06b87b3c3032b0b4cc9ae
z90437495c2e1feaa21da9c24731b9c9a582a46577a8b314688ecd77d643a95858ca9247e42b0b7
z8d0bbcc70f627af24bc7f280dcd9cbaf1e332df9141748ca6140fc4ad8a26fc81d5c8cfa7456a4
zc649b2f833c352ed3c0ccf705403f9a45bb3eadcbd38fc2821dde1c694c08ebf785c1bce5786dc
zb05cd56f8ebc6c53b79e51e49aed37659b64c61040e197e650329de54100298d3efb9256688df9
z0e7d31f164d6f95b2f36cf257ab25363b080da98e3671445667c26492b09b3c3e4b539cff0468d
zc5e58ad1f7a8ad62903ca7d12d13b29d6ad5d43dfe1ddfbf8441414d2787da13ac6bc68256b068
zbe0d469f8f7a46922b67fda899952b188ab73a020006cc8bacf51dcca065831376b18e34c4a539
z4dde0a1e517ec915fc57931fbb167e20e87c826ae36fdd88ef5613b70e64d9b15bf65bdea62319
zeb9dbffe75b131c284b8252ee51f0bd11847f6900504ed0277d720178fc74a031c5e41c19c7ad4
z1f44295754dc5b76fbf9e6b0be6a8f2b46691f5746397471f6a8da05b61a0e78e64cab7c468821
z9e9a8be360e5799f24db9b2eb0c43a7f1c04a2314f821196d59d3e78045feff4ce16f1fc5eb9f6
zee110e96c5533830db256bc972c0bf4370821b0ca2055671abcc3162150c5444fb71bb9f342085
z9677cf049a97466f2a645eb7b5b138bc47acd80883bf104612b63c5aa648475511f246650bfe23
z2c092de411e5b55d3ba67a07d86e78333db9d2485eae1301385e471252da24ce3ff51a0b66beaa
z5787b0d0465fc8cee734c7b35b55a4f86e91157223530bbbac83f4691bd855796843c4a629c50d
za7d3d7241e1c925d83fec64becd22ed467e4e9953fb9a26c91486be8823031f943ef8fa4448bbd
z7a67510b1512dc96ae916bf9063e741c48b0d276e19975f3ddb9cc58911b892940d91df802f918
zef827e83860ed4ee920882762962f7137cd31d062dd1ad0edb018f4f226d05e2e0a7e71b1d6aec
z9bb54ca40cff4deee8596851a3b31217873df24fc829b00e40d4ed0b9d1ea441b77dcfc8c7ea9c
z8f38629c6b7d84ad78ec22bd214fb0da978a6b7923c00af6b398640bb89c365b39885dc8be9c9e
z9c864c539954b175b7bfc8dd21b02f6c31ffe86da6efcdafd70f7832408024f4a777e9ddccb08c
zd196873e2b14c13425ab481810856f1b59dad341fe8d5ba0837b65cd676ee034bde71e159c5056
z64458368b5f31fc05d9d89fb2353aa4c0ec5516dc10eac3237ffdff4177255b70eadc369052ee7
z878951b76859348a2a1422f95327bb6c9750ebdbd4da1a8ebef06954f8e2eb27c875bb08e037f6
zd6652d6e32e832c3751352ebb339e3ae5e2750816e61e847696055cf1fe2c36941a500bd9a7527
z7bfefa78d5ead47bb63847605b9c6c827f1dacde2287ba21a48a4db02956a0b2bfe51d52de6c49
z62417e82f4a1159d90bcf34ee93d9ec004f13781f235707ccfb8bb5c9552b93743cd34294948d8
z8ca56e448b168df339b9e3a4cd95635158b3b16af30af523cf05c2035c8c0dab176721dd61138d
z8cb2b30fbb67f35bf3c60aad5b6a69dba5f899f6c3d375e7b1443e7a5287208e887d03c4c94e7e
zc352161dad5aac403b1cb4bcab8f69c91c2a005d99b290d0d58ceb7e04e5efb07c1934123d3dcc
z6daf56d42f42463ec8226df08b1563a715bd033d5f5210281a41b89ace34973737740d3d8ca8a4
zd2b978afac8e3ab82241998dfc82e91077c7557aa08989cb2c06d2e702ba558e8f5eb0505ad155
z966f5aeeea83900de48e764a4aea0d94dc1a15b5b44985c7ec3f0f668e1a37bbab4ed64b5c2616
z5db6c1d5376e565f3cc17bd78069ff1a78a94d834e2cfa52dff62738f25026fe2acab8fb9b26d3
zf76154fe906cd57af79f72202a6d6771e6846ba1871e4d5fc329cf6fa2fbfaa3d0ff7c9f63c8a4
zc2770df1c309cbe8b0e721b5279acb8a239f15c3bedb722d85fd49bab347907ccdeb0501080ccf
zdff9963eb1b65538553897ea4dc523797095b3446b0ce4c71b9e089635f10f29876e59da352d67
z73910e561499dcc75187b7739234b3b0cd665bc72f5873aed9301031264310efb1d92ec101cb60
z5a3ff3a62d7b6c52d70ae3493dc6fa396f63023f0d2df9972f0e24d70dbc8b3c157a8272194f0a
z5e05e8eb6f7f944773aa17309a0eff2772d41a2f1e2b667efb95c5a5c3187eb0fb64b2f556db48
z01baf35dcc0c70db6e110d0f0bff623890bda1aec7725ea746f9a9541abfd3fb90f4ab5cb91117
z4b2463c369ef96d23c30a01f28b300a633c3a44d5c1c94007d0bde93364d091540265a10b500a6
z204d89b00461b102e4dd3cd1db1d3be11934220a4191f84b62b91b78adce70f4ceef6e6c704596
z91c933b9cbb846a5038f6539563697525285f0ed9f47ec24acef22618457aba7086f9eca2cc7b1
za6e3056853de85b3cb37f144215890d4bb0dd653a04150040a8bdbdc8b185574e23a552a9fa7b2
z85b7616e983b878e1831b5202fd72de609dd3c219f10cf8f835d66a1b5024fc3f54627a2c1fdfe
z6b6c92dfdd42af07162d73f09cf739fd2df4215ce04caa25dd6538f3b008a4b37b807634c33d81
zbff04e61a57b9e95904d8d14c8a4e1d9728c138f0823077d994d703c72c43b2090e74eadc59688
zb63838fef9ffce6b76a897f9f264c625d4892c4c7dbb1162d4aa849845ae8e078783bc37e45710
z85781f2ab5c7dc22548b62f0963ae0ba46395dfd36614959b7922a88487f0ae84eaf5391d0c164
z295f492b5959d233b358953ddca1f87416c02d27d48b74cc3c4ebf2db507fa19f35a71d4e235b3
z02aae89178ce292867880fdf3cf579d2b345d01f1184e7a1802f9a1674a9b0291f0d819c84362e
zed0178af8f8a314100264b438639def2316391b29d63add41a6511f3fdf2ab9065c83c02133862
zc7f701733ff102aafd90e49d31b4d7b2ec54bcc65ff8d6f4202ae6d9519f18ba1a3792d1ac386f
z3324c674857708121eb19dfc87d36b8b11059f37abb99cc814e8ff8982bc6ab20626f915935653
z9f056703e2b38e78c985af8aa99f040d829ec2d975320feddb1bd3364ebb400bb261ab787e2089
z1952f2098fad931ad45c8476e8bfe2dc0965ac010f2b1b6d481a8ee44be28f4fc64ee9e71f28ea
z3ad8a5c0c9d56183c8dc44120bf67fdfeff0a8e322bd688e2035bcce61b4daf18f1776299e4f27
zee257d00a0c0a2861a61b34156d96248e2775c41cf27c8dbf16a8cd3338b999c84265d3cf5e477
z35892e5e3b4e79fab026bd306b62e2b405b6828f10805a30eef109085c5e90b24012f9dd708dc9
zcc080790f367f76619feb649bf0cb2cda6aca63da8942c845902c84bc54e2ecda3db3121917db7
ze576121bbc403442c0cbb11d9f88603d50a05364e4e084f1254ba5b88c8a527a59145b19d80153
z23a36eb84ef0469444545c2a79eb6a028bf8d55f47d2408a0ab497a5bf8f61042c67c3937fcb1c
z5b54670457fa5c9a8fae1e98d3b5d459294fc440e1577f99205738d5e39e1e51367516185149f6
z67ecb05068ca019342367575f5d218b9afa2dd1874cf9c34329dcdf18f7e205d443aa54fa6658c
zf834a41d754ebeb555b8bbb0736fa19be3bf2574c28b438882c7614f961d6518862a0a44f881f7
z238ebf4057e835fc2eb18e4126f37176c766fd46b7d92036333ae90b8f8099b17f5050bdd5443d
za7c9a99f9e9a6e3cf3aae2f3a78906aefbd2e10892b5ef6881470dde07489dd1163fbf2304830b
z1d05af02cbae3a6a7a73a1432b897b6404f6567c55b2ee10c62b64aa81c1428bf4cb1c2c961eec
zddd3031ff40f0fc8bc7fcf6e2a6f5db1e0b38c1921c6f827555522dfe2e1870d3be2bb12744fe1
z2aeaa40dc92a4189a91c64fe8fb82792d7f31ff25642c9456de8fb3d747fa33972c5140ad6c20d
z23ea8791c82b991145a13830393ee2c50ca4af6c52b1d82bbcde7fe3445f3a968c2582cce79878
zfe268bca2e3d826e5824758a504ab2cab686390960547452e5f588692d72cc8dc7aa6efa6c7ac0
z2d6ff3da6a451b379e2409920ae386c301a2511be54ef376f394a26f3fc40280eb2e64066ba05f
z6812713e6d607223929c2e81783b08f06ab04835e61a1eb3a3a104e320f601200ac3c979293f0e
z967997edb12c5b25827b60004a424b0006d082e38bad82ad4eb59be7208ef2efa2f2b6b02afef4
zed876086589a8cfe0735eb7243c9a8bb3ae5bdf9a2a0efa4b35bd8125cee36bc1aec4fbf70b289
zab143afd1b3731e819cb49abd38d0a8e38a8fbe806f4f166aa2e1db58b7c347f3c134a60a5c33f
z4c5b0fbd9f88e47af8db16ea4b8acb6b28185d9b96bba368cee24aff3e612ed45fad8cf7cdf220
z918477a7e6b5a8009946fe14486240e730e2dfd038adf02418f688e91473c0881e79c342c3d117
z179d983fa2703244cf1b8fb4d19c587d13ea0b62fdbd0a8efe3b09cdab0e83dee6ac8efc75575a
zf92d3b5f1bea03f82a2f95a2e0d6542d19ccdf6bb1fafc3742493f39d37e35a21091cc963a8456
za6ff91f35c00ae10dcdd63fb833435c6c3335826e7f57f7bd88984b3ba717caf917c196b5d6398
z18f6a21c88a5086e975c59db3cb3c6745e5bacfb06e58a4aff0c89473bd8903f4eae9148d642c7
zf884ab756b58cca68a92dd1a4077bf6eca9896705fdb55702fe42aa5cc1cd6efecdbb657bba10c
za53d43309e30d14a29228253b7e23f116b2089aa1d17bb92ace137fd76d8c3d37b14eca0d6c521
z95e4d1aaa6c68a5b5509b0b4267db266eb420a1ab588ee3bc97099a09fc78f706e22998edcaaf0
zf1d76dd55a862acae24fc16091168142281ba846dbdd226228d17ccd2955a1c341ad2338c16cde
z6cd5ecd8b54a55d9c21a436b2f94b3db3ba468137c1748eff9cb9fcc2360425f69ee6391203dc6
za71acae690325999acc36bf7bcbe075fad2fff882b01ce6328dfa2378867d96023c20b5204793d
z7854499f4a67c6342fc65ecd693c326c089a52afedaecea4c34f04965cf33121ea2f7bb02d356f
z7821dee19ee2d33993e423ded94d375c223d74c3412d898907a4a087071e5b467bc907fa2cc31d
z7f05d8f7ac14b50b9d6fe88d68ef67af9891733694082f40651163e9be87b38ab4821ba489effb
zc405459b796bdb1510a09c80aacf7a93afbbd2060365dba21f39fc70b8f40314c70f9d1927f5c7
z927f138bb525756a7d5a362548ef5e83873f5849fed045fc5ce971c51173555977fa28e5313d09
z0e18ac757e3c38da9bbd0c01a003ea09b4ea04fd7c9e9c1107543438a12b45237ff3d16aa95edc
z3874516220c676c2c7aa5016f30d49ddd22bf412e1e97da09c4c893e9c61f3553ca0ea29765e3f
za8f0a85ad44d6f38c8eb3bef55d166609f42420b2f36d1d4dd0ec81c11918725d370ee841a8355
z009f0bfa83cb84eddad856d018945bf6ca1bcf03c22e88dab684d4a3ff56057673f893e03a1267
zb690391f49d106334e209d0af78201cdf13aaeb9be1a8288277aa859c6b59f93857b8cca6ec831
z6d0b906e3dc9d3ac1113325b33490f53bbb103d415761787d1ca54aeb460d96c11f0187b9a75ea
z22831bdd31028faae584eb26136e520801eef0ecf5bf07274bd77be1717dad8e783e8a8135b96e
z3a82fcaf6dbd382b26d28bfb4f55fa76f9f1f43f0dd30da9c736da65b9ba80b99bcc8681dfbc98
z744e2bbcde1395cd53321cd6c5ffde32309ec7cab8393e638a197cd417284354d067eca4d63ab0
z7d0076ac7d404c65e1517dfc33b2672d425da1cc5f54ac4df46cceb5f7775abb8bd9602d105d9e
z2ac40d988e683dec85372f7efca522acf76c926628a81236765b7489bdb645ad41525f69bfc182
zbec5f40ec1bfe4370be7e920aa7d03893c827fc0344e5a4dda24a350eb58d86827e0be8f1b8224
z07240d00fe8114c6713e0999c2f8f463111008b625ad7688ffa44d192b49ae590ff9029c0e915a
zbc1573bb266918d34fd17f05f7eada5484d8b97fed163886c9f6ebf09675ffc26e8620e955595e
z64458ebf719c75f4c491771c3b2423da2c28f3b6996613d0aea917ac284698d980658299995fc1
z630bd92d52ed11222167414d5b51038029425ca80e8cc09d9143caf040f6201545a804c968e68f
z186b942d0a5a6d2381290dc022d6cfd9094acabe295113f2d0d8d9286adf0c92c3bf8aa385ec9c
z546a03b18c41bcb42e9b40dbd300fb41940cdd0b7b5acf12f9b4b4d688392876665e252b03fb3d
zbbd7d47585f57277505fbfbec50caf64016175e5594d88b5358b31ae58a18cf42115516bfffe56
z03f08e05ce8619ded2b398f450efd204a85b4f9b5f4b66851c29afa337b8cc7641a6596ade9518
z32050c7125a7d5a5d05f7812f722509b3e1da0154b599a808139c4c7f6f9b1afb01253233added
zf9fb05c322e2670fb2898a0c78eb0115b0a8716a4e173bf630033d1d8b378db145dbf31c072a91
z73ec777f6a9cd9c4a49199be3ed43223384ba7f2d1c6bdfb7976e03b79bd23e835f8fd8e186d5f
zab05233338f5c148cd1490668dbaf6bd3992accac667b4a6da4b78ac83ff307d6f5f033dcdcbfd
zacd7eae1919d5e4c1133cb528109fc04b81d568c06a56ebd3c52d75a633e388ab893df58c5d1ac
z4150e241dfdb1827747a56b670dffff72eb2e881e30a0ae828660dd75bc3b5fd51d24d67f5dd8b
z11789809e6a022a85bd51765999593256b5e7e12189f5c764a827464c1e949bae76c0994a2cc9f
z3ce8dbdfce722b25c5e36b9b535b97e7481eb7f84891868b4406e0cf4a29912865a6e932c70f83
z610c59f699e55e6609c9fea8458297b4cbeb079c33dc7b2b04e8bb2e417837b6deb06a54dfe4bb
ze5f4228e7519d055fc01cb2707799edfea4214d0e9884ee1aa260e39d691377e546473490cb26e
z9f46c4dc01030a5b11007ca9409b0e9b693df500678a481cc16753aac35ac4e63bd575885120bf
z2a8810a315c8cc84e4764534146e7bed4c4041771b3e41971a57333b662cbe36793fa73459f8df
ze522b3ab35dc4ce8f52b04c21b0cefa7b7c70400f398431d58170b0978ae2c7915115ad49f3417
z06923f64c649032fd262ad8b54f4974d0e64041894a6966fe0254f072f00c232a241df6e86d97e
z028add631901b3e0356c0c012cbe1ee8d3ea494ce89ecf11f85660cd714c2b2a22273d88f7cac5
z18f128b054543aa53b42f94b2309896975c9494e359088b58bd188942bbb6788f0b2eb74653ede
zf7734415172c50336c8ed1ff86ea94035b86cc475d24b0e2a9ce421f147cf9ca43c48b8c97ac4a
zd3ac1d04d1993c4c76ef180763008fad0c22b54b7936c67e88e25c15b3bf85204073395415452e
zaf62699e363301391e318779fa6528be78fda4bf20f668951d92daa5cd1239c9f0cf35a5e5c987
z1ecdd172bf706db54465d3d592b76c834633524b2ea42c17ae2f9e613a69c4bd62529dd524fb1a
z54052feb332cf3c57d1f7d90ebf5a972951f0e012872fe69ab236dc0ff243a2809058186f25c86
z8309f65fc3c09d6c65dfab3d4bac286a80faa9d8f2997790a3c3267fd43bda7143ca97f7691e64
z4771540583018b41305d3a0d8d02fde592d0cf52e9b653249134dd23fb6088df2f17ccf1ef3dd8
z749312370bd7f52562c5a945dcf5a9b9da71037a16017cdf538df39d05a068b5800b7086a42292
zd8d82be4343f5a32c61c6d124801fc3808e32585c6e29debc33b3721522d9593e3f2d27dbd1d6d
zf27c7b3968efdfc3d862e5186a8ab994e11a3ec8c45b91ee9e8d41d425c6f79c2786b759b26c80
zc8600734e6e457515132d946cffac2d2b2939c91a8b2c3d815598d984909912442adcb59bd95ea
z340a22809eed82fa0ed50f5fd2939128b7b818f09bf21c20352ac1416fad1215dd1614389e7a07
z522c9df4add5749ac59516fb42e1281c5bfc6f6edfb3b240f2dbfb33cb9cf5f7353d8ff0c3fbf5
z6723c6ef85def74fe185f597e9f9c295d0e92e1cf0748b1916dd69dd9c9e2c51c0c25598c55821
zb4ee6fed9f77e5c7ce42296e012615009919c544194cc4310f832c26e599b7f64e8c3796f8a8e0
zcd0de21e80112abac637d8cf9636befcba7d193619b596e2ba1037f2ddaf45b501bbc000ac0aa2
zf374187e84cdfda96fbab2e66581f5a6d978c04907c2c5f578a84cc77257d92caa79b9f80f1b03
zb34853f03f7dc1e6193a8d1e11a4f4dd68dce96718718bbb1e7d6735c812e42161687579726876
z12409432aa60a9762e49de60b0c65f00e67cd6eae88c7bde84684c932748adf9beb1f50183540a
z2599bbb86a9a0749e34471879d28e0a4da47b70cd39f999907c430c1d9317770248239bedad5c5
z85b813daaa6c20f22b55f1248afa2615aa50382a4b47b95888060f2150b6886ec064cc49b97beb
z69649610436ebbf7180ff5c893f118ebab6d6a2461720d989da3c79d89923d1d1ab2a6d049089e
z0a286225f26996708ffd4fbf8c8f7f6d882eb25476ea10ebeaf098edc49999efb894e683b2843f
z8d8fd4833fcf9193ff06d93cf980ca4e8ab5b00aaadf8080827bdd4393fd1bc4be466f58a58d07
zb7dbbd75c29058cc4a22dd5bc51fa2918a3bacd0c6f8dc3f81a79c07dcacfb9f834041a626d899
z883747c88c2c1d551fd841266084a2366e00b6426ebf2f2b04ee0bab6926b646b80373cd858967
z732f3ae54ef7de56d4d7835ef30354e692189073aaa1da07304572aaf5b8b9a958d7ee413e8e6f
z4e358f20b28ee212ed5fd70e670cf111039d0f288535447215a2f02aa5795507260509f3ab4f83
z6879881859c47e0768c88f6399fbffeb9fcf2e06704ff4e6d7291eac073302fdcd483a27b87564
z2086d68a02acd81416da4a8b3dc00469c9f4b71a8653949682e1cf566e30f81f85a9d880e3cfd7
z234b5688067bbaa5d246fc59c5d44631a80b47987572d339cbbaa750be55090e74d5959a80bfd9
z1f022258bd18ff5f080933abf2115eaac4c7ce8f497cbe57e3d7c7b4d6149957c03174c4f1b8c1
zff4c79763d07a4b06dee4993f87c7565ff74969bcca28058c5e70bac5f2c9b068133134598b400
za3b13e6e71b8919661d1c4bd1142003073b799dfa06a28bbae2ad7022767f86303127e09d53860
zd6b1a1cc5fbd4752b989f9fc8f994039483567d05240861f6663b1b93ea73ebfc4a4aaf8ebebd0
z356e1def6dee5403f00af52b3b4771062c730b4adae450a9e0d50f9c75f3968e1eeedea6b29023
z6d7c2adabc68ab43111afb24bb9f132ab8f47bcf7274d6f664441985e720ea056f6c22ad86d52e
zc5158d1737ed08e311f860d99c54d2f5018213a412db3e464dfa59cf9c280c086aa05fc0641a8a
zab2c0299a92f0e9336bde52f2ac20c6f8841f55f3c4d430d0d7f249141e7dbe561206c1db8ed86
z6f05f9302fdfb213b572949503ef3aa45fea2c4a7ca395e3bd0f03670a68cce62a29125f52a1a9
za10f999b340bfaaae725d2798001032c79716689e8aa143083c5e7c7fb4a6a8b593f13f5b6a0ec
zdaec309d452ec8289fb2786dfdbb3f706dd9c01f1da7b9b22df6deaec756237055cf47a8ce1d5e
z098cbb70893e1d0f58a318af642c66ac61e04b55c526e452b7b303d61ac0d118aa3ef7cc87d4fc
z0d7d91839d269267acd058e3830cf2220495018bace25c9afdaaae23b0161dddb6c085da860061
z92e2478a77c73f5b421fdbcc38138eabbdafd98fef454fd352091e98ca4cff8decb59be72e5f11
z2c2ac760e2813e59b41e3aa677d8fb39d4099a4d80a6c8ee25d0fb3b812c21c3564298f3ad8f91
z7b07ee96b9c4e78df1e981342de2125684910f87597b18c09a1d7c50aec6dfa1a7ab6bb11c5385
z4854fcce120a9634f92e2d544da464eab4ecbfc5f5d8c4c441824f6b51cc1e7d8fcf7b3bc0274b
z9bb247cedb99677b41f9a4e86abd9dff47527191bb5afa30f9bdee77737bce50c491e5cd21fa03
z1116582f87114f2267b3daf9132aa331f3bd6af2a58c973850d8dcd288c418e009556de3c604f3
zc763afe6adc874e3aaf22121d898e8a03839d057399a7931531082ba4f3951fa62a6334bb5b0c1
zcf3e784132e7cf611a15cc5867bd71edd39622ec0dc87dc74908926141ea1d5e24af7070933a81
z59d5360796aef8815f236de9c59e7db09be76bd5223ab24d8f102fd6af74d8db3f763dd8343c80
z45d5f32c5ee72fd68a19df713e7c4b6ce28d2c4f1f2a6acd8396227c0ca7edb06a898b90ac81dd
z544fbd907026683c29a7092bf29da67bbd2b549079cf95fa11a66d4271852b2220b7913da341f1
zadf459b17b39c669928b523fca5b57e617e4c8326a27b7087b0780ad94eff9e7fce99065a318a4
zfa00c3096c6e033dc17d4df0112bad6d3d99a40a9b9ba80dd0ce577adcd73e37172eee99f3e043
z15cd7013918c74d827b53a27b825d85f938fba56f6e052c7abf62e25cd2d3a1946799743d729ce
zdaa1ff34295368a70d0b6bd98bfd2d11342f394572d091db5068cdd20bb2540c01e38f5e3073ed
z0cd591ffe5ca7c9294eeb4376d2a922031094c16d7d54b13f11a120a07575e7463c3793c5d79a2
zf9da29558c09942bb0cb99f01a523c95e68c95ea5caca66a2ea1ab89014aa2be5ed1e116ae1890
z40477830de2ceaae2f84aa56352345fca23e1bf037098684a355df474d3a9cdda63f3eecd037a5
zd82c683a07cb16cd8b2e176bda2c94f3b15c8eebd9a0e000c0e0fc08c16801679054b65fa56d7b
zb3aaad43def95e48bbdbb55754a71a99579946185f4d18d3d7986005350584799277db1ce2a6da
z47e5b5688db93027c1535a390a7d3e5cb1a1d24ccd1a567ad70193818b2a8b9604d9bfb5d30608
z7953b98d5b614d7b5e21a9868ea9b13c466752ffafde38bb0d638ab6061b7134de43eea300ff23
zea5049218ea7664902f39ac77253413941c5628d66fec41108c493d4c1553f35aa55d826a0e958
z6dd8916f1423c69e03242418b87c7762e4933e09a16494d76d132492275ac1a5ae6543482953e3
z48b93831c292afe15057e98934bdebc3e56d34ab8acf826d84212fc4ff99aff866de771dc2b701
z51afde59351a82d37ec99dac2c9c5c488f17de3ad5da623ba94c2c1ec5bdb0c4365207f45a9c77
zbf1ca7564ea54a5628c97a730f873239add9566c1b641c6a5da802ec5e0d454b839d6848022281
zd5c517db81f4c6be8d66dee0f5fc6efb5bc58154c48da841f1630af95f4c9f353c3a0ee5a1a824
za7eff256a28a6c1058e12aea25477371aad839a5c47447e5babfba2b301820a59c0a53ce763bc1
ze5754209270d4bdd089e1242ec328c38d438fe01d205ef4337cccc07cd1ab6423e63570a3edf26
z2494bbef59613f801a541c868975fc42b690c2c735225ae94f307bb979bbe296546a49d69f7bb2
zca63ee366becb2419b448a47c2c53a42726d52870e9c5c2d780610ec9410672eaf6851eba5b278
z97064180a6083499bd7f326fd479e19d4d6279e2d7ff068ffb0a0c8a0d0431484d91a57b561658
zeb38b4b77b1edd87f94b72f5a3eca2a7344afe07fe6d4751ae062ae77ab73421b867508b19f106
zdd9b592fe26f4ff16cc9d1d9ad090d598e1ed11e6afc80a0fbdb096a8da0ff71e4be3c1fc4f461
zcda58caa07ae6a6cb12b03fad38a22523b94557aa1421ab34fccf5781540308eb5789152f73132
z3f4e9c96f788aaff1aa5fee210e0249bee859403d1994305ef296c8f220c760b84a93bdbd4598e
z841845867632fb308c57d3a3ba58535a2592787a814fc766dc580954e131b338ec7da9648c8faf
zb4275ad3e454433dd7350855d9394d6b70cba325c26bfc8f55a5176d8e308107d6484e5f37e1a7
z8881043e65cfd8cfa07fad7cfb99be818316bfa1e90f472d18ba9c4e2b232a226e58e2ef744d9e
z03e67ec74c556e85c8c533efd0bd34496d92f55796143c8715e1ee8e7a8e918e935063c9b45eb4
zb2ff7443ff7b64cc4e12446d801053822ea20442c4326ee4459784b1216fdecdc234ec96a858ad
z2c32fe3d20f930cf63ee240d2f58fb7ee003dc24f6dd53d6606b99786478543f2062958a47aa0f
zdbb1fa1616c8a4032a095dcb35bc263d295291987dbbb42f685edcd130fee9c6bc50cde28f280c
z0078aab45f4eea2b9cefcf2d385ee964d4cd9f32c8b74f68e7a3a85623a86604eb18feb03fff14
z1be9ce3a3347b4b53ad6e4cdb305e56bac8f1303f41c09e8366c1cd125946d91381b67fe827847
z002f61c81144f65f866186fa082c1dda5f25823ad7cfceff4b7f79373613000ef9f01006671437
z5af5b1c7fb7c7f414fa694fce347e372feff7c7db968f3995f838a9084195cb653f2a949ead949
zf743c8cabbf1ba62869ff8c4c69ddb146b1d29c194eee49a737867f2f107604a29f0d2ae943f2a
z189d144aea632c73f60818acd2a88bd52a606ce9e86a6a7862bbe5cfb440ab67556e1fcb48f2b6
zaaf76a05d58ad278799e25a07b5e3432792126c2008a6450a68ed024b7e90f44a6aadb9b5b7161
z45fa4e3d6fa33120f0bdb31657c0d1aa20e29c5d9ce87a487e1d0017cbc7a7aa3a1a69973c8d6f
zbf06a7a0605ea10644ca3fde512a252dbc97cf7c5627e0992e9020e4626f1f3a1526713d41a77f
zbf0564a9dd7976db8e7855e755c8efe4bae5d3c2b1a3fcfda23d6b3bcec77edda4f708a3e96d99
zf637c6067af1052040e3a1761ff874d875dfdfd36d456be5934a821aa6474a5e106c20ab5e577d
z3d90161636036e5d4497253c13caefd746cdfd8c24346e461d528158db4f88f8a540799e775ad3
z0c65f4a90922be3a8522ce329da52166c25b26c5e3376f9782165011d3166898b1ce6a5c8bf334
z8c3e46bbc4c7995ae1680a28eb35f4ecbd211e1a9410f7fecd72bc6dab399e9c969f6353e54a0b
z69cac5c5d3ff5a927e1d0e6279086e003cfa6a68422a7a28b7b2343caab69f30e50ed4b6441671
za19df30e58c0828eb322c798586dee3987a820b0ef83cf455ceb6af7b40cbc32512c7037299d39
z6ef1405010bc29a95278e64e2bc4bdbab95f81d699b236b0e7aadbdbc3d9ee8bcab165921a254c
zf95e929f90e5ae5cce81298b392159cc60f992d1df23668e27ce0916ee31c9bf08af74be871ff9
z3ff62f9411988aabc6f61aa082ed8764e76ab11f633d7fe1c9ae770f64657fdcfa9e5c4a8b621d
zee557d21422c8cc577d4a565bc9a7ae694947048ac084e228741df2f27792e3aac2db631038f21
ze19d9ce741f1884167f2a5f374f4ee6b02ed7ccd0f4faefaab4e02c49af83cdef3ff46cd29ac7f
z6484764506ed9f7a2a56c03d744a923b33260e9584cdc64fc308a74945aa2d9a783341479c66ea
zaf546aec28675b499542eaebf19a5692e729bed4a7fd1cf9c32eed093130d40d9e9d4a9ab78255
z55cc10079c353d3ea5ead6a03a26b8b63d43d0173c502197ee0e1d063423e113b65d6ba67c3f14
z92489317e9c9b098c26a6dc7e6ea842811b70df2671d4a9ab9b736ebcb6bab2ccd2a5e7488699a
z6f9c1f32f14be80f069ace65a0bed7fb04591e99b5ef3f47099069edeeba0dc7923b75dee82827
z29e1132fed9569506f40df739e2d5a8e8cc25a23353ccc485c905bc1d955fb8da304573bab558d
z516cac27cdd1e6ec66bdd302ff959fa6fd33e2e22d6d31c06ef4f3c1b403098160aa3ca3052ad1
z3ac7ed9d9be94142c10814202b9816bbe6c6b937e45194f2cb9c55df8e89ee401873dde98f505a
z970b3d8598eff71ac94745fb228083c14f794e85a6c977e5ac009845a7616dc6c50ada59b787b6
z265f7dd1ffa305e91ebe2411c5204bc7d2c4fa89eee41f754874242eaa91507ab956cd07af0a32
z5c42d11e4ebd51cd4bf3927ae7fbc504964f81096c1668b48edf99154fab305518cfe5d86416e0
z4c6f1ba5c473ae01fe3ee5f7ff069b21ede61c223b9fe8f8eadc9033f188ba69095d6a4522f8f8
z589fbfc947cb091ecdaf9520013d83532cdf4c27c417776b7224bd2743974456475c04ce319103
zf5fc9f0a4cd7d49d87abab5e65cc51e1b6a3bb3eb5700133aa1f134a59635a78133f857d43e8c7
zae2dd90c2de0aa62901fcd670ed772b69c0f9dbfce4a7079e73e503f887b9b97351e5ecff6f138
za0b225237981ed2419cd34817a6aa74ec4251510ddc00f82b0dffb7e6caf678bd81deb5e1d9cd3
z2502cba883a4ad8c635441d660743ba0564e3e4b2575ce843079a02fe32714057b9a6d6a2a85a0
z8325ca5f33777cb63f4f6f540b56e486c08d2be2db90634d4cd743730fc36b10e1a876d640ef3c
za5025fb55a64bb48bc5d301e72b75c04be8b98cd2e3abac96b23b1aa93677af9aa36e3e0e58d41
z8f677d9619fde828efbe927c103928addb062214ba5099ca1ec3ec141b53fad10204acf6eef6a7
z4fbd1a35d877a33e6924dee344a516fbcf0daff4936a38f13a9c631b223a35b1f8844c6b0c7951
z5242e757fcb5126770c8f10b83f3a2a6722d82e48d15581896abc52d87f8a1a2e5216ddc941e64
z124f568ea9e2738262124bfbf98979e24d9feea36bb44620008620dcc37f8804cad0586a6037fe
zf2fe8057eead5bca2a914da9ab655af28e9d90e9282d609fe2ba455a7d19e34d13d937cbb84922
z4e82bb0b0fba3c12b30829061be0d4e7de3dbbb1fcc2003425e06c028fbd3e55e5c6aa1973e9ea
z8b6e6edc4a30a409cac522d5cbacc4222191588c03f70ead06f4b232e6dfcdc9f871b65a7fb3b4
zf1eeba6ae217ff9cf3c290f50689b1de875e6afea51db0274b26b53071e383282d2e79997710ec
z54dc542605878b9145081644643a5834953530524e3f8b8e7fcf4b14d4a716c4051e1fdda143b1
zf673acb0938ae415406e0b760244c39b0aa493df07cba84cb58fefb463aea7f2cf5cf49c6a936d
z1a8a191b76b94e577c22b249aebaf9de52c3c925b8b90c8fe8447b9d89ab3f8ed0aa82e5ac5e12
z8855a86d8e6eb2655a8576d9e503e64e4818d05a6c06eedb7f5ce34780011894f00b13f8d9b8c0
zd1cd8f01de74f094ce328fae58764d2a1d1cdabde6baa12415f8949809aedd106d56ecdd54e1e8
z483fe270760728990f9f0ec207979e74ba58e5aa40f010e78fad2de2a096b4d8c24881ed004def
z8980a5c581b555fc57b2e65d52d50627c878b566dce0ce3d00d53e1d5221c594927c7ace7737bc
z5feec7ae1ef42409c2888dc29c82482609732f0d349de92beed1421c36d4b0fb1ccf9be2a52fa7
za2913c70c41d18b7ca92d9409e828665c848ab4432f256ecb8ba2e59b9a0f90c27743d8b676397
z9f8582e7a2265b1aab301f946c8707c392a448b3fafd078d74d35a8d7c8f48777568284ae803de
z20ad7f27a45590ba02d04b12875846d5cffa44e923329796e3b9c614c9ef08ddb3977fc224f47b
z61d6f00ece76b666df10462df7cb67c7d22f6481aa3423cb66749a399af59ed77a4dcaecc4fd29
zb70a9557f7a7af590ddb8616068d9cd7fdf05a3f07e70f064b96ceb80ad1f90c4e827d441e94bd
zf92e444c674c9cfaea0d76a06bbbdbcf3b8451fff465c007fb65ce461b291d1e95172cc55c5931
z49621937319e6d9c6cccd71e520dee1bb1a6ac611cc32332986f67b0fbf6df5cdffa644b793c87
z3d217cba68c995cba8ba51826954316ad18e5ef4d872720246e48bc1d79e2fb214e73afd9e5f91
z771e8636de55866c594a6b25e9f73c9d00348fe86d03ebcd9e522f5efa2eeb8de4b9ce7387b195
z60c04a8a6d4453a051961bda4e73f80acbaca89fce685357d16c00061ae90554000b19f96d677c
z4e3dd0f1b40ca6e63a7ecd390a0d8657325ff2d362ae154af0f6bde475a903dc373aa29d1cd218
z2e8e6a5bcce1485ec14989fa2167328224890cf86536bcf729c845cf597bd368526307243dce19
z9f8431db996f9e317963e8eed27085ba6799a4d99582250a8000591e023c8a91f9dded77b2d212
z77f19bb3d5b22381102c963a30de96db765c7c51cc0dc2e186293962673e25c2f97272f729dcce
zd02a2965e04d81d0d76a9da89bf3c2e71dd5706bea7a3ca03f759f6554d9476081adff660a8acc
z91c646f300b892d23c92e3adab3b49472e3d8f614f651cf7c34983fac7fb9335680302df7a1573
zf6c3eb6ad36ceafaaa9a229aaa0910dd1e7a20eb4f7e6f323f5e098a13ad51dec2dc23b0a83dbf
zbd40f601c9535259ec65bb8ea3b581a0c2a087623a13035ae0eeae7fbd4c0f2daf61b201524659
z98edd1123251092e00d043142ba77428903ebc1d9da9cf85aa39a4601ddb482f210f2ad654a602
zd23ef9ef2c31a8cc84b7d99c0b65793612e4553991ad0a8177a802536daf788f4863eacb9f1fdb
zed462e0a4bf5d77721db5b57fbb1efa33649cf5f560b74b1547fcbb6765a58e4a58a12934a10c7
z4d161986b62e678b5a4df93ff93b18cd1c2ef230ba35c0f8e515ebb3d153338aeecb599bf8b8c6
z4bef7682341c6559964f83134d4aebf3fea06181752db4364cf214703812bc2314debea728cd94
zc9cd12faaea8905d76f78ff41c7c55f4d3eaa1f62f5f106a26465f308d8abcbbc939c9aeab1096
z92a88f0a6118a0e80b8520e7190280ebe9f9ca140c73534f0c2b11322dbd4e1395a3e210e3e825
z40c6ecb647ebdce235211c2c400483e6c3e9cea17b349d7f0b3da6117ea26de5de6d66de4f2b3e
z47f8f562313fdc4bce499f0ddb18e02931999dace2c09749a1b84323c6c7b6b702f68b71271365
z7d8cd3b4a2dc2b2ca5d7d746390719ff4ea1b41da6392788a2c484c82a2425e58f6bd2e7956cf7
z7a532536d491937ee692f0a1c2a7c4aedce2b2a6fad6c13e94acf628908a7ebc2177a45258e06d
zb4279f908b85379feda0fce6074d86845aa26a57183fb55dbd181b88ab6d1e318da04ea09ce777
ze73dbf0a4b74432a51b912c04fbe0e599af43f4079e371da186a45ce572d69b4da1e6b92a33931
z3103ad3614a23590d6b8d727aac198be1d40494b352ddd14faaa8af32d55caaf09ae69a63b7352
zf266bf456fd596a79d088705298502635f39d737167d5d9a97443ffc3a8288395c8deb447937e5
z6b0f6478617718585bef8e563b50bfc291dcf52f8e4ab8fd23a0fd0b5b8beac984b554e6fdd80f
zfcb5e1fd1157a26e0f54d0ab411b7f4e71f64f75bf86215bc349f8772c113dcd33e292df87fee1
z4a2f7b544a5bb5f57d64a70d9ea2cf5fd3c3a5163cef536f3c9ff963aa8390f71c9dc68cf6231c
z1d4d40a58e26b5ca3ab9b2c6e916d5aa2413a114baeabbdb36d1b47e3b1eed1877e2efe38fd1d9
z913a4493dfd64ebb5dd5c1d43732dadddf00e535da288d8d097a3570698cbdcaa83dedf62ecf3b
zdcea22cdd450b8f0a39d10f402ab6a1a7650bc841e311da761ea032acd892b8088584cda882300
zc9ca5432a0eca5d3bf300ab40514b1134335d5b1fb1acc5c68b623fec5192ad232fa6ec555e020
z62e48d8329960be013c299ef9570a6cb42c8b61496b41d55715806080c6d69601067bf6d7f2838
z38b3b88d55a14ad2a24febecfb003921c11d4175888c32b70a54ffeb4aab65eeb510bdba81b4f4
z911ec73f19c14c714dc7ede21bcae7264661a34e97a32f972e2ef35aa90e45672bf23fbd3fb042
z850260fd60c304edc53a3965980b5061494cfcdfb3b124831e2288812073e8224da247106c85aa
z34f13c685277c709ef69ca1b8c908cd0b0ff48a4586bad5a011d7d14cb4cceea1efe710485ff7c
ze1ef4922b70da0134c04a04e02d4a98ebfc0536024c22c87de7e9b16ba18fd60f648685ccb7606
zc6dd304aaf10106f36df8517743048561db316d4d6f5aeb741a6ebdf00aaecc592a85b8ffbf42b
zc2f3202379956b188afaf380ee6304e0430310107e29819f0abeb479749e2778f0c000d971277d
z817f44aaa136e158376f6473abad1670c5f99fbfe509a70c1f7121559cde2a3a8c7afbe3ec1939
z5d4744a5fa54b2bd2bd7a48b22cb0edc54808a6a73a8b87a8a06682c4380331b3b7109897b5f38
za44ac0f919a65ad6ef345f95758663c15f8913d96e7c0c4711a20116c29bc8a5aff81bb3ea27a7
z2c5e3adf85a3c4086e28c9c3da81e13451c42c0556e720114168ef87e3c4598d8c00ee93d1e94f
z1c42776be7aaeba34af431fdc9c1c466c0f22be1bdd982461e0bbcef24c41fcb72a1c65ca95b94
z37362c96d67e3b160f6fd3d6a2073140a454b99aceaf6c2789780acb4b856c967d6a63c2db3413
z5b788ab2be31c65f085d5a03fa0b44ef555dad36830eec60b14c8b482703b4f10e46572bce5f9f
z6da5eb54a71999abad6f86f67aa28f85c9d0488ec87137adacc79a1594fff9e3f2d8ec014d4d90
zdb3c5997bb3b7191f4af2d078dcef5d7aff0a7c2a5530fd3037e690c1a2c0a302592101de00590
z538e309e5d28523b1d00984b76f20aeaa92acc8ac7fc107ce99e21efe73a64b568c5d43b79aa26
z80d51318848dc243abd8ff311e9167336b744e9dd319ebe2af70f1d20853b92c56bc37411aaebc
z8f6f9c037803ac700cf5e36a1991151bcac210200e3a5bf82b46b08580e56022a5767813381a10
z2b2e7465461b3803af1b20b465f183f04189db3b119b77dd51f5e6643482888536b5d51e29315d
zb0294595f900af839799dab1ce2e0861c8934e2068a993a31f872b9eb39b261e0ad4a1d0119e43
zc2e9e466c6ad7e7fe936f121a8ea7a6e52357fbab1723484f316ac79776fe3753b2bedb4f77963
zc82776b75b823e5dc132f5719909da1b833275dfd7dda6b1c1f4fd2877291b986679d8f4f6ab4d
z5b879624001848e87ba74d96ce70899177f8d9f73037e656f79bd4209505759fcccde370b12927
z02e9499e93ea598248ea9881f7b73139ba3d07763f52cc97e6f3e5d1a1bdefadf6e488d4a6cf69
za23aa3c76a2e02fc8e7c3af73bb3374c9ea702825cf577268b240bd99c6901b1cafb4b01ffd20c
z423994984443e68445f69997b9c7bfdf761527f2555e40ff947c2f44540de929d3881eaa1b9eae
z78cb7cd8fd958333f082939821812bf395ab1490c91f84a47d111138ae0d29947018ed49356ca5
z90a47df8799e1434303a56418104c6049c3a36b157e270050ebc491af290ead231bc1298287a5e
z16e1ecc38086ba353b97f1473c9388d58aaafc312d96214ef543f6759f514e836f8590dfcc3742
z5f553ac792713728edf4415249eea5b8d0115bf633d8c30ce577448e9c0a47e57284d13bce3b92
z730c48e1a69afc6d9aa931570210ba5863861dab510751328fb5a2dc54c4136b79678456f040d0
z2cdf082b27271edc66bc13017641a187fd0da0d2b20becae4e0119ca54e28ea952acb35172de49
z435e2fc066c2e70810d29edc24332511d00bb2db2c085393a5f9230ba6f11936f750f7801f2a6f
z1cd6b60305a5f76e08ba29f55a0c8be6d381e16cc3be9ff363ae9acefad0c0a7ee33a61314ea18
z9d9698a4140e51f11a0fb643611e0780ee714a0862b7d4ba1a14600e93e3663e435caa98d3bda5
zaaa777a9f5df39eb6160819232704d4dd6225386d14e8971f9170d6989f6feff2af58fcf4e15e9
z6c823ef3989e03cd7c767eb9326acca5472a52ac1869db3a91066b3598211b2ef70db820894c85
z8529f6df846f857613747dab12e4a3cdec82d8247d6f7ec26bd7082848542e9e2042e2bd97269f
z0ab9dcbc54c29922a8c3104f8c3c59ebc93a4b35eb65028bbdce5d03ebd0b7e66ec183ec5cefbd
z0b9ccbb95ed8e269bff7e1cdd259c5746fee86ccca979c44c263ad3caa2dbe53e244e2d93b481d
z0188af61c3a79c0e6f43a2b2376152c933006afb3cc900c9c203bd29a1465f0e7a4b9568e01353
z70734afaf3fb610e934f724243e5d1c923f59e507f5718da7426ded2c38d5af652b395cff4b298
zc0cd2d89e8a8d20beaaa4e4084abc2f22fcad02d92bc374b1ae73a6d8ebfe07fda27e38ff98dfd
zaf28f5a99eebd0d71d892d684d2538a7888371f96bd69ec821cfa768ec75c7f06b282f7b7e7477
zee1afb95dd26662c8d5f8a93403952ad21b01886ec107ee70a50da7f80ebea7508342b0e2d2413
zbb6462f9a6d334d56f4d007d7fdc12a5ecb5eff510dfc604db69d8aa170c6fb51a9e24d5478191
z5f38122375416e1f1f05ce17cd7bf5b8fc6b7a2e70cf549a7818d835425b94ce7050c6ede4b8ef
zf39e26cd036b55aada3191d5706c087a12af65f31e2f205189d8fe210e816ac5ecd6b86d66cd6b
zb9d71fa08a74ae70c031e77ad9f6410eff60fb9731821926889da4322061679c989c907773d190
zb9cbc4c65d1372745359f4457cbb2661b621c99f198fe800904296428ccd267907a206db6aa742
z78aaaad40a37e53d7872884f4618fdc5ac2a437c481d79aa8f814e5d81e7cbbce9fb5306700801
z75db3a83782ea945337410f3f93c1aa647bdc12383de7d82f8533e9eea8b50a132560e890a5914
z887f2a22242f0e1a250cdcb2305a88e92c3d2fa0528d7a4f2581c662eca2de8d25ad17c8e06740
z442cab8dd642db888dc1da3127b64dec4a683642c6ca57bf49ffc8139f4efadc2cc3e3b775040c
z3253f2b4c80569043f90c95522db2468cb7ca2317f2654c719a88f11a9979041a468962fb42686
zdfd3a183f860bacb5c35ce565539fcc2a9759fcd14856d8aeabff5adf494fcc271855926dda7ca
zbc7e7050f0cd817474697623f20ba4dfd9a0d17b668ecf08020f3f0e12845571d067064728e0e7
z64d7c0a5938a040d02039a5829c368902379be4c88240483595d6f866fb03882dce7a49c7f24e4
z3ef76c0036ef01cf26be57fef6b1be48e09c5cf749d1ac1ec1371e300efd25e514f98566b21c54
zc1285fa3193da511a64e4d08bd3ebc7fea5155d0a51ed19ebe5c97b4cfa3f3b5c28d0a65564fff
z05cad7275f0c9b66a590bc635b96ed3cdac6f61294cc4d3a6f4cebfb62056721a931e037ca95d1
zbbe1d87b1124ca1c2bf7a44bd51f0f89c89b12eb9d5b571632603b2222d4e9788193c3aedab204
z8d9ca1c4cc8e654b47d540419273a1dd2dfa3b7e617b396ed6ed1fd4a607cffb033b334c53af73
z7086ba8833c7b683135e0f62dc268d629b920f6ea2af8868d73018f782a129740ffa1ddddef8e9
z7c16534b63f7eafec072f10ad120d4ecd7e1053a8b323c450e255ddae906b8153917849bb45ee8
z606ae51624fec00387280aff65f9d39d6c697664dbbaf9714ff2fcd6d1bf1ecb28270ee800c08b
zb143e66b6f682a78c5f5bdf5f6333aa1c204a106e1f7400eccd0e603c7f6e268365de16c0f4f8d
zf39a7ae2460bb2dc08336568bafc7d53926140f229c4ace7f470a9abf47e3efe357b2716745865
z19b9fcdaee9c89075bb5fd8be41dc00711c41b5a60aadffd52f0a9771d8b8f15d6478c61e6f810
z47acdcba25b06e743baac6bbeff0789953fa1a2cf883f289d42e8cc294cabf8b6086881b76b811
zc04938232b79fff9df5d64bb3dacbfc13151452e6c5fd3ed935bcee4c44d50f5c616e24d2d5b49
zb21abce6da62a442217decaea8b68227bd0a82c169297f1bc662e507b6b8b5edab8d67d651f1f2
z98091d337456ed4120abc386d1d3d3efcd0bf9855dab6f06203e123fb1b3e93b1985cdc786ba63
z6e9c5452d2ee513a9a042f091c56c0c4ecae22aa3817b270ee966175945d3bf5113db799d64bc9
z08c550952de2f61741de25aa2c45c6cd1064e3ec16120b20797e5d4ed58aacbead2f4e4d26ad28
z71330fff4f84e37acb30452acb5c4ab3902f130ab1d8a4a9a84dab5ae313b88d7384c84cc86cc3
zbbace8769b4fde824c01585ce567499d718bfacc7ef132d877b9c73f30935473ad2d1a9c6bae3f
zd87a51ace33a1482105f8c6d8bd1a72b39153101b2e1ffad470ab48213ae80d951db74a09b0a92
z6f5431d46acb0ea0cbebe7f63362136884b45ce52f90bc4d61ce81fe98b35b67be9d7684988665
z1464f3ac301792a0896194490282cd09329d73aa454a31fba0db20da1d077289571a0717d5b223
z1bbb67d6d536fe4a216518da6056a686e5b02fe76d8ef2fde9b34cc9b0d0bab26c719f015ca49c
z079be34f39508187625c088d35737663d228169a7d15d9f58855950da00c2f544a91bc25198cae
z7ff26fe98c185d14f10209fade3c736d3063482dc7dbcbb9cb36af2bf115f31ffc66de3c3ee4f9
ze3a860e6f1f102547f31af2433442ea8f125b7fab8d9416daf9c6edbbf34bba435f94ee3c2e33e
zd09220decc078160b2d69eb1b066e29f65b53c526781a70909274172c9abab7021ff7015305d8c
z8926d57ff493b51b32f06c684124c72dc8ae3cee6b0bd58feaa61c545f2db03c928c288a5bdead
za2c0f7026bb86555bb843801a39437667af5aab2cffb8216f1c93c4fdfb0d35976d4d999f5c147
z0a8102e207cc9c34b410026b1f9f493ac62679aacff2f9e3d5740d5dbd77dcf55f627dd157121f
z6421bb8cd8a2a9f166edd7f4dee79e7debc60380fd28783d957de7624a4e04fc2862db1ef4fe6c
zf662fdb294eb0dde8d226fdc97f0aa8a64e3892033f8bf63888c3958849d1727a7a6ae7cf7b80e
zab03240dc00b8152c752496a63e277d4b00a1e40e52dcb1d609a1867b2ad0e0d0e6cadf9296910
z2d19b0cf2b88b91a146f14063667da588fbf48276a4ce11a3f2e918f5fc9973921090618cf3f9e
zffb12d66779de65edda0d347be564d4684be610fd26e607ecd2e2b232064ed6a247f1f6f615da9
zcb5ac5adcab6a5b66c9bec5f7783407b48e7593736542307b5a4d09b2dc123d519a9b880f861b2
zf46d8641e0d34ae36584ff41ecbe2973203d9e25bac8ecbb3e1fb2370cca2547efa73239239025
ze8f3def4143d45f048ef749b3d6cc1141e91c55c83ed13dbecb650875044e8a6a1de39d1ca6486
z8104e06d0924076191dfa44e316ec35bb252d7312439781e6290c7d33134e7f0d7d09039a52d07
z9dfd117b49107c871d059b0704b6edc13e184dca14861575fe52b42ebc03f48e68fbb11c8f0631
za567001306fe2911c9750e3a8a995f6484713cf9b84946ca9d18c8deb711856ad27883ccd5c021
z5dadadef66b752fd2f1367edfdae0ed82482a81410b756889f751d5546f3174b7950f532d6766a
z51d6fe1744e1a8c389d31a146aea990770a39b84fe09027393107840df78597bd4f62a34c6eed8
z076938006dc2e2a66da64027ad8d7d97d855c33e72d001ac29c7c9ef5d5184a3c71f03c667e50f
z458bbb14c6d4862a285ea949cab56916ccf8929970d3be00fb80136a45cae1e4be6944f18d1d0a
z5c4d7bae567c2e2741c92d3aff1aaf893a86c17f49150ae95aac1b61c2e482fccc3bc81049a7cf
z7ba2a4a6727145a43fac755c46f36ece71919b4547431a14be66ea39dfdab7c8847771b10ba6ce
z4d1eeb6445023b149a8b9c1ae3d29b8314b7988cf927d3ec6038443849215ab5189fbfdf3480c4
z3e77c520fd1704b191302c6017206e5d7b2608cf0f7b7c20082d1db0c4a013f4af139a13725d48
z5af51969fb2cd9f28e7d8e533e5c8af45c4df362197d778d6eab21904ae05ce21baec7134c55c5
zd4579ac1935d5b04c3daa5abd7a00b74a4ed32494a20321e2110b4d1e95c16c2b764ab6ed01d7f
z3c2462ebd7ccb757a252e0f98c2bf81527e452ce483c722a9ff7d55a45d05aa9cd8d0d822eeb19
z23d30d89094670a2b48d8701012467ccb97702a6f5a3f6cc25fadda713e48353f2169fc5152955
z2acac8cbdb9f3f76208cebb92444deb3b9f5a0207bfa956b55ddf7676e70e92639c301fe5a0d8a
z612e213c511f340888a3850a7526a1b1d4c67fc7d70ce776ce8b145b95496cf818394b110ff62a
z4d2ccc9c400c6d43386d18e364720e4d89c9b258210af64d05735d9a5b54d49f53b113d238ae1b
z673e0065fb6e4d46fa98b9e136dcba9e2568da09cc60b296d10d1f7f571f95a588e756fd693b61
z87ef9c0cca739ffb30d85919308e4167f6d7b014dc93e28bd8e3455d388230bd148b7fb564d3ab
z47c746c381c3412025fe757746fa455da6430dc9fb3462ee0a797c0d75d683bf83ae34607c5554
z009f77b3fc88101b1dd8d1e39e47ebecc231830571c28d093414564bff6d18d0d1a7cf0bc1bb91
z91045cba623f100bf116064fc36c858fab323d325d00c4b0bf1dfed998d37c90ef917b648ce41e
z42cc23fa636b6ec7da5aa44cfef804fd08ea774ea21473eec5a52f702b0f27895d7f01995ca399
zb73c6d092e88d53e7eaea57fbc7b64d57bab993b7ca3a70244f022d3f98c55bc825021b721aaed
z2967afd3b117b2384d6b9e727a0d797bb2ebed1fc0716e90e186dbabb020b743c33d4c316cafc9
z9cd5e1c68149cdc73287fb584b1a41e2afc3b986531edb7010ca120320240bc5a9f8aefe6c54ea
zfd22b7d7a8a3cdb4e73afee6ef990032006e7d63e465ea6fd0c28407b71b34a62906035e4de1fc
za63c3d8cc5a7be613699218d735bf99ee9efed57b1cd21c206c82e79f4f6449cd8b1caf9a8df1b
z6ed3974c17cecceadaff1b8dff8e4e56af88afba6a74c256368193edd76e0a356dac13881b2980
z20dc60bbc4dc9bc0f826387ae468b7171bf301c8a9e7bd2b67d9e22a12b96040357825d25e3e63
z53cbff1b062333cfa61a3531f24752310651055cf96139b0fac3f004ff59703bb25c2922ce9dd5
zf4e4f6b0d636b7b0426ada1f74c8433169d722d2aba7d1fa630649fcbd038e2432782f19b99bcd
z91f45597c82e105a4a31663972bcd96c3b936ef3699dd19348c67632f5772bebbe668fb2db8d0d
zf3deb90da8d3e9c3e5e8bf90868a6dc523911e373576484edcf830beb679c8a126ed230dd6a431
zb49fef5dfacaa0b18fd6899281cb6d85c5987365c90b9b6c28803a94427d3559cc658d4af5f82a
zc48fa7019f279d292c04ed2954262bb10ecf3d43a018814322eac4e302f34dbc1c441d1e4f09ec
z7de3993e2db71744da2b12fce97acf935592659d6546a20c94550b56750b2825220a19dfd67890
ze6af5fbe4297b86e620aaf9881b00348c1f70f3da06a0d9240c5418732dfb2ebf2fc54233a137a
zb3ba914801a290e8b0acd085fd1991ad4a50548f0f8b19b7178e515b674c327f6cc33fd629b1b7
zc29e78036982854ac542bf3e20d6909bd048a75a0c08ac60004df200095c0bf946f513c6836681
z26a33baa60449ea9aa48e5409ff0aecf64b89926b9322054ffa29f0c1a8ef662d7fcb29a52b24f
za9f00786ce3555badf0b80446dde00defffaacd70cd9f77602361b587aaea8fe3ac1d479cd037e
z4bd0b0f0306ae431cafa33bebdc9fd64617bf3cd60d7601d21b71578fc4f328db69e248e21da4a
z4d8881fef17ac52a4f5eb334ef5ed07cd500f1f9e31b7b66b3ccf93567ef25580904d69b05824e
z2a528ba50c69b7a15ea99d4d79757fed67979da8e09b3ab8a835b5e05449e6d04fb3f1bd4ae732
z22b0dae3300caedf7fa8a39028378a8d74fb01a6264afdfc20af816ec4130f54042337ead0cc10
z0c7b8ebdc1c3181f8c9c0b5298a0f944f0e1e078553f35fbe47feffbcbf4cbecc687e37a6ea63c
zb894e0e49da84c136a4e2092f693defeb4e1dd74f4da844be09069c4a17545ea270f0f8aafeb9f
zb502724fc3db1beb4e5634d4ef45ab88fad68f3ace265ea17568364ec1b6bf204689dee27d9bd4
zb919d14b96c4c8aec92f66b675207f73c364c22b863dc57a5d815d849b6bf759b78b6769e7a6d8
z0d5ca5e3d7eab117dea5a99bf81c4e3a5fa29b579d2be464270cdb18f1bed9947b0297060b135d
ze28c5637fc9d673e4d90a9022e9736c17cd8abf93ede023f30c2d1235e4b049e780902a3a81b7c
ze0ad6e0bbb8f15562aaf2d44e5d2330900285e3fe2a3109fee3c15bc4ed0d881c559a92c9db592
z8266cc8c138f4754afd1fb2eb52f489df8ce0daa1310c37c324c5f4ef21fad7cd9f93d92ef795a
z32619df1320c31f74f134191a7e0658a58fb524989f45799695d88a9d04d91e7c0473271cee8a3
zf6f266c6d1fd7e93f28ed38c584acf6caff74b50d539dcacef97fe6570a7d7dfac8fdc5e46a433
z399fab5acf68736dcd14efa6da7b0b6794441f26c8429bcfe430be13cf6bc1ce0191de0657d947
z8824b5d0d57e017d47f86a9625d2f4703b5b579a518d5d29dae12a64db7f998e9424fbb4d04101
z3da44add6f2805dc847f62440744b4adb04ee3cf8d2dca19f47ecc9430e98b2fc44d1897034bba
z16afaf52df3b5beb065e9d79e191b104377d795e507542b733a534cce4a53cdbb31a038afd768f
z4ebd912419c7330bb6aa6be4a623752f18edc413f389d6e4083fc2866f1555b7ec58f7921eb0fd
z762599aeca5a6f158da2531150504d75e54646de73586646430a034374495dffb019e67700fbda
z3a03b96786c7fa545077ec1a6e4fbb1dd8f3561eda1f370cf76ebe082fbf33b8e6630f223a037b
zf47648344ed70d9ddd79c62ad148b5c48f681e289b1f03f62b6bd711496d8b9d9ddfbb69a873fa
z5b732527460025a235a5c8093a2de50463ef6bd3eac946382d4a12e92315f598cb8850a4c33a8b
z5fb5a1ec5afcbd59a3f4d26461c012648746afac494b5d3c7f184f6e9589c3c67bffc453d412a1
zb58d5101a968adfeaed0b810d5a06c2fed0dce941df1da868f1f7645f600b2a9345f507e103a9d
z8f1c6a4381cc7edd2a6f1f4df65641adcd784a0f0c9de876c49d2447f270b09b13f53b4e111641
z78ebf4733849afc1e72e5d9956183adeca1ed0b999821bac9593acc1559b509d37a9399684ea3c
z4863fbfa94a9aca6c2342250cdb82ee9a40d33d425b908b342fa4d1d882788d76028aa9f392708
z158b604045c92bc2577c91b94db4d9963a877a3486bd0e0b1089f5d2cf2e246e21a337c00201f2
zea40babc1f73ad487eafd6f3119208277eadd39625df39c180a81264740f6edba3890870af5b22
zd2a4c8b85f1cdd3deb0e8cbd586a1aeb10f7d8801cd384a01d8dd9e758ea56c2811330c83f2a08
z299410aeb98a6867d296a745491d70c38c90edb24b312294dd2ddbdfbba0138a64fa56caf0129a
z1dab017202f7c09aa502b594f2001bd0eef8fdd4e9a9f788b4ebb78368b9b19f29875d37617fd9
zf51397cdb58df1a08c7c97f591fb62345d40190e62dc3973617b3edab839fe2f019ea590304bc7
zf08149addf083c65ee93ae349bbeb99e1a8bafa0f1a19419744674e9e626e28db1803ffa07deaa
z7732e9353c6fab37f621800f149349e0d7850e464d5ba8097305d21d71af3b92c0e990f2b249f7
z4d28a3ecd27cd2c08f79861efeb36c0a1558ee2c89944c6dcfb8f0ad67f86af9608f74edb49416
z503f495719fd29fcc2d7c9f9e732bbec1432c71a34a16bb8433e80831ab2c105c678dcc777ca71
z8dd71ecc83596ebee4e0f99bc05076a6e9b2adbb81b430a80d0de6d5c5ddf5b226fe5bde4bf81f
ze24a44832f7deea096b9615686b134eda25f103b592cc10b8ba8f30e21ef6418ee64030fe04a41
z9bf5d66df22ae53f47dbd12c2f9b08a6853d5add5d225b224814040e9261b501f531a7282ef0f7
z04e80971c7bbb5f05d7668c19a985528fb6faeb2f8ecbaab0355c8af35d50f986db0d605911b76
z490088d2c0700a28a2f24a754fd65690a675908592b85ced21f80e2fee191b97791a2b8de4be63
za72da9af4d6c72d33b71a3a3e0dfc3c37f148a2fa293d0f18ed1fb3817827dfde92e09b3ef7c94
z6f304825f7b6ef72ec721fca6d9208df5e6f80e81a593a631a474dfaddb62857d001b50395e13f
z0f1521ca8261c00107260660e25cc356187821d28bde0f9e8402c2be83444123940fa71c5ef4d2
zf75b300ea0ad2e01d7c7b20bd6874e4ebcb61fbfeb7e92fa445e348cc2c3f394b9ada2d2ae34f5
zbb91fa94346d35efc260525f57134e1c250ff8b006ea9d5bbd2bd9a76aa18e30ba148f251bf8e0
z3f1b08ed622902a054f8a400e005083ae0dca95b9f8a70b2dae623e53504f5c60d968366b5a32d
z56ab4fd23a22bd59a698046eb90040d5c60d3b68ee2ca8b28e0561e4ed2893935d02a61fb1f243
z020de52ddc0ac9caf3e501fba64058a2c67689c79acb5c870bb43f8db03e2e94523482224477ba
zc24664b3a1dfa960ee2dc03af9e8a9d507bbc20d1eda4a1055999e2234b7ad0bea28d50a0bde46
zef3067a52f4ea3df75dedb303d9de1b6eaba141258331459738f0fb9729aaf6e976ecde89b7fa3
zcf1dfd4338a2437e5a53f0b25d76b06cce9c3b5690010caa66649988246987ac2c4b7687e3c9d8
zc5f6fa1c697af46faf46fe6eac864d9af1cd2d642af30287d67ef24128ab8a8f59d196d74ef6b5
z0c8b68ad9095a6787a58dd101aa0dbd6360507365d399662e60599e030d323057423b4f696d415
zd56f736bda25205a065ec147507fa4ef4a26c07b57830e816c667eda763a37da87e5ad42359537
z2342e3f802e08723b728d2102e618075472b39e3d16a93b1edcd22d23c123b74eafad4097edb7b
z7f19b58c58a18301c78e25701c7c9efa09142a77e9481ef10ba13ae20ecaf59d82feb949cbccd8
zd82fdaab06a5975af88272ba32d75597cce58d8cb934bc8033a0aaafbb1ccf29990dd59a11ecd2
zfb5ded8c69fef6bf31a24a66105f8bb5a37a32d6ad5d1b2dbb3ddffce3ec0b46402f2a2a9ff49b
z208815a59fea138c0cc4d29956ffde86d752464fc3448963a529472aafae2beedf8d361e5a0280
z5af938d09747851039b3b1d2dfe5362d86c05d4c2bc77fc818d47628ecfc56cca25f27e7997e1a
z7a3c6d527d393daa83afa570712743279dd0c361ba8d023786708210a2e13cf7bc988ddb337cf8
zc804b34c8e42b5f0507fc906e7fd671dc7ddd0e6c59727af417b68f229e953b5b9631cb696d9b8
z061894da2bfb5acf676e1676c1829b7c980ab85f908e6a25a0b34897a52790d9a3dcde6c31044e
zc98be11394ff4d9f02b44215f217c4835abdff37633bd96ab7aa934f10052aa0759e44020a240a
zd48ee272939551d484296b1363f89990061a67bcd92fbba0f7fb5aabddda8b82766860d087c8b2
zaf47f88181fb3ce1c626f952aaad9e87c0ad1c8d43c6ff66d76aa7a6113e9fb0f5f315f63b6e7f
zd97760fe7149d8ce2c41ef4221352704dd0869c4e91b49842d94a3b47ad3e528b1295f2e1cc4a7
z1e37e00b327aebc9a7be9e40b6de975fa3b5a09114b1b611d96db781f688852c1071bd931ebc7b
z60763f3bde41ef404d26d665bea1731b5dc9247a7944aca9e86a1c9b8aa544b5158009abe84db9
z8e5d296eddcb14dc7d8254d3e41a6fb8f528e7bee4e13ca87451dc6189f4714971a2ed22ed7243
z8fd8adc66cffb446245b28db52ed64cddf93a8dc424d2c41b0fe5f0e9d5f5d4eeddc45d0dd6982
zeced54c12b113b836bed8b8a4ef70673313d92b27d69ffa75ebe7872438145c1ab1adc5a83f517
z699eda31a25c95bd9267a32b6c51ae52cb494ccde7f464c36a0f0b9409754c00a91a0d7208fb0e
zaf082ad2e0f1ac65ad114caf8755d1fd637ea991395d84244e2db8d76c4068b89027f8ebfa21b6
zcf0f744adb48efdb66502ac2058ec388b98abaa78ee3f2ae6b803ddf614fc120041306cfaaae06
ze788081cd2e71e07a12dfba162a0689baa4c08fa77771af6ad78d83162002e26af416250064874
z44fe9065b6be11250b4a0b6d18351529ca726844ad82e3720bf9ad4395e3ebf124089fc7348240
z6c8b3db8d77300ddea0e3882eca5c53fe6d4304569c6e69401a85d743564e8df693b0e5c60e19b
z4f888f7a09c31f62a7a28aae4274890e10f8b384a15d8c5077271892671eef07afbfb5110c58b6
zeea2df06372f926154644c5955bdc4e9d41345dcdc1038cef475ceb30c2a957c85bcee827043a9
z51137151232ec53dae71f00851797d0f0f102fab6ed514b81fac09a53039d9d765921354dddd8a
z125bf0e90db0e18b9cd40abc306ea1f0f093c6508d08217df63ccd31cf3012796070693c5da312
z260bbe41f876935afa93cb68e30a1b141c4938cac976bbd2932e60b23e6a447e664eaed0233d26
zc139ffc4db1576c56e5adbc60411304fcfce2adb8b96d22d4b4a4fa5b58d95227d8a2b4f277f1a
z6f1b33791a3891e8e1935bec9ba554a3f66b52959afb988f20973ea53f887d7e30504e7088be40
zec3f297575a52fe28c2d27fad65cfe71685603279e42b228bd65d37acffd4c0562b8c5328277a8
z3aa77722afe98ee1b108fb1f1c1615f2853661e93abbcceadeea7a5ed1a6ea4b165a229e0df261
z319b3da17f2bb1de10d178b4c6704aaf7c01f4e411af675f337ff2b129b43daf5eaad5c2730b90
z9f031ea1559fb859d43e2f0b579d2378dfd476d7cf31247948a22f6a144d04e636cc475a896533
zcf2a694dfddca78238b9d904ddb9293d35fa86bcf5d68fa81bfde767058c00f9c4e67adf01d433
z1b6cd6d15a674ebcaa5d71bf2c6d720d03e9cf2e5cd60ef6b1f5b50f744069ca54b155692f3e5a
z323bb1810d78de5806e52887fa1269618ae09174621b0292b0167af6ec66b502222e8624c622e0
z17d38fd2e7b512f154805c4a1e903a3cfcdf45769bd005b71719f37bcd2d8e9aad2dd99f457fd8
z2b05db571ae768c20894d4cbeb25891eadfb79dd398843ff9a0f7dd5458f46d4c53edbde306cd4
ze617a157cf4410ef92bdfe5523c4948ae882495c37f054b8e80a4f29d4d2c3269cf646c0c7c7ee
z2a259bb08eb1cfb236b5efbcee7b080d083725359c7ee7971759149e14b3b6e9c4066bf2de61f4
z62ef298fe4d2a57f6faf678f49471facb0b854d270f1d3e84fae9b7e9502ee40fcc6cdf4b0c946
zd39b360a9961d0d0b859397cd2c5c9aa13073c725ffc2fe16225055829f387c50f52b6a0e32373
z0c4dd962ba3086d71c6d8350d76fd24a265358aa1d652425b35be81ae131e55bea3ae4abafe35a
z9e2884dc8d9834b13ef89f18cbf9d0ddde9b2681ccd91a37bc8241e2efa14ebee61e2670b3d279
z49d8b98a87e74528b92a3197d4795ef5d7eaa06514d35ff35e5fb089395884a369cf51317c80b3
z51f22d95cd11c459ec7cb90d87ac1d960ecd74e19d7a9a0388b8c52908bcdc3862547d4f3a0440
z234221923029b635eeb85a949af11a95d6f3524bd39cd2d0fde868b13a63c2efde0b8b6d7671d4
z5c3838f7d0b0341ab2f2258dfc85b4694c03f462e0f5bfcd25fed475f40c20cbff837ab52e8c17
zbe1f3874f4b4139b06fcbf548ae5a002bddb38ac4dffa960a7b23e626f97497fbe3c251e11167e
z010479b879185ddab55da318bd79dfcdc49f6508986a5822f9d6865e594f7eda8fe1ca76ee6efe
z45020d3d0b44a8fa4a793cf43afb3f3943674a5b29a225b4520172c5027c8d3cee1ecc3ddf9a0c
z32572bd1cd73afd74fada4c348eb417275d6619929bb567175a7a57ad80b67e06dea9ac10abc64
z5ed2cc04fc0d8510eb350c6363be878d9535ffa33538b797a31c2ec449ce64f33ad2662c740ce9
z8d26fd69acb5a6cd16ab5183aef85fff88750b687708f498100b140a54c504b2463e63ef7e7d3c
zef9bb37049a5ae1e3c31bd58b87f448715928d3561527ed6323baeff0117f9db5ff3fa93e99a0f
zc9a30eacd1474b9b7a523cedde694c8d7749b146b698aee41b5fb4dd1febfb3164e1adef109b7e
z4deff875d39fc7069dd9fa7cdbe8aaa62e9f68336943a1b77d52dcbc88fc8596a85866224c7180
z191fab5fa7c9d8b1d3bee7c4cee63665d4afad2add787d8b76f4d3ab02fb210cff13c29c7938d9
zef0b4fea06248520a1a3b59085ab82f3256b498b310907484de49e2e132eeb83999fe2fdfb4368
z2d2687dcb3a132e18ad7445bb40c04f7242ed5ac7b60273af52e381968347218045e239e81b0bc
z9be8dc60c166fe19c8c417677d3c96a048e012b01875218d3948d37826cd76a66f72c338a884b1
zff6f93d00e6fb75b4553bcc488cf98274553d2dabebdfa5572271e93d13210e664d0988568bbfd
z5715b4a3603713f77f01431a79de9b94fed2602b87a8f1635dc5b938fbcd288dfa69bbe9f569c6
zd7d92ce9684119f275272ca44f0f181aa5554c0cab40c6e60c714830436af8112ca4d4867b4388
zc399e98cbbdee0b878f67e4bd49d611867d31acf41319811b4c8ae798b169e2a29eb44e779a7fc
zc88099a38790cf4cb02958833fec761a5b6d7846bf9ac392dd44a73e719e42269ca273f18dd443
zc790e312ca02954db5cd3f924d8de1dac609f62281cc54b7bcdbc447d980ffc22aa25f05415651
z803c06b2be564f74e14ceed5b9e1fbffd7b967816f0bab17008c0a5abb1d7c64d1eeaa4c96c477
zf10bc033df3caf81745888d857963a05a58c065a371377e8657e4aaed0b842fd525109929a33f2
z48c66c7a29f6ceb7965326d55a0f066af81b0720985b4b8ad4600a8e4dfa4e6acfb4e428f8575f
z6bcb1b91870b550b311f941cf91c2ff141e2904b231a1a4b50ff9e8ecb2e283d39a13916439fbc
z01c2f5d25a361c7894d59ee577cd785912af2b370c60c5ecd6622856bc37653172113a272ec8ec
zf4677eddfa4820bfd813866fa3e69612c0990a1002f263298aeebc3be51eabf66592c047527a7b
ze90268f03a5b0c7cf975c8f8d7cc577a7a26cd06cac10fdb2fe46b2fd4cbd1728ffc4bf2298709
z4d3cfe14e57a8174b8cf108bf47ca10be6cdd38b8f40e0746318100c1648e00a2db4d7654ab2bf
z35b4e92d6aa53f0f684f7e1d090ba1545911a81761b3518f2f8034008974dacdb41b5fbce19574
z57fa32cecd78c341d00efc2c81ff4b44a2c00c40ed34e326b704afac4ea77c70b36910e461d189
zda575f3ebe6b97e56d8a46f668a977c13a0c0b755a2ce76889b1afd8829864d0f068a12445bc61
zfaef1a384c80fd45dfeb41d7bd3b990fc463451e103386e220990af75c466198119433b17ba98a
zbb27d91c377f6f436bd1699ad46583805543fe6987f958cfc6d6245448dada6887bf3c70913544
z771f1b06437366afef76acbce43ef3ec2a4096dc0a228e6e0f5af3b5f5072214c6b018ff6adb75
zf5e563ff0eed72a43e56d9a7dc4616c4ab2e482dc880ead71f9be8e9073e957f7029643ed75fbc
z585b4ff6bfd0fe905e8dfbeb9b7405e7012d0f740352e2cd323bb32d6a7a1688e2cb669aa905d3
zcc3732951875df038a080f36595a6a47be6da40234be7b4c9a839a8fb5596e4b659fa1efa8a6d7
z404809c740b83a7be1a1116c4b547be62a793789a7451659c0149b5aa072d528cf98f4051c7aa6
z8a704dadbbfdcfdbf6adc557c6a4f80c04380c14a9882c0098c21af138493135068d8e758e4491
z67d6092bbe875364c7f0cc8a803f43db58fe69f7e0decdb5eff10da4a02c8c72242b2eb2706111
ze4b4a4cd568ea51ea59592ab638a3e934883d7f4a8326d1d173ffaed55f48740826f251c7f04d2
z546ada12bbf89bdb75a7e7dce44b9b83176060b954e8fb7bfde1caee12848068c69cd2dbcae9ec
z57e7af53b9d3118e04a442d1938c058000dd5368464aed4d61d072f458b66f5466e0fcd5d84006
z3a0b69f2dd3b1611e2a6845770264c0ffa06cf95725c3a544278bc367e4fcd7bde83eecfd42309
zd98ae575494bfdc93ddad54c884739f53f7373ede1dbb2b84134bf41748ee464e2f14972caff81
z0e0a317be30fed1edb3ecbc13a3329032df26a5fff50cf3fde3517db8f4db9680463d9e3be7eed
z164a053d6b73ce6ee14e0113a13c0708247dfa3b15e9084f9928689143e98aaa8f3e108c8b2b73
z927cb9de7718547193ce309ecd8b3726903445d8cd6902ea902656ec5e0577c832327c8f96e3c8
zf9b4c7bd3aa25d782b063d0043728f8c7552732c914174010c3fc664f9d2eb15a05ddcce33b0d4
z10f5935c73869f67e777d6200c611a1230306038557706c42110f4fe422ebfbc2f5a057523874a
zc28e2dd327045a7cd43919668c15eddabfe942e728c6441fc3f8a5afe9a63ab824a6076929fa8d
z2d22290f92c4ab89a79b5614761f0fb8cec24033d1ccdef9a5bc6f68adfc590094f980cd1e291e
z00913068d9331f8bbcb5da053611d57046edb8848fb8fee40a15e53a9b20543045fe9ef8e95d9a
z2cdeaa2d6203ae587aa142b2881b46284b91f381555980f1dc4cb91cb567aaab377daab653c73d
z9614e1185572b40d9ad4b2367138c1598b4f514c59b204a3edb68eaa3179ce15afdd3dd96fd7ad
zcfc6c312ca4d49744b23dbe6960d81d1138fd7181a3e869f81854042af9aad3715dc2923ec4188
zfdbbb0de1399519c89c22f76a671f6d057e5f63ebb625b7cb40b1341b8d6dcae256bd7f9eb89e7
zc13cc057dbfb26eaaa4d70b90b8300ad4571b3d947568544d9148fd83d5cd3c8622c5b2acc8d11
z59ca21b6363915917d861e6b3a332e262483c49a05fb0a5a7389b54793400cc88083ab8e2d61cd
z3f9ee6310d62a36d7fc4966469892623520bd8883d5d427c415082fb0e3b56ccbd8ef259a32288
zd15016929502dc70cbf066a328f567d376ac8eb7d3031dadb026d6326012119f938331694c7c83
z9667865c2f839206ce700d3ea671310b07700e3c33f010b86aef35cf2d07e56285f24f310a6968
za911647d3ee07d06f8ecd319aa7fdb44f7dd0e1424284610edd512a2a5239dac2b31f3edfc8ae7
zdcd182af83fb93218eae29cdc7bc7e10c38e7412d5da7b399de421a035029aedb53942d21cb89e
zc89f2ffee06fcd899a17f0ffa0db16994d4dd5c6cdf48b03b56bd069e6ea9e120504b18acf7300
ze155a477606c0d631a93487a61172b1832fcf558e0c74e47b8719291d01e9fb808ca29b68fa3ed
z616374c2a1cd3155a387b688ba6f42c70cd89b58376b849293169e530dda5072a9d753254675d2
zb0959c6f1081238bdc6466af807ceeb1ea099da10be1c8511d4284966a6c554ac5ca27e16a327c
z8e0ea92a53214c19b74314f898772e1d10731fa5cdce7ae9694718acf933208f8f54876c6be4dd
zb3a8c17b28c9a5a0ab9a545c87f8d44cf15c6afa311bbad3a2d9a0ae8ecd0d58add05f299bb9ac
zb9177784c31814652376a4d4a7c9be10d3c69bbcf390b3ca58581d2874dfe5c8eff3dfae641928
zaf82bc82472c587479a8732e915cdf2e17085207f07b3f73ff5628ab567d23b08e822b567c17ea
z62c41cfb03fc7ee5a919673d7039810f14f475ba1401a06f06ddbd3afafe717a50cf30851090ac
zd7c300e4407668188ba9f9c3efd34d39c7796f5f82bab3564193626307d950b4b0b961975a653e
z51e7656bd32249bcac9608aedf46358ca239f4363fbb970135b36c5f92b99bdd28675c6560c151
zb4084b3407d8fab880ca905c2bd3148d1131f6d33baab7a9aef64961c4f5d308cc4f63a54be0cf
z66fe1802698c1e5c24e0a9fb4b8a24e0e97584bb41627d0d824f858a8ff9089e8b041bf20486fd
z19b6650e791bef7e713b5e62be24c8b42a413c4d5108373c837b2481045fe1e32ac6d58a1dc37c
zb3aff02fd99bd66932791c9e10b6c725def659948e97a6695b611c8a53df37c4e84040d1c812d7
z9bc0e106644a0cc147727678bbf272e14b3d3a397422ca76e48c557b4a998010cbabe04f760683
z9fc0aa30796b9c6ad067ea56d0bdca0ccdc75ea451e7e0dc8b46dc2adb37619a3b6144ee6cc539
zc7f1b538a8893f787127443dfd47c71d64908d70926e10fa576acb788c6850b8ed03db644e773d
z36a23564a8c849fc9c1ff70d6d5ce13296567ef34a97da12bf22f356e8f8b68d5f0d62efe37ee4
zac150253eb0a4aa4d8cd40a14866fb494870fa86ea94b97f44e360f98ef33874edd0e3aebe10bc
zafca63f8a9f0860a20771c04968808200f15a49ca55f97ea52c7a7be0490062f808e62ab577dd9
zef1e5da92d1ce692b09035faf96bcaff9e3f7c5f87ef4d9dd31f7e7efbc86405a6351613a8a737
zf1039bff650c8448705f7163120e9799933eef0dd0c4060660718f899d07de5b6a9832bd20e9eb
z8716e9948334a0ffeb0ced5191d6d9eb4c5447bd27dc03709b9db0e471ad87acdc98466fe723e3
zf680743c3fbb8b6ca617c3c736c4cf2fbcce956a3d2366da84a77e3eada4a7fa93795eae28ad3f
z51b7cd0f3f3bddda9c89ba096928f9072eca52cadd310a91d31dc7179ff64fa931c3053820fed6
za336208905dee8cc18e3cd87d34082f5469bd6031767d49d21856f5860ca0a57e1b711ac945910
za5065abb65a87416b20b194f6d01c00ebe640a936c41d2cf86a22757ce0974fe3be4a0d1ab9751
z8d4dd926bde69e980aa066b6bb9a390492f99d81074443fc2d2f23bae85378d6c02112564478c8
zeb7a96d03be187be53021b1ff4aa48fc06e7c0fe909ac991695a08230cc5402551dba284e437ca
z38a7c8f24a505f1c5d70478cf7fdce98435ff2296585a113286416210ffc2fc6c1775a1c362123
zdd6d8ff888c9a6d6294a4f98ff48cfc4e80c6ab6fa23c2af904d8b8167d8665c167879e81008cb
za3f7393dcee78f7d24c76f09ccd9be550d9ab11810ce38ce92a11cf684fe9959037ab5d08555c2
za89f464c4ef8cf248154d84b2cfe114e9a0a3f2b229ef585a0d78f850ea2b796c1078e152237eb
z218c6b337368d2b6b8d7390b77a77cf93535c54ef2f23c0adb1417e9caa25558260dca03dcc251
z3d0a9dd0ff400d11d0753b8724416647bed79ce5a87e895c49f738f01fe22bddd5fe2b96f2d7d9
z7dd3c32b58ed9d5135f927a670328ea449e27b1b6a0069c0de83dfc606cdb50ed0ad970859672b
z82a1da3d1efa8f4b073c3137db20826fb98bd4e27869dd7a17f3d13927dec346f78923a278f04d
z4271e40b4aacec3097d594b51f5cdc63d58fb753894d4f183c9ff658b75f2cad21b57783edfac4
z6c31639412a67903c1689ca4d9408ca8d659d9e9f89dfc43a4e1021486dd38c8475ca43b13e036
z3123e788994e83eab0be80c35ff077fc1112f47f9cfef7e956e40b4bda80bc7e0a88ef3def0a4e
z6097593f76b20f238633804a3fc7b62b300580cefa7eec34f731b3822f216df5c1d596a4b9044e
z18049a71b9d443616765b3d13abfd2e1baecae2a43573167a004470f0593726eda1cc4e8e195be
z639c6ffc92dfbc45ed3acb545334a13e0108f42cffd25b0e53d73017be4dc65e6fcafecc823c78
zcabee987e13a042b09256ba52e612b65978c23dfa054596230e020685d305d4c172b2ffff23273
zaacff987a787365127d01d6cbeaaf60e2017e9719d8365feb46f9b2c274302264e6ede76c09da2
zb76cdcf3adb4b1f502750ac7a7f2c2af908ee3d2f095d84e716d878bdb6b39e3646ca67ffbe2b0
z675651c11cf1a98450e550f76f4aea6b6526e2452f1cbbd5b8ba8e0cb5e8b75573d6ecd62c614a
z53951342164d4bdcd397f6f4677f7076d288fd323c5d4afef90884ba2a4f7a414d9bd43424b603
z2c0b0f9acd1de799fc8922c442244bf4238d11d13dc8f39ed816abb4d1c7cdf4dcfc3d0af10d4d
z18ccc4ca7862d097164f724bd4f8f58495d92a8dee572607a535154ba59c48158635026bdad0fb
z722125842e4fd283297ea889ab5f9cb5a40f28f5cd0c4cad400ff61617ee2f5cb7928db1767287
zbff6a04908d434fe8134a938b709ec79dc6c7fe98d8db77c6e55bde289f0ee3e43c6dfd3521c33
z4d3a0a6ac3b30631613e453987d3de0c8ee823aaf53d2691352ce803939c45d692fd86cd2ad95a
zcd7857b02ad3451c686f549e22fcbc878d7d845b1ea36464e577b766b3d2ab8984b141f69a55b9
z32e30b2665123ca7a2f5f53c0e2f781e3e415dad301ef1f33a03688a1d6be33aaa766a507ccfb0
z1b98cbf2ed12d87831ae96dc75d63e775da0e1b0d3993765a61a4a8bd06fc5da83ee2e2d4571dc
z29fb355ee44e92b79dc74ed355ce7c30eeb42ea867fdda622ae4d626e537162c562159aa3bee91
z4450f712453bf281ab961e50909c77c7712fe66d50a2020b7048c35a56e58a8e7b4357467ece21
zbe2beb8b5f7686a8318a3b4a4fa4a8a85e698781b8061eccbeedff1806d62dec0fff57a9036a3a
zb8af0061b6cfebf40d121bb3df38521a993cd46f6927177d7afa4894f2688ec4ee11f85527b3d6
z321f92423ed753457e70d1dbbb16dccf8825a849031a1b281127156c7f9e9d25f6d2b386a7ee91
zacda4700e77e7de3afff059e40fa0948a09aed5b203fb4e62eaa8e31069d826772df274118efdf
zb8a2051f5e0564bdc64214578e4f49b631b49e3db809444852c5f823f7d1052487792843637ef9
zc7f3ae8de7035e40fbf6543353b84c78f5aa71bc5468cb49d81bc6ac35dbe22dc552322bd9d5a2
z158b7fa48fdc483c690cd2639f6d7936559dbb3dba9490f40fbb378323ed05d013e80d2906424c
z570b658bee0913126426a24d94505eefd81d632ef7063731bd23c662a4e707a06f23b25673009b
zd3054ad4529527aac4a70cb55e1dcd1f24306aff7ec678688fcbc209998bc87bec1395a031e16d
z16ccb11e82d3e6bf2059f09d50384c96aea6a1e7fa749f58c79fb5bafdabe0bd058ed6f2b46e95
z345d422f90e3a573cf3c85b9bc8b096b982c07977759015fbf10833315f5fc51e4aca216f998a8
z63d1eddc8f38617899e0d2f0e7354781c6a62d773032b9997d597847e7cd26ab16c4e6d04db5d9
zc1e3fe24f78b8ea5e1361e6a1c5845b96d7abcd4def09a721e36a4276d161d332d7b99e21a0fea
z4f2aabf182d2ab0ead7c7010e3144548a3839f902bf33e55c839cc32e226f0a7c60c2f8f1335f1
z89e3fd609ee3cd75ad01d4e9884cf270233f3b145149781f6218bcdfb73a55b86764fdecb25ce1
z4ff39d8673d5277f5a1c0d32f97e69dca8970e049edff7f3409d95db9947d9c0647f30c2ef7df9
zfab36b125231d18a0939ca6df1e1cb40b2680e2924d43752fc2937edeba98bd6899b7e5c3d9cb4
zc4e09ad6b6194a7da2e9ab685b270db88fadd0c7ead01915fe463a688d11b7d1e0a770c5e12ec6
z3d4760053e2b269847398f397ac73f230e8b8c1a76f96b9ef10fdd66448be2704511f18a2aa564
z739377c5ee4b423194919d90a029e00c51af60fc84d08b4a37204cec5e5f4f756d2079b5954ec7
za6095f5fbec730867e1ffcc3cbdc08cdd0545354e3a15147e2214dbaa7dad95a33c5fe1552111c
z520e309f0d50ad511fb6d7c7b8a14e0c248825d5943471793d089ab932353a029c0d14f9dd3204
z43f496f0bd2541211b6847d39ba1bcb502306932596d3f2460e5f020e4fc26c324fb91cc7779f3
z4dbfafcf14591c6087d40253db4fc7e34228a771732d87abb68ecc44de32b2ac6a791f911ff92b
za9e1e1e90462dcb1b277983988ec5d8ea2e9ebf1af61238a5d55d6b79ba87e795287eaa9914b07
z511ad4c5a8f82119b1513829f733b02559c88926ec87959e090a5d79d28fcd2d91855db47e2fd8
z2c038a773a59cefde63234d7e8f4629dfdf3730cd95fe89c4939b79b9a0693b62c77a50c42062d
z31fd873ceed7f05c6adcfb94f7bd7a2d9ac7ca74c436891af5b779eaf029fc210528dc3b7f6831
z22c4f94323be770ceb165683453d99149b9d75611700993f8bdaa4412158a0c9f37bad078dbc90
zc7b4211cbf71512e17bdcce9b9e0f3b96ef6358ae38d2b35d39417ef7d661060d0a545d527c1c0
zf0fa4f1721b808e360a2e3a5c0fb54de100090939602e948bb2def318a63e35ac48a0fcdbbc06c
z3f72f99246e3b68bac3ca50896500a230b32723792835e122ca12305ddd446bcadef50008eed4f
zc934ae0d711580ea88028d7a98097bab29f5d24d5c56906c4a1d3b53593efa2d5619093c8caa67
z04097fb9c458113a444a17ea44502ccca099fe0669e57af1bd69ee2447b078dfe433aedb36d496
za63898db8eaaf01190b72c97a1a8278b5da02dee6901f26c281da797f6bed78c3a9de0d5a2b28f
z90911979eed598cfa3ebb5572e43c514e05b8b65097c3dd958365019da0ea141cc18c89b359b1c
z0cfa70a6e40444c81648d63c255be88dc5d7a13cec160ee351c50f821b7fa556e9f97d030c2e24
z96d1839c8f01f99caa625d5398014666d5d707973db428cf656b6f900d0e1c61e38532ab1699f5
z539a063853d3abdd5ad69501482a8d33fe0c5e3d1e3467c2491b216351d7f7f7d2006a51a6d0b0
zc599818a616e2825fa3a1fbfedc66b2b491f0cc7a4fef18fddd16415e53608f2f3deee5ba9f87b
z99d208fc97ad8521e3ec3ba525f0f0485f6ee3f77063dbf65a2a8df2da56cb86b03867a6d99253
zc2b1d0dc988a10ec8964cab903414891f5522747eaccda6ee025eae0875eec07361bc586ecd8e0
ze54ca95b3162cd93cfa991d215aae556f61368ecb9979ac74115f65565325e5edba3208616bc40
z05d80becc733258090a365acd99f94fe00e859a02e4fd82f540585c0add3b5bf959b457b41d147
z20517f8dc495228c260f55ef4ff590cf17663d7bd1977cb805b898e51c27b2b04be519dc7341db
zc1770557866569ebe4e0ce6668c784357f3168b984cdee3286ba7b06e1091ec81275877ad9e25e
z46f4c146d4071cb735c775fe5cceefb86b5927e009b2cbf0831db2f20dcea8f281f3258a8426fe
z520877e9e91db9b32be1b5d4826d5c903908cfcf200ac85b2e5f736a84685543b36da3ae5fcca3
zb30f11f95f6e0f8303b42b85971e647218ddb01aec11e9dbb0bac1be533fd12971c167b721b30a
z6f947cd8dd253f80b1a74160f1d9e2f3b072cbf7627c4b5ecfbdb5b6920a823e485c889e03ed2c
z7b6d78afa59b37496c6c6ee4d9f7342381c37b169a4da91f16cb6fad1002d4bcd1eae5883d21f4
zfcb56705955851d8c52ca369b69885d0bb380d027b17219f3ee0388ba144e90125e59bd4d7e683
ze35d874f8810c72dd4e55f8bd50d910483ca146029500cf9fce74aad5bfdcb5263a92c6138b7db
z44f388a6287ee70be5cb7133b8f0d86cc385b70f0b4f88e58bdc167beb068a44a75b46a227181a
zf8e226d8bbdb9dac08453172230c91ee704c70120dc2f0ccd5c6ee11837cb613c861b3ab955298
z3de8bef6155a59915d8f7a7682d726808da2c79e19d42342e48463d30d0c2f7173158e28e163dc
z30b973611ce366f57987b8a6e5bb21c23503afd5523b20d822e24889192ba491fd59c5d765b0e6
z80a31860e1f555b6c6637e0cf8f0bbb5b13701b43f32fa18ee5c9da3335398776ad4971ac9fa91
z37c5df0ee32dd3af7f24992ec6a954f5f8b29b89eb610c577bc10d4c8b91b09ba49d964b68d23f
z2d85d6073dcdeadd307ac445a5443267e988027e9f4556f16c87d7c1c5da9ff2e18788ee5b63aa
zac3ba9f1a4455aed876b5bae20b38f900a266cb7ff312fe745ae9def67076fe509a0003637f9d6
z0707e15621a241e32151c5574a5d9d441177e2428c376a9c9bfd12428a541da62b81008dcb4eda
z50a2afc3bd6f15c573679e1882ebf118ae32b1d70e59437686625971d6ad09078981fdac6184d0
z63361386c843d103ca89e71aac28ccd0178ebff3a915f4276997d5bb88a147e4f73cb69cc1e134
z9f74a02ed89a615ef78a4410d4ffa73d28ee9a20f8cb93077a227f027e919011fe311dce3d5b19
z91a948721d2ae91b86764518a6f5c09ebc394509fe073a9c6ac123eb2d869f7a397cfffdd2ed1d
za71e680a9d702c53ea454e79829932e337f80f0a94c8eedf7493791e2a8f36fd7dd646ac1f31f6
za2b6516b98cc529e885e1319ae97fba77140d4d7f34bd86f6bee6a56cac18d22f45282d3ab8609
z38ced17405ce616f0533f65ff0ba2eba9aeaaa105da1e933a437a865d9d59745c7870324083354
z1fc1dbbc0a450d4bc7bf2620d28fe2fab475c6cc1c3eac1ad75e0763d82aba4eeb7a6be157e958
zeac270bdc833d721ea077dc04702e780aa440563d1220adf679b22ddb9d243b8e9fd51511a42dd
zef484d7ce4f660dc557e3066013d6fae3f944a84fc688b27c8ab4dcd6f2e0fd88262d37ccc47d9
z5502deb2a442fd8ad82b53fbee6317c3bec484aa40e1c5f6de4681257ae703fb15b1fc84665e43
z2712ab54fec06860909020bf9df1e6b807df0224aafc74fca97c106ccc2ced2178e6efa0b09e50
zbbaa7c01ab98f80a9eb240c4df7f9b508f6f68d6a2139d0891902b2cb4c4eeb9024ca91df51535
za28813084e3039801b547b3f908fe282d3a780ef227432cfa405da437285add42c5de8eb410642
z166b91c237cff1b3ea182e552b3b6e2b5eeb5eaa294bccb344e917169c398d5a3b9d08df52a1af
zc6869e0f739473b5b5fd6d41c0e7b670a1c422286156fc5e47209a3441a33ef66f4e2706ea4d02
z1e9e79a933564ed354f75c95c1fbfe8200924055cefa3d5b8a1ab62b786f14688502ac532323ca
z068f95d21fbfd92e0d5e567eda577885b10cba5d78ea5cdffb21e005a70c0aeab55a3b15dc0567
z679d1c3896a188ac37fb693aec935f8415009a4070c02b5e9327ea7ba9cb296b5fd46037ac067a
zb79d5aeab95cce24a0c2aab9ffd3bff78590b8ead06348e0968f157ae17024a6bb98d17d2317c1
z66caa5184fa16938fc909b8f3763be15437aca83cb2258d34d0b234c867e936ce08416e730ba52
zf3f8f2285635208e5260c5b48d95f917e46bc78b570b2a3e763f815a54d241e8404d6df973e395
z379a66cb734feaa0642007466eefd6091af8c4acdb9f44b7fdc0e993dfc909c6196c68a3425fd9
zc2dda9266c2d681a0f480124084ac4df2741353c29c4132bdd32ca94aa84d36557555c208a4706
z8b0353666ae152b65fb12511727575ac229b2c6797becb8f31a9ad56fdf84f414d0839b71e2614
z387c3258abcfbfaba1d09723e7956ab978cbb67d058ef0432affc8a5994fa769344a1d5b1dc172
z7d620b696c5f39b919466f2ea513bce677c45c999bccf79be11848f51ce648a3305071de3a4ac9
zf20aced29bb264e2d44a3055f3003552e0814f50e0670cdc3563f4d40acb5bc7359acb17120a9a
zbb96f4c12b0f671d750ba81e13e62e0b8ed4c76c75100f290b7e205ac0f03e1a8b2817ebb728d7
z269573c1a153e60522ec149f6e425952b30a99d32e163dcee0fe95a2fb1b9789d6dc0abcdac98e
zc5f5f7f746d676bce388c6b92f2e99e7f1231c03a6d6ad23f618a5ad690c9f4515f36c3e867238
z416efa7333fb5491c049453ec4c20538ef9588d3e74ec39a333fd9150ff5ed7bdaedafa340b0b4
z7c46b1ac2a25859fcbf19460ff1957846e372d244e5f567b5b28d5e759570d10202176f0a78791
z948eb16086037dd2a04a4f5adb83976206ec119023dd79043c0fadd46bbdd1635cfea2ee94127c
z31eca206ee9a1a904953e1dc16c72d98de5ed499b0e088c375e54552400c5e5ef9d87052080015
zf6148d295e9af3720aeca4e6e443a6ac2ed3832ce8c53b05df499d61db37908c242c936957657a
zd94114cabb875aa37d11f8140d691ee05b8f0b8204406906972001f7e964e39d39a8a05b15383d
ze9043faa7a000f87d4edcaae2666fe0dad24d9e1979a7e1a0b06539883883a47f1a067f1665b5d
z8a7ff5935929b5b8f0fa37700e1ed887e602f7ee9458a8af2cb30371cb63567db08b5313fd6c43
z291a7f201fc95c43eb1baf0708514f8b64e9d062461c68b8e44eb142e68559e77a9084883448f2
z662d7836b03fa57ce735005afb19c5452ee5b6548e757ca7106adf2a37f910b721b53b102cf182
zd97e974272e091a05978c9759aa2274a9f3331dd613f7f285dec1c19c8e84261701d595d46f56e
zdc6df660b8d610565cbb11b0ae2b1310391c40b427f5731b962605f3f9c7cc9a76040d2c4a98bd
zf8043ddf7b8949169a0d27e78e8cef629a242f0e943be69eae8a3e93f304c525946f5448a1b97e
z40b6a1e065189c6a1ee729eb14209f3b1f03288cc1847ed9e7195449dde656845b2e447372235a
z4d377e645698c5a3480842852edd734f034821248ee98396a80938eb19be107766ae706ac98d45
z591c4a2535aac5c703d1339f3e6b99e75b059c80e7779a4e8ec9e31a5f8a70beee179407646b56
z3ec3ee157b5ee6f466fd0fc0c31a05c6c7938f268708d5dda095e7d5cb2bbc0facebd88c5b5e26
z500411ecdab748586cec5d3035949a27bbb28f603647c5396474db5d5ff89001489cae1253909c
z7fffcbf6603980612faaad642b64750ef189bb446978c58e07bcc0470b336b50eee0fd9b34c3db
za4fc1d6a83c6d681d1ec53cdab3128e14db95d21936ca514ac0536ecbcb9664fa040ca383b9fb9
z938955a04bde18a4ea9bfa30a309ab5c4e75ed7314972f76dc88f516fb9afc85af81cbe8a68278
zd14a707fb63872f3c1f5899564feb049ea2e0e09fd19d2b1e61f2a3b0a6f3ed8115092d5542e9a
z42861eca1be03a34ac309c0b37c4090eedc511cc82f1016d9c421052aab0aa2d147eeda2639e14
z90f7ffda5163241d9d9f69a391e340ca784f33f6c1f08f3eed55bc70edbbc7b2ea0a82aa0b5522
zf7e024b13c182490a1a0bff1b39e2958843869cec5a140b57900778497720e6072c5dc3c174117
z31bcacaa0b21c4452f00509196eae804b8bdd8c5f4fdb5d7e6b312ec227edcbbc725008f08d018
z6edbde914e872c45b9572c42954a3a5328fef17baed7f8065dc5ec8300820dc446f0b10066a9ef
z0ca9004fc87681241d2f7ac9c2894b442548fdf5ea6c9927a9f69f8ce1ed15f30080b1377ad07f
z4a11201f9b7a29277e473cbf2576dc73e66920268eebc51a1eca1881a59d4cb847858335bfc86b
z90d9e2923cc13b7b959f319621891c12ee74b22329ed0fc23a4f002748eb08917b1d90d9475a23
z3282c6e97277382ee0772ae349f36051076b8ca3ef02b7f8eafa5f068a29bd077b583ce16bdd9c
z4a686e61fa5b61f120805741152d30004f57bd82ff4b32ff75834e51d700b9ed7c006dda0b371b
ze75e5d4293071babaa87bf094d85ff1fd512d28b2e8c81ac1da749986bc37b8e567103ca5b6ccc
z22cdcca3603fe25c95fa98082678789e93e85a3afc2c35131c15da278730e5f194475baaf82b0b
z54395119b8e57417b2c90815c07db07bbb37f127df285611b09f2397b4851ce780193c190fab36
zccd19a574f41be2281a40486c459bbfd1b29c8a142aaae741d53b4048902f55cf7bcbe4e48acd3
z058b3a68cd216bc1f948ad7e6bda50fdb953885e692ede536da88a2f87dbd8efc561b64eeccba7
z3786611e167ef104ecd73b7f629d8eae0906f33fdfb63db3dcfcbeb66bf37db1c5ccd7440d48e4
z231c5823169a735284c5f4b8f34fa176ed3dfe5d81e137cadabfdc6297f43cda5a7fd61872a293
z3f649a020dbb3cab864f6ba034bb237cce6067fa77a1a650063d92531677767ee1091054b73bd0
zbda4b8b7abf766182f122cc56c270674caff51cb9fb05952dce3b12f47487228bc781cb3563f6f
z0167a2303fffc6e344bbf58c664b8bc2bbc5f28ffe93f618a1d7a95af646e6e648b34cfc6edde1
zfcd1233db4637860159d259462ae707979dcdc1a6fd673dc0be73e68ea0dad25dcba8a318a939d
zaf253cc3ace6b3a3c766dd7475e163c0b4a99dcc4902012d1f6d1b49b303308b0c78ad0576648e
zd7323db7d85c4f45f2f94be9e486064bbadfe19bf3369137dcdf51b317e4fc0fc0491271011aa3
z5a8e694d2d448c258729bd1780b7de1a01ebf280dbfbf5d5f8b970e57c8377ce38a05a4ebf8a8f
z14ad8c0c0453c293dd89d9d24ee633079b2f889bb482f6ec285629b1da812e8c8fca603f37e743
zcf0c312cb952e82842be95e361f5b0c75271d7f6d022056d7fd0e387d5400fa9a446c56c6b6b0b
z0befb704682a625bc5db71f7441c2315872d95e5c690b05f66d9bad7177efe1f2987d134c64e03
z05f1357019d610be0b97b2789ebcd60bd849b4a648235d9d9aa4d191fa5ac6f7ade0f3974f91b6
z3c87e04395ffb01a43bd92d6aed3ccf833d527270be239c058397be43802d9c94f0faf5bf5216b
za9be912cce0740986c03155ad83d1ec573cd0493e614b3e42ac7d84ea0e4202ffecb98c875106c
ze284bf06e16c2c2bcda1cad2f1c97c2844c6f407f99cea22c5e24d19e112042b6944f6a9646221
z3275524c4c3f0eff0a532c187ba1caf57164829f4db2db284bb610fb9328721bc7c183989098b9
z84e0e19dd1a31f223456a930baffcfcf2bd6b2d0c0a874d9f18e89b6f932276221b546d817e49a
z6f73aec6733ddaa0100ef0b6698634726c04f4ed566f6365b599ce2eeebdae85a7e89fe13e9d06
zf5356551a3a0d56cbf6d4c3a96402cf8d1fe485670266d35fb9affd7448e29d86d1c509d9ce504
z1191f3db8312396f00fc7e8da310b9437c5e21c65d29d03c985e6f9ba3ea90cab76c5710271e57
z0d49fcf4e5eca2fbb21ea6cfc4798e2cefe69ab6587c231acfc83ca20000791843e7e72296de32
z351934d05673d8858d08614d1555086b8bc31fa1a1000577406744cc8e67a0c53772491c49229d
za560ae9a1dd5666eb68bab8d1857218558e8c855a989bf58670f0a86e8a8b9919519dca879d421
z0a4a767bfa54bea2d9e98aa90c6886a5e77f7f7b566143cfe0da132120f35852bf4ce06a209b3c
z01a360b6dfdd4a330d0aefcefd4fd083bff67fa1f0b12deef5467facac61beecf247a7192a8185
z5226342247203d2f54211ae0731cb754213015e00883cd6e7f5579ecb7292afe02c11a15864dc4
z90a37f34f155a9c14cd9efd5e1ec591e9f43dd3cc2381818c09b90d666a592b3114d786b03c497
zc52d0295b69637db3f1df94427c29d75a8b62607fa959199ea6fd463a930d57ef26a2fecadc8e2
z674e0032471b00e321e3815263f88e9bee2ea6e33b1afebb9c532d112216842da64b4c9c986248
z1bc76a4c9a526f75e082456b30df6bd5f84cfc547ae58cf5417eda81656cf4fc8e6ee55f8873c9
z87c06c97775fcd1c8d7896fcfc0e66540a4b085f20810cbb547e61c97b0b4c290d85e03aed99ea
zb22a1c5b1272d8a572da60cd4bdfc9b1d1f7dcbcaa302be9c73c0600ba053c739a8491fcb2e722
zff8b5aa4e7bd7d9ca9be8b004033ee91c3944e9a82a14542dd011f735d51bace5155db70b47b13
z91236653ea1af918325c3d2284ffa36f077588ade0788be599a9f239a7f49ed1c05a5f3e63b886
z7c38d6956986ef0ad4146c94e27045463ced6e90338ca386dafff81fa8f9221b2b9d5554b3616d
z44f24117ecac3538679a4adcf49ddb637b1eef54f72ba06e874c9fbf9163abbdcc4845f2417383
z5ed4af2f9e23e251f4857394ef55070d94e60bc6402c0443b33e5c35190b26fb1bc3be8331a0a5
z678c4ab8ddc06536db8d30caab4bc8364950ef9eebcc7ff2951b5f9a47b726e3357b6712b55a6e
z4a102e0a930948dbfe22e1f138e6ac7b89cbcfb3d28087b4503115bbf0d4a85ed04950978fea20
z2a2fde56d6e637c786d7fb980b56c400cb2e7dad6edcda95748d1e5622256a57291893394dc35a
zf0b0805951050250c2c9fcf0d3aac3d3e326a54bccc6243670ac07e943dab780eba5168a452e98
zbcd43f7de896ca0cdb1e967b09b11eb2a9e688a72bb0bb62c3b4a5fd294978bb2d3f81cef491aa
z9b8f1076af2fdefce087c1125713e060315b27ca3cdeae965c851c535642f7c3963e25535be754
z6abcde2be909a1c25d4ad55051c69dbe1a4ee40de59a4b49ba53a393d8500408b5432a55f7d6e0
z1da8443c128d1d50e9927595f8c72d2e16b61918db3b1e9cbf74b9006a4e4b41b8dc9a10077a8c
z672aaca962d017603422e24bbe8e9b1d40a9803edd5b99cc0ff4192caa0a56d3df8c8083805d4f
zb8c95759363aad4bc3431d0f8ee809f3247e2cea091ad0e3e46e9f31d74c1c2330eceb978d1610
z2388e9b3f316ef9f1570846b52ec46aa09b165def4ffe65a4d40cd9a9238beb9db3d2d2aef4c45
z8ee2c8c91b8acc722bff255b5e0ac2b257a94a8cc8f2db5280937d9b9d32233a5f46bda34b3bd1
z620a040c46f0f1e32fe151bcde8b303bbab4096581f6182e0ec3e9ff367b842983d8a97d1be7aa
ze383f4e79652a77d6b4f4d61185a50c3d6254a2cb049de797b2c272ddabe597f15a7250126b7f3
z936e7c007c07eeea02ff552411f410b4efb00d429e4528ae3f1710eff4c37f31f9861c5fa9c463
z1f191f48fe2a2feb75628054566506bb44573ff9b847aa11930095d6a1752e50e7f45ca800f74b
za361d8fd7d38c21985eaf4067b88ac9f05b54b32221b2f1d2f5596109fa5190c487ea28cf67b9c
z137ada07a80c72323c387f80f8f73d0606447a91431850b89645c572afcaee27ef6d8996fa126c
ze1f64cd831e7d470ba8b3765e4722cb4c81ac990df671f3d10c6bfd38f528e38dc786723dd9f41
z339eb2245fc05fffc9119e7f5ca543a7191b6f2475546e0ce9ce920132857c480a786500a42200
zde717f27b6b90c0e7ef625c09200ad708a8432722a54b72c1e9d4b83129f9423b118dbf499da52
zb75a14e6b26badd35065cc001ceedb934a52649e7ea943afec2534e40cab532b210478063a566e
z9ff8d9140669462337a3fdad7c9d989fc911aee9ccacb81d34334f9625df3acf660883bc790d4a
zc0e01e7b3e66e146d631249b124ade12cd5f3f19a9cf228788d9cc66b7989844c03b7bea4457e7
z296eb66df1021cf2884847c2a64b4887afbc2ea69676cf1d9138ad802020a68960daafc1f2e420
zfb427d2b0e85c05b5bb0149366b733338bba3721f2982ae298937fd8d186d4cec06d04f4ee6191
ze791326705ddd2935dd95ef51a0e2e202e88d7040435c84177bf4ea729078ca521ea86d356813c
z93f8d3a191d141fbae8729b67b168d5d1ef37df4a10f935774f62e2bf6e871999b988e7ccf78ec
z407c9079ff16b87fc64725e714b13328b525518d23cada31a980580be6d8ed187b2ec77146e960
z77d09725e217bf477fd1ad7c3ceeb9882d89faa7adf162f2250369202fb936864abaeb96736346
z873a6a35b4a436591ad27a13d5c179708b306e88b0e68547ac56f459efb6cfd69ba17867d7aef6
zb3867fec15ec7ffe0c2dcde45b7bc7025694562fe87652a8bdb77eb24cd93553e7251c741c7071
zf9d0fe19ccc8e5fb7551cb0bbfa32e73b1d8106988e8c43c4a20922fd34ba4c3c6706258a8e80a
zf6e0a4e67e67d35ed0472b6d1d88de35dafe96b337bb6bd954f2926df7cca4a8e8fcb619c085bd
zb7bce7334fe8e975aad630c74ebeef67e24a78ec55c15afa59073d6f9b0dc739a238637e58f104
z913ecc93dbc825e042e53eae00a46594484e76637ecb135c13e58d6d77635742ffc75a29b9a2e2
z961ce917a2de500c540d8fadf58173683bd78cb1f50603fd408ed4a120efbbda92b403c853b209
z88a201098a9404381376bef3eb76af03d25fcc2d34ba6f7407aa5be7aab1c33f959cf53ba1f5a2
za40ad9ffc99bf3ce6296fb4065e183cf634a19d1d6a4d9817ee75bde7518c17722ec3022e754fd
z09ac3e17d355d9fca8f88eb2aa6a73a0b478d163764608f92c45de5a0e125cc117f79368962367
zce502adcb8f24f05bc62156defa63b706932bf2425dc845a9956d47161edc3d29b74476decceae
z4b276a710c98d7b85ddf0c437af666b1c6a525b1f9a00a7b19fa0d1e13c114967f6feaa5adf182
zbf49815a4ff85add29b143a98f23d8d2e0008fff0477b1471cb908b721dfe41b4c688a145459f6
z22c80102786a3f7da9917dfe9e895e529ae751b9cf5824b318d97163b2a7786bb0c07b9a3ea0d1
z49b2b62bc7761c514911d79305db5273f663849a9ad2aad7e94389cb7767880335ebe45f5e2a88
z99645e3d58de98b39b1d91b629b4595c1eac1c083f673dde40c752d1ea3b548bc51056d2c119d0
z11fcca2cce01f884b94ee42bfccdd84b80e4894421b7e3874a86d90650aab681141af498e0a439
zd8f83f75d111696afb1cdd90c10f07ebf37286c29427b4791fef440d45718431cabd2942f2d687
zccadd398d1630763a74a38d7edb3e567613a206a0bc37f040799927b659a5ba8efb22c5fccaff8
z782f154ae4973f26eed44f20b01782c9f3f58e7a90699ddddf8c7dbd9b43254f74c37e2f0df094
z8bbe1fe55ef144f9974f7fcb9c1c27b76bbeaf35042bc010de557f39ff8c1703ec4b7f569389a5
z8f75d2f9f2ae006c71322352f97c32478b421343eff9e78e902dfe51fbb4e1b4ab0128c2e2c869
ze4be37c86afbb446a2b4d638634b9b4c8a50c3ac16aadc276c88632b761190132557476292a24b
za888a9dfb5e7283aeb922e2a6b776a2c93b83090639674088246f7464d91eebc535117e174ce65
zbe6742186f8e2d7341728eb47af5830f9576f8c88af914fb885c1ac69aa4816af4cce3b45a898f
z2abeaa5f995819bac700f91b564fccbc8b0f7642ad85c80a5083f5aacf302ac002b9ac1b0c762f
zd3952e05ef979e3629a856bb63cbb27d120a73209d4b65fe8c1fcb6e8e9684c8d6d6f992dc86cd
za64bb01ec6f1c9ff554ddd43e8bbd0e4d0f3d2831758c3dc9df498ee07cc57741c68f8fb112268
z554d444f27864559cb9452f8fee33002a07bc0952211f8fb73b287c5673b881f31198e0852aa48
z11c1f064b9a33d6e5153fafcc2b5b5bcb233ed2a7fe6c15d30f87305f3b11597e0466ef92cb028
z53e3b736d3a3bf579989e284f40bbc4a7310e3fdeb8b98ff7990dded545b070627075fa10fd60e
zd4b49560a93934211e9442f539ca3f18b966fb338f4d37edead687f665690aa1481de18f677c3d
ze78b581d485346d41aa4757dda5ca9e2ee1a4480a2c38dd586f1ff0e25fb378e03bc386b839d99
z2ec060055471d1c6c525d44ff3dfc58ce5ccc418046485a637077da4c60258a7a6c7fa77b768da
z0b6fc6c80474ee41405b8d7d8e5c8ea9f48cbaa2c2be93e585608f541f83f6b74abedeef965385
zd83907dcf1d914a5cfe0498c36980075d2f46759123a7fc060bbe3091de057060f28be8c4ef7fc
zb17ce65e54685416f052da787e7dc35d6a2b018a93a6e576b9312448472d5c0f3b7acade2ab8d2
z595e1e05a65ca3c3d68c61b2ef486ae70f2f57b032587e28666a3ce661f1ba9e2dce1aea578e1b
z316a264af6c26ddf394dff37b03e56cca272d3f3398b6dd8fc8a182018ca7395f8989c2e69f0fd
zedf9d649e242a0ecaa6a17ee20bd39ad214e970f3efbc3024be885043eb7bf58be5223d30b71e2
z351b3de67054987ef65119ccd199a48a66ed1c101c2cf72a3206bb49794fca3242a9fc021be124
z26940d519590b0722e59b563e1e587afa41e04b54c1621f2b8761ca1a2f5498edabb976446bb48
zcfd0cbbe5c3402e9734e7862773ac0d3d62eb1d9db0306a5b6682d11edc31eaca75f42cfc39727
z9d5d409b0529caf18ff590028b1000b651640e9a0e56a69d9633e0853d4b64b43d28d3cc87b3a3
z690ac34db89e87867bd24a05394eb438cdd49fc1ed1d7248b4a29c78f1d626497cf3849628bb68
z9f27b2e0c7687ea74741e71add703ad36aacf33ff489e4e36762960338b9336a83ef3cc36826d5
zb10fcd2d4e58dc94d352edbb480db8425c824f40897af489ff714982bc9a88fc943bf9653c1aa8
z63658e3cfe802725a928eb3a28ae892b1168ce2e1a8e8bde0f8998439e49c5f9f2d24c9c872e6c
zafa7f8157f6bc1c98a6064d4c92ea33e89c19d3cabf3f1e15f81fabb0b2d9172489618ca7fdec2
za07e7f05f504d3b74de002bf689a5bb8d8cab4b7c53139108d3adbe3bca50a61f9ef986f2b4e06
z575f8e7bc8508237c906b7589c79c4379f572a1a011486d093be610b7c666f46d787bf7cf23bca
z264b44fc61d55dd41ede971dc466a0eb43f8c6633b860b355ef609faab175a9abbf2bc7a090213
zb674f5fef45af00fa1edd22cacae497e1e73e3eb5a5b789ec65b6065299f09a7a7df501873b352
z92b7906df5a39b62d03d8a156f02d455b4972b4fda1ee701c76c9aee619f0cbbb6f76ecc4c7346
z9973bbdcc62e0f515d1440e92b1a5fff6e506d589a6c2b254b3c9b458519dbf336584386fb6e3e
zb4eb9ce83bbbdfc739b552aa8af3d313f2e4434b2f2ad6371053c5688b8c72752474f73f6e28aa
za2c44157b8a7b11531efd94b79fd61fd3e27c4c1579cf9c465c43b13e797934eadf4dd09b1431e
z01f123537561b24229dbd574d6db56f598d0660a7b41c914a7186d1dace98aa5921dd1a5b5967a
z96de708f2b38367b8ca93c778e13f843c21429e3d2861a82f2620f035a8dc8c9a93aef429379d8
z6166b863ab2c79b5c123bd5df4fd1c5b8a6da2e3c1e4642e062c50a8e21fbef6462ca6213f9eb8
zcb410d44ac98ae6be6e654f0e1e9366a093ed79c31837ef8c7c447e47eb880a858ccd524a12414
zd18b22f590d9fd2372f2d4de83656facb575e9f4d38aa75dad24fbe7dfce3b0590c068a4cd6d42
z1a3ab1ba3dd076578c2339a59044b8cb3632f2a01170229d4612bf2349c65254da57a0dba796a0
zb7ed4e37919df48f986f97b15542293e1d1a443cff81328c991a35bc7e81da2885daed5552efd6
z7af68821390e968836f4f2f7cf918de28fbded3c28db4a3735df580ac0d2967ed8f9690ad499ef
z6fbbcd9f03e0324e3cbac34fd0adbe1925814637abf5aceab8836f9c1a5e88bbce47a8c0ad26ab
zfae4be8723f81b0175413adbc7ff813f25afea38cc02f034669b21ea382dfc641642ca1b601c3b
z05f32c6629f1df6ecb9e59fb5bd8f958f4f947004a1244eaa28a2d475c513df91bddce21bba00e
zf1394fe37cd1dc26c0b54961e56f92aa66837f6f43dde15026b259a603b87cd841738188322982
z0ff0be03de19ed60c054c6429784962db5c354e8f3a9542fc0c8f25adc607ddb45668de342891b
z3d93d8dce97af689f99d42466b66517937bb24d32819a2a230bda4331521dc0105f930968ff0fa
z7ac00f212868a0391f26c85b06aca3ebabba9385c2999dc01d6b0a1b81968636915868cc1a22fe
z78f9482b49285a434a56d8eb45c354e51d37a0d7c85acb763f09306824a437a5780d12cfe0a40f
zbcfad3135d7da908ed4ebf48e4296091b8560a8e896ba0722d5e97c6a97ddc86200a7ccc921208
z2395259ffbacd11c08cbe9fafe1a39bbbd42de9085d27a29d8ba9434bc3b23678feee75babd954
zea45ca53a63b6765fcc0430b2a47a47a13065cb76c9be5b44e7cddcab7f01208a0a2e84a68f141
z3f794395f4c531e4de2b76c23e05c116f8a47f799cb0b2d0a5ce26803e12f45d8e6d43e238c319
zbc74e62cf5fa54e6e6f4f8dc900f96fa185ead0e3baca2a166714a54b2c2dfd47a081ae19690a7
zce9ef3344bea7e7623e798b1a7c6aaf2e02cb04af59b6f3c5f92eafb71d548c3f0164facb1721a
z336327937aed90e1b85c178c61b11c4fd5a5ccb7f96e18fd40530380f9a54d99dc202ec884db63
z066932aee4744ce85d3bab6b6d335cc46a6f5bfba27fa9ae61d3d141d59be4b9eb33d12e093d19
zecf0ff82231ac2a6d89565e6b8fd7a153934e530d97c70e610e49c5856e61a67504ab70976a172
z79575cbf2f938ed54042fc7eb314be89afdfafcc9adda9ee2a7b1fd52d3f3d2e6f3df16f2225a5
z90731d3b1599f6bb24f83debebe090f76e8ca740a6dfbdf8829843b32d4c3e78a82b12b54cad88
z0f0c1804d4c0b303f9807a9adca4a616c97e9187d95d81b01f8148292882349e6a4234be1cda74
z268e48dceaa500ed8cf7da20d4fee047efd2cb0f4be8cec6fc0fc3b3da6ad3cabad1053174818e
z2a4666ef630e7ff8ba8608405c1364270ae3372212a90601bb9163221099c86ef073457ad1b558
z0ec0166561375bddcf0830d429ead1787e31248867f27b83347ec72607bc3703152c8156800b07
zd85f100eace3b3ba1c1bee97157a2c42682b97242d87a67a7e5222d2d152c890d2db350a237f42
z7bc7c7f68e06c5884a9e21fe908cd959495acb11d683d156e5afd41a6f6bfa86e45336724daf11
z1fe102b0bacd9cf4b385e4a79870144cd8e85c039999faceceee7095119a4ac475bbe4df1a8de5
z07fd6c368795a4ac7d795ce01d4276c887794d583067f1054349ad53ce4830655fa6a6f78e7222
zc308f0c9cff18b88aa08b80e055595ecd89dfe0f09d1ebfab635e3f86933e6475ec91c70335726
z24b121d68ea4d1db25220cbfd058d04b9a372f16b4a2a7bd04eaeeb377bbb52413ae8dc0e04b53
z38857d2c46c5aa74539ad0f95383bd1982b04e123068e3ddcd99195b694e3917a3b659d2e66b57
z0fb8b1b8b4450f05a1a647e8b25aa7376b8d18b0a20cf764d926b9b4415d1bd15795ba38c15028
zd1cd1d7c69978ede099efb355ccb557511b7e9b2cfb5bea903097da0cb030b37434f7b01fa14a6
zf06b56d4a450f4379325a5e960b6864d939be887670e084e2d7194e3f5f04f5f0ff7ee4d24ec3d
z45a6a760562fb5f0b8dad1c05d252b7e351cfaf60d0fead5ece681da86dec2dbbe001a41ce523b
z434d15df829c0f0b6f9fd16821cde91845114342f507b90468d14e0756aec225611cbdd6e0fab3
zd9870eb7342d08e6fcc99e14c23bf7362c1e51c14dcf789df62637ad6b777f3e5a2b1e453af60e
z5ef63710c7440c511dca3dbd8cce98f9e5ba8f711d7dc30e347ec622c90791297581414f59e7e6
zab914c5b20fc1be972e1b981e85570f6c640f45b120bee1c559e72830112fc3dfa48e82c1a3392
ze145c40a0eda130f95cc874a35434a8d3a8c0d12bf673314abed4b99426bcfafbf720df708dd56
zf318b2b0c7341ff9dfe09d033a8797f41c72b0ebfcdda937195bd6e56f1d9fb1b259ba1eac9515
zaefc2c83b7f2a154e15816700682e62a9ec6e40ecd27b06e3abfd424d463c3c075acc370767f38
z1a843508244e55756eb6ae9b6755074bb68a31620dcedfabe12a3c5c817ab111ac613326e3dfa4
zf652ae653730a26f78776d3b493982acbed69d538fb3224ef844ed93e35e4453276d23e1144058
z38021ee4d1c9834341486fc0155181a936c9c22cb131f30933255df981d2d164738a7072bd8648
zf93932f5a9829ad60b00256bb8692e5e394e206f0f05c06e4d10161820b06969b58339ee6b890b
z081f3047655fc20fbfeb925939a6808917c46142a38684be0b8bbb6c8314108cf03d7df21be929
ze89cdba0be09bcf6ef1b7b3f49ecfc5653d0bcac4a66e1a8f2b1cab58ee35018e6ac0cf26f4ae8
ze24cd7c3f7f74543336ea9bf31e1abd343ac80f98140f514b6498ffe708b75b3961549d60454b8
zdfd4cf2df1d4211cd14b1b1f2d47d6153a07185bf0da4d652afa0c07411c97b3319581cd41244b
z51b5ad14232e5ca06e1e6188f35a7ebc96d54ef3c7423ea38b347a7a4cc502fe8d11165136b40e
zf565d56867097cce73d2d93ffcda95419088390f73e5bf72ab7dc2d9f9acbb364dc4110827758b
z061874c16b915f4155ca822ad2798249ba3229f31cf6284d1fe8701d7cf06dc952b5e23aa15ccd
zba874d7226dfd0787dc1f7c84daf5616b926cb985f8f8cf74035c227bc138d2561b331aaac3b5c
zd49b72a2b8c4b8c05dd62ef6f404888eaf89947ee3172bf4829c3e4932ae3bb984f78ee591aed6
z42d5f05eef44fdae01ff9c71c3727c489f00e659152533045906e5b47c0425e8f699a41938328c
zc76c8060f54ebcef8c7eb175f5b543b9c7e8cb0d4e8cdc85dcd296bbc526c3abe94795af3a002a
zda509be9386d4cf93d9f4f893c11c8597a8572791c957a8f91c48992ee50be40827f92d072080c
z1cb3c6b2ccc4e10efb8a8181ffda6284b89447d230bba5d6448215c874de1f72a44f5985246c4f
z3d16a698a895c22c45a0329db3012eb0f2dfb8b132b343e14a8a25cce60ecd239203b1970c89bc
z63cbdf3dced4609491839f89a2a140b5711538d6ce950fc37c61eaf930c617b54ea433790f4358
z077ff063ef12f2912c3fec966187f9b441a562701d632d56d82abe6bbbd677067454551819d03a
za4cef06d771ab73dea1487b0c62a566346e6105767cf80c8fff1f17de293e35870902f7ff5968f
z01ce66ac44e6e881b7de4acb86df95194d4f4f71403307916553af242c8d41e17069e9401ff33c
zea6c6c269ab3a09d7b42dc114d4036321366e40ee5728b6ba169cffc5398d52869091def38e0ca
z3d1a8f99f347f9cdf1550f63c69b2e0e8f9f6f6817fbb2ae460568a807bfd01da3b3074ce10720
z677b6d022b635a93ea5f095946f6248107018f5c7a98449060ae26aa2fd35a9841793603b5c32e
z285f102d6a3a879138040fca27a768dc72f152118cf7a397b256ad9b272531145925ef87fa6023
ze309232b00da0cb2a69ea25a6f61575ec1f438910932ae1d510794d54dd46ab4830691174e169b
ze847a6f6b5e89d98b57fbd50f721e20c5910affbd6b659842d578a2ea57c004fad54d66aa957f3
z73436696c761cc9f2dc5479243713ad1f8fe72d4ab721166eb705ced98b21cc3789182c325d091
zaa17a67ac1ecaa00c2f941391f0eda8f95353c73a9073614d4777dd7b42c81b4d02df46a153519
za0d4b17190b9e0dac4cc06b8e02af3c365325784490a13438ab4bd9ffe14e562416b45263d3f36
ze24ae958e5c5d1e9394b076a925dd724a9bae74364ea7b717214e3bca55c0749b31bc35c5395ed
z0eb09ff56d17c9ac8e107c04d87fd222c8c7070a8406536a44f33a025e6503fe0509e6ce7a09a8
z3b4361d89d73905cb608622f01bf4bfe8f9f780767fe411929baf29c0b05742ccff0e8be9943ac
z54ec91418f36f7dc864a6a2a31e5fc3492120ac4d33aad731fb1d11e81c712a485b8db93ff555a
z3576985efd753b6ff4bc6f25f86e68cd11c115b717f6a5abc9add23487a097a40e1d19ee783b1f
zcb8d12aa2cd3e044daa56ae07c4b39682f62109fd1552be48cff3a6f1bfd2219c9168a6b560c77
zdcc3fd2ce52c99b1be1c5d87f4520b79b78b60cfb733d075bbd38d6b9b7fd640b7fac87a43dec4
z76c67ee3479108d0dfc5a92787e6489f4bd0bfb3c0bf5999b419fb2157685d7548844027890827
za4c32778a4aaf93b19c053079e18ac6ed599f4c05e4050a1fc379fa082ad45f88ebc723e2e90ba
ze6655b58007a75960232784a7623e91877bdd21084e45fa6dd07a0435ab5a765404dbe3406c81c
z18ba57373e5ac51a50ceaa5b00e3405e298fcfea562b8e9410098e027b02d97051fee9537f1cca
zbe965cf261214812d3bb522b4374334b8f75583a2f3a546c9ca0139de5b927194e90aa8a5aab6b
z3124a72ee8796d96879fb43c7040614b763cbf8a45eca54c29f9ab90324f07b715f499eac30da3
z69ed8202d2b15da9a1e4723fdf89256aab57f12a7ac278293190a8c4fba912e12923c33e8486c5
zc6dec4b55f82305e64b7d7a40065d407026fd79e3ffa81478c29bfe89609c4f009c36281829512
zcb4faf2d228d456660122fe95713ef67a1c613269853d8a6840def02e4a1956f2cf802a5e59bb2
zad34107446783eb4b81b5e4158e337a2f388e303ae77a65b27702e6fd629c81d97772d5718fa64
z8374abe54b029cabad8dd097fbdef0a9d0a28dc2337aee4a017168f17c5172ca2be57f64994fc7
z2fd046a6c97334d2053d7c57dd990e179c74a885d514102cacff974359c209c6baf10ea3cdc9cc
z0e2866971b10afbfbaeb3a0942f7e354f44a0c818ce1014e05d2d6fb104d6f0f677d6aef9b5ba6
z2b2f7a6348457f298fc4c0a50d85a32fc173058882292ca30e1dc8cf227d0ec4b22fb4688a2446
z84ef36ccc955e37f97479cf479fa4315b5909bdedf701e330d1961267156571619bb51a9fe4cee
z64be624b667e194f755f8fdd71b36cac0534f590be4d82d97bf5f12c2cdb5356e11ec572e1131b
z88ce36aecc05bd8b0d0d0e9769ba02adc440eb642b3ea3a841423c572922b8a238ca6791e6bcec
z6b83e73e7f2481595961b1ce7da15b4aabbefc2a90742def69b53c8c693d8aee47a0a6dc1bb638
zbd5e3cd41107b7a881d0c401b8d48ab0c71277034bcf78bd570c6f1425de6101e48f12ed1b490d
z6e628cfd1c782b518a7794accc8e77a1ad7c0ae1433739274e5792db31f1e9d9d018c660d91b80
z3d1295fc4afd8d1f248ac8dfe87db0350cf8ccdb03a7ec060b1059edc9463c238f4d60246b7b68
z8c0e9a04460d724cbdd1c8322f0f0d8587b3884a7c3ebb3151b5825016d6cebc6ed54bedd33bd9
z0974db376ae22be66720d57b5c8a5c66225779b9de08c4b3fe49d2ac8ea0405252ba7d6241648e
zc77476c57b205385c088398a70e0f1d07950029ab7f3e69304f6a113f2a8f5581c6740a56e2032
zc889765a8acdd31fe4eed3cae73f9e567762bc2cc56e294626b0059788e9f4242be1daf3f94a10
z3401b6752db28d3ea776dd27bc838462e6e738744eb9fe2ff489ea1eaa03668765aac6df0ad34f
z58374daf38f59fe4bd19318728f1f1062e29fd6339edb6d0b9d43b1ba75a0fc18ffba24d20a48e
z5f179da7959083ad1a684e3d67e4e28c9adac8609ef3b4bff7f0516e82b5f6df74981c493794ef
zd25a442524060a1563aa6a461accc7d1b7d35aa45b4caeaf3159107a6dba88bcc5a123b0fd8ccc
z90e96394941bb7fa032a5fce830a73cfc99b181759bcd402a000214b7dc71c839a429f304525ea
zb0ef4de6acfb14c091ff2468b7cf6effbe229381564e38a389a111d598058919c305828b233ce0
zd61d50e848835f6efad84d368ef93d10dc3ded3dd71795195ace64cbe97ce5147a931d66b81d19
z5e60aab04f742242e168ad1b51cfaabaae3b57bb9c1dc80eae24e4483be9c0fabe7a3dd8ee9cc6
z4224ff3e4a5786dbe144619275be57d7163519c2e7d3928e5fedfc93eac4dcbae0615c8eef61b4
zaf94a306ef2639b987446ffb073e99808bd61e8c1592633b667759846e00a1147636acc894a246
zf03fa01aea2a2ec1a65dc49b4cdc33c3faaa1236f2d10010a9f6fb7231b0d40d528ecc9bc5f35c
za64907b1345dda3a5644d24dfd999e1907c789f04cc3f7df30031a802ddc80793551cb48107648
zceb971a551485bb0f3e50c876d5d1502733fe2e83963db9092296699cb03ffe93bd23718088508
zb61ae4685a7f83f726f4953f49207a3c739a4d93c6623facbdf4971304460a561efc4528f5c0c0
z1945fb6e879d46be81aef7da00f2ae208ba826e629d7c61bd15594c1b787c35f2d0a7617d1a132
z716e7b40b4c408fe61b8150bbb7a9afcbce96b79fcc936fa490ac5d2e63b70539564b9fc903685
ze050b3021fc53ef9a6e70f9d4f24609d60f01d463fb214841c96379abe01849f7cc434b6ab9d60
z80da4d9a7edd543c5be0207893f7dd05a8e860aed804197cf2d12fb5a7c3de2a6047d26ec0e95e
zea02e523f0ec8f6a08c7acc51c3255981cc15054852893cd21e9649d8d4507d7d370173b786ad4
zf1a22085e0c9dcb21cbffbb27a3ad1678c6929b049a3f3aa9592f48366d4a9ac5c393b8e4ed991
z56a4ac68d7774a4ce330fc9b1b109898b69012ece773b04b847462e1bbc9bfa6b3feb4d7acfa86
z31b859cf2d7f501c5c6f6c0d5e5a5aabda356f1e96e1a9a864517de62d03f69969e08ef20a67ef
zb246e6a2169591fe82403f429b05a03d5f8c65ff4e92e09a1ca7a5b8347ea05f4e3e09a329be60
z2ac6f9410c567101170c9062539449870da8aad0b792b66889926913b7fde20871d673b5038bc3
z420b405e9dbafaaf0f3408eea0343f5e76b70473c82cead2d6503d620bd34c56e3b5ed7e02e5e3
z9b911d6afcca561fc6eac0bf5ab8695e223350e0cd6777463f9066dcda737f458166863dcee6d4
zd6baf71e62509a084b6732674f6e7b6dc5a5a9424e81e54a7cbc97f3cbf7ae3c00bb37002df769
zc077324fde2e69c9ea8e8cf5c871fac38ec03d62315521c70d938e66cf648806ac6f457934b11a
z2264583be0b4878b559a7fe82ec30f716ee0443f1a45a849193768c30f9cf35b91c9a9ffa2a01b
z89f08db8377681a1a0f52bae77942bdc0064a3425b9b3e3d3550e3387e0440865de9608642a62e
zbdcec6128054917ba09f9984efb2cc8867490702ecb2deed429b05dcd3381dbaa8a58ad00e106f
z38fcd420f3d1b4f8a2d517471820b7c3b81495895b9c85fe89d1d32996e9d6ca984b4b3de27ab7
z3b13729212e1a835fe440b79a98f9f456bbe148354ff92bf49a99b9d628ba765323eb517f14a04
z4fed5b097327c2eb5537b13d740f853e67873e5a287e24ec5f3a57140573a75820dac4be9eb2fe
z618771fbf5de4c77aa7efde1cf13a5291ec946e6b5203f5fde2fff6767346bd63653eee1f0e30d
z6ec4ab29216a14953ed5220c3bcf4c8689dd96c52c94a629db835e1e56e02db848edc3fa5fe2fe
zfe26a9ee4c3f7b51528c5c3fa467f01e067ec405c880abcfb5bd886ee411639487cc5cd2e9f791
z5c88fe78c530232d805b7309f1d273271e7e96e879d5f90dada37093ca76d6f57d8e9dc9cf1aba
z75b29ee49fea07af505bc2ffd55a2e86f30a2fdebac66aa54b7ed46534960312e885960c7b971d
z6ab1648849bb3ca0ae093428ad916676e1429264d16bf3cf6807265c1c36278a5fdcf070801aad
z8e398787394bb65d1f7efa9d99430aa0cdc8716e17e7f6a417e29dc3f5f383e61dd5bd43269ebc
z44a55910dfe2f085382178130bd90b9109d3246bae1e36c5e71a48a009f9f1f2b9616ce2c0bbcf
zd9fbbf0b4697955e4dac0ef73d68a91dac7797720e8c34af85cc610f6b685a201e0d0caf207ca3
zc24bbc86d604fa90298df1561404514d66d0c77470682e31be684d4a9ae181bce5c4e015f68f37
zeaa9e7a65d33fd85e8798a9d7f867cd9d23a1a71275f24c6130205ce2f761285621154329194f7
z7cea5289339781d883159ba693e74ae9f9c8ebd06473cb94c437d98bd77ad6acfa58e56510b2de
z7a848d012ed750077e92f47033f2a4205f588d1df8d13b74518cbb4d4f7f6f59f2a80c8dd01fbd
z2b145585562c6d7c7a9e45aee8f1a21df0d524fcee89fad6f075ad2bd8e82c365bf6953aa94318
z226606ff8e53be01f72698211b8ab748d27a94131e844b20f8c1bcade6facce7c97fedae0126b5
zf4156ba3dc4a81bf36e8dab002eef7719d044fc0979708d86f4f769bd138a747b0eafaa26afc34
zc6838ae98574f116706e7b6a197f9f979b7aaa513304f5d0c25710fc906fdfd6cbd559e3ac63f9
z956999b6c77bc057041a4c0db3dab98ce303ebc919a32eeb9eb833c2e29c870018cec9326afe19
z3cb791838e63bb4a5d874a501056eec10831ca6b848b1546f2e973e8e451e06585c10e5f8fd875
z5b68698bd9f2b1082a26836cf12e235b2ac17976b11e0923035ca568f1c0fe184f43d4e93f6f5c
z59898d07b71a3cd6b0a86429e3a198537ca59f6b0ae88a5bad7bb6b55eb58ab46e1ed200c66bc7
ze01aa9f34f7b1cf4b1b5f72edc918a9f9b4346f146721abe5e250abfca41066e8d9cdc65719eba
za11897a532cf7ba70373de2da29072b3083c3ab0949377cdc6ce1d4e35115b888a3889c93ef162
z55f24e9fdb61730bae4804afa35f4b70190fec58b51620eefe0a589bc2671b4f00b01a18e9637b
z1e3131ac03413694f69ff038098cc7f03581e98ddb2a859ee6538e44c52d2a3779aab111e2f7cf
zef3a11b3196f6b99c2b2779878f61db3be8690b08eb4049fc41bb554c5de0a687926209f0c55e0
z8fbe85b38220f3d37f2d05c0a411bee00d62d25ef41ec42ea01dd7c119545e12ebd5db39bf0c59
z26baa40d7cd0c607b308bb0356635b7a27cd8186c89091154086f798ef69e266b394a2c4f63310
z2e3e11a58ac677eef5b44da58931302067a5f3f203c508dd2a20c3851453b2a93af0caf02979d0
zac622fdbfa7ecd95b2b9c561664ddbd7f1d68569a1c93e1427781ba48f8a13e92971c2ca30cd98
zecfece5d3befd65d926df4ef1d1c2abcf0c8b99b2cf31c4fde8fd31e365e2e42920afea0444d32
z495a7bc1c2ed21ed30dcb3fe1c82b0e8b72c4dac22cdc89d8f4bd4bf35324838f1ea6541faddc8
z4cb75ff6cca7dfffbe5e68ed9cd8bfaf9e8ec9a4926273b3db859af2e50e8953b3b6934feef906
z1d6a412863d001d4c3082e59b10534e056a295dc14f630beb9dd5fe2eeb05c5a8ed8116439c920
z27c1e6b56ea5cce040a2d2d15b03ab6be1d7c65107e0b8d9c3e8c610489ab4deab655d10b41cfa
zef49263ff03473a3bfe012840aea7939d207a4772c0a54808cac459020d220ccf3d84884764a1d
z96981c2adab6f408478156593d1548902c6f1fbd6ccdf7aae6b78e8fb24e01a28ede0f3bf9626c
z5f323e4558be14b3acc4d4f052827a2c27146a2f467bc4b8eeb7d514a2eeda71b6314de6430057
ze8969cbadde142efc752fe15aaca997358c411c985dd5777b9adc56ceeb39c3aea1ffca991ff2a
z441bb41b21a60d2841ee208e4a33c51991941e5b7f35a9f61899884d6a8cedd4eb89c67628bcee
zc2390e4b0be7e7dc258e6d0232d7b3237461d530fcad758a8d8bf985ea06c4c526406374d592d9
z8a3a6fa22e6eea188976ab6913faa77458585a277acc9f25c76b65ca7be5918e40929f416dc2a2
z3568e19b515334d0ee1eadf17e60d1ec36b7bd9e9126e3d924ccbe0a7a7ab60b1e16beb33a8200
z68b821e60e0103d12cfb278f8546e0487623177727997d147ec4aca9242a403baf5922f5b4e26e
z525749a365772b18696b508d328e31073be5d3889e3b2d42da0ff8ed4dc291e0299d56ca104aa8
zce468a972466e96dac078c03f47608bcad42a6410b7369312298ad996fcfe74d410f750f86d977
z8abdc19a19612a8cea19dd29d4dd212a8e92e2cb35694a142a5329dd7f5a9f311528fe71c2047c
zd8e20ebb6fe52e102645bade199a588385c35350303192ff39fe8fd6219e033c799bb500871f04
zd02a5581144f1bde2b07748b93292f9d7dcd0f0e61878cdcd5fd4625c22d4fafd79a230b19dcdd
z97adfeb6e9e176ed0cdd6d37759542383ef5f9a4555bba68b4644b93841b3561ce563f01d31742
z235b73b46266bafe26ea141463d5c7f01aab24176cc965a4a8babe9aa165c660cbb055dc7f492f
z1c908ca576fe133d1edcdb0276fdd0441cefb174a7259b50c0336db7bc2ef2a8906e2510cbecbc
ze630782ed26fe59e741192a9c5af42a40d0bec6c4b2c665b3a26e865c97926cf0bbcc6eff55260
zbac932d74acffe140eb3e92f6f42d222a4165dd77b10a059dbbd7c67514a44d99a8b0bd4b63a3e
zcd5db10013a9518615f1a8bf4514df18bea85acf43bf1ce0bdda494b292dd96c88f6d6fb8f443b
z0ae076464480eb314d7063e9dbf7b33365cb0ab91aaf4da7574bf6a41f6e2b2a9b0fe3a646ef8e
z2f462d1db686d544daabcbd4965caa767c8de872bbf28e26237f464e38db786af061ccfee95b1d
z60acb6e4da5f0c7d6e29cf94593ce2c72f2b9154067599251dc09163f0fb2c7f151cffd433ce2e
z9e7e65d8fc493383441be2be5473591a77df784ae70f1f0610692d443ac20d1731a1c0bff9b781
z4755495ac96a8634618ea38b46bc509c92dab6b5f54d7a5464b1a88aedbbd057ea0d1e340984c3
z5e30f59a74e71f45fa431302a208727c85a212b49095eb3538c0b274daa4c7453d2a27dadd7af8
z2e290202a8488bcc85e00c9b08ea191be02e2006cdb224bb4b12b390938f5c4f1b344c213f69f4
ze537a03bf336d13979e721d019669d1fbad52c774f058a7b1d3413ef84494d9fe4ce87cebaed05
z776e7891514aa3b7093bee207997620ea4f6ce4b0b38e4449ac6885c4932508b700e36d3c911f6
zca614189c285ea77adaed1f282a300cb27debb7c045e04cbb38747394a4ecfea8db40b9f653ac4
z12bfd60470a42172e0150f866b22c6e64d7d0f85690ec6e0a4273d75b4d18d59cea7f38cf1dfdf
z61ef31e906a37400b4c2c27c6ead68764f3e3566e10df15d73b48749a1a7cdbd6daf2d6dc9fccb
z6b0b0d03ae9a8ab375d1fb547171d864285518348476e82c9e7c0a370aa6bc51bf9f36f610eeb8
zb3de76515a4b3015bb425a95a39ee027843b429985f18ecf43237a7270d5f77757734bfc37a7ab
z369e5b7055fcda1d6ac2beadecafe5c97037e434b1e7a8f40ec1611bd4715c8ab15976c5324bd2
z59dc6d3ffd56bd184baf827b4fa82e271b29e92188f0f2d34bbb83d7c6854167fa95f5e63f40b0
z21b1c12ea383507143e747c3864b11894bdc4f41deccbe4221b7e133fc21b726d3a6700fbf4c94
z3662a592c5444f072682010540053964d43d6d7f1e27d09fa7f1fafcd6ebdf07012d51ce1ae645
z6103d98ee37b8821d668508f80f7e96650fa08cf188b10c638c33ee5780f2e515d31aee1361bc3
z7c39a52336a2586f02bf910d994ada7ecb4b3a9db3086ad9574fa619ae128da2ca8bcf103c21fd
z223279d8e506cc5a833a373230beefad01bce465e4d88762faa270a6545d143906aa2785fd6b6f
z264e6d08469abffd1c65fcc3babece440d6074f17c64ec85fb5a5dddd761131154ff4b7f6d95db
z99a7774fb9a383e855f2e13e0d1eccfaa223a9dc94092a6538e63e64fe3be28fcb34a1f4c71a56
z49d5872d968683e901505b273e5b60088c320e6ec9b6e471367b06ef4462645ef237be08333b57
z65bc910385351d0c1c5a452b3f9366e2d39eaa95f2ad46d88da0169c9d985c5aa5ee04f43d57f9
z5d82e1a762d3dc7bf2de7618ffed5b5208d0ede0341a4b70fc38fab82e3c65b42e86bd0a265a1f
z7f7ccc312385d2c7990dbeab6e55df88b59549a5dabdae70e62a89a53a995efe6fb824ce2117d4
zeac00f77016f8905396a14a9b2ba17358c47b5cec3d6f5957f6fdd359c3ca79008d8259d1bd306
z3d7ccbb859f9163ed32dffcf8b91b7210473853a3a414b82fe4d7a8de2b6b2814ad86aa1b61b0c
z74d3fe29656b00aa2eca9d4d57343800fb1d1d0787d6cce09294e60f8e7647bedd5095f274ac74
zc7f9315dfa88ddcd06878f194c5e2434329bd07ffbfefcc50f54b5676c6f3477b0e814486afbd4
zf51ead9ac80f9496ae39c56f68b80e13d0846b1aa058530eca2f591810c84997ba9d83d68c5657
z98758a0f3e786770a7c513b1333e1adbb6545ab13181c0f1433780b32e7d79df2b99ed65f0b0fd
z3314be739fb9734e7223080fb4be949e3c3e3436563d4aff7ab33b6ed6c1aac876a41b0aeb93d6
z080c8f35fbd78a0242e7b6658a11ebef1473633d84bad8df028bbf0a521ca31b4d704432679b18
z4c187ae5d7595ed1914ccc282eac42d27a06e30231bc2ce9677bf8fb895eea97e17d1c27831fd8
z71691a1ec1af07fb71ed4c0cf5c514a960bcfae55aeb8533448139ef9067243b5f20cceccfa21c
zcf98b3d389c7967ac9d3dd1b00ff5bcb1f5bc6c7fbda8e093dcbf6d85ddd9d4e74857a59b32b7e
z12f8df31918eb34e12b5db1c341a7e9cfc43c6ca09520c4a9fb668195631518cf2caed66e40b63
zf1ddc8ff79818178c56a3409eef6dddc0371a5af9bfd8de2d87da787b331aed6fd8358f0ed988a
z2a6886d734bfe8c260a2639c61a233fb1d4a6931e218575859c06456f55a1c9b8b59d890b3e81b
z0bbebb0a973bba0e6c3434e1e94b1951078f92ed920d1802157eea53face3467b7ea0ce2eb1e6f
zb6fdfd523c94d94ef1d4fece6db6ed0e71583406dc554781d1d4978c9f52aba467e87ca75d2772
z0af5fdae3d8842a65f42980ea03dab78b68faf62baaa820a81782ea42e1b38ab774d96695fa4cd
z29d6474148f826642a5f23b8f13119385cd7bb52580f74c6494df6bccf262cd41103711e6860fa
zbd1bc826b3afe4e3ec60b09b6faf687dd8755c1a4648d07c1a6ef11ddacc2def42cfec48a24116
zbff7b2aaac40bc94b001a20e76d038348afcc56d289821f6a61ae20c6391658528015d2fcd2eb5
z2fb48680509c31968e5ae0e79284160077eb1f4c6c26a8786659aef87d4d0495ee104ee58ce946
z9f19b7068c459228f955541fe69f3d14a6de44f4943d94f41a9de73a01b855fa574fd61cf6811d
z1943ed94572a58803b4398bcad24fb643be3e610f916a2465ba6fb1bc059bae4f8ceaca6622bc5
z5925f87a2e3236bf81a322590ca0216e230a7f3abdb85c7d89c951239145bec7f2099681dea7ec
zd9748259bf6d679eaa5c54104d0fa808d75a22935b8a6946a70c637e10de6c3e157dd009bc0a4c
z5896c40e8a4cca8b18d9f90bcd2ab969c8ac16241fad059fe75150f0d8621b39b6f5b8176e6720
zb39f2c4d030de5a2d2e4d53ec948d8eae13e8bbd6d10462fef9e3f8604b2877af24d250438a0c1
zf0968d2e127f28fc62d61dd164ef676e4ea5ee34d7e459a1ca806876b7c5a4b9133cc5d1c8613d
z9066ebbe457f153ecff3c0c01bc6f5834f4bc0d6eb099c225efb0aba5de0a3a9698548e12a1645
z9626971d5eb648af6c4f3d8f1dc3ef6d7fe5c6c3a7d3612814654ddcf9f2a3406760658d0c0617
z9119973bcfdd5b0c1c11d370b6297686217f0fe0356426deafd582e287b7dc80c930cfc22fb19d
zf8baad60a056d4b3a6d4289632581b0a486bd930ec084736513b1c98b129ddf0c1503f5db29ca0
z5b2a80abcb406de1c9cff07792cb8ee14e0d60da6c2d1d43538bfb5a84ef5b2a0a1a5ed58e5127
z68aa4c6cf0127abec7e8571a44f8cd907d899fe9ddc3bdc933552b0a432c985da181b765a877c3
z662f4d011a947bf48df974a616b3eecaaf2895f7f3ea95ab84cb441726071243a64526c5fdc8ce
zc37d2ccfcfdfc98147da748b9b119b1db237f2726ed5173f8f29079170acd78948e4b094534ca6
z578d62b87da079aaa4e99e25abe5198bbcd9b9381d32248f73ed87f226c1a1f9eb4dede4bda223
z4a5afdab166867207c7696bfea8594f963a9adeeb8571e64f39da5f87c1a0523bbff5cf9d9e74d
zea52f56bbefe4f698a315b6eacade507d72d3fc86571b2ead1590fe59f35746a47a285827892f4
zd80c92383b57f42b52a2cfe3685b5f0b6ad1643008ce7eea3cb6e3ef657e7640eff8c7fda4e631
z81582a6a144ba891ab93b2c1069eebe9e261fc97e500bb3ae8ef4cb0a6cb91a7154fab675329be
z136543a34d550dadb4f631fb169d59490c9aed9449302a256b21cc106aa0cda089b238979740bf
zbf8a2220da810d2cabd014f59ecb0b54fee08ef861b276a864162ddc5bd0ad57134ff6c1e5d1ed
zf8454edaebdeb6636390ce5d9e6a1db970dfc214d709b2b224a521222855f20e8d5c7376496c28
ze28b2457cba24e2182ecd85a9354c82e6027d43ac73c92608cd62288bb208e1f8fa605a347eac6
z74222a64e999af4f95d43e052d9427785cddeec490d500fd409d08703c14634ecd76823f075280
z426b28bd99f0c86a14856bbe791ab6b69909fd8c044d95d5faf193e014ef4153cee1bf0195bc9c
z0819661ea8cf9c7a8c108cee577921d9b92c908e4d08a94e43a26959267d227094ac03ed8be2bb
z3af26f5896bb632ef2758da68c16934c5fe7965726c8eaaff52e33ba0564807b483c15f51300d5
z71362b8d2442ee28f7f9cd2f491826f833840fc6f037c0dc2a850a600813f009e6296d60f4addc
zb50a04c7cd605ebe4402ccc6c44b9d1cc0f7ff9f7e1b25feece1a00907117d27d520f67dfba99d
z2b61fd5a113debd7a0454658702a354a0b14a9318250904ceb3eff4344a41f5018b09a8eb8e6a2
za4b28409e681a13f8610714ab65d3f03e4cd903d3546291bd4ada64b254747700e0002c504d546
z3d8d3953f1d4386940bd96b48290d69114d6fb10c77e664523a765fd70365432bd2771c4b52026
z916bd589e51535dbcdaed80d8af36160d60c434e4564ee39cfce0b6d0b0c91973302d5c00f07b9
z9c4249ce013423e41422895e6ee1df73b03ff74f86fd6c0afe2a01c78f601c8792f1ebd5f887be
z83fa0d9a69512db1a977e6a6c4913be8d0f5ace636023cd285404a090b17120315ddf76a39037a
z14b17c890d04ea5631bec6bae2be8b7a856c3652edf05e6587441f5f5595369ff674c3f54e2bff
zaa7191a80a8bec4ddfa7ee863366446de76989f76620a1020d21005754d2ef911fbdc3224d1a63
z5c133a521e54b02d033d2d46276913d377e2df7c04103bcd42f776cb19598a13bb5fedcc5bad2e
zd259a73c4a04d8774f8b4ec3b269c14933690f17be2034a0d8e6151a351643ad4b686fe9fa7366
z94ea1457794e6cb5ecdebee6d11360f7848c1d714cf22ed96d4c655ab1a7317bc1b113cb5964dc
z9aef44133af272c91d491e11fa7cd2475e07bc293899fc79e0a51e63137db9a9ada38b0ce705fe
z22ee0cb56e87d9c85b096a17ad7a5c13f7a102f66be4d8c78a9c30c82f15629d09a35150a4ca52
z41c13411bb6167b23b9779f98820aa1dfb062559d98c390a55174e9f2eb18ba54aa9e3f2ebb30c
z45686c42868afb2e5ac0d15c91cf8b27f892be946756e32825c59c1e3dd4e63a6cea6ba0a9a217
zdd3f038d857cc8bf157b3ccdee35d6c4b6e14d8e72d28b6600e793c8ef19b5a3f1900f06dc1690
z9acd7a42b6f49d0ee7c43a53e624facae99f46bfd556c6725c0b980e166aa5769caecb9cda3824
z529cc6a23606efa01c5cc67537da25db09e39e57951bccda729b6a1e3052d934412a453439e3a7
z4b9adc152f98812d11f4c107de995099102e345357e62ea87bab4d362f577d1560a24a3f426fa4
z0f948fc0a7e29d7627d1d91dc0e01a27dbbc5d00e1f91017079333314fb5add90183189cad0b85
zcdc99b008335dbb53c559aee79922ef9baa0110522681b20498d55eed765fae6aa17532febe10b
z531109ab512ec6234a6bbc669a86a3698ee2930821a8dc8b5ad0e08a976e9796dd03faabeac43f
z452664eb9290a30d263ad7fa8f19f046eaa4d63245b7f131b4fb5e13452b256572faf7e0860736
z4c07fc937782a9b719649a76537f7aece3486d2e2b34aae55072a5acadd57af8814ca95247eb25
z41ddf0eee6ebf2239aae2bf913f2262582812a6dbaced3ad878d11036a39d12e955b7113975264
z3a5df08b618f844bb85f2088e7a8157fa1c5a3c36390cda9235701a4fd572aa4f3aa64e6a8256a
ze5de18c98021bea6d023d1a4d868b4e99e727622dc2e214da841f7dab7c8a3481d3ec96e878c21
z806eb3ebff2ea738588e82e3392f7a09a6f135ba0e22f175422570c7a6cb14125f47750ba0f347
z0fcf94c021694deacf11cf62a69047849c1f0b5edc31451a9ec01f74868c77467c2e8d0dc08296
zc587f05db03660b7533ce2689a68e51d4dd8e8f4843cb4c489539b7774f4fc9bfdb525fd9204b7
za1a4b5cbf6a6b64e6fbab2b2608c02002ad2d8f8e6f8aaadb17f5419c37566d8868b3a0ce85a32
z32d53c907ee1451ed4b666c5bcf4f03fc3ac66b5fb893d494e3836f3b100d91516ec87ce600327
ze0dedb13759b23cc65f6bd35929a1af11912e704b19db79a18222745a28bf5b75babd5aea8954b
z71fab8e9f9d975a18a823f87ae6de5b2579238c1fc64d5ad52b65ba8a3e300ddaa63c90d3242f2
z268ec5c76d42ec88046c8e21ac4433f06f4b3a0f9569313985e96e31b144d7773574af4a6ae548
z279d09a599e433bb2a55e788764dff86b8b6bb5d7f12a1c311ffc57a57dd13451b2570135af101
z1f26e94565480f177cefa68c4d30870f319ab6dc1fb7d9020ab055c479dc072ba5ede428268f84
z764e2a4693fc3456237255e99a2cd012c3c3d0a9e26fa79ae81ab763af669b39d3387ea79a1cd7
zf7980d453663c5b2a0873ba0942b714ee306f6c51698a8b952c0f103bbf8e4e72c2dde05f235c5
z1f74134d0f90265b3beb50f9ac42426fddd6424adc52ff1b2868c4d46d0d2de8bf55e09666dd6d
z399368d1ba9bffddcbe2bb501f7a01aed572f2574da3763cd37807b182de68a99cb13c4711d84a
z5399754f1e8e76adbeab98838b778f05a306e92cdb7e41b5ff01b0475bc4151503af7847843670
z387c5664e108b0c4dd195317f5f563e10f02364cbf59b93c1f344dc7ef381fc63588b3b6148cbc
zaff437352c383ddbe9061aa5860ed08d198319c0e84628b9d36fa5b6240e120eb00414ce7dd4c4
z0ed9079fa3a13b2e7fa260fe201732432eb392b5122df8340fb39f70ad60a2b645f774fc83c205
z0f4bad8d9f24efcdb582d076155efb8d094564ba8ceddf7d7697e829d8fba0ed5929bcfa92457e
zfc3838698c8fd62fb4ff53894023b29ad48528bad47c17be1851ed4ebb1934d5e39c15df789c36
z8ba895075aaea40eda853230bbe3c487dfe79825c2be4dd08be5b4cd8a26cfa1e75ba78d1609ed
z314cbb98ffb2dbae08003b9d528b1b0ca3857845974edd44a9e3bc4cc2abd60c321dcf9b745b85
zda56cb57f99454ec71b946e9c6e58838497a3edd1e5ca76dd5d4f2d3561510d00cd25c44f37d58
z0af1c07382c35310c97b2b90074dd2ff952073d9eef44f6c07111cbb7084ecd98f1a511451be61
z7d3b77bef98013d8da704c83a9441a19eeb32d1a70dc3f8825a0971d0d5ca4bb2f197b0bb42baa
zc7629f88a37f76353afb41c358b86350d99c7316e93f3cf766c4aa7f0566bc951297ef5fc28787
zf107635f7b7e732db8558a50c00b55ed023529e7bf85f9e9b2eccc600d4de718cca9e58a662201
zfa75e2204d7358c609b6aaad609abdb0ddaa391ba90665d5765f48a3c4fcb32cb18a0bd6379e03
zd720d9d94949216d73cd7ab584a48b29539745c3f860eb4525dd7003c328ae074c46c6940037fe
z7c8785da1633f354d6a73921008b55e77010177ef9a39bf3ff192db8509b5b55d2b7187e287c11
z9224959023787f4ef98e5bce9e7a83445f897f268742f48979133ed4100ec16e309d233b346349
z32747ffebe4e8a82a57d85c95bb4f60fab9a5733dedf8921d26378ace9b3dc037a3b34411ab5db
z0e5f60a2804b453373bbb860bd767d5cb49c48696016c787244628aeea3843e3626d36d43a6ede
zd43e53d44f5e91db45a9afcc066abc80f42283d3eb3b0c8d329270eb984bcc8f7e0b1d7ea7a513
zb1bd97fcbae67847523375d073619960dfa40a2d77163f60a3a284d014e0bf5b10588326d20329
z3598e7fb99b3f2ae9acfea3f1bba752b196f68f76bccdb48751ee567a35a28bf82f0974b7b07ed
zd7987c40b7f2baf7acd1e875587613828ec096c4cf9c313abebf2642cb64e933ebf31930643f08
z64b51e4f87477bacfc8db2e30a81b8c3bf0f72de9a18d510144743008519ea1a9a467b4947fbc0
z0ca4779ba50407cd574615635fe9008ef40c1ebb6a4a28e2ba84faa5a7a5e5f34707a94d6a3043
z1333bfdfeb0c912cd5e5f67487424c261a0193655fb7749fa5947ea3de1de3e44e6b322538442f
z6e72bb76efbd3b6dd89c4d57d1e81e77e98e41aa91721490fa59f85ed337dee82852809c33265d
z59b607fa0f4915f871d4fa498d5d743657da79c085f35a15d83616db06e154e97cee7feece40c3
z42f36f11796983f96ae25a756d66c136142a9f09c59f0861ba3673ffef7e8dc6a31390d4747e04
zc0cd8eef217d12f5b891f397a8f88863d2812a4e41e09d1c1d9af0d8c8e5072763742fc23b0336
zcbbe426790fdd69ae8ea86bd42aa74bfac416f5fc190a829ae7b209bab3aab059b6e92792465bb
zb3e0818ebc9bf7084482cdb671bcef263df08c07780ab4ed523123cc2a0502f0b4194ebb2b49e3
z37b4a68b8078b19f8e97cab59c890e0ceeeaf6db42e2ced8638ff306e70402654595d127f5c047
z71c51b6232a8c742abc7280b0bd52cb8558d3ee67cf56db5107d8c6327fb57e0910391cad4f68d
zc9015a7c83509fd71f074cba120aa88de9ee1af0d3f746b36df2586991bd5709fdd063775a88f2
z557f464fa20a30f913b42ab7f54ab5f3dfb341b1a6965bcaf38e3c8ecfd0bedee79e7c17e6e03d
z3b8052efe689c5cf36a1388da884fee8935de668602b050700ac3cac16722851cb71a419588461
zc8db83db228f72cecf336973bdde8b63c22cabb7529cf31dbc2767d7e6512c5eaf87f53d679327
zb6d390f498aecd44234a91bd44cab8ebedb9174fda7200a02b118166d5371efc56d275c002fe85
zebdf44fa0b5c6bbdd5e306fc3cf0282b13a86fbaa225785b99df02d94c084c2797e042d7c85015
z6ab0d3844e314d99910e3e2db49cf0416e6132d593bd579eeafd25b02e8803ad6925247730dd05
z4832a5298870022f63456c57016f047552aaa87907f23ed1d43f711c47475c3a87079d7d8200b3
z894b86a69a3bcdb530d06ea8c91ed32862a69fafc6cd79e0702b8ae32d7967e9d9b6ba2b821a2d
zba4754cee6fffaaa6339286a65e6bcea184b3201ff9da99a24460ef10b7c24165a4e762d0001c3
zcc7689db8b2e26e604b930697521bb30618c89621aa1a6e07ba2865d21b5b46e54740cf743e102
z70fcc7f4be0fb3c415599d05d43b7eb797adb684cc5cf063f6ba3836b143591ca2260c1f87facd
zfd71acfb6d5d64cb634bb7b733bfb9d59f444c7677bebaa58630c2c1b7bf5a4a555a91e75802b8
z3b705ac088afc0e71c516b4af142e6d199f37da1dc24d6f5694a2ce1cda17b81e25ba05ad6c470
z6000567aa08e8d0d0e884b59e10cbcb499ea53f1aca5dc2144fd8ea59009a7e364b50190eec20b
z0161b238f1a47cc07b88db57ff422bf26633052e972a9f44d6d422cc306f6aefd629b1e075f1d6
zbe96277b12dc354bab26300021e2c022f3556e727a3ae8489976abd5c13839ed94b48fd9117670
z9a28ba8c2f4ff83600b0d1d33238fc530a7392333368fdad4f811e1486c8956c4af424b48a3427
z764723b60a3cfc3c592a88c8110b542ed9e6a927c2c3d42f452b9b1cd80e16b404f7f6de548bf4
za67abdc211d1b7e9e1248a415d83470b235344989740f4d055be4c7df661bc257c13229af50c5b
z9940db564b6b41fafc2f44a75d83ce29984942c8dd8f2e9216d734a305e627c29f7bf6c6cd2214
z3f3761c025509e3ec44a8b7b21eb986e3c0206de91be68691d18b1bf1fcc0b8b2daca9fd331c62
z11ba366363a00010b04186220c8c09343146bb00b1a990e1f86f27b5f8f8e93a80bde1f6c592a1
z00976775d301c244c66106a03813278b44ad126fe0cec163722d05570d05ecfcfe1ef91f9b48dc
z8b26d8fe7642868d5652e36b887a32f47064e5532abfca966df8e1cd502d12a554d2d04c7b70e6
z1246c0e9c1b43ebc8526b3a8f4a264b7c9eeaa71dd7e43753df34c33b45e6cda322148737c7fbd
z555ddf47ef59a0454af132ba72b835aa58648c4b3cd19d0861f99fc160ade2b4793cb0217d2b88
z6b4893ada4f0574f1c59910e15431e88894fddc8132696d995a32bb0f7bb851bb664ab275e5b67
z709f534f7d133638b962ca36a88414d3d843aca556bf37dcb02ecf9b832b69603480f0077e1af1
zc6fc0821299af24ed106d08c46c61488e60b40d56e83a9fd6c44373c203e94c2d2effbb523cd15
za7c9964eda4b44fabd63b3fa0a0d8aecfe608b9372a1c5cf938be7a05d977700cd56180508dd77
z05bec3bccb865a94e0611613de9249f854ccd073f936f4fb6250d3a381777c6555d292080d45ac
zbd8eb608789df9847a74b3e43dd24b800f33113b015f37fb99be9fb549e81e47e7d1fe1332174f
z3018803763cd1eff5c33b5f98df4ef89c061f92add5e53cc619ed6bbdfa8119733b2771f80927b
z14b57436f41622fe86a7ff6c5fc889f8b9e60366cbe36ba1a34fd304f5998e0b0e7124f2086ab4
za5833a751be4f618ff4c5c88e692f03d4f1495fe8d7c4e614ed936796a13530898dfd5809ea766
z6719ce600481c30bf6c346bf6e2375122ee713bdd0027adf90c3002adf06dff1627e16ee39ea4e
zef9d47e9851dd95ed9d9fc6d0fa24b691dea1758d92d01643ae313c9b8b9d8d8d830b3fa611c91
ze14b86180fe1e9fb669413512ae046f55ee980de730c34f5b8adebba350be06f19378db08df93d
z1134c043f5e855feb1cbe5e8f8aaad1ae7a388b301dc3288b8ea9d2e619203146462d62aecc3e4
z57cdde899cc1637f1086889407d901d14175b21180944d118c6cdd6207c2cbeaa546c12322c521
z404915ca646c16c342a10dbcf88b1df89dd4d2d10e8efe13a6f884071574837d4b23e46df8054c
z629532914beb57fb7846fbe0476ff8a6605eb3e9454fc2fdc579ed9697e53cd0410fe217516311
z049acaf38c6d11e9cf2002b4468fceef62bc0b5a63273b6d424df5e1ea999170bd155d8f95be8a
zf2a162ab8dfe41adf0368625826992a580978dbf4495b69ecad2b72ddbda004946831a8a15da4c
z01f05cf2a69658aafa8fd5c800dcef79353760ede38f3823289456b5b3c64ad4e9bdd863d66b36
z7eb2da75767cb05adcc32d918889371502d10a5c69302200b6a4c237e49b6c8eaa53c17623cb3f
zb43cfa609dfb9b9273d5ab9c0262ecfb2a242c7994864408a4cf4ce6d2d324966013cef7d4f942
z28f7bac99a2877d5f66c851a52cd34c429c53a70eacafea4171f5cd515e2d1222bbc1185cee56b
zd2a367ebff37dce466c9fa0bd830819b9e5ac04640590dd7e9e325e57c36b282d6c7fb05a1c315
z3f0a9fc008d735e481ea97a6c39095331be79f49e51835619d4461802f47fac6de9faf3419bf9b
z6648cea050774042d66216766b7585e63451637eb884d102b764b34473bc0ba8594a93b48394e3
zdf45f3861eba37ff8b7a6cd3930087a7ba94db8260774914a962eca62460780552102728683590
zc485ef6e23c051341d554cfa461bb7833d4491d5ed6fb1018734b032c1f7c466512467b263c608
ze3ed100bf7feb5428266747d85dada85802bf5c7c33e3520c30967f3a1dcda12344711f97a0fa1
ze15f69271200af4045e22738a71e6c1e3901d20c179e87962409287fb1eadfe82fd50b980be8d3
ze15a64e03d141bf444bc057458e483fa8e084a790bd597dae8f369e7e7692beb24e18022716fae
z25d460d9beeb49e5db608bf072fd3383b00c172d156bd6792db6b59e0d5694beb5ec970fb93fb0
ze360df9e6e5acece5f3c8863a52289fe7a8916d9593a41e1767ccea64f596271ff17b4f9f50adb
z4baffd5c0e0cf52c473cf6f6cc4a32c658360da2b9f9c67546a534e3d9be7d7e3dee7a8f9fdb9f
z959e2038d7fe18e30671b942cb267928861b10b83d0e65d4c3077a3a685637bc221ea87a8f62e3
za74c1a06d34299872ba740f4d5693da6d28b8c3e57f0f703a0c34f9ce7ff6d807096aad4b98819
zefd0afed5f52ded5948a266576bd2f725e02bc61868fcd79d8e7dae79ce7d69634dedcecb23b89
z0ccb99781d05786130892fc6e23d229e3f0dc7121a8f0755135581562c2592d2f0bbbd4b4478d7
z12b3d8fa3c0933f4462dd33a8ba5e27238b8f04ef422fdd92f2f4778ce097c7bc2700d02979969
z0cf0ab12c74e0b55654b18d0c65eaf9b87bcd4ea4853d5257fcf0dd588e7d675949fafe693b66f
z0bc7ffaa15806fb7b0c19d8bca2cad48b2cc92c889411b3655783ddd8eb82fdece6218ad95ec36
z7e43be8c8a8b4d3d558ca33bdd829732038623fdbc27102028f2f16e7b16073b5618369d2b065b
z69354150c2dad829a29be12a2f007c9bbbf2cc7db2ea893fbc700bef51885befe2a7b93be082a6
z276f576a60fe3a21946c3154b97813b078322886cca05565d716e2ce79ea6ba22d9861f50d6c4f
z6c9268e4a76a0e8cc6d8059a3135f19952916769341d0e354e15ebaa5b231102750cfc5593f07e
ze4eb18dd75e105bd3e7408c6f300a876e1f9e23d01d30363c0d15fd8a180b85d043510dbc8538e
z28e4fd0bb1beec505381339ca9f7a31ab6bcc9b87d4c0b0fc8f3293e1ea1aaceb41d61eb8e558f
zc47b99e0070f3573342be450ce3e427b829e1182bac84bca56eab6173457c499aa7e47d5fdec7b
z4b31de8ea104300716b01401845529926affca86d3221e0d347496fb17c22e2d56e32a8b23028d
zeb787560284cefc319ba8d1e9eb2b0e1febbb0782de2f7735b9936742d45a25aa41019c760899f
z7949275571018f2da6300328597c73985aae9a590df331c0223644a3788b14446ed82c4e5f019c
z42a664ae24bde95c38e99ef23cd17e99189ad986368eae0b0d4319e676347540f078b560038f14
z00101c552a493eb995f72adea3ddd175fa77c21f23352e6fb0bbb19654dfbd1b349a6e453176d8
zfeea76f32588b110af240821715de331358402ac9bb6459ab17641f8e37dfdac1f7de39427c108
z8a02b98379e142f5b211aae3932673f992b86b9e45b37db84d684383241fac1419315334eabd27
z48df6cad29f3a61e8b440ce5a10447ac976114f6f65c91dc655ad6fa55cc9c4c2ef492837ba116
zaee147a1803810c0f0add22164bd66d05b73c896e1ba89a6d39d21b4a431b7686797ff555a2485
z3f78f86cca8c082aa0105500871f3e8ab1f3dde5ea76ffaf5dea42f135e51b8b337e7bd9bf71c6
zaae923c555b994fda970d9d81cbbfed196954d99489331379be8f741e3bdb06c2ea08d60761415
zdcb4aa04166cdf18ca8e998d788003fba50af939105855b0ee98b70fc9bb1c137200c79eaf608f
zdd448c7ed89ad14040dda4c22a418e98ea300526e9858c7301b95ed36cd1a2f31234568a02f4a7
ze37c72112f5ba1f30a6ca972215ba389e05cf5bb5c88555befdd8ff71238a33611c2122d0523d3
z5acbc7b30ded49e613e040a29bae9337acf616d95dea3e0b7e178a070154c5df3e0baeea3ac2cd
zd44228f0aa0f4f8f519d55ebea29acfde3cf15a91f64a36970d3729f59f44423de7b6f7c1cae24
z784e755bd1ed442f88e9f70dd6fbfc8aef12ef706ebf94d7a4b7f6de472f4f82056a4d5434c03f
z7b7c5a15ba56bfc9718fd86bdebfd46e832f139f2441b0b551584f924178c21aff6335a14aa168
z8308586d3c96713db4a31bd717b82bc0e15be2462b524b1aa8958bac1bf01c069ed2fde41f8407
z2381e27fae927206
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_express_rx_lane_receiver.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
