`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026255b1a67613e9d37e4cb6285056
z2a3865dd3d7f5f2dee8dc0d96d90b314bb5e4192fefb2ea90129ca1c488110fa91a0d5e66fad09
za69199d8d5d6adbfd86b99c9f9d957ae4993d8e0176004a73e7e01aa19ec291ca4fd53955157aa
zb3fad11e63a96ec68408d8b10159ee1442d48a983b3b26963a12b908efa5f1b7c21f34c589ccf4
z4af08af789ef62d9e9daae5d0698fb73f8791a34b7d429e15e7705873b9789071021aa1d5c0be7
zefcf5762abd9a379c2d4c4b354244e003ba0b1ad8b9b211d0f9e9e5b3b649b85a91cdb7cabebd1
zb362f659658bb02ae3e1303b2904948346f3446169868e2cbef9552a347e3e4edde3f6aebee5aa
z5439502afb1aa1e572f92b73d4ba473dba357e9fa9fea8a0775baff966d555fba08459ae2c3c1b
z6e8ea463b8ab1b458f732db8105cebddc8f96745ce5a1e2339feaaba5985fd28e97ffbf8226c53
z3980bffa99a9a933b93d660ee8ebfc05fbf9c62875956ed26dced7f430937ebad06dbf4840c670
zdff9b327abc7298c5a59768022d4a2bb2ac7e170f5bccb179f1edd6ba4840c2d3a35952aa15465
za25fec5a8f99b2de321394f2832f948f6c5f3db1d307ea9561d3f0daf1c137488d53a3329439b4
z1a1d5897ab07ad08128e9a7a3b98da088a74daf4343622fe87658652241cf97f7407b170d4ed90
z844f51ba353984ebce00a3bbc3e7f5d89b332a1ec2891f4addf3a565929510497bfe55b0048f60
z10f7bb847ce741b22f134cb1b9bc95822c5e91308df6d51b4c0ad8b0efc3c871e06fbcce8f71ae
zedcd6b9f173ef32957c2a90f4430abaebaea7997d22e580d3a5b798194c1e5944ffdf688419ebb
z65e0a0b3784dc1a62287e135658907588e23afa33e2b99928f2d6274952cb044dbdee4c24e7c73
zde1ecd7a75851bc8726e7678ac295eec858bdd0a6659b74266ec7f4af16469c84bcdc620844bcb
z4a4412083a0905e260e19544b7f6c9a1b323f8effd92e98ccd26ff56d133f5b05cd6a70f1cd52d
z92961d188a60b3b8456023668fa540b5199a17f97e8d812309e67aba0ebf48d8b067b14c366711
z170bb793f7e9e82f784c137697a18047c791e3b28bec000e9cbda3663648348e09ad04f0c15625
z925d11a47bac842e7b5732e2a5d548a87ad797617568024f479c90e802c96a57b07a7cb9e8dc70
zc0c5166ea8b32fb8c4bc9f5d764679403d8f8fa9b60838e9c1c4683e912b0a7b60f7ddb6975770
z5967dd988cbed6a67d5a4d3879f1916fa55ab5f0d5d4a13cb0066895f1edbdbffef5a5724d0426
z0e60796c2505869e211891e6965a76b34265de373757dec3e20ce547cf78e5d3b368d94d2bcf05
z4366443b7a6f2c6de235aac79a8a0588b69ba42d742603ccc498223a28621910352b481148edad
z329fcabe42f1f14fa22a3fadf80ba684e859fce72c0b5cf727274a8393b269bc0ed006684adc56
zd29d9c1192f4c2f9612b79e74dc76cb2e36a2163b2320e8e95e573caddfa16e53df1dd6bc3668c
z8d59e3cec2dbe0733b556b2d3bc8b70d3a827bd3367e22b8a4ef13304308ddf859709b18f65528
z724670fc88f66f1c23fa2ec7470734f2e8ffd3d234a4f197a4d393cea17908195a05e907d4c8eb
zc237e3d8242b9c92b8182ccd5a6967ed493da15e2f62fc646f1ad908c2d22fa90b7bde4cbcc93f
z51d7559dacbef63778a2024ccd74eb24ebcb9b6eb253d55338215a4730d7be1ac2ab6a4067fb9d
z94d5288ef890b60a8486dec91f6b56878736e0304772dced8c4f8cb66da29b6950ded5c1254726
z08da1a665990059c072566beeadd52a648c411362a2df34d21661b57c9d6f7f9b2543c6e5ad89c
z83fd5c8ae59a64c2a1f2dafcc9b0c7b0db1ff508efd3015d388016531d201da611eaa5e960970c
zc3fa4a982e8567e8088a6e6ea6d7cd871eb7af2fef253f75437690bbb3075037fcf161147ba2fb
z002600d8643f33dd3eeac3c1279d69acfff5e2398dec31137afb5f5977d9dcb1d1846b34520f10
zea76f34c10e9799296b45705de551bbc46331fbbd2971d1454f0aaa4de71e4962ee824b1a84ea0
zda493514b558572c7293d10ed74a8628d7149a3f529a75cdcbaa0efec50edf0890d90c9c922ef9
z6f8b9e4b1c8c0d4ca1f155a41dbe5d079ca6b2cfeb9662db1262f289cb105dccf6d767033dd56b
za9611e09608d243abd3b978d4195dad0c01347ad1c046b7f3ef71970b852f9d92f021f2d8d26eb
z8d9f5879bde0903e2d86fd2d9143b23993d161e24396cddf816ad6729c50863f4ff5e1dcb017d5
z9e4f27a596177d936e7732609f044a4468a9fa898ef91dde946c61ee7b01c121f9a1391ea9e318
za1605b1cb69bb0cdc7211ef9b5ae7520032c491ed112265f565f5c3b05fcf39f3f2cb1638b983c
z75397cc1dfe06a12220463868e94f5bd511ca74aab2ba901c240ca2d2f105b72bfb14ef92484a6
z966dc91b5a62f0385f711c053d2c01c9e151822e5da183c4b80e933636e30325085671433dfb12
z63475d65eb784f49b457146b47927ed6a0360b21189c93469bb00fb05d5b10d0a43b768d95aae1
zf701f9277ee24c9730918c7edddb5a2239d933c3840c203b1aa432f029a3a61bd044c11eaf8bd0
z96e83e63916dda346b605d31dd790492bb52fc925cc38de7e7776833021b3faa2292eafb58e036
z6b6aebffeeb4e7a844cdab0af620bc75fc3f5ab36bc3de8e433ecd2ff0e4671601fee2bd1a870d
zf8cee53ecd28a2ae533cc9a10141365ae4d500a3d6c6469b99b896a935502715ebb0a86c790628
z25529a3eafda0ce9537fa5e362858f7a8c114abdb1543fa0be492cef2474c4eca30ac79462dddb
z143bc933d3e0bcb9296e1e4aa4130765a3351e2bdc8c2a66af6f4fd1583824b670a0695c582458
zea28ef498186ed6e60fd59e000c77b4273186c338573ce3ecbbd81952fc78649d4e8ea4b47ef7c
z66db95c6d22ad91e2cdab358bfe2d2dd10d97dd9f2c57f189780770e765e10fb79b06be2abf379
ze8231fd8d6047ca90db216e9b842763cf02b1244ba6851576a2ea8897a6eac934efb8b2c5444fe
zeff092258b0207928ec385258718bdf2437fdcddd4e86cfc86d2f62e3307d3a9bedae66b808486
z683622eb0f7af62cda67f849695a939d8292edf2f2c782a6ef657bbc15d6f65971bfe89fa05d7f
zac65ae86cb24af13035bfe1c98338c788fab7cef376568824be26deabdd89275a70c0d4735a4ae
z0d36df55a76944c384a8e06ee60439145e4633df7619a63f51d9506b0f966094f0a5f7bdccbd11
zdab7a54459c7b7016174b806913089d8f3115b7ed4d0f2e39aad40e7711ccb72d425d58612f07e
z42f429a439a60e1d96177b72ed742c9bfbfa823ae3c5b6c197cc4cb87459f393f5f8f56c1c1ac0
zba421c19ca1ccf0aa59def93a3ba4a26106ee2a3bf2b873eade31488aee6f81775b9abfaf863e4
z1b74c07cfeb540329ad2ac43007c94bcd1bd7afc0c173c5f452356b591716f204e138edc7e6558
z04db99fbc6319e51c04e8bcb9004e5adcf213f96add8d772b5e2b7ad8127a77f39c8c9ca933907
z2adf6e22ab9b09375dcd7aafe3b942a365f970016b2f5d95e94b691154780b682138b66afa5bd1
z741d40388a2946eb7ddd5eb18d61fffc81e3f91d994287c5c3dffb949831b5db6a938be3708acb
zd66e2886d916644878b3fcda336615b2f827624cc30736a5e5f4356ffbb967da2379ee74ef2c32
z6056c80cc293030ce7d64e8dea6272c450b8e97b5aff205738b32b3f73985fbea0ff252ef7acec
z7345106a2421e66400ce843e070704d2e6a126c37ec319e52ff15a18bd34bcb016c3320a91dc6d
z82332979a5bef02bd7f7ae69559b7a200a583a9b8408e351bb1b07fe75946c9e78124823255ab7
z786cf785e8f7858b11d8c464a563ebca519d8956acd10391c76565a37dd67877ae7be33d622c94
zd98318c729501d419f4c4a02fe229d300c5a634d64c4b53c73355ab852dc69de70ed3efd35b7d9
z203b2df7b7c62b82e534d37c2c485496103663cc91bab0e18c76799c05e8a3a33d611460d19d88
z1e7f96126e9714e036850b66d625254ae60698780232e16cc173dd82ba6ba0647c99d78a826192
zf5ea8533d608b8eb2cf4236efd274493653b5f508e9b519062c9e078b85eab7d03ade5cd60c2e8
z5096b60d4202186afab510c36bbfd5639f682878ea0213898be20c41e11f592b29fd68136a8257
za2e4c90bc5e0c2bd043ff421cbf05991ea4582b52c2bc672ad4f0be2295808cab22ddfb862e0f3
zd77b65505c592af9963bbdf98886c579064ff08210455089fce1e8c88a54a4f5075863de9f2966
z2e3ce72bb78209022ac5d0fbfb053448818eb7ffc56ecdb99495358abf2f6d4da2cce10e3ef98d
z67f98d6c36de570aa61d7b8642ae8dc9774b2cd02de230d69b7da9d278576987bbe9b6c7c0c1bb
z242fc482c4e98b52bd71e9265180fbdd049f850b4702b0ee9bd520f26dc15e6d7ce2feedd6bcf6
z55804e63936cea5c6b39cd866edcf5fb83b0e8c467b5ed1b15dff641f05f40eaa86d9c3decf1b9
z39277bd3dbc2403bc4f5c2b0aaba119244d8477239868cfc0a37c3736c114a58bd4879a08a25a9
za5dd43f0b7ae15dcfe5ed3baa9aa6d5e9e5e70c7f7572bf6ce49e778d688012cf340bf097ff4c2
z58edb35d4f15a069be79134c9a60d8ce415e6a5590f8ad256b0823c0eb5f0b3cd2ce4df471b9af
z83c4ff78ec6d6ca42e1b1cc35ab4e097da7487a41f6de06791342238f018e5c62508b5dfdc5898
ze34af96ae017d73b8ef9d1b549e80221ec0e119790752a3c4b1ea1a03a4633bda04f48f8afe5f9
z8b20392c7819348a57cd8771be8e2c9fd8c2be47fd49d9b9315b652eeb723d7fd92c734703efa2
z6512c8d77a00dd498b8d014c64aa284aeb0e7f7c4280e21aaba3a855a802707e2a0f14906915c9
z6d9b937c69e51c07d38107700af7a4ae65d64d83db23f55267c565f6652580265d5dcb7e8e4683
z04be09e3afed46bbb10241e2876cbbf06324c21198a4afcd6d7318c830c7f354081fd3ba0da92d
zd785bfe6d50a14b13a5141b68e67191fcc066f95548892fda774a2a9751bf805d79847b210a432
z66579d794fad92721e77d84ba35dd26211d4a0169942a4f71c29f30111bf3a7f43160b960ca922
zc7b21c7a577644651059fe01039031fdb9960b8a04831b29f9e906b0b0b0e53517399645f220d3
z5995eaeae9c2c04fe56f697ba8ec048100543d7f9235ed22aa81b92ddef87e3ace35871a82a86b
z7d1856fe121c97ad223c69fb9a9f5d1bc40d013b9ade06a47c0cb3878dee9141b7f34a0427ee79
z29250de75d0f506931fc6ac8a21b5aa1125a96a94b99234f1aca858d27dda92c69e44d81daa62e
z823c4abce4229bb8fa019f44558182acfeefb5fdcb7b17e1327bc758ccb7c3ff443e4731a57507
z63cd15c915a5e6264dfaf92bb08b5ccd727679044e14408eadfa343366f9ffc9791afb434f1f07
z0a08c7ee32bd490828ed011f1118e32291ff1fe88c4e0ff16f888201cbe75c7a1c123a2bec3a6d
za7ef7611cf1e1e004fef30e1e2aaaf5c862a3c339994ec8ef388225a2616af06e12ab525bde589
z46147a800e6f86492932bc7f31c9fc37b73fb7bbca52d3233bcfa3f80a2783a75ab6fded0159f2
z50803853139a850ac643fa1e630f2859b06c378d2bec9e9f325adcaf62e133903a8a43b2e10920
zc1d58b63ba608ef49feca2d0a0d60da5f0e713453de4a2bba8f165590a7268a8f65e184c5ac7bc
z81e7b389a2d75c8b1b72b4f7f7409a12bc91a7222b371aec502403faf3f1ce3e54f1b0f21c6c47
z6e6a3cd51ccf92fccf4de638197dd758373af20e93efe495130b69e3718164e1d8caed8c8569a0
z0ef880095bf450d8c91b9d2e353ffbac80ffc6371f89a1bdf0743b29c26097e9e3c3c5b6c3ccc3
z5570c9ebceb48f8593e9070dd380e903b6d41cddfad7de5bc7644fa3c561b9813af6574f80e3a7
z5fed30bd9cca8fd6ce7c35e154804d85eafc6cda80074935ff2c8309293955ec0092c89da1fc05
zac0b0954a9ec58e60a21d641a87a249803f2c29cbd65e918086d64e6cbc02d75d89415c3b9a911
z6e0cb7f414cd92c91971b400a193958bfad0c4a827c123608bf69c40834ac4c489c7f17baa42a0
z79079ef83ae972e4823fde3594aeba56e32e4e78473fb0d99a88236987bb78eafb92334d18a44d
z8284be1a04d123186010bac36da9f9732a7308691a40d2aae4ebaddcda0023197d2febd376325e
zccfdac4a81309322ff519a268a4c3814647a59929c905cf4352465be5ac2463c15cd3630b5ef46
zefcd1a8184cca671cf05615c7f29f3403570fb36ac0ff2cbade676d46f90fcf821f0c36dfb00c6
zf2852008fbacc863807dc1aa3f33291ffde365717d33686befad303b4fef51b10af399cb8f6267
zf564acb5b09671b8be8cc5af7d1e7848eb4f905eac9cb29d528fc157cc3c3cfdc6baace2941704
z95dc8977d2d26ec08366560eb8d730779b52a050056b253d41a23df3b63dd574b37a77ebd3c596
ze6e973a62f9832891081e752a6c9f93e2f5ad03ac4f0de0b6f94fd3ae5b21bf91e84d401825ddc
zeebc7e3e296e13b46e243ea256ff6ea50c9851f17c5b3793e4eccae35873d0994010921ca35886
z243a5dac09fa07a8e0a41181c4bc40fe7e6d3520a4f4db9a637d3c2b09d5657aa4ca3466d2f952
z7b4450cac1180a63ba2404dd57b0ef1c3c71a4c5a1e4ea4b0be4c1bf8ac4c230d60c75f53a3c1d
zd305b5b390423983da535834c98ca555c6ea3d99cd033c04ea193817956b3bbb55fb0c7e63538c
z4e442666eaa5712da64048a66cad31cd512c0d97aec09c6bbb3bfc329b3f84c76a5679ebe93294
z6cdb3a060ab7ec0b529827d7669b60d1b76b414b042c0aa5c08a188a799ee80c5e8b87d5489292
z02d7f62f5877dd57dcd33f3a2ad70238dda3b0a22a31b994f1aeb83322ddbc3a9e9ab8f371e95c
z03b240d2130691a56b89e191e1a4d26a826ff34e2832040cb571fa8336e7149d6e218deec83102
z721b914274bbeb2c5b7d35b589980ad26d7a540b1bc76431a306f1a061dd5eab4f973fa1e24a8c
z0142d5e709d0daf6ad95af25a8b922327955c5cea57c02c53be3faca2bb2cd6447b0d959736501
ze085843d89f02a8451bbd0716862e3393a3b046b9796f10b9bcc41789e668d49514a18cf9b8a8a
z970bed1cb860e4aa0eda8593505ae538ec996bc63dba9c32f2d48ab4a5f5ee112d090818ccafa4
z75f4a9fa5527a55d33c4f7e8bb8f2434a26c7774dcde0abef5122b0915af680076b0d319fd31a5
zfeea8826d5305e26c6e442909eb8b3789b4b4b34cd60bcb226251883380a8b0a3316a3f70450ce
z37526efc1b7777ab036f7298c1e460ab77e93dd578f20d27244c1567425f17196aa1b139570f65
zd1b847ada00a1a3f09854e2c84ae35b0189a143b9917b86183bbcd840af5f57cdd87ef6d7556fa
z5001eb8c9f3febe786408a003b6aa2b1cf3dc936fd22f6894f0a6328de0889d7cf42bb1ce3b790
z070be938c4b785e38ff853459fdd9f91b648d2771c3dc2a48fbdbbb7eca170fb3e4e0852d5054e
zedd7e2aed555b70c75f5f1703736d91931ac1205ecc49aa80241113f35929aa9e6148aeb2d396d
zc2fbe5eaaaeeb04e72c3e0f79d2a06780041dfe243d81fbdba193d4743159bf8bd60a545e6aecd
z3636e2581e846f122f4cc27a2ba423dfc54ff8fb3c79be347b3446f8cff959f84f7b3d578f5d39
zeb1eff89be255cc61867f1906c2d82acaada8321e5bd58d0331c5326aa7f97674074276e03dab3
z61c16cf1ea2ce36596277dec2613b65ab5a735fb0e2d8f7079dc11f940381299de4ae347790991
zd1492b9b8a8ef5998711073d709a1cbdb2b29bea85001f9f0131e6f10bd17a0c74176718a6df21
zed9db984ed1229ef1b97b09fcc00b2597411f4ef4759fafb9fc87622727835085cc6a7455ea94a
za5717cbf137ec5cda29e21d0de2b57972cc14306093a5856b54558ab564e95f6be55af26cb1a3d
zdb901cdcd082df1862aca4acb0868259252cb75b34ed5db4975a4f8ad654fa3976dcc9789c77fa
z103874f253515e9c76ad489784ef8c10e3638c604e76a5b2aa936ccad473065f59c11cb22dad4c
ze7e7b46ced87c7f4c69b981fa35625b161175a6dcb0864ccadcee0ec8d86c303aae2f8bfa0c726
z5f562734eeb39856490c601cd22d230713f4e4ca350f8128c9f8131c7afc87afa33cad04c0eff0
zb203d58c3b417574291ea3bf6283221369b0fa7272f0742d2be8faca270e4d2cacf2f21820d0f9
za5b198242b6be38bd535aed4117cae271f368674431faaa2b41f07903d2201564fa6b91305298c
z0c7bd94a19d14b23233add8fe9d8b56bdb89efba34cc92b70e050fce17705046fdff30f43ee8fb
z0c0e1f4ea8e72d432960af9f02f2396ea288ea651bbbe366c5cbf03dee7757d81d2dabf76fdd43
zcce96cd9f9aa8f349eb67df24107817cca7f91b3f207161303332c769d515660469685c2d917d2
z63d41978ede6408149449b0354cf996a0eb5bb8a690cd5c74f766f20482c2a00313f77e790a393
z3eca74a8785491a56af8317925ba03a2b9ef5c7def5994b99a29c5aadc113fa2eec3fed39a6bbc
ze225d8f5a2e8c66f2b015500b2a7418366e8e6efd0b347673953303598380143bab6f2103cc174
z20b85544aa53527543374ac70e06ea058a94b9dd66897e9adda89d1ce72f5ed69bc1bd4cddc2f8
z44ab8583809a9bc6d7e4920235cccacab88c610e96a64ea255ab4bf7e09352029956a8dff78f90
z8d63b27bf5fbe51e73f9d6e26aa81ad7a5d9453c438c55b68b060c5c9a0fb45b7707a169863886
z81589c3439f3d5e1ed9c5a444a83231e9f57c0e285ccd3a959748509d7877def182eb5c0a76f57
z517e55b98db720949e6fd18ff34cd8e876a4f3e141b37874826709177447435d3b36f6d19aaedf
zf526e49f9d68fa6bb746492cb69b8c9e9160c6f2f52cb322fedd301ac12ba94658967b90791948
z3f9fc2cc3d7f762c7966096d4377fceea911ba0eada1eb33818e3dda9713f50f037ad1ea260d0b
z8120c7fdc5ab5f2f52e668091e31a149a11a049121ee5c4dbc954a11863e5678473545856f3424
z0716d44e717f0bcdfdb79dc3183baa57cdc84b79b43b94f21325a7a2f5e422d99b08462fab741d
z92c0b69ec3fe57e901519b8f30e365444211cbac01bf5c7a6a989877f954949716582f2f62b3da
zb28913e52ba814745c6d96c6255f93b1f1e9d182dc5da4728009e202db862dd1a8c6d1a1847c53
zc97d55c556dc39531e1de86324771a1559a55f79ef2743ce495b14643c02764afe46017538a77c
z61915361b1908e23af85a2f62a985b3817aed1c05a1fd437f9370a904e57734527b31252097b69
z19a822b2bd3ccf24a88a0707d486643cbed6189f5bd668a580eadb8c75756e2673c38139b50e53
z731b9a4d8a8da587c675dabc2f1c8678e6cc48841f43f3ba0660eb30eca73c370e5edf6378c691
z84bbdc8be40f02e0f3806630a082259a1120fcbd2ff2f10c022d9da28e6afc878b442c5500f232
zd57b5f22386abcdc951925a25d94945534adb886fbaa93449a25d4e604b09cfbd99bd433a91502
z33ac53ffe03cc716c771342e687ae9a7e4e99f43ae43a142ac7b2c76f9d392dc6d00109baee9a8
z511ca55de42347c9b23dcbffdbc9aaecc7d6ed722c1c76b8a5aaaa55c60f67d280c4b652f80003
zbff732dd5d28f55db3527bb6f7f8d42943c153969a1a2fe76c1c82040833476313807d5d5511eb
z6653cce7fed946390eb53c51caa9e4746769cd3b340f9abaa12d318b30f8e22d2b8c2dd8a50383
z9bb12215dfe2316c17c9127c131bbd135cb16e3e64c1270f016d28ae4148c400d558c22625428f
zc0bb8e12b13559eed8ead854a28a0bcf5305209b4f05b2fb31151a38c97333316ee51912b759b4
z78146e9fd0c305109ee47e660d6af97c08b016f4670a7d882cb999ee7f448dcf964a269d8e746d
z62fcd6010550276b8ae114dff3c27aa4cec3a57415f0614ed2a1f50aa60a9a80368c35bec19db5
z71be07d59022e39b1fcd822f2e9620f3a2b797f72dfa2b370792be3e4f6caaf7c1c86dc38a4471
z470bac0b43677e4167e183d1be0ea16719b9fccd2889ecaebe4edbfee7197d607f1619bf919210
z2f261f9d23740b5e2958b4f6a2c34e0c1257da032889af91bb76fb9f46da17271595c551bc7aaf
z876381bdea0e0fbeade7056d1b91ae1632992b11b8bff30806a3cfcb3dc44208407832b19fdc7c
z29eaaef2ce9bbd47310ec0f16d9ba32f580ac357abe3383f4514bf1e9b6c26ea73ce07f75ce5f9
zd7774bc4764a532289a033501c6c0bf35e8453eb62114ee72537a6966c7fd7a9b90e9fc18e348e
zd5bf6d88d505b5209da3d4e2f267ebb5879eaa89505a9673a65a7266b2861d1f444e6777d07367
z9c46dd5907b89ea05a55317cd46c566446b9d0c374cd997baf179c2f1a1498c995f9296a003344
zc25023f155e829108a7ba2a121950818b4403ac2894d0a46a977f06f6ff07a4bb94f2a8e68b530
z511bcaf1bc6ab268a97871452ad4267d7ca18e4696c7457a249846285c809a7ca06080c26fbc40
z72e500f049cef325b1a18100856a0cab7e730ab0292c683cbe4640d1247cdd1add353c08dd2c27
z9313aefc79268435fffe2249547fe6fb9acd58e2edd93a2f343983aa94f013f3490f2ea2342378
z0717ab70b4773b168bec394c169437813cb4fe8b088245ce71c49b05c066e0be07b7185aa48dfd
z27b080f710a6dde8a17ea5efafce95d67b252418992c50cac8e64b254035e90f9d29c436e670c7
z2e25654c589892a2a64e0e9f43ecdfc52897e4942ac910446fb0862059d676b53da069f6711edf
z429d14000eafe4be854d75bc6b18179f18604b11fba958b378bca2f88de9962074fd8fc5a801d1
ze21821ae3bc3ed1e16d88ec50b320ea710e7b44c945b7e15702dbb9f6f2a11c289b92d48803ede
zafdb678910fa20cecd6f627e393bba7fce2e7ce179146cfadf6e1652ab376c830c44e507d26cd2
z49a87e4db6073c35a2b799a54ec0c31f4da3531fdc0c891f9961822568e1a4908768fbf83ce170
zb6e0138c47519baaabd8e32a10f8ca1df0ae78993f518d99f31a86b7f3bbc7fd6c58a3600d1a05
z9de810203343b975aa64fcad41d3f91bdde5dd785b6cf68c6b1887408dec0ce1502146e5354364
z33f8ba23e9c534556ab3529d180e5b3bb8f2a80d47d21af5788d6d211ae8b0e7f58f6a674d38d3
z37d25fb8bf7b8922e4a77576c53bc9698a3b55903f0d00246a29b2f6c1b7e59904cf69f99c0077
z3e07347b56d92ede560f68cbe5d333b52b50a3e0d3eecdf41fb5751f65305664e43a3c47bcea3e
z3af5bed11b810b1f7fc308064276e3bf6ac167fbbeb2ad29f3f48b810a0a8d3271ec3d1ed0af4f
zec54ca14082621488619c7a49651e60be5c7b37b10545b0bf7db2db3cde7bc8a97bf00d989e343
z278b93af0cf9f3377a9e722c414fbdd1a7e8b5c933ee79864cf5a66fbdd377c3f816768890d2f3
z76b9cc61a03404d29038329c7a04b2983fe1664813fc67696f5f44e79ddfd1333138db091dc44e
zaf543e79f378b58b879c073fae17edd99a1b1da96aa16ab2c28fe3912f85fcd90afa7d7303a58c
z45c2ae413b78dfe5fc0a2bbc0615a68d8e6f65862d10e42c4780016abe6874c9fdedc71fcfa189
z119f577259013a2703e6832197463822611ae987699ba7cb4acb149396630a521a60f996cb330d
zaa1279bffb844adb5a59ac1792068d3bb561a7a5fd046157061f8cd1a6781b9c683675f4763211
zf4d81568dd72a4f6953cb8ef03c9f060732142fc450bf0841572ba86298f3dd8064e272fe684b2
z5637cb60aef05d88113507a219434319300b12f5f6aa1884aff8cfec908cf255e19b9d0e203f50
zcb26e61a47fce3dda46bfdb7c3ab8b248a3d2d834fcc88e1e4a1aedfa6b62ebcfadfd8f46f47e4
ze8c08ef107f8d8884abf705b391b547d95582b42f1f1b4b91d70f95374b53cbb9cf58c5f03e3fd
z8af2d02b5422e848d779a8848434be32ebf1e8f790434e380d163df66dc4f6bf14070a7fb7515f
z8d66c6fbea8f73b84a1d90c038c60055ce834ad81a1b09c4e6b38c413111ea6e7dfcff1e71e441
z9ce9d7c5ab1ccd412d238043cb55e185eecb16e5c56b794e2adff2852fa80386108a5be55bd3ca
z61043af8ec2b05ce3ab19606445b35564d7a4fce508f5f23b5ffc04acc7f3ebc2b19df95546f3f
z5147a2fe4e15034f9285ff7c03fa2ce6b7c7e351ea4b6a09e99dbc15924c6fbf1f10ffc0622484
z5fecb5f7da87c0a59570ba8bfaa706d4e39db0ea9a8394fcf0e63922e1c32efdd7b6b9a616b853
z96d5ab68ca79da0d0d9d4afc525bbf7c66e611c055b9fe3e03bd741594c6b28d32f16a4cb3e718
zaa324a146387c470ab096bac4b40722e9dd531fc37cdab3623a9ce687c584ed5c0a9600cdb22b2
ze26f063fc4b55bacd4ad5a86281774ad52f4d6a4c092c5fee69b5af21a3f003ae48dde88993b79
z39162529cf01a37b4581dc47158ccdf4f18a1841a8192e2de7f1405d9bce4e80f668f99decee5c
ze4ba366b6830bb7ce020920b92d2fcb217c8a56509373129c1dddaae3d8b8327b7d246202eadcb
zffc183c75a9f13bee4d0570046f33488e3b8e17c1d78e7307938c1a3a2c0335169818743806544
z224658f6de9ca1e231a78630d82b934957618dc20db86664e9a69adc86edd8ff9f02e9ebab5b4c
zfbd3aa17546c686baa5fd37f5c05e12be525b1530c44f65d736a9395f1922a25443e495f4bcb3e
z606ab3730c1fc332bd3d0ba69cb05214cd2eba0f9354af444607ce9c678694d7e104272bf30c37
ze4a61de4e3f906f550eac3acb391cc38aec80ccc0933cbe2e0b5490fd189fdd7ecf6fbb61244bb
z1b73063cd8ee5383f75eab419cf3150e9bcf1fdecf36bc49a5fc590a7d6d42db004a67370609e0
z150854f6d3f9fa66f10b5c7094a45861ddf389aef9a2305cc314ae08eaa36c539f3011cf26f490
z149a5adf7099c3fc903cc027353fbc2d4b31b85b5a4540fb547758037fc5801fd3f97e93427d67
z47022158084d568aab026549e1aea932b3d2be889ebf999edb9a14b3d8f2a5df0b42648d45944c
z5e84085326ced0a7529a63e19bd2f8a8349e16128690542db1442a213faf4cf5e0b99d43f7377c
zd90cc5b939c872be4311daaf8b7621a243efdde15644b03b60879cdb9c829f8caf102e84079d98
zb08af4b10b64e7fb9deb5ab91bbc6f5b7b30eb5d2c5789a2a970e656f2376f3eb52bce401f9c67
zac9b99e11c324d8ed079ed066978db914b132c5e6e268cd4f205fa8c8c45b30bf931c62abf31e6
z71f341ebd33ef9166f770346ce0b78058fe8fc94ff5bbfff5029874f0035036d1085be8ed80529
zb1b8e8dbdbe411a6777f7d3f9ab8f388f24940ce4cdc80ac6e6f9b05cf8b268d8beab93e20a8c9
zcf160d6ae314f9de877a9844146a4971a53509694217d0d84e29417d34203ebefa9b2a691b5ccc
ze60b4c697ea42eb7bb27ced0e609ddb563096a15a942be0a9297d98f564ab01fe3b005effc02d6
zc56ae2743cb310604c945eaa6dc1ca04c135cbb9f25ce6f38ad51dc16b4698dcf84ada1259131d
zb449453e7a4ef660270293a2768516a394dfcf1e05dba9a5063044d5fd46eb163fdd4f86bfdd70
zf67af929e1e2fd2fa1124fae2bb100f96f461ea10b9236526a1437f0cf1c55651ecd72be6d92f1
z99efa56dd7536826b2c0aecfb59011bf70e95220de7ec11a448577e6d01c6050ed87e1f21fa75c
z8960898fb61d0e59f1ca81d49f1bbbd5f8a6a9906f1ea9c542ee4b85fd2300f3c9f68e4c077624
zad1e796da44131c250732174c50bc8f9ef872eac97d7a5cfbb8da8970e08429f44c1ef810086ba
zb13a136b3e38771005bea137713407b3044ccca16d98bedbdaefab388e49ea05ab17b1772172ad
zd7a255550d2a2cb6c1767cbcf4e67f4bad55f8c43fed7bf626108f4e0cad93173fcfa3279b2ffe
z86f12e2b953074ca6311761d89e6b9aa074c458a5baa9f77f6fb549b8c0fd593fac54d7e3e1051
z2fbddbdc798be21168c0319e36450b3b34e944c35a8fa6e95ced9b791677c5de22e10a7452eb85
z61d17ad0adcd84c6aa042eb837c2858028bcb6189fd76af86054ae0a539497e9943d501e81c7cf
z236426e2d209c8be71e321f9e40a785fc17e90c7e8852498f522a1ba7bda20d4a71c4b14c0dbaf
ze7a723229fd9e4d6c1d73c145c15a76f498a2c5a711ea774c6884e91ef67e6022fd58603f0b384
zc28c3603bb5b1ebc23c46bebbdad605186f17177452460dd1b7787fdcef0124c3d878d401c1d8b
z1fee0d759841cb35e3f20040b79dec6a81fde1f6c6e7b3d80b5dd96f021fa787770816f2490cd2
zf432d913158231bda4cb9730f29e0f9f7a4ccca7664d3b69b9981e5ca8d60c7ca8e02276b03641
z504fe959a03c1f9bd75331c81a8e8e3ee42d701cde517ef14439f299f611df340865edc84d1615
z1e15a1448da4fd44586c2529073cf91269a5138e4287d5595935dbd3ee95ee0ee7ac4e6293d7d7
zcb1e4d65f910f1b4df075f5ba2a9844bd5aeb818f253350df01f63ac0685cf83417563307a6a0f
z0f73510b328914bc4016a9a82d9541e25173c7e602ad4d8ddb3328b02321d0d7411fd161bf511b
z130f946f1447b3b2c48126f64f1c36369261f6079555c7721d9a2c2a912dbbb693536e1118efbb
z9619990baa713647c27066bbc6dc42f8ed2e6d1d82d2a5e7225bec95fc6e2db8c0ec3320897b04
z42badaa4448ce8cc9a804927c3c935ebba3198fdf85fa4f92078979dab2df997aab72408cb92b4
z1f52b6863934fd284bd165923520ae1ec0873d5d506ce854011b0dc102a2f4b7c7b748e31777d8
zb1abc48288631df5d6a53484df2086ea98591d92230dd2e2c594109bb92c0dc2fc480a39819d73
zf34ba1b8ee91a664f4868b8b985bbc1b20d6e49807e20dd7f9cd7e47ade3aec58ba1139c1b1767
z3692e827755f9dca3012d67abaa8b58bd4b6d91dad36ae4de42c3b1c2e0b06fee5dc9277d20ae6
zda4de95e67bb3f903628b36a70b1a0db46672f56169c05b9ac79639c9ca78dd9098547610a47df
z0787c40b42046953c1948b2b9825b4893edcc8847342af8b5304d086a2e5db02adcf404ccc2031
zba5078f1fd44b81bd3852f38d035d81f81d0856fd6e80508a375addf2409c5f154f406b263e86e
z2181132ef4161d7c5e76ac94970ad06cd214653f365cdfc26d9dfb5298331d35930042a49289a9
z805bb9c7f4f71f733433d842ad8022d6aab123e233c3a0fbf55a876aff754b41bea5c474519b8e
z45f83ada62a65c3e93eea7f579fdfcd5fa6be016e3b32240cce752b8d563d41d41fa2920011397
z3dfa023dfd3e3fb25e579b4d9e70bbeb11a68479faadbd6ff296223bd1ee096c713612226eee2c
z7be68dbd82dab3169898332c33c909ae0ed33a9aea4ac5c4a854f6ab5611ec660d6657d9e08a0d
z4502c2bcbd4c10ef9a7e737035a7676f60f7ebbb92e4f1a2deeb71c1ada4b3bd4eadd05966f418
zbb77b4df990777edcc95a936f926bd35f1416bde288b9dfd3cf75c1bd99ccef3cb0f75a9ae0753
z9df43716d2cf1f3a22b17e6c7bccb1583a65b26a0d8c1b01288b485b6fc93c6f23cb4a4d04de49
z8f3cf0ebd7cbbb9c0b55a3abf4ccf6b1ac8ac3b9a261ad53e089838fcda4e212bc68eee00aff42
z23e563cef1c1ed25be89ab5de7ed4265410254491d60acd908e6e370784ada07b7d735cfcc8b42
z972947976fb895a0aae70617a7ff151f27bf040d9f514987c6b92061218e36cec3574e0ab8034f
z335e5a4a084ca15dd0f1e1b2e3d95efc0b736751227628ca63798564bb4107e896f717ecfed5dc
zf205000aeef66e82612ab74d91331f5f14adc0f915705cc723b276d180e83e694d03587f2d6ea5
z53e52661ade7dce51c8ca9333bda919273e09748580f50faff64c406736a28d74aef0998ffb0a2
zddb3d5f492fc8935950bc8f48b2af20f9cdcb01ce9cc0cba7fa8bd9f3c5fbcc20e74db3b044ea3
z0018191d5ad20be26c74a6f6cffab7f7ae70de4b32c3da7ad7b67f6f265b6ccd70b63cb256a16e
zbfd6f1ea1dbcadefe4f54d27117bb892abef7ec0b2000edbceff024fe5ca82f43beb93e68996a9
z1f0cc159feb07e48a4c6f7db3e81d0cfd1a1d75837a4097503e782fde6d7b5ca58a673a10f7717
z598fa3926330550a000fedf00eab72ac3d3c695b8df0cda8957856835def41cb99a6c493651a79
zf3d97abaa873dece6ef49eef91327c96eea3d4af8df073d291bcc49b4092eba2b858fce8b9b913
z6cd54cc05226857dbc9894658d4009baa6f39e47856da6a93904c36cd7475604ccf5ebdfccf082
z509226e2aab0ef3052f2d7f63355f905960704c71d099eef6520c6ed5b5c4e95a316c4e22ef215
za8df48854fd306f6b880a5292c26086880284db78381f41aadfe94c8bdb10cbf91dc5098f99d19
z4eefa2b065d960e7467136be795cd838706a1ae4e868ae5f0ba365df842d620746d7c9a97d4c4b
zc6b66c843257258c8659eae043ad0ff5d710b9408a76e24177ddce067182cf99877a10aaa8e081
z3ee87e75cf0330b68fd3f5aa60fb1c34aa51615a4b17c86afd304074ae8c133888385b84fbd7d5
z796844e3e7b6b43d0cf894e397903622b69353196dcbfcfd13e7a2db5e6a91e91e5c4d10995eca
za9ef2f42009455469383f6fa8855faa9dca6611f4b88c232ec61d3a7760c6a347bf2c5e8eb9856
zbfe1df5fdbf19b0aa8bd7fd0f2d6bfbd727bd984eabd08d4b57896143f8604df4c6c7bef2de852
z6cea8638a54a8ca0a9889f234561b23bcb0ab8259dd970d63ece0374d62cb5f25b754ce764eb19
z2296d833c5537248ac6a0c9fd4a13e171d434fda99dc196a78837b5d10aeaf8bf28c10c877484d
za6f3c8a2be4a0157dd0ced403a920063ad796a46eb23f22147ff784e2565637c2c456e17a0863f
z06568b1e548ab6715ffa2f3fd9a3085c3cf78999e92c0d68a3ad942ef0b1049fa4adc29e2df50f
z09907c169293ed512ed8c005930bb8dc3c19fe1612132e80ea175fa4fdad7fe0a0880f83953b0d
z6a16f4d1baff16402972ce0236fe7dfd25430796c3535fa639b4a4fb0614a4d9e9a0c4ac2a7bdd
ze2f8f8afa2c5197ca75502a913f71d2e99ae96dff78b221c631c174e106ec73593b8cf07b66af6
z5612edacd432ca52286f55fae19190bc65f2ba80f3b3bc6d00ff042adcc13b2fda888e2c3ff0cd
za87533e376d15b7cda401187339d69dbe603f6a1c573f0b04df9f3915bc2616e8c9234c7519931
z42e343ff17047968fe21dd0c234c7d7ce4ea6d71d0a6fe6e9d01450b5591522eb80523c9333297
zb591503109f043a4268a25a5e7968450699831ca20ecd5aa4a904659de86c9cff3303c99af2f05
zb3993e25532f6857b112e33f0848e1a57627e0e6273e0cb08d1a468e306eb841f9d8e78c7babee
z120573912bdd718c712165af0acc5cd764c091bda79bda6c13119c33f00a0408cb2706a9450681
z9cbcd393010a9e4f8b86e739964e8d613db47ddbba8bc2fab1b3885dd026a5de1d351371f48637
z9f8b5bdca8a17b3e1d879619931be476dd9391958a8206ebb96109cbb543bb7df753d73fb183ec
z81602f1698af67746b1067acc6d8729ad1550532282a9b2fc3c7c23ea61b93e8115a34d07c65dc
zb3e7586e55cbe44d69273f9ee4305a73cda939ea9d63010738ef4919d27ba756377437cc3fd74b
z8d6af3a8b541fa0e1e8c9a84daddca5249e115d88e82634a1dce49d9ab072a37a2be96a76e76e0
z5cab476ebb33aed63cf8d4781ad588842cd8f34696bbc2d7a333945ce3ba7f75a2a4b10c072a4a
z0386dc71bf93975b89ff3370cf5ae703db960d8a2a9168e1692ec69eb3a0b611457cdbfeb5262e
z7a8e025125739083841edc53e6e43d5e956db1c43167d5dc78194014424b0396786f964741070b
za0db2327687ff6584ba3dad1a8bddc69a93dee7884a8034209c22ba18109694aeaf29efcadfedd
z808995c8c7a2346f90ba39ff077d6f19adf686f4d3ef63c32cb850fe7b73dc45788bb39b48d942
z49f4ac21d68d148f42216a84022d5c8c80e03f023208ba6a18864f84fb9defb1e4e744e9525bce
z17fe8f3b67bf097b8b932e420a6b23a9838b46f564ab838e451977cd0075461926870594e41e54
zbf334e5b6e4526dafd8e1c426ce4ac80803382202b68b73d7755d1ec62bdc7b8ead48c7a8d6802
z379de339f5cadfb2d5eae0755fa844abc8152b4c5d292967a4362eeab3cffb3ea06ac01c1c5b02
z445fbf65a96c32b0101bb2f6f56e6d67c9d9116d5e87694f047636a78fc12cbd1ec4e6d8940dee
z3b562562bbcab7fa2b43b6a1e62e1b159856338cd6077d686f2f8fd84e815cb0d6e75060ee6576
z396c71a671ef76d7838166209acbf29e57f4948de365a755143c3c3e0f6c023275eff3e41509b8
z020dfdbc729e8cba6430e5089774a039bcbac695062c540e03d67dce0381bd3e17c5101df6dc43
zf3c52b13421b939a08dd32dca413026f861b481bb1144eb242fbdb38513131618c19b21563d426
z070155268e5c275827bb32017b7087bf1c6f21d674e8b9e8ee8c854afb2b64eb16f7f8b1c208df
za4b2f3449c089691b66a3ed57a25b4532538857cccd4fe3287a782251cb5b032165911ea57a7da
z4a8214cf44ac28f7e301a6f0bf413f1514c6aef6b7327301044de9c491a5d1c18b9454e449da67
zb83481ddda6f05cd275b69e42dfe78b18c315bb324ae1a15a3a4f29e98bf49c946102bfffdc0d3
z4e8de10bc58790196c632115b2031a7d5c3bd567acbcb11db28fada650ebe57a6c118f27392d9b
z1b7c0551305528d6b0bd2a76e6f36b0cf8f288bad329299f606a8e542fa7fb8574dadf9198297e
zb785cc320e127c9c651b93f202c64d419057cf9c70d8ca99544d71696cfe50aee4bed98769d1fa
z01ba1f42d40d128ada4405cd346d46a01a2a04588be38411db3a7dd54cecbda463747436ff18f6
ze056d4bfc439669bf789afd8cf90aa90ddf78b5329d0f9126db96862c1ec708afaf066de4aee4b
zb12c7de3bfc975f91e9f1542a8e8c71ee59d36bf5ab84316e3e359d57473e2a492f214a46e4a6e
z1b9d1f4e872bc6bddd502180d189e2680a989a342bc0517f64a0730eba97
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_encoder_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
