`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1bf3f153bd631387c118a296ca10cbf0349426
zcf2ea5eb241fa84c8ecbbf7180f10eb9ddd4966d421e6ca571b198ed195474578ea51160ffbd6b
z0f73216703aef2bba31d04f6d0877540c760cd2535de4136d5bd477110774792da6835e634764c
z9dd137305fe30c578d9f560107e20f590b4eb309f308917359e9c0915665f92ca16e374ffd3213
z5882ccf3f5b11090d90e8eeec978eb04933b9cde5825bc780072c8a583515260f27d62aa9d03b3
z6f3e04c10e3836fb118cdd46aea7f3299c1d41c7b27b477f1090e204c6cd392900036e6a8eb175
z65cb01f9518c42e024938e18f85200596d0363d006eb9c81cdb647320cc07b54a7bccd5ce1d4f7
zda7559946b8ce85838d9001dfbb2d7a30989720d68c9529bd963202f9c10ef5404bfe96c71c37c
zb07f8dc7c87ca12b1ae75d6cf5f3b1525bb3c128eb5652ca59a9c62fb3978782d5955795adef03
z0f8dc29f07f11fe7b992412b603a751495d07c284658c31df21e34cf67abcf2783edf0a4d91253
z23d6950e82c2f87931bdf908d532d4ec53efca335f59c40b7475fac935e7cfb248edbd1b2a62c0
z21ed85b838ba1cf8979fb72da43e762384b95126a6e2945f5b191c9139a459e1bb0a291b5efc5f
zc0753284f869f70e22de227fbe3d858193f5c81f39d94d02c87b94871c7def62dcf5c5d98202d1
z3340712fb72f0439ccfc0d05b1c9b675da1dd92642de4f9c57594edd79c8727fe05204d54dc065
z509a1bc1c362e7fe15aaa4a681f3b32888cbc019881ec8268fc9fc9edde13f702ee84edaa2c567
z5ddfb7d328eba12159d923db1b5ae4761e9816fec0b6c95238ff79fbc9735e447fba09633da549
zf0db51f078987ab7dd9ef7cb4ce2673c1fa000e21263ad52799e2de9ccc0a8f4f8d2a04a16b217
zbcca4ff1005aafccbc0686e0a5d1ed743c20d096403d4b8d39a5d092b54406625e7a348578e772
z26d6a9d8f9dbcaf33d3e95549a1b6580064bacd4b7ab6d5662f21ce418518f91d4ed2099a10634
zf990fd8f163228fa1398bae94fc1d693dc5c6102be2a8bfd0d2de1e75db890cf6de52143340fb1
z6e94ba7539848a22d536d0d41d17905db53632b2391a2870ac9b9274c0cd0636f8c229908f4a13
z1fe693f35cc3143f115c4cf33c49219ab5d2d1cf34a21c30f9ff077e3384779e4f9dbaf6421cb9
z14a06a4ac07db33495e3a185f4a2cc4819eb38702eda8ca4cb8318a2cecf071cb01f0854b5ba7a
z8f3ec9bd7a0e6319d0b83694cdbb423c9087b8e050eaff2cb15cc3323dc1c4278db7c1a31abfe2
z63c56e3d182de2e4f5dfd65f17c2e1f6abb66316ad0745b75f2803bba2be8cebae7ccd9712b4fc
z4c0340d77dd4f808a42f19753b42d6155c40fed730694e81212171836258913706bfae44384a26
z5a50f68140500d9b66a45f02a78c78ca65222ec65d76401bf14089a729821dc50634811971bb70
za093eb1d8690c420148f8e618d43cb6857cc1745a5099abab1902e6855d1bd3f7643d108415f2b
z13ee9fc02bcfa79815f8f67d31dde0e5452a1a51037a9a62b2d1928c5000e21214ff678f073504
z7eabeae56a270e8896c135ea6363968da799ef23a6527627c7adfbceee7e4d6f667d8d4a5defe2
zf90f8de6f4d4fc5827a4d5228742f24a8731b2907957129a827479db13f906c85767ce3b8b04fc
z97ff689aeb184e84304bb25b1473ce9d4a4aae9845e289fccd633983f6628d8a7cc28d0bc73c3f
z38a18650ead70569b77be45617d075a36f6f7faad3d6f17037232aec2392c440e159198709baaf
ze165d558164e97753b205ed01b4ddf096c2faa4197f4f5b4687052f72a4f5b97e0d33acad2c610
zdfc4eab255e985b7e1e3d0798bdd30de16054f8c16db201d6ecb2087aac5cf00515f16fdaada04
z03c0ac9753d859f399229890e4f4935f216822f8b253ca24b921f9a9e72e6f6c46393ba8d5f9f1
z2e8f4e3d46bdce4c37b8a9e9d646c475edac8c97fc6dfc08c29ca0b20ac350e2ae7b58de9e2c71
z6314bd2e9489c51cc9193a0674ce6679a866d141152b1f69c2a3cb3bf55c15f2002156145a1690
zcaf4ac83ff7750955775a72390ad868efc2b73c3652c9020df8b56e920e1837b6f1d4d8f20e06e
z9734c55b9b540544a14ca1c5146f3f9da51936b58d20a80ea5d54658a174cd8ac4e31a324bcc4e
z57e43db4cd14cec0f36c129a3dad273b7a6b83a76abc4113fb36c9d1e4ba9583092fc10b18392f
z1486a4922fd5349577dc696416b998932ee6982635edfd3a4ba7998bf2d73c65fa33059dd5e98e
z3cd9206c5c0077fc736c639aea2a74efe4ce204555753a590339ea3f7ee6d406e17c5db371db51
ze6c554e24e494a9fc74b469eb6746b009cdc392f022b96463a4fd0a649901d84153eb0688f1153
zf242e4c5fcf62129e4d30c2651e8acc94f100bf0e543999ed5530b11839f9be54a3348f38bbf87
z6b685381d97869f347a5ce1e2714fa7aefe6f6b5603b3498a7a6bba6a237d8f11a21c13a16c28c
z21809e88240bee9362b78d5c601a809aa627f16c5afb35da85c44cd7292b91e7726fa25bcdd018
z20f72a776724347f6393b0d7f64e9a09bd58af8d35a9dbb2fd5882a40a1f7fc6b66133a3a77afc
ze09b674b6ff3456f7a59e518c9bae38c6ca1f7b3638dc10099fd427b9b38f9ee49feabab741ef5
z8e03e678607fcada86b2c5bf9fccb42acf1a56efec3fba7f251c8934cfa536f17757bf196fc1e0
zdaa952a844a5bb9822584de85364a26cfeef8dcaa19d98ec7a4e0edafc1f784b58c1ceeda5e5f7
zb5cb50048c64c3a298fced31eb1a6bde27211ff4a845b1d85ce359468d9909b299c4e7b4efbf69
zd897edd9cc41dc9fb97391748b371cd46cac3d0d56c57b9dfcbbce8cddcfe37d8b89c8224e62fd
z9976938f1bc1fa9d3124222722098eaf54d8d369003232e9f3afbd36b3d5188ffc0ebec9cfcabb
z090855a02a5b2cd279c79cecf4af0ee4947dc32996373bb572c46912b350641f70580be539e5ed
z578f27c97da8e961171315fa25a8f5f9112bf7eaa315dc0c22fab353d755835987f6e44d697754
z8dff4923f379d5ae9ec7b6c73deb0642ab46b0f8770d19fbf0c2127354a96643251e889854a4c4
z392340bb9266e5772acab586e288a5b104b1bcdcb4c93d8c715952e3ebcc94d9204e0a4852951d
z1608a8c3687ba2741b1ee8cff729902e438d3e0022856f921f9bc5013150be142fc8ac09f9349c
z260f7835deec7142b0f2154797636c000d6e1a0f8c982251bf985113faff26bc662c9688d395b5
z4456c62dc25897be9d6d890a54f389fe57792a0218fb757ba8356def59f5ec9592a77bca2bffd7
z9021fda8f61851b74fc70a53033846c229995175f5d5d22360bcf399785889cd2c3130f5edaf85
z09f87819279e248217b74b62a5e7781f2902a240837c3c48b96ac5a07dc3ffd482eeca40b17e28
zfe00f7302a71dceb3eca25f2ec48f510bb70b1eb94f2e4eb844d21b86209ee7670dcf8b9701399
z0d4e52c23d4b7917fbc8a465830c7a1c234aad5ded605db499dad6ffcabce43ca5f5c942e51f1d
zfe70fea440a6b912a9781cb83cba0d1d59e64ba49fc70c9b8553a22830ef53707152bfe22046c9
z1c407198105244074fc20d757ef064950e9d184857c865940087a0ed752d3537fc1d5a1e86c84b
z42c84854773cd742d855f04d1e90ff921185bd03533aca9258acc1fd6247d8d6a3ea258cb6e16d
zd9b339e480fb56f602a6f683319d62dd40f59b4711c4603f7d79cd0ba57e288f2aca1b55005760
z9cc6aef24477090034c6dbf18337795150324c9b8c0aaf2cd11a630e783ed6368da966a9043aaa
z431ea97e34b56d42d09365b08d98cea112c760d5e564d3076a0ed37f069a4ab3cfd82c073135a3
z518345696da5db0965373878b85a120049b9364550baa525d798ee6abbc8243023682960de1993
z3f5191726c2935a0dcd55ccde759d56284e25ac0171cd3bb9e1a235e82a35287289359cfa6f4c9
z94ed09257c05a400cda36012334594a27126bd473616a1c3621b97a81ba38d86317512c5ddd5ac
z3226c8a28103113589ded15d58eaefe0560660270d5b74ecd9dae8a30dbca8fff256f6a15444db
z7c1d1510f136d248b6788c172889d1f220050f1363a08c7823509213a333298edb6e11b07ed7d9
z569327c63b5b5cf2de0c6b7dc62ea778fcf176dad6ed666ce1a3bf0a248ec206af6728701a23a9
z46f8e212c2015dab93f320b0b5abfb10964b3bf717b4479f18560bd1a5d59d8cf5a334eeb8e11a
zad450403bf9cc4a51533cfdbd715615f471e050954442b10e474018b231967653aa13cd1b0c4b0
z060d041230039a05fbc176f76d9911d864b1517e33953bdeef2ba5d656d97cb487df32355147c4
z6641b4a5a595db1d01251220cdc400645641a040d0b1c0c51bc80d115a389f081fd67f67e49f2d
z265634c31c705f0ae4b9bd747e6e38a59fc8b48306d32a19d83c6de31c9b4b9ed48073cbbaf88e
zd45e08d8631e09195e26ac8f7889646721c01fd5eae0a73513bd5cc706995150df24242af95faa
zd342ff0565c312b9578f025ad38c1f9de51952f56f820a817ee259718fbe42554d65738c505a89
zc84b31c85818463beb76e60f3d7da0a5944e4457ec8862bc19483b73c32bcd3eb9cbdb88dfb336
z5db512de8f8c0a9778bd75476a38e53a20aa379db7c6ff82d19bed64ddab24df984c9a472705d8
zb6eb8537f50109d536d13fb3f056293b38d0c638836f6247978149cec6cb759c28f6b6c1e16939
z02789b080a963ef15b843664b73ce7ca520e8f25faa64f8df6c44990f0ebeab130c912ab6762a4
z28a5296a51590b1f5449b7bba784a7ee1cd6a1a86a365a26212f2354142f0258b191777d24ce82
z0f98edb4191c127a23f7feefb4baabd96022da915467ea17d13e7ab1dc9b7da66b2da7e534ff5e
zba6a8af5773b22d4bd485643d271b71e8ef847f2f946a0fc73f890f886e93848270a521bb6274b
zea82f2c82387e81baa08909085386893db35d26af4d0fc968aca4b2974549ab953acc5e8c605a0
zc89e7c400b84e8b830d6bb7150ca220709669b15882c57e5098a431b34ddf8ae3480f7126dc393
zc7fe2b14f21da10c3ca481e1ac56d660c88b168bf8677ddcd05971217062283b712236af0b9415
zcd3f78fa197c0d3bf9a2e3d5b00f9572daecdc0f3a025ddda3c733fecc50024c3feede8aa0b760
z0cd977850e178caa6cecb614c1b83b9309f6dcd66b0a807a0c2a8a0b9d50e8e8e8d6cdc6c16aeb
zf438925b8aea28aa841d9b4ab7e2075490a325dc28bf911727d72a56856a2f0eef0f77ba65b646
z92756720151ff3fd725fe91599aa48169ac5fffad5d796889801d71ad489c907912dbe42019709
z207797aa498541d72adb6e3dfdd51ddca767f7b5528e5cf55997c87454e86db19aff257fa43511
zfc879318d54984a0ec6c9099a2d8e4c6ffae12da3dff89df9504e26ff1cfee8f2e75c2afafc0f6
z9af58e0dabe1b5164b7c2e416a17b2be8e8e4514a8d1fccb69dc262ba2f18a4222a351550e859b
z1a941a3ce1a7f63bc4bcab843ce51410ceab25ad4756a55b49eb6ec8bf3710838053f79ddd842c
z77dc17349f0d551434033f5d22e59a5cdf56970776a1b52bf1084786782cf9e1360371f1998971
z21fc943d4e312e42e84cae3473c89ed847c48a05875db0cd92d259ad7ff3a7c87bcc5d9c88d747
z16ba2626a80871c3b662f898de4b894e5ea4021ff37b4bb7357bde38e0ba7300f6e2df42f8dfe7
z9d5f123af9d8193fbd1fdce8ef8d4ee26ceb518b82560b9b6a428024199c8cdcdf0af9dea14e40
z0dec15a06446fa2316c34c5250ba3f79ffbe8339e87f6f908ee804570f2c8a7e56af33a94cbfef
z252ec7c81778edc222688282fc471ab4b59ba0665ff91f887794ef9eeb8a4aaf95caa0690f0735
ze3766cbb18336f6216c21ad052bbba79f35d2c56d17b568d25769ace5ebf049179be52ce150e38
zd74fea998cb3a5510b0ca7d7ce0667a16b78ed570b752b88ee5d0f892a6f1e8cbd0df7366aef62
za7673beced533075eed23291dc510a7cf803c0eb35bb852b30ca49cf4e289621ec31ad71fd5b35
z9e89171a6799af4986c61711ac84536a35966491e610a2a79ef08edde0c30679b44ecb5f952675
z0f67abedc8c8845dbe19b56ece954af9ffab8370645d7112bd5bf307f525abdc59ca110a4ac539
z85b96f0a244e781548fcc5eaedbcd2fde05984cb5f6718148f4d6a013ad102b12b6660e0d832d3
zd12ab9cd78d34711595f49b9da1eba23d9817f5db1d6de19f270b15e0c757c167e020be1261929
z03b2f38c745470f3a6b178aaaa6348d18833fd211db19c96ad32e302e6f1a7553ff50e8266af8e
zfa3ee54eb9baea45f4d155d26a5de96e100db5390abe914236397e3759aadfc4c1e87ae66e6791
zccbc9a95171634d4dab6cd64714081543d6b3ae7820522a60b13c1e8192f9ca4a6ec4f721b64a7
zd40102da2d2862b1a00086665d4a2b0940f95e11d03c6a515bb8bb268520f4d1d7cce9b29f589a
z25f258a96754c84105a430c1d0b1e7f0a7fb28ba647a40fb1be93398a173b8c353aefd349c9972
zcb849d1ce442bf112594149a62ad7909d50877b104d7da56ef80d43782565653815328f39306a9
z7400ccb68889c9bbf382a1af04a7aade1658e7e73b3ee7e4e2b6dfb4c02bb1246398ade4c7f4a2
z18bf708244430a8e50c000281967c813ec0091ec32fc990b13c2f7e665362dc5e66f70d2e20c63
z192280634f15f4939f562bbbd1044065492966040599adcf2c7342d2bc31300b3d7b560b9a82c1
z28c6f027702f3b6dec7c3770665f0f5af2624e2b4cfa08fa3d68e611d1a4dc312cb9c3f0b667ad
z0f7758aa26ff2ebf0441a5aeb87d9c49798abee53cb9d0dc2fd5c5c7d9e660613653c80c03f2f2
zec056bd896cff0aa380a56912850a28ad36967d0bf8eecf1b101c0925a2268df4e60bf5c701198
z55b4112245d57355c1429b38b194c227f34bcab3078cf1562d72eed5cf2bddd4210f028d9bb0fe
zb8b1c09da49c776a718c190a1df3ede97b9aeff844baa5430e5dcc87eb6f07e1c2627e70669c3a
zcbe79813590422b9c12abf53de7567e3de6ac43879a683565cb19ef5829b8fd61d4f12a112885f
z1e79dfe7f794231651efa6559ff0d6e0b3b4170d226431e47ad48f7ae51ab071393334acea222c
z74e9708e081ebedc1ed4a9b869510df36b32d2b27e72f60a4f0fafafe9601260512ea0114c6d2f
zf42b003fcd946f5cda114c7e64105c6be67de9da87f8ee4af9d7f9df2e14199a288e100a1e6d49
zc59f75e123d01476e288620988e2e0d0c119e2b76433ccd21942eb040dfb6b7deb53d078b21613
z8efa792832d395d055eda78948f6f3bd9feb0f14dcfa79adcb9a5a6dab0bbfb3c211d7da09f956
z8b81c239ce79a34c7e83f147ce1b7a0f5ad15ccf3a1864d5ec30b0d9575c5bdf48985e26390ff4
z16c871bb589fcdc58a2fee253deb0753f2954b4919d761289af971e1f6d0c023a13fbd4066b7ff
ze389dfbd043455d259c83fc1251f41a63665ec31dc7791c0fdefe96560503e2f7e1a54845240b8
z4975c961c7f2d97970fe07c5f68b10c9594da77b4870309714d395b66c1ae21d399a9fd0460e9d
ze03d0d7185f199787ef637c2afc32559c76b293edd9fc24e789f29d58b1b6ad1c5a9f6689d5e21
za35c9de3c68ef498b602bef963df34d09e7d5b980d9cee19a3a5499a8cf83b7ccb6b950b02a148
z6ac5cc464646b08435f23156c4515e93ce6e298ab6f6c49a6d1fd6a12cda4c3307a8ba2f559c45
zbc72cd353a5e5118e18da91ac0f69c24f6c977449a9933744e0a0b996e27cddcc506aad3556402
z30fef8bd1173ce224a891fc428d19cae26475cfaa3dfa0489780b19c861555619f20e654802345
z1ae4e3bd1d7efa8fcb54464826b0c15795b4163faca6bfaacb852008ee975a10bc04b3b92839c6
za934f866ac9e8f02f80ba5251ccbfffcf9236a576da34b9e1504d1b45ba49ecfdcbebd7b2a9e37
z0117bbaac3869eb7f63c3ffc15e0aebdf7037928a3fe5939b16c37238d96fbe3bd8b1a9405987e
z28b0a9951ffabedd4273d6a26c09bf2169c1cbd87bff6449091f50a0de888003c9f5523168d6b8
z5c78c8992e1a3481dfdc7336d99436bc016a8d29de247298f5c76bbfddf8d9f14d523b1d66c7a4
zf7bd8fb4b20e782eaaa887312de93a75a758aba4b623422bfc24e150b23932c40c0c80c96d805a
zb603146f2b4b397f80aa7ffaab8108c9e2ad2b5112ac7f19ff6335d104381db9a0f7021cc280a4
z250e503bec099b530bd297e75f7caf2de837b40a92a50310d2001413295133e47d0b8b211d5df3
z9c1be9a895d84b40052a79f0a873d839a680e6602488bde89bd51ff1f55d815b4da4f0b2648ee6
zb3e15f694452473e99724b47460b99b062dc30429d99fda69e15da5918b8bd158a07f26e74485a
z3ad363d114341b83b20542cf597ead15f10d35131111c72f6e7f301040bbb77021c268a662b195
zb18f69bb647743b9604bc38b6a2c1ea99a4603d9cd0ccd1e0dc3eb70e3f73afe8f89cfedcba37a
z791efda718379725c795b312192ade26984ecdb0e65ff9396890ca8a16182614a14872ed2bc2ec
z4edd1183e96530df56bd5f802a392b510eaa7abd4aeb9daadca7e1de90ecb352bdbb382a36d18a
z63574f866762f564e025f994c00093514750155d8e64bf6bd19c2a072b98b65a5473be4effb79c
z1e16a9bf11123ac0aab11656f006e9235a04de9607436377ec813c1068696ac9681316eb8d421c
z970fdf7a0f8252f96438c65aea0157378ecb6383ffa7ecefabc4e373295679a2b7ebb351ec198f
z456889b4ddfee0bf072595fb7b17335582a7fe754fa8ffa6b2cf13133bbd230c3612052ffc86e4
z9db7f7e1a2e136ed7c8932c263c5af1cce9b38c07ddb71c6f623b5eecebd43d9ef636f8bf513e2
ze86f3e9fa5a90b24164370c1ca5a4cc16adc7459ec47656f0433a47834a9a6c2a646026ff1bc04
z784d878672c711555e5005929a7e0b5444a76e67b8eb326ee332b589b7efab93657116b3708b34
z1a9c5d82fc74c7c54034f81dedcea69ab0f7d9328f7ebb8b2736b66df0807fc7d136c9d5418c4f
zcd993aaa1bd410bb4fcd356d7e8edee8f010201a670744c0d81db1e8314621fff34d967b1bc826
z3e8a6f5d3f41d0ea4e23c6b01840b09a83807658106cc970df9b093b819fe37fcd3c6393cd6b35
z7282156fa24e22dbc45410c468f0620ced2309a5d2662876257c5ec2b6fdf6e84c89f4bd4ad4f5
ze3db7cdcd7ff45fa77d08187d33601403f1c7656a102779621acc2023efae71f2f1dcd00fc8541
z42c0b1899b250dc802391d3f51a4e45d77e19e52077e2a4611f22340808e5fb2bec108af0be1b9
z9021e55695fa3a3843136c0be687d2cfadc5a069c54fa2e500f2f83edd90240bdd2cff87275776
z0e59404fcb02a034388c468842901be09f5d2fb885df166ea9ff8907d87b3075cf7d7751663061
z58bd4553b7586a38f158ad216780b7f1b29627e98079f575fdb126ec8c69fce3ad1a97a51a661d
z01d28920bef8399cf4dc804dc0e832c4eee09ee25d09228d3c0dfad0ade363d1492e6d6af37b64
z7bdf6d8e91d3ef9c54b54527d556c7e7875b532a6ef1264f90688319646c0d8947a48731de5a63
z76103c636f647e52bf745e56e7e3b08339fa8ad0d94d75b8320e97bcabc3ae7c7c2ddb0f290de1
z46aec3a93afccd375ed380fa61faef3ed1aa67015bc70e58c81d1e1919e5a4a0dc9c6f0973640e
z0f32e53f15fce8dee2b3483787797f5a32e48e48810b641fb5b57c84feb0c33d2a55237e9aae4d
z50df7140e8411ac2ee8707b0a91162efb7261cef7552f4ed16a88d26a932ed2e533499ba5bea60
zd062f2f977b4974d9fa5130177858125dd437b72895ce61cbdf4162f02b27a14e885bfcddc3343
z978ce2b535a999de592a76de0b8864288ef089a8946803c9579fd21c77b5821b0a526561135fbd
z506d1e070eedbd2274781b1a3063423c3ac50f1710b58914e1e3df535859ca8c8595f4a55ad2e9
z02e2ab9ef1d835776335163d35917ff33b922c566593183a7d7f8067c566c3e9146fdb9b2b852a
z7892ecf0473a40f9ff4fc84b4b58856f9705991161f7c7b580d32293a51bcdccb61581141e23cf
zd03b91ff8dadab4787289596944ec0046ceb8de79c66fd5918e0d86fcfc48d72bbf8b43cf5fdc1
zd0c5a57cab603c3ff3690d7d9ff761e6fe1c2c89d7e9337a04c02ee67add949c7809715b8318d7
zce47f0dab0c81d818af1cce571e2677b01f0e3b4cc9909f963db15b1707a578d1a7d656d43c9a4
z6d21698ccdc5ef002213a560e3de481aebc4d95d0b88e0e52490250301c9037f38b1d05c9b920e
z391abea34e5297ae0406093062cbd87a68d395b882a663ac1c5f36839001d7dcf25c199e38e76b
z94f02a3e8427c4b430c4f1ea1bd201a8667e39a78fa325bc04ae1bdc93c2cb87bbd4dc654fa483
z779c4d222601750d4e405970f036f719471db31b8f3a15e711b062f9e346740cf6cd915cf5e801
zf121c12e5eb63b8ffe7024936dddcc2e63e7d6f3dec8078f44a36b2f55a3593aea3770d35ae606
z5ff0f25e294a4c9037dc1ca51be4ecc02fc430bbd425838fc288faae9729a535e980f54f4e4caf
z3e0f49137c45dfff048eee27df35abe1b9f9ea92ff68c31cfdd46d39cfebf89e642fd09cd84645
zb596173f34413c5b5ccce1c5e44f1c762833ec7cd5004001d67ed4f0c180d8f690f8996d779b75
zb67a3735883d516df8a9ddf42bbccf0928d132b38d3cb783eeac7f902038e589910f76a1161e30
za81d023f8df90763ffb525389fa7fb7916a521cc2c87e0237ac7af157d216696da66a4015a6c60
z7c12b043aa75a6fe8f34d71151c7b331b03498c45f7f5f55138574cd1f37245b5cf445c8b21cd6
z0dfa7cdbec8b40dcb0ac5ad8de0c510a7459c5c907c9310516fdde73dd3d6e0fecf30d63ef0797
z7d1a836a48e9511a49424ff23c7b4b6b5ec396e1e3d54b5d8b296453dfee06acacd51d083e2d0f
z5e481d73188dcad2c623108dca2677d30ee12a01091057c58e8739fab53295e3411d7203879c50
z4c0d18803462d0e4189a4689ba1dc6584661ef32168679ee88e0660712d64f0ab09172fe41c312
z35f715249bef25758d08c06016aef628bedd6ad9e0ccc9e0974da22867c4a61a95555819bb1c57
zaa5964494e9e8af0960168906fe8262da18cd10ef7e8f14ef061b3f69d392bf7571d1750c19908
z7ff4e4a5193325dc8c805cc934c40670570bf38cc1ae00ea4fa7bf37469dd2c6c50b691e493630
z26b84c6bed9d6050617c9af9b0f5cfe816128d4544c9c92792782ce804547ff2e549121ac5eedd
z5551b374cf11d8911b6972c4dca9c3bcb9683e7b4dc51e8dc9b0d06e8f14c68c1936f229152719
z08bd333e08ab64d1289d7eb71492705f624be137ad8346571bb854a2b259dfaf7c173c66a9aecc
zb52e26fb4ba5649e8a6a554bc884c3e5fe32014a5596c80e7b498046afe55bec5486cbde5cedaf
z6638dbcfe31d7d1cb43100476095104459022898650d608d042d832847befc3d3a569236be3fc7
zdd56d9fac976d73b9ae72254b21b0bae1ffb48a89c95fc445e87fcd7ea351544552a800897156b
z8ba147759d6d1076de969a89bc90f86e69b6989b750a757aec3e2d0185e5f4cbbe2664155cafd3
z26cbf034a418a08267bb380d1b56edd60708d19e06d2de01c9111d78c609c7ac8ec13c8b99ca0e
z4f1a5e93e6de1e88517817a7f31e2652d363b1f8d654f24e003a483a80323bdae607f8e990f733
z257a56dc182fb8f8e3a64e1e9634244a0e32ec2d4b7f0226d453590d184e4a0e31028d789b4bb7
zc1d368be6cd852e491d62381ea16cc06ea1bc16966dda935d866870fc63a4b7c3521f786b769ca
z2ff0c0150701a903bf7d01f24bfc8804cac47b7f252f491409fefa48c29a236fc89c84d3525451
z97b8022c303be1c491b4d2fe7fa4f22e8760bbe1c26841b808286effac41100530a6f01b770b74
z96a6bf9567d505a88d5eb3b2322a37bb37324df925e71fccb7c192c0ba005bc166dd728ed67ccf
z0745a80e2ca8538802490b5e222d982a514abf935e47d6a12e99bb5c8c75c3b68631166c50c909
ze44cd499f304e3e39975e35d6be7a2e9541dfc1c05073a7f1c73bae9097fb97ba501aaccdeedc6
z9a3514b3f7d7fbbb31e6a588acc35b7963f6079c474c5e56662082a5078220fb6601102eaa36dd
z5c43adfab4d5139820649e2c26382b57a5a9c57bda076d3e7107101cde00148d15c05fb286aabf
z21e2b9ccf7590f3b419fc3ef762402b7b8673cc4570fcd2102ae286d6e5cc159d85ccf80731905
z2e913d0f08158c17060138a9fc898ee048007912f8373f3d548d0a7cffdccb8dc8faedb5c7cb0b
zaaa68e5b72924548c452443d5dcac3ffee81f76804ca1112781af75b4321d167a5334edd2cfa48
z26386a237baf1d49710bb995ea150182f74bb3ec94f6430508e64372ee9cae0dcdd5c226122014
zf5769fa4af832c947576426445f1291ec5a97e36294691d60d2026fc16c1110b2a5505fee61f24
z699e3ce207a67339efc1f80b7a66f95aacda46c969ea6c6056be1f43031ae26deff9e8fcd47113
z35a7e180a9a1abd229553c5b0f73bdbd813a93e7668aabdfa587f142c7ab2e1731661054c53dc6
z24142f676a036d98bc8df00f60d5399f02a4319f08a1aa7e9b24a2f8e050eadc4b73eb1bef8785
z9ff5ca581fa5d75c98409a0cc03d46deb76142dbd7aa7d0e0553937b31c5d0894da08b9eaeb7d1
zb983b824885e98691b1b662f0ceefa9cbea770f4e4044f7eebcb2c6a36123f8dba8be13bad13cf
z00a76df71c8659b36bbac4bb2d096944670b88a99b3734d08d2655c8a39b03c068fbf9794f3439
zde4e16cb5aed1f305949b669405bf307c48e3780dfe69dd7e40f4dbd60da8eeeb0b17fa85e1aaf
z10bc75262caa5809e6d319534de2f29bd520f03a1bef309cae51bca717b45ad21efdd394b3dc9a
z26ff26dc3e131fd61ba909d474ed0b45ea271e18959639c4196db138167aa665178b8b1f8eaf40
z18113e3e4d857ddd225a94448fc3fd0b62cbe8f1b425d87ee2ee0314be1e6a0d08ffe3839209dc
z464a60e0e0be81ee53f6a0a7f3976c9ccf37fb353fcf581452b7cbea647184ef6fbe339871ecd0
zd76ccfba65647b75bc666eae28c82c8c3931d3d9f628226dd317da62c8e4e98ab6253993ffbbb5
z5d826ce2bba8d7dcdc631cd942c1eac2751175dc11d2089c065a480e61a4850ce5f7f98f2c2dc1
z552dcd26bd60e98b6367ff6b2a832d277b5ffbb4fcf5af41b0267d41da4cf4dac6c2599e69aa71
z80bd7a671cf577055944594fc6301bfc49e7ae3091fcf2f22d8aad70d1a87af02c7351c0161ad0
ze06968e4be3c35ebee49289e5a1f7ec5de7e59f0be5c1e263139636b2d41c050201dd22e95234e
z8c0aa2e9fb4b4dbc840d14eefc0234c19cf8e9ef336338e5f54a42394689e814c4568dd1e3e2fe
z6fe3eab91d92dee58a9eecd5e0e473899afc7299f41c42bde8ce4fedfc76e368bc6ee20199e8e5
z61207a0b502b147e4209adb45e07f16944cc66857e8cbb97551a7a1c4f02fb1f7124628561abd3
z74522b1e10779b545b1c925e5899723c58aa4fb22bf632a40d18b98b7d934ee6d84a615af30136
z55e9bac19d560280df1d196637bfe9fd7cb9520208dacf7ee1a4deeb4d6479cb2963507a32bfc1
z76a630aa128949f518bbfbea36a3f7645f9407ca927949a5d831e9b8d4bf48420efc48dafb1145
zcc35ef6766cda21f3ace8b2f8eb4ac5ff23d15ab1f5e9928fe6a6a748108b13be39744c681ca81
z9596dc0f9219a940a9a8a27fe10de46c57ad3e385f233564757beb96e009dd229a11bf6d5ecfe8
zb437894e8f8454652c836945a0d1ff7908496134fe1e1c934acca3162ee34d11fc0bdcaac8d3e4
z33f3fce839e8692329d731f2717b85d0afacfe394707501bae873d2f074c3e97e95c525fbd9837
z2f4c5c01e9b92c7a2dc6dbbbd59840da5d3db59459b8fbfbe185387fad90da78c12d792a0bdfac
ze0226d262b03289ee2379dd18c8c45213546d66cb5650502f473ac8d4bf2c9d398a98953b61e0e
zf01e63b88d5b5c70c94ec13c2559bb571a2ae80743523dccf108ce73327466a597aefbe87e7e40
zd68a5103a8cc1e579491c7901fdd3811cd047498a4ed7e61527ec6f1e5b780a2a1f77cdeddbf6b
z892cb3ffaa40113e1832da35b760c8ca9208d9b4e0f1aa5426116faf8b540155861e3578eddcc6
z24c0ef522e931fb1492b3f8a710446556d1b57a8bba6a75e6affd815a73353dee8adb33293b09f
zf72a9699ad7dacfea3f0409e71992a78d0b5e9fafbc61aaa62f0afdb44b3a932fab12e9dbd30f7
z5858f1444cc735783954c371d3eb7fdb18547e854642c08577f4ab8252e056337edd245033091f
ze523dec141d21270487130c626e3736a4e3c39ddf334269954a9d3d1ecdd30c8c7a03458543b71
z12029e1a5b3ca355b222c569a728000c667e2f94e319b0b2ea354d8abdc4519c332050805be64b
za8e28d0fdf9d481b5693db7a7de5a193fed01dbc633afa004c3547380eb847d1b37160930508ba
z01f5b6d3d3bf96b6864331efb6bef5f34a96d7959e65d24d3df97983a2292e1cb8d926bbdcf1aa
zb4a5540af513b520d78c3789fd69c8b32698cefcd9b3a5b9061d8daf115e8f4005f99821129c89
z82785f4cb51c47dc64783d0f22522ead92be031a9c717035aba01a355753eb051454317db9dec6
zd0ceb689f69e31d605b43c89128e217f12512f7568200e8b39a58fd6927aa07451992a0c1c5a78
z6811cecb81616154cea2064aaed5ca76d3af643a173b4cb3b86fae37b305d3611317500b0d6de1
z0a7b0a18eb8f7f14656b50f7b2e716382be04ab1473d5a039baf7fb069f1b60d45b9e9c026c53a
zc943a408a5f453d25dd69456c0c17207df06edf35867b892737d0fef60c365efbe5851dbaa8f93
z4f921b6db6c5c68f432b04884ab1d1e3578347cd5d4b01597653b05dc86609c88299802f64a0f6
z3a56d621426a35358770b00f8844a37acf8a2bba24b3c425d1531b46b67dfb1d62e07c6c74d618
ze02e75b82223e73c1314836f5902cbb1bec4d1786c06d265d129a25966ede56c169bff3c4afa09
z7b1d5539b488717d16bc110b263d4c7aa2a4ba13868e52cedcaaa3a1fe038ae5a84c4423064e36
z0123ecd3d077850fca28fcf8df5087bcffed5a79c568da2c9de620e926b8d71b090915782bb84f
z7615e9b228f17e04549d31b0d43012e1c1ab55ff087953cf186ba808cc4c04cb74eb10aee5b780
zb938af48cde6422b1a7602f63cf0577fd3471426dfda24b2be38fbe4c46a25401ebb512e4628ec
z16689d2f99c97e48152b888289c5ad99277a113e4197787e6805a600349c934bf460c5e09e3460
zf7c30e46cf9bb23e31ba63b69f8c331a53f32fbce2c8c1c11eb74e1f7a3e6fe498c088c054ae89
z03274d709cd5ac95ea334b9e32e88a099b62b476a706478aa1dd81351941bf75967a43ebb2addd
z499c71e9e30f05983603aa4e5f2637abbc7bdd9b2a2b74e863c5487871c2ee73482995d6acfeff
z64b3e87d76a99948a68ed9ecc1e8716fbaf66a3418c9e5be0f5100152ff0d804339c10f7dcd470
z69025f26b52893c2932d89f81d25388b8a03cd43ce38ec55f02be31387b427242cd5675e2ed534
z93b6c2b55ba60f5d88728be82a622983426bc6dbad0c3a487f9c773f456fa28cb617f7c2ca968d
z14fa420feb3db6d2c028954d103b12fd9c993ae1a2737cf4dc5f664c21455bb6ccb33070d04c44
z811d174f67047e3545d612ba2092f6280340a0a2c985a25af889c34a206ccc3528fb8fc3f98013
z2197a462137ba0d4621aab41ead6ae9980b64cce52bdb55310e09847c113b9c0ee7ab5bc7dd962
z38d3a365d9573696f57b84adfd6050e193a9645472e17e2c9d947eadacd3b5c94013c0df87ec91
z83e2b295852873054ae7978be3fdf03923260cd5c873e939daf957d1e6e6522cb98b825951d9e5
zb2c8ac9a38d3b7545f002843863bcc6de5d579d3d6e52ff7a901f17c17c00be3fa862f23843592
z6c092295478255bf842d78aa581600295ce937554f1e17de5b5f17817592029634792be7386106
zd8a3095fed478ad61ce96bdff3ca10d893770af7d62f0c2ec1271ba7a630eab295846649ceea60
z4481529efabfe12b768f703f6604ee364269c3c403cded18d30ae837d8af6fcfdf90b0bdb992d2
z99be41412a09d9090e2a544cac6dc5876bd1f24bd1ccb302f6bf94aebd2cc3f83184bc8e2356d5
z2e2db70ebe33e00a3b231eedf8b818f4e3584bfabb308eff9d0115391d7c456c7ab4332b6c53ed
zfad907926468230221324ab8ea6f112a226a38e329031168b073e4353d0dbcc346da6d3c339050
zf4553b928f498586d378d81a4a4421b10b7309bd8ebdf86ec5e71db9c6c7de3e88d8c1b7a50d0a
z4ef2c36069557ebd45701bf088116dcdbfd6c90c671378aa14f9fc0720924765fa3fdeeb73534c
z17e7da9b3d588f023ac7d0f853e77d715bcd680ebd34ccb379d13266a039b7b8893211f58e3996
z6cbbd9b92821a9635651241ca9ff8a0482b6a41089f745481ae57819509cee94eee565c3571167
z4e341c4062a3b40b49634ae1211ce011aa9fe51c28970ddad6a10aaf429b3574953f8533c14ae5
zd8da14417eaf3ef072b747e8b7524fed0bc1450ba22b8f3928a906f1bd504f87aaf2fa462c855f
z46a8559781c7ed26a8e36abb5f6ff8f3421980f36d058efdfec51075b760034e3dc3303cac7929
zefb6a3a609f42919928b427aff7e43174006f28c3178aa882e3558222bf471827c7434b450c1de
za8b3b7915f0642ed57c2c2d5b2247b3abcb63b17b41841244b3d05f4b2b288aa8fb7f63c7a93dd
z7303539dd3c547bf1e536c25a647b3506be86aa6fcdc553be6d95d8b9791e1d6f4e9f5c727f58f
z7d5106f8a0c5ba0621ad159e85cd33f39f96d6d641f4ab443c20ed0ace1ceb52ce34ecf3297ab6
zd050e750871dfd3b9eedbfa4eac794ad897f2f15e0c0510fa2455e0db32a8b17e482d2d252556c
z14a74e4270b08d7e99f3099f1d62fccd2e3ab564ad0654b6cd18f05184c75b8c04fc0d9f7157dc
z5aef40b80c040108d05076e904bf3022252d06f1e848d5db9a76deb51b15da5ff006a9e8d26ae3
z4e3cc8247c9970f165f6d5b5dfafacf6343e18ea444dfc6ff56be3c02eb279af72ee5ebff3dc6b
zac788422e3819580e73bb62e08b11d4298ff95c3487c353fcf0faedf94aa691c8c34fe7cca1141
z98b4b186af7547ab5a907b8b31c1a4f7a31d540d971fe829c7abd9f0af238b87b606c0170c7c89
z24f0b49b2065b52af290091164b2d58e2fcc2bcf24787e7d8530a882edc0fef0e194fcf91dbfba
z4fdfb0993d07c3747ca2ad44be64f9e77189cd75d0ef8d06e6ec9f51a7cddafa4cac5544d07462
zfd0f0043d855b0bff0ee6c9053db4e66aafc00922a555b824f0ef4b74737c38779c472e4690050
ze0b5605ddc37021795f3c1909b67f8300acc244d398f1acd957e52bfbd920219dc8a175b3a94dd
z20d7da9457004cdab4fd66450197793061c9ca668cafca13608baa94ce8f898a0aa6adb32b8ee8
zbf6e89f4ba16d981f082b922dc870279610272d3ce9a3b8a8abc3f12cba760cbd774aaa79f719b
z139340fd256ac9c3dfcb13f9e6fcaa479e93020c3cf34ba7b44caa16dd99b13089fa0b027bc900
zec481969990b286ef586ec9be3728c9c4b7191f4b0dc6d110d6876fcf61f87064c25e63ccb8a47
zed74a500e35272a899a391211969358ccb4c797fd6eed097fe083be4db80f64d1542d9b2b63522
z6efedaeb7a6643b60662736de961cd1e470616a3487d04417bd659e0b190d7b3c9c95babbb3eb2
z3404383e52ad189675cd7cbf12396f57a7b453b326acb31b32fcbe5731b579acf9c7c0dc669552
zc501df3af1ce676a5ad2d36e94c2f5e0136ee3a7ef24747483977ece8dfb6ab827e3af26fc9862
z5ba4540e18c2d5cccc3a94197e2c739b4e91087db8c02e5234039afcae494eb498298461c2785d
z13b5f6350124dee1adaa2b0d4a3bc4e64197fb064374b192b6117043a43d6b6ed454b19fa4312d
z5e2b15f563eafb3d4c8da9a8f7d2914ec1c56cb0a89829da9bc05af70fbb56bbc81868f30c1856
z2d95a5508d3fe2a4966d45453a410bc2f6d59e89823211ff7fa0347767669f6fa9f18b3dda22cf
zac02d728a3a940e3c46541c573e44b44ee5e316d45b9b0b45769217fb751c773f756b3f8b662cb
z7408b33158eb3ca4dd6eaa4ad034881793784835ba061e6cf2786bddf3d8ce628d7fe0fb53a2ec
zfbcd9e1e7f99cae969579a462afd71eb3034679275810064333890942f826228037ccd5a5f3de8
z68b09fa0796d8bee794097025741616bae9c6e052c832150101394be5b2592d066f39f52f640a1
zb6056fda28882034e2389fa51adc5bbfcf990a7452f0dd72566ea0aa01384288bc3998d7976b2f
z377b66a966ec9097d66de38e33d25ce1fcfc2175ff375e9c10d0451805fe5d9ae92c9c72b5aa43
z016eb96e215eeded15c25045dbb33ccab4cb2d27a2f5b1f19bbdf65037a44837eda0eecac6b986
zfe6354df429aec665bd3d34dc817d215b0ffa1ae2bdd46f143ab05a391d2a6922640160830d825
zfc0972e73bdeb397ac8286c9c311bc9f893d58d7c4dff4512846b8bb71d7a2e187b4898849e1bb
z1202bcf48b452966475fb1a6f27633bbf274a7c170c2684369d62f6cc7f0a26a27e195ef695554
zbd52603885644f718de69ee626901478a3fc9db13213b4a5f5db10887cab5b95ba4fa0a763ad03
zf58510cbd0f01a5e40a065ad93dd8dc1cf6b12e58a9c6fa32f5e7fac5160f624a7bd95d3c798e5
z8939a47baa1477c10b4c45f92f9c1c304a9f1d6c20452832037c7c6bfcffb628014f39e64ae1d3
zf913ee4791680fc7e957d4fa153c4eca142d4d9dad91ede9c317aac1c33b6df97caeb593863e68
z193a61a3ceb763eab362b647eda874fbcf39b2ba06c46f7df4390d4cf36f384046804fc8c91e22
z75c29a7e516293de584c976f069cd07153af3098823a48bb09517e329a2f4419b55ee9ad96963c
zd70d037c02d66d5f1d101764e2ddd4b599322267cea108389f168c162db45a6a2597e4bd2b3575
zc644db84422b7a0ed8c1268921a8fa0bb661ee4b4d1fd914323cb990be5a63a542c9f89415308d
z6e28500b3f1847e005f066dcf6119b77c8c209771123d2605a0ba2239073fd7b46ade821dcce6c
za540326b8bf5477bcc68a665482849f6485f569878397f1716b580d7ec52dfedd65daf5fa107ea
zf2c99957327d71d0fc43e7212248ebd43399803db54c76b5778730e3fe566eacfa962fea0f9a36
z4574f953d875f4fda0ed052d4ba5dada428923a1f01cb26e627ea5b20a5ba4d709952d71c4a8c2
z3f026cdf6e7d4e115a8d42abf9a66bbcfdd83b377a85028dbdddc9d3ada033481b55a11e1bd86b
zd353504a515c9560f73ea7fa54e4d30eff5f9af41ac5062c8886a3fcb371f6836917eb81143cdf
z0980dc6e2557edca74c9c2b30d51487eebca824ded07131c0ab27d712ce5f7f9a2d50f64b23c74
zded19a5c9821ebb4bf0d1cb785f7f84aa731cad44a5ca9b81e637fd212e499e3bc0def3ff19feb
z1981aa0c3abe8fca5655881f9544573f7f657f3335597c60b4cc4ed16496eb3972bd1f3bf8bd0a
z061b2f0c72ee0559906dff1de662759477034d549dde545f2effa34671e315121d91e27e9f9682
zd860e5dfbffd3dda8c0433a2487a96829027e61af1bab75087fc684f97265c6a731a14d61e8f9d
z9613d439ca2ba79923fa96489700c4f77ac5188824a86d6f1775919664ea2fb052432a54e22587
z9b283d6b3aab38237c7d9e59b682c2ca7913328764c46a1039f2d1479657102edb141a8cbcec50
z36e990fcad6166a64dc8e3dd00341f5dade1b9b259cf68bf8170e4ee3ede5dc510dd66bde48cb6
z3aeef9233a307a0541efe753e4f0b1410faf9140a6a738ca0cfc3d80375e8565bccf365af5cfcf
z7b2a479f4658dcabe3f3d800000b4711944e61e98d74eba04342d870d86e52e43e2392dda01e69
za1978102a8d92bd078fd31f0fa654db8077b3ee847a3b3d2ee9d7146f7b47a6a10be94e2589269
z05c5117498f4df17f3d7a3bca772d15debcc7dcff7d33fb2a7ee5572a31ef4cfbe3559ebbacec1
z626fa79e35ba1dde76210eded39c4ee0e9d3f4d65573c0f3962bf1f41883fef6e5dd117a217e61
z4397fe0064a3f12b62839d1eb87a732a4518038e7d6d3f7ebe8656ad485e66677e3962a8555ad1
z3693ea3aa39d4e254a57c130c5590a54b3add25560ed9c24f45ace9350d54f4fee7bda29e1e090
zddb9704877ea6d18ec068c106c3cc7c9860407bcd949f11bf0b992ce8a246bbc91e69a83ec4284
zd265053de7b484e244ec56407e444227e55033cde87224e6b6ad626f3edb8a8776f62dbfa782cb
zd597d80473042be629bb5f53b6ea09b01f58553fb076a8ea6cabf8356f702fa971620599c7b987
z9212301f90c997c724179284a2762de0abbeb136b3e810db63bb95f9888d5f8331305a454b28a8
zd351921fe8526a32ba5defb9ddfe514b8d6d88de4fa4a1998dec94285ad3a04002297813933c06
z5915bf135cab02ff72ef0eeb48f83b2e48f28e5b45f50b1edec317fe1afd14ef9e6f10bb450ebe
z370f32a7704f06f637cad6642dad158869c75ab70b7bfe40c96017726998de2f38cac3ddc92921
z2e494c74d0e02ac3b1d810010c7573f581980fd91e2d5fa8bc2b80761f72902918956a0a953aec
z6a1154d38f06d3e68e020dab27d7ed7b891a859eab4429debc7844e73bd4f1629a81fd0d8b05a1
z166f42abb0eed10dcf6732a534ab175918d7d3b110a9f97dd4c5ef15d87a5e9890e8615370d361
ze7741b8f763736fa4e7abae3bc6d2fb6e3ead7dbd2423a135bdec6e5dde36223b56435a212344e
z1fee281db5bf10bd95ccea433ab7b6004c8cfd4bc8e5245c5f8ae54655a1983953069c4e179808
zf87d51a17d25b660a6d46ac325ca5076dcea7ebc04469dae9fdd6df7b0acf7cc725ea34f83214e
zc5e3d334e0d66768a9af709cddf8ef2007c4ace05859cdc748574ba880b7656a7f5e79fe4a0070
z7923dce78de7ab395861ed17e162790ef76452720b44a8f9b758629fb57456e8a7a34fd8933660
z1833760bb36f3dfd92dcf9becaa8118ca952f351ad1964b6a9eb0e61f57efb22b9588e64c1815c
z5ef5663c8a3b3dd03682964c01c56b69d2a617e060619abc561c0ac23d376eec9f613bfe3aceef
zfa08943989b7e86873419556220f04d065cc6b45bd823049aa641415ceafd1fbfee7adf142ea83
zd3510b2a1d4cd0e542acbecc7e64e7e670566f092ca3eb348aed36357fbb4c317a21f2e9ea2542
z54094eb7815b5fd38770533ee087f2e1987623f68fc01a0313f48a576d6dc9ec17340958d5613d
z29a9b0cb12f926292e239522e3667d9f9dbd1fd4b098205a15b55f420f189d9fbf65f06408e832
z67d2350fb0021994cc43841b7113393367dcd96aa277a468c0584556d0d0a73cea46fdbc6d6d28
zbed4872b5daac46525881171fcd9817dc91275c88c9eb0687eedf286f6accae7968ce32b98a571
z6fe2a86cd924c2f788712d3faba39deabcf7a83aa4fa740548a0c8fc18724a6e5c09d6d1276536
z86473e685f3138d85e29fb251465c7ca4c397915d00d1c183cfd4c04949dad58413ea95e5d4f2f
z0255bac9d98f20334fbcbc75003be5b85b2d3f450cd4e7a6ffcebc7667f4f3a4835cc7ad092e91
z422318b346468616458681975077c8d4ac059d64761fccf627536f04af60dce6a992936eaddd01
z9bf97fb04ee2d56854600aa83976ff38222bceb412deac1be5cc05519aa06f83a293db92b51cfa
z404b0f842b9ec3a5cb5a9ba25ce2e1368a9c5b78de3875d8ec08ad58c49b19aa95b47ed3390e21
z58e5bb184e1d0467a7654ff61489bfb18e36a66f0e006cd489de30d62d3512cd54b3fcc2b01721
ze3f2a0748c27c3d234f012160c12df717767ee13da7646c0cf5b5e2b6e69a99b5d78d33bb40cfb
zbccc4fba6c1013932c44fa87628449d3e3207032342cf9e541f1dcf80c168cd92722c45214f9c8
z1c40eafe0dcd8940579a0d4d4fa57a6e3d0726a87635a92d5f230c67e2b55baa20039ba8b07235
z8426d3fd0e269dd818068e0fc62a0d0256a87b5c256af79e14628dffb251a2d32f867f540557bc
zca6045586640738c800548bbe9da05b6be4f0220c9278934ca3c4762eaced9f3413657a79084e7
z5aa8a4e8b303bf85d72c2e221f2addebb8b9f92c7b0de305acd35bc6619585b601bc8d655a4194
z5152816993ad615687d66c3bfec50f32f05a33a9c173b62ea75266e3c1dff44f734a41a53b9e44
z8617d608a4ae7efeb1dc3b773dc67795182aad44359ee0269f7d397e7fc4acda40f00697415bfe
z284e063b359c44cd24b2e40e2b3550ba8459042c876be10d8c0dacc40515e266014c2aa4b13c5d
z17203fb724e91dd0c430c9abe8b7d30c5f59b29be1ed7ec35f55a82fdbc31837988c9f123a72c7
ze36661073f886285b8ba379d5f9672c095bd836768b5fd862820408296353b62d6501259da7db9
z5fed7fac1b6488826e564c01eb1fe82292a448ccdf25c674bd2d80a3281848a60bab8a47949c7e
z0722c6c41d8664fe1fc5a03e8b0a8bab9fbbc1bd71f2b71f49c5cd606132fd68aa7e9c06f3ae0a
z7fcf466d3383a98eb45a515a6bd0ad9d13c0af0017e885e4d173b6b20771e1673e2d5ec719dcbd
z181563da4764ba78003ddb7beb1cedd098ed49b9aada7799836476e09b21e0c79b632931f93b35
zce9e5c81df5dc4479232a9625db4168eb8deb443a45550c4d632aa01d2ee55cb44a1aa23a99057
z03ca46e32d4474a5af33cdf64fc7a084708be6159a1b1f04b0afaad71d47c3453aec13985d2244
zf297bbd7d1066be97b450cd26cc1e02d042705eb2c4643a216041d2795e73202b3eb55077021c7
zdac2bed8c5789f2eb3dd7b95316b7693f6784ec9dcac0386573e555227aece56ce2e1695f20a7a
z005eb0c92e5e2018226e529875034e5600623350f176a9f4934cd778bcecb7b7bcaeb00fa8ada3
z0293f3ddd952a50d7b5ce8b51b996c6a04898b3261204f8f9cc7bd65a1ba4b7b3c452656088400
z224cac66c9c585f3d2c2e8a4b504aa39c9878bb6af9a7820bf973e46e8b5145d93d3e99c929900
zd5ac9aeb1b46c92716541028511bf7af36ef8a98f2f5444c509e4d35bc4e22b959b7cbf96ae621
ze6b0e0e7c9164ee51da4d870a0db9ccde88ae08d960371c5920eae541a46bef6fb74cd3c584d5d
z8ba9ddde25a2937d48dc8ba8e71d54e485f13fa548a7944e615a33d1c19e3531f763cf7ecb8373
z88546502538da4a9ce3f0f9fc24101187297cc4f0793c8ac16aa425fdb1d9988bf8198161bfd30
z4cb40597161704e75acd271210d6cfecaac9d373d6cf04b4ee5c92837c1fa4a0fc921f5cb55466
zc84ec31d91dc1541c44be2c071e313724d5f9ee45f44b42784b2de47d9a8c6d489e4b31850d571
z0453508d324c161ecd6b875b3425709448c3c914ff30b96e8b808d2641d4cf7dc75cfce24bebe3
z2ea1083fe8b1844fb1f7a1389acc6c4f6393ce11334c3997b6008ca26cad0ba24a56b60fa0391f
zb6abbe1369fc4f29e8f94d2f1068f140bcf9e3cbbdca022f5388a44af67eadfe4af5a54babfee6
zc27f4a415a71a3ecf7a1896516ae430eb98a16823c95ccf4ff343c85a7866a8e868dde4bbc60b7
zbab1cd6bf19729a6423249defc4abaf7373745a4b22a15a64d50b3ad2dee46b7ef52437796eecf
z5a40eace76bfea0f458e7c7727152f2910ec7cc8828c6ec7ebf2c0650ddd1075e73331b9c3b4ad
zb18b68fb5437e446520712afe8654341cd33efaf57dcf4a6fe093ae49db48588ed82062c280fc7
z3474fbecc1d88dc453b4461c95417935ff0440d852fdb4d8440eedf6b40c8b3a031e69b2216699
z068ce5f80036c1c2ce35aa69a3fba6d165b83f630501e8e7d634a055cb6cc7dd2d5d04ece71c85
z00f2055bbd904f1a56830eb033da8c9716c1e358e4d5507ac12989bdeb40b859c70440db8b9581
z25da8d495bae003a70cef75806ef05ba732f5c56b4c8b7d79c07dd4fa2c817c877c30366055a08
zd1d7158e00d112beeca8dcd9f32c48808a12cf61a2f96dfbcbff37af817411704c25c25cf30636
za819ec67b45c970879b86f2dfc09d81a3c408b42373dc434a7673086b1f9c0d555688b01b37078
za8451f1e845aad5610b55d1597a3f62880ac4122bba0fd86af009bd476283b5e2d3af2ffa755d7
z1f282f9ac01ffbcdea9e69d7f27724ad7abd36ef0de43803383b3101c8be246f1b46c8e6d84b02
z5ede546fac4bbeb8e6c530baef557f1824ac3c7478949109cd1c992496ec3dcbf095cecaebd684
z13e46ae66effa01c4f6d4af4edf4055b0c0f5d1e8027cea6b6055b308751f5f0c6b211fca7638b
z586944a773ba35158252b4c4d4deeb4edac76cb5cae0365463b13eb9b97732f2cddd9e17ef248a
z7434e27918649052d464523410b9f4326bf208e0d908fb0f115589daf6d85a4ca01f1fa6b0ca3b
z5983527a1983c430bc4fce2b47cb34bb88a3bb05f716abcdefb0eec6e0e5796ec6cf6f0f42f6f7
z4277110480cff5de0e7dc111d871afa97d4b8bf3e30cd6bce53c9490ae3bf56aea051630bece85
z3c946d23e5b194c441f9e60bbff796228f758ce849084e533a47bc17a457405d707cabf46593d7
ze903b7a0abdb54442f0b93aa8a28aadcc8bfa08e86450c9ef2ceee56ec3d02026a83808912b3e3
z9081040492938d7d4704f46c2157bc89dc5d443b78c35a452a1158a7de9fe241dd6e9fe36c89a7
za87072db57be4af5780eb99287151579dceb3a0e3420e18b04a314c10673a46b1c9466e0e4501e
z203198b05bdd9e64526a52f31e10f5c3ac62477916e62f578fbbbc362827e0df7dffad6eea0d59
z2e586c44a5d6297dd76e45c5c7d77197a4ea1738a33db44dcdc7d244ebb7cdfcb2e178d822fa29
zd8cca665dc3773d7676d8e4928c0b35d3395b8a2bbe261a6b6ab8fc0380050ed7ac9ef403241f1
z2678598089db0cc4dc46172231089f4feb47a0fe0958e8a81dc1113471d421577470a519d3b3c9
z86532d5aee95b60773930b80177a346b2a4d4583271ce0e0a2a75c72a6b9eddd88659e2b803309
z0b3c095b7949c98fceb6dffe8796eedc5558e066684efbc4f614b70ed9fc357b003eba4800c41d
z1a830c52caac4315302a3ca4a2808572959a66974bd9d8b34cb9440d1e444f19a6a3c71a477b1f
z810defb805d1e5791056a392a510413ab3f5c6d5b173d6fa3780d1bcbf8d918b562847f543b606
z3d0053d69f84bbf04d57e4023cc8781b9e718ce156cdd47d2585812d034f1abad589c691feb982
z00a083c6b15aaa169f1666448c4d93fbd2f53479386600d8d1b11c9d306b5e91a5113df51779ff
zeff464fd6cb5e27756ad6f949de8d2e2ded9650c416e9fbfd3e84ffb5ca8a1468bcc2590ec079b
z280dddcd0a0f5b2938f9953c6c5aabb3ee7d97e6a7925d497e63250c5b39cb5c6852cc228cf2c5
z42557f54a02f87c77a6372d1722f1cbd3871f749f454ea89e5c796ee1fc233c28b0c9f1ad1b9b6
zd6484842d960ee27537db218954506d42844095e5d1ed22c7f1135e2e4b2fc8e7d85ce0bebf942
z76a528826a1e28ebec0a5d73d6a3b7565e916ac2064a637256debdea818c2ceab0cdb56d84959d
zaefeb2e8a6c63725b5825c5e29e09439f389ec42676eaf344ecfa259fead79bb5c9b11c4b60d1c
zd6d3e86a52948dce97609c59ee6569c3126183e0dd2300999ab9a510fd15f13f6d9b8f7dcb53cb
z5143ae555c38de45acab1e1fba8b51bd2c526ff7d5de534729ed70928e64d44b62aedb5ab75fe3
z33d8f18bbbd9e979b60907d9165c25bfc78b15c99cda726a3bfb6bc58499367613d2273076c7f9
z843b04a24d85001d1655170d6741eb969969729e4e455f569f524f9954666377ea9bce711f4b14
z2b450fe0fdd55d318ea5e5399cfc92005228e36206c13861ac3f5605cd2a00bfb18c7657932c9c
z8f605b2437570b39e696ff86553704230ff3592e26e6271fbeaab18be74ca96ebf0251ac04a076
zeef90aee629e117696b7721be3cdec5a9097b6d18f610c48bb270c2a69eb56f62d765e68381e68
z950acb4a59c9852a07d7ad847496c61a9535100efe2af2e01a604ae523239a534f396bd9b44eea
zdd250f0684e90d6f59d8f96df1df85df3b37213ac5c1375d986da49c5bba79da283ac9b80a4b9d
zffe387f4580ff71431a2b0add9b4d94231aef13c05c256e38cb7dbe7831765809644c89304073a
z8da8a03ae081db8cbd7f5e9a809a23336327914859c0579722627e3f5acabac68d4297082cdb8f
z82144f60ce19254f84d815e3abfd94be2c71d2245a2daf61a7935093445cc0a23d1b90575ef0e2
zcc1827721d69698a90c004d6e01baeb0db31bd52d0861760bba7e1660f5d8f61999333e041ee74
z774d63aa17a95bb6912c9b175c6a7f0ed80d6bb3c3674bada41666e505460238ecea40f1399d2b
za7e4fc19b811136d7a99f401b793f16c4e37255480d831f0363d08802b0ea6f46dcc41f87267b4
zb6e73acfab847590e31e67c7ca61f523f671ba518f57177da7998aeb18109de8bd044a7e16f2ca
z4b072f1b73377ffbf4024c2d47d7b68d27a4ff0e3475ad27b8cecaff778db6b7e851868aed9804
z3093087a4f2b2a4a2fa9989ad68dd666cf134957fd2507a5e838d3784d4418c521e3d174bdabe9
z9575676591040ff98cc120f7587b552dff5cc1343ad14da93a4a04fac2b5fab1596933ce321f45
ze3e010145061bce74d0a9a1ae532ff8c758f62e2bab9aaaa89a4d9b76aa61abe55ba9fcb46d1de
z32b709fdd7be49fc115fac3efa87815b07f03ffbf731f3913e1add2baf08d245725552acb05e37
za6a90b45e7e1fac966dbac8651da706d50bad6427c93b710a64389efd0c6dcb4318e7984ec64b2
z5e204e432b94ff994a5a259ce554b104da97432b5fd27753a812598ded5a406c1a1495b5aae3f5
z39ce8769dd86165d5cd60f3b8acf2592d55a3eb4ff7121014e5749b6291b14a1ab4d1f430d4ae3
z11201b15ef095df63cdc25258a6c5e1cc9dd50c3c51e60b0442357286dcb1e299f3efaa041f0f9
z9fae734cfc9191289e61b2c7e5b7990fff8bc1056e6c04b6e93db5c78b0b495bfd913051af54d7
z297fa02a8d55c0071f787f6c72b1f0cdac6678df2cb5e3498082068d106abab437ca80c26c4cf9
z9bf85ec8c83a1f34aab723ec8725c8557d46e5846a4a7306be4ba879229be73a1b84393f58e599
z381b6aa73da99c0b014f20f74c4b5075eb1932c1f7621f1aba4792a535a613f351636c6b8f4e4b
z3b9a702bbc4c738ddd524a5833c3ed7954a83d0fc1f37fb00c688a3d23164ee44f77423ab14c3e
zf17710013ed2cff644032ac72191960bd7bcbedd83343caff8830adf96cab2d85760ebe9199fee
zccbb311d17f953d2b8071ce7c20c5d04de2dd228fd8ecc5bc74325ab4317bb23f75b7269ac3dec
zf7d1e0f5c09028089ed4a5499f8d416f1c2fff4d6df5541147a1ab524cad986ea453dc32179155
z71c702d916f4d06a052fb49c32a74a3a558dd53a9e45460f8f703163bb8cc22d32cdd71dbf1a3e
zbc319c9edb40e5c100845393587b096787a56095ef7c6910799ecf2476a07f32b0a5ade421eff6
z288fc994567dc2bbe0f798beeec3733ea2155c987ed5fec30e77835efb5d06b12f9ff4f9af3d17
z4be62ec7a5ea96896eb4543c6ca88039ca3551f039be5229cda15a06bd39f6d44c353633828cd1
zb209713f38d0b4f03528db98a4584b735536e208fa8d39c9a4755f1024a9695f01a3e94a0313f6
zce908098dca14b3ffdd942504cdc637cf17cf6a00f3621050552537ca9a53a749e6767afe25a2e
z224bae6ba81ab13f4e1a8df33332f35216bf65fa5c1cdabfaece07f03fd3368b30eb080158cf43
z6a3cc282c147cb2e12ed1028aee33de404b1ad94749f166d88d78c743d27dfb0860134213ac698
zad92fa074cf28718631d9b5ba9dd5cf78261e08a3eafc091dee0f53eaeb6f95d88cd0514cd88d6
zca4c9e355140db909f1029d72cebd5c3610af4978c6987f71cd32eeed1017bc9e06e3622a7b6f7
z79b7f1a590a7aed453e8c1b9bfe019f2e7d3116a970d6e32a5b8f64cbe6ee04457c0dd55846cb5
z2a80cab573ff0a09214fe200685b351035aa30f6fb9b00725accd89a899cdca46a81e2f37d0f27
zbdb017f5cb9ce13ae52fe3de0c7d6c1e9cac28fbc4069624c243056ea1425ad970df01269ba4d5
z013750c0c066a845602dcf611b298edc3a231123c7a2b09dccac544ff44d1001767d93b588e1b0
za60b6bb500f58f4db4d593bcf4ded379ee88b4a6535a7989701f06c2da2c1c26dedec4db31b4ca
z84e2fc0cea6e35e4e946d2725b0cb110a3906ec88448d127d35e651fce2a216456f6346e3b33ff
z15f60f78c4a736d55420b2b4af965f024e042400e0d077888576378de77288db38a897f7d5483c
zcbfd3ddf686f63f67a453c725a09e40eff3a672625d12f6ec4c914e87eb891de11520ec0344fc3
z398272c203a47e36143f34f72800ccf48dad15fc7d653e819b5baa9b5e7cf3c10739478c0c9712
z208aca16caccea6a905c0bbd3332ef5f893b1e987e829b2859fcc9d41117bac3caec952d02dc48
z7e7211a4f162d714d2ef98c4f5c77f2140308139d9d53fec415850148b3c46722066a71ffe0a10
z4ff903fc4a0af837d1f1384dcfb80f7846d196c8dbcbdcddab70800c8ff05ac7d08a31c3ff511e
zf31a828c26dc7c12b9619b33e09cca83afa0a9e1663c3f085a21d3e1bb8940cee732c16efc8c37
z9712f676e3af7f42c7b04b9d2ceafc576bb781494e9e083618252b05d96fc3ad59fb7cf187b819
ze96624d3415b4fcfa4ed57d0f838db655700da2fc6fe2a4496e1466a2b83b669491122d80a4bf4
zbc3661d99d80c6f49d2132b1c244d817e890852aeb393c739a6246e35701b1af9a6e66ed8bdbcc
z01a0eba351b5e10679d799478982741bd58bb73494a8bce4f5d1280347f6000f46cbf73f9a9ffc
zfa2ca3b442d56ca38b4e77eb452ed51cafb6c296ecc6b1cf2a0fa86be1ba1f8026f3d7ba1ed23d
z6a70cced3d469a87646f46484622041c3f091fdf93f6db0b31ee300d0ab633a03272cd456fb8a2
z581eaf5c16964e6a8816b3a55dfecf68477bdc253c266640bad0fe79a39d62d21b39b36173e22e
zf464de95c47f2a0f967755551808030b1cee65bdd1878d55c9d076488224e9d279611dca0ae69e
z5bb5e5536083eb86e227b8572c4e6cd28b6796f1b221a5d4a20ca8903d7cf8e364c8ae26e47756
z0cbb9bb3574d922486a42a2d1e67c985f815523ad629efc04163b919a2bd7fa0024f8bbef6b970
z3111c069ae70cf6a7a9139c3fed8e2a3d7827b3a49dfade4bc23d20a1685300c5cf0616d6aaaff
zf302e02d6c9e6c4ee4b37341531b7aa10a683d5cd39e794cd764809b8de3fcaaacb9851964c96b
za3b1b0572cca1e8e3e5286d37ed08640de94dc3201ede1e6e228e3f4bb64313de0bf0aa2cf9452
z725c8ec9e49a3ec638de8fbc66101035bb11eed9305792ed01c311732671eb202fd7486690026a
z55fbdbab43c656c82b08a4de7bfe5ed2d2cc3fbaa013ed5458a3e8249d7d7336efb5a76d459e3e
z25fd248cb9c75bcb3c4bcba509ee637cb88b5d7fe123f2102886919ff696968a7cd9e27fa598b5
z68c8e0d699bafb5b52258ab5deb1654cd3ab2543a1db00e18849435929781be8717a3d848226a3
z572a4743a3dd1538e4f5821f4b8f79b550611ffdc9c435c90e8450a47debbf578cc14cc57f0a3b
z01458c9298d6341ffcc259a852444bc95e4fae2e1d3ad63fa4a286cd88538768f140b9dc7d5b9e
z624ac49be4f52b6962b78d211e78fbe3593861ec7aae6638947a7f29d68e45e8bd49f2bd31d4ff
z96c3de8d803a1f2aaf164404664d789a18dd5cdec2efdee3ee3ea74fed3b7236f59c9408ec01ab
z06b88e357a560befb6e1ebeca6bb1f7f3618b6bca5781f678b9504809764fd14727bb00c0e4acb
z57c64c86a8dcdccdaca4d425670a92c3eeaf6a3c8df637e842070285f26e363c751512d63c742e
zf989bf135425596f7caea4bed37f6c276c2b0e491360af39c8e7d8029735a0cefeff24f4668499
ze691609c5616fcc73f6becfe887da6a8de080999de6888ad45dddb95bedaefb07c9f2e6d4aec59
zfcfdfbd9db2c58bc5a8a08808309af98e7ce7c3e77bead954450ab06855477caeaa73e7aa2dd8e
z8675c0fc2d35b96116b10cd26f7040f4eb9c715bec964ef78645e1303353bb687ab733d92c9408
z02da65a2e003411472ef0a11b6acdba1a05a8eda3b11923312394c4298dc504ef97bac1950ee36
zfbfae1cc141aaf236eb76ec206732eecab8a7b9c52f6b9db1d3997a2a665e035f84a328807517c
zb8ef5ef148f977db33189febbf15d03ebc0b5dea1f85662805e33e1e8e6fb1517e0f59dae938e2
z110535e2eca7756902d32615a75c27cee2b2ef58eb89c55843b488996a7308a0a2320bddb62829
ze51f9c978fa3fc51d1635f89d71459d519a89d51ac3a129005df9001f5dbc64908662e030ba264
z0e7e554c7d7a3bbb76e873f72b2051364debd1d5c578a84ecc2f05dbf7c24e031b18340a0c2f2f
zbcf9e9f98045eff53139dc72a7d2fd3bcf7e9dd1f46e1fc6978a8f58128e05647a8830a8570075
zf5bf2c7624dc1e991357d81096014f020e4dc84d26b91408d1bbdb5affa3b903646707a95e19a4
zaf3949004ff5be55b5742679900b8240ad52f1dc8e14215114a82e74bb2b8b3433e307272c80f9
z1195639db694c6553f9f65beed10fc118e329ac3776facfaef8c8ca083e1a17f81ea08942940ff
z590339ee173f22795121c135b2c8ff369e279aa0a63c7ce9018796528d1798000c95334a7f0312
z6274f1cef7baf22de148d87253a1b9a44d10ade114c4b1184d4dd49262b26d1f3521683c9fe1e5
ze5e912ad08f20e036a81e225f66843498dcf84c2f3a568b37faf24f6f0663ede2c583bf3760959
zb3467471093e776b29ad7fcfe5caa8b5b86f00e0300e2c83b02954bf340b05fb804e8317996cd3
z8005ad153557ea4426cf39e369d8e8e850c9639f1e6e81f41d7c811380f8027e7c74b0a37fa866
z5f3630609af6cc6c30f0ab2faf23bd05d7cf63dc2ebed632c7910ee980edd5fdb7263ce49bacd3
za6ddb2e8b69c5eff4e1820878977d47068cc9fc6eede211cfe9e837f3779a5f624aa610d97c3a0
z0067532bd15bce26b3cb58a89ca923abd28415d53ec9a79cf61f6f7a6ad0a14cb9e12906f3985b
z59e8f9817cf403d90f09334c5b3e1d6d349276207862a4dfef65e03d46d3c4cbc33542c1a0b486
zf67502106be5ddf624f13a355ed55221185860876750e57b8ade11425e530dcc50b61d36559bb0
zcd7abae02594b09a05e9633820a8f5493b08ae91ab4a344d23ee8073ddafc3f540d7f0ccbafd21
zffd0a22cdf7741aa160f50d9d0231d10bc2ec2dfe47e4b63ea187b1093e29cc5b3d53f7fff271f
ze7036de552d75021c3a105008d188d150e611dc20c6d72e02298d5ca717c4fb4c8d5294c0e3dc4
zef60509cd0e28d0bc0dd5087cdb62d236f85cdb7a569bbfbc47afb65e598f3d4db544650780c04
z753fa9a2918e20d8377da16b36362580a593e53bdebb82c7930a6800dba6818c73158874575f09
zc32ad419353d9826098c9c58f97e4a1ad6dfd5d18d117e2e110b6c09fbf2253713e78efcb5df96
zfb60089f060806b2e75e4325bb53210a074f5bba878359c407cead9c50895ce7918f1fca0118b1
zb36df19834bd1792d61677d28647e653b80106fb4e77da1e038d01c5264e6050c791a6bdcf9e6d
z9eb92261e8f1fcaf66c92b3197e3b8a6f52856162938ea806cfd60acc2a570a7c7c5b107f974ab
za767fb7ece94e575a6eeac4bbee6a26357207bed18ecb98d994ebbadb72baa0a3390598de179ac
z079d4f824ef5f8230ecc48838dde70b3aeb24aa7f807f9bc46375b90c5db4f1d3114a3ae0c047c
z09fc8a567c2f45e7230c44d860fd9fffd55163fc2b1f783a3ea4d2031092659cb929df2fa427ca
z41d5c549978c48aeaaca6311c28364c56d52eb34239e254e141529ba93004c9dd29cedb070cfad
z8332311062f8606ccc70c334eb68a29534e885b91702e662b916f929a91b21969edc4fedb041bd
z73d5cb0d3bf9341bfefcc5ce25dbb10f25ce1b21ea544cd98643351326fbd93d0e49edd5078358
zc9912004fcf5499b57e6cc29cb83467f14941805ceaeae68760edf0cc386d4ae3176923b861506
z6ca89f8e477cbed0b89fdf640726604cd0063da505202ba32a0d78960ae926190399bba73dbf48
zae3cbada3ad7451763444cd454cb430c751e88a8641f93f1599278415644a3b4464443b5878966
zbdc1cabe745885e1c2df28dac18dd6517f4bbce4efcd1f49427fa29dd9dca80a81ca0b9e2c5775
zdc07f70960478db2ef487a96c34831503e7fc703b2c81da877e66d6b4fb9f0c36dc03f3b8bde6a
z836540bf2aad6d0cc984789a041050f879c494d334aa1d1ceed98b316b71d41079ee135d29c260
z3b1025561fe7ef8418a76380f280b3cbcc649cbb60955663ed59e7a978c8510e7db5e7a1a10a48
zf0fb678774fa00905a52413b3f068abab905e80c859ee42651840e44c520cfbf2333786806a8b7
zd57b5a65d980ffd24f368c1a55e1a6cf0afc297ff30ee55f502c2aa138ffa3374b3e2b80c54399
z2ba1f2c60ae5feb5f492a0852035e11e602cc8cc0596008fbd983ab79eeced71994e1ecb62b580
z7aaec90584293e79d95b1d79d4f646089a3d18c4bb1a43ef556ba425c26f9405c64c139217f7d7
z13f526430139835d6e739d0154a51a3fd72f7018e3603853ddb8531993b43823b330b5db4a0e6a
zfaf87c34d9be79394f847f3994f09b6baea6db215233d9a827fe89f48344bef74e9761979c6b48
ze05b82a1fc450264f71b6876300d5a9a5b08f78e86a1c3a7c22f8a47800eb669fd6e2b71a3b871
zd54394ca7b324ad88603607fa881a464e4aeb82e7e65921f62248c975f51721f94d2c0c33d4dd2
zc05cc961182d96b3e4bfdb22e91af908f8c6a5b3aeca8d3c069f6357c8a0b44859b66f1025ab75
z6fca8e8fb045be00208f5fa6b3e080abe4a7addd2987746a8a8a4b09edaa575236bf3c6ff14071
zba45d1b253bb962888f163c65d1498ed36365d65f4363592c5487d42208a7580fbdbdefe75b9a3
z03ddba3c697140a4bbb03b4d30fd148ef04b2f80171ac66a46f9adaa2ac805a2299c2b65247bfc
z6f6b88865d1b9d10aab744e5a18981c7a6b3e86c3aa9d780a0290fd0c606e334fe53ccc08cbb05
z44e0f625171e2eda9059c53a7ab70baeebc6b0baf57ef6d98d7db759d29fc901a9f1cb56680994
zdc95d68bafb45fb2f648ab6c7fb22e375e2a4c93708a2081642d3d45dfac2188ef75440a197950
z4534a7fa85dc5e1fcb6bd1df605835dc95eeac52d9e878d5c1c1f6fb33304fe9258ae5fe98edc4
z514b8c4fffa28e9958e1ea2134570210160c291c6f6c996392230997e2ed51258241c4721e54df
zc1dde90970027f8d6afa6834e46601420127f78e1363a0ce9e591a20fcb5941efb9fa723bba9ff
ze4416da546781d5a60f1005b51db511ba5eded51dac9392fdb5c644b2ebf4bd3aa3dfc8565c160
z8bc0e8642453ab880d74a0bd22d5dcff15ee212ce00120d7f1f9faa166b4e4f8be83bbc40ff0c5
z11e680603d8a4f069a0b7fb8093dd654a9e53ba648414764d2309d3169f5bbcb0d32bd1d6eea00
z076da6f62536f876f247ce9cecd0d86227e6dc1a80562f11726507e93f3d0f93f80124f89187c9
z4e660a91f78977ab272ad337d224fdf3f99b6373bb1eb922d492aa82337e200def2a6a4067f3af
za4a2d58b908f35019872ea4272004ddf13b7c71522d3cf9fa32c2b956ea55e4ad7edb376cd92e8
ze8daf16430e34632a76c2a74f084c6bdc984dbf20d921389829786a26df65436b96670acf7c132
zbc34cda34e406091f5c02f1dd6e9bf2f46b7075495f59280722fe66a4670ea2cd2237238860b18
z45037e8d8db805646c12db1413ad237bacd2b3541ef3501934ebc868dcd1b072ffa54fb3e67883
z066faeaf5e4333398dbc7ab6229e1a0be760250f43891ffe9541e8f5016f15c9cdbd57b7bdb524
z58b51a56875ec7e7332266c4776355195e903aa6d6a3d707ae60d79f2d53112aedbbad4dd7a508
z12e9621c7382aa112675a59bbcae2ad15ad63ec2ed176c4dfe1527c10360dc321fcc4c1a2df602
zc6f6f56626e19657a73142d34e57f4a8a6b9d02089195c9c9ee36d3a3eff6d8a93222d322ccc45
zc4b1c7b3bab711a6c894a25cbfea8a7fda835584cff4da9d08c4232973e0ccb140691f350bb678
zb330b4926948f383ce7a3cf3bfeae384e816ecf640ceb73233bb61dcd069e2783b754b4b94d5e0
z8f87e8c6cd88d4bd61b01d27b45f2fb734be866b06ca78b86ab2d6c4846335365743cdfe75740b
za17de926469ba07c7b21837f27e8ffd84eabfbac184d1d182ec546186bd4fe835edf84c35a2133
z4781b0e48a2dc36041cf6d30177377d1bd423563502f5c09f43ebfa2f2cd0451f942f6daf52227
z63a8fbd13180c6626cad7ea805c67a8dbfd7792799d3e3d4162cea2b271b69b3f5cef65997e34e
z4b3f8ee6e3c2256c4a282737ef04c6f9a858c5898bcba66c27172b483abed42192e0bc2eb2b493
zf6444b7efe2a6fd57571fba50c71b0eb4a1166a189c27154e7b3d5dc206cdbe8990937f5f6c00a
zb0e52feaf5e5989829a872e91a8aefe6f0d2dc6b133f4a073b4b4134c6e2018ac1856a0e455d58
zcd5210f93ffab9fa1d405c83a291526251b1eeaa1b19f65cae940cee8d111a28511e6aafbe61e9
z8dac3be92affb842fe823e7baadf5342666c2db67b86dfb971bfde4b1d54be478b63d750d85b51
z7cc9498489c19baf571811cb7e1c963fa3b56aff44e5615ff4f7d7b634c7c6b4f919c95f72ae6a
z478db5838472dbf5be0a96ce6da5c6db6c96f9e5d8a857be2cb45c8b9fe21d23f05e21d39b1121
zce4b2eb715c62d0809e206cb61fc6876a7bb8f4a32d03f377094e744101d2dcfadfd91be0b890f
z270e75f9deb0298578f8b5bfbd9ab2f66314c527908df3aa34f5c7350b5771147ece99c50b883d
za74b23b10b0e01f4a038f4a9eee885749fd62e2e866fe7c9e36cff7beb8b8a46e6935e5bb5deda
z78d168313025d88301a553c3549486bc41bac758398c52caab654eb409ee66018da53afd28eed5
ze7ae1d5986147bd0fa7938f878908c1a316879e0d401d61041ec23d18d83d8042cd7d8d23dd170
z581904f6cceb2d72e3cc5bb476001616e1271c7a8ad79e8016b9e60928ff61912b959b5ba4a252
zeaf01a59992baa4c8512c437084cf9c34be9c9b4e2eadb89a651a04a390da9c573a434e8a7c3cb
z25c33aa757271f46e9f8f7498e05c7eb39b3d30d365e2e171f82cd2acef594230bb0e482877a1b
zfd61010baa025ae6a99eb45ef3be718b1332bbc0b55a6e02344d125f834993ad7450b30c83800d
zbd2073f7767cde2bcc1403d5e5d2b7a49ae7f535c4506a593e08c48f98a77f8f49b4b115dfda53
z17d99544409dbc4585cd6848534ff3b1d25a472417533c77747f02fb93f899d007b6b8b68e0ee0
z18780dfaad9c6a25caf06821f89c7f8e823e7ea494845febd009cbdf1582066b53c85f75442e73
zc57f02bd62f8260543ab2daee48b608791da3873e3dccb2173f4c6facfa57432fb0ed72559c617
z8f02fe92cc30c4091187d72fe3031e2a35c7a26879a28000a70d0805fb0839c5b20ef439532a08
zb7e4c4252c297d633bed897f48f7ea5fafd270699279361f6f11c7953fa142b640e1f42cb7b63f
z0763c85287abb6dc111b9206598b3bbb19b0601ed5267b7892572bbd3374ca7b596d3c85f7ef2f
zf927cea7b58978d5727dff082a82535b054ae0f32ef1dcceed570625e3ec70708b853bcb9db941
za2e1db9f9f55fd4868e25af31f293b93d0029a45436fafd5e0ada324ab221d50d1c04ed8e97590
z8ea9bb34640dc8d9f15135e2c638dc2f13c74180aa867b710b9c54cd75460d9b0905e3af1d097e
z8bfcc9925cc5c5ed4e3ea7034c584633313c2bcaf1dd0f52464559e853fb756429d33c7037eaeb
za70c0e4e8375bae0874a69580438329ea5b1f5243a905d3910d80f746d91178c0ee2d4e51d1431
z3786f1852237b28ceae272468c780528c91622a0e9cfe2e1377dd7fd8d0ea9b20e1d1220f26ccb
zc5aa9893c66b04d0860d633f0cf89bbb43c04f4a511004709ec1158872e41647ae7e4e04ccc3f5
z65530472d55b202a78ce21a7608a94e6a77deefa5a32f8289338e31c3dd36eecb6af8e4c5a54fd
zf6e11139fb5a9b0ee0cf97ef67c024838e90706f63bacf9bb463c2d240bb571794b53d21108fa7
za97762e1328cdf9c05ff592ae728d924937135da43f4e9108736043aaae8c710d8d4c3d3e503ee
zbca58bd18dd0be041cccd5c732bddec6539b919a2d3b4afa8c242a329e8d6ed8e055ae9480610f
z79bcf1aabc265a258a9acc71848879bc995f5ba37232391c6cf54f2ea285932ad658c252cb8ede
z763a5cde8ad9337fc2c837ed24f5ab68d91237efde386a8dca07c92776334c16e54eec036c3c8f
z8f8c0787dda3812ea10bfa76ff229e5bbc63d3b7d55f9fe0943bcf800c344002c6102aae2ccec7
z4adcb36c0b1a520fe9ef71a49a3894a17f95d78c8d46277a7cf62c05c72d2a8eaf5dc80f552ae8
z6089d6ea077a9bbf275db6bd8ce6783a4427ade562dec608f857a8fbeaca32ebca919532f0948f
z592b4b815aead3c66cbe3d736290836bd491e4db5b84e24bf652dfae1eb4f26e58c12ca044aee8
zccde2046729bacea49dfc33e4826f92b08e6ff9be04061095939fd2fc83829cabbd6a809586b73
z5389c9bbaddc19a710233863af52fb5b95badb86670297a90b2dc17ce46d1b4d39fa7ffa36eb5d
zf936e81c70a291095b66fd1408bf6f0f31da8334215a7664be0314596c098b2b48966121d23cff
z44a0484285cdbc2a6628ee8408e5702261fb6223435e0ec40b66847850cd1246aa6bf1f7cbf55e
zdb709f6409ac8e895de11c27bcf07dd99e295622255db00a49d908ba2163cb7bb57ffa31bf06f7
z27fc9ab328aa0b002b21c698339fc3f78d7a7732f1a00afa6d10c521dcb59f7d94e627edfbb74c
z05cc1909bff42cfc3f52e5b4f2ddd5871c5baa8394b73a658f1d77539aa6880e62d0e125ad4698
z34cf77f1a36ea4163c0817f129fc30707c2f59051ac0dfeec68840f7825f7a21fc8c0836daea39
z664e9adc69ff8fe8d55c2887dbef7aa4a8f453ecf4bccc8bc616ef70104982c4d6e8c27cd0ca4e
zc7c7d4b7137724cda200ce5aec54f252ba5406683c13968b81cd22b2459bb0d81253c27c4c8e73
z59b40ba967918518d5a4b2495533b1caea195caef9cec426516123ce711bb3aecf343f74d1096d
zae9292d1ff0895d06243ab8661a43e2c0c69f63feb70818a4ce1f601bd0a7e17ffd9303f465169
z0afa5f49e990f087533bf8289d95487dc84906c85cd996c15ebe8ec5ab86d69510e35c0ae1da8e
zefa9b1f071983fcef0f934de0eb46a4e2d4f907f24bb5f6ef8f2a47196088287cb0280abbf976f
z0315f6582b5c648e5556f8fbd769711ede27485c22d1eaf0c238154c460ba5940d53f4399902aa
zb91ce62df531155b434666b14f1eb63dee605fc7799fc8db5de009e4ca657f474d1cd09144c787
z732381895c534a2b72c91cb1086c0364f337b9a389b59a7898f8ba2a09886ae4cedd97c54b347e
z488f08ab9c72f40fbf3d1e5fd8b7502a952a4e6c4a2d67c04879abf56446fb39b4c474dcc64ca7
zc0fefc76dbb41acf81d8a37308a503e09cd858d442a247c45c6198cbdb864a34119fea92620ccf
zeebeb27f814895ce4f72ca309e1c5174a865dae62001d9487b38a464ac99afbc6b453237bbbddb
z28e2305b16e843e3d9a9fc0d5f036df303f6e941b4039a41e43871dd13219c3108feb8e96aab54
zecdf424250ac9f2b9ec381722df2a5540cd16172dcf6d05fc0a52fafbd19edabeba430818dcc9b
z59e907f9ea3c4bcefdbf7fb52b503ae342f26da38bfd698c9d65d5c00a31a9225fb20563c0a69f
z494f580dda5b5b36ffeed780ea9844d6933cb6e57b1490da8a28d97cd08ba6449485f06cad870e
z5d5fe88e7b46365974ae174ccacc4cfd72caecf5e21114daa8f6d7ca22f8816cd5817b67d5b01f
zcb72de290ed4efa05de519bb5f0c257691f9d718d5a86112cefd895b771fa5e30d13dfaaec0297
z3d11dd165aa4e9e03178a6f23fff7f68028143d613101b80ad1d13c15eac16cbab1e2eb9105c88
z54849c49a4b7a0382ec3c1f28d04e5c5bde63c344fed73a200924598cb23427146a5e8c4574fda
z2b9da1dadadd1697c49e0027f618d9deccc9706f7f7dd4f7b0647f616eb30767c5e5260d679614
zc668c216c562be72514b3b5442896a6723c6c01bb7643a43c2e507dd3e68a8ddfb5b74055d6d7d
za981343632e0f532ed0603c3da36c49b4a44e7e1b91e2038371f3e8efd4bf0df9847aa63630c69
zdc204eca0bf83331da8bfec323b4d06875069a3336761a8ffe6ccbc91505070e9fbbf3b5b472cc
zcc655aa1a838288d4b9be5e21e9d9fcd759dfa2a6e842b11c4953b7058b8a8ca5ccf02bc76341b
z1ccfce77b6f39eed35a33ba5c1897f403de2bc6aa7a0bac521f863ba805700ff46fe7a846f3ddd
zd1db6b0314e8042f42e733820519716a0f6dce2125e3b3a702ed7f82d54100e596c9cefffe1fd7
zc8ecb5745c3832696eee5ef578e7809844c8188d0b0981cdad9e23eb1de1ffa6584b1e325a6d94
z27e6ccda35e4f3e978a4863c844a0ad95b20b54ace286703574d6bff4e1a7b96a88809ab3c3b2f
zd25c6bc5eed62f34e11a16fdae45c2935ae8acdb07614ffdbeccb6a93282ab5d8414e24176327d
z7cd6d0029a880f1a58fcde904e5f34a7346e532be63ea8b6400a3179a4b85e61090e95a433f6e6
za63361dd24fed17477067c0c83a699a296a1c6fc7db9e5abdf0a399763867cfbf5ff8f7f603a02
z72d4d7894eee3ef0f8cda2350c9840a5ac4b3bb86a6d7a34d2b091383b4bf1d3ec901ec12cf0bb
z34c26184db4723ce0529106997b9f052d89de371fc0223ae3f0dfdaf773d795dd296cf99aec40b
z3de4a4d781fb7737216db6cd60fd6cf0de5a3bbffe88f8d3fee26803048e7cf1cc9abb505e1e6b
z12d91ff23d166494ac826e9791638f43c7750a07125594c5c66b6728b67888956c34d9623c9b40
z8aead015095d743ff7a36cb25fc155eb0f0579d056e939a1be8f053ffba3b4d2fb198f1e465d65
ze85a0413d8b8ad63d939cc64c0834bce80117ad1f6a8132ba41d16d4740bdf9a68e45639b78b38
z048653f0abd0d369a78e08308f5d3e8611255756fcc981532df24dbea77878665ec2c5720616da
za0670ca4bf9f4d01e9e4b6d6c0d355f79756df73ccb1502e002c74c55b64d4dcbcb46f276c33ee
zff3bd935b3aa3d95038a8ceaf2fd1bf2dd2eb78a7a413db183c82ceca12824c27ae98fc25e2f2b
z1b18a2fc42cda20401dd55e66c0b154b8c8fc15cc6f0e0e40503bd8d13bda5fd97a60126999cd7
z12af1f18833c2b776ca2b8fd8943edf79a8df8fd2952e6ae6dbc4eec2b6bc31a004ed301503f01
zfd4efd4d2c6e1d97678e29aad0d0ee7ebab6924bfc9b809829116c6d42eaae31cb698aa2918c5a
z286f5f1d4450436a909f4501b4c63042fa421fca20660bf8e7c2a7da04de3d1b74ea9aceb236be
zb6a52643a16f188842d8f52f11c4cbc12e171a73a3fa91a566553808506bea32cabf523a3be066
z711da229bab761fdda475448f3ccc7a8df3536b11a3375a24499caf86f464ce64c915eaa0abfc0
zffaacd5fbd91705ed77300a58823223a1769f758f7001ab56e57ddcea7e1ce2f0dc81100f5cb44
z400b02646c04c416e1cb1263bad489b57ff71597b6f876fd6acb71704e85ce09e730f3475f6768
z36db862a6866a62e90a78b66504ffe5e1ffba11d4c83c1e8b1c58a7fe9e5c80c77e3ab01c8644f
z7a39b415560bb7adbe4a7c492b610164bb251bbbeca8509cebd122eb22224a288df08a51e4caea
z959042ec23011794bd795ccafba2816b6f7fcc495f6388282ffef17d613fa1a139cdb25e60d106
z73b0ccd08b4eb9e21fd7bcc7aa22eab6f6be1639b383bab4562fe31ff8be61c81a4dbfd60a0049
z223c70a3abcf725120d88a52d2ab235766f182a5ce2402da8a50fdf1dcdbb2e872a71223bcfe87
zb7d1ed644d3dc8b1b1aa0a64493ee92a7427c3ca1230c85798cc46a5950334fede77b893888774
z70339d560759a46324ead49cc3168e45f6a02fd81956f103b7a0d090c48fc32cacadfc475b0cc6
z97c7c2b55ac3a3d2f6b11b513bc7bf1f6d1c152cb5c12cfb3a977f04e9edaf278ac5481b2d7f6a
zf9116523a3db64e43fa35a0e2c2a4fd63112fee70fc46ac255dda59b1ee856840d866b45302f12
zb7e12fd38fd026620a75ac7097724d7b6c36528626aefcd781970d84a1b287e686032c69a9096b
z2e04e92d39983790c9ef5c812776633b5d680336966f9ff2f0cea119a295e09420479cc0e50248
z9f1cc658fc998865888161ce883bd75836aa1a5e77bedec465e00320800a4d0699d2acfd76e300
z1d6b23150c5366ccabb8c145d982ba040e01bd1499ccc60939a5c9dd2b55ac7056bc6c342c8ca4
zbd60e7c6081fb007d2ab3f1aa3e5d90f66b0885ae4368071e53ee59c53dfe812207d1740ee2ad7
zd934f99ac410aeb95ada5c8db11a95c38299d037acbaf01b318790be984287913a624d9ebbd110
z7d5fbbe9e1179306a69f10d6aeb896cd72426f3ac3de9c4fc9fc71c80a0360e2a7f2a1f0c24797
z1d7aeb31d6ef97226e684835e2d5739727ae9ce44fa956cb55f23edd9d53ac5a6bfe2a25cc3397
z32477d39733126017081381490b0b4d422ad30f56858fd63805a2d3f613c9f013adcb673e4c591
z2f8aa0494dfdb3c818ffe3ee25a34322576ed7579134b68b1f921a45e641efd543a2b0dcb843e6
z411dfbd08158ee03ad11bc993b6f2107f2ee988ec6db395e5619baf5333a2b3cd3b4bc2657c0dd
z62d49cb7475f817a8ac962ca1cb4466ed09d207d43c2533df6ad671d8b9b268254b66ce5023dc6
z3ebbbea885bc42c12c2b19605db8a7153f63df8e24c4391455ad5b4a8881f0bcb0202d1bd7bdab
z8cec8158459f8ec3bcc84d067d0f5f44b67d71dfe298f319593e96cbb678e45c301e7585daad29
z33ff81317e724d38cf90f88f1cd6583bb9f53e928f94faad31b02d04700cc05286e583dcbebd96
z582182f91ed11411da698f5e02baf7195e3271654accda528fff146b196c99d3541aca3e1fd993
zb8b8a11a31f6c9eff212a34f2e245dd57f1559d4857c85b3d0797018cf6b6fd056fd56fa7e3327
zf61932040d76262ecb610624fc1d891651d0dcf2b3a5f72492d23a7416e38746462864838f5c7c
z0e34b67674b29a63d91867ccfc59797a7a99cbd361f1b064889fff60071010ff364497feb74bfe
zfca705c1f4023c940912273ab949fd2e9b7a0823ccc33ec5e37f9db29159ea436fff57d3d5cbdd
zbf81bc0ad9cd45aacad2bafe44504dc34225b15e425c162aa87684e20cdf27095c6222830f6bd5
zaff28134968fa55e8c363be18deadef7041d08e4fc7bf55a96ef6d1b30c0b6e07beb5c206f46b7
zfc10ea2ff248e9ac7815a7efe5b39c78431bcf27d3a2c5e79c105ebed86026f58a023f6c24f266
zd76dc384ae6bdcbddb933925aa0d55d12b264ac4d156fabafa8c53ac1d4a5f51cdbc7a4b3464f9
z82f558671e1554c254fdc7bbe851020865795c42717fb6870f6ca583ed964fdfb0c353141744e2
z33a5a993540536350a23d384703bfaf5971d872d1da944b63e2db2b73908e14b893b3356658ed6
z2471ce77606e06a4d33aa5aef7474e409d1d21dc38811530f85af1f375305fc38084f63022402a
zb2f676fe97f903faeca3b63a576e4331a0319c98ff1a6dcc61af0dc97fef41fae2a15736aa0e19
z013a2511281a6fbb41a28b1c779c430842ab54a32a6eda2b9ec9c33eecb800015d9a9a6a5b3a87
zee6c41b9f1133398e18e5f2ea8414829ddfc4e3d9d61db036cf76d71219201c2a3d8f04e787c71
za4a98ae7911e589967ad702c812af30c1e4d00eb83f4e9f0a847f7d0e3c8f8417060943fba5ba6
z9007eed36e9a680f08881e6fcb28577e47fe735958645f7b41305a05ca019804c431004a351b30
zfc1496c6a0828589efd9652c0086607a434538a02bda5773d9d0c38c2143dd4075a705ca4495c4
z3e099d93191e12fd576f8b0094d420bfad0841a71a56c63f190da5c10431d141ef0b54b4ec1c95
zceb43810077b5482ed418a9fb8f787522324d2e7fa9ec98920c05510ee3a2c4e7064c4ba62d2f9
z7b33c872e956890168e26c563d9b269ee18a89670fb5fd8c2fd5daec5dbe881d74f1ccf2477b91
zdc7f8d1010d0d7520945c07f253da50933d8f72304cd298eae765cefe2ab5d3fc0e621862dcd5b
z53f657b175335b7134c799c10f9976841fc47c090ab43b969c5baffa89e4954bfbccd55fddcfd1
zd813075a5cab8569df631a795202c8ceab70131746e8c93f71ba2d07c031f24fb475926924174c
zf4effcde8bb9bffd01cfd8867263937ac36e74c04fbbed7e82d9d6d1749bb842e340559eba5b6b
zc0289a60a3bd267455d92771475fc0936261dc24e22bf9567475b75c9f8c7509530207467af2f3
za102af442a7c7a609ef111b6ae6548848661b892cecce221a8a3a4adb302fd29ab04cf68024ded
z3e22f21d6406a3799934b409486c4bd991e197208878eaca16ae0f46d15b889a5888479ad74193
zf160be42d09e698d72896162c65841a73ea0eeaff80dcc7348e6fd376df6a290cec5df6e2cbfd0
za4d3cf7323e6f51b782306274bdcc1f95c9fe6d5125c444ef51f2b2e19483dbb1faab1b90d3a3f
z0e9f6055d930774c0fe597dcf8aefa82a9505810c0c6b9793048b951b6fd3cb1f7fc2243dcf237
z879f56e518a242ca3a9e393c02873bb337e41808e0262d87b9a8f177835c4425af47138b4649cd
zea955f019631d3f2b15bf35b214f36fd8bcb4dbccc41f80f9b742bc33ba56e2516af0c12cddb13
zeb4dc085a2e91d1f13013259e6e4606ef9b9e6d61362534dc55776221ddd38c0a9ef6b3137709f
z7e5328037e8888f13bbc62b40077c2db47afd463c0309bb2c83e00e1d37edfe5457fcc06c88ce3
z738bc014a7e9fe2fdc0003fc2a294af76c24df68b3291706a7d034db16524212b867553913a8a3
zeb621313cf78bef3436e37309d5fa36be4329ac41abaddada5aa75cad89f2003f1f44ec1acfbde
zc2d049672fe229acf3885b817a4cde7a3bf2130abf1aabcd9ce6ac0406b5efff0f166bafe511a0
z10e8afb9521bc317a3b995c0e6ebdf67ce600c965d39186d111dd05136859983b002ca7e66e2a5
z8db5260aa68504961b0854f4d093ffc9c20e9f34410c00ad49ebb075f78dc8fdd26bcba46275ef
ze581b61f822af01c2075b55978496ed6c3c543c422aae148a0cabaf0508d665b92032c1bc7a203
z2bd922c1d03acae5e5257d45bd4b93b3177880b05dd92710ea729e635a0206194c83c869f37359
z4d3b5adffcb37df877dc1bd6715f0a86073f182cf4ec55e33bf3116cc41f799069d456a54080b3
z99a40a7089bb0d34a0b3be978b4c2641db750cc2fe80225315ff36858c1bd651747c2d90490855
z130e55c687354bf200a9fcfe5c9826bf2c8a9e1bedd52c58cbf398bfd2258eee8f8bfa353ea103
z048d81dcbf862a3d9708c165ffd4e14e99558b4b82238dd89a5428e98b03eeb15685f67e613dc6
zfbf56765ae15378f6c563706793dd27011727bac43d2433ea7215833e97c19729687d9e59cbefd
z326c8a2f70be2dabf48d9fd32eeaffe04000c3373553399ad4479d3028e8d9ac3bfc123d1462cd
zff00ff6071f7709ca04de7914cc4dcf8bf76128514b260584d8c0c6118d7649d12f28c099467a2
z6f270930ac33cb0f68bb319f10b897f46759d86e3c9cbab3b734936bb80604385816a9396506a8
z547b6a81ec00c3122f5c4cb0ea2dd73a83569d2d33396494e2e7d1e168da8a427e94fcfb4c28b2
zb7afd0375e73961f2da1a2a500597614abe16370bc304c63fa4e27a0af6867ed9e38e9abd79fc1
z11e64d4ae3ec4c3762a5c690ab96454189b90c06a67af6b9bcab449a1d9a7d74dc2312b1acf998
z33bf241094ca0a699113cecf37ee77004e79eab3dbd8122d1e8fd540ed4569fc189322d945c8d2
z477790f4f189b1fb408f563b22aa43e9c8ec2bba0ac941ca3fb42d56310db9735b59550bacaa05
z51821c53d4967e66b9aef277359d81d1052d1646e866bc5891521e57e45806944a7f7db0fbde8a
zb85f3e929e1973278c4bfb92e7177e829412af194d615b54cabcfac372022908562c2d13fce2ce
z0a6c34c4ec28e3e9066f29b2f0d4bd4dc5d59adb51d08f4e774773892b708f480415ccd431bac2
z65b9f4dabd401367e0f67778b889b0080b2e4e16d285ff54df04102d2e4050d223da402ebabc67
z0b5a352a8ba19463e8402106fe8913372a7df96c1525dc7a2848156ab2c5d235bb5e6155d14665
z3aab41fc84645d2824459a4ebc13e89c73816de00511ebd170adba2016bd036e6994e15e5380d9
z4911b8c8bda3af904a50b028c889920be06989c7810b4cc63852457cebe32313cf11fd00fbf22d
zea4d3ad323a0e7c16f1c200ed9823f8718f52e26140e6402ee3eee6b3e85bf8fcbed6c712c44a7
z94873132979abb45e1cf02f436ecb5f4293c5f6e65956870e007ae32519113b5e554436acdaabe
zcb58172fecd2818713a31c2a81527a1db9736f2a0299d401eff2755f3025f9a8ef10b2dd1a48b7
z9260be9c14885c0d5cba11cebcdb2b25793d86135756b683bdf3e284a7f0139ebbe98bdc909ddb
ze2216aa1a3a2f291e0c6a3e2af4ff040ca2596633127ff67141da3b9ea1852654ccc7f018b85e4
z4218f1d9f0ffe039033f45f256fcce0445fde2e71c3badcdd4ade56f00cbff8ef3b91ce5d71e88
z1cc0280463de147547615b452b2132c393d38a923ec21eb9a11d82680c71438ef452059bacd89c
zbf4cc68759cc3bbc9386cee30e04d38cf3601759ba9e025ea7ec5025d98e46f3a3b5f9b36a6f57
z159ec38230af8c846f67525e939da5d58695b60f69b325d37357eac893e0a87a0fc6aba77013f4
ze2f38e9e9d8990a9d6f44893207fd8214aeca0d93ed04664de34238900ade1dcb0aa299909f1fe
z232d8c22ee33197635a4996f42d665a12086ecb858dd4bf63ad252ff8a51eefdde48bf2241ee14
z2b651aa54481b2cf6c03209e9e0ca2d6cc0877f97056922aa272985af4b61921648380e8cff755
z7322a2cae92d2328cd1f9ce9364a2af4c8a6093ebd9de6b8c0c9a787ce0fe444bbad4e4aec3650
z03e48e9b903856b6818d2d5ef5b8dc749d3b78ab64293349d8e8dfbb52c3171c891c8b8bcacc74
z5968cdacb471a45de06a34e329caf85b39fabd918fd7c86f55ff2ec55eba6160e7d5625aa9e53b
z8f539743a3f571af8b873c870d50b2b9c025497ac65baa9710bd3938accf9af8283e68f21e9413
z514c8da44f02f3d7ee1e6a9df64e17b7e2ac88274e787aa9e07d54cd4c354c117dba80ccc8d966
zb7a0f39fa55eafaa7e883cd3e8a9c4d1ac20a85d6eec0c595c999f66a0ab95f0671c1e4aff4404
z89529f719e5ab158ceba26db7828737879c114c67b512edd311eb6bbdd7bb7f60a7d70310f6517
z867f273766a751a60e8cb1f8ec7b4a8e4f69f6a680ef2e414135c395dfd1eac6f7644376237c4f
zecd20fcfe5ac7711f182b3f2f14b9b036224a32f778c5ed23fe866680345a34e4a13f5c310e976
z126a3a0338d7f03c94260ea67414efc3cebcd2f10f7eb8bea57a95018b2c53a53c5b881bbda799
z168891b7026b6c83f348e5285df9a6670373175b3c226a6e1f0bc6b510316000250681affc0b3d
z04606e6dc0cbad59baccf0ea3a4577ead099ef11194cf5691cc29cd7e104cfaf24a2d39e35a485
zb995760c616b3f6b810be69fdb6963c208b18477a059736ef862f357f5266f24110425699e7e00
z8644c4c64abe2433e8ee2d694de33ab64c25c941f3f9938f5a160d7d9d02928c95d58cee485790
ze99acbd028c0ddbeda1ad13e22346ab9753ac1bd088319941cd2f402d6dbe2ad60f9222172bb54
z905c6500170104a93e6d9afe9d4897f5b5ad39840e0da1bb7ef496d3dc144473289716173b4811
z219a493b09a155226d03df8d05e446ffb5e977f21a5f633e0789b4287e0f09a8fe7ad444411384
zef3bc4c492ca1089e1f48d0e2dada95347f44e25eb6ee47730f1c22b7b7cfdb0032960aff86531
z2919588b748d5ed41739cab41baa3158b2d362fa6c06ba80afbf154369ccbd5ba285450ae88704
z1210688b35145e20f78651daa56e2bc7be5f76e8b591f231075413ed656b5a078b587eedd3b3fe
zd6fde0da33ea9dfef52e0b7f44ed6fdc68a3788d0484c179f13c38a020ebb20170a7ddacfb9c59
z7a7f53964eb593039a1b676bf8124f8f5ac07dc88f6a33c1ea7742e3a9edbe64ae3045bf571dd9
z7fd8de4662cc2560876cac341aed39906180bb6f18cb3292cfda675bb55b1b11d85d38b2f2987e
z24c757b72f5ee8fa73b03d566a04ea5492c7c25fc8eb7c053a0aff892fc6be0c1537bf6aed65c6
z5104501733cd83dc4c9fc53da086a43b30c7d53bef9cae1421b3fbb36dc9d4fa99d68b093c9b46
z236b956b6f212b1f0a5397db330b191162d21665de6430513b69cc7ab0895fafb80f236adee54b
zf491acaccba79dfeed0ed488be7e68591181c17f56a96dd672b5107832154bcf83da67fbfb1b66
za6b694c50a9d46dca465c5af3374f5da4b3cc74201725775cdedf485197fe374aa903d21226957
z712ef71c36893e83887ed85cd53309c36321fe6f5271c6aff895a75b171ee8301a91127a2ffa65
z99bca22ce03a94dee52cfc8defa51c6e09f99f83d2cdc57b96870d98741440fa70fcd0a2c85eae
z05e03d10952fe00e88421987dd72ec11b85c69fca60ee74e65bf2245c4068224f2568490665848
zd75d07af95782681de2ea6bed64fe3af01f6b1ae02cc70b98f64e3a342da7404d2806531aa740f
z99e6c149e2227cff6fd59087c5cb3fff8506c09cb62b11d8eed4715c81f54d0bc573b2ec115986
z37300e20e065fd9d39e36ce0d3ce92d0e2a4e97a008d187aa6370a97ce4799772a4dd3c63b6b5f
z05cb6509131a348a51b7f1b59855bb476b57df2d4f6d2a555f40d22e44396b84a3d46899eb2a58
z4f00b19bd8172f6cdebc820e5fd675a341700c5f7796ff4b1385b51498bafaa7d4477ec9d93cba
z474cd8a5a178a5f54781947f7e9b9bbbdc5361ff577fe791a25f29d2cded52d3c19bf73eaf5851
z1774180b0dfb3d980dc2b65586e3723d86955e0a99a6f5c370551e79ad9fa19a7f9f5dc4387bc8
zba46eb194fa6723789d17d083eac5b0810a758db2dc56b9e1e0bd524003b36eb5557ebec6a90d3
z16165334b6a09dd2ffcbb66f9d21c12d9326020281e48c05d58a8558112a66ee20b1c75acac263
z2cc6dc548b3382b92a1a087ad2bf78a10bb1577601403deae9ab11167626d04e1225f24b54b841
z3230cc648d8c4e18f5206576a95c50781af51e040094cadaa494aa0467003676d74a591ee5949e
zf2c039ca2d4066dd54802b1d551f7cda408a9d30f59fcfadbdc6c9ed6c4e0927126572526b17e0
ze36db488c47c459eeff8f5cf277c38a706b4686560d449b1c749de13a59ad75b609647f5c9c8d0
z98f2aa56188ba549ed6688fc268d9a87c761f0cd9f33f9a7add57bf4e3126300487babb04529d3
z5740c41685c746d7d7c6cc097b14653b61ef7dca1a83ebff300a9ae7786e8ddf44f815bbc36cb2
zffba76419912bdcd4e291190bf456d1d771efda9b3bfd53c50b1c32cd8a42e7b4d9159063b4b4d
ze8aad4cf16a342e8f80a9d26e3e9e64518228a31f626319446aabd3fe6011c956e8cc0faf1f1f3
z5507486b5cabfe67776a72b529b7f7f9f5138fa7c72b5b43b423c2abfa135233dbdd8b0469d336
ze840248b6131fd39376d47efe414d8b1e125422feca9a9aedc38b26e1150a025f75afce45417f1
z795398211fa28ed124f682369afbf54909370e547ea1d636863161e21a71bcf0cbe7abc2740db3
z608aa2cebf631da796d51bc0666d83861eefc42b39355d1b3de417218d285f3c57ca5f6175e27f
z1ddbb9e4b02f54616a778e0c3676a5842bfb3198b1a24469b4e82df472101f2c12884e97b365cf
z90a0be9227e174eab056cdc299b184ffdf9bc1d8cf5b0a914232c500395aa83a8db4bc0c105d2c
z2369d491f8edd0d2c08bac8f452afbc7da0331f26e7e5961654c4cd1a64abef75ad7905edb8289
z2ebeb150e0e784706d69df2ab86c34fc1081eec61e11e4b787e8c33a2f76c1716204607d0a38cc
zfeaf7dae719f3ac997f16a78cf4dba0169346dea7407ce7dee1acf57428d4ace1c891974c54a69
z5136c06a4dc085f0cfad909185effc837d8680624848b3b3cad63d1260989e3ecfde6196fb7995
z6df49e3d2c6669bc97dc9a915d8cc7310ad746c504ce9fb3900b6be7eab4968c29059454562312
z82a84677abee90ed8ded75a53994f32f505076431153e04a3452f5d8a96e1393e6954070282b70
zb23eeabc854ba5eb51dca69fbc0281ae1c0a53dd0631db8eff52b089f3022e9999e2d903503b7d
zb9f52369ed6de1df7660ff66a46aff236d580eaab8aca0ad824ccd445e53166e06e8636dd8eead
z0b6bb25ea7e47e4d13e23f0d92bdbf814cc2ad0b3bcd760db88d96d049a52f61da2e3711449b85
z2947d29257eb473d0337709b3bbc0180edbea714b9474f602fe9c290228fa111d80f5f6d5fe1ec
z40d8ca86a7462902487589b0d9bf87872ef719e2ecaf0c686b0dd0199dcb7218075d4b47ff519e
z0c5c15ef4a996b294606b61ab4688ad399115f607d99bf4977b33e56f1b621d1b7d145b5cb31d9
z9db1d29439a79f1752ccc041fc809d5eaff7b3943a942cc537463bad91f0ec816c9d2b7cb18b48
z495dacc9efaaa987dc83a1443ee15c15d0c2acf386cfbd0640dd6fefbc78065c14b672f154a8fc
zaef10bdd207acae29627b25cfc7417bf5286cf794a7aaa5b8f560963739a580f7b054c5c793862
zd5300402ddd8555c826deb7b0baf947ae726262f920a043e868a5e740246942cd5e0f9808be56c
zc5798da257eaaece0e521f43ae208f11ac95c9fb7407268fba130ab1995622e3eda591c99cb263
zd540c6ec83c50ddad947572b43db7546da5981fb919d754a090cbeba57ff5a16f72aecc8422242
z4cce20a3b0c299b5b8d0e3128b859bd7205ae766a624bd3f8a629068cc28440a3bd28d44348dad
z2e7d0f834cdca5602c5fa2a3b803db6c80d835a59b4424c95d97233fb24b997da5d5124a2ac1d2
z6b8c7f94eee8350d94965d56afc43a9834aa88defd94d5e2675cf16c82748254aa5e7ec4e8ee39
z19c868f3b736304a42798ced2ed3c873aeb737e1e92d20eee6ad15c1e952724a4293cb58c32840
z2e545d11ba612d83c172513e21740381da3fcadfde972a0005dac502cb12f1f18cdaa21895c7e7
z296b20bbadc00d7fce63d0abcba8c2a81c13310e86c64e993c0df8dadc6abe8ac783e6657ab5c1
za459a0ab12fb9510679579461e07f3d0a055591fa144729f12afc712df49198829ec70b8ef3d35
z6214e828b143a73c5e521c3171c73278615db42393b5c3c42cb22e0742e79e8ca65788d1c15abd
z219f6a414297497baec98906a4d81e32d98fc774ede990d78bc6cd80445ee2eae67427dc50c34f
z197af9eaf349176b964b0fce185e926f5f475b468420fe1630b83ba490739cc243a2456a43219a
zb49eceeef89a7220e685304a2a7f34adab0ee396780d63d824d6c87d26eb1afc982d3dbdb22dea
z3cd84cb025c2d10cc365d28772beceda7b8462f772bf92c8350754013f422c1a80f38de9b828cd
z979ce9706eba0a2ad2955954854527ec48b05e44904eb7ec6aa11686288bf9cba8a58ca723ea96
z1679ed424dab84ac7a35676bc3ea7e062ba16e7769d53b9a08fa65ad5ea42c3fe6b9752692006f
z1ac001f622239b657529e73f30b6a2e88377ebdd4bcbb6f38779e5430e0014f0c2a8fbe40605d9
z2e64d06808868204a0826efc32a3ced927f5b00062b10df72437fe99244ac778902570cca931c1
z38f902f84ccb321a738fc70c445d9a50440d7be95c0e0831a7f4eda8dc5ddaf67628d07ea4f521
z3e6dea2b68e9d027611974925492ad346056ef7414786f68326c4add5cae7ea179ff798a233d56
z50df51481d6e754ed38cba178fffdd8cd6035c00714e50a29fbaad5f0f4fda0da9cc34db54652e
z7867c73be96fed0e00c426bda976bec50e3283e01af08ba46397ba2601c365d027697a452b088a
z04bf2ebe664efa528b168db17b3b091bd83887ab384caa38404a75bdaeb2365e2b1ee6542034a0
z8bf5e9f30e5d8be6cdf95ae39ff2583523cad215155e8afb6d3202620d3d70dc2fc67b38f38209
z00da8e489efe8c4f4a7f8f36369fa83b1e1d40316fef5c008e20215f0a22c75fe7e16459a72f69
z5319264202f7fedede6b769178d492b4f309ec2dee9c963394c580ac80d70d9f482ab25ab4584f
z577228a5654e4737c5d4f60f567504dac095bcadd77ad5a1e0f67b8b1c05361d3f74a97c25af09
z127f5332186cf89ba1885a3aa426ce088bbce65b7beb9689d2083f16feff3b7bdbcfde10cf0cb7
z571bd88bf40ce807fb58d1f54034bb94c6842ed9d1fbccfb3dc408e3d5cc44b9ed2268fd67c61a
zac6668cd15f8b2e4ca3f0dc473f64b7ce435bad8d14d1f77888291dab4966ca3ee33d31240f7a8
zde3c57fc7b5cb462fd21e48ac2826c40d4a22a7257d234a67e905e2b20aa396b94c8beada0a54d
z630dc97025c16e4dd118432dc94bda35b866b9557744a993492424687e170caf13c5230d6d05e5
zb8644da0aaa55b77c3f20afa70560f6d9553d6375e091ced15ba3ff8da07634a565453bed7fb76
z5a55f135c8a24a8a5743c6ea91de11b4f1897f5563ef71c48e0ec3466aed137b97c2303fbe2fe3
z06c2f2bbef65063cc080700d6494b742e43e6b44c95f1d17e93ec3fcccb4d4c895967048722f31
z6a41f6efaf26eef6dd088df7138bbc6d227da249091ee782a4d5d8065e88a646c942125dbfffb5
z6da18ffb8c229e67f5e4cc966cbff64f8ef1df0709f724fc8beb702679a594d32995d2c6bced4c
z830dd6248257d7d35390abb1e7fedda82b1f6420a05eb07315f4a06482972b7a114934910f13b1
z89127f1e207c9c86e4bf01c38e49b32b1b1494997066ff6e14434984db7541cb1c314b69d14d19
ze2678ec7999fd2ad0e90e7a13e1a839281dc46ccf0ae7a7d0c3a6093148ae5bd9e2239e4a2f793
z51d893b04263e5cff81317646793d175276434dd3e4aad3efa0e520d9b1960929ac50d44e8c654
zaf8d5d868af48399cd0fe43f3ede43f1935e0f3b4cdf1ca8672fdf7a38eaec1eefbbc90794f66e
z51e25e6120e432a6a60d78e164e4af0db96acdd064083f9a1899b9a70e7f2010fb71c943221ab9
zb298fb152c67acc67fccb5c69f2befeac5d4bf36a7d8ed80739215f07d4fb4e9774a488bfac666
zadcfb6b265fab40a2290cfe06c504f957809d2171f870824424a9ab7d75532259d8e1d44d4f5a3
zc427ea0aea94825f8a7f5cfc3803636f4513e48f8742567bab40e1f8c688a07d32cc761d6f82b8
zaaf3c44789501b2a601bb43d56d73545356639700a85128b882b9e4c5e5f010cbf07d21f90a407
ze2bbc23e31be959b0e1560e280765d7c1f3a232c1b1630a3604fdffb96d2558ab5942191f9c986
z5644fbcab77de92dd3793b0f75877016510b179837933200576f06019b60ed051a6c9b54db8f40
z1a9cfb51f05bd5e16b57acdd81c472a10411435757d5a972b5bf86cd57ac6fbc56218487f10e84
zf887eee08a1793b431a9a6cc6ec7cbf9b74f39edc771232e12cfa95a376a2b2f2e3192961667a7
z611feab142bdb48545150708923bfd72b1af296d2e9e9aa194c624a3614492b735b799a47864c4
zad71878747598df5bf0c84f0581a97f773dcea5db6bd51b8d248499de5cfe878009a71e9123b3f
z0436c045690ce3961e66b849ed865f3059b11d43643d98b7ae97a1e170b65009d7e781657dec64
zb4a497fe03a77e3f3308e5fd31881e5062c2632b3a2e37bb861f4a9ccd02f61d8b96d9e9738bfd
z471c1bc1c55942ab7596dc6cc3086488804278109154a13b2afa21d4e552d387eb92310c9fb47b
z652fc155dda87bfdda6ab4e99be72cf2355cab4ae52f85f96d800b02889a1ab06046571e6bf4ba
za34abe79ef64193e66e46563f3d2d71335cdfbcef9b99977e8190eb9cf5af0e89966adb37f2af0
z325c1fc1d6c5b5e0ec6346f9df220e75b065193c11f7796512a025d4882aca3017339bd737b1f5
zf89244bb8b3253226208d0f87b258436ddf1ae0e6ffbcdd38c48b7586bcea961d7d856f08a6b74
zd197e3c5771da8569b40bb1b0b5b3a7dcbab9cb49ad7f74d5e537e1d7ef85471dd1b25031d2011
zc888abca3a26d1cc15ce3fcc1dd14712f7184c7de5288dfa859ab8910f41fd8d31b4baa952d481
zf6c48fbcad0289a2683dceec522f399ac8a8a65bc81efa139acd8eb3dc3338689346acdb91d507
z6871b64b5aa57f760c6c44b1afbc4e441df9eff4d531645a8ebcb5cca5ff72a8e1dabf3afb245d
z741c2bc2ecebd37acd25441bc5577802c3db5002fec580e538aa9be4362e48fb950ed280b778e4
z1d6aca478d7a4d3d1d19be8a251904db164a8ac32c29441bd32bf8f9d75368465289cd53963d97
z30498c539b05f1bfac895e464f9148215acabf0fd654b5aeae30d7d9fc7a588f7935e2f0a3acb6
zdda838231755d5a8d71a4f767b9ba97b34f4c7c5c1e802acdd235239b50760fcbcfc9db9b07d13
z4c8ebafd9e840613bd0a8a9b3add693c59540748dda322813903642362658c8b4bbb266b5463a1
z0dc7c71f1473067b2353c7c4b6da7183d742f24a3abbb47a7b7d79d617d3905726a9d12727bd01
zf441153be525478a5557c038d859facdc6b7a3cd66529d8c8966bd6f6d6c44fd6ab0f527d72041
ze58f8c8f2c6e55d0a6fcb4fb9adc472a2536b2fcd76bd2ccd72d0ed08d9cf4f48198d1bbeb470f
zc5167e9b0572681ba049a193b122e4fce3b2f8e8a81fda821b5b589fbd9576f3dbd09831553ecf
z467e0cb5f7e2dae1be1e949c85ee7c13b6b4f2f4db61e39f1334efb96177e6e8994df5e0c266d8
zaadcbbbb84170fe98ff418320a84a3d84039d15536b5d73269d9e2d3377839d2b64a85275af07a
zd70f0fd380e3a74478b3918e12e989f01712db64be1ec07a24c2fb34643abbdc1e0216443445d9
zca13f7f0a8471de69cdcba615abdadf1b8ccfdec135b43e48c8a5d13f69c1e2853b8c71a6356aa
zf88ffa7a0c0e2d6b4f44164f2cf0f3d55610e9cb488e99c14e46ad2d04435706cb387f8fb96396
z3247d7cc5ba193f569b52d68bc3dde57dddd2ba135c4c7de4983db77aba3f4d7642d86c20d9992
zd045b7fc19da64d3e692c8438fba961f115afe0ce0b60f89f90209a9c646ac72a280b093710731
z432ae8539388710bbba126d766027d3e1a07f3dc72b5caccf879fb005e7c82817efa42120fbe6c
zffbda4e9b066f5d33fa704c40bd80400b5f2ed18f98ae6fdde78a01f9bfecd133bd05b57a4cf78
z04b50fcdcefebd666907d45ed72408a8731dcc3ecbe10b680ce9757a8dd92afd85a3d48656c448
z43f6540be7b1e3e767e82b9e3e9776fd3afe2325853f81dff03229a66f81aecf612c806d73c530
z66d31928e05157ab426ce0bb636d658f8e0f4dcfa855b648258b355ae7a2586155f8a758906e58
zb221b90804548382387530da0b724162fdb72985599971fde396b9e4fe3f30fde71d6f4b59464a
z1b22abf568151b3a04382270584c5dab4104bf34c0349ae2044622326abd9e2652f396ac3a8553
zb12bc4c6f6b631910603ea918570596ab8504abbd0bccc6b976ee60c3d64e4c22b6faa50052acb
zef0b6f4151d4cbecbb3f79b0957eb748ec6f8a24136cbcfc90b74ae9ec977d42419f18e8e3ba59
z23aafdf0ab74dec45cada782fd295233d8b751bf791ce80aca7cf765ff12e1e8c75d36b0aa1294
z224d55c7c0e90aa5517bbab1acd910e753f1c38ff6c66ce8d508fe1ba5b859865a3d1201228d1d
za38307ae885ef5638509ef96c615a1e381eb9731fea8af331f456907bb59bb2f08e505da1dfba9
z7ee7414c009e112b11fa3ac0b5bcf1ff5d5099d76e492bd926f2e5a27eebdf75c47baba19f5dee
zf9c3bca309f1694138826097582cccab49c5bc5b767937fa6e737367369f47080c3c85e206b484
z4a5d3a32b76e0b3d33e88a4f5456598f7695d51b265fa9ed89842c7255565a65e6c6e186a4b773
z7c5aae6a004f99d9ecf30beadea2e80982c025ca312cf4eccf0e310343bc2a8e5f4696a7068f89
z853e63c1edf346f7b65c01314fed3565a8793bbca8ae3e07d98339e66d4c6ea0edbb2945a59810
zb3bfa5d82f7960d1060694c72f94863f1e8f30f384653e833f07b8f508197b13dc8e9cc94eb2d7
z0b2c9db2a342ac12e92ee2b4fe2fe678da70dd3698fdd834f8d9779fc693f2510127c8e85940d5
zc4be84d960f775d3f9bb361a39dba9086247e4a00983bdba7ca15b2e0fc3f83b20bd8b9336dece
z37494d0c6fbd2df758d5c36ebe663d390777b2626fc67c281cd62b08cea2482335a5d924bf6c12
z4fea54339966a197891231e90ba923fbb8be4c6309dac526283021f38e6bae47afde5998679078
za8e59e745b35a50693c7dfcd7018c62d86f7fd68eff9ad802fe0c8a989b4f632d9fbfc2741c564
z801844adf1992d97aeab39aeb80a57e4d2b96522cb677689611037aa45839e94a9360559e469bd
z53ddfe2fdeaece98756b3d802f4620239556fb775e5c4aebcd43a10c6c2cd9143f46a62c4b96bc
z5aa194ce3048e0a1a7a4243afb6cc4d2de3b024d2862dc6599d2e760ffa1dcdb878260882f5509
z0e84d6d267a1e57db494701af34bc32ac3a58703bacaff7fbb0709f7f14542ac615b56a05c9085
zba6ecab2ce67a74fb874dc4fe996631ba8ff4951c3f5b007a8d0bd0f03a2a99fcc4cec823eedde
z3d1a1971b509d9d95c021203fc7b5ce37955aedd3fd780a0558b7d490028f90fbccc155ce3c936
za9c5e2b0716d274a1495259004bd1fdd0569dc28d1afd78d965a7f8f701192a8fcd259c2f5fa24
z3027678939b874ec842336f8e8277f35acb578a67c8c598bc7d1a7b7624440fb5aa9cfb1b5a5a5
z725320b9707358f5b5f1fcf93ebc67cda0e559baee5ffdfbbcfa12300971feba4f6725999a629e
zdcf96e901f5de1f4dbf35aa25f8aa9e93ea2f12deacf165639e378c88f2b67f807fa908a554a83
z32436d4b614a0a1f817313dd7332419ec4d6ca9e68ab578b3dc18e307054b2bb605a3c94ddbf39
z0c6c0de0ffd6bca2bfbc2613f5beae49bec470afd36d93aaea596b373b12ab82be36a5df1ba83f
zb2c790103567f5c40d27f24e87f394e89fd862d2c9ab3720e2d6dbe25be50f7bd471250b2efbe3
zcdc5185aa0d07e56e2a0dff1bb60b62ce67810440ab598f0b9242de9d38fde0cff4a2dc749f8d1
zc54613bc2642bdb9536b2284170ace9bead7e54422162d9bf4abb1311b5630658e2416481b61e5
za2729dae7cbcfaff315a0f6993b7af3abbbd1f989e3e8eccbdc11b184b22e603ed8bf083cdd13d
zb63025e2bd550a847a5f8d2c151e93dc75b403a0079a1326bcf7587b06dbeada7eac46d3d69bac
z058a0aeb3ed906e1b3717e6509f86064020e0af7c6e689ae95d26a4c173249d09f4930a54792b5
z68a0762e2d902b0cdaa46b3e6f894554ed4ff65af4903a72c947a44fc3738305f7dc0b66263401
z5a994e5ca5d250707dc7bd0d6e84c3261d0eb55f2455157de1aafdd1dc34084f9ff9d9d7ebfa71
z682017e9284caac934cedb9b9703ca60fbd9cbd55203c778cf6edd19cb467d44afa82ac81d802d
z5ea85889d88b673d7de383b33e5d28b469d2d26383f371e67b3052db48c59ba1a67188b420a146
z6fb3828bb00e75c2eea0dd14d45c9f8806102cdd3d96d2aab212d54fe7b586fe2083687aea76cd
z46d20d239401bb0bdddf1404e4841b13c13497df38ee7d92537b9fc076b78c836502219ea1412e
z1840a4e0bdff7dec47fe89a5e21561074ba9f73037292076cb8835803d8205cecb0818f868aad8
zcd6890e6d7818fc454980885e916857f933f9523c0a193909c874eebaa01532b595f9f47ba6c9f
z3c754ca671f1ef5bd49b7fb46913057783dcba22f132c901bd5df9bf7eaa608c53a6e28ecbf8aa
z305855a21441059cd596c2047222ed3bf7f0e55d3c12885a7df8b99e34e1312f25ede658424430
zcd63f59210cde7bb374e1466ea2a6c4b005327f6d41bc465b7647acf5f777eec003cbf85ce4939
z784599db3db959c33d013ae56e0adf106f90407a91bf5cdb305516e422e5e8ebe0f27161798130
z726b5c1a3addb336a31b508a479ad9642649e23ae9e7feda9dbfc09fa01bc4dd602876c4999076
z3491dc44ecbb28ce0a37822d4102fac27bc2077e129c221a38c609bcb223c96f4d4d0cbef2c41b
z9a0dfe3df9b886c4ae3e83897ec4aebd481970c572c45354c358ab752d4a5dcfd277faf62bf817
z6f0258c6f0dce55ab8ea9619915b2a4d01d96ede1c460463b894983f40a017bb5b33126e3434da
z739d6312c31e11c8d8f2bdcccf074c7a86558a1e8fa5da430e2cb172e7d536e0a823f45dba5c17
z05f96c4c5a2bfaaba35d73fe61456792e3023e5b97db74a8dbc4327d38500c0f1a4f679ed439fa
zba9672394b004b550c8672d5dfd017aef255d316a208ec59551a833d1b54ade15b673d4ff18fa9
ze9c4c8c1d046d966e2a38ca5815aa3dde8fcb71edd169f4353266abf1c4c2d6a914a22ec6bf90c
z330cdabec67fce417bdacc0b3a3655e62286188bd032b9d8f77797f3c75833b168f539d0ca9ab0
zc7b937961ed89d112a4e74f3596ed983b04a136c4b2044dc05ff81a833d196c14ef8a92693b5a0
z6fd8ef5a8e47bf16be15d1fe08426d2932c022cfc309c8862c17567ac021f0a054ed2294f4c7d9
z24bd935d2fc68b5edededd58492660ec7d294826dceae1b36d6449ce42a2a550a0856057c954d7
zef5aa90c7ceb4593ed2c1386f86a28e36bc1ba19ba69b79449363155df2b92215fae0871088262
zc876fbf8b92cefdb22ff6c2c5db50f789682a5b3f40fbc5eb5e0f275b83286e6bf5fc4c7aaefda
ze0415a48eff31245e6f23a1ca74682aa421028327af6e35affbde65558f4b3f397cad1f9ec6aa9
z7c27c9406f127bdf1e6d91ddadaa7c36dd8f3919cdf31c3b311d3d0a987a5ae06c9c1e45469b18
zcd6dafb2c2528c49533e50208b6e2043a1df11ea5d932bb2d1d9cfbba34de3a81662a43a7c9c13
zadee8407567a2a450eb2605dc0308de13ddc1c16c056fc98a7e1d63e69fb5d54e53be00dabc1b6
z3b8a6e32c2ea5983e96d77270e25998ca0a5273a1ea9bd42789dff09034b45b30eb9f5a331df6d
z5c646a587d52a6baa58871da90e9972f80871ce1de5143a54ed3aa3a29d5dca82a623e36095f1a
z6a21e10d7aeaca9dccf28bd4e6b37aaf6d4dc3f8c31eb11ddf42767d4999278ccb1c9e789e6b4d
zc147732b7f352baa27719a3fb055d64cfc55962c6502b3051a2986ea0624c1e4d931e9d391c452
z94002d771a75ac87b5e5331091c91cfdbe94cf54ae00603bcd4b819ab7d619d99d35adfa986c67
zee65fb8c49f18a4dc5feb4633c6a269dd3b9fbdadb248675768c148a5d3ce3a4ff2abc12431226
za0928cd138dddcae84d9b31ab76185b883422a3f9d9dd4a5ab5675ad1df076d98290e9c21e822c
ze28d5baebdbc217f6d9fde763a2df969a7c67182524fc0d4f81595ed00dcabce5f755a114581ea
z258d7e5779454799df9fcf2ec51e0e8d19da8fa9726e7ab7840d678e3d32f17571c11b2f1b669d
z81805ca89e0dfa2e769c75f957c4633b6f3fb5ef834601b6339d87d612daa707e3e363f9620cd7
z1eeba83012d33f8b29833983f5b65f64d0a0ec8b0de821d689bdad1c30dd2ad79fdc7ad33d8b37
z65b058674a24ab968833df385348924705d904b9ec7a4cad6dc7ad9b9fb7c753f8f81e89965cd5
z65ef89b643869926a3a3619d31937a91c39c3d101a174b2b34309025ef4db4da3540e41123f03b
ze995e66d626d77f8bc37574d20a60d9ae531575448939d66045435fb56f1b1b9d9ed9cb0bff601
z68ee1a42dd8278cd290718dc4fd073640fdd78558340cdd1a2cd38271bc6053fdbfcae6386294f
z064cf9b73846f69649fca4dfa832b6b29362db9d6eaa0e600706deab8347a6a10871e9d6037418
z87a00ff81687b0739e95ed90026a2bc0ecd963afde90518560f14c740a37c5d4544095d55e25ea
zdb951d204e75a4496bda1bf1526aec6c62509243169b3cbb92d17e47a73410aab7d9bae86be313
z08ec45d4114884f2f6aee2921bf9c77eddc522f55fa5ce18de921e44cb3018cb061e855bc8be07
z62fbde62bae0386bcdda510cb59e3cde0ae6f337522edc8123fc2b8448f170b0b18d8dd198ae91
z16a389cfdfc832cddabbd6ac0d6c51ecbf99c6ca2b4138ae945a5f9f61c58729db882eb9f0c008
z32dedc050444e6bc3e8fe9bb36315b09ee76a2f60a4a52e4d00a95f07a8e284261f79bd8d30514
zee3da5190f18206a34e5bb6c133531091b6c23edc9341861e45afdacdd8999db68d58ffd94d298
zb1aade617b8e7a593773d4697bb6cf37d35660da51866f0bee4abbb0f7446ee239dcff6dca780e
zbe84d018fc43ed48780c02473e27fe76ab10790dd45accc4a4f9260fc4970a037a9fe76e26f3c1
z1e6d04607130c5a392340d034bb4a576949a6df9c187577385a9da2c5e76a0791bce707aea3003
z9b125afa79e56bbc422b9cd0083cc853f159dbce0d30ae8405c4a974b59b77eae13062667df8a0
z38cf5a6d24de038f4fe544365194a7c0684a8f6727f7e5750a7589fab6150e07679c96915f135a
zc9f94912b08279f1a1c41bafd6f4465ccf260f2f865533e488734bb80558590e4dd6584f6b5635
ze2af165ddfd057dc718692e61e8ec2301cf2efac734a59faf5897f47e95f855a3fa7bf5d3d45b2
z8258af7acf8380a871a8e37d0d2b7acac44bcf7af53c816a9302af13cddb8e9ec5444d7eaafc52
ze81175775d7824b81f280362b75c9768b28f1094d97ecb29131056180e9159bb38ecfb409e0012
z4dc524efb63137cd919d3b63c494010a23403aa39f509d361cef8598be8cb267852f6d63f764d3
zcaf0cda26b36b19f90e1836ce0f3f55078cdb94ae98908369d99fce7e110e4a9dbc32698441b4b
zec758a678867555362c7e5ac4908f3777299744a161bc5014b6d1a052628817ef3fed745671639
zf8736b0b145683bf15a5bb038489d139ddb1ffc1f2f2510600582d6cf3c519677511a60e4b9d32
z485ff36b95e2bd104a3a914b7abfe0cd9b0736669f2ea98017198821162fa0ec73a91c1b8ba5ad
z65331be860543e9134e41fdc6bfef50f26c50aed9c099821162efdf60d11af8515826f8802a35c
z2a74a9b788e96f22b82bfdca4829002c7b8b5574b26637cfc504017d9c91153db8475ee74e2ddf
zc6b8e0d807f8620825dd00386d0da7e0662b31f0114700a7356219d4d58e0101f5ddd1c7eac013
z40130571b9fa2aac22fa7c0eb32f971f2c1718de4f2a6addf5f427fe77dd28a508076868ba6c5b
z17c8759165b11e64df218f86e440281f750651f9fef73d6fbc73ebe47d4787a2b4aea262d42d23
z5a08d119a9e80e0719e34289147cbb888dfce1d68f7e030fb8519f9f582e73696639f1651af7fa
zd7a5e54ab58c3f0f3002279e5d927cd2198f823284f467f9353021d215c42eddef5d2d39ad9cce
z85a63fa927889ded954d9f9767e98554ab8b856cba56e6a1d97693f523e22f5c975176444b291d
z790bed3ab47b8440da03fb7a1dd6544b0a11450f6ddc0bb08103f1f8ff1c31cc630462b73363fd
z08d243d5aa62146c143d15a7260a571fed584b696e1688842862bd4721be4863e19b17a71fc53e
z5b7e4f2e54373ef64c4e94146366ca610879c2b713360526b971e7e0b009bb2410bf03b3019b29
z9ef6d9b3b96c54a6450f7b700d205785fab52a474c11f7f66fea201030f9715d55eb558b85e4e5
z3162ec244f75e82d5e1fade78bba58697dccae1db082ac32f05b0c945393b216a4bf9deebdca6b
z2467d9b0c9490c9be396f29f80f5ea695c0e35d4f32ad526e59b99c9c0b1eeba692cd57e541021
zf23737baa9529fe65f543554d58979c13c30e4b661e90e3ea023db0b9ce7067ce3cf2618ecd2fc
za1f160f8b2f48d2dd7483a719c1704fa27097a3130636dda0716b9c5c44a9e5b1353a9876eed65
z3278a5096b32372e115a967acd7e4ef1aee3ffee1a2be5268b6617e8914dace617563b2e867901
ze8b3bb76209f14f623f418ea8863e6954a19187a99368ca0e617f79fb4f8849832603dce497d34
zb69a1225e7e3d5db55e77c39218a375a5c6e1d5db6f2da303fa244b9d5c054a5eb5963c5c4eeac
zf64d57be1f8950de00dfe2be546cf8208ba08a3e4c3c1c8e1682ed63025b8c582f3df86f885ec6
z0005fa02f4cfbf17c829ad03e8f5bab58b4e9918916a40fc21cd9ccaba0355fd7a2fb297650f51
zeab50314c9eb20ffba6d95a89002c1dc64f5a09a291db15b966116e0f1467ba19a4c43477bdaba
z10e673230f64baea0e25ac83dab1ff1e80e34579bf6461d1222291f8c19213e33deecbec4ac056
z013680c6a8addbc03d299c9283999d895cf7ccde65ac12734ec58b6f7217ef7453500718299193
z24b8b6314beb6bad88caf9594a918536f431505e814e120fbacef099fb2668ffec76b8464b38fe
z2b19e979d988d407c087fd4c3bafde3e5fbe1a4ced302da8ca1a66ed1855c2246d348d3c2d4516
z34857a2aa446b7288b1688251de170b13497653d57f41eedfbf6acaceef9bf1dec519d00ac3993
z2b9e9b3de91d7511e9cae7796f492e0ee343b5fadbd246c02db45c95c971f515f52c13c9c6a67c
z550aa7825612000468febc602222ead4f1964ad4dc294320e6e6267cffceabc515ebee9e8dc139
z91be60163d934bbf64db112643e6319bb38d391d16b05af62db11fabeb75bedf542277c8d40762
z1cd1a73d7f399901ebde55564ca7e344e9b886e7a5b7b8dffe3c802f99ce39ebbc8571ad3fca1f
z9c19907b33e3f4c65d0e45a8fc7201cce37d0377a2cddc46c1bcaded6a64843e9ac18a942a7c3a
z864b3c6aeacb28e00abe201774f08986b624a4fe99a18a1430f75ab8d7a287db2feb9bac4ea714
z2d4f58d82e0562b5cb2c3c3eb0b8fad8de873b123d6f86d20e691120eeda41b95d2d664778364b
z84da13fb00a017bf107cc9c4c02fe75d951ecf5723093529ccb6b53e55e7bcd59cbab8d750a572
z52830e7f02012098a5aeea86ec6a04a6eaab587e130794b0437d968623bd3d2a9bf5d31de5e1c8
z2c7f094ec23e7957c880b341e586994ed0fc460f6c59a339e9a518dfe739550dcf20f9dbe6cca0
z9081308efdebe52118838f96fb730f81077824a11b6b902af0067e69b06a3cc400a79323c2fd62
ze9032aedc665cf477844c6f11f672ce34fecb03310c8056eb83cf004bd06f24fd34f02fa3937ba
zfd362453dbb69fd6955403db19a358a6dde8157442046dce7c3cc6de060a90c62637e3a7b115b4
ze382f98b33a9bc87a7c85775279e9dd24f30415fb81a4efdb06956aa4984319e6a12bb92e4f388
zb4c368a59f53205996bf6f2b4a099c9a2f160b8e1826dba620398084852906a9523f7152ceb922
z81035ea0168e56934dc8b25c05cf28ebe894dad4799b342785355775889f0e57b67a998ad07ddb
z2d0ea03912c06d337b7d53a3940ef511d1001a7579b754bbfc61bd914f99d9e74eeabf9e9f75be
ze54cef6315cf9847df4d5e7d5275800550ab6349101568fcf986734f1d1da596e5693c98821492
zf6836e6bffbacff5abffd30fbaf64a9e1edfca6e5cf8956bf2ad302dd46106a96cc998b6886b9f
z6cb3adedc862e833f2594babfd4f3ec98dc52bcfe88c14411cb09601af982026769751bf2f8cf0
zb7fac84efd52436e02bebc9d5d95cd2797a1ad887829bca657a4a2845f3c4c6ca7d9dee3d59423
zc6e3fdcfdc4c58a8b563d947d924527b2962a8e7193505c94ce162c69ab5a01019d5918720e118
z28dac65c906ca373a7e8dafe62d08cabde849c267ee10a2830c3dcb9e77d759e70a41a3100e153
z66952764051a3a3028c90eeebf8bc03551f18b00e7f0ca0dfdf9f899029a5d534b69705b6d5768
z37a447de249bffec46a3732e600db20889761dd205757cd7973251da315f9459733ab5a9635db5
z823688e7421b114611c079a62b197b27f9726ec6793f187aa805ad80bb2ff501c1dfed7fd623f4
z6e0a7d94ea9f76bfae142d6ed323201b52b48e0092298721a90d2df7bafd17b4df095a1e32df8c
z02861ed2489c28da43460ba731786cee90d44aa66b88e3f8bed0ddaa256f24f734bb312d94a53e
zdb6f98d757d74a66f6dc383db384bbcfc3b7da7224d4305f36c438564df873dc0ede4e9931fec4
zecddf8ce6b135e6adf1f2d4844820aba376ad971d4db3dad8126d6aba13578aa93903253138c8a
zed703023331d4513ae4b48f34011b8b41b191fd8d7b281269594a6966a61b6c7c36955f0854ecd
zc64cd33c87ac5a68589b9a99d8e43c8d2b4c28e6a9bef41b26fe9945be4761e0a76b146fe88116
zdd5628657a04dc51049c7f81ba243a540e99c51c352998375b6f8ab42847a30382cf41869e5ee6
z7d874e7a27e9c416c34712d9dacb628694346397c2ded1f86e2e752195e89c8d11ef76a61746f2
za312c791d6376eca39b5f0658c71bb5e454d051d6dd1589c48051887d05862ecc922e06930c54d
z223ec9d39b0f76344fa6819e12dc8d87334736ab68b889ff6565ba3658281cc39ad72de78f4366
zc22c332d3319cbbf999b3a4292c117588a8bac0357f33217e0e0701d1b4c89d915a30b32286680
zd584647a5ee018b782ae9826d4ebe5b6a4ba72a72fea62532cb4ac41534aec0f05c7a59fcf9681
z7db19ffa4bbc75fc7bff3e2b93fbe1e452beff901478c9c736ba9af801099f5e23e6041adf06e2
zb06c91fc331037fc521d4222cef6cf5403cd63fb60e41f795249757e667eb9f9e9fda8300836c4
z85f8d65afc28e39df8cf297c17ce25187e19c9f23d352c96d4f0b66182d174932d6c7408f24639
z0eee0cb0319f78e7f9cd1b56c10f5330aa82bf71a5b29f80d4316e7f9ba5f1f4c1acfee9233282
za08b48d5661f6f1c0c515b5a2f7bae49d6cfe30d8176c230d2f6903c311315a90376ae5728840c
zc843f096ccf89d539785154b3a210502c1206e7f5e92de6f84e27c6a5a4703603ef7b6d195f607
z075e3d7b60ab22bde5a4242b651b368268799779854e2196dff8d3f5a036921d26ccf219d9641b
zc1180f5248a9856af09fa02e59145b315d65c13c7b2ae58499f9c6e4640bacb35bc9fc03a87baa
z616cb48ec4785b516ac5d3fd044204b86b855aa48724903222d3fb4e84d8cabf810d2d97fb9fe6
z8f8d5aacc5899953fbda4d343163c3164ee61c882ac4bbacd74acb0256b2f7a6fa1ce5d09daec6
za296d8295a3b6726470150ede951fa06f7a2d9e68b1c357b9c7b1c708c5fbc2c477fe7ddc36523
z632da823bb67848ec74275425964bdd775f81aa69d54be2241721abf49e6c59171bbd05d8c44c7
z072ce33c11b82df9e03046d53bc6a70c1125b129e3b52aab9757749e6ca345f373ed0f3dc50b77
z5005e4b1b1192108c7b421b50983453365233af343e1f819904f5b60005bc4fb70fd19476f6acf
z648d6e84fb1c4b20f04a85a727500f8f5e3bda55b19ad3b31d6fe53dadc864b85d2651be94990d
z214e1c6df18bdeb21db9857c0f799252ed30ce11835bcc02049368d00b981449d5eff40a559728
z9ecda25da9cd8c1b36d205b0b17c502035aaff1cb0b7bbf284e743d483d14346fe870ff0debd57
z029b68162b8492c0690ce8505af87c5c6fb981569a9749c2aee5d8fdaabf84fae30327ff08d71e
zdcc7d5a9db8983f1ba87b284bd1774118e9b8a5fb39b7c6b19078c8e35d1c77022410b5897f041
z7dca47c6e6964fbfa817f26dab6382c247993877149e440177648db51bdf078936813e60ae1e16
z8acef6ebc9de9a280d9e3a205f4a1a17ffcfcbc27e7bbc84a9410d5972cd57f64766df39d9373c
za2a47eb89bb8dc40261f9a25ae5c5dbc9c8407f25fe46d6c77f2a35173957de76e2d5f4240bf3e
z678db36f219b4d5c89aa899d111f4d4ef1d0681f41fda96d25c657bed9551e8cc722ced78b4b89
z507336904602306ec58518f1ed019777b5b5ca3c343d94260a1eec10abe79b8f69f5e1e07c0c4d
z532a2d9970fbf31a6b5c86914269fe2d2dc7f860fe437c00f8ea1a4c24b6ab3879570e3746b046
zad609b4d0351675abfca46077bf5593ba39d9a5318dffa605a2dbb35067a063e9a79fc446e2468
zb5ac81e6b9693713d50e0b7e4b1a01980982021d8b6a63f15a2ec48dbcd721fbce6e226b43a94e
z050d3cdaf710588322675cf62d94b1a37f6d4711b9e2f5dee8b83d1f0b49f79dc3a1926cc85640
z1b12e010d2128ecaa4ff6a84238f2c04c79008373ad1fd221b0b47eceb93e74f2973e97456ba2c
z5c5ef0f7ec17a4c00985b51a2c795c52ff3d069e29cfb64b8f58780afd7f17a46b6b960d3a22f5
zd1e52ae764054f432b944545346d494ee10bbe1a4cb9913048bdd15cdcbf93bd118418c6ec6f2c
zf526486c4eef38ca4d145d23ed222097460cefc6e7f4b97da8a9345cca456a41fd26db38641978
z21c7b8d802c394535b497581d9b263b2c9eda9b86d9d636ee7bd6433a60a097887ff4d1ee9d0c9
z2cbc940fe47adb87a10ef2e8088140526eb4d4dba70a1555cc00b4b45e4904b0150579d91cdf83
z1a743a4c0675e38764e6d89d810d92649b64849c0b68aadfd9a2cc1bf93d3a1a536715357de545
z271d17e320242d3003547d1d5b47ba000a5e5e83cfb97eb4fc2dbaf987f9a278a042ca6307739a
z8ada59aa34fb75e973c75fdb97d69184fc4dae5080995c57838bc8a9b3592b110ff178832f0388
z65b90d1cf09c6a629f42e76a22403a8ebbd867f5f3036102855687ebc94cae8f7ae8a5ef94ee04
z1a62635422c5a68576930d4c7915f98798a51bfe6e935752a3491bf32349e7d28de207b2f5ca14
zad3a7dfc69bbc8704d65e6c7f226bc60fc057be6aecf3faa6f3829a04f7f569eed4f9f2e1c235c
zefdbecc1de8ee47a5c14862a6f9ccd8b66077b822703f77947bc0b8c3b986e1acb88175246696d
zc786683df9ab81268f0b364c69ec07957ab4f88dde035af11064f5beac5c3771d0b45eb92895c9
z3e83997a70f58aed3905db316d56e464034ad2addaed31182f8b2e20096562f3e812d9a7815a73
zcbd27f1ff49b82730c24d94d912b7d1ce2cb818c2ec95e6b2d3c79ad9c7c7c7a0a6ef812ccb8bd
z2b173fb5ae79da87f4cffc3ad0e77a4fed787f8ddfbf51d4c1fb22faa6dc7820a8b75738f6d705
z8b917b3a8337e018e048961831210928acae9ab474dd83de0e14cfc6fdead0be85f05c0fa70cde
z7dc329073aaaa1a1f0cf536871a0ab58cc3ab8dc585bf92aaf26c821508a1ba4c45c435b877985
z055c0d68810e61f0cc7a4fd76df602adde019556aa990937fe13775856f49ecf0ea4a4e2a660df
z7478836903267c940b115142ad2282050ed0e2578465c111998637aaef25c1add695de125e8241
z13d8bc0debf9e2216c70ed99ce40fe46dbb30bac7a4ab2f9ac0a61447d70b09ebefe34bf2ffbf8
zf01f0b19e6d47ed8e2340e52bb236e22bd0ed3fb00f1e2624e46564af87729c6f388c90cae15dd
zcfad384c3a172ee451d408c635a64dc50de0771e8d8dee2b19c57c3b1d0ab25c9c60bd1f94de9e
z3e91042b06a2f4ba5b63468d49df048be3b1397408440eee35da90e15d9c976ec4c3b72f1e2f3f
z349267c59770c953899a52e6df0699c6314dee01dde213d2098a42d5d548bbd74cc52bd8c87a88
ze304155ad1394a461e19cafb1d32791c00e2144c9a30db676f55ffae6f1643b114a12b0a58e9b5
zc735818b7923fcac7d3dd1391b75fe3525a0744a9728ed6d4fb9440fdfdbf98f8c22c0b2eac5c7
z9559b2cc4bb1e5d5f05947d81fedd072cac284c3dd829be477e0e7f0fe1b22b8cd62c51c7e17fc
zfa689cfcded06e8f95fc63aaa56bc1e63b270de4ac3152fbc0a272c0a0490338965a824c792ce7
z5f8012b0c8e6e0b84ffe535b2345074d111f0f08564aaffd40bd8c087c60311b2aa1f94fab2c43
z37798b454cae44c6c49fd97af56c7aa9f393c13b6710be27b7ca61c34f9b92ed3d03cec34deba0
z915580a083276d18e517e6a039cbb6f16ed63549376778a0ec65ecb6a0b3376fd0a8274b31e9ba
z55c302fcce5bc91d5796b7d3c389c21b6c251c205657ef130a0ce91d70a606ed164b232c8f31ea
z1c504b02d4cecd78da0e8f80500293b3d1e64c1cdf4863b93eff87e8a10b411dd41c539b2cab2e
z75dc0128a2920dd5e152f8b0665ac67275d03c500eeb63f4ce2f4a5e72dd18af22822fb78fdc27
z03dd9f29aaeaec910ad7bfc2eedcb7803c6eb80b0f406a96c1470e3e787fd6ea2934422a1f8d77
z5b4561b471c4b6cae211d2d480f518449a6dff5c10adcb2d8b396c30947e0e97889464bef1709d
z0038402acc6e8bd63bf8df9d1c8c7d352c8ad097456524b7d645451be5a4222bdc2f1c9417da38
z7cb01263a5325fadf423502b5272d62009e19904e871d03eb95531afe87df1a927bed80e43f5a8
z85c7070cd5f27c180aa1243d24659a45e01676e0c7443a795df544d89f89369009835592f6ac56
zbd2e225a20ad4d542c2619c041a9f94d7b7420a6645ba42464b494dc1fe8799376d0e7623d67dc
z622c1a6850c42126adbf28c2349d071d22125decd2c3b257c4aca81445238c69a3e9e2405c42da
z903e2ef5ff8902f76d8f72b2a68d722c37b8a3fdae9be4b591bde1cc180a6e501c643e1c465166
za71ffe5204bb3b0275f7394068f3bf165d4328f0a4b3e7e68364b2f2f11d8604ec85891419de48
z6f68f9c9721dbf9f65a83044d9153462c66f9a77a9098ca67e653db539b43fc5668d28c62e25e9
zc9ce4f0a738cfbee84f08ed62a5e5c5ab294c965929218a9e92915be87a17d4a6f4c1b8cff4c40
zf9ea8aaac23c591fc0d33fd5af777fbac80df55124b522b01222f9d20bef77fcc8898970ee8d8b
z3beb1f27f0996682d3315fd58c38a8edd79697e22701bc7b6a7fc131f5d7d8e8f006782b1e7ad4
z7a03f1475c6c38b9b65520f83e29c8d6b13f7ee9f34841ae08e8f3b5f0a026576e72571c0e175b
z10b9302b545deb69853f42fdb9f51e03a91951b0714edd53e48cebf4cf48a026a12dd43b16895a
z337af0904946581fd40a9f138bbd20b6c001d48d562a80970c5a9803400a147e89ce0d7cfe134f
zb1851ae4c3f4d4ea984c623af760608bdf880a28fbe04028fed5283e628549e5c319ce0504ee2e
zec03022645b01958aca04e18e847dddec204e6fe3591868738aa30df66794c6d90b352513325e7
z8dc6011007ef08751232deb2d0c30a142dd42b00276cd4887f8e96933b16ce6090c3e197f4774f
zcc2490aef4c676a9ca48deb8200e827ee42f59757ccd261567091a2a0d102e6f3dc6775a142180
zca38ece00afab7139c467c6e510c4fad8c6d55056934e886b7c1757d05926d491a0c028a2f6e9b
z22d6c07aa0cd6ee934d89f64110cd2b580869971cdff0c6e648a80893357367fd9e996f4f8373a
z9a178690c8f41355c9a1cba8af2af8e25c35a01596e14d2f207e4d2f530a8ff271969f0cd1079a
z202ab8740834bdacb02ab513b9e7cbe1056af190e82de84b8ccce2bae234da818b07a74708991f
z555d84339ea1524a239c1f35b28744e4e7e3505dbf207e6b9e92d875a58232df6305d2cbfdac95
z048ae90e8548b2a4f62201aaa90df87925fbe66ef64296d6b4b447521ab3360d6f1398fa444aa3
z6a50f672a2f982d751a1a7286c335cacec27bed0c09dd64e89d4fb0b8f7899ab75894e6bb3c87c
z5f9c13e5c07e90c43413153edf447b2654fcf2de40f64611ef1d26d47911420bc0d9c745e5df2d
z34809e3e98ced4cf75f3f53b009893dff143c5e5f7c2da5ce580ce5e4b3e40aa0b2310828ddf6b
z7c74079c19a51825e04e5885b206c7ca2fcfb0d11ad29b30ad3a0de221294a967ee06b3a3294ae
ze711bf345b92b4add5db6e75eb2004da497afd226ec19ba7db2c069b9c268241b0253d5a3cd3e4
z5322d4b27708de9fa46571b69bdfcb5ac422a746e870c101e7ea954c3d182d4c11a0ad63836825
z8141879ec095ada417110fc8a169ee4e20e9f5fb62edbe79cde81ec22eeb4895ffb3f1af86fe2c
z5a1197fe1451f0a5867118149a177d4e262e56cad9f3e24380d202f8e51afc60847fc5397ed0a8
zcf0a409bcd823a3038959ec6d56ad906244c6763ad20ee5b15e97d054f38954db314b55e7202f5
z59b4f2f6fb6e4dcddd15509d66c0086c9c910ee31b6c5e13704bcd33cf18b5198591381d73c23d
z3ec9c099bcd290d5574f3cfa4130f69666d61ed5269fbf86757350385392b68d4ef88ef7931491
z1d5ebd7334be8d94ceb41c04e8139a7f8d1a5f9fb79839b38df0986469f9bec45de46be8644d14
z1c78a9b6518cd2ab317d22930e152f6d2ccafe902c7371d6fb425322f2b6ad5e8bd1406f96b72e
z32376ff131facbea7cdfeea7782de942b030a8d2f7c77f3cd14db370c3293112d9a65b566b790e
ze64954a2f7692c44d2e5c9a05a6799de729d2090bcd40cfc6fc9e64a53d65821a81bb920e6f075
z1e2b3aa40825216259aa024514a9d3d8c5edfbdec4abcab4a093d9a27d6e133997e0ac1c21bbf6
z8106e76a9d117b2f1d8d1312fa905b26b84f90f63ba0b329e19fff7db4124d49cad4bf1f9eba36
z5c59cef4c20a16f15a5d0b028f2577060ca6a36ffb0e085506c9c8ea57ce946dc67068831d105b
z474c971f3535ff300cd055f10592bbc03ba52c075bc7078a1fb85fc7c6d1e72def19b569272b41
z6a905c26820779b009755be2cff9510a10ff980c2631d71470e5b3eefe0106928e49fd2064fef3
z05190f27f9c726daa8db1e46e02ae3c946429a7f74c55790f6cd64593b49a400099b58673f6a20
zcc54dc93711e406929cfd78379c580bedf23b8dd8a1789be0bda0b246c089121c1c4f8803a6810
z74199cfb85230759b8c7e96ef8d3ac76d899f7b743accff1881b7ac4ca10ce32d26e7304d3947e
zb93c71ed080858b50f3a2e8d1e371001effff3de9dd5ffb4aa12d0ad7f170e91ae64a552ea0abe
z9dc0830bf1de103ddd10eb778ac50290b9a882b03012a09d015788344bbed176ece5b032dc322a
z46487d155f1e39155a781b859045d1f9d501650a9fa1fd64a1b5f92457d9b586ee9ec7db110012
z17a19c758c9aa4269321bb6c669370b89eabec185a9633c3c4d22bb95551b073275e8b7d4e4c37
zb060ea674279a590678ffd622501e52c94d4d278bac6f49b1a5028e5895baa3d1205b6aa99cbde
zc8f79010b82d5edcde201af1588e1e82798c500ff73159687cae9376db37453f089aeb940866d9
z0e4bd571a49d388251e9f81371257c86622a9910c49e5b24e070df3be84817b81b31d0bda30ba1
z81ce2f2e42b6c1ec7538e4b4fa6d2ae924015f04639fa21fac1e9b10f27ed504b1b507e88f697e
ze11a9beb8399aba94bd61b9bada4e0e4c9dcafa058fcd8962b1b92aaa3ca9ceb9e4673645c1bdd
zc63b4da8a148cfcc564c3ce76d2c33cb1c5c09994c4ebc09a3d90c179eb5960e12130f826784e2
z83116dfddb313df1d42d178829ed9637422bc8c2f05037692fac5817fb01d24122da711d642ddd
zc73bc1e8aa02ad1368752c9bd2c49f60d463553369214a581a798ac9dd2b6464c3ea79c842b7fd
zf669659978a5fb7b42de5a4ac1bf4a2fee43da98ca720ae54d830d3290cbc32aeba562f3cf7dc2
zbc5f212bb060dc715e65fa26d416d4f981dfdf9789f8ea16251435a08320825252da447351810f
zb6d743a53200ad7c7b20e9184bdf6a80d93d746452acfd2f380dabf416748cd9ee55c21e032ce5
za548425b81484585fb13949703cdff54b85fea166b8238bda47272d33214096efcae35d75aad66
z89e3a08afe7e3cb9c069d30605077b6370def92d1b2dbf3a6ed5519f1db7887dceb79489e94e09
z352781f2c6b448bcf59ca7f769d4f27cf8fd98dd60cf9da875f2e87ddb5ee620f69a60c2769c83
zbd974a47056ebc18551dd3da01c188123ae58197d26ae1f64f013bec6cac3ef0ddd83c86f8d26e
z0b6655dba682263620c4783dfed329761a2daa1ab451a05586f698a9baa26f1fbab0da5e0c7716
z868aeda76181258f2290eb1fc38842d64b29e800d5fb05f70d87f93f5809707f4bcc981bca9636
zfd309ec01a38fe3d1261cbe93c4c73f5d99bcddb3793eaecb938d5026b118f8da59aadc0ed45dd
z1fe442c499871164b53129893e9322a4a1a41e4f9cf35cdc60b67efdda4cd890d5e434dd1a5d03
z019eff62a984578c9291db53126206f37868916a4d1d9d8bea41e4feac0aef8d1d72d8033fb605
ze116d933bf10e708cd67dbb507a1444d588dc55c4c1ce8b6d73b44d4b41dbcfc03250a94357ba7
z9de513bb387930f160bb3173aa9b6b088cbb048840c9f54f22674cf4d79abff30f2c96576ed203
zf5e633126bb6d6231b3c7d259586f913f5bf7cc7b94580e51dd7a162b03fd8e4a66431fb09510a
z6b973e2fa778b55f256010d0d14af5a2aa09e89166f21bed4f36932dad3e9a7e7f6cdebc8c8026
z5155b48d25bd793d71dd5164fd77fdaccb62687b9a6400ef0994dec9707eaa6a8c823dfe196e66
z747d13a76291399ca23525aabca086520e6a2b95a92dab34bf744a6b1bccb541951b62d617e442
z459c6e2756a7175bb3e1fd407e065bf8006d9ac931a0bb430a89fdf2288aef507b67b99bba915a
z70bf39b63fcb018ce93ad877e0f1deb0e83457fb3f9ddcb1526608dbdbb4dcd54756a2d2f6910b
zcd1528d370d4391985d708f115f7891ddf75f8b419c53685abd837dfc60583a523f7febe4bd49c
zaaa3537c29c078c7b98aadcf62b783bb09705f424d667d391bd6490ee35dcc3741dc3fdf553fae
zb7275b72e5010b16ea73852c0f59dc368d55ac8561da16952a0e55a61554ef841597ceaf51c6f1
z90cd5157fc7fd7503ab2f804da8bf6f04a26e48f021877043dd2e5c31796258e25a2a9dfccc2a8
z5ffb46fa489ac0b483e91d3d6c3885eba975f5a3906073feb5fb54557b5a5304c9a0973e8a135c
z44ba832b4c2b2026382cadc35b97c18e6387a9a36fc8b5eccd4330b45ec86b22a9049b50a712aa
z81660afa100215d3e61bfb0b1b3ca3be0c622d8b2292461683dc5718280ebf848a02d7a169d7a9
za0069ed47d6e5630ff46a3b90dbc7a4cb07d6638c119846f1193488e73628dcea8c4d0e89a07fb
z69f7333f80664f5a6621fc7481a5731026a21929a71782d8cc815bba6f25f5ae34af9048761a23
z21eebf203dd7c547e577f5f6a4c4edb411865810ad84739334c7c209666db7543dfd9c31c954b8
z91d1d1472e1a73afc1bba7de4216d8e1d76e4e186ed59a3d98d40de31ac2f3bf808893d83e2d26
z69c834c070a4ae7033985b6b524619ea960ae993d985d34cbeb155f05a9a36dad6dc8c1ca0658c
z9d91913a937bf009e3fffcea52a5b1e41dcefdb30111b775fa2c6fee63048c8e8cb01a186bdbd7
z97a503b2e248314cf8583b81aaead0a198ec628d03ba484829c69b185918314d1ea6a058de6aba
z62b94d44c62b792ce6907bbb223ba1e122f3e59743c3115fc541c299b631a0365846381eb4d667
z0f6283075c1e2890315c9662646fdec5c935bd9773660abedf5c90b566f5e23d7d831ca54b6d61
z4fcf601c23c68343e8997ea95a53d3eddbf116f2d5cba4a79d541d6361d666d7c81564e24ad6f4
zc218b55e0e7cd2cab789ca852517d7744b51f9624633222e4c2655e64cb32c41308d62bc34f1a9
z4a53bc3bf19a14f6a07a9472794e7287e4f623a71dc72d9077f7354e07d3df880a4f35371aa5a2
zf26b5e2f6a3ce7882e789a2bad4310904542f2b2d426730ae9d075c92a0c0ce38b6450a05fb010
z13ad3c93294956e4c4246c1a141c74116293925914ba1f59c5ee116b759c1f2fe834a744fbf27c
z17b5200eb32a003928ed4f34316e24da8b6372a26432903ff5acf3efd418a5fea49067448d438f
ze942172b66c9ddc636264eeb9b28a61befa59fc9972f4e885e2165c4e7fe4b6d6d84b29a1887b4
z416b7c559182031b9413aa09172e060414a530fe7be302c6fd876c1dd9d451ba24526897c6fe22
zffd3b2c8266f4324fcea56b14ecff9a8f6f3b32530ebcd572d6cf0dbcb78722772714b26748528
zfbc2da18b66f5f489d63850326baf774821d665658d9a5c5fb6e7229dc97f5497075df708e62b3
ze6587791b84d227e2c1a992d2087ea99e372b8841ec3c60b56ec491a27202ca30df3439dab8d88
z5fb429ffa962f020fed1fadfb3511a54d83078d82462fa6b584a41b0eda3dffcdc11b153120a3d
z303e91cb0d9e064fae867524eed5d75c56995678d4d04f062f8bc3737bcba26ace475f5bcdd314
zbb93c1310e2fd9bd80a3cd94a5a1e03fe4e4e4a5a9eb9cb9ce7dd3bafad6f0ace9d158de08b68a
z0cbde229f5b36109e379085339f017cd8cd8ab3b3cc5541a5002286a6ad24742747ba7f25b6a2e
z1373d7d95daa6ef3a48f0d5276ff4fa33b7764f8eccfd44d0b83faf08bbe514b9b5c66138687cf
z8927d669e06aafd67b358b47d7c5f47ff4559ee304cc0ee820704094c91a7503c7cd4b4ab6f0e8
z6427da2748c7dd921cecb0de9594c58871358979ae49b950d5608687fa136bc121d568378147e7
z737de56081cb53d2674debc15d6ff8c95310a4ca91694e418ca1335b37d3ee501661d3ce3cd45a
z1978a8ceffaf8897117dec475d87584f34c3161ed521065fe5cefde258d160da9c1142285ac098
zc042b8e1d13e2456ef1ac26a10b72277fcc4e5d5410a34ac5da449940b2c43923bb61b04bbd1bd
z3a1425853f883881d946792beb3f2a55ec13ecb24c4672ae7be6a7fe0b6b75085bf7fa0b8acbe2
z591e3bc4f8d524510ae67ed8f185498ec38feb35ebe25d3e69f39bc4112d3355297c9fe6d4e914
z9a27dbe47390dcba391129bef7f3be856e6ab774775e70aab00c27d9de6cfd33a14337be18547b
zcc2daf4d548f3fdd81e57358ba34418675c193deae88821a09172893b73f38be58ab6c97348439
z7e2ab5a4b0b1cf48e24190179ade49e224e489600fafff48b117e6fa3e158dbc292d6e29dfe01c
zdeaeca31b79e54cdb8c5c5ab3c81ea1b58d580dce36a575b9d991ae21da07c787a6874570f0e27
z310c6bc709adf778ef0b71f0017657f1b1e4bb0626eb17c8ad06b07a4374dc8dc5d8ba32dd7822
zca44a62430c019553e56ce1705e855bc3bdb5bb8d14a43af55b13c06cd05c4fea884a3cb3cc2f9
z77ead2313389df6d5bf4f958a050d277c4adf4c98ed04c4f791a29449e72b96623717c202d5b15
z07e52fbf1bfc7af562c4a6b492e7197a6d106e1f57a8e357a742c3c769c4a27acd652ba2725850
z727051ac9816889e411283ebef1e6c3c82a1b70cf89e128cb86ac45703baa0d367341555c89c27
z30cc7e77a4520821b08946c79df6db232101c0239a7c1bf0953094bb345d201ca41cda941e3ee9
z1ca96e66f6ceb7f4e2c048dd54569492d326c4fc817b6f5cc60e518464bc4430f9ea8477efb95e
z41821e8bb28eb7eb175567bb56eba18dba234986d98c411fa510fc5e4387778a7f10de03a3d8d7
z7b2ca13825d34cb96739d7bb5b9dc7e49cd1f4eee6aa1f2db6f61f1be582fa8377bc94e7d8111e
z2413bad8b5147e50e915ee733a6bba21df1cfbba7367f3fc4bd621fc1b15e96706c480d942deb0
zad3da72bb5611096ca7b950b459ce726b3cc41ae901769de3b7d1c9f80b4057abf3f3d6dc54e97
za42afd14fee9e1b376c4ecf79c45bcf50906b145046077cefeff6238d4fb0864a43e0bb71ba57f
zce4e4e80e03ccbdff916dfb51d92f25734459e61061dd5fa580250ad21e069003742939ef749f4
zecc0838dc2ce71eadba67d37898d621d20a6d57ee120509cd33f7d8eddf28998cb9ee1a1236436
z19d76dc38ca00a85e49be3eccbe86c1a1c998475f0de7fd1ae541083951fa50bbf05de829aec56
z7961dfa309a9bb317021b7ed9e5dfc2e273143425f6042027d7618fbd31575a5c71509c0dcf188
zc72a453f672f76d87fb9c0b89ca715fe4be027c8c5cf8c909b19be70232fae3879aaf6e4155c25
zb67dec210a75a9ee4f0c85a43bf23fe4de1c762c61ceab7cd0bce1e143d71c5b120e490c23d649
zc27f3fbb74e0776b86df0cf88943266a7952068a1dad4ad8e8efcc3785cf5a3e244067e7e23259
zec5ee5e5e3520db8a147954b6fe234c5ec30d2b08355ddc2d3954c7e8260b1ce4b44bf971d6182
zc07feaff4579ec224f9406ff8b218198e0819a9fc7d0e035abc884994b0c502f841890bfb6750e
z1c1198d4a8b180a927e3851e8b496aa7084ed660ab2cabc2e36ef1a609fb2b034eebef3cd92fbe
z98f4a3ddc99ed4fd4104f0e436765f321769af7bdd53676ce4781f649e1d052390037184092b87
z427476e339a4f47aac3a3a3fa19eac56ec71e08fff7878e90edf8be732f4397771287595dabe3c
zbb71c6512cf2134e7a998007542dcebf9f96dc3e0a48e4549354eafedddb3e5336b2305657dcfa
z98edb5bfd0639c8e7832914b912d9af4d03951a96fa36ed02143295be374236babde07536b96eb
zfcd67ec38da1802ad27bab727ec9b537961495c0ce46d472c768975f1176d7297f3a7b3def8b0b
z010aaad164627f379c6ec2b67b19cfc7de7fc436b37c9d20343e1070d42ec59c10fc9bab3b475d
zfe436979e13c469ae432291745739f7a846488462ddbfc2f295f815f3d89706c2b4f19d596c715
zaf0fd2bf280fd4c382f37ad3104ec1630f3fb703c882e3cfbb8abe918c78e79c6ceac5d97d152e
z89f076886e86e3ac85e6ead6d9751e525a8a00bc77e735cca4c4fddbcd41c68b19bea5d48db3c9
z90dc6979be6c9d4869c5e6e7d8ffac63a1254489e45987ba78ef4ffa4a1debb8c62e8c3c538f8f
z78d58c79cf3ef5a0f8c87efee7663488e810171b6494c56aa65a67f656381d776da3ae219b1608
z645118d03e9d44cef9d4f31f9dd873388cfa4a360d8b4b50eacbadca8bc0f783a240df834dc406
z080c87fb447560eb889aeeaa2e97b11df46ec095111c8a3d66abe452ee6696047d375cdde7c698
z70ade10603f2cf29ed704464cc8da50eb570a8f5279e02ae792663d3135ad40258088dbcfaef01
z28ec3515d4bb792ba9d5feec827356e61e1bed0c699b554fc4f16a44c33b1c4a45b817abc32923
z33ccbc473ba1a879700be9d19930283fe79f494762c10f16af154b6359b098e916342f61561303
z6a67c90eda1825d501c807dc93b04e5df29566446efa2149fd777063432b6dbd165cb2bb284019
z3bfa15c3799910f68ad2af3f433ddd87c53534e7ed51bfd28ac417d97ca66cc0a658503a0dd20f
z6eb33693ab197259ea116bcadae07ae99c8a04856d153df2e0162dfc7df90fbe48d52b7afba69b
zd683eae453a430f0abd8a804a3a83ba1153643ada08b865a34b2f6870f93bd07442a7f941073eb
z1d6703c19c83258f7586a5f23dd90c0fb88a6081b3d444f69f0bab5b7e436b60ccd95a49a74113
z8c711f7c1795bcb5ff9bc52260e2b13302f8ae5ff966aa55b961ca3d7e6b3d3f90f236b4a4ab28
z74b53d824eb107c2fd565e992788fa8b9a8fc93c80c2d77bbd4c9dd4a45618baf153889e4b681b
z48f94866da1c557bf37b59cada029550fbc292e4cd6a23beee94179f8065e564479cf6e0837dca
zaa6f1615e9f824c97f5997c2b122f9e0da50c2062ea634dca3b2eb1a4e693517cbc5c843fa6992
zc816bdde0d27afe964248e2ab95fcba06914a5a3c29a8741bc5e937dfd957e5d01ab61e33b6013
zcd2ac3909c2ee7ce786d106e91f8dacef02303afda9189cc313d7f9cebc284d9d5a409920c697e
z8bfd8902792163424d04bf9f0173c1ee8a64ba02008020af6ea2823a8838ff4b9e02e195faac95
z19ff784186e0510033daef861b889cfba3e0ec76544f7d513ea7fd2b004d311addbdf4e4218452
zc17a7f993ffa69cfb79d7b3761abe5b8c5913ea91ec1258c103b4b8c010932d430323ff619ce35
zac5f53f59151d6b1d17b0824a5b2cffc1dbadc1dc43798a62053e83d0da218f73136cb559b4cc1
zf6e843f123a5d037fb9d6fc2af04be162b7cbaa30113ea2c79292a92b6c5c70859cd85364bd624
z23925473ed864fb66a36ba7d49f6c6c95f64c2f7ef5d2a6b2cbcb8c7d70b2b9d10328560af1b36
z05eee1de3fa130eaadff7d08ea7cc129c3aca1980d18bc39cdfdc64c7d566140a74629fee2e896
za12ab0fb86a500a17ee76dd4dfe487621f4cd61af5dd66083f6c570675f26a7b4f273f8587e560
z1a6775452e1645f0368ac789f694a0a9419749a890851e221726905f341154b0a56df7fe795a60
z030cfdf826edf5b4c82f4839ca83ebfa10ffec3d4f1f3f952821e022c59b43311d3dceb85e2729
z82a5e4462244df8684e9d94466c7fb8e1696280af2dde8e104735cab83d3c2e9f16b5b12e76c74
ze1f0bdd607d0365b2db3384befe03ecc748520f5e6ccf55c72c9f1b26a17732974e935fcb2dbc7
z06b76af149861c5071c662f6df54750f682517e16c61dd483ffc5e8ddf6a3c45ec12607128b1ce
z74c77e03d57e6937e2c153aa8ce1390344997eebd2fd9b23f46c49a4b5368c151144009d364a9d
z0e3ae3f38571e8e3d43fc0d963470d66ef7c9d694171f1394bf90c4395a9e1c9a0c2d837cbefc8
z367c350f8f5110b4b791a78a311e2d8d83413762b1d354d74bb71f3dcfa67b49e7899aee15a31c
z4c88172e0d783669eec7221c99a9bc5becee282486e8adf107cbdfc012def83504b0643c99ef5e
z8c00fb769046007ef3d7f4ba3279a97622b3dee4bfa634f94ffa544c2a26a23fd965f0a6f260b0
z469b4b634408066f3bf70dd71df92bbe3b943d268d750f11608d366fbf7104674350fbf462c9de
z1a228ddc2a26284b4c5c69f2d6905b073ed9c718e06f831490af349f00850aae4c7f1fdeedd928
z9ef1b28ee389df9d6caf1ec32891b11fad488d841694d3efb90dab9900cac133c974e82083b66b
z90b4c96eb4d7c9ff2c03d407972b8eaf271d7294cd4ed99af1b14a822f7632b09e75b71a4f2a62
z45ecf115ec8d9fde6782328d501dc556b643ffb0bd597d4147888bd44f8e2c572a86260e2749d9
zca103bcdb7056758b6b10f97e3540c44407c2215a98a0701a1df66b1221fd87d304d89d2bb4d83
zcd5b2857b72e9cc70ddfbd44def9bdad0ca850741a9b906f138ee2a5f44452b6a01edb12b1deb0
z5cae64cc38177c866b942e88e8cf60bdfc5b07cddbe84a64c4bd16b4429ed02a34c283b8d21008
z8a244e3c51e23970b14453ac20d4afdbd028b4e3f001e77c77e188ba65e0334ce9934cda443f53
z72a55977f9f2159d2addbfcc26ff4d5128df931b39acb6c7ce42807e31f4c2c18ec001644d5c6f
z896a875d0fcf8415d51b46f0fab81dd9a2d9da4d2637f2b9c7ecfc6fbfb168e1a5788dfefa39e2
z09bc3f54dd6ee59544e125a506d5159f719310a28eb01dab72d25c6c84a6127bffe89f60144834
z02b3eeb05c6e3895834e11eb01f42cd959bc0c780311eb9530cd5cb1f8545da08980f3c769d5dd
z7151d41d32b8c5cb8b24450cc7a5e9c5a2855b33eb9f82f38ec70b716ba61899590e4c810771a4
zca37e23f3e67724eedbf385f2dbbf1ceb472cb96b4c60db11951479014473b046c404189b21de1
z1c923fd942abff0f1da2181c3c279ac87a35e62119caa7655e297f7877ecab9f93d64526ff4ddd
z64a1254a2d2625a3002f2bdc625a0cd3135cc3e555b9aef76f16b009f827f48f312a84cb16f212
z98b6ac0f385fdd020e29f7f0513ea9cd1ea9bf4036c1f90063f125883231902d76ad005691cc6e
zb6285f585d10f443e613ab188444ec29071b54c9efcbe638793bd55a0731cde9295b66927bbb2d
z7876b68f8c4f713f44dff855604ca6e052ee02e30479cddc5f4968709bd65c0b570e0757629517
z626a9d594881ef82998d58591bb9205787207fc4bee4f2ec3ea983377c849921e99b9f5f36bf69
za68c893807bb70367999112ffbf18d7259a2dfa430678313ca7d326b5a8db465e761ee1a326dc3
zb50b59a47e362bc218722b38928a7d2dc83e558948b64467a5556d33f2729fca687e4e6d041412
z25cc3a8760ff8b409d49cee362596bdfb8442643d61073de4eb984e7d528eb3cf489bc4d383b0c
zb665e30b1ff744784619f3d670b346542b39652f255e7e20be287d099b87ab300d252b99ceb1ee
z36a50267813f2227b7c9325ff2d5bfac91ce48301bd31c464d08ce5d9e863f381063940ef273d7
z65da6d797dac6ccad2f210764cc0e0f8b569934b63a7df8116a2003907649cdcec7887256bbcea
z222f2508f857623cf849112e0d58cea5624104d630e803096869681f1e53107923effc3d73b231
zce7fceb27b3935034434a0a4b2a789a70ddbce1f80a2511b17e4bfc58cf541201b418c19c276f1
zf912036208d97ccc3218f2655dab3d7b7f60ffc2972de46e46dcbdc6abca0a5f78153e156c97ba
z808dcb50b4f2070da1856069bf56edd830cb9260d7a848776b7637f860ba931ea88b49e4ccb2a6
za20e713eb293c5144e8576b7584afc6ed9014ef47f2a2d41d23c66c02b06afb647b893ca715eab
z2ec2cca699c49bda642e0cdc871e934fbe064a78d553c604b8ca039c7253601866c3286d0c8c0f
z7ec461ab9a33fe6321ddc1f563234652f251d6467cb56806154b3947e49ef9df76afe0ad537a39
z4f0959ae2c642008110f9d4daed2e962d6b08d0ffeedacd4fb3a97e13b61685ffe5738087b35ab
z990eea8aea1451f9e13fb6668075fb66f89b4dcf0250863169bc4f60d201a0c252f6f79f903979
ze9b974ff00d8a9e89aef45bf245da6b70a879e96aeed0ee9a96582914711050a00a5bd8ff70c59
zf8fe204f59d760cfed14f1e2cd868b65810da4cac42499a331aa4d6376ed5dfd7f17f588ea763d
z8974cc745a2ac9e1cb887373b45bd6dc5548d5910b18454d0db6c56c5ae2c76abf010c28f5a24c
z90caa820e12a24a0de258b8203278475776ab0bd0af8c31b4506a07355351e95e4a316e94cfb12
z16bb7c3fe0e1d41324e3b4c4d08392be07c83129e1e4fb9ec309cff4203c59f1f8c6c58137c175
z798b804083ec56b505de9b6b35f74280bb5e58b02db217cb271f5688106b7c77ed96a59e8e49b9
zfc0924254679e4c686da29c18efa5802cd7660a359dfe2906dce1070d0db47b210e8d977a44d6c
ze7ed43e5146b6146dd6ecb93cad04982100a9dfc81d66a5dd49767d0b62fb7f4a610f9ddd4c7f9
zf75254174c604bf142a8727ae9259266d759624e2006cf92f059c9f60f5d3d9e6cb3c0c5365b8d
zda7ddaa475fc6ca136c8f934e858945881f526da1867b3cf5dbac7dfec537221c9ca62f65af17e
zf60771f4024248a1e80ddec13ca6c7def985fdf1e48bcaf033d0ac4163396288ea227b061673d4
zcf2a51375068266d0c4985f96b9266c27a517377b1f92c6d34490f9771348dad85d219bb13f496
z59f098fe76b5aab6603b74460d3823930fd4e33c8aa0c21fa1b90521b75a645591cea242f1252b
zddd0853174f1d3ba1ba08469e6152caa091d624a7624bb7207374590ccefbb86c3da2ea1eb5610
za57773e36828ad0ed4adf253c7491c5a32832862a2866ed2ba864b24403714c3d44851b21ea45c
zd0595e9a5b29ad9741ec56a69ea87a02a67a334ed4cba37297843a91481b3d4c614471c6e5c8a4
z0c65a8d5fca8eb2e6898688742092cf6cbf72ee1909f82e47ccaa5f1b6e92a388182fbbc73bd56
z0f9951a8058aaada5f5e2a5f28137caa0e933b5a869033b3018d37c4ad22e4cf2cad88c37c8971
zeb32c63bb81172ea5dbda9988c2231f7ae2bf826ad19dfb94376b80b4a6370f071630bfc4d67e1
zbe1d3171704f9be0e6c2599d0e8d10a42e5d7ad5f980e1f0d92b8a2f89e4ab22479488282d7f79
z86fa78e8b13f365dd841f93d5e6901edb814f177017cf17efdc51553be02bab769fdf647c27cf1
z8f53c229fd9e7304ddd12a012c9fd25117af36c523260093a10096e6c54bf38cf85a6f9a4bc570
z8b348107f752b221b45722de41930532a77ef729286b3216b982d3b1c637045929f791ef8b477d
zfcc07246c51d8c1bcef3a8bd2ba8f9723143e11038f892e638a89667fb661325275701a4fbdd92
zecb90e907c6b3dba837c186f60938ba8e91d774262722bd15ea7da226124c769c79f705ba428bc
z148f8c8877a652e67e22776fa175fb8f47bbf92fc719345b51ba1a5ccba25a36bcb328fb1ca76b
za970ce8a94ce2b6387df567414dbf2d945f19f0399edaf6cbc4dd8f23eaccfcf2448c5189528c3
z5295c19372d8b8b00981557fbdbb1876638be036ca690e1cb1ebb635fc2530af59c77fa43e966b
z3038a6a92c263b1aa9141499408d39022c4c4e4bb5517f251f8f6b406c264a2db6eb0f57a12ac0
z861c3f8fc1d4c5a477ee647f3aaae081fbba5f10fdc82c442b0b683bccb5844c9ff1f4e1804def
z3d47b6edf0ee34cdd195d3086df7261672441196694d77d34d23405453a7b75585f203a336aeb4
zeecdc3769d5eb3d7088e8f4d6c20ebe2bc803d42309101a4a425afd0dc2739afc6813f5c5fe461
zad094300be550e8daf177780f89bbb09afeeccea3e069102fe6c6ffa02580dd526a763a6849a11
z2b414e1775d574149241436aef08b4006bed5b14b47c355718b012b1af629f1258151f6d36ca04
zf1b0869c3ea1bdde2d85a1d98d85457add9266ec05e4e0004b11581f87f0aab232da428607eff6
z5c547e273fd0ae45d598ca324e154fab12dc11d3c209b09d4611c499de3f457a968d3c1aabd5b8
z1c90d5353468866a976d9b7da8e8c183660a1128e97656a0ab8e41fa748ef63a8856f508988f46
za6c6ad9085a1dd5f00f37b6348c9e854e44af81b03a4934c8c7cb25471a1bdd6a6b8a717c88fae
z3689244d4b05b8407c923568a31436d3cc32339391ac6ff98c8181a2fef21a1e7722d0f030bd58
z687577536cdf596ab1ebeab18d3f58c01460379a834b7f42399be4e5701a4e90aab778c5ddb2e6
zd8448a40dbb2947b4b5ece7dab4725b8b1201199c1a17284228c598d751f6f8cf5f5d231cdaddb
z2a66fe8757018551976d524a9d9695f849ab4afafa930d2c940fdbe9d0b9a2730f488d08c84b33
zcc94d497f08cc5741aece45132fac3cb2c04a82051d99bf182b2280200bee3af2f1aa8173577cb
z88940f43f968ae4d922d018c7291cad32a3a96344f4687d88be3cd8419cded1239391cf8d820b2
ze806c5dc9fead05981e6d45ade76a776072415ff0783ab827daa1ac924524a58a9ff94c7f131fa
za271a540aad9824e48e87a385cbfcebb5925287c4e5401dd9ff075a0bbc56f02a98f924c37dcdf
z1343142982dde60f931ae508bf4e3f98337e238515fdf21f822aad78a2fb68a34b0e9e06fb9256
z9f99ca96d2db8557a7bf9f0964ce02a2e6b7fa0f84e6427f055983e782b2db3263b46c762c6e49
zb4bbc548165259cd86128e294ac35be874f0687bd1b13c13d02bdc85becec6d2a5ffb4df794392
z23ea5bd6ccdac2c2209aafe7bbb35aa5ccf6e1e78205c46faf5c06279210cb9cddb4d61ac788db
zda6e6450810992aa324b7a8ddc527de2fd74bf39fd54ad54d8997cd36e0cf9cc9b5d0101c41424
z9406fed0d4b7a146a4982b151c7597fdcc3a4b4307bb92e3c525fd439eae71f424dd7c01e37f6c
z9397a13bb145c92e708bf386c84ed61da5b5e4e72570403ae7331d8641a19887bb33e7f7b6bdf3
zc714f72f609a56f5c7c15f9641815411948e262294b2bfd6d3c7a88a11af40a63f75fa5ab380cc
z1c258b414795e3bc0d7da3590968f1584ba0edcc714d30bba52727c3b02c0150fc7546167105c9
zfcb76ef424dd71c5778d8836595acb67db7e32b1edc1a87a11fabdd1c863034d80d81fa9bac9c0
za6e7a5994a33c09ea2a854b64ee811877960771cd0fe2a166fa20a0e275e5411c4e0a23cbdb454
z70bc39e7493736e41da0330a50d3aed76530be7d35aefc096483ea12b3ba1485d3a9ae1dda92a8
zc6fa192001378029c3101acd6dafc96db4b5b2cf591e37ca5a653fb8b33bbea6ac66c1e7f38b15
z0f556393565b797da4b27939d909b626521e714e50259d84a4ea539183cce92e1938d582fd7e12
z4d6549024542065bb78c3d36f0c2dede6b5bd1e898f216e55aa4ce66c66dfee0c2cc244671598b
z14e4c5012f88e217c78744ce0af2e56d0c9dfa0b2b45008e91ac4c75a6f0698e3dd8d5974dca96
z2c9efbd240f19c83ebc0be1f4f491428fd9850f37f882534758c6325d614d7ebebaeda768d39a2
z9530fbb35363808220af2c328298f7a72ff4c0deb837682e422df8b3d2b6df7b564950b16db9cc
z0f02c21ff6ba035b02c990d613619dc22efc46338272b378ed6d39aefb90ee56ba751f96bb62f4
z03ee9114a7a305f7d856a0b4a3c056d1e228ba4765d14765242c2b0cc1fcedc823be9b2cb7dd4c
z9f06b080475e717d4f1afc392c91b9a156f9f6d9830a374a3c4d69be18238253bfeafd2b878c21
z675b10e27ba7c635989b140d4503f5e0c48b422a547f5669d925d03bd467a86bf29bfcdb5e7444
z50c5adbd6dcd900b10b20cf9a70dfe1c7686b8ddb3afe8f61023897b828867cb10cdd9c2faed83
za33a251e29457a7afb4f78f6eed83861b28ed858c733266aa8e1e37fc4b02f921cb5cf78f214d7
z1c90b1317ce52f80bcc328db1ca272c737c86da5c2fb09ebfbd7b4ea128941ec85ebb977071e79
z59b49749dc939ebb2a5de5c20cea8b403cc9dea5b0aa6a513c27ff9f3042108ef59d4d6948faaa
z3a5140a4c65ae63c8df339f93a7fe46f06171b2924fd2ba7244c5bbdb4a6fa196bd43fe6bf1c58
ze5bc5b3f1b960ffd6bd0ad52ae3e0078c6e7581e231138e072b97387eda2b3f7dfd0ddf79f4f27
z630bc2583f32270b246ffc0eb4c33bd883794b9c18e6ba8f2ff82bd7d80a96ba3d0d46a2a6269a
zdc06913c76ee85e9848ba68f0fc4dc6788bf9b0f9eebfcf0e5ebf09f352761bdaa353bf7303d1d
za1e50b27abc13ca4695d1d88abdd57c5b383c911efee6b9a1e02405706c4f048dc351175ab9637
z7d1f4f5a3fa0786d45e8c58610db6192ed436e37329103c84daf1330567c0596c11ac596008993
z0183e1462745e18ce34781f67e76fa01cc21a38777144f22117aae98164cd1e7047db39b155d2a
z228747548259bb33ac7f604dbfc23f0e2141ef289a03b16b45704704ef0cf8811e7e9d3672b4ad
z53472b720a83d2d8e285f07cafa952ce690c45c4a585cf0c66449d0452622b090bc0a436e19626
zfd5773555fae5c9159534e5453905bb1ccc193211fad828b3ae83225c86f9edccaff6bbb57bcfc
zef8df9058eb863dc31532b1f406a59866cd59230bd252427be9c62ddbda0b1eafce5a8665f3ec1
z31b22902ed0dc8b965f3b0bc64e98e8a09cf62340e1e32763e6e7bbf2812344c57e0f093442843
zb983526724546233b9b2c8c372600366e294bf9752703cfc19ae3901c993c12f45b4e122963995
z66a6f3c7dcc3abcc2d16dae3a42c3675dc56fe8918a6f84bc34aea160ecb5efcd6b201369c374b
zb6c5ab297ee50871f3700c096be7757793c1fe8854e886d29be17f81ac0c06c27a97bd58d082a8
zf41312317be543066c25a058fb7e03a66bfd84e4a506bc01d877060caa723258741c0a44496e9d
zc36c44c153791ce94f2df37a200da5f284b4527a072ac7f2dd1c64da989b45b13acfaa9c446285
z101d68e4405457fac11f4768373ba3665c2eae4a8e64eca1b63969e5abae3a64308da8fc08c35a
z2f48c8fb65524f0dbc3d0d5595e7d2898195b82ad7688825b7012d74662767038077b05a322d97
zd4d5954b43f90893cd8efbc0f8fcdfa1bf394531dc31176c450412061d8f2a3e2c3bc818758747
z35b4d7bc4e4026a3bc2c002521e9d2578d84f4dd008451cb77db3c4d9882a5c5cccdef3ea855c5
z770e0adb7aea1fd47e1bd11fd45a886c5899d368b4b37a7205cb7704c57eb4f5540473045fc69c
z88f65b3a7feee78f1935a6a30212c2cca48ea6e14536b2fc7c193a65bf3aa422a266e5922c5929
zc2d8c7529166d40b051d3af2d57b21dd875b4d77bc4300b113acfd5a9be0c466ce6ff2e6ca883e
z063d74060429cb4420c4f9f7e80a15b977d470e8d5e763504663e495145dbe3845eedbacbe2f4c
zd509bc22ce2bac30a09dd096cc102b8a9f9c4ef076f3ebada481629526cb8daed45b96112ba8a4
z44bc336619359665f53cc9833e4849362b645ccdb2a9e32668fbdee3a66c124146c2de0fb437f8
z28c4d791ee2aa23dfa4a6920ddbc7c4ea3448068bf852125270a75bf7e83c67e647eaced8a20b6
z7677b028bc9bb616fd5a1a1d50a81dae1760abb5fb010696736913594f7938341607f5b424a57a
z90b451dd4be2a57339393d28ad3c23cb8db51b0e754849fa45c419b002de4b9b0aa76764a0a706
z90510c36073e661def8e50168a655c85f2893a1351cbec762cdea000c0b41e86e7b3b1f3ea348c
z8d681acccef261b444c88f3656f86efcc606b647eb90b157fac72361ddb16f68d394227367694d
z47d1a8bdf779f2c663a30afb42ce3f3ff32f1ff5c034d81a756931d3e77bdbac6309b741d96ec5
z5b436d01fb3df22df83b433da77cdc11bd503f5ac27a54a93c4936cefd4c289b321078c16e1365
z17e9b4a5f0b9d0442e2a9971fbf1712f8feede80c487368ab1412e531203d7084c409d7eba82f7
zac035c7695f1863351ce50acbeda5da0895e5cbd7ac94f04da3f66cb651c7fc87dc7dc0d5250dd
zbc483a81e75a8c8bcd1c302d8fdca5cbd6ef70e7626914878fa3e9d2c4e05f916f7247fe452768
z63be40c0a9ae2d7e9a4432d1395e72eb8be7152111b8557a4be0743325c45db3fbffedfd37993f
zc2dfe7faff177fd593d7f104e1119f46b0f5a92b14244684050984d768adb45c9c7270e735e8fd
zcc56cedfbec932822f8b01882e613cbd2aeaedcb248e829f755cb89c1cdf39b25e74c6f9751718
zf8540a963b0bd817dc5b6ebfabbbd60f8806cd99f62d005296482ed8140c0dace97b8f17a070d5
z7856ed5fc35a670c6102378c319a1ca57f3eb0182d1c6795ef8c95662046d74a86606162594e7f
z837b9fdf6e0da7411213b1cc9050f5527034c4ed6d3f664f7459c35b4724c394e821e27c41d1a3
z54523923882dd752f41dbb10442fd743aca831b3bca29a940da985bcdece4001ce51f3f9d837a8
zad2fc68d204ac5b5eff1f3df4d50b9d90e53e72d210c9697c0c9d9542754bef7bb847860e3cb3c
zc633c6ed0bd34e0b6a59bfff3b882cb69947d37e57495b2b1fa29608ddfe9de82a9ec1e5f8c9c0
z44ef26e0b9ae222735a130783f6e4b4633fd8be87314e794ecd7a0dd2e2875af25e2ace5db7809
zcf274a67fb7c7cb37e8a895a8db30b3acb2557306a971550ff53ccad608ea52d23a2bfaa9e5e75
zfcba713e944cf2ee8cffdced7cca9204563b3a194993a44f4e02a2ffee258841db37af4b887054
zc514a34ee6115f4b33c898d070e7f15fb6beaf750e845cf8cd73d7eaf0651e78db40316d15def9
z52aac4b58845546016204b5cbbcc9b15974c7c425c140646667062b24d9b575d2b3a99a56e8490
zd0d7c8880bda8270b904d8ad73d7684b0c93f2290cfa114b638e42dbda7be4ae1ad1d3994989a6
zdbed2411eaf141893f619d12196ca8a364b9d8dcc01f7a70628642df4652e1e0679d7bea930371
z85b7088691731b4b5020c5b05452568561bb1154aa7dcf9a7eee2f026e12fd2531f65c8e40767d
z3c270a8b0aca32266554e2a99747dfa9555bffa1e9ad878c76334eb591755006508fb43920a7ed
z192f375fe7ba1b939513970c28f5a31299961a0d248329656385dc9196c2cb084a107ac54b34bf
zb498357139fda1dacfce30fc071355b900e1ba8891ed40e29790f5787abecfcb3f94956ff3f956
zc004e239e90354948391efcc92389718f6940391cc661ba664009ca5a509b82a88dea1d940b334
zb92429cfe070816f39a1fd6b16324447aba08af128e49af903046a29bd587987bca190142c6272
zd42f27dd59027690447977c70b5d921a4bb994d1bb6de08300868fc5c7d27ae57de03a9c666e4f
z2057b46a7ff89da349a99d840caa3b1941adab795d503ae3b329ac49ca6b4ecf4937abc0ac55b7
z9b5837515da9cb54b956d981ed913ee26048c465162279e11a7c1b2b5c802e8c50e7444cf50288
zca65f56f34241e29a3de8ce9dc1ea02d8f1583c739e6d3dd9821d6bd8d451efac8ef4784d978dc
zb8b6ede94a6462f0db5baf52751954a566583e83d967e3776ec169f2a75aa9435f6ccd10d7d5f3
z8a1ee435843b1a3fa7078edb1416db8bc2501c9e307cc3ce92a5a7e226fcb26312eb75120dc30d
za477b5fb547f839c56c743b9cd1e8b3108d33bf1aa4b099aa7b70083a27526763b8fb9d8429376
z96af37089b428e6d3d56f68788dc65cd6d2b6c7bce1e09e3509c81f150d30375f323659d4760a0
z42879fdeea1403a2a39c10af2d77a1d96923ccf389166cd8cd1fb97dcc399a844c14ce908c47eb
z3027675ce2e44c7bfbaec6ed10a0e66047eb8bed33ef7d34aac0a56d1b4478a8d61da469301d58
z3ba4d3d4df64e76957d211f1f91cf12a42ae91675c70561459228b5d57b8dfc4e0c960f0f322fd
z41cd38606cbd338af4b1ad5f72319ce5591d916be602b66f2a097978be6ec904e627e6b3913df3
z39e5a6eeb8799d0dc486bede2ae951182067e9193a87f9d0a9129a1b7fde18dd4c8d71418c6faa
z742b5714888597331b9f62ca72fa0738343f9a0805835e004f2f9a73144b11172c536412451e1a
z2bb77e0b1532b7d0030620dd8a858167f5267958a41f870e994aad2408f99a86c807935f1218f2
zdc5c081eff683a0dae9f74e894e02ab8a3d7a445d5446737971eed0c092fde62f0b740eb73651c
z85a1829786d92f72942f075efffc191ff0c6808367467d3a9d3f19366b5fbeb346ba6d53846779
z685e3aa7da294461b10cf34d261cab63ef5fe4a44bef84e441e5962c69735dfb7bcb9bff718e87
zd531a550c2af17cf04e0d17ee46f62d4a269b2407d9cf2b1640cc9655ed822a314e7fd6cd88309
z49f90cc3a7687237110db23afdc0f49262d72ed8f9b7959b52d754e04c7747b19a6f6d744c1c3a
z05ae7aab540c02409df3085b23cbae247dc76b9b37865c2e8cb6070f9e25ff591bf5d77b41196c
z0144af0e77105b09ed8e0c65a39c027a76d6a7806ca70ebb40d2c1213fe32cbd8fc152bf75f813
zb289b62a8a64fea9fb982829e2aefe82901a23cc0d6bc2184686fec4ccfb3f69ac1ab37ed04d5a
z740099ecb23f270d20fb2cc2f61a193a50c10567ef31f01617987bd2f6817ab44b30a30883cd4a
zb06cabac02ff463d6d91738b4a4502b5e57b670bd8da51c64a1aef55ba89b344a746827a497205
z1819faf7c7930bfc60ea92127d1ac8e6254b6eb929a697b4cf508f2af8a60b22b751c1350eaec6
z29d1267ab89d9e5e8daa4fa71a957799d01a2d2c50baeea7385aa3b68f413a1b4a0f7872dea417
z4b9c454fb2998f8b103f58f329d8bca2b0c2895ffab57e9074b2d88d6437b0d80c6ce18c42f8b9
z7e575b3ad26f8fe346ef73ff773a5f8c995ecf92c3c51e7a0fd7b3b0e13c0b6c2dfed7b80148d5
ze70e9dd0a44c489eabdc42161530972e5f96da3f5f4ce948f1b6d89b9735bb55a99f7d2ac3e47c
z3a4cd0084c9dd41beaac6f7399d61f366f6c06f6d7cf0f0b77f436cf02c3504b53c8a6f4673561
zf8c3328c0bf6b5c0879dac1edb39ee9904bc571e24cc55a7ed1c6911799e996e76262ed0d5d875
z9d2be1f54e3f494bb16368a377b073faa24070488b22fe56977290d24bef714712e87caebe8a09
z6689f4747b4a7d94b31d5d34ca0a8538314ff972a4f8a860807aeaa3dd82d1c637629d5479786f
z8f56cfc7ef11db97a7f87e55804962e97507378e50554d66a976a1d47b11cde292a007fff4cc06
z8b79d390f8a970f7c8225f8f22bb2aa12d618460b0e205c1a1d52775b69150cce547d6f65b5cea
za1312db72e690a2b160ac14c717e499406d546876339aff86cbd756d1372d0b6a65afafa56af7f
z9d876367a3d7863f5c2ee91ffe3057bd638103317d992be0b60bec91ee5a9d92d3b42917adc505
z1589b3bb0463efef43eb376e69da1c49c3e48410344bca6bcd066ba6339d73b879d2dd42c81bec
zbd432879d2bda86b8246b64db395462b3274a5c30397a00c0496901cc681fc6b5745acc469a1b7
zd88c107eddd823fbd04f118ef034373e31415e302e3e9220eb8f3588eca547de278dfc64196fb2
z77825dbaead7fa06d31d4692b2e539cb69d12a80fa3fa766b20e5000fa21ddcd239405c850b166
z3860d703df89cc983daaa11accf6e0c5b9e5a029eb8d8af6906c02c9e6340ce1fdac1470d80459
z19490d1e158119fd3f218142387a9749155273eabca66e9fa771a577c5cb1623b2230925c2544f
zb5f5809bb03a6536c43320d3c8623d9ccf73e25aa492c6479345c8601fe9e72760b3e01e81074b
z149b1724bbf0972c91fefb4e8f0221054535deb0b2b22a7fcb4dd23225990b1d8d2aeea2f1094b
z4edfb42f55796256cd998a41ebbcd23d4639861db5e22b06547cf828dc32a6e5eb5c6fb114b569
z0b3ca615cdf458cf9dd1b7dec2384116ebf0184aedbe0a6b406a47aa19ea7af3f98d643f96a088
zf56dcd38078a03dbce863ab6008ecda4a761dbfaca0d98376f3de7a7f3194f6dc246e40e3ab3c6
zeceedd9c8884991364d3cdb1da1e25a265022f0330772a6dd2026e6d33c5aa085f243b979e9e64
z0f2bbead2a07225de52b23a22a73fd96a34add8cd1ea155964f60efcae4a3f7ff7f134f2610e34
z57b0f252a140e45fc51fe5363c52915a7ade6b8e05a0ca9bb67de6be96a4b2a27f2130b206fb66
z0667ce5b20a5dfb872556b31edf8bdbb7d53717c5edb6c4f5cd2297e3c199b1af6f9481828856d
z6000cb39f87fdb82640db9e8fc613ceba9927d427840279a10478c1b06903325e3b9275fea9f40
z23cc435e377db42ceb4652f56180da8d97b4600967158789c3046cb40a834f16b22d4cc65eb133
z920a75c79ad9e66d6bfdf562282f1664a15342f9248fc6eb793d14bd01c347a4caabeb5315fb9d
z1685e2ec8deec85f89c6412a1b98840e79457bb48c87b3b2003912d034b234a45d70aa4d75f0f1
z45a7d504ae85d227f151a422289129efd4c7b4cc0d14cda62b574c6de27ed8a20a03abb603007c
zc63a0bd78ff5d69505f64f3b7798843379ecca0a2ab8509d30277bf8c786b66a505ba36921ef0a
zacd66aaa877444e91bbebfe702cfdff9c301b77341086e86c7c28a9cbe54d62eb80150605b8718
z181807bf9e33dbdaac7f0eacc276f8d29bd479790f550267946a338b947806317f9dc0c31f6609
z2d51ac50cc6ad376766ff2c8fcd6aa4bc5b6aaefbd97007cf52ac246e2faf5d40bd5d6b20e92da
z411a4bfbe912d0f6872c4b3acbccfc137abd5503202235c6edf1248a97a3cbd1a09116d31746db
zec55c3cdd4c06e0067be169a42fba4474a92923e439d71e0fec6852ba3c3c624a85ecf5e2cf8f3
zdf4fe49d4752097126f51883c8aa371fba141e0ca18b07bd56919ff71c08e66a94ae7aae5930b6
z4b3d8c00d13269147191f148abbac8c94b3382e8c9d6882f08ee98efcaf43865bebe618193deea
z398f7cd250fea3c6c5f2cdd06445a53f0aca1f2c08bf1924523489c5805c47258622dbc87ffcab
zd14343607e388da8697ae47b80ee959702b18c704dd1f963a05b4855dfeda12a7aebfbca1b38d4
z71e961144d39366c3be26df3f1063cfc0f4d07e53fb71dc5b32dc755445ff4752c64121840a6d4
ze1ac54f4538c6562acb3da6363f7101e09064036c7517aea4ab06e121c5943644139ad097f035f
zdbec9bfeb7acaddf1d54a952dad660de05742c0ec1cf33ceae06a5ad3462589463ad18fed27e55
z7b13a3b58735321b8c5eda71a94ec133e0f4bf41a3ca44ae27c5572bfabddd95ce892e667cb573
z2deb5252088c2f9f2d7aec5db80e6e527ef52985022bf509caf09a030c9732c54a650360f50245
z930ba4a62d9c6c09364d83cb57552b787b33f797dd0d448452b1a11754383646e9612bf22dd8d7
z088ea34746c3e35342583002d03488b40607242ff2b41a5e62310643db75843594f96977201cef
z1288c1351c56952ab7a4cfb9fe0dd778824d70c35b1ced493f9de8f6999bef9983a4d0f0e20dd9
za9e8d14636d06da12032d519882de02a04fddb8fdd4e74c62151951e0248b97e4274d7e6247701
z25e7cfb499402020b147c82db8766775f70658d46c5aa1a6d9937aee2ce14ba0d21c2411776e57
z750f6b050877ee36b5126297b94de5cd541dd0fba8a7c204e034fd1ea09f1faa22384997be3cde
z059058898ddf228905ab8117bc0044a6edbe849282452eed31c69ad44192965ad783f6f7ad3ee9
zb3cd66922711384b71c4b843be0791ed339400013fa7b742b1246ce913bff27d977cf21b1798d0
z1258b4e7840fe8791874c126e16c88f22c5da86b34cd5ac47917ae461b0a758ff4f18511536d45
zc9a6a663a3af2ebe34ff2174a4dc57f11e4c830304904f6a4f49abf5df7ad848f3a1ba9bd6a11d
z2a39cf90b7e16a56d70de16f549f327538c05cb187348fb2d2cf11dc19397932fc914888322c1c
z93947e331c46ad7b2322502c8721bb4066906b4064f83265fd4b2de65daff2a19912c7b046d0c8
z5364d545c65b4e5a1365db9da77778a16ea2d23f5f8dbaa027cbc6d9433dfb56d8fe64d580dbc8
za9527e70e7d6282cc9075efd5461c83d950f0ebdf9831be2100f57b70f509b17e1cc44eb1deeeb
z7e69ca1ef94caf2cf96e89ad263a018b58813893c43953017d62f1b078de48da188b364ef4cf80
z6add57c72d35796e71831334b2637c00155cbb9faf67c4712361be380eaac45685dc64060e5026
zd65183d7f8530c67688c5b648651a7d23882663d753e533d25936aecf117e8159319c1d38c13b4
zf866d5dece64a949e33f502e735c40aef64fe18eae3eeda1f9729fa75db2623c00af410decc1bb
zb9b02d5a5f4f63c91afb04aaf08887cb4aa9a66164fd9763c28550e426ab40ad3c48e5bdb8d3f6
z9c83a73bb39061e45b007420de7974ba14f1f6c986c13fa22822a9eba004d521db70184f3016cd
z2ea2ec2ae06b559eb6a473abef2e3ee0a9752232a3e4768f2e5656b56bf51beab55d2a87bd2a7b
z720db300cac15e924638d184a4cc13ecef30bc39f5724b99569a7ea27a030c616d40204cc71ad7
z66e583f51f5b2d0da9d09fd81172962624fbeabd2a74b98b3fe0b9cae8c7fbbcf4ef9fe000f9de
z81205279459f481ff2951bbaddf10cbabdeafd8a4e39d6646fb7590fc7c82ab6a1c4616608a59e
z9d0f2eb348d708691974a07c172aff55b692b1677b387717f4850670019f57d40102a84ccefc92
z31c119d41867210ea3b99d0bfdc2615732fc595fb9a46e04501dff94c3a595cd58aeb0c504aa49
z24ae4b82b9141882df2590fa273904e386523e42be6d61656bdd33216393e044132f46d4e82c4d
z09fa73c27f87ba3f36016e17b7430360ec5a42e96eae81b70dc8beb0e05b79be9be5c7344ec7fa
z1f64589bec9de58c79b487b42ee073522bce383f08e5f020104e31746c26659b005173ce5215c8
z920fecf76f6147c5d81888949cdc0da57afbe8fbd9f8ed33b5ae7a0ecf4f3b57cfd5bf5ba2e756
z919c74bdfae46cfaf04cd196ccabf229c28df9798d425da28b7a6610c6baf355dbf2ca0490b701
zdddec83b758346c635f8d2f1fbd450c9f6fabd2005e1b6119d007d528894c387609c392174f42c
z24d528e812f4c3bfe0db88ab689b160c0a7133ff25a29583b16ac8de4f5069f480add4dfc81bb4
zbce2ebc98bdaaebf805700832637a28f4b6cba4d46dee984d9e9b279ae4d87e74a1fccf903fb72
zb3ac1518ea058610d8679139766590742199271db72b89c8123f81488eca68b6a11941e8379220
zaf54b92ba645810f63a61ccb06028d9a136323f340a033af93e896f9e73634005232dd337f0c9e
z20772cd237876b0bdfc5d3e84f05128f268ed1382b6bd7ebce9e712a80efffb45095ef56d7d75a
z4fa349f2b777bffe8e3ee076a9f07534ae090baf27aae2d1923c3365497a74a35288a1d0a17c7e
z7190770046d9a51f131868dfa05e3f21f1ee28aa005156166afb4281914cac6687622c708da02d
za914ccbdd4f512cf606c9933117fa5f3c6f339a3ede532815b6f33da3fcb33d8995b9a80845f02
zdb814e780ca77050a7018f37a935ae46e18904bfd87f597911c0260af843873569860cdcf2149a
z6bffe32019ecf35a376aeb7000d874cf8ed835e3ec796c3a1b8a0f63a197e8ef8ada126960336c
z1f8eec49fbfd7b2c235d18a5d24f9b8c2c061f2867f56adee4f87954b1b6fdfd8b0ab665a281ca
z0b262cd99b0611d94c2596bd453afb2061f15dd1ae17d7e703648a2afafa7a369151de0639eb02
z5338c43bbce6d52d97c3bcabbbff56d63c0e3291eff8ca6ba36ed25218747af1bf0949d0f74999
z94a9e5021f3a82d8f9b135a0791528fb154db197bde4eb9bc67459643f931f61d8f76a166bda1d
z82cab8f6765b16d2ade7f0ba305c1a4a0af81e88cf4beb24b655b6a6354318bba6849575ab2b9d
ze099960c2345ac48ca66a517adaed27acb78d8a6f3a510db4710e04d3905ea14a6ee02b8b4ed31
z07565e2b2536bc1145efcf9b60cc181fdad3aabf7e94f91b509aa73e200ce1b28d22847c50f242
z6ed429887f9372b32bf98771fff25e6f8f90e11d55403f29937bbe9b27954ef8e988cd40a23968
z0b1f2358c5fd8d42f4e47ccb40aedf91303cd5fc6f83880827a285fa84d8c40ce25139dee5e0b6
za3974bc9531df78d2a30bc907b0a9d9456e0fcc5460cbd128c40e3a6be9a6b2a941bb990d4f84f
z41c390b70a95e2ac94205b7dfc9ae763e45624f62ba3b26e1aaef834abe2a815dcf0c46f874dbd
zfd0cce4025877b452416c18981a5e73a86947d6cbac7dc302fe0db53ea003f417f66d11b6f841c
ze279e4f35ff98db855741a13f2ae0f0f4448507cb27fb3b65efbbd30142e6dc50c27ffde779c71
zc9e30af8bdc9e2e6e7becf1c30c31a812d6e3e714644a13c4719d782ef21a9e5ebad6a42c83e00
z26015666b4690bb3e7d4490b0334f5dc802ed90312a637e05390e84deeabed3d74a62301633a32
ze18aa7a3ad68512590fbadb16e31fc92ced44a933b6ee7c8c6fec68f7c9fd4b94a49238e7cca67
z1032c6531026dd405052ea690e85843b23505f33a33f85e27ae5da88890fe9cf901cc09a0f1584
z7063a62ed966b4e1b4303685e70c9004465935cd228cbbe412c0c70375e5cf8a8ceebba0ec061b
z1f051a1c221c33b71a6861299f9c6f4e2f359142d6fcf51056c3b9f07fd06eb04199bed9ea67d8
z9f3a0b15cacf3d88f3b1d7454e79841a31876b536fb0b9cc1da7512c7fe68b83f5f2d6ba581b84
z04f7599a56a7e0848834472284d20defc698deb1b36a975ef329afd962086b94c9caae18c949ab
z167bf601506a86ad923d6318a8665b7ab26e6bcd0701ca4310ce15d6e6dc910f896816a02ab5bf
zef840f3e30be885be3a1970f4d33122aedcfb1622b3ae08e87ad79c5d9b3c185bc308fa6066f90
zc51480100998008d89fee72adc4143fd73cad18d84b17286d7b68c3bc879fcc522ffe14d31f060
z62a1df7cf75275c6b7966befd55d59311bd484e3d3db165603adc6f21e8ce0eb29ac5146398694
z64db73455f0375b91021a824e6114cbbe237079a742293e923564d6e9f661f3ebdd89f9442b279
zca3b973396bf99818606afe52b6d87382cb88003e617bcbd4e7cc5193539a30ebf4f621248a095
zd6d247da6aec36f8797ce3a4c0561e0047011fb4a5d1ed5993452e450abf759db4c500584cf4f4
zb0eb589bf2dc2e9a1a554325c4e2d436c835ff23be73884de7a0a2047c4c226a4102e6b026e7dd
zbf48a25cf0933f47c575f5f55e506e1a3ea9f17f8f4878aa1eefb4b648e0e8d8bd8ca879d22426
z76ac43c2739e58d63c958bfbb336d7be3566b61523bee8158411dee0de45be244a507f2187b7e6
zec82887ac631fec72b36394d4cbaaa4130ee9992b9083b9d3f36bd079c26b8d6ab38f2cc6385da
z63652d54a394c34514162f1281a817c67b9f2ff4b4ba8034aa276738040a2f18a736907ddd25c5
z4ab94aa018e8eb344966c7e82b429426b1c1472dc178eefa3e6b660b579fc207a3856abf96ea88
z9d61d8c26bf21624d62999b12d1427a55df14a2f777317ee2bbdad9b890ba8ae26c04e8efe629d
z381662edfd52b148762486d39661c28da5a9bebd1ec2b153686e87785589bd1302a7143b604a94
z9631163b01b912d3142468ee35a4caa3f4bd0c52f6c80528245ab6eac9d31cd0f0a3a2a670620a
z62aa39ad4a53f9024f8a0ade6401aa690ac7b9b33578ce9c88c784c4b369c94396c4cf6793fb60
z58d0fea6e7060e9640eb35efec6eb2f4bd28592207468a24e426383b834e66ba28972c143e9e26
z70424232baf73b0537135be255b0bf86308fcf663a87019304138069becf3be7ac5edfbe3bf57c
zcfb99c2867e3456bb2608da8d9c5d07bfe81ea78e8f5a69aacb69beba90299051977e6c8833b1d
zb748eba7c723e9e47a49af43f23a4ea92f742427825b63ff80ff0694605b3929aca92713c8cd7d
zf93f612f25a8ec431d5567f2e9e2684124915e297121b8566f2b1a2b4933a700d156d58bcd0bf9
zde97d3a8918be4689ed25b859be0e37148f406bd75a2307825fc91fccfce628dea456360569305
za3005de7d7118b999478a1047ca22584e2e179d357be71716d1cb394c50f04d2007bd63c8f3626
z9619df7ea6f49992ff463527c4a5cd1893c893babc24c7514aed78034680d5001c00d0bf7bb43f
z1e27caf5a72357e459c482fff7a9bfa36210d5ffb802cf689364e40a5d23058f8183d5561980d6
z874ff33c385382371c02eac9a771852351c681d81761fbf20c70e6a66af4f5472e8105317f94f3
zfcefcc59ea8766f7400e30dd27727488d1d42f10c924ce5fc9abbbdba17cf41bcf4604f021e7c9
z06d5b91e781952266f9b12f18c784c7e5df4a1c75a63ae75ae6c06c52ef1003452a8e27bd75c24
z0d0c166b7ed6318c42dc30e300e8b790a788c5999d0c2627147f8ee5541cc15d110b393e414268
z7d66c61ab9b932af3b6d31f95afa9a868247d042be936a008268d0e9a630f44fabb7434187a29d
z99def21b0ab1c148160a443cd86c3e0dbf5c8e35ac3635e00f104c2424511df305db6b7944ba57
z97e829e966c44a6011a055ba9c0718e9e671897e57a322f52681b9e59c86446503a6a9b1de2fe2
z0c6f7d2f277ab670ed65ac9d42fcc329175e2e0dc695b4000a56e349b729c35417599e1808fe50
zeb903eadf86ac564ea93897645fbcf2f2f7b390ba901ac97426ca92c226dc551dd2b4a229ccfef
z4713db2ba9d070a5ae59f9b3338526a33b1c20abc1031934b1423a8f1e5c26ca8240f0238cba09
zc4bc326cc1d6a4fd918375b02a8f4929f82156e3385dd75821fc84a59596650b37efba9dc8c84b
zd6bf66ed380e1e016e710860f4413e8f30e9f8d0df8d899fff77aeb120ebf52613cf5226c57691
z9833959d7064d2b1cc64ea99c4421e7c25b8a6ee26da832d7cb0f55aced73361f5d36b34bb8e46
zaf1cfa9df507615a8341cd4f607be2d36e447ae38f71955c59bf67e7950d078941ba4b1d3b62c7
z7c44ba0db29071a501fc4e0bcafe868ce8f0fafbd18045c782fc1e27f5f2eadc28f14d37bd00c4
zf9e1eb456d0110967ee72e7994ed10adaaaa6dad8dfabcf835a4f639d869458b4b00cd30fcfba0
zd81ac8665807724dc84d08e926aed99382e2fb74cf504e2b4dc674fd67d7410effece3e8000f08
z5d4ddb1f8e22eccd133e0cf02bfbee97fc38fefb07cc4351c27f760049b8c7ca1ab8dcc4e34fc3
z48d659b28ac1d7ab826db07b5689d527a78788ff4506f548705bf79295221aa3e68586e8f636ee
z36ccb4d25010780a4e831edfb421f989f5342abf56cc405a7276093c2981bd95491cd3f31ccc5f
zf41547fce2b9d789e56a0edfbb76818b7bdbf961140c893f89721e5460847ee72e5ca72eaa48d4
z3eeac3f724d924ac75517e3f56d7b919f32be319e1db2fc86b5c23b01bd2529cac23016980577e
z5036882107c3d17a17116b5f25b2321fe6e2285afc8c5fe29b565f738c44119608cca7788e66f2
z5926ce24f4894c4f8e7d703b5273c5a155a7a29b3cbbbf1254c3ee13e1c939f82454046f1bd5f6
z1422ffe91b702436ed4b16d16365c583b58a82e7a9b4b8dc5203720469393e7d04a1b70250936b
z11d3b0503e68a7a2c123b06abe206f8bdfad357b628220d9140a03cead11bc24637054162ee101
z56a234250b8bc343fd90b0d5949e66fa2cc26e047ffe62db14da2cda5a6e82c4b578513fc2318a
z0259e3a33bd55b6e62f66d67136bbb9ef202a9524d1a101cdf97936d34636150395babd5f21450
z1b5f4e37655532c78e85e8ab786b16be94e5e7c88aba53ce72c663f4bb7d4a7a8390b8e7790078
z4b3d7a0ff0bd0e29c00ee64d44596de061a959cf8a94c590351f074bad5cedc5d851fec86d0fb8
z4e8c0b91416e0ceaf03017a16c2864821a287ea269777c7acefb34443507764fe95b1ec05339c6
z2d04ee576ecd9d2b20f19efa8ca7ba155e46bee0e89978c0af82b68eeea4f58a7563e562008f4e
zea9a4bf1541ccb8db1400a7e216ae40aa87312d6c683550aaa021af0fdc8a1383aa32dc863002b
zea93b9208bab0fa7b03380d4e9f3d5c535672e8f1293379b8137b58cf525f3b82c0766a5252148
z9528e5f5d084c0ea54c2817650311f3c45e99fb84e8b7c2fb3563b0ffa55e282db3d3c28457c31
z93e5dfbca935b20e45b6a0332a81921b042e7eb8d7e0ba6412c64f68c9b4998e8c835838834f64
z793875dd90e981f7eac9fbc77a139cbc01db82a5042eb4ae80eb322d10dc3e5bbcf77cd85972b7
z59784d566c5a10985cf3ef1dc5f9d3e17d149a3f61c7eea4711a6726ad66092b9d79a0270617f2
z78cd7bd5867acfb3205df4239cba8aa107dd2d5c91c3f048048f188e07132c68ed9987d583b28a
z0c3da6bc483b9ca91897a72abc2b7781b0c40402b71c3352bb35c9adc3befab6d957007904d8f0
za42e42cf14e1a2c4e9f6d33933007db5841a62e1da40184d45027a555562567d9f5f5d204d2934
z2e32bc1edf7459998eaf4c44adde6111f0ae76da78dd6e3e5f3f2eb165b3d563c21a2d5b13c815
zdc38a043abeff4e11a58548582e9df0a3273060ebc497e9a36f69f0b3e4582bffa5bdfbe956ef8
za64e9e34f7b7fa674e9b89e7374de9f89b7b1e9082c5b56725c8326d7bc42b62bf033a667d9be5
z17f1e1182da9503f272398ef7784af8ac2d85755d177a7e13e76146d91a0a880faefb5ccf6a9a9
z7cd23065d67d96f5a361e7bc1265522216fdb7f89f6d254f0659414994add4f60489c25ba54cc2
z172ef2d2923b4c29007b2d851aa1ca0f165ffe34353503e2f26f47f8348f7ac967dfa8f3cf4bab
zc2d16b1cd092a9b8217343f4309d0b05e3ae0b6d1aa395c82f243747ce22537bf311828c8984c6
zafa2fdea16d9cc85130a89c36c9609937daf9d51f1162ccd67761b4e8249529237adadd87c5d69
z1244dfc1a48e5b0ef180151aaf37e316bf652b29a1301d7c7154ebda0a76d32cdefcb3994b6bdf
z7478f10a3f23a678a1dbc16d204b1a8b4cfd62fb21d745dce59d73d34d77df6fbf38578e2af95a
z0c731f0612302ec1f8511cae8a90fddd5d63ca083638b2c1df43abb69ea3b449c0d249ef691728
z280b3e2fc3efc7c2309ee4335fb314cbcb778f84b46e89e43e4d8ab5e721eebba4e231607f6aa0
z0f914e052dae59e32ce1762717b55b828091e609a039558081b918f19e2f417529351972fa9758
zdd708778c5408c80a38b13a3e02dcf8f57433fdffbc76cd18d9031725cc77093482aa6051a6323
z6d741e9b4ac00e9dbb4fdc088e5c4adfa357203ba56d14ad823982ce8a2b657772788015e6ffe0
z489714d4845f9677a305da28ec059356acc40a295f9e8a6d704b60131d19afa3478fb28c0246b3
z8844f77ef91d9b7436bbca9275b171493d074b2a890556cd84c553b2c7abc4917b7f415ccd6086
zc655990f2fc71187dcc586334835f6d08da5f13a85ba559ad7d96acab5681296dfd036607d2bde
z0ae25bf61c72c6f20942b0e8b25f078cb53afd7a356406b1275b2d206158e3c0b8be6f99a07b73
zb18f9dbea312ae43344a94ebdd72c7f47eda8bf6fc7bdb5850cef8992e0434d530bd9568f1250d
z8b07fe5bf6d268b67958161fc0d2f9424e8ee551c7d9f8f4a308e68b265db02bb33771f2e01afa
zdccad58fc4706647c3515ab4ca0b2fb1640f5131bf61963cf25e7f3e31aae341d6772d13ba0a0b
z5e1dab9aed401625a4c790ab9aa7e183bb20cc0b47df7cfc1da571be95169220b69bec60c88cf1
z624b19fe85783f167fe612d32c8dcc83576b987efbc7cc669dac0a2556a6fb7363e04a802b58d0
ze15445e226ba39da17a24a1fb0f24030f6996199c44d3987c0cf7c149502e72302fa6aea9f0601
z4bb3b985b8cd623f69c213f2953d6ce1467e234903cbc58aa2ebd5829ed109706bf4da189d4c1c
z6c04cb48e2c33163c36e0de209288836413372e96c0f67fedbccf8ce1d9fe5beede84d2e30badc
ze7f2eadd0c1bcd3a1f4b300195e5184b73ea61e24b98166b4e0e728f4f7042130be418c9519f34
zb67a3d79e281addc39957ace05dc68d748449da6e096069d3c846e896789e582cf1c03f3c2e97f
zc563c9e7e33b51672f8ac2974b6aa46a437aaeaf60964452f16b6ff50610b5681241c99043dd83
z2d06aac03428e385340648dfec7d4e2b5a6070feaa3b84d440d5f980ddb39b6a9e78d9ce61edd6
z9b10667221b63fc8071215c171eb468c589454c551d7b168d5cbd54262d53e12dc8332df5081a0
z5f6f0301b0820eb9fef34d9e903942bec5c2cd027e2fbf064377e6baeadbc6d788d029a1e0581b
za30411b15034548ffd2ca2c64fcb34b3cb304ce51e3bed7002ca5fcf6f5e1121c62479d3a50284
z1078dd64fae91f10147cbe707439c511bb8084f5717d7de8b0ad8ac05ac7a214b83314d11498bf
z60af208f2298e39642178fa2d85592d3e814f322408aa0f435208714df4c6d5fc4cb3dfc771978
z47a5d77463807f514096d6efe4f0a6b65feb9f5369b03f3d6ba026e5d6a1b9480106b7797bc65d
zebef167daeca6d981d0069bdb6a26e37ab7259d42d617a0bce8f2c01f5537cac74343b7468fd90
z7ddc30265caf910d6e41b869c73ff52fe112018348f875b705d4a8cfec2b4c0348f31fa57f22e8
z5f784bbb1030d24883379d9a84b97c02ca81997b3ed15f29d0665ebbf8b2082ac53de2e5220dcb
z19f6ed58c8e30b2cbd1a428d408fd77203a151aa7fb18f98537a928cc23bcf5d703754b2a34a51
zf5f929015184c7c78a5be08eaacdc9bfb5829c273d4be4c69a509d88db31a75031dea04d5b46a7
z7f9c07d8113fbb5129ba027e9e338abb6e0206cf700b96d1685ba61f585626238b0b3bf556a59f
zb7811e30d1302c46e6f685408a357633ed620989961a7863196c856a3afe6c8974fa9e10a7112a
z7df650b8d581072edcd74cf0bae63189640d3ceb0b9e32c46276de0601e4aa942fc29b5cc9da44
zf0993337fe50fc9b775f3faec1758c889c1ecf8a0c42abe89f0cd3ed0246e91c6825547b3e9f0d
zcdf4c165bd42082bcd5ca656be5492b29c3f6f5c8b695580435f1ce95659da3c25b4161feebeaa
zbbf4638ede20bb9e6b55b0d1185cfb755442cdbd471c0ab08f876c975336030548726b9d55bc26
z17cc342a1bd188e24f5d8c684fa627d2eeb1e86377dc6017763f3ebd8e6af7e09827c88a6505d3
zf150433ab290be8b7ec77350bb4be97c4ba60c2d80f7e8b077dc0bcd5c5f90c046471a87900e40
z16bb0efae06c7fd4d48eaab3bd6cf70777d16a73bf89f32e1f9511503cf60629d0ccbe37e5f1b2
z2f0a0aadc442c2e2ea5bd9d3e5c9c12b3b946c3a679f487d2eb03bb461d0c79d9508a17697dfdd
z0368f2cace704c02e7f7b55c12444211148f9422b7aac4096ab7f22c33cb51c57dc00ce46bd4a4
zc65a5b7ced092a0e97c7cfb00c9feea6192bb1e52235ccc0a433db9db45fb1d28c65600e274cea
za08f49ae228fca1bfde08790140e88b07a5fa36363204e48799cae9bcc52dbb3f7c6066f0d4160
z4e9134800198fa437d21b6c3842734e14c15874e884eca2de161dc5deb68559e2a190455a86c27
z02fee7fa980327c0bd18a0e85b2b1771357955fa6c4c1337be3971878df0560093cb30cd9908de
zeccf2918866307d2d28edbf5653d1a3f7c98f7f8a28d25898fd78b2b8b71c74cc591f7f1df928a
z97176feeacee3cd50c611d1644c118521cc3a682f01797ce87ec621d5daa4e4474161d8a13093c
zefd253ad7bdd0c6008607323a558e1ab841d3ad40c98f277256d904923cf4c54643c28cf4373df
z27526b5df1aa7e971123229ad73314c3d7ede20a11fb0d85c79e5c6b9460f6724103123d103161
zf50053af911c53bdd84bbebe8236ab941b4c6861d5318b6bbeb3e8932248e00f4b2ebfa5bbe734
z4a9337ce53bf58b15dbfd4a83cd3b4587a5d46dedac5c8304187a93392e74c74b94f2f631181bd
z0593f6022616feccde2b463aa696b176b1a0eb1b031c2ecbb7024277859895ae3967e93a4f1580
z4ff49e8cea899251c57e73b55e0ef52eed2f2d0690c85640160e3bb0971ab20d600355d0a8ceca
zd793e2f68f232f8a2b0a700b1a4435349e06e24acaa6451eeb6c949293a0bc353ca7f4381e0ef0
z4aa8fdf7c1981608e89b562e8c8bbe3e9576bd4fc8749b6ec8a2842f4d38f5b896783950e9a98b
z9a3e2bcb040bb08aaf03ca2bffa17e89d9f578e5e84b40a802f141b61aeefc5d1434de12e8167d
z1baeb8ceca5c419fa7c1885650ef8db100a4e6503c4d5a79aea47ab356d2f6ae724d64f2b0ca9b
zb136ac00bcc76fb51daa337cf49e3ad05fd7a35c2a3623bd24abb8adc7b9f1f560e993895dda5d
z1301b3cf60a82c5e4fbfea41fe1aae479e034ebd774470ca2e55b056dfb9c4b4c9a972c3ab55de
z904c3a15cab003eeb7ce48b2c15dce544b37b08c7ce406c01f7dd6b071043b6a8da15016c03514
z29d05834eb6ab8b32614cf1b9e4432fc1d59b3ec88424c98f1ddccad6998b1e6bcc9d0b3376db4
zd76e89a40b327443d8bb67c5d1f5dfb70ac6416038e2544c85570339dec0913066ec4d172abaa0
z6f38bfc16da230a290691a4a925361ed98124ef7ed0898f976e92b88ef320174cf19fa46d16139
zd8007519b673c3a48e55fd5ffd1d1750034b2476f1d05a108c6801e48a2627fa1d12bd35da81a7
z154a059b5d6b28e568748c5f62c04e88f4752783cad26279b2485dc6e6745fa94a956134d98491
z045d06a6b74bbce53ead48344114a0cd243cf1d995d081fcbf5cb4644c3f42ff7dfe6ef5cfe957
zc9e1b81e5a5299bbc56c64720806fda808074eee1278316cc6cc64c1c36624041c266e64b270b8
zf6523e1481b175b5011c34bc65e6ee0745b9f45a2de72ac2d0d0587cabce874cf728ebb6e7134d
z31dea16b8b502a9b99f34d733678655fd5826b695a9f6dc620d32c23b31483c5531fa127674aaa
zd94176a355e0956a5f071c25eabdee22512db803fd33886596d6f55a5f52e00136ca5b9559b296
z468c170af38af39e1766be28d8e1af746f3b8ce22a56da18b302206de2c584cbc3794ccd414aaf
z0e6672a872140843adfb65fd28b0aaf0dac986a9672f047f4784a5e24d532e3c8c7b0a1f1b1334
zf90133f8b58ccc1dfaa2f5ea3710354ad8809dc785c26ffac1075fe2d7751563487748c10218c7
z7ca872e36f9a147cb074b8bdccd3f6995df83ad19ec089981a96988c6d1354c1a7fef7ee64ddca
zc943fb267ae48ae5a9d0a45aa31a9b98a3e1da07cd63dab73b10552fa4a52cc683d264ff8afbd4
z917fc5945c4a3b8cfdefd96a32a96fb2417d09def9399ce2e43b7dba70067beb316a8259e96d0d
z0be5485c45ef9a6ab417daea192fc77873dbdb7b663b7c2d8431d718ea05eb7d856cc258c1325d
z200b3f13466beac7d08e6edc029dbd5ade4a6af7128aa14ebdec947ce68fa455b8216e7823172f
z3efa6ab117ea215946eb42313c70dfcb4bdda758024342d216423617b3fa30256781bbdce63319
zf5f4e0b14b2b3b18f2426ec2618770feda3daa6437ca94b1b16731506b15f858c702a2c22363d1
zc4f4d96a233942e63c0b8a465150c7227372f31853b10a701b9c715666e7f0228b43955558106c
zffc05a9ca47712972722d4fd2de042777ae9eda4a9418f24cfa28bae5bb5e1863116642982f281
z66b01ae20a76c92935334d850e079d3537ba68d4dbbe3cbfabc0dcbd467437b5d7da25e7bd310c
z062ff03cc8fc86af35c218a6af23e4aac3a07c356c46ffccee0f40627f60451536d8556c813e97
z1c4674753039b665f03cde8b59add85eba1f31d31927085652be76c9428c37fd61cf61580142f2
z352d922c0248663a470e597ec2755c78534da00c093617022a0e7f590be922498bb8ed89531166
z14a094b5033543e156f6160f32a40703306b717dec556c4e902093df89a876463bf1cb25a424cb
z87aeb91ef66f3aed9687e7715e18e9a32855398c463cd38357747c0f79293140d7b80556f98b66
za54aff22e54b585cf3db65232299473c05cc71081dc663a10d80c22ecdfa4fdbe320dc36a57af4
z2c758ed71c56514c02df3aefcdc2f4426e6683db6392afc48b16ef569d3fb90804deb5e17ece4f
z2d1a474ccdc2bf952053370f1d7148a5f4c6c882a2d495ba30d520329ebb91e4614423b8500fec
zd3506d64a2aa1b1ad2a537239c229697a038226a636f7bb13188fcb62c6649fcbb9da4a04785e0
zc2d91c08ee79726ed699d0e1b16803827c57904fd891e3184a9a5c5f440383c964410c60525612
zf9973765d990b025e297de7cd0c9ff16668e56f37bd5c027866405c2f6ae9593aab376a1eb2cf5
z666842e405f259ea9ced798e219b35208f81dc881cf4d10531be007bb5eaa1e9a616380c4fdbf8
z9c9d7f3300fa1c17d5697922ac190deff63b0499787b08fbb3ed894f86df33a0d25c2ccf994f60
z490faec21e0a7660efdc33df3eed6d65cb27e3d1ca53c917be49efbe17c28a70e5ce98b50ce044
z24e2716e2a9ecbd9fb88706c03b0469e4c2cb42556de078e5fd47e21f190dcf21a3abe66353222
z4da170ea54b2b75b24ec9a7b7f3f1cc6190d68654c53052aa6078da70185e700edbe3fdfdb9d53
z015f84c44dec6365405c1587e191fdc49de347e777595041ba43dccea334883b8dab83813f3e5a
zdb61da41c2d4395f54e0931141c1fd9bd0db7f2188a249d7aaf9a046f14a73a0d5781ec3fae451
z45ce7249e5ec945b9caf4f2ff0bbc0e235f2cdefa65ebf8e364fab24b9aa16d27f6191b20f7f92
z6de277d770f021a9e7b3f0bc12601df6745566165e9f498d0efba2f4ea5aea536fde676c659c8e
z1df21dcd79c69a5756a0e0e6decf7279fe6c22233b85ae01ea933fc4176599ca568bd732787167
z928c7ffafccafbea096d795e163facb93732128132db63e552247a96f2a9395c5f5037746dac90
zc22aafa8237e158376e324dc2f64d521fde11f2dc7a3ad7e2e6ed6a403a734249209e7f80d5bdd
z80f62c5aa2e88daeefe1c177c39ce983476dfa47f616821586bdb7e6288b5503d59c93e6056438
za99ab81fb6eb091709a0f0d79ed436169325933b45dfae574385584ef4c3f8fe8580e07c54b0ce
z6d14cda7bde6c2bdf80c4f8e40a661f86672759d2d5aef42693a0a796dd7a1bad81357b9ebdf3a
zfe90bfda1a2bdeaf83bcd850a7aff1fb57e016f9484f57310fd597e76a483bd1b02e582b603bc8
zd61c57689bebe51bdd29021539a03bdfdede70d64ae3a632ce7118a1ca29ccceb2f90fa9bd8c00
za14483d916361d1c211b254ca1bef63ef0374e3c9496eae864648eb1c2a225b72e41e004d38f19
z4f73481ce3b97153fdabc64b5c4b4313f175ab206f2643e53b4dd958afe9658622621396c5538c
z621ed7fa26c4b35cd71bb02bc11e6b8a5ecbf2c2263576a3673ef137dd83cece79688c4361bf04
za5c6a3efeaf6686a014f313f1860b121a0fdce5eb66cf9a39cfdd99dbce4d7298275f539b1465a
z4698298f130f7d65d11b05d4c8abd631bfc6f4d47c521c300953b9587d06c4c7e38226f90c9c0a
zb0c8469193085f1c953c87d269fb82facd66aa15d0e86021698c9fd56596470a0d2ac44f1f26b6
z0ef6d051570f7e7a973e05a52317a7d64bf9331fbf15ad10635ada95031d337c8c4b272187bfd0
zc6bc9e491ecf37e0e85fa5cb9c05c47a301fd5cfb4ca426794f13dd22b30e9356f14b6289af701
z20b854a03cdebe8fe8bddca1c753336e12fc92402c7f994c6e4c840c40a52d5c0e6c5cdaacd841
z5df8aa4004e225257e493b24a64c9d654c8b48e0332bf1a46b076916962c948226ff86baa11323
zab37532084ff883d4320450d560eec168565b8450da8df5097483ca4a8c3960b2c7ad766b72b37
z5ce4d4da64f3fd4f9edb9be1ef55f435de49ee787632889636be22995cc1acb4337d50f34d28f7
z27ec679ef71349067f2a31da9fc3c84560d6c2a56935b68ebc4b25395a5a2773e73ef9084ab7c1
zb3cfc17aa6a58d7fbe6da2d72ac3175fc7374ff3e158cb8a667c13f952de50ff154055e5f4e939
z790e0b3f856d6f874c84e601cb4898c1c03bbe439d4592587375db157235977bd8682754d249b7
za6021aff6e4befa7b80541e5de298bda4353d0eb041fa04ddfba81eb119f2c7fd5373da57a1c13
z7524a28f1f6cf59d0500dd06b5d69a37f3d0f4cd6883f20a4e70d217c15b7e942b51bf8bdbe057
z23f1f4598b44e3b12c5e2569bc3fd09da95c8405ee6967e85d2e6adc8ef305ce394c5edd66ea49
zf7755e9f62e916033ae7a80f53600275533d67d967da508296e9f634b55712ecf9439b728c786a
z3a5cbf405978ff18577628052b565c5caf03ac85320cf0faa35482dea3e948d0d7b54ab95965a2
z800eb522f94d93f3727bff54fbf682ffe398f0132304226a852e05c534d409fc23cd5aba487985
zdffcfdba9e86808a78ca587ac00701cdf5a2c594c02848947eb9551ea7d721c51a6f4b6b695804
z631930cd8c2b670a75ff697edb35c0a96ce32e2f7008c074273c383f65f141693279931bc20fe6
zf4ca90c1dbbd3e89cb664e39f4806625c8728036575ae28677e89c904fe04b00845955d32a7c66
z5bdb72c1b4ef1f64c9afe34bdc5cd5079d0d6a48c5d7cbcfafa52f0e1fd1859cbde21d6c911dc6
za24dd878d72fd4acb368be7f6a4185c9bcb9567c665ac75745904d4d78e75f41b202a77cdc59a5
z1ebf2836d43afd4ab83864ef777f0f1ac7c4f73edba2003c7f23ce94e02bc2cb53742eab4a998e
z7c5ae5ec67e2bca0ab207ac1866d5b6eb98d07440768f98c74a9aa680af231d02e0db3c22b5a7b
zec4dc09ef63fab8f8914c3b813dac1d56b214fdb824ddb118f846268658eff7a28592f88a64891
z89bdc7c0ade63b448ad0cc7368217a8cff5df0a6d56d551f719bd639f06f39c92d59bc9fdb7ccb
z9542436655cd9a12d25abcd4a13396950c7328f19cd49019829f38c34991a4518a7e12726ec91a
z4464916257383de5b25b4f4055ba2299b3724b2019f5765ace2f93d278ed920b0d2f954b5ea9fa
z2ad073c8de47c8c1f88dc44560f63719cac701394fdc6304117ec9bf03750059f338a40b84763f
z29941bd93d3ab306bae7272ea09049a625e4caf2cd685dbabcf35d8df00f0a49675eb0a60259b5
zdf2b5c84f087a68179cab55827c9632913412133871c53ad8532c86676926af351625711fde46e
z150a3ed4e99f713c8fce72a31522d35a50187d40ee4a51c4112a0dba91dab67928927405734cb8
z996a2a801191bf88c62acc19d02fcc3c8b2ca0809e2e5187cfeeb235162ff00945fa9831d1140f
z209678aa7125836cdde7aab8e19fb22d0a491eb94732c5975b4d3af9145936bfd75256fcc04342
ze196e31705ec4c2c909a3c53a168ff720ce2212fc677ac5b3628265d16c3ff4e00d23425ca93af
zbc307f59952857d9f960719f2a9b1b8cb56c6d98cba3802895daa851e69fa37128ab102de05a8d
z163d123121246f2017ba5ab0c81681d7dd65fd82f4f72dcc130188f38ee8503a81b6604001962a
z7a0e4a6e030567f4d0250421a58f1a1e6ebbe3b7bd6d587e79b8ab65d12d7f50b0cdafcd67253b
za2449948e49a8c16baaa4e860bc5a65fb897426be39b75834659311963d304b5eb902f9a36a3ac
z5428aa3df2456728a734baf64d764c4f8168b31d1388d6c7a80b74677378407b5d30222ba6a69a
zb5eda85ef411d238fe67bdafbd3a5558cd86e7e9cf47d2e51e628c784f4fc9a3269a153cd8f9a0
z7bf217b5d5f18061fcbc20601020dd82edb634143047185083e7af4d6788e59de96ae0478e318d
z42ab5a5e88c664a335966181e74cd4466ad3e2dffbaeb57a16a80b2e98f5cb72c2304377051fbc
z5870bc50852aabec8c9453e16110fc7b5361ffe71707a145d2dccc14c200619eb9fea3073b398a
zf860c5eb5b8633a0a1b533cc18b61dace082107e1cd2209ed1c2889abeefd0e0dc07780321ffa8
zea41ec165c0f64a993abbd15caa2d0d86d866110e626c9ed5250db0883d3a089882123a6716837
z5d98f5b9b21b9c8e1fe6902fe30e1c9e91a1302cab609426783df3717d12635b964a275cbf19a8
z444ccf864d70f241058d5ceacd510f18a8f58b2af07241ef6b2321ac1b2371d33db318ecd2bf0d
zb1e9d51fae3083f3ed2cfc113a02a03fcb2d91188c45c76fe02be042c2d90c7a0585415ea1e684
z51668c1514ff039aeab041a421c99210216a1e4147dbad02930de47b601dae9c3736fd68def385
z92ca32562fd2e64777c8cfd69d0c39599385db15200ec994db1d715da0febe6dc29b6915116c1d
z2c2449736395b6f65bc2b3388c858a94ca467921064201d040e78dae4e5b5f756786cf7dab1ce3
z2ab67cfb53301fa5af065910eafe7807b8345038c196b456e5290ea9bbe146ecbcbf17905cee32
zae25faa13f670daa1a7de5141116a9d3debf31df116063644e78b8e7aa8f547b244a1fef6a4225
zbf854491bf5305acc2fa471c1be17c9634bec9f566f41b3ca53a8f12f2637f6ccd21d33297ec16
z818b46d92d121caaf55f8fda9ca3e9cca5c0affd46a2afd0101489bf54dff30804d99a6df1844a
zf15144d1ef8da608df0e29a6dbb0271f64d4465fe78d2dfd7eaf23888bdf9a120fb5332ae99fa8
z0d5a69a3e201a1156eac59fb84d8b411cb97111a3cec77a5c24ad4d83a18802076f1b3fa166919
z32458fb43dcbe7c127b72eddffe6e49da8819c01b0333a5e510f5c090cba589c5da2c999169342
z476ab1a7ac6d27fbc5870a5690d97f1ce4b04874930658574cbe859ff420cc6e740f9b65b76473
z8f3f72dc09b35d677cd17402c4542c0301b7172a18101a725e9166a6668e050fc43b2b893d453c
zd897202e75718ad927eb5f0e3254dc14278e841aac53638b47d23f1d4e41737bf79fbe6462d045
z63f004b33bc92e3093b5d32b2f932f7bec3c48ae6d7212d2d6e5a7b03322a4eb7e2c169e92cea6
zb966906d8a70582159ab4433dfa1f90ecadecd1e2bdcdf9f32b30f95f3afa7f0037eeb1ea754fa
z639a16ea476f627fa284d6e7c108ea20f9df299a18b5e5d36cccd7a0c34b3145aefeb20a4d9fd8
za79a10e0d4251b9ac845e0bea1a6487c1ae4d14d43761b6e9b94af9fab67488fc0ca100e0dc428
z5901171036bffdd1271444ac80212715545b2ead8085762af0c4ac993cc18f509c5b7ecff91047
zc699b29af03711de6b49fbaac929d84815ab915debfc3ef633278502f835c2714c68106edabf29
zb9a3cf90852da946a29d347fcda7127ab9b3fb83afe84d872b91ae519a7a2957a2d776721e391e
z5490c1f8312087374d1c22614ccd26070b7824fe411d22baa4836f443d6beef073536687d8a6c4
z58a0238074bb841d75e80c95305ae67fe54fa884950b584e91917f8ce1ebe6a7fba746f16d5d80
z2cd589745fdb466025957501d0158da964bd5b730c1d23c64ac12b644bb7226b28e29c243869c5
z31713241e5430159f51c9d4ba5d1cb98c40774ffd9648fd8b9eeb49c43a027e832b3a1c1372906
z85593feeadc6da0a399b98ba49f1bf2217ac077119639a9e431f46cfca65f621ddfbcac318fb54
z587e221678513d588b543d39e51e2942fe64b7441bd8b0c344975568df93b6ce436b66097eb864
z3bcad03f271cb4ec628bd38eb72a4be183233e3cb43e92be78df932a67e90172be0fca39a9a972
z532645bf9e13621bb8176e4952524e532554646834c7df26a6cf0f56437d91f3c209fc140004f7
z05b5fe5ba73cbe3680a75cafb9cd050c762e992a4a4ec2e8111c9d43895043e88ce7150491dc89
z340257c00523cda4da7bf7e8f675067b00ad5fd0f480088fd06ea4069414d31943febbc8666850
za9907fcad451167fd12dc8d7b39aadaadeb6ff2f9cb9b0466b22a79f7767dcbb1a5725c5224657
za9d32e327f63d1508b37b9284a59f0095f490d4a8e31164eb89c8c218b835ee9ba43c83a2cd679
z64866ecb3e6bbf930d796a77b871f0da3288a52d5914d8913d9b7b2fda67cc658bb99b82406d7e
z5b0f87fb5f0572220e1dd15e7515bd39efa919fea52c471127efa46c7665d3738ea603e03b2c94
z135fbb5d5368fb9b233da1ccd90f38f5fbd7c83387acc65bd07cff8ecf8dc3bd87d1a40c0f6380
zcea250a8f6fdbff92425f72f379d95007b2dbcf7973f7562df573167da6cdad40c6e70acdcf02f
z3b0ebab5c0e4106358ec1ed34d153c0f312205b0e35ff9b2988f2f4c901c6fc0da55af46f51b6d
z5e0073cd440338c8b34884b434015781b658f4b4a9498c759d0f2c8057d3571cb303fd2a1962e0
z0a23e3d5de2e2c6e6d8ff151aba05ed85c7eec36bf2ab33adc79d55d2733a439d8872a8e1adfa6
zff9b968f48958704997302abe2003cba0a9e2c17000105fabca5735c11d0c108213a2f8c7b8247
z31ef3d64d4a8890ea968b9297014e5090debfc53d80f0f0d46c95240c9751477abf720233780cc
zcad2b240cc8cf4949ddc8440ae48b99d02958fca610fb45fe09be018989e26a744544004fd7563
zdb0496d5fe88aff3a9f13cca1bb21923f07c421a1c11874680c55c55949a98612ea6d8bd745f1e
z0575b447baec6ad2847d4fe7128c1bb6b32d6b24e486928092f1d5dd9984d8ab7cdd6350714211
z07e67272f8262fae9963437b8823968699c0903095b3d2be20b535f224ee80eb70a87efd8344e7
z8b255127413dd2ec219ff55c674881492ba2f0fd0738aa1eac97f706d493e9246a5f62655a38e1
z971d9b6ce12769589bf12763aa5414276a2418d72b4a02094b28866c9cfe3d12bee90996d7165f
ze074f8c0e64614aac26c4e477a6293168d7663f331e3b8bca7838ab9f36a946b62b255b1cfbee7
z565f9a10dd9d64607d90992fa5042eb5e6e314cf73d27a807186ecadef3e2edab138d0177da526
zf1900a1a0258fb5146ffb61c73a705559afc1e5f76ca44fdc5519e1a7869459a019cdd292de46e
z98ffd6fa8784888066bf27506608e5810bf4e2ee767bf8e48d5ea0aeab0f09ff4375b2347f430a
zd84e8e6b32c338f47bc044c5bdbf7800730a36a892172fc35c27678043334ca5163ee903fb2d2e
zcf6f59755654368df4f4903945b67797dea74f4e3f9a02f3f142f219ae9deb593a266d5dbc699a
z0f4ac0aeb3502556ad0b9eacfd9987b0a5df5e061bdf492dc0cbfdd42b54dd886dfd4f18823363
ze0785e39ed33eeca7201c08508bc15027a2b93f5b1765e9a96c3debae5a169400ab5bec20d93ed
z617e3fb5355d218147311c52e3666ed910cdb8c9d4af918052c5f72b04236ae6311a027208a26d
zb8e94f0e2fb7611bfc9cef59ec43d0fcd1b82b63b15b5e42f377fbcd8d3f04a3eda65c93734b86
zabf437a44ad538ecfdc3300c4f9f2d7466ba0c1091af1c03c09b3a461b389b52b342788926c56a
zb61725c5db66035f830790812b98384721ce89b6bdc0a8d02773798d195dbc8267be4e32a7749d
z9188d546ecd18549d1fb9340b56af9fdadac68453e39c7431a254b774338fa2b5af198660d866b
z7c4e2fcf9aeef9ebe09455a071c85831ab0e1c8423b3c0cecbe7058b4a6c3b0141b82db8e7adec
z6a44648cf1e482c94470209a3736c9f0bce7332b1bae0c42b58603c52854b09193029ff7fd1fed
z180a7992dade751a23b615a7e298fe0bfd87f274c12a50f1c7384e414c48ba5893773d8b2b35f2
z1c123b279ac1bb0100b641f758a87dd2850758a73a969c87f6e30b254fc8d4b7b1f47d2c92afe0
zcba8fa5e09f9cb371812acdd54ea240114379799465973afb5ec77a3404bfc83775da4fed2ab75
z668efc0014f5e9fa5590e9ae6646a9a916cc6735500b23979fa74f3cb4a1f4c053d4f9647183b1
z8d997475eba060d8508b522d9c63e9f3f0e656fdcb8e5b0722fc429b13a3d534013d8428936708
z0f0a454d4cda6c39d1d47d17d88cfa0caba879267073778dea20d54158cd2ab04758b694a66bc7
z94d06aa7adee6610a3a65668b1b7dce6c51874cf6b254c65cad07378fbe0faed9178e41d1203c7
z4201b182ab774bcdfd3818e817c75c4d69e44b93e332561959fc243ade3a8ca5a2d9a97148cb68
zbf3d22a75b4f438a09fb8298cd618796b650f36eec7c7023796d21487477ee80c0161610bb8e63
z65e40e189e0ff4b54186cc0439902d55c68f92cbea62115922f087ce5d2f33d46c28372cfcd6bd
zc800f6de9adb26e60f51a5315a69e081da88510c4cb04c53b73c34a5634cee1d76cb51e7b7172a
z06961ffc30d423f9a30b3a25c6d4f04c103c43a72c2b3401abe28fd823d8aea68a2ee3d7708d0b
z7bbb74af8198a9a56c1adede738880466c75583158357a0e4f080084d9e96735174e897e972a45
z7cee0b6b9d812b8ad4ae794ab8892c5283744abd732bdda58a9ee2fc06091dd36654993ee88903
z12cfe29c4d25b6831bb1c91239d44e790a76e9e9acb234f47ae3996f4947b504e0d8d6d72aedaa
zf9447cd97ccc781bca4b59b9b9f480979cc2b1931c7f15f36a7797655463a4eecc29cd08113b0d
zcacf5995ba81b4ffbbf672ee6da6640a798dbf73cbac9021406827ffc84b130a3570b2d58ff05e
z00d1c553c90d396e49ea4bb3d28dd9adc95c98a27fd69492c2198f17f5625f7d7f592ae3e3526e
z53e36fa0157d2be7494ab28dc7513ecc40a9dd294fac4a6d76eb731e16c838bc6ff8d88e10e416
z5c53e4f455c753de79891e3615ef5094849eba9f91e9b7682652f86b2d4fe0cd9ec32f1882e11b
za2d6fac7ab4cd161de5fb560eced25cb94736261ee157c32f620a97450972173729ae4019e331d
z5fe76913be821cd22219d5d64bbdad286c732aee9647440ea078db711910d54bf691963be9fae3
z6d2490d5caae8ad27cbbb47ee7de1cd2a58458cd51e31b6bce66fddf41111a0dd62c61ef3c92a0
zbb185a65a680f7f8011673f65c3a8f2b2ba36ac530155507ca507022a452e89827e300392fb9b6
z3903fa71655ebf3311cf1f1c3818648751a4d6db2d48c8df35e325b7f63c8d9dc1802f7649b4d3
z07e0cca985f94617d2789d605dbe2958d13ac4e673dd1b79d265999d98ad8bf24588738b8893d5
z7915cb7ad68c354c033b042e7c7e8a0406ec681d4d2edeb62e7fe4aa37fd98db13dc793f7f5b06
zd369021936ad44ec6fc7520a38516f0166ca669bf5b29a3ca9ec5708b3715e2bdcf13fa0815f14
zd00c17cdd060492613beafbc3c79950da91bf8d03b34b28d261881003af89ff918484c1fd9ab26
z5447ee36a1a56a4462a3289a404b3e55f79f689a97ddb447f7eb411ce4f3c833c8556e0cb074ad
z4e3bc8904c9e5d8a937ca0faa71eab3aa2cf73ec8d339cde2a9a960bf0fe5fc97321a5e1ca9922
z3603685baf732f73b37fb820180e14b215e00e12be66b9c8fa0510e70ccd523de0e67bb339dd9c
za3924e63080d5a7452ff328be8cc2be352f83506f6ee2038d0adfc894a92d74d447c825ae482bc
z6101dadba7761130b964bb521eda96c504a314dfc909247c1d9bdc6507b62104a3c5b72e97730f
z7d667685374fa22b54762d8cba3f81a4ca971859ad6c948173305c47090f652eec872294831a2f
za1258dc29bb27fd417ee9a3f0ba037b2448281c530df0a1c83752c98000c541c46807ee33c7d78
z3c348da436c4e70b97b9bc3959e3e27881571196acd97ca487c022f57057b990140eb93ea98051
zbc65d1d0c269fe69b3db68b73b91e01783858441e6bfabc06625ab6e6ca8515360be9ccc249c9d
zb91b181770b1102520340c15aa01af0f42ff2aeb1fbbdc7426157c740fb5cc296e832a70645560
z30f47268de8ea5baccb5bfe8f2f393da0ae24388986f7b639d1a66c452668b0837993fcfff57b7
z1c17ea9c7e93c3954bded881a9cdb999586e0ad8372733c74b1c7b57e941400b4fea9e8a569c54
z71854da4252a179345e1fe92f9d972158da8972f5d2dbabf60dc14331804bd80abd48390fd8a03
z21268e35e18e2e32fa6f8e59e0e46db86bd0ae0f1afa68cfe0099dc988657bd6bf3f6a226a6dd6
z911293ec4c180202787c113107fca3771a800cec50bd74febf38d3938b8ca8c432be4c366da35c
z383a2d18c20d832cfa4a99949c720b36bab274ec89bf7a367f9800a7257423280face6ab8c0ce5
zd830fca651b0590af06d2331298e67d8483bc5b75bc132489464188294c05a0afed45040d0c624
z1e28f33beedc0e75741f35359a8156f91be2c692cb8eeb745d1d0671122746dae6008b6ff9b7e5
z24a8600638d8632cddd89024be85f9e644830e1ed33d8636d4cd2aeed5fabe5daddca726594832
z3acfed1a44e4e6d8f38d158c1c26dc24f1e5be9c8af7410d95aea0dadff706b91a6702b8e70326
zcff9b8a6f6d27143912b78bee319c42a23fb9e908e58bd5b8f94dbbe59140940f2c64ba13b80d2
z0b5f17d7e65a85e22e97c2f7e3e2d263532fa947527deed04e085cef843176061da87a969075ef
z1ebb974cc2fc4a570f657276db07d4ebceb353ffea4259d89a2ea9aa59cd570c8b1e75b797ab95
zc07b026424080f4733448f9fc166043e2aac9632ddb06e5a1b218f2eacd9c17c25c699c01ec9ba
z25cf243ab4d625c93eccbcb0d966063f86ff411502d8ab009737b71239b6e284b9d7aa6c600091
z18b1e910de40e167d551a1ae00daac5b388fc1bcda79e95d35771eece9a7f87d6b342cc254c370
z472203de3cda6a0c2dc524c956ca64627f6a0b54df57e29a6a30d56d0639c9564922f4faf4b20d
z0413a78c006fb741a66dadb998dc18e388d860b5128e262dc5a4198e654747a1761577f08a6d0d
z739bbc3bcc8f29f7ae2c5475c10b6230d2e024dbb9ecf03395f2c84b27b29533a0b777fb8d3169
zd1437030ed651a4274fc7a982d028c2b62c34a1a203d66ececfce831740fe61cccaaead84941ef
zebdc3353db3ab8eefa3254ef3e324f0f293289ea19d7bfca8c8771986037d8037d50608d3aed2f
z919e6203fca7cc1a685f982fd998e388f49e884cdeb097a790eef45fba1a4a5d294c987de42569
za058bc19734a6f6d9980c42f74a1556143892e702f432eeb62d9714392b2551d9f95feed1a4945
z3468cee56f681a938cb8520652cff7338b38e0f30300ee35b53cadb4b98986417490d270c8540d
zd4790178f96ad5251d313fe900d7bd5247f2a14df01d378a31273057e8a44de5d2258992278135
z1e97326db6b4859d34ca0e7efe8401088b67e0753c06a901afdab4546700bb0c093a3b9447dd9e
z521dd48c0675ed69fb2f44c3277e06796db735cd449f74902a3501a42ae2dbe78b5fb4cf2ca785
z370ac2b0c272fefb227da8a2593104405680edddb1cd64f79c08503122c1222aae49c3be02d915
z68351b0373913649f00e342589732fb19818deb5aae33003dcc02d4e126b679b797602b7ffcf61
zca62e750eddd98cc9ccc2100dd633379bbb8ad1006d15047aa9d5ce70987181e5256cf50788599
z5b739f9902c4b34bd7ed55c3159010767a73d3b8d0e1749fc1f69f1d88901df9fc4e4985b0e3c3
zb80b9eb10fb687ef4493eef1c9215e958b51584e71d2ab383e43a3e386693dc7ead2fc49db73af
z5ebd99a99b7811704afbb4b60f31fec1f314d9905cf5e0b88d58206ddb118b3a78b383fbc421aa
z7d42b0dfed107d6a7f9a12dd0b2885f980cacb11d742c80e05508d0d48551773512440d0888520
z898747c5d5a63d49c32937513adacca2b5d9cc6b5e7bd4b7d75c70ceca57d94bde2b3ceef9e1e3
zdfa8b29fb455ba874b03a2c8d4a10e55be83d62c4efcf12ac50dee68fb677f0a1dbd59fcc08393
z93ed39a812880576f5ff5387c2ae8f8c66773e2de23e3c65e26f73782fcb628a858aaefa559110
z4aa54a938ef8fbca3ac04137fb1a277423cb8748ea2bc609e035684eef29effe3b0e0b874ee435
ze097027ea97efe8d0699b63d818d4120284379b39d8d94235090a98ed07af9929f82fc5856cc49
zf1b329808bbb3345a27398e92eafd0501f77286fd74f531f9362c4ca97a66248868cf46a48562e
zf3ef43b378d692d200c8f5f9915f06601c8a6fe0795e7a341e296051b88450e808e0f8bca90dba
z57f583d964742bb8fa71f336ca0a5af72c3f92df3ef41cdcc567bd6c138fcf0895b40847043823
z13c621f66f37914e72562c5bc2a4c29eccc1f8a080473467529ab62d84b03dafdfd9bf455bdcf3
zfa4efca03614c05e44dd24966776caaf65aebbaf361bbebab6dd80935f51cf86feb299a7563c40
zd0452a05cb1d0ce917af828b2abd6b6c4c5d41d34be757358c8863cf7eea6c5644ffe2e066365d
zfa09893612159b143a7f6ae8a98c739643d4bae0cabc93382def1e867a28c9ff45acca3934063a
zac69a5c3ae166484b0a267803cf89995a8f95823171f52cdcef24b896b9a5de1be9f6a37ce58ae
z0d0276a21f6b6eb11cd5d50ad56f129f259e644b1042be3875ab2fbdf639f7da60c99504717719
ze475dbcffb3b369c3894ea1e0793e227e113c6f8a675a2e8433728d85571b1788f8e6c13cd6a32
z04fc15ed434263fb2103805c756d8a057314fda3a86d6fdf55601bf8d3bd1daab0c125b55fed4d
z0f52d85cde074ad1ce139fd35982c33161f2b9f6e614cbe55a9e110073041ce031ea661fdc3375
zc30843139ebed1f2eb2419d706f54f3842a85e890e8858795ff0d5cbb0e2633f79b8d4ad3e0b1f
z1105e2f7b8ad96f430998245104903701a31b9710c8c0894dad36a42db09e9b4a204fe32a572ca
z6eb39745d1aa1063268e779f78f799f84398cda0cfaeafce739c5a03be7e4ad09c504024ea3a6c
zaa204be128ea75a68b3be25143218fc2df3abe905fd3b6131b40c8d25a3ee5217f374dcddac4f7
z3d0f1fe24aa0bce381a5efc62bebed5b3ade9b3e5f54a12042308e18693fd6850d0bc53a3ef716
z8a273f48ea2bce3d2278399304c2a73b6acf0e795f733be05d7dfcda6ee01f81609a2eec0aab10
za19e40a2f3ecfad40744468434ec84e4fe7e6fb5b22395ea275f5ef8dbf567bfeac8278d47e43d
z1624a05121a67532c2c8ab61b9061424e1cde12202cbbddd6bb22ce1ee67f32cbfe31d513d9c03
z1b71e9391cffccaacf9a2440ca3362d9088111a4c763049ee11855f7781d3bb37cf7f65598196b
zb28deda51a171154709de2b25d6977f2adef4435e1d2694776edffa5a328371639154938a16200
z5110e78262fb3b7248985044f2eab9ff0f7f41fb7330150ce284463fa148fc7b7185e48d8ebd95
z43fbaf7ef1a69767e382caecd03a6b7dc760ee12442da5e8e866c04c25f942a7d80dbe5e4ac112
z2ed037b0a3da434c1009bc905d20fb700a3d57297f3e5b0ae73aa9a82ec2a74419f3128c41c50c
ze6e269ce11813c47fd71a9d4f2e0afe64fe40fcf06f57cce44de4841f90137184641542edac8dd
za14a86b8cc0b81b0f4ab6dc13c45805bc6c7eb25168b36936d20be57052ae23976c38036a4b83f
z81ea57d7543df82395c730f049b0c9d33757ce707357f99fe6dc057a87595b4ee530be8e0c3ade
z12c242de2f4456c287b7b8c75335f997a5999d15561ecf3ad0982451996e50d225bc41ec3c1ff7
zb927f9b116217b81fceb5be948c3cc2150a7993305d3b111f5c2efe782b876ee62a7c4aa06b3c5
z85bc8dc732954b34102edd0e81c09e70ed44dee8e990a4869e17c6cfa4a5debba94f28a458ac8f
z08b3b3ad647be523686177b5a6d2d28b160537e22556fc4583f6a21433231692459899668400de
z55f9edadb81ed7419e4857f7f1187733ad0e240a0d7c16b5dc3da87c44267eddb0e9bb9e4093cf
z2a4abc385c9144509d1cc1bf0fbbcc9055745d95e0bf3f0b388664429b54a138e66314009fc4af
zdd92ad8948e8d3dbbea2e786148b05cd15762dd5a3b3f67c1a82cbb7c064d90b83664e9987e923
z43bea11833242823268c0da1b3231aa1d44481d95309684062528670955ef7b430e2c8126bf3f1
ze497761faf3d41f7c50b9fdca486c77db0774d643233e67383bcf774cb2a6e4e79f2ca68c9eaa6
z5f7b405bbf2b751128232801e23bb6c15c2c3b84f9187eee632fdef6ed5a7358eba714010dfcf4
zfef90254e02d527b0a5ff2b7ce4164e10bb89621e509b83a8c6779149aa59951aa0c729d7a3be5
z2b07e4381bf6f28c95a69736bced0a7f543c3e850e9f17d1aa71e0eae1767fd98a54e6e046c56e
z067174e3e7e04a1a8b4462fd954eefbc5d54672f42ae9f29aa9f8864e7ce69cd207cd56c753e0e
zec3f60e170035a9222706c2371062d259122a7814d563e56db9033b2fb8522bc3c4fea5d706437
za8ff0b35cc34a9cd99e760e285f46515c0b06fe8350b22bef518bf7fb9ace3bfe826f69ba949a8
z693c8912758ae2f560b006fc532729a78d0df2ebc5c8fb94d2ddad01e1243a4ddfd3d2cbe4d008
z0073228f65a05eb2c7d3af10335e422b9e9da08718332d50b22eed6e70d88e943415076f66a4a2
z3e56247ee62c26fa217ffc823aca29ce0c99ea48fccf749255bb3f3ab295e31b131ce5f11eccf8
z611512fd027f82b570c53b6246def3b8e11e885d8b18964592462f300498d75ddc07095125b267
z343aa03ca0e1253a46d47ee0fbba5a762fbe79cef992641efa16117f579b29742c7c78eddc6593
z2f8a6903e698dc2a344d5cb245c28167fb279abc82516922ac8f3513551ea25192f3848dde6326
z6feb8c5d5bf1afe41cacbe0418790d45a68289e8c291ea4c78c8489f2acceff1ddbde5397a941a
za78b840921ac2fc165536562a9a433ab55070b0d2c86abda38e55b853aeeca1c8ca702174d505a
zd4ea9beac66a111b094a5302d6a2989bb0bf6936f30c36825e9bbd661dc6d0d22ee5bd88706e42
z12c522fa1dbe431653012ba647a8a7c267655a18ffc8e392f75de85bd6f4b4fc9fb55e9bdfc6c4
zf09fed4894f5b18a224b604577d9e3df91d949bbd2fb44e71a5a9489de9c640472835ac4ef7b38
z133e66bedfb0097a1df15d3a7a609c837632989d4d4dbb5f2c1098ac3c32af3191bbde7cdde8de
z93e17fdbc65b8d2f9cbc902c96f4707e6763aba964d1e86fdf6c9fc43bc8c577ef460eeb90311f
zab12f399dc948db7bb210de9fe035b40ef95a07a87d7e40492545d456f4d2099198fde0f0e623e
z50132251c28fffe76684186898f75bb752d81dae1f9a0bc14a818d0b4f2720807a48e006e33489
z67dbe9d7634d79428925e2ebd21dfdb130287179a3c1bc5ae895c724fe6f7167efa333908b3e70
z128e7e79052764fee98a190243861eca7ab99247c48c3f911982f0616e6b03cc1c48c0b66a5815
z96a7bfc21c325aea4d2eb4be402efdec2b83cc9e1ea0f1dc1cf261d1c41623660c598fe51fc6d6
z6a031474cc6a7b2e09e95a9a6f0a0a7fadf80fcb0e165e6144894f57e94d72c7d3cf886ce9d15d
z1fd082cb0df8f41396b3ce97abc93454a12e64e8fd95971c9ada5dd7bc320e44a2549d4b2c40e5
zebab18d93a5eaa6192e9734fd67e8411bf4ac6741afcc5ce87bad3ec6b54b602690f3a6be732e1
z612792b6f59a78eb9c0e94ace214503c7e641ed22eae5a10c803969cc4eac76ee26e084d1d43c8
z3e5231f525c871b54d6518cd2a4a438490b34208fc7a7b7c4a71ae2e56b33f99190fde2b3e3537
zc8d12331b5f5e7fbe835404ef1a22bddfa6d72248397ee64f0cdd0530ca6c5c1282ff40ee885ec
z5376e2287397b669ee60f2eac5b7d74432b85f71cb0c24ec54ddd7024fb8cc6a8235de04445279
zdea6d530ff8a8fd99c6664d993dd7f38b1d3b16a1f158e9097d4705d4a7512115ca4ccbb701744
zb525ef15ef1bc0614b2d52252c0abdac75420e9041f016a4f4b191be2fc11fef8d40f4d89a4a47
z7e72df8115f9897cb13e17c4ba4ffb3acb9cc1b4bbc9a68ca099780685642bba9d831ee7e689f7
z1d0cac7acad93ffc43e6ef31f51bb08598a31dbd1d74044e5a7bffeee413fbb1b71bc8c1950085
z7475fa04f25ddac9303ec8d56b28c2de48c42fe1ecf0ae28fab0bccef7557d87416d463289b953
zf94d2843911beddc630924df274b81370d58d369e9292f6bbc7cf476caa7ccbb92c778e5adbda5
z507dedefe8930523ec91c04bd8c8ee41280cb0dcd7e76f079348247b1f407e7149b08d14f28a40
z5d5400091349ea1b76c9854ade8b20dccdaf3942a32b99195bd4a64837b1e19a0c048ab0e234ea
z8951a689ef46b0ddc08f2a64a3beb435fdabfb4efa56e02528e140575f72e2b9afdc809080a2af
z0a8e7ab8eebcf87c3675b1b04295d9644a429284df01e824c3095e97d5d8521f72a6faf43f6aaa
z08316a099471ea7ea28be124c7ac535c70175ef99ca6ced8fe8e58a5470d823b807f1c4f7b380d
z92c9be013d4f5d1cdc926d951b57af8a1451c3e971063cda30ab38748a24c58006b98be4947499
z7a8a8d5993f22a49f8a336150e981f0ce88eb1432f8da13a5377a155082bf199f763705256992c
z45885158d0a3315b8b616593d34befac1eb238d29e9aefe64d972f05bcbb0d27e86adab4e1ea8b
z035d44ba85e9d082a255531ec0fe321aa49d35bf62f5c1637b383a1391a870d488f1286ce40ff5
za21b75ef7564f51743e9aaeae4d37ad5d6a0f8fd611f92ff5cd8aaf760d831ac1de1a2d9e7d728
zc4b56624ae882a901ad2a39215ffda74a1a6bf41176968ac03f2f89617eeb2b20e790b1716565a
ze4a4775e0e887fbabfbcdab718f90644e1be6a8ce72f6b43a696abbd64c04ec853c2afe5f15b56
zf5e274c9bd1063c194ceaadd37bef800ee8bae3cafe1ad375c9350a7b0b50f8abe828ccd5e5f90
zb43df8a0a838f115db4fcbdbdf236fc9a37197270722309ca025e2cb94dc89f24909f5b266cd64
z555cbf28dbcc19967c8d3048dd7ee144a544e6f99ea218e5fcc5f4fe51e10f30d4dcbfa6a91588
z1774136063420ad4d3f9f67c326d15dc0f7dc2cb8d7116ed2c79e373ccd2e182e42b946e75c655
z90edfc6cea20c60c33809f670cfab49417b18cd66d2e2b0138e324d33dfed1a62717a3b8044dbe
za4b4f57694e78fb7635167b695acdc3e799efaae90a644d9aa600ce49cac314cd4608631ddbefe
z4ab4565ad3045cdcc00c6c03480878367012383743233fcf90473a51007e44050bfc4fbb240dea
z94e129f0139f97e189f6a34029f23d53394e2d1a4842fdc836c695767f6616129ce69845c1f373
z34a3ae8f212e5c17f53a0e60a95c635943f649fde62ca17d1dd7ee13f7111a9913bedc84bd4849
z1f5c9677260709d33667a92d3a27679bf80bd4a1a3aa609a57cc283e8e8f1601d6fdf1f272d20a
zae8923f5b9700c21e10b2442ec4702f6380c16eeb8ac69415598f780385a7b771b0a1a542dd3e5
za7a848de4e9c2d988ae013b8d447b85bc5517502914d8fc3ee9cceb13f286b1f445be0d2eaf9e7
zec522cd1afb22a92c248ddd5312454c9c134925e665e017a0f8ee4131664403839b837b3ef175a
z89d75a2f1953029ff23b5698be0c9622d1944537e766578848a135fc1dc64852420e455761e410
zd7162e4b7af08022968b4297955abdbc52a4a200e1fabe7952741dff9cae9ee2befbed17692160
zf28def895e5add2e0eeb59d7dbdd521e9f04707aa8f30d381b415ce243cd782c572f2928dbb805
z3ef0bbcaa19c82528b1682d91a3641310204ecd5c3802b172250405e9601908cc6a57433e014c6
z705ce53632ee9674d78e08eba24e9cfeba0ecc8c97d8dfb2496ca321b6de67e43019382bd1a770
z96e5fab6e919e39070cce563526d25e39c6278b2f19e97985f35d52925c533bf69a79585be68c2
zccb2bdb936682cb7b327b5e20d68f3ce832a9ff538ba569dae2182b2f99f5e541faedab7659847
z8e26398ca5d3ecba7775b00797f822f19e4c4d751dc8f47229b295e44b8edf78bb7a659c5ec2b5
z41fe17b594ac0ccc5504845921883bd3a6ae3c3d1b88e0d62be83c74127ad88e65638f2b7b3150
z38bb4115c0a089617dda2584fa7faf568ecab32d8457bf86792344f170b7471c3a6d3bebf52390
z350abd88a271f5b3837449c15ad719666d992a50a39ee1819f4a0208b4c36a47773ca9899b583e
ze2e9b34d17ba5a28e9d7f2225212b271845ecdcaf43bedeb19a1fc878bfc8ae346f552cddba9ad
z9ccb636b988b9b8e4bc16580ccc5da6ccc436d4fd516bd7ad7ab3b6557869049e8fdc8c8e619c2
zab4763b23980f717d16df87052501615cd73094c7eca82f022961dd62c24433046d56e3747f27c
z37f40595e6b3a1231dc3bc6eba164734ac19707897387dcd4c7df87d3b5fac717d81ed41f8172c
z96e761eecbaeb7fddbe9ca7da2e2f83ea70ac4e6143ab7e452f21ba9079795bd5b2a48f0049aed
z437f32bb529e4f10663c8024b7854a183296882ce1570586181f3cbb8d546a52efe5bbea0407a0
z363d8b2a78fe5d774048a484fbd83a5e1e2b14162941c1c18a76fa93880d78758cf1b3c1571f81
z1802b300e8fae2076b938378a1cfa774f1ae05335baa20a34dc02b2643637714970d88fa9531f1
zf327990a129bca2cb20da1cb60aa4d55f12e15548c90d9a186c2d1e3b1f152942ee41c298ba08c
z06b9e93ab352c237101e6e45cf42651158908557f2286cba76d780b03b47f99af79fda3631cab0
z4f2b8605d812dec3f2096600f83565a0afad45938a8b3f6898a753ef1ee7c7c1b7c5ffd9522411
z7c98171521fe350de2f1303c04d04c869155766a96a21c23bbf8387a62c566305709a5ef053ede
z7b4373d40e65c43173daf388dc0f6797572155a7005746c467bb5c7261246962baf59302016902
zc13bf063fb6d689d4a30054820744632d052ad24f5ebb2dbec38199e6461255e61e28de648682d
zc861a00cab09be5913e3d1877f0189c24c342749732fb2017f713b1d98a522b8420fd7e7740428
zcb4e98651d2a6fa6b8ea9e263dbff63e61022fd38e76a388023bb784bef7d971a7dce5879434d8
z72c9c7043153dfd0d0e1d613d734ef4c9b4cc250d9d0dd5f86cc2af825e79448a1779fd94c0032
z6a96ebc7674cf7718b885027fd579647f366446c789083d0a131357e8c4892fe0df7356e92c22e
z1d316494ec936f8001068b8c706529583909eb6e32bd806d6051f295d7596431ff98a751d32765
z0568c482cdfe2533d89f130e6b73dd3b24c23b90b286bd07fd22e4008f93ba3cdc01408b67f05b
z4096771cd265480e68c54b566ab2d3b8ded6298e000447b883b7a61671952a3acb4a496a182691
z8e9cf86b04016ec24b398bf11a3e752b217e7658b823a0f5792cca5d78c561abf4a658ecd29ac6
zd654c2c6a3778e1280ea2af9bd104c876076e7e34abfeb6e4b4b508529c524b8372cdf41b037d4
za7e0f6db4ef37a02fc24afc4159deb472d82fba0c9992fb16d75dace9f301beb71ee1c33ff4d21
z68c061f8d3996f4a25ae8a754d2f11228d0eeede169727b6a4d0c0bdf1ca344f50b75c738215b9
ze0f683cf7231e61faf1c01899d11972666481ff96777f1b8ce693f78d250d24a8440508363003d
z0055d2c6d5301c93acac1df1a98ffb9125b136751c28b2557057244ac8d7cce26521c3435d4a47
ze687aa3a7e776790208d60e39f902a7646a74a4e11a7736da0259323e3dd82fa98f4340ddbc2cb
z6c7f74113fba650a83fd7b901f88f5b10359e50dab635958be4ff7df776b0b0237b5c66734f9b5
z2fc1a87457b2235c4b4e2ddcf53dc29a871c66238a4423713d56fc1de1b0f323275a932461a247
zcb58018965160f0987c10150746f583c8bb6034d95be6b8dbb3a878a6730fb781f0c22c7687827
zd8d91b1a09d4aec431230f2e74765a9ab59076911bd156f81d5298ffffa449730493b6c2c12d61
ze414130205600f8790258f5eeecd50a89726631367cdd014d95e07d41de900c9714691a64f552d
z7df8690366ce432d94a8f6f15a8713253dd9e5e7e6197000e944e226958c47b06f6fa28fa3ffc1
z5ec691f129ebf33a716243fd709de0d4217d99726de7dc896249b1439454cad56978ebd9a7f325
z4bc744e75af6b3c7124cdc87433351e82c276646d1ff8c4255b95928d7da11473cb4ef727206a0
za83eda9d035540aff6380cd1b51a2b10b2d39863aee369e903ac62a6e9d509e1c7ee74e69de2ed
z33b3ad9894d66db21a1c4ef5238cdb012119cdbaeb516effe4c3278bca0dd9ec330db6de7d5663
zae6ff947e4f9e0505c100cb5c3f6b51b578d8812fdb547f813e1a30d120fde2697c8841300aa3b
z4a4dd0a55f316806f7f81295466b66012b3d961ca63b0a3987222e02c825f2b777d3c4a6abfe0b
z912976c92c67e693ce8455d6ddf34ec3f24fea1f83cc057f6d23b0b4165b069fec8fd0c541e7a4
z4827fbeca36a6b2e1e68373b38bc0337ff3fd588705793b7a0718f1afa8d4b4d0f59c370b79c7e
z75a680259617d9e38c191fa3a292a9e3a3f3824c989484ed1532351dab163b645d3cae9178844b
z9a474887336dfdcca3dcf809934824a2dd824104b35a489834a88b5b844ddb4d164c6514b60014
z4537b19b15b3367facdd4d84cc966471d5510cf6831480377260b5aad45ad1893bda71f70be1ef
zd286a849e29e9e9b92146ead93a24b39f092690b8042b2a6c4fe425f04dd74eca2d0f5f97b4aa8
za3a1ec5193b69cee5ea474f9e5f01a89978a2dc9a701190d22a913297f84246b72dfa7358c451e
za0e103ea04ecfc7df349f524bc36291f508c1952d6a6864b259491baae2621c3ce6c78f02598dc
zad4deb2cc854dd0f2ccea87f634239e75c9c70a8ce3bd6b53f15ba8f307dcbc7073a1af029fd01
zf2a7028d9c13397a5a2900bdc943661dafb5e4630d373b3a9696612cc6d215c9e1d61f3c0b0449
z378d9b1fa8618c8a287538361d6bda3ae1139a1b4b2c86ffe4aa394ae653044e7fce92aa263d38
z9bc9f7976946f48999462bda14cff2d25f202caccd9f00f121252d4ee79fead2e2c3b0dbfd37d8
z2dc4e62483bd782521eac3f63ff73e9bcae8ee92da1228d775562e69b0c86b6d938393f6f28535
z4a3241bba171c89bc1c2777a0cd182dc18976cff7af505bec7927a6f2c29767b26e05ad5707100
z13c0a1ad7e843dd470d199538b0c60ae70325301ecb1e797bfd88aeb248217fa8a410da12284be
z36ede6fc7ba0e255357713f2545350fbbb9330ac1601964ca7c25185b25e4be72467b89d96963f
z8ffc34aff0615ddd6193df3ea24673fc404993a12133f3d867872dabaa7d600e6fb9195eb7ef3c
ze3b4c111c7bed9998f8b26adb4f6eb095525600288a637bd78aac4dd88cd1aa38e63601739e4d4
z7d93fcebc7fea33083c6bcc06b528905450aecdb24fff087ade5c21533895446b1c4f0e6d62c03
z6a82ace9436eadf2168aa15422691b33e64b3e1b7ee4c92efbca56b9ebd75c4a970b6c5d98a54f
ze18a1b785ca3c9ae1c23a7d127e72981cc1ea1ee641f8750ff61e187b53bec6100b964eb3479c1
zddac5f35c574b1cb68d3a539731d47d2c5cfdd302d685b37781e93936d060a9acf91e467964e0c
z68b2fe6280c1133a0ea154d4c51192f79ca964dcb6451fb15cc9dc111f648afd56a1453641cea1
z7621ec0d125b6324310a3d7998a4951c4c328a4ad60f55ce5fce86b84a7412f6ddd8e4056286b4
z81d1eb1b4a4858570e813d2d00197fed1733666f17acb052509d158b3f740b9566ecc03497f7fc
z59ff4803c28d29838fb01b941a3295a13dd019ea2b9daaf91481c6226a6ad543f5c843d89ffba1
z130095224b9466ffb0c40aad7aaa3a3f4b0d50ec157376895892e62b8a1783fe5e7791f4124cee
z8c3f41fbccfdf7668b46b4f6783a08bec26c5842dd85e7a915376b53bf780132e984f437c3575d
zc05d0536bef279d095ab1885d78ca72656d7795536431f7f97b3b8dc3fe1e45bc4a1aaa4c1bab8
za243d2c8a63a7428a25055212843f3f941288c707dc87276997e7ad5aa1799cb9026b16f782c91
z539ee8c057d4883970ce7cb9a70da3524afdaf749b9436d68fd63a1f6d3977336ec0faf1ec9cc2
z7d8e85264de5ba403a0b3f94ced29b0ed4ba6122cd28b5268847c1b83de5df06a485e9e1355be8
z7e55ddd5741aa46208af60371514ff25a168a41657e4279e2455f463a5642665b9099d3278a589
z072ca131bb3be36a7b37c142bb8a401d7c42e98807dc0998c8a8b0cd651d85f3910e46b69246f8
zd72d77052900d0627c771216bcbae0917ee2c9306df5ba8c6f681a5e65c1ce7add96b6d9f75bfc
z3e534717acc6a39c5feb5f8744a472394413c0a191a879047176eee34eb38c8932e66994762cd3
z9ac14c234829991c9a3fcd2d9b2ecc31853a0e57f753079c336bc56872e4f5e9741166c361160a
ze86d1619a95b324c6ea2a43650ef5287a653e8f7e20ff9e84484f049c0b398c958bd5d181642a9
z06aff0ca5d385e17ea5b38ee3cc5f56e79fff8dd490344070cf78b590f8cb92386005788678978
ze5bbd560a316e04e528f9782f9fdcfbd40847af680b072b82da35f627d8e6c8952e5f703ee9a78
z6dac4da2c3c725dcfe8e97eb8795e0d78d67b2452ffcf534fcd54d332a3c0368f904351f7275ef
z3dda081e78a54123d829421b012b78d5c87255d380f1dee490afe492f8e5d3c598961c879fc56a
z3b26be58f9d34efb8300d3f0fc60d7e94167e87253a4dee8f5fc07f651c4760c35874c9b4c363c
z68d246aab7897b3e32c9b360296f064af48568e1415c373cb495587d688416f29ef69291c08bc7
z2d22c1f3cd83121b8ec7a77f3ca586ee33278286f46a0f2a8128bd234431437678b72d53061c87
zf7399120129b8cbbf43b2441545146e7a4f0f6dcd559eed7288535b201fb01141080402f1bef11
z58c2b34575d38d741f3b9030edb9c4d89655dcc9c14c7384d800a7ad1f85955deb63d21650c361
z60be4b1233f71be6b7ec4f6d4ef2687b3811e807c5e68281c473f61ff161886fc30500718b4ac8
zeec66971b3fd2514168015e883a3f4e654251fbd3597e18ecd947808c8541c1e5f5f3cb5177934
z16b8804521d67a0256d7e3ba5af91ad31fc9afad99149b79ce1f08d6e84c94fe112a160857fa2d
ze0525c653d1e5ee340608111655d23a9933af121da57e89a48bbb7f76b84b8549e49ec15efaa1a
z3f48df3e5f801afc32d873e1e0c5a980cf7ef251c468fca7f21433c1a5667f26ebd5dd72c064e5
zbaffed58736357a2335822948207de51e0a2415d610cd97002c3a5b9ec88fd0a02983353dca97c
zdc4880e55ef2c1016eb3809476569c98e47b3a22141411b07938c2bb9ea5a36f90c6827b2a5ac8
z832c58e9213e57d0799750e33a75069a3db6bcb4b83917a08dbf2c84d303358b7d230125cbeaa3
z75871f0136ac7623dd5ee17261c3543d65103668f54bc0f82009f459d1f3a3e3e867d54c318e6e
z0b889ec0fd02b27419c698d4a2306eb5ea6270ed8e06560acc32ea249c67600c966bb8a31683f4
z23cfc1d3d073ea9d8470a4f3cb1353b95a7b419a9e21ad9933c6eeef791a5a98e598b42f3750b1
z049fb32eaec3533997d18d69de664316c51fb8b0171d328d863a17756d786347dfec2ca5804e22
z008089b801ed22cb6f937a108ba69bdcee3d8d0dac24877a3da71367a3ffbad314f10702abbf39
z2815e79f2ff2b6b06fb3caee8094743ee1b81449884635be0165a07f4abbb751418a6009ad7c6e
zbc15bb46e5eb50f3d3e83e3bc8443d82b472f4e211d1ba3bfca181bd79689b5908c6d0e79f6761
z64ed04fe719bfd1d8063952f2d7b7d2b3d45bb0eef903dc3b5d2e220d7d5a84b29626966e4b3aa
z06eb4bed17f256a8ea9074be18d77ec80e11e67d1b04af13e778a5f973c76aa43ee4c6d73f9b17
z88929dbdaee36667332638ab70db93f5df2c89feb1d99f7c847f30fdad7e8fae86e389c16cf9d4
zfd18779f6027e56a9f8b7bd051b32765847feb75a054fb8c1157590b02a1dfdd52b77e686492e0
zeb2178f0e0c05e88807a2c4a0fc148223354b5bbf9535bc1b27e09bd050f09d46e9a9fc7e1f65f
za31eaa34002a5b5f0a580ab1d79c43bdd403bf05b808e25ec09878eecbd0a35043f091b60305d3
z5839c713de9e4f06a4a1654c676483ce4395ff021a9afddb0748736ad2c5cc44f931f273c0e0f7
zfd3dd5e3cedd55afa21f22c7e29b3725f268721954a5197776cd3f5fa2e0d44655df0f008eb5de
z4ca61a6a452c77a2c1d8383767dd2514db9119ca113c20bac6929364528bc6e8e5383084c786fd
z499e3ea54dbace0810274ebe31b063d15a6d1a6c1f8b63e66b9090fd0be5e457076ae58414fe59
z80e22c94cc3fae37ffcaf0021fc45411c60bd783b02aa1c535f08a29435fc05f695ac0c583f382
z9bdffa1cd4b35f8680b96ee695b68b2108710592fcc25a0ad45ee0674520c8725eda4133fd982f
z6c8a75647187b9e99ec8e153999a160e8e2b3e99144b95894e89f8e9bd493b65367359173efc56
z2554a3235ab8bd5f75f599e8c8e094bb895719a9952723d84d725977dafe7fb24ba69155744ef6
z20bd60283da153072131346d96d08b712bdc46081358b3463d29ec94bb7b796ba01fa5ed9e3677
zd4495a8134fd945b622a58c745b9af72402a4a3b5ed1a70f31b196dcab7995e8e2bda682374c3d
z552a47fe2db292f79c25e8f0baebe7b4528b0be5942ef93681dfcfc7945045e367121e7effe083
z4dbdacd669c282d8a1cc5882444f6f77a79f82e5b60e28487d8e830b4686e59e79a10832a1019f
z944785e196e01dc68f1c4d8aacf3c03fd657f3b08ba1a9a29dc4caa392a4646d6a7a7046afd62d
zb6dcd70e7e6b0668556016c294a5bceb087cc19502eeef03d6f0e56edcb169bf58c6b0cb19a9f0
z9a71f9c38cf793ed020625025b47bf8e5ce173e88062d1ce8818e392677ec8d2335a32e56be081
z2ba358e2ce61ca3959ae128980dd10a92dd3e46cc6db9b87e1c339ba63f3788bf39688814615ae
zc21d18ceea304ade54f05a0bacd31279c7e4f1ba94cd77e1c205dd07b02d86513177df166db3ab
z3de987f4d5c5684e03275777797ce7ab508867a92273607441032fe87f862bc48f637a83f0b667
z2386bd9a660ad75247d28c64dae2623e72ebbfe5a9e363d0c32c472d521d0b193a2dd95faa426d
z1462a71706dd446eff8dbb208f18217af5d2009aeed06285f1cd7aa667a7303e48b1f36b296aa0
zc7919a56ad3fb597edfa7958cc9536a2549eddfbb7c2674f4505ce5a8268453a9f09e76344915c
z04a1c544bcce75e773c0090e2c0ff5076d6015c3d318389ef037964db8c0b19884a8b9a6da7755
ze9cd5b94edb92b98fef1c6d34e67896379c2378c3ff6d6ce089e8c9738a83cdbf53f27c4187fef
z4149e75346c78b6b73519221f919e11ba19fdea8356ddccf532d321060c4a14a2b256a4153281a
zc5580343732cc70bfc2fcaf0ac4697653eb6bd712ccbc2f8467ad95e6ce57d40be2c47cb29be1d
zc96dfb92f282747fb28e04eb4a9cc1ba26bb17871a949bdcc280ce0f972d3997afca43c333e7b6
z2271bf2e70c28caa3a24dbdeeca7c28cc2e0d805414a55d4a7703474fd962b537e9f948f01ceca
z9cdc2d5659563c0e304c83fb61ea9f48d68f4d3f08350c892327cd2947a6e90d570405b3302d1f
zba904bf97e2b987ad85a2e9843017a1740b114c25b0026a472230cb4ed331ca0856c96d907201c
zb97ba2971e4206bde6aaf80b3acc7ffc276c8ce358b62c317116d1afa6a536b775a9aa7badb1ba
z1bd4577bc099fc69addab8bd785ca378457c07232f33b63fcc21c5081f11bb6f6b777e82a5bbf5
z8374399aacd32b86b86382f23e338ec519922c2e952afa7edcf8e6763ac02f2d5cf9727d286c24
zdf13bc9507343c9d2832cdbe1abc02c5497a2da06a360c980d28b6a5b83cd62f4d061d0066ce66
z33d7d477854bc61e2a9b9bf72119004409127fb26fe995558bf6152c03077a4161bb9b62e24784
zee6f1d339e7e76e80773010cb08ee8115bedf56fc31a12ee6e78c856e444ad97634e59176e62d4
zae7abb75238eaf282f570d53e41ef5d03de6b742992410466439559dcb28d2fca33e68bb793e35
z172163999ccf5dc38d3624d9d217cc9f4280f2631e70980583c1c24829c3bc0a73feb9eee2770e
z0930908427af7d2c9d413bfe589acd63a01ebaa53aafb50abb9f2bc3ced187da3dd8fd656c4ff8
zc822ff572ca5a1f6def6551b238ce46f3180b60e4a681dabd2c30e20b1aaac36d5d23da99e829e
z89529267ef15a7fa633fc5c6cf09aaae5b96cb392223726d79f4b37042b7434cf2e85a5d243525
z5adc8543d7e0a29da113f4b81c4394fbe432fd5eed10ec28279931addc6e9d8b6d063a87c9ba57
z67d740a53c9154ce2c3b855701057049a82aa7048c564b7def630f7958fd0858974289fe1f8084
zdf6297ca00e5ebd97bd82db181f9cdec2add60ee782926cb8f9f7f1cfd53f56750d50054493ccc
zdeeca2f250b42078984ee954aa80dd1e32a860772c7ef9160911ab1b46a11a63dc876a6a19e603
z00be83d88b88fad56335d9f92ab2fcc72b40408bc368710210a3c1a97b1b1e12305149f50c5e6a
z6636174300107fe405f4c6b6a0996e7623c6f163867fc1ee7c75f27f95df4a10718111196d0ce3
z56d6299e599ada74f95ba3083b42cdf85b12324a39db61babffaad0c4afdb5f81ff09de3707ad8
z412eff0170cecca93f5f341c02235fb08740d4a9aef6bbf6b5dfacbee0d829f839ed974fcbdc73
zd1722b9478c36464bf9578a5461b7e5964bbd21de4b279380b3c6f207d5195d24c05484032206c
zd659ace4f62c23fcfe250c0d10e69a77ef890ee208b83292223bc211b67178029e0a95d2a1c7f8
zb53cb317edbf7a83134a3544a4159f4d813b0fc74b6b5f9d778e9dc85dce863e93603581994c6e
z9fa9a79f32e136d8bd253450090c72f9709312c0296d3af03f4b8fc140152b19e2bd459819c591
z1d4fcb13567ac556b04890e1e7967195c41908d7273a4a52a24b15a008bd3b2200a6a32d484429
zab829118a05aeeb3b151241d648cebf5ef0e830e28d68a2ec63de37e028efa2b99ed915bdf61e2
zf922f82e0b512bf4beda14c6885725a98235e7cdd62807d1bedc517289f65504b908a138bf0274
z2b77a0e6c599c2a6b071f30f3867d69b1cf3fe1c1855a805a0395443665afa48b298fac1237f2d
z29c1e1628d26c65b0d03f4c4f0a61af7a37cd1f01f521a9ed9d6ef24d4f6d678a9b964f9b455bf
z81fae9bf62c827b305b50de2708a8c69ede4d9468384f91a3d61798cedf87d8645272f8ee63e8e
z810be2fc6330307ea3b2b9f1d0d674a21c32696a6cf40e31ebc3673976b0eb4b86dfc0a123e2f9
z9d30e9eadd191f86b37035288c032f668bd2585b43c3944fd3b43944667b14092427801babf5be
z0c29fec9efd5fb4283b56139788fd6c603dc1930b36beffaa2bd5238d73f38eb27a09262651c3e
zb2cbf8f1b531282771c477fc9c12a5eef57c3306729aa39656bc57b6ddb84cab1a8c8d4488f53d
z91e51c22ffcd7d0c9ce25fac05de7367e2d1fdb4a1e8c60d2b1e3de0674b692c33dfa252e23f2d
z9113aef9be347c7a33f084751473c56324c2cdcb638023a103a3f2eb0b7e3d43b6fa5c824e4d38
z87fb642af6c7d69d6701bfb07e66cfc5098d1f75916eff0fa9c122d24095a6e931fbd386057a93
zea0bac7259174c8a29096691c1f462d1bf9dbcd2bcab2d4aefe12e8a7db21cfc96c404ea7d0285
z76fc4d9397e4005b28c53d5520be7e2bdfce43cc738d49120a4c5b4933167908e71864ccfd86c8
zf5dff64eb5a51095b8aa2a2ec95abef958bd7b87fd843a28fdfac35a5b2f05515e33aa8e88e283
z3bba7a1983b0465d80b52f5cb807fc4808c8e71c0363a9b3147552f2a7d196cfa66ba1fd2eb98e
z397ac7005a3aebb11f3b3495413b2a6fbd1ee85ad7b983b8533f2c38d947fc8c59c455bf1e019d
z4409d7507b9a4fd1e03cf0ef507f611f728ecb30882e63f5eb88d5ddddac917f33dc1e63a37b7e
z61381554d02087662ba5a83adf2f7e8117080ec89f2bf4918f9db1376a7e06c22c692e0d31f836
z308628028de389ce09ead5cd7be8f31a4ec8b0f5431eace457db13ba3c3404593ed644b27ace56
zb789bc888501e2dfff20e1bbd5bebd94f631a3607214d7ce36a5ae0ad1cba2900416f53f6b4757
zaac3b9ff2d994d0a6fe1cfaf5ce646f5abc0cb9b55353cc853d521e696bed1c819ca0cf5ad8315
z71eccfe8f16d31626b6d8a92cc9c53c68cb7d3b49ec5e77124d406aee4e7b4ff970d9ff8d465ba
zc6889537edc2003086bdc7d907bf7e192a502f7ed87e9083ec00a3074964dec42be7fabd6b56f8
zad699c7fa1ef0f8383974e2d14182dad81f5c70c8cea5719d2edc2264f17e52dab7d50f167ca2a
ze6fadda3d71d9411d92423df91bc7d655d11f4b0ebe27c2263202b54b96eb03b567a736b21a913
z3c83d9e06731c43d1f03406a5a8a73665a71f571192e92c5b4936bdd8639fbbd045da666d69710
z40121c9c95378204a9fa1c6d424b5ead67ea90aeca7fc33d88b8407e3da265412f208e85579d87
zbb41364cdba283b3d1f4ce521f597618e1cea783fc9f5e8061c148ab600e5da44a497f3a79c2b2
zb4a7b69417bfa652871434171ae8441ef65d1a2a25128ee79d39973630c5d3193f67af77d4f02b
zbb7460e37f653a43d150194666a07293f69b14ef524a590291cb6e7205bc0110a29d708118b3c0
zbbba004258c58faef5ba2ccdf7bd735cb1e81958c8d51c849ef5ebda3b35db58041c285fe9d650
z82057b7c456addc1e19b5e423c0ec9ca1d2bbd65932dfe375cf017bc1795aff37e0781d81a4da0
zec70a6935a9b9af3164fac0bb2662897b1da5c00170df4ae9cc5fbd4cced556404617bd24beb05
zfd99c26a11f0650100fb0a7d33aa1b8ae7b316a0df19df6fd9673555d03392b0f984e41cdf47cb
ze2003074c3b71eec8502ca76d68f8c174a0a354a6acfb7f50bf0f0c5c4980d294d9eb625fbcb38
z715feca0fcda879e5aed58d1ba7b6127c368cec646a1fe3f99917f7588545db722c546a40844d6
z7a29c1ab29f309fc82048bcdc253c5905aa8d3bd18806106955eac8db9906e4a10cd4318aedca4
z2a67a1d21336449c9a4e997d2a6f0624b1567fde29ffc1e16745acf220d42f2c7b9c4d2c79f778
z73e9d3a58f49d1c944181ae54ba08fcc7abc052037725cd45383731e76f6c3896de21c37c4b39a
z8b81d5c76d4afaffcf6eb5d225f8c19b4ab03c84762ea86996636b5f1d81617160bf20663635d7
z63ba7981a0904b22467fdfb64c412c6b05e28c241709392cb76ac73ac2511822f1c3f79d4d99aa
zf52216487cf66e5602d91e457643ae9f5527374e641ef4fc2cee8abb54928127e1666c0eb78a28
z4ad8a1bb9bc36ba5e7d3a881d47731a972598ec62514c3c2ff568b35b6d870379ed3f7e89b1530
ze7c2f86eb445c1f723d3fe208612c26618240c85064d3077fe2a8959880441a6f21ade3695f12c
z64d95a5e455068e1b90965bec32001d1ef8a958f610ccedf90141eb0ecbb1971e1ea0ebb7e0dfa
zf20bf0061fe6584c30b569debed5ec3e81a66d07b61ad7f0a8baa188d75505a219dd445e762d2a
z3cc2a769bf6b4a0ea31003a291ea6b846edfbcd2c96e654430d88bfd7a33ea9533c012ee900e01
zea9d31a13ecae79b1015f090eb9fd0ec29059818807cbd319cf9e220fa63ffc6574a99f97191de
z6c859c0b3b2b7612cbbc6ae00657a39d6f7d7b3da6e061cd47eb5cb9dec17dec5e3e1c1f1e2995
z7a4678818b7da77e81b420288741462371780a54879880122ae55ac200ab65a66cb73423c6168b
zc15835527971f869a39ac458833fa0ba8e572da3621f5b36bc1a3ba76bbae91019a25a3f995a32
ze8933993329a8da75e5b2125bd4b199c90161308961ff9790c3c65dd10d875f1b8146f383f5af8
zf69dc5c419d5fbe499ed6ffe6217ffdc380d1cbbb0d527cd8522ce3e0fb7d37c18607006fec962
zd42aafd70f503670c0ed79d702a6ae044968bcf67fd21bfc49a585176a307fa67c17c25635535d
z8b134f33e8bfa414c691cc2b20212afcb429ff472cebea6552b94c9180f6a44fb471ff77838a70
zdef02c54d9bdf9374789fa4fe9034dd90e7dcb082e91cf0cab06e033fbac750bdf4afbad320e8a
z02e4b2e404b9ee836dba69d9517eeb65e944f74e870ab3046b830cb11505757504e1142219cbbb
ze27707211cb5c4970f43a0c316ac4410e8a829ca86cb6df27f8c9b4648a071b7c67b60540734eb
z3a65d2971211a93822dc1f7c53b56b9ba98a9251965427e61a1920b6a1927d9cf0f1952a9dd0c0
z8f142175afcd9017b3f37048642c85c349d2b1f581bf320bddd44e83387134994d94e1b0a15e83
z2abba672442b772fb7d1b1a90b7364a02b93622b5236062b53709d6b16b3c990ad28c77714e526
zd24aed6e035758634f000640347c5d7122423acac788c03357e1aa2c805bf967e6ac6bbfc01c8a
z7f557681455338fe3b4df2739740fb443660afc75fc40bb6f3e38ee9d8a43e7180bcf4dc5c927a
z93948846485b86c7a125c4b9509c2ed5950cda9d31456609b3df95e0232d9511fee7bfc8eed775
z33716ed5620c8b22bf9a83c45ec03d96a8c7cd8afdb27c7db6d502307e4e764bb51302e73cbae0
z703ab0cb5da64dc5a07c8deba2fdd16bffc9fdba35721eec3883aa69f344fd02444214ddcf3893
zaf3efc33107776a5030560257062cea923db99753fb8f0522fc12e2ed98121f24aeb6b2445c81a
z505738a578b6a1e3d652c4cf799fe98368c09252faadbb7a2669996ab51575ea6fdc0f181b7cf5
zdb9d727ce233e277b89f3a6f0a05c05dbb5ee8598eb2f7e10fe8d7b59187c0bdc979954f78c7a4
ze3c3ae4875d93fbd15433c690866444373b43bbc170c77a361aea3c9edde0fdfcfeeba20f8d773
zb4b5a62004c48b29b747b7c30cac7caa3c4ab4b00921edf3849b6249949e4d8fb1cb8be91d07a3
z3a314b5f64c36ed4c5aa31088793a4148f082c47cb4cbb65291f2534e0c64dcf7639526d06818c
z44835563057e43410e36f01160e6f9351d0236de45a4afc8681ca6ed6febfd55ffa4cee53fda48
zedcbfbc95de18fbd0904fbd7441f3eef0e4130163009a768080e016aab60b957b7f11f43a1d2d2
z278d8c4ab8728576bd081af36113d1896de5b479a83d65350be2f178df3cadb62c4229192ea455
zb526f0207874ee615d4f96b419fa6c76587bc92975eabd4965270d17c3b241fc1c121ea491136b
z5a0d87223b85f4d36f76ef11dac2a24f4727c8f40cb39ea90e997f95995d5afd0c09e2f2d3c7cf
zef23ff2df7b334e2f8900bf7abf071fcc28fed1e42a0cc1887975db9021f24e1f123b2b3f259fe
z4ba4cc81a899c04354cf218771e65e26ff37cf9ba3c182895f94bf7d6ec36861eaf13614b0545f
zd2763d6c3a158eeb9b02c97cc3a324a24c08029e22c7ae88e2714b8447e5abac602a429e0c5821
z102d1fa8792904b2c4f5bdaa4cf9dd25e6c9443fb8584b26195edb2f843a120330e89d510c1182
z07e18fc3be7556abf6f52a56a26555ec3298bdb6cd89822a74073bfe3152c65dff4ddca5dfd0aa
z00ab677094cb204d8a9acef4b7c777fba641ecf32ebafdda0da499910867670dde0dd119e5c8f2
zd71cf7e83d7f2734c73dbf42705d366b046ca292e3851b45a127045929db4728875b672cbeb562
z0e37f0beb43c0d458698dd7277b11a6c88f8b5fb93e2cbe9068304861fbfd37a4a84f6bc54daa4
z4d8a0be30c7655f4048cf223bf920260c15502885913c389c3554ac7ed6f943f7ac01b6fbf42db
z1034d0a1ba637395a0fcc74323762b759eee97596340aa161af55d21923c55a209025cb57a8cb7
zad664b0ad47e85261252167ce9485c278635cf6fdaeb421d2c66682fa45608e23ea22237fa2a30
zba27b8b0d342e5e1dd2ccf9ef609aa5ae580faa697a4def5d766ec8e78dccbd8a57458531853e7
z513f428da6531dad2c7ea2039f809fdbb29b2c302e7fe67535ca059f249f519422e4f1aa710aa1
z63a2cd4939b9c9f20f1bcf23e0a046eb93977d2f9466806faba6b24382633fc9465da2a75f6b34
z470465e203d9630473eb0959ef7e35133382ddd7c387e9593139db6b9fbca0287e52ca093ab198
zc6d0d3b8ed5b6b55174830d51a733afbeb74bb5cff3e66b99caad4924da3888704ec313630a29b
za056c7db9ec70e60313fcbac86ef5aea4279206c26b964cb5646cc435f42c36edf6a0c50da83ac
ze59cbd311474051830011da590648b986087d300d67f14dc3d35214ac0b24a5f44ed3ac1d70516
z03df7dcad314dc063e32d9d744dcbf4e9f578619e00a4e22a8685896a31eb5f91738e078d2330f
ze5d46c33358c32e84c7c828b9dda27498fac098910855d3cf9f2920615c73103a3ae5f55270d33
z5875adb1bb94396100068baa028c0c93d15e2a4c2417eadc19461c8c1e20cd357bfd44b8e762fe
zf6d530ca13d893307e3a132b647a4240611a8894f74d04834c61eba1d9de48500225cf901b715d
za19d13b61af0787dd555b2dacc91d08b8b0b1f47f0fadd37a4f4e81c95e5690221fb21536e4ff9
z7179f0fde94138284801b29b2f79809a821fd6f34c6c350e8b2c238e548b23e08aa82dfa2beacb
zced10b53a466ea238ec986e76b1ee03a65f58b4f7708c859f926f438b57620bc40387130371e0e
zfa83aa197489ec345798ca621d7249b688b648791a9208c207d9ef023a8b978a4be1431787d91c
z4ebc13979f3f1fc0c1b8ad9c70b7ccdb488f5aaad8938b6b3cc4b83cbbec571d4b9099066e0f79
zcb7fa788a0eea0ddf72a2ec9b3c56041c9fb0903623c5f6a6c87cc1393baeef84a9cbb82b0fe4c
z7c059de704fadab80c7c5cfa4b4deeb6cd5b7afa6c1be0a1813fb61578d687013c0c76c867c083
zcd2fbc6e1a878ac7defeb12f7d86dffb663a3e5b9621b40d5f10b5773d9123723e3a590173510f
za79a7337b4f24397e6d69fadc40826ddd05560e8bc4749693d3888d0e7f3e0f82050a39650ea26
z907168b34fc7092c4f9c5597e92e9ba5b4f165896ba7bf2534b7021e25f430c114157bd1060e58
zce8f3b4ea8b7f901e1fe04bfc21984e458a8f53e67cc8741f34557759bc5203dfbd35288675720
z22a83c1dcb1e9de2530f1c85cb99d6c6682b865f703eae6a98be75ebe292a02f6eaa7452ac51cb
z474ea98be1b443a8a8f938a32467af02966cc91c17b878a678f602b35d0367e94bb14f193ed88d
zfae192b292f560c20b9d91689627117a52e1ec64163094a46d2b15163b19811c022aecd00f2c8b
z22bb037c59b7df4eab64119bd9797ecd19d3fc9ef36bf751d315810fbcb594e8f506780a438708
z57f186f729f8c8df03dbc0505f58cc2eb5d4c3e30659bb1bea1bc45daee11600cead22c4c260d1
zdc26b308ecf32806e1865630718d6fe5dc282c7869fd709d42532ed93c235d3cc6039822166f8d
z4e9c887f02fd5f862170463980b7c790db63c3bb211628c068012155654374382236f7d1384ae9
z474f96b858ed84717fa4fb9d4f132bcba947f21d6a951f3bb8f72ce3ac9a92ef800061fc9c82f9
zb735a6c49efcf5d8ae4670d2aec40af867f6114a0c186721d06a07b1b2b5393197052d24698f6d
za83be8ea92b8bc561ed41f653388c1a2b9573ff02c36556f312cd4f66bccecf98968cdff96fc1f
z64280b9bc9691070ab8296ec4ef6519fb577f320b78ce7d5c5d2a1ce266bdbdde48817d97388b7
z63cb502c8bbbc6b084304d114a9fde3d3b1daf8f86d304463855db32cc055c3194c26c63011011
zcf868b5a9bb268e2ba2c35b4636ddc43dae7c3165efd83c5c1ac623d8f8f700f9879ea60ba798a
zf8b8924bf5ebc760761cdc27ad5f941e36c287e0c54d030b2b7f81368d9f31120888aea133fa80
z342c267fcbdbe5ddd47c1212c18376fc335584e7e420aa07e94b7ffca4f5bb27e50b336fd4401c
z32169ffae7cf7eb94b79ad576762b6ee3e2b17e0103d523f8639e6d100e4c6d410800389408200
z9cbe67e2071c67787215ca55060223cd0175ed51da6e24e4c0f2529faa4e9f8ad6cbf4646ed1f3
zf0588c10bd37a1ca8fa07a8045ed55079c88c1481f845ae7e2ca2aa847fc4e6be26fe79b6931e2
z0ca20616dc09a4b8ea786dcac12602d87affd429501fb0eeab0b87230f82b9b9c851374f4e9eb0
zd55ac3f8dd9f0c43b38f3e75c7e90c76e58cc8a9a1a3e2f0f0aaf3aa72cf392062b63455663046
z7b0160403f6595aff40f5038aa67badf10665c41417f105cb9b7c0654410c0b4726055f55935a6
z6d0ea0213a9713df80e696a7eb36d9034c4ea55dc6b7d57c6051dc982435ea006354471ef2f019
z75adf7b668d44987ef38a5efa3bbdbd6a2d602e30b1b367fc376e39942c26158e4c4002d53f2e7
z01a037169753b6e61f19451d6c2e87412be9aae95f0dd38444d53da253b1046ac99847ecc73dc4
z2da19d63542dc8525fbb7eadad98a6ff34cbd343123df9b4c34dcb7235c0278229499503648441
z88a5ea340d55cad184ddca261951ae7a777e853855dba17dbb477ad02b074312c7f7e94c34ec13
z7b1ec4ad0ca561e66c677b34ae04c9adcc33ff0953d9556ba26572c9a66e61f1f9fede2249b86b
z464f290dfa8d7523c658b210d936f35fbe300d1ef0858b610e093e1976e4d5f119ed1a2923b201
z39e19d18a1a5fda5782106ac8003a2f31a2e09ed8463aa61ab07f09d1d9143f17a957249330e82
z7f9cd007d7bbcc616a29cdeeb8260e55187f0e9708457bc5b8cdd3b36c2c8d9957972b78924c57
z0ab62a747f37e698c8edf54efc192e0a160a165f8d2760f1da560cde9ffca79edd688998ee89da
z911ed0e892d6ea7c7dcddf0f6f4f0636bdccec3a4950d754c7f23f65e849858381bba00062ef88
z133c93281ae74bad493f5aad3b9e7e6396829c2810f658a2f564f21ff2b7dbb6d371433c2d56b7
z6c8b07b8b2bd723a7916c7a1ae367bf4f994939e3ab2466789811d4096b6eceae7e203737bf9e4
z820459aa4f329a34fda15b3ac7ab96091be7ba05f9bce95a446e69b2ba1d822819fd2e17b31bd7
z1c7cd05de3554eb35642f428b7888c1ec9d53bb7b9fea2c08b7c6157fef902fbbdc06d2b4dd76d
z9071cb12c0ad5dd152c015922da3ea99d2a676d9e4487a0e407b378f29f3e6c03f68a83cca0191
z367489a72f754612d48a9192411157daa1045fe26203c24a569cad6875f189dc6d325cd9756e3d
za7b6ad7e236bf60097abc15911af8d76b5f04aafd4f481757ad4bf5b9fa2a644190dc9c1a1ecd6
za0cd0609e989c42ca690878b2278302c898d2aa87815fd1f8a6afc650ad60295e4b218cb467d44
zdede1c43ec70eec898620eb50242829826181598922da0e7655486b240414a35613f45104df18e
z6a51330ee3d52975ea873f9a3b437a71e40afb60e3c61b15fe03633dcea84ddb819df96bcf703b
z8cc2fc56a8bf9735d5a73feedd8b695177e508dd7e8db37981f23932644c60abae7643b62723f1
z1cc57f46768e380fb2eba71e9415c54f9a27a2dc2ed2a6abff56316184a4fefc9d1e6059220f14
zc5a1c01436a3615f75120ff3f60ed44cfc623dca41ce9ba29e5f6852ba3c783b20c06449c9eeb7
za571af22361e7599579f1509618b276687f74ad07207718a806868550156531a7474d39de8f2e6
z5848c040a3b91cee2b55e5e7e60a8edd1058fc64e0755db45fe150893014280bd6ff08a88d07b1
zda4a01f948a338d7fe74ee1117635a48162b874aa7c452abd11405cab2595c3113aaab3ad89109
zb87a7ff834903f3c163a2fd3af36c3cb96b0fe7f9c17704571d2b5e4991a3108ef5ce394bc4f0b
z00d586e3b1f82fadb90fa6462747d98c29b2941f1eec4395ea4adeca9e16a81e0ed80f8dd08cf5
z12620c3659c71bfbcc56b6ed493d524d93805820410814436792b54b89e5ee63cb6e81f7639561
z417cc34270bd9e5ed3c5a15c168695715c317f250491787f83e4ebfd5eadfe3a954d8b3464a987
z20f949bce5b1ee141cfac70664c7110f25ae32dd6c529336616025a9be11f1fe0ef8e7dfedb064
z2421aa27255e24bcb38c55455da52fcd0cedcbd98cead664172d4b50dafb1aebcad53f4f5487b4
z43c11510c4f0748c12302d3a4a90d495f41d48f990f3530f358e2561d4e73ab1f065533f43ec32
zee644999907dbdd1a59000afdb7ea50694c64cb5be14e6c6a2624f509b62eed8a03c995d217e05
zbdb5f36b964d929deb1c9d9a52b506c3d8ab04070fd38bb53dada55e987ab015c7c423b9109b3d
z7db0d4b0653d8531559224a3ab83ed675a4af79e2835fd789d499e9a920485250ed4ea69d79a7b
zba2dfcc3d8de6b062b589063d153510f926467f55df1aadb97ed88320d63c6bcb1eef63b9969be
z09492dc7c71622c74d70ae4cc9c882bd6f5ebcd12cd04c1a384ed40f689784760f2ba0f90284b4
zf39122eec4e07ab5ebcf79a1f5d7c03b12c6601e6c49b15e1240c5a2a2f712d1df104b01d851be
z64e772ec4bcc34ec22df29af428728544c74546ec1c354e54a4ae30442b94aac6d30e02dcb41ae
z0c3c4ec930098b753773ad381a1ac6e8a2c97ad84ad1aef1a46f59b1c9c9189be0f4229a53a82d
zf1d93d77eac19a177ab5b246edb2219a6c19511e168e23bfb7d73197d28c140e3216989aa13654
z8b250163199d69c14a1f665b0789f378b05c00f644c851b1afd79206f1e57a56adb419f81f4190
z7bf598383b08aaeea42792142043a8038c53b4c2be086ab6d22eec53eaf337c43024bc521512ca
zd30bde1b1d28218918c7d82f8bc4d09cb31c8dca470f91ffa2c3c0b8763451671064ae91d374a0
z341e88c18fae1177b81ebe66b1d54589201601748f43d0ac795b1c5787025f06964f9c1159f92d
zafe78bdfff4e571180010a81bf4d5596c0648b6c4c89011b23f71d5cb1af410bcb3e0baf08c2e5
z18157acceec779b8d469ca18d582ce9b218ddc4a996d1f3211b64ad5f6d9d307da7c6ef1686b9c
z9d61b5acb67bf8450db71e4cf0a6802454f4c7192a88a93e0a1cbb19385a52aabec7efb462d766
zb5890544e9849035ae99c5ea2ed1df6cbcdcbe4feaae33e442ee0be15f14a84a8f797818c8e6b8
z0b87b2fe0004d16696cf7728218daf9ab7d6f92d1b0d099a78cdbce1c6fd362d6ebf9bccc51753
z502ee6e8609509e0d563bc3f1e21e9036ea04a41d2c16efefc43de4ff17eaf742c6ac38f10c79b
z7eae8e27b137c11833b4f00e0a04ab739f40b9c800c49db23f4001067ddff843b8c0a48332f575
ze74f21d8f5078ce2924bda38e144e44a44af669684f5f6cb2da71ebb14bc80c84f355c406fa789
zb5eaf5ca58a61ac61d9f6bedc8e1cddda53d2682a1156a9c16e8634ee58749ba724a844295997a
za16f4c22f33a067865039c8f6b52614c552037f4a614e39cfce3ec18bbc267e20e1112da919056
zf44c1d9a37f758c94c5b89e1a3a02d064a77b5da98aadea604bf03100d3c3898ab4fba409e4c54
zd943bd6d727a8bfd726d14ad99a26b96233b94f10f8e6a45cd869746a48de5af87704941481b1e
zce751e34482b88d7ace06d77bc2f93bbf0f67fbf6b086e7d81eadba88b15202fb35eecbdbc3675
zc2edad0a3eec66da2a2f51b435e1dc323c9bf9bc2e5c6b6ec9bf2cf88f0077ba892464cdf13aa6
zc67139d19bdf19a208bbca5e82d58c6b7994e5d41c5c62ab3a823310479fbeb1433f7510e24666
zd61c137adc62b21b5aaaed2fbc31d38fabb16985a3de37f7cbdc0468f007f9e959636f3e82e46d
z3af5f83214aa9f8f36b67fe5634148b2bbeada262ef7b5170b5812b2518dd9d6437d9bdf91d9a6
z1ca46f4616bbe81f123fe24dd823843114f56e5fa4b2609495e6a08da3c82647191bc352dea396
zfb8046336b10d59f58d844e28559acc18ba6d5ce91b9100109f9be2eeb35b0cc23f61a76f9cabf
zb0dcde7ed88645b15dcde1a08ebd54e37c6d1a67b32bc89ab4fc1eb4d0796c1d84765f786d26ea
z02d0164af7d4124e0d4a331bad0864411eb3c7a4bae69027f7652ac5b284735a8fca2eaa8d1e88
zdc02b244d97ff0205252353098cdaf977771146bd6930d8c393ff96244b9a2d6f9aa4079b5ac25
z3bc6be57b0d1821f6d5b7fa3b65feea984086d25ccc13282fe8b7cc376cca3e39f5482c683fa9e
zc0b64ebce2d48fb57ad113ac4f7695bcf3b9bb0481e92c2c2df3e7af9f2881c316b6ef67cea8cb
zf6fdb4baf01c701fbdca38c3993fdadd0f367099077d55dd98b58841c3a4117da0deb615f4de7c
z2b207191b8069f8a3469b8747ee1da2f9634d4138efe31fca07ff0768955f2f49d08860492c152
zc4d1ce9f3284f5c6e10cd741a25a2e670d608d86288f4fd67387e2e6ac2aa3c644737e51eb18b1
ze862cc611baa2223d1d34faf173407c3986af8028eab266b36f70c0912d28b3463c8b7ec3a27c2
z9ebf71cf25baf1b6ff21b3695d6259c9f3f643c588b390b6b84bfdc938f1485641d12e5342018e
zfd476405ffed2cca2b39bf7607523ece285d8b400e73455c1431a47fbda73cc80f9bbfa31e9081
zaae161e91d9070429fa41315b19cd8be60a3e8ee95ce3ae215ceb4e845a97385e2b965eac42056
zd2861fdd2d2aac4a5be862f38b6e0c13d1c1f6dab832206bd6bd253c4b9bb28bee6ae76e031bde
zd2923ffbb6b61cf20c841800ec9c97ee059ed98b66ed4202b3faf6537b4545f9e81aa079c824ed
zbf289c47f89322d2324c18eefeb53eac1f9f99992f519f034b61d6ec05303879d00c8a65563867
z2cf0d74909b5200ceee589049f66112f7d0cf58f20226a90f8e0d162c29a25d9860c0f43fc5576
z2845744a5b0e8906ceed8e523893e2d8ca65df483ec9fc12afe72d8680d975bb52171c20075460
zbff7667c477d4ee183eb45129293ff8997aa8d8a16ac3e0cefd285201bf63476aa5d883a7a915b
z30db6160f5972ae1d6582609a5379f8a93daa6bf70793154d889ebcee0292beba5505838047833
ze4fd5127304a2f21f1d09588545c7eca94aa1ab383ebea1dd5a8510cb3bab28e5386a8985a844b
z192a7fa0c3cac903603a3019b3a31d517117f3558d9d1ce237d954b6e4da1d5127776df95cc8f2
z22355194f45bb6291801eae7b08a74906144a75ceff9d5874cfa99f653c31a16017569761acf24
z7a4664e204fc00069d4feca881a7011626985eed107c18f73ffca68595b012f841693adc8e2c0e
z7347b13ff085e3c091da09dfa5c08bc4dc6deac4828196bc4b3e42f0ad5178af11d8bd06b88125
z663cc09fae86837828a71e39f2d9355103019ea7ffa55eaf736a749cda58661fa3dea8e362b759
z203603074cb3f44feb241577e23f1c2adeb5470a0f89ad9140b4722a3a66c10f413715b16cefc5
z5ef0220e02d9bd2c8629aebb0693932812de4d09379791a6c95c2238e7e240b07e93ec1f2df65b
zf0ea594045381791bb531a284ea8d1eec126ae548746b6db2359631864e1ad45510e85a5a3bd92
ze80f54602fcd0edec015f9abaa237332523dd140d9d0b22caba46f41b7e7e79b73a6db1c223405
z1ae0ed59d6b92ffd3586f0fe18fdb1b60d50a539f5820bcba9256b5d4ba1a4fc75d814c03f168a
z794513b6f524c74fae972fbd5c751511c336158b11551a7fd931d76f98f325db53202057c8cf4d
z11aad9495bff5e604a0656c1e8a1d897348c503f0ee806f04bac463ee6aa3475444cb7399e1e68
zdc272177e89a8896f3e4244f5b588404bb48dafa15c15adcb82a295fb7128cacb2fec32e192446
z33be2c7e8f51802360525fe43c8c4d17f26da5b6dcb650971ec4c57e3de05dca388bef0b6fa64e
z99940924e4d381cd7265f673e75836230523018459efac282569531288ee4c14ccdec8ce197e5f
zc9da4c48292d5c6750404e2daf2f3ac5b8f8dbc93ed9f28c575767c389b738956fdd9693a79799
z2218f9751a9b2936e23e74855b7b3b3f7d7ed3689df4d6b27ecc041f0b74830038be6aee5a872f
z9da23fbc1c38d89da91a145880655765f74af1bb8d78e358a04ec493045f03413679b024867b42
zdd6962bcff54a705be202dfd7642220d352737db9a0c95aff24e3fd9cb390473d0bc12c9b1200d
z83056e13813025c05673a582ef236ecba92f45c1338cbd4abaa0cf34f8e9532a11c2a8f33e75b4
z1b5972e4b681b179595607d057594a4a10223fcf23083d81dcc7325a631bb24b758a69bf0c6307
z34c8db55b99b182593574e4b868249f23e997b476d058d836e2c4ae54e4d295d59459642c13cb3
zc609f305ab7a2daa2583089dad52198bb85859033e8f58415e8944204263c19094f8ade4a1a755
z172aa1995ebfced4a48a0b602549b9907574b8a1273aa8446968f61a3a7cc97d4190e13c5e87e0
z6d555a274d115cffba1c9b40ce6ad397de210a0a59dc9a7b9eef11c4926fd4d10692878c69ade2
z1d79f576460dbf40625d27d92d6d67c91e070b954d23e0e32f2e1090c6b39e735c6764d04b3265
za00dbb630f4bd796576b845bb8e97869246fc62a6510a0078a40b2a2ee3df4dceff5a4f3ff8ad9
za07720508059b7d2725145895f81dd246e64cac1418d93e53676af12cbd9a52fba4e54f29c3522
zda75e7cb5e5e8e2e609b5ecaa6c890e966c6a1cb71182fb4258b676b386d54f1211cfc715cf39a
z6b27a6286f663e1f8dc8a55e014ecc10186245b38d51fc59787dc2e0873664dcaf472778a4e2b1
z3800a32d0625122e3498c7683446ed3f6fa026a83044f15e51a7c857dc22335a37809231505bcd
zbf1680e64c3b3c6ecc00cf82bfd303bb303f76242c578d08918e4ceadc5f2fc88464771d7aa54f
z1bbcab3a92d9a591de897bfd79aca3e27810a84813ff285dabc1bab02c8feb326625285c504217
ze534ca05aea936256d16f5dc7baf43305bda81e4e8fe367912d33323ba4f45328c0633537ddc10
zb81461a39fce5527afbd8e5010eaa71accdf3fee322643af0413b1e88267f730a8dfcded7def1f
z6ffdf78e0d5e3c6b995497bdc1b6a45c881d4dc4d611f30db180c7f1d788cf5c2c67b3ab2c7319
z3807ad2369e44790909f623ea003f344aa90c03f5ab0747ba0417c578bed8812d19749e775f7f5
z8fd4f56388162be50f602503924e6b9e6b16bca3d23d56b8d40e96aa6742b35f70aee45cef13b3
z45b6d99275966d1cb91fc879055367332f660d323475a2f4b5840733e04ae03088f5b9f233d94d
z94e8317c12f6c88145b42abab79e2a0888147aea9dbefed7bc45e44f01f989e74f63ab1dfce3b5
z8fff919704a887eb63614e0de06f39181d1bd25298c4cdda15df9c720783a7f5a87a52d53887fa
za32d6407c337fe1871cfd8b8a50edd4e317ace53f5ee452f5ae187e0120b6067b7ce4a6b113a63
z74ce4542581e7344db59b2ae33f2a306554fd4b68a01e3d7ebee1a2619708b65e9cebb3844bfc4
z60ccd4b947e8d56abaed6ebd60151375c4db9bdf8d71e9e17c70b3db8c4f5d4ba4ef13120f4529
z32db7cb5b4a6a46dc70b7ffce9be8465bc9ae85b8ed31e5439f541733c42c90e6de7436e1d6851
zb0b2a5b1ae8788e0723aab26e4237ee41dcc7534768bd3ea599b2a2819f0ebaa04f0c3319f5e39
zdace2a51230272716b79e9bb90f6e1ab1af1f6fefb96ad57123a1251102ec099d378a45bee833e
z2f5f9bf69f170c874c47ade67b7ceebc48ea530a44792b9fd9c85db286436a5588f6325d3d6e5c
z0700b4638dc2cfd26ffe956a43eb0f8900c47d6c995b27d41a50335180d8baf589762bbf178263
za053063ed6d1c9dd1ed050a34c7217fbe3ac014fef45739c383a3a96922faeebc5452d0ff6d84b
z19e0667e98216566150394a1a15698200faa502a25aa09db42a65d5763998512bc14f904d54ef3
z6654b53b5ee08e855690f466f10b7b83c17c0cecbcc2819126aef044732d89d3b97cfe9492d158
z6853dac39cd8cceccd709781e4a0b732a151d86d8631371273b9445ac81951fb725f9e89627106
zcd704fe462651579fbe9b408bc7c5ebdb48ae5e963e1bc004a7fad56f8f66e5efb52c50087ab7d
z8b19a9213e21940f8ca589932749d9a165fce6bb66d95bab08d6fb4bbf6892bd656151bc6a42ad
z02a3168b3b39116c4d0d96d8197331eaeed2fa94b3b235aefc1acf45bd531cf8e6bd944523cecd
zbd9342a9967e0a0d1b4aeba680fdd42d9a5d1407959e2f7f8b50d35ab590c254bc4da96909ef94
z597aefcc1aba693d0dcbd25effc3b3c1b593e2dbb7c002cbdd29fa15f0898eb6e23af81e4f2db8
zd6805decc599acd61f369aa2ff9dd6ea1e3684f3695402de82517f25b2f58051f4adc4fcaf685f
z190787e072294b7e85ed478920792f122e72a897948b589e1a82c76dfa3ed44cf6495e00cdf25d
zc5b20f929c347f697ab884def808103abf6ac83a7f32ec95918c74e5ddecdc41472a25b69a0e40
z01962188a4dc604030342303a4b385c452c096be3dd5052c800b20cebb73b54e7f677a449bca61
z94cede3498e1b9c3f9252c02d7bc4bd7dfd630c02770e2c70ec8c30623f1274429760589c88ec2
zd95a6440538e0273af90bf1754fde50bb989bb88ee4383abe14956bb943df7b41bc7c659ee54c7
z1baf413d87be28f8a9eca06840d16bac55b7df4537629f2108cd8cdc8e02a45730cf10e99f0197
z9de2737a41900d1303c5a13f93b2cbfc48c148d157a05ee550699f514cd0cffcceb8b7b3852a08
zb58f8dca1e470369ae07e568841442b59d9fef5893a1599b928e63883aa877d7e0a3596751ff22
z68d23c70659edf99767ceafd72143ad414331eb5a8bc19f19321ab0f1cc9e47bbe4013430e3b79
z4e54756de8880bf95c03cae89f41196ce5315d84bba52d5ff0906b6a813755729716c21f62cc05
z7698b6eaeb7a481bef75d541a056213c268bd483db7b2b03e9e4259c6ee955efc39dc3bc8b6f72
z283db79509d3361efd883cdbe14a8837c1977c716cece03f1a0eeeb38676c5ca3a5b46c295dc7b
z02bd81452e723fd897d3137742e8d1d21c06e89fa8ec31e44b1500007c213bbc133499b9dd8da9
z1e2f23185780c70ee9d1fff9292ba1290291435dd1637f44e94abfe156562092508477ef7dc871
z63942c2608430e3190c1221c6714706154a87fd7afef5771c5f6e8448250e8057abfcb3a880a88
z96399cbc709b8eb940bf2ab7a408a4180932cd2d7f85d6f03eacb87dd9997809deaeee90388889
z5ce23797f741e7014cff38ffadce9716473b4d3c05fcb1fc839978e4bdacf83ab7bc108e6e6a70
z70cd9e5fff34b9e93f765e5fdc30ba4e8821e4f99d241f2dd882faaa003f393c3064000e60bb18
ze437eba499f05f08e8ad1b9e5e629a8f1938a30cd0e4e0981a22ef02f7ca9d8f7a18392e2f216f
zefc58a96be94bd37aa5a74b0d916a485d7487f9d4ccba44bd87c71a0a558b01b252175cf24c7a5
zfd62058fa2e011a80e2b643c6418fa07ae06f025b1dbd9fb8d5f7eb1954f0f8a5879e8791b9600
zdeb3c8481d2e136093884e288865d7fcae368b7f7aaa1fcac192803d33a74648030b864c720702
z44946ed09a3692322672ffac4ee4c8e4e95310b0620ec4c1a1865e8da2a3c4165064496cb2e7f3
z415e9ebc67b08ffda41412e24cb004876d18cf5796045f98ab8acde9fc9fd005e51ced7d036fa4
z035f0e665acd17135956b4afb9282dd5d2409d20c5515b7977cf541bd44ce42f6999b68aaa5715
z6c595e8eedb09ce4b7f7d520bca9b93e7041aa9b0d5ca5c35e2390181f88757c2cb0c18dff5b27
z8aa563e1f39f0c49fd2ccf4f8ae059aaae778df340dcbb739f6e5f1a80b0af4cbdc9b15c7bde6c
zbc65091a956bc5af245fd3df395ee4c30aa78e812115f0db168d070dcaf7a85f59ff56dec28d5f
z607af441f2d13d2f283b096cd0292af46476257770318a2fe283c7c6de260625717fe6979bbe76
zcdb85a9dbbcfcabb0c4bece3e80c79e87fbd18f46783c9045276e9d2525e565367b3dfb4ea1c4a
zf8beac12159d282ebd311f6fa47e1fdecd1e7b04da6104cd36ed1c63b90918a1351865f9c99827
z056d829f2dcf6b21eedbdec27a26249a6716cc51531e56172ffa4ee5febd63c000c171741a9cba
zd5eace69b9a3b6c04e45b2360580478ff1719cd53e44e5df19b5d0485d2d348dc2bf55e2ec3bdc
z5a02ce6d114c747dc52f86a0a671a23a25b05d433fbb188bbb2bf7e468cd616fa5f6f1acbd92d7
z75c76f7017b8017ab6dd2ddeb1ccf2d09517b6830ca102e8c2c1eaa24fd7745ef803f66a24ce40
zb9d9fd5238b621de7425a1ae547b183fd80136d88aaa4cdb793b5919abf4e33e8458f4c800a700
z341d231776862b12213f3ac8f1498bdd9359ad37a1196aeb8a9a91270d6d1ed370ef713455c00c
z7e8c5234a33157ddd109f8f2f4e7080b39b0539924073bc0be32023d4ba2cbcd0ccc127f5a6cbf
z7de27ba9e8640c84125fc7d7d59d4c4beebe820c65d5ebe0c959f421d364d2116a4584fbbca064
z8c9f45eac3a4ea00be14937c460a5e5b0f8851fff92c979a51221d4eca2e0c8690f3e7131898d5
z60a882ec4b23820ad211fdccfb57a0f6cfa4f27bb1ba814c04c7879b14bd7265d3c602da426d50
z7b49de7138a97a1a5ee7923b8e3b0b3308ce65fe1c9fbcb9a2d26e404f0ef86779e1b0cf3c934d
ze9028e57585f1051cbe834b03ecbafa4f5a2e612c0150611a4ff383ad00ff742dc2fe2e308a422
z08f628ae922eccc8aef78aca7e54400dfa83329c27d2e64607b06f11a83f2b1a48e6ca87c27207
z425c85b66f2ace35552924c0b9f8c232081a07d3f82ab40e177dd4d982897c9b00e3855bd9fe70
z2563a191769fc5e23e0895973c67690bdac2df6dcbe1a63445c37536c77a33caaca4ebdde80ace
z2e28900c42c4e49083fb2d50ed3206be0534b14e8b1dd140d48b6fc14598848269a69960cba361
z51b0c531ede9ce14c606d388cf46f605c425760f14a8e58945af94fcc13a6d43a2505c5a0f8e57
zfa774479f48c817483b15e475fa077716ffaa82eb7d1cfc491215a6713a27fe9315fa29257c24b
z27fdf123ffbff6451cdb6c037000fde1cec634e116219f08819d487932219c0173797143348670
z6bbfdd25a9c98dd8de2fc0221784def8da3e7dfa194e797187f1d97786cf37a55663cb40f5593c
zba2d4856843172e44dc55fa6719edb1d5b4e5063c15d100b037d5a52977c64a206509c2aafca90
zf8b45d91d567aeceeee2953b3794b0a50c3b5035e2f21669bed78671e0b3046039f16c31258880
zef0ee207f0b338794a6630971356e694adb5b59811e39ff5dffaa63851d7600fa362e27d82bcbb
zfe10526a6c66fd95aa4bb9d409083437e1fc4daae878f06b66f406500cd47693b135863da19a1d
z48885fc40004c468aa446959fcfd73428a257eabf119e2fa4a57f4df23695df7ad5aa78319b43f
za0c2bf5d3ddf920b1140f54b4d18d37397ff871e6e0df3775c667cd235a5c0c2ade12bdb000343
z2c13a6a58109be47bc70d914f09cff3c53f629f6b42bb6e4ca795aac55c63c21a214b3e0ee0738
z755ffe715ef9b93099a2bc21147e322d010f9e35cbfb9b2f83d652aca07e6e09c455b800db3a65
z0abe63735aa220901e72f2584b0e2862e8e8f167fb98f1dd10e3e3a45689c28ca34a2477807fc8
z7642c19cd10d5d52a2f743b0f75f88858c4b34380b0f3ee01de709603fd87bd1da400e5b8463c2
z50dfdbc512a1144930000748c3ceaea2c09770f0cc17a2082e63e056dfdbc1870e753e4d60cb26
z3cdee2ab542244ce4b4b0931cdcba1b31edce3aeda34243accb8ea9c1ee6b2ce59183d19f28170
z7e809f1e35a5275642e958f8e8378962f876ce6b827643c5a1e772a9708c9d1944f48fe1d5eb7b
zf20adaf1836af8c450b1be4ec0238b94778e2c84cb18ddfae99871e0d312fe82e1a1f389248098
za87279ab50564f59f25f3d4ed97f2e374e2a28aed7375aea4dc1e94e9336fc980b4726588577b0
z656776dc48619602c290d58c8ae600ac855fe02baeabe00ef46b829e89b1af1b0bd51c7fef9283
zfe9bb3a0ac14baff61c864bfa16cc98627aa6bcb9543869b04ea674414b14e70325229f9fcdc20
z1c56e8eee4916dd1e881a996e47b84263a404c0fa8443134b85f7d186389cfd9c504a1b835ba98
z66387122c3337163141b8634dc6f47bbdbc3351c10b8151c10e8f48258f4542f42d511dd704088
z2758a21db92ed9576487d25ff2d1009ca617efd5c0b4d793d0051e36683f1076c288f6e695bd63
z1ee307c443317bf8af8bf22225807496e7cb999e1a52d14176e0f6ef46a20633729620ee2dd11e
zce9785c4db827b0de6a994f8fd939b2aac08192765a295fc3a65aebd0eac7a49e2e1e31c3b1ee7
z911095f3e645cbf07fc62ad06a1d9576c58b09600e23f3e73a895a7aeec555a19b866e0c8602fe
zff65b1f463d1f8095f2559c4b94613006135caa45183b991368852ea8d507f6f6be9c24becd5a1
z13f6bd7fec2ecbec7765476358a8b5dc65e29d7bbf84d51c03e4a085171a820fe4f9ca887c4424
zce7182dd0ed2d95da852d41c342474bc5eb2d0714aa1b0f8a882c041f27df6ee5f187602fc2578
z72fce686c48ffcab6d413e61fae0c3a880c9df5bfc2f09d092aca59fe6718c5c6619c4560189d7
z5e1999cc8f1242b2a109e3c4301ca521f9bcb7a9e6e3d63703e6a33152c0b9461cb30abbdba644
z295cec715805e9c0205df5fe9beedc4ae37e7459c77b88cc7cf1e3bb17ac9db50389ab4508026e
z00be6a14b7013e3a8ee915f06263b7ff4a2824267ae02f3ef94e502ece9e0ccc8679a9e824d47f
ze43c85b21fec50a0ca420430906ff3479178f5b26fb6e883ef06a9143a2fde1afb32e5c455d053
zfe986ac08532493f08c03b1118a013bd2b89bd73245f5965191aff210773ab72f0721cba9d4a85
z16d864731f596d2647696616049e2918117a64bccf9a6ca976bbbed14ae05c817a3792a17d42b4
z0c1dc12330365438ca764ccac3579012cc40b15972fd215c2b8b184ade47d73097fc59f5cf7e09
zc775cd49dd7e1d5bf08dbe51d0dc203900626eb526bb8f3dcd4f3a5336fa587b5f8dbe3755bb23
zd804d8a1ba136794fcb345d6fefc3d5fa55e3ba998e6c8fa8d9ba3f67b2379ae10a85b9aa5d844
z624e930c131e09d5654cae6fad49e284e75e7609200befeb8b49be4a955d882cbdb4723faba49c
z4b609cb2afe12474245af3d0b115d07f91c687c112aeacf1712944610ce00c560e169b81aa24df
zd48f5a1f79b8b99583d5271dd036f144715c70e537ec3a456fee0d319dbbb7730725985079511d
z7ec6aba37681c0c6c82430d937489df191ae32bb24f40e7a4905e3dec34d3688f8202e788e08ef
z78d9e5edec68a4e79a9e212c7cb9efdcd8fc638779f1b5646a76cef247ae6ed10640db2e18e85a
za49d5ee5bdaf1834791b87aa17522eea26110f6b998d08772c995800691d9bb99a1f37bf2e109b
z81b8da011748727b5bc0641d5865c0bbf858f75922127e1611ad5b1d62d31816d88a37e8aa3972
z2b4bae82b5da76ba3d54a889bb8bb4150465c67555ebccd136b8df8a354c55341de7beaf6ead0a
z5cc5ded1d0e67abf7e0aa09c6bd6cb675c8b948be89545d8e63668a8c0a10ca3d6d60c201b174c
zde02b0ead0831c29b56fde094af3ce828218bfd722542e75501f7d680404d78fdd804e2db0d0c5
z84bfc054ebf4e06e4ae8b5b2ce510de35682aedf0a35dfb0b9f29174c1af57493105fc9c0e0eb8
zae58b0f6854feab2c4c5f7dc1b6a26029d80f8564949eaddaf3beaaa898100a4f964def091641f
zd363186fb7b645472a4170a28d5b62c75c8c7ad19bfb02030e777d82e6f9efd7818f1825f73ab1
z2e65404f8070dd56822c1c9e537dd4e509e0e834d95f04022bfd611a0228b26df05f264ac042f7
zfd48671e74dd8e31a50dffbe4c3a9aba17ae7318ffb065500b2c5178e66999d4217c744172f39b
zeab31fe09718c608332f7fc878a91591eed4bd89ac5345d37ad59f14024cd65413aab9863422f2
z5581967ff24849ba3dd1ee37668e53514ac012f938a6f78be81c78ea06df795e8f48411aceff74
zc5e51f7aaaba366905a52eb62e141c048b313262e05851066238e0246c6a63fce2e1166262cfff
z47028b5fd9a1f65366dab69feb1fa9a4cd663151a135e138d5f2a855ba862c8d227a6c7b651573
z25cd5828e0bb93225a40ec9578cfec872a1cea50f079ed68f83ca4d2896e4dc1b83c297a4a1fb1
zb7b630dc7c3f7f23fc9acceecca2393ddbf16bb5e54ef42dcf236d4e866261f209684d8f736950
z9ee99e54e80f7688d591988c1424d306e250c44820d37d30de82878a3d237ab706b6982aec2c59
z04a5ede0be131f1ca49e8ee34a656361e387c87662f099934c55978d1e9e9494dce1f49af51da5
z9d64200da5a31021c8b70cbc0998d30e64d177b71d696509e5b515dd49126cffba5f41d3fd848b
z4518320c7fe844d19cb562e22be4b9a2658e9a47365aa23b2253b7fc0d6cedb7fb5f8f4eaf0e8d
zb64ad5df0638af4021c7ed585fe8564db9294311232dfeb86cf61694a374e1fec3cd2447f5f762
z5d89192cf4c4840f5727003eb0111ba1b13f10144b4a9688733cd5e886dfb2eb84c4f4269df0f8
z248c27b68f169b9474f216d8dd59a046d607721f63545ba348fc607b54ca84524b5dee9c51e0a1
z15a2542c284deaa14c630a5c63bea57df7721aaa8de6a494712dbdced6bb39ec291c40c049fc18
z433971cd776eecc78b7cfeff84e30fee62297ab60008b019371dcfe4cf0ecdbb0b5810763665aa
z81aec95ea5bc05631f77c1f3c30f7b5c48382f7d533f247d80edf9085babd51e725f4644a74a12
zc571dcac49061fb39cba5a7f82a629c9d9651a01ad9af3d7cc3853acedcd0466630ec61261910a
z84091c82d39579e10e6936aa3cfa019ea6c7fe994582f1a9a0fe02208d4374913ccd96edd5481e
z764ce3604e1fe9b323cb888b3a9a653bd50dbcc074853a5a818cc86bf80309134679e4dc054d5b
z43da335d262056b257a56a9dab626d8c089e3b143c020efd45c38011af8a1e5b7a2fac1ff95f26
zafa7405259e5e19de9f819cd0f89021b8bd9950754d0402391c2f3cdf0675b22a68d0e688a92b9
zbed26f654ca9343a84c25217cb5baf9a3766bc5d247103a8a89f8684b4cdcd776668dc412815a0
z3da46e7f11bfbbca859334d06262280904d5a3751f11c78824f4cc02cbc74fccce153a18eb9dea
zb089abf8c2f29995e13480983e4efb3bb5da3fca0cacae6f2282be22b0a64770aeb70a1cd1ee71
z778a8d0f350fa6e4b498823c3271d52d5874df37f35ea14e85fe7e53d831a3aea3e0fb2f53fc84
z4c6c40ced47cc199aee27c242e0b1be5e20afc3e067f17aa3de7ac1b3d047cb39726537f8e50de
z44f09b18a6ad0c102ed10c9ae79ea6c5cefb6719987190d8ce032ff584c34dcf64a8f5bf1b9988
z4ab09a1ed794e1f61ba5593d6a0262f42aca06d94abf45ace81bf1f6b1b2b4ac69b4b3f2605072
z346fb17f3cab1566b408fd7bb97a6019d239ed0cb3d5e773754cf0a9e7c06301ea6b668604c3af
z402b4d6cd78a6c2776bd50a674a8357b05caeb65c12bc2dcaaa1367c818e84cd3aa1af9e463415
z22d5b7a0f78eb5922f1fa00102f9fd1de299287532657d1a5bf0d092d26608ed4bab8cfc98a2cc
z706f63e0af37182fbfcd2bc46531c72ac9a3fde35d5e28de4438ac509606f58092ac1c8577fb7b
z4b9ab440216583c6f056d373bfdde2b2b52d549d61ccfa65fd22adc16f7e1d9236bc898f3962ab
z07217fb1dabe36792d0d0cc010476f98791461f2d3223a938bc3f5372ca0f496ab0507473207f4
z7a08599cc2a341ba5e8bedd5a99030eb7ed9f982166714fd1b7ba9eb3e2a229386b161ee232a86
zbeed85238878aad70ba042aabfa0bfd2223b5b3d3acaf2d898b7d5fbf3f0077257cf8f942883bc
zd3f81c31a7cfc7bd39c45b576d5d4b163c1f2a157f6e63c2e655ce524aef8006df616663812504
z5f522f7b68e1d0149f718cacaaf7596fd4efeda56f68ad29eb2693794bdac4634ca12b8512c4fc
z53219e864ba93e7b715e1a2f889b83bab44f9e53c970146ed1719a9a7d0b4623699a49171e81c3
za39f17ce028d6040421813b9c6a70f9e52ef8e5472518906e6ba1bd91f1b3dba37a0798f8546c4
zc18124946bf17eebb620c4941f3b75739cef0d0c2f5fd306e4f15d990ead4eaa654d4069acc3c4
zcccdead1c8eab71b27f70567818f16a5f0a88efe577a38d342b838df78f56efd121f134008e847
z35dc2399f498f5e4705cea2e23401de548a5da545dce1b2c4df11e42d0bc7cf2389239512f2ab4
z62aded5dcf137e6b60a8919dc1766830cf84d136a5bdd51d8b21f8bec15bbabb9f5079101a44d4
zab293883240449ca3127b9d7d54e3aed8b940bebd88d5e35121c382ae90d46e79ee7edf445653f
zb14705a3aff307f1f99e8e20194716f008bb6036a1d8cab8ea6ade603d0e00422954c007d1073f
z1a178c9eb5ffd0043f155f69fbd27eebde31d411f57944c52f97bf0c4b75d19b005be0fdbc8a6a
z2763cf0f60a5b70556662294323b4f532ea6ba64ca9267d0fcb87ad2b7fc5520ca1dfe6168af83
z4cad28a81b29f26b934888228c7bb752491ce4d810bbcf75c748e7cb2d7fb6c5ddb33e94e5ddc9
z03eb4e72569e57a4d8a6e1822004d6a8f9cd8cd9c6ea60d07ebf124e81b23f61ce3f8f25767436
z20efaab898be3df2fb58d3085554e441abf27fb0e2acdbe594e32eb302345c5c407ea64fbb6fa4
ze578628b025f955478d9fb6f9520b455f675ce32a50569f3ecc1be72ed023f5438f377159308fc
z2ee6128342f0e380d5f70699d49bdeddb4391d4f9e1ac3aaa40447c5fd3d3abfc49e8df96c147a
zdc310b90539c6b194c5fb14291a3b54f8b9cb674319203ca6db928b904f84eba13f9147e94a571
z496604483aeb02bdc8e34a81fdba91bd7efea9702a424ad84f64fbe07c6085b080167d6d06deb2
zb0574c2b86f0b93b7764c42f39854f368b6c464767dc4d4b0941b70cf3c4ef2a87a283fe57f48f
z3894ce5f43bdacec4d22b5a903bfabf018bdef8688405001fe383e789697d6408e059bc1c3f323
z9e8d99a0904585426a3fcf29a34c3cc2c6ff781722be7104dbc5d0f8826fd1cf47a37bdb773c07
z3fe2c3dd2bfee9f659a57292b5e6ba84a8121ba168c4dfc1b40da1b6ab5c91c5a296eb7cb9582c
zc6997ba57ca67caa83a40de27d3a39a152d2a71cbafd2345be0a811f303201a0f1a899e0ca5982
z6a430ce863e7c20e3167645e20bdbb4d8b5890d736dc3357308e093c8be487c951a25c42c4b03d
z082d3faa4367c7e487a5340130eae2e29b1e5218b5ddf5005334f574391ebd1fb02584459628cf
z1ba0ead9159195a671722bb3f2a50c78ad2e992445a19f91b3785b5aec45d983e352290e2d9893
z9be34106f3753ac91af09116138a7adf62d171d1a1fb397e5a1655248479d9898e2ad1d0652afe
ze44e71737402ee6d7282c3a45cb1d07734a59e20709b915e7fe2a004694b67c0360c6158392048
z6ee3987c2b4580f237336a6f91c4b5d2a49fce39e88657ed1659da611f9f3c87e6866c62c8762b
z945b8a78ce0e3ad04b380601f02302b56129a0c72adf56f0c4e57abcf0cf8b2b945d5ad7178c66
z6f87553f110d40b8703de48b131948061338496501d4b02ec50da2a3be8ecee3a5a5453b4545b0
zad62354a9a0cf465bff2961a9fe55a2d134561d56657a0f4971b4959da4cdc2106b4b746b34e60
z1e882acaf2936a2ba655f29b38e84a6938a0461f72da6a859b118f103bc6095de979b9c39738f9
z0606f977c072578462da0771beefb3bbf06f146fb0a4f1c57b6fd426ca2aa20eecdb58e7e56b3a
z6491ce6b0e0146a89dc9d9ade209a66736e9ed40859e9fa8824e0465df33ce73e84de37d2c8aa8
zed246d33b750b853a1636da6914795f0cb013024ca579812a83d25a968385465e1478922f1b7a0
z63934aad427eeb96e422fda559535afdad71a44bcbccc68fb5e99b0a18d35c8a066ee6d0374fdb
z443c715cca5d901ffde668227ae0102b2fb746f76eacff42dbbdab25521bf51e3bc8ce4126c7c7
z33c318174748c0b1e1c3ba93d28093c820cd2b2f1ca6b44163d6a22b4b5eaef37763cd5c225e5e
zbf2dd48785cd281c99d7f6bf8f1145da56d8b4fd85d84d6284c1ed31e7e3592752defa57132bc1
z54846c1a121e060e06dd7d87f6bb24c0f6148604c8579fb52978c42648500867c2de6efae8bcec
zb3281d368070898d986170681624a06f2a8b93b17285a5b41cd9ffa26ecaa61f683c57ff5175a1
z1f81c8ac9b2166b7f23e4f661d1e193e915ca61124997a38597cf863ad23904289f14344cf6f9e
zba3df65c3728d4a80e8747760d199a6397b957c0397749a461ed253f51585316c598de6e53bfaf
zdcf66f48be24860ee82704767443d982ca4b5ea86d3967a86d8dbe69512a877415106627f4f102
z426c5d36537a18f70f47948202a9a16010a5f9bd84a0f54e5e9f6132543cf09645469b51d5f173
zafe248d3f784fdf75444046f05f99df8077b3e4f1149e874bbb99c2d041a62b050df583f7cbbbc
z435b414bfedd24761d4ffea9b88508c6dff7458b9776e2d59c5150a2c973f567e2a76580f50002
zf720ed1ead12be4a3201c9f211e8c39a981c95322527909e4b1129b4bc7f40a0a9c2b37d93205a
za7660bc033f50d6c0a24383c6cd047dc83a4b871fd36983d0be397eeebb83f18d16a4ce0c05d24
za503a24ce3be0fdfd459ffd879f8df120e7c1af7b47e84e68e7b8ad7742460925939d479a3e6a9
z9f1df2ea10d2b8a181b2091ef3d510b92e0cc0a1e3acbf82637fa56451e0c1ddb6ec3ecacf7481
z934eea823a6951247550be50681d7c1ed2c358b5976414eeefeacba6e2060b05befd9fdad3b8e8
zcde5dcb18e2f2fa7cd72d8a8896706cb75731c3f0a13d169a7d5be35161e2e4fba3b38dcc9b865
z10124aae598b878a1a45296b04423cad32a915fd76d9ce68355a41f55913c73ffbe401da39906e
z93a90153e6e56edabb6c0f16adaf9b2878cff6e11a8d98a43f0c6681155c45dc80f3a74c37cac6
ze4383f70978e4a3b6fb5867f0b4b78d7da37841a40f30bdc3bff38c19ccda3dd2ef50545de98db
z5d02567233b3042b329355cf803f657bc528423dd01fba73386b72524477e8899ae04eac2ee013
z029b4119b631f31f5903a55b3e4e372588088e9ecb64bbfec0b92e10dedb4e666b93fb0f07f5cb
zaaec0921e12eaaf470101baa64e1a306b4e7e00f5e323c9a4c1dcdaf07a7157f1b2a63a113ea05
z3c05f28c0670ecee0bb6852d17050a0fd7b5e150a91cf7af56cad29c2b5317421a0d301ba1ca32
z8c4a4e5854c51b7d7edc5321050f90079b7e4e70772d7bb7717612cf10c1e95bcbef16462bde16
z19eb29f8b7a4b6764a3da11aeb37253f2704a4ecc32827af1d7734f74dbdbb01276848dba0ce82
z9c698a646399a61cb1d3282f69a69d6252133dfabfef320305dbb6d4d2bcd13fef4befb6de4ca3
zf653e4709aaca028af9b844ddc3c04864db1914909c163b4fa8c42699c836631db7c363f18b6e5
z0efaeaf0f9124efc4cb0a996d5d6dd1caf8cab37b790e693ee02d365975c047d443dce1cb4a331
z8750035e24fabd75ad517a8bf78174ef2315c82a4b4cd975bf9830e66447a8f531c729886ce038
zcfb9f5550d221525bf0e1c37d5fb1f9970083256e7f1d5a83510da74790b9f18db6b300ba4d5f6
z1e7f65d3abf0ef74c77aa927471ecd7cb74660161280f6d1fa202e76f8c93a32dfe2a4b69def27
z884b38c62c83b842ccfe439e721e6b22e50a395bbe4011a2b1ea8cd989942245bc00b25043b531
z2c214ab2f325687f3329c17edb208eef9f6cc70c629d4d2666a8ad22318a9ba7a41d33f3adc1a8
z341240e8b12fad22f01c1f9a5a6985b73ed3b5db4d439f8ea5c947390e8a1ef07c2cb2e0af809e
zeb574dbc443a835bf3cdf0a0171fe1d6b569f436153cdfb2ce9eb117335ae5fac560108c44d547
z6cf5879d36c242b76b8786a977ca007e1a323eceed34d11da630719911c7ab27f87842698effd0
zef9dbb2365d3f47ec9642a0be65587b3b8c2cacdc7232ed4ae9a92a5eb6df6d379461188ab371a
z5b715f7d85154ca4fbbb0c1f37dabb549a02d0d87c330141eb0d94c27d3a6eba8c23b90eddf367
zb09132756be7babfccda0bc56622b714f27b5db1b02d03115a39fddff5283353ab85f102a1b530
z0306ccd7b7dc832726572c7664cb5abd962b83469ba6ca3bbb20d4c72a255140b87ddb234393f4
zf8fb6b676e39285741742defbb33b9f7651b2e00027e914243bf49453b27fa06e748212a85cd67
z24b4f7168a270147366b844f4ab0adc5d121074c824fbdb7390e5e1c9bd9dd32ff964e99e7a4d4
za610af7694976d8adc7af83c5a9b60187022e55504317972e8b3fc12aa4eeb14e75fa1da8b7e9d
zc38607652315b85344e697e6374a22ca89b1df83b6ea2355c64f12500be023803c83ad54549795
ze672b8cc4f1e1ba168e416e9463f004f7a375eb79fadb670093d3daf5091b557acdf899d87175e
z8563a48ee296cdb2623c03367da7530ddd31597f719996835ea2acce5885d588cc0fb2f65ee494
zc624ae93d416aef1aa735dd54b1b680d1f07c07dd3111c61d6205becac16ba5793e10b8c1b48fe
zc3a9714d68251ff92e0f1ff3d00a360ef839c58a84e96d4ada22d61ea5736ad64a252e72ab4add
z6d88a33e982f8baa6749a4f7e9fa099cf7551d7d5de031e1797f476e93c608e86ded4ad37efccd
z3a26dddb7e0cb56b4cd82fa059b8a5b40b459e3e12e48ddcda7e2f5a36ca0b250b0f203d4a4d0e
z3d70c4ff22d97bf407c6f16fc0ae417fb8a50079ee9bcdcac676844d910ecf1515057f059aa821
z1a637263f134cc5d4126994752bf1b0846336f76fd7bfb12d26725e6d7423f6cb351aa4f434a1d
z29441f40de85f2c6375d7e6124f553fd73ac3a796dbd8883a5e7d11b4b3ef385d55faa234e5b3c
z4a0aa79e516825d4a1adbb6bd615534caaa388db36e78d1ce1e5eb3dc4ea4ea4af8cc05da2dd99
z7546ede376d39d42f582ff2ada12d932cdbbf3f0cb8ef51fb9a38db9276afde797c5f09593126e
z9b3b661086fe919c4eb489077541b49ead2eb08207c6cd08916a1f44c8fabaf76b30e9dc846308
za6edab392e5717c36f2fe8d66c43c6ed7111c22aa8181ea7e5b3827d7d3ae0de60985cdab976eb
z63aa6d649f4584e6261e3b2af9b909d03ac3c4c7098a2d911885fb9c01c48d5b048948e6ffda7c
z08ce839b7670301b1066ae67df152c14f7714b9cef9061f2d55aedf4d04008776356f84a6afb6c
zc7f09ba4d1621f846485329732a6839cc3a3c29173cb7981141adc1420cb9b16a894c36aa19512
zb445646ec9d90b439f33e8636280cec21abfb0a859a01379110b9627df27ecc81a4b72fc1accad
z95c984eb3b883c8463a853724bfcff715f359d0fda7be43817cfcd5a022e09a273714ec2993167
zbc0b3c779fe82f41ab806fef782b11f83665ed5f6ee0bda1a37e8b3d92ba863f6fe07b87fd3849
z71ecbc42ee915d5e017f05892058a4ce207c478c363847214c54954f03df158317e9c9c18fac65
z433e128b135903336084e0d52b65b550ce79c5e3f6b35fbe4cc41af55c3cf6c12d982e5d4d602a
z7944bb3d1f1fd4148b1cd5fcbd3978f1e0a347e7cb0e04966385bc24a53395905c7061e7037f28
zc90b8d645a4a1512e6540962fbef6807a348eca43ca8d0f641916239bf4ca9730f4833f536789f
z51f97c7bf67e86c94d1433ba2ce25f247dccd44f00562d6d1d8da657290f2c197c49e862dd6a36
z232dc72323c2d3ac3a5f1d155726bf07cb1eb6399a9393dbd9c14f9eed515cb93586afa90b8c31
zadc79047c670e1c97fe27743483758ee3569882af5b9859a1e1f035e8d775ba4fa82227c8b112c
z40091ce69fb05011a93979c6a51a1ae01c24096f811c4a9ff1e3cb03b9b02f0e72272f7435d115
z29f4c361b1cceb1dfcc3710959a06fae37d339b5d2fc7d2b9bb589a1d4daed73e73d62a87b4995
z3768bb5ff0ee27251804e82218b19f861040c9c97b7ea484179ef5fcd31a5f30e0adc7f94239bd
z92e4c64dc30de451a8855af6be021023edb8314d7dc4173cd6264e640cfd4c7903a220721ee3c1
zfe275aa199dd1aa77e2a719d2e7cec20d7720d3b7624008f3b83cccc16e70cd4876d03c97fce8c
z2bc86d2cb03d5684ec37845a6e08b6dd79ea94fe5954aabfc5b3e89b7d16a561f3f2a324860674
z5ae3e4034b292ab1fb5a08d7ab38b68d24cce104b5bd56659646ca0a654396a0936c0f229d223a
z9cb575ab8390916d037ef5febeaf1d6dc7a61543c79f4584ac11f977940692ebb5c8c18c3e221a
z8a06aff57e7aa097cf27100c961cb8ddce13436fe9e39ca2971ec164ea1db9f7c9c191df552c5e
z0306032aaa35d66e557c37cb733f0cabd8e51f7149d09d2338fefeee0f413a87ab4fd066634c04
z75645e128cd141b03ea1c1306b672a4ae99fd29f8057765bfabe2f5efef8b37cfc61544bd6225a
z6b7cd661a36cb629eb4eaabd725ca1a3c0e1bcc49853d5a333716af757f804406c6278c4481396
zdd68fa96fef95b436c01eb647cb348d7e472d14ada0ce873a8ec6d4bd65a0a60df6c6248e59301
ze74234427768f3a06e84773631990df3c7e98c49938cf53179bbbee356ce242c46648b04a2638e
z94ea574ff88010d2178c4f642e14b969c045ce745c29365e340f386db3a9483075064a1eed46f4
z30ba50b3982240e3bf4bb5bd3076ea6a4900b1ded68d1c4e19ce92babb27cee8e4ed7bced6ea47
z67b5f3f22715ef66412d963806ff5e9beb60781f9bc9317a78f8feaed3256e2393165e99842dac
z364ff063f97140034808450a7037b43c157bb2d8b0b24981c08631409e3e06fc83e9df2704a91f
zcc35178b061b11bdb4643b02554c175e6054bfe5968c1582c1aea3f77a1d2f072b26b1efa7a2d5
zce8fbfe95213c48bf7eede5c51ec7040158b1067e4b8e9256b31c38c8563d234ee1428053805da
zd9c790f7364ab800f53bfa6c0804a5a55c11cd0d3aaea3e88a719bce9d0d7000051ac64cc0511e
zb79a2292706867c5f67e3b0774a6692fd857bb84d6bee990b71b5a490f2c4a836fed3c521a57d8
z5026fe1c61a569b92d7c640cdb5a93dcaa8de9e957ad29cf7cf6f6cb312e0e393ebc76a256d82c
z73af74b38aed545d322419a73f5d64b58b10424c61803a11c0fc707f4818eaea92b3abc1059ab4
z432ddf1710c32d7f05a851c86771a300eaf81ad65f20436524b8fbe34d1aae661c81ea8ddd2f1b
z202c80d0fac2fe16fe64b0775b095de2bf554480373072a8e0209037bafd8f99956d50aec97aed
z49421d9bae56d4d6530a8ceafaae1a10d8fb7c2ad18cfedf73fe8e31fe166e728d2f1c083c56d9
z49924fb5063c72d4cfbd283475d9e7877e3d4a332691eeb5080267c5f8227a18fb5384afc60be8
z8e64a6124b767e38e6420bcc4dbdc7fb79e5e58143afee7dcb68049b6dc843a2685b39421d2c49
zaa3dd60e7996f14ae9af1b0892c9f97f04096b6c7e2932925ef33bba824852743c769c6b1ecbb0
z023bff3d7c4609a71cf23dd2393e64117bbf58a24d59acc9f22bff93f233d334046016260cfcc4
z7c2370097dbd78fd6d0ddf889ceb13666cde837554bbffdfc73b1305ca35df1fee982802b6c111
z991984d598562be1131227fa54778ea97b187e727801543098ef651d8d6fbed8e848da5e4d994e
z38ac6ac6e2387be885aaa9a4aee28d74da6358288b28e810b05a82171d394d91cf2eabe6bb6ec7
z8e45754a94022e1a5a25a1febf705faae774018711ca40aca2a6e258c139b54ea8a2e417e5fe92
z94817269846dd144b8af573f6d69fab9ba34c3506392bbf482646b4043cc7cacd566bf85d4afba
zaee783c4b6d2c90f1f1858ff6dcbe70a1ccd01863467e85f9b11acc9bf472545aee5a97f880f71
zd1133a2698b347e58cfdb554faefac7f689d666e9edc87dc3790329d79cb449ae1a25c88e25e92
z7584224b40a8e423b5ccdd2e1e1d5db2a92a7a1321e388b7a007956cdb86c72e091f5c5fe46e79
zd07ee271c54276c70cc80c25965832b8c545193383d562755c4a5d326b7787629258a9215edf2e
z6cf6465993e1caece6f57253ae78e542c501f469a7f3767fe4c0a8053f45ce164c695945188b69
z904d5e5b98d018a57744b74d1ac2f00e9c984710893509c164192c71098a6cda3ea47681ef7de9
z7f0778fab6edfb579cebd7506553f26a89394ab416d1f63fbe0cda6e8c564ed3f1a7080cecacf0
zdad3c7c6b7843f0a83cc4e2a4eaa8c0996d0ceb51b2191b1fc89a7111cfdefd1866793f1bbc757
zc143a107069590c430a50dc5ec2faaaba0e3881b8637c6deb1a7e099ee7103b34f61987ff4b1cc
z3e18c7e0fb8b5dcc64feb8332d1eaef65fa8f57d6a2602bf599cfd981c9065f1511d6561d52595
z179ca650a4cce16e457729b6247007cca7c244997f3e88af79ef7bd42f8a8d1cf42d35e63841b6
z46776bdd28d18ba597a20f55df9a43c79b0bfad1320ee4c825c8bf81b093885348a3084a16189e
z38eeb65676c36b132dc3aabbde9820b15fbd76e51af4db2ea39e015c536e0f0fc82b9cd1b06539
z7cf79128c34bccb9dca14528d37abfab49843a3d87c7371afeaea8337884e12eb684fc2f68eda6
z61334be2d81efe206a6a470740f7619ea2c3e72ac3e3c67774ecd0bd7981b1074cb9015ab39701
zd9f82e5d0ac01d747ef1802ffe8bb5fdd9f98a397cf5bf3ebdc15461d74b13fedc96589d557767
z6fc61c60cc6faf4467080c64cba1029fa16c54d649eda10cc350fa7ccd816cbbc9a7c41db430b3
z1eb64e6e90324aa3df6f854244bb7dc89ae0ce2bcb75d2e6edc75fc242ff03e47b582ce91d37d1
z8afe2bbc27f18843840d8006d745bcacff7be1a71c583dec369bb0d1ef93feba27376c2cd07589
zdf97ed472aa7608c408294a74505773107ed79f7b0b6adf8b17bbb9c3f81ba8400f8bfaf8e0977
z112a499efbd7c7c07de29dd0da2503d5da0e33ccda4a623b504c751ad91d89e696ed571eadb802
z74c3a4120d204094fc726302f277bdf4305d8c9fa9af9a95a5a16321fead721bb726b387977e68
z3a8ab0b287c3df8f04c648dfc1c23a2e8c893a9de5b7774361ab16e308c448164965469b4e2aac
zbc0f9a3d0380dcce159df8311b39136eb4ad7fd8bcd4595adafed58ab3fadd72a140ca7073ab9e
za8191fe4b1657a0d872bc39f2a8c5caceacfc86fcb4bd53725477442e3804ed3237b3449d402ca
z388851ac371af8bd91f527b5dfa05a288fe91cb9d635ac3e340f644119aec4bf2eb88097d56a8e
z1789ee84730af6284954591e86df67c227388b6390f5ede76a9367a832eee0fb774d2e18cf1e1f
z7f778375243bbd5d42cc43fd4481031164788c5e9598896037727635154d8608495d52f40c24a9
zf44c9370c579c0f5375f1742cc0c6f3d164ec11be621001fdcfb4646103e33c466529275ef5d19
z77710ec22a8a51684b30fdff545dc7766a29d19545bf8ca143b78d59506d71f056eddb6bfd6e9e
zd03486fc141b293021670ae4e62da5f13d0286310365b186c8e300c15e23db67ae51cbcb806d9d
zf57a8e1879a708f089f492dc9f09b55fff30211c47a88da7d7d209d556198ddf6e780c912d9211
z7d4341c9980018a422f5cbd95c4f5995829ec61b53c7e428b5ad1c282c7411b7aa9dc339b376ff
z6588183229f6018989ccbc8c729db2ab30590bc498d74a49bb17945f3efbc46302770c51036047
z4f1c014d753e6f890a5a8bb938a43ca85627c863d1340b163ad497b72a9d6a9305046295fe7d3f
zb9ee81cfda93adc58ab11226babbd53ac1d6b4462196d77e77243645d9ce7092a0efc8d5c29469
z880bf706881addc3574910cc12c37655755e9e8cc05309d03506a12f2fdeb12feb24df332397b3
zcadd32eb6e9c37dfc12ef54833bc7d42a21b9e82a0aad62d5e69c67c97562d190fcd23759e2b51
z91ca4c0289c27707a0b3f2ddfc3c6b24038d919d1056952f0e04fd82394bc667308d1d4fc7c4fa
z9c16bd0377f3a78be16289e86026bebd99d868882eb93475353489bae31a72bcdb641188d34e41
zde1548ac8351af81ffaba89aae537cc2d1122593c9fcfb23e76c895efd5f620f6dd2a04d5f1f5c
zbfd6e5f72ebaecf9a0a2d2607fcf97260a7c9bd936abfc9ae9f13ac721656e59ecbced1df407dd
z77cb143f8f8e0f649a630179c1991347cdcf9dfc51444c64ddbf0c8ca2c120cc1f7bc04289f053
zeb753a5c43ad64185a8584f2da6bee90a8e4aba10cc7e22797dc5b7ecae2e41ebac2d080b2555c
z7c33534e22c1aefe7109e9a6be10d2cd5c6a3fccb4bdfe86c08c8aff9b100f26c52057f851dc52
zdf4c7733d95dd6f71befbe737c4afa00cb800c9f417bfda42053eee2f2c1e0ce5106734e17b6d8
z421b7109cc501ac043bc9945b4e31b3bd3bf7e58848e1ec02e8f777e4c6900062f7c9cb4a4ed83
za79e8e3ddcb4029b7e898ed7e6fe2b8083261196e6a20ed88d40d26e689de3257b5946695ed3df
z01c651c8de172ad803ace4d6144e52d55c0f03070101f3754ef1ce8559f0fbaeec599d380af860
za7c775a625b9c7937f69453c09112b01511080a84c17bf6798fdb54c9ccaab183c56bd430b77df
z2e4a3fc340fca4e8584d47bccc2561ca39b1972c5d293c807c22f2502878daf6007dee156ac4a9
z41dc0ddf2685e04ca8da9028876c667d7d654fd97b3e13ac26330bb84c876009a6002f5e622bec
z35e0f29402106c2198d5e01c37a1eaf1c8012264e817b637012d1d9e73c779916ea21210cf2b0e
z714092f9d3eb45f5f2ec2c197dc7b2e5f8060fe45511ed87cc308e83d2b12aa42bb6c035bee02d
z2acdaae8d2e2d4ee9b515431ac04b574c09c28165fac7747c80eef6fdbd36aea1f527639234b28
z55a3162912870098f09f0ca520b25ba95af7ba6f9e7a133bffb31b93eb83527834222b358d6ef8
zb4d645cfcf22859ea841d4fe5b841aaae02b7d2d70e1b2cebc7827fbf4b1f3704d3f6919453a24
z509816e2222a82ea1b44c4c54165c87a228baf400db8055ec98aeadb0bced4b1cb21d1fd2d1fe7
zabab39f5ca4cdc62a45a85c529e875811205f3883588320946b2534d232b400f3ec2a06b17ee45
z45fc260b29644c5fa3f64e995ce55c74dd89e61014367dd0911f3496f6d26dc454cac0e0294c85
z4a96151c8a74d2d8bce08fabae45819ef9e6e97bdde1cf0d2bec9230306ce196043ab22f33e8a2
ze458fe6d989c2535200ecd66d626fe481cf270c77f3ea7b463e4b3d27302e962b3d106ff6996ab
zd404a736f9bbbcefc988381c90a2f59d5949f2eb2fcded4bc3a9961a8e5a7ee89eb027a4cda205
zfedbcabf96746c49c5f3c22109d3b717d6413843ba25f2d650bc00c940467cd2d5c50b8e3884fa
zee402bc51390d712416d635d1b633e0d761a18002aad8115be872931948123e12fd9b56f5d7b03
z2aa81e2a8aa790f08b891a2157aecfdf38086dce54d93899f5fcd4871f46712b19a93c78790631
zd06ad2b62397f4b39d4752493d0e90b4a7480ce77d7adbf99a9c42ffdb602cb97f91db2f3fe65c
z6d7d1bde3be3fc8cd01e5b58cd99845450f431ac6ed075def208a2eab5463d3bdcc4a6551cdec4
zd051087c41ef3f6c0323c23b2e9cb35f760338027806a26ab27b69631e9ea8d791a134c4d43d43
z9fb292f00e141323ad9132ac80c30d9c78c48346f7431a7152ed7ea529574ca8af917e925f69e9
zff87776fc8d1cb1c1b0fb0586ae0a38829370ba495bd6fc0e7c093bf105aa69c785574989ca138
z116009493c94261da72ed4d1a2541c8d0cfe97c3cfe74eb6b1ac9a10d5303b8c7d28cba1631695
z6091c4da3b80ac6a5e1668f903f944faf431ac9bb3f537c2f0668129fc913f1e2c3a80739688ad
z4686a9c5957c1d85e30c1228c2da4a89c288c4e9bbbfcade5ee4acfd668c65415af1a72c7d7f4c
z1765a664ef7cbf2326764d867e3ed1941d148b5f5a4aff91caa67391d4c8ff2c3ffb3b990039d5
z7d4e85e0f0a0289460c265e9ee2056e97045cbe22b1a8be5ac227509d1695fdb4502419a9ff500
z39f8a5110439410b6b36d63a9849d09c3b4b0386657441540f82bdf4b4edd6805f4a124d9721e6
zad7060c44cab3c1c381ed09bf5022df47042c1883162667f682778ad2e41307744872f9ce44900
z208ec6a3d0cf185521e317040284c02b8a9f375083e7d55d4d724e392094d7b6edfe8b88aaf0a1
z658636c4d95c9f4ecae36f5da526c794a9cec224fa4460b6efcec3b80a2de6179b3239a36a00e7
z95b270ca114c414268ce7e587919b671d29b159c8d7209df177bb4efbdd55aa2351a614d55bcbc
zfb6285ebfb4396c8625d293afcadcbcd2fe2708de10e365d290770f372e13107cbb2c3f5e86f2b
z933515c21833987c0630dd5a8517c4b1f03b1830b8fd4812d4a6a0262d058a2e23645a55144c4c
z80d03598cfd1e1e3c29f79cfa1b8d2cc5b2b704b2c91fda5bf7dcb9afe7d75e43adadedfe712fb
zd248afde0a22ebc044bb0143fac82a0518ea44e0fa4c7c0b8d5aba6b91d2efd1e93df400f7a0fb
z26221fbd64e3eb2cd3907cc22da147ad44e8cbb9ba171916ca392b1a9ef5b2c55604ebe320cf16
z77e66cd5f1328c2a62acc82f7497c79c098b697487763ad23bab3662c728e0df8f90b8eb9d968e
zd7374066404591e2056fc4db8af5854b42e8dda44e6e5bb30efb79079587b4dc9c41cdedfd8588
z8479d220824cd1ae41a4bca73ec809f3866a89fc31dddcfbf2800584d49e9231d400c45088b06f
zbca3d3d16a0c43ac2df55cf91d4bdb3f4125bf3deb0492aa3a809c985329451c60fa326f2a618c
zefa966f7405549149d291f777a89ffffe8e1c6212cc9d6dc461fec9a8b3f716a9f12df1d1845c9
zadc733070f62c1c359c3219a664de68445d2728026c9fc98903b9aea21021fc872154a3b376c57
z0f7f637503aa5c2217a9e7530cc466d43e1a3194fa298cf85507020e7a227cee026c81f9b7fe5c
z4a0325391d2eb9d25ba8b43be8f678f975829c48ca9d744dfec63d0301bddc028248ebbe2c787a
zbd153b59257a14476252da1079d6721737230ae82c1d648209d32c4ff2de1bccffbf0e14ddebd2
zefb8f55a1c99819effd03c931d001eef409ad2713c3742bb74e59ac8d6a58d4c228ab928b6fce9
z4c5351bc76ec084b108a0479974f7804957c587352b3c1ad99134786051bcc0c6ff6226ed0791d
z8ed6cfa211a5728969617fe58d3958bce8960297760365d55a674734c4056b583428b7bf08fe06
ze05bd89d9d5d63960d35921ad73d1ebc716c7e9ba147f7323d6b149a753449245cd9bee96f63ce
zd71748198577b361ee488783bd0647b4f401c8a53c77f8259a0b0ff1ec17f49e323ae2a13094dd
z24f547ec66acaf9793eb0b7032a2a03cde4ff406b5649f15aa1cd7c1dd759e8e773b85473c5e13
z74804e6e187772f9fe2d185fa43203c9cef7ce4b7cfcc9bbec63439f92b53ef0275eef8917426a
zda759ea98e1483deda4ca23ebea73c64c07786a4128d7e9be9f1f6ca6ba19c8923898401498615
zbcf14a118d619094e8222ce841b064ee48d67eddd6891567cecd8f6cbfa38ba4c069bedc985d72
z4ee6da8db72d30321c01766d65dbc5210eb9d3a5960212607aa62b126dbb2e25e5943a181d1013
z624b649f834fc3c2dc332a9aa616fce9ec2756e5be3bc924c4adb14e9cc51cdcd07419d4f95107
zdadb0e5cbd97c130771addbd04fa206269a80458ff6d06dc60e9cb5333f6d6f5ec7d8c9930a297
zc2bdb1cb06ac1e105d353ec696c1bd3159d9072cd85c93c8b196f68ad8d5d5c9ea3486642fa099
z815a9369f44d205b7680f594e1f932f8f9a19292a75b0ed29a2dff2e4d771c0bc6d9b02fbe8579
ze5681f6becd6a73c223b79516933b9794aa439fcb9c7b33817f82b67d868cc37a537aef28a09ef
zd4e70bf2a60c418726df88d590448d7abef5682b38b644825cc338e4cfbd5307c0bd92216d2ab8
z09ccc7751dcde954c7d958eeb0179a1c9b8dc64131cbc9eb9b8effce56804b79d35c2cb9ecec2b
z8389c8c1d8bbb9d8c269f15c780a2bbf5b0e4e06443981b3818da99cd9eb0fc709079251dc7da5
z74833b6d4792992f45e4efb74e231029bb9c7003e9f502967a67bcc69e71cdf6c48b05c9febc2c
z68b33087c5c8d3bf71ca812b4cac58c714c33233dac415dc48a6aa359f236cbccb68bf015c7f0e
z78ac81bc869c86df11feb62204b908a593ba4b5023f958bca30d8af85949f795ab6cff6bcc9fe2
z8d14f6dc4da8382596866c96101db5e5081dbd69bbbebb33ae127a5146bd8accd53f7088e81699
z26b98b81bbd7bf72d28ae22aee4078e4f769cc1676f0aff738634bbc13ee982a0da8689bdcb491
za19f0bf330c24d5cca5f4fd5830648384478e58d850b34afc94bc459f04eb3c4e2692120061494
z6ce17c8f3565f275e726fb61c46a64982f9eb4c24b734b0a90c15fc41d67ce1674efefb45ef81e
z633e77c56e7320114d88b00405d8bd82800bfba25b67bdfb5a421f7e020e0c7723834948bcfc24
zaf55ae637ca6bba34c0f4c998dba02f5a5e251b0d4f13e3ccedf1db3de28ece9d1fe422da99aaf
z9906712d3968feeb8e795d4b3bf10e291f93283722b1de8dc8d215cef85170e2a65691a6910675
zd2a833eea71e94555f1d3e9344820dadd27d48aab4bd77c51a7d3746a8dd7aee7570f54153a772
z2eb9f502e2d938c02501b6de162060b240a64a8cc8c1e53f32f4ed23d62e81d71a6304c7685edf
ze89405e12c252a88f6c1b93496cb79e33c3975d1cb503e0e4584aa3b1b8d799ec6e38df45a805f
z3fc1d3cbd2bdf803ea8041c9c06670e84dbe67c993badb50dc2af9e32ba2746657eb240adeed5e
z0cff08504e0c43c7bdb44adfeb344681d0fd34da859480a108a87e9b1eaa961b7776527c35d215
z57f5a174ee1897a686039c38e142aff53cf62b88e39c8ee3377cc4e0daeefe7a301a2489362a91
z63b1de6c3ac7dcdd46a632755fb945e42ea1ae6363b32064adf36b043666f14b98b2358228d1c1
z84775fd8132fc51ea1dffbadb9fabc04d71425116adf180e8714c62a5b658be158e8c583fafad0
z82211a07fd0096deee2bcbc6185b0d589d186890c4334ce2bfcfd10f1bd08bccf394584ab1c0ad
z8b1d7ba496142288e6bdde564314c8812bfd6840cf8f8681f04f7a61c55ed3fedf9a430a8015c2
ze9f1285109525c044ff04685e7b5df8eff4b0be5deea6f49601dc0c1aaab8c4d12a897fdf7ac77
z00382d09c7677af535d0550998c33d095cde115305fe6277e25e03113709c6434a80dc1646fed1
z4800a5b0fd944042a17a359ffceea1ebe2edcea9f8b95f3647ec458905b481f4a31f1503bc3c17
zc41f50973f79f5ba351619c6d162444d7dcb9a96529213da568a2324075bd242343963465b717e
z5457109bf1f9db19d098303a74308c69c6378e366f9fe7057e9a79c38c469bbb60b44ffda036ed
z2bce571516512ff88c332049c3674624321c5884ee87ab05005434ff2aae6231724ab877a26574
z88254f5c90484805ac3bdffbec6b1c4d9ea43689ab7f45f73616f2a5982ce9c9c74acdd4fa56aa
zd1830f5ef34b37cb672fb00f831e631117e6dfed6ad955b17c7c23d5ce934dd71b6c3c0d3df64b
z8abcc0956335fc1e8cfc8f20a8fef1af9bc9abd4fcaa604a43a27e98fad8671b111fdbd8da72c9
zc5fa0c3b22a795206a59b4447dd2e3a07dad666012f8275c3d7bcb16db7e6405fc718b54353b72
z90ab380d743f4fa486fc49dd68456f06909fc01ad6d39e8d5b3d1dc904d28696911cdbd02e03f4
zcc278859e3169f2a8ed4cf5474759c47573cd264624fd6bf0daa8dd2709e9d6ed943ae1cde7388
za803dca80c99450de369cbb53e49b540f412bca94695d54b655cd8e6e08cc4fa04227d4085f010
z1152606ea4133f3799ce874a6608a41e80874f59aa4c92de73a2b191e02006cf93e755b362d5d5
zf1f2139d6b319abe0bf2cb79e39df2849db4dcfe88c96d61557cadd03c2fcef5840c437f6e2c91
zf938db63f3feab509fd444f8c1517775d8abe6f7106585403aed56f0290b756fb7a620b6bfa8cd
z59d441839799e2c46083161e05acbd2de151e8572ae6f7864cc0857b314c05ea094ffa28dc7286
z516c58c8351793680ffefc91e3a6f20b6a84675c027a9ece288638eee89164ef06ccc7d5aa5896
z9a0e038fb8332f33703eb7dfe2584616b6e95d89708f8014e8c638acf0ce5f9ebdab7c6c4939c5
z66c4ec6a93c97998a86a544f17c0a8ce7c66be92847425e176d997b52662953e674ffff33a8971
z2e5bfbe977cbebbb7635d494f0ba4adcc140c65347186b009745af89d6037803f21b37b77f01cf
z2f98e326d96efb80e97773113db60f5b72b6dd0e30e52aebea921518b8b7e4113c1b58a12e310d
z2f032fa8b730b421e61bbb2b3d19defc7ab50c398f34ab52484a7ddc020b3f63e1921bd2479fff
zc8f801773483e54561659ad87f922adf8c32fac21c7a9f517a58d4517200a1153f32799c6ea3ca
z09d831ffb7a0d0dbdb399deccf03734e623c4a3c7c06cceb56807c135dbb7b5d45b5e11e504b86
zc1e29da40d53a0792af3497a9a8be4f61dceb2f44a75349093dda471ffd22ddd69369dafa4d64e
z781406d5040d1e5ce775a940b057ff3c0cc470bf1ca56f0baa6362fe1977288f976a5373137568
z2a9c4ab904f4e9a465e99890954298f6e3ac31e7296010e89ba02474411509384f88c5009668fe
z9f0afb1be0ebb91fe48f50f69268e9bf6874746c130edfec6fb5c5ed7c6116f3fc17ed579a4eee
zfdab3a939984542e680db037ae3312fb0b7e01d94251d5cee043697822854f21c8bbe371939b5b
z6b1e82bb08f177d6efeb7ebef65fc79d6c3f7a4d11cbd5c1760ed98554366461b7c0a3b812d797
z1b87276a9a4f2612b083115c311a0317cb122dd6595eb44cc5aa06b4e5e5e3642cf758ca4192f9
zf69494458dae30620669eceb60ea064d6776a21b475c0cacc87185692c9414dcdb768238faa3d6
z1e4a5484a549bd1c5b2debb647132263d973078d27d324ef195d349c57b29a86f61a187af825f6
z0f1aaad5e56f220264971db19e23f762195d3b4d4a7ea8a783746573900ce16233f7c4d7ba22b8
zaa9d7b8d3a61fca96264bd8cda6dc1a05bf1339a5c8be98296afb47d920040cc1b506b4d0d175d
zbdff9009b9e45881542b94378dc7b33c7a85d09efa5ae609017deef17c5742b71854f93641a8da
za43d45eec15220beda117c03fd891ee5e0f1683ed1253cab8c64858621f7e7361c147e9c24589a
z5d07c4086d493e455b8452595a499cc8c4961c5f09e3d6b6c63e6aba08d729dcc8a42f3354c25f
z8f5fb05da4cbe014498a42575de0c24d3e8cfe3650e762674f7e9c6887d0bb4f26aafd7d0867fc
z76bf218c54bd8df82c1f4a2f5e498bbb458ed957fa31804d05f09772addecbb7c5a139ee62703c
z668439e6e84d919af2d3941f636a361cdb9863bcfd9d0b24ffab5182692198795e3f319ca5b5d3
z754972673ce9baca1af911658a2ac4d2f0de9fe4c63ea73cfea55f8ecbcee7c4070cdd6a93b092
za730d4426cd94ddf17c15c91d5cdbfee3b4acb11770002e1a9736feb8b66cace34eebcec0ecd13
z400562268daa37e3eeff19eda7e615a961dd7cf207adc8025937d070f630d3a1700c558e30560c
za6620a25419e6475be59c0da636c06f0356ee90d241565d9017bc4265d68cac2a9230e6715c435
z20e9403cc9e268ad7d11d46346f3002b768b1d4ed4cfb351ef28263cd57690b76e2d9e33d9d241
z9f7b057e950991a7739760f73207813be8d3fda739e71ed385eaba4cce6c9c9a108a77499b6bbe
zd20283dc90b26278d3f9fb94d1e424602cbba7326ba0068e8a1ea5abac2347cb235a49fa956502
zf86ef8ca70405c0b73b331227ab4a1522e6ac1de6e29bf9915c935994e927a658b63a71e43f2cf
z942eb0a4db9edd651a3335e8f916e7e29f1550e701d7a4fac85869c4b1a5547a6dd5a6eff4d8d7
zb8641207108fdf2ec47e62627f5e6ff6c4156a7d01403e47fe4ed92120a2da9701ba52d50de92e
zdb27e4b28bc1aa39d5ecc95375cd8f4a271da6ceacd7b6675c44b849f4102a0d50e47b0ad40e72
z162e5235e1598936f11eca781cd35c02ad3848e3f88c0098d31ff99541538e3f3b009647c4875c
z5540d360a28d1de2ec4cd043819c29a3365c25cf3d7d4e4769284b7ccc1c691575736bd1f458b7
z2e84137bac434fbe0dfd2a8be1fc151ffd55bacdb573c4e8b5cc8b64469da8a110d9e5097becfd
z226ddedd41b1af967a8b5ee8f36663ae953ac2d9fc04c6e370bebf2ebea64a10ee9b2a2c1d7eee
z82460a129f2ec9f183b0585d038c9f2070eb95dc83422c57940373cf5fcee2bb8e40b98dd3d054
z6f16f2668f193496c0e0dab9b32445d586135a5fd1369fd36accda1594272b7760d451116f7409
z2eecdbfc232daa0dccd577486e20f4768d7c4520d22f6f09a429559aa94de1bc7c99834fd1547b
zca8535f3f587ebcc530fe2fa97c11b52879b22f0ee0745d200ca1da2e4102c2de5ce4970dc0d7d
za78dbb68e1d2ceb066bbb8575944d91ca20f0990dde703ea41aee9a8cbb08b93a78dc1eac2f2ba
zf24a75a2d94c762579c8ba89bd723a351052c8550e5d979d7ab28b3c2c0b2f6400919af9b9b20b
z45e917a671dcb6f97fff198303250fd7b9e53bd0ecda787af8cdce335767bbaac5fb74c318b3e7
z04f8b81d43752adc5548672fe0d7e6c70272c1cc98e2bfd98c5209737ad16aba693397a6d15683
z902d245fe7478f2213cee6af187c909aaf7d075f7ccdfb1e79a777c7f0a8a70246729cbd65426a
z90b30db01116f34ff2058dcfb969c0c7903149303f935884103eb2b3e5aa944a25cbcc062b78b2
z76ab4afd56bc893ce36d3bafdfd90c3cfc38e5b473297a29280b9cadcaa7f149d0f2311610431b
z889d8e493da09b442ec08ca47e6fd0ed22ccb576f9bb238dc562ec8c49a8d27c42d32760ad884d
zdea9b01d9545963e50cffbd4e73372f805489b89306dfab0a449066dfd4c55bc6827925a243998
z9b90bf2c8cedba3d5e1f2133db5e722119f72f5620b8d84e49119dae53b9f318434a30ce5fa350
z779b0e186b02a5ca579b4868730c79677e5d083e2c6e56c60d1b55c1280e4dcb45a33c9a092c5d
z5d0085c7b7966c36be67ea29e9c60dff7699c9e440a0925626f8a007725363b6689829ead1fb3f
z03573e8df15dd26032b20724fc8062953434db3e2c80cf73391a7132aa8ae8cd3a3d56b2a79468
zd72f60d2881567b15c13a736a7b106350a9580813b7f3bb4122873e28968d438ae1659d84a082f
z82846e619602b63ec7464124ed4204d596ee742307cc37ffaf4fc2c3fd33f5d085bda63ef01114
zf7abba4747fa8820aa9e7f6208853ad6df30cc2817135d5428d397d28be0b79b5264e76409a30b
z7372e9819add92d5b276d19c664d1436ec6021ca4ec8fdd2f961fb01995d4acdb523123a1cc93b
z790ac165b11b66d8c09eab2dcead0dbea319279c71376f817cd5e6ac7d2debf5aaa3b99a58a085
z960c8dc530b96c3c1cc60f4532f7280040d51729aa49236e8264278a1f99de0b81ce385ff53f15
zf647ca5ac8e2cc4370029f695fec3716a5eab41986fbcd0d6ffcbc35269c31f7024a46507f110b
zfed4519918d3f5d30fe61096a9124df34ee417c206df1a3406f28f907dc2a07ede1acec3a63a5b
za2b16d3875add713c46d251b65c6fb520f2dc1164919ff860b562cded79e630548c1562fa92c9a
z9155828c0c840ba698037ac802df09c07ac37975328b8d3e1a9279fb7764a2a222fd2335fceccb
ze19ee64e9472ceeea4c55fff6a43eb0d7143ee1e27cd0660844236a1b40ef8b8336af01812f373
z8a9696a936164cad1e9104277d7fd00a4d637b6789716d21cbd39af8954daca53c5c398e7429a4
zf2f9118655269fc8945db569284f3ac964ff597234a02d7dfa4e277e92a19038b9d439b2b0f127
zdaee23be84c6c0736ea5003e3627f892f46987da9c23f2c24a2321eceb984316a01ea800d23fe8
z0d5528727f627507b80c594770433c66d8283bd1b9f450a166a2bc82b251a0998c06ffa0b503c6
za7bdeed880b93a89ed97e1ed4b815135fbb9961c8e4ebc40b867b8585f342fe3d643cd04593f93
z82244c6ce854701cd6cf274820a7e75fefb099bed56e6774a60e408196056aff01ef83f8e60681
z730390d273c6be61ff39ac5bd31aecc84b28eca5e6f17a5b574c48c5934bfdb3de08f11b816df8
z6a1dcbb5b391a525c43c536dba35400d73efb0075228a9d9f92c35eeda352d338d8b6424035e15
z05447ae18bf56b6e71b2b38ae523354f5fe2eb723965e05f03315ee773ee7bc4715e739971d067
z3d126408066abfff4eb0ebd8c7bba94481c8cdb1b82d17b89c2aff22f5a24b8174119f6adfe02d
z797970076025301b27b20eee597cb2a59a578e5acef3fed1b024e30020d861e5fb2a1bb4dc7717
z9b2239cb3cd6c1c1cfee9ede59d3f64b84db1b32737173e8d8dbce35d87ff744f74b1a8e83dd20
z63f84ae3d4403531a2a6c403f08bc1c9181b1d6e20f7764b9892e25fd490b00ba10b7a8e0a4cb0
zf7b6868b159113bc69ce9d4dddd55c8a3359f91ca93d788769f9fbebc9f0b7f3f176bf4d55b13a
z34980e112b9da4ebe4d060f956ee1e0a93f4cf360fd81ae35e9cae7d7fc926b44bb42ea1602b65
zae52ad3c8b78858859576bfe491b572beb9d9d7b98095a19d2dc9330142df0add40b2ac8df3532
zd5e177e2b23d8248b93784068ce3ac4b8865ea4d37ab702ab244d43e9a0dd370b9543f2c442801
z3e0751b9ca38c80b70abd56435815d2400cf38d7d23204105410910450b97ad9e958bd80105090
z43873de6fe45646a4c5a00dfcb2a6e6b5d7191853d986d677e1d01d9d7006054b276bddcaa13db
zed78989ee889a913c19d1b4a192fdb58ea9b7f0eabdf6991cc53bdc61eba89c8ae6ba8a2be1223
za562108009990136f8b7966d351912590c9c397a2d99a628a2809b7b3f678402f894b2d205ff73
z0cbfdc9c5cf8105127b917f11ec3443b58b965c0a8eb66372daf6347a7903e1d233c598672fa08
z5c6c4e81ff11504a546a41a2dfb41e5524dc251af0417ed8708f3e31281babcc5b7848696b09a4
zcb7c2811a8304475c5eefd0f5b96c73208112bf0da2cb790e59c67fa6027d5ff6441649c623ac4
z8c030bc598d7398a3328c8541efa3974011f1723d45a0c3e75947d97fa06ea88cd75e2f223f469
z75d63b719cc1d32d7e9601cb7a58c37d54459834f5ace39103dd54b96a72865b71144aeb273cfc
z2a0d1cbd2ad310477b88a5e310efc525879eea99e7a3ec74c45b8ec573204325e5a91f41d02197
z684507e6206321f1ef59562b074dba0063852d0957fbb93415bb77367c95c17daa969e314aa56f
ze45bf58fa3492ebc70f8dae308e7c8e7ea5915db272e3e509d73c266fc2763d9d7ad91b015d1c6
z4b912564530efe3a7f1cf1b847ffd5d5dfc619c124103fe015d468532922db7179ff432b50443a
z4ba7616dd6e498c81501eff8ba2b0ea10aeae6df98fc3e05924f07e8ae2bf06bcfde746d139cd0
z8aae86e0812cbc912d706a1ea6f944a90b6fffac25c425c1f3b8bd96298d3c4d73c866e7388ace
za6650fec7a17a31b59dbe53e4f4203ead132ca93c70a0f33fb9a8f03332da1b81f8683dae8e20b
z0d6b67c725005cff3f409697409e37d4cecad46ad2ab33041725dff90300aca6053d93b63a02b7
z6cd0f501211eb58aa7f452db56f45d9e89b876a96484ff56a33b9d8639256ff0eb6a472a84bffe
zfd41812604d88ea1e7a5371e16276f9e4dbd0aee224aa53f824d73d2f78f06f6e07957ea1f3ec9
z61106cb2f6f88846b51e047ec2bf1720a1a28e23c7f41a9019843cbbffd84ac721499355f0fba4
z39852ebff4360509ff6748349f2e45f6fc0ccea4b45f2aedb6c03ba4848d95753af99b3caf3b2a
z6270b8ff17af2cf1f9477a57b0b957133c2da2ca67c21ca2085bcab56979205a8f0d1d546e2f32
z2138f831d9725d98e87aa1b02f168fb2938f1909c3f2a32f10169d4b55f9d3b004058e99518f98
z649bfaec5a7117f7594bfd987a70d8bc5597341fe50816049d933b0e08db37d3feb37dee6dd82c
z7cd6e79ca5e97c1bdcd06513965d964c65794c162ba6b37e91b98715beaf278f402efdcd8812cd
z27ba3e0c0f8e90d80ab2f634a25f79e2e3610078d758f47f38907ce0cd631fe0e1f7095e7de8ff
z6a7dc28270bea41974c8186fedfda7c5a1233d7ca0673611a0108f745d337647625cf5756ff0a4
z84b3486f9fddf4130f2e598b547c7b97bcd654c6911f34a61ecf022c75121ff11c2f640ef1823e
z06421b15208b6102f07da1075892cb41afa819a5f06f294ad435fa0f71128823447fb6522bdec7
z7dd81aa7028b9863ab29fa5e3904a14fdb4550afaf969cb3e34d6ff38c4eb2db8d5d34dbbc08ee
z0c236229a50897249489e8b220bcf2160b66ca6ba6e0c5b60febadbfdd6ee66a61ed4e84e1aea2
zb53825083aaa5e27ac87d2c2664520f7fecffc4c147df8e547b30df23de3028573ef17078d2ab2
zc4b046baa6df112f1a4e1e4e87c7ef4fa11375bd1126627cc7b446cf1bd1aa695ac433cf61b5f5
z1681a93c32f525410662bae89e80056beb243735d4e35431ce88c83f75c88d0969553afe5c5531
ze6ed0f58909193ed6c43883898a521acfac97051bdae8e92406d9381c4bb12a2fe17e71cc6a059
zd6517cd3482353827a858b0410a77e3dd8c63a040507b35f5019c4f8333c0a6351c8890028cafd
z994028d6eeffbce0adfb3f74fbed69163e915afb3c2590bce9132f6eb0dc68d9d8a630769a48a0
zc50e5bf47e34adcbe7410ca1e3245ab9f3c5bd6b0072de3770b7495dc8e968bbcd407f45606ee8
z983c9cf94268d7097fd67fe1c8162d1def403b7bc6af9919744523cf86f65fa270652b8d38c261
ze5b0bf64a4db1ee02e59fc8f04f35d8a020e8d4366a14a3c96b3bba7d28aafabc4bf95656e16b0
z3e1cab78888074b1147fcd49244f0d045c3e312f8f4a995e2113668b69eefcf6d929d6d9d42efd
z945ba1eb0e104e915da2117ee5042d0a46a96f97dbff2d95ddfc1a6090cc384931ff18cab6d70e
z97b9593752e20ad6bf1ed86b1455bd6f7d22a6347e8a0d2f8eba0b847d5ed9c13651346511c946
ze0a4c7b5715d3c57af512822364b202b1fa5018dc5d5aa40261c2d63a6cc4313c4f0b802d08764
zb416c5b47f2db675052eb888831b0e4ac4e4142679857b187e7ea03871971ff858e60d5062e973
z447a1d947ac695e2c7f5acac93d591c64275f458c903c024a975b3cc40838c5320f3eb863bd7ef
zc5f3f5261897d1e5a2b9ff27897140408b28e72d6c3343b88ea43627c60dd7020651e90121bed3
z2b4b5fd78fa460ea713cb57da68bda0a13e7746bd66777e5a0d783c13d41863821b041c4e123e1
z5553904e7cce73619208a544d05719b8d5532a8bbea04154d598d6ef763c49acb73f4401fe31ca
z3672ebbce5f96eb5250c387dadafe4bbf11ea78a5ea3a339ab047c0cff2a852e357e92b56d2d42
zcb2d058a5faa5b948e4a52bba87bb208ca7897c1761f681e29b07102797e38759fa0b62c962aa7
z469afddfb279b95a20b70f92c33872ba803aa921dc98002e44c42f5a8811bff22eb4bb3d929015
zbcbf383525de55ac1266edb8860c47947974a0a9cb86432d133f42c0bffed2a339a9d0b4160d2f
z5c666bb211a69c98fbae7dd31384feef8707a4eb9c8a4dbcb9842da2b9eb77cf09a07311917d63
z553683ee4392cc4c529c43097b0edcb7c56441f9b4ce12912a13028c898095787811de3c65aac2
z32f86feb8e783e4fd9a5cc6cc426e880ddd5d655ddf2d95fd53344b0f82d6afda3a5a4e0242d4a
zdf840875d5a5b887a0c250e11a85fe6189946c3b4f89d8a60529faaf4496422b2c9d87558a5033
z639db8798653114d4cf2a6f09470274ffd5dfe8ad2a656fa263c9d3b65d7c0e48777ad56407dc1
zca92a2bf41e30247af9ec407c674849685d7e572d464d45ca4276153c0785b57feae49ddd1b5de
z6e09d6c6fca2a7c29917b7e55a367ecf2de90329819f2e352524dbb242735854cabc2b364a959e
zfacd9da6efaf0883ea8c416cc38c8b299ec0eec446ba14cf2ab7f5fdbc77e2f4ec24c73540c805
z821bb746f382ce3cbf0da8a4b1421bf97f5f2032a2d3ffc75a21b53ad396652d60dda11819f95d
z4d39eed55bff4e6007c1639c7cd9ea385ba5e3b0a27a815e754fd4a612c5602ced40e7a913e77a
z4644d8cf5864b48cd5e657c57864aa4a35c84c9eeacf31f6f9091e8155e86ff735d77848d850b5
z01e20340d4d174173bcd62e977ebd31a3c75ec4c376669d44f6aae1a30c2e14c5c4387687a7367
z26428e4982515b27deb90acdc99bbb6029b7ae375175bdff0a24dedf93135178e1fc09f051c653
z85be8aed463b8e943957199422cd03cde3e79de870e1d47c4459504c5ec42c366973f826bbe998
z88650c1635080b3cd41aa2ef0970e36a6a92802a82ee96ae12cd1a8c92595975ab028e7b54c124
z2bd1cf74d12191a826b2c54405b902dc66b2d612fa487c48f38c98735d4c1774f23b898a6ea291
z181841536e3df62a1199bf5a42a7c9b67de33580f78c8f9db961efc626ddd935edd74ac5654458
z5d75a1e8acd9ba9cad663ad03abbe348b68bd50b5a9c27ac4389e70ef3de288fd180d4c207c7ef
zdc564f6480968d50877605615dfc41be506dc0401bcb32b008ecc15daeefbfc027aec3dcf617a7
z43de01d39096127cbd87ca97eb3d032297a4017721bfbb26768f20c4c961059e2062d5a65fb019
zd693a04882442cb7b09d5783fee8feed2ac534914882a642cb591e5fb754d98cea67b4ef2086f0
za7cb1eb8d159e4eb7179da36f73380b54c205fe2d586c234756eb30eda8bde4b6954010b7ff115
zdca9f148a28e04a16baedff11ac89b8c0e7ef42919ef25357ab4ad79cd7b1871eabf65a4229398
zc12026ea742f197699f5c13ea0b4f6e447c033a5697abc09a5961ccaa4a5424901977cc99177ed
z6a884c4968f6451fe62f75a533871e86d5400685ff741f4f6a6a0f0ec76385f955cc43e9334a5f
z26e3ea001b180bde69adecbd7ee88827d5f3f3b436beb3c25592923d214a9ebc458eb1b2871344
z73f0783dbd1fa2cfb26f92589b69beb3646230376f3670f4302cfab4fbb68f56677112a95e0890
z14187b54261a39182e5f03e1d3cc1c1c4c3900dbe8f28fc3cf0d14d66f89d4c8e7a32e06e5821c
zba83a8463924576d7611100f3fe655b71dc91431b5e66cb4791424f2af00f0cb8d2da5053b68a8
z4807d6e386098a07c4b92ee9dc800114c0f01c4cd3dd471f20ce3f624d49370366f651d7df8cb3
zbc04d8926d085b5a842db61a7b393c0e0782584af827d7074cc7332096cdc6200f5202edd15366
z8d20ec51166dca8319953bd1258e317ad33c9b701e61746bb264abf32c8ccda1e09b2966fa4525
zd82f3d719d28cb11d3bad02e979734685877d22fa8b5498af2afcbd9cc4805ef4ee030c9f86d0c
zca13475af15c2ac0180eb72129556bb125ada972ebff1d41ae786684a34edb714b4ef7fb4fde6e
z41ec2ea08290593a7c8fe3b71e590d061b2a5a5b279398e610f5adf5c8ddc3d5dbb59ee115eb6d
zda12527a8aa883abb791ac8dff5d937ef9715c42568204504d91c6348e12379e1663b171657c52
z62cd6f4bc73391c8e98ec9a351fd44b7fb04bff83a778f4ef8a237c0e63231bc0f1fcca56424ea
zee6e741482b29e63dce70ce2f845cadcfaace04225febb315f64b3e2e9431d1481ceed46104b0b
z66dc491f272b47f4b90639451b2e5cfdd8568f50aa41f1792b4c5f8718f8904c9869607dd2851b
zf8d929224fcb412ba4b11b168af0ddceb3f884472c98529e454999799b3c41685b68f53a2597b2
ze87e393d036356ac7cbd2bca97fdb28c79ffcd5222ed239766eaee3b4cdf6e44c3e7dcff8b417d
z5a9960764d0211f97771820611d536fcf33bd853cc4cf7818861b0b03f823e2fb592cdd63a6d51
zba741b69baf675e385f1a985f0fd5eee93dad4ead3cd88600a15614555e407463cf58b65e4b8dd
zabfcadd2b8146f260176579ae3d0082a4c406885332486fc81611b8e7253c470b719ee61f5156f
zf805d762f086f9cba9aa26d6df7172fe7ffa9c7c48ad3db3ea5bec9a4d2cf2887cdf9f71cfed15
zc01ceb24f70a96db63259d54ecb856db99a2a0a4e4f46ee0adcc708b2a8f29b61bc8d0e8bf5c17
ze22987c82e38efa6f7f3984da790fd499e20ba08951122700331d2da8f8de04d3d264256947bb4
z9f5433d8479070e29deaaad9e41c1f903539898488045749590c4fe113adc39be03d6c1a6a3064
z6247c7ffc2df48bf820d9a7eda9797925438ed225efa339c7190bc07abf7737f833aab3d650005
zf1c7c3d166baf653ed6ce2b3f24a05db9ed1e07a3b5259dba565f56d207cc9a7b2f6c872012903
z59ba45033f1fb821425f9f1fe4ac96552ff9b71a176d8b4ec6d01b610084c12829e12a098cf542
za3d77af0cfd04c324cecd39333ed3007bc864d2934a6c8156c24fb6f26fba69eafd4361143046f
z40828e2979554b1ffa1211b903f206e50e5b7fe8defb8b3f0bd66143cff72d199073c2dc166381
z684065fb93086c2f3f7f4377ff0944add13b81419a094a05c934cc5c368be92512d52e1d3caf77
z70d730cdb8fe557b053ec3e63ff26536e155fac180688291fcba1532045dd2a270a4075bae6a2d
ze2c8d7f234aaf228e613b21e3bc4e976b99df15f0d44368d90043158e52fb97df1db51efff5fe6
zab495bb1aa84e6d7fe2fe49faeec06b28e012c64fe44bf163dcde37c43ea933cbd521a280ec9d9
zd3ae4311cf6856b13a1830cc8f5405fd1dcb8797d435fbaa9f9f0e37c49ce9cffdf05c51192e7f
zca45bb875089da030ce3cb209b71ae990671e47164151cbf631184d7d14228d619828dd9e1e688
z0b9648a0ba03e33eb32cf790db057302040424f57ca21c57fae81fb76cbaf1c8161f2366e7b184
zfbd9312bb75e69ab7058def5a6be052c16671ae777b11814a0bfbaeea6fa12a20435f3b6c313ad
zb757e87acbe3d43e3de04280e6509d3135e1bf724989acdc6790232966eafa93a22429000eb5df
zab1d76c406a44c4cb43d48b580521b66d176d1f81873106bec64a6a8c4ef344548a7c37b7f21df
z9133fe4cfab094b5e3c5d77aae3e6a76a0fb85c8fb312ff8d7ab413f5e94ad0fa7aa74b81a6b2c
z2beee7fc87ced00bcda05593ba8b6374fc433288f3a78a992359049cc2dc187f34a6f92bd3d438
z354f01f7ecf400ed6fb3efceb10e66a9efc0f6e4c2caca50c6471eb95efcfe58eea06abc876818
z90ec904f26427a792a35284ecdf24266ebc54e7c714ecfd672499cfc69b0a77e3d01b27ed4f486
z73a3acbab33e2b4ec2d9ec30bd0ebcfcba60832a6cc8efffb293dc45ac48de19c2b1a6cf035582
z56513e0c2d4c7243a945bb0d069b622674e513f0e8e74686a3f40af3a32913c186db455e203ade
z9ab3a1d6e83198b91d9059f3fb1b363dae94070739d75374444c87468060e0193c7121a474dd5e
z4cd446e5d02e560f953a93d8513e5db0733a4ab1b2e9da570b6fef95a252df4fac7bfa07e8ca4b
z8016a55f1286dda170529391b08fed3148c7c5414b1ed2b691fb2ad41b2f358f6abb760ed94d90
zf390f4f23df48265952b3418c8be06a2a88c5364e793bd6a531c0fadfb03e18a0283e62f7b9149
zaa31fdd5b8061520ea1feeba006949532fcb2a2f44ba04ada9bbd08e5044de5ed162546b21eab7
zc9a2cdd050e81a0193b4d3d588272240e08a0239fce449ea4407bc9a7e76fa93dc43ae193bfe84
zb9527e4be8f2f07cba308c23ff84c82ad5710b7ff82b6834b6ed8ae3d040d62efba5f212a7a537
z51fa94cee16019ba34058035a1f7b79e8fabc4c6f00cf4a91af4ef5bb0b6fd64a6472c8e08db5f
z1465ab8d32ab7410a397267b3c53fe8b26752547530d93dc407a5e265cd1f461c300663ff9dc90
z6a94f0c2cf3418c069822110f5115106bdcab010f7edc2c1e634c01bf2f46685f9e00e72ba1c28
z50ce71b280da8b55a8d6c44c9325b634eb2cc1dd2470b6438abe300ed82fc6ad0f8ce3de331351
z99595ff888d267c5fc5d82ca912154755cd44734ddcc50c87d9d3184dee60b1e35a7c58a39020f
zde3b27a2e03c787ddc3f94972bb1620d93932b738a8c13bad9a0b70968e9e0c106fc97ddb1646e
z9859f164a9b089852cc096ec2f2a5b194f3bdd8ad9f0fb69289a9fbac438945f4a6d4ae93d333f
zf5c9442b958a897de2956c7733629f51d0f97bd056238012b613df06a09504afd2dfc076dd6c24
za42c9db7d4a37b2d780cc3f7f94b94a99579e7ed7661a44c55c034b96f2a00cd615f9f940b2cb3
z766b9756f266c5e40e8a390d9d5ce5ae0c594d8fb250e71c8f28daa9ccf46a070ba026349662ec
zf815cbf6559aee43febfa117c47ee45f8bdfb797b79986a3d752b5a2e45659f18b36adb061a1d7
z4f36204eafdb43e0ebfb6d0ba10a4de24479a33b23c4450fbd8bf30020bb5ac092ca4a537daf9f
z7f78c2a88596953e743057044e2412634ea5fd824b3e1de4f94af9e267da979695fa8fda71be01
zb94a9cf9e4e48f03ac6e4d8d5999c5c54770893342260d9e30f8fdd16f048e0978f60fd5a3b942
z8e10e0aa86982de0032e482a11e85d2900de3f4ed74af2344204e3c0655d5c270fdcd248c77513
zf6544656880f8e2b654c7f0edceb97b072a9af8cb940d5ff41fbced49d152967af8857f12745b1
z3ca5107d92dd5a6c2d97210b25735fc849ec4315cf5e726adcb9229c5bb3dc2f7f0aab61f2f2be
ze4f077c3b2e4c8594939e5829ddc96fdbaacee4bee6e1048bd7dde22ce08922bc8d6384e917bb6
z0aa1c410e87864655813c016a6a2b217d10107019aede03a8b3e9f6f95b32f83b6fa2d66c91b66
z1bf3ea34b8e4391ed14e39cc0e0b98bfa1dddf0c2542ae809599ced1cc584f20d22372526e774b
z59c210d5b0c5a842c5a000f7ad48c2653278677b87d4744231320154850f1cd650bfadc0f1d640
z2224d0bcb4e2e4d5a59488664b64f73fa29448acb1cc440662a9bb995381b918a51f2cfcda3188
z4d0a51b9073a4146d6b59c15ce7a1e1ffed19d10d874975d8f4409728219e2cfc2cc4d66d796e3
z2c779c459ff58091a2687e7c0c97f1550c667ed860f3a0acdd0f768ef07b4cbbb3d7e180503b18
zb0e391b5ac7f108b21f020294dc3f19b88ce6a31ce52813cb7b348686da0c43b9cb4fd7ae61749
z1e7e96809840135c06b3c54c24502f2cf05a2d834e42766705bae87199b9bd013687efe0108264
z44fec4a0a5d6de7d92f0ec2457013f418029985b13844132b0c4da50a8a8d11f3ce9372ca86a27
zeda21119c3d05b2d06a57fb85f32b903cdea3d2164c1b2a7c01e1503bf4163adca922ad8cb609f
z31a8b43bd97021764bd5604abcdbdbfc7af38b8f514f5034158b7f12754a872c12a4bf3fba3a1f
zc9c34acd6486dc02f9209de83e5a006638e5fbedb1378f85a006e4f3fc51346dc4e849303c01ad
zbd94da7cffcadd42446eb5df4ee4b7ac2db2553ff1036c2e0d0f5dac739f5d3bb64bad9a7dc4c5
zdb7678676e31a78b9fe31480ead66f70e7224dbc849db9092d4b9d04527df3d218224970591e90
z2427caf629d763b637a1494cd0c3e0b1f1805130f2cbd28b36ee7ab8c1101862fca9896814d3cf
z909d6a2b458059bdf747e7a4296d0318f484c9637a5c7494c1f2b7ce52bdaceab7ba96d2b22aaa
z8e25e52f83b1e224f271ab585e2b928905f506b1e6cdf4c2b3a0a88186b769eb31643833a634bf
z567628bd4289525e009037a74d46e3f55a4890c0a996f350c68056e8e9db9acc232e20eefdcf34
ze6a963a1ad78c168829938d22e92d8b4e88eee27574e44368df76d82c877bc7946fcad51735491
z13a941634af8ce916c25732577ac1cf57e29217934e30d3663410f4971239b1e64360f34824fb7
z09ac1a14df25c041ec42df7b67ef44fa01a704b4742091d8bd29cec8f52c2a082bba321580e6ae
z6a6620a8c9ed2d1248916c8c186449c833f2667b18b44984e3e8f834425aed32cad0518103ec1b
z062f6d53aea500214399f095e4862d98deca06cc5a217f8b251de6d049aadc83a13535e0537c20
z55c49fdaf728d17445b5fc00b94c891191920e0f97c26f72b972d18b21c97688a2051fde47ba74
zb61880473aed169c3f5751426bb9fc58ac44307770299de34f7d4a7bfea12624fa88e0f97522a4
zd07bb01836e56f8fee1438fec94fd80b6883474a0afb2e2a5b99dac7af85744961267ddef4b483
z62178d1d2df3b6ae83d1f28f2536b6ad2d1d2c2b4237649b7b124623874191cd591f830956ed23
z6c75311c7580ca30b38d95091579136ae5365622e8a5e337603f15754a543a8f48be87677ec059
z0654fbfdc3a866c9d01dadb69b17eeaf76330f3dcacf4ac7cbbafe3bd0fc4afeea823606cd2577
zbcaeecd35bb549b30d5f13f1ebbc485247554a3ac1bdee1f9dc613fb916feb27e00986d7926d67
z1acbc2e2e5eec316ea696ec182fc948ff2abe975b5682d084bd3edf767a7fca815fe5e8544d5f3
ze0ed8538f0d7cdab6c745dd7161217948d212aceed11d7716305c5b88ef32bf0fd300829b5b6b3
z96fd1a9d6e4e903e13dbf7c0eae30330d50329c99998cc8adc103637d0b65496866dd7088ac4fd
zd00fe77a12578893e2aae8b949f4ff5efe7194f8125ce37d083f51f31d2884a117a7cbe4a5e843
zb519ee465a2432fa2f6016a153450bf2ea0712422cde41eb52ffffaffe62170f8fc41ae985fb75
z3dfd6176e75811eb97d3676dd206eef0f8ab71a36ad924fc3a2089943235954226d0e9e8e3f61e
z5f1885a0822d711876b153dc2d05f071585238a8edf7ff9957e8423289f51a22304938ce9634bc
z0cc765e1e18e61214f4d8e122c58d0c8203556dbf626eb5a7b7f256bafecb637d81709705bdfca
z54e784a9cc5cb20077633555846348722ae38acdc020a1cb90ede4bb2a99e6c107c1b1f1a44103
zddea5831585eddde29eb2c2145246d0e3b1d2d26ae136955fd6cc0b6e6c5db502a11ad52284afc
z78506a48a9b58f5135c1ec1adbfaaa6c581cc3643cb1b44f61824eda68b2f6d798018c93107c8e
z71d6ea827c681b1552fa6519b1b07c1661e67ea0031e3c51efc08079a5d3228d96b710975a7f6c
z3f4c98a145020ad34418a77fad09e7865452c5ff6d8789840bb287d32489ac423b45062d622d23
zae13823efb773b14d6eb459d3764b37a623a3a17019ec6f6821c1135c6ad4ea07cc1b18a3bf688
ze2abc476c71a69ef78b7099cb49b4eb7ae9fc83c1e17dcb27b8a7412b77b076846d81c8c61a0b8
z5dd4a8c927ee8d1abad3bce095a530dc12322226de61aebaf9c74c4113831189c6f341b44958ef
z3b20f7950913b7e09a024f26e9732548677327f1845e125e7f3258ba578765f337e710cb8abb80
z4e051fcbcde03a0bceb865f22e40e49d00e2aff878a440d3762a6519a68f94e50b5aa8aeb6046d
z12b46f06b4dcb9260896737b06955cbe5f02c8443ce4f7bfef48e0f7ddb8319ed701e734ba3240
z8188373f62356ffc81b2a3559326ef5c72387aebe4bb94d511c7ca967d60b5df81547a3908da93
zeae52b31b26e478373e72fb88794fb7b6f49bff28f986f72ffbe62e8b74eba99268b1eb85b4e20
z070f255ad10380bfe258fb5a113e23fd151acb8f31bf7ea376eb5d524fae5acba722470d4c34c9
z4b995501081b69a445109f5e52d64910b655d82d566ab835358d2f9981b65bb258c07a30b56028
z5b0756430e35ca87131a2075b23e6960225fa63797234de46b3c69f71af6fd16eb203e726b3f7b
za2eaf8c59536023477afa6d50baec1ffd75c6fa56ddef300e00d65123f328fccefa63066ce16fc
zaa53f7a7bc2919c6ce8400bd78b16950449e55a08698e6b8cf11045da6f5be1e61c10ad7dba16a
z7026901508fea3931cca77740d26f4ca65febf10c2f2ff53b8b0c2aa59d86eb6d42609d8c2be91
z74f2fdd983cf1442ee34cc53b881b1755c1befa619709dbafdda8b45dccf2998e28c6a50dd906f
z103c6743f789ba5c8fdbdff08e405d2ecde5bea893438c6fd15075b3e405996b28c09959e7cbd7
zaf8f65c3c7ed1834f51914edb562f1a38e6c039a5275b3722806dcc274ee7e94d9580ce6b7b743
zb11caf7e63086c7a39b3975f74a9fc7d0bc6d7861c012ad1275054990f3065c6943b4b25218507
zc2bf1a404ef56eb4c8a9566af1567326bb6432adf6f1cc3a286217daf5d7d9c8296879a9cf8bb1
z209d979978d17df0e066ac7ba60c0d76de9ea7e9eda1a7cd1a963a9ef1f3c4185b9022e8aaf2a5
z3fbdafe2dd7461205d46389cce34d9c3ab0b4bf7c0a370295ab335465790de1bc1cbce018dabc0
z87fc71f603c310d203a2ae8630a0f54452302e6ccb80084c2d6af15c69dc8ce7a1e6f4210fa6e2
z6e8dd976fe4a6d7a51329f86fc8364314b8c94555739335e9fdc58644a002358ecaef90f9c8030
za6d9215e1d07211ec0f5e9f403d4567da53cd11e0b05fae40fa1174bb2374bb903723fea70ae95
z4d8bf7ee05af2bf409537c216a32eee8a6c92c321699d2e91fc6915452e4ef64e774af65ade309
zb8d5d01307c880ae0f5880c4d1f69d54830ea47ec2cc56f694b7ba930df0dda8bbeec07f9ea675
zeece8e5d42566469ee1b019d2741d0285442c5d9e27d4d736ad40f844fa1fa793cb1787dee2e2f
z184d76d253088acd0be76a9da0040fb26662c7103c14f74bb280a4f61ba1e813ae8ffd7d02fb23
z0ea01da8683f49058fe5f968497255e61bb265686bc35fc7122c6167946441b249a1ab4c420ac1
z7ee2aaa4164f2f1ab38d530bce214da80d6956ace45c8ce855c1556e89367329c272c9bec19169
z42a5686d0fb4a5f58160e1d33f4cf520a2060d729585465f76d31a4e7ff2caf567f5e6e66ae1be
z7e70261814717a15251c467af5b88391fc8ce23129cf6addc2174ad83cb773859c8e0b15167b42
z16d4a5422c580be22412e58f4041d497aa1062b7141165c92779cc240afb2f7ba891bd4bff8aa6
zbec5d47b4244102ca5a8eb170460941bb89db2a354f749a1ac18292bf5e1fe53708d09072f824f
z453ab28d2857d271f2b689378f581684f58df0951cecf866682d27a4f82f618d7dd068e97c1182
z0f0b28827e3f24fbc59fede0148b8413600f9108bb6fe7ebcd2fe0bd4ce2c31bc85e457552f96d
z333d3bcd7deaaf5c6e85be96c0a430ee36c9f2a4912e622ac81bc8a92a5af63fa308eaee7d9c85
zcab0bd29feb33902063e1858918cba3ab8742b2715cb2bbaea6c408a9b2c1a84f97e67dd78d873
z0aa8b6dbd061071f075c879b0ffd283b712a4184b8514a02fc8a93b5c0eea835d6e87378f2f902
zf8c7c3780cec039d619301914fdfe2c952b66dfdf27f26ed9bb84229c42115ec207125d631fc15
z5a12d7f2d4603071e252fab028de455e633c269f6b083ccbc71aef69edf0d6652a77114bff7f6a
ze19a96b47bb61eb7e6aa64551cbaaa006af7615ac552670bcf13279e9459f058d1de5be508eec7
zcc8589666196b2fc7aea815dcf07c08b9a05b6e7f56540d813cb635a288eb9810c59cecbe7c872
zc62cddb18990a8917442bd22f61caa17c5480586c173881dab8020104d4cbebd6c91e9fd388048
zea005b9149b6eab60d16dc5f4cb94cd17a4db8ab94203f41fc74348273339a6d4cdadff3346bb2
z44b6aea734468e8661389957bb64da8521bcb8c0f2291a13d96babab1549700c86b235472ddd3e
zcaecd7dfc7c58d8b12a0802189eed0eea1652deedd8f2f8a476ffe6a700ccc605ba10b62b585c9
z82f569345d938413d444d4577f33916972d4b8964912352b1d978d0ad6fb32c71b2f0f6ebe6904
z3ed3d10092d6fcdb8ef01e3a371d893bdfbda13523f1b62bfa339868ca6bbda1f38d0cca987aeb
zae44abcac196656bbf511048f12aa4eccfd00a6ff08a7cb69bb4744f038adced036b9ecabda132
za38499bf1ab2a1230f701a6536bf97472bf6c5f8d107f328fd64350698bc8a0e703af47f1b977a
z73c365924c4d747783d0e89c07c8575cfe588b4f37f0fdbd87bb4a54b87e2da4a0f6b32fc8818e
zf4d95824059c07f460d0c9dfcbc201f1b1168c06c9c81eaaca20e2ef3794cfde175201fdfe1bed
zd8501e41a759e73c91b3c61e4f2feaad5911394c1b7740f6f95c09bb2d979f21e82c5928c96243
z94dc22046665a51cae0d18b57b7913c2d6748796505a04c284a5de7b82a8ea0c6bd001366a05b8
z42e325f88efc2e782b3ce8e83ff12aa2a131cb6552489b4954b0c71860c0de9f10cdaaf90f0544
z5b7d1697f314489b3ec41165dd1ea55fa79da5c4cad339c9a07c4d3d6bdf54813deff7d15847da
z008a7cc435c55b7e813790ed154129663b349e0ca38f2d02c49f1270fa952ac4fef51ae92071cb
z40dbad152501b7ce43973e71be80d21eafdcc710e4f2c6a3bf0aadd15249c7ddf1710fc5c6aa2c
z38ad716491f89c50abdac65bd0ae68a64b57c4b79e0b68975db9c7278b6744e4ac129b16fd18c1
z7c909bb5b27df8a4d6fc172fd3c1c106be487f4f97c3e2fa7558290c7f4b6b583005604c095fab
zdbfdc612dbc3738b42f857997b881ad4d50ab4b643b23fa11e6810e37e89be5294957d9fb5bfa0
z2d48eb12b29a3ab25c759a5affc69ad19d1994aabd44bce5ac808e466b20213e3045c84110d7e0
z077a56c833f6706d569ee57f63bf80d2493bbc5c27acdd462b48c3bf736d2310feaddbc95ece92
z6d8f03b3b47dae6d899f4b54099028e9f6f22291d5fa91a7e7eadc40a06c3aa0cfa491c8dc8438
zd71a38839bbe04a450c482ea26c6f21cd92d133e49cb88a0c7d5868f46941053b4bc7839092fa1
zb62a72878bc169c946a491a550392f70eba47c49120c54248c5ba768061067c36151845d2c70b9
z0a102e4f3e4ae6f45885d6d5eb0068620f8622fb024b4c1aaff33fcbb92f2ced0cb7159dc1805d
z81f9d789ec43cf967870241d25f3c62db6eac0059c6d692deba9ac138df5c35e19370a3862c965
zbc682030fceea9b7866ea89bfcc33a364909c7b187bda873dcaf28cea4d9b7ba30c64cdcc7964e
z187eda5f9b5d5fd8281934a309c4168d61d2ddbad955efa6970bb50471c31479d3cf6eaf48d8c8
z268599767d42eabef019ee106c68d1b5d3cf425059d2c6565d9f3d5335ac148b8fb88b2a00fae5
zcc2a1a3f8bdbea3bd4d9c3df346f6cb16a36868a97189d3c9404165f20333ec8c7e06d5f80366b
zc4a6b2c2362022fc2233d7b9dcbcfa4c23d9232768e3b962d8e09086c69942c9faed5abf8cba81
z4a54ed8ee94b2fc6fa31e040ec4906651f9ee6208bb814c3f32461ce4d5b0579a91b43d116015c
z72e1c4e773cb33a7a4481245e01726f395b06b2888619d411059b3d89a619a6876c2c0cdb8594f
ze95efb1ddc2fa1c0266955e0c248ddf79b02165703209deb9aef4ce7b5603dea0f07f45fdaadf9
z6403e2dcf92fb4054fa0a3a4192ae6c1fb31f6e48c691232fe115e69aacbb35587f3675e44f1c1
z70a5a2903443fef77ed6703a592de0cd305490aabdad45ab32d47c0af8140cf1c382c562ccb511
z835502b9aa9ad61a2f51ed194764a520d958b0ed61e79e02de89429064d062e5f51e94738f6666
z5b63443fb8505ca5d2a17a71a1fd26d40cd23a6d1ca4653b56a2cf76d080c8c2a9053bc352c38b
z7475e3aa435b59b208a754cd56b5b09342d516fb7f50b5ae718b6779113f89c02a25b27eb94f49
z6e10476fa152e3e799f1a00425f5b455cb50d59a4b0c16c8cdf01d97268e413736148eee15e75f
zca29c1e61fb5180b2adddea46a5d2c57c83fa3960eb3f0a3896bd86cdc408cf2c02cc857e83abd
ze983bdbdda613ba82f7a91ccadc4dc9aafd464dd1125cd457db148c8cd71a8c18651947b991242
z4bdc5a418f69a8e9ff983768dd8ad97daf06ae17548fbf6ed0510de6fd44c18198976673b98d78
zbe71cd1ff5423128531977a3821117e746985ab68eb80a01b916e2280734249ffcbaf063dcc4fe
z1a4ca3a472736852589b18165226642eaa5b5468eabc6d1a5d5570a12c8c608f50781fa61e0045
zd7ac7512608ee708d19f095ae9e68b8165a5893fb1c5a95beb9ed584761d8712c9f7ce840b821e
zdc2828c637577817f6ea693b679fce0c827f90d4f23f6be5cabb9a3659ac54e9b9f571b38c2571
z1a6daaf6f2b25236980c8b4de58c5e5ac37c6ba42ad0276fa6f21a7a5de04f336a5cbcc63a6c78
z6fa742f003ab2e248a4c62aad16a03eaf934f12cefe107ef481c9474e2c092156d7c1960a92d38
ze500e4d3b5dd7077899f2930bf9ed76c0bc55449143c6c9402729c0deb1e5cb0869bb1f7682a9c
za9ad3fbea5522a4360a27b8188f41c57076d9bc73fd4c39be2e783f323e8790d99aee70c2cdd20
z42abb2a189e2331fa87f34197f200dfe7ca4414dffbe4009e01f1076b186231368a891c900ebf4
z05168941be01e2fa5ebfcb57a40e50227ff4778fce5c29aa4d69bb23388ff5edc01506da5ffccf
z4ca69dfde228c74ecdadbc1b904437586e764d40a1213e2e8b45f2fe0afdcf3fdf72da63e49658
z6a0e8da681b4ac401b5fa5d19d269771c049d0556cfa14697ea28a10bbdcf3552e60df8365de5c
z2346476e3cd9a246fbdfbfee0e54dc59946f7701457d40c169029bc3f9d7e0af2d7155c6e8d0b1
z0e73a136846a58f16dda418cd4a5c3276015900baea915df0bcb9ddedac657b50bdc3521ffc920
z7d91656ef6a1fa08ad63fe44e5b70db8be61f3bbb560579322e4ca93ff13b0064ea7c7d375e99b
zff1e6e86c09e3c5ae9fd2b415c2d1f19302f85a1a2e2c123f939e359b0e9fb60e7d1276594c915
ze59d9ef6633ae49f2cbb7941491bcec0040bc1c67b8c0ae84fa6e550a0ba73d91db84768179b26
ze6d490711e5c3c1fde13e07b5b0d6ce6e1e7d2860d9c827aa039b0602e137b894884a87ee943a7
z955c9b2fdd95c213ae76af9220467387fafac5d6dbf01e69f61c06f654021fdbdd6e6fce9debb1
zad8b31057f48dc7766361417d0fc209d9bc643033e9812f48649a028cb1bd8dffce586167e170e
zd860e5436a7695607898b5c668d2ce1873513c886a6e869c3584f6733bc30daa7d8da9e70369e9
z37e74f68df827abb5b75fd0899be80863b289072121ff72856e0ef6fc17ce1874d10160b107607
ze10753b784e96c4ae3c0c13c134801a2180bf7fcd51543243bb4bb29df8ef7677ed146f3ba9d09
zad005754aaf2230d2ad3ec920bea0d4b8693b1636c97667332ebdc3a38790e44b12d5c24df5ec6
z52d35e3951e0c0347865862af904cf7a08d93211e8cff32e62ba931602a67895d9698fa236d366
zc6aa36add9d1b51b3e933db981e08498774a82ac816c22da76ee4d9d2450dfc656c0ecd0a507a4
z0c49acc65b2b07d99614d50410029ac48b23d5ce8f38d26b71b0a6a2f177f4fc29a745b58deaf6
z507c105c2b89ac45d15edaef1050c80fff57f94e892d4f871faf2a45320ad1f932d3e0f0e37a69
za1337c4cd2d6cf5fad2c3b4499a15b6465e5ad165c692938700ee6b6cab0aa28605d147fe34a0a
z39f1007c538adc68efc3c711dee7e406ae2e4342bd300de5bb357833d902b2bf29336088aa0a11
zc27f3761370e881d8ba5db47b172a15041ea70a86061f0793657351e1bf668e728efd6415f6c41
z1749a715934ce74efda6a60ed9628c0a7b487d6290ee4877ec85821a34e587397bdf378d5c11b0
z5995961d4f14c72cad5f96f0d70de8bcf146765ca34373a6ef8ecbb460d6b389cafcf8803bffa5
z4772985b1ad8af79bbac363f6cea793915c05a79c55fd36698f1038fe97dda60cc9e1f728c6665
z3467958768fee5192a6194289e6e2ba97698b619c4d9f084075fd1dd89128b49cba9ea68f613ef
z45b0ffcf96d4fdfff78bded9a231f73756912bbbe06309c53de64fbe4a3e16504d43e6cac2cf83
z23aa3dd4332f697011350d4c8ec51e6cbe945b719a780ad841ddbdfa92dea44185096505d2f073
z55953a90c374015d1e3c6e45a0448f5771ccd161e42e8f379245993837394b654165b351deb916
zab307ae2b88320bfef90999f71c56a9c35afd394f533f83f0a9017bc3e35521dd85cdbd0df1820
z6b19d1c8e04e2ac2c80a96e5ec5bd7cfbb324c571dd5ff3c8e56b7d77158544b08dbbb984a16eb
z7358fb60c0d531a81d090e1c8363ef2e30c1c4a61c69ab28c5eb0b9e67012a4904eb62496ead4e
z0d1664a79790d53ea49accec486e3109f8a5fec50860bf881119a63663be595b4a61438903df06
z7222a26365d5b6d230d4551515418846fc9b3a82ab7b562cbe67d3c15e5558bf0affa7bff404e8
z4fe863e655f5309c0659634b903af3f9dfc7615cd1b2252560b6e062ec9f26c9059c0372b72fa2
z3c7a6ac4e5464516559f3bcf120466c44dbc9446a37728b222015d1a2335d511025f52fbf3f05e
z7cf06d6b539b3498a676bbfc8bb5709b5f78935b5adab6fc5d6f85b239aed694dd73f7de7af346
z4fd60d411da607650839b4a0a447bab40bd9845e8efdd9c1d94d1730e5a5d5ce0afc742ef52688
zc325e8db7fcef7b1d0ced1e294fbcadde5755c70155b4ce2144901fd1d21fa1454a140d60c3bc3
zd23d9fd44b5e222e3e64adce4e09d5c1027678955bdcfab98bc8db0b83bfc819ee7eabf8ee71f2
z4dd588e9ad33f3da848b34ca34c4435c4027b6e7cadbf66047303b4e75e6814421e844fc10dd68
zcaa3a6d285a3604ec1bc33ac9da982897406c2ad8e267c4f4902201075c2aa4e44127099b757bd
zac73565405189139d571695d51b22084dd11aeb2c343fae03599d6819a6973454d86e993d53101
z3a3aed3b77a1e4b026705b0769fbf6480d3d940d5f2ecfd3eb203006a8497b8aadf3dc1a9e777c
z16bc4260987d345821840f58e4c07f4f9301ba9b67da042d3e9707616b19555da155fae79cd9d6
zcb8b6b2e077bafa446ca9f0bf07760cfa48d1a48ac4f4fd8946abda1eb677c942a56293616757d
zb0ea420a6b259aa4d04b0acad85a2718c3f3ef6e58a946030e9c3da2bf8017b9f50d133c142ed8
zf0f142d9e4771a748745659f80e87bb90aafc5e9c6c277b29d5f2784722f5e3426deb30aed49d3
z1f3d5e183bf1c42edf50ae6a6e3e2e9fad3fc5c37ffa77599ad6af7b0cd2617c6234d75a8d8f44
z0a3b97d47cbc3b947736f8ba34c3086d26f0f51bd5821f35fb86f0c72250a05f1cd50cd29f6b5f
zefb8af249f394f39006e5544fc58c9128aac47ae039e6443d5e8f546f15928e1bc78b24e5f9ee8
zefe69881a147d21d2ac702161c971964d9e8c0ec30a54b52ec1af14cb11d84d6ef44eb7d2a7055
z713f7bf95b798a4955ee7d6db050f9aa4fec849b63c8f17d1504ac03a87888cdd9a9e1350f72e3
z1bfe280ab69cb4db44f4109f12f74ef0fa3ea7399181573465af45b7022959948075e7ab18ba7b
zd735838b957c38706a3371865bf76a0d21fe2e0d4455ea392ba673ec334207190af5105200431e
z39aa549deb689058692d2f2b4e2782fd904b3b1e2f96d3bdd44c37082ee7e1820f056ee7ba298b
zcc2f7461f5ae97c194943674330908f27c1b657a5ecdc186801624048850e39396d328503aef59
zceaaf790cb4c26e0aef09cbc3bc25657d4f3cb02185586321bc25a43938868031eee97329b62e0
z7778b321abfc3320d28f330f2207f8efbdc5d227b53106194c915c13274b3a1878100d55fcc3a1
z1774e30eb9e8fbca57d1dfcb3c6f1aa347c00a26652954f87cc1be51afb6a67132f73f81555583
zff1209365189941dd4cafa3f8eec5363b4819b389076d96648b99c00d921dd70c4b0d12ef496ed
zb9e77a1c1a2d47702c5b78065e31b09bcb4a7dc812d4969ed3072e63ee92dc4ff182496bd5982d
z519ea35fef28bf5114849b3d04ef363a86eae248c907036a73f1acb0e44c2be714712c55335057
z7207026e614c4c9dffff31a1972e37e52710cc2fcdb0fd6ff23a7d4212716d138a0a04c3de5cf2
zdf7691a176106786c03d8ea28fd71e2fd726a8bdddd4f05e3063f63dd6302638ca500b9c0364c1
zb479129f044333cbfdbc6c4dc558f715c82ead4ceee5ae7ad842ab51b7b1d516ded48d1a60a234
zae35fd202b0c3c7966ea1f8bf9ab0e038a460953681f5054c11f28abfc388e8bee9be8249384d6
zecf6c8187747c8682810cabbfa75e7e53d1384c972e56248cf9d734c279c4a8a19bafb8a6522a7
zed240e3e7a56fcb818ca05125e51a348a82f04f72b2fd146a136bb3704f5be267ca28b6ca90fb9
zeee872be27a7bb50a64df4ec421bb1788da28beeedd6c712b1e126e8bcb2b56ff4f931503ad45a
zc4c6a6e0ce82e7e29ae78700205428b19ec2da26ee27e45051c81bb05266dae27a14eb96582280
z0661b0201c43343cd3da105d660fddfa6cc01218e75b62bd10c0a2baa2e67ada6e761ddd45ccd7
z6d8209fab98706bebde6cf3080658c26f0fe148a993ce5b4a9ebf5c1e58de9cfb29fcdb0ad8406
z9c58739136bccf18bfaefbb2b2b22581aed625cc642936b8ee7427648fbad171342cd53be7f6c8
z78124b32650698f52e27a7b475ae1904c415701b4ad0befac8e3dac48b2b7a46bfea0beddb984c
za3e9bf1438579abe0bf9024c6ba7c2b4ecc058ff11cd7ff2a6b5bb3cdcf02723a4fa5761b563d9
zaa70748d18da17397d15af1431710a772b5790e042a9fb04425d09a2c80bf93a98dc3f9a4a8a8d
z3cf7ef69808b5753a33906ecca9159abc495d14fa3a781e90a9d6b11e4371e0d5fd43ace6638df
z6c896951fd94b007da3dd1d68efb1f2e20d7b9cab90658b280cee6e101d8ab71ec22cca4e8405b
z7a9373f1642df4c51ee5edb739273605604a651ea73c7b1aaa0b42053a46f90430d4902f7579d6
z07bd35de12e9e4b0263cda174b9511945be2e643fda1d4c5a2db4460ee90e225516b73a65189bc
z08f6aa1d28dec8bc5954c603d5cb748feb0d67610300fd17c4803a5c82347f71f5a4f7e257ec37
z16445b524436863e7b692f602c12933abe0eadb98ee3e0c084b88c80db832666ca2a8ebc99ea6d
z3350e8f56769a377219e5dda4cb2e75db3702a72400b6861084155438eb6f265b36827dd37cc53
z99df9440282c2097777df8a6251d33d9bcb881bdf1468005736a8eac18f7c30c3562e37e4b9821
zef1fc08b6d5b6fccef2b412958cadcf7ff2119577ee79bb9b071e8123591b1d7400c7844189e5d
zbcf46af228e7c54603ba24dc763dac1ca64df899355f74a207e60d548970fd1ca01966bac657b6
z097a2b198853a25fb0987840ea3570f287e80eea30f2b7bf786af964bcffc9a77349c8c3670c70
z450f5a5cef3f9665538ba66a9b8acab28f24f2807134e33972119906579a2f11c14c3bd24bd16d
z76720849021b9467f6f406e1b5f37be9a27fb18d6364e890aac6e0a0a2cf9f5684ab9648c8949f
z6fc03c6d49a8866aa09982619fa4fed88bed5cc98a8f15a61cdcd067a7699037571bea55aa73c0
zfd4e05dad9a75409296534ef348961d137d34843a67c0e7b2a6d8f085a4683739399e9098288bd
z7ae98d4d93295936302dc592e3054400326f2bc6cf14cfab03e9520110103e60acb434f8a7deb6
z1ff4c8b956332e638e3330a1be9f23f1f8faeb20b7d42ca25e8cb7704ba1bcd06fa9625e725297
z9ab941698788c0e14ec4812bbf307b491f23339a16ae66fa117d88b30a7f2916d4e19faca8dc46
zf95961007a130d081d9318bb73a93029081401341ffdf83d4becc9ae4d4c13cd7d0595c5abb488
z74d18666dcb597803948adb8269f61c32e8e9e5391616456a81163809522ab039d75c094e2e49a
zdc6266372233fa0f43837ec372351b8dd2b7937cdc76d23f64936b49aaf556329c2f06e30178c5
zb5ecb1d5f8956b315ea8889de90791d3dd6975783cd81b645ed443af015be37dd42353cb1b9dca
z398f3fa3fa674daca598791158b2affc088d6146ba5988860268fbef1287b1169845f64139180e
z639dd017f225154c8ed24fd79b453e9b80e5c65081cc8ca3f04c7f4a43e46fdad8e0a9679e5fcb
z79c7c0d029571bd6911e585eb348e0d240e29c76166f4946d969cd1ae1a8076fd4cc77e249f409
zb4e4d24ffab87b50aa6e8ec4968fa878cae63ba99a7e5c42fd3e235a0775aa17322ebacbd84418
zfd1dcce3bf0c737ce97a7484087cc0c3865bcfd601b1d40bf4cba546c9506bbdf1702cb668b07a
z731fc19babe45879a0ac84e44c75297f3ba2634d9bc8307b5049e2a5078076c677e3cf8cd51782
z7c00b013d762e38d9a38a23aa4e7bda089a50357b1e60d62cab596b5b6bf4eaa199ee76f15dfc9
z7907aca1496e9d3b9dcf546a409337e6b397cf158ecc619d0514031999e17979ac24912e206df4
z9fee0473dfb134c6ff5223b89b9012177fe7c78a5091a5f0a3ddf788979a536193b1d7c0dfde79
zecbe38b93431829d9c37c4bccf2124c2c98f76a488c57f08023806989a28af0d8bbc080cacd7b5
z902f42062ca4fef0f0530f8e2ee89e310a8cc0b6452ddc50ae3c6574042265d7cd3cb76ec6ca6d
z3cbb34cfe69ba3f5d489ae79b98b6ede94235a3492bf29eb1972c9c7aefe0588bb65be97ffa995
z881ef87c5730fc6f5b527b713717eb74765a1e4a81ee65c3224b8f60ce595463b06c18ddbf96f4
z8e354b2c680e22bbf1db8220635f4192c86f3f13f61403ad4963e1e7949dcd54f465598ebb2c0e
z50ae45352c0b5c76f647a75da730e175220e8bb048d23b0128a8cb66f0001fc2af1ac9847a4cd4
zbd3403466432782b2c387aef493f474571af36f5f45a16e4eef5fb2c208fdaf26b885e6101edf9
zca64b61a01560a0ff43b72466a8f6d728b13da36bb1f8f39d4dae86cd3a3c956d3065d64fa2b42
z00327a8fd9359782dc0cdde84edd4a621a0877ff36b4616e66f5d77b6499aabf45ea800e0741ad
z74c29c68b00ab06f70385f20d601d5665a52a9b1895eaed3acab7b2b11eb2b256a42a428a65c3f
zcc80040d1f66ac13cc6a3fe1c0218cfbf2259daf738b3a8e60a5e009a87bbe6c6e924fcf4c5d75
z5359296cc625d6e56114f12945b027ceef6a43c6fea31d7fc064ba3acaa7771c6d77f3807cbc62
z30e0e1eb1f82f77b464ca045f3d95a721264b344e71dde65dc00703be97cd99482e3774cc3d772
z8639049fd9ce19171a0c5c87bd1ca48c35e23ddba62340edccfad797d498030bce88b89f81edac
z503194f6dd152677f23f84ee397fee3dd5e8c8b18283de6c6c161164fbd1b1177ef0a9c90050aa
z7f52c24406ed965b0e68933453875330fd97f9740990bc3f3975f8ebdb34af4bfa961458988ecb
z2ca9e80b70e196764cf4e0af6aceb12c92965b9f588aa8ee5c5b4936cc90e2765128648a59bfae
zef1739baa7a28cf296d830d5c5c33c1295119b686b2d7e0a2a4209dd05a389b1452c2d9d24ae31
z33a5a7266b1bb596c16445a6490390a15f8e473b31200b255ebf5e28ecea03e1afb86b800cf085
zcf7eccdd15a4c4f2c0e5297416b44124be2a27c51710ad44d432bdaba391f399c785d5867d910b
zc6fda6c7ac271cdbef9488d6845603d3ba3ae75a636fc7c3e60c9311dd9e8ee4d0839b7290a39d
zf7f1cd51f63e6b9526993987f9d16ee765b3492c054ebaf3016b12a8fd6247d41b960deb5ec3e3
z5a0ee552c4c52898e950ed57c469843c84bad34350fd9ed8a1e680d2e1ede51995841b79ab0cca
z4a3645d23f56ed01aaa104b45555cc43e95ee46aa421cf01aae143f8f9a60d2efde1fe0621d513
zb9cd1083fd4eeb1592c1136a9e897d7ff334d1b2142fcef8184a49fcfbd17fecaf3b116a2b07d3
zc20f45797c10f0cd0fcc286153de939e3a7efd4ad20d86332192e4d27fdf3af6783869645ef7a8
zfcef0dfc27bbe6af76c32359e36ac9ff53b61a7af023fed224875032d928e4cfa3750aea9f14c0
z23e5c00af2d15412f8f04485138f6d13db74bb1a01f7799aaf7f13829981b282d88de3a7fae92a
zacbb78de3b086f379beb5b12f9f90f0c4e60d7964f95052b891d195704d33e0d139f5b4816c10f
za5dcfaaeee277106ec362ecdcef2f334a502be917d02f8946a0d0c48cec4aaf57f38a52b7e7fb5
z0a012f604d822ecbae0e68270b9cd893b51d2c18931835987e72a49a76fdfbd14d142713e7aa4e
z7740f84ca30fa06142a3a021643f14b16c66259198bcd770068ef7da82da0e8d498043067a3475
z2ad6b9ce60043bb142239a2dfd9322b1fafd8d785b359fc24f94822b9844d8ac270f4465b5021f
z9e1a1025ce5fdd104ac192405e9d715a6ffbf74f7dc0ce6b232f1b7f7f963f473da65eca4916d5
ze220d39ca3e197bb1431e6ce7d1bf15204338235d2e42fedc426537271162602f8916e7ac01b6c
z2d0c2f9a8679cee9084bd38bd049b8e41c9c88d4929d6d1f93c788db973d451fd5b8571f4a45be
zb32356a5c64f3f5d2256087bc9ae1d5d025c52d1c4d23a5f0bb1692882d412b5ddcd9cfcd5f442
z304166e2f157edefdf9c2c9d45a7c13d91c8daadfbf811bea92066a15552df20edef4a97d023cc
zf65c0694db871ceb5fed904bdfe2ced51cc732dec7ed6c5211b114db27e41a38f0d98ddd12deb2
zf7eb236f8a27618618c1c8f1511d2f8e7be7c1cb4cfd79b9830f851ae452a7aa4a4dce927f8c68
zf9593e675584893882f6d60ecb4326c6b23e86ac8e13400825504b5d618b53ed42ed11e7fa6273
z8b65d62c497fe5caec37fa435895ea752454777e9df57da431c10b47a0e57a3b3cc8307b697aea
zc628eda949efb0bada34bd2280cd0c9f03b470cfb3fe934e467788ff322a18fd8bb1e450947f99
z4d3470d0db82cc6e432653e99711576df23be5f2676749c946ec5b9a0d3e945ce058a1bf1c0edd
zbcf7a8b2d877e4b8f9f34a57e85bcc1ce206b376af88af9d6d0754294664c0c92dac57f198b281
z851a079e1ac055ccb69e56b398847f0c2e5f67b5eb1dea1e36aebffd8d7e016cbb21f46233e0b4
z2863f14796d4106dbaa16f699245d0cb74419269e99f3d9751b9ce7c3d93e00f9ae047285a92f4
z9c72175f2a476b4ab9b3202ad6f1deaeb9588b75609ea12821037c3ac55316f7ddfebf9eefa892
zf1c9609f2873afaf5bf4e755ecdc8a2dae689e7a381f04941fae31e784ff8b1c875f2b9bdf87d2
zb8c8b856b8628db6010b9842294c47aa8b35516e3a3fc20f9fcf507dd02e49a7c73cba12be7766
zc5c4994e27d33a814860afc3e85cf338437ca7c75f1133797e8895643e32b6eb051800466a3ca9
z4d7cbf1b4081dafe15c2e9eda4bcc2b81e9ea5dbaa6b6ec0f2f81d244b18abadf24a22e9202209
z651b5e05f596cee8151a5fbd76840dfe4eb7b656c62e5b5a9747d406c523e384f5cb917f3095db
z5abea366b081d4a69163886d7799fb07d4b894f1a30070a2935de6e4e86f068ae79eb055e23aac
z4ae96b00c164750b1b15e4e1928b4a258c894a3c6299afc2efc0a6c3eaaa9e5ee1384ff6fb76ef
z3cb1437b7046aab316b3ee2a4c0582eb2cd2a2c67606be58f443a984d891828bcd477e5fe26912
zea3c968b0135d11e19a69f50c46fcf22f7e0036a044233027e52711e56ac1f93a14290728f5700
z57ea3ac7a6316fd6209aeb27b15b5a6167d97c099b6817c8e0668b1407dec658d4df5fee045521
z4417bc118808f3c1ebef1e1fe848f1d29a42fae160a14226b0600254fc49ce907db5cd4e20fbe5
z0d0ccd00e7ab589e043cdeed8600484abfa73d791393316f279fed97f8cef1b473ebd20baf4395
za3995d933ecd4cae52d68717bbbd6794e29e8d1b7209ae5c2053e4a005e8c85e908856c78cd7a4
z82a28d96d76ae3031c9879dffa641b80d1214085c9fb646c4fa3a6a507f8e16351156635ffd4e9
z42d3988ee4030e4123e2c57b40a885cdf5c4402681a3d408f37121b2436735f2edb5880ce0130c
z7d554c59f45b9188028a7f4940062505267dc0bf529891272c1af2ea7a7176897edea34305fe15
zfbb0a86bcfcac3219a1daf5a1d8d4dc02714930c6cd97dce4d574066ff2e39879c12fb3764eb18
z360246289f73fffbc50fdcca627b3a1cab0ce360534814185d4e98d61fbad6f50e350daf6662c3
zbf004814271f70a44f6d3df80b19331a48afd5162b936a8659906459e6245c1b09e79c4532db79
z3c0d45cd21b42b701cb9a192ee4ae1cefe9a57c27b030c8bb68db336d2a9b96a3f7834c327be5e
ze99b890567dcb5a56c720a2198bd5f78416745e38163f007c12014c8c967564febcfa7084843ed
z2a9ca93ab205c291b18a9ee90938bdc42825265028ca7a56d383564374e26c8a6384637f03ea26
za1fd193a4597b3c16e5f877ea457fe64a30b7297ff5e936f2cac15dc741f5cffcf31d5ba75bcc4
z1e69dea36e460cafc9610175752a3950eceeec21258d0826af9ddd8bc529709270c39cc15abfc4
z914d486d67b6a50ab34372a7b059b62b0b958abf2aeff5c55c950e68513e03458ac1b0e33c5b7f
z6bb03a2abc06f2f419ee783377ba20e1bddc6b8457298e71eb746820ebc0291406e2ce4c4a143f
zfe93359c218c293bfeb406f90c32ce831ab904855ab29bdf93d84b808ff0a6c43041943dc3a316
z04aeb347a31d930225f838f6b3527280f3da649f83b0e84029c05db90e90ae6217c56c42a59d26
z5b9369cbc05af3c2150fa67b59b759ba23afa6f051c5b7524af55a33e47b1f099bd4335fe6ebcf
z9b55b44e7c25ee2604b58cd6fe587c84658032792a3f5de8dc761100d7172b621cb479471c860b
zbf23e7ae7d3d2c3629d26449e66bbb482c912146f5b3db0746dac2739f8a025f3335b98c0b0547
z5b3bfc0c0c79cc819b0112c1c1d8721f69c4c6c1ce1d4ec84b93e43612cef3dae160e439f23b5e
zcf65a499d8c67dd3bcf193337429b7a3fe75d03985b74d2d174d6155e89a352504add516e99328
z623f494e5a65d54fa2bfecc6545123d20a435e343f8bde76dde48bffd45c916da4d348edcbb675
zc61c21237acf458487503a036941b89b931b010d5641c639c9d80dd6df5890ac8a8746f559fbaa
z598926d447a047a954333795f62e23687dcc37e5c018523e430f717600f8b0ca1b57ff6d598d69
ze6764989b656921e4b936403844b4806d25ea1c7a1668b3e237999b43b71b4d9cdadf44fd739a0
zdafbe5927cee733e3e5a90c1614758648638f6eed0655206ef052eeea9eb0c79185c6fca5802ef
z4c1b6611354ca51caacd4aaccd6ef35889b6cf3c25f34a6510fb5b724ff9770b8af13c72b721d0
z0bc8b650068f3136c6f220faaf7358318fd25ec5994457ecd63b786072289c1ece4d3a94deec92
ze0bfeca69fe8c63af5f21b3e01d1afc5544eae6c6f2fc0cfb0f98048243d080c6acab08045a536
z4cf3a3f77070385d78a384a721eac4fe3d2d7e686b903aaed1b6ccf1a53c4b8d8541af09ec1aec
zc8948f229b16f91ce24e47d87c314a57e0320e1ddc6a4bc0c9e0be8de50ff9b26bb4b3582f9b3e
zf208cafc511ced9a9ba354cbdf573dcca7d7b68f452e1a7c6df387ae3611dbdeacda15432f2cd2
zbec6a5bde39f7ed70efdbf7a9b013388a505a9f23764444e552d072cf30e31db53318f73fe4b3e
z956ae8a0573097c913bbb477a48f8385adfad95dd15ab7d43ffd738fbc3e545e44b2786f06faf2
z95997616b74109470e6f40de257c3adc5e8b569cc61ee62c83ee0f56d3cf28b56bbbc51af86374
zbc3e5efe9db398e58ea620a96b9a49f0e1a1b1060dc3bf1696ff88b43b6bd70e71a376cac56b2a
z25415f02c8a2fdb1744e547e111563b1410eb58f722f47fd3a9ee6427d702793235d7f7be6c8b3
z5b20d2196e4b5a3c1c5dff059a31dc405a5ce97230f8a54f58e7c7c3c165014fbf2ecdf6a4e9b1
z613128cc1e301c4601a7f58831d76d42f3d6414cf038e04c9b6ce9366c39037a2fbc2ca2fa5202
zcf7b4f1c7b266e3f4ab009f19f372f4e93e8aeaf7460a2f85c8920870471dcc0b2c86c31a17cb3
zb37d79dce05f8c207e69dfb106a3608297fe9ef2868494ae621993036909f2ee296afeee131576
zaa3d788c609ef1a0f72ac71669e2013a7ce1ff894f7f2522a1fe43e3d6ecccba2d65a881daba77
zc0543d7279de8a5c7e4b8a88eac9276e14fa2187b3a76fef51fc2726596afb9818947f80ffc2ff
zfdb4163232147960b860a82ee43359422d24a3738915d62c1201ce8b5c63ea524bf587cc6e8e0e
ze3d7bdf9f2714038af96c97a8952a6fffd938ac7bc27f7998232960f3d6787dc48f766e9d848bf
z4985976984fbe4e32d8587fe570bc6666f5b9017a14ab420df767dbde91bba5c98832724220b53
z644db553d4514260c25d4e30a9c06e2fa61b5e21fd938f267bc655a38aea0c94a87de7c8c7ba5f
z33ea0c098e1a9c32cbebfcb3d6b092d432662d48cbcfe32e4c2396ab448149b3090d0d9d785832
z63d16f2d79a086d2dfb2da3a2567dc938e97aea01089ccd0f57eee216ec158fe451ee4812c02fa
z0b3bd8e92ea275113e0abf2fceb8c2dd1f406786ed75cccd0e52317abd03ef55bb4930a0d4e486
z47f93417f21734c58f25aebeeeda4fb29deec53e5d69f1c2a25033580c7a9ecb5b54d81a138a50
zc2338a987b87c5918c7435227aa30648a8f4be6af545c3f89b42e8c9e77bcaf298e9e89d3f27a6
zc31849618c7e9f10b42622c399cc1e72cfbb1e6a77274a9784e9c74ad34660fe099b9e57726ddb
zbf0cf859ee27329e88f4a587e9573d2a8929c713eeb8c09c0f236fc91737b9696cbccb9ad1f71d
zb9bb1a13e32099ecbd357caa5a0a200d9c459a2c615cc12e5126e98bd2bc63ef333cf29d50859c
z2bd44fcc983b59ae283f3fbcf5165ced3c3fadfafeb5bfd2b2b167d4adf541d3fa02565c83d7c6
z171dc98524ef44fae3241e06c932979c96d1a27b6af36022991f6d78d3165e844c41d8ca091521
zbcb62fcdab7645713c4c08d394d4894ee30fd96e7cf18358b520c517e94e2c669e8365b96d72dd
z1b3a68baf89cca6e50136b2908b72a6e301a0363e36609fa35392760631254c2fa5d0898cbd875
z02c590e0303c22773458b9fe623fb1fc519ed56a1b2835412556d9a0c0223545bf77312d62d67c
zf5546ca6fbc634b19210f7155c9432a41c238d4986b24269b4be0c99306c9e840ccd1267d5228f
zb374f88eccf3b06d9f556464ed042d224f9a41d1198bc6b86df47c4cad076327f15c8b7fd7fdad
z96f9b3611bf097976e4f9e56c9cf60bbaebf5993609fcc97ce08e970867c6c3b2ba25a26674a2a
zb7cac876a5a2eefcea161692b3eba86dcc812026b93574e1e1709a33065190c54785c05235d7d5
z09ae26878ded065378daa5c82ee060b9e6dde8f14aa10adbc5e8fb81beaac69529387c8c84e846
z14433e45ddbaeff7118de23511be9aeb90ba2a79ee4dc0cb4e0048d328cbd7d325191cb33637c6
zcfd5f63b3023f9a8fd5477a87e5b69b005154333bb8b098a2e306b9787ca438ed7bf4411d336dd
zfb00af39558e0c3a1e3741eae7448bd3650ee63d8c5b92b559705e83b3e6f725f28e3ce8e5db2f
zbc8cd95b8d54f84fc4ce1935d044cbc48aa34df28eaf018e95a114a77e5901172424ee35a5a58c
z42e6b53a1a79807dd85b12f54a8dd10f9d331e681d0e4c908228b475025f0cb293152066adf451
zaac1f3a2595d7f937f36f99e8b0926f8f7d70b0a4f7bd066499a935a0a2287bd8e68776cf786eb
z4f6b15be18b0372f0232719aab1a6a60d5f1d6cf114ad1bfcb543fcc73bbe1c61972030072d762
z6a767687954e180586c75cbb72d529bab0843fac33f7e64813927e1c567b64483a5e0447825d12
z8400edbf3c33950491005cb6bb3abb898f6985f184c5bbecebc8dd2d2afd6da79c1a3911653771
za8d215fddf9a89c642d54fad3dbb4d3245b13da509fee843088477c1ddc5f04868e1cc5f307972
zf7dd609719cb9aff4bd10cf03fdb9d89abec2ee5b9eab4b8aa84b0f8c8daa415e9712b4ba3ddfc
z65528bf092529ad1e0af6b966c0b045a3ed2fcf52082b0eea380c5dab1122db28719060f9ed5ce
z80b8eb6f04f462fee7252df4319b321cfb6c890dfa6c6ec3484e8aa851fee858023caa976569f7
z6b37155eaf41c28d5b95af3dc96403dcf86c2b6c24a9604254aff3133c1d354478fe088dff3f30
z165db8548d28e3260ed345eee2110221b10dfc4fbacaec523522903619c039ff805ace5269664b
zae3637699242ed7743c4bd38f4ab55e1b36bb745023f1d6886ea6626cffcc2ebd62b6a81c0d72e
z43f0fcf23531efe2680f0464f618f637abb571919ce7623652ebbaf86ce0282c8729bb6d88679f
z77bc619f26a5611ed5d9e01fae26f46c6049de467d466cb14c15ae6303e443faf3dfc50dddf4a3
z11feeba86aab5de94735c149bb95f54e746035b81d4aa030831ec280f15b0fdc7d5beedeaf5c8a
zd3edf8ffb0f494cbf19f41b6467134d68870211e53dae1b7aa801081b849c39e1939efa6be7ef4
zac760546fefa9381067313d988f1502a01e6f4153dc97fda4688a919c003ab6a748fa4fcadedf9
z7f974582b62ee9bad09eef2ffb0ba0b1a761e7fa89d7fb50958d60af8221e795424c4e6a8934fe
zdcc07cbbfde46467cc75cd296e2ad745ab8b32c9e539bc69b7460039dfd22f8c3ca93377f836cf
zb9c79d830fb81db2e16784b842e85ac1b8c0e1b0374a6a9e12b1efd2b64c952360806c97223d7e
z5500243e1a70099c9086cd77fc423b1da138b52411501e44ee5105150dd50a829689ee94e97da9
z999c94e5dd5ee56935e5f13c86ca63b4da2ae195e162836ae9fec8baf9f1a1e986f6a6bb18359d
z755170b89c5d140616b5a8a7f46666954bee12148f1dd4e0798a7185d8440fc907747f59f3108b
za56fdf4fbec6cb97f1c1742a45469e65989a164d87931f7a6d3acf81302799267cc2e462b72a63
z2e2f3eec8fa8e5e51a0e483aaff6bd7fac9d14feb84e5fbefd0d5744e4557eee7a2963d069d703
zeb38c23daf2274c1f8795e720339b20005d10b825726481b81779db93ce438d9569173d25c0d89
z71f6ec449b53b5d1f5ec2a6aab2a2909c6c473305719dbd801bca64f6ffaeeb9b65a6466748667
zcdd4aaa4b0e5a0c5c830598f3a356e965808198bae61dda7785933689aa5a85bfac9499379ad5a
z2f5126e10d184fa29a8fa795bf9533ac7ddf9252fdeb346e4b4fd517125a610840c983a595bd81
zd9b2a748b47c71a287809ee92a70564aa41b601442a708dd1ac17012d3ac23cfe522157307d65b
z516c72f38a45e290e3049f4b5dcbf23ec232853a9547fb7070b4a6c179c302c85795cc4756eb20
zfc266645131f4bd11598bd59ebc446a353f8f640618adc4999c8183a515a53c94d11cf21e4abce
z47d5a8ca0e188a77b5e137fd194bf4540ba538efee3a3a4c4e861f432abd502999bf7a7fb32e7a
z664ce226f60e96219f73fc4d073ee888a940510757eafb76588097208dc0bc6fee21e32c2958ef
ze3834767e6c9f273472b15c52ade850a01a5be9b6b49145982f060e4d8f220f066461094cb62d6
zc501982a0dd828387f65f9a058dbbee483e123c12ea1dc6240586206e4fd196bee76e71025e0ca
z4ebd8c30d84313782832a5c50b94bc28af33fd1289a2f87b19c1e1cc6a41eb9968fee80548098d
z5766dc9d9af55ea4d67de909e7bb3de2df20d720506b7c11030f27d38506cd10f0eef13467086a
zf842401b4c22d2d9e9ed69d76ac5fcecf5c1ecee4f0930f3238b732fd5340c3084e7008ab10483
ze1513d55ad2cfc5f2266db9245e44f4000a4bc0cc8542e09e8e62f0ff6e9569e65014b84c53ab2
z73ac62dc46245591c6640a9fbe1d0ab8491e1c203663d00654753047f8b348de301ea9aface3e9
zceff8bf4dc72f87f40c5caf3186257e1234ed30fd7d5f2407cd716a3bcc074f74929250c47be93
z61b2880938f50d48c48795b24520240554572c23759b0acf066bc31b8e8c0c39b1abd9bda6002f
z86afd104ada506843f274f12edc8e3db2dd5e290c3de85e51c740111524c132d2da4ebc3772520
z9c99e20f58c0b3cd5f338ddf8df087fae13007a81c3bc59e7472ac85877a31143e1e72df560eee
z52db77e202e0bfc949dd156334dd0904cc8d475cdc2bdfb1024449c24b31581c11dcaf28a93860
zf2ece15079291701d33e8223afe96b54112b1a9c5d70c3c7edace7f2284ad450a92671ba9f32ab
zffba4288ed4ba91ecebaff4718cc76ed45e23be3b44b3c624e3183d805afe5c4b21c5f0180c2de
z00b35f97d6d432cf56ec8dc646531bd70281b339e65c6bfd5ab24e04b7013a82c2923e88d412e8
z802299e82291c51eb525413c3bb98e4da672aeb3a02c87d97aa7dca057b4c0b20fdbc10bdae452
zd647b83b6a0b8d9f3d1c545807431e84020489d56c2df931f0534a629dfb327de90b4d7b99fc07
z5be27f752bf0c64cbf0584623098d7257c3538cb048a6082f85aa167c42098807886a07c8e24b1
zfd1bc8566759bfc43acb4b7019f6e0c52664c25f6e2ca7a19e52130aec098ca43ce317b461a0a6
zab212b420a6120d50c49bae1d25bc6574282e094214ab52b28320c0a5304223d71f3b4785baec9
z4266d38461ebc7f8820a355e96044457dd1a69d35a287d876a54798fcf37830ac395d72b3d128b
z2fa31066f40d62c6a7e81249666070e8657971088c1c17273a21f7421710854494756bf03cd4ec
z95de270c44da674685bb62120445dd030cd242bfc319d78295800eb3840a1e0eec705ac6e3ae7a
zff42efcbaa12cb0c92f350e3864ab0eca78aa996cacf157b20c94d6511925b4ceaf4e8962708eb
zafcdf22b66c928d3a326b93af3f9fcbec7ac5e7c153dba055804e12e59f4a60b030c89b6f073e5
z38eacb162608607b32addcf28257adfd95fd6a878cab97fac27622d3812985da0e76003ce62064
z645ef27e886c1d137574cfa1175e45892d193f9cf6b1c54269f1a51c45faab7cd944079642f9e3
z8d86a257abd263ced3493286d5316f9ec837e5d478598fefc38db484dda3438d70db30944fd3c7
z91076367288d87cbad51eeb7037aac4cb78cf7372969ab0f2584b57348c285401ff47ce9fdfbaf
z72dda50f64bb8168006e4ad9ffb8e08decfb30560be73b250f83ce29f44f4bc67d39dd8431ac0b
z5dba7017dac620338f33d32152792f6271e3798ac21b816fa35cb4c23462aa7ac9f9fe7d05dcb4
z82227fe53a105658e015384fb65171b3537f38044b466236ab631a530bb084d5a3b1d707b9f721
ze8819fcfd1323c574a27be346d2bd6de206059d346152e9d91a845783011b259c3765bd76fd2a8
z49b7674753a8fc11c510b0223293fa1c8d4896edd613e4b6a2831c485eecfd7d97d644284c6237
z284e27da742df0ac7164ca3a8a9444bc1e6f8b07d927bf5cc8d03bdfe1c867ab2f057393dff4cf
z5d8ff50323873815c32e7cefc01291b88cb5507084520564e3df3b02c630ff89f2261b86e824ba
zb4e5eaba56ed5cde179bbe3bc69cc322de6ea0aba08e24c2f1ea926948fa5e9215821bc8142ec2
z76508fe5ae8473ed26f7912b3b3074816bf47633f96d31bb5ef0e5fcd3c66558f114a92726189f
zbfc8fbe6613d2bf1124835dd3e54ae461eaafd3314170efddaa599be8996a54ea2ca7d233ced85
z2d73cb2815b2dc39f2b905e4dbc61f8849a0d295ee0f05d3a8d14dbb60e5c398e22b4b5779629e
zbffee945d68e80b9aaaba62cdb224ee22d458dfce5289f0543be428a9aaabd4854dbc69b048e5f
zfd2c9e44e83a1b7ebfa5a6dd33d46ce9c9ab40c551ff427af62593e905b1c040d5a51c7a4652f7
z4a6f8e4064da07861bded656eb53ba858dedfad65197a4660e20df7b6bf23b5f6ed13c8933d5ba
z3e7d326058addfe41d015923c2318e7bd0f07c38bf354f987f11848c4d325e732b04e6042487ae
zf6ebfb7c7fbfbbc1a5a8aecfb9d1040ae66c5bd5974a3e8a2afee4a8783d7406b44b9e1e07f241
zc4ed7fcfb59965b532104ac3b60342ff67b824fc470df22d0176df771bcefd5c505dffc54f3fd4
z801c3a462e5eeb0318f3fd380b7baaf004e5c5da10fa84818d3580eb568f505260b192d7de56cf
z5a7c06e6b9307578eafd3babccecf2c1525698680ae461936a72370c33a7de32845e41f1b9835a
z97fd7b35206758c17539939c70be4983a749c2d9afa9e990f792b1d8f1113d259635133acadc69
zfff5e1f4065f1f5c1a65d11aed8932e4b544b9a4ec949c977e3891e07a2245e35e0a1371e38a0f
zf31238b26dda4225776cba65d41b0afd37884baad30b9bf5f964833856fbd68cde6533d8b85dc0
z1f35c708515512e947b7d42ba4708d66f52f5af77d7cc5381c819842e13ae7155c24d68e7d1c62
zfe1d08ca0d969a0bf4707e325532d4ef6e01b41a62c60d24f9468cc688241faf6981517e904cbb
z18cf10fa2f1b1349c163bb5efc1c2602d06b1274aaa759ce6218636e949e868497dd54681786dc
z1a9b57f8c330c4bebfc8f2db63c84206e9d84ed1ab6d994cb8ad5e423fc97d8a2ec9fe6104dc22
z465556317eb090bf3192f2402065501fbc6bc38d57ee0c68db9c1f891068a9bba918513dc1534a
z8aed7880b52c21c86cbafedeb23ba0ad820276ce898d9d3d698211a361ceb6a6431fb4af855872
zadb04b9c7d7bb6780fbf8e76f0a1f810c769db6bb66d8e6f90cc4c738187ff48ea87e058dfa237
zbc0f57bd10c91034b71224b24c7182254029b9582253b49a584fbd5ed3be8b5bba6f5c8a2ac12e
z36925aaa031825847073a16dfeaa03714496a29f8e5747e11e5c93a8e83599f507f52d06bffd44
zef014fb2039a4b12c2f8aeff45e083778ce3dc21e31b76214c68a2b4aa4fc3a788749945c93f46
zff2ced127938ebba1de4bc6dccaf5741a89267160c5e50522557b9e792520d9a276386dd377073
za9d51dbbc3295d1cfc99cc4ab5452eca7fc022305f0dd9e5d6bcb00084ce895e4ea8eeb9e5badf
z71ce8301c292e008f8a248ef5d1aaad03180d219022a2ea97b90298d88a891ef04328ac59263ae
zc096041f58342133065407bd6f6957fc10baceb36da0c7d1302abdaff188876a578a26c8a7440f
z1aa142d8ac1f81df306db6633b87dc23cad3d8b171c6a49caa50c19b41bec0affd5c2285edb525
zade22caf36cad9bd5a09d1c0ed53e58ac63c8ba86f3180b01d3b2a81e6991d2dc89538d0f4afde
z8eaee96184b195830e203b4bd62dd1579c5a929682a38f2e2c68d18c6cbc74353f8e4e1f794c61
z66d3ecc128034c8f281bfe2dfc374fe7d4218a1e194d65cdbc35131e87cb269c1fb6a0a0a5c99b
z01ddd9ee33df2b550512bf45dba77a11cab717a131f6b5d02a8b22c44dba690df19d1d3fe6ad2b
z5a62a39cb3051580fae4bf5168f1d3c7610499b90bfb68148a09254aedb0079d8937927be33123
z5742802f4ae9c772e98d730e34fc0c144618a725cf19e3cba0eac2d17b9233e886f403439f1d4f
z61b6fdf666992bfc0000df28e92ed1c6e09dd3b021ead408d24bb4828152b40298ee13bf78ff73
zcafcb6dc3b22c95f3a642662f41c29d0fa660ef3768abde45956c76d88e6f006daff85667815e0
zc765aefe0372fd3674340503f563d11fabf47ad81178598a7b176b9cb177d70d3122a9cae922ea
z9856687d34c971bf90f77345e758f4b6dd00d050a31b5a2101898f3e81cd8300686c9f797c9dcb
z23779e47506dc4b08c340bf1b5eb5140e90e13cfb3913d546cab29e393232f48d9ebc2037bbe97
z11f4289a124d944c5df312a19fa058325df064d144f920331fd24803de11267c85095b1fbcdcea
z671fd1eaad47b0ceba3cc14023d22c3ad6c08f2c8379f54046a9d233afea55117531d8a8f942e2
z3bc0adbeb6bb7896abaca4fe27bcff3d73588567581b06c26c72d21cf2b35c92bd9d6b28f9f851
z84b6be3f91230152986f13d4529317259ab5c1491befb9fd0ef2240ae7d9221ef0a56a5c33bdee
zd5adf50eb12a41489166a4bf7403eda50bc710ae740f72e711b4dabf6345f53f0a6eabbe43b06e
zde873d45b4884f6fb019cba9071c3884324c0cd4f186c29b75208c814388f5c3f08ffc34ca86ae
zd50037ad78978869654bce282256cafc7d659d5155a32fff757e770357cb766a902195e29fd2ce
z418fcf8ba2df33cb32b0b78da98468501c956bca3989a67bf028977864ee611ab33eaf48050008
zbd36bfe5eab1486f282ab3a97f0f46ccffc515b421de734eda6328f9af94eba6ad5fd4f63741b7
z60b31953ed1770fb7ab470051e86022b0dd1341677a98cd24fc736a1d7f8b8e8784d2dfa82853f
z4e9039c8d22966ff4f251a504b282776483e87a7c11a77482e2a56ae790ef906d1adb781fd71e7
z1cdee9496bb468388864ee0380f78282e478ef009e59837896550b91f861b6df1f36c61c1056b8
z1ff792e89fedab6f1f487189907161421b209665b1cdbd8c56335c69596359d654f373e5907d2d
z574976d47d3aef01700b2b1665617c52495f462d46b8b9431c2618248f6602f0c38b3d68417069
z6aea110174a4e1a5a94247c15027f33337ac81ed711900a297eb056039a4e60bbd4b7f17417bf3
z7cf382cb7199e51d5bc4c01499c5029d98e08d04f65bcdbec246c97a873e8cf16220f27a8f0c7b
z959ab9107313796aeae30669fb254f3bfd95bc7e35b00a447812735d8502351bba1f4d912ab55d
z690a3bceb1fd1ba4b6aa4a499f3cbe04ade51a02a1e32ca361e9b229720577b16f55cdc2691b7f
z456e45a4e71a1d233ccdfbded6a4261207ea17a4f81ef0419a26ae907cf69298452836451b2f63
z557a97fffd43225482512083f5b87d1c65bd0c4a66a19ec9b9731c969523c6fccda6b315cd5120
za4cdff3edb48bc48c387c830eeb982c2995e489e7d87d6e59985b728fd4e7d396ddb51f63f6c28
zebb7a0c99659389c4a7724c24366ca476dd676b0e82d8cbf23b2d807928f89bb322130696e0d01
zc441975b6103552414fa29486d0d252f20bae6816374f962d00278bd990e3aaa6bdb1544699b38
zf4a6855978cf19010b0a394f5068e95b7d76db5ee8559f8bdf6cbf245762d90dd9952fce53d203
z7441512f7293779925caca54b9170af0463cc0173a4289dd87a72fb7bf8827772c865cd2ec728a
z49c3f2a27341c2cbcd7aa6cfa24d6a1da6451a450e372430564fe521b8b40d259766e1647c6d26
z5104d5ad393c6b85d00a2cb977f220f6e5f452e0c12d5b0dade5d945d1c73081073a0e6d1127cf
z29625943cdf5128701ea8c40a849179a66f5fc2790c80f7d0a1c7990717cb38d0aa05d5d3b08cb
z67a246e885f97f52926d33a2fa03a1ae99b860afc41864c619f3239e7fb8165836957e4fc4926a
zeb68ab71e6e51b6cdc056da0d2b115c2452bd70c009581ac90bdc3980c32dd7e2985e65c3c2c36
z0517a1963c22bfab87acd69486be5fba8cd630b7d9bc828cf5dcecf9335a83ceb8267f3119ca41
z808fd5f8210a539892fea17b4231b0558d2bac276f05275e4395814d2b6784a517c0699f5079a6
z55f898ac74884409869ca780f9062f382259c83b1cc07e332324e672731bafa70af92b5fd274c8
zf44968b062fb3abaf492c0c5ca9ebf05b3d9c05c68b2d0a2d0c4743b42769742e2386323c916da
zf34f90a457559cef13e3e9325b5ca685982e4bd7d3840c148d2abaf77f31e8ff96a9c66925ab4a
zce5e110245eec245b1fda84fb516ed7c3e1e89f9a983f4be07f4b26acdca1bfe96e74be37e06a8
zeed9734c05af828d1f98a94ec73f55e2ffa0c3c61e0b2affa205eb1a12a1fb225ff8d0aeb8ba50
zb881ccc2b94919b763f11c91279e1914b090b53355413024bf406a93cfcd3ea995e28cc3e940c6
z836c80fb403aa16e53c702e0d802c0b766f3c1f72d74d63690db89c48c23ca5bf578acab6b90a9
zd172eff9eb93820157bf039ffe4cbe113d1821370f2501ebbd4ff17548b9386f937e0f04b9ad0f
zebded42047c779b8638714e9e76a3dde4ca72e7b10a65886edfcf0a333ea6818a22c355d42ee90
z9259ef07e7394ceeb54c261d1a4ed6e7668782b18ca291ce59b0935eef670882ffb4bed405bad8
z08391dde0521e86c21dd6aaf639f6a5b485d1f9f60cf2291242a474f78a0ef70623673aa8c110c
z4d981119c9f7e3d1a5df2db1673f819ca98ed0ea397b8723e80f49657dd519f4141e4614230577
z10914ad6578812fd6048eedca3af4952a49ff6e0956f4fbd11f5f4d3d373bc6eb6749e2f8f497c
za901d27811d81667971e9805b118f137fb62433131146d108e6ca261921a0276baf7ba6faae1b7
zdd6c92c32d11fed8ac589338ab61da44f4dc803a58a86964a257a59e9863e779350689dbad60bc
zb20d308e6ceef301fa0f1aa65f6742ff282817f511b77064d602fc68fe3efb510c9ad41f9366a0
z3664d7eeba7896a82a1a83347f93f7d946747d0a4de5563184971138b499270cb6815d76c7f4bc
za96b6a412de7e9e13ac31cf6bc4038d24625192fce3ab37e8148c212d6769f5a20e4a720f1b259
ze311f91ae59cfad029437145d1da43c72afb4d5009d420bf9368d9c56972058dde2d7eb9462713
zd9a149227a8056e6de7b353b13b3f038728142cc777a1c7c39ebfb76b362889f64fdd32ce6ba7d
z6d32fcaa45d7058a58c037fdd3f0f1ed644e81a4de2e99c0d939dcc1a2bb292f3aa196cd87c259
zf5de48077ab4cbf3c3c9df08a4ff57b9cb6f9ef786b1a261e9093cfe8f13498dfc7fab0b48813d
zc3a6bb6c5de5034cb2ca122b366c9404802ecc7f71466db53af0ed521f05b929d33602dbc63358
zb3d6fdd6e2ebc816fd16364db262aaa262a719b08c29603d364dd1d07301c0fbff9a80353ac9df
z96c02227522329473cc2307ff0aca495ca945e7b1cbd081586c596fac90ab85d07036873e46ef0
zacdee01dc69e914a41d39c54594094c500152e43c0100c5c8fc1585ca9aa0d0874c18170ddc54f
z7552999727f2add18e185f4484024941b928fe2d302a0df6269a0edb69a8bacccfa91af08e1572
z5d4059c8ce6cd64c71205c2ea13ac8e4a112554fc93c776f32f8c8ac4a65745baf059f1e58ae56
zdd3c24002315bb3224cce44caea7de7178da6139ca1e989be8edf29aea1320d3493e36b2a797a1
z2ec0bb96f7517638ddb105b726e213bc6a0d9e0d487539ece6177e21a45ac4417ca23faa6a5840
z93a077498c52366c3b8ded4c3839c93a43caafc033c88f8612c70261abf5e685e8d95a39ca3bd9
z69c67242a36db7c59e823f9b46ce9e2eee6067d32c9b7bf3a955770aa7730bd496050c84ef60e3
z4f7cb2cd80a675b07a936eff4af2c45e511ef64602c969c28bb393b32f46f45be8ca00282d8474
z45b0caace70f17f72f4c087e2829744de86e5789da83880eae208da0a0b9f8c6c2c90005163c84
za3a5907ffd83d501f778e09b0804cedb4bbd4d24248e6afe8e1d699c12483c876e5147545ee00c
ze2ca6cf5d10abe8deda161624920c24157a235399fe648dc67b2563adef21f245b53c82a84fb77
z502561bcf35de25c86947c9cbe8752fb0f30bfb3c01fa59b7d6736d388ac489a1a2f63c26bf706
ze1b02c2100bf6bce6c33ea60b1f423451dad16cf713bb576fa84d95317e0799037329d7050a524
zd86c276abb58c0b4da78f991c9b77c4e4ea6c78843ff7fec11eb73cd743ed9adb91d1fda428c4b
z677aa325f27eab92e46e768da19f38e1e6ea6cff611b9b3186bcc46dcf0596f4adb6860483f49b
zdabe47d9184ae85f6099a776cd4530319645e44fe73e473f86241567b099bfdb9ffb8b1097a0d6
z85ea57434694322a7875d17941c466ef9eba4aecdb7e2ef6746b4559314e588494aa9f0a97a6be
z6dfea36d3aa74195c028aaf2ab2f645e603bf9ca6cced23b6b99fdef89bd96200a9a924605f04f
zaf046d4adc202ea52ea612ef92c3ce38b5483280c1deb0960209d97f5976f04bafba2b36bb894e
ze019fc872d7eb9a6c95187e11de2bb59b9c4bb3e006e4761f47a41d68df9a274b01583f92d27c3
z5da2c7f67929d00347e278f157fb8275b114e2f56419dc94e449f3d3eca19cb2279a39bfe95ac7
z6b8a250dc14ce125302925a269994353f33e9323f430b5af7c9c892dc632fa470dc63b08f40d36
zecb6996fa76e621a02185e6d673ee63f94ad3542c6916d5041a93b5486d434fdbb7c612d1d5574
zee24472f0da689b7cb42d12f258be5d6b737ac393ab97cfb6239ede854335e789242538a12aa7b
z5349d12b88dc7271c44e7b0bc8296acc51f5f8d432ba327f4be5fbe4bdfa9a7ae81670263265af
z081c49294803861a9ef7c913765b18e204f600bfc9ae7544f586fd1e24f2037df29cb56574fc13
za4613fdbf3aff5135d9059c49b437269cf33c1c088dffa178e7b0151264faabac00cdf61461def
za37ed048c4a338be1bd1f42a87224ff9e9211ac099b63196318cf201c20b4e52a1aee2db40acf1
z5984b514f736a398f700aa8fe79de37f3aa4b68b884d094a2004a70bb3334dde635aef83edb008
z3152446d50237faeaab41d7e87a55c9c96a0b44819884f627a001480d86b1c79f81a1b99d47385
ze78d6af750b40c9ed6bae39b658e35285483cfcc1af446bd3fecb9710b9216733ca4fcf3455a5a
z4572a0a8ffee164592522fcc5c406c066629e332dacb85a79cc1f49373aa3f6a691e71a76ef647
z18c9b592b01b4ed16dcfe3413a1ec2f6e5ce2ecce80c3235242803eb87fc6d2859c18e75cfe015
z8c860d891ceccb2b0c59a9a71e998c10ca0962d474fe7f57bf3ad1f2a1d0959f5cedc7dea46818
z61ba062dc4eaf9cdb722768744be00552d7a504c846152eec654ee25a3317d6b0cc357ab8bdac4
z046f463efa155eb7e70390600785c550318932305d87a7182e07a24bc8201d64e05df6d03dca96
z492333f7808509867f7d4b82c640adee69e2f65a34c7048033e0efbdcc00013e539200ae015f1d
z7dbc7c8fe0092b1cd9b653760797d5f3711d62c157d49d38d6233820d5620c1c01c78c70641a1f
za8dbbd8b267541b1ff1a27b7b3ae38e75f35180b26dd345b4530d3320c7d59bd37412f3faf9dde
z9cf5ac4407a7af341223aed365fb1cd27fe2610b3ebb331765dd3c6b5c96833ca53a3c2780f691
z75025a461bae0c58c1a879cf338281e808b6bd89515346cb436bcb48c89e2201f161b5f821d0f4
z6e717e531d83f24f8759c6be169df75b429f974b19baad5f46ea948409453cd9b6902ec881916b
z23a670216df0c338d87f55474ec7dca23ceda25c276ab70d4051de7bea0cfe1e33fd16e54f3e7b
z37a527faf00c23fc0480e633f0ae797c9974a3a11ab8493ab1be52acdf307652c63f7a3a2bb38e
ze726e6d467cf869683162d7e31632c5aeeb21bf43fff7bd8448278b6c570a23e867cf1333f5820
zf0fea4fbb969302096d17afa66522e486d7924b248f0c2fe0c588ebd40a69da0c24dbd6253f212
zc70b8eeb42b538e51035ba815fab4ac92654cea908731541b724176a2aeead2e36100293e934de
zc49b948051fe338ad54488b946ac25bcf25da128618164fccf84bd9f7cf737c3945ab840efaef3
za879b3e2bd7f7bfa5a09fa8b4cd275573447c8cae515608ecc131d3a9518c3d736502c421bdc33
z0e34cf33f3c1a5d0fda8d750fbe038b2abb37e446c94ff25394ab373b2a3d6c271d9fe85a1b302
za1dce9900eccd2317d70be450480fe393360dcc078cfd7bfc3d56c2e4d4eaf1fdb4d05dc028b6e
z2911e13895b7be97a1023dbff16bf560332ba2c1a07b70be57aed1679745556840af97dd6d367c
z44f7789f03792ae3bacd83f174c4d5514bc0add0d467b36ebe28fddba2d44dcfbb26acd5b54482
zf58ebf4c3bfb387d2c2c0e953efae348c0f650a5207ab6c611170db741b33574bc6c418c4416b8
zff742398e09364047181ca51dd9041838d1bf0d5e95012876e49a1094d44fb1168fc056d8e087e
zbc55d55b266ed8c92af5cca868cc3a291d13980599de8a4388637961c73b2078c72d3e37fd9bda
z7a8da0a6d015556d85c80b8da8e6906b9d32d3c0b19e2dbacf920cd6fb0dcff6d071ac413cf820
za4ca90243ec607c7db12910739933d0e35c90a3d0a211cfc0f9b094e4a3e511e03972ff3fd405a
z58804af62c920cfccd93e37665e43fa7eef1e7f34a79ecfa60b4d46b33b6d7009719d4798a970c
zedba723f771dc7656a10c3c91cfa2a85dd57535d42cf7bae8f5cea25172adaaf5280edfa00717c
z600bc4245ecfaab12d0409ff765368b57cbe17859bd1225633106009859c20b81a5508d6aa174d
zf62106737b165d704567f83bef83cf407319aae1ce0261e19dd305b22c19ecad9437f72af3faa5
z8f6a60818fdd36d111ed986f31802cc1ca8880268e47490da30556dc4fa0e4ccb0a01fda45d7ab
z750092d23ed05c12c26291305290e77c65a2b9fe31f183ccbd837417537f5df530e0e049dfea97
za8f38adde0be72108525c70322de96c791428bbdc25d9b971e9c6fbb1621d927c72f4c96abfa73
za4cf45d4b0c315f7672b6fb80d3aa9f52400d4fafd08dec2b7f30a7a4270fcdeebca4e791fb4c5
z4690b67aded7ab8935af644091d0ec360ae1e6bb11d8c4d66078f43ff0d41bd3d30a6fa3157ba5
za9cb5af7692022dd250d360ea2a7e89549272334abbe01543db8ffd568f532d8203153df45966e
zc81e91c07e6cb2c8a7c2c49654d8778e60d1259162de7ef90b6e647c762bf6e0c0d4722594cbeb
z58f06a2dffaa25da89bd15dfbdb868a33878040b7517eca565d41b4ceff4216e941474f551ba17
za35daa98f75800f8d434acbe1daf30e409153b5f9f7082b32fccc3a1598f173783984273af5bb8
z733c5d05ea0ca48c364d387d024c81746414b095dae425bc5c249088b3ab5770dcf6ae60ebce1b
z10eea24dd34b29fcd538dd49219a8ba892a6b4353fae9d89f1b9f5b6338d9113aa6aa6f37b7b5f
z73968ea8e67014cc1e5b5bf0d9aaad78ca7267585a04f8e9d26bc0fd7c49cc6bdf54a2125a7029
zd73478e14d37a9f4bf4ace018d63f528e190feb9e4afaefbb2caa278dbebe083a01a6805822c58
z1e2147b71391be963f93f93508f37e5ac0645e212706d662dc2ececd7d8f991d949e539499f556
z51e76c0ca51b9dd0ce7f4e5e5b974edad499b67235bdde9580a83aa156bd1e46b6f97eee3309b3
zc6a5b360b002c9690c7a23a081b3f6fb976576de43f70c928ee72d667b1772ab7182fbffc1a1f8
z014bba0274ae4a537d15a9d543a5783b60afad4b9879249631e7634141c8c8cdb8ce816917fc4d
z421db2f2813422b2b3a4f57c5f91b500267d0e39e3a0b0c4f9fb69dd761b20ab172ac314dd1b29
zb335703c95f49a045be2622ebcf760b7ca2e0f2c30480b1fbde72ec3dca4a7a3331507e42020ee
zf5ca5ecb0897d52f3686767859792d90c58657326bd65ebef0f88ddde867ebec4dcca54bb66336
z0c516bcbecd2be3a523cc9b9202871a6661af94c031fd3f6371c1cb91e81021b0d5a6b3371e5d7
zb3864f916a58674cf5fdb845d3223cf6284972752483205f02c6f7bcad257952574f4c107309b6
zc7a7da5eb2d8031d1bd716fcefed436bf7688fdb9134f172b4764108f150b0b5236a4e3ac6b013
z180528cd5711ddf75364bb63ed5ab451361b704596596c92657b69fb6aa11d0625e989cdffebdd
z2f08dda67b1bee86b2d2cd3ec638ef66f09b439e2b3871a6385ae3bf45e98dede9be7e3d0491c5
zf5a6a0ad54f7046cabca80bbbee57337de49102cd4a66ecdd79d5549c256bc6deab693fbd98290
z66d462812fb2c0c542f02465b0f8cd3f50457216a9fe23e4e95644fc92e3dcf642d0e089ee35c8
z4f0ec931ca772da7e8b8933eb48b87ec094bd33ed712c894036b35a93f74bbf827c641b9ebe25a
z9179e1c983368620a3e3f745be763d3bbd1f4262c2ef6d5f40a85be27375bce2ee6d11895e345f
zc6bcb82be6043e43ef30a2ed5329ce2f579a177b4c113ebd15796a7f701f62fa19f2c1c9138cd9
z91258fd0fc581615442a4cbca31e4e6fa380ebc317e73a68e792b26cda80fd2660ee3e5fb83d7f
z534432d96cda089a664536ba7bab30f631d7947638e9b958c3d44aad20f1e0158f0211e521acb7
z68b7ca2bd8b8a07d5767c7439a70e85002000d92866c6becf82e7699e307eb8fd9a91292404c34
z91afcb490794811bf66f4185ccd29c0792aabdf87d740e15e3fc89cd758fca6cfadc4805e3a264
z61497cb5b875273c7438f6b3a8fd7017b8ddf157cd249ed9cf31bcb0db17cd219068cd9ca0cc1f
z25bd16ba4718da9ff20a0e5e712b89fc3c7359813f2885a32e6c4ed84ad75bd4b8bed636b29440
zd3c1c71baaf3507017be213a3bc19cf586fe15ca7c35ef565f34dd62a5307c30062882a3272f05
z388bd9799f56ce56b3bc781ae6c4a638e36df54912d2eec65ce8e59dcb15e1b1c03cc3ed30dfd7
z0929128809fc063358e00f91c87e98bb04103f24b02f90240d617795e5bf818bb8551a41feda34
z953a1808eefa56b32a94590d7e5d0ba3b1ca5048043a5c4267a19ac4ff6270431c5f4cc93d1d59
z0a66b428ebef04a4d79b269f5a76d17b857ea87bbeab96984591c839ed381afbf99f3ca445d55f
z7c5b70ac1aaa130209d4e05f70d1bcaced834fc71cd53a329a586e08c106507faec177316e12d0
z9b86e4c9af42461cdbe6260d6f4357d3f45d23a86ccb9c9ea12daaad3a0a0cb3a5babf8a28e23c
z3b9723c51c5127f1369b2fe3c51168e67cdc555972d50e9b3dc1f4941b7aa91da8f74df3a6cc0c
z8059e546ab2799a710057edebca2a6f50a69ce4f31f75f719f28ca0fd9a387a7224f5eab3d5fbb
z3b84e810f25bb01cc2ddcf8409b74ceced1347d954c6d38bdf0863d97151c2ec5320a8b2def3f5
z76f6ad7ab11e5acfb67402ca71b9315725671cb54f79337c6a1a937e17247dbd17c9a52a0fa041
zba8ef977c16aef62308cdf256de0afe8cdae2e13f7d3562ff9167b8e252fc3048883cbd026de59
z94eeb0746035a7905e3b38ccfcf51ae2d8f6c1752e6a417b8cb253947fe891d357a879881701d6
zfb0ae51fdb93e991cb50aa27e9396b02d11ccd27f450bb401575bfd689997ad81b2acb9e424aed
z76bae24d10b6117c6df19a4c76e0b085e10118c634ceb26f895e9aa69fa42bd4f7d9484d220808
z149f40b21dfee752a706b356b1c899059f524dabc61568810444a058ad75022cdfbf5cf56553ed
z10ad33e89e00e3b8876d5741768d0471f9b3971b3638624b70a4d2fbfdaff86f6f63809a57d6e2
z8431f287dcf0820cffc925159cc3fedb589f61ae8c76326b6102b5e74dd37ca7bbc587c4035ea4
z4018187378074a4466ae75d1b455f5597d5e24e01d4e320c5b16863644b757ba9316f3f98941b5
z071d432fcc38f0e7b44a557470d4b48af41e86c45f728cb3e2a22bdb65619ae5c1b1b15e0bc6bb
z8689e842c68349f43f3bca4c240e10db058a8d95f9db8ea0532df7f9bc765c05c560e60c8d9f4c
z1234980d3ca24f9f8bbe033498747fc44aac2db32dd03533066f8d13bf4f8acc80af3f3f61c9de
zac66ce022949419f39339d1eb0b933367227cc1e19c51803bcf1b37813711dbddd9b81fe200f2a
zd0bcd685c3e66f5575bead569223e2f9303d31c1c9423f2fc82d50085e0b22857fa61ae9dc4a46
z63186e0f69a9b47f5ca6a39fa31a7d2eaaf5bd63e0c92205781491222edf148afeb09436bd0131
z5e69d0929427246518bd830a8990eda9a39582f56e4029493ebd1d329eca6b46fe8f19495c8fea
z2193316a049d3299c9fe24ace48907800cf8a7d5696c5a87ccee5c9f9263d5a8d45193998f0ce6
z51831331f4f5ac98010059b9d4e014154b7e9d40d26e876a0253b22673e8dfb2911d85b4c1f3bd
z37f29593a729c53d0301c87496b37ea9d93e271512b9c4c98990cfd092e1b76ca63ea877edfbb5
z113ddc885c0a45680677ac4b89ef3bce22d1aa230236cf66660282a2cd26f9906f7f3feebc9d98
zc226fba6ee340fba1930e254cff1b5392837eacdaa4725545565f72cb489c33c13bc325003ca28
z27c88c48d188528dd513fa30bb49a08df7294995118f979a92a7adb286475b87540c2cb65cf75a
z858177f5bece7a9fceef68a7317f2116339e093963856ea7cdd814a14a107c775b04808433e987
zc9c254ff52f7aee7491fc7b68abd8869ea3359b6c5bf4f42f0c8f9b901c7108e9d7a7a2ba8e9c2
z091c8596447b3be0909881c1aa93b85401c22716dbc6646f176f5e928c4cb6b8e21eb44c43e763
z13180abea146462b8e4e494a687debea59fbe4e9a0f48f6621b75f251e3962ac55135f34d78367
z384dc79f03a143115b7767432b99900182615b8a3f5ef77df87589b518800bee07129ddda93a4d
z9c98774958b79e27aecadc6c9c7deee3bea4d28f132442a01e91804a3a08386ec68cceab21b308
z1e96aac08d8060066347ce3b175bb659da907cfd9fc2daff4decf599c16f03d91e7ed0c27ec0fb
zc01f6b96aefa120c86581ebfb96c78a779663e872ac7b8d973440a826e6a198a907e512dfbb52d
zd00bb974a8a069448e068de55568893effd094169a3cde349a07806f23ebb92c33aeca80afdd79
z9feaa42d755d632a7aba701bf48a9a414b7f47f0abe3a3eaf1e5e5037774bcd6b8b08883a6ad75
zefdc3f8d50703b34c0b57e555297ff0d8de25917e5405634cb1f5bcbc6061209f4bd77903a30ca
z66d9b3b4ffab6296023264bb6ab022367303746793203948cb5b7ece7fde7e8701c262ccbc79ce
z6ac6774cd69cb603731ef8f7613f35ab7e2df0fae0c53a12cea24206f0d75df9a76408c022e916
zeb1aa39ccfff80d40601b889e5dfe1ce995d058336977e17a5d9c0c82c6124c9df1c0b6f2d053c
z4579dee4f8801cf277c77aa1f341bb76e717680214fc4b2aa89d0edc3932c4bade7630dcd1a2ff
zfd1d657521e6cc2d8f0c66f3c7e0e772192f461da745ac913ca8515244a9440a7302623e681078
z773caffe5899b45bd9c11952d9dd64975778d2f9bf1d83401339f29b10880b7ec07d3c355beba5
z939d1fba5900493c29e7d68b70ac11dc38ab87010aeab4b657eef2823aa07038808ce6f109445f
zfa7613ee564d9c1f9a2e94df2169975c06eaf5ece175e404623717945f6593a25a7e3a40002ee4
z5298fe38b2bad6f930c681b37303a3105d895e26b410a098c293b618eee93d94e269e5ac5a5cea
zde95e2393c6573ed718313213a0eda25c1a6d6046ca49cb7a01031f991d4f28e8e4c363ed9873b
zbdea396ae296ea57c72f38582696791e97dd0876ac861d2ec60eeedbbabe1a914443593c81ea4c
za74577403d778a12dad7028883dba0c12b411208337f1bdb76724cc53f88921f815414d340cdb2
z03ec5486aa087e55985e04dcb461e6fefb73d847bdaba7caae52c82cdec4653a5fc30ecd2c5051
zad09adc9447576696f6894fcad43f9d80db4ab70e5e685618077ca3385c9e04a47cde0b7602a4f
zbb12102cf799bcfc1a06115ecf2e895b0c583fe19663c3e81bbaf78f11d922e8ffa0532b872961
ze0d4946b69bb2686924b6ab3200aa315e2463485b8c462eff13b6a37dcaaa941068cabaa3bf897
z11693114d5af4bc7f00074497c2d43e7423ec9162e35896b8587f58215a9cd97327bee96bfae61
z8f81743197555d05082ac930759852b1cffe729e7c3b7f7624dbdbbf43096e41f1009a2779e548
z2ca522a8b9e5baee134f76aa488312b39e4677d2d8aeab0e702001422f6c7233d2656c8f41139d
z53f82c8275676eb56a5f9a6d04b7e6432e0f34d69a7fc0eff116b486b8fa40a80402664b1612ee
z221a6db30c82ff24c8c7029a0ab5cd1846170f1e27953da35b8321e0bd50884bdce241924b4a28
z50f0cf0040dd7619ce20635eb01750a6ca415bd6c8abd7a896a7022a36c46902dee0290a80cf1b
zd2787e23483d3bd08cfc01b6cee93619b05673ba0c0c4b61271a61d6b6b744caa23acaefab994a
z253087df96db4d8a86be66b88b348a5a3bfbc40dae81d15eef1bf0645bef13b21210bc23c18f22
zb26f3097b778f4fba4c5107ce37c68f16528d8fc439d2a77c2671e50bea228ff2c6aa358a21b39
z14b831c8c015218268c46201335a04b20232a4c77ea1e1ac72a1913186a96bf0883559c6e26d52
ze8242d95e93a304d500b58182eefcf165d88bddcf47f0e3c5a4149bcd9b02c1ac02355471a8181
zb2a49b65addf7e30e17f3920f4b0892ef196ca5c11d996290d54d70b722eaded241899f3e09d15
z9f8707ce1536ba759fdc44549c7fc674ba0f10b51c6e29936d9bfedebad4c4e3838cade4e08c3d
zceeb040f8557cc91cee253ff7aeff2721e9fe2b1ae9a495ffdc2ae19fdb01fd4d787cc2311c5d8
z2a78737293f640c022f4e30afddc51e376203e61f62a93ecab88d955024ff3dd1680d921ea1bdf
z8cb22af2e738aa1a835bc91330d48372d18710f7a86e7b46223345e1d53efac0ae22d0ddcfa858
zc7e3ab91560eca534f454f033881be4d30c3a7cf5202bb1cbde6036e5ddff483b1dbf4c287aa6c
z1de6dfc367fe9d9f0b9ee164733d5ebf3a6feb1a698a2dae3e6612ab7dae485c7b1069c3824dc1
zd5670d77e3c562971376aabe90a3a4158fe90346e78a174b48c856a4cf9d2a6688318c7c6af744
zc7522f63c74832923eed5ca50a8f6515312d3f1fba6c54421cad973091ec287b547af9256cb163
z048fa99fcb362851be1799e1c439aa9b4a39fc1f9ad8a50361f9b30789859bff89c5bcb1c287d5
z1dd6c8813311c0917180efb282d5fa747e7e17d36582c82a2041a9f47df4225ed587a99bd0a9c6
z2250b3c881ce1a266c42022e5addab305bca30923a75334008a17513eba5aeb0355507adb00fb0
z2ebf98a5e719c4f94696388435d3847ad2856b85b024110e62109ce43e48867e49a98ae32dfc5f
z6e09013c07de576b6d7093de718fe87228dd3241a6667d4d96155275642cd073fc8f021332b035
z470867958ebf7744692dedaec778dfc8a236c22e99febf557293aec0b65ccd25ba0331a8b4e9fd
z8cdfae97c05fa2e85975139cd3bc9a6937c861c1aa916373a6bbdbdbbaf0d0aa5c1b7766880275
z5cc34b35f7afe767b112fd4324eb97be5ad4fed0588d2f35a4af1a20d6563db4e78213070a2514
z1e2ae11802348d379323e878aa84bc2aa608ba8c8e69c8703776cd39104cae5506e68edc9aea85
za39667851b0c9a7ccef46a3515140df13b31bfef564a137dd66aa85982918ae675634f19e74ecd
zceda57f75eaf424ad5756a336ae891375ec380bd4ff921cff4db6c5889de6b986a31301a06de64
z25e0ae6cc7754dd5e4170e80248164f9beb6fb030e637ccb01353e1ed5637a87ffa85ebc7856e1
z80fccef211166b339622718630919b201f3568303d6d8b236f5c81d1b89d7471b21b41363ad74f
z4f86bbadf1ec3d7e89171acfbd3853913205fcefab50e22906cde094d10072712c095d5b612dc6
z3840ac143224cd5f43439324e9d6f8891ca5382f47c136bc3aae382aa9bbdcfd068cb7d9813b01
zf4c898534c7d5f1df294ab487343804c2068d01e0bd343ce590ddf19fbe97650f3422a558ab9da
z954787f16312ad185e6d73eabddb722ad71b8713772e0ee4475994a1f80668a1b86cb9a2893fa5
zaf65f629a5a86e41ae31170233c45cf701823b24d231981890b611214aff79ff1e8278c1f68a76
zdc5e0cab1031c1265f16e9fd18f67c65e58046967d92c817ed47804e462dd14aab72ff6ec997fa
z69d75e082c37beb43b1bbe0b0e91068a644089d84362436ace61ace839eb765209cca7ac0b5f96
zdd31ac206134e5cf39fdd1eecd549df22242674e8e6c93ce962d9e47006f34cc02cdcd19a5a85c
zfba28aa8110eaea4862b2a9c0ad766e532df035fe52ddc5d5c6ac764f9a5f877c8305586c632d6
zc00e61eef5cdcccde4f0f0aa3db8323334cb48c61b5e0d99b4de78d8bca62f325a5c80b765cdb2
z28013b5a5f7528257a13dd948572cdf4fbb3fe4d00c8da88ed545da74a2b6708607ce29791a670
za3bc635bf4df39b478ae9f48675f427ab61e6df76829d471385f2ce7f86cbebf19fe51813db517
z471c58cdc37925c1bf22c6d6bb8a476fbab0bf1aaad768024c13c279ced44cb81d891baa3a82fd
z0c766ce564e6162da531b431a4d702f9013e22e4e7afd560382221ea49829460de2f0e5128f3e0
z91ad295577a4e71e168080f7df019678a5571ac45c87db45a1fdeb9504d36719ed6a8b6c768d1d
z0a0a9836548bccb6b8546f1ea19b7053551d9e234726cb952d2b645088c1c7124fed6b06599409
z763db4411af8eb345c24d975e723f8d303f4b6d31f863b00d7a712839544eb0fbdb81f113c6b71
z6bd645fb36c6c029e96582e2650437622dc9bc618d143a1df5dde53f0104ffa87474b284ca9442
z1df46c18426fb680b749f96c0d3b9a894d6c7d812aa96ab1d24174dada1e8a1ab5ca9e3765003a
zc29f7a594a8af64a7ff226f4b1167ed218f5fe4deb7fbe8e0ccd2cf11761399c2b21069e49fd28
ze3267f71716543d65376b1ce6edc16d92b28078e6c15238a6a7a948c74801bbe53e1750a49477a
z3aa68e1b95ad93ca882875b959cc145edcc232d8b91347f92dd1fc036931ac910fd9e64c01e00a
z40f76191974fafcaf99050fc8873e782c9a4af0c65476c9df5db34f4a6e688ebb5905ee5a04f77
z6b55c13862e6576650d349a3d47cff10db68b41b9cca39627413c740fbcd8d9b507d91890a82b1
z4d00ec1c43926438bb2dcd539326cf39cb3ad658918c96cf1af1ae7f0cfb5762db78d191e5e70d
zf13b6f6989bd467883ff8a832307181bc2683f598ce66b71a0ec95dad6aa679600a19f5dcc0a14
ze26f156b4e8792e559f648be5a39b6525e87561b13b62e9d3fa7cc1cac77b5ca3fb54d73793eed
zaf4c0fd0ea24b940321a847153ad35c4af4fc4dec101a3006914b0f3a340071ce7bcb01026ebfd
zebec051312e12d590212685754bb6dd973aa53d3b1ed6e78ac4baf2568cf7c31ebea03a8006db5
z037a2eaee29ff9c9612ca1abce2f9ea7516e550d0deee1322e1e86fe6aa1a6c8fc1b22c6ddbad1
za759aa37576f4726db49dd8654bc4a398b3b0ea854c62c1a33c16036b3620c6bf17e0e64b50d99
z3a14a290c8b74a887af1d75a8f535770fc565863118da1792cbc8c4675c0dba83e90757aaca13d
zb82739863b4a8c644ddf0500b361aab901c0e967ebbb34e522a3daeea84ee147738b69f5595074
zb9e35c923e746172fcfbd8d6a46841dbe5ebc7f3438bee6f7dd65eaa25f0186b6fa9ce25d98e81
z1d8d823acdc34190ffb2108c3666269686ddca1b26ba59375eb2b46cb2cd4b1340e0f579deeed2
z69cfde8eabc56b1a22de4d09d89cae3a0870dd83b6d1126984275b2a154d24fdc7caac3a5a7666
z488d41b6f18adc33ea7f11bf2ae26d8d9f083e5d96c49ebe8d56615dca93f1db15247f86f4cfa2
z4ba16f99b4399ad03379383c22df91c842931e4751460dfc4442557ec3b3e76f5857329423bd3c
z8a96a1159952eeee54672e382ca395869ff3f70c537115dc1ec393866cecf903acca25cf0d19bb
z2a40890bbd03360f930a3a9242d71e71359aba3b85c0568fc42b6c8be185527fd9add8c51006af
zc8a1426b547c52bb1ea2d453211472ed546b468f61eb147d380429b63e1f990f45637b757f15aa
zf0c812b2a0eec5c904a5d27d169e68caaeaa74f4269dcdd5afa54d187f1a610ddfba7df840fce9
zfb8e74242526e16a6c7c3301e72c62ef5d7bd945f5a10e098465d4462778b61767d5886e4b4801
zfa588df040b8fc3a01f07fa48fcf4e9c7711b4e16bf7c29efb5d327f3f79e383961d02418c64ec
z496c1adc58e2d81edff323c207fc07cc6c0ccb6167d4625e32e044f7a3da2f15d0d30bfa5254b5
zccaecd043d7e1118b605fb67ae4171b42c2f7a07c4bb86e75605415cee97080494206a2ac8f4b3
z6d446c40b1db76ff23f684c7c42943786ebdfe4e85e0f7377115eec83a06c4100951e8e16b8172
z966d230f64d93328086e1abfa4d4f3e8fbdcf4560bdaeb8b8dd83b516e0cdcb997a8bd1c4763b4
zf2a69cd2088de7c502a440b1c026d94adcdaf94542cd58192e49b265e0b395151d36bf7956bb44
zce8a44c080f422e7c4c4f3eb348db6f3e4d2d1a40b58de9942b3d1c7c2658f9c057d291a536f4e
z743e7b0470488ca269e399caf0b35209e0122851a49488c45ecde85d30d5f444026a5eebffdc11
zb33feba4fac0124a5e06e23b302af2111ef0076167ed9294ab7be0e0c86de1671c469518f78c69
z6efc389d3e7055d3807fde1faff97ff22ca255e7e1d2a8a4e36bebdcff8e579791b4bbb98b142e
z4f8ab39917cabbff495e08b6f013b1cea7dbdfdd887e121939eb9eb4e739fb7bb4933f65774dc2
zb07ec47c1140de9415f179a004288285579f491f567845e8142eb42abc1b12e2d5798848198449
z470149436c29896b2380882a3c52a66d195b43ce49a593f91670332513b8feffab81d10327fad0
zefff1e44183cd2bd12cb619e119d59d5327f416de6efe7501e92a0762765864ab7f2de03482484
z44170bb313d161dc98387a9e44f74c72f8e4713a155fc43daeed59a128bc1a0bae0ecbe849a1a9
za4316286afde70d265fd0a14b3d9fd531e70c75db7b12f854aa9c8a2a6734ef1c509f48458555d
zeaebda2b33814d0dd157695e613f6e6505f7830706e897effb9bf288385640d71ec15c27123344
z27fcbe2d7b29aa05f89067cef683a234145efe71388ccfea98ef22a59bd979ac00eb7b7c128a54
z72fba0722dfb1ad1b775f3994f6d3e2f576dee5ff684e186d923dc534d93fb43aea0c6d9d3a655
zc70e20935deb35bba1f818fa10823249a95ec4dcdbcde90dced2bae3d5c6ee83a2f82fb837f85a
zfb57a6efd67984c2ee53fdf245264dd3bb0a03283c1389ea5409946eda78ac5e3940d5a6cb4f55
z344f1567c72c13ebb7778ed57ed934bef501fcbc0333d5311c40d9df3764a75dd88e5e002d8ad6
zc8f4146fd75b0a6c905a32c654c5866a12ce99d26838cba99c8e0facb00133635b18ac33cf20c4
z77c2f3a71e0a8bac8357efb94a4cdf5e5c712e511f97b904bf8872ba5c9de0af935f585597461d
z19dca41b84013633d39786912c339d3629ba1d0a0513c8d0b3df2fa4ff0361c68944caa1bc22af
z96fbd7547076d9c1e3e1812bc0b5fee8a402a6a11bbc909b515b0eb120633affa5a327cc116b2c
z9e6ceb61bed2d02154eb1bf748d57229a2c906f400b9059d7dcba818b25a4170fc8f13fdf1dfa4
z97949859ceb9971c30ae17a29de8ab3fe510f553cf38b1720e02c135f040e08d577194bcfac4e7
zdf4df03f444af1d3441d90a27ef092334dcb8f9180f51eb8ccfd8ffe4e209d083c3b2075dcd7f8
z2247625f0e24936dbe07d7f498f802e0a5c6e774f73ef094d27f5ab96257ec5a58d7080f5a552f
zc934be484da3a6a7c0c29c724e0a4f54ce25ce0bfc37645fa8b71bb4e571c3db58884950749c23
z1c627938c1bfa4a28427964fcdb9e793886f142aca7e005270b90384ee58fafe61b33c2c1c1d9b
zff4c3f58b682df1fc16c0645b6dd2df5e5afda5c2c6f2c63455f7cef794032067dc47c0db6a715
zb0c5ba41d255ad72782269a5b5672f2d3d97f7a9d9f7e017a705552547b537894c7a92b88e437d
z5697e627c4698b1d13636c214aa8f6bf6821f919e1d4ce426a86f4c8753508cd5665898975b5f7
z54505a99926a738f8d6d5b6dc8314619962353c6fd6e9976025f4428b3560f27f65e5f2288cf02
z09393238cc5fc1e1e87556220fd9c94212c6b84c7a46d13a008c88c32e4068a4ebaff0812d1ec8
z09c1ecc87b58f9e14954dbe2d137453399221861443465383e983de7018473b4d17fa53d073d90
z64e562cf3985fb206626a8298c8068082d3635fd47c3eaf5a5fd1f07769fccaabe960f1453529a
z1a29204122edf92c44102fcb6d1a3342dcf39c2809dbe8d2593414110f4881ecf14c81216d4c44
z3f789cb7c5317dfd882825021f644e69637a90890e7bd99072b0f63814d71b8976c555901b7fcd
zdf585673bd178efd86a56b89321d88c8c3a47bb4cf45bfe19be9fdde8bd0e8d1f70f7088643a01
z2a12ae007bf4bce07f6bb8878d961ebfaca43f6fcdca7df1e01531f1ba04cdc4a41688adac38f7
z7b76d0637f29585c5c815ec4aabd5ce68e0b4492dadf7bc12dd1ae8c8958b0f31f375747ac4224
zb181b114a1778650f2fbc41666c7956fed885dab11dad61270756687565958881962cb347f1225
z38aef204745bc50a8203b2ef015d74cb7aa08bf3131eac38362a10d1231a0ab22d11a7932fbeb9
z932f39ebf6e1e5f51313030d10a83a961192d35ba920eed3e18faf510c93417450b03511893c46
z32dfb021b4dd55dfcd17cab1a0713a54037150a6da38bd572589207c88bf6ca34602c9ee5cddee
z186a304027587fc5591d29cac42e356f1ceb1b5042d31c208bebe24412aa10906b967d3b98e80f
zd7e92f93405c9d3112b60df1388beedda42b06a1d43570c79a2827957d6876090eb78be42c7e70
z92030c6f696086b582cbec8828c315246e5e838969478f2da0465bdac2b9b4f8f347d560aac6cb
zc5280d3d7de837e9a979728be464c2c7605527d04e3c56ec4fc8d9b093fccd8eaea1632fc3fd00
z2084ba2c73510cfac2f4a58ae13c446e2f0ae7c2bc923b95b8316a50195fd98a19182ac59190cc
zae9f0dd3ab3939737d2cdae003d15c9ef32951d8309a10bc59ea682077d2f0abcdc0bf0858848b
z6d30aa40effb9614a7162fdf016ae2ab9ffbb31acbe734cef57c738257087109a4240c54fd9a46
ze40af33211fc2aab66c817462ae35c0f1c6ce6964ba5b4a6f15c0919db6435cd29c4499b241b37
z9f954497c90bca422122a31c656a1ee4615a3b3aae141ae06bebfb390ec4d91b7cff384a836b95
z607aa5a8e04d98bcc835efdb362c1ce9731bd4fb3e4fefe895f4561ec52dd7dc254f5a5e09a960
z51dc521a400ce3866492b704aab9defdb3367909c3163a8f9cd49dc3b01562e196f0364ba776e3
zedc45e6209ff5c44272a85cdbff74fefa267d72ed24db3965a971ba889192dabf20d0ffce31611
z05806c1727708efac3cf1984b14255856396d14aecefda54fd888c617ff2fe3fbabbd695908b1a
zec714930bc9655521349acd790bcfe10d716c37ead3e37c82c5f740f4c1b9c31b3f6c4cb077b3f
zdbc1b6582ed3699936b11224df4fc6682188211af53e0679f6e3a0296f5c5626dfa97475ab6fd2
z157eb92562b6eb9a7fe3335bee1b82c6575080b3ab7854fbd5aa0a5d2cea40cff9710cbfa84b5b
z83f3fb771967edd62d22c4c3e0b413ee89c26e866ea0e8b2f6e4fcfb6da7c90e9bec60453e33fb
z74cc0b2371daf908601c5ed067a10997652210fedf2c023d9676973ce9f98c9bff88161d0f3be9
z4acdec2bd7840b16270fbc5a9b93de1205625bb02c53dd981073792d48f80237f34026b8b7f811
zf251f7495d1db88e7cfcc9cf2cc7d0cce816738d98b58b75ffb36c1f3cdedcf8eda9c29f7cbc99
z7bd08799a440cd12e8ae261422221e55eb521331413c08b464f45d1dc9597cfba5574a4c5c0360
zfc89b162e744480322dff9fe53e6d63075df4d1c06cb666d9914ebc59248664c970d15ee02a82f
z9ce205e6c93e0dd9a9582093c970bb2ef9b9bd14039ec2c44553070e39735c80acf7e8f8e7d885
z35bd35045c16157b9edcd03435a6930bcf84d9a8f6ac4a074e4456fff139e789d8c762efff4aca
zfa09bb575a87057e90520c4f33be1022dabf7627619ecd2ab44fa64173d3425ee3bb4d10cc9805
z9d39a2932d3401bec457b5e5caea0b00fec465d75edc9f81dec96170aa95e6640ec3629326eea5
z5900d2f1801656bab4176e8205e74f3f932e6ded6d0788aa427cde3fce7da361a9e6e23580524d
z86fd7cd297ad6dbbfd3c4809e8c82a1075ba30f29743317bfba5992e60683636aeff65e66116df
za977c0771d3818105cd881e5542814979cf80675fe92685c11f532e12de314c05c5a49d98f3067
z4d087040cf8c3ca2f2975b1249de35a0c737999a5d4a04c3d6b72a928e0994ee8b456e91db83a2
zb4780c522e027a7a2f1cd83905faf9d062c7b8ada6218a9768677ce7200b3b959db75042123c46
z330427462268a42562a469c5a127315f6ee88ac8204becb4ea6938bd3426b11741b330ed5056c9
z698e21eab06c7e967a46a3f729b16c27fd15c29618666295f3c5e82940f84d53954a1afbecbdc7
ze3ff20c576500dfc4ad2c3566373505774cec780c92131bfc8535c817b0c3dcf72b4be0bcdfdaa
z307f33fee3743dd8d4a2ab0ec82c4b0d822506bf7264d41446a3825319b5a38b2a1784ce19c551
z2bff1f16ed6317b1074dcb7aa07cb9c9b8613565c22c9b93e3aacd11de558cf29ac1769dccc4a5
z9ce804628c4c6a0fbe30da92f45593580576b967947c78d726c4d018bff8c7e4d6082be35b9f51
z0928b1e95e8e21a3f9755e992c996fb262edde30ded0a6ae426f7080650fe26a312fca09615a06
z1bc8e20c7b5a83ffe8cacd450de9a8f0e74768479130b74edd981c307f65e3960632f583756e4d
z0d35454c5b3105407cf49122ce832056f99037d308905de3860571fc49ae6fc43c923da7e4db85
z40c14876a0806cd07530d4580914b9b941406c18521276c4b500e75f2199900dce557213e1a25e
z2cc88b880405b2afd137c7cb36cd995a50f85facf559f5a1f3eab63f433ea740bc24519b50b9ca
z392b4f5e5569de9d6211db4efbf505bc094b150711850989a6663a56e01959a19b58e2632c761f
z58aeba0d07fe9fe8c5749e9e51c23b1b765880a7246057df323b21b5dafca56de3a06d21d0943a
z32d53e704ed7b8cd39e5271ab183b76e46ee8aaa0918efd595213fd5e3150083ea9dd93be79223
z4c7bb1daf02f429e7879bc31c8e5cbf20baf6da594b72a84f5262008d31afbc04acb11503c4533
z7e6ece64b35cf4ca41e2f86221b6ad134083f50ecca9588d0747d786ea4a7472651a3c7655b734
ze440ce4209e28c22d8feafbb13559c374f721c9bf3b7551fa7aa72840784bd1fc1be6eac66564c
z5041f0ee202f89f5b89d793aeff78a868d8584a83078c95ac314334ed24907729c3bb88f6ba142
zc2cadae3caf6eceb3f95597acdf254da1cb243d6d1ee2bb4a21e5c8e0f1e4440bd8fb955a16782
z4dabc97aec4844940f3bcab05d7651dda68c8ec5384f39df50746b373bffc94bbc58264af1a65c
z2c45478276d70b7f30a2d31cd4af3fcf267fc99b4426acd2864a20c403be87f52fef09a7829aa1
z33fe4b8b494cd28c4f3ba10d678dafad4110e1968f30add232c5aca1a47b03989c45d8c401dba9
zc4b0bb50c9601224878ed4a72d9332ce2ee2e40499ba97a9f3157dda489b6385b01b11d178d45e
zce2c028e706f6c09169290d0244eee66cb5b1e6d2e4a650d2baeb984e8112124c0dcd0716822ae
z0a9340f3fe6231e087343e829612a854af7ca378b096248f60417bd76c96a5cfbbae0664a89fca
z1260d46b464293a32b2d47618aa0c96e1863656b9f0a2507625f60e64d5118a4d3013ee8dd7e29
zef689889f151c75d1aa52db336d321d93514e6e467e23ac2681e4a2eb65c57ed09a9dea086961b
z98a22fc03650a0d512ac61e44a01b1490a60fad344f5aece0a6d9127b1e0eb719bcf772560a560
z2a992380adf2b7f129fffe11824026cd71b1944ab28cda6f589ff4a1d76d9ad2b8f9ad0c0e790f
z4df33fcaba4bae690ca5819594fab08f5fc2d3d541dbad67e6ae5e54c62ccc059ec8f82ec2af70
ze3f2439086d63523052fb116627108b50a50aa3280240d4434a22b7ce4f5adfbb1706eb64acba3
z532a7b570aff1c82986b3eeb6804f80c01a74790943882a2f9b50bb4af90b084ac1b3addbf10e6
z6aed784e3dc4f1e5d901f361315b3a7d9220d7e80f7a0e024181574504a273099bf642a1e493e6
zed2bba735e2cd7bccfcce08afa1e8b654a13c0b622f2f9a3661540a00a97fdc504b7c27b1a5022
zbe0cf734ac6192015c4a8412c45a7ad9456ad624408b1b83b7299409c22409d7c4ae05a849201e
zfa5921c7a64937805537fbde36f2de592990a4efa1ae1eefb39395039971bec2eae3a8cf534911
z6df07e64943ace2015a73488c3f31591e4e510b5d2a1b87d738a6a77e7dd82a35363305cde4ccc
zf6d1333f295d928e1f64ce4da14cd33f7d3edd6896041d67d4b0bb7e569c0fbd73c87992ce6719
z00d438ac8f201407ab5a3e62c01e63f2e3dd2408c26efffd1e3f0f9d5091f089e55ec8b4bb4726
z79d1cc4da6bdd73a4afad0b5e4ab06b593ae312200516e3e8a89c8e0286df6087b71b7764dea66
z93f8d2f159bccc781f2a551ae43c343354f62d3846b093563cca220a35d3792cb5e93f0df132af
z90a284418557dde3919900f2834b00156232b497a4364b8ac18dea4b45e8dfb2fcdf2673a366f0
z6a45d6f8bce0a78c7149e507a30d9cf0306dae285bd64d96db480b4c48cc9f7b137ae0b119a913
z90b5a0fde0bda2c6d85ad5c8b36adad27147e42179226e7a9f98ad45a4bacad75aff96921c53b0
z037d6bb09814a291b3702a0672c2b2baf4431b943ef60d1ab37d70f0564c80a1d017882c82e038
zc38f471e2b9fcf33f6b76d36b011616192709433dbab2a0ef2382acb0345defd4d269d182ece83
z3741d61e766f842e05e05647d2a75a8dae35dd8399506fed25e4228752d8b944ccd7edaf627678
z261320dfe2d9a4aac9230c0deb01dc314be953b0f139f314213b223cc6e90d2959a2ef20a7e9c3
zeb8e96b5cd51f98a9da509502a6dedd03ee1dbadf84443ee2b6db8abccc0caf15da381987be225
zf4ab23e97ebb2fdb5185f6f93c39116409c84829792f6ad03b1364e2453d56285db746c912c98b
zb6840f13f617a9e092a69b11013fc792364e00c415f0964e03c027a2c1d5e9db551707b96aeaa9
z8e6cbd59203ec6f42a6ea3c53a389d3a3bfa6a044a1d0b7c738ba5c648344fe37db2f3ba82815a
z793399b977d0c870c5b512af938923e6d50f8be734ceb5a91fe65d5d9cb3d01e7082d22964ff42
z59dcc11d6291bfbe5f57e2520ac48f57fd217e667cf91106369a22c77d03034f87c81484822b8f
z3c6f3f7ae5c359bdb22c109f94cec841de46b3279d5d61966830a96e0caf44c6ac3a9a3ac5dff6
z383ce87f8f731d7c9ce2d4192b1a8896b6b425e3d6cf9eaf14d846b5e97ebcaed309335d16ba27
zacac415c498f7b16de54aa2e7417ebdcba032c6339ec1ff05e55ed091b67d8b764cfc5f86bd1e0
z958346e6daff378645bd40a7585651b2c79d46d7450bfda0bd7b4785f9d2b4507da08d14f97c78
ze7cb999d24a0bf182f98c261ac46e0362d2792487d075a4b5781559cbc771a936ed78ac879e33d
z55a5129efb1a1df9d8f36a2e63efe808648d13a6f948a599ceeaeb694d0c4024955b6cb2289ca4
zed8adc8570c4b7a29a302f81078808febf64ab6843659639ff55703bcfc92001e3604e33bc44c3
z296e241052f80e86c50b5bd32ac8244c71dc704a4515aea23aa646bb6f64ceefdc832428a0d14e
z1c04beb47a0e92d0f23c045e131986e2d2887cdcbb03e481f424970dfa339548cfe9721f99d7bb
z5bfc9f2ac0380d4beddcd4871f3e5b4a2883ca0d2deb9f253130739db01799642410906bd34d2a
z67b9125fed1acf4918eead0964df1c877768dee172eb09fe8cd11e889fdbb00521cccef78df7ed
ze9cf725516dc5b1ca0c944656f4fc3cac415a1b98c7b667dbdd5ebf6acfe0dda8a4cc085064ce3
za8a93e3a3dc19c23ecef54c7bc5dad3a03b03e32b0ee9a8be91217f605af0add287b3837428402
z43e88c7885357adfd6d0bc359061967759ff92700e6c8dd7a233baf4750d4a7e75a7ad8ef24830
ze2ec9bf5fb734f829003b3d89eb52f3e8a9863db2d4b9389d2d9e41580e3aaaed9974187a461a0
za01684dd1411245592bda2f60a8045716865773acf279bfd204b659e50780afbe34b3263a4f253
z8e2b98e4fdf9dac1724b388c5654e310acb28d0efe96e76236067040fc67b417497387a7713231
z244baf57c0a9866b9af86c9ea4432fb96e857c6a82e360769c73d6179dab4911a437ebcd7bfc9d
z5eddf461bd415b386485096e3885d26b5faace5416807737ea2ead6aacb1a71408ec15a9822a0d
z99ecacce7cc34bbfc9d27fa3708060ba00a49b656016f5329bb0b6fcfe4d8cb1f0e69bf40636e4
zdaf6997668eae046572f12b489810939d2a5a05d137bb1d8280413fb150e4fa25354a27cc42fb9
z073944d46b5ebd33aa046bb693ba7fb4915fb4e85a88c79d3937c6f97d42ec91935228c18ac29f
z23d40156bbdbf1e101832a701ed1070421381768f6ee129ec8e57a7224b36a4b01d79c2fdef3b8
zc79aeea9187c4ed62087a99305a820f99bd8af54c01bf8dfd50a3e15fc9b2e42633daf4de4db62
z2646c92983da98b84b3b75e93099b03dacab7602a9a63a8db6289d904c09f285c2187daf11f4e1
ze507dddb2c1e8284806bea8532277525a7219c14a470cb07075822f66d6088222acf0ef033bd41
zbb051045d0a6605f48d5f49e746005cf7c0d05fc588dbebf848faa36b7306b4b2f969633d1d2f5
z177ba8f3f3f92bfafab730c2beaf97bc0e6552a1b4643fb56e5a01d431af40a881022da22d588a
z2aada1bd9e61d62913574ab85c5995eac5c9c27268b81b7d4f86dd50c234d4ab198d3c225c6b1f
z41ac744165ebbbcb6e27816bd6292392d0cc7e286685c571bc1d5802accdf0a7d76a22f12a014b
zc443ac3db9986f4de1559026c977beeaccec95835da0dddad1cbea6bf69a8b1db094cb20613795
z49d2b6b64a76702df67c7151ef65f6971da2d6e6487b15624338a19779bfde9ffd22d710b5ba32
ze3ef8505d912495c3192b65ea9d6fa84d1e01df53030ce48b4a9d44ee2f57b4bb570ee0192d4f2
z97322ece2fa59e42e17de9bca3b71922b46d5b7440dc26c67fe41adf1b7010054d9230887a93f1
z75aa9a702d127941846271d6287c3edf55a453a5ac4002a1e15ef44498e05cb08f37ede461133b
z58fe6a5c521c901e5ff1897ade0b2cfe24e962ecfa41787d73db7928cdaf8fc0cc2714a9e14d1f
zb5f4aca92d504fcd337a2d374504320399f47c780b032958a5e104950b8193952957a86609debb
z5187629e56b126e4dbe6bd0d10f2b894624c77466f334fb6e767d20783d45ae9f16768f3fb88da
z5388be903eb285511461e1775305176989d32f8aabf4fab20c256a12dcd501dc4756591add1037
zf8719d3c39e1302c7514aa1630e09d0a1ff035a4c0a3fb3ec29417b99491c5e1ce03966d2a1068
z0642bb64046be7e801b27fc67adff95218ef432a3fa5b19f2a54075016af5f3fb213cc88670bb0
zd44dd546a827ee204827b15a276dee63362c8f50b5249aa8eee2c42453329317eae13b75fd0ed8
za1527c54664cc77f916374075b1e3cb69b9c742b07ccb6244b0d618cee583888c39dd0a9346bd1
z330c105f6adacd550906d5504fd1fda125e8c51774b67aa02d0ecb871120ad33790f9685802e43
zc7ea34bc1e72eb0e8cf3f231e9f09b6b2e22d637ff0b318b0f7a69e9f42236b551aae0f01acc18
ze2c49bd00db4d941370a0d49ed8a18df920c7763f407c207f5ba7cb69adfa56137404b2ee254aa
z3e02648760625ac78a419fbb5cd93cd91a7cc71992669cec6c3e503ea49c1c7be02d636a051ba2
zc2ea554b3eefe84d0eef7d0ad6ab31328899a0fb14ba98966eb542177cffb518ff3c66dcd4de1f
ze446d65f258c275da635e10586dffebc77e1c05254ab4d0c91688493660d904243a2d7bbbfec4e
z50e9421ec5c336f1a223421fa4b0a458393296fc50748b88820fd4af12b9e3192a4035886799af
zf914f3fd15e41147a167e7942421c670c083aa3d1fa94ea2d58b8c2cbf4ed6070f5ae1884c477e
z4df4b6dfb88bfa1acc5340922ce342e9d2c3301b32d601910e34acfc37ef46d23061eff28ff24c
zdc41002c5d96eee6cec705968ac60dbd6ed0ba9110dfd9e53d8068ce3dcbc3e8865ba481412bcb
z86f45a2db034df7c0285d52203c035bbaea07c750c17a4b4b06585a1f3e5a6e495b4908af4bf6e
z1dbc50ef52e807d0f008ae2ae7ba4e370582fd6d74e9de62ed53e4d850f0b56c78fac0969c77da
zef10390a05a4a89d482d121a919495129a533f8472c0ebee7055eb431dd6cd9c94ce4bae6ed98f
z63d5f632f53e028e6fd45d2b1a602820d43b6984732b3b1ca8bfe0f4445b8391bef1a325eefe17
z039fe2d650757af29dad79046f0b47a0f09391ba740bbf175c3f8a76a4edd5af1d521ed4c1e3ad
zf07f1434683f5991828a0fb437271a3fe22b9d756e22f9e1b405cdb5b2e29b3c4153adc90b00f9
zb89cf9cae0ab2a31e06c5e0d5c8b0fcee92a76ea396e09fa89446a4c1fc64765ab2b3758d2881c
z811aa58645175ed951f1e22fa372c50f318a836516c1316b8742fd6eaf9cea5f259ec516840add
zf16fbcbc192470d7538ba583f4bc8ec4b702001fd5cff90f94e2e0f120a0475604ce20f947755f
zccf7bff9127263e8856ff5223c792d2173523d3169cda80252f9a93abfcb692dd413ffc7b217c2
zfb43cec03b8733f8f4aace46136d1cf6d054de7456f19f5bae27e0ee79e5c9a81fcee7a6066c50
zf63bc0ca235f529966e64022a3bf9a9c07dced584489da7c91b23bee3608e35eb6d93b268fce23
z31b8f680f513f41ed39e619d9386ace52274b70ea7f69fc089f08388d23a5fb18a58c843e61934
z800e9c2dd5a58464b92bc91ee68fab7318b2bf0d8a201e46075f4fb2def553781e25b7ac8df660
zd2eed5502056dbb498657c239d6b65958334454048743896869c72ccdbc9c2b5802d1db22df6b7
zb5a72d3eb2f9568eaedea8344a7b2d4230b5585c4fe8ac56382148311e900d048ee7138199a395
z0195a05c029d7d67ca88e631e335cdf652c4dd8039acffedef256d3e57ae57f735e6a1bcd61e0d
zd16a994e02f0004ddcf8257b2d88f8c122ec780b13df6def86f6680073813fd7e077370d7b7b25
z00a39e84e22e56196bc47cb6b9dde8be200b0a993aa46eb9666b4094a34538b42a58ec686fe585
z738f8a39c0b8aaf7148935ec2c37b7eb870658fe31fcc80b9b2467cfc8efdb3f68ac298696cdad
z7f70b83e3ea86edc58978581924b60fe361798a37586a785b6a8ff4c40ee069355fc1edfe600e5
ze5d35b8ccb6bb52b5a1c0ae6c74d9de9073683db16483048e968dc0e1f30169709d9d9a121fe0a
z3f6f1eae24d5ccd0f349932e20f8d5a29856a63b01b4c6286740ff89b289c6ef89077cc9278f8f
z07221bf4fa3b7e7e1ac9185534a6df70e7519872ffa50e8d95f157648d90bf349693f216690342
z93262d1e5c4f2f5c6acd003a996de99734ab81d67fb7ef46d20798dd432d52ce51d4dee1c25ff6
z191a3823fb72d7a476ebf51c0d3c89d3c5a99925bb53c4705c0e8825f6b2658814393e8cc5c2a3
zba1ee9ba3b5ad1dbdd1aff252bfdcfe0dafa5f1b1c24b91b3f7b9059ea9795c540fe0e22b9a97f
z06ec522f0c6c694a9ef3c11eb18ebd25a298a34e75c8864e195e2bedf76d084ce9f2a33bb3ff54
z38fa51456b94cda608d9878bfc1bc200f73cecb441d92488cc83221387374c331fbe23aa7d9bea
zc6035340ded46eaaa6de1d4cb1ad25fc1699fa671eb30640eb5415170262dc2158fdc320b73283
zbe92cbf54a3bfbbe424c38ff316fc50d5e08c5ee2302d0dcfbcd310ea55d6266a3aa38cbafd77e
z215e17a924239dd84f5e7c870c102eacedbf83a9fdc11ddfa47aab20ab8b84b3846b789c5e2fb3
z061fe87601d32271aa95cdfd9d670b8710da00e8eb1f06b1a6805c2cc7182118910382516bea2c
ze9dd7cf12bc40fc2d8d583f71c55409c7344ab189b006c04208949830cd5a7f4cc3f3d56319e94
zfc9272a3c048c790d1d92d4741efb71c9854ae13012978f67536881b3ba0c75a662daa48b781b8
zb6ec5434bd28ec10b9ca4c5663b13d977d7d40ee9ca89d331955af3ee61a53722955f636823c89
zf27d55e4a308143b6a9186f223a43cad5cb8b2ec23cb10e0382cbfabd21c80f17666fb400da050
ze17118eab684989f0d40e20d48700cb1e5bcc984d4a46ce46ab452563127fbd4442aa1df5b9763
z08a9725b79890eb072deed21f8599aa90f53aefca186a15dc153be3e72ed7af89333bf11a19c09
z45fb7508d9f94988db83b649315fcaada809eaac595b228c522761b7859d75bf3da889ea2d068d
z81721d7a091b836d27adf1f3a2ee84b8cd22f63fd9b37b909c6b80539a305000752ae334944d29
zaafda50d29773f82fda4200ac30e8e0109ecc343743caaff3fc394f464a0c95496d2a1a5b736cf
z0baa3012f07c337b89dd9634c666f0042bf4166d9704c737eb11b0a9da3b773590b8246777fbef
z633d7cc545b6bfaed364373cb5103fdedc5f3ac86202b28b1732ac518565048db2243b60011863
z0b800136dbb4812e864b37f56370ff57f07e9f08e73e6fef0706d7357f1c890595e00749c2d554
z5f0d19a5d89c113ce9c1ca4410c01d3ed880dd3845045e02dcbe7223f76e1d7e371bbdba1aab54
z93702be4961316b99e3aa3962a08123173f81b617d91d597be20faec289e299dc205a82638aac8
zf3d3c4b35d693d5f155df155f178d527317f71b54b7381fd297cc4be8fe0af3d43b70240940939
z4324786fdc139f911f905f0c8968524b4c173d72cf60ef3225948621d00b09f22fe75d0db75e2c
z47ee384ff5588948fb928113809ea32a0a19b05d52b70452dbba6806d12d5231c953af1aef090f
z4e17fb43820c196ad74cb2c91ace87658f2e6227a3b0478ba6ec7eb02e46d2e9d16070495b4815
za18f02206e8af7501f1b89a78a32dd352cd8062f306274dc01fa961111a977c214146a0806bc2f
z353d87380d0ee127cb234b1f3ac6b8a28054d2f54e1c9fbf25281b3ee47155be88ecf3a586d325
zdcdac8b12ab00eeb29e8f64ec552f96a32698a61f0eb0a39b8d63f791308836e66130f50e66b96
zdb6bb4e825b67bf276fdd6bbbe693d89953687f94fa2bef49a59e1bd59da8117f621e1a40d8b0b
zb143e1c702d4f46c88921c2bb9c33ae710d7a19b7a38fc3ca17f07353579223385d84219ab8645
ze8a1a988aed0179ae65c568bf58b466c4bbcb7f142a22dfc18b00f8d8de9772ca4376296b1ee4d
ze76d06ef17a364f414613405f934372cb360ec062bc1a6346e58f7503b34eda4bb809fcf7add8a
zee89177b4837f54f69923c4d3cf396337c3d00e07205243098a2a2de30b37e55e3a906c55e24bb
z7a4fe7528a3deb831ca0a42eea9d8b98b80588af1888da99ce0d5ad7c3dd5f6f25fc16b4e23eb4
z202eee9c2470588d3ad40f9e788bdd1e176f82592243eafbf71938ef33eb9d7bc611ff77ce7d19
za50dedf3dd94b63682a0454fafe775064b0f16af8dd287a6011af3663dd6d83cf913c0ea127d5d
zf5de6085671b5c8109685762188e66bec8735533f73f300b88ca60296985d4c10bd28fddc47a4b
zc5e165b5aac5a7fb0753183637a6963181cf669718ab5a27c5dd9a2332790729f0db70c0e84342
zdea6ab8b0d2a1a493d9b90b06cfd40a7080d290578f64e77b51aeb1a850333827815a66275d98a
zdcaa7a423ffcc9c25beddaedfe7da52c124b0ea2f0a17911d80a7d70f30d831122c59abcde768d
z20a2058af66c2d12486cbdf62a29ae4d1b95688ffc672d6081ad291b60c2c89dcb1faa65647aff
z9ba2b9b7b67fee057d76db7efeacab558dccfa77bcd1d7475fb7b58aa12e92026458aecb7d5969
zcc656e21d743f6758aa19bfc0745781d2e9600990897046a7c8b61a6fd376f7eab792334ec578f
za5a6a16fffc36db7d33a9842e65cdee5ce1b4198b964043c358633a05652288189cc6a61e5ddf7
ze79d6f370d5c49a62867d8be20e401ec97e96332ddaccd70782f84e3e8e8c6fe1ee0a9e546eabe
z040e3fc29266cae0a7388e1c2e608a2a73f4eed8339a03ccd36656eb700c16db09f87febe1a2cb
z2178028e5f1acdbcb832df99ad478a2df9946e7a82869f473355354618485ee9a7b386248ce993
z3e161e237c05473fb6f252c2ba32b6bf7575176d228e00f3c7ff98c0e1394cab51b7ad395c5815
z2711a4c7e5b98409ea62c7ff533975eed6c97efe04faabc4dbf730f147ebd44fd7e30dbc842b1c
z85d7843c4603f4968a9b1f1eda4ede87bfd918f45e3f3d7b6d2f63adce43a456d6730c6d329466
zc471dfa0ffb3e6ec053d1762a61f7c4d888a8e2385b72dac64b85031563a73e3fe04db0107ba32
za15a003c7e9a98bcb96a57edb646a0b1f4f780a2c1a02740b7b006cc4132f5d3a66f0d440ea486
z2c82426a298194f867531c7e543de2565bf6fdb21a64bf3629a51b6d5ce63513157ab8d0817913
ze53c5dc2fa34f5acc2e01cdd0be339af2545d9b0790acd8dd0643c9e71afd5316511696769fcd8
zcdcab43b1c388b2cf338cc7868242d963c49e2aca39f4d7bb816b5b5bdcf6eabdc160f80bedf42
z4d51874b4d7f16b52f4aa860b5678bfe6d73bbc2433933d99162f954bd5bfc9ca12ed142a64d02
z068a8628f69461560124353fc782a6140f3aa3c60f1466df84271522551c3b42993c4e12c52b2b
z17c9de0e2fec2cf11364f5f0495cb7bba45cbbc4f867b8270139f436de118da00b5d12c9a7bcf8
zc3f3dcb3a4d0840d2917a1845ffb4c5da5fb0754ea7092ddf12c3bb93ef23ec2fdcf537de25e60
zb50a235de5286d4a577e12351961c5135d62de44409e29bec6242c5a9c105191ba41498085b8ed
zcda1c20e8c3dddf0d009e5f49cf8cabcdd2fcc925e9c9c5da5b88512608fdf749921548b9b7d8b
z11f28cf43c4c5fb79ee6e6f35e3bb68425fac756afa76166fa40be26d21ab53dc4dd08f922cc95
z6b8b6388f7440931c98a73c61571351dfc30d4847b809dc6bcdcc7faca23bd9c0e3b6fd60bfd5e
z75897dc4a43bb86857591c01d0d9edc3e6c18be560419fcd31bc79b877d8823d6709214711ffb1
z6e2139bce732391d618364090f52b82ea25a00933eed32e32855a46b9ceb69cefe989a48922beb
z773c68e24489309225889c524e6fb15157fdbb4d2e4d05060ed92d7872055c40d05b82aad5613f
z49f664a816f6ae7eb9f940f2d3cae4bdb34cabb63722555f1c2c6645a8646894f7f4342d3e16eb
z124ba050b7b11c9b8662446c49e0566b92cd2b74cca35f89d30fa86470d64a226655f5f1fe401c
zd26ffbc2b0b361e6b4bf3cb6591f6f88909c33949158c4b9af1a2154764709f4856bbe3bf37c4e
z9f212e812e7aa94ed2670524f314552da5252fe7b418ff1e54248e40b769282c091b8ab17c3c3e
z8f5d4dcb6816adc30fd7c9974f070e92b2a32e35fb6b3c6e4128ee1ae73ac44f9bff278bc58270
zcf5c2af5c8ee35b88ac521cfa9e0a910225b3f8fbeb18cf1c5c13c80ef6ad64f8fd24b1578a827
z144be36e769e938e2c92bfe60103ba1f933feffb6fe5020d1757a3e1fbfb9b9fad4b65d4fc998c
z8cf93cf36a5302f1a7b0c9eba7f87c459ef48b1601fa4790652cb4f1b6f4148da99fa479f89ba8
z3d941c9b04719fc567aeec583c6b461a82300794db1e62e17dccd2b0d5148972ef4a12645bcc15
z6de0fd02cee94c1cb831ec5a3fbe661af9d279b233657357702ea8fc46a360b9452526e526f7ba
z001c3d6ecde5dd80a865849f60a8ddcf1c8ac10646d1f9c5ad94d0ce68e36b3f8523da10bfcf76
zac301b5add323f29c2b19bd810e429d089064d2d010674bb52b0ac205fc478a17f7ee621ebfd52
z743174a5b8f00deb01e5417bac4f7e880360b31df5898f057b74bac5202e792738fcd1f18ff921
zcef48be4b04a95eab7d20ed251b639642280e484c7de9294b973d6799bc181c5dfd7e6355a048a
z46645fad09d967eb88ced5e724884b6ee85060ff2423cd7967de6cb440ed6ebadbf7ac730262ad
zd9fa4464639764396f155637a141832c025289269fbb14d357cc8116a3ed545d015ba384ff8476
z2c6750de3b543ecee1d075dd368aa9a80d7df91057675d8fd3c70bf73728a9d846971573c5dfc4
z766f1ba29e03f33bfce1e7958b53c3672c768be7cf026160616ba2bc83bdfdb8c3ca641e6d4a57
z1d5d552f67259fc4c439aa98a0a56400ddc17020ad2f064e712bb191d26788fcd0f7db6188beac
z1acdb03c053b07ab7c34a661c864bb0f89fc4fdf9411c3c7ab812a51f87f8f953ae68e45faedc8
z23872d09c9685257c2abb71a32741710774efb64112d7415e564630e55e7ac5ec6b578294d84a8
zf226554210182008b2df28de79c2efd004d0d04f128a1db5f542a0e87f2c26274c4fe24864a4de
zd16512ba610afee6eccfa350a9a559630cd091f1046472e526e883f32bc66d1c73a607f5619302
z20379286f8677385b7a94dedce994449aedf426641dc4b35e7cf06037d1b56c591689841516056
zb96b9fe47650b938ce6b841969a84f84d0bbe6678a60a5efdb27c3060096e047985b81a8d6d808
z91df343da0e87262fa73432b740baaac194929767c3cb8e15de78dc5b5bf446dc0762dadf83ecf
z3f906b199e8b1040013b6c0720bb0386a5370a6a72ee9285273e565e4264322fb4157dc8cbf6c7
z1eea578cf8a89b4c0a55557dc7c027f61051deaf09ceb0a40ab1e39ef8e874843d595642c48716
za40fa9ec3719e6871c1f4b1a8be6b44380903b1571e2794b71c008a85ae34b6dba8fe08d05dc0a
zd34cc64c8f9ad56d6951792f91d22c818f4b4489f26c897d8a0e10bb3f10da9a2efd607c31ef16
z1971aa6f1cfead0166d349f65bb7343696f4708ce3ca7371fb74d8dc9fa4191db139ec0274535f
z8e3756bf4e341c328b4b76a8c18b7e0afda865ef8d3f342e77da5732c19547c6c4aca15b62519a
zf6bcd63f0c82e9c8414b4280044eb98d658ddbe67feb8f8993f3ea19a7b6f85fa8390f5b7ad14b
z327f9849a7ecb08c678e6cf9ffc4f18180b7bffe469258d6df8c9c275b1f73194b298c4de18bc7
z17bf30d7f2f0797ecddb102b621b5b45c677bd1c1ad2236bd9b078588aee328d43b2c0d7182116
z11305fea6529110efc78c63a05d5a1131258a50546540146fc0e1e70fd837f94dfd434f00b9270
z3373f912674e31876d091e93fda070f706f9b6a23c2321a42d1ccbda6935bcfbcde4509197e885
z7bfacd25d6263a09b24d47fbaafe5ed791304c6596c5af763e7928abab79857261c5a9e9fdca9c
zc26904804e62a35d61762cfbdb037c25bd51f9c5a4b482c55aa26ba4f05d54f172447ee7a778da
za76ed62c1a3816a80244147a006a380a14065eebe45767381f7019c805242fec2db77f6223c951
ze7600e76b6f1c2fe8c4971b3dd8c332be48d4d1d03a9910adc1f6052a04550c1a664525cc02a13
z57e8d5c644f87c42ee92572e4e41d8cf9046127ec03a6764b80d7a2e707b05e03b0ac3ad0f39cf
z6954daa40c78cc26132025834301406179308185695e778662adf0ce7e286f99d0240c7eb2e1d7
zd60da01a3d45e43de2bd365d4a0198083c7420146c6292130ecacf10815425a23fcd52c7e88c5e
z691ddb033ad74c490070043b4e410a8af63ac05f018385f6f7b080ca23fdf88fb83df53d43da2b
zd452a218a6603c3d935dc6287f7415b7514194cde679e043b6156ea742cbd3fac0c0418aca4abe
z7ac25e10810a5e925e0153bfd247da1c0bd719665ecf5acdfb187d5c729f71614b0c8a3f210de3
zbc4d7f9438968f5eba3130d21ceafd7c4cff0e9fed53ef0b25f023ab34e56341d0b006e43d1ff4
z42719041ed90a93a01cec6b0275889b8b44c62d9cd4b7ec5c1b913647bc2f23936833f69de094e
z75cd2cedd3cdd6f65be470cdb03a1ac7b55d7fc4aa161f7d9256135add64cf8d53e07a498855af
zb370767b4d44d76485c356e54dd9479d1dc8da3a3d64da33dc07555c84752ae6433b1a30c11925
z057b6013e6a069808061f3768aecd9ea83060aad3a44f7c189f464c5bbbcc26f21affd42b7c2a8
za1ef4cd6851e1ec6db10359470756f89757ce157b17d3f57cd14519a45cea0601f34ba464b8b0f
z888459ca4c289b1c9020d41bdb1686523046cba2141a38772acea08681b3531b86490695bccd8d
z011732ea30096766e77eadc476d792390a312550170bc85235c5651d5f6bc7cda9fa6eace91d0c
z3c09cf8e7c6b83468d36cfc24f710f1f2bb2b5d43c22590596066e899204665fa2e27f6b42da95
zf56e05a0d02c0c1cc03168ba7b0c25307a2fad082412862a730d61db407a906a2d798131c27d6b
z2eb57cb10f86bf5ccd3f22f1cc89dcaee516867bdc6e31c0873ca3d568a6ba42b3f043f018cd34
zb67e64562872c50ee9703452a2b8d688e2936b2efbd17baf24e0a0f0c9032fc763ab5daf150c31
z9098f3eed048356bde0dfbf44f841fa921971c33545012493e4b5777165c9fa0adfd30a94fc2cf
z60ee54101fef1c2245c183bbd731b862bcf603d4e3e392d0d07940dc396d3eedcee99ed6acdeb3
zadc4d5638b25fb1f21d8c9199d0ed5be35510cbaefcfd59b0f15d83a99f9e0dad608928dda0f04
zc08bc5f7a6cb43d02d62ce1425622dfce0c8bcbf74403f42bdddb559489900d820e70abab36e04
zc74d8160ebd0ec0aa0abce68e27d599df2c88fee5e015e64f6036be816632d071cf1afb8562034
z0a86b1ec5bb74b2a4241431a2db358104be95459c0ec2cb543ab089457d0f487088326258b0c72
z10892a988976c228333970809d22de758d515fefbf7b8b36b974098e68c296f53140eb6c50a1e1
za066a3a112bf54c0d4198fb8f03d00065a3e8d2d6b9c703c114992165c9b4dfbed8e1f1fb6cacd
zbde36684408afc9f8b15f1039776117396ee0ef41688598b33b7cb0c6e613c098ec821f5adc13f
zcfeb3b9a8385b94834608724497541c9c19357992a35bc007d04454189c367f7f7358de739944a
z7f582b8bbe3a4c81ee5cfc7e952c769a0ac2aaf9510faaeb7c5636323692e6e5850068e26303dd
z0240647397ddbe0dab6c6fd771ccfb411916bad24547578fe5bd6ffd760e22cb9dcd44966d8822
z503b418a1bc1e043dda5ae695ff914e7d712e70dc6648da00fb2c8592945f6a8d9777cfca80c75
zc64c5ef23eceb056e721b112add92fde38be577ca2d10b847124bbd52fb36dee47177ba6b201dd
z1cd770ff315f59480f16a8dc13d1fe30a664c6de7d037db3e117758ade8467a72d5090482f1796
z1e339469c0dda7eb7df544c33284f054eddb080ed3fedd2cba2c51e4232ddc2e5b1f8660171c50
z748cf2c25985aeb66e6d70b40aec48c124ea9859228a5aa3142e0c63495cc7a698c77d1c4900b4
zcad237ac6eecc3784da711f2dd5708d4164cb3e2798cf24c83f1bce712c09d3b766a9ce0538e5b
z4b8c69aeeb87875681e7e12bff071755e23fd435b1d291dd5028bef2087e8a37fbe61b98fa5e22
zb59129da6605dc7d2a48f28acf3c061220c51b13a4c78e21e84653f566852fee9e4a5fbbfba1ab
z22e0fc091bde6b7a73e525d11b51bce1365ffce3b2ccbbc1e91e9703be03880f89d3295464e1df
z6b6aca1d4220e679785450ea2a1d8e42681f89ad8409c568ff380c32fe1f3b6dabe6b4e90a4deb
z0a7db763964d517ea17eb32917948f646d0ea4849d503542af025ed672cfafbf9cbb13cf90c3fb
z75840741b8446fd498eee4227b8745bd3684023095d286282e0912f89bbf551c590c28a17ef3f3
z3c7bd1c1375e7668f3997ba4a038903861ceaba255dce57ecb0b93c510b4e8c1e03f8f321b94f0
z47391b094843881f318a4266f15be6d3971aa7a6e1a7f9a54271f5288ce67ae54ce8fa19b5b7eb
z3da755f4cb13cde49217237146b2337661c860605840770f885b6fea7ca285d7efb39824dda267
zfb31bcd9f90ea86701e2c3fe7a280f5d63d1ec5aaaef49349deecb1343205ab76b1a91eabf3ae3
z77cd6cb2796ea141216807525c6d64988616e1eca5d2532cb75feee4c082e12ab75653eebe65ce
z3606a8c21dad7fd5c3cd6a48300485426a6678d954963996ecaa5199026d4fa8f9d7061f855147
z8cc2bed89287875f66c8586bca931c08864b149697d226242ca90990f8e0e68078d720219b21ae
z7086655563830593e903c62500ddcfab085f31ba91f57dc52500b49701c8d827386ecbcbf48688
z4ed08745ccbd90a8f848e3bac68b96f95302125fcbcb08aaf18faf38ea568728b6deefb44ae68f
zba57a0a9b835bb21132d60df420fea967403e127d931809c21afab74b32d95537d58e1501f1afb
z790df4f970482338fd979ee3532fcdeecbbcf0641c9bb3aba994e4a854acc5068b79d149b8d307
z843f9fcdfbd4b9cb92dbed59ea99b282d67ede4457456ba0ef39b6e4ee878b4bffa44ba7a28cbd
z1b3a6bab68b95ac29f07b915bf07a68b931bcd6d74f1524dfd18dd822d2b6e90dba546524b31a5
zbc6e8a106475613ad6ad9522b58098b0616b14e84f3d608d0d2f6c0cfd6ca1e7ab2998f81f0340
z2f66947aca8e95c9334cb5ae09501fcd4f4fee8a6d066901f0e272d336f1d81d6a9b1ff67f02c2
z270491f61b163b15412a7105008b2e2ae8aecf6bbc6d0c40f83333c1d91b4bb0b2bdd08a5d0fba
z5f8ee323c1dc5e56b11e7816c1d4dcda2bb0ffa28b9c155379d3889036236cb4538288b9b0f6dd
zbd50173e9d9d10593c40114c54ff275d000d5691ec14bdcc174d7bd8a6f707a167c9cffc56c75f
z7662c5e27e8437311c794d4fee0737f56ea37f77ddbd9fb5e97ebf9846a643c6529935db454c50
z5f561cb97113341962f1512aefa6708da3c52519d6877f7b592584489db8ac2e547a81731799c4
zacb89bbaf753af1d3032773136d6a9f6cb25e82dc27cf3036b1474f0cd42e34c8a819e458e924c
z89f1b6ddff674ae243053a7055acb2bc5bbd00dadbaa9e9ba1be187dac044665b8abe49777bcee
zf96eedbc2ed29d74b1e54c980521948a120a8e44d29b6339ce8b5a9f79baa762d2f077435c4db7
z4bc7a4e897607517f7ff0f3558d0a952f301205489dab6151321026073568454a65b148d682483
z8d159c406a5de75a21296a31ac9e3c7a6c37d034c4f772578916726be29f4bd109685488ab6dac
z6ed0847a62f608694a9efad6f1ac7050eb492b32c4d3885915d243bb871771dc1b7e79d3f431ba
z1776ed08ff03d1f49175f924e2a4ea5e1a4d86e3c1d478691d227f2b7c972f3816aa48494a8b9f
z00efef3c99d1714a6030e14620fa925988ba3a8f54708c6b1c803c08409e170e3a41ebaece7aa1
z8c857105c11d79b1579ed4bc2871a8bd6c6a7ffc22fb6d1c6088aec8ee27c4321a255a00166844
z9ce69c0cf65edfab1ab7543da1192bb9ccdc152ec2223bec9f2dbdea53fb347a3afcd91b9a79fa
zcae68188631ac159d63ae9b4b23d4e9990024214b4cdc3469a8df677879d1a87fe39ffe7764c14
zbb2bd110ca204ca533f593e2de1263cdba842b926c979b8bcbd3a1fde85f4f77aeebb0d0745d89
zc52a4753344481aee009eae20f16b0f2f07fc75e0e6ba5a781ab94450534cef62048eb9a35dc9b
z250b47d00b2ad888157842742d32af2cdbdc645d7135ad7b716ba22c5e75f025862441c29432ab
zf559f0ba35f3d899d50c14568fbf9e49b71641c15705af2751ce85d5cbdec657145d6df6244164
zca52cc23261689e8b4508c1f891fa84a9ea359555366746949865dcda9b61d34d5e38dac75953e
z70a0c2c0ca037817b0df86883b0398c0d9223b844c6cd5e45b08cbd3d5269ee16ba256c67e0bcc
z2c9fb7f899aa913990364d26fda776462cdeef4a1e0d50a8901c709a9a17086a88de23672b35e0
zec1ad43ca5239f6f17df0616b25b7a44480e2609fb2ee7a6d4a585fce12ee3ec2ea5e111070e11
z6cbef123425b779b12af4c228b2d5dddbf08ee6f2f07587920927005d8b4a2ccd56448adad3cbb
zdfa75a730cd44254ec2c0a152ae0ac040b793af3aeba6fce032bdc1e100b3bf268a7de83b46fb2
ze2bc157bc3dd852797f4d77221fcf751dfc70576cd928804416fdd1e8b843bd13c551e74993779
za0b3f075e430d13ca3c089d78b6aee16b96fbc96cd1c903b2029d3bd4ddb7358b1df6b09d4ef98
z8630b4782b4bce74f25468c2a978419adb89a175c78d8fc8a7cfacefada2a02cbf4351912784d0
z9867fe754a92683c254e70fe7babbf7f722314596eb77216c7b34797b2925182f39eb6f2e9ea05
za8c56190b2748a942ac65cd666a8ce9840caabc7f18308d857b2f0e0cc3ce773eaabed58237e7a
zaf8dc99855c18cc5473ded2da3aef58b13b8aa2e9b0dbd56ed58ca2649511d9309794e1a2d74b0
z6edcd8602fe1774f86f6541a182919aa65229fa5a342ee3cbfc6c622d3ee85b4560a3d68de5278
z35887509562edaeab2d7f22dfe1ed8d91b1e2a4e29f2b73bef8e10bf8eb4b49a1a1f6cf2d40619
z3e62032390a54b09b3160782643c5399f6dd472c80090ceafa560e3ef3f6143150b1a69ebc80a3
zfc97beed15abb1b6ef90ba53db75e075e764db8f0f12ab8904a5eb5328f94314614c3fe03a145a
z46e6535ea47303a477f0bc8e163423d9c23fe4feddf50d913b2aa1a0d290b45ce46b9399210224
z0041e8ca62f31d9907511252278f04f7d5289221ae003d45fdc763b0d85e941fe167f6ca012365
ze6beaa1f0925da050c53c625f9f60c2cd469156b96a4a680c474d6371171a7df4bd17004fc14ef
z0796fc0a1df4bd4634c1ea524d1e8b99fb0c69398782903882e143d42a1866c3296aac9a733bdd
zeb81a023ecb611c84babf03728fd4bad2b1ef3ed6ce1f76ceeaf564d2b371e4f4e4d4de3dd7baa
zd1d7a7dee6e94081cbe4ef4de5af33ec1d974a18cf772a232c6b84b8eeaff22d7a1494bdae560c
z3848a021dc31265ca7da5d50984fa36a42ca33f29b84f09cff5e36ebd7087e1836c9d6f9c8944d
zb2e0d6ee6e178e07763058e5267e6c467ed3e7a8425699185d794ed0dc637bffcb21361f8f780d
za2e9d291ff1040cee2297c636ed4c49892c30349e0158e415f854973dd6a919907584b0e82fe2e
z572b57945c035daacc28dc70b8a7fe0ddca0f66c0b4327ea719522b866debbc26cc8788dacd979
z163d504f324367e554c21c1245443d4acd5627705fc0103f00e69342a7001ceb6af451738ca44e
z9f768907cfcf2f26810f26fc16e0f461ec5485f7255dbd6e1d94521ad6a8955d81c0c578ce5cef
zf67917c4fa36a54c0d189e51d86f873ca7300d38f127240d966051bf5a17732d48a4e5d2c960d8
z316f4aa8b0cd446524e4d35bf412b7dfb545126e9a5edc56e5304c7d59b152bb499bc270f434fa
z393cbf659c9a9615f05f0f1a51e60602efa56df612e5fa404afda0fe75622f0b986f427fca6b1e
z5b2771d7ee85e20caa2116879a43cb68fdafc906f8a578e53ac99300a7a728f98cb5b43c53b4b7
z10ee8bfa9d0233c0cbc4b6b426c2a36f19adc734491768e57a08e1ca09340da986d2d50b7f6bb9
z2a526c2e4b41168d55de58340be58fcc4f293fb8cd97bab69154e0a7c00cd76d0e9dbd1d396112
zf3114a0b58796d48fec405fdb2c1e0c9f74e37a24f214688cdbb6ea64a7195ce35fa370e2704bd
zc014fd5b623019e79025104594b5972cdbca1a07aaf8c09f7ffc218061537b6aa8030144f18522
z97e4bb9c59b939da619ae762791bc586aa59373381247f8f3b621dc5c68f13a0c26e89e311a93b
zce6f7c36381de8267371cb1c484a3d07cd3d05036a147086c0c8a7e51d60640765f58e96a6b1e1
zce442c4527f5f1c415b291fb28467f7d965b2b2398665dcd3313d1014c0db43e98fe29f6915c10
z82d7344a0eefd35e1f4bbc8387dcb17bbdef986ef3644511cd6a56b1695b9afb7992b6858db6ef
zf64ac39d052f49feeb9656b39ae36bd765fe3d19ce5de73db14469c17796a90c7971a9a0d8b348
z0935086370722a521ce2933da2b93b475079bcd863021ec91031b6398be2355b4a9df32b571e8b
z82907a22aa09266368463cbd94d1e30d1af97b9dc9e09131e32ff16e8b36d4d98fc8c8c17154de
zf1b41b34ec498aeaa0408428fdb18f5944665574d99aceb721034aca9fff837b10895ef1643b76
z637f6600bedce2ee117b0723c66ff7ec30c20da1bb28f633ddd076489160ad8a62bc0317e6ab60
za455dc1e56bf6bebcf8222bb5a35f1bb758a5b27c5c63d3bd966f468ba61bff22f08831828fba3
zd2abc19c2a2df279de2c91703195da06243184d0e7cf223783b954c50024ffb382822d553d0f76
z3f94bca82a83505e732b8c445de07ccbd427c05a486740ae86861759e78ee41b1b5926b26ed172
ze15662177e065f6d30cb75e0cf1286b6d011bbdf83c799f77cf8f98b22a87167397859ab9000ba
zbe88ddde5d1158af540ecde56ca8a4ca0858ec79c9e317d25c5ecb036e63636ec902ca9868c2a7
z23f95745219711ee15ff2b1e1c9583e925361e1eaa6434d475da98f1e1b45287be0b2f924f09af
z4b8ead92633ea448792820ab96a649e0167aa6e929d4f1609efd3321d7796b27b2b542863f22b5
ze810d422af46610cfd47805e62fef6f01e39dac02019d99dbc62663af63c03743a5ee34c3e4fd7
z42070c91a7f7254a9607d794d933f81ea034ec23bc46ce1a3309a6ba4c96646ffc355c5f5d8004
zd662fdae0083f04b3c3c86c3a16e539bc3749ccfcc0097c1cc228ced3d327193f9ea50c31794f6
zf3c009200f77df78f38e790b67b05f9347173595d61359d332cdec80ee74122911efd4cd19e095
ze9b44c9670992ed028235fd04434c8a7fd8094d73b3e56566480cf90fd44f38e93213d35e74841
zb11e53bbe859b60c854ab714d3f0f018ba267d4ad402ff7e16a67ce6038d9e8d7c3f250cd23ddb
z3f868796fd85489f113134bdc9ac0b659a57e5b18dbd9c8f58099e75a6a34761885574227875fd
z61660baec16c57196b3ee94643e08eeb031783e69548524466b1f90b0d3333d0720ecb41a3cbad
zeac08d6b45cf801656d6460e9352e318fca301a031d6a73e87ad906952d04ca4d3642e80736788
z267a4e443d908538da4f77ae564531551955017b2fab235df11511f1b8b314b7865e0b0cd75cc9
z0165928714c76d11a5229c251506a04378f461dd22f059fdbe95715eec5724e96bca90e111f6f4
zf4023bf613fb0b1ab86b3d5dd6fc7cb27b041497d06e1b2b790e5a5aa956671551fd7a17d35d7a
z2d6fc0487b9b469a16ed9bcf50efa9938cba784970828efed73eaf6accefd7369679b9b376cb2f
z5fa0b6a40ff2e554f97f6870da9bda30697738f14f859e6bf3022b686f4b034955f090a1546a1d
z31e1150246033307eb6b0f65577b712f182fd9ceccccc9de9d9bae55a8f9de1b841a8f23957c0e
zee2d9da82e3e0a1245cf76859ccfaaf4d79346efa0338a8615282134d5ed329850ad67ab5b8243
z62d3b709f572a6b2f3e8bb619f8ccb318da1c1ed4a1950544c763d88dc85ebfc8412a7f18cc236
z236b678afe71fc67325dba95d4f7d0849fe63048cd296d05da957bdfbb6aea020e0012ab2432e3
z0bd989e6d7a98d4cfbe294d81530ca9918320a9e56a1b722e89e69d0693e69a1dea68a9ed2bffa
z9a21cc7fbef1a5a8bbfe7c674980b5f0968fb1bdbf9c0170014a3843dedcea4adf3e3252b44190
z7907a45165fb929e9c5acc75b4ae7ec4b4c1953cad694152f1dd1f1f843e5004feb46c16d1bc18
z257a0e43905479811405408b73e869ac4fcf761a46c03edb16b1569e0b896281a4524c2f4a427e
ze858d8b8038b3ed3fa41e955fd45d225ecffc4777986ee746686793bd3cb4a1dafd870138921d7
zbec56fe52ad7c2b3c695a1ec7de308318a794248ef050609ce325c84657eb2aa73b85dff75987b
z0de5a369b923b555a80cfcf5ea9648aafba1b52cdc58863f137712aad42550f80ae4812b13f67f
z38581f7f5f7e0f6d354b27c3d717d75cc41278d63a0099a45b55b107660bbe0854e302d50c8bfc
z04af0cc1998b9c6bb04c2f55668bd6561d01514bed07c600205b54edf14f5cc043367f13acc723
zddd5a760b5636fb1e6a821cfa3dfd14f4dea1199468a007bb84ca61ad4394cd137530d51ff0c8a
z17c60c5cb178c234275f16e4dd3dd791f28f96fd689eb0e83a11d4d88ccdc5e5be470b48edd482
z86a2914586ba4318283867258c4e2fcbccebf7402980a9e173485106b1c2dd73d875e7ecb2d79a
zcacc410d8f0a0994430b50a3b3feccdb09acedd0ccc4f3779aceabf67706cb6f11a662e6cf7fc2
zc3ca2d106b604b815ceb1b30333956922722774d33aa34bbfc0538b6f86de0712a8b93e257db99
za1992ddb83fa8bd0e5ddc165b275410742eda483cda71ce7ad0a3b4bfb15c84f5f04832f46957a
z37c54d4d516a01f00878e27f02219a28e3da3f3f51c75063580496a95bc8410548312d63e98098
z5026bcbff626be6ee535c3ad7a9ed82e66345aaa8cae5d446ed6bdd0a2fd7fc4dfb72786cfd700
zf98d2b318274405c5ae94c642eecb64dcf41dfca704f1ad16891032e38cc4803e56972c53c5374
z91f2f82d7d7e7bf16ab547d7135d944da45580fe5b3955c51aa41787e87965fafec41d16b1e140
z8ff9282f6e6c0ce2770c421556b2595430d02b25947668163c4ab9cfeb00f3d0e23f53db5d6058
z0891f600f39ccd6355a6fcf9ac6c0ed3794b89546da330fc81d27fdc745d81f17685e3fdda644c
zeaa5ca8238cb2c21cab5d18080a19063b0a6bfa0e23c14d7962a257c83597241ad7d5b0053a139
zc2216194773e29243a4475d2e3c1a963d3e103f11c3fcb23a4f0617b61d218cfa68b8cde678d89
z6829a829bbb1378d59854db5841c313c8b820209519af0c53165ff7ff62196c7d4aa772e64f10e
zcddd9d8aa57f407d0041eb1b852fcbcf23012c5eca05e328b9730ffc5d7ded7919070b69dc17f3
z2b22ea04d4a5d89a0f5fb544a6f04a6513ef8b659be302d6ce5405ec7650c9c032903dd710095a
z8a1df40bc7c7c6fc09974de8d1ee2e9f82fbb61a8d79aa41b89fe443bec0e49a6a0c1fdebc2493
z45ad5d6b1d49d53a2d86521c59a08db0f72eac27e95626b201933c5009e3adbb9091f6cfe85e44
za3a2dba4601344c572e32f916d366bd66175dce437256e77818972cc6f1e127e1dfd3a7043ce58
z27ed1545f7d173da0021f06d08e11c1a33bc12dd169754106a2d8ce0b271e288d1a7c4ca68cdbd
z11dd76d3201eedf96c9dc242a3a189b75cd19a61331788ac6f02963b1129141a42d0be1371fd3d
z22cba40db5bc3f1b6b7fce12c78570df90832670536cc8bec70d9e33e16e78df139477a48f28a9
zf4f62f46560ec6d832ce346a8f30f5ef04ffdb1473383be48a468b59b010cd7a2722f6178df9e1
zed75a342386af3dc2527940d615d656ff51106156f5371010087bb16d789f5e6b5752af61e8952
zd1cd3083440721e813937b8ab9a27d2d74673c3413af72fa363328fb9e666ce7b10c042d4ee527
z99eb9d734812bd52bc606750fda2b31d35cc196811929e080591619e7167ed3e14f92fe2cb6f53
z2bca8ba74616382ec4c6a23fa6f048152e4dc26d755b5eeefc5fc7b8f5098b9087c8d4eb07805e
ze65a2a60aca43972940fa5d6c5c650a6a760ef448bbc716671e586e08e80bddcea823dc6d6728b
z95eacb72d1e192922daf719d8d546efcfc05ace33d5180eadb5c8c2ad277437c74011c89d2c745
zbb0e4fd4eda1ff79379d27209365588deaa01b1b5670620828a6513c5f29a17002feb377c75c88
z498239e7857ecb6646572ad11e52ced6ccfd0feac5832f36925184e0518b1a12b4d1654d1c9d56
z9b5717c6e75122773860fcf2aaa019bd68d1632bc1bedef84570a98d493150c69dbddabf178831
z15387a17fe4fb40ad41fac1de715576fb18701a91874970a020bb681fc407422c63fb2aa32667f
z2fdd7bd00df0418fc57b97d14e2ac80ef47f0bf0cd2038d833d61ea935868a7e8f739cbf8e1b97
ze952f0f836d8ffaa76f7f4f4515ef9c42d825e3f0fe6c1d3236f73798a9b85735e083911d09ac1
zb46fef94f60ed8f0de47e2500c826104ea4075243691197b02a59f96a30b490601ca09837ae66b
z4245c2d4057f5bdd72a431e070d1fd0447359f7bfae3adeda721fa2f3cd4fbf955bc045b131e40
z7c3745d7ad5b3b523b9580c1ccf971a4a7699ba6bb6fef12fecf3a147237255c0b1d1ba00a9abb
z78c775f7fe71ea9cd65a26746e2fff1d5cdd2f96a51b8f33108fad1abe1871478e4ee0e7e33801
z06c440eb2502ece1f4ec27ce62cf1c0bd0678e29d7c5b18c8a7e85bef63e03572cb2410571e9c9
z9a8de869522975f1a765c399d99f101674aa6addf07844514debbd557cf3b866e1279cc26c4557
z26d2bffa3c86d7267e6ae2e57c9e35d7266781c74e2c4b09341c6ee0f449383dd30161da69bbb9
z3e0d581303e340a224ea53939fab40f42c6577425d5bbe2472451066d04bb44957425ce273a590
z4418f264687cd6ab01bf8b3f27dd1d021970c1cc6086b6c1d2bdb7a7b77654551dacf8994565d3
z941241f6992a1fa7693d470b68fb279934e3861c2afe1379636fef647f0ce647dfc48cb52ec761
ze9f6e4f43b651c529a9ba46a32d49aad594c52d61e7253d8649a747bd5c89f5ef0e2a217aed38d
z07c7ec05abe4f3ae2fa2b0e9ac9c1333da3afe9f63f235261d6f1681dbd7e2fb232b22666a7928
z6ced1b15e46a4ab75c525cf526c8022b542a8cc36ea21849396cf89d489537d9067f76f5ebaae4
zdcc972c4cbbc8c06b46418ef627be5a9ca4bb943642ee9b5214e40c09b3d3c4e3b115b151df4b5
z94529408df2dc0ad6e72243021a1fee5303a3672a68d67d2ba85d927aba04cb47a6a2d96719292
z90e8fa542f2a5efcb7b85397329ab3348152e98a1f1906ceff68595d9e7a0875dba1273d045d2f
zeb8cba29d4144ddff4a4f98dc232cff7bc7fdfbae6c7338035ad529bc62673c772ff1408ab0de8
z3faf417dbed2c03e861b7a531533838fa5c4795765f178940ecb4ee961a24e759bb076dbb3e61e
z1fa8891e5050188cb2ff081006612cddd03cca9602314d7fc08b783c2b394a7de8da53deaa8910
zbd09f296d1fd85aef111b7cbc711ebf08fa1ae527dae2c571affc0368e547df8675d9913420ffc
z34aa8e7957a7683bbd618008e70f030d7d94621534eb145bcb20128e8a02667fb397380b758b03
z784c266589dd7f2c6421d57f72dc26a6bcdc5c0be60e9a588bead99c32d6a877d6588fb8f9c826
zf4bf3a964ec4e42029a5426b2bc7e244abede32016e6f518828fe1c50035ec81cabb9d9c8b8b07
z1e235ff503391bbe5889cc0cda6fc36ff23f949abdbf17d890f754d7e55a01fae2b1b15f1ca897
z3adcebfda066003fd0287171264f97f3bbb230cddd437fbcdcd67b8f8bdbf2d75b313fc6f870f0
ze0997e20913dbd4f26c9a3db5c09d39d07a666a6f1b729cbc7267f1109ec53bd463cebea9679a7
zeeefba382428d2e23d1aab70a1da68896a770c47c42e3ad324fcb796563c3a7af0b8988a32a750
z24a5aa7c5f71ea87663f27958b406e29cb3919d1ef4d0f7e84e3ba08e457295c2e9f1ab514be78
z3d2e1a0572a6d706650a3c15290ac0f5b4126f237f9268237ba083152c7ee4f6819b902b1256e7
z1a8e8fd2f5bc9b679b6be43c6897b2dfc7b8aab61e6c1b1f6bb14761ed91cb86dca5b50a757311
zcba449199487514da1fc6dde6adb78942be3d2445340d854ac406ee42becb9301535eed86949a8
z3483dbb8260ecc4087c0f2aa8960de068bd992598b95bfd2ef379ee0da01549e805520c2d35c77
z4d35263f0e29cb46c99a547f6007e561b2a1ba51f3e155c4c03b9e73113847a9f86029d857960b
ze347b3da4d611a8bcc31efb1ef267bd8e51beb027b0fcd6559c43847f9630b2b007cfbc3e68fef
z916691f6316ba706684bbc1bfbe1021c836d34197fc5095ff3d665635bdd233c48073551b1e242
z1940787291d2bf54effe6ea9a812eb52fa692562d594fc75431e0d4856ef7ee8604ff1476e967f
zf06593c6f6a66baec277cdb362a268e29260a6c2694fc89e07dffb0b55eafe39283bd926238a90
z581d6f3533ef78399aff4cafd003555ab4b9d6dfa7fae89009e14dd13f06bab3b829ca003f5e16
z7d220c96154e55337df755108343f2b5c76c3c5c3824e478961515fcc74e43bff464763cc0027e
zb256a99014b5c4bd9351b51f49067f27f1a169efda283aeeeddabde8a3d2e212701f6407060df6
zf1ff05d28d290a69ed7c67f76abce2e3aba361e0dda3f1e5bf00ef7f7d4954273d02317cc0156b
z72d18535cf8973da6f80600dbe7a05ed78dbb0721671518dcc9c0760d1baa6f4d05a9466504d14
zb39b7fcd9c1f28bec57ee1b353a0c51b77a3e2574b7ea29e7739d55b6be9fb8f8d8d74ff3b7285
z9f1f628a6878d875d85bf07ae0f039cfa1d9123d227d7d556dc5b0492caa84128461541feb086c
zc16f9bd20372ce2b8bc91e9ab56eeae7181fac88396816c99514f18c0f98e5447127c8bcbd556c
z92264363129a56ed737f0e6269b61f8d514fcb2e1cf51910eaf6ea331801c335c3f94b4409811a
z8bfc8e0e2b6e0a69d6a694a798feb4dcdb7466411e402e4f2faeca561037bd91160479aef1d2c2
z59410234e7f8240dab7d4e078ef7f765027f2eb99c4bc037ac1517204261a4481968580ce475f3
z47fee4b4f2fcf24885d985e680693abba1bf5a4b3de007fe02a9d398c0ffdc4979eeb004e139b4
z76d3e18625f62e103c0513711f267be9dbf5bea4ccc233ad7374c5d1d002836cc9a83945baafcc
zf2a06034f3a66ca78a4f3af6d7c1325b99eb58b82ed84a169d1d88cd6f1639047f00b4545a4d78
zcfa422f22fc0ae77f822f86c7c492297ea49dead9692e61911959347d45580d4a719c9d06f29d1
z519541b2f42f39e52cf0c42d18f63be2af118089ee037ef077a305fee961e422e3e7947c154444
zaa679bad6db12ee11e9d0e289c67f2b37857cc80914da7b04f4d9ea1c810b6d517c3b87e3a3b16
z93606ca2fb9308f58ef3081c16301ca0c19a7ffeb871cfbac98b190a79fa3ce2bfd82266c26c08
zd004bea7fd9db09054bf4e538f2c5d6742f0d245ff45650bef794dfaf4d8ab6cdcc2682d7ead0c
z528279ac07c9fc574ee73acb445bcb7c5ef560e04d60886c1c76fb63b75262ee304c81d4626f72
z656559e705478aac095fc321df6ad51e525a087bfcc06878048f0cf87efd322ddeed9aa9f07a10
ze560e7b15c6bdf9b5bd46c8cc5e69f32b98aabcd0ed36663d9f3f8d4a0b8118ca7b81aa0465ffa
z5518960d1eafffff2b7b71a21561318c01a328ce7d92c35a55f192c90f3d0c8bb85bf01701f5a3
z8a510a94290959c94129453221756278a55ebd8ea37e6cd02f294a286899231bb709a2c4574e40
z439b18cf7d9a06012b597275543fcc4810c528f6f3a48e5a2935831fb5e314f7c24e7df44f8399
z5368603233849b1a44db747060d8951edcfa82f5b3a30ebf6bb1f7f452efe38c3dfc5e3cc8c162
z877a9a1a3bb13b966aa65adad00995952952aaa0d9e4f8c793f3bd5c7834af43204d38bfa67c81
z4b66846249a8b49404149510dc0ec9ec8e6fb3114cd8e53d4fe052354e1de11184de131a6be766
z70b1d982de66e3bdbbf7d132f30502d1105705c5fee77c987ef314e01cd2b9c6649439fabc2962
z04d0dd1dc30de4a076f5b5d9e8efd80cebaed07b447b58f0669234650570a2deb4fbc5b32ce76d
z849820cc3b4542c0e4cfbe049d457732f673ebf3d0b4f59d94ae93f09643abedc29147e29a1b21
z6f5a09f32e83ff72fcb628775806e9b34655b9a737bc043269301bc1a5061c01ae05d9df7bb84a
za382a0b088ecd04917c11c1e6c1af2021c6e14e0205044e5af4505ed7ddb02a96c63e33614b546
zb4594c3d86830743e8823c743eb5ea007a0496a540a1c3629f74f23402d76f14a393fdc90f477e
z8a0ac4e15be71cf310084ca569c16366c979bc1ad19999e5846e9b5ad9ae998ca2b4168203725b
z7983c07289f3b5cc9c8c885478afbeccc4ca8f4e8cbeb76279ac27eda73c7462f7a6cfc7f7f2af
zb7c3d3226275c13b65c89caffdd0cae6210e2a48c54aa89f131b633946204d8b9e13a75443472a
z893a1f1f6b34dc8edc0cff3650c91a72e738670946c11cabba7590a3eecbb41169eb1f85498d84
zad16d7877027862aac9a3becc651db1959ac8b39282a6c997c2b6cd2504ca7999451ef54965ba5
z1a11a40946917640195c42cadad2befc386bd727556cf5fef07ab4afd0a6653296031eb0d95711
z2b1903ea1b99baafe2a8f725d9ad9a44d4d310c5e24159a74226137a2ff2122b6b7b7cc33dbe85
zaade2fa4f4d4d97815bd2ee54cafdfe476f63f740f8c5d6c67253fcf55378f5b7c3328d68bfacb
z0cc8349c246ce08f23dcfb059eddbd23aa2606b61d585edc8367345d1a5a96b28405b20401755b
z24cf11d014b9aa06713721d8d599634b5a0fcd71037edfd88d70f0a5f5a4a4b5db2ceec0c1adc1
z9b2f12cc8f2f6d962f03c999273e251ef5b6bef0e3ff9144999ada880e480ca91e5341c0965720
z569726712edbab54190fc9d44d4103bca423ae49f39ebedaf9426dbcdd8b958f0801388f1e83f4
za38859a787d6e080888d0e6b824000c56bd6b8e628ef95a18b272cc809e9a4e4ce14ab8f16a57f
zb26b1a4b6318683696a362409fb413fe5ca09a87546450584180dcc2eac68eca4125d238f5efe5
za910af52f42e07fed1cbfb7345b7957cab4d81dc48af0f7a60d1c575dccb72c9126ca274dbb7cf
z17714bb318be0f3bfb2418d2dcf3d3fa2129e7dbe59d4c31f0c759b2262be58762a239e0acdcac
z370b4b3397187f1b2166e6594edfcdc479adb5f298c809a3070fb2d40c62b89977be692292dfe9
zc56c7562aebf9200219a3aee981eb94daed05ae9dd904ff966d5a33472bedc70bd80b9b087acd9
z97013c67e823e253c6b5d92b078f18deb218b4c315a463ad7b39b362815e220fa0c916cd14b956
z1fd0031063fbf9a7cf3403046279dfc22bd3fdb258f0d372eaf244da3c2885fb49040489db43f1
z8778b8bbafb7dd685881cae347336ec3f45957cdab5b7158f7e9e9df67dc649e248dcd23ef973e
zacbd7092336e472bcdd4cf621ba7c2e7a1b5bfe01c23f82079864e6d0a9f3459adce8d8246ad49
z78f46f5f3fb85cb541a6518854109022e446bfc153b4885dca1b23f7b7d000c8ad2ca63355c631
z1d1c469c22c2caca20f42d4f827a0824f9b58fe0b93002c04f99e1cb3e2859eff6bdb9647ac741
z592bfec26bbe700336a7ca76259deeccb1b0ab7791fcc24fd671b03d62bb923a2198abddeae0c2
z1a0b050af54dceab01a7ce52f1b4971ae04f64f460ad4123d52181f6255cddf11eef2ca09617fa
zae8c8a2a9eab06d2319c7351abd755212872c5b5b9d41088bbdf9d5d4ea81300b82f4ac1d0ebf2
za7c396bc72c3ef9b96ae668fdeb04cbaf181728b3136b62972333f628d80dde7aaad2ac878c336
z78d6541c097c6a88f6de7346c636223a6a7efdcb6d18a4dc6225846d8005e69fd2798eaee62f8d
z5217a861764b51b716e31433c3b0bdf503087c3eb6aa0f9f093f07e86557376825054e0eaf4f22
z9407575103a297ded48304ff4af4ef269f264a460fd750de8e73ccde14561b2311e29f4f0d8c76
ze781cc11c913f0cdf77af83239fc05de5c80349b7741d93680b57350f0d6c184ed16b97d1cc810
za287ef2e08356a5bba2f0f7946133ce8fd895614cf5a651abb73ca97b988a8df44ca3c6add2282
z96e30a4e17d4e10b4d85627c0e5a3a7ba392c748800218382b40ad2f8a9ba9837cccfe8846bfaf
z86c5d8638434d49f76c4b54b2ac5c4203c95a33c979b767e8e27c8287ad68c04bcf8bed55679e2
z1011bee9b75311c3c0e9ea086e47f1a6c1db965ea35e3c7449d0405b5cac4737ecee4a2f001ccf
z828db2358f6e6b175b7ffa9582ba27d59488e07837b6630c435cff3cf06225f79826202289c661
z0b3b716b3bbdd6150245894a35313976d1ae7dd0a6a2b4bab2423b02740bfcf01214d1d90b5b1e
z3a49d92bb5e1a26c5348235ec4cee3a6d8c2008f162598c49bf941a8e440e45dcc0458826c3baa
zbf9327c0c38c9bb31d050a4a501ae0369028bbe59f4e0d976f674ce31a8e06bd4e441d8ba7654f
z2317b582f5da7da3c7e6312481590530e829ba1ead2691db8f936f646238b5523791db5160b83c
z164604213edbc28627d15fa2646362d3215a8351287facf4b8e9d7efccd5d019f48f8c44900444
z09047362fc77d0c67dfe1d5c65281d4fd05d5a02bd99cedcab577624ff0e68e9519f3882f5b47a
z3b07fed3900dc89b04e6c27b96908b57b5d5c5d40b7ef1882301224b4e57ecaee8353cdc80b7b5
z967b8c5e430dd22f3a773a612b430dbd09f7b396283088807e172dc936ae324ad48962456274e5
z30f405c53e1316fcdf7ef342014d780e9b75c68d1f647709a23f79028830c882fd52c6e393bf29
z42f2ea5dca8dfa0d3215eebd9d54e483d096766582903ec7c1a1f5e37dad95aca75cc6b042e55c
z935c07cc959af4c805144b14378a83950b6f85c1ec603791ecca41d08429a26571b1102db5a74b
z0607edffc2cdd83247179daee6c7e4430a90d591074943844283993c349b4fdcfd133b50733bde
z3e5e5f81389e7dc4f9b04b89549314d783aae81c18d444907a08c6e4e1d87915c0c7375b7b5ac5
z59ff1c46820f79cb861fbcb23399aa96e33804448dc45515d6f63c39f793101b2f1057469fe107
za2d325fb81e8c2d8f612b6f9353f07038b70085ab81e1926e12571401705c248d558723b7863d3
z2ef388c58c36c318763b4ae9077119f5533082026a00e7f316d6c64f64d001606b421177a51b7c
z23003ab333a97731b81ecf9a6e880cea931a6e4b82ae41345dc8e050fc6cbd9f4a92e0465653cc
z559d614a5c4819a69080813434b7b1e6e56b645781257ce2db91492a70edf9d2af866aefd0536f
z2d16c53260083ccb5ff33cd639bd4fa2ffa68626e3d381d37f0d5607e0d764f89718454bdb08f5
z97c2d65f4af714c0760839f9fdca62566d05e2179fdc5a670359fe7abe58901c6f8673a764d710
z1e9ffa253fa592e2ed2806caa50cbff304c9ad640a702103f90d432d5fd1a888ab52ceff175c24
z5222ce04d46f8ce68c40d76c53232af99ba02cd8f89f330fb3db8a823283043e651a1ba81ef821
zf02758a5a5e38b30448c0a28dafd6e8a5a4003206b3f23082fcc5be0e6f31a2d550c8a84eb5e4a
z80f4e91b119890df34359f00d9654954128fe931c0a2d84fdfe38fccd33d3aa3ddfaa620b5372e
z0d9fd6b11dde48773ed62162ccb58e0ee8543eb6e48b9ba626c3c2a0976704b0e9b88ff28d1477
z9f60668f8a2f60e902f99707ce58ba3f3044f360f79184b69de678287d156d0f06379b6ee5d944
z57db0e7ce8d0739c586c67ecf869519bebc050e22774328b02cc7d2d8fa4b9783fd6005ba23d90
z80418511f3bbc65cebd91136d682b8463f6b546c029d99558bf9b5bd79df586da7c933c8d46317
zbe3d38c0ee12e1e665b763936fa35cca8857e4194823803943d791d5857a0d65f6c3c92a57c9d4
z736d13219950f34ab5e75b9cbc3b92371583420119c56aa071a083d329b2d959bea0590668dd73
zd9f66ae1592622a3aed6d158cd487ab692671a8f71e4c97fce9080f15d7e35a2994b38b5967f18
ze0d21d12c610e8462973f0adbcdeb369b5fb170fdcb1b7635a3dd9e7659d58958743643aa173f2
z77ccb31db1b82bc16a3451a112f4318c61df722bdf4aef4e2cd1a050510d0df8862cd13f8c86e4
zc98705518259a71bd605de7f2615e153346a8e8322b4d31c685d3bd57ad38d8474222d9ddfa2d6
za8100175d9878026119e8a92877b83ce0395abada3835bd56fa2ced8324cc6d0afaa442ad5b9f3
z519f14df9e67428bc97898e90123e1ced92d379f6ee005a1f273928dacb7a0dd093f8a6bb92d40
z528cccdd93dda1afc4c94b31a86847a5da656e4564188b7a4025983b089409d3b98cca23cbc7ed
z316002399e61b54f6a8b747948bab85b0736fe6910816b2d6d31447b91558b71f8f2e24277e680
z65e95f61a25cea53c6fc8a19fb89d89150d55c10503d76c102ee9f464e46404d1ea5f529b98c15
zca3e54d2b1ef7e9fe65e9d19de247cc03c1d0d0cfe658138479c6376a1bae854622f996020aa6c
zb4381847475c2f1a4eb11b42720d4ba0d76eae3740e82a9ab42bd03ec53788caed79e26b873665
zcfa381f1c975363ce496c20c77766c8ff31535b08a780eb10cbd2a8d57019539064fc08a902a7d
z222441d1401db95404819465bfa4ecb5fdeb991282da97ca6f829b11b53e5da34edb41307ccdc6
z862735dda2920c42ad2fa4fe42425adfadc54acc8c06684e8e1821c3ff3e39c0e129d81706cdb4
z03160e50343f94d94db062a656b29bf0f3e85b9e0c38bf0d2455921cde8571515ba646d94070d0
z37b4792440a2ee36ac7d6723f49d9d731dd437c771414473a25f394ce48cd9c28b8934a9eb553e
z494d003a7b9765ca1e3d8bfc92522dac6f7dd503773d9d9a49228683a229c3511e77dc0b8d0cbc
zecb5639387622a14615ac249d9004f1a3f22c9179ded3400b7b02d950382a09e09bb9203e4e140
zd4c9e9e3803829d93f5c029108170c6eb081af2d9bccded298ca0f1fd0806e2e4c6f69be30c219
z37409d1a65989d5f87f8069aeb1e6efeff7abc93bd79a85c5cbdb7068ee50f1338f13959dc6ddd
z090abb150315ae31471e939b3f37133f74ba76a85d4d35119d430a47affab8139c1d0344800a17
z8f864377bf66d50af1002c9d8d728b3135ec72cb525d17f6eda06106b84d69175e4531088ebf46
zd7416192f68427acf142a0916bc063b5bf00c317d3bbacf11bc745b2795f1e20595503f6851198
z343e8e7643fd4b54f72d9bba8dcd4638cbb7a672147c5af73e349c2ed4b6fae64cf635f7c94514
z3f1d3438b9801cf3659accde4d3da8a410a383ed669f517af1ab7da38d72478e9bdf75b8b97816
z4be13f1465ce102a53d1759b5421ce6046e41d98a32bcac6b2454b826c8924697bd2ad99253b64
z4dc7602f00bb1136198bd0c04f0447444d2665ba8ad7d1b0aa2b216d11b15296fbc0c82126d0b0
ze66ab3fa1d817ab59c86b8edfa9857d866939d3d9427cc69dd00f717d2dc3694ef8666792106a7
z51775bd82f8e83f913f4d4395e505ff31136170d0e0cf5c691609205c7cff5487fe88afce1fb8a
zc6336aaf653ccb64dad61d27096a74ed03f3501fa0bb875f0aa8bb5e041cfb0bbda56285cdfa6a
z6c9c694f3f910240b554a5c1dcdc0b71a1956159d721effc2d756585474021c9b1bce52cde91a1
z936d6d6e6d6d4fecb8c9015e07abe1326deb1841b2accaad98e585000a1693ba9d0cece147a62b
z76cb18f975ad69ce66e398004b7a58aad313bd3e20e8338207f0dbb0b62bd721e656c923bab21d
z43bba3b1d8e9a441cd96887b2a4defd136fc229bb69e764ba7042ce853c7b2f075ab32f11e5667
z29feddcf46d918b4bfacf216044273b5ae3904b0d4546797a2778726cf2ae50e3e1d53bca361d4
z292dd634a72b1097dbfb2ea387365bf6ed3421b1f7d767be49bd17cb92b43b30bc5be891b1948f
za338e49fd148791c3a267f01556ef01fce40d400737fcca038b3e52cafb125f336f110bc217ba7
z1fb5f6f2073e1f18ee11b99a6ff5de1300559e2f4d2bd5de97a28934bc72116cb35a0b58be20f2
ze78d7154121fd7284b048389d9a1c24ae4beb2f88fb28f4e9ee81c091fdf0ccd5917b797ec4180
z059884959cb6418226667c39be36af1d86648a502796146f966753d0a006d217ecc7ef653ab6ed
z64798bc59273816cf1c24f1e3f8ca0049b0f3fb43ac82b9be45f1eb8928788e648147744d5a331
z8312394ea161b7a3eeaac0c5752ac8b4f0230d6c6654565618b3f83fd74c824e7f32f19c87307a
z5a9decc6f9797097dcdedff02d82fa1b1cc7cad153c54ed53322cf143e8a0d3213ba39e7f704a9
zd3b7be07a16b310b60526f49e0c910ad5c9faa1f05d284f2b5a996c40900d59564604721f454f4
zfbbf0d25b000c0334471a95172583ae130a467c55374735548b6df7b30c9be1d32f8172c24b609
zedbf5bd50bb441e68b67bd1c6f97b1e1d3133b720fcb65e3a74eeae1e1c9b40fcc6ec8137ec8c1
z80a68f4b38e6f503ca783e8b10d9261d3340848823fc3bbb77eede60ebbac53748e855c432c895
z25c35f6b08ebe631cb5acd339fb23bd889a008b5244519f188c34bbc7b16ce3631b9d8f1004a3a
z67748e583034dae47d8b5082abd85c209109560ccd7c9cc5058c78304b7bc02bd7fc427568ea98
z0fcc41296157f8cd3b20fab61eb4f51af7ba05bc7cc64e62255f08fd3f8ff9841b3dec9fd2843b
z7ce5840e500f7465e40a3de2fd6ee2df4dbb3a2ef5f39068745c0dbad2b1a08ff5bacc06a10f0c
zfc2af59c73d5afe5b8907dd9311fa1cec6c39826b5bbc754b9e272766fb8612a188883923f6e1d
z20fbeffa1d45cdebfa13c2afbac8bcf54a35aa1d069f906abd96ddbe6cd292e52a83903f6a8604
z2a6d6670832511aba4e6b11b35e04fc2e53681b6ddf1dc3df3925510ed8b681162c327eb3eada1
z9fa094e2998291bd5ac6176b89bd76bd1a5b5bc5f7d9882cf77eeffa054bd7b3d188f4630ee410
z0ab1d7e74f5c76ccc79ba44896d01b5ba6e8f36d8b3bf4d2e7645b1ff48880ae8af794d669ab5a
zd9c4451cff4f47d247733d472fa9d84cd65fd434aaba0fe03af987f2eb7f7c6b68139c29aa54e2
z77197519aba052c98bd5e2f8c04c6561748866ef58835139a578424c0fc0f742466aeda32fd130
zb4f920e5377c801086c6ea36b2851ff988faf352f35cfa16b8d888e4597c33bcbb0997a9e7418d
zc270f22e50a63d9d57c0838bec1a5d66c8ed45025449f76ce049e4aa4404d5b0ab4a283cbe9445
z6fcdb91e1d1a9a348fd86944d51250cd284c593c2a00380f9f27c8bdaa95037b62470a37d0289d
zf8838de62d26e89292a20830637288925b71c425796fcd9ed34219ce1c8dc231f787667783a088
zff1cb844fa93aede3725d22faf02840c5db65a03fa88cef3bf9bb0ccd7db47ada53c820b151572
zff4e8e19fa0dabcabd8803d03823cf0a6ecdaf61eb52045f0c117cefb27769a03d6cbeea0166a2
zc85ff74d9700521502b27a1fb3fb9b42a9aa0f7fee1227c7fa839fa2b87dc6dd801901a2c390ab
z41e85dc958948b68ea2c90aee5cb1f438c8e0d97b72d66c589c46859c9128403925b7d1cea657a
zbe48d331532b2f7f6c5b885d3461fc5c72b4409beb8acec6c0de662bddc277858adba28d914763
z04823f0ebc3e724a03d4714c156bf587f020baa9717a4157b7881cf9614853c6c3178d30f45f50
zb34102d18d218a1b1469826f0d230283e92d839f5250ee0640f4b7ad66b90fdd9e99efaf45b6e0
za3197f84f1bfc933a3cb919fe153555f2959a673f656ae0bf4939479fdebd4bff0c7e1fdcaf950
z68452d8f486d43385bf4b9c9f4c6bf88a7c5db34410e24cb90a4ad310c3c07cd17e5dfdba4236b
za866de3912d07259df72f92fc58505a04e46aa6aa2774b7076cc8cadc9692a22d69549f8839351
z7562490311d061ac48f7e79bba8c748c66b2ea10e113a22dba46f3544a2f9c9d07c36d9666b014
z8a941b3251904ca4d23ab370827e928e76e3a5d41846c485ee3753e361a8ff654c7499866e5f02
z7eab2533d4105fe2d3eeb341b0eb490ad4a32c620c4f0240a954d9763f3abf458b99764eac5975
z32884529bdc2ebe046675c505635efbb1382e8e64f3699f5ea64fdd104f6f2abd25b1a5159e3df
z1fd1a43d7330cd81030a7645c21de0920ccec51c52e482bfa710437d12349c448aabe32a163528
za7a052d95956ef761ac7e4c97f81352ec7b217ee59daf5fe80b0af86ff00677efc5a827ac6fa7b
zc9e6eed047fd6a7ca82ad8accca4d33180a15e9bcf210e912a6bcf17a49cd9acc16eaae5961fe9
zb7082e702ce880ac2d71f15c6d28e45260e00f16e0b997b440f7c94675d1264d298379bfb31cd3
z15b88064548ff40ccc2176eb9649c79b1fca1343a451645de114698a130254d30c37d2f64ab6f9
z0d1ca675871008f2eab6d008ac3bc3bd42e929cca3ba6d89d0e0f0bcae0b304e0f71dcff5e49e3
z057bcc3b08315d16d6fe42a4c25075b3dd30fecab9f924f27e78a1af9acfcf36d930b632d6ce6f
zccfb337b920c111920f114b9144ee6a72f12424c94ac447c5e9069edc40f80734300e600f4e4ae
za418058030865e80fde0ac6806097335a5949c1096958a8eef71a83d32b2c63e8d566c168106fd
z9ae6abda214313af59ecaca26da9c1e9b7b9fcc192e1fef52e96c4888b267d88558b8f6e7b13ec
zc0f51ddff1769e2600ccc969616e3afe3ef3cb0e559f8f3cbc582d1274391a123f07c2ecbce1e3
z6e9228681aa86368e8672ebb4acd7e23266c45bde5f9fc05ba90a15680b41c792c248ce85dfd37
za5eb28899200e054489b6c4a75ae9fcff5373bdc55e5309eff72bc986e5144a1b8e15099bf1cbb
z71ed77d9219d7cae8d078e7e4e6a27b21f20cf639d1fa253d5ec18c983d5d189048ad9c4d95458
z3690b34f14062235986de8667d82d30ef098518203ba6fe9f171674eac30443a39a5a7ab9fa605
za2595e5e188ffc4c179de391a79585710b11af960361e305faae572e464bb4576b0a971edfbebe
zb319d0d9bc5f32581d33249b346ef7773f523def80eb85f7a0df1c8f4f0fdd74d43cc5b534df33
z28c01b951c02bc5455a0b083ac67751725b91804a37d7b540e876a14e0f5ac8fef72b157f3fd1f
z02912d2637391e6b234244d19258bc52d7f36467d53b15935500ca4a4261ae7c55e9bdc48668d9
z3112af68028803a1612bc4b436429551b359797036cc2e55116bb4edcc6b2d9b9547f068834fa6
z8f9e58991e88a9097b0fe717f0713d24688027752fc10fdb5d56a20efee8ec3e59174fe1fe264e
za8e7c61924fc8d49b4890e54c68071c7a04d046535e2faa237f453ca7a22022425451b5ca32431
z2685b46a9ea59804c3ac5ebda37e40f27c8d95a1ffc0ccbc1a14d038eb300f6bdd12124960ea8e
z9692ff414f8518087527b458d0b78c4bb603abd8dcc91cdc5e033f88caa9a1e6b487bd01c4150b
z5f5c081cbd1d7e9ea705cdb08301c800b74f711f473c9f271f63c2ffa2d2b6845123e63ee717d8
z32e5bc407fd0a77b0022336a48eded37944f0fa0425a948a3198c419bf1b5c8946bbc712e36616
zf54f665d4254305f6eb00fed7b93b862304f2476c11d58f75f91d3387fb75d477edb714ed4e2d7
z9db13d5125288fae49ceb57b04ecbe34275256b7cc86436da7cc51d74263915ed0962f85b8712e
z3e10c8e5572bc9c2b59c79e48c5c629793a1c23509df38afb54c8e0ba8245ea255324b424c8063
z127e8dde27a557436ddba6a9a1e75efc3f154af7c26589554a19d793223ba993fb17b3e562a0c6
z5164240e1d483670d86cf94c623211a040ad1062c5066beb2e6cfd4933d210ae282285fbb247c8
z5cc889ff52bf6c8f892cbba7cf9706052385b2e15c3187369124e14c076b451f7b3d9f7c5718bb
zc2104a07d0b2863e6f6892433b1e5aae2fc134b027cffbfe9fff6c2b1e6030b544365d8df40f61
z8dba1a672e000f07a5992dadc3b54ae7dece30b4714b59f94e67a1d1097382554db459b4bcc79c
zd2e7d497b682b57c2ba16530a389d794ef5957eeafaffbc63afe1ff340ec1ad49a5e68186c4037
z522d20df64cc3d9646f738f378ce3e1231155d365752716b1974f1566371af8912d52184bb7e58
z3fe47143fc5e5c7cc347fa804248e213b6770fce9aa0e935308662439ba59e9093212beb24eb51
ze23613436ccc97331c20e8693a8aa07a4a4137196766b0bfe67841cb7346d5e962c3bfa7cb0e0d
za9f0e651a2e3caa473059186231a93fbec9dd618e594f9a1199a71b3018d73bdf53b77d1e739e6
z171e06c3f9e0f188ad88ff3fa2227c63d5a73349c5c16b429d05180f66dcc40e62f288b97ae556
z620ef94b9a4c1dec5768abf9bfce4640f75d4c2b6c4c8df9253482bb5841b6a705f60a5dd560d6
z60469f393950137ea0b286380221f778591ee4c74765217ea08929c93133900e4e868857050fae
z4ecdde5b01e3a21794f481d94b45d4c520e67819becb78c3aa41cd2064e7f206631a432d847bff
z37f509460a2e7e9ad927e2ffa644d311cac0fca0a9571bb55e8744a7cba68878d594b4eabdd96a
zdfd5377797eae1420165ad966cad6ecbc04b5a3b06bc797d5d646c0170d837463d18dcad75596e
z684864bbeb3fcbbfb9be9f37e1c12704e78af99c109f249dfafbe8ba1360938eaae400636fcea3
zc475c8c1dca69fdce3123f12495a3a7c3387eb8ee14c9aadf7e506bc6d4de21edca35c24130635
zf02cc9c2d54fc7866ea7c3a3183c6f70d06e092c68e057754f2328a4f9ff3893af69a5f30d31c4
za475f611ac964a9729381be7d34a34d8a88b8586323752e12daf7c2b9bafd0d490e30f975dcacc
zd18009b6c898361e5c9b8124c32c1eab62c38f78d25bd65f58ab39b26f42beb718e317620d13e0
zc86d93b9411953dec3f9bfce6defec28f0505266ca32cf1e84d592d135447c0078bdcf560699fc
zf2b937b92b6f332a5242d163f134f065c604f92d81351a2f46626ae25de13b3493240d15405200
z880bba967813a8cd2e693994798ea52a0a1b1614b382c9a66662b2d936fdfd3f7fab4f7cbd6d37
zf5548c84cc7a7e67c16af2679f9f3abcc68444d96c2d278cd8e0c8fc0159e625a431f8aa75f097
z57f5c3fe7bddffe8ff3ac67e0fa7e31530017d0d341c87cff048deff489f23c72d412a7e0569be
z57999e9c3ab314e04a3a1c74e1ae6979ad3615bbd7430446471586970a83a684efeabdd14d0b0b
z2300adf377b8108db2999211e2e5e34323ef69802baf0e0b6a27f28f4aed001f3e4ef1b7e1ad5f
z3e6398b599cda3a08585bc3a22574e49c06bb613914f563ab4eb4affbda9d1a6bb15126e9bedca
zde36af0f23503425d87f1fddab50033f5bca5accfec7ef7240f39be2f45fcc22d6d8ddf0a36c63
z77c372aad696bd8b58c15ad40f03a40b9c1673031aa9c2b68063c20f00501aeddeb6582a806e40
zff58915f8cfe4a41194b1701d3f03d5758d88323a78da3b6b3c6410ab1162024b7c5dffc8e2f2c
zf1e7cb045481a8567d24c0d5a4f4c9ff2f35bde7a7d843f3a304c197f8bd05714a0112b5b210b4
z78fa2ea07f79a081fd61ecd501e3b2e645585dfba5b229cddab54f5642ac9af64d7248eaf856e1
z745432ec870cccec49555ac46e0560facbaac2f57673a52f60593ea9c3f6bbeb4bd1990a2446ed
z4544ba0830aeb7f7eb955d5c874f402202808c5edd479212e25c56bf34c56777c91aee42ede2db
z1c262647654dc4b78aef37d3c6303bb18a89843ee148b2dec35c151161f0fa47c835d155f15c1e
zca6cace59bc6caf9b68996c004230ad3e25c0eb19cf62b06adbc039e0b8a7bf25d99a3515ea9ca
z01e827695088370e8729b6b802d396a5fd7a44b7b67754263702555e4c1e164efdf43a31cc5442
z159cca8c42779246a3022afd5e8ed64aa7e5a1f2a6167b09584f714f792e361b5ed1fedeb7f8d0
z6c2963e72603f3ff1e00a51c56f1e80c14fdf44b68045b79e55a339268e9c526f8da853390eaf9
z1daa07e442a481ae9eb264db8a931e6bd1527239e3484522ed84e5084de5b7c72866269ee21820
z6740491bb10b3c81b0d3b11ee2b9acccb4ef2a35a432b141272aa569a44171d94f79bcf550529a
zdd4c9e195b8f690be85c32435563f0b06fafcfdf1eb64e80bd6034084d79daa472219eee84cd78
z7c1b8bab4868e335621a20c4d8e3511dc5a9be292fb322ca36a5538d06b9646a7f552ca688c709
z57ca736098cb262e6eba51a384340b015931af4176e7a694bb0891555fb19e57887bd84cfafdef
z8449db523b39bbb7fee2494c4b8578339d3ac25af9e25680bc84f071c47b7288cd7483e26dcab0
zfb2b27e569a870f954d1afdf4cf0d3c5450a3977ebf365fc7fd58f5cbec9cad30c76b0372e1947
z01774071fbf440ad07c77c63a2f1b3fa65312d02c72d48c020b34b6f892815c239757b9fec5a58
z9db30bb5d08979789191745efa837a8581499425bd112d6fe260a4ffcdd0502b708f9fe649633d
z5c9379267de0f89dbc1cd31fe7652a51e1b58d9558e8fdf07a469a34ee689654237e977130fa6a
zb255af1d5415981ddd77cc0332917a5c531fa628a13d61556f3535512627f53d32a5922aae75a5
zb3f86a813ce08fe12fa204c1ecbfc2925fafc58526dd1908f8e5556ff4e198cf4849f8eb6c187b
zd6c287812da0109d5fc41c513073e1cec0e60c1e8d0799a43e34b29e3abdd7a0b182fc3919e018
zc0281fe5e1ffb474a041b395e4ffa37bde605bf1c14b9b15b61936f4fd4f9177492adeb06e79c1
zb4a047d0e5575e32cc01f715f28af58aba58a7e8d491eff8e8bed7c9a5d25322458ee1357b1b3c
z075ccac7ef19b7aa144a2cc9424c8dbd01c83ae73f81174b7c2714be06abd89d8a34ed0a827a82
z8d5f3a979ce8fece38642895ade51a2f4ff292ca0f1c4b23ff7ca94681a52fbd36691ef42d7aed
z4086fb38f08c55519a3f247b947fa2b523488b65bb09dd8ab0ae5e3eda62b3301a4917944a4c96
z0b9104f2eb80e9b59a2fcc695b701d191f96f2d4876c3cd8657774cd740369f20f47aaa67b07cf
z67331dc1da54c18631dae43646ae98a7bb0b116cf7adf1e3f28089e9051b4adea0a3e7be91cbc6
z0520afcf5c3a1f4b16e2f2c678c088e60d58e8704dfb9fbb350d238fbf8531722090b944d937e6
za3f4235ef4e0ff4e9f09b335764271c68c16755b5637cf2b2a4858c7780ede5eff2cd039f8e80f
z01b8eaa097cf4ed56f2ba8fde64264b8f55e39c1d428c1b67346ce8ebceb098c74f884a55a58f1
z597187da9abe86cda8561fffaa31050221f819d7cdcb675e1c2ccd12c13befa7c6158419a7c5ae
zf7634ed545d3757b4954dfbe198a08b2a26b56405593abc1e5bdc9716c2eb3f40e12be562d334b
zef4be33ea5582057414f6c3d330d85e321abb6ea2c6f22ad0f26a418f506d491ad2912bd1e4430
zd572832abecf50e26fe78ed503f306f8e114503b01ec41e9c6e08c2074c6b367c93d6cf1e8ad35
z10faa6e678302f3dfde92fe9bd1f283f57584ac63250657818bc0b377174b994ad57b0bde0fe84
z99142fcc1a804a66441d1f2d01e91a81875264452e70ed0bf73e6733685ea189375d9fa7964afe
z0ec7c69b1fd9b9c02d90818060946331740078c1e03852912b2d23cb74e8638b2453cacded3d5f
z4627786078d5667ea67ae947ee77c7f2c405269caa47bdae2f2080d9ae58fd6228925a605a5053
z490bb8fe688cc2fdb3a3e2dd86ce235b16c83dc8aa60e23c18ef76b21f80bd90847c705240612b
z2fe234e6706fc0977644da958007389fd348645c330887668da52d790a5cf35e40417f173b7315
zfb490214d4d6043bf7b3ab0fbff0552613568749625bfac60d65c0ed64892c57cfefbc4be9cb2d
zd90f2108f23ec10b9dd0440d17715dfa06a959b5e35a103fd54559e904e15e0d68f96188666759
zb9a48a26852b8edb4f0e61ae75d93eff58376997408ad0bd7beae382af7b932a5397e1b8e1432f
zb40fc36c14b4c63b7b38c1c31c9f425be203094ada75437a8a950c186c8d7c318044188b9d8749
z86a8607ed46a0565e91c83baf29a2bb4c4c1a03517b0bc4e767a5d470bbc18cdde94ad50c517ef
zbe2006ea0cd0a4c9221e48b06472559d47afc2118af41aacbb0da4ef66c589c5835d27b9dce92e
z6b613999b1813cb232f18b1f9f2cc3370340ff64d6be3a8ad028215fd148456bb545f6f3650b9c
z9c5dbbd37139664163f8283a7808da99f4c3aac23fbe7d0b8f2ab7dc4e570efb861e32b0e2165f
z40f4d5518782a3be390b64faac70ec136931a12155a4400c98466118d7ea2723e535ca375b7c16
zbd8a868aaf6a3cb5e4c7163e605c3dc4fa9254db30f3090e24d7631e03bf0bb2b96dc5d3250670
zdefd0bb0524fee4c6a811b7c5dc7a40f34bbe5d39f238511349ed7e5138feab22599f792b0e1e8
zd1d5f28480f47ce2193ed1926d16a129c6e0b8769795dbf37249ec72b8d4efb0a1376b70e58b49
z0ae362b55067c7fe2bf1baff4d209dc1a0321cce906639d20cc98ee838bdc13d4597b0cab87e28
z27de62b8e12468e5ab3313e85bbf322ef41d1e06991b550b5b372036726e63f3eead5d09528535
zf270374bf8ae422947e56fc7f7434304d5a0c7be24bbee73b31f130828f2c12f6e70c448d0ce4e
zc0692f6cc361cbb0a7034608b58b6838d84fca79eec8f2a447904e8fb2e40a975885118b2a8bec
zb83c5efcea7230bac3247de3d4ef22b6cbe1e951f51398a4030606cd3556aa592dfc1b4cc6dc71
z3f8dea426afbf665df99b5954bde7fe4806d44c52bc3023060c7b7eb1f94f9ef5938498f55bf5f
z427faf4c1c792981f5a7917fc1171faa170a69ffb675af4417c325848d5281f47774eaa4316c10
z8eb847fd74194a4ffe98bfc5c6fc9585cf8b9645306a1ca3d2eb322bc5510c11a711d2508b6c82
zf528e4c9deccb56e423bc954d21c04e154a88f9c87f2e329b01eafe96ad05ab395252b4cca309e
za664fbf2923369bc84f728c91336eb8d3b76b2ea5249eb2a9f6af6458fec0a9c54fb5cec8a9d71
z01e2ac643df9ddec73333ab0a65f1639c3301803b7d0552bd93ce2d649e8c8ea41b0cb44af5b39
z50398099056b67429648f3d594d78e0275dd60fd884337f5b5e90dae10230f535f5a3fe3551c9d
z65553744588f45e0646b226c032e379274eba13654bc06170da191711c38d1a72c21aded84b194
zda1f0e70987d93a227f5f314f9cbd2de23e658e436b02b31ba5dfcd407c8052924443d94233d3f
z1d9248c3f7890dcee3f132b3171702ab7b7dd790dbe7b1282a7328d65f0f89c07d3850a1a097c3
z866ad57920906441e88b8cdd57f72a72d800fce3e2a36addc4c31b6658b6f413fc30ec2447c5d8
z65d6d8e903c9cdbbec717aa242d5b7dd0f0b42898bbf470d8333ca6c58796d19c1d255761a83e5
zb72664adbeb64f1310baad9856a7009deb8c88560c52a4dcec518f571aa3075a3f362a12b45c32
z2f6eb37b98fd2e2861140fa4d6575b817501f5e77b8ed24d245dc1edb97d6fac7fb110b2e81748
zed8ed2aa22a20af9f0efbd70e5ec533f1adf96b0f826d1106a19291fd525ef6a07f181050d8e57
ze5193989a156022e66e58fea5f5119ea47b4f9aa6632776a221bb691ba392de5b820be9cd4b8d7
z5083a04d2d33f7e36bb844f77b79cf236f298cf7af2ac26f659cf887a23a93ee2633cce0734ba2
z9f6bc6a025d048f1dfa3e72887209256745aefb63ee25d350ddff02e8e9b4fd575449e6679f2cf
zf5dc90516dcdc18236d60f2a998f49c6f876752d89837ccde69267b927b2415fd077df8baa0662
z9e865801f1dddb59c48809e602ad0326cb1f25f0de0ee77d1b8d9832bbd237e7d6df54417fad00
z4771db87574e4509e28caa16b11e4ab134d386bf4cfc2c7d74b074fbb48da05466b5aca521c2fa
z737af081e162a84a496e0074120287d2d41fce94fdc8889b5d757acfa431b2ba6c7f3115527ccf
zc8dfbb871c1db133ceadda2b9b45e064836d304197af2f639db592c77090e2650670432490cec1
zed27b41afe26c0829904b450944e065c7a95e913705388c19f30a24a91dbc731b12bafc1187053
zd68a7d931249498235efd42a8acd8cc7a7f5c1a6f6f82109053b29dee5e037f6b8ab30994a29b6
z704c03d69f6790262741c82daa9cc25f83214f6f4cc552d653f90f0d7696046265d1cf52f9e91f
zc7b9a710ef43ddf64db6365203c4f86e1c9c99f7cec57b0f9e7fe1bad089bb144e21b40eb390de
z879d4cc27ec0bf22eddd1b84e23e0cb589727c9f3d3561947eb04fa82f55126b8b1766ab258540
ze3cb4d3f97778800de950561342c5f0e89f4cc16a17fcb4c09ddd1651b1229e410c3662668be1f
ze03a6c12e89a1683da20a2ff3d7afcaf1a0645d68f522edd56ff05635fb303ae2bf3d0758b5851
zc0b9c85d42df2b118937df8c150c1f2b03a985fdd4bce7ac160387625804890b9004a9537656eb
z6a6d4c08ecf15c8fc0ff1aa0abc9a80e9862e14c183e1530c5807c40aa575cc70eef83c1ea23fc
z9b74ed3d75b13afb9271deaf7c253eaf59e9b66a810e17e9e8bd9f042a20e1bfa998c6028a09b2
z62ebd2e7b5bcd01233bcafffc20b53248fe4e6240f7cdf6a4fb4bd1f6a3830fbda11e66c4f25fb
z50c08bbeb26e875150427a36184ccda69e3b04c2186b5dd33d0f935a6432ef9576c3b9d6361989
z653d512a38b0dc8d3c74f14dc4ebc422f3c0de667b6dd8f3538fa7acf0a8ea86a2bf4fef91a66b
z85f3330533830a25dda927869b98d4c27607f912548bb0a90411a99124a28cde36f08d50dfdb5b
z189dd062a2b49f7efe59acf8b3b94a071df58a9b91b1a7986dbac169ec3d61d98494f728682c28
za8552e91eaa057366a44cb6233d4593f8a77b36195819ef2a685b0fecb9779cfd7d38694242407
z9323816b7629671028a3341460e7976a55f618774f1c6e42d37660b85d4fd4246d0dcbb5c69b05
zdb2a537fc82d248d60138e01a8664b50d353e9daa045975342129116d75cc4af32b035ee8328eb
z4231b4ad47db05051ee50cf224cccf0c53af3dcd139946af359c2b930035fe3cb6531de7b23a15
z194246cd28c2c4b54fd90c34697ba2588eae15908eb32e7329fc754b6c1c976f37171b2b851e8f
z98ac2c541c3025d754b6207f82cf924a57fb0a06bb923f2cc742b5c6013c2fce9201d9fc3c1027
z584071db5e4d5ce49bc0e403a21757d80d787fef9f04646babe832e314736ab16088046fc2cd29
zac700172c1f74e57113abf9b4e50aa537b9be2f61890ba5b995db84cfe345c663bab81aa86c58d
z375fe3c0b3682dedc4e8c2f02b92c3189c3ca982669d1b57e7071cd094eb347aef950968100515
z45405e4f784482203d884098731bb2f4b38fa8581164aac3f29872172696e282ef7b27c3b9c4ee
z6a0e82822dc47b3a28ef9a7af1a7905defafe818b95cb651a886f2df46358dd685fbb38cbb1567
z6921f02db77bc30b503671175919f2d271e960fc078a53f1a1898e2b81d50b14851d830290acfb
z442a631b7ca07a5b1b8c99335e9afc559aef4718c3d1a333f8643e8c3c0a32553691a05b09f450
zeb6d70713126fcd0448df8722d1119d4570789e75293962dece94fb087f224cd4226a6edbee778
za2f3c8e3f508f1b5c24ac660444ad0f973d3376821617e04d90e3f3e8e9157f631f54c80d6c050
zc8f4aa76bc643a8006085ea9f8ed8b34460ff2dbf746bb9bd928305fe9a0463ad4cd6b6d4abbc1
ze1f528de22f6f460122628cbe2059e36584c5295b472f67cf282ad2d259d3fd77cecea79110bd1
z6d0668f1673eed6c9110fb6ec4a4d4d3fdbab0a9f83e738fd7c10ca4af3dc62ca2e5d53ccda124
z7635905c872a8eb7785362a64bc3ca1c1c23bc3f41fcc9735443bad57b5eddc59d520426875bae
z8aee98de642a35019641f74aed9ee8c41739a57b2055775b044b2b822893426cdd2cad607a9895
zc2e223d0b4ee77f08474e118b6684a1eed1aea8f25362c2857df637cbef99862cb3ff284f1ab47
z429b519e5c011d866e1bea63a0f51c3f422b4e4d734bb86b327f35a4bd4f1cc7c0e343efa15bd5
z72a844db9a0fb5ce5478e68bf2f74919a23cb4c5686497ca7ba63097de96294026df2e2d1455cf
z3e0885e76101c1af748768e522f66b23b5690b77a6cc24a2a5f2976221e19e537a0518f54cc822
z66463d6c4ded781d3a8e374d2ffcf4fd232502bfda44d4193d4644bab5f55e291b8859fb6a57ae
ze74feb203a3be50080c036e42dae50db1f85bf3fe99dc1a9666dcf0673b25ea5f70d56ede51074
ze437b57e5c419ca3344c2440aace4359e95dad0cc7a4bebb3d2a4dd7c8881da9d650eb1432451d
z140793c345dbe09772d63b14159890872915836a58f3e8441f2b6048c993decee7c3d406089a95
zb373d816498c2cbcc9f5b6bdadff2fd3c8e8e61607b9147654846e31e7d63c7934ac452d4e40a2
z050e93d6d08572a656e1c448d0cb99fdd65f85773d742949c1ddf0a1cd9cdf7787a7252b794935
z36a3c2f63187e7bbbb8f0fdd5638932288f5760b173c3d51d354793409913b59a06bc133375d9d
z8d09125c7ffd18a1f9fb40eaeac67fc19f84ec0bd6126eaa7757bf70101205293aa6e1841501a9
z328611392853a6c7f7e66791f5a60725fc7ba3274055ce5c8b2141c5c5ffa268efe9741b2c5194
z5b2b97e85491ea98da75b7b63698cc522d909cd817c75a4a7198ba51ebe71da6570dd54b50dcb1
z860134a9c1a4cafc7fa6d8eea055364c7cd77a09b7ca48f1bdab63dcdd4a0779c6ce2fd635c9ee
ze045d90e1b4ca16e53781dc887de43b96b6ad3c0be2581103cd8eabe0283058961f1a267535459
zc385cd422d3482537218d7a2d0777f064fec891485e46a9e71125e6eba51e4176de3aeab47fbf9
z3013bccee56fe421718f998db2cdb811bce4fe2926a2c698d2eb0f6746abf55c761321e3846f4e
z51713af83d6acc5c14f333a22c863953762638c6faa7f5b2906950e174a86c4f56af9ca9c19812
z574ab3ed9a4d95c4e23afd2bb37b6a239667cef974de8fd39f323dcb92df3689dea3d7f6cc71f7
z1592bb0bd5f8a72580f99a40eb5316f327435fb8b8e52e868b230eedeaddb87f369a99bd599a38
z86af1a29483fe0ac80d2bae3b985ac4a99d96948dc3b3aa592e6ec69ede6ebedab2772dc735b27
z587c2c5ec8eb5d85bf6b8d7db95fca956b4e4dcf82dedfdbbe203ca33b4a105884f3987a1eb18c
z1615e3026a8ce1a43fe4d46a6489b731babec62739b1f03a7ee3b5eb66ff4aa0a9bda32f29d00b
z8be5037c3b6948e9e592c91f79e245c0430e012e50c6b7613b249daf67e2e436f74d848906f622
zcaaeb9501b74590bef22ef8ebd00728e1967d02fefb249cdd41df35c7526810afd80f1f7548aff
z13babf5bd46d2913c63c2896a4faef5dd11c16e4b45decbbe164b21797c775a9a669133514d073
zaa91b05eefdcfaa196cf980a486a9bfd15fadcd8502226dc738d57d9430bf5ed6472d0d559a1c5
zf87cd9d6303b46985e5b06579b824848297a5c775d3c2ae3058fa529a1d153a5ce7b6d3e33c040
z65c66fabf1d24508f5bc9f1ba6108798879dd2b6f6c04d554601c2258712b01f9466abc36ffc30
z2c87d3fc67796207110c0d1f53d8a2be8d8de2dcbd3a2a1bb6d731aad35b90acfb6ca62ad399f4
z8e60b0f5361dda1690bcc6d3b4fcab56d06bb701d09c307b6084e229d6a8a6efb06ae03e6fde1d
z2655298d332806dd2ab5621c0529ab2e02b46da99f04fbbeb058c9a350cf62fda900ae2c44a78b
ze95824c3cd69fd44e1ecba8bf204bd649d553ef7a42149ba5e4ac3aadf403f163b2d2d04cab4b7
z31f04b6a5ced7d427f9612a424a7e8d972efe24cdfa8de50a12de806539daa410f279437e5f9c8
z2ec06e953cdf0e30e4452c5b9eff7b80fae37d3357f3641516355cd4e0110a68c995bf6416fade
z0982e392904865433e8294c28f3644020da4996ff721e108637d330f20667a1ca962bb01bed631
z639c2fc38e998f78c430d152b778d07a3160eaabd499d5b5bf2439977bb74bc1d756cdb9419666
z8e6049160d8d6cd09b120e3e46fa313711857db031fb4c0aacec02a0ea890a2f35d6a58b83fcd8
zecb1aa30444352f3deee3d578b288e14fae3a4335b3beb70bd17d9d4685958e59baf0eda87bb78
z41689b88627f4cb77243da88283e6378a2dc1ccef0762bf234ce46390322aace6dad261a0ee90a
zd96eccca87d3b890c8705a13860f4aa924dd73d2965718ba70a71e2ff29ea96bb34e37192be317
zc1789889a127f929f03344d3be49d5def865c61c590a1e769b6f9fe73ca83f0f20afe28ecef2c4
z373d98d99cd95636b649d774b08fcffe9d32f7307862a917827d7f9e0dd557f7530b7be72de15d
z67d9735a7368e51c3d7f00915611cbd2e9213d9f37d87eaf83722700decad46b0abbeae73d4d52
z6004c9b73f32fb2c841d30b7f8b13652c3d3a77c2359c1bcebc525be903fe804101a50dbb97358
zf760a8147268d901d84d95cc25cdaea4f396dcea6b8bddb6480ec32ae202f1c97dd0f566c7087c
zacfc0894798d9c67fb65c93aec55cca6ded96cdc2f1a98dcf9b7d9da108906d99448db4ce11be0
z9ea7d75b4de5d4d8c32ec2e904baee3813ca7e8b69ca9790ad6d53bbaac023e70e5cf3b6f25738
za59aedfb25ed19227d2f51a256e915dbdb266b38fe57d1e234a97a192a29e374ffcf7c6dc1a574
zabc3176a1ad2061b48fdae2bb645b9d31cf3151fbf3c5de84e423c17271af71015c81d45b21cee
ze938290cdc69877123dd39ea5dfd05521b4b722d47f8ae32499f14c49c128fc452b45f579fae5f
z9afcfa479a5cf0b2a79d1b37ffb602d6af9df7992b329e9cfc7a0f489983b1d324691b2c163c1a
zdd500d61da1a4738a2f5374b6f8c665343d875f823e23ef0a8dd99234db26e93ea4fc3c2935a8f
z40278c2d1d7d67008bcbc1edfac8d963f01ae1d0e04c8a2c508d4f53e7f7e0656dc7005a497e86
zbed1db60c848d5376ef0bd3ec75e7e840287851ec0f43b436ac8aa80395beea58a48d465f05006
zf7462faf6e1dc70d8d36806947ddd2b46dd575b5324d9642ac7ed19ec94c971c18c9e91e6a20af
z9ef4169cd682e944af5b9c6ee61562315d8a0ccb16c2bae4ca7e119f72a9b01a2a961ee560a046
z2527e890a9b31bb7bf44cf930fdd014bb727e61a5cf3b7870d2832070e312a0d474f15264cf9d6
z44cb5b464395cbf8dbc86c2a6ffa6bab070e55024f4eea3d9ed43d8fb5cc9378e38073ea4cac34
z2508a7ff8c6dceb56af8e9258a4ec5a20ed3e1b96fa03706707c721c44918a04a7003d055b8a47
z373ade60bfae4e5979949b92aa3c78006aef73c23cb6d9e05db6f6048a7d427fe6124451fb9c6d
z5efb63835e6e4100c2aa8aff9e50f599edc5232595b665ca6a3df2ffdbed108b78751b2235d896
zd6257264bc21867cebc6b75cc9b651bf74a24fcf2e97be98073b3d87768d69094ea6afb07111c9
z068c866c26acc06be653f3adfce0dda6fbce8ee0fb0bc6516e20fe09f96ee46584952ca5bd018d
z9822877356d81b63e15302bcc734bed5702388823569135db67bd07af8a8aa73a11ee30be9f7fc
z09ba013c3b170ca2e716feb4230f30e126d15409e4ade67698a522709cdf6f177703b3e9f6d162
z272de507f1f6dbcca7aef921eac03f0a0629151c649cde2b62cfc1667ffcde7e10e0851c96ffca
z058e0dfb0831d4cb9efbbe0bc7fe6841f62ccb88366158317d1ac52c2ad66ac8e35964e2d6e7ba
zc38bc2a48696c841fc04975e2cff33292dbfc9c0493252bf61d4d8e4c3ece47ad42a69e06b4e65
z7184b26e70b91e61c463de740776b0e02bbacbc555c2d905c41b4ea29ce54688552a0ccd02d647
z7472b363a8b760d5d55c4457228d389ea5956a7185061676e220d2e819a120bc6112192e004ca3
zacd4ffdc4846b541d24168947ad2bcc4d3c3af8eb2330c0c5845ac31414f032de9d20f59690b79
z707d1a1c46400cfc1cf6304541f81d8448cd35020440e7ebb1ba490463872952e04587a78feeda
z4387e87c7c6c6da430e9ddb223de1de410f33a53d000cd6949d317b2da37e46e4b4a93afcf43fc
zaa7843f030ad1b322236407369e94ccbeb6782b228f51b4182c3fa6ae0dbdeda3af987dbac6765
ze3e8302dd93ce02276205488e058591d079d5c091169dd86654045ea28fb1a5909c8c5f893c5b7
zd25038415eabe8b0d7edb4ac000a75c338161d570af710fb608f97299c5bff4f4b98268087849f
zc85a6f42a12f236cc0a3e125c26683b2118dfdc6bd0c972ed6e99c58b45c618ecbd14cfa33222d
z99872760b64fb61ace7ffc936415061d61de6550a899fa842d413ddded774a2f11e7efc9d0e194
z4d0097e89c4bf711431d8c0e4d15b1cd436606b0e736ee2e6bf7200dae7fd4fb45108743bd13f6
z6c9bccbceccecb77766ffca1cb334fe7cf07c7608248ac026b2af42c8ea449a77b845924c7ddbe
zf887e342aefae91260bfb08427144aa5bd9cb8592a156d2851a8986b51c4c1e89d6a20147b59ac
z29bb0df57c46ffb92298a87b7091d989df48cc2811afa0278fe17f4d4dbd16be9d3a33b8b76748
za8ef46d4864e1770561258a17a58351593fb47b1f2ea4277148e0357c9bf77277cdccaa836f19d
z0f52118f70715894aa69319d77ad70ca0d7ec9c44d6ed0842e470e075110d45c93a210dbb37785
z5ad66d8af02d96455985ccb1ccb3cbe993360919d9f38033d91477b7faed7f0db17fa8bb1d7fdc
z39532142a57dc37d961fd8d4fbdba5d04ef5fd18b6cb92f858d2f4551eb0571d77d03a775f0d81
z291389483b77a0c1c8b37bc7922ab4e89de634f55f5f8689a96d73d5d7abdcd08a478a3f969fd1
z7bd9dc009efc0cc279a185852fe695ab9237ee4fd6c0a1bbdf5c081f6f1b3be0b806ef19f92026
zd63b9db767359413c1efa8bb1678418fb1ad87e918e900a5159c4b2ad977253743f2b23705bb57
z41e86f56d9b6094245540014d68689a501d06da33cc88a162db3caf6a3c621a040aeebcdddfaba
ze5d766e715c007d13a78110369898e0d095fe0a0a735695e5f3ab1c3653b09dd12c134e9d2612f
zcce1c8df5eca6cc855c8ac867ff472172662d21f8dcf5ec0628adb184c00b53c488be0ebc1c878
zc76fbf5bd5e2fe7348036d9b3c7dd0003a609a4f1cae32e517e1f47180e149133109c27ae3409a
z53a4cf9fe1a25d3b1fb011709273248d41a230e13fbef5492c4ffffc69f1798443c51af4ca9e27
z1379b3c59fd53d3741aefc73bf905a5dfe40c98d35a898edecacdd215f898e557eaf9f052384fb
zbaa17231225fc7c7a01ab0a8e2b78bca3c2196b2bf0bb2eed2efbab944299ebf261570e1fd28a2
z259d71fb8724eb9a16886cbf69d702a31366ccb6620dfbb3fda12e25e85ccc96041b9e60e16bc7
z6fe977e676be57badaebe09d9d635fe8cdbdc774a3d2c945c6dd40675adabe0bdb2f48aaeb771b
zd81177fed024cdf3dbc6f922b11252f9e574f51912f25b4449553f28f0f9b455dd3160e0214d69
zf86e1c2d2eec0252a6970a9633e178cad01c6d4dc0018cffbf3038c5b61f7b455ab21d1c517773
z1990e814d9a44093676b19876e71ec2602f9f45998cf5947666db745fba79967f7328a2b37429f
z34e2b5064db560e1bd0753946319c198439d0473a24d5a53931243bd08475b43aeae51265f5d29
zf5283c2e10f371177871dc7bb366b68eb14b6df87855085400564c518e3a084ee5f96bc2efe322
zd481d518003352be82c7b6f0b9bb666e93c1ddd31dca072883e6df9861cfcb8faa0cb2699f7251
z1733edd69c61dfe87bac23d4dd2a3bdb5d0f076e33932db0b7f85ad178cdc3c66457c7f885c219
z421b3239579d00ac3303d4c33bc2621c01f40728c71ac2175be5f4fc8041f4b63bf131b3d2ced8
ze62b46f548bb9e4664814a6e70c2aa0ae9de7d22b8e87f71c3c087d2bb8a29e96139c6b550c12b
z9405b1c8f8eed3122f2893db1ea3dbd7535d84a1e76df41746f8eb9425728dad3e28049766886b
zeb7857721a3f2994b4ab792bcd2aad55fc2e8b1ed9ce0f90178ad67ec16451a51b28f32235c607
z4855e67a3c178419e77b0d8a0804d3354c677a656f16bc1d82fcf398fc2db65c340359fe57dad5
zd4aaa9b6f7677af89d45743e7480b29449258f90e646acdcafbf3fad27b3b2ec101b9557fe0e83
zd6a774aec1c1f6eeb1ee07c43ba68f453fd5f49d020e9fe9eb6f308245780f22493cd17679e954
za8a194be14a445ba54012af5410e5c66f398bf02ff87ea2776d78f40b834a084fa229f1115d20b
ze51a69eb7579826d3eaec5f9d95e3db600a57a70463b756d71aa4b777e1c380574595ee035acb1
z49f6a74cd1d3a490096f1b6cca86ee7b09d315555f6f20db2e62222afcc11dcd3ed5dbe1fb7c4f
z241321c434f17edbc7c32680c057ba92ac89f9548dade1ef907c820991490ef12fff285df7298c
zfa6a8a02821746f4ab0d75fe69d7230b2e7a1d7ac6f9de8fe1e3348cb53168ecb0f3992a6455fb
zc448600f747434ca6230ed88f3ae6164330c8922f9289656ed4503bf95ebf048bf3af850f5deb2
z14b34ecb7c23a4a55530ef8a086437d1fe465041af5a057297a2a894d5f565de6dfc742905422e
z0d1f1185448becce926be0dc9f750305ca0cd7f7986fd5255707d681d1a889b5f1e99d8c208a8f
zca5baf5d598b65f076c845b52f3d2f41869139b11253b1f62333b5893fde6997a6250e2b06adfb
zc1ed7d18fa3a19980bc10a9cdfa76da4999ece6472a6ce45b0f4f650460a0ae1123b6dee915b0c
ze1c7c9bb663d5a23f219200a10e9520c15f5baa7b1d18d512dd59f15aa887762abac73ef4ac2db
z13181ccbc0ab983dd4872428da791005ebe6717adac251213c0fce8758d89be486c6e7c9492b6c
z4cad8ce1c1823493eaef77d58ba4a5e9dddd997d0b1631988c1dc494272af6f8644114199a39bf
z722f7d7a39b36630392c583a3a9a53536c73e967baa9fa7713f793cfc87cd320b3e2086df43366
z310154344da289014580dd7ab73d7be6ae2dfba71d2f4aec38e2dd781017ba5ed032311b80e386
z3f80a9e748ea743424f86bc5efd3176ba8da66324cc4d8d7e6749c6621862dd4e3252d19cfa5de
z16ae55b67e56d881f70272536e20fdfa4976199c374a83cb5256c4491918fe70c3266cbcd783c3
z938df6acfa1e652f600e9d577f5c0183a86d63f74e86a91385437081e71f71d48c0626613a22ca
z57d995dac98554397038be52daf5cb5cac90f42cda5dd62abf7c21f6c245694ada42d2cfc6c469
z3d50dc4db2c2d4db47b69b65266054417e4e3167a3496a306e0a9630081b7528ef5dfcf7fd4c42
z858b170b18fe2686d35cd41cf2517ca6261617959af69a61143f935bcd65af0dbc741545b2b654
z51c8f9fe2923079ed3bf96d8881d87b63c06c68f45d01414b5348437602e06bb76151d58a87a5f
z6df93a2060f081af23dbc858100f22f41628cff38257846e5172aa4a2888353ea31ccedb01ffee
z19584c84b4c288275e0d710e30c9ee159f3a6c2d6591824c7201ee71ec02796b867ec1a92f51e4
z87f6bf8eca98d146b6c97e77a966d2e57a5e02796fc89eff0f0fb90fe97b264d7fa26d2eedba52
z5e78fa6b1480acc1e1241379044af9d4d3c0ec3425743f7f11dc01b2b09136e096e538f36cbf7c
zb6c4355bca625b12ae3f83218cf8c72170c04f7ea050562a906b2de709a1f21f53a1131633f74a
z4b2b7d479e3c2406e405e62e9589fad7f13b4378fbf53bed876f4bfc0bc7f5e3d731b49eca119b
z3858ad65ea3ebaf89080cc467b7a0503dac00cacb651914d391c78263ae26d59c94b167416cb5d
z072ba4889fe5889b58b3b10840f60007752457fdb9a36f52c270e65024d540d16311b48d40fc1a
zd2072b5977531e97088d033e1da774fada70be0af4ef7f37bf7999f9845ff9424570d980c42f7d
zf5a07bfef1dd3dcc63e8b90fceb16dc6ff7eaed1998ac07865e7b5cfaeece72ba3cee8b2b3c987
zb8e05281069a68b6661effeca91c6997d276858938bd5ebe59ffddf7752ec61bf59255086f3c5b
z1fa6a2e19d1b6c73d66e227ca9bf21d1aff64eea692f65e49dc6dabe15801034e119371aaba37a
z155cb8a51910f1819ffecb6204b071262ed40481b2e5fcdc322940e1bdf2085721d31f05f89875
zc1afc683d5a8eb1bc627db66629cbd0d62de32d371fc368bb0dca3c79edc70ee56b7cc7faeeec4
za6e08e5200bc912df61a656af018eede34677019536736c96d6af0ce21acec55b4a7e6bcb72b0f
zd54255cc54433113a62531b80a5c8b5904346a283e605456aeb85371d80203507fe8653912b1e0
zb5af0c87b3cad9444164b8f0e98923efd58c4910acb6df0f92446bf6a712a926867ecca8f6b82a
z96e4dce2afd4628e55f2da5ac9b4661f6634aee4d6e20e0eca0e27aa265ce2e0fb1608b6395712
z0854abaa9f2188a319177a12dfcfd091f295191a7727b0d36fcf949bb87e258ae59cdb3ab38eba
z45363b23ed36fe2f8c9614d597507983b0f06356e3c0f10265b91c917ce857f337e8dc37cf5d37
z95a84647c8b0fea05d81c11598ee4277b1f4ab72317ca055c5fb35c31cbe8229b1dbc1bb4b348b
zd756bb8eac36d3d68f2bb99c2de0ac487dc0170a546f5b00d8464a35269f941a19d61d0f43c1d8
z5122db2e7840bce59012d7a7d436328d4605c047ff074a430abde1df2d0c7a05aac9201c10e514
z4bb25dfacf50cda1111a2a03fb1f88e415eafa7109334d760cd269771c3a586ddb4e415f9f9b82
z3c219a6b19075e2056f2b88c5b7ff0bf0f752105d714eac07e00b68886ee23e9f1f174ea70515e
za7672640e708c0809c038b769fb92bc76ced417290f208a391f2e527ed33c3bc01842ee8f9863e
z5997cca10f4b851ccf0f243e7e08b1c64739fec856bbbcb1e530f919a00e21d01a8cea308aada1
ze0bfb4274ace2b2973352c23ce40b1afc3c7a046b192b0dea555fbf948f98f9ada1bfe4af342a1
zb851f0cc7061b3324b513d6f2450afd90af8bb310f801232090a8d8e477691e4d53e582c03e803
zf303e6aa63652baf23189719d9323791e7920497da2aa4406dec6a2055ec33cd5cfed4591462ec
z650ecd39d1517a36c862e593978dbecf84b3c3953e60a64aac09f7042d07918c9e2b33594c85ac
z2f4378d7b2897bccdbf86f80222f0bdcae5982383ba34ec5324d0e267e3bb2634ab967adcdb1cb
z7606526bda785da64784b7a14fb3f0d279c2164de7efa582973ff8655f3e41c14732aed5b71c2a
z678e7ca30cc4ce9875570a93c9a47f8ee822246e290383acb6479cdf52761d2160d545d2342d8d
zd6fac95848e32b31de623039ca6defa602f920ed688ce9c725cd5700cb89607c8ff188a45c9414
zacd9fab13bb02dd5892216e356e05f194fabf3ce5873863a8b4f69e171429b053c52caff30fd5e
z09b4807265ad314b9b8f51f7d1f70fde7b2d6552f1509a270dbd9658983413611c04326ab007ba
z8415bc5dccbe33e04a457bba9ea1278070517655fb669a030537b33fcc9b679df2e8961dd4af60
z7b15ceab43346bda1103106aab42548e10e1af9dcf052575bee7875fc0d024f6455f7b6b56026f
z8f1c8def6f8a7fcf52d6714797a4285983465c6a88f68efca27a43ef2c8c976ce7bdc4f47e4e1e
z5a7cabc5295e983901cffb23c3bf19368e94f11f1ebb8c063c750788ccdf57a5254b9057795114
z266309d638927efe3ac94531d415443a951fe64f2cefd258656447233f9a84943d2de3424b3cec
zf9fd9b0f60793755765af9b53135fa52658e72a37c8aead7d11258139bdb5525b3720446a42a94
z203f5019a34429a6f0a28d0a0ecd889cfdf28f35bd0efa2533b30947ccd514bc6d6e1bd98701df
z7629007176cf1d19448938a7b166c9e02f073f0d73c18d11857fd35c31caf62134420664746796
z1710c7dbdbd8b4b271c2d9981b7fea6d1d47f89d57d057b4412a5a074f234d58cf2059b633d855
z42e4151f789b5cacb53b6dfca2d910b64ba2bdb179e11ee32f942d10013636f9f3bb8cc0eaa6e5
z10ba67c34b9779aa4a3dc5c437664265e4db377f0b00ad771daca5bc7702ed2e85da53476d9e11
zd66e46e0b296a09f039c57d790107ac065f030df3429c034e40c2a84c09314ee6d890f6755997e
zf4c44572208a42ab41d2d2197db5b83b1a54f47373a6b44a71eec3b725208cd18654aa9465d7b1
z5ea96de1b014c7a923fc7e31807e2b6f5c3637a41c5f5a446d6c1f0fd661abaec279d9be7033d7
zb14e405d7bf99a4836a5fc3fc914543575b4db4fa776ae27d277d80a363a9f4507d81dcff7349b
z023571df55029eb42fb8360b854f576df28482e46ad1a4f1ec9700cf08626a43652192ea0d9ad7
zdfa424fb350b34cb9b02983ef54b91993f6d9f6f31ba298baf614d726a4f03457c71d0698d07bc
z0d79c5b79f19feb3476845e020526edc82dda0add38bbec07734b38aa28dd2f407ff51d85c424b
z61d4cf636527da2119591a3b9812078a8d5ae6fdbfdcc36840e3a4e0f1cfbaeb3e5965f1d3f36d
zb19f09865a3a3c2e1d2bd76fe9307da8da3412f4d8aeeb93f1016f2f1276245cb3afa9e3317c8f
z9683b4d9259dab90d025a80999dba14f0287e9c5c9a697a731ed940c092001dafc3198b82d1dfb
z9c82cfebcf3e31f711ec9963f35b12041fe9785e7457b85d083f306944e20fa67063f560b539b0
zd66530154f09c7c3b6b2c0f30e8ccbf4f1e2becaf32c4460358817125b8c138bdeec8a1e6974ac
z4409c0d90958d1430691e07983b0d95bc8168a5c4ee7a611d32eaf04742daf2fc621a3d24012a9
z9e76ecc2d2b05d476415702b348fcfea47e561d1a1ba4023a6b9185b912cfb5368a9f350d27670
zba4751a82b0db92d9244b2aacee20eaff70cd1df643740b158add794494ea4e56cac44db115763
zc3d6409dc539404e91aeb5384fa603b4c3dd6c99cab140e3dee1a4a3e2b4a58e0e4808c7d807e8
z80d470c555debc31068984398c15fa14ea4534978f592ea79a85513da8ed086af79e511ec4adbf
z4a31ff971d81feb8c4b21153d99c45fcb09502705adb3b65408f6ea96505ac309573635e08788e
z324d2af0b6c6da255459c71d632889c6019c1c5b0966f6878989561385714c9b462571877dc4ac
z5895c1dec2bb8acddfc828891ed535c4f3c7b57dfd29d2d47998a7f279abe62d78385faab853ba
z21bdadc7d5138e8097b921c90e1c5e2f5a0e3b156ac3e516b9803ed7daae609273ff155c6b78e4
z81ba3cc88a6ad87e2eca8688afdaa8306db02a7a30de64065779ef2c474e85fcbff77e2d46159d
z1c1c91a6c8af8603e650ea1720425af278549d898f67dad79d0189daf4425f48a355486383e137
zda1db7d38526338e3521d1b1fb7951d2f4f224fb74693935dd56e5eed8c70bc6ac1d2f119ab746
z55fbe20c54572dba763224534123b631975f9463097ca27a29a3e43e6507567ab443b353e3994f
zb2cb34760a2df530464a44bd4c77c768b78cfcc8bb0ba7b1d647d98c0c4237eeeb190388472a44
zeeea65d5b9e55d33238dfaa204ca239d949cba1bd099b99b1c94252229f904473acc8b5a76c5a9
zf0b05c4ccfd700bc11813e71032b0f6c4bed7a28f56e30f8a62f5be1caa43429f1f472c33a7e1d
z9576cb6a0e91592af064076dffcfefb9e7cbdbb1987042aa905939db3c3f895735c61f7f301f7b
zbb22a06d2c4ba3d6832e51c3094e98a22eabf5fc0a1cb65413a801080cd068798d922ad26c60b1
z4a34536b17514f82a216c0b537a99c2da6ad8d1e2f787116fa8137dd20c82d9e962b435597aabb
z380bd955fc9f5908dd1ed720c3fae0a16fc83658f67105f05b53b2539820a02edefdb178c6543d
zca54f6e896cafb61b71b67274adfd5a10d1489dfb14569dcdb5c1f1200f4e96eae34a6da22b141
z09164abdbc63e62f3db8d6d0bc17bf6cd173d5a87ffc3e5f98a24b047d23205a33036f22904e44
z7a94f4d5799b0d7c72333687342e2e9b4d7bacf4101baa953cd2bc318ba6ad400860926d7390a6
z3984099a679459a03581d84e94744c3c324883ceb2aeb148767ee1699c12e83d3d0034c5879e41
zf37a3de00d4c454043920b9657dc885dcf6b4f682c1ac6ac52c5c212cfdf557f6327960fb064d1
zeb1021e7637e28d45fdfff34dbc2adad936d010b8a7244410ae8be1c23bbfa659a7ce766c76e2a
za1e80a62caedca00954800d05cf96cc27920140553aba2deb776438ae57ad5fde868087f304291
z8f7c10a4ed3a084141e4a00810f21f7813e71959f79eab93937d2a782af9942b732535a3df47fd
zcf0ae260e6544a8dd79e7dc691a76a557fb3f793fe706e8be6e2efb2cf9434aa3db37c0025103b
z8ad5a641b3035284168e39031d897050f4ba85f8e22d3bb2b27750a4f82dbfe645b979bb68c636
z8143cc4de6079350b9c67350666daa2cf0a9d4e0190d3a0347884c40efa4773c6a6d2a18ebba0b
z6c0a030529c924aa1674dd897b6bd7e68b9221a75df7cd649c6a9d0b0f4e0fd09d2f637e54f878
zbbe5124c340f0d39c5d1b623a848367489c6d8e2be8b275a48b5a55032b343c9a2b627343c84ba
zb1bb962f0fedc00af51666f5121210cc91dc31e6ba56a689635a0d0bb801965807732580fd27fe
z7e9fa17a138cd219ed792cae5046ba20469c7f5d89d05b5d08cbe35a764d604b7c2d7125131537
z075453c93dab059163540e0d586bdf99a8e7cd726b0eb69d2a90ae814cb3018b6817c150e6c17d
z537674f6e20ae5405a98e5f10cb69ec3a9225ac18ffc0caf7ad33dfeaa340d60e0cadbfb8d495a
z07f9e152d906a0d100169c5e5c14d161f1cf87780dbe193fa9e340efae177fc0c3f922ae33a10c
zb7097a2643d9fc537c2dd0c0e978b5d74db19a12f36a8013bb3d8d3989ced23e2f145c19e591b8
z82401cadb124ed5ce0678279404b26601cbacf459c52126807d1eab1d11f8f1ee11f825833717e
z84b4fd9e3556b90cd6195c7bdea64d311cd1ddcb4348a80d53cc02a983d3b0663ccfa0077b60e2
z3e88e6dc59399d7ff1260fed29dd2e5b3059d5096e751a963099ea6b356894f2422b98b00d00a4
z8745ca89d3ba06665a9b979bf7d6d279f5d3e9b49dd0ff2b4c9469c85813560c584547de3e58f8
z1b3203265cc801d2b943e1409e93ce937c81c0db619d830f2901311cf91b7210076dae9f643e78
z5175ffd33f6a8d085fab67c4e117d81fbdaee23bc0abee807ebadc60b241aacc883f089bef86c8
zc92834f4211dc972d02fb9dffc4451a25b2a39bac819f5b1edab52692cec124a4bcc4bafa7e7e5
z28b805353379fd28e1f3ba014e5ba19ddfa1da62bac2ed1fe52419ef348c9538120c7acc3144ff
z5fc9722d41b4df03baa934c4648b1ba7c8f2555c62a2dba160f00e47db0bdb1917cd73dc9d254a
z79727b1ccbf6941c820d20d636b8f1bf042b59c12da655864bbd19fdda5bf294a33654a47ecbf7
ze44f25059e2ba7c960193456b2c7d7a824a5196690d60f8faf403ee87c116718890b0e63bf3074
z55d649138d3f1911bec1c644e2736afa31fae4d63d5901c74b13d742c11982defcd4b26ac3ef9c
z0b34575d1cafec40fb158da2afff9da39d1ee337d196b223940f46d5014f8ce0fc5afdcd97194f
za2146eb4bbfafd085e3b7091e2da83597e9d8a14edeffdd3e3edefcd15874d5625a624ad0d286a
z5871bcaf61fcb26269b16f86bf1a814e04fb1a24b37e0f025ad9917116a83cc3875f2687e391ae
z97bb4ea3d353dd3230a59fd73ffd453d9564709c4423fde4169ffbd9f427d97978bf4b928e8617
z4b49d7c9c185f3d3b1eb05a181b0bc35700a4210fc6d29b4154ec7fb991f7a0800e13d96506a31
za5ae4b8367af9b8e956029af1f4c2094ee14e1cbd1bb757cfd7f629e7e9ede3ffb56d91eeb6cdb
zbb373d89221185af2a60ab73be7fff001873cb5a9150162b8f2bd5f60c5becc0163775dd8fb9f7
zdd7f52a64b68d82c9b2a30f6621c4ec81354d3f99d35cfb47edb83c0b1d0015c8a830bea8fde2d
z49727fee5a496df0983881da9193ebec5652097622981a968b91659119f021cfb96fac38b6fa00
zca4924748db62c93baa5171a68c1f512ff76dd42ba565b339d616bb674d8800e6467e2ec21be72
za25740907089bc3094d01782e4044a689fe150f0043efe16bdbcf4e0f46356f8e7c5fd2f08f78c
zba7ce9e0b1cb71da4e04a7d65d9465c4bf887f359b2b55b212ef537bc9df3709fac73fa0b770ad
z048e8d80b647bfe344a73e130744112c8437b9374371f16e69731410339f86e92eefd71261b27d
zbff48e46d27f4c353537af4c6dfb9a8b71d7bebee43d77b18c28db3a339f39c5a529b540595819
za275b50ce31576fa01fa378acbe7ac24ec360f935e8b5f5c25b914febdac1abcc820ae4a33f7e5
zc5ea535d1a6eb4d06afcb9f2041c91353c70c2be60f65e26f73901983ab583c9d16df1198f7ec7
z8e3f24a12b57419b8edeadd5945cffd201a069e583bafd90897c2f554b54e4291e51eac7a7d41d
z9d0f65251d932fd2a8f7c8c2d6579fd4593132b45430cd4ee3e16ba6b019ab23e14d41d766aa9e
z36960d2e2cd3460be44474bb51041ca0988b477f586b2fb0bc634d5d7fa266ebffd2ae3a40d0ad
z7c2f3013d0c88b1fecc427948c434f670d427c7218d1d977470567f736e96471a3236b71c96e86
z55479d6e582540bd186332f18833dbcfb0d5fe36a52ebd821867274b15155e549e99971deeadca
z9fe9142cf7099f09ba1e4fee7e53413948c7b2a1ca321af210a2c1e17fb2fda3efe7e982db9164
z49ed07b36e721ec5528415b29b9b7218aa51120e750cb0184fc39972f4e879cddf31610264aac4
z8c919c5ff3c4abfbb0532bf9bed0381b9d5781b2aa95020f794e63f05fea2b3decc26d79d11417
z9e1d7a15b6e41d40bf3e476e08dbebca1fd77a3c07ce251b79258140808347c1761909e1c890bb
z3ff2162a52c6121a9e2784e80ac7a4654f7927d259679015aa4ede800e8390f1d2d8177b5088e4
z33da60636ea646abb71ea0a6c7e70eaf171dce0e86b1bbc7a96f0283f0943a00f12766880c8042
z380a43ee551d8370f9cae5f37e00564aa22bf0649f648db68ab8b10f66f24b1eb8da9c9dee2689
zd42daaff772da21179d8e86558a1d3991a8f131741f7f12121d92f2c6dae39e9959a45bed500c9
zd2192f2b25e5918e7049d693da48917fbe40edbd951154541474266c1f65460ca711fee35395dd
z215813a38db9b87d8233fccd7d86d834c4ff7e4c7e05c34d3b8fe9709947a09a7b5f68dfef006d
zad479272f2495ebac384aaeea6801453ad434c7a4ffc402e85748163400587061df41ae20ba0da
z4ff7923366d8bd90bf92a1052d917c0698299725a3a1832fde36811457082cb13d132abccd3bc3
zce2c2fb01b730cc6f7061283815116e619a1d16f6525d965d98b2e864b604ea3731a34ce7c25fe
z4c6cace225d92e4b54b85cff7693cbecc1b8b661563858299ae2435287e964b282d6b5868f56ff
z0ca6fb5f0a02b56ed86fc086bc198e39b8cd683582055379fb83c8218166337f08102a43bd07fd
z733eefc36dd7b28875bdb1807a7445ab0d9ab9b2642eafa3f8d1f8c0f4604aab96b9f96d318f01
z693b302f521c807ff4e5441ae41465053159a803bd350175243a409836a5671b8b144795adee52
z6b372ecb4c946d1c6cede6fbbd12d709c20b1cd6b3374cf407bc1ac522a2d3ebe9c272f3479434
zad55df153ac81bec1bf2ccd344f158df857593a3bf6d851552b7dbb86d34d51bbda35bb52c1465
zbc23234f899649d01bd9a036b5618827af4719ed44bcb73ea2a94261f2a37ad1bcfabe67219888
z96c9efb83479085d1a3d37b94f533ab0cd586573f726dc478f3606e54099c7916728a9ded45f66
z206dcb83e3dc508a23624052e557bfd30b21a1f093716f898b485769a21e8b81737c068c3ec414
zd64cef25c376068acb8f8d0d071c78326f0a209d2d3ecfa8cd8bbe75a108b6062c4ddbb8ad0044
z66140e4498317532e29f385f3a60a36ccbb98866faae09969318704f8d16348b68646bee620189
z40707be52ceee50430faa8b5d1fefd7512e527d4dc56134b1ea163896df53144382df34871895c
zb4a0e4da5e28979c4dee1cef70841a0cc42314190d66e92f229b97e21fe9beb2814084bfc96368
zf2bb9e83ef9194e2a21909356b10def6b23510521d95892d2ff682ed4e415f54e4b883f28b8cd8
zdc2c5236e33e98ed7dd918d36fcc521437f10383e529d782adf5dc24917bd5e8496cd9c1d26e5b
z0009beb538bd5be866c0d342e7f11562b28ecda84ae1f2222cdf22a3895259d3cdc2f578c491be
z350d2511e381b740fa7fe44558bef53514c80ae26af57b500c68e65ab6d7d62c64f92347e54d00
z3c31a03d43c90c342d8094d22b6ef02cb344cb892473e0bc20f164f672156387384e17d04a7772
za25eb21cf2c4ebfce8b2d4d3c4ed0d411a9883e0c4ffb6ace4620f9c5de14dc0e352372d0db036
za2e1a221d445fe8a3b62e44f5955b8d99889043fef7b9b9a913cebd57a9dc0a5d99ffe9daa689e
z050a05b3540b3d86fe635b999f05fb9790db07993f9161ff3269a783d32c5b952f3348656a8eea
z874dfec6eeacf03e1a843e8c40d21cf2f189e2d5e544ae6d7bae0d0049450527131aa69ff8a12c
zbdb5d4e897766ae40f84e52012bbb96f900412801f826c7640e1a5b5e39689c0ed5fc3391d8e20
ze5e62c053d2d191873c7dead61962ef4cb4501fb4f74d256649b85a142a1d3a171b12b7636f9ed
zf96d19d535a99ba09ae3d7a1b35132bd9c7e63f55da1d79fad739a456fc6e8224a80d26c6c09d3
za180bd8e06a3a2d510915fe6d3758dddee024b48a05ddf095f175f89bc6d94846978ffbd5f00a4
z3630e03de8c864d09b10227b5bed19779a17e9b9f6e4106afbd3515f41a77ccf503f1f3be32955
z31c7ed79e75abb9d1aef0bd9b60ec2145c2123395cc110b976d9ee21fd911d51af3df255f8ccbe
z05785a91f36a116bb83fdf6fc3884303e6b307faea8fcc6c4f5a9b79d0741669f2671712be953d
zb281a1630414b11736fa583e6246447692deb346f617a7bfdd9c013b83f11f75e5ac4cf92b0435
z381aab02439f51a040e6d0f1a0e2a87614ef7a8199e486a28f353fd765a0012cdb55f49d11e642
z2a19016ed058a2f91b7db5068990137b5053e5439cdea6e1030b50070bcef4219913cea6978394
z1bb791d40d5680b5a81c0f3d19874007f127985fa70a2ba65a3176c444e40e65c32e5ca0c2af60
ze5f923c72c493be2d283683b0ea7d9a11ccddd72fa61777bcd223e14feec8c680b3d073c8d7984
z4e32c6a52c5f27d4f846464937e9a9c1c88df6f68b87422d3e4a4fdda07971bb3d0dc265e5e847
z18180a4cde005ab1e38e6bfcb1772da9d81d4c2b429f0033cb7c1858d5fe11c176928a03e2f5a4
z1bb3a0cfabf65a1bc9b4c9a504699e7ce353bca1733b3b6af2f0941c95401b45f73fcc4133db42
z339f301f8b97afb3f0ea2e8864942f8d3da0053276f29d0d06af75a96150dd8e974df06d3ea626
z999841158d354341cf42a2b5bf766d842d840dedb7b30ce5b86b5d8b33cc854c22f28c0c64a37b
z7eccea55b1b87d195e14270927a5e3deea13240812ac5a995aaf5ad5c1b2b6b4f6da92af286b30
z446a0eee936c16aa14afe433c4d4ed038de0a48970044f5d92908accee57d9be7b03a661a4241a
z4a61805735ddbff1f17c09571d16776750b83615fb1d2d1434ccdf370dcfdd8c58a94e231c0c2a
z2f0f0ca6d5f11b5cd3cd5df31543e7fd452e8773a7334ed524c66b71b3f6af137d7054dd5a6220
z7fbdd6b522bc0fd8ca6dc68a851bb137026b40d7154450d57c73c2ed361472e2c1fd86eea5bbc4
z2778f3726f37fa3f78b0848ce108de0bf1df0ef579c3e385cc865b1d667c82109957954cc5b3b5
zcef1863234b56cb7704407bd61c4fcd8b4162db51fec4734aee372c13852fd59ad8dcbf9d5ac9d
z97aba6b9514f5539ecdf6fdbd153429dcfa743be585c4aafb2f1b0162bf6a5d59dfdc4f86924c1
z5459cb4f5de1f391dbdb1c4f7a1583065f17596b1dc1cb903f17ea20830d0b244d8cd020d4995d
z09aae48c62f1899404e71c1de0ea56001ecc586c945a8efc8830688535606c2a8a9c221f30cc7a
zd8d59ae431c317f748257a0a0855ad100a6712703113c6b911bba1f904e4b33361799cc6290dfe
z9c5350f00c1f452f674acb8907e6418ca577d0d9aa715b601c445528b52832a71fb5fd708522b8
ze27107ee9584989d86deaafcbd582dccdce84bc737a779f86c1d2cf1ff25227f863ce439e5ea81
zc63a4d090b00e0ec24f2a06dd3c78c6b14fdf893cd296d0a55a12c7d2d3dc21aae5ed132feb269
z302cf0c6d74b7823d42bdc1836f2974ac7efc255a16b1c185adbb12b5d589ca6dcd4bf3d299256
z948f2a3c663d1df5d869fe5d3cf7856d60b57b12cfe2c37364b5f0bf6131e5af02cc2a1db05342
za295dc1cde44064829e07c13fdf12ccf3bc76cdca30350fd5c5f62286d80755ab4caef6989d7a1
zbbd1a134dbd87050e021cb66ec6448e80b869149f3ea28dd9a1003a7f890d4e494e244c6933756
zab8d4581d2f5264f337d7732d77eeb3e03192630616106c927dba35b94d90cb86647a7af47ab71
zaf53e7895fc4685a2914bcd0d68e66a015c83f14ef7b7e8327e1af7d4b727aaaeb62297cb97b19
za28a764062e1786462d98cfb32bb5e0fbdd548b103f6188536eb1ad97a5f867b12ee4a12d21ce7
zba6a716bf6d7cd49312321094b98c6691e7eeabecb4886d6af5d7509bacde4c18d953c57519070
z253bbb2c2561cbb1f013993c0d1707e7a2fc86e98013b8f3bb47bd9321adec472ee5d3d9fba32e
z03872e73dbe4c6323c9f4e82c32720a34ffe9212e90ba3efa41c4fc098996500d2945ee37f0d8c
z72cc54471360cc5c133eb91694c3b99663e2ed9a90c1d7c0875facba5de756673ccd790c28bb69
z3e7456acc551862c9aafc00e2b159999f0487a4b4f87b9f8435e911f2d753983b8da2c445874aa
z7c84e78818dcfd052a734bfdc7ff4e927d187223f5a775575f047bc522c4f4d8c2253e197a3147
zfca44b90ca6f97c7badf2ac8c508580d6a691aa925dc2071b5683c62a73eb9e5505ab88d490892
z984cff3a12d826af7e1460daa24f11a9a75e6d2f6ca920dbb7dcf3bf0a637094dffba3508641fb
z245e56194e11dd0ea3bd8c1ecd1c56f7a1e5730d3befdf213eeb069ac1c9bec060c81c393d6523
zb8e46a05369c9c5241ea86b90a96a5082114c925b6a1e7b6869a6d5b50da007667f2420e927eb4
zce548b50d6085bc5f8e906bb05046c1bc01d5edf17336f516ee572c833811029c2f5f8199a4ea9
z1b8fec212cc93be2d62f5719c56395c3dd2925db8a201aa7cf812aba454ddf02e7aa368a48f377
z553df652bb86434fd4215280cd7bb3e75ce9a7d9543d8c5dfff60ab6ad8404a6e470bf1a9b7eb4
z7a81abbc220d6d08d7ed06555fdc336f834d2186928828a90c0571f5be1bc7ed98cb0c98da7205
z70dd0565325fb8b108099a4de5d8392bd5d827d1d2a8e2b7eea110329725c919fbc28cd8dbf1ad
z8c5b40ddbee3cf4f3c50840ae6d34392586ca63a84687eb9996e82206cfeef5276de5154549a94
z3a938eba246741432b31373e61ab2ff99f158a6f460e95cb14a1fdfb2f530ddafd9fc91be65b61
z3ecd524aaefa837dc1579b65b0dbdc2fad777cec0005fb550fa0a7944ab2294b7fcf5a94478e45
zc8865d645bf21054bf9a37f22e00d6bb691dfee494d5bac963a6b176fed31da43178075d4f778f
zbe400531e7563d8868163fd0d40a866c24dc724b299b5ac298ba7e2bd070548c978f742bd012cc
z66e000bbab1f679da147ec1cb233d3396090f1a6b2c677dc3144361af57dab19e92e4fc18ee86b
zd3f20d1f60a02a01ff3bcf72766cf5d268478cb2054da796949e3037df3b7f1e978a41d870eb51
z159f26efb4304d139c4f42fff266d350319e3b73b8d710326580384529728a1e02ab52b6f4af79
zd4bbe5e2eb234be2ccd5d556da411f8f09206db49b9fedc96a26225965becfeb4614eaa6dc8e97
z7457f23a9d336bc60a8e97e0035a1cdccfc8a0b4671c9af692372a3b0b0027a3f47f798f6e6a5c
z1f7223197de5c08006cf30802df8c7ddf0a920f3e7e85d18d3d6ad62b490c804bec54f97088865
z27cbba1c0fb6de8c262031aa8b2d0c1d2824b199e8fa683d6c564b7d174f69222a28c58764fe67
z21054b168b1b34a797b686b85e3cbd39022cea9c28a6784742147e0276b89dd6b8fec690020382
z129a46253326ddd3ff2698b3097a74762c62a72d8f1358cdf3595ca04feda62dac7b4b92463aaf
zc9c74ba2a1212ffde9e163c39a6461f25f811aba60030426e4aa3ef436383deed87ee181fe1725
z2057807573a4cb9d9963ff40b3e28dfdb7dc08c20150d593e0a652cb33b36aabfbebde4cc5ecfb
zbba00303c66489a2253f9fd2428232457b285ca1c3e58c7655068f25322a1ba049922b12c7c57e
za96454a6685c85946338e77e417cbb63ff8a639a4fd9390d139f03ebb936af73a1ad4af12559c8
z670562c27d264be76a41b2a85a95db45aeb45644142c3fa21dda036ef3692e64319a5aa5a0f98d
z6c60b25ef4c41b75b15ab383de9596e20899a61f1e705abe4ad497b573d8401c600daf6be72d6a
zf33d41a6779fa2e184e8ab52dc698c0465948ba2f3be9c5228ad7735cc14112c4756cd39ae3c87
z3e418d9bb97b6c5faeefcde7ab7e5adde472f3fa37f1da34e101bc9e2a436b2187f2a5f002dbce
zb4d2be5c05ce69925467de63fb9e1a7a4ed69ef3414dee9b7608a5e0d787b01b89377463bbc754
z4ffc3c3d97e655fd84004470ea09ff3983e0cbb1ee11c18181c55775d2c0532ad0d4c395775d9e
z399dc1da20c35e7b648d6d087a00bb54cfa1b0b653497b81200c7f29d556d098f6bc3478d04200
z2441f209da6bec32f096fc3877f719c35d47b2a33e34b34bddc794ba22355279135d67ad51ffae
ze427a750cae1f8952852d88bd00f8150716e04cd9020028157d1bde7185c26237d2acacfda6286
z642e4da3d22d37a0fa1d9d204ed5e4a229cbdeb54910a0b3e427335c927ffc8f9d8ec0691d472e
z3df7ce395bafdcc080f187e3979d6ec11fd6bf3f00ae5ccc748f64915ed7ca10bf714fc2e23774
z2b7f16340027b9c91b3764dc8d5bb688bd9de2d315b7af2685117a7e1bbf795f88ddff38c0888d
zaa4a29e3af0220a53a74c85f75cb69899d8ef24c37c4bca8378d09a86e4db8fef0f6549e0e138d
z520f5812877929d1b3ca65033079294338149132cc1b518143a8eb3fc590a000fa54d35ab4f819
z41c060c49fa94c85b9368fe98ea270883029a18f01d312fae0f593159799f2fdaececb18e81cea
z683952290155840336c37ca154cd7c50f80e228b417c849c7871266a60e4a7aec2408644066b47
z7e51018e011a73a30126c9af47beb2d6625052ef46abb02a82be430c7ade4b68f7f1c552847e72
z16664a948941651b0bfd6db7683a589b9bfcbc39deb2b6b46388d310f27fc530f2a2d7f14c4e40
z7126370f0983febf1df5f382d72efb39f76143e75980e0d95a3785cc0c89b7d7b1e0875a6f6a67
za3b608ac6cd26b08481b77ada9d9903800e834563564b6a28ccc62ead0b47382a57e6a615e03e9
z7bd66d1e15fd8950239e89552b7a5f6e6408f6bc4c692e6fbfa83ea01fe369bf05cd79771a8a15
z0017abab301da7ccb6b5515d7bbe65c68a4747c88fb3e4be73663a5caa38aa67fed6ae473fa3ff
z44bdd85cf4e19fcfb09de281c7bd0595405104e5881f91885db28462e9dc6cdd0f452fb189a596
zdf9125fef795d4c78643aa479aa3560df522f9db1e5abbe9b97956f24ad84e369494dc298ea4f7
z54ddacbc1ccfd7ea92980a722960ebe1724d3f613df617100b6a78eab7017021cb9d03f49e9d4d
zf73cd925172c7c3ab9331e37c4048b219ceb82b2c3b30b822010fae81187d91160889b50a3b84b
z327f569cdf395d4080d0fbaddadcb0950708168e82c5a2a9dd6d5fce562e7f7018bfd25a54eccb
z70b00d9618451bad4f1823fc698dabbd93cee668a58dec479535f6e9b40b5102f06675aa5fde5f
z45d8d651c0d688e715537fb9c0c3af7dee0eb3ca0eecc6e6ea18c33b793b76742dd62622cbe502
z4cffd5ba11094f85a91352ba5b233e405c9aa63f55a28a1a7eadb9fccf76697e816bf35bb74ed6
z1f934085113518adfec44c5798d9a7c9f588798fd649e38ea478fa679bb3e0bdd253c709fe987e
zc667f49c6913ad74a4cadb6d8b245861d8026d8bfdef53795af2c0544fe47691095a05ad0d7188
zd41295c1890e86fa11b15aac5f9bed1e9c5eed695b8bfdce20dd3b8c9f57b1be1558e88ae471c9
z85a3a910181548b2d7cfd7747472f24194d5ed9d9d3cb70551502cb3f681b63b260fab010191f6
zd4660b798a83e9541c072e32ef493942082c2a7777dd67583f5124cf6d95152cb98c66e764e275
z352bbaf122ffeb86152aad59e4fa74ebe88df40153abf2a835ea710018d651298327d3ec9cd7f7
z856c8f55b2d10f96f4831c84ee96d8bacee8c6dda672781be8b5d120d9831ed368ee9cbf5af667
zb8bd7645e062db0040794347698e8cf7c18dc7bdddd95ea042943c71b394ef1ad69fab3d800f9e
z01fa60c1852dd010da74f9ff40b7b9865e175866fd1d6812d9d887d0e2dcd3593c440a996c0ccb
z888f221c36e118a18366907f888e69bb33fbac3f86036a5c5c4b1cc1ab474d773b9c7aa72bb3e7
zb8735b0f95cd7b7aafe57982d67ce37573b6b69a004ed4553123b52c95c0f21d684c81d235439a
z8ed4c27e7325fd6e28550c5934863757fcb664d71e7c88952da45c421faa9a810a1d5831cae496
za6c33fccc8036e3401f0280c464017e044a067c15e46ac91b006cb542d9ceaaeb03f46a7a27f86
zbeb9cb0f2fb69e63425222ceb58b1bcf5637d00132ac5a2a66b86f2a35537f7c2129c8f1ed9ca0
za974f436ea3a03af77d662d2ffb07cffaf007af9765cc269b00a1b8657028aba0efb0b2b53718e
zd14f362c9c1a5a52e591dc39744ff6e198b46fd50842ab50bda79fa083cc39baca72ecae464296
zb80661787c8ea9910bc6b020ce266326d526811795d1de997e60e45bdeae36768dfe4831567ee3
z0c33811bcf7226e888f8dce2a45b7e7a59751f209b89124e11822d912bae2557a9ee6387f20878
zb34ced2afde4c32b1ff10fc71299ed22502c444fdfa3d23a1bcd672e3e9fbd029a76c5a0696327
zb4f5f05a8611c05d75b7e025987bb80fa5819263f3813edc82f950adf42755d720b7c5a07a7cfa
z7fac70f89b3e2320ca622b5fb588dcc368903ad18d5c95c00dedffcd5ec4253e2a11b6a29dcda6
z4d3e3ca4e4d02649e911989f0a6b1556c25ea7b19b0344280d1f1acfefc3469434fd7c35d2ffb6
zacda52da6012276bd6fbca6862dee3df26877d2ba868712f586d9c69d1c525974ec7b3fadc072c
z407a4572d6e55016584fa3a779f89462f2993de94e328165bda48778f36791f19a1f21b4e6ce7a
ze22943c4db631ef11e51e121130ac7941e240ea2cfbf7ab62cce6778d375ccc1f8b09cfb4daaca
zd2645519932787427c0af048f3d36f41a527df5a12fa8adbb00df131d07ea33da2be2ff9845280
z43899cfec5345edccff408f69df4d49be6910e1c36e87fbc655a6487afade48c5fe2c886ba27b4
z296d4826e5b125cf1af45b0f4c802dd343bdb69b7d1dcd3a40b59c7365f8fe69c8f8754bf5abf6
zba0b6a71e754f0b71cb02a34ac34e05e701d6d339f25694c28fba1c4aa5801fcd25e6801b5d6cd
zefa1301a6e561bd376d8d141387610353e1b2faad266b99969df198928e469c66fc0f73517fd8c
z4ea2b6048bf81df80ee98b1d7d97e05f3cd445db67bde73c9f1dbe93efa259d80dbace19a6446c
z301f71c6feadcb745665623ae54c3647f262715b846066f62b4787bbcc6bf11bf6ab5e824db11f
z15e724422d4cf85002c886788f3f85c0b44141935103cdd238b5845e18c9f580b94e2d32ba0f9d
z52841c7d553bacda9ff1b03e523447fe7bf879ccb81a576453611c5a49ec6ffbf8ad1b8e3fd3ab
z08df64e5eda056dd3fd1de94cee89696fbe17a31057cfb708889e7125f0f837c76918ebd074f04
z2aab8d1a8e0dbfc13c34507ee23a918562b466f7bf360b0da9864da9f1a42ddac7824140f6a9b7
z0b46d8ff2feabb98fac160e14de751b70050d72e73acc5a7204e72e7acfd68688d025b1da0512a
z67478f099bf0c74668c09336536ac79b6721650e1847714928ff60c2fce3b69994e834e4cf7671
z3b76b19f671cd419b164bd1b43c0338ec18a8dccf3f65d4c8be67edfa352c04bcb23e399273cb8
z64a6faad619d59dc5de92fd513bb3780c32e8e623f7faa9460c26334d0bfc5c0786bb79027c8a2
z1734e9aa687b11d24ad649e1e54ac8f6f3c7e595c0f7f997c44cb43474df093a088373593a7b74
z58d93439735a92043ae09b97d0a89b66cdea328daceb4101752bc1afb64c59064dc405ec4e1056
z09bb679a98ee8499416f77323b9c18372e165d08962d8b9d874996fbf12688d941d83c1b41ae5a
z29c6f383194b53834e69a962ac3a4bc16e7b22ae3d4589448a8e8ff8e899f6d96e3434f4fbf122
z71964aaf74842fb38815b1a09276e82526b0f1c3dbc56115e3fd4197ce185f4db0195956f8dbbf
z11de360505d2316a5f80ca98160530029d533831c0cc024f4ce0a7561248f3f2374f55358146b6
z91234461948f6166f53cad7bc8e748c9b1f82829af4db22797db42bcd997a3ff66e7258b515c35
z325696b1c314c868ce0d4eb90eef5c6283592a59a7f17d4fe7a60bc516ae8a995dc365cd819dd8
z7a3c648a8d74ec276b24402ab5460eee8f326145983b733bfb2b26753e785e6479bb5d40e27b1c
z58f6b489d1482ae0375f20d7a3b5ca0af3e251fbfdcbcd462ddd4fb95df62adcf227bdeaa0eaff
zba6a58a531ed2a10042b2d0b492b7c94cdb4cd295aa870d1721ce94272d1a28c91ddee0c3cf1f6
z76fa667608fe37144ea3c0d4f1696745cd7d7d6b971639342aec4ac35b5f7914f446490f96efbd
zdd5d5c92d7880e2a08afc2cd8098255ca341e9ff3068fa1707b9a0f9cc4640dbd3d640129751de
z9f36ea676fa0647ef66fc789077e81334e7afdcda905b12809792f112d1153946c7a1cb5b948ef
z8bb304643f970f1e1f7b653ee4f2e65bf91322f7ab87980f56539361c30c90582c107dbb0eb2d4
z0dc2b763089561e1904d7503cfc84a79f55e39b073b80180c6c76dcb577f9a92d97d5d3a12af59
z6d34365cf70b76091b657dd3594c0dba22869cef1e113749f7b9466259ab6fb581c6ee55035b95
z04679e03750d65ad76bd5ba945ba9b6ea3eb08335149edf42f30e2c17563022866dbf894d0f816
zb0c004e5955e7ac6c0f603eed3643848f55aef4c308ec34a74ee9e2ae94cfbed75757e6b615b4e
z380d6b003580ca600ea06478550a0ab7626d3e423f93d43e3b4c5b429e6aab23828f9f31fb608c
z7da8450332b692a16c36c9c07124ce2ee6e1493508c40597c4bd5882eb5931d490df863daccafd
z9bf7dbc82f121326c1d24cc6b6b089237739e05fe49e7340f12b97f93111bf80ec0fa1496689e9
zec96241930c7742bd90a6c8a5203f4c11742d13a6e7a72c4ae6894c32129c8f86a54ceabbbae6d
z4565d5099d3a6936a3f54387aa69410317ce30002df90ad1ab2b90e748360d478cae10d1d45c36
zc12cf4f9589fa1351e6237d5ffba465e79b786e44761b18ad5fddca1d3790dda40b37ce4b421c5
z2efddc1a485c19c0fc0c99d33fcc415870c460e4c90599ac0946d0478a8100371bc459a4f20b1b
zfa5381e5983a456217085bc56f37bc6795077604351edddc657209c509079f5b2c2e3c5ef6d9fe
z7387fa1bd5bcfb4a3a7f127a7d01a83abf3c98f6d1424a6381461a4ec243e83d7973ce363e9196
zf5dcee44a9a01f81b8d10d5ac1ff1664647c9e8c4dfac001daf413d3f33dca1376101787ab3268
zf7882e2c95f8459173be35743e7f33054147cdfedcc882023758bdbe9ba92bea4e89da592d1d7f
z138e811d171e8baddf8eb9f52a490a78ff870ce5245958f37b760f2c537355c171ef08d8e1be8a
za1282e5f2aa7037fd559f31905e152c348104c5b6d4d178663a31d5a0a7c77f9f025ff3f316f24
zd3453e9047543f3dc77d3e0d32ee82430fe99df75771c0efbe9be520ed5c78e1454b7ec2b8d395
za2f6a4f7fd5c5f123493849416058079c2b057c766ab664ea5a20596683a2dbf9b84ab9371f720
zf42d6b3a181cbbd0ea839eb3a022cf1450fda8a6c4e5402ebb78d6b79ffbe19b9f2589c9fca2d9
zba93953a568553da97eb4b94fcde97f5b70a49c13eb1180be861afb2707c64b2c4cb8151f66a68
zfeaa0b4ad6f40ff8929a12202f25ca60a4a961ea6be772402f9787096a891e3dbcc89517542db8
z472019533b86049571878506cfc367d8083a3339332af4d4920f691bf8ddeafb31342c21b95223
z0e4064afefcb91959a89d3c2e3926d5b850cabb0e07a8aeb0903a8d35d27089dfbe6727c848b1d
z38976216a2c7ffb39283fce2e0ab631a8a48961dcda66aeef085ce40bfc97953e31f682f40dc33
z89cfb8d88bd8ff0bc2b44c7c9f2033398c0d57692825361ac8bad649a829cfa7a7154285542cda
z2168a82f03a6669c019a0ac68b56cfd63b547493554713ea875c578b01f4fff2a984ce3d8d900d
zbdf3ec7500b64e800405d5c8ef9a94e2c2dcee971b932b0ad3780752b5174d3a9e312f4919984e
z7a2f9adbaec1c88dd7962c3580e326551635b457a1fb04d504a7f84d5bc3284c11d19b24bb5c29
zef3ff6a6e5a829ffff266d7c1288cd8e70c8940383a1bbb56c0a29f0ea63a97e1619103a087948
z565cf2736dbd923e59caa1b4508fcd8f139f28bcde33a023bd2e8567c89050da4f9cdb7108ac1d
zaec11860e30212e1e7360cad020995a4fcbc8326b6dc7a60813e0a0d2ecc37a51f0e6b0ad87893
z79d68bb3bf6cf390cae9e0b683c7c687e0294b6d3b15a247e838bf781585fc7dd89568fadc31a3
zc4fa8f811691cbf37f6f5a6847cd40510ef93016471a153b1a843e811d10807dc1d87d7b252aab
z9e60603dce5edda295009c4f5449fee68af6e2abcd462f064085433d4c949e95d672db1de8aff5
z5297c7623ce9d7f6ed7968549d58fb826ac196bf4e60973a3f4813e23ab0ceeb73704e55dd18a7
zf6b874b4ea0452463bfa1e110280e30a877fc6dc877b7611ff72d6da373a191e7cc298c3a259fa
z03fa9c09884588a5742aa2c8a1faaccd7f0c63b2a11ffcb2fffb787994ad8d991117527b4f82a0
z8138d142faf26b02bbef24da4124263073c488ba3370a4c36265b26b7b92c5eb30b5164c27c584
zd46b12f21b0fde9ed3c7c71849b73f0e6f372fdc4794ccd47607e01674c29eabad00b087aa1cbd
z08c5ce994e881736f29264255353103bd11f731cdd47be9a0e099dac34e6d33959ca4772ec73e5
zdcc0c82c605561ea24bfb8433b1566f1299d129afcf72a208580080f192cb90bd4ae7bf98b8fbb
z99571ba6474eeb6b2cb8da17b28a5710bd41aa45357fd6eb2843bc8bd366a5e422c556c09bd392
z2c7575b497e5308380cb92380b3ae8b7613c482eb200e2fa9f6a5dcb7463a4fafc2ce36e9c147d
za360a4043626cb9c3a8a2e08d7388dd6c0e084bfc29df752b1443870795207277f5c45bae70e20
za41c20505804efa200d7aade1b068c4bbabc23d2dc1b07f21200eb79e387625556d73ad7ef6130
z45a2dfb3123bd58949b8157f0b58eadede8d9365841798f924fb4ec13e53a1ee7d4ae72978ba03
zed1463534b58b0bb4f2f28b8bf5c7e2eb7c7fae1027a68189b5017c15ff9b0754562dec00d720f
z33e7d634e82b545d032ca9a9744c18d48e54bf8bc8682779579408b4560449ed1525b94f50038e
z04e1325a3aedcd3caedc1fae5c19aaac35b5b29ec4ae183863fad41b417e28c317cb7c4eb7fb2b
zfda492987b3d1719dd2dc5c2d27e83131d138b89d75989a6eabecd59a544036fb5c3b69f24c790
zee0974b7a170125b7574921ffa55ad7231ff97dce44ba91493cfe30174edaf51f79a1d3a231a5d
zcdec629c1c30758e108bb15b05a4ca6e39679c6be6b9d991dc226c3c9ac52ce2410dedc2d408d4
z808018f9549af2596d90d093b4433b4ca49bf53c684216639f0512f52d2d485f39d5edafad1378
z18dfa2d735970d4c5bc41ebbf85c5022bfa75a170a0905807f4147c7e9ff312a92d1797cac0808
z8be74e6c02b90033ba1d19d1b6ea06af4f8815f6a9da5477c9f8357767a3e951007295647089a7
z426d685019cf690fedc41d90f694baf903436236febd1a07c292809c5d9961f5a3ec073e95da57
zc9335a4a211a510d4834290177948c5251907e9e9da1f21cba9ed2d5fcd5c1bdc1097a891d09a5
zde13e1865e274591b04777b66e73fc48ccea0ae166dd739c12a3b9f213881818f8cda9ccedc032
z2e929b83b7c4a123edd02d3a6a43057ac0cd284d5ae49628daccb904cd9d11cbd1df923a4fa18b
zcbf4e7593d09e292d43bc4afe444faafb6d05d9ef9dbd41fa0e1f0dd05d31bf92b72172bad3fb6
z9ccc0d7af2b30971e8a7bd94064c8cf714e7cc726f7da0a849aa925324353687b66cc4cb8ba4f2
z06982d3aa32fb9b376a73bbaf9ff86a28576d80cb13bb3c3a8d6645f74cab9297c6b57673cca77
za8aef593c8b89b8700c383a4e1e7e1bc15af6e0247f3345f1b613eb66673c0055e7874cda708bf
z531596398eda8af43a9a4c75ffbc1550f6c461d19953f0a9031d02792834ab40b2024254eedb2c
z0667988bc355688f5a882a982acfb3ae80a904f7fe8cbeccb69c203989f3d71eb69d889e320d22
z8ab243e65a793a05cb6bf6743d6d2767a2179ae8b99f212d7682a6b785cc29bbf152d2acf75b06
zc6143500257b7f4da77da992f224b639e3209c6312e50bbbecc95fcb3c0574e181f39c43361ff7
z27e94dc459c4abe075728f2b4e3024b00e9f1ffdb0c3b0d7cca2a2f9a8a16b7889d865cd64f5b5
z85bd3078b97726e23c629724fd4d0f2a7cea8996e4555b1b4215b40b6c37359f0473adf45ed241
zfa8f7d1eab1e74f0ab03a7d214ea4b00afcf39f2fad40a80d66708313644132dc08ea73234f10a
zd08f25d7669db9453c8c1cda17c84181d945924606459c87c76581e414e5dbf74db16898c56e64
z9be12c9d777641460bdea01ed2369bb3c9f7d1eff32ebe47bc68c4c93a382bc9f33bee1d2a8843
ze8f0898aaa1d37cb279dbd183ab4c6df1a9e046bcf33a5aed6e391dd728494dbe2cb6cc7b188b3
z90e17b48e5e3cbed8c502d7ddb1efa6500a6fb9270e1bcdb2ee0e1ae3b2ad079db56279e289f84
z947cbeb88e9b2e4b828d12d8b713800eeb92174a08b014afe13a1db7598da8b360bf299cd0bca1
zf23a8032acd58592766f4bb1b1a86d69878ef45b0b0f0d38e77f099bde71af07fc8e068ca776b3
z38aa54ee11c6455abd439118201b3173ff07c5a8c57ba006a770f71ca130179984e5581bd76062
zdc0087f90938abc36e072bf88f08f80d12609b9b316f9599dbc1dce2d0162e8c604cccbb4324a5
z08810738b10299d434f34738e80255dd739f0e87dc6ab74e97c60106b26b2fa5ca470d23fa916e
z56595514a2aedb84414da8eedc52543b3279c394ebfa463d417cc7d6fea106a3112fd2426210da
z27d8a214708457bd27d4627ad24047f01a5e380c184d8ef8bde1eaa938f4ad3aa1a1cc95a1129a
z1e34c51fed508b02f0825558f0757a2948fe32c1173a0eed53bb20fbcc2da94149bcd1464af344
z04dbf3d1876d088203d819c08a25180ba73bf92295cff195e48f3c2b585a60fe474aa12cec3514
z3e22f4cc9c1d9a55beb770d1efd830c88d1a13fabb53e070c4423c3b0f5ec92f5c38a94573c670
z1827f4a4d0889b75aadde5036366c13696293dd1d1f11e317a3dac955b92bbc8f06b50a05654ba
z2cd3b938dfee1ef56146197eeb8b3fac5481cdbbcdc0fb3902a7353484d8f8040b54ca4a738756
z243e3fc5a7e56770fb67b93c33fc24eee9d068bbf671d44b385355472d17b76006c671e2c046ee
za5ab34fe6c766134d9f4a1dd8784c6e0412168a24ff744ec22fe349cff68c65d6879c4be2ad5bf
z1a5cd6c63c174c6116033d168e78f308df40321970cefacc391b8585069c1036fb93fca096f0ce
zdfae0063ffacf697d96397fa697469a5f202b80ed7d3997e6562ec1ce5a09a0dc441e6fe5fbcdc
z340a06c1e4ba7ec9f21e4bb1a39edd3575542434660252edc4a01ef1fa30b909d997eafe0bd209
z6084c9752d137c7a5645f1a405ec4f9ab8d45fe042ae47c3d4ba6e9ecf04df84f43507f0dde6ee
z29af9c2f8194dd37da26f42d9b3c8c58a4023f7d7e7a0217750fd43d9e7655ed8fb3cb06da9da4
zedd898697dc24aa205a1e0a3ba599f596f33462cf457021a12b67084b5290f0c5f35024b87548b
z5d615497e192869cde65d0ef4e9d080c051d126170c89aaeff4167428f302863cca91bba85dc6d
z04e3de778831b910c7638a03d98c73a253f3db4c939095cf79b68cf00d440296281bcb4e4907e3
z5084b24a5e07a80c1d55053d1514eec4223f24383d5a524119c751c5bb282b7034907436e5e072
z6c9e4648e39af4c7353a6e837baf602b5b0ff07949b8541b7de9a29129de29ed0d49d065f359e0
zc2245843d51ad880a1a9b87b8f8fd1a4cb2f495db838c1dd35b6de30e6e1324ccf03de62130157
z9ea0b508327c0c4b8be7a4cbf41efbc2a2bb402738aefe4aed49ded981ca79436db33480cca24b
za79713d379b95d9db2b53f8ff0c532f17b28034f58c891a9b09903d859f944c00cd159db0fd719
z14dfe12f2e0eebe1f5aa7a3a268ab33daa6e1ec35eabd644c9ce22325089448b6cfdeedd8005b8
zebbaf4014214870b7f43df7b90d98f93bddbb7ff8bbb3c4bdeb147df0c2fd7ad59525bff10a8b5
z4aa77f841993b648fc61ef3f0d98d9714f653fc777a504e1907743c11b837c75f2422b34f33206
za2821cf95985b9f0fa10203abd10f1522eb66f3b41cbd7e3411a9e5f3145ecac2c9e86f373f7e3
z1fdcdb071c65f5525441385154e84aa7a9b8113bec1f8129d4a5a1dbc0afd72bedadb06ad4ddbe
za8f57f052b0bd3f0ca23205c1233fbc44f46a093c7e1a974ed976915b4b1f4ada6ce3ce04da17c
zc360f6e63cbf7cee03b8b0847a3170449952a0f6836ebe1bdf3b634b207d197c656ef4be717ae5
z8d83eb017443e6599cf31c62ededd0d9d38b71624283201fbdbe012acd6065a9fc7340d000f55f
z13a01914642892e49970571ddcb9aa321bb11a59d5672969a0e20fa9642c76d5c6e8a712f52e79
z26ff20b3a1f52b47e47427af775dc01982813590e0389bf88d686f74534d27d369fcc4b6eb5dcb
z4045b590657eac01a6173fc787de88323c7d9f52d4e39f797a0d7f07d6f8913d62b73249634f0c
z8132d77919082053031a0d8681055ac33bf79bcdb2ea8e7b1a0b81573fdca8f32b3095d1337905
z76957d3ebfee094ec33f2b0f2f975b1e27e29229814e2bea1c1bccd5aaa76428979ddd6b1e42b0
zcb3299f0a9eeced55b98e10d93594912c451830cbfb2f5345374f20a65d1adbe629ff51d8f3fc6
zada41ffaca81f029dac17ec1f3f88004047f5d5e4cbeac7701eb998f8e1cca046b772012fada90
z72915d61d0075c8dfc8661ae11faaa1ac17fe0bc78a5f8a838791c1685251024ca4e123e9b66ae
zb3511096c2bbfcd8a40f6c2cafe04ed5a3e5368dacf81068276b79a61db890ac35c8fc48a6b37e
z397b9c2ddbc82a0c6d2d15c4e0afdec03023972425aeef8cfe95321dc3a801e311f70b4ed6ba89
zb71a5723ded7f8a7f1b9d2173f8842dc86af76c8e94a454c9ba95c1b47860dd1cf17ad51320daf
z4a2c292f96a823350fa0f5fe5bc7da32fde1347a29eda8c815646700d8b332715d1fb49f8cbd56
zfb2db3f103a9e1ba11ce3a1a3e35cdefee0c16997692824bcb956c23214e5c796f9f1d1f74ba12
zb9da248dd8154e021158dbcb50956f235856690afbfc71a89a91939cb3802010d46f1c021a66f5
zf41f6e62b4f1a3fe0998c8eb401b7472530a3ba38a4efb7384b19c349799ce49d8b8229cc7108c
zfd90ac93665dfa29f1c49eca1b8b7d4f8abf40741ad4c67a17d98e5d2ceafd33d84320e48346a4
z1605df2bae5f88695d97e25cd0b1fd5810391300edc956dd9cc41856ccd5ebb577528646d13306
z36975c7408bbf3d12e5a1a564029bb2e34306f9c50e4a1267bccdac4683ab4acbdcecf7b2a2edb
zabcfa610b6122e4f173cf8dc672bbc3d9dc46e149bfac876e019cb707ead0f25fba8872a795a0d
z9ab7422f906b964a21f68b99fdd9a7042231757c2f43ece394f4417ef40bab3c1f6858c1f88791
zccd53113f66b672b090cdbbe1456c49473225832c3f5294d581292ac6db4782135a65293ee46bb
zb4687018d13a5ca068a4ef1a07e156312f1ad0ff432762e2821abea7132f3252294d562215d71f
z4d6faa2547a47ef1de160b48aebf70e1f51c1687741af46389da003214f8d18aba6874edf79af8
z1bedb38d60f783528cd48091a7cd2be438d8eed2cb5ba29374e4bd588bf4d14ec858f626ba9e01
z952f25d81e5692f3591502224b1e48f64e16ee192574dd9c6a60add77d12068feee90a05127361
zcee625ed2f0cac2484edfb3299ee3f99187add5aa59c1bf4ccc9f1bc58c2d7af725253ff3ed780
z66381549abdc3bf62c6894465898df27897045597bb7e06916c1d07f06b88bd474391c8c5af9a2
zf53e7bd22fc5f64bafecbf3e1ad6d94852992631319421fb6dc66f03f2c3eb3bcab85d371178fe
z68766a5bcf82f2c1cb7b4889ac997f662ae19185388383468a7a6c409c867b7504a7b27b106c39
z93dedb5612fad76ab8564c704135740291d8b19a566d3f2ff23a2be14d3fd661f5086163b2b6af
z36d30b5245243c9be98e7b818e07b23be8a23632ce2ccccd01836ee815aca0218320b1cb423abd
z05137bf199d74e425e7f6deb56659fe12e237a18679d3f3ed9141abdfbda167a70bd2e2fc77a93
zbb4ba860bee3f14179078ba12be30e8af425e508bb6ed2aa335cafcd28f2d84334dceeb7fbaa28
z3beabad34844cdbaf2f0d849017f89b58e4333c6411a3b9268fcbe61fcf1c3b90d281d7900a68f
z50bb5dad6067e7976ddf9cdc55a26e6c0e2373085286820c2c172cf42539465e34559d95d7103d
za1b7db72e516412bfeacd317efda1f90d7177d8374b831052c854251ed533231c513a59504b108
z07d73449ef8e940c7aed804f9023833d330f26375bb464a797a10d5065dbfce5291e147f3366ff
z56aef06d48f848d19c3b39554b83a6b2539353cdc23cbc140f196df6edf46970a2622d1e71d19e
z7417f3993097c4237be73b259ebd03192ad7ab96ac65af211ec22e3924f34558a551e965749be0
z207bc6d0b7fe65672737f790df882731078f85ceaa3adccd010231dd9f29a07337b7fd7a3c1034
z33e30061ffd78c35aa88af42365358cc8a21aa1712da7decf9ea28566281dfbbb5582f54b0c078
z573fed807480e89edcbcf1ed92052337cee5d6faf75aa06a66b03652f16da32fd8e52e7974a1f6
z5eb3b802a9995cc37c7d20fbfa125caf21826e5461a048371c427c1ea93ed96ad2c5014caaca4f
z2ec47dd0bd09bb2b51a378dcb2e2792d675c460a1c76ea4718b51eca81f8b49dd4bc2a8016cf1b
z1f658682fb73d45df60a564da4a5c911f1177413651e6f41d022f250a788c62a1445ec5f3980c8
zb05dca617dc6500b958b604eb29a870086ee8291e949724ab50afd4db733f5b336694dce32aa44
zb960ea0d14501877ac270a8b6f0619bac848680ff7525d04c10715716aac4293ef59676090fc2d
zdf37e2a1b9c0bb46c469305287a8a149a7469364788d96307c584e01b88369c8717b719590164a
za24b74c032ac00b9a6c9ed8bec0866de500626e411e2356e01e0c1bbcd8922ac8dc5c22866de06
z467449a167ffa2ed0562ed71df47847bb2e469dc3c988e4cd69b9be7fe11993b7aa4c9660f61ac
z81ff0523c9cf458c2c5342c2937a5cdde90b051a0a4b463c69e102396a496b5338fb5d044d2360
zc3bf1ccfc83e0277d4c9ef753b5317821e5f66c7a9528dbbf3cc4e60eaf52c3e24bc11c13710e7
z3fc3807b894727651a5320041551b2746915386039ee900b39f4b69db121692941350b54b0540f
z602f34667b2e9e5e01b4dc0fc2ede50ebe8aba397e2746d89f484f1448478f5daf3110d751857c
z62fa76949a8bd2662c5ef235f0c2d10f2e63970128b770aa7c508ff7dc1ec0a2bfa2f31ee11a49
zf20c57a1f00495a11a1826241cf0e00dbba46b3d5e18b6cbdf1b9c926d9ad93767b95182032753
z80baefd8e1b0202696fd3f59ddc8012890628dd207b3ba3710db84e8fd039bcdc8e9c2fb83cfbc
z55b6517b7057a708125293eca5ea0be81d83f82b2baa7a8d4b950c8d4c2e58a70fb17251f3114e
z1f20c830e9fc1eb788edbb65bd67a54187d68d271a1a6b173c7108e3110659eeb8cfe102e2af3a
z6071c094a47ff939c5a990f4033bcc2cd0fc0303e46197abc611f0b8ea5667b826c7d17b25eb41
z05087931b68ab36ea62e3468f34cd783de5972dc8d2d6f8ae53c82d553c6fab43303cdf0675c01
z1b39c1d6ca551f70900cf319c74224edebdb7ea3c479d28a98bba68b422ed15b125674de7ec7c6
z759e09d5fca10bea398bf724c1392dd7caa77af4070bb2e6ef1348d751060192e29785aa56d49f
z1d75ee6f193aa8aec7c674980cfdff67ab21eef1d905c7a2c666c5c77bc0f059587231e85fb6df
z3e0e3b7df259b28ace7fd75395b12ef9e4ac7c58c6cdd7ebb80b43d4a502c107f5bf2ee497e22e
z84ca6de2ce68fabeb35ccdd124323298f9dc063e11585430f3fbc6169a2dd955e8ab424a4a1c49
z13b14cdbd0b0abab9bcec46cbec21a7c8ddea9b685202b4dae0d8f0311c2b8cad37d35e75d6c3e
zbadbb20f1f75411242ccb5efe9971fe4cd46ad4fc87f3ddca25ee0877de70d015f1b55ced57a09
z80b5062b4d4c4a94f7a02b8cdbd34640620a0380636269145b677eb32f3aa5ab4bc13d7b6cc97b
z33fc9769657ca6379e499f3680f2847610145cc1ed55e61e38c7a7f431bcc51debf74dc35e7f3e
z7419ce155577dce4f71f32be5c4dc46319265c27622a6f6becc5685d7c2ba1cbbec7b65e7355fe
z4f9e7143070babfb055dc6c9c13518bf84e73278807e9c37fe0bff4b0137db5097eb1664367b67
za573d2abcfd4f24efae1d73806e61897c362320f69d4800f367054e15543f0be02dbd3fab9bffd
z0ff7dc8b8cfa4cf2b02a5cc51412684eb537ea182909a39237b2b30c6739516a7c2a0e6788172b
z7126cf3a3c0bddc08bfad401ca6ae006daec1f6170dad7fd5e19f0566c6c1f27639641ae302e08
ze508d444b40237d9f9f0344053ebe38e99e205c6fdef53a24a5ce9a748cbc73cc61b5eac98a5c8
z11129826737ce9a3ed3b7ddea6e1a025648c4421a342fedaaed250a79baada8bce951e7d4a4492
zfb46acaf4f2a5f1d67582efd0e2ce5c824fc524b8ba8cbc0c3983f51e72ea6f56e8ed422a531ee
z3dc437232d996043019eb8257a1d82bf2ca0ff23c57cf8f822ca15379b79b83f52f5b0734c61f5
zcd20701256f85f2f7a924e466e909ef5fdef62e3e6ad54d18217b78be70cd75aacb79b7fb42109
zf842db8f8be3074d08e98fd388a5a879f2140840eaaabf8a829a0dfa0ecbbc5009441d27bc3c30
z1b20f079e3e21333d775cd41d222b3bc7e454c15c7d2d47088ad2339d5494ba3932a4e544c39ba
z235a99e5b7f86d76303959c1e7d445be161898c35b6551a25a07654f9985c9ed53a37240dd1984
ze2bb048703e0c2571580a96dd8014111cdb1077be80b57ec858160d407e2a110e72ab8db523534
z2830f0a1fef55a2b9f1f333842991f88277702e5a1a85922f971956f50b096ecc4cf6e68a24468
z68e869b5c32c1376ed9fe34b5bdb18ce0ccaf1346bbae6a50c6b29ef6b9021b77cd22f04496af4
z6d24727d47d9a07bfe9ac8d9743b618f48ca5697c9331aa12df037cedf4332799b08a651b7b398
z393083a920186a70f658d1718d502c36a5b4f5541d6bfd6582cdbfcd337a403d961ca6683e355f
z1a3c3ca9a9e1ade54286213de94ed3d3780588e41e8e9b42e587606c71226a1d31b18bdd4036a7
z784fbe927d47ca245b5877c491b348bce1f99b7ade520c6888e3225e2605a7a769f57d83662c1a
z29b5554376281d9106b8b6d2c772651b073ba3d1273ff47f98c8e1193e87c8280cf1a24f07de16
zd5dea7766e1b61cc332a5423cd7d386e2d949a97dfaa9e75bf797ace968b4bf04f57a5e13fb247
zee2befe75b64143453b8aa4064d8bc8927c8c5b363eaab0fd94b79ca671a075e45d1ed6d7249ba
z446ea22f3d1abb659322f18d471d798f06989524344c4c688c2f98de8a890c061ca664ffa55413
z70224085b29fe9c6d42c301ec24da0fe1ed14350e8cf7ba09b64ec2181f4c5f3fd85ed3ffab960
z534aba2049866d88863827050e8234c77c0d412c602d56f355e2fcf1665e349e899dc36db9a3b3
zd9cdd41a97e46bb200b5bb2b228708751704aff1077258dc90012521cab8373c09cc265a536fd1
ze8f3c7a068a57cc8d0ff353929fe1ec6e1c05aa903bcd87fcc0e0439fa3973aad131e2fdfea165
z1d54ed8f49e288a4d4b8797530bd0199718de0f7659aaef5fb91ffd5d761830d6a4d97ee3374d5
z05462dc72960eaa4c4c7b26ac304fd7e94fa4e1dd95f43592b650f0496be424dc5fe062f2fe1e0
zb92d3aa9d8816a0449ada71853d8845fb1346b5fc68c3940543995f47ea220524c3a04d1c0980c
zbaf3eab5bf303045d7ca27e04e4d125098d9052334fb7e5abfdb020ab992ac8313ef17b4078003
z97a1a0fc6a8e259ca889fccb94033da0bc9baf0ba6a786d88705ae5c227ade85d045896934b57e
z197550fea781bde8fff21d8246f755f333db43ccd32765581396850415d4cf927f32ebf63c5695
z2dd70875f9cc267e06526d3adb0aee0b63650c4b558b1885f9124baadbdc576c5fa02893585583
zbd51e8ce2a678cc9bac37deb8a64530b3ef7531225cf9e2ab315d74500c51524266e46eb2914ee
zc23bbc95d37012d62e1c81e73d0cdb06ceb42649bb7f4d2f85dcec94b7897a86fdd15fc17e56ba
zcc7eddd10c87d2f16cda63adb229033c581e117eec4cc0c32e3217c12a552bc4c012aab7710530
z74c6714a4ea6031d28dafde3261140630b1f9df686ac4ad431fff9ebe7558f5a66c36fc51d091d
zeacd2d54c7106eb0e46ccdc84cd49c96b11ba36b38a02a513984f8470e87f7b3da8a09c28560ea
z15efe3ea17dc4ec6abd7b5ebdff07a9050a75e6d37cdd0983f4873557495f2a7a66a02b6f7d985
z5392bc3dd8d3353a04d441779b697d0ff610b8546f1b2013c155723c6dd90f21727cceb554e421
z0b36cdc1df7095704ade4b010df5d2fd0899a091103679b50de549268b40637f2d41377fd5e316
z90afd9c49b51f1e1a7a6f6498d3c86acb6d0afcb0b283d031cca877464abf0be4cee36650d5342
z0ea144169cb8d5715255893987c8a1f33f090288de50803ec90238f7bffa13c05b88d510486688
z3d437b00b4bb779ea8f20c0f5c7a643f83d3f3afb2f70ca39bea5bdda1ccbd8e5e4cad6d640616
zc2cbefac8664d33d23de5080d197f8a5dcd2f2aa16e4e11e6d29cabe5b08fbd130e5c9b8465bb1
z5c643ad491c85bf7af22e165849c5fdf9cdd9d3faf262b866024cb1ac95e9ace713c09bdc6f47f
z44d99cce7e82ec195c2ca05ddea1e95a46e4deb86e418552d66c69bcbdf0a09178bb187aeea125
z4d8974aa63b762dc8cfdaafb696ee42fc1d79182f7aa2e9519561bc39f7104ddfd0cfb8d4f285f
z2a2bc525e9a019ed0eec395c81c72ff62adf7354032352eb789f8da70d1a40e68d22b77263c174
za8000c015cba170ca61a4950632ddceedc75b0a7c7dd622de2f8f75d03c2011178720e6cdb3de5
z902d95fabd4b08e5bcdce949aab9e41f04bd76a5efbfca621f1417661cb133518c5d908f950e1d
z58d1e4245022e8d0500386943458d71024f861dc70889d20887434d16b2e7df26d43782d978113
zcfe880769abe647d6bf91081793e511f4901f309072f26527fe2db048497a10dfe23e6cc54d6e6
z5b505fa4613dd4853bc2d1e140cb7af1c17044a8531a6d53d75d51a725ca4c1fee3ed90908aa86
z3c9a5f6f73f56a026a77033737aed3773d4625fe6729e61c06c04e839e558662edad168aa41cc9
z9877eefd6215610e9dbf67cd8c1ba7bcc49f3d5f9b165fedef069b178c67f50ea1e159f0ae6aa0
z648b19332af27dee4a0602fc6bad960875a173aa5d7a69b426e458df7e41081a0d13424f72640a
z4f7ebae8421404f29b8da9b4ad87a25c3fb56d2d4d7a4d2303b5b27d89109da4d64fe173efc37d
z38d06b66d071422dbe9b7092cba37a1bc761ba1ccb6d5ebd9f73e2c6b05a5b0796567326c332b2
zd4d0585b58e9961b59537993947b9aa32b87cdc79cc70c28992e0eb4ada3f4451188ceb9f941a0
zf17fc8c35dc82e6c85b6592a4a5ab598bf7171e0c3c0f3f6ff61069e7c5849686f8fd11b843d86
z747da124228d6ee0ae5a0392b355aa3b636a00c3161fe37671f1ab056b9c7bfb3689024a2faa44
z923683dae804b06f7fa7f3841ffb28d125e0edc54ced78882e58b6967964cac625a84a5d654626
z7fb87791d3ed097099faa1795edbb304932fd8223a417c29d2de813e5e2b241e9f0e92151a6116
zd31e29f258955db6d26a2431b8c68b002d76e5c0d4b7aa09f643ac4ee3a403ac1f1ad50fb715a5
z29f7fefbb93dc361c73b113f23e469c094022a28a44f52ec6a95272a61f175de7fb5403896f221
z7efac42912f35ae3964f92b2c99e57295532e866968b3679c77c4747647ed79ed10b3a1e15c4b2
z5840bae9b3d9126478a3902b77f21ec7ff84b6601d1d3aa9e22b0e4bfb908e9258269eebe78849
zddcb6410d7e360a26a0600daa328b78fa0e0d9b2ddd17cba72fab7c19a5122e5cf98c6cc2a4a25
z3806767653adbd3e75e7b8bc11ce3fc4334a7d9e97db92e8f18e5a55d1bb93306b99abc5b9e4ce
zce7dc3061f9ed513c01ea0e5f87e9c0f082f65d64679a2575372a1cf012752513b1c2d12a28f82
z02a63994a7d850bfe5a436babe7ef98db91061ce265d8bb0c5a755e23d81e78a09655390d7bfde
z7963c1aca9dac5fd465e4f0ddbd6c91a5ce6a5d628e0d731ba31cfb6cc342742eb6ae8162704cc
zc0ff31011015ca77cfbe1013b365d73eb366f88c4ae7ef9fc4d9926051f881a6a5a1b65bbe9443
z316b30d37a3699c54e6ea87359e838984bcf4b8109e76e23a23304a8932f3d119845791b01b92c
z34eea098ffbd8cc6ac005d4a93ba90a77187ce203c251df8e71a5d12ccabda8f6456643ceae5cc
z0e212390b0fded875e604c34cb144b7a53be3a0d19b39db42e5fe1adc98ff0d68b45f29ef19264
zbf6e2ce2521c80b4381d89ce3a1531c7417dda6bbab2bc23d87149eccc14fe9f0dc92c28aa1b12
ze6cf2a26f1868c12310ae15af19c5c599860fcdd57ad8ab810f5053cb666796a80774b4cf73ad9
zc24b510260e3937f376a009b0e5377d27e69784c8c91e86f376c6e107698c0c607004064c67b7f
z680622e04a9ccfc32fb6083f13b0c13b166397fb096275aa6e860ad24250758e5d2cf5556c9fca
zbc335b7375b2e486893d65b6f309ca0e0c1544a3972cfc37a953965632b74f25017bfb5e4be29b
z3b5a3b2226a55a10c758ed9f0768fbe0b72591db9fb4edcc53c5c4a2a380f54d8054fcbdf2ef32
z5fc35b824dc9a88739599b3100568f406c8814200019453b83f37da2fd305ced349335682b04d5
z4911a52f8e92206fd0e8c3f660dd4685a19deb94f04fc786509793cf02834c034db7c34da2b8e5
z22215863f74df18669de7c190a105fab9c55cebd9ee5aee53d00b5d96764af814a394f2d805af6
z48e11666bf7a3fd33e3ac0b4d151db469fb2f489534883b1abe25a3baca4f1e8a6e9615a4063ca
ze31b9e8bd9422057daa6a521a5b0402bb58a1cb79b423f4c7ad8ddae58ba5a3ed88599e6b9acf4
z585fe46b74fd21ffc6b5bbe8a7dc2d4aa72d4f674a3776edbccf903f81c4a41066f619360c60e6
z8a579bfe84b770b123ea5608f2252a5c87d47a13ff2a608fa8e8f8213a77a1a6a06546c11187ea
z3cce1b4e07f47eb1ef14292452fd8d4df80b01c1cfd1ddac63c0d227d2c6e1835ac4d3ce972afa
ze6b307632b294964ba1ab9267bb86ed374cdf730336a904a02115a92a6586514b51fb9ccbd3f73
z52b59ef81b71c76018a4765b9d623b263a0b5be0f3db6ba9202d3bb6a86c4e6b3d196fca3a886e
z7219b2215e3ef8bc753dd97d6ca02f73a6f97d0e1ac92e022593d5fc028f20b531a731cc1c0117
z5a873243aa9f597e583e0771fb3867aa44d8c26a47ec851180974ab185054f532993bd41016d7d
z77144ff2316811531aac51ef03c362084a2fc80e39576de81b0bdff82ae2c64a5cfaadf9cc03a5
zd478ee1467b14d63ba6c0c3c94972f46eca7dc7f1021a419fb6f2f6edcb215cd17519b5f0d04af
z368e9a4ce3c68608ac87da6f79a38ae71bba27b764fe55507d437dc1c9f7b5bd530505678c8cc4
z85f278bef787d0b253aad806fc0cfe017bc634b373837a2c8f826d3b85892f9b259a71490f6d2f
zf5084ba5bc471a93199c650b5f098ea5bf1f1b56bdea7bc5b6e25d9823051b49751a1a46b81585
zcb5237bf76dbffa315fcfd9b0070b43dafbf5c7f3ef02abc17e0a118d8959a8216f7b3b32c3c36
zf392abe8463caaf8f69adea4e026348ade665746f711ecf079528bbc1f324750adace55b33bdd1
zf467a00bd54d9acf786061897d20a2c3ced76998cdcebf77ea09cae8d7841e638d6364c05354c6
zd8bd9af3f9879074a6bb74c8040408ab57ad7fff97d57f5e7ef5b677bfbc0baafd0f999bd663b1
zae27872616828bdfcb6a4d00ab3197787bc7aa3e0072789e6279b5fcf17695f3df12ab87683f16
z7cf5db86f8712ac764ae58c97e95009979f8d1e1e567d506172abff321699b508ecec5c8445ea7
zc8f082f1cb0451595d23bc2d5df8195d0fdb155cde9d8cfbe58869ef59875922bd5062f7a37152
z4f5cab8a73650af734beba9107a0305ad5d6329bce0db02c500a9afcd5078d6df0f8566fcfeaee
z73ceae7c422c43be8c826e5c5db83ac790aa3bf719982cf2754d8c27d9edea8d849fe12f02c98d
z0c4f090d00f66fe8798e807c4eb46288278e8d5da0d96d512cb3110325bea172af8dbd038a452b
z666b42b2a9a65ea12aa1f473c857261ceb6cd930e815a4fa83e4857c4c61eae04cdcec5fc02e56
za752a10b3bcd37a6e02d3c5337f726c89e51cb2e08425740c394c00c8c1da9820fa47b9596c2b6
z911300522b17f3a556478c384d119cbd907475085a06d7956e1ed36b54aa0f7cda5a47b15ae0f2
zd97319b38425b82c426384ad8751b70268dd69c56010259d25355002c1f73aa4ca4ce5f623b769
z959d11d0d47225108a9d733545b733ca1213443c3b1cd510579c5d3bd84f7cb0942a192ece37a8
zc9234c0acacff223326502fea829b36a952a31eb2bafb01714c8c56dc0668894e00c6da778498c
ze439d30b727663a5e4ce45e431e0d72d598c9eadd7de443dbd216bf40eabcd350774e97eabb803
z8e70501219cd2729258078d1921f26dd4af050b81e3b9f2a8c0e98c12cb9a7359fd1abf53d7882
z781e3ff71fb86c961c61c6d0eea2534622a00ea1fe6abb8881c1116ad799d581c8050b86297702
z09c79bc18579f36b422581bcb1957232d4a3a5cdb153b7e5a0938b6a2cff956271b98159c1354b
z7cfbecbfe31129de267df1f13610b8684c43b5cbd96ab8a990fcdc2e3d02193fdaa8f5b403f283
zadec9812af74bcad470d2d35f90bf78f13e78b99e8a643b78a1f6cdbad81703bcfca1c5c84b506
za74a2db933b5a02cad952026ce91dbdbdafa26dc4df00125ccf0c1d0934764392b93fdb06f22af
za3d9b1d44100c4b87e94b4fac10a8f1b8a85a62a40ab6d4426e3c9f9903592f9333250737bdff7
zcf168175a57543bbda5d1025a9084a3beb061f6d7ce477f90887328e626766ff5bd0546166697f
z2fb484f3953fb2daec44469768d0adb39ec09109151ac517fdf743662c431faac4a0d1182cbcc8
z5ebf70c7f88559727aeccdf344e2835d5b9770f329ebd004cd74c317cbfb7c68a20535b533d064
z2ce62bb7916570715fcfb3c5d851ee9e1bb74d0d9f7fc70af19d6a6bda7951de9ce6ba51f4aeeb
z0f7f594a32e3861d6ee0cd3600fe3a03a08a644a6fe40d852ac3ff3db92479ad1d7863179c9040
z34fdeb07634c40b339217df60b9fb890ef2dbffcfaa552e8b4d10a73712a82b4c38538d4c6b763
z1beddcb3023f1b1e306255c8b9f80867fa70bdf880a98a1f403535735417bdc51f800595099963
z2da97009e0b3378198e2119574c4180e346aff5becafb50d0f4003cce1f09f6a64516c61ce0c16
zf5903f04e65925b6fed07c9e2cd92a09683828170a94fd7faf9f6914d2452b5a6a3ad10fe81249
z23c50ef330f94c634d3fcfb65aab098c2b79822fefdf7a60bdb00e55e64b3fdee29a678313c85f
ze621be8d715192eca65d587be05ee2a4d70325a4e1cf1c9bea42b6631350e745142e069ac4df4b
z66ecc0e41234651d40f881a045ed2eb765a4cf0a361f39ae4491447502e296afc039c5dd7bc29d
z60936d9ecd8d9b638c8447d0355cb49d5a56c5001f8c57d5e60e6f7ea26522488529c088564ab7
z577784025e5a43fc38ef73e71454e93b6e3e5382a86171847e36764d0639192ed0797395df9961
z7eaf9fcab5dc59a682993d46ed573ddf4c1e03a555dc39bb2fa2acc54fb13c41ae534a81cb3f92
z72af05e1a4c9fa82305f1d29ed85476332ac5512f33efd9b6a9ac243a4b8e4d8aba9a15c46b9c1
zc7e404037fffbc958e8dd5d3dc0c02b1d448638ec437f677692ef931da8591b48a06d4ed63c7a3
z9358590f7a40975ad1c7d440773189776e11bd671a362aeb5a401f17bd7a840cf78f64803bd0f7
ze5c937633d6d37f8aa7cd40c127e410d5e5ee17a752094b2562ac88e7002d4aa43ee467411bcf1
z10cfea878a5b1da62f7d6f85156b2b7a76daf69095a94790d17bf2e0db3de1603746ea0cb06807
z2f4c4f59894471aaa4a4bfba3d13125831b6988d502f38ee4accaebe57fecc0f0c292acc30d902
z19afa22fab51f0bc62834a32db525c885abdef3b673d3f18c18e8a7bc12551c95737c5fa9fcfe2
zfe408b162e07031a1f11c243324b1cce20cb27a137498a82e80a14ddf307e2872f3beff0e4b00f
z57ea2d385ec2b8632c3cdc6628324ffff7ebbd1c03166b95b7f6a186511c6f03cfced183406bb9
z1d4b6e8ef15c3c9221ea076ed7d0724eb393a95e2e8015d420e6f1c4d498da4f3af43b62a1ca8e
z6d070c295bcbd623bbaf4b331105897aad70a09fdecef2600cdec857915ccfbe8dc5c9658316d5
zb57ddaacfd508e4ac4d56065a1cd3948db480c3fa48cfb3dac0e11255edab86fd97988b6b34ea7
z4d193ec4c97d06a143fe3fc261b82803b76545187c6e6847f3a9634e86e1724fe450580b80f492
zc588e89ed8587a8985e7ea6543ce50325d7ed4803a7c0d071d41c1dbd1a41fecd94cfcc3a88350
zb1e85990e1643712fd83b7c8160baf858b9ecdb183956decdab14192243f4ad0b36f4eb5bb046b
z9d4921d4c04999b9185e4d28b3cf720be31101afc3b2e1c553d675b1be267d04203f3d080c7fb3
za78eb47822ee162fb9462b12db539e4ea6a9562ce15f956db0be40003ff1e402e88351ecfce0ad
z06d423d73d4bff2ad6743bc3a68e3256d718ec13bf2651d16edbd8a21989b0a8d16795b7f99404
z50ae0f343b112316122f5a6684c670400b49d52b70e04fd58a7eb64d0eb3e1edea2b8c212037fd
z240226f6eab4793d49635afd7fde8f9da30c088ea2233420287d50b1ef5b7449facd355ef5d47a
zc49b9e504a73a051fa55b6eb47ed233e02cdb984cd0462cd15b594ed98a614a164d4e4a2386ffd
zfe5d57324ebfcc55159c90371a60659cb51ddd44a8c20f1cff3fce8058c905d8071fd45179a26a
z49c8ede053346fb68d80511acdcc452707de1510f71190ffb9794b9458c21f3a7d9b300ab93375
zd0b73a7b894b617593ef259bb4b1605c4f1bfafc46ee0857f860d61459401f57c9e12050f3f27f
ze99ac07db85c7491c5d28772ba27715ffd9d9111f14b9d47788df958acbb0446208aa802915990
zac72b2a576f6bf24d85887e0a7f18b6a49bad549e50b450a832485d1c5e5ee39b4004a1a255943
z0688d6bf5ecdef2b6da3e80b1e1c9ffdaf4265e90ca13597bc4913d3573cfb1d5395ef92360339
z34de6b1ef0e65aaafa485f48630b085b18786f899fcbbebe587cf619fe085a3c8c0e9999a8efa0
z4d00737b83f2c9198db103b5d5ad0d9df365b0637aba09cf0fadf8d1b29d457d25e989fa4b8cd4
z1927cd8e7031d59ecce3e34acdf30204564375a5d1c73406a3314441081cbdcf1d5e72c717fedb
zfcd08e39ea290024cd37510fa865d454df47ac8293897c635220ca6f188d5d3c188d64fab54e7d
z5dd5f11c39d3bc58c92f9c001875a963dd627aed9fbe7f089f63a0282bd8336f9db704b3ea0fc1
zf666f0623e7ed56003ae233c79d40e571874dae4a1cec5e296fb97260744813cb24652e9058f28
z43256281fd861c9f6394d347e6de5195f60450001a5b85146fc9e44fda8e51b3a82c7e6503f6bd
ze9a782834b18eeace6caee77efaa337b9a2517fc1b3bc9e9602b1ce2904897bd7a20f2d418c96b
z2ff74aec86d1057a5ac75aa484ae141a6f64febd466944c0857ed51eaf368c8eb222883cd4c8d1
zebd0cfb39b8bc521306b1b06d9eb426ce75c0476b04af46145d739f176f713335e11fc5eec9f97
z1c8670f7e18d45411f963431af0835293bede9cdc930e23fc568ea31cfec4bd308eda43974d50e
zfc58512d7cfa71385c7fbc59a00d8043233a1a504ff0d67a7e2c79b3364b001f5e907aa1271584
z91ec6bf43f621da5b54b38847e10cee4b184bed381e8861de38d5cbbfb9f26b03e78fc0f6d713c
z434251c918e10b942eae48ce8458c894af4b15668f3c844d8090fafce814983d0d555f30d0154c
z861e8b9e533168c534205eb80935f91e82eaa3989de4cb7eb0567ad9550bfaf4ac0d531fb6f1ea
zfbe5d7e33ed5d1c2df254ebf641e73de8e9c812262d4dc23e07d1705b94ec1ab445436ac798bc3
zc0303e5b2f65d66854d6adc1ed57fa0afdcfbdfc5cb9584e02856e1dcc065fc37294addbb77135
zfec9743cbe4d6235cff9538069c066405692775ab1a1a53ab13d55df6bb38282ba4109ca54a75a
z3cc562d004a96296d2baaa549774dacbf6c3f85c0e9df0f42d486af94310d52b301e698fd8f422
z9cb71bc86029936ce3c8d66d3f8b46644b695b9d68e651a202a97caf0786011e99f229996315c9
zd8fcb4c4260400a9efab03621164ed67a4f25acf3a80bb3f7b74a6d2805b77afcc48eb7be681fe
z0ec7913ab710509b083824898888d9668c9a73ac0346a3bdd211313d55da65a513aba67390a379
zbe3ceac8ccb3dcdb24928e72b5ef0fcfdfc0de1b14ee412a3147b5096efb3de87d00f5321ddca3
z1ba6ef6d382bcde4bfcdbbd7315804d7e4c8cf0e35aac60e66fd062395a6840570fecc960f9f14
zf4876a8a20f5a08b33a91e68b43fd579aaa514f50bb94a41dd23f49f3d738d15579885c1e69829
zad19a11010a1e9fc9ae2b06c7ac7ebb6a4d1123472854bb3c0b49a6586a439a71d55dd19ec4ee9
z3b0ed034b0d53b4d675c80985cd1e02b4e88312a775382cea7508d60b5765884f81ee79af8b253
za8b6ad9c86e8a8154ae35a88bf7dc0db00606e7cb61ab8c1a60488476385c7852d5ee98905ff49
z14aadb43ff2f73305579bf2b9d88f97cc4f3b13c88f3152bf65e1f5d34a2fe6fb82b8a6b32e5c1
z2e35969726269eab883bb276b5ba5e26e16cbe23743bd6603f5e1ae42ed5c0b3868db44dc62910
zfd00a8e75e8f6dc007764dd32285058f0e6b4c9d96561d96902f5e3c19ddbf14bb7023ccba56f8
z1b7f04a4e94e11a5276ee62b45e00bb9fce9298525b6bbe5b2fa23019aca2076555f93fa7cdc87
ze98ed345d0754476e860a3625138ed095a55633390d722c128c463a1f92040c6f0ed192c03f42f
zf7594c5749429d8f4b051b301ceb1cbfe2ddc7f789478da214b6434f90e9c5668e43ebb766ea51
z04d6ace22f96e3fe9c896ea147dc108c5d03d161463be325599a6fb0dac8912b5af48e2248a4b8
z5bee6d6debae58462ae2740977522d880f5ff37d20f1f2800d6e2a7a0072795a23ad09f9fbed08
za00da709969eab874ae238333bd5992937897afbc18cfdec8ad818a7a0e9be111b16719e3f3041
zc24e54506b72ccf1d9264a8badb2c201b878c723ed91a3644a59f8fb3111ed1dea320152a0b804
z5f904be39ec43bfabb1b34f4013ec51fe8e63cd2ce2644bc4df6ff4d26ef75324321f0abdafca7
zb52fddd3d9f174c2a11194e97b277d6a4b5b27173a2d34c33e79c72af4c1f1d291401088dd6fdb
z3c535a81bec1e37b0a11e809514fe7d22b646372d736a64577a845172226587c7206cd7cadbc8f
zc34a21ae4b856d57082df128199dbdbbfb6b338ada2006006e35fc6c7cc4b8485baa677b39733f
zb641f127bcf31c5d7ab7a7a6cdd19b2200ef7c1a708e1e271ed88658db34ef542110ef961da4b1
z7e05da68cd5c3550ad26088cfd89e84e76cc458e42a92a03806fb0676069c15ec2be413fabd47c
z47b627581edfd972ef0ec6f10a93d62fe8977869ca2063269619a32efddadcda07bdde53a1c1c2
z2ee37c94e500fbc9469b704e14978b1b2db84deac57b97af5513dcec85d9d1b0ff9f7a294809f0
zc6b34a68b09d130a0fd99f34d7ed7a4635f71e57b93e983a0cb937c104da70c1ea9b8599a9c2da
z47dfa96bc97f537689cf23a1f0c602b473a87761a910267eec5eb93f214d7711e43df00970acda
z07f863b2d6b08c23274abdb384c97c9dbe6de14f2ab9577e7b90e1fdef885e97c5dedc12c205bf
z98a264b445fdef6e93a69dc646949435d92b4927649655ee7f552370ec1dc818a8c9a6866ffea3
z0287cd51d6c0432ee0f72f44d6198d176914d56e0888b96a0db1beec20f137c004e42c422d9c09
za61cd50339feb6f176d121faf953896af860c8ec9c5507c726a945427af3c73d3851c3f1152425
zd509ea5438a0f9200e98f54a80f5001cadefd0609879efa2dc8b48238aa8e1c1c921cf56b2b3e5
zf904c15e53e56e5fd207850e10bc89e88951455544bfd8d4e79492a5ad4a17cf39f048b2bf0813
z0cbc026e6b2895598608b27e4c151aad15487e62e2f6f2a2206894292c0ee856d48a80993870b6
zf9acfdea73295f8aa68938ca368f805e97f16ee4e49e9ce3294219ca9de5172720179933f28e93
zc0e3ae5b43a7c9f75490800959ddb15eb3c42193a13a9af09419854af3634b0cba01554e55eae0
z39d3625f3a5b5e0345f0ec4a8e5dc728b54af81f59e8df56739a15a695b08e83a44eefab96fabc
zc2d0e472822020bc1bb81351867faab3a6d272b4be31472f59f30221f03173ece0cef19c8ac04d
z1c8cccd71ec74d8565807c03dc9de230c6463f6318097a169bde09b5fcb2cb94b9b39ba6bbdd06
z031ab13c855d08b4e9aea55b48bf16a0777835b5fda32f52438a7aa570b8a3d989b0cfc1201def
z29cabc4d6830429c682aa3e524f7f50e933ef1a4b19462ba37077da26187290338ecf188638b39
z87085c6dbc4356806fa11e2486c7b1d41d48d02cbcf2cc52222794b2378cc4ad439d550ea39f33
z6a5bc3249e5da2a1bd177f150a141ada82dfaf6b943dc824da42414abb839ccdcd53ff94cc33dd
z88774f18b4b6190635ebf0392963837b30e135998590847ef053e670f87a5b165eb57319f560a0
z61c5121fc5972734746a7f74288ae927088818a48da22c2888b770cb1eaa0450bd414ddbb045e5
zafa65691d9b0f8e5b6c221d552b4e00c0b771b14aae66c120491f9a2acb51b3c17f7d3a17c3f0f
z740103249b716f2ad905e416bec197b68484ac9a86b037aa2325c531f43257d1c7c28345bcef08
z7218b095a1c85d24f366ecf22f5420b3c14f87a76dc14dec7e63c2a1047b3f05529239a2258361
zd9923ca5fa0954b2a2a73d81a1969cb1507205273d9c1737b2b2ffb2315a769d004620c9b6bf7b
zb700b0b7ac39c4a37d8863707e6d06a802d35fb125e5c1764fbd79f0254d8c7f0af9e6ab06ed1c
z3c69431fbd92a3145075be9a429c4c79847339193a6b0e2383579901a1eb2068a1d4067893d388
za8d61f0a4b36aca34edc855f2aae40a0f5e2c358c47573a5b617b483329d92d6bedda2f94539f7
z9a39d0da170914d6b1e294d15b3c748612a470669521eed4f98a078fcdfefac80a1cbeb2c5f54d
z50bda0ff62ecf025754f6cf690e76700c77285b5ca56bf2ad4550f59ed57b6cde869489ee68520
zca0b34669699c98b1c8d8f66411f382df68a50f6f2a6f05e37639b81ae1c8b8e7bb2811953d352
z08e92d7b65749d0cf64314062d35f342b4f36848a64b3916a3309a72848ddb4aceae792b519771
z05a7ebbff3f0ea753b4c6ba3f030d6c3fcdee2c3cb59d10db659d592ec65bbc459fe14d2851755
zb1958511fb6983ede27511e11f0ae0cb3d816ffe39f97ec2213cf963f604167766b00782d4bcb0
zc75fbd557b74e6458de576f2c6eb3a705e18f69816189e97c357b0c1451fd6608dfe275e66a2d9
z80a8e14998e05d6097f8c50cbc81a495b46d4c65601414689c7532852f43ac56af07bfae4b1c11
zfc215c001d049b39bfa798d6b69371a956729747872fb5d666353f5c6fb786a9ad2a03cbfc1aa9
za3d130b92b83d56e266c1380c602ac7d6a2683681fafc45f64a1834ef50e9cf9cb3b734a3ab84b
za54e3e7df1694d0151d6824916c9fcc33ee80d7af6fca2d38d62e7bb8cd49b5ccb9c5f25789466
z524e3069ed07b3982e2e13a1c6419ef9b0ed91527224e270345b836f532533f100a5265167f5b0
z96e58a58c8b799749d7c24ce137d1d2cb541b268c7449c06cb1e69e4d33c22fd5520bb9c54b790
z540bff924b59526ee46cbe5690c2fe0ca31f0999a92f901bb76e958463241aee202c920f0bc84f
z4bc735cdbeb8b5fc17e6c5cdef4c13dd459977663f75a28c6e9e461806dd9f6689538244456147
z5b8c0d8c21a5eb7624b67676f6a84989f409887d7a5cc2ffb154ad4a6e97c74ec32de0e219fbe0
zded6fa47dfd0e9178270859d6de13f2830391ece717d3ff231e0667d24eb399432e0de6d8fc194
z4239eee9824234f4cc9b8babc4f3f389ed654f65d00c5c828ec91eb8bcce4b6bb5e2b493debe85
z202509da10dd9d29b2352d3e3cf39d5543ff33418e8a91f406c8acd7e9671d5b0158e9b0a6cc17
z66d2321080d334377bf6dec666229f506df6e26ddf2c00893f1a00741a2cb14765319235f87071
zd48631a73a00794f5310e73cc641e1c5c98736a24f4257b1aeb4aa572a790b33320cd60483f888
z816c3624651586fdb1e4a28da164af03f43a4f46f42f6c3e4e97a23099199f9a07d1e151b09c40
za1688fedc4cf1d409e48135904ee7bf1caa8f67836d1ad4259df5cbfa72a31bb8ea6e606fab900
z066c0df568ecb4410bc0e00cf912b0eab131b87deee900f1bf67bdfadcebf67d850260bfde61d7
z24b97ec95b416f3c494a992f20437de9119a98e327f6d9f4c614068cf0cf5903cd9d2e6173d685
z009804ffec2c1317204590d8f4bf017dcfd8367acbeae2338b15bd6a18388cfe39f8940111f5fd
zbdf5b198916e21fda1fa627f19c8f37c0e13aa2a3deb77ab4a0426a3a4b2b69244cb91cdc7833d
z55aac9e0e564435f1e7de44b91949fd85a213f9b9ee5a7133fc80b0a3eccabe8ab63ae7b1728ed
z9ae6a309ab7ca85bc7bb3c98feeda44690f924c61da6ac92478964f4c857acc8850358f130d28a
z7e655076cf8c3f30d0c2200a3e89972544dfff384fee85e34b08fadca9e65eb6b443440dde20a9
zed26ad7acc1cd0f3205ea4df0fb2bdc6ca37ba8c9b127672cf3f2d90076c0503161530441d78a8
z2252ace2c093541088bc3d1c1a89245dfd653252be76e0b44faaedba01099a3f49f9101b8f8e76
z7b3a45ac961e80f3d9794980638a99e1317daac56902113ec20fb7b496a41696221b9959a30499
z84f05e419e07c4a95d2c78e212f7abc38774a1daf73d9bf7bad07304f5ed9c1013ccb6c1d64926
zd18e7771a82878755773e40958b97fcfd8229e3a3b688044fbb89782dc3b0007571b7481071129
z437aa05536a1f907f909aa7ce0812554e5e00148be2050edb305f7a56a4ad0360852ec7be511b7
zd2a6d6ca937a8bcaab7f7475a0f8ac6bc3426f82a36fa15c41e55ec890b5e0424d7d6c89235e1c
z060a7e4d9a1bc9f9bd24800caa2e5239c65f828c91af32e058b06c7805d4b7c036c7ad6ce087c1
zd26d88198300a4560b9ff43ca01a4266da193ebcbe478b41a3b4cce52230d05b55ad991187879a
zdd60792213c6f61edf57fea17a7d47107fe3d5aaa43fcf2d886db270426b2175910ee5a9981148
zcb2e0b5619851a255385f25698007e58651dc35b40dc4901fae180653060fcc6d6d5f20630bde2
z6782edbd419f31cddfa0fb1c5df9ff209f06d2a4b38f766db6760bfcd212a34dd034c4afd929dd
zcfd034256d2f50e7a0465488e572f573994163b0bbc68157a1fd7b2e0ed24e9a81b2341676b362
z7db51e10ff4da95e8332cc2b2d796a11d05b9af1ba343d2a5344381da818c695f4b21baec552fb
zaa1e3aaa3f7822c164124e3503c2561bcc1bd96a02acc985da655f5afde01fb3ab93d854ba0c32
zf4e67514e64285f57005c369808dbe1cbce845df68140697ef62d340b37ae3fa8d99e281794621
z2205cd6c43dcc34bcc133cfc1c01b155d25c3432cbb7a448f8b25bf1da3c3a18f6956c647e40e0
ze26cb7395f5e38813b1c9181d8a037cd67ac0dc309e633ce616021eb3420f82c557469516eaee0
z1694548f256d521016ddb3d3008e35d78b1b8ffc8543a32083fa100266126833b55e6cbb514286
zcea78cd2f0438c00489541f5f13c0572cbeb7ea80937b209b4fdf8314d92e1e261c6aca58d0868
z587c71122e7bbb0a6c9ce8d8b0cf08b94036c759b001df6df88add39c75853faade4331fd60004
z183a8cfab07bff50f7c916b1774e62295268c243878e32046c78e85f4c972331e5e1e490a91ee1
z361a7a547e964e00f6057f65f62ed5d6c232433b64317e0ddf07b6059c98653fba733fbc62b0f4
z677810138888fd5a4821eac395d9c382fe84bb36a4414f4fce939ae4bf570f68bcaddbf678cabc
z739474ceb99fcb9746c561e0e0e539f73c9736d75995915502e48a01697b8c86fea511db9fba75
za798c5fd1ccccea4b7582f6d14de5c34a12732b259b9bded239eb79d0d0a9c9a875135540a41f8
zc00f995783b42153967a80369cd36538817ccb3d1085a139eaffe63f2a1101b044d4e3deb370b2
z0dac9a387f8a5fc751b14d8c8c88b52803af31df448bb3cfd3d9b5bb89160a08ac2187deedac1e
z8e9d7db124dd0f1f4752dc8d2ed8038c7f35507f8fdf76b660e07ec490b1236381c3954f8134e1
z14636528bb7210dca9e971f3734ae09ec51603d5bb63b53140e7be9f33849cb709827a3ac071d8
z7f90e4a38c2c0b83a86c73cb2dc7d5473d5b49a60dd2cbce254f02d3548fb8c109f1b273a3abed
z9cb676681aa66c1eb97c5cc6bcc1772879ad6256b41a69018ffa532d5a38c48cbe659d8354e6f0
zbe9bfbd1aaa177dcad158b4711eb9af5983bf97e17dcad1f195491205e8dd10a06f7d1519b43b6
z69f463262fe4142c3579cdd187b6f0167dcd56e1a1d5f1328432a73b5b9929fa1a308242b54fd6
z37a5be3bd50cadfb0c3ea03b78fa2995175deb62e1de8f1ea5ceecdda1019317e093f2a1462e9f
ze1be6267d3771f1b35ee89cea139cf1a6f5639f1d5f530053bc5a794a01efd5b133c544a7aa677
zfb4dd30f9f7b463a667fad2ff3666dc4429ed63c52edcf58b02c113f829ca2e7b9a5041e4fee3c
zf5f2731b37ece7fa96499a15353175317903822b40bbccf9d7d511ddffc7e781c2ca9c0ccbe06b
z5e682b14e907a0ff898c6c29988e8855ce5b3a0315d0ce357f77e536f4540c7916520af8a301c7
zbc57b48374493faf98f8dc2ba02d41dc83778099e3afd4e90792305c4e6da99d2c909aeccbb54c
z3dcdbe3147720e054f6119ae6cba6ec73e437ea82bae73acaa8e8bb1f52e79c444e13c9645820a
z6b94eb36a557a5e7541cfba435db549a61414703095751ea6ac1312b39697f4552c6a43e5b3878
zd5767d7ca3b38fd28288d7b56affd4b40cdd5b2f944e70be9f744b0fadf02e7a61a748a140a34b
z7d1ca1755d02b5be57b2c2356fbf19ff5515b5df71d6cde45cb2a4581a3310c216fa041c267e9b
z6afd5f459282980b6b556a74383b5fdbc75353f43b24d90632dfc49a235ac72424f09775d9182e
zfe8436e4b52d15f4eacc38f754f6d758f5aa0a22dba075bcbf9f6ea60c7762523dde42b28965b5
zca61d19625545f9e37b55324da47bb5045701a55cc6661f4c78510da4d1516004db099cfd97f7c
z05cfa3b2a6379998c04e7ddb21a537d3e9d460a4a82c13a505b155bfd369bb8e3769607fb1babb
z0139dc249ff4155c07374a13ef9e92224f80eaf321bb75787ffb4c587bbcc20f0d66af77e5bf21
z81f96bc5a864cf4f97273d4164b76cceb2be1b5f8d6f906b25ca5880eb4aad516246fb34fdb26b
z3e2031db0fcbce7b2d5fce3874ec2b3db5a306f0bb54f85e42479d9f6f6d8e1f50bd11f647d81c
z642e0b58290a3e1dd840bfc92392d8994211ea0630ece0ba01618995ffcac85ae04210f6de4799
zd215c0ef55f730017d5274849868f5fa4f66518f237d262d1470ab4b9a4840c4f3b5e143e1fa63
zbe9345afbacc85c74da8e583d5b026489125b03888865ae8c2e76ab7d918263860ea7a814605eb
z3d8d3b5556736d6ddba8018e160e0ecc1edea7dafb8092bfb26b6ceeb44cc9f1c226462c3a2e85
zbf1c24d4ad88f7790d047206e46998340661de3fd389af8278ad77e743cbeb0c493f7580548180
zda06ebd923f32f21434815bc09b3ed82819c25444a435b7c7c6a59a71a6866aa55220c8cf3b8e9
z61b9b629a97bbb2b4f8719dd583b8d9576544b9b4f27e51d7556d229b6ff9b43d4c2d9c718f1cd
za496ca3e1bcb695b738a5af16a52efeadb97a04aa44c5597a160ac13f958d941ac74bef81723da
z6852ee8c0e69a48958d52b36891b86a31aef5316923fa499ffb050ab15273803db72d9f54c319e
za8da83f3271d8f4e44a1ef24b126901f53814165cf4df495913151f8e07a7ec8ac5aaff7f0f9b5
z754706b5181f8e4ab462c2a9c30e19316715583912795b6a94824c894805a93286b3b84f26d702
z16ee85422761a9753ddb6109c2cd7e05f0aa0ee8afdbc9c30f9c7705cf623f4a9897a0e8a4436f
z85a0633206d47c4ec29fdd73a2658ae6d09399f3052a1f93cb444b9805a71865823fd0153cced3
z3a105b1a10a8bd9c9eb210ccc54b480066806980db20b14a303bbf18413d7158f37b4bf4cd4043
ze39c207b6e14b72acdc4bceebe7077eca394ac62a0385b0fba9794ffa512a58753e84b382a6444
zc98874f1ee933218805919a0273a62b4e027e3c0c1c72b2bc8c638fd70489b0bc16463fe7b3aba
z279f9cd520f2921a081de9c1fb40438fb08eb7588402f908a041e689c9365e924e179cfe98973a
zb7a2c787b72df29dcd87f595af13b414347eb9c3a373700039e985e350a530b2641843c1ca3352
z58164e77cfc475cf198e95a6b984bd3250184c51ffb888c80432f97f55c12b787d1715c262c9d5
z7793a7c77d91d4c8aa53321b70b4d33c8c62001af80cd9164b3de10eb684d4a9f876d5ed0d9e5c
z1e0613c2336fbb3ee40ad7a3458b6760c3b9b173e62a6f75501966b99ee3657b84cad1494347d8
z1993ebe09aa1d42688cb56cd0094955e8b8ebedbe27642cc2fb7793a5bc128d79f7c439913a744
zbd629bde3ac2da63718c2ba1970f2f540f489dcfe1daaf98d1fdb5ac66005c24bf786ca7ad8c4d
z8b190a2124911ab17972fc87471596b3239407f7e79b240672c8dd1b3dab399cf815a13c98e228
z770159bd9132beede03f5bde880c788e573126adc0fce720a569dd4104845ed9bb3aa5157c5571
zfd9a62e39c53b660dce28d97926ba895ce14dbf480cf138dcd82ba66d388a7667b7fe7d5a0559b
z5977b6ff30e36165546920e1c8473a78b8fc508ec1aeda0ad4ec4f892c5a2a1f0427f04d122aae
z618e6182a36d0d78d9f129c9b1c4dbbecd9740b3ea7933bb2fe21f57a0bfbd91710cb24d56d9cc
z66b6514c43a230417fe131da717f1a5c8455e39b5e4449e785d4d2e459788a05684efbae0aeeea
z263a031b2bfdc16d2b93f5be6457f7f21cadc7142043ba260bc895d9420d17dfdec101988b3fb8
z068784639e56f81ff6dac3e15ef0757f99799e3a848818960c2c6f9e6270e5e715e92a70b6e788
z2085ac9a46e24e20a150a548a17b8d974551be68652e074c2a5f6dfe393ed28450e26b53e06094
z12665017e6d23a04d184fa63f3a04a96316e6856d80f225b6145b588819480b8ecce318c70565d
z7be73a8ce57a6fa2d695b0268f8896ad7e9262a69573cdefb5fef945fcec8a3d1367a8a25fadfb
zc6f91ebe05e5b5af11c252abcf22c6ba63281c2b1180a72abe4eaf60e460a2ba5558d2b9e1b0ae
z92bf4b9c8c5f5f9b6ac277565b1d114362ed83636bf34e49fd322674ee717b78e2da04701f4bc6
ze6f07fb477eed5a7737265b604528e2c60b7c381a3a2f8688a00aa3d7e0b23d308b16857a3880e
z74c4ab65576149891a6977517ea924a7d99e5df1fb5d1831e551f8dcb3778b9ca3a76db128ba13
zc86e9192c02a5d8392c61c6b209b07f4b08b4cea0feed4fe6c5799923bf87b7217277b52a20ee5
z3167119a2a6f131893cacd2081902cfeb114fd22b9a5db7587c33ab5ac90a455d3f828f754018c
zf359c00108e5e44cba037101d6f95662311c6bb2a0fd1ece5b8c59136d09ef6f493b8d703afd2d
z0f91a23477f8006d2c91313b48940e5a4768aed7509d8389740c6a65e71f4305bb487d3dd8c1b5
zcf55c21987116ae322f2f1ed228fad68baaf01ff4cf9946af5394dbad2c9ee37402f2f7490e6de
z6444e56d65cb47b425c5ada99ce4f43b03a85867291f471ae8a1871ddc5645f89fd2fff8cd8112
zbd4487931673fe9dced7955fefdff8b5998c993fe2b18c042e82a2cf33f7c8b4047b305c94d431
z2a76dd9a08c4fd8cf5fc48b4be6dd92e883b95e2050ad1942d305eeefc7e020d0c7c21b46cf476
zb2aef72eeca9f4f56c3fc9fe2d27f275bd7750cade24762e7d8f84891067fd86037fed3df3a2d7
z46eeeafedcb6adc79a02fa3150d8be35b9534d9ed9205ff5cf9db39c8803842a1a86d402db54cc
z4d46b5f6395878caf3378243354ed6992bb9a9d0e327e16d88b3f6e1edd5b79886dfa1294c7c3b
zf82bb0bab735bd8ecd603f067e81913f6cad5ea332ddf57d101827fca1c2cb02782839f4530262
ze85269a07648da003bce954b3e19fa35cfb7aa156e6384413059e027f4acb266f1d1b4887c26cf
z338cc55b2c29490a04feb4fa81237474b5e7911111dbaae4e306d8489a7ccf9d586ee0358d61aa
zd59ba13d422259b3f771f9c7046277af89df8de783ee87e33360b3e8e10338c13d13566dcbede5
z0b0a9e3b3c5691068f9176ffc5b6f7551ebe63d34f62f21d4902fb3ddd01d83257430e7811585f
zebd82e42801f47f35f8952ce719ebf7e3f821e97ac5606d3f0da09bb5dcd34c73bda969287f78b
z64c82fbd553a103f8cff4a4e231c0411e3d3592f17f807a426b6de646c78f9966ac3ab9c6d99bf
ze8f25b1d6f31e91daf9008184d51a7f6c3dc41570df21e9f6132d0f761cd6c0a31cba13e684567
z3191b1e28f7b66535ed6932189c1ef126cf22efeff44bce3343a99b7ed763fcb8a8635f1c14519
zae272c2fd539aeba043d193cdf0626a5eb492b752b0702917ae7e4a93574672c2aa81a4b38edda
z7880e0f5bfb708ef35a4d3c8cccdd24b3aa7ffd9771a813be3b147de9a8781e429ca54db2fcf5f
z17ffa676f2fae85afa4c857ff42b85dca1caea723775a5ae8fdcd90cc235d88da19d97e712ca0b
z7bd133a0434369b1e3d1db58eed02b7b5d33e4bfe1b74ec35cbe0e6f55bde74f93b19d7c43fe0c
z36213794aad4e06b8576e529a37bb989c9db5797800245072012197ebfb32b260da1fd14b78e59
z19b36ec52c5305081815cafe0bd2a766773e3c809a02b3671085a5efa94eddc4664a1810e8d556
z725c0688b271a4ed69b6a5b9a60e16ebadaa1694d63d169689affdeef6dac2e4b19a913a9afd57
z9806eb0f2eee09a0516db77bf071346426f53e4be6df921f78a5a8c2ebdabe6a21a0c07c280596
z6b3eabe4c4694b5f0a5d6b408e9e992528c0372157bd7c80dca5213cba72506faa35a9dc3f1ae8
z3bb4d141f6246508796ebb58df81824f17fc5a5e6ef816b9801ddbe4283253fab82056186d00ba
zfdc72b5fd7bb5ccbca4f8725e6f4198dc4850707825d7551af681715f312695ea341d4a3322aa2
z7002941c7e1d016fdb6b723fc6cc9da6846a5b9362133713aa598c9ed1fd9cf85e9a6bd9bf3123
z17064cb79df123b21339b01a02e0255eb21454da5d00c5eb61849c711601c6820e3ad7120d3155
zef20a3c998c1d50439b2e0a78cd7f1704428b9f75736c0c727584ccbcb780bb3f9ac01ce4ed8d2
zf83d3e3700ae034ae372e7a81f02892badbdb5660f8a1c8709321c90384471c99f24d5ac281efa
zb4b359009ca1c1a8e293bc00bdfdec224c7a3aedcea3eb379d4a9d9c393707a6e759d2395cf36a
zc3ff2c9877cc285ed3574514e18bf64f3a8a1aa4755c5681758d16a40e31ccf243bd7f87a78003
z7dd347bba0abedea0c2bb6bd7a2bdd389b704854ee57817fa09ccc909b28607a5ad6e8fd13b87d
zaa8d031711903bfaeab267c2e436b89abf4de0e1e85e61300612d7d9650164159ba342d6e5b06c
z09162ced0799c10d37fd2a029784bd2e744c0751960e7c64293168a17abbd20c5f8a0b5bab9e37
z585a65077d0d08f8069bdacb7dfa8abbdf1f77e34e7e434776323adb45a7cfd07b51a4767ef9d3
z4da34d2aee2be1d92fe3b3a69deab6c06ba568acce97ad399404165158cb7758de710c2d1e5626
z04ae28a74e5f61083fb6aa3172b8d8d37a840940c4d39d6a46f6761efb263d2e9630747b30f536
z8f251f5bc487bc34655e0ba3fc75c38beabfb9baa9865428176ceb80737fbcbce8aa8f0f77fd45
z5b48144cdd00fddc48da26a22225fa96968ac21394fe9d5dd8c17e1ad9b05bd609a4f5fec92d29
z8d3565bf6dcb4581a268c705e9ebf881ed54e94d60825efb1c0fa75b46a82c45f59a286e1b8cfc
z7f8c53a00e1f6afa97091faa3153f33198ce5be0beae1cfa65e06b296f38a8c4254dff1c5f53c3
z6ab8d955d49c529d521ddf5c6249d4568939e0d3807da9dc977b4b50baccf85ce159d09ddc6dc1
zfc53bf615cbdff32daf09a193d64c9b83dfaf9e833b7a7351f13c1afe2c8a0fe2be64397526008
z17766cec1435d561a47b211c18bf308368eef668143bcf59868eb7be38353c3c8f19baa732b38a
zf79bfd01f13b05e10d14e836de880fd3cc323e8a4ab9e95cdd3cb4deffb3c21492fd6f6d14bac0
z1fea38cf52011aa6ab7bb9a66035a7e678be459977969b28f0f2a94c88bfe8e9d9f25d17b13b8b
z6defb3ed7c989fb9d573612b26a67ee9886e8b2e6a46db994e5761bf25f47763dad3b120950d48
zc5f47a80f7fff6a60be7f038fffc1680295de911dac4bd4b18eccd653ad1a8b2fa6e433ab66ae7
zc8a45f2d071d2dfef62c673e46abf9cd74bd179d2ecc598bfbbeb1378a2ed3a375287f21153d51
z4890fca0b3bb780972cbe2e093de92cb5b75368e0811368c2a934f650bc0340057d0179f912a5c
zfacf5522cc21f6a7a368b4479da79e38f43d7392311ed66681ff6a03dcd83a343fdf7816403090
z6c40ba9d4fd9534206ca220add71c7b74db5403c0c6db2951593b75d4cfd595b8bddbaf04fa2d3
z29ec542272e2e59017c899f260f858ba417b2c5c5389e7fc35d90458fee1ec109c0303f246290c
zfce1080e1f5400dfee9e115e0b4c67eb13efea0dc95f78747c6472d68489d14a0a234459782db4
zb586e417119e09230cdcee1e6c590db1b193b4a5aa7a996c16cf59c30a761f04b29cf46d74874c
zb389fc08b0e9bade2d329efee2f40534651a5533d09cd1d4d4150bcbe56072e81cae716eeafafe
z068833ca8c23e0fa6038be7d3d3005d6ef0f02b6dddc669d9aae195f3d2e249217d5fb7b3dd57c
zda50014ac7c14cce606e941a31d47ba12518d4547554a2050c0914cab71399b35b5921aee83e01
zf0de101a7dfedb55e3ebb90f732610f38daf492d0acebe72e6c64200ca1dc93c869c850d404ae7
zcc9a377d41b9eb7e0e0f614b9c13584880ac0a85303f25e4fcb4e4fddc770b8620c60297084495
z23d1ce8a69ed442fc914a168d34cde31d825cf0b15c75be4484811265f968ae48b6353ab10d707
za0c851f57ae6a11013a2dea150d9900d308217d79da3af93c0639ff64eabdeb1a7bcafc5ac7455
zd0687513980453f70181749913ee3e3800e004a9648dc6f971d4b3842baef9e442935eaaf5c330
z5679d28353f6b3d92c043b3ed62b2c5d1f0c6a516d39e752eb97f001365ac1fcbedc67f32aa92c
z0c6be39dcce3707682380748de0d5e12a5cd1a5068272bfa4962df2df0c2819b80b766783474bd
z1f7358f903cf2a561de22303223f8a7071aba3f9f74e7038ed775d549ea40b4291f82055cfe45d
z576aa6edc17116baf1126d48fcca49766377a52f1ccec094270460a538a19c19896f520c7bbdca
z7b281eba9f5bcb436a7fdd09a87a74ec59b591ec117e908a2a2a5aad486cf6a1715f534c3cb1e4
z7ebf42c15445fd56fff7eec065682fef50b640af9e8a7e2c7de4f61806eda282d0aac3fbc850a4
z1e49b4dea4e8ae3d83ab8eb7329c24750bf3066a91aedb5d3217df9adff46abbaa41a9668ae1fc
z9a9768ea676d72791bf7d87b3556a8b079033078daee814f2a102ec02846b7913e6cd60ef517ec
z7c1abd4933179ee63dde5cef18b105d88f0948da7b9a2a3ce2ff2abd11db2c519078a7097281e3
z759f0ab423f6a3d35e7905b20aac14713ebb298bcf89135a5cb1675410c25a16edc6b6ca72d7ab
za22e7aabf78cf0893c4a50aacd040e5fa9339b3842e5073951c0987893ff4ed451b381e9c09f26
z9c1b8282a74d9447b46cf1bedf6dc98ca3a44dd4bd804de2fa0ce2642c16ea3ef1890f908645ba
z857eac3d21735adb280bc080e00ee78e4ee0dc231e9bd1604d22bce97cab8a4f40d476691d6da5
z65b70f6b0a7bd02a5bb76300024930d02c5ed9db6a6674b66d17d0bb5d7f4cf89d3f81f2e2240d
z2f355a9df70cda954d3238a522e3d8caa4bf57a2f4f3583efc9c9f4e4d533e2c0f244dc825dd26
zd5b6db8d0ab28e62e13ffe41b500567125b90f63e3f6666c30585ed9a88a0079cf22a8c9fc5302
zeda2fff07285190418459d889e0d954282e46b4d57fddf90e260e7d9daa7e0b66e9b3af70e0173
z8fcf38728f958b1b5191312999755dd840bcba2ddff0911e9dadf0dbd4c3adeb5d7bac84ca45a7
z6c6d5469d83574b567e1d13f91514c545ae8a94f5146f8373bdcdf267d3d23581d5124b72b0b5d
z869c556b27ce123229c93745462a61f3f787a102b8d3b827dcf1681709182f71682d8fdeddfde1
z1217925e029eef460b4a8808178e2d256deef4630c265c67adf7d0fb280fedfbcfcf6f598dbf40
z221b1f57ecf7ed5170accffb1fd44a6b2ca64369a9d355460d3769dfd811abc5cdb407d69aa8ad
z449e217dd1b833f56ed4bb0fc9305f6418e73c66fb5187229247d898fc2f4b87fad164323e735e
z77e2d93d276d1bd9a577e715a2ae513b29e8b14fc738544371fd43b25e77e571b4741d91548487
zc7f16daa55cd16202643fbff16b8143a6102d01aec5bc6813cbf611ff80895c4e7ee852de5263a
z625e0988b142d20187201464c076e6b65d70b16fd5efb198315ff71b99f286767f68a0283e3699
zf0266bd16b5e5dc559380f194691397977f35c05293ee97a5d1e080b5ad06ddd425306c621b87b
z9e8597f6577dffc627248c470f03aa68b3551f896b9b503a3f06f27eba19546ad3bdb57b8f81bd
ze97b0d9622f8a8c74a9e309f8753b1192228e74266c9e4573192a1c6587d259babfc773c4c488a
z03e1356e2adde8158b36f62553cca796bc5c3d3bb123ba563b3ddb080de0e1d643d8c32a72ff4e
zf9345edf4d314478735239e6dc2e6e454889669b11e6b7ace866997521dc442d9f0b0937a04cb2
z17054daa745ed10897b04b93e5c21af4b45689a3f455321a91f03124ef4dc3ea1a3c1ddeca1fa4
z81d02df308917639f21515f4b9b0ce1483aa6a58eaadded82c8bdf27dc3386340b86265d2b6333
z65792b15e8eed5b572bccd45999ec63747e73c2a851bd211a3c244213248bc74827d05b0e27578
z90dd49f5f978a3b6ade7495580200d93d056c88a7862340e937486a401cf8dc67a41bef20d2c8a
z1b352765660d44799720099a4237c53aee282935c3eb4593e48d0966a99ba26e6fb9f964c1a2b4
z4a70b15b6a26759ce8aa6cf6fac3518480bba448d163e17eca5b85e7a66f232152aa48043a688e
z6d75cc76835682bc4f3d9600af6a518fe5191a4e0bbff17bbcac95b6470916c8d14608b029e055
z7b3ab38ac25a49b051c9bc59a133fc588072dbc213b3ac7786507fc629da277b6a1543d769babb
zc45766b099b29bbd8979ebd553ba27237c10edc2a0c794ed5784b038d2b82e34d04cbed50aa528
z4cda905c59c8d1767437db7514ff3d15cf54c0b74e7929d2e9978147e800835f53aa350f95464b
z271923eb4e35f1aa2cab022cfb43a392b6fa925f28c07e4c5d3d6a3a82d51cb9fbf675420324f3
z2b3a180cc4376d02af0f0ce68e27fc048082ad62664630b504b80983b2185fa3c095d1960dc10a
zc2b889400363dd54a042aa8c4e189a47ffb40c2631604404a914d70087a8edbfd8770efbab3715
z0fc85dafaa2596d01ae577987e24e903ffd0ef8b0765c3cae3d070dfaf53d132266e58ec179c6a
z4c38e0d4c02a9392ae9acbc7ae77f7f6eeab90b986755722a9a275b3084a4488cd57b1c8c64b65
z45afa484bf0bd3a21b25630072abbe3771de7c69cddfa9122cdb9c89f0b7720244e9fcfe890240
z34873094af0f6a6ae9397cdbb07cc1ce413297c15b8c2823b3569664353419c7d3e65a2cd5f1b1
zdc761f5ca5c6567ea8c2a860f02db314da0bd951f121b7860cddcc2bcc4d843fa417c7dbee4c81
z773da565423a891521ee618e232996a45322efc9f996a98146ce90174ae83eee94e2cf13bd2bad
zaad249dee83164ab4f09b8f92ea7bb127b80a0ce86eb23b86a80fd25d94506471c714dc09df3a5
z43616c5fa57a7dbf8a9a23fd67053ae64b3ae7d9622cdb63ab8422458dd204a82fd297c62cebd7
z8087273bb8c68019c7da48c63eff5e5aec6eec413703b9cf85d39fe15dbc2ac1e8a16fe5bd39d9
z12fd591f0203f8193fd07d33786d217f323ec470605500f57edca8c9322d22fc98606338971a35
z6de8ea064d5f3db171c720b0244c2e50017ea416b28422a7507bef491926b820ad9256985acf5d
ze02db6bd67825d6ba84d70d35ab60ef2df502fdf75b50d12acd65f30128fe39d6747989976ee21
z4b9c13739501af325a7a1ed19e131608dadc24a8b6b161555fd793d7fccf5bad02b3cbe5aa25d7
z88b182a772d7b127fd3c2ca03599b1c58514723711cc9dc845a520aa117820c2615bee31c989ab
z2ac87b05b5e2458ce0988ea4609767c2d95e72b044327f0429f6967da75dbb6b17cf21f56a03c9
zf82dca79368dcbade5d7b4773946f4004c2ffc42efe5db485e5e18aef398578b3747f818780855
z34ce6d3be4911e82623dc165e5192e963d4f6201db91e6d4f1d064f18109f2370ddb760dc63bdb
z05f63fa6b5735345c4df7aa7d77590619bdbb59fefc40a920ba20d20a2006c0e7633f457276f94
zef4a9c825451db9665c3fbc8eddaaac191a61e86827d8d3e55fe08e1c8394d7f77fb6d23376b99
z210caccda803842282b94b4f5fdece71482898818763b0f2d2f23a4cc66a6dea04afd66f7503d6
z0db7465fa83ff3af614cb804b076bb79f4a694279027f97b9b4a856fdff3396a2538d6374242b7
ze4938b10acdcad2ded1806b8c1cc96d09b7b77408c3b834e7338ce7d1c4e3ca05a2f7d8e938cdd
zb74599df2ea68ec2708c52fbb71f25dbfc4de2c12f51e619eaade6af28b8fdf5096966c62f30a4
zb81fa08e353cee403b68b42822ca98c76d3928e54ae85fae0fa7f6cd9c1d6cb1e2f95650f244f5
zebcc33c2ca7c6266a3f9ab65970efaf0a9b134a2df47911d14594b1299815bad6a9f9ff1904208
z304fa04f6e4f5a9ae47a45eab9c662a001ad82bb7a67b0d7471ba7a452e07bf5aa4a9a25869aa1
zd38f1913d9fc8b125a12bd93d5ea1118870d91c20df48095544c03dba53569aefed5e2848537fd
z286ce89662e39fb062e0d3b053d3e59bc5aad0a66203fddfce0acd69beee4be39c939285ea5c70
z492c88391b5842e1a459e2286ef02cd0669c3867dcd91a2b81aa33fc44a0ca7f1e596fddf8f22c
z6842dfb9e4f01970951907db12e0cb79f63a09e47f01ae0d3262d44eca247315504955df059e13
z8078b76b4b99d05605fa9d4f841e5f40acf47d3ed1b87db4d62ca76d1413fe752db49fd50ef732
z203d9e3672f0416d47f9e310a6a13444170ba3937a4864c2597383cfbe6c30fdb2618243fb4010
z2ec837b4445d66acb2a39778b466f0cc98b6d38ef8d547723f646f6e568db8eb58da7248b1ae0a
z8f554dffc3f3a24fe2db02ab9141cf7e2411eb81e687dcc3b0e7bd249e45b06a1ae7f7aa1f8ce2
z20d4fe0752d4ec1159363d5c829b1b52692442c570b25e74b2c7a4e85ac4f1ed778a68b486e5d2
zcd1b8dd7479f8f76bc9031d15efdbd79d8d4e63b38a6b02415ee5c594ef4e719ae8bcf1b3aacad
zd37248247b00faed3a7b98e6722cd4267543e98534ac2e921ceb36f0efab92270ded1440fbfa4a
z624712e522a024470d4398350715a9aaa534487cc8ffb5758301f69a5c3938cde457678131c60c
z610a4d2f4c373f573c72a79a997c2d7d1bf23117eb4ee2fe946ea22b8ef7c92f6e334e867f8ccc
z3815fb2f714581c303b3ffe704002b5ff0b8c0eafb258aed4dc2fc22620843a615cb49e6f966e1
z4c69cc9a434808c048ad5def8ecaa459402f0c7c688477db05da5d1c3692b0141ff2853d3e45e8
z76fddfc4bd2900c3f2880e17de624ee1295a27d10df6c8007fc8d2d36ae5822c7bd9e9fa7329e8
z1ec772ccebda50e1b32f88d30ef88a6c8b5cfb9026a31b4367c660bc84b08eb8382d192eaf28cf
z071ee9d486845abf9f10bc8d0a0f7909d4b48c0c7372992659ae8dce8f9a372c37a32bf4c93831
z37ea4c0783fc52690f377f1b06d41d91e9e15336705b398c2b1c74456947a1a6ffe66acaebca28
z2fe86857a80b8e6fd6f548d125cdc641106b7d18783b726592b93fe0b263ce569e25582fbd4d58
z574536b654d9bc3e4b1fbd9a0a6bd9cb5f97b2324a339ceff572ca30d3c6be823b5b3f01456f84
z047497d4e4b51f23340df3b5668a5b2aeefc445342694d92917f4c49b6d3bdec151fc7ce484123
z4d22486405eb7a8b9647c011146ae03cece48661a0d268cb91dc20e384d1d0421c924cdfeb3feb
zf0a0e0057562a8a6de1c273aaec840c9c7c7135e7158e830a886d4dbcfd8f085c6c8806843bbf3
zd5c4620490734432fb82c2b2e1a019eac60298ebf9b82b97bc4cc43785a0131bd54d57b78227e4
z6d093c4a7efd64a08754b2baac4e6917e3abf80d8d704635162c94d76da7f2ef92a11d691533e3
z7d6592cad71d2cddbfc890dd1a6043176b94114ab454100c8c4e4411c9666a8402b330b8785bc0
zcbe3beaface69251f9425d8e0e2034e8b65cff7a6014b43789baf51b9e7dc72bff1a47dba34f8c
z059a6e4b23ec1e1029285f0e031481067a7d7628d97a3e0f8a97b6fce4748226af5ab8b05bf514
z148c123d9ab758a30c2c5a8e9503294faa10c263832025a317cc0477a380070ad9b16a38ef752e
zab3d25cd2abba12f5960dcc5a78bbcda6b7629f24b2ecc825dbb94715ab3b1d24a579130572e99
zca0e36f04cd512f9e29047bc44b39f1a10001d6a15214749fdc2436554c9242658ba91551402ca
z161145267073837ac0d9859560f6f1876174d4f4475dcbf9131fc2cc696ca8d53497920dabb935
z8b5a46b02abd57af5909c3636252a09a3b28a7ac489113852e7b7b002d35b41e479d7e628e451e
zd0f36bf5474252e1a594ce62e50e3caf49593dfb5babeaba8b14ed0ec9a063ec59c54332d161af
z09b193d11ca880ce10e54011fd9cc5a96fc6110f00d4870ae6b2e2d52f9a9eb22fe1f2acf2bb76
z138a19b62a96c9be6a9890a82324c56bba330f85b92a858bbe0606992b379315500292bb6a920c
z96dffe53ac4bc8a18536ee51b2816852cbb77a343480ac1d7306fc936810e6cfa71476460a27fc
zf71e0e47072d299712f7bf3c71385ce2c8419731c09eea248f2ce2b9cd1c46e7bbaece97da6ce7
zf9b39e55ef5efb06455351d43bb03e5a97c9b64167fcae8316bbc307ad740a9eb7ab1496aceaec
z852ee8ed4dff4851872dbab1f6e893b6608ee8afc47d8e98911f324d780be50c7ae73733197260
z5e1c1ee9e10eec53d05a7d9051fba8e9cafd1354a91dcbb5b7e95f9acb8fa71736ef38241b16c4
zb2ee171d1193f3af84c354a45a00541374a8dc6fa9587b87f362722958bd7dc66b46f37377113e
z5e88f1cc889b3c813f5a892200f833e0766d532e5b974d8ad27ab6b165ccf36b8dc6fded9f8cdc
z7161cb847ecb40645fa2e671c508dc6dfc073dc2a7589d59d1e5717a416e76be4f1e2dc8107784
z583ee223fab1e1efafa754bc7d58bdf1f48e1cc962121daed57735077a354a45cd0b375d47f9c5
z76f6d6ae8d46c6490f12403d838ea57b8f480304a62b3c915b2d8fb2e685847adc80795077b9af
z13c7758f8ce7ce55d3f9e58f98e07999b2094f2523e7a53de2d937b8b2dd1a461e0f8b4a626001
z7a8688a95a7d3514e879114f811575ebb6dc2d0e13b5485d73d368e4d1abd2ce3ad0d3be16cd93
zcff3bc1aa3ecb30faab0ca64676a19fe6c8609453dc573fbe99dcadc2f6180d05a1976bc4eb17d
z9ccd803744c5bf177a9ec9537237187cff915a2c6be7c770251e6a94cb6ea2527e0fa86dee9b44
z3cde36172bc6f2d46d297425e5685f5546915702c51631a8e78e101d032bbc918120cff7ebffd4
z8120610a969f5341de1e90e19e953403e2d94687a2d69fb33c9ebe7c922e55e5ea531ea1922138
z95a4c43f7285b68511ee2a790d34741794ea9521df22c9395358c33001a01dd2bc0aba1e6f6f5e
zb7541fbea63ec34d79b6649304f35c69201bb446f8b1abfa55b5130002c099c01c8ea511ee9746
zbe548f4b364d505064e41afc43100b133b53cdfea68a81ffe472ef85f864e182dd9261dbaca930
za6279a33b8b37d48fb11dccd8ccc556f46882f88ba6773175fcc9d95f5077c1f5c18eb798fb2c7
z6e4cff5db4652a08c8da2eaa088f5d901c7d71151f1095e56c194d4db3839d25c831ee1e0ee4fa
za6aad79591adb03cb3fb983400dbf420de9443678a86fcb26bacb2dd4a817a71ce596f431f9bca
z8151076a0efc34dab082024a630c9c1fad28d52e77aec21bc840dc8d266edfea66a1ec9b6eba90
zdc7b70e083616a0881a9017631f39af77fc680a1c76795e01032e405c3b55a269c6e89154397e3
z2f7cb75c59c2a20d07f852affa961dbf3c6d1f7defc39b287bd9141469a4b55e239ec155988039
z9311b2bf85fa21870d0e1ff3a29774c06cca617901291c73337128cb33f1ed0eeeee23547688c2
zf44cbc8bf74f32b8d6ad93f5be2d8b59a3a33c91753c0183f923514bf6e04c673812a494505dfa
z70d720d0fa187ce854bbd4bc80c397c5f307d530209f0affc34d2f77e99c4ba377c24d61830d2e
z2cad28ba9a964ad9321b783bb8ae2dd9252096442a783c066046fb3f9303912dd5c70fbd1c9281
z9124048c6f23d0b9808c24d1f40aef193a5ee186857b5d5ce011950a97412d5d898ea2e1048f56
z1630e10c60cc0a651aec41f843c1660b232aeaf5fa56c239a48c5b8be26295970f6fee4d7c4d2f
z2cbea46ebe7d1a34cc2d4f244a5030325814fe20804a6596b0f8e98d359c35d5968ce8e582968d
zf6717d36eb31d9d08391e84681e5813b7113f233d2e126d8cfa47caaaecb13057fdad71f59d868
zbe3ee46b188db7541dd02f11abd4fffdabf1a46689e84f4bd10f3d8fce27fa6586d95552638f9c
zea93436388844dc297e0ca969b5d551ce60a4971eb49048aefcee9c6a2fdd0e07e66f585c84e68
z31b5fdbcfb8160a10c2edddf69263588f592cd1b1b000a5c4eefda3876083153b853b6d9aee84e
z2833de15f4f5006ef9e217d28439095e18ecedf510e069230c8e4807fc4abe66da28b266e713af
z8e110e0752452a8ab7e28f22cc5d52bc760cda7094365731c38ea024837160a6ad02d563e9d17f
z5410e600b4fab330b05c247161c52fb3f91e775684c1dfb6e3b31839995a53ae8acc40d3154385
zd3735902b473d9baf2c370962bfa40a630f9f2aebaaf02fce3c525858c13f5babb416a184477d0
z0fd15ed1bd98dd270ca14cc343b4ff7fac7de38a1fe50e0da9c7257fe4f941f883eb7b6817a544
zaa4127aa427911664d97ec942f984ec3fe427fe67a0d0d9536783c71556e802951b27d7767bc5f
zb56d63fd5f606c931464e7a83569ef918bb6a771dba0937cf6ba440d820b7cbd8792c60e06c270
zf68103c1d515ca6d09d627e792c3b561c420375684bdd6bf744b74bd565504179ea892d3252990
zb3df00cb946d91ae16158465a735440ac238a60dcee436533c5a66dca36242a31bc514e091cee2
z4c382babc915f070beb0d7ed3c93e78b2cdada17ddbe522c3de2494d9fdadd7e7941d0e8682697
z431f12ac9e0f42dbe023cf256c5e75d3c8ce32563e631dacf226fe6fc4f84589b43b819ebf185b
z123d9d48a118d7bf76516e37cf89f358bbcbaee27fe026a088091a5f65b0c9a9db587607005aa7
zfe29b98ae524eea3ae28da231251776b1c1b5f3c80c8d94391bcc1bce655dce4758b709497a3ca
z5ec93926cab042a7244a5c1ca5dd006b3a1b0954957275e1ff780f64f79b932d43dcc9f5410108
z59c662ca37c58102fb8153dbf5798a43e8f76184804156d09a2a0b75bab8d9c0211ff9457344d0
zc72e3f87b34c6d911a3630619ae96297b9c22c8baaea0b28d2c4bde6d94dcff9eb67fd02d95e03
z4d2e1cda51fcb46dbe040329d6a98606d4f5627ca7c1ff96575b57f03bfb6f48f32d4cd1034915
za1a19bdcd6fb8f72ba0cfda68aa006300a0c0f24515da82084fe26b0f1e312798fef8a979d6231
zc1d9db578b390a98ae2b727e50cd3cbd7e2870d4cb3fe502153222eda10e6edcf43ef4b021acf9
z15aea519a4851f7164c490c5bda6f22711465ea4ffa71a7af81d7afb241ea02872f23b78c77748
z84ee7953da89a8ccc5fe80e418d08ec9de1efe670fc57bcd71b89d9aafc9cc91e802ba0a0d5c90
zd2e954c6031f15ff26884f0c0c8454d61ed6e4a7bc7bb2b71e0e4bb943d59620b2fe581f404b08
z291c669da3ebb9003d4befea066d79b4ed954aeef713b1d432751d84670c828fb5043e5a7a58e1
zf4d848f530023c727ad968c29ccc8f4ca8d7b2c3d62627fe5f82f91573c530ef84c98baa31be36
z61fe40aad3f1bcdaa9198833eb50a613c73a2d94238b60933c337d17ae97223dfc2eb51bc3d569
z93d8802a5f51fe26a6e76751d04d1b0de2e38cab5f0117cb314581a801549ccf0a44acec67131e
z1e705a5d50d9fd1e1c67e90af867db30d8f771f9dba9f9affafa620a051e4b23dc0197ea81828c
z444a857a04cc88b2eac81c2cf111b8b90c0682142e34b0625db4b708841b13f3a08512558f6173
zfa77647f409e6e874c60b0c934f1c0f2accfac9ce083bc68de325a343f2efa1da65e50e0a70ac9
zf341b63aa8187455f943a63a432395b214ebfbf5aeb9559e47e6eccabc31d0f63b9cc9c102c231
z9c6d7966f295b66206d1d70289b41a3384352d923246b25d4431af67daf1b3cc36332dde40618a
z7b31bcc96f6839ca43c8b8712ca6c3edaa412f6db3c5c67b9e9e043cd3b067b68576751eb23bb7
z0bc6001283212f8c67921ea1fabb4d4aca8cde915110b66000fa6960afdce3bfb7aae1d2dfb698
z0654bf9578491632d86053d3a8f1b1720bf4956e8acf6bc702a9b4d0bec020155c0a8e43e6cba7
z27e64b9ffb193169277f25228cef3d3a6bfb06a4ad296f7ce46d8f266593e561e71c054b9fd9c1
z3e0e21a0dc0b2b6d56ab4a104ff9e02db3a7836daf027268d9c66422f7d6d089e9db7fb939c659
zdecfb3bac6a8c448272db512daf32c167d3185f03d92fcb29637910f813ab6534bedbb9a1f9a90
z34c7dc4d131934f3e56681ca8c80abf8b0f6bb82545f2b9db7f635a58b6dff2ce314f3d7e1572a
z1f0ad139d0b4865489c8c1fc6e038454cfc1b8ba3363f7075d3e599f703ccdd4c1417036ed25c7
zab7fce7277a0fee3600a15f02e026308721d177ec7cac17ea562ee966eb9df7de39f9869391aac
z1421799fe3c480318e98460275e767e38f98e7556faab4186d4415a3cb3c617b5ee0fc0b4585f4
z5290a081f1a6c56f4da18a7d6c503750651c95f39535de3b62ac7a92a4db0097cb93f7f21a4be8
z99da33c30dc9088b7bbc8e01800064801d5fb33431ae4b01c9fd9aaca3961545ffa78276ae82ce
z9a207bfba4b987aafe28ed91b1020f81b10325b31e69a24a3dd444184c6e0b5201832a15c2a7e4
za9151405ca6e3cb1c7a7dca97a91d617e2dc070b669bbfb7a6103d77f9f8b2bd6aa2acc833856a
z3d5357e86420a719a12e292e83919ee77d769dd705797a0a298fa7da9a1165afd2ff69014d2b59
z90e5aa2dd9ce957a69592d0342d1e06b300cd25114fb3b30c9a39345be7b4a058c914c14f35362
zaf3c457521e42a1d3f0294032ca608653088a7bbdea654e0ff49eb16c599a491751132dc2d1ffe
zb587a94e580d0b0180ac2a4cb2da5e8ca7c8c2b61277ae9be16bfebe4500615736890c43dce53b
zc7ead099fc5ac3a2b53dfb74aed71bc46174c98492fdc09f3af563b46bd6acb30315d38b60ad96
zcba97de4945de56b02c8f4f44911aae8122184147e2ebeac3b952c8f19de16f55c1229a96b2ad8
z0e45d04b0e2818d1e4d97cad4236af0546fdf5c5aae54f658dbae8b79a2f62ca6ff4e031322b00
zf68515ccbc335130fed8a02d5467d2149a29e557d5ad9dbe6a52ff325546d8e3d90592ecb7297c
z6c0fc573e9c943c46b46132f7284c506cd5ca3c44fc227b3c78ea0abb8fc765fb5594ef1794423
zc0980b027aa6ab87b81757ce3840cf2818b2ae1b0916a70f7b7343f31f157db03852676e0f1dd5
z883cbd1c37f86ecb23d083a2e07443cb8aed8703eb511ed59098887f07ef1e307d4ee17780928f
z97789031aec8eb3c3f257037ad482a4a880045fa1d94b582f9c65bc11e9fd84f142e3fa6c87a94
z737069aa1e7d426742298dd85f9eb6351b0fbdbb1d2c82b1f39bab2eeb2d9cd505e7f930153496
z32e2cba5cd27692a15dbafbff614f9b2ce81f1536bf609eba9306b254aaf4ca47335dcaff8d64d
zc183e3ba262116677eae4c627295977100aa21820b3c8b8ccacb1264f16bd220822327125c8464
zb0ffac0117a07e319fe2dde49c3d2612b689592ac2dfaaa277cdd7614e2406407e8d35921fb22e
z9333284c7adde673e5b12c123b3c05c227740b4ddda4ba9fa2d900f2662e54fa709ab3a7a49ee5
ze2a9d33be1766193caf0433a02e222f11e105a61e163b2f5636844a8285883ef5adbd51d71dd82
z1988f7d2dd15fe16993ec707b725fa7456f78961d6dceaba343b9af18281f3143e5263c3db06fe
ze6cf153315bf6be773f6c5d50aa834d4e275e2c1dd1e0f1dd878d250883bb78877068ed1b2d3a1
za786c41f5a825a5786c2e67b5bc3475aabb3e69af5077521c6314007304821582793da55997601
z9fa8fabf19d058d5106f6b3935bea720cef4d0012e89295d55747ddc47272bbbc271285566368f
z76fc668e0d9596ac607df4169d702b6efd245a2c3e2302d46fa2b2b56aa93f4f0ad71a1f2f99cd
z2c8c1be78763627c24ed6259ed65e1ab2874e9adef213be5cc406da907c5f425bd5095cb97ff42
z60e25da224ecba7ddd0c7155ca3c97c360d52a94a461b6fae12b23234c779f9b0dfb74827e5c1b
z91214e30cf1be33c4d6800b126d07a2b0020dfd0ecbeb2f2cc050343aa48913439c51bc91b422e
z54e5b54a562b3495a51bae05bb65bb589da9cd08499c22d0d687f554307a58ca81d029128129dc
z61f35fbb01a312b477f3aca09ec499ff10da867df19ac027c1febbe1e0a752a12fece42f8887e6
z49be8e5d4a7fa6625aac0bd98500f83107765362c8c9970c66bfe55c9bfb044daabe0c01565766
z70d95e4d03b194feb22c4503f14538dc2c9b32321a53432ea06031171664ae3f273dae34fa614d
z904839d528b8f6fd74f213bb42f9f35443dada5d349d1fde878964ccd5dc52760e7ba79bfccbec
z465c411aa755385eeb106f3dadc257f44bffbba578aa2b9ac64afcf461c5a01261f890c2fd2a3d
z5e0fc3346f0743fcb42ae9ed4f88151f930a8362004a6352202d2ebcc35e3b3ff831259026adf5
z46ab3b10a798c7cd0e811120e002729d08b04fefa73578c17346b775bd6f2742ca4b6161b3bea0
z8b0b8f1a5e687da37a151e9f5bd2dada888d79402c2c832997e94177244cc01c05a37ecce2abd7
z82125c25cff294b36a27166f577cce2fe37f928faa1382e089c2e7cef7259c848f8b4b4e956a32
z5d26326cd4e03fae3cd37f47a93deccbb324a7f6c548cf26774da3ed5161d36a95d3a99b10aad4
z437621bf0694af5b670fbb9b0db0dd9257183c96a0a4173140bb129278d9f69dca0d92ffa1cae1
z0a1725685b6c19eb02091f9c515ca6cd31d69064fbe5e0fec2f855bbb33cac7fe0b3bb1322bcfc
z59a7d9da2732e0055907fd33dd9b385ee8b041207394b67215f1112667b9f34e2045ecb5d82ced
zf1207604328e1bb008411bd64b7c6202f2f6220bfb057d04d69cb2bb21f29e9792f583c685cc37
z66f043692098cf116634fb1957c0992080f9e0b6a314ac9fadbbf605d89db6b13f73b90c1b565a
zef1ca471624521e85cfbef0603282421ce5fa1b6e2187eff795ef6cca00eec0ffb4b37fa14e41a
ze919045275fe2189b6dca9cf0fa5aced3cd19fd23116f75c3c0e8db12ff7045319785529fc722f
zbe7cd00484d6c8397c9dba8b536da3536c2010a98a5a926e73060a4de74225db4df7343b30eb40
zb6e71fd6e789ea058157411ecca51ecbac020a4d95e2657c2a19a827bea25df04073154bbf673c
z0668f34a82b543582ce59718963927d4f0601325d84e8f0482656f2c8b220cb0d85e62e95f821a
z8f4d4160fa41801c4e3b2c4760c173af193a11555c3ccc5ee33b8d2356ebb578958de2d6c3e0e1
z546bdf44fe04189191ec8a5e458287412b7500817d92e6b8bf364e232beef8f359a2bddf31e2e0
z44857996e08a34f7a8ede879a71166606f45fb420d558452a1d87a2ec425dddad2621ef52a0225
z2da82f54ba00b4b587ed68203e8ff206cdd4cb57693fcdcc2840054185f8cd4f288e7a159730ab
z77b47862d11195db9f8ad48410d5d7ec4dd568b74794ffb65bba461176f4d4d10671cfd8f334f1
z0e718ccb8a2e53578bb3d650eb966d4f51660bcbf8298bc3a68c1360287d8f9c62e619e6c16e51
z2420440b0bc56691dff5f23818471e41d7cf4fe9e267f739f306368ed6e2e7ac60f350745006ac
z2b17dd3f33362de80998c816e29b14a836c421d46cd4c76667cbd644bed9017cc2f90d198cb6a7
z03e5feb33bd566dac36c3acf8a5b441732b6069728f5ea24542c064120f41818bc08fce0a7b3b0
z70d8078e385552eeff41cc108a3f1daf95e1a20ba51c0a1dbcf5e6f6f40eb3b2e744b5442a9a94
ze7bf8006d42db79b3f0ed1486cc4a910310aac7f37cff16f4c06debdd5b7167d6dc153367aa30f
z67bf2c82125dcd8105dd252f15ea2278899ac54a24e3bd3d8a7b2895ba3f1229235c4eed6915ba
z9fe34108739c26f01ff8f610c09c3f752bfa1ea02840b339159c7110050b4232e4f3a23956b7f9
zc2e51fbb213bb892e8f62abff5cb3f55f07b21271f3c8301acd4d4ee6ff11f86d17f9b0d18f2b0
zee51f43ee14f22281af3642808d6d6607752252115f0f1d94dcb3320df6faffd7cba01c37e03be
z6f2bb5e5ccb14eb075b94ce53cc3bdb93a0a239f56ea419dafe2bc7493069227d3cce5776ca11c
z9ab56e961b5215b597e75d29ef701f66dc99be2c07f1c1f978a8d371c78c7a2713e9c28af4978c
z6a8c2e073796c87922236805e071576898ce8837d59189145fc15dfe945d618ed2da38de4db546
z56967e69ef166855b1d22ef3bc2b9c16b1c8294d834c32643c23c49803f512d1079583281d96c2
z85f1632e2c2557d5b7d4a48e99096aa37fed0bebeee8aca0774da52187a1614eaa674dca5a2cb2
z4e2c98794bd47ddc190661f8876cf1849bcb24345bb1e7b9d7a5762f50d622b6c863988af40f5d
zfcd3a530487d3e27be9d3ad4e07ca83c2adc552797f35f0f6a45c1e4bbb98be43f9683aa1d711e
z61d8464f88b2f2abc8a030e45f7eb14c75597e06ce671220d58fc2fac94eabf9453641d1471b35
zd97643bc0dafff5f29e029b82af4ad5e266fa5f2532125f19443e96472c7e7fd9fed6846810116
z02b4370b73e560577413c64cf64d413e42e18a99cc8e48521633c11dcdf24794cef946a90a5c16
zd3b5276f660b508f1cc26e7e2a1c2d263364b9377321b4692b51896e0b5786958349bbebd77244
zabdb0c50c8481eee8ab26b85e56dfab53743c22f6cd7c4f1c1c2c5d4b03fb26da1503d2d77eb66
z19490ff684c2b3c88db9647f3122ef0ca8fe6483666ddba77411c9e32c3016a87a0a3f6a78250a
z3622c0d26383b9e83c73320d1397d2c9211cb5cf28ebc0c069999f452ad01e5fad3469dfa29fc8
z35630fc58ea9723593c924193503564d48cf85d5dce7ecb225327bc41efeaabbe37cefa0dd7fc0
z09531d646ffa0d672604f4186ae4886b8f97ef4e6b73ae0fa7526a319e6227717b57fc3eecd845
z22cea5cac132586454c7c3acf7168b756a7e8de57424f6dd149dbb72027e2fd4f746d090c12181
zbbe42697d0d3b0bfb2621d3cb0f3e59b112c600443799e784547fa170dbac310c70e0c4235d62f
zfac5124e81af88f67a6ee0f1bafaf6fe134a111bd2beb6ade64be2326f23acedeb0cad88775282
z23ab675ee9d434cfe79191425b1de140b9ca101dd8d4adf86cfb42d0611a3b4ff67978c34c2b2f
z1a695b679cbfee9b57f4104e9994c7a12a5415371a68844a378c0c090219657a5d0a4da956148a
zc1c8d39f1b9578b92b21df45c8f5e174f67e72e199a847ea9c9c25c24d2e9247592338a9d6d000
ze79ab09ff526784b89eae094275ca71602ab469c7a18443685aeacc6721606d357caa574cd73b1
zcf1fdfb2ea9316b95efb4182e3fe36a4ea62fca2f48d950e0e5c0e769e71484d6737a830f9516f
zcc50a1aaeae9504d2d51a56e9fb4f24065afc197883e2d2a92b4054446315314ad72f5afb77cb3
z6524870335d14e52867d65bcf3dd18a5a84e0762a4e2d83790c545454e4d1cf21248fd4e756c4d
zefec89a784751f9ff3f1944866b9d71b4cb727324d3b60cee49d79a654d032c574e62ab82fc95a
z883c20c1adab89f2dcae068cba08516b33e6043b5227e1fdab7f1a024e6aae9078b1ed7d284337
z176e3fe27d76c5270488b23707edb3da7bb80c6c5fc8583cce41727486a99f1cc2d9759d3e8cf3
z2873ad1b72bb63352bb4e48c12d6b7d69e34f9005409067c1e6fab1c8d309bfb3dcced993ecce2
z4f5dc1a75a069f548f2e066cb6b9fd489666bdb0a52ea9e28b2f411c154b6d72cfed97183c62ba
zaadf0589d67bdd99b1fa6d156ba6d7d6a1d81f0999fa819e8742cf1582522dd16c0dfe8cee6713
z5018dfdb5a322c632cdc70fe8475f11cd9a86b4c70650f21b32d9fbcdc541f3b2cc919aeaf31d8
z54fd1206b1bfd9604f939394d61a7b8002bb8bca6bc5164aab5f8d28b2e2fe57f11e9053950737
z0f922a3aecf2b7598b61b29717747fe0379e5cab933bc7f4f77e81b451181aeeac345b2638a3f0
z5906d723a61e9ad6aa31798f07c84139995d6d20b8cc906f1f6bc2b382549d51cdc10f053f7dfc
z3ce097d5b0fe13d2f80369566dcb22b4dc1e9fe1dd07c1dd1f4edd0bade46e0dfbdcb97ed7e8da
zad24cd54f0a9a86bd898218419b8d95a614885ef2d851903317cf37ba27a613ffbb048a63c2b94
zdf00ab8e22b065d3350298cf3cbb6efeac9070a6b951dcdacdf60480de4b5b43536282adc632a9
zb93c65aee144c68d6edf50089415217fd2fe72931fb30071ecc1bcca9097a2c65f3aca85a5ec63
z67d54d8ff8e9c7b4fb3770eb5315d4c42ecc18cfd2fa5548a913095508c936c06518a75123f628
z505abbddb7ba7140b5be491cedc5248a06e3b1190201362a0ea9f87645e0a24c1ab47948433b8d
z2c29eb12cea732cf7f66983a0db6bf7c139eacc519b34d4a1735dec902b6793b1648221ea6b0c0
zc80bf1cbc2d5765419b96d6401bf036987c0788b2b0715760d44712547a17c6a9af7c56e59fea7
z9f66ba23c2ef88fc3d676e4b2f61c00a295a0d90d17ae9d3e69f0e42472c84acb8d7ae18a701df
z02ddd24247b7a7736500fdd33e6a82c28c9d7d1af8a053844dd26e45d6d5f0355c324dfd6980c7
z422295d834edd0b1ddfaf30606566129ede0e6f35c25ebef6c2bda39547450cfa2ea6bb480fdf5
zdc18e74a936c3fe51c277a6e1f6a4ab83db9c370ebf3c29b5f26d3454f99cf942e710367d3c8ab
z8e12655e644fb0874dc336976305f9b6370be35134456f34ee94853b883769ef0819b17fc0dab6
z461eb208a2c10e0c08c29c609a92217d9e115423adb84cf0d8f1bd01f967d32e1c69d6e6c3d874
z7cab74fe3b4a8be0197e242f67480afc98ed6060d942a1ab7d3dbfcd311aaa43b824077cdec788
zb02548c54fd8750b9432b21f188061968c153746c8887ef608bda47cd9dd26a1dcf1577d89ead1
z75f67bca50ce29297a0bad554ae600ac0371b9c0b7c56e22c9b93ea7b1a869b8bbe2cc531ff5ec
zcb5ba417e736f796cfeaf0b6572e059fb873424c17e296d786151c40994feff03f55b0ba736a07
z5764cc6c8da184e1325f17efbe14096562497cadda3633c075a45db1115f2760dd8d0618edb0c8
zdc18986dd6d6d5e5848e7d5f493f219bd84ac658b15912289a16864fb1c34d83df5ff64f34e37c
z923389222cd4bce7bfef649cb89f9c905102f08e3968e704eca286f59c4c1d9bccabd2f3d47a34
z9a0e92030511e076c57471286e7ddd1f1b63548bf537d2f42c49feb8e07a7c61a357a8d5166386
z6b5ce601d7a43bf248da58e7c8d5d0e68fab9a1b8d9d5efadd3f5924c81aa165b26960fa44e0b7
z2a613677be8f94c81ae8f2b293e24dd766567275da1f47f64ef0111b17b8e4b6743fe400a65ea6
z57fad7530ee1d728e314ccb489b0dae9e32c08aaf70e52260332d88ae044f379f450ebc99baecf
z1bc5329e675a62e145ba5024cae9e3cfc2a34d6200cfaa5c3e02b2e823845987e614ab69636823
za6394e2f2508aebb898f62f0ea61a456108affd5c8774c5f3ca02b369a42f01ffd6d96eb862718
z36532ff9ae2ba838a527e07ac537dca6c4a50810d01287e4fd583a61ee6075c14e3791ae043fdd
zf501f4633267ddd6e27683e14a9ac23c3dd8ef6a4017f236557339785161cd598b4e162708ba4e
z0fc1fd257b0f4035ee8184222e8972eb0cff09800e8124d7a7cb38fcd28f071508486382fb1b58
zb5c608fcc7a93e1b18e0aaeff0a131f5bc25b4b36ceff30c261b2ccceae772913ca4e085d53bed
z10dc605a87d8e8be673521606fbe44873a956b17b3a7bedfc8ac93dabed86d956832f962ef786a
zcf277b9e79d8d6ce3926905a5febd6dc11085e335eed5567cb9d7561f92a4f5c3ebbc1986114eb
z69ab8ef88019264442ccda3acc2978583e3242c2f5d808537620c8d03a9e3b9348df70cea9c14b
zbf8395d02ce77cee804d5d3a9c8db0eb1638d3b9582db91c9dd456b4dacf78753aba13126049ca
z61b2bb1cf10d77f56028e15b426d8d176fced5bc0a71405100ddb312fc3f75b6955ce81c9ca5c2
z3f05fa85c671f398e8db23c19b4ec51baa1833f09c5f4715d96147ac5d109763b7b79dc8bbe473
zca8b32236ef694fb77efe9fc8f638241cf4aeb7433209077edee08114d59121443ca1c12bf7b73
z16fe5731452e82321ac353d15309b1df70704ff74cfb5a40a595c9aafbbc201c849f6ff5e37ed7
z4d8af5557c8e72109400fd71e369c22e0eed1fb49e5ff1114a7832447d631e98934733257b3cde
zb89c7a80f67becfe79d9941c40e82e21d5923410501df6ab2945a05888ac163a410092eeaea85d
z9d39719c3c883f1c525f272aa6b10e16c02f6ccf3642a9a42eb2ff4fd2eaa98c8fa90b75356bb2
z58e227f33244b854ed0eb517758b88e76f061c2aa2e0aa033d005d494ae4e358c2f89eb0f26072
z3d371a5c3078a74c7901da4bfadfd208cf576a6e1458385e0dd8dc2ccc2ab72f47aaea663d9bc3
z4e3c8d82bb2e1b96caedff9b921a9594cace46a455e6c29ad59cf68a18ccfae6f26a61a0107068
zb7eb86951e2639731d262df8674ea8ef4c3d106a08b6e8c44249e1ea69f8764cd00b544ff3fef5
z5a5b11f44c7a31637cb44acaacb85c9755a8a4b6dcfcd556e9bcd7854c042a8abab9869dc5740e
zd5cb28b01368a5520960137b096b3996ace52baf6179a887ee6a1e43119a997b6a81c736eddf52
z426a8b2642a81aa3f0a05b8e8e4a6d6077dc3509f72603fb3ff52395a9830e43cbe01fb2f766f0
zcce0ed38a5405add1d7e038db9ebbd70ac251e5c70de370d9b7f423da0180bcc1bd416560c19b8
zd69321fb017c70d3cd7c922dec872c09ba8bf2922ff655aa5c2470b140dbb48204c10c88b4c4a4
z4d507673eede462ff6159a99f8ffe53b68fc7019b917e8c438e6fc0bb1bc06c262ab9f30f5d6f1
z557b88750a054abfca64f15e144a4ae600c6ad77443342ad02a4ea71137dfd9053553928fa8b23
z662e05b5c318bd342261085ae8e758fc4fa5ace7cb07568205bdc6b09e8af1d9ac9f55268f7b1b
z272d151e10bdd1b9c9ea2d63d51d0e008cf3811b476e05e1565dc7d8b1605266610a59c5b341d0
z9768727ba1d06ac4f99ad998a7a59f4dbea50b4ab69af3115e32b110562164380457a9cdc77ce5
z4929a52983e37f80e61a62ec81c434f7d601c85013195a33b815020d308a37f1e5f77dfb1e83c9
ze8d7693f47663ebbdd702d66524832181413f325816e72fdb04892bc64cc0bd51343b042e2333a
z90f675dc86b89cb0424bebb8ba3fb4bbc17d6e25578a81174fa6967f06850d3b6c9e7ba35f2f19
z18d90bf70a1560802c21e0638ef259ab3c1f655ead61524a780c2b6ba4ebbbb2666911b00e9923
z93505c1678ecd4ccebefdfb3d0b129b2bb38df1c5d7c811f613bf163dbb7c45b21ba7c920d01c8
zab050ad188780d242cf177bd0acf322d92031eb991057e17734f0f8c7facad0f0c4c149aa5ed41
zb5adfc3b6a67c6638ed0251d68137a638f4bd664aa50bdac174a218901486da699c26a81cc0414
zf18d3ebbea9a2919dee3017097d7e1a8b7af30c3535f910646ac124717e9f1fdeb0fea07dd65b7
ze16cc7ae166e14aea0e56bce0e8a9307de0c5b75754736d381aae2ff60d09c0941236a73b0955d
z104a478ed22e720060b9c61f30b4fb8be348e9053154771a3eab185f03413c6a5e2eccbc4c3a2f
zfe87292f5e4dfd64f2fd7fb3ed33ade5ccbef3d1f94cc148210a38956cd67a5ff13af00a00b2fa
z3cf541663f892fd36cfac4d2635758f6fc50dbe83689aa2b0dc4415d98afcd545dd7aba78b3120
z44720e75d0b6ab9c49fc4743bc16009ad5f9282dbfce1e796cf0b2243d3032acd99d58a229e1ca
zbb3563d33551c9a263d6d42bb1a969f55997ebbf6679938eb89a0fe2f6b7b3766ba58df498149c
z3feeed054f1682986cdabecd57ee4097434a23c1699ceae9f8e65ac67acf5d2b3c09d8f898ceca
zf6a41fb7fc2bf338d0600fbc4510faf5de858e7b77d147ea349e40308690b27ed05039c91ad3a2
za905212861de5fc455e616107d898a5b131b7777774adaddbcac5ce17d9720b8a466399d8d956d
z9e265913bc6b95c13f5fde2785c46927c6dc7e7221da7791eb5da39bd84e1540712007bea58a59
z7e61883be748eb22d3436bb1f1d80c4405fb36af7947e5751d1e1a06b07c1537cd8057b4ece4af
z15f32b7dad67aad611164bca1fa4e496afaf28bcd513a9e0566a28134852fd0d66a2c5087c35c4
z63185f772136532fc3d15eb14fa9e71c1eb2f51b86fc479ab813cfc7cbe867fa6300cf5d7fabe7
z7e014646a0dd2c647cb7661c202c7ef61027e8b4014939e63283c0d52e31a1b53153cb3b2fab36
z8137aaa7828e31334165b04854353184fc372273f047c98dc1350ee727f19d3ed2268b76c93716
zf1bc89d64a4c17f740d0986e7ffbc7716008ae28040713e94c4451c03c2c02677fac4baaebe0b5
z484ea9fb33b3d3c51a257c04f600e3dbdb534b924e8639ab2a6ad74a4c47f476a9a18941331a81
zd82be6ffcd3183cd09cb5c552f7bd50da2d17adf82c70c7af952eabf773b734b5f617b94d5cbe3
z8303638bc0a76fe7eddea645760060a185eade44866d8524fba38a9f2fe9cd5f2f85656add2b9e
z5df319201004973993b401f74978d5502a01f0979248b944b40a93ab433a1e7466da46017c0d8b
z2df252f466cfb618bdf1ef121c9a56d0a46aa0fed205b9447336300737ae3ed61e999265f188cb
zf5fc9cace1e5b0efc99207b9ae549af0cad9905084fb88b347489d4171b2295010984d53fc9190
z6f0fa8bb809ebc6fe5f01746678e1309b639dce228e8beae23325af9d40d2e2f33c9e8c235e2f4
z0bb44af4004073e05a3145f07d49af8a322392527ddd1f7e3d699ec347c01ca0886dc5b1e0be37
zcc950436c51e40a119c8987bee601ae477ebfa9b4a2b6ec5138304ec07a31471242fd5db4d474c
z010823c82cafb38bf164b11517bf8075c52eca76c2ada6072de1a05066ae9a694522ab8e7b6bad
ze363edb5bf784926765f7f5a1f9309778442967b8a10e34f156f3ac87390216ade93eb1439a5b9
z94d2fc385a370063a46900a62c0a76752d8b5f9bea6f076d1f58b2c71d7ad5a3832b2855ad8f9a
zee2e63b7571bad124314d4541374e8cf9eeb4ece0457a242ebdb1519ac63f589bea1cc3766a4d4
zd350ccb0d8261c8844100dbdc80b7134c6446782c6e13cb9a48761c4db78a91e08bd83462556d7
zfa6902a6c2125cb19b0e4af2742d152b3503149a247de4f3f0bfdb7d50c88339da0fc565860e89
z11eac90465010cca6369691de5c606d6034ed6b64b8106a64cfbd815c33025bcc1625630aaf3ff
zdcf0801af93226bb63fc7a04bd786d4156bf51b3dc37b3393ad6dfbff3770004bd4365d02100e6
z6cf784ede3339f94d813eed55ad4bf0b08aa5df0898dfb35d149df3abd9d9d85081fa59f79e834
zc16d1d1f4132b3bc2ef1a1741e7747cd10fc97449048487e1daf11fbb22b5f329b52e6996f98e7
zf4aacaf5a547124b9fb2a10384529bc46d116102b0a28887bd88b54af15105774b6eb7ca431847
zd4734e2ae5b033ca4a7030343988066e27f886b05e42c23aca30a6e3afaece5964c1ba0b52c4f6
z602d48c8cc3ef4aa208658ea6531aba5608da4797be3df26cee3bc0ddfcf40edbf9021ef5ce617
z0601fd93a5aef094350116b9083e771e9fc4e0809b91d08e8a413bf29858152aa0f4e4d9e4d7a6
z7919d37670e11d7617666f372da530d69b940dcba37cd5c3e3866d9658eb555825e4c269bf6f04
zf8f6d154cb8f3dd6f6f8f6fc816ca2416badf1a94009fe7dc97353ca1bab95c6d9a9c1aaffb453
z45b9b649127286201f209061ad56bfb15fb3068d7c94ac8eef5bd5b3749d945a2bfad06b91713c
z6b37d491da8b3fc210ffe357c22b6adef495315079a953d6314c3a2e21b6a40a9c88730be62d84
ze14c3d4dc1ffbc1931fb27990669b9aded1af6b865a91e7bc04470d418dce608bce88149c94e07
z0e7e8103505b62076bde14369f1f18fdd178c297190bff27f91b0bb9f7dc5a19f32c98f1c19a3c
z6404fe42961f28f3490e5f34a1c7426c5e8fca41a928d5fb8ddd6dcb895f64266da6d2d7a2b091
zc1f6707912b753c09d991b8bfba02b87fed39815dc2fb4515b0618fa711d63a5c4ddf8bd795a01
z6528343c1f0633b0ba1a191ce70c2199079324e6c5c8d788a1fa28531356f2acba6df23b630c59
z2466fe0ee9a40b0d275641e289a70a87d9c0f898caf14a9a5981b7170f3de5aa00b0c6ed9ccf7d
z99ffa61ff3dffae175607c29b9bb3140682347ffb30ef030de0748975c5808729b5c3521260701
zef515522986ac8bfffcdfcd479f631e3b699ff2bf244ca9ba8faacf38da0a0510336b8c720a625
z90117e06f14ba3f80bdf7889592723bb83a1dbd76453c12fe9571c0234cdbfb43e9201dfa56cfd
z41acb82420a53a76d375e228cdbd8c3459da1b1addbe00eb34fe98be9b6e01b51668340f782ec9
zbac9e14fec105859c26dd9ce0853500451f028c03dd2ec0058279fd58e3ae69eacbcf5726b4d32
z1611fbe0b2e6ade3e6aa0fb3a6d1422a5a3e9bf9548370d997c2003ee6f8dd02fd59fbbe25b676
z63d548583f0d5f972e3f6fd4514b3b20d1dafb0559aac06bf49d43263452881db00a7df65f985e
z5d2a28463bf810556e9d88a7a3c28b4b3f8d6a7f9e2420ce3754956f97a74a3254d6fa51285f67
z4e4ddfc18956c2a4addfb89e57038f32293eaf79bd6f067b30a514b86dbd1da9eff1aaddf341bb
z350b71ce3f6aefbeb48a10863c66d1d7072ba4df8330778ae9d7aecd2fb0501219e447094f8d5e
zdf5881c51689b58ddc5a084fc4ca96fb37c3b2a3fce6b526e89c340aacc7268f6a0e54bce34d17
z549ec77764377dc2d06e54bae7c726b3b1a31ad1380c6e28b7c2d5cbcbbd368a639590be16ab4c
zf169a168602df576f26892ea98d363055b46b58da3e089c687a2d0d1edfdb4d9a0316723fb79bc
z0e8a23c73d89233407c7810dd616b47b63045c4e67a29b89de51b0e8ed74113b9ea99853baf7fb
z153a691b222379f4f808198229cf114ff80b0c1cd7983a2974c3dceef68f29e6aa5244d5108b2a
z145b79249857003d2be8792021a4a3a66eb97ac2aaa03b81ac3e1593155e0de210ffc64182f2ac
zf04c00269df20d7c8dfd91e222689d75101db95e815449f0a9f2e9a08dd7e81e264f72406e0981
z1f3c8306c3c5aba17ff03014e908671fec2616c3d796026d6f56523ff4530329df20001d8dd6bb
ze9776d03389f82f1726a4f589761bbfdf67bae2ff9a10b03d6f1d481a513fe59324a308e0ea0fe
z07a2dfab079ea907351097472204521cb6615632bd74a970ec7f55ec6e14fc86d2bd3a819247c7
zdf6e9cc9d95ff072cc0e7ad5cc191143a840af2304ead8da142f4c4e8d6f0b0c531bcfbcc286e0
z8bf396a921f5120d2f08a859b0d6441be83401618a243357488984d162641a83f426b36a1e40ae
za9034a4777e917b6ff53927cdfa919cdc48b9b482b8dde10ee3f9376321b92943c641af297022e
z506216192fa9c0b16b5ea0b04c5e5c0a7db4adbf6a51a31c256436add531fea53ab14f830cefc5
zfbd40a0ae0878751d29cad43b9a7a610a7c5be87cad13b6e5480be40263ff660d337bbafd71e99
ze790b71ccdd1f04b03bcde42239f7021c9a0a7c1a6f53699b54e274a8df61529bfed377ebddcb0
zf567761777d1b8e7e4701f05a0c5eb6d55a616ea1090de34a5e3808968773576abaee09a9c525b
z00ec5a37d4b1ea9632d7d9aef6259ca436fb16432d6375177350d4fb20f4a7e6e72bf8876a6c32
z069ce6be6882020783b62f4365660c10ed577db53faca22991419e56740e9e268ac588f14f9eb4
zc4ad84cf301560b55ea0d415f54f2cdb769fbb870216e153bc9547387607da48f0388d9c2f9374
za2e38a0b3bd4df6d1fe48c6d61ffca2736964f2e87bb9dabe8411f2b8ccfd4bb5ab1a9e7e7d54a
z2f0bef891872ecdf31d3a244b729bd4037d7acd349e097548faf987358dea6a43634e7b7ecb6b6
z99f274e28df54dc6377951ec22f8dbdbedc0ede0657b787321210b9c342043269abea72d587e97
zee1249b2a745e3cc50c92caad5267e9c6afc1213853f7cbbf7591cbb1c8f17fe1a8c6a3380a331
z03fcb97f764a4cbf73372d5081a6a08a7732bbf9c4ea286ad964959f204a80b46189849192d2d4
zeeda7c60667a504c6c9befa9ac4fe6b5f2c45b48062ae0028e8456035120001d42ac566f8c23d3
z717aed1b6c61d884d14e80548347adf2fb758e6aae2edae6f91848faaa3fa1fe5feae16d1cac9b
zc0c6f9390bffc9ddd71edbedd0ad3eafcfbea4e687779b1a192fdf45df2be202d039c85ab4b11f
z8fe0a1b460916cc10ee51020d2c23deb04cc2e0fb43547c4bdeabb6aa318c7dadf5c3d7f14d555
z060ad758311e1c485a429056c596e8fe1888eab7be9337e113e3f8eff22b316ae48a6c6636353b
zcc16adfc2e88780a1e82aa454bc3baeb2906d083e6ad22593d38faa4598272e8c3e56fa7212000
z7704ccad4500f9f1f44a565823e004bf668b50f1921c60f14f9000170e38f728bf47d8491f42a7
z339633dd02cc07e42c004f81e5345ccd74e2954bfdf61fa9365113157bd5498ec6606e559850da
zad52934c265b1836efbd23a043d31486c8591e74c3511601ae560b12ed56142633d623c8633cca
z920af22b53b5c8d23d9a259c11074a5bcced66ee35a1e603fa67f76eff33f023b130aac869e833
z7261c02d6adfdb8727d1f76cd04f8f897045a48a2c579f65e66bd0f8b5757eb09e8aa3861c306e
z4531ef3907c6cf21af59cfec246cf76f58374c538a5eb194c2b27b32e46bc1ea2738a443a0bc91
zbce8e5072824c658907f3e8c6e5b56851d39629b6ffe4e74e3461d0d0dbe728d23720ba0f0544d
z9b8fc6737087c50cabbbf1754b2374042916d676d6ad98998092cb23ad29c9eb53f47f85fe9f9e
ze39afe0a06daa48fa3fada2e0ed3b1ed5c4cda428751a4eca23b0e97505e7a9909ffb5f0ba82ff
zd1529954f7c73f26b6b7e0b9e6d19ca97176fb339602a94289d4e068f2090eec919aa2453a7ce4
zcf90112efa7a6e782e5d6f98c0320e12b1d7c57f72c7add7eb9247666e46cc2b0297833e669955
zf7ea046443cb5250acf7c6b1cee585e85798fe36cb434c81225681794249602d513b4e46fb44d3
zea845e52e72b98b510f6ee0ee7525e580df725b4d3c7e0549896f330d581b8d100052012b3eb2c
z9a383d4a71bbc34b46ec39138995270592add8231752feb80574d027b4d2640a736444adf4dfeb
z09f0ba6152c2cb06334628aa7160ab285502b6551e551faa2789ace2bae2b2ae40e89d5a29b6c5
zd24f39faeaff0787f3f3e55565d7c876396983265b905606f903e1840ed65db30b8d85b0ba8b3e
z34bba9c3afbe84b98fd75abebc9fb9fd5e6d1ca1707314fdf7174ea47d4920e727c8b40aa0d28d
za235ec94a86f4e39d03e13c8124afcac4c4c4fe92e6788828e583ad81553b45292d0ef472ebff8
z05db529194bcdd1cc3c391eda50e0c4d3e55909aa2a9fdeaa9aeb68facdd48df2e470df400c0fd
zeea2328afb047a2812def670715cac1a4471a5139808b9c3939ebef796672b0b215f06b7f3ce95
zef055576816a1fca29e9e211c3dce0693fb88e444a03832c9700d1e4d813e4712dee4b9d07e2d1
zcc07fb3fb2682e48b43acd09e8392ca6d8c8b4508b5ccab5db0d3ce5af358d2f9c7b1b4eeaefa3
zef3d231d9dbbce6d52b757137cffd25e23d7db88303b7465a2b87954a6efa2ced0a9eaa748bec0
z88dc87e3ac7ea886b618c83e30555716dd588a625f8f9e390a2ca4d3d3e265c2959c0994dcac70
za756141c1ba3a2f43439cffe6d18134ad404c45b4ce211cda08248ac649d163095f8128628fab6
z35719500713d7a98401eac68fb6bc1936013c8960e2330c66e27d80260a999d47e78e70bb652a8
za9986f9b7c9c694a5bbb31728043c8f23a1e44ce13bb20103582952ba9cd1647d0556f0858b3c2
zf4dd353b24d9ef8f5523b8399ff636768f54c9d0b6bbcaa59905f33fb23b1f469ef221195e3068
z43f7baa3a53a3201be72df864715c76617a75695e9d459189b654a28d387a97bc03ff77469e5fe
z4652fa3dd92534e4a222c502cff5b2c69211ce29844360cad1f95da8499b7d417d807de5687c92
z511bdf9ab305cff6837d5fd7a8909ed4e690e161a47fc0f352e5dba2f67885bf7e292b2bb786be
z950ba535559e0e60061a1720a3e3a747a7b433b88e4a8207dbc86e231b32001602202c09267676
z98264bbc7a476eadd985812f4cb81b41496afe0edb12008ff000f25ffca86de6f4a95258136fd4
z72e4d06ce1a7bed14bcdd75a5570aadb35e5a5ebf30751177c23b3168fa87061698dc0be4ccf51
z5d64a39e5dc69c03222a97fcd9d5e72344895365da8cd636ea56f9f0ea5ac3942c7e256c2552b8
zb08cc8d0a6cc0e650b704cc2f03c3e20b296acdad22bcf90732131e38a75df44ae90b08d68caa9
z28365b143166bd21b8394586257d9406208b547a4a8ac22d6f87bb4e505338c8bb4aef69528be3
z2e16143baf4b65bf77024be92cd48446f05b860cf739a87eae7f2d53cef2811628412ad9589bb6
z03f3df62c7cf07c8ad9d7470b4922d6a2adf2d12e4eb32d91718d78a0a5ff2ee8a528a6b984956
z1fd577224ee35b333862e83f5348c760245912b248dc6a3a7efa2b7233c6044ce010cf6d8d16b9
zaf3332378d3800f3fdcfdaca3c227dd31532ed082fc260776614832c9232db4062734986f0b23a
zdf00fca1887caad762c5767fbdc083624b2c3a71d85755837f715d0022f9b8e383f43cf076b3a9
z6ee669b1de61cc597f20b2d71bf04cf0dca0da8b418b038334b0a94e9a2249c3411b66e3f1e816
z4e662d7c16e9c0103ebf4648cc7db0e83d63765ad458f5a19ff2b41b0d6819de2db1af0f3b8126
z80d966177fdbb1a686945d05da44da7f46146fc2b45b7cf98ab400120f644c8c4f22504576437d
ze38d62cdf9384a368ed4d8b8a1afd935bf0e0b87cb5e6270b1508effc7b9b080ba57ec369e2bf4
z1bcf2ec68db491afc83074914cf31081add6a0229f9bc255fa08323fa9dceb7b71be955017fa50
zccbe43ff9bd46536bec847b88f5cb0ce27f3fab13099bda8161ffd5d61290637e1012dacc1509e
z90f8eba5f0c2821db6e84c592e10b082b153a905bdcf73bc65f543472d477cc1a0f4ddb0ba1a94
z76d3eb1076393181bc9f29a20f5f28cf770e40454952926de7b38ed316652e32100b7532ea7117
z7ef6097f236a0c7fa155e43bb6486e8cc1cc4e7b325ed1e615afbdbc5cbd097df9fe0492b223d7
zf682cf09a3d00d10ee51560bf1dff858711b34f818f1f66813af22c06049161568f45678e4797b
z1c3b82f45663d7730dbcf084f1a8dc96ed53b2b04c752d8566089f2b5299a5bd2160f7e36d8cf0
z4c436abc33f1c7b1843178ca5aa73fdcc13976c5f01e855dc5d8f3762039da33324a3f935bafe0
z6e915c974596a63595959e295206af0d8d27e83936ea466667489ba1cfed32eb042dd83cdfe153
zf26c6486af08fc385508c5efd10cb5a7919731f1ed0bec0b7d3c457a3d45b6efa48d97a56759aa
z43aeff563a45fe0918afb7d2c16b6eb05f2083decb9efdbfc096f22f16bd0da495680122c622ec
z1a5a8fac1d95b78cd7cc757c5c6bc7a0218f82e27bb775099e3891f298114faaa2701aac1a2b02
zcba7430af57e5e5923b7e2f3603b3ca729b4204bda5814f3bb8717ae40130d143f0d1fe7d64915
z8d3d218c15f417b836aae49e2ab06091738d570125a06542bdfac29ec76c651d385119800f4b2b
zc592cb27ab49114f0131f48062c2823ba36668b8a60e8006de961185f68c9067e6a36f624293a3
z94a750e758a733826cc1a02ce1be4e774b2a163bbdf7cd6ba2317376acaaee8057923759f9c2ed
zf4ba7061801bcf3e652bd25dc3177f016ba27f369bbe3a619d1d21ed35b4a9f2da93b85b4f7437
zc517327fca52d5ad36daca982668da70debf7e2b70b2fe8f58293b3b8c2c13784c61dbd9bc118a
z36cb21a09cd88f720ad3c4a5334c4556cbfef3b1182b43119cb29b582f353c29e7dd0f9dbda0e9
z882434c72d935e3e1ef336e65feedb62350c0f6bd18d97613db92c8a5deefa656b53c0a270c54f
z996690f3ea38cdbb1acf9bd34584c20d4177f0fb8b28455e940018c17332b9c79131885bf698b2
zf1e09efaa17a74e57879d75dd58caf7c729f7d53d3c5dae06c173fb96f040cf142b073a07bac91
zdffb4747ef58e5fd0393686d70863bd4cd966b825cf054c37992b2b40e2244b6952dd1e047cff0
z91e756d7a5624bc6e820da6d4ac71e902dd60192ef60d546c6e4c183788245d6766e51c8f7c2c8
z9b59f83a44e01a58fb51145f6d0117c21278cb49bf53d65adcc00a9f2484616d5a6b917a55239d
z0a986e658578217ac363d5114baf94dd5ff542d4df10bc516d0ea12e866f2785380d8df18e89cb
z679c643525589628c0f7a12cd9fdf4072681c1468c0a6e39b07175a6647f65ab3e7c43d1f57055
zf511b1bc5304f9986c0a1f9702408ea87ea33067b9a42143b69ae2ea4da20aaf31a2e1912a9487
zd4e4133f4a82c15e5c8a05ba86647a08be48cc8be45d8a3fdcafe19d099b9101100706a6f5d4fa
ze54216ed640e9dac66f759ff3ea1fb1203d902e44d0c6ecd6a3a275a4c3c923fb240ed65ac1eb3
z757c64953e08219c9aaa5a7a0bd49ebc9d64e7008c589dcc4a85c2890263bd2b074f918e5e0c63
z114bcbe7f9b82cb534f698fd8b10a90b328474bc1d04bd9e7f96acb92844cc62d3fff7967cd599
z4ec09a6393c517a79ca2de377829ad450f280418e67f8c5789c673439d0b18bb0dff6d86a69852
z4032370b2c56b91ce915da9b06048bfcbd926d16b6d32fea6ff1f1a6b7116b2d594fba987f2922
zaa7310b11a109323059ce008f2c31e744e057fb931b3962715213c04db21323f9d5f5db1c15361
z42a37801eed5210b82ab2ea9b36e3a154ddefb641f8cdb16f0cef924d405373d2807fe92327f8c
z0344c063c32253e57065fdc8cabf8f77ac62a99aa8c9d08c1510b7021af4524050191f372682bb
z748a07891836b2f3d7714fa70a60d6a4092cb009a139985a4086d73e04668c0206b76282e1377e
z622e177edb8c5d03266cab0ed4d554bc1358c7580d6431f5338dab7e720459ace3f7f95267c0c7
z28559b6e0237829a86128e667eca2efd38b21b97befb66745061fe315485d477dcf30cd491a6c3
zd114b849c6d62b0c8b023393b0f8dd1e3dc7176fff14aae84d3b3fc6ebc9ecbe5e9d4e0b73ae38
z6ac11586580f5956e12a1d49a374881ea812e3050bebdf3b2bb77adee6f6415c6053185d4f9be0
zeaa43d34e30489a47f63210c250e76ee52f1118533e0be99f97bcb3bd8c9a93a6844eaf7f39dcb
zd2804a020c29c191c2ffc8e8c533c31a235a1bc12fbb9d771e3b16fc43a70095cc0ea1d000735e
zf78458bc136cd4a8bd7136e5281cf32ebf92ddbb7c70c38b9bd1be2813b6689748724529a2af03
z6176ddcf042430884b9281d03322226f316577e932493d4f083eaed1201a31cada59d79c116d02
z9dd619916b8276af258a269eb039487d939af41914542d48efd2d4601fde023258a77d0f0ea31b
zbc509c597aca17e97a6e40493ea0992b0865305a2b35eb4d38729b22d8fc845776b922978cccf9
z09285674c817732081a30fc9c012769411150aed1123565c6390c66afffa7aa14871692229b3da
z4404a6c98dcdc8b654af30dd75d0f8391b2b7b7da73091dca84de768a898df701c84450650e796
z03c3ce6e6e7345ae0a60f946e1f7919a4261057e00140294aba245a3bf93307209d09cc3030f8f
z8686a0430412275e2c070982aba8535dda243ac533c77bbf8e9e0982d7b8c1611d639c549c2019
zc56558e9facdba3c17840d924653f57ea3e660751e2b3578f34383a3f09a962a393878d6b1ddf2
zdae529a375a7118219041729d0b81047289978285a5b382e17574b6dcdb9c4c60ba8ae256de449
z4b581d79ebbb09cdb4170ba894b96b243b52c9c7e04d560a168404b75f944434bb2291d7ebc12c
z657dc61773104081fee2af0179ab7924c55bd2b7646ab6d6515e920147099d4ed3fac89f46df20
z3ffb4f51dc3bea145b36e243ef3340f74fbaac84e4fb9cfb598fd35214d0f55b8bb5b7b06db78f
z3c1eacc1e78da6b34e29127f2081c6a47e621781a1b97c2c8193b0512cd46b42bd6c8cf8007778
z8e21b756ed2b87e3674b4ce7f54c40e57ded768e9c20672917984c34e457b609deeaef1f2c1cbc
z9d37634bb44c588391ccaa261a1e397a3e859397b65b18068a308455974cadb29dcb9c291421a2
z03b9034ae93d8308a9fcd10e0dba4d40273d02709d298bc590467c687992c43f0bedeca1c32e91
z3186da838fa0fb0c8f410bcb1f55b48634fd6e8e1eb7562ca107d4eb484eb681cf4a9a51021c72
z31dbc4ff763599678fdcef8485488ea7fa7c0d0c75791aa5e9ef889591cd3b622ab8af45f844da
z7bef3c1b77ce7be933ef1d51c074675feb8f15bdb56b5627d89b86a64f47aeccf5839fccd9874b
zc86a248756f8855f12ab13bd47c8c41fa3d0cf87ce35cacab4f4a6bb1fe80d872690e4be482674
z370fa65d061981fa8a625120190a8daa6d05f1aa8810b45faf999ae852272dcab3ed3e6e8de2b4
z6351cd5d12c5daf854786a4ed2b5c90e7261af85fac21a7a775c1fef42da5968c5e557127b1180
z669aad4174d01b23165e4e44ffec90d7444752fe3a62d9e7c632f0e0dafce4aba680706ee38b4e
z6e32d2af99d71a78b4d67274346a8b6634b78bd0af62c7e243a018a666db2b8f69153a897c64e4
zac5c6134a44f49b804359cb3ab9b2508081d14bef2f21674e5f31cb4e14d17e12a120c486f9977
z2ac0ddf314490c6921435e4fe040d433dd2e0cc11998ef284a21ab961ea1e8895c8d741c63ab5d
z1a185ed8780c1ec452d461bec312721d3865aedf19e614b270ad313609e08dcfaa6a21c774c1ca
z7b7b65eab58121d14765c85ec6dac3a754bd4e5994addf8694b19ecbb07228d99c2a322dbe380b
zca6e403db408b00d21b0ee42db56b632a1ed36ad179da765e52a34f02e8ad8a3e1e85af654c82d
z5890c29819c05faf41dfaf990e6f39c42df59c62699b2e2ac9422f96aef64a805096dfedb00a2e
zdd4da31f9d0d2506d2f3c3644eac4922044d86f5ae2ff1c1e6e089767ef118d602f9d1c5af0115
z6a6f9db804c7c75f3c4f8517c64025025995becc377ec47cafa18ecb1bbf33f1ff3aca3942f905
z14a000383732b31444719a369cb194e3930630fcc06cc99f0ee7b7d27868d7cccfc5cf395d7e14
z1bb653512a622d155900f7d3a85fae3eedbf331c91551f0bf1c93998c5ea9e4d3c745befd97d41
z0ce639994aec7266e3315816237f7e8fdf9987829de8d91c5257adc44c7c8442bdafeec2d2f9b4
za000127d46649598d671681a1aa8cd1c02a6eb602eda454474453a5d430edc2123e501beaaacba
z7941a154196b67f06a346d880137fd51db0b31ffda3d10349c11f6143e2477862829ecd47eb9fa
z9d4c5c2822a4cd85bfa009004f16f529fc79207bb3d8821b8bbd56d6c26ed61d4150005994760f
z8617edc9b6057850a15d194e2c61536d655a4f52bd40e9327a396ecd38f5a39fdc2f921640fbe4
z19051c73322e678441e72b399f9329afeb90f3b52b4cd4ba55ddfd49865a13eeaf57373105193c
zd32f8ea971bc1cc9d59493565e37a2703d8ef0b56b5363e896025170ccec9e0dd292f6cdd13979
zfad80457dcec88e9503dec3cb8791ababaf6731b8d31867c97bd4d26735622205c4e277af53dfe
zd348f249e496a5ae6f2b99f484f70f55404bb6920e6e0c415f0a288a198daa1fa58a7ab668bb45
z8a05e825dddbaadef7dc39d94b74f9e64e6a091b3078eb4e83b8e541495577033e03628eb86576
zccb5157b7fa9162f2ebda2aaefa73b5ac1c41bc94b96cab2efbc93ac4fb2104b2ba08029fcea20
zed03e262522fbe6d5965afec2361d2c4e946c2d20d84018b5a5ba844b3fe73ae1ba12120d27dd2
zbf02859df5bb2c5f53fb0116769e111ffb8534dce23b49099581f6c437c303fe5451fd09ea3459
z3d61262c76f1981a92d5182e0110fd1b741a1d8990b7ed82d5455eccd8085448ca22d015c45121
zdd3603a68b53262c3dbe6a98afd332ceb43019d91899464c6404e5451d887069f85891707830c7
z974003b90dad9d3d518e2ecd140524ef53e11fc39d3a6c6c6b71443432dcca36571694ce6ffff0
z30d9d3a4af68c315bb65dffdb6e4cfd2b581b3a4bd0e9ff9faae2d6612f5636485e69892554926
zd65fc0b874e9df9a270bb7de47e2fea689f3c2488299f44dcf0dc378243ac241e5e6a89745a6db
z8784af3db783dc6390937dbf4d9f71d1f3975259e29c47af60ddf8465d681e61381cd8ed6ca289
z023407eeaceb41fc887aa2e8dde2511545b939c4a3bc97f93ca8933ce2852bb6bd9ea54e032a0b
z8b695c89a7b3b07cc0bb87e0a0d3b92b4af2fe63e3f970f717475d085b72f1000dbade3f700c5e
z85eef4b3765ae87b91b8bd3d98413beb45a5ab43c2ee8991bef17e81e7f8fffe39f7f927715265
zd41dee4aec909d1d0289a778577587272b95711e5de9e66a49f7c57593bb0fa17a232cacc25e96
z0bceab00af05df10153ae0a18bfa6644068eaa678b7cbe84792b050ab57466616267f4b30d8412
zb62a304948f5715e6f064533bd5dc7a1c562c72aef7bd627f6cc6efb728b67d719d502e5095b63
zd4356f0c11a0d2dbc1d8a7f83a335c49081eeea0875b60c4da0addabcac9a847caf8eda249bbad
z3628b8dd337bec67ea1b7c13eb80cb1db1b135afe77de71d658bfc8213602bbd0241aa79c0b782
zf6c11e111a59ccc4935452ac3c962bd8da4f4bc7a275667b7d2f653b5495598beaea7545782795
z1e9dd4c437de58d4c78039007f04bbde1f0e6c26568874d3e8a493d55939e0d31c1f93da569190
zb72aa2846b4293c6f6414b49fa18258fc6105403929baaa2650b2f08c478c9bb02bc30e24ef091
z01857e638c301129d24fefea848bdd2ce07ecafc9e9a47b7d4f74973176463d01b7872dd5a6fb1
z9988de098f9ab1a86a856c727940af4fd63cc803ae08427531b64ad91b2321f118f14d8c28a9f6
z10b22cc7e48fc737ef5c25902eca7fcc0713a8c99290ac04131556decb5150bdd04b0b31a6df01
z8dd3c111942628465b1fceab2610878f2337d688d04c7dad80f1eb93e54dbd76b6f8f893baede5
z457af0a9231138b9f3dfb920f880ed51c47dba540f90afb182028de1562d07c7ccdeddf0648b88
z5a3c2ecb1c9b4cb6c332288fbdd94489d925c146977e66df80038911690900b7128eded6b03776
z3be9a9467b7eeb16cddd4075c306a7a6dc8dc73fec8c2156d9fe85e931dd64677a828439220934
z91784c3f81ea2ef8decfa125c1c36db056d8a814d9bcfcff7a9826c675cba03c14740f655dbca3
z00408cb29051517151c1d9b1888dae4e4c1f3bbace0be725084807db528a433bfb8676b5b22746
z1dd5206a704410de1e36785d2b34f2fb7947f64efeabc6e5a4ce9e8bf61a217f3c5d5b90e91ed8
z6639989dea35797cb3f4d2a87282967deccb08ae8d8ccc12494632efe4741e4952c818df28f1e4
z6a49c8f2e0cf893843d435fd0c5937cd9a779bbbc4bb06b7026141a33a3d8e2defdc8aff587186
zd83eae374a781c5948eba8057b7fdf96b2e8c5589e93d51f0e2ef1111da42adff0b791c612cd38
z1f2d94028f48f877843cc7f6df85d6bbe951888e0d1f5caca8ef933b8eb36a35fe2172c4bac92f
zeb6385c131097145f00863ffb8ae6cc8b7209447c67cb37e44fc7dc6c17303feee45f44ad6d963
z3ef8a22441284d061d60c662deab3759a4a57a9adf1014311746821b75692f9a4e6b399e821219
z34e733de198c9c9ab705ed801ca456abbfb2a54c2a66f2e3e164cc19d806090710538774501ae3
ze3b97d2411692f9e52bcaf3f82fe036f4d8da1582bef3fe635c2f4ae8c775174dcccbc53424d83
z614a07ddd1e425ae38d90ab859ea5c2ea713eff011f826c33f98bbc3363751290e544f07e045cb
z0bdcaec2b6c4dc2841939594e75665b3492955387e7d7d3aec81f6ddaca93cbbebdb22cb96cb9b
z5472f3b87f7bada0fb52b625ab1c3de11f8cd44bff30c46e68b1ccc9fd675f24277442d9bff5b2
z71b976458f1d3ee5957fd00a53b556f5bb0459d6cd35b361be1e30bb496f45f9e2082d6cfe11f4
z8b86301e3e4ec1ad21a63ebf289bf1d97efd00ab722df729174ee269d701171e159c65be360724
z5ab1e05a8f2d77e0768836ec7221599af68de603f2f2d01caa18c4dc120f526866145019c592f0
zcea010322afaa83ea2dc399522d2e0fd9fa940f0b77b5e5208edfe00d0444f84708eabecf1fc62
z110aae5b5ecada0886efdb8607aece338a08308bb35c7ee35ab8130ec1d4cd5af07a4af504dbcc
z8f61953c95a7535624b3a5a105ad11141d9a02d79b24a822977023a5836094aa4bafb8a016eac5
z19f5203c0269a945796917a5a49a7f1e059353e2d72d6822fc8985fb6d10554383d9b491e56dec
z486d61c9a8579666726a915a40a73b29f3d50bbe8d47bdb09b5922afec9557fd30c9668b636d50
z5559bb958e9671482a504660e18100706a21fb07eb64074d0cde8a1ddc849ea9cf939d3a017f9f
ze8758367927ea1bd04593dc472e6ef415ae87eba561651bbc158fbbc2e430f5982102847550969
z821a2a89769da9bf644a62f12ac12d77610064d4fc50407b3a28f7a9308f1d6604c506868e5b73
zf03cf7101e0d18fd4a8341180f0cdbe4e241324091ee5e1b1982e73538faf47618f9a34773e58d
zf59b599bbeea873f52c28637bb0c6edda9501e5a0a6b0cb3876fc5edc396088618ef1de5af5365
z6987767acb8d8848662b30f32ab36b8d380a175683fef55f511c5320bbca63dab53caa31a28ff7
zfc58a3246aeb9c89dbabbfea29a9fca54ce8b3a4aa097ee52772ecd17799eb694cda37e1875f70
zd8b6060854647455d16f39b6e388761886a744ec9655596e3d3dbc8907f28d7ab2d63a503db82c
z76342dfe236fde80d1420997774f1a989c2061ac5c95779bdff5a713c2dfb0a8edfc33c7dce4d1
z5c74739a3c297239add3c624982eca5da8689e6f55ce0b4fb2e3ad0b62ea245d77ec703e84aa83
z5d4a6d4605fc7ec016ddd612dabe21ffdd4e8f35d99bf5869686fdf60c746d7239616d14d02dee
z1bfc90896edfc9690626bcd760d8a24eca24c23565a411f8894d5466ba0b933f508860b98af50d
z105e7bce910f25b1030963f8d9a824707d085c99b3ef262f024c9ae01932f21053efcd3b629232
z6e342bd7bfcfad29a26ef00493070936ef7a4c5377f0261e8f3dfdd5bdc29a5f20e74fe9a434d2
z4ec72d8c31465049ef932e3e7b0f0e09d3695fc831d01787286d837f315285e4628c024f427815
z65dbcf774f8a13e089da42008f9c8f3b434cd2dcf086207c32d18d96275609b8b8f81361d4bad6
z748f0da1c9f0ab4ea1370e551919f6dead4fca34052bfc35c6abd16948379e5a12b3a6705263d0
zefe58651441d36c6252a5d9856d738db8d20aae0ee5434160b81c66c34b0ed49abba819186fd99
z6fcdc1c09f42bfdddb9fd89dc48b62d977786292bf699491156fccc68c0b67458bc2bb626b7a14
z754370ed3ace9ecc8eb1325126ffbfb8bafbb51efc4ee026392ed43d1ac4c3b7823f2956bdee1c
zf1b081cd4a659fa618e189cc4da269a032268916208eeab915ef9e6a6620f92c62aa113f2cd81d
z3c258f9bbceabb1fe1032f22d5b5a65fd2791cc7775dfa578eef3701c685ac370a1e7401214415
zb6f39721daecf0c0d4538b0acd1396d06092d6dcd9dd7f02e1e887f04be03fd3716151aa3a0d7c
z2a773098e1b9353c0520a2ad6684bb815944f546fe25b614a2dee28ca60e96f171a55fd2f904ed
z31e3f4b998eb84788fd5349331b22870769c7e74bd8a05feae3bccbb1b04eacde1c3efb6a9e929
z42ce207636a14c4b691c4643b82057b0a6f9813f5ceb70dc54ecfcb54f17e265972d982a922bdf
z41fd1237dab63912aae653d3941186beb1e9de3a4cecf29f4b1e4ac4b461b2a7039d6817158944
z44b1ef7df2e216a4528d2e5f9be0771ef755dec51f546a1313904b36566986bde8b583bf8377c2
z55f9f1cdb6fdfd3b4f9bdcc370a4f25cea9ff17b6ce5cf70664f1e59b275171925a4a9314e1f2f
ze5cc317f024fa606a4e79fabc70d3b4a3225c1590489834d81ce866255002d3720c7386b558410
za1ebfb2718984e383793dbc8e54e47b4faa3bbc617fca9d168b902d66faff89f67308f396a9945
z352d4a0a814086f590cdfa71d3539060e1af3a2c93551f8b4398e88ed9e799a85228a30e05b9d2
ze316dc597c30671f365f9994cc0d49e3ae8671121b7f6a53510b89b2ee12c183aa2e2cc73b07e6
zb1db25acf032ecdbe8e00da3a7d1f0e9f1e9b81bacb2d8804ba54f073bca60caa0191899c7b147
z0ef9ec3db7181e389e40d539e523bab6dd1914981df335a1ecb1e9e26ca7ae4face6703f944337
z492855f3ac4f3cf2be82e166812edeec89dbfdcb8cb11de6e205ea59f98590710ca15239b108ef
z2ee99c978e36ef1a7115480c3340abff50cbc9a54b88dd87841165dec51e59dc77a69e82e73af7
z7db9e7605078a89ce4af2af0d12f36c36d7f4531ddc61c41e0e485053ee5f328c0699de50ea28d
zd39b75b2d6f7145af742ed0a2a2cdc3e392800a1f349aa0404f6fd01b4a18e4185264507c0473e
z68765be8f05b0c00336a8f299c0a55ca42c07b8072395dc13bc92060d75efcf83865c6a54e6b5e
zeb2c072d79af2632d56f4e78d152687a0488dfe5ec3f1f1413618dcdb1f0924d8e8ea53a06a7fb
z4142278ca844774bb5c5478d07bb67009f7b6e5ea0973cefb5d5cfbd3a4d186aafa2afc32ed028
zf9b0bc3441ae1f1fb6e3c72efabeb9ec7b3d017519f04358fc08f251a023ce5ce43cb6bf25ffbe
zd0d256eb730dfa0bb3a37fd7e2fd392b40c7ef22df9c129baef58be08c99eea0a390824ac2816c
zb510857fc898cde30245f26533df870fd8a316e7bb1a2d5ea9cd36d09ca9d433d527069fc10cad
z3a86934b8588c1c1db95453e511682c0ab977619e415c8821477ed355eb37e6d4f72a25b006190
z9cf0d35bedfceb49ef0dc7dedc13eefd0c2090dd9a543fa901b7c18ce0eb3883b10e658c6c4759
zef86c025150eb9eb4f5a635700f3c53ed1790082cb8af7eda864e0bdafe0801029fc92bf22cc5f
zee7a319015e87be6f4e4c496d798d51ab170469b6176776b336af90b654009a10dcdd8e6dd883e
zb7f76a6f5560812643b6b498ab7cfdc04f73fdc7048447d47b154be81fda6d5dabdaadd4436784
z14e9e699df4dd814e46233f90f501bd6b797e280df3d3a4e65abd2ff5dd72e4080fb1958baeb75
zcff8dc2d8fd3bacf85ca2ce95ae8e453969f2ac858c5b3a510d97347b1d812ea45db97024b7fd2
z40c9e88ff6516d6d1c099b29a7784f2717d3c4087537d26e5b84a8bd4d597087649b6ac5133177
zb938ee20fd2e11975b4365261fefb877db9f3bef99d21f39bdf2680aa8bd6e9a912f4bb1a2658c
zee430f13b472f422fdb514f56968b918f3b76cb167ad49a8cd3d24f4f38ed51d5b1bdcb5ddacc0
z23a9f0d968dac732d1e6580c563ecdfd07dc4e2be80e2b1572a430e779037c309d407d725dd933
z0c609b954f2bb8497e5f1515dbc3fdcf1079572404b62351cde913a1419b927517a822e8b37176
z9c9375adba8ed3fc31552c9fa8cdad41666248f8669e113c0a2389fcf163e13e9c6bbe280502d7
zaaf39e9cc3d62e8be78cb6d619ff4575a3c968261242a7d83d309febda6385959ccff7be44b33b
z56fd3fdc0e5bb0180652b86cd035fd4a1f14c382d12f7e30cd0415fbbcbb48a533648d4f7b7611
z2850d2aaf887f882b47f79a7b3ad34c04b2487c9a34f7bf538260e1ed9f1ac20bda05ef45e906d
zb3a96bfb64f718b5ecc8a15739eb90deee71bd259980c9430af4aac52f36685b0281c86b8c0a6f
z8dd7836d7dcd6cd45fa29cdaaaaa1ceb6a532ec716afbb90dcb82e57070771650675553b38909e
z80cf303ada641cf7eff27393b1c88f5665f60c1f0f1a380f60494462b2da7def8cb8a207395ba6
ze8fac9a0e7e4896a6822dec4726cfc5ef111503fc7476383adfa5d309ea77d422d96eeb72b61b8
zf2fcaa500413039beaaf8c56dca9bf93daed89677184502aadd262db3da8594e3ac8d2ba82bdb4
zaed4c3755d6dd696fb955e88c153f81f924e0fa1578acbb97ac13b8b8256625ddf3f1417952906
z72b3f72c1d8cf0bc4f1b0f1c09e252bf74cd4656bc7e630b96963ef70f2771749eadeed2eae154
z3ab6a144c6901a6520bafee05661bd34ee5ee370d8a5eec520efe168aadee9da9c90da9c1078d1
za4d2a31322524240f44c07a0b6edd818031204ded01bea102b7c33b4e808f40266818c081da961
z1b7b260eef482c409e9054a78e094708efd0def775bd2c0c493c3cdc41c136d6c4cf505240a711
z324c538e4dbc3ba3961a9d0002f5960c0ed4c3ae4033395478ffac7f2ba30892975b85c118e253
za11ae9bd5f068cbab7eb7acc91dcaff6918a29b0b470c9fb36f32e3093e72604818a2366ec3183
z91def19cf941eb32269a6d3bdc040a72352cdea47f034349c2a468c590b500c08f1e0d4df8f94f
zae16346e9b952910906fc774396e16ad17c72f9777f80dd3e3f32a0198dd0435c502104dd21a60
zae7aea0d1ade0d7c95898624ddc60ba236c0677935369b807e47880190344ecdb120b018312022
z5fe0bc3efb94815bb10708def7f8e73ad6b9c6a45e63d403a7ac3cde6961b7b709a9616845931c
z62e3e5232eab70e70bc1b72d84b5b0f95a33bfc19af8d860b7395882d000767453ea6b4d4c6ef4
z72f8c1c5cf1776da1b6f1d028f3df3c9061147bbbfb62d1f32c9c3b2de4c31b2b7820fa290e20c
z787c71b4e78db2a069fd2100b6d2b96850b264cbfde108041c07ec802b847d67eff0ce2d1347f8
zc8c1728768959eb949b727928f3c4ecbbcccf1e43166a7c8853920580d69d888b43f17b8780ff5
zab4cafe920f50b1dae68b3c73a26aa95407b2e4f4e66fbad0655e846a56d5323082809b88a3374
z96177b802feb6d68e4a3804d1219796401bb9a95d285ba6f299d40d92cec1e973ee96628c4ea20
z44a72eda5f3385718ba01a8b5b434021087b4a54e6f90d630a9babab473e792ff410fed290b66e
z5bd2371863d419d1e21a9a977c91fdc889319de70f67df2a5250136f69420bc0f37152cc6b0fc0
z8ded0799cbd994a871eb444f59692b3313a0771851ff16e87a602d81cd20aedd26357b47a0ba55
z6ec8e519f13947b686de1af46376d05542a714bd4004a925cc94ab529f8c3f87b29b3a919a7d8c
z8676897ad4af44b50ad0e5db6abd2bf089d922f1c350af70be000f85af743b4d2af562a0de2e90
z15d331cd4e44d0956ccc2298bbd99482361dc231d4c4328a2a81915ce629f71765de471d2f7cde
z66b0c43f50a0c38af042fd0dded20cf91b46d5110b7d1a7d8f652791e33e0301ebe4745f6f34cd
z5da2b796289369c6cbf0545e833a50f0461ead7ef956e69a24824cd85d2afd52ce21ed8c3a7480
z364b451028cfb621ff1085e58f9872caa6990fa671f19eeda76ebbce0e0f94786836e2acc9aea9
zee04a8d8c1f2c72890fc5c03c4199e6fe68d3d340bf6890218b1e5440779bd02f90bf77d634212
z80af4df514e6efeb3922755be7ec43d91290ddefe7800975510bf13760b9d4e26ff73d3982b7c8
z664a32c4b15403e9775a5c572d7eb3059eb79c05134dddca52ba611a94ed7e6e19a4ca59c73160
ze79a8512667d069c1e2f1efb04f0caee0455bbd480a6e6c5d1a8e7e438adaa41db0d9234940f0e
z2b8635b73b18dd1e987431519300f2b59ff1fb75bf91fbfd024adf6b0b1f33c347b78d953424df
z3ab1dcc3a9f96a1c0d4d377b25a7d4725c9c095eff958879676da5829bdc39051cd7b182a20545
z6b72d2670cd2157f154a5b7402b1bd68fbbd7c174ae501d5262073de363fed5077dbad95870e5f
zd566dc058474cdd6cf9a5b05d2ea0db70465a6f690e3b7f140255c22d28ad060b05b5d607299e1
z75373bcc98009a2cf62334e1964d306b98a3298ed673a1d1a0409d70fec181956bfa559fcc7462
z6dc9e1e73e403a2baa3e6bcfdff01ed1382181fd5521753414fb43653359fa5353fd1d8babb08f
ze029ad124618c316bbee6d855dc0285da5a81021e6a2df157874e7992c823efe1ce01bfaf166a6
z118fd81a00ad3bc55143b5a8137299946de41fd71956b1f726b918bc14dec8c6b9ff9127493d33
z61f85a3482c231b32cb0c67d8a0ce5e61d80aaf98c92986bf6d3b8370f496f8113318add4e986d
za8d7df70b033b7ca92496055a98af6cab678cee844e146dff8b01ba2ee34320e235fd4e031ee42
zb65bfba588be172a2906b6fa6a9ab8a896e0a2b1405ca413e50cc1f5d88f028d193c9b409ff4fa
zbf871ecffe66ed91001d622f7422079f31b6f61b3afe9a04acf0487d13b93df38c9fae1179d4b2
zaa2a1f3d61854b1240fbd77b794f6a4fca60aa512aa17cd88ce71a25f49e6567ff2a931c0b9498
z99d0224bc0639d52acfbfa2d340fd5228be6a953793f0357475a5b27b5869eb838ecb42f67329b
zeba8820038724a65db847c596caa571de0795dc4e6503c0af65f4697578b8cb3297102704cf492
z864ad04cccbc99cae20cd9a17f809c62b0f0a16d4002ebb1a782a946cdde0e9d6ede9005e2def5
z484fa700f34d71df1858856981934ff7a1da6e9ce7bd81a50e721d779d0a8e72a49b925578d139
z9bf577de5fb6da36f50e60bcc9eb568d5be3df16ec210a4ae95e25967ee3a363e6ba1c387c9fcd
zcf18acd6a31bdfcd50188b45837e33728e497b56035f2d57a1598811ae94929ddac517f6acbf40
z2ccdbf9f0beaa51caa5ca9cf60d823d1b1fd870945ec43fc1069185f0f36a24fc33d4a3bee0655
z2eaf9362158ad9b6386f64bcd292e40dac48278177e6049d9719e5e4c111e61391f9db08d123e3
zdac4b2f50a514c08efab76ea7683a92327983f4eda7dd0d0b751ed0aa775b2a32f28553198df1a
zc966e21b48e675820e14bd0984c82a8fa9fe47c03f83123b2d5079d492edc9be12cbfd2cd8fd10
zfbe5fd32dc5ba9539cf7b290b4c1ff19b2022232c8ff96bbcc04ff35389a3d9884d62004955e4b
z57967a7d3d11d3389504fa27a73991f45603154409123665b4e74d3352997cd051e4f1ef7a2379
zd97dd5761eb1e17c6c419fbc05a127957c19fbfc94057a47b22148ccc62c8020f22af7957545fd
zabd349f7c6ad14da12005719d2600e5c2e3880effb84ea547979964cdb30a07563ab9957de802d
za3fa4c6141801b260d823f141229d5bba9bedcfb5fa23f2cdfa35dd6a29b219714a6c67e64eed7
zd8d05513b2dc4860f89393e157a596313acf51d2c76e699d706acd18efd6645d800a72e6230399
zf106e6c05e0219f219f287d1896adbc868a3e42617dc516085d030e3665c3b1838aeb046e200a2
z818b7922680865a9934d57cca1a5fa045c0f897dfbb3baa75fb89ea5b87203b89fafdc90ba4600
zd7dc787c8134b0c32c519b9d904c3b6304f09dcd399c869c518ba36a8f89e8f2e40b30dbb7b494
zc8df0be0dbea809a56c023be0a896d11b9583d27cbb5efe6bf8ad0a3e612c186c9374c61378a7a
z5cc8e2392a30046726cb2f6687f7b9d7662ebcd17cd2be1e4783dfb051b6ccf9e961008f62b231
z1f00cea95b8a1de5caf14d41461de990bd73a8c581d33265325a8fbc459d857fdc5857d8364023
z9b09d3e8e3cd74e5eb217e88ded3c0b00df655625221bb61807fbc7c452a2c20add07134bcb0fd
z21fa19a15417485dac58a349775ef657aff47391d3f2fd553c8e308e07b8310658f2a5e710a793
zd0b570b9cca26e67d73d22ea3601a9d6374fcd8dda4aed063ee59fadb1f0552e8386647db05809
zda242c944a300fa668bf5783d4013f65feb3e3dbdafd27175d02a0c56d6cc336892dd60954f042
z89836bc2f1b677d06b8ae8e67c2ea6ef7e4cb53c41a7197f7a6deccfa549c4e05515e6f5ba7edb
z380308785ddf6abf9a640ac74769bca4105431cf97d6d7d7650603ab8bfd3f4cab2a7ef738110c
z129d926110565ed82babefd97b00018933bf101482c14ff53d1e369114c4f60e7e96b20fdb28b8
z7e97962d70cbd6fe4d291840e10501294855c2842502aa9ccb4135eaa5776bb99266cf3208d631
za644eeaa883a6f79021e44e56d9ea76837d780a7e6688a9bbe2946a0eb899fd4804a48bd44b016
zc836677df39bc9981b843748b92aa0bbf7ffa80075cce1151f1f7ade300fa8105823a46ae81b4b
zf520af550f06d1b35f27caba4f9390d476c77a54573dc6dbad01d22882708263eb17eae440ebe3
ze718fd02ed9189d1fd1beb03e5ddd8fabc492d6b2271dc702d292b001a30d5e5dc58c8fdcb44f6
z1236b8382291504ac38c6aa927fcd2be2ea4b29ffde765b709c45c00ba11d01a46093e7769d7ea
zfd2202b80d451debc9b97efcf25ef4aaf9b3d6ea5b98fd19570482fcde8495ea4854ae80c28043
z91cb4dbc4a3d541c011d05ca1376c146aef140341e05c2dd769481a4283280577b199af2a85b90
z5c51c4e2d330132def6487a68063babcfa15b12c395148f39d481be841c520deb96de3d3a55f2f
z5b7efc01c4ae1a529fade9abe0f6369d3bf79558236deedf2ffb2af903a0e8b8b66debe7dff532
z8f9a54796ca905e87c36339853d72004b120ae927e3254ee77056b99f369cc8b1475bb550d7b77
z14f1e389ccf53c5fe54480ad351422a78f6a4544f9dd99e1ef55b3694d5f6b99b54c63b71382d6
z5a4a69aa310643bc39d4a6a1d7723440165dbe203fe8367b4189828dfc532f9343965db003bc53
zad2f8155928917a327b8ec5986851de901fc855ad1731a721bcbf4c1f6da5e886c76aff1c96a93
zf59e244774ac706ccd61902c4f326416f2625dc15abfc1393b8aa17d397ecd41c57a3f1fac7447
z090efaad842b9ebc58ff4abe97327fd9e074e3440eebf18cb5e497a1d7665e832298ac7a9ebe89
z1fa6b2cd14adca3fa1af912bcc1c327ffa0c487b171e093b7d56f08abeadd2b67d099d05b34b27
za63851e98b802cdd265095bf69edb37cd6cfdf3fc8ea54498b09cde487ce4f61cbe158abbc2da9
zd0007bdc213cbcdfa91ba216d3445016ce9258404085cac9b390d5e5e8282bf9ef9ff351110fb9
z496a74104e3f896ef407d059ca45d55acab6e965d658814a2991a3b54d1a4f618cdb419a1746c9
z1357a0cba850832a52e4dd27de351f8ae965f5c6c45e841d10f2f1244a3d4ed31bbca93f121772
zf0d82dcb491fafb4e96321d27398de24dc24252b742dc94503086715b1fdd1bae8785d3d2bb8c4
zbfe6ee443553e42123e16e0a5f3bc91b87c4113368ab2bdd3cb34814d0a9e52f9547607ad57f98
zf003491bc845abfabaa804885ce3f95a07063fe3de667fa4e5cec490ef5c74ad057cad513f03ff
z178d22cc3cc7987f18d25968966253beaac20e636a714ec7d9067d7393ccb4fa3e3640dc1a5173
zbd5444f86587c89c56a7bf3cf10a48dcf327cc472eb7516b414570d7de33fe7e977586e071101c
zce955623f1e0d407388114a47a84d9e6dea4741a1ff2af9be614ffcdba63931b51ecdf8e3438e3
zff0136744238525141f83edb46d3cc698158e29f0f29cb1524cc8a20ec5c4f78d713e1ad4f2d38
z5382f8918af2e735b4d43a7581ed1e80a21529b622bf448ae891d2bb4218a690195dd1a8f53888
zfd683a9b8386d827b18788340bb779d7293ffd0fe5c3ea868d31020ec6523ebda58ba914094e1c
z03d80eeb0a1ca54621c8b5dd85b39b0dcb130cdaf6f24ee2c8c08cbefb6260b2c0b63cb9662a2b
z56da60fff950f47fd72ec43e50bc57ecdb90ad205752e99d31a614cece9e2f767f2114138e3cf0
z3abbbf21e6047e9c3df0c21311cf9d39e7743457be6bda7a2aba8a00c7b6cb1d82a5fe8e2dae34
z66d9c00b25da11be369075fc848b48bd4b2e63c02e4be5bce908a11f46a231ef27051353990a0e
zec4dfdd549f4adbc492402368c556168e41ae3ef7f41f0eb05b300e94ae0e554470192dfda81ce
z01ff7f2e2481090e82517cbe1f18365dd218a0e2f844dcb12c115a80248ab8a840522cef72b681
z61d3cb2e6e1c8c7932f3a8764debd4676dd8d2ec749a0a3e215345c4ebb6a489cdbd1ad625d0d4
zd6cbe6bb5f35dd05ccbfe44fb2ab34b0650e703ff9f3b0f3c371634d1f2b4ea5f2863c986372d0
z799ec9a73742e7f258625bf50db37c725b5a3ba1d97291f288cc49beaae376bf6402c8deebf758
zd3089d7d7a4d2965632cb2d35c57f3eec84d542f152620a774e8425ee9633ce6eade7b9b9b5f03
z5f3f8c1b8de31fbd4adc734a4ee415554e1e16d4df45068bb956e98d0befb2530df11a1772faa3
z9c17c9cc8c43973ec9629877c8048c0356d46bfc5b1a799b4f1951b02605515bf8117df6709f97
z86399c02ac47e5a979c43680a9d503c1af049a4faba4e1a8a744ddfa4a33dab28bc189a42a55b8
zbbf737f6a4ad72a47528e9ac72652844c73cab93e84080980f3100a0b4c4a165f3be1eaed3c37f
z7554b733e604466d5751c476775d65911e2030212806946b9e0a2490ed22c591345ceceeb56bd9
z3cb4cfb522de781259f53507d73b9615552e311fdb796cce7687ff383ae6aeb373a8c750f1b5c1
z80786a847126f537ddd8a211831bc713c2358ccefa83e67fd9917df4ffc25f69c8f86652b0e23b
z0a551c675e172474d5818a872013451c7e984d090f4a8bc7036630671994c86c5f04f82ba3f929
zd547d13dd657681fe75d521293fb6e0dd61f4f7443c1236025cb75941da4aa776cd1c1448762ee
zb5ed5d236fd19b884ee50bb0b225691c20ebc95bfdd14574d9624fd87a335c4eda72891852c9a5
zdfac6ebb1a580da3081c4e8f4894a1a06e31cac5d0bbc7a404f8db19b356cc70287624732723c2
z9df85a4110c6a74e7a4f310c8aaf0542bfa6132e5e805cb95016b4040e73b60a626136fea353c2
z2ca223c6d80ff993297bbb8b29c192bf20918be7e705139c135e3e04f3b28c2f07dea28c3bbc04
z37cfdfd23d1d76c2b32ee803422d987d3ca04193d55a34e8bc2c964519a4c8e595d93d64964d6c
z862bf2c0ff48083f43344797a4560d426e5f5bbe1c951ed0b64c15d80c70e20a29b56d288da456
za0ee909173a0dd9b94891a782cf5f94c8762a806a1fdac9aac86cb47837f867056ce1c9717130d
zbc475afc695f83fe910aa40bbe4ee36bdca301760df472be6ca53c1968134b3a88acfd11efd129
zf3cd07f612e1acecb4f5d73d7b8551902929dd38f3057399c39dc470411dee8d4a0379e320ab98
ze75c35932882f18a1302bee1e12bce7d623a20aec802338e35422b4ec988af782e4efb111d392b
zd3fcd84c1b57fb9248a11befd96065c2ccfc02c5485e781d6beb4711f085f28819642180ff5dfd
z301e21b705554c71c405b464c704097bbb297504f8144ffdf0a4ea1828d934355949b839564399
z12fa3b6a1aee881a9c7a0da54a4f4a0e8f9534aa6ccb89275e8b2c5555c55aaefe418be27feb9b
z104f23ce341aef951559fd67b6bf7af24fb935e5b4df9f5f82b313c0ef957b382a570653389889
zcb2287e715b307d93f283e48f7d031f39f0957447180dae2a9449a81a6bef372000dbb2bbafc05
ze19af18c59e036902644fade7911f77c201f919c16d450afd10fe9e569b1f528c00d73bedd0c15
z07a7c4efb2cceb2c93e47980f6ceff3df1590985d5c8ca7f232d886d9dfdb1f26feff148d3fc44
z7edaf97bd6f72d3c6657816457fd7d5ea4cbe830dd36ae215071d72ee42439bcca26322ab126dc
z4e38dbebc34339f5aa60986dd0bdf55f5dcffa9961551929b0a5a29828f3dc6bf318e8980c7d82
z4d494ad3a81c57e8ad8d889a6a85b0f176f0fc30f0cfb9fe4d83d8c90ccec01daf338eadd7fdfc
z3dd8c7c2272f92b6769e4e9af589694d964b0e8a6dd97b26522cdb666c02bc02e2efb11773e9be
z10f7bd80094e9c0109ec0f3e2f6ff38be6e571820920acf4335244af72b10d19d627070041699f
z9eef2537b717069b583253ff62c7fcabaae070c4c2e5566c8f808aded32c6981aeea0777c1e5cb
zae4859a196610f825c0d6c86ec1d355142e32638674165d32936e9e4636d71fcec163f17c197cc
zb4bb60f0778db490b0a4b1769696c9b7f57807ad1d62754047ae9816c9a44979918d488290a402
zd750bd62e245de36d9fc268b9a121a85177fb9353f467ca01f35e7848f1104db4bfefe374764d4
z520171d66efca41727c8f62fde73da1080fa4d714ba1b1675340152e9080b18f056d65800c04e9
z40db824d692c4cb9e1e145f79667410ba75d51ecd6a0e1b439b3f86696430af90c46730d94ee70
zd5188260647efea8a568e4b48dfc8b76737290a24e0250c796a6bae2c0ee12c41c3d88a95dde3a
z1f3947a0a74aa5fb0efbdd02d639bb2057c6fb87f624d71e1c4898e9904dedf97b6e93c0e40deb
z3403c02d6b467500463b8cbbc8fd12c8834bf1d4878578ed41db8eee20889ec01345f520a11ce7
zf33f01ec4fee21e0a4b327a2854444db614904e5e555151fa5274cc226034ac67a48c924ccbac2
z230c8b8482a3797169b34b2ab60c825607377a14fd6e1ea77294ef24900596a9d5cc2068c2a31c
zcc305e4fed359e10a6402c0e397507c8525a7af1e2d59926a186a7fa2a89b44555eabab30445d2
za857c34320f3eb6264a45d079c969c0dff29af3ad618ecfe8663198a73d9c66ffdebf0e24a5e28
ze5082057d50ea82ec58441b35612d1f8a415cedd263df0be966de21e66f05367003779ad1ae263
z1517d3eb456ea919b20c93655bb410bbb8fdb8019ccb11f5515e2693d1af44c40aad44e57505c3
zc48d28a77549079d9f7840e17915193d283bcd5e26569e120ab797c94d924cc67fc58c1dae2ac9
zadcbb805ccfcf5ffd60b76f008a73cb793fcc04f1758b6302b6fa2fd4c7d43ca5c25fe1c62fc14
z0b6806fe01981d5ef5149b13e261d50a4df436ea98e4c272bc3bbc4b7668adef22758176bf3659
zf454af2bcf986ac3df3060a389b6253baa0b8a016297ee0604852a5c6ca91075819fd78c7866dc
z148b623f168fcc02f1e2268ad15b6b6858b8661e378a32a31da098f3b06d1491aaebd43b9d0e23
z34bb4d4faf61f838a0fbc7b3c8a493f988236bd12702aaab15d042b91953d4aaaf46c33e486cb8
z2c9865473971e5471f6883d643bc22b485dba9771405411483da9865a0694cf8c130deee816cd3
zb17e03316c0dbc9e8e9feed3e444f7b1a80f22c9a140bfd8a6784bc764f70e8e0ee33abcfb4e23
zfda0cb7fe6c6331f61c3180ee40adce2b39d2e869665d26fc55cd1cc04547ca0bdec2c9075994f
zc5a907072462eeb6e422280d473cdd4d31e817b5e4811e9dd289623aa5a1b60da87fe096d891ba
zbf2ae561121cf70535e6f6544b7f6721cbdcbae056dfc083b39703c3c9eb5d23616779621e30be
za84a666bc6f46b49b669b3f6ea113b1a87e464c50e7b05c8a500c7262b85575235a54b4f78fccc
zc72d1f9a5d791022351e0b5e1db9859d614ff134ab0100a055034eb3bccb26480fa198b917c156
zadb7a69e4edd91888e407930180967a8e862b7c56f424da29ceacf506c1280e071b148b7ba3dcb
z0588d5294c75bbce8ef792cff928891f75d5723553453969e0b376f07a8057b137296d43e79da6
z257efc1b455cf56bfe49484f404e5793a0aa5a2309fb542802b9514b6843e5396d8b6c53172c58
z3c28eb48e0f0cb943d5022951561c71a68bf369ae7987e6f03164daa28911c26890f269b7e79c9
zfb220154b5a8c2e6e81562ad844c6fba7d9e1549f824e3f202e28c89b1b606915347385df55c77
z118cd0a28842830d0bd559bec8db163303483554ca0d33e08ba465e251d324045d67cff174ee3b
z56585901cd75f60ac6f77d84400b94a71728ca234bac349106208925d46bc08c0863720c3320fa
zff2c93393d264d7b8357553ab10fc895a5c7ccddbfa07a229b3be51d771c1b9762087911f534ff
z1c38574dc0f5485fe2875adc80879339008bae5b2c06f4a2c8cb18f21a9120762ec689f310ba9c
z39bfb40640dce5090d4093badd8ab1e26ade9439fea7e2f60b6f0f57b9025143768b65324a4fb4
zd2e72a1706b2a275ffd479a6c0be786bcde8b306c8d4e1bcbbd79e35907bbb2bb127e42558c302
zdceb6e4a08403429c045708e3690be2fd8a366c1951261b0f5b3f85e4ca2ce8c74d26b1f657d4d
za6643fb1446539279a50d01e2050e1e8f5b2b5b0411b9f9b1c32c69343048a4a6933446d36da4b
z795afd6d82415dff52f24cf9bb6160bd0515f200521251e1d2eebead4dea2bc8e654c82147508c
z81ce949d4c515376031f5ac9828dfb50774888a4d6f701a2cf870ed6fee8c134bf30d99e55d42b
zba3bd1a031eef3f17989a884ebb55b0973d014a68d6c32c92ce7f305cfc7e78a5927db77b0730a
z27b815f34760004f5fbed2eefcdeee542c77e7e02f95cae332a9b0a2d166af6cc93e031404e760
ze1a5b6476b4a900936f7a4099129a10150ca8905cbacf33d2dd3a7f4e4c84e86f882b9a1553935
z6e6948c3d9d6fd84bcc492d9b50412a8458704ff781c7d2fc4483909f8091d02b264c42844e372
za794439e84e9433d2c65f6d864f1711764198c37ea018aae30ab51fe4c6366ac30ecfd95215c68
z72749d9fd37b6a127540ec20135bb40bbb44ff76ba557d1b09575e02b21790dc015a5b105c5f35
z0ace4d5ed8a28582ff46676394768b2c73c449dee72fe3790ba94b2e5d29fabd48283fce65da39
z592a8f52481d155018c069b0601db01adf80cc2e75306059f2e376e4f1e91a094496ae24413ff9
zef7e3eb10bd48bfcb2bd5c082a8310d03642ea3dfeba65ad73d394fa61685d824b357e804c963d
zd6d54578345c519982760ca51adaa30f38a44f5529ccfeabbbfa0616751e6763a796d067c948b1
z071795cc2eb21f3bb3535f4a00dc6e1648de32575b35c50cc15909adf710b6fa474088aef132e6
z0f54e553b802234dd3b86df3ca39b4776978dbacac2b91bb0d089143244bc7d4826289f55ef933
z87e575516849644db8271ba5bc10367e76c4e9a5bef2926db7e36a949ec58e90718e71a37e979f
z8dbd070014504de43c763122d6a9510145efccf5a9975b9c08acf105cc19bb42c863eb84d0ccbd
z67baa80f845d4cf9be5a878bf36fd55c3e9a4fdcb49d9a89d2dac77ddf7a41ba08975417df0b1f
z559b2c7866e41be535572681b3ab40d402f5f1edeac041d35392264c23bd04b3c66d3b7560dc86
z951d37d28a87b8c065d81c9c7a82899820c9aa5e16bb7157837d23616a1063c7bf7c1991614309
zb19ce9b8475aaccbeea241cae1429e211ae32e4d9c3ec48e31879f3a5263706bb1b46599601335
z3838c973fd189ba6a78a258bc715c97e7217d359b0861b126ca4bf6803aeb136bfa89fa2844e29
z5bbb4354866435ff206979656f503237812e3b324ba4050968c406d8ac69256d41a86681907e92
z7a212583fe002c81e2882afab3c8c4b9c0ba2ae1fe0f5044017719dd10decceeb1cac8408f85c4
z3e8dff17f67bf2fa0fb7c116198df3c95e2a7831cf4eea654644d399eb04601524e1c6067a2f4c
za719895578e971a1f90d535957e840812f28fe2f25a17967f8878c2dd14ae665b948e092fbaf78
zdb8378373edc9c010373825e1007b6bc0125214ca14da68d7af6338e39f50bad7aebc9cda18293
ze29820feab1c4086533497b25730739439b80c9c56f062acdb9f2fc7918cdab581fad8d8e91251
z0b47640b8301705dd9ff4a4220363b69623c9350795c4808594f8283102fe310d975a02e3b0270
z9c54144516bfc0faff427a706e56ccaef5c593179b00bcbacf34c5b896b2caaa7c55011411d33a
zfb1fc0c3c0940b43822fff2bd6690839bd2588dd3bf5984b5f97f80982895cfb6f0677902ac871
zf878bbf2a4d7431fb7ed37f6097afaef4c7451feea2ddde92946cfe75b7db397d0cf23d215db0d
z541e8929a12dda35cd1e6b1bd547aaa246bad363dc4ee6f8c62db6013f19111f1fa11cb8ff3eca
z39a1ede3ba5a8f6ccbbc01e5b337f5a3326c55c6afeb8b605b2d82375d5ccb84c6cdce28a3ec56
z150082db881d140482f08898d907f54ec2bbfdaec060400934700fb4349705bd34cdc6c6e4cc85
zf422616ad810dd0b5cfc873a6aabfc9ce05f22130a1d25c8e73c74d4cfe418ee61be5f03559aff
ze678bf834d5a813eb6a3eef603ddd4d3fc23b9b0387ca02d3cfe2ab93dbcbc0828e1ccbfccbe79
za7fec6d3294ae8c3c8c8efa166f8796d07b2b5cd30f7bfe5bd80df75b999c61e35f20d74c08639
z62457f7d251d8d43905151cf3644fb913a5521f299a366efcaccf78ef0b9d58517663760669dcd
z3cd37b5f4b66e6efd70b62c1780309b6923d7afd4bccb2eecf58046bcd6961335fb43681caddd1
z081f46c18c816ac02bb2e06ab41ebc34d8c6e83d2d0d458a5cd48dba7ce42214f606613be00b34
zead009cf7c8006777eb99af2ce51f77cd795dea35f44763d5dd336cd5397c65cfec56711f72346
z4d3b3988958c84c282b52077930ef81e7be4d4a9d275d0ae68601c22f735d0f22ab798305cfddc
z07319e7dff58d2c9a1713051a25e31b180d738afbc1890be73f673548a855ce8e41d60b89900c4
z8465ba491022b189e288480cc278269250c3abb53367e931c0d542fe6a1921c45fbdcddf0b2599
z0486e4bd8a6d2930ba23f7cfb0ef70427c1a2b45dcaa8d64432caf64736d2356dfc566a78de2ad
z4cecbb7ca3d051bb6bdc48eea7d369e21e27baaf6f40b16ac51389d0dfeca9b7e86f16b2343ab4
zf008b69ff63ca762d905875f049abb97763347264395aced4817ba2281f73d399db418f5904620
z5cb2bd9f5a7d76a8b2ef42bbdb0e7ddacd1726b15e042ff63da98b20c0782f2cd0b8e5e2590187
zeb6cac7286d1a2c0f2765fdd506ce523dffdf9bab5780c4cc3f63675b0b8ff1188d7f067b734ad
zda4f579ef5a85b89f91bb3ee7e0b05ef38ef7d2b71daee363bd60ae67b7f53217f8025d72910b1
z687fb8ffff51fc890c23c272e95b98e112ddd71c579bcaac6b76c24083fa9b24a7fe42efb19855
zb2595a6daecc3481d0e025c8042689f4edc484d712cb64effc7b36fc9b2344d62e6c25f4a8feaa
zb0e92ae1aae884e9cb77cb92106669f57396db3d3071c4ed3db6459fab0ef62df747328b399496
z737100470232494002fd9e7b8e54dd473e859fa7ccb36c6dc900b70e250264f1065c6433281e98
z20f3c2ae9933a14d02b321843bf7eb8337ee626981bda08f775ab0b259e487acb1b1a0eb03f8d4
z03fec35058627096194c8665cf255fc0a2df82090a6f1e37d9216b388b17f252f41a160a62456d
z7f3128ba778f696579007dac8363ccc96b8e4f9f612c4bbe9860a5c7dd4336d377b0ab72b69c81
zdcdbdc9f07f1bb416e3121aa14ddeaa1b1d9bae29ba956e377f8410aa12a216811789b0dcff575
zdaa3e8d6d7fc0d88803abf00e3efb487f0217ef22de322f14b18751c9f38b5594d52572f39b26b
z0ef3dd6a8f66fe20f51f246ecedb877c0898737b795f9233fb8a64c33ce4085b3c150315bf4694
z418293bae42bb2efa4fa718d9f21682500a334cd787d56f6632cf1faa6d8319e4b824ae9faec1b
z5a78e282f2784299ff1b159fc8290b00900c16e9a16a1a89b02fc7c537ba354d55d215791a9d0f
zf95f74ea9d88ac5545748edf957c1bc28ced903dac24b5ff8527c5bf57380c08908ad98b6a14ab
z1a74bc5454bfa5b8c8ceaa0eba8699c21313a26c96dda909eac31dab99328a1a234f68ad9c79e5
z7aefb514fabb53ce31017c1089a503ce3428324b21d0aae79a653334bcb98715cbb0c999c8520a
zf1a2f671dbc2b533b94a8bfb1325ce7d447bb207b73e6345cfa37596debb93488cba78f82791cf
z17ea694e0b2990a79c283fc02b05976f665550446867959df97015042520bbdb1a3e85b5910dd0
z559805c882fddd8224ecf12dbb3bbacb1e00cb176382709ec9df64247a6111d10cc64e82fbd03b
z4275246904603c8e320b045730cde86b4d5e50604be53983eed11fea5b529bb5cd20e47abd6f3b
zaf1eb84031979e2289b59f0b598a7a639a7510e799bb745b0fe29b6a9769a7e3e5ff41fdc51666
zf3b513901e9b88471db86c527cec7115d1e4bf32e7838a7161a11a0d1bc49157bc1d299d40670a
z873ee737fac1fcde5e379135389e6a662ff0a85c1fa70bb1601108c7cd43432b84be2580f04ad7
zd1e72236f87e352cec7974a36113efd1a0dc59f92c04bfcee18fbaecc0587d2d87391a52f39c82
z8208368ff0c3d05161593387f30234d15118f506966f8b180a32c527a45dd81d2f65c9ce6d633b
z320fef212d423dd5a22cee9733d8972bbba051193445883b2db9361af909f2bd85f7c65fd4b47a
z7a2123378ec0cc302c09598e1cdfbd2d879e675e1214eded9637458d5188180784f3e40a479cae
z2c4a107c7ca50512a8b8f8439f832aa35f5066f35da3003669f4efdf9229a2519acbcf4f7fff8c
z45d6ab977de90ccf7624f37683cb3368de2743b315201143150b2cbaf433b8501afbe99c75ee8b
z2f0979167bcda3b66a4f2c5c5cb8e6d80a17f20aa1fa94bf8bfd2097f4e47fb016a66d53d25462
zc0337359fdcf9372eb4c084c24b467e61d1be5617164695cac0ed7dbd3aa8c165f0f14f7915f4d
z2a28f20ab64b7b455278c090fa51d57a4f223645c145815f16a43c9b706b926e3b5fb1afbb4890
z609d9b85abc87e64206a401bbcbbebb28d9f12d43f42725d82f347afea9cdb775d825b80c74abc
zf3e46d28004f78b298f660090de64b7b86e890e0a49b39c486002ddebd71d6b12fd234f69652bc
z6153769d13ddc7d0d92ae3e97b992850bfead98b93f80fc2b251fe5ff9d87042344bfad35e40b7
z0fcc684f50b098a11274cef981b315e98f9fa09c3c08918b0722032a46361af7a69e54f5f9d1ac
z12771a179bb0b9462b9013e4038bf42e6f1ad642aabe2f063d343ed787c2a46599b1deddb9ebd8
zcb2597279310827966b75ac3cc9efc41e4024e2a46ac922c75cdf7d70c9d5f0ecaa5372b4ea666
z1f9f126232eddf9d544fc744a2d22a25f35bfa2f209995f38197b67803c857379ff3efcb3bba05
z899eea03ee575c0d0eecb923d98fe90745be89abe7b0e8c43279ff2c4066c2b3697f9bf4d53a68
z92c9bd3ba85e67c46bf1b66873ca74decd9e607238f797e5c11e36b4c15c3585d4a4c3b885bf18
za9b9bf672f78bb5aeae30f7fbf697ac3d693ddc5225022090bc8a1c2f0ee8b41b6fb960c9f0f21
z0b937d938e5a5a7c9905821f1f60d91f7e16505ddb683f6fa752736161e6a8e83b79824d2ddddd
z0da336078f3d648f4cf652113ffaf362e40aff9f2685a61b8157f696d7acdca228a685d51a502a
z5596f9153d9c9a6f8e367dd78f87a4ffcd6018049cb43c36a09b0cb8d88d47fba30299f35e8fce
z0ec75ad237126815a59516aefa48be84b355e2e69b4d91be7b3565720ff8a187e7977c36a280d5
z418f3aa787f09b13c7fc585c1516025229eff91a5aa7b1288614a0f4b75d57040067802f6fbb40
zcf7466cbdd341f8215aa3ce15e7b467de8d4ac1366b2bb48946fd19be59b7714f15770c1b68bec
z8b64881350a6defdbd1e2ad8c8b215901606d7e501f60c0a8611c1137634ceae863f8ad479a89a
z0f64017d8f273debed5be0bdb0f1aec0740d4b36cb39f73531e988fce40eff7e57eabd42158c6a
zb9a0bbf68911721e1d7cdd0b93e8e73626bb267328182d1b340993037d2c194ec804150e6b78e4
z95662db41daa162fc122ffc3803244996d54936600d74040b18a55ec6ae85d1859ec26957ff26b
z569831debb71ad7346fc5db986bbd14202f337da09e040e9cbcd0926e649dedc7fe88246db9c67
zb47afa8a1633e2154575bdfe36332a6ad5e1606ab7797a1854cef65df6bff5ee79810c970978fb
z015f02034c28c91d3ae32b1355b2da39f9815ff8316ef03672880b4700804bbcc2aefe520c5656
zb68435c0ea5a1269fe36187350adaea647868bfb3ee8e1fc32ee67b233ed7de91cc1a33315bd68
z5b9464b4a9edbdbe24d9a68a2d6bd5db75a4da5bdc3bc47b89a1b6d089d0f72985e5bfe7f9254f
zf4eee18106558c880835a3d09cb3deab0c0d4d72f6ec13fb6e2b187ead67e7a43e7eb5204729ad
zffaf7c7114d5e5cdaa98b2a2b88d257c1cef29bb4aa3bdef232725f07b18530cd35b2d9fd29149
z8627595353fe9ce6f10f31af8eed2512c1d665f4de6bf2169f757e59acd47646153680ee6c51c3
za47d9a84993a93b6180f6f9cd1744ab81663482248b7bbe846999f15690e0caa1688d530ffe6a4
z0e26c8a248a63a8c6d66f9ad8c54bcfc0169ba896e2b29d0ea5e248204dc0d047883188ec8fd2d
z85ab12c9188bfef9614fd3e3965a1498fa6d02bcb727c123db2e57fa24248963c2de822ed48849
z57104f47145fce27a2b1fbe1a087e61b7b82e4c437f1350161c0bc6ea986333d07d484d0b21590
z08a0812f92611d3a4dfe72cdf108501ff3c57003defd53c76d13da997658ff3e3c35e15aff4837
z9366acfb3b8326cf063a913d96704bf5705f48b83d5105be5b7cb0ef8645215810ab07c123d095
zce7c0bd280f0888c75093bf0930a190c62c02deef0ffad9ea841102e3d1bca73d3ef5ae78c037d
z1904b5a4f2b9ee8b5a35c97d0391571c5cf9a584fa220f9fc4538c6587a3bb90e8a7fdf40f42dc
ze46c485f8c15de536620e05190868895938e5d4d8c139d6b865cfd6e10ef25d31dccaee5f240dd
z19075bb91d6dce34c414eeb0ad6cd25dd18883910c92c8457f363b108550a018d3e48857f46a24
z8d21a0f563031ccb5749c4db07b4d02864346ffcd09505fc326e4b7a9b356f570a294580640ed2
zba27b7f8a8a31ca244939066bde15ace5393f7729565c254cb4c23113844cb88a8a555616b7ea3
z47d73235a58eda2fb9c07dd59b6cf089cee4d7cbd4e1d468b29afbd9f977567b11a345b97d34a9
za06b636fc204f2ea71b87b671067492b8ce79dff985d08ff7ecdd68170ef3e1e735a5c415b3d62
z56c34e30e8362066f915cf28262a281d6d6fee4771751fba05faffdeee5b142cd6c4e70c8e223e
z9c3639bdf998edde41afd8f796531a54f46f5acacef3a489676da54d491a5f09e995837bbc5a1a
z9d1bdb1e82cdce832c5927fb08a52738554ff40ce46aa5cafda7fe060eca466751c1f429be35f9
z399235d2a50edca869d89144ff98c95bcbd5249ec7a41b57b17a3ce30104a524fb02aeaada8ab2
zd562c4a7db2258599054a865d033ecef7baf3ea64ccf4ee4e655f1e9dfbee9f1b7c6de8bf4ce92
ze39ab2af44e8a8aba1b9d328dcc6702569269b4819298f26d979ab7922438818c7123d4b12031e
zac939c9a0050c1202ff9f0bc79b0df0a1b439211f9b42ca8c66cd982c99edc7bfb89f42faa5a01
z7a12fa10a9d857fce6ce5929e8aa57cd44cb1f7ef94a116005c9c8eca928728c6be9602f97f4c5
z9a7a2ebf21387f8c0e27f8a182f951a1803c83ce911742f1dce789337ac79623cf7fb1ccc31405
z27dca6ad681a1b769e2f66919e11ee65d5b9fa19e913bf33a63edf2d227e7c9cb48fa533f016a4
z45360b7bc0d3a619025e4f7709f5ee46c1c500d4d0d0b0b4734635e747505fd7ee63f69066f5cc
za33cf2d9f0c3836b17c1fe3d4133964104170d3edd475811efd329a426fedc5908f4df563657b6
z81c4d21f2cd0589c634bf54d7a687e1d869b33240f2add36f81d3aed7c2a395214128529fa97ca
zc539ef9c26a9c82db9b33d6220a99ccade20216e341abeb570f10410f0f9de4cf3b6365b1d3ed2
z6c4058845fbf74686817711fbb26d15881dbb01b2676a17996da94d0397f245260e5f883c310d4
z9f7eacc68a5daf0a42a480b982e625ec6a55bcee6a35c1342d5733505274ed77abafc8329f0697
z178a0dabe4f6eb83b7384b62df47c586c67ec93c1105df28bd2e4a17c6e335da97af835f90b246
z2a92d1f3c9ad727ee7a5e8582f8ec887507a4a7b85970628b1d85b37dcbaed1d47e40ed2336738
z817bffe0cbc9a52881b2700a4b80cbf5b47c5765ebfb37b0c2f972dc934b643be5f4f768069a4c
za1949cf504f071e2694f7721d4b27d9a753383ac6f8296768ffbdc0e238cdbeec7447b5037e424
z0ef1cd61f6760a0fba50b83fb279c34aa6b49b34e363e2be3eb6f3de21ff1f0a2d7e1cbcd53ca2
z96e200e545b85b3c1bcfee237737a77c10e0be09758f56bf53b7f4b8fba89cc06a70c822a24707
z69a6defa0c3b8d12b3b41a80cc389ed43f588dc8dc746b388528d34f5b08ee26b5ff36b1252505
zd08c3ea2d24b894179a5e0d76a3020df664f2d870e8d7f806a1e2c2d15fa22ec40d3d23b355f1d
z60306aaf3a484af3ae92264105a37b5137b602d0465e4d05f5785aca31237a8f69b826c6e9b3db
z622c4b38fd9397ada496f33ec0063d5ee9bc233227437933aec2a4cec75990027a7993c4fe7ea4
z2c27afd63bdfa74be31db2742309e92e238a445a74d913dc23adefaa9840520a2d9535359dec58
zbf9300eaff80bbd741588147fb68867e3056c97579f7eb5d797da8d6ba5b87ebebf129a50886b0
z94690bc11d1a4c97e7def4d1e42a97f2933aadad220a318ef2f1983969aeefa1d35b0571e4ce72
ze8ec2e27479056e1896625494125704495131da168d45ad13175f0693fd249e5ba7461d07f87e6
zb81880d44b88b66deecd7f3c3dd6d2c9bcd0a3deb0eb37d343325e89ffa6aba527cc64ce2a9b98
zb58088bedbcfdcc382c24ff939178e76bbc454c57637b6c71c793d5600744e05fcffcc85331804
ze862b4e44258e7af15b5f93d9d39daa79f898b90291cd22bf1152e15166557432291cd22a1b408
zecc8bce3e09e63982bda41290f7b92bbd254a49dd1cbbdae3c240df46ffb44b0fb17b17cf296e1
z2eec712b1942eb4144f3e45cdbb23cccab3f8f4182a93ead7acc013d3eae58cd277b75f128aec4
zf34062c645e33a8ee7cd6f90d5e8e3bda09d49e0176706e2e9555e5baee58bd3057c9ecc80217f
zee83613519e454153f76050cd62819b7f634aa872b233b990eb0af047a416476f296a8031d14c8
zb9085924bd261a33534ffa4f227e8d8a2163d4d1770e674f2fc1651bef4d9bb099212c9a1b25cd
zb34b478ba4e96543e52116b3d425ba781fcc51414d172c492e8d088384739d5d1ee4861628326b
z808f5c5fcf749c14bd9146f160b166ad63ba5ce263ea8148bb27a8112d265cb5036c375179ac56
z5c7ff31e4cb4465f8e6991500c9ff97187f03be8db3643ea5d993d4e9543b6b2cd8a368846ff9d
z465934c668a796148e56cbf10040011f6f3725b7ec578a9a504434262d3020d59e157450370634
z9442c6e2951cb198b26116f31a0ec447a6b42e8d62cd02afeb3ba69804bd5a0f52c9a728ed4663
zd4e77a6bde517faaea128cd6bb4582ab8b92ee173658ec1dde03d11387b8f7ff30c37036ef66ba
zc41ea60e09f957eaddf57259509036a88441f4320477959b7c824f6d2fbb1a56d84aaca863b435
z98e16e8bc1c51af67bf91bcffca48a601099126dcdb514077b029e8496672e2b8b9e09fe094717
z2edbb9b94688e54ba4f5cff7fd5b312f9a8e2b57223be036258a27909c594a456b553d96462542
zedecefc74a3cf70ccad93ee22e662f4c7c9583a1f1caa8c3dede5e77bb6dcb29a73e2998f37323
za849437d0b075e13babfd64123136156a9b67e3bb698e476f10a794174f9c0bd8d69d613957822
z19684201cb1c3c1485220bbc0fd155fda7f6c4430a56862b79ca83b7c50d1cdf720bd8f1699e87
z20bb1950ac611501e19956327a8badcd4b06657c4d68395ac0211ac5e29cf0ac1ca0857ed7b9b0
zad0eb91c3e4f775b38683b38dce586757c7e15e7a6f77a25296aba92640217309478d3465a55fc
zcb1c18a891a2bbb36f8b4b925cb8a7e5a22ca9050a168b7bbbe7c8112b80ec458f207830cac69e
za58ad93e9461741b4b90e9ceb5a31513a7bf9c573bda4513055b22ffe780457f4d4cfbd4ea91c4
z9d2d3a2537f197347805b5d465254371b3148a1d5c160763db0728a0530631adf61b1be33ba47b
z9377763c1287fdb01e7010996068bcafacc3bf3d459af1d95ffb861024531074e352158fb4dc64
z6b77d9d15514681f0edad80e3d4f67f0cadb962af271cc42c7e01a18ff59e15ee4a72d6cf2ca81
z6595cd45dd47ba8dc753ddf5a3bcfc20d666f07b7b01531894a85ce392753664c6618bdd1091e6
z92078305a3e62de0e7123c5bfd292ce2bbd350d182b9f876ec5e652a03c05f42030c01b869f2ae
z773962d1ad6accb7ecb266276e98b2b33e064af688083e3d1e5d069cf8ab8da2321726961318b3
z75f3363e9b1d4b7247db6b801fb487ee4f7c540abe67d4f3ecf1cee2acc5253a22d0377b57a304
z8356b5c0c3986340935586580dbc5d4601c1d231ac74b6a45b52f4e62665f0006f18f8fdaf9f5d
z944b5aad977f1441a99d1c1fdad816ec0effd47209ac22c40ffaf77d2af8714fd4bc27d1158fcc
z1788445a9938c9a7502b85a82e147be74d255a3d855d462dcd5aa68f822279a6193de2d44f4ca6
z7532cd6fece58896b5126d58a00a293b759617f04260e69302e4b6bd49159ef2087512f3bdb155
z7901c38db73c92d80a53549f1a02c848402b171e3b98e9625988536be511d452c39dcbb520f9b3
z2b8cd028fcaff9e03b3be20ab895e01831ba6b751d99ad758ad9bd26c2a1bbe972a1a7cee2a0c9
z82a9acb0315aa0c11122d131058f96698f10f312c457b84374aa963045df9f786a1292e8198c82
z33cd3796e777bf52fd1f35eebb5b8d345faf833c068deea02f6eebe93f0fe5d3ac2fc832c1a716
ze85c4bff84703ebac4a5a34362defefa9de8b34de33944735fc66408371831323488480c761291
z0cb50be0ac9c08fd93af997cef9bc63a32a86ec02f201b970c80615fee5603b4b90ad7f38e0293
zef13cef4ca3b7a37af4d35a0e9249547608c9d20ad01e61294abab2195300f03698ee1c9b37211
z053757c9d769fe5fc741dceec32a8720417699022e76697044724fb68ac32a5838d2bbc487eae6
z4ecf8fa4c2f901fc33fb1549a4037782035a2d56abcb343619de309cd126a27dd36de21120df1d
zd6deab25c0ede2cff317fbf98dff281a6794f2a17b2321b25259c0db88c0d6ac330d39f370bf63
z0aa042cce4de48ed04158a7d38bef198d03ae18e51c20b93d6375cca04cadcb84e3f397cd9f776
zf5d6474e93749af0af2dc04e1dfe22a7a0fea26493a1bbb81d45fc177eabeae732ec46447a2b03
zc2e5f4b59ce2b8b121530b8062eaf9e861209b3287009ac81326624184bd1bbb6a0eae8ce74272
zb14e3b45915714bb64814c9b2ca76c158fdfa3dcd81e566637c7f55c2c01a7cf466f42170c9e3a
zb8e48f7e379f25b8d0f6100074a8eb9c04c2c7ac5af7d351c18208a5b802d06be5dcd035fe74ec
z2ccde619b54e5f28c8ed08a6eab8d4550935db20af05f93c74ba940f355a46500f0c4f099e8d63
zbec8e502bb58732936f3a817ccaddd75c771697cede7e8c7893866b310d788089f449c7625f912
ze9bdf1d5f9b66d9d7a1b752ec3e7ecf983e0ffa5ccbc694c857dbefe1d3d15d348af74ac97eca2
z068419747f96406dd605813b9684331a553e450eecda0ba2c15955fe4d3b99c8c672fce3f68961
z56f58e9426e9ba1d5e16e99089ca2de91dae99052e635cb3dd2c64286b9ed2a935463e6e3b4b7d
z5fcfd5f8eba47bbcb0e8360fd99b8922dde5bbf1593fcd376959fb0e825775af84a8eaf4270832
z66586c1e19e5ea6a1875c8bf2f837926b08d589d1a2aa3c31d203335c072a9afed036536a0c4b7
ze338630802dc918d05f39b7e2f9a2f399ba4a30341d15d5b2113ac2b6a9932240ee75266312896
z5d5360253b0b5a4756b1c8bb00411e458edf562327b2dbdd99bfc9cb6b1b4f2ec6201c08b436a5
z5b2b36e1c85c911c882bfeb37f0453dbf585d77091260403ae17ff1dd5b4622b2b0c58ee6fce96
z97522645ce87ab0138926c845a8adbf171e3dbc5b29264627eac02283edcbef96b08f7ea38eb8c
zef72c489d2b59461c80fa29703b2cd72b02bb75bdb12864ebebb828615a9be7cfb5bf096602378
z0d50d13fa150b09f37d70ffd7d9e2c67264005e17b3b296af55bc49575ccc5dc98754a117a35c9
z35a34de54272d1e3a6a26932fd4b0cdc337ec8d573cdf94ccfc9ba6d06f84185dd421bb28b9299
z3948db0e6c3352ad93cbf8824f0ac15f16b2b418e186dfacb4a40d127de1857b3bce0154d58900
zf4e5d83ec826720b1cbe08e0ba8715133b0601fb663c57e87daba16cdf22f4ef9fc044436bd350
zf4e2162f776f46ff26c87b7262ab7de13bac63d7ff815c15a3ccd749a75eb031ec640d6aaec0d4
z2ca02720d1a9afa76a5c845456c61670619536b32730c288bfed175594b2a47c04a3a6a8ad94d8
zdba9939b79e5e453b22b73e94975f2e63feeba48c3756db45645977156f1a2507b238b30bc34e0
z1d5af3d9d6446be4d04ee4d984dfb9d6484ea340139cfeb9a22d121f1a15fb0639a610939cf6e9
z7b973f18273b2407c300414288cde31371b5f4108ebeb9605a0bcda4f901ea8d8ad09c7e4be30b
z02abf731b4abe288760f399879a6c34ecd84c8fe3b40c7f4a04cd17318e1f225c7b9da45a40e06
z6e7eb59cf6ce5b5a332ce0c0ee5d8959cbb6dd728dd02ee3562c61a12c92c6e944c983092a8b0f
z7e650343fb180c57ad6ae68d91bcf13c4fc9ee6785dec9f18ed40b0f5df138d56e8db1a2da450d
z8648ad4cfee1162a44d30c3b5ee1b259ba8568b1d2dc942e47529099abcc9410edc7a90511498f
z18a57ab155ddf41edeb9e7055ced71d7e69d06775619e15942775a60d4f7deeacbe15338bf5d41
z7219f594fe7c3849412330c7692ff975ff4f994e7845c4692c9772761ec05f03f32fab6289e5f0
zaa4dfb4294819da512c06a6fad3e5c2ebeaa41562bbb80fa48c0fdafcadd9a273548e6dd1c2343
zcce394f6b0949faa351474b985ea541ce68a42126f991f2fcaa3a0de890bedb3aef1593c1d27e6
z12bfa39a5ff29a3e13352b2a40c41953902389e10165ca8b2c7c92d7a8f3a2827e31269119ccb6
z9160fd4e3d4341ed9e61ee1fc246ff4bab05f2b8a74640bf43529c448744edd9c0f8122933c3b9
z6a4c56392d8f63a4547db9213b8a7e06ef7b22c242fd7e41036b2ca3d6e79dd68bc1a4b645ce5c
z927515be1d161f0e7dd8643ed778fe4874bed981596465ba52b316a68981c9b57d85c2e02e02cd
z48352a2bce2b4225ce7bd646d34be8f6a9e91b2e19830079f1d0a12203c1aba1fdb0ed04567535
z89a39fb232093e9643d4b6e9d54e6722c1cad1488a5331d0338e686dc8c1ba31533091e2bf49f9
zcb2cc08236a1e57186d09622b8afa422da8a0a12233dfc9eafebeaca7cabe25888c59b9c8ca5a7
z4e9e5e5f9c6e7a713302355c1388a960dd8ffae3adc628be5cd8e556643917969382435606cf05
ze824d786b0e03a612f70cd2e5d57c3ffdaaf837ecfada3f297cb1771e7b0556e61b7252d9fd509
za4cd8caca9733586a9b52479783a639edcd0591d4eab3b5e5dd1da6a42d981f1d5d44bac6ccb04
z9e4b17c7b4b3115dfd61ab8ec54289b2897596068f2d056e3a232d665a41c55e142afeb84f9048
zb35a7215f9f0cae53c48781ac134b97224df0bf698fea79dc1d77af4a29446e628f4e131943244
z7e35532565c14f229c5a65b19dc3b19076fc42518a580d1925f870088bf582b9de49d5985a220e
zbf31f8fed56ecd9f85fa671ae7376f2466178bbd846bbea48dda0dd9a385eb70cae01dec5d8911
z5fd8c550f87d5291b2fd0c95cf332121494adb9602111c2d0e9a1fc569151cd96c860d7bb5b008
z889debbae758afcd065c1d850a4485cb700ae4a32747d7863c24b5560bca4538ea9e30e68ad899
z01ad94704c66836f6346b5c4d15854e8a59fd20388052749036b2c16e8607fd99fd52c60df7f13
ze771914a6ec617417acd87014f470a8c4d143c0afe94573f3e66be15c56423ca56044972a7689a
zfefdbcd40a4eca822697929fc80f6a6bf6d1ec017430cf86bc200cdedf521ca262f60b4f08dd9c
zb440eeeb3d7c5974b18385714698611476c877aef7ccce6d09d4f1d509ed5994255496b39fa9d6
z3db64d4907875599c20c22557cd964cc2af3628fb2c15b472954ddb252bfb92f490e659a53df5b
z2f4c89193de9b03d27dc5c24beaca18991cdbb3305e5162121ad617ebfbd359574f6546f129fce
z1978323953505dc40bbb8b5a409e3ba4e11d801373c12c321f407ad70ded3827bc9a0a7d3ca44f
z7dcf3641c4b0a3c0c78e1695f77c11667bb5728207e457d203b13dbd57f18b9678cced202380e2
z25fa5df7a41b71583043e96e09fff6fabf1fd73497e194b44ea63709fbb9a254af7b1b6cda2260
z4aa525055001eb7deddd707829fcb11ff3337333f8ab80ac80459e01baf21467289ed6e5719091
z2b95b11238baddc3f79c8b115c603e324661e34b072b725c673a00c479ca5841fae553948c5bde
z28179616b0e2bd84a171e0e54fa4a2745a3df8f014bbd4740c5f69d3d10fbcc60bf09da0e3d52f
z6223a4538752f17f7bd6a0befe61703e1ec20fbc34291ac26e4ab60a333be0717febd51dec77df
z80eee62ec5c8da412ee99ac5287cbff713a99a1cfeda6a8c45d02c61e10f9013fdfc82eb5ed9a0
z08c9d4fe05c4fcc5c31c397e4d1dfe416ba1a47321050965e857fe4aff405af6b9b94a86f7380e
ze2634d3e6d18be390cfabeed901b98dbe6aee0cf2c760b5be577b842d2e5a7ec99c751b09f31fa
z4136ccaf757d7931c6077b16562c8462b3e3873d8d32cfe7ee7811ba503bd025f08e138c109d89
z1b2d7000ec84dd0b322dabd9de4036a5fb36f894a9c33cddf2f73a18dcfa7c5d751638ce3138f6
z408760c9277908c48d6074b3ec0623d3645c58579e063d7b4ad12a189068f42d60f252f75551f8
ze261d7ac1690e7486463b9fd748af75129006153df0fd054b85c82eed68756af435cd92a022683
zaefdfa58d0ba433f0cfa290c23625cbeeb47fee3926ef619a4d59123887648b022d1e0629c789b
z2c57778eee878fc113c27d791bfbf56ccd3a7c53eabdea6221c9595b4077da2f13ce169bd12af2
zbed494b2dc79a87631b67c22293cbe75531d75f9bd78fce2bb05ba2bfbcafe50da1ad9efcc029c
z486280a25dd9db130bb25b2f2b23c703120eaaf8c2773002ee828048487107ff6863644b8659c3
z9e2f47748e3e49d8761cd44ed2fec2dd6d393ad84a8f95f09d936d6255692357075ad6fdfd2c4a
zecc594d8d83c3d61008d3bbd0575e0401cad8e55719c715a917d0cb6ba1f8230b004f4fbf63357
zecacd8cbc77e86182f12c5a14ba91d7d90614dd8f37ff12557b180b6e78816d0181b424256ad53
zfd8b0f2a3551474b2165f6c1ba9da2a0c17b5ad568902da34123a97436d0884a2c7b8127ebe0ba
z8717751f71fed4ddeb29e3f3b89428b762b97f2637bc0287f6f5484c32daf8e8ba6ce06e2e6906
zced1fc0b7e2af6cfabdbf194d17461f0e9fddb4030feff1ace4fcec8ecdfbccdf357f538fc57fc
zc45561f06a93985f4c6c442ca99fd38816938668dc89d580f9d3e15dc9d7e0b2f6aaaae424aa61
zf85cd28b75a1cc85c9c28d9ce26bd4b927c16825ba8e8ce6e1bf21f39a1975096b0f69d61edd2c
ze06fbe33794c4a76eec9ee965cd221b37474cb8c7e2e4c35a9099c906c7b714ebd6443e8aa8303
z6fa728fb4eae305a8645101813bc16841fda3eac20f2348c8cfa66a6e6d0c1874e613759dafe0e
z13e8e3066b55418e28d8ec5826aa9d44c61dc00cdc59ca5ea850d6f2ffa3135169f6e512f5018a
z8282b76a7f118a9a5d4487c6ed19e20fb8ab85b98127a95228e731213aff7068603c6013d9a13a
z9193ae9142997c72b60cf3aa009c520e5dadddaf24451bed8f16a26bbc4defa99fb303a0cd9997
z1b378b9dd478e28d90b9ed7c2efa040fcacb97a3a3743197e35942f0ca400e463de04f99502c39
z29dff605f36408f14cd47beadccbebb3e4bf57acddcf791bde4aecef6f5077c33dab9b47f7780c
zc44424e90cac924c325f8668c3673c26754b2c50b66ae76ea73d8dfe494ff5035b19ccebd71576
za0c1aaa3c3e7f44f9bf19a203c9fcec63c6983a9447c04b5b7dc7fb06e237befd4691c5628b7c2
z3397f7f95c1befb30b08117773bc5697581f23854a6cc849c04bf5b05b2a6c98876c70fd20b2ab
z1127e45df1cb7dd83c73b1621e729887e0120cefb809f9b4ad5ed26e34fe80762e8d9afd1eb032
zfe74e0a01051938bbdc2464f3ea9a727a2f0f7c4994e4b467a7cc1feff3f13b4d45c7202024bea
ze5e7c5cc6e0c6e8cd2dad1fe6361e327f9886d9ba5cad3d48ef62109490720038225add8c4e610
z51302d7b255f6de7c5d1081d0e2dca1299b0fcc49183a2e3720a01a29a3a249b7471fbe6e25b16
z42467ab9b9360bd376bc5bf2672a556eb09d7e4f4fb98937a24a4361ba5d3d29395b27e7789c4e
za5c2dd136bd0c89ca9c39e97ae04a26c7e77abff724e5f8f249227b1b575b3e6a2245dd6d28e3d
zd06bc9c19ff9442f0fb180771ed5a80d2f3d9b56b9b41ce55867d5c84f880ebda22af6f0b886df
z48809b38dda90a9c7eb0148f96ae5a893cb579131140fc5a494e702019e1b23361c310957dfe71
zf60339b4ae2eb06d6d9f8b991cfd1d45b6890ba51ab77ef43c302b5355d0f4527e8b63d44884c7
z9a793101e466064432682a0ab164653fb2f5d19b3be263380b447e28aafcafb98197fed9cd08e0
zd68f35810094526422f1621446ce21adcc8e21dd64ab340e3360071ae402a7217f827a371ece2b
z03587a9e029bb832f9454527b6178ae615dda25c24960ad1250cac9acdea08bb2d0c062767432f
z10bed03628c58d4c9fd5c7f98726287960f49f63d4c18184027b11a936d2d1f31de7aaae29a8db
z820aa5472aefb75229501a041259071224eb540d80af6c444c717b622c373a1b7201a464e2f346
zdf449aef8b378d78f513c639c75e034753126f372356c51002472cbfa982e1fb314dd9eac4475b
z3812784abf3de5e7171cbd41a980d69137d62f2212f4b060498b19d384040b1302c12f5e9c3de2
z7b920c5f179002af091468030b6d868ebf936650fd2590f7e284a031c0190a920435b441b7120b
z1714fbc7a12175f8f712b68bce1cb9001d310ee9ad00c2a594461c106615766a6a78ca42f37a52
zc5606158529c38416f15caac95c1afcad3a77e271387d45a4026bd37f833e8731819c6effc7e38
z546c455c15c84d8c888f0943d0e54a9a40cb55758fac79da738c307c71b1be301d9f655ceedc61
z3fe1f0d880c1f766760a17f74454c92b307bc0e148dffa78708b03496f51de8578f0cfca5aad55
z86d7ea6cfe599c60b1a33a498aaae95317de35fc4316c7780d2058ab26564e014e19f058716faa
ze5bb82e45f8d622a7642cb0e5c2a1f02ca2461b2630bebb315ec2ae558b114c26441167aad244f
zad4c3c139930fe51a090ea730e09b336707ba019aaa04414446d14944338a36e15d6c2d0d8e4d2
z9dbcc386e27ba3127726967ab7af3324f1c67e5542a0daa89d426cd7682a930ae02a2005dfefe3
z8f4a4b3abcc0e48b8286bfc6daf1b87d306b9a1c9d99e785a94a707f166bac7cf46a0b34383928
zc069c8a0d9e85b1085424db9b4a0df939771c0c6106875098f1aac44824a8fb64d5a59ce3d35c5
z8089069da32fcbcbc51f18c69efeed444aab3faf33a2cd0977e2f6e89134e2fc87a2e81784092f
z78ab26d97b5f45a0ee2dd0c8b2bf9e8e3ed695dc606d9a0a475c6df53ce5e561e098a4e8baf34f
z6edeeaa107d2fc3e3b1c0dc2f6aa01c298cc336911437a3d20ddd29cb983ee5f61cff62532bb84
z43353b1ec41939d47257c179c5149b0ef1f42eb3b80d08a6b4954e9b117677ffe743e4c4f77bc5
z9c2145ac0614c967d320623ce67b0cd49cbbd5ea67e284ea37dfa667cb67481987220b3ca161b7
zd160eaf54d206e2132b76761d2545f2a5afbe70c44680f3c3523edc555933c2bf859ac3644cf72
z8f9dbb3dfdcac44999525ac1b6797c12b8e83361e12430472bbdab641de232a6ac47cc56a89f9b
zb38a38d96cd9d28cf2eaccf1ef0ae1a230648db37fb963dd34030d73423e356175f68f4cd94970
z013312f01f7682b59cdde369b68a00c54da04089b6aaf28682ed10cff1ab1a08ab0a0013680824
z7221d7908886124a6358a7533938e4e1b48230c8b8cf3a919d6fed5b3e3b944e4cfa5fa87e8a8c
z01c17daf7a5e9cf889d3a05688061c78744035553b0b51c1fb1672b5ace8866553353da73762d8
z969ee56309dbd1feb4bb544cd426a2efa27147995490f62e8da349124ddc3979d9688d068131e1
zd695079540bf5d6c232830a9eedc7ceafcf97bf649eb0f1fcc49de00e3569cfd46795fcb2c43c7
z898dbf5a6e70f1220e2bc840ae150ca98a212ea7d5aa7697b276d9c83feabea2d5f912f03c500f
zaf6cb8851d30dd61533d699abdf5bfe49b4dc11baff8167d4f88eaac04f7dab077e67f45498d49
zeb25fdfa687ae427c9133ac679c0c685c38052f3b236c39d527c024ceb12156232170c4c7f738b
z46568014ea9ddf33956f5c064d418f3e1a97fa8efc17c85e69f2cb744ddb1783c9a7f8ebb76b19
z14cb1edb48b03c53ad41053f7c353f383ed986f2d31f569a80a4ef77b6567fc812b3bd01948e01
z723f7cd9175dcc19395790c22acf571c98cfcc051975f9575778895be82361254c9f2c9ff5f14b
z420184f94da16b264f65d6847972792a31ff4a40cce3b2bdd1cfea4ec70e5b2a9269b04f09fd5a
z3c5034b4a6412f45c52ec59ac1aa169e3fe45b9a80c4c740cb38124a33f50104680a86b797a0c7
z6f6952968a6353bcb69d78c766ac5aa876d5648266149171901828289cb31bcd8b24deba2eab9d
z205ab499c0482efabf1e171734170e40cabe2369396052303bd4477f75116a6fd28af67d8e0a8d
z0b8388e5dbf6763bd7d48a36b4eb885c46850d8a1137c52584306a42fb8d9e792ac2927927d6cb
zc8aad48f1386e5911ba984f8e2c9dc363ada82dc9de8e1174a8f03a977187474a6f36fb3623e21
zc3326f2c41d28ea49d962b56bdfe9c36763773d0f3deb3a05aca5fcba93f108f8a819a0df47a79
z17a3bd7f7ae00c53cac737f5ae228ab56aec9c08176e8cad9de25540adb675f45285c15cc682ca
zd86855f6ebbfa60420c2ed203ebe5fa645322e573a4892ea714db7bd460fbeb87058ec1286fb51
zf85d336bfcd36d4f9336b05c10b9a5ff8c1dc5faa379278a490c2907ea868c63e10aecd88d0f6b
ze72b2779f3b5020c369fd9509c8b646f26a7ae76a1563e153025605b485d3fd756136cdbd30b3b
z52d483714024097e99181d2c7413a112aeee989dc5b25544f1bd4ef97ef4f17aa948f7d197bf05
zc353ab259c3357d2880c4e523ad49785d7b94cf1f0bda78310b69704ed60cf4530608a233b9f4a
z1fa6e7a51a5bd62cb9da87af6c2bb25d8d3a05ef537086f0d355886c91aeea6b6ee792e623091b
z0202fdfd9b2fc34bfe76ad767590df37f440e0b0077cc09fd2b46bdd3d676046bd11db9f7fe7e8
ze0c1e93bb90d1d11a6f47f5ba4fac2c6e735872596e99db9a3ef0b30dcbd528252d59152884d77
z8ed781b07d2d34542031316732ef54c272a339ae42d9f92654a4ef094566bb2d930ccf4790f609
z1886a5469b596223e81ac90baa963bc65b8ffbe012792ee31d1a382c8ef700bcfae92b65fd6a0f
z8299d18ca768a758955a85eb2f635ab215a52498468ee79af5d827f7fcab9ea29aebde1cd0903a
zf47707b9c817c518b838e3670099a881c8c64608f850aff4f413f7bb95929ff372c0be611301ad
z4da9f37579eb176ce5192a04b6a41239e8e0e364269e45fa9c5ab5830f4cbec28ac32aed0d1e31
z129b3d533af99539da1db7ecb8b827d3ba51b3f6fafc2e318ad4c148f254f1147e40631cb358a4
z5d60a25f2ab250e6fadfe404f61829b35e8ccbf78549ddde4999526303a501109db7e9d8c84b5b
zc154b6930a5d27d552e55386c54669b46fec3a6caa1de9e832a9826c68b2739de44042019de388
z9c9aede476c3f925d5aa2643f5e8499027e95fde0098449eaa12ea609fc39d1564af634777fcc3
z2a9d2a56e3cfeea1f8211f99dc95445fa50c3b313148427dd05e6472be946d79af8c25f43f25b1
z5d4d89f9224caec114d0e9e19586047e69d0dff03f7b89f0f8c1a0f3fbfda659a57fa06897193a
z8c3279293e470c13dfe19b6ddf733e598886f3bfae6753744c32934ca80eb31f5e113a7b761bfa
z8f126b169de2ce55b7df4625376b720d84ff2964501accda409b48c90af99a4d28875aca0f2587
z76c9dd0389446953f931f0252a0137696d85683c1e34907cf43a0b1be6bc40c4f1ab0793664ac2
z4833b23af65438357b9592391692e833d65650be38b0d53cb9ea315942738a33c9e480fa42b57f
z986b92db417d6fa013f5471fa90ebb6da26b2cb6524a22b624fc413b5ba7f808c760b3471294fc
z0f53411b235fa46d8a12ff935a36d7f4d0937fff1ff2714e911c02a85b9a2ee6cfd135535164c6
zf672aafd9033fae0f32e5b68cae4b21acc2e6d5ba49c6ef1f51cd92ab7330eee099bc93a15eee4
ze2e03065f14ca1ef0d6a98ef2233c6d307d42ccd3f90e47b730a8dd1df1c84ee668ba3b8a2e1c9
z7087b4f3bba484c8e947925aa599a0480a3a60d4326b89a403d20e0938233942ed42fe474881fc
z4d090b076c0317889e4d2f10eb6b3924f03524d0514509a1a786ebcd51da01cb9e6799c5352ef0
z76f54830dbaf0e238f1bc8dab9bd7b1de1bd9b466833dca309602f30708d237e8ad4872032a810
z5ee317306593e64e85bed6c1f7b7404140c27485e3186e8111a3f6d7613f3486434034c69f8b9f
z655c454d89717ada29ebc44bffeeefd5d9e7e8fe88b3532abbb8d9e8942b9bce81df127233176b
z99026e45c91e7a30d3841b8ff6d124d6d61ebc0cf57533c3ebcc615a1bb93991766d7f00254f5e
z3b18b8e360225dc9db5c65ae6abdd0928b8c452058e1cf4355f8b72c5bca9bec6dfaf09dbb3481
z44001ad870cdf180b6758aa676c8b808777bd0d64d37f79b7b87133898361f92faa86ece72c4e7
z7fc6ea4d42f5068cb49bee2c8af6cb97edd32e5521efaaafe5d851280a1e91813e7cf4af27224c
z39bb12691020079607e79e7b5cc6eda1f46a39e0de87ef6ac667329f3ee8439d478ee9a41bb0e9
zfc4de2d797850976ac290d7a36a8ebf9c8bd92e2a60dd45a5db0a29efec03f7f7d5e7d88a17bab
zec42e276fd28d8285795cee6be00a3c4af70831dbfa898eab66453ca33d8e29515bd6c4615a5d3
z8fe5fcb0f691485375fa56e4274fe3b87a27796e6579088f063aeda0a985e054295db2bbfc6919
zc54b94824e827b0ae72eb577f742709aee0ab46f2b5046cdc162e315c0512d064f1cc849985e7d
z48b2768287c7e5a0db3f7681da6df421bfed3649e1db6594e5f3eb1da6889cdf05e1eb09351fdf
zf733ed3592d66dfd88927bde3c367a681702602dec73e68efed0540decb64b6da803c2142a2390
z96d5c8b5bdcc0527a3aba51b5ee6c9f0fa45fe7e176c57b331eae90087d0a3978f36e26520a1bd
z1c72a8f44a70df7e7dc14de884bc2f449bc35dbe97c5c6e3ac4d8cdc0886b91d282a860ff5361a
ze383239fd484debee27216c6b7bb9ecca29dc51f47b45fa26fd61984bb582259d4f2a8215327f9
z4eadd5241e54d724b9e210365c48662e0741c5f909372405dbf161a466e6931f3e2761cbf4529b
zae47575dc5663cc941b8e4d355f5a5b13c4c331cdcb735b03d0246fb9fc4bc34e09d087623775a
z495825a0be27f87a6bf62992ebbb2fe7d10b9a9fa5a130ed58ba02226b74dbd46125f8a5b05ca6
z517159347cca241e5c6c1dc289c9562e3b252df4d41daf7aea1dbfd4ed77fd5ef2f0440723fdfb
zafd7c8218d1ee491559c7f4314e299161d719f65c150cb2353d053df3cab0cf72d7d07bb833c67
z4a73d2566f37fb0ea6e179cc0442f1323b6a65f785b974d14a8fa48478f1acce8005eb5dd3b05f
z1cacfcec34c9316eecdedc541d298e4e7bb6ed89dd130ecfcb2d1517f9b8a369bf32d3d3b4494e
z997ddb096d730fb82703ad321b655081500e429bc2f9604703b3c5dc46530d8b9bc1a2cdcd4667
zf71c165a48f0e90307c068412358b8dd7aa0cd024ef88897721a340775c57156b6cd7d646c0dbd
zeba91bd161c5097afa5a4c6383d0caec0f56c8e0b871b617b58551dffb8c4dfb5094e09d768291
zfe46f8fe0fc3ea851f60bd6a283f040a1b5d46ca0bbae418eddfc67b832c62f51e8883d89b40b3
z983658449e6445f032ad3fc3e5f19572c81a585808ebab0868a760aa449a9fc64b96900c5f4159
z6d09306e3219c3c4e1297a1db2a551b61c348a254fcc6e5826af009aebd64d0f7497a0defae357
z6de849c80491842b08d536c46b4cc0d62c127ad645373062102fa87bb5c12b0801073724163645
z9e3d646e046b2ea3a5258b3f6d9b2f2f18b6ff61eb33b282a213fa77292e85dbfc16c90fe5dae9
zbd76d6681b3112d7c49a5d69608fbe570014e09152600fbb5a5ba90d753bfb7de6c6d5a1e8560f
ze9ffdb592557ea8ccc5d98564d5a73f22a383424509cb3a193744136a8d56733644749608c9a97
z2b3edbdc9207be5421f104abba05cc9ebf7a77dadaf12660b862ec3a26a481cd7b1c4541f3e587
zd26bbe75ef5b9cdc09b2171e0ed84c71633550e9a7ac4f1b0c417571556375aae5c70216e6edfd
zcfb1aa5fa34fda3345b62b1a703052340f0c464ee4d29abf19012b76b7d581dfe8fa1ff6e84f5c
z2e3cfb800cabe4831c3118f4972cc4f9795c6ece2dc5f2122580d585f741e8bab61c9a9c2e3990
z3514490cf53979e1dd7fe88855239f0737c1182fa2e26c99d5b347cd19ed1a58c1d821a885fe05
zccf0c4da321cc92bc133856bd11c30c452582c32561deac54ef85e0a3b2ad489f31495a3d4d2b0
z770131a7ff0b887022c81f41a9ddebf835d42889045509f319a77a07fd98894ec3845efb3c43ad
z8f7af3c91abd0dcc94a29715c7591fd846edd7bfc20c3015c221f7733db7d0c66d7acbcaeaa57a
zab7bbee330897198e26a94b05abc57e9947bc98872d1093c8817d875575eced6c71e8025a49d98
z0e86a75e3e8c2e7eabb326d8b62304bba0f6933b90e09e4ecfb5d19284b305895cbefa4ad593b5
z6be2e09a5c80937a5cfd7cfc886eab13c24f45295f0933c7b7fbd65a1fa207f02d4e089514aab8
z5c17fe0a59b10317cbbd12c28938ba7a2d8a914370bdb66024d39eba0717f8a63ebc9964dd70be
z4763104e869161bcd0407d19bb8397e1f8ec5ce9fbd076ddef23a6466750d44069325f57c2d0b9
z2fc916f193dd50a8177b1bf3ef9cc353ef4a9dd73cc78566362e15bc8d88c71e78fa767a51d9dc
z085e1948c154a11dc804b780aedbf76fcbfeb12a6aee884d381a42371c024f94155b9dfb63e06c
z04eda94698f713b64ddcc39ec217fd43ec5ddcd4e0615f9b3b1ea3cce2b3b5d868565f0deaaaeb
z106f96b931409109325cab6f81a104bb0ca15a9762cdb5b7232b4fb134d4c32ed811b28a21b414
z707af525cea6a6a886e392defc552804549d0f824e88b491d72e2d097c104eba983091deb5ec53
zec7aaaa10fee5d50849cbf190f6789c5a323e9f04bc21c0ff431784db8b5717aad0b1a3f2210f4
z4cafccbace4e188d814a70e4a5666a628b1721c8d55c7ddfdd1d941c2776c3eb0acebeeb29edde
zdff481cee28ebf488bc70d68114fe866acf5281f3f3679344bd297e055a4f000e8a81bb4d9c258
z3825fd703ae20ee506744598bef0cc54329f69d9c31ff0e6fec25456416efdd6fd74c329c4e9ff
z6f6b901c19ec00cd796925bdb14b7ac6261fafdd615e7489d518509377496fd336b6428ef74757
z44ffb5936799a8a68ba95521cd87e2cf28471034dfe4f800a74590586a6fb9f902c925add1033b
z6a4312691bfd3dffd77ac6cd0638b160a7f72d56f9f2e89828350ca3b9fdca4c1e2a75b75b47f6
zf91c5e7e1f753ea86ada3065f114165223b4a61d4b981002bf4a56bd78515764fdafa8f1d717ad
z39270218aca07ce638ac159e8a2232be4470643af0d8e751dd9202cf074a9a54e5cd490066676b
ze9623690f00cb090bf8e5668174861d2a3fc6cf1a81d1f42373aaf17930e25611767f6f22f397f
zd945d2ea37a72e8d25e77a833a7fc6b51dc69e387cb4e5611a8ec42decf4f49990e427153d39e1
zc763fe22e3dfedf014160cf58db475f99a1b90418559c86351a5ba861e50cc388a9ab1b0d4356d
z6d90ca055fe962b5d78c7d740c15de894bb75d9aff7cf302ad94763b45ec15e9c7b0d088ebd75a
z3e6ce34e55c4e7e4a701e9b1f55bc6d7a0dac8d5e1ffca892a50757936398e18631fdf70ad81c2
zd0b1075b2f3cda2e78b0b5149ae72e012b81cfaed7adfec5fb7506affda3e2e7a1d9da60a2c382
z478bb53fedc912d73bd298b43a0aeed8f94e17ed57d3a31d58504446316c161bbb55016a47ce53
z12f5de3259a6675d5e3f9136bd3d345cd82451a348d9d898b68e0b8a28b92b30f94e1084d0c3b6
z1a19f830016cb6a76451fe6714c1054016d8dd387d0182c1aa636750d4cadc37eb9ae340c0f877
ze0be7ac9a7526eb4ddd5fcc74809135fbdccb085092b75651004d5bf6eab97f6f43cad2286ff2e
zdce91dc8af2bb851bcc4edac25efd58bfb624b3d4d03e580faa2fe06094b394fb05600478a7140
z407c086dbefd6f4ba3a1a6149a94f73b762302c0d12648c7043e64e493b078e7993bf552b13272
z68546b153ae1b5e14eb5eb685910c821bceaa72072f09a68f06198333df3a853037194fa508c0a
z17165b378cc3f729e1be5d0b7311370a592904f9af5a9c90c6ab86134b322ffcbf3c14d1ed2860
z9c19e8d8f938045d022179405d1af7f991e89997a13242792eda320e57cd9351d611dc870ebf0c
zda53fc4788d88b8258b573f8d5ea4b2fdcbe94936e27ccb2de156c1b3bf2f3dfdfeb09bcdda32c
zf874cf851fed09f840dedce0277ea75a87471504dbb42ceb00a71b43e7f7800a9fe88e44dbb513
zabe2775809603d490a65b8de5b8e59921399be68a7127b844281ec65145419e2d20a70c5a43da5
zea2a57a700db4a8a75a07e27cde05d91a1dc82fa366e1393ba250ecebf7a42ba2f41ea5dbc1bb6
z7ce55870e4b5b574323e8fcd40e05aa7cd800870e079cc476176f0a832731be9197164db0bc9a5
zeddffb7a9d6a3e3c9810237fb99b7079d93a21fc12f29449eb381d1e821a18abfa1480803cdc32
zc9bc71f1f9553441706a54b41397377e33a229709401cfbb8f03e4a1dc8ee418181e0201701d42
z1879de2fbaf5befac1ddcb195677e27e6512971ecad4e8dcd5398065944a9ab1c6f07392358761
zf2e5422c084b016fe58a8384dfb831169339c9942943f07a4a1175f656ae6c50acc12082156f24
z93a270bec1cc9a9cee06f89ac9c6e08ed657e47f7456cc124a34e8c2cd456fd663703dff759719
z431c5e53732ec1fd00ef481aa62d3e01afb5e473082e4d4d6df851e09ddbace9ed627e34861214
zaeeceb1cda756814833f843b333cd09112cc5d79e364a97a88aaefb52199e389c6097b41d24f13
zec963142bf2a12cf8f2a1d3585be5a78ccf726916d2588b14f8e575f801040cc8b5af8e4aaf54c
z8bfd55d0dcf66cc06ab8b61e566ec4a2049d6bf50874e860a621aa5310410fd9232ed5e5a1d6c0
zf351efaf40bc96ac01a4d0353e6c72413c8fb9ff289ecb42ad4031724d10ac71f612df12f2a925
z9045d9bd176645861ff9a10410f007a5b53700ba3ddeaf0a762514de24e25abea686c5168c3afd
z7e74cd63063d3fc32c47b3e1b10e943b1f98c4dfc846c59673e1325a457d35a557c1d23abcf37c
z3115de00ed81e2b79eac285352447fedfc06ad1b2c84e1cda47b3d0b052e0a8c8d3ceebec57382
z25eb8109cbea3055b54a058c718317dc92a14848f1d89e36d0476f1ef9dc89961e65bb6963b581
z20b30af45651ea1d379d60d55a7fc9487fdf0c729078c89e014fb1d533adc00376795c60279941
zef9a233a9f272c7f8c903d69864de06071a74e64bde74869c5ba55f566b258340d982473950b99
z7f1ee45ef72ee78a4ce920707ca8be3b9f7c039900bf330d9ffb3b9b0036290a49b364127721b8
zc8d5770621c77d2e50704bb3f3ce734274ae90f4b3119eff2b640d358ae9f433b6818f85bef30d
zc7ff2ae15c8f5158335c77716c800bf797d9fcdaa1a4e23de09633d801a452813a663ec69622fc
zff587b23616f75fc05b7bf7b92990c64440385258ec0fdd8f84bdeff3ee80511f9146280f94ff1
z685a5d849ef012e6b1138e24f4e71e7fc00dbff488e64ca84ad753cb97e5b3e693ebea78defcad
zea71bdb9f36a4711e35f13dce56da88179e892198f39ede9c20875797ddde67e8d7c696714f7c3
zd801e5c02809fd6ac060fe93cbdbad4c4d04a83d09a8cbecc82d7fa90d713eaef1ba711de6b079
z66c29efd1bc37158f7cde5794d2641b2fedb022a7cad2240ec22ae14c683a00f1b42a9ad55f4ce
zd5703728795b79c044a14ad99e8899689e0b963f724a13278404daa589296bf5d922838ab88611
z98b58b406bac0db27845e2a4e3e8b0ec7bd4507469ddc5ff7a0812e5ae372a527773fe51b5abe9
zfb4362f292c2f67c3092dbbd75b55d01ee44e23d681f3a7a3c32672ce97e7b3f231c6e6bc28570
z4582300762608768c0b9a7a68c85b2a568e730c41f85df1fa643a1e1da270b3775c10f782cfad2
z6a707e959b0615383d3ce71487d762fbda439734097e1ece2cb3654803e01aae29e36cb0a955b1
zd1b2b3ee9140279f2ac66b937681b14e7a9dfd0b6136bf698ac03f8b7c542adcbb7a5e40d4ade9
z99e4d92330d2159a4064ea0c936e6d1d8ffae7e76f1b9e88c362d0bc0338c5d4811cc0e443f77c
z519b715f1dcb8b318f2193874f3c0eb23c99a9b0f9aa243e381695a598bab1aa03e68d2fcfbebe
z7d685f797dd83a642df95303512f5134f9cd610947a2dff078ff69daa8f81c82b6055da94fbb35
zb239b85f682a20241ab7316b5df6126a03ce89779f5a072ee2ba8cdbae6254e148b3d5d221285d
zd2bc73dad62a72d81955e967bcbf2dacfd4ee10bb81f1f6081b00da8d073c9d1477c1e72ce8c0d
z8fc15e0cdc27b0d1493a2d6791abdfabaf17e3d49edb1a1699240fa0c2fb74ab611bb5d9e2dd84
zc68b137fdefc206b2579654f92be593414b727cf9b697533726fd74cb716c9a75c8965d797f83d
z313a4a6c0240a8bdcd08e025e0ac4980d7f12458168a9c814cd7a079f0d64e79ef10ba082b7f9a
z3dbf9bfa6d6a9c1ab1d1469a50334fd286782ab7cfdc590ba038e71083f22fce5f47c446c61dd6
z82811d97d9e7ce831e4f6754e7afec0715faa2aeb028541ad76679c2a1c8f95b88046a5becb761
zbdd5dd22e32834a553f2bb675a32cf9744f38fb718199317434be626017c414b32d1adb55b56a6
z9bbc03b8fbdb0b65df222167d57fbd386d59f4bad56f5229cf90c5c72a3a846a8994455ec57a45
z5b31756f871ea635322121b18797483fdf45e7a5248380659533238885f3a7dc197a76560bb09b
zcae1ce9298fde939fd1517367649370264422f26dc7a318e4be6055177ca6a9877d0095052e33e
z484bdae91a07f28aeae4d6b9f399fe6c611eb8aef60139c2095758976ddbabbc6b1be4f5fcb032
zf9d6a34174a22d8a7b20f822236cad7cbd6b23b25a90107301c2d53bd142199bf5a2a6de191ee0
z4f6a2a79691ae98bb76595d287bcdf5e63949755dcb4b2b7d6aac940bc5160f1469a51cbda1c38
za88c014ff1b68769e2422a4c31e56c9025c1dad5d92c27dc4cc4945c2c7e62a771f38e7ed2f03b
zd32759325c58f277a1c24d0e15aea0b47f2faeac0148ffbdf79918ea231c8532b7818e01ba77d1
zbab530512cfac8852987b161d9887632b757ebc32d233fa2b425f2c51f361d9bd816daedf99fc7
za7ba4eef301f450976858db94e8742377a2a171a5de1ddc817353a78cdff692ed9fa6ef770b27f
z72447e3dc815a607cfbbe5f8b7f3db69aa73ed675ec540919f8dce34ff66788fd8298f2e907956
z2f21368b498b54444200f9b29d7b3ffda2a751fa58ad92dd741ea476bf5835292987b5db704b88
zc3ed68352053c4b4bf3b3ba160bf5089e1584f534edc9c38814b9f4d707eae091f0e755651a477
zb5c08d2d7c12bfe81f637bd68043db1362687373764d9355b7395285071bb62af171d4ae799069
zc967e2047e62951536c9bf6a9faaf95a1d24389d9426e9ab3da517b42943a24d85157570505d4d
z56ce2c6faec3808b58541f7c76e750dbc0ebd853d01c0b45ed2bf938e9658fa095e4f330e8c650
z114d7722e27e285b3a660e7f5e167f530e91a9f770fd0b51f7442b195891c6113da1de32a52649
z081d2b0d08b4d84655b93c8fc72175a58432276d4d611850888314b442982fac78c7c7c7cfd5b5
za39bdca1b667230fcf7f5f5b4f9178fac5926cc15353ad562324e90e8203999018df99c56a79fd
z3eebedffd8046510ca3397cb4c29ca7db9e067b13f240186cc27d113dc6b9a388ea6e8d01e1e9e
zccbaede39f792d5f56e47c0e02780e2b9f104734dc3de31cab86f89a9b3ba47448ce9f8797a465
z39f2ef74a13e3285a2681f1dabc580e647552bb93cfeb87e000fe3bee3a5564434abe95ff10af2
zd5711b9f3e8bbe7dffdcc7061cbf812f5165829c773c7c3848e92b62cb8659e25432fc8c6d9bc5
z0622a32240a0e196c5e63863609002639163734f46fa2c184eeba61fe43c9dc2f1158dd641f22d
z2a9472192a464bf6e4a84c308b052ac25201d9fa343b682f97c99cc0efb8b4c025ead4f52de615
z7cd4ff191a5bd60dee67f8dfb406c519384d59d3c6af8561ce0d1dd334e2b32af3593eada481eb
zeff3b3cdcb8cbeaaaedf318e5f176fef1ee1bbf9aaf5076aa5c7e3da67cc48c8e59b431a98a3a6
z71d2ad02d4ada7c902eb00b885ea313a6283808c21a8077f7360fa47846de181f221e78b7e4186
za1ef491d981ed64c39289abc73e2b432a71819123a2b251227b46fdfff62afbfe5f7426cb8b4ae
zad2e97510b56463f54bf28df760ced30b9d117332a1a4cf177971aa52eaae81ddd397288962d7b
zf4c31c9e382494a643b1d9ead281cb46cf22df55e528684b84b00c09abcc264e0334aa1a5db2c4
z84dd49789de6db9b0fe96ded1c6f32b753f5c3b85cd4372b9501f309d1b4ff4cde6545c9ed1a31
z30b9e791ebadfc9d31d2998badb0c1fd8b4cb897da9810e9de7d9bd7648b1f121f165d47fcae1e
z7b5751dae77546ccaf2f77a74cb9ec91ee8db1fc8050820bd11dbc199d6e376fecf6dfc4c0d186
z824c2b8d73f9b19ed5f7106c505d0a38dc71b05287c8be047afa92f56a5b1e5dcae02907dcc2b8
z833dd5732722e02a0b7ce6a3024e8417c800d3bc2d64258783826d4dd1ecda2b25dceb3d418751
zad493a02280d567a5adac57cf1267907e0deb488fbd39cebc5a43a087fc4b4af64228e709f66c4
zfee8dc0884ea4649787cf1dcf65239faeb2f6d8a28e9f2522532a0ee0d6dd0e1c08a39e61af933
z010bdc0b723299e705bfbe0f0fcf70f95591b0bf85e9e30494dd6d0165ab40ac46756ee61fa7bb
z0faa6ff44368d3dbfb7db04759363a4163240a7595d4e7e1c1983d21520f2bff736d477a32b931
z386bed8bb3a4ab50bb113a246f1d2f4b74e18e37132f5be7bbb7219d5329412fcea67879d5bc9e
z1247eb6af02a817af9ba02fbff5bf2d952ced8157b227a50fe1e5037adc8956c0d659ecbeb7369
zb603d2bacef7f61c2f367684b4d13abb56fea2be2161323e76b8f4a08ebe235e725c92123449eb
zb39f8649e8221c8b9bcb4937598225245311cdb367000dc17307cb96aa12b98fe8a95a7d059828
z1587650175c1cd5380f0313040ea2556f5858b11218a72bb84cf4ce09761bb3e4cdaf12c1c71c6
z4b4153499d3b3e08ace38971f7079b55f4d01d4090826fd1d57094deacfa446589089895f5f5a9
zd37622a01c771e7bd3c99eaf28e169dd35203311dd145eff3cbf1c34339dbd663c136f942f68bc
zbcc0ccc3e0fe9a1ab9572d59d05a3695834bfa225d599cd7b675bf12e2b3224a35e5205174251f
zd70cdde7ff11719791a6760879b51fe06d30f045ee8a7f5847c102e51e474a1de6d0bf41fa3ee1
z277da6403ab3a74957956dc8fc68d32972b80645afebd74cca6557d9b9b9cd6edc5118a0902af7
z5c9bc6d25089c340e2abea983596f123ba6017b36ecdee564b4d57f3f46a953d586e8b363f40b9
z75bd6063081747b2f0a115ba28a21acc705d36d7592c16f1733aa95d1c0eedda5a0e3d978c56b7
z7c2d97ad554aca1cc28d41d9c1f61016f345e64cdb46e6338f07dda9da1b84015a1785d26e5546
z3fb217a4634b1df2e89270211a9e4e0cfe1eda263c2a4ecef1bd60fa110de704b068d70c05dcc6
z1d7f7a4fa5213aa925b3244fa48e3ea0a27a4969c75bdcc2e3cccbc0163ee5ffda5e9430590077
z23938c28687b905596ca3d278745234337e833c9bd1bf4ee790de71a2a3b5a1a34e69238248ccd
z2c55038eefc27d63774d0e48d90e3a3faba82557646d38abe5bd739b1018c98e8a8eb8176fc80b
zdeb90d76ba7e72a0aa8a14785eaac0e6482ce38eae062bac8f63f11571bc2bf1e4fe61e27440cd
z7865b4a6e2be99e180ef6d451a27aeb3305e6bd26c655ec7a79eabfbada5c5ea9c7d560edb08bd
z3c949402789191a86384a163ae21a9c4ec1ec12480fa925138fa7a12177c4a4305804c19dff2a0
zda99ef8eff98ee86e736876dafd88dc6b2ef28b9eb83f1bdc3c156634209bc4eebc73a645d9a3c
z67b1bc9d80a06b9a4f95f528c193921a154100955b99ecbdd03bea7746aef3a9255463cd1055bc
z40a130de13306101bf2c4edfa37be103a3ba7415be3119394ec5a3f0f16fe869d1ac475ab294f2
z234abf3ed4a627781757392a8a412a9a0f0938cf256e72ba4cd935c588b7eb1a20cb7af6f75f2c
z97fd5e72d72e49dd76977af66d4b0fbcf2eb9ed9079f437e26fdd1b4569197949ed8a315e443ca
z8bc158aac95761dbcd48f3e514d555ff0c31f1af4536159fe2a44da9687857711140e530250929
z60b3aa739fd74af0e38ffb473b3aff06b96af85f07fc9f51b636c7c25f13ab9ab570e52f3a94fa
z07c053a5fbcadd6f739ede068a59ddf8a42a087dd1300bf34bd27fd7f866346fe48a40e0aad0b4
z03c257f30706765916e3063d19fa43a5dfc61572931a687494416a63556f0c46a57bed91de189a
z6ec368ba4e7b6e907eedb65d2fae4f1b30962f37170fcbcc7e3aa752f50fa3f895db9aa990c6f4
z9cd7d16859a3ab7d4b23213c8c55afa9df8600377d9037926eff36e644ca59b42e1909e567e372
z0c16d8f4ad0d5548ccb2d433ab42b6b91fe1452bf74492b8c7ad644e70160b11214f66d5da1e7c
z51996833bbe0483814fa4d7890e3eb5307264e6fb8e4b3fdae9ebf94ee09a1e9c5fd163f9bd06d
za0266c5a39e73d7223ba83c553777b5b874b5bf657ff40e19d5031a04a6916381740ed868687f4
z5c9ca75524800ebb7d11527e23e16ed77973649f92dfa6fc1043006bf79d2a15520ec7abe3cc13
z129d70cf837561ac3340b3d6c7554c549cf49840cd39ca09f441559e2058ab7854320aef4c1985
z0129f03ad6e14e013803de8556bc58d60e675b92b1e1c1daec42233fc42c44faa4b62f8a206037
z9ae4e076526ac440c194082fa88ada6240d7785a0b9e878725c1cee68d38451eea77a099ce259d
z9611b3490081e05339ac3303fefc0a13a692571dea9963c2ea85f4cc23a6ff0ecebdaf8c289bbf
zf4fe239d0c27d3620e5ef5c38687df2ea7f4820e7a67acfc3ced8474dfe6e0b5e603ff4d21346f
z5186d814dab6ad59ee110c87c8ed5831e2bdf903a007d559960f3e0b7c3d6385c4beb9a33138d2
z88eaefc3617b092d1cedf9b0b35b3e67d5e7c339a9a6c3f31b550379d8cd60334c651902e93f42
zfebb1276551bac6e16fff7fc4317d4360ba2e3d27f7cdff3207a68a1fc6ecfff9be99611480037
z46f70e8a085cd4e7114444fc2775e583bcfd1cb7d0ebee260f9473341d56bd8c1c7191b1d13a9c
z8e04a181290723ff11030723a561919c2585591dea03b2d49d5bd6fdaf4739c141f5171c7c2390
z4cee081a47a7743a84dfcc49529208a3b2b2d0cb775bd75ed09435e50c8176ef26415b8efd9348
z206f547b777bd6e23f445c62c27c4519190de79816d19dfa8183b57a44998ae7b87d90d7f7785d
z6e31e02e15cd2fa92c159566c75a87f5edee4b87ada0ac657ae3eff3e75edc249d695c0442b789
z4e488acfe9904ece411f3d3090daa25616b1a93156d418d33b536821338bcb77378288b2256215
zcfbafbe44c66ff0e3d21d4ce720c14ef00d798c2ec1e02ece5bff5ed580f0fb2ae7435c29b38e0
z5ec945075c0e90e936ff80d522fe5ba766fddad7bef325a5a8c622e4bccb154e29a6f716c8012c
z5c0aa6abdc0627d1bd96340c66a12ce5812508b6a13f53e95e7c0902780ec302224eadc06dd999
z31211d5eefcd726279a09866c67b47c1fa4bb1a74399b990aaf1d8b2e7ecd87c9946522f2bc59a
z110d704beab9aa567d36e5feed327426bba4747b1aecf86d2309b73832424355fa137bd727c2bb
zd87680e1bebbb50d8257838d6a005468b44fc5f23e6f63674cfc98141b503764128dd4de24cb59
z1863c0ff208ac4e5671debdda33f5b7968ac36bf22802a9f288658484a8ed63c2f561f052f8fac
z1fe9beae5d19b476c31f25b65102cae7915eca96ea8161d49ef4015468a3c301bacd92e2a83639
zd8aa361968a24bb7592454724fff6df7b6d9b9188dec6ff2d09f359b4c1981ba15ee161bc1d8eb
zd45d884cb466a7c3cc78c934a2c08cdd2aa6c5ea1b87c6985d119ba964baf0f24d6aad7ff1c61e
z883d29c992d77de31904a65b2dc9a32345bfa61c066822b128486fac9a3d6cb1c14cfe1cee29eb
z1ac2a4bef3af9d42342291a6e80a8bc26f57c08adc84c62bdd794575705bc8911bd7ff899128d9
z8c6621c4bec9c22f7248f3229a36035eec21e084928c7902baaafe5ad24efdc8cb02473af2f826
z89b9312212a8ad3e7e1f196e8ab2fd69613403d70cd72bb57bc5b72599d5ad76587ea09708ca30
z83cf812e816830409995e7e39b79c1cbd78d47ea46c2faf1abdd1d31eafa89e67f7bb5fd2fe2d1
z4d8119f745dd4576ce62c956812d5e76b4f646306dee7e6ea1c32ad4f19a2ae09044654d0c5f11
zba8013602a830ffcb485646bf65dc48fb299b9e69768dc30463d01ca5b321ece4421f66e40d2f9
zb21b59406ff8ef1b1923ba2c432509ca6ca17abadc6828f1c4b71f70832095e259e368a04b8ed4
zf57dba1b1afbeed3072b2b3a2c270c16f1c90ae7bb78aae57f232980c80d2300b4b55f91e7c067
z3710f117682a43241ecbda1e76345e956dc39d04c07c9d789073d09295b5f6ee520ca8a133fc86
za0029a4242f15410695cae83aff9371d08b2b206c9a59f85f86cadd81472cfa24b54a39344ae3a
z85be71a5e7bbff4847dac2f2d3fd2787ab53b684893bc9abb5c19d3c7893d8a9f589222ade205c
z2aed55bc2608667ec91200026ea625fe21e648f947c41f79059e5d12b1eb77606a99c5c157642a
zec4ab7297d254a5dffef5659ea1f0ecc1fddc6e7189a764e9eb3b7ed8ae91fc8922594b3e5421b
z8b01f7d682ac58797f3c568deb3748cf4d3433b5edba7a7777948d38d033c30940a950a4ccb193
z0827a6d325e57cf8ac15b902e67496130cb0dc97698fde9668d0784dfe468157cee138b91b6fdd
za81935d91793302ea5fc208021e5e742301186c9458c6c9a4bb4d0a9783c5be8c87a9b01160415
zf6199e258d9ea134897493101c9b588a0f7a34b945bb56cca55f5b0133a881015888deeb1d5a93
ze13317c8cd6214c9bb9e7e7d8bac9f0fde958a6626a738e8d7ea68e3a401fc79f59c4b93572b5e
z9672ed0ef5b851bcf13355548bc04570bafa8117cfff98e59f751ce9e3cab17b17f2c8f74334e6
za78acef6bda8b90e489ccab2bb6c3dc9d63fdcfdafae37b4a5737cacb264670c96dcc9f417166e
z216ed3c0495dd2dfff41b99fc16b93e2907b6eab0df7e72454c14586a647989bdc0cadb4fc27eb
z3b294a37318fc6853c4e9d0621923b776a493343691ed6de81dc8849272e0bdc3ea9f8322ab72f
z1fe8a780eb36019222e3872cbde4a2fce53be3c9745b7452ede80c9fbe708b53a28c611cfbd350
zaef4dd7da02a960f28189e34ef0ac3745ebb35eff7b12a7442e165606e3a8d05d4b67ffc1e18b1
z3bacefd208422c329f3838fcc78cddb79e62b9b97a297e080285fb71ed1bacd70c6d031082d5d3
z342bde4bec82b82db5d4c7995664bd76f51c4066326fcd985b98adb38f3008bb7388bfe2ed1662
z3448ee711dc16c751ebbfc754c2df96376b053de68648a862090c4514555fb350a834faf94aba5
z346949dadebab7882c96c4684885e1b18f788a65685a3af9da4b5776007bd505762cce193d0977
z667622f9cf682d656d3c14641f83b01ade1b7cd21caedbad6b3969226dd954ea033467f94ddd40
z084755dbabfbd492eb14fb54979fe21450fb24b76cdcc23bf4ce1617d1b2ed130497f902b61177
z685192c9c177a04036d81200b33a078a21706be01533fb2a048eb0a5ec016c84f83f632e0e949f
z6bd40c0aa159f169f53c8ad300535d3e2e517a6625caf0ec584a01ed3094b7d1a2510e2fd35dde
zd672aff26882e2c61e2c1ec72e45578d84adb1f7ae4e509d51eb215787600e63ea78809c5d8b34
z398ea200d9acc221611ddd2555121d0dca34eecb6bbc9c450476497f712b82c383c821a5b2ba69
z0114e4ef6c10ca10ab726f47d1cf80b05e6a1df1e7e5940c587d5579a0598accadc2a5f7c4c084
z1f65aef26ec3b3937db8b700eb1aa110de0e0bd96839f6269d47818e3d184828484c1139d51c31
z21ebf8496b0770a6557431db21900128f5f3ca3d8463278a39b2340f72f5c893ed613c0c36fbc7
zbc98b139c7f8b50a95d5840c7957bbe09a2a23217e11dcfc3eae67d9a7d71aa26d1c095eca01fb
zfbeb79acc70723aee22712c1315cff2259dfda7caa02b3839da7b9255f5fcfb6d32ab3f922ef73
z4ddeecfbc6ad5d67b0a86ed7254250f2585188735b2d3fccfc3217d23a9cd29131926344856f7a
z06abab25e2f50aceb957414841fc30867e68634f8a57644cff80311ebf69fdf1c4fbb1be8c75be
z27da661ae58d7fe0a405e362103afa0b8988c768e7c69f3a34fa8808a34b801d4a38dead6185af
zefd3fd9d312505a9abcf165951113be03d25b2e923fbf23a24c88bbb161f65bd65205650cee936
z4770de31f08a7dc4903931eb269e9098cb437148201e9e2c08291de44a2deb8aee6c0fec695a33
zeae6a686709d85e0ce87058f35f2f9990af5bead9bd4acc9bf8d5fe3d28a32d77968c0e92bd13b
z78e472da7f014480afb770fa494c02fd26e2bb2259827e021f238fe06be2120c89a2c9a90ed0bd
z6e4e967f430b449dbaa9be1f57a1d06eec7f0c91cee2c9e23b20fb707c60f3e36ecd228a8db2d4
zdce0979636306a9a674b1afff1edd21c4b26f854b2911e08257163ec7de81874138b71bbf21ef2
z613bf9a7ee53c04bada3e3fe631cb090c0e5839328288003453a5080b29f219bf8e9c7b5ca1533
z39afcd846013ece9c60cfbc8e1b7116b119dee17b86744ba564d184b744d74f4a8d4adfbd53dc3
zd9ba65558e9622b0a23917026f6b16a490d8ececba988ee3d08b81c9f007c1fddf65c1e0fe68cf
zc1fe69b8dea458bbba98829d73fdd49189ed41a0bde9adcbec24451dfeb0664eb0688fe45e4c23
z511f3efa99d599e7f8886226c5076d963012adb74916af1fa392376d21834d4ebfde607fbaa773
z06e6d68fe59518b4ce6b301c4011a43897b6f70fe1cdb29719ac95c34575e0790600b6c251f237
z65eec50e205aa462bbb49b4bea7c4ce0af0365b5485fcba56486fbbbed6617dd0a82d58d6a90a8
ze26f2b7bc418f31a33c602b1f0cf68720afca5390ea4a7a6071e03b0d89eb8d12599fee8caf1df
zb8b7cb30d7b3fd5be6802d49a77bb040996160f42056fb0da1ce19112cce0003d401df45cef292
z58c86e1737165f9500b6ff9f806ebc79f268f64239c792dd1cb669ee4693fcb4fe3bddac311dd7
zdbba900081dfab1e6de35f32404ee54df4dbb91dc996086dad2df4dd268ab7daecf7094051232f
zffb9ebd7f9fc341e9a8679ff64a0240df73743595617ca4cbc31ccdec9b3fc54bb3e3855a7e8af
ze73134d7f10bf75e9ae538201edbe57fb40d04912b2dc6ff01f44f4f60e95c84b410242963a10b
z7e7a4e9a79b1f83e40adfa5d125ea72350c9705fd094de9c03ecd0114929c36d9403f51d99c2d0
z5357b418f5c7125f9659fcede585cecbef0c0e2f2b0db54f92c511181a384c106d36273a64d7b1
z821591ee8825767665393a4a5dd55146cb29db1a5afb14ed55e4821308d14dfba5247ac99b8d68
z5919d3948275b2900d915d64ccdcb1d5f7f38cbe84bcacd13cb99cba5a3a40d80ffb6fe21e2519
z70bdf62d8bc9c02b45ef51bb222eb1eed1df4b4ed2f0bda5208f1d764e9c1e9b8ade95ed151c2a
zc15646d556a41ad9763b09607952949992c4ee4991b7753982959699c21307094383de68cf266f
z7fc3a9dc42a8945cf0e4d0fa97b06ccadd3e13bd9b5239ad959add6f7717c7b409d6041b8a45d0
za570f0e572c260701f637814d1daa2e4df7f8756a79193e4aa2dd75e0686c231088d2feca64f97
zb1a0432f34a8610f93bcccf45670a161bd68e297397f8690b0e53439da1557a97a9be8db318076
zcacdb4cb6ed7df02d16807a85aaabe3e8a5c1e2500f7b2af160343a4b605052edd0da3a85a0b3a
z5439627a3afbfea335a115b931a3ff6db56a067811ed068baf16548676817cd04da13d6e6447b9
zc245a3e612b26825a4d27c08656150a393a4f301e836f5d6c1eb8acf279c53583db0946201960d
zaf7393d652eaeae034aa191ac78f370af876df3370784d901fa160bc995cec702013ee6508d0f5
zebb270d1b4254eb7324c6509366323455a19a898363f8b142d48a6cc2fe049bad51e296f7a7e11
z77ce6ad2c844c9bb6c0fed8943d47590a3158a8a62b9164c7e4d6628afefb9b906cba45a59eabb
z373453e662a7dc93b0bddfaf0110161e38b13ad680f4b576b5a3c1b28907fb75c6839fd8eaa613
zb3ad2d0a97ab7b043de0830729833fbd11c28442524b0a4f9c2e3ece1b31ccea1fccf82be67474
za992cdbf3c9b60e68ba6c9242e8c65f5589c7e3c158a8fa312de8101dfa5807438ede7e2588085
zbce7793c4f93a783fa4f821648dd929f1bd0de2f1969c6e3b7e8294bd5322362f388ca35fe823a
z6733ebf852db9b5033be5ab9da474711cf3f5065cae2695bfe2024f150d7dc299ed5c2cd790375
z08f9b448e233236351b29d679cd016ceebb798dc117fc25e07210a1018155f97f74990ff6a2590
zc47082638bcb8eb0e81a1f0aa889a83798b78d0b062157204fdc8df113cdf5dfe32f87add23c53
z37dc4882225a3ef8f5e2462e4003e57179aaa2b6d5e9bd299adaf655288612d817f122fd4bde1d
z99bf18bbb217e8110ceb2e07e9b6abee60c051fd8dca04301eba9fd1ad3ec00398ecff07b9bae2
zb711f8ad89070486677bae8ee8e4a00d861ce0cdfbd48a9820f0663e34323ce98e37af226fb4f7
z5b3d32006f0eff6ef61c071aeb5e401e12e3287920c2f51f5583f27d4e9b5e0098494308c985dc
zc38797cbaca304bebb86747dcfed7ad4cafc2ee1c21c14ef993eb6bed050c446b80c6525481555
z28bad873103d05fd62c74b4b9c605447daaeb6584c1327deab2d8bc782852089a0db9e0164fbd9
zb1f0f244f2c59f14432c9c994b7e8c0873815a4682cf3352b5b87ba7b1998264b112ba25f9389b
zea8f85cd71df0986675308d3b7665c1e1407f9a0e17e682934d0f05d80a9a45f96d0f892d7b82d
zbff92e23b22ed2187603961aecba4440fc3a751ff4396f5638f7934f27f2261d681d846d96916d
zb935d642a1500c501a5813dbb801bbee266b50894954ab1b9a0e00996f3cac45459d5e3c2abe81
zea6c482deba7e9874bbf0fcc206bd4fb0d969358fb7cafbb1b306db28b26ad34a5caeaba1c34ab
zbb7575edb633465f5a96e1873b4400dba8c0af3503608a33ba3604faeae5189576a2987502b520
zed7277cbfaebca2352aa2da589b0dcc46baa05d487ea573ca109cba280162c41bedc1ca256e55e
z7dda3fa4c847849211accf3db2e344255a73858361760979eaef8e46b018e507729009541636cb
z67e401b022207646523de5b65c6c08746a117d544d8367883d2a823afc1f04eaac23677a286b86
z0a7b60218a68f500155ae13e1201421cbd8167cfce5a5490398fa6185e709ff7854d4d17a24497
z8e813e8d1d549e1e9ae0d9272b7660cfc5d7e302c11301b204e4fcb960fb22f7fc42c8665285fc
z46a9b3fda958bcb3604279f8de8f1de0c90294fd4d9c0d7bb08f8f8d41ff134d10e8ca014688cd
z656f29b8c6f110110c6d207795d00cc2e37bea48fcd1d722d35e156555c350d29a5fc33ec5c4eb
z00fc34dbc1f84661fc7a7671830c46662aaeb3ed5e85fd10e50dbe8d9ff7b1d594284fab9511f1
zdd7e737e1ddc910b78399a2c054d228d35799a955f3e78b1eac42e6463292c478b87b8bed4bf38
za52bb4ba3ded650e69b9698f45e71a6e5f5f3861ddaf561b7cd0eebc2b98134b488506b15c7d99
za47b5c1ddc153e28181c26cfb4aecf743b4d5a9fd31766551098fae5e4a843d7bd810f2b62428e
zc348629b108dd93c59b5f1a7708c8f13573e0f62cf067c7e649d06a2189e83abcc5f0f57724f59
zb2636c99b6005c159745e7f8f8bfa62a5ae9fe09cb96ee959de446fe1eb157e6f0b460d0e8154d
z88f0a714127f81631f9fb03163b52aadd39335369291018c961d9112c34676956b2706a6391ad2
z395bbfa6895d21aa026b322c70ee46e45a3060b3b6a2dcd6276fbbb63dde738106a71b0e05c959
z1d69755d143c8a4c72d889419e195dff4a19b3f67fc3fd26aebfc0c5f4c3e3dd3fb5a33b8743eb
z9f448aec7f26a8000216475abcbad767fafdc099dd4d3e3b80de1efef1a81529e9859a9b94424d
z440489c011a3a84e489ae776b555ec77e84b5f0525db175963401f82ba55be3cd687e2f04cc905
zc8eab19db47486445eec0321a6d7a5070cb42e8b884334786878385c6f4e4c0667d0085eeb17d0
za50716ccf04626ef290c4b6acdf01603a04377fa34aa749f090131da79983eb5a0029bf31b4f0a
z6ec05720a07340da9b947ffef8700c682e3f4e48c3b69df28e9dbbc14dd78ce1509d6aa5f6552a
z2f592aaf67da1b3111c261d607624a5aebb05c41b9f224517209378d720ae1ffcda58a43a3402b
z29b705833d8be012a1a0bf2ed3b0a31d356ef38b154bc511f956eb037ce878b5fad8f44773ff21
z96bb39e1805ef43ed9674d06fa68ac02169e73163a2fab06f217145aa075b53275bed266121ffd
z7602da3cb76767d93e6121f12d65337811cbc14b257e8e02c8c13b874fda88ca74f030692c1006
zcf36a2ae4bcc95a5ee1cfadd660993293dea2d1be436293548bd72c6ffe78770d6cda6b67eb9d4
z70059741d66767875ed8189b9ab1e4959191f4625c19e403bfb3d0c6db187914e323c01883d364
zc97e5ae0d4d7a5a8cfde7760ea7c94cc6ab91f76dccb6055940e8ec5bc4b28e97dc5195964703d
zd8e48d48ef2d83fc12ed9d2767ca060e0e939acb6a2e2d54c44916d8fa3fa4cd63400abc46b86e
ze72b99cce940a56424c3a0684b10cb806977b69b818caedf218644772eb9370ff983ff05e1e8a6
z0d2c2da2f01e397fd7190f1b19c8fff8d99fa50011da340e33a0538deb52347652dbf8598f51d3
za2e6251a85eaee41dbb16d0847365df1c70f371c102422f5713c0bd55b226409e052511684918c
zcac1e57c3071ca5754c2e9f5a1bc985de7f909c72baa95c8caace0924a16ccfaf07b1b608f3e89
z6d58ad8c182ff9b780bf7a15e9c2a96629fd31590d06d13f09ae5c30e8e55babb3c35e6c8c2f55
z0b5f9d92f31480a966164b80a8aa997878c39cc61ae5842f34e3c93ac3f5849eff5b6cceb607fd
z25145e3c7c295140b5ffa2a476ffda48bda0615fb467c78d1589905473a238b5ce4a2b6b51f5ee
z6952ac1fd57ce020d6b972bbb1ed97e4f7ce337d4da74d0c5e853711ecf12d1ed03183ae26ab2f
za1a0bfe4ebba8803fb3dad9f186f38d0020735726c14d3e885d0d9dd925ea7b994757b3fd960ee
z7994d0e825f057c31f0e5e13d3ff0113223e865881dea79dc68852372f279b071f34f2b502f7c0
zc3bbe6737e3d1653199a6971b21f040cb1e936fce9849664743f76d988e7030cafd11dbcfe6939
zdaa110369e6070906b204fd5f5563d545b33d90dfdc6d650ba3aba432a2fe9ab3b4485da821ab2
z612275ab72601e0167ce0e7b61195bb447621977ec1d873ad812adf37645f3defe45d4f3867bdd
z137a448450602493c974b989c97a42b7ebb0de3d189283ba810273767541dc7c3777c77fbc28cc
z2bb4c2ef31d54ed6082b2d4bd80b6c3bcf233632759845d0d025441d3d82ce9113876f654e778c
za7e9c2042f49d0a84781f00b4bd52825d351ca6cc2d22ed68aae0c8d856a9b33fe77d2f1cd1c9d
z4b9b6d627521ff458706be74f8d92c42283b20e7a74eaeb22946dc5d5c9c0853337dc46846fafd
z580052e7378eaa89a66564d4b8dfbaa989b54a78bea1853bce43964c7a48830216ae0d46f829a0
z557e1392aa38891f3d70f696f2b7050397e2c140885196a544ca1d976fdec08295152c8cd8453c
zb6db2c798adcbab59424b59a072052f463d334eecce623efdefb42b6526a4fb214cef0c2e9157c
z586a062feebc4d97b90d43febb8fde28f518a5e17feb67bc98e6330d8223ce71d1623c6876868f
z3753ea44c27214f7467498bb53b788bd30379743e4075e6b9624d67f628244066d3de943c0c828
za1f4c7acdbce8d2e23f79dec6b13bcd3cdb254b0e541e2b0b16d60433d5e4c66e73a0dc629145e
zcc1c218bbad7f25e95bad9697b6769fb7c7194e7af70987a2c221108b85ded6d50cab4b03b2229
z243555185dd9f006fadb3e91d65c16c51f12e1e2b2d09e0c8d80b4652f987633a2c0a65caf6a64
z50f691079b6e76d578224847a9454028062e173fd30af4a4aed0e3dab4f8027088217c12bf29df
z5a3a4c38d97cbd2703be21ab9e537915cf39d79dd4d642b871264ac16524ca9ea61b5e57c32f63
z29a1f2b849bdc48d5ccbf06705a1cc5efd040c5e2e4f3e627dc294e20b90f4d552000ba9838ec4
zf5e370d8a26c80ea12e151a1f7d997c71fce8edba5bcd43a847a2838826a272ed870038a7fc9e4
z22502cfe7bbfd4dc953ee9e890fa6b19a131dd7b2986fda320e81212c2de198649b0be0bac5460
z359ef405ca24cdfad6d2c6d30713f7405302d134ae62eaf100a785d7bcf30d7f7a4573f19a787e
zb2a3b5b1e918820598c45e6ee62c81566a7c0e9e481b0c55e8cddd5916eef4eac4481e04e604f7
z66b3cd17c90f6ede90825778b22421ebc5e2cf1fb733b56215379282ccc2d182b8644581fc24e9
zce3773d400c0f04f2f4000c542efe7407b169ffbb4aedc43af80711c45d8c13b2e0f4df116879f
z56f1368fb2f569f171f0df8c21f86849e87c0b9900f0b85f669150cb6cb3a8e5cd4cb233bc5450
z4fa2276376a5de80f4ca713c0b4434d4be07ce30aebfae37e23d643c865361e142e86e7d23a9bb
z0654fa8dd91fa1cf5c43ee0dec8bdaaafdb991e902a7d94f828687c28a307cce37167cfece1443
z42371f6340faa1b37568e9c2c7a4620498c79747d007f0907ef389d02cbeb9216e8423f3aaff26
z154adedb79b498e249524cadd3f8793ca51fe3a21520db69152cb46f45527b6cac861496a8705f
z8229404fcdd1ceb016c1fb0fc61d828e2928f7eb903be54c46e931595c3b0fe5a108a9c03b2480
za36e123f93c322c3687b24523f635f601adbfe715c098f83abb15eb3803b421b7719931df5529a
zab9ea730b0208372bea80909ec201f1092b19ee66cfc6aeb41e53b798d88aeb9ddd70f8acc3452
zbe1dcf1d29bb09668a8e2cc16e2dad4c548014fe1175e856b0466fb2c6ef1105689be4fc9249e3
z77f0292319c5d9b9bb4b53ed4de7e65a3a90106e17bff6e2d37fefd5836d9a6261dfc6b12a9175
zf6399f843543a916318a535f24f5b0df9af10d5044ccd4102faf91ca8d1f4816c140c7a84c35c8
zabb3d9fed7db13e4ccdbd6f2f80b64463906d24de56f1ac91f0a42460761b270f928db34ebb22a
z2045d695f0ac591dfb922252fbeffd4d7fe10b5ef6fb6e530e8b714b421dded595fbe64b15f8a3
zf2340c8ae2600fafb5acc43065f60daff9b2e8ff310f2e6567628e24166eed80bedbe1e03636fb
z98bbd6b97179f06feb51a2387ac7bb782d201ec69214658d4e85adf448486686ce292d1cd7c7ac
zbfbfbd8736ebcd0828ca99a175dc25fc7a59e5f7fa9e700e506618bf07c6d1d5d102bc1f4c747a
z9d576671d74eedb28f37059ead43af4783753699ae091c6939696b22992d7b2489d59085c8ec13
z6a1f029ff65b22dfe622d9e233ed98430fca8455c544b79f1043041ef36583718b64b91a71e216
ze4d79b491803c432af53d3e49fa76bc699be7ca7e8be075db14d262c9f52df78a0e1d10bb82200
z45987c91ebf01d6405c5bb50bda328951623c8294937dcd083ac6fa4936c7090b93aac94329a6d
z0b964766133eecc8f0080334557cc34983ce04b6c453c90b047b02f5208782d58b74fd2cdda059
zbfe8c3ed921c071e98056ef156d5a2a6212ebdc4700646cef1c7b05ad63ea4b43d76a6601ceb01
zac19ca5533527d03a4138058def059bbe57462339d5019d6732e33618b68e6ba829143a93662c3
z38190114f9da322256a0160a80fdf31825b24c0946cfd48f14f17aa2cad589dfa3fd107c15890a
z81aa089af7fa381aa62d035565bfc07eca52c392527aa3ee263b7af9f1dcec14f87a9ce00a7f1a
zefb076127ec94dca5808704544ebc2c3b7b4c07ba367108aba3376db76b09e6a892a44ee5d16d2
z05d00264296bf01f05d4d0015875682122fe5f3b6e10b9f2577cace2abf1b2fc18bec811533c76
z3d1fc98471584738f4f9ed871537f361afea5983f72e6567a9028e46ae341851e41076f47532ce
z354941da510e4a08aeebabb3f90c9cb417c3034090f2b284d4de26cae11b6df521fafb1b4d2d7d
z9f7c02e31a4dc5710440027b5cf3d50d140f516cc081dfcc5699dab850283bb6284122dbb2f701
z285c421a29fdcf4dbbe525952377564e27b92a25c9893b667eeb6611d84c7dc18d286bae36dfaa
z3251ff2f4a6dde4089e2769cd924e1eca6a487292da6649e78c2ac22b46c8ebea23948d932beb5
z2819754d402be412bbc82ed1373f890c354b2bef43f4f78d2373779a957b8f006f2e56ad2f263d
z0b4bff615e035808a093ffb2e1a633e96e6f36bdb0f0d6038a044ee0c68b338f54751fc1490982
zca9f57ed7e0813c809e25f525571f638c7b082cd88ac0730973c228e115eadc18c800f2ca2a705
zabb403b816cbc3239b8c5fd44fd7916f628a1fd69850a2e1413b45582681bcbcd9b7e8126fed20
ze10dc992848583af13ba838e7eea81ad8791e0207972d7d8776586bfdd3b9459042456544acae3
z8acacd400ff62ab2d763c040133a0b555ce516590fab730dafd80f5fab258506e2c649e6426c85
zf8034b36eac3be6d1d13d2a590e27e71722d446134a3a99a30db78f6496d494ca3ef5662265c93
z041403d5d1d305459f14a0b9a1c588c88eccb153e2b78670626baf2cc83915971ac30069a67d9c
z155f672939fab1bde0bcfc0b05303591caa5219de3ad9bf5b46d09878f34d14834b3b9a3fb5fa8
zd7320b5966520ff47a1b1eab4af44fd4f306778430fe24bf779a20f5cf355b8ecc40be5b8993f3
z27b07fa647daa4242c8e1157bcfe94ed7f8933a2dfa9463a3f2a1fb13bb6507ba8ec67bea9937c
z95049d3855de8717878a8ed4f2e320587a5449087ecbdbc06a551451dff9103d25b02d711378c5
zc4ceb15f89654e4c4ff23cd45a2085098b42dcc011b73d2aed948db9808ace08c58567fe159ea1
zb44bc49bbc4054b647592621433a1b00586c6500ab417c4e47b31938d6df160dff2fca03d8a09a
z23a3321c86d40ab0ac5fae0d69cba525c437ac554bdb6d37973df15de191db69e89fbb64bcb9c3
z4ce57f0b69a124eda093ab57bb4df6ad4431694f5aa3047b3c2de780c2c305b2d6fcf9f2a8afc5
z82bd477aa12a39907ab55622722a3b92a7561bb760a5e80a9193ab7f00213d666a6a3c61610b49
z40cb21bb2cf55c4d3b377592d4020049cf0adfba19beed0bcc68cb0b9bd3e5f5dd4334fc91fcc5
zeb5194943f4a3d5d8efe5233d5bb7bdc66cbf6988ed14ee0e586cb9297716335883e56f7606260
z69d1bb03224539512491d52bb15749751cf5e5c4143d240f7a512fc29de95b3acd96c4ebb31a7e
z219cc4f93a76134f439f7ad78966b2d7cb52b8b40a5c71814252225dadc88cc4b67d1540118972
zf5abd73e481666ac6af152d8c27b00742b0aa5a3a2c6061e264a93c18cb728301ffe50d5e0ff3a
z7f9265602cb83e0593a5caddf61f51603d8688743e72c82cafe36547da13bdaec0f98667d6f65c
zd13ee9ba66d6086b290e2c254e8cd07dc67857c72da154c8ec72f43fcf424f851a6bf6d3202a19
zea6994d4c15f790ca9e07418bf88b40783aff450f45a8f1988146aee38fe1ed348403aac7f7f38
z52fd4c38c2d6b410c8176d7f5ea5f975be79841e448a6aad249d224d97130fc631a4627962b820
z9cec30740a47720e2ee8f70ca732b63f439deb2a8414b411697decc086968fcc18e6836d71cd70
z2860e0164620a6ddeaccd44ddf451428c1c5ddc5aae3e54a2409f220a968705c355886741ea055
z388c2013ede7c86f6bd19de6919d72e19c9a17f50fe5288bf6eadbd899e4ad41ff4888d2abc0e3
z18d2ce3c127b3c2b0d24930bd5116946a576b2b5f9d5c6af531b271ca0cb84e37953c1610134e7
z7f9f5ed040c09f8ca3d2b64541e67f9b94fc73c45626991c19bee1fd957817afd0e9c1ec1ed2b0
zfa1bea741aa20579bd66d4a02d25b1caa70824d05ae95bb6d192b7216d077a05d0305687459f15
zb729d5e372385ef0ac44be5b526d2450545015b32040fcf79124a6deac4d31c9116e922d9f912f
z22ec879c553677d20d3e6411d9acb45a5d5234394b0833a0dc16abcdda0463604d3cf9e9bce78d
z3bf99f00e39abce1b6906c8b5c4222aa6ddd2699ddb9766df36df5eb09bebc47273a21d00b9e2b
z1d4cd2b887f0c46aafde9086c74963eb4ab2e34da0e0e85165959a0d3a97515455b3ce8819057f
z7d0d4987d8464cfbe7f5d3b27544559170cfff10e4320ac3fb0e26bf78d7f08c8920b5a62d883e
z4d0da518a3f56057a1e251f4ed484bac785f1f0778cb727ccad4afb2205b4bcb855d83ab9ab991
za7fa95733523041a13db9517d6af3cef5ec769295e672cfdc4d0d525c94f08e24e463d2e1d8265
z7d21abd665cec8e72e7f4c213970e969a9c25282a3922d26e6e89cfe9eb13457612281e976b40b
z5081bbc67c5cd7a80a906d696d9529a73e219d864069631df32339f4ab9469d5428f8eebee2789
zd39c62dadf57bd4744057944df7bc1eed7312cb49e044b8220bc2167f9a00d445f6389dcf840e1
zdb0cac1088a4ebacecdb16b873e63cc744dc9f6b18a422a6b353b5cb9a05239d2b9acf1d53d388
z5ccd26c572b6a8821cb23d25c5429850420cea1d593f1b0e00a8e41aac71f12be572fb74677f3a
z41d61155073ddb62e78edd2942dcf631c4487152c2a7f4a72a2c11a1f7f6e7ad301051fdf828d9
z0124d027469ad488ac72cea3deec5f6811dd88f7c94f7998d98b55e113fba8145f22e75a6650db
zd1aadcc16a4716ea0ef2616781b964be5a0ab43c6d0516239705704b7014ec4af936a3e27ff02d
zbbdbe3adea757cb461e3026c571157aa78413b09c33edddc106de117abb58b09df048e22c1eb4e
z2dbad96e48f34fe6a9f5c16b4398b5ed08dc1dbfc144dfe7d6286c7233b69d37d54dceb1dbaf94
z007a7354721817d71d1b60af94422a8c193d8a70b13d7a4cff5daeca6962fa073214827bb1bd01
zc76dbb957a4bce919300463392ae971de84769045e730c4497d40601da1861896bf6bce6c90e94
zbb25f006e50ddab0504ec9c156dda40a64e0defb26be97404b5bea63c5c0650bd6f32333536798
z5b45dc333829c1d32cfb0dff4bde71fa08d74ccece00ed4469ae76b6b9cfc939d032dd29bd2441
z778d4d15ab6665ec5fbf1262c669e4610dcb3d5893abae8bb26b8dda393ee1cd833829c5abf4f5
zb757d46c85aeab5bfb9f89a539414e533e93736f34d99caa29cb0145eff9efef58a9db2cb2888d
ze554cc801f6333fe7e9e580c556eeec45094f0a3fecab460c85bea58d9b832ec50d79dc8be4799
z8ecaa63b8e294922f824209cb497d4daa42d28439083dfd194e8e2b0b5700dcd38a628ef4a601a
z6c20fb0fc50decdeb2207edf2c5b0a48647788350c98465df16500f5df0c9cc7ebadfab4a62721
zf64f89a26d1059cee95612dae70a7ef4d098c13e3b42e8733f1bc007548f38c268a1e681c9e881
zce66b237bfe7b30d031fc78491b7bdd9dc176b1ae9dc46a689e1673f9aa93d4379121edcc9e935
z88c62626eb2ac9f2b4b48f91a71fa932eb41ddb22f6313ea4021418f2655d460d6df3edda2d667
zf334362d472fb434596cc469e273c44da7a8fde04c2993a317700c4d52afed1a1c5d001b77ce1b
z1a09897666ab8ac4aab3a081fd94d2f76e39a6be22a23fea6652dc7e46913f94689fcd83463432
za1dc30f7cb6f7480d8c86856448f9c816ce481a318be27926f5322d2aff53d76c259aac37fb9c9
zc70145141274c0aacee219430760e732f5714d91b533716c25b7ee0a57ac220a80ff926d43664a
z43b5e822a042bc5046b20f392b5c3becd478f2af0a13bbd87f8ab36ab31c4d96e86b919d3427f0
ze675b93629e19889af7f2ded8959aca3585cb9deb1c342a56dd4266056c65f60563d6ad57517a2
z94194d090ca03def12cdcdf2930e3c4cb4e497d2ea794c6247b85de6024ead4d12bfce0e80f242
z9aebfc74e61c13bf3126dfa52072e8f894a78af4f2be59673d979a1619fde317c3383f996599ad
z71332c0f0ee24184a0bcbefcfd09e0eebc53a06c304a03384996c1442ae70536b9b9e7b3db7806
z2b29c388c808fd8d668e3e728cc9680f5a2894c87ded7bc83e25c3171179963b28c49aafbe9064
zaf80984d291933c964a9575694e15bd7ea57cf6ffd667fdc3cf77f94f52b3649067099f1e46003
z36d6d58431ba9f5d71b96b90bfd13262055b6ba3bdf07ffcd21e282e8c0c2c1bce87fdbc5637bc
z9d7240dc3717ec7d0f76a4bb0d85c8d78825e649de50845362c3cd64c06b9892f83c901f1a0b1e
z68c444f4ef02b78923365f11df84e6b99a7485580bb5cc98cf11975ef12bf1a83826cb5eb2a558
z82700cd641479f1087a3680ef3e2ca0500205afaed1d3f2ab46e3a7fc14f581cb97273b4e9202f
z130a50286a76a345ed452e2161c6565adb8591ccf57fde017612c8aecc0644a547633c217b5d7e
zd7d36115db886a715a20862405dea9caa528f47ba077e91ff208594469a537d582285c12561b24
ze0e8274ecb8c10765f9ceef59269bcae2922fe07c7f9d16e9e8159094b15f9a446cf54a6cee4be
zac1ee7411721362c1a27497f4425eebb98def2b544b51978e7fddd0bc6bed81a8dc4d9015e01d8
zfca5d34503ed4dabc985906e22abe451410c99d32dff2a1e81730bd468a196f316d7030940c870
zff1fd7b00b987953cf34a6c8778490e52ab37e8e195ba39004d3211d4230182f7ab09cf851ee32
z42ddff279dd3f645bf5d1825a77af80e49218b2e9699a488b36ec2bb1e41e1c7f77934b45ffbf9
z3971718520db59a54b5a69f7e241404d175cd02a231ad5b9447e2908690940b420df9e50a5db0f
z0a1caf9af90cb035e762c170a7b7a90ac4060414dd7d4a3edc1f11054ff5dea40a1830d06065fd
ze48b6ad2403bd934b00a8710b6f2fd7ef7e2f0df483fd2f2ed314a57c13232cdf0976ba8d5d4eb
z04eea806d575e7e62ec1179b34c61a7155c2c8b8bffa54c2ca172e5e839f5d188df61385db947e
z7efb09a58aa151f41a9055792f0cbf9ecb3b360b3d147f6ab0f1ea33c79ea8e8d501b241ec9e6c
z32d8f7a4eee0ec5ae91ac41e0687dd3b0bd3b755bc87ff6e5c7fe8fa9906a0c682db0c457d46e1
z81f31068ef1bee6d0b35fcb1728fb255de825e41ba35ceac5fd309736ef395f230c83ba8cb4e4e
z8cede0d80dc45f8e581b4a9ed425534ef0d0da9d3f1145a8366f8cf16d7e0eec420cbd14077b3d
zfba97ba8a60fb4bd9d800cbd4f1478d4fd4019e7700f0448b9d8ecf66cb630c3af127dcd13f975
zed235529d225a30a4d60957f754def34d2408f10e1b932304cf9c52165be580104a1b09672414c
ze05158cec097be1c2157be7074811e2c92e99b89573d490b527423b26e75221f23951d0287db64
z150bbfbb5c08839c87df4435a7de82d837279457989339262a35542672df268b9797a1ba0239c8
zd61872334358a6802c681dfc1c1ad4cac0a70b0881a11b1ece2bd671a3d4576ede8f655aa40447
zf7c976e7ed437eab55bf4138eccc18199d567a84216f5527d1a68765628288877ce02f2c1d8dad
zef4740c2af0084f35c39fb41601d426dcf354d624581bac68686121bdc435f10b3da500a298a1a
z48cce2277288b4a6959cc488ebfce8024aaeb1bd4b37315b5ca0d67c00f569704f6ce6f40a6031
zabef9d9c0c36989c9ad265ad1cd0c809e854e93cb0cad404226ce005ae75b20730463b159746a6
z4db0f6b738c68c0656a43a65963eb5b3c92936fcb39a48fbe2cb051ea2a9bc70f4f36ba8fe787e
z6fac0b5fb4f4699e3ab5d689ffd97bf76d3dfb6da6a7cb1358c809acbde61d19e74a77ab7ee69a
z819e7664f4bcc7d586bb7c1f75df2a7bccdb2360e9387139d82862c0e5e6d8624e454541675cf0
z922582fc98d94c7d8451a86e2387c5bcb83bc1206e82976a5cd3c20bf3e389692ff3fd9d21dbe7
ze31b3549e51362d43933ca0e8c9102ed4d708667d5e7db3b2c1322f06226980a1a66dc8902cd99
z5334972b6a6b54ec887724a9bbc758b11b11c50d774e58013694a62789c47d136bf427dea6dc5f
z88feac29e8a8751789ee9853cee8e7edea8eaaba1116e429d66b4227831aaa1b32c50c3d355714
za344ddbc87b9a3cec409bf5f1c2faaecbd9eb43d8dfd838e7fefa2e09c252a7e8b1c6f0984f894
ze76b14bd868f25d733af9e3a1e8c9b9d6a51ed3cd2746fe72b7f8852b903935db2e9f7e5be0f9b
z20de7273ae8927207940b960951675fdcfd73e70fc0925cc960d8c793a450774ca68ca7b738ffa
zfe362226cbfe579e324de86482087492aea49a0478012bf9bd41502dc0d63014f4d557c0b3d088
zf22c6a052c003517a39e731934cc870789c338d48a01f7669d6c71bdcead74e0d0f4ba7aefc569
z0c0d855c92842a1408fd8d82224d91f12a79f10ca3c3221a6daf20fccdbbf4c81baf3aa266f631
z4605ea42f4793d06053175ebc1b57533aa0fcb15817b3f114bc87ecb623b1500325b4523d7ec07
z19f083b0c4ce8898323710d70adfc95ed0931fdf65f0d6ae2eca68abed661c32546d4b0bc54a70
z1e2cb35c9457e7eca49500bcc72596e4ab5877e4d68488548c395ed40629b539bbf8a98d5cce2c
z20c624d1226e845f3dce35e0fba18fd347926aa83b7527021957fa37759ad5492c50cf9abeb1a7
za9f461d7d72a6d2b1ab8f2f80ba502347cf1e2aaf3a4bf75f070ff584b3bc11ed693d905db3b38
z63bc27fc376ddaa434a6efc6a078f46ac260a68b0f2d3fea98b0fead9212712ff655f75d592cbf
z1b49a1a5b94147413c9a815e350441dc4b3625bda252a87851c8c5a9c735a41ef29cbaef43f457
zab34cb4539ef455755e47bb0abdd11cca195d7f2de52545b6bc43c260282ac2223ed62c983d9da
z64c89c87bd6ee73796d64d1d83c03a91abd181aeeef9b3c1b0bcc34b46c2bbf63ada700be61c2a
zc95d2c279e212b19000766b4af40b5cab5f804fd2a7044376061c86ac23a394fa3e273b5b87d7e
zb231f7aa8912998668dbbfc88c002d400673b97995e547c487475cd8b6fe9900559e29224b9607
z38d3e147db2c4a3cd0fe32306bb7f493ed133730d6e2537f06e8023e3e20f57432745836a69573
z1994c55c2cb17294c9b0a4bb310f6aa6399b33e34900e5be99531c50fba730bdaf782f0dcdc874
zaf2099c2dbd1b69bbf951595dcb742f3ebeb1ebe9b2e20c2a19650982bce246d59af172a9d1cf2
z331b9f86e4ebb96e5f48a030750d7a4a98d2d1fd0b93b6258bca7c34f6e7a96026bd0f319001a2
z20962b7b698ce2503daba929ec86d8140d79694235c0fd9ffa1704ebe171f580a13dd544401a49
zb00b617074be7b24f781e00d7614896e1e2dd9326ee353be0177eacd0d8dcf37a17290fe2479b3
z1d997cfc19ea11d41c04a1efb3279b877f6c214cfddf87b458edfe232c5eaeaeccfdbda4adfce1
z61afdd580f46de1a44554be47679a88c041e66674d6aee613f4246be63b3d742348254087b77ac
zf89e05fa7cb1df1f798578cb0bca669a88f84c60d4fa4808fa5cdaae54e219162cbafd9afc9f43
z43109123890f07115c5d365ddf820206a9a03a2e8c50dd6f2fd757887a81d9c353f2778a2cccba
ze638394d0eff8a75e04c36c642dc48afcd59816ad7f756a07b299bfdd89d66111810d263afb469
z4cb9d5aa4a8aed7e7c49f371cea38523a99201d813695c9c40082c4bd3f15e20f7244d06eda1c5
z1d754eec3af5ea010bc3aad55da4ac63ae74a5275ff234dcb090b5f6f7a9b0fd8ee46a099239c7
z915a0b8f7286f274a8dca0982c146d601e64bbd5107c28f3da87584b6c1b39094be5ea628c9cb5
zaa7c85e5b11cc3b834f83ed8926712bfd59614550b2c97df09c58018fcc6c19641900d3783cff4
ze01db559897f97635178c587940a3dc09fed35ee162a63a310a1ff6bbd150fdf86c963f8d5ead2
z4c75b2ada613e33d6cfb498fc68ee116cb885d86a7839b8b87457d18f9aacd11565e5b3e1cf538
zd6adc5adb1929e6c505f3338cc97122be3dedef31330fc79a0d15180e41f1583ce8dc3979d2c38
z6a79eb6ceb3dd98527a704b853361b3e86d681810a891d4118d68d6137980f89d43400668ab716
zf696d2a792d22cda23f87ebc96f3ee426503b50338940ce64247e09abf5a3ef7a020e57a7370ee
ze39902a4a7429c0cb05797703e63283f9a2b85e71d8e154c6c6eeda3ac169de1aa1860facf2a1d
z7d5dc2e5ceb2f393608a1a6015ed133466ab48e113269d6b18dcc238abaf3ef99285e424de77be
z900719f6080718d1740847b60f31a0c9554a6f075ec6cd878fefcbba39e18ba07ede6d972118a4
zdeda917a8091c9e45bc10221fee2bf9d4c81a57def6ed5126d32f62b072ef01adc473cd41bf732
z89176f29072af6e8ef3e4571455506719b0d6997b08f9d14984e7351fe1925d420279da201d1d6
zeafdb95de535cf15e1ac43d8318af3d9d880d14abf421e946e8e1550d653724671cd684d6ec458
z71db52812b8a1ef94549d81eb08daa300331ee02ed0c21bcee11bf131cc4d65d10b74069a4adf9
z593bd59363af620aaafe8dd1f3127e5da7c2f2a02528b6eb269387f369a1b57f1931d99e9ac994
z135e24284f8a6bac5c2d2e303560ef1231f4841864aa161ed29c49aa78f8b19d9d5635f07c38ea
zc199d9c83c0dc37cda464f9c9a235d9942ee9702868e835414115ebe46f469e7333d35c8f87e90
z41f28be1b3acf6247272cd72ad5c9f57f570fb8141d9608eb3804d0f5a3a7e7a14c8d0d1378ba7
z961bf2331f1263ecd63d4a11c758f8fa90f68517c4586872897f3c5eb8b631c1829ea5c0d92a46
z627aa0512095e6a19a592027a36e3c3d07093097917687425d09902da43a45c100693e18806f57
z8770e76f7df122a17673da6fa2fdc930158bc6013e29fb9efade8e2886b8b1546eb800f1ddbc65
z959c718f6a21a2bbe3b96b16ba729557e733a327a06d6db4a2c35489dad4627b0576e466778255
za281cfece26837d8d54726f59e5b5cd34f04e87581a33019561161275e6cb1d1d296162a6509c2
z8fc6d1b8bf8ac2638394c73f504e10cd93cf35dbeccd1e5f0d51f27a6277e29506124a6123fe03
z69d40616cbb42ff7b5d17da3ae8fc22a7e957bb85469efb296da08dbf99799308b53c64f76a5d2
z12db9f5e669764bf849d4d58861c47ff5b563f0450cf807dab0629e0bce5478a448aae1866b861
za3c6417b00bb68a325f93fe060c2a3d0e5462a9c1d9603142be7e8d16be36bd7482fcd1127e59f
z789fbbc6920af7fa9e1a0b2ff7fad633133b227ed1b7a1bea8cced86d1ff5b5b4ffb68c4e62d85
z17683cef750c27b06a3fb54a7be4a5458a6d5fe1a18fe5f43a361a2c2beff3bcfff1e9f8189ed1
zd8c7e4710032c677b3f3e335fb77d95d6d7ebe50123b18a774eb7a105151f1d0775ecd9620c855
z063084f5060dbcacca78bceb91b6def4124d4234be57e41753e0fb69b3a11ced1dc076173231c2
z893f90021c06de04d404134c9577fd3c2b668a418c5bfe79628112dc356eb20cc4cca47c0be015
z195979cd013e3b892ba0ce306c79b87f2710f611eba0052f60502d1594c2fde2e52c9683884528
z4fc298707562da6e6a2fb9918ca23615225ec5fb1becfa6b2aec45738e063ecd88dbb1cb83caea
zd87cd69bef5e9a7d487e25b457701268e864e2fdec456ed4d9d4fb76b9eadaf7852d6dc45e12e9
zf3c18824bdb606fe02dafcf734f7ccce3a2ba4cf84fe44da69ec2e3e25cb906b07947aeb2d10bf
zd121c010e169bb6af641045f05c859060301d7a2ed5e9248509499d8d8c6e8099e721896ff05e2
z8d07fc20c26ff327db7a28b356cdb78e070a64ee21effee16f43e9f66bc6965b6eb11568f9c479
z5f2a6cc25c2334bb56b3d0cc1d84cb48689256223737c9f87f5ece0b8102c15d34fcb21cf34bdf
z6162a74733d634889a2757bda26b5b7161009ac490821b425460a27cc04f806b2c22ebc1c66d48
z0c63bec92e1e0debc26e77a062bff32ae63a2931371971f7850dd0b674e77c2c1aecf3f5a543e1
z29ad6e9e089204628c130d840b977a2c69608d900e9883b936f7e524babf45012d431d46151994
z6db7acf527c39c7f58dbcc4cfc9f4a249df52491b8eac6340fb859b72822fe4370479e8a94660a
z913061a33d0c8725d4c7ac10c1647285c555e89481d3e0feefbc26c19027d44b535056546d58a7
z1051909820cd147d09203231c2a9a4ce3eea635fe2d4f5a58d703f70cf95775aa552136c2c2757
z661abb07303413e67b67a1e69bcbc9b7db1e13f8006bfab864d68a31d0e21db9fab8766a00d7f0
zc535455ecb1f994a5f2d268938b7a7b65ca48e6c72e9dacd0b3e194f1e7750f4bdcceb4c6f7628
zdbfeb2d872611c237fb1f082aa052f19ce80abfcf2a1a7e518a76a4eded91dc0cfb95220f9199a
z2d93c43571e7c931c3dc3c615028ef52ed4982d6acbb1a89244d6fde16528033d75df18b2ff9fb
ze9f196d4088336cec1d9a7808e01f65c6f138f101d1da0b78f78ec7911de5869c06192dfaa5b99
z3653cc2c00d60d1d2fa234e95171b2281f4089670485441ca07094dc6c3d192b38f3881935d0b1
zaa05bbddeca84c4a65f42f19894d175b8ee98908e7fda1813fb5bff4fa6a510813610856751fdb
zf73414e00aa94735ceaabbf6cf1a4f5df9ba7bdcac7d8a6ed7c3df43e3e1fd346c29dbce215742
zf54567a1c15753b70e0fe85ce15a52eb59fee6bc7824873e84abea1db6b33ce185fdb7cdd1c433
z2829d80a10274ef2911bb2c418ac5b24ca87a49c8cd0367f9cacea44d8656ce4a3587b7518f6a0
z52678cb1b383224e60ba9e1a53ad3ea03132120d1c1b044833a55f51f6d590bd82372897a6adec
z0349610e73e82704caafbb8c6b4ede56886cd8b951a33588d17faf5644d7319701fb91ac89bcf9
z354df0ad497e7a32e5503f6332b9f42bd375bc0a26012277359365215a46f14017bec5f1985428
ze4e3c7221b7a0e039d1849bb49766cd245a1d4718a91f7ca6ca22acc856295447335373529f473
z9a7d0cf1cb55fd930d40f8da71da5821bd948c41eff02824de2f5cdc0121c54a4be634f46091d1
z796db53a4b461f6fcb74f870883b4379c5828e4d42849dbe7842ae7e26d2c800e0e22f5e2dd783
z05f506df405464fc1fc3451b703d45e35088152307c27d9fbac0e92962b8e969c5f94a2c3828c9
zc6ef57163004f561983e588eaf47e742ba7bd14d6a5256df7373876054ba246fa0a42981fb0ec7
z02cd9752b95f4069cfc6462441946d16092f7232ebcf326265dbee374ca4180cc3376b96ba0182
z9b5452da99682730c0a27c35b4cc180f22722474ae68946c319adf52cc2bf90233746968de8406
z95ea58a04eb83de4a8b5fe7bb88a0e6adef907d01d9994f6f10bde8108edd93e07037dd7979e76
z8937825a56687dc4fee91789a0679a1a9841888d17e30271d02b36de0749cd441e988ef479729d
za0bfaea36b8a693d954899efd6af23d7612129c2e97c8f0bfeaca893600664c3d83b4ba12f7bfb
zf6a9258eb699551551487911a3204b8cef40255a0b112fa40a7749fbf72e068a2c9e7ae371404a
zeaa9c1790d98b81c5d25b9c101fdd0a4ef567019a0e3cd177f0ab3b8f4b382b795dcc8febcc84c
z4b2fde224e943750ffc0e412ada911344175c8525f7d773d7216d3cdfdc53ac1383d476a37cf48
zee990b2cd8dcc27139cd79654268548527f21c175833f96242d50befec5abdc83ac153928d826d
ze2b567ebeb289978d8bf64f5e36222695aa1c562266804db40df10b724f21b2fc55c7739b1d4fa
z85a059a8bc92800781f5cc9c0d0dfc5fab68179b7ffac88bb61303d75ae66d3011fe070fbed6a1
zce43db6bc1f0430267ce1b317ed7c1a7bd285be43c7be68b6869e5b1cb3a070348b5c1147c723e
zb8d2c6c7b7b9f3dddbe79fbf5221f814c006c03a2e01c86d1e1015791bf68f13d00a28e3574af8
z2537408b6c4ca28772844a5ed0192d7ac5c8df55d169573fcac2b86c65af16665f4c2087c2cc0a
z36c8f3738dc038d3bc2064daecada20705c83a7d1ca290fb5b58dc76e73231b69761ab5399a564
z312d808aa4115811526a3463f7fb88f14969faa35f385442e1bd64cc3bb330af7a5f0d20f0419e
z9055b4150a8de89632d3baa211730cac6ee189a9a68c07235de6717abdc69525ecdb0e6ceb57f7
z182eadf015505a04f861192e3efc84d055aa9508eb6a84fd7b86881724c1c7e09d98999c11d935
z1bd1ac7ff4037fbe2bec50a13f0788c859c7d13db5d2db0b9a8043702fd8f1d90e4bb58c24dd23
zec7bb104b4316441a1ccec0b853019f2157233fef9e034c1702b3f3a537e39ca8c0e75a50332a6
z3ab8d6c1a2542c953bfa52b4f147ed9f235082a05b82499de3fdaad8d4efed3027d230bd48ed0b
z158d459247391cedab1f3d9e5356c61bc787a2dd7b47297689a68632e2334171cfd1970ca772ab
zfce829480ce31371dc7762769c494e6ea01c5cd927035bfa43dc3913796b74d557ea2d52ab8db4
z71ad0f154be075d84827b4d574099aa7ede8f72a248d77c0a1fd2499f3f52c94db6964389c65df
ze9c85a3549f2eabefa1b46d3a034c3482d97cf828a3dfd7e8eedf98af0669b56e03e8fe76cc14d
zbbdba758cbcc7ae3fc75333766f2adde28bf877f58197b9eb869da36c3f78bd3cbc01a1acf4435
z1c1382951b098e5ba0f24e6730876ed727b2b47968edb89efcfd97f8233ca0c869f5f80ae63539
z664b4ba8884ee50d7532d9e40a6b42159d060f2671753f29069534e2fd1f8a04fd76cdaa589a75
z4fe09e8dedbe4e978e610fac0e0cff12a14ab039275118fcf10288d97618cd01439fee0480f5ee
zbc31abc4168ae24658d77643257e7610d6aba87c44ac109f9f16ddfd7443e358c6fdbaed5041f3
z786623d64781dfbd9b7697aadf82ec636a7c47f922a17409a31dc84239c96a46e9e279b3214441
z7a602700086f918660bef800ce6b08a1358d55d4049557f6c503f04c5f87d2736176f33d2074c7
zbad2c9b199e817600ac97e8e306837efb90a9151d8011c54d85a67768d172c5fc56d50e5bbf0cb
z4a8721905db103d392db093f1ea00811477b2e0473c3859bc569dd43988d31904806a71b51e44b
z2c5bc54294e09889de57d0c58817e7a82917d5df1ef3e6995a4170079c88865e2ff2afdf8c7122
zcc8208a53c5b0817d0afa0a54ba055c739b5f33919167b48c66325ac6c9ad99bfbdc8334ca2b53
zaf56102f1383bbe643696b4b7fe6eba4fb18fca9c6f50d68f35de93cc764e5a571b1a086bd892d
z0dec3a8e66c32b99862063175a08b73fc39f689308278ba41c836773ecc83e735264f38b99227e
zfef9d159e208fb09c3eb732c60e5ecfcab44db362e05ad8dce845e430ee10641842fb82c72e0f9
z15dc8b1cdc724d8d8d60a6b3ad29b455e3927ef53380aab165a7ffc339faf0aefa655f43db95ce
zdf92e2a595c54941b9a8e8240bafa6b58d7504b763eea673f24ceee304fd6373dc600f66c43d68
zd2f93f2b27008eea52013764a91db471c7725b3417dfb9735f413a4c3264bc263ce71824759cb7
za1c6f952443e38e59563e38fa7ff8cd4da6b33c77e11fa10f79b6bae7629f04cf5b88d0ee48c93
z39119cf35d6591f1ba5d996ddfcb09371305c84d2b3533e7548ac979ee07b8e80d78a33cfed055
ze0e2c246314134015e1525d02602b6e84c32f0198d2fcd4f08898146c99094e17a6675aa1e12a5
z757dff13950872f4cb757673bfcbf6ebdb0599633beec4b80f8794a51929f4650eb14fdb0c8075
z66760299af4147a4da5c9b0e7ae20f087e05e0348ef407f3cd119d1c733eb4e75fb29e76a73c49
zee90e617976c0e8a17fad5193a87d61c3279a9e7a46dfb83e2049ad8b4ebd7131868a423ce98d6
zf963f25a975ff0196599542490069bb81c1261d65bf2802838d8aca94c5be8273239910244d309
zbf525118d77b55bf22cf3150d0e62134d8745a714f596c6a1b7f35a7a7729be3b8aba6f0a3390a
z0747f7f0ca84fc0e7029fce50e9fe364de9abfcc571714fcf6d7e3f93449bf21ec4e486ce85ccc
z18e7508012d9b30118b29b701dc4feeb61d93dfb4bbb0b369a28efbf4ee871d082143ccc7ca1b9
z1c26cd33c3017357ff50a964da0b94f1b7ab593c1da8a29bdfd6b0a62f8a3e0680b1beff89b1a2
z4be158907d25acbef50d6388d926820dbdeea0c8b07ba63908ae2eaba28dc6f2b17f769922e7b5
zc776d2fd5751204de06fee025828cde8defc9f86c0341bb28cef7352571c1879b8a15da7c83d28
z4c33370d8d3fd503914dc8bf8192649c8ebc1a26084377dfbe5c48a14e07b091241817735fb53e
z4a94cd54491db8061197281f1cc59911a5736f090d5cd87c2b1df843eb01be4031fe7981a6d3b2
z96aec34ef859819ff6e8271038cf416e0880f7f68048b2df694811fd34da1a99f992aea7490624
zffc1c3704a836d01aa2051f4f591c110aaa2810433fd3e4fec2e9ec35846d6caf95f2383dc237f
z14fb4b057c3f7e0fac12b82a3772e987d136c2209f25d2950398747be82b2a75882f417cf82683
z3475a1d4e8a8a7a3e0c47fdad425659dd59b2af27316b35d4cb159170f552d3446bb7b8c2226ac
zfb3087d130b3d1b66b7020d4e37a82c2201ac5d5f25a48766e48b5a914647ed56a0a84f6a25514
zacfad832d413610ec98cc94883e6f15edf8b3ff5b27050735136c3eb30a3bf0bb71be690f5913b
z4d376210685d5a0f14f3e86d83b306e1348ac2469713449f2ae298ca70d642b2c636977ef71e42
z7728fbcb217dd939da4ab45aab5c1d4a4acb81dc42c727e07a6771bd2673dc6543f3424847b236
za4a63cd4d7d89950b84fb0b07493aeb2866ccf56e86a8a9b371aef5b87f012c602fc78aa23f65c
ze10986edeb50c35200f9dd1e5da936a2deceaa8383b1d7ba46e86aa92a168baa114d9048a83ff4
zd718cf0acf61be1a895b955578b7ab57de54f0cd56ec5bb42c16ebe5b79a88dc43f78475be14b6
z7295319ae7de5b75ce1e8d4c0748976c7f577c9ee333c2f8ba1cc9214b1a2af45bd4ba34b4ef1e
z8f79700f658c8079dc5db35775aafd53e33e7b91d79875ed2ea239c030749b91e7d3fee3c76c33
z50cbd40e6cda01f464847f1db696c75c321a9e7fc6f6e03e9074487b6f94366c927f6c5bf36646
z7223ec8b947096d2f563bf22ee4e6147ea57fc35d8e6aae82370b96fae7f042a68040ceebff586
z908f29934b293581536743b8dbead1a3e1b81007778e258715a5d9d04b803f02564674fe9a6f9a
zc1045620d6786d5cc00f2b6a5f3b69fffa658f6606832505e065a1f58b1bf6ec59adedb3c7e6aa
z9b59d34b7438d3f642a01854e9fdc1861a12324349796862dd450acb0483e70da4551e22438d93
zf17449667cc58a1b811d0ca4e642763627ac8bcdfc7aac2c07a6d266a201c2b18d7e502da7cfdc
ze3e63a6b1bea89fe6320f4e3cb19a7564be67cf673ffb57b73b0607913b91f3c273430a86fb573
z08b3225672fbbd7f835aa7e9ee5b6a59af827d17b4ee68a2d43159f40adf1751e96af3b25412fb
zcac05cd1e3432a54e24c4a7c2f88f923aa8db3fce013d6b179bcf5090cdd62868c86f8d405153b
z9335dc5c8007cef8dbab52e5028400d4febe70d08857f470e20ef24337e7a7fbcd74f79b186026
z9f1356b716db335051eaab4c53795ac9e574d5e25af2b329598bd9408b7d2451f9ef404b527123
z62dc658d30559d5b6b01d86b0823171b815ad30ecad5291eaf7d3294703d2ec97f2885d7513a64
zf684158ce2510d2fe0a64f6f8a4c3db6b8363863fbf0bb7c225f0fb5afa6249c89cac6c4605ca3
z39c4b9d37f223d30aac964aadaee5a63bd2807ab761ee53e41a8b2e390f366d2c765b7cfb93ee0
z4f47452109f943a83d15ad8acc3e5afd1b6bdb4504794c19dfc8f2601f0cbd346850c1d0589d82
z237ef0075fdc07c2922b30f5c570393cc307571977fc63483573c3982527e1df890feaa0cc44fe
z9ba17dd896d82119a88eb69773c650bf079e2bbe8c3e198fe7b829370838cf7f9b7e53ff936c7c
z0c9b52a752e1d87a912b381151393d985ade9ce227b73975d220097c2d6e0a4029b3a52f6226ba
z2c51389d307e1658202e6f95dad2fcbf11a7f7431391d46c55ee34207be5d448b5cad4c40f5264
z480249305928a244a7bd227688efbee1086ab77a42358ef164827fb398ec77f54eedf26a2eecb8
z234c08b0f094f95153215641f12e0edae887956d14b525914cf0e1809ea4aa8c0b553002715c3b
zcb7e7b63a52b0fbbaacb5433163e372bda43de74e300a0184a7cabd1b56ddfa3bf7928e531a6c9
zc94ac16ddca57e9bbdc14fb42546ffc61d517837fd1f27f35961d703f7efcd2f5b4a2840a36bce
z196334f1fb7d320b96e6e8e9804001c5f8f185408aaf3a09469dada5216d1b150d6a810a94823c
zfd41331faf156767a6e54524d0fc5d06180c4e72e57b8b02abf8a733ffbf1333615fe6293c1fa7
z1b32f5ee2d061fe2964cf2ae233fff57537fb86fa8134db252d1941da1034ca83d0d16ed0462cf
z686324d3e6be3bf4032b7658c0995fa7889a2fd11109cb056c7cb752b6ecece9b9b6787868db0a
z55a42fe6c9cd330d1dff7f594af547a917df120190ec6665d7d5cffde14350e9023b035dce82fc
zf920b2a805d1d38c9ca55d8b0cfc5cc34d11128c1a658fdc478451178d2f4cb6722ecab93e4edd
zd7a51399ed430973e05c78c82445ae3ef7707f19b1fec3bbb0ad2520b9213e6f44b90f9497a43c
zad789cee3ad8d849dea04e306e607208077e0a4c0db60c49624317222552c78cdd2c4606476db4
z52c528b40062a97872c8b29c35d4d600111cfae46e9614ba4be3371a6c60d4871e2cb8360629b5
z555241396faccc52d3aa72fe0575e3c9f33249f86edfacbaf61bf83de31fe07c7cc8873b34e5d4
z95439b0555da4bee581fe9c7042e2661c151d32d6166cae07a7af925720b273b57ec258796aad6
zc3ba4bc28f4cfc0a42e4e3f5aca8f23f7bf22a1a37a500a15ed2f26e630ef04ca84287aab3cf93
z8de02ac0c190de044b3bedf85e2350f34c1644bd44af7ac0da93f43e7e16717082f1f4eafcb4ab
za35327dda818e28c7b9ee93e8098b5fdd735a89684690992d0bdfe217a26120c0f422c93f0d79b
zaf7b05e07e1f964fbe34f0037689c59be101b481920ed9a522ad2f00a09e20b70ad8359e151a76
z01c853b93359c11cec9441a0a9ccb75d210be008b32c03280c9a807602f6f5929c788a50de0d22
zc7ace5fc5955aeafa18d4adb2e7463b58b7134a633beaebdc52d90115142fefe48a7b9f6357e18
zd2b99871fc77e0c95d9449a59f502c31cc98b7bf60577804e3d9a50123fbdfe35593a14cfdf1b1
z50275b3f3a355d0bd94335a6b6d836cd9369674190d4368ebc0dbaaa89cda9344d424427d063c3
z70906c41fcdf89055dd9629ff28feb6db45ccc6d05b19d108f75b02e7a972896c7315c52998329
zf7e75dc4c36c3f0c7202adc73c8f2fdbd66548517d1cd4293892c9af92a6972869c933c2bc197e
z14800b404f1d7f1891774688de39cca6469c19b492dae7b50256631d5bbf64e921b8807a63b37e
z39617fa3fa560326d101b8b5034b21c5c16259222731721021d32329b824171e35b30c8efaf802
z040170b29958f29da527123f7c053d8caea83e0347dabbdc19cb5c390a40e4ce52b94eb472e707
z27d5adc7f5fe6a882a1d634b5f40691f1005f8746b076b7b6314ff1341778069ba8153c3b5c200
z01a07bc29cf694b35f42c940d361d3f4d21213f904fbf7e99e6c4494e7aa62bc1ba3c2d98b439a
za00673e29c178d2f6439a6a4716a65674930ab6d074b584f05181ff17bbb03f6d441ac545677f4
z098a6ae6178a9da51727a7bf01db5506f53b62551acecbd619bb8846f9929ecee5b661336a940f
zcc9ae6802eec7675759ec0038cc71416a5ad587157a6f421272bd22aca0a6b1ee5c8fc9a6c3544
z336f810d12622a4401d9c05309578623cb88f543b421fc44268766b7a5dcbcf7c372bafd4f64c1
z4afc01426e88cb079aaba355c71a3231e8dff2388316e3dc3200af54e29bafff88a15aca6544a4
z935c244e00c459388c986770c60717b394ad20d6d8cf04c9fae675bd92a0dfee115dc7e10a7c68
z6fe6077fca78857232716f445ae3da05995adf41c834e8ecbbf0214836efe6c1c352e4eb070dc1
z611fe7f2b2efd32f581daeaac92497b84e34c314b837d4c5ef449f78aaf10ab774db3303c85ab3
z4b0a7847d2db86d605e6ae8284fda85e54a8ff816fbe03655876b09a3dc24f9923e6ebd9b0f53a
z328ab6f08ba8afa5757fd4acbb877fae24453e3f6dbbf8180d52d55627c524ce52b61c71fc7c5f
z3d9b43de9677ed6a62f27e6c10895ce02223867414d2886588b49c78e9eb931737b3653732d077
z8441a1eec63b85fa6b53f278c5fdf2cac41f1e64c4c6763ed54a57a9da60c16d3fc538db5d49a5
zc7d2b5a9d5f08f11d534eecd1ca267d8a88d02d767ec7350a6e2802165bb45034981c98b23c1ad
z18415938898e90eb76ead237be9a0259a75146b5df3d103110367ca32297dc4d213ec7b7ba3a3c
za44f5600c49c110cefe2d09563fb8a67b65e523a213470c7c803949c899b035d01d255add93087
z64cff8ee8480becc56698e7e6d5a75fc0a8c163654fc80f0d84629c62046f35c3429cb20690aaa
ze0fdb6ce322a7d22a9bad2c6157f3d96ce0ab5808f0cfa92836336defbcd2f3c5153c7a03e7649
z0e362921dec7277508561992d0406061ce97a80093516bd6ace99e0775a8d38e9f6b171b62db8f
z22d79a7d3e45c18d5b9c11741519bbe7cf69526e39966f555adf6dbb3eea065927eec221ae6e63
z2fab3b3b708f96897ea8c3f31c8e015e9e4ef2504a3d0c30ff5b58a514a8764589636c76f2b54d
z3177c6419e0218e9166ce8f73641157f82c47b4a2e2cc97153ffb20d0c9c7e506054263c91f03d
zcc8a81e1753c20e3e93f10466aeabd729b5d2bb18c440e45131e219917c00393bc00613aa6b861
z1025a36bda24afad55428ac1895e7f7d317c1295692ed28517d9046dce31920e56482ed2030345
z9107fca36f1e72e58426995a36529dccce377d0c07129fe39de502225f392242eaacacca8c89d9
zcd884d858081f1cb36ea2273ff791ac345232dcde1c9fd0c5e2c21b4cefe6b448f04409214d6f0
z25fa2d0bec04b4177f85c4c68a382e1986ea379d853caa45ef032cad4e84bdf082e4bb6e760371
z0419ba1fed6394e50fe68d367c67056aa835df39d19fe7ad693892e4ca5073921e123b9bada88f
z640a97f9e23cb1291294282d50df37b33146f639018f2a2425611f07a12de9ddcb409cd1d119ef
zb351900f77f2287f54c15dd523e87c2f60527e8a3d17118b7b1a9bd663bacf3f71b46c6a8abb93
z6bfb10e1e1e66eabc9b38b3036bc4ff04452748718fa09360fe4f6811acbf8a808619c75ead38f
z9cdceb31ef69e7cf0ae6e6240cd3d498b6087b732f8acc18fc2b238daf26e534dee339929acf82
zf3f1f831ab9997283d73f2e1e73da4f40c211e1ef64e8209b4c34ab569fe6b676e2b930009bf05
z3b0d1a8fd6818c371794dd49d14caecccb81d8deb75556270005a697f5d6d802744b4dcf41665f
z7e822634a1f2ceba45ea3ea18e4b9f1b3093d0b575d1ed1f06bd14de278e727a83cdcc45644aaa
z9edb5562e215dcf74b73ddb2e044eeff0a07f60d36aef4951911fc11fc6435a30916e3e4d0ae10
z33f9972fac0769a6c25ba5a56537050e4eba8516515487d42c386634acb500f3f8e5959761a187
zca0677cf101b4d689476795886f6c2e7e3f601fa5569fa69fce43c068e1a0006ad5036edaf3733
z1c2459efbbd9e47f80a518c65a810c9d65ab41267201be2bbb075f7a8604cb372adc08161322e3
z36e3569113b5dcb7aa5ff63461ac0c6fac0d9400411a501da132cc729b549b53605d4b55c1e7cf
z2a96a233470bebb0062bb5332bf99859ac784cde3fda4621b4807e1aa6c103150364c3eaacb5c0
z427d1a33385da3081e63cfa76fe2b3aee711eaadb53721fb5a274f96da0a0bee1608548439c650
z93195d338288b674c8f1cab3e43a67a80bef528652c13d17f6202334e26a9648fafb186f51c627
zf4a826952c4d588efe3d69b62f4dc31430a56ffcd7c3b79c205eb894df1915278210d18ba4f058
zd54c8127f45cc7d982ab4230ef7a38ec38c37684b20d553c64f54f60b74a92798d797ef1ddea8a
ze3519bf86fb6f519119e8b59f10ad8731c56790b16be5a1411f51d76844e5f408a4ab7911ac5b9
z295f17f1438c2b197e1991f2c706b2fb18a7103ba30365d977ce42eb677986ab788228ae839463
zb6b85ab18d496063236d983669318c7b9073c3f75d3e54da1d1e885dc58f202675d79d7502efc3
zb6e28a74f390c923b86f33e174f3e0450028cdd3f80e8ba72cb5ac4e1804816c04c4d9cfb5711d
z59eada0a16c971d34ae6f134a634b5fecc8f33c158bd8358faff2ffb22eced23be0e1dd9ba3492
z79eda126e1e377ad0f111d6926a6b92ea197ad9e80d227a0e05e6ce2a8df3b5a7c700a698f7ffb
z51153f5ac375e5119d88da34670a525219b85b91d907708653b7492f2938f4bb9920a26fa68ff3
z987f62220c171094d09dacfbdc6873c8a14927a1232732656a3184a90a103ebf16f788621ba460
z0b4fa35857f86b02c57dc846257f27fbaf563df919f73ab8ed63cf6ba59027bd95c7e082d2c4d0
z5dd88c881c9b587b59efb40625655be36a947d495eaf2b1453843616a2a5ee428a3137eee255db
zea215b3a69fa34e59cf9336d5f3f19ac96adb08e200efb642f9fdbbec7d02f13a19c0496373e9e
z7536d688b03468aca35478735bdc371681dcde7bcbcf7455966e28b5d45a214cb7085590746ec3
z063486ddc474888dd5214d3b4c7864694cfcb889e45893414cdfa4527bff65c75b894b83358142
z1de4858f4797a90409e05429bdf763e59fbfaa31fb3c221db87748b957de5f5626617058b2eab9
z84a39d07374ffb9900ab24a4e88534aece12e48c8ce182934f634d9c222c0fd389dad17b07e9c0
z56e69b6f9867ade8637adab322ec69ae77ca144227ebbec2abc0e196eaffded7fc104d14e6abc5
zbffd220af27e8f80efd98259201f7b420016193de112b78b3e9715c816c9a5930c659614f6db6c
zb587abef23f48a477f154b106b59b0125ebf01676eb2da777e49b698b91107d58246680c2d3b45
zb066e3a339ffd1000b61f4566d999c3db58b954a7513db9a23b61899a12ac674e4bea329c54089
za8c5bc0fab49eebc72d7bd220150518013cb7de9e53f130356d0a3e16126569fd73c1f1bce18f4
z3ed46718e2ff2e6e557be37b8299aacaf8e4a07138f05c17c8f96516e7e3169161fc66237e45e3
zc567a6b20417ddd8efe19645f97c1ad826077de2a52854e5d519f3ebc304ab5c357d1cc8458122
zf650699190e31727562a507528a6a5015f040551601e5b120ec3797c71428979cffc7aeb696b7e
z28475a1854b062e25d77c1a13af741d4c3421de85beb9d9d3f075a10240828b582046c2a4ca6a5
zf23898864fcf7f6d40b455913222099c4edc6c34deda976f044c79ddd31acb919905b5dba1d680
zd26a844a0ea907bfd72e0ea6b3310a6d4c2c8a1bd251615b51d3b98811f3a4eacf260e9410288d
ze9ad9651b280506adad19e9c3fabe5549d0090e6b6a64ff45bb90fa8ddd09f2498615376e9d4cf
z2d22dcbe7d5963b798dd1f3991128a736f323e7eedf5ffb051025dc3a27a9bf03913532b7967c8
z48811d1930269d9f7ae5db880c5251aec94d069ea118b7587c6bea6df98af801fe0c24f74c2c26
ze77893b9fb64a73875af141bb9aa37cf471a6f70f971908a19cc4eb47ed56a4560631ff61a443d
z2e26db6d7c08fb0a17ac5aab0b4bf23dca4a15a35477ea2ace66749b271ded05e9cbc73250a7b3
z86ea59bba03dad328d269f38ba4f8e07990bcde6a43cfd63b66c69bac44dbdfa3e1aab29802eb5
z0cd0e231c9b170c1b3f2f359266afdc7801707055161bafd3e7f4b95bfb5e2192ed3bcb7a4b1d7
z5e5e9be7e2b68bab5077f76e7a72ef683fc67c7115c049e752b0dee385e353cd9c099a726b61f2
zb4dbde0e0a8de415f711dc5a4f063492e072a27483b33aaeb83e9c35660a17b34d3525b8958f78
z61e81ae8eda7c0d4c3ea67f9e25b7730ef70a5de94cd70522eee088a10b5065dd258681d49b617
z002f252e72b0ad312b3d0bde97813671b9ec278a1a5f5e1d94f5de20e19b61dc5ce5f17c4e6466
zae9c10161d92af992ca45a5890d6fd79d2037047fa59f118bcc7b60fdaf11fd532065e52f21f3b
z71497911f3852aded35c3d0de57362d53761ca4b4723c068ea1a3fafed869bca431c5cd01f85de
zf87ff09d350effc5eac18983a9ea1a09340978a7b486fa27d8fe8fd34b58f4a903eee3af2d1ce2
zea2e82a5f77e87f1cc7112372f881cd20fb8a03343375547a05e7362b917dde106b4a2b3822955
z5057898775fa2f7c1d2997623ed758c935fb755b3b57a66caed2b9255b6c3b72be2a723b3e8560
zd328601dcaa1d167094d9f81246544e09c05bdc92699d572bc20639c12a2a0d9b98e0c8097770b
z2e8df0f875cb8f7ba940a72325bb7390eec46a53588d69b6bdaa849e1fa31a5ad28ad9ff2315fd
z5f85be5fbe1f0c9bb53dc3f85432e217cb46235c53df38465bb4b68701259c1647301124c4e4e7
zf48cfdc827272242418bfd49c25fde40a4590ddf4e770380b04a64827c2eac3e8fbbe116387683
z23e09d0925df04a4f4e0c8d358e80d29d88774a37c75008179c7f4977450ab4c524874e102d278
zca3813ddc5a3e9f43d377c5e2ace5d714cb584142c262120ab58ef589f8972934c0dc79867150d
zb8d3e76500a7011152cdacdff5023b3807cc53a45602f5ff9b42186627173b7c43032d940e48ce
z7fc132e8873290e5c289daabcedc22eae3d7ee418cd8d073c349565a8a8dc45e44c7ba06d40180
zfdebb355d8f1df00e5eacc7347e6ec0012ef8ab079c565b300b00e26959cc8377c841e6c5455cf
zd1cb237d0eca535c99c3bb17682fb8584e9fe136265c7564e043ee969fb2339a7a8abe76605962
za9cfa5eaf1509d49b4d022659441f7b6e3bb60dfa3000e46c22bebbfc306a36c1d4ae60581ede1
z87b80602e3c09ffc41ba8b00f3faa52462bcf3245d1e03ee7875505d06f993024c3a80a9913c86
z0f965db88c04bba8dab6c45e37479b404fe03f55c373ac11d43eb13721f3fbe3638a934d1d20c1
zb601bb1f9b8403a17580a29a70edacd9b80052ebe9cf2fe1cb7825c9006735a9c701395c4286c9
z341694f0de68247403d26985e5343afa3d8d71210ed7983b9268ebdd34aabba850d381525e2d37
z60286dd31422b1a82089b40eebaee2d6eeed2f22b5a35b9500d0273b1b2340773d00c06ad44f54
z2236e9b8196cd60b55af05b9b2ed2d367ecca9c78ef6c1fad2e7b55e94d5ded77dad67793f8c8c
zff0113f4ff12f7b8bdfaecffdda41cfc83b15d68b436b7acdb586315aa0c58737dc1bb32ccff68
ze08af8d4db35cbe677d4dbdc3ab80e57bfb827dfba67826c3d6a0e26dc6415d7fe406ea175d68e
ze0e71da3b216abc91fe81dee247912926851c5adc53fb9914241f68c58276543244821a2d4309d
z037a762fac1134628617c4e113bb2fc48ad23f0139c31884a0b8887a966a62f2ff3b2888c46a72
ze78f3a8702191d2cbb8f48fa991fa59bf954ff78f6af5900c9d39f8d3129b1c7a3b2be1745d900
z66fa5f2a6e06fb3e0c24c4cfcd028b43e4280f4384aaa3c7e2db8c4e8174f2f7b5b6d0fcd2392c
z28b394a131e87544b7c92efeced023e6334b7f18cef4d48790c5c3754f6528d5a3ff3f7e2fd896
zffd2ac9d20839eb1cedc1db0b4e86bc101b56cafddeef86f6d15fab943ec57b8604b5b83b54b92
z2c9c621c4f3df2af11a3ce2384601d0aea99b96d1cce2961c96126fcf29a9dac7a8cac47c19041
z6d0c135fd3474f24ee130acc6be0945f94486907639a830aab19c962adb6362dd189a065d64901
z2447ded3adb100bfdf81580af9c0543b3a5c2a43d7ae2e4f5694219393d5c0c18af9e0f8ddbbb1
zff5368a5a58aca4b76c2564cfcadc1817a164819a6c833fc6047ec5690c823d3850b8bc771f2b3
ze0f2707fc9c094f471e35159fc60420ac6ebc4b615407d44510968c5a13319e1ea847f417e6550
z47b4de52e3e70995b9fb63b6240455d288d41c31aaf10a879273332cfb7ea16800950c4c637a34
zc37ab236a8d9b5b2dcc82beb35961f81be29194381190016b9bc600951aae9be262dc81d11e674
zea1a45e90c52599bc54252d7ba86b7280550acf610ca9113e98f9938412935cdda0adeb6d7a6cd
z3e2e08c736794b6a510861c9baff295ed0ff169df304aea9e84553be526507723c0a777b231c40
z07399dcb00566e9d013ac4d54384904d47b09650f0731232cde8898e5e39ca05fb0e198ac1cf40
zb4c6ee4d0cf6a67e58e41ef2de381d41d483280b6a0d69c186c217295d8640f3f54aa32f7ebf6c
z04dfa3e97f65ba40095ed6e0ba971317277ad7d10951eafcc938d525886bf8b761ccd091a71cf8
z488eca234db244249f290a7d126d61ab426081c5a0d37e8d87a8a5dfd5997e39d70a3dbecafc09
z90eacd305a2cfbd106b4425358ca0f5bdb9db715a8af706c761bb896739a49306f700fabdafe20
z2f1238d8ba01efa82e5170fe572865bcbf394b54ad3e8c461b91a868fe038164afbb2a92a2e23a
za2a921b848e940a2631e94d6c32e492aa3403062576091fe0d5f820854d850e32b3977a5a70a1f
z6c75aaab382c5b76843b9314f8b53f63ef2d9eaebe1bce56840299c35ad5200851c26e94395d81
z3c42a01995cd2f65599fbc2745cbb71dcc073eae42d1defa560a82accc5f8d8993d7451d077b4a
zb687c6121bcf86da06f0508c2489ae65c69ebe14b3765f6acbdd27a198ef02a7c57e4b7a919060
z5fdd75104b0b9132760cf3892d961d967a4c41ee38bc6c735c3e6932919f7d6bead5a5b0d5e2ce
zb297abeaadd2ce227cb39cccc0ce913cd273fd8bdd43fe4205e8233e479b4251200b1901bc67bf
z61c5a73ed8a0015a8069c359dcd6f00231f5d46e9ff237663daf909f7af607766be7391384664a
z0e0617f487da18eb663b7455dce10d85986acfd71157f782d0efb746eedea35c7d872e49651c76
z73454ce400da9d03b54e435119267d1eb7c84cb7ebc983618b3728ac85a4c2bf6bfaaefc8a348a
z1e6d48b1893782c1efac4d632b667cb8077a20233353bf6f2c763698935711dcf8fd852faedf44
zd33d144f8ef7305be90c2ba0a7b64f57e31f8dfcc88b7b8c9dc2a2f5b0abd8ba5b98cbdae2f68b
zebdbb41461407820cfb3689895fa7e297a54305edbd4ccead4dfcbb58a1fa1d680c1d1598d61f4
zfffe133d3a04b9111988d32fc53573ae5a5da6dcf9b220dc37516116ac2b930f3c61fafba0ed8b
zeaa288946b99b1b14a139a818bc6139afa6b2899128ecb62a4ae4ab57a8106f3fa83ed23dba4b0
zd49f7501dfa898e65c816630ee4b7acc7fac49fab9c9b7e5e4cd3716db3388ca9f606541e178f3
za4dd7c6e23dfba0fafc96190f7bffdb04455812bbab8c1e21f6cc20e69409b71588c25fddbb425
za691fa7f9750338f618b29b4877ad97f84115eb433ee3dbdf409b417e1cd350b2f4b8979b967a0
z99d00fc3e90691a4a056b58ad0e2ded020401438d6bd4069480e219c4585fa372cddcffd927269
zf3e5a41f59bc4b1e0768eb3ff5c35906be0e67eb7852ff5794e03bbdccfe111621da9e72d5f412
zbbfc7364c5306a1f8c66ccb5b555cbc20afcfb6fc01164e482c1da51626457fac202e8886054da
z9f82172a3eb6b57cf5e933c5c0f6569dbc50b3771380686ab7d759ea6c5691b5dc3354758eea42
zc71f573e29b1231eb989d8b55faab45f9d5c583b42a79ce797978992d6b735580ba351f8ed107a
z39185fad45e550d04c96185462f7a40523b77ea278b62396dff9109a22a18b8e952f4a06a11ced
zcfe38c51b602486fe4022cae3a7806a81c49152a32487880be9c24a3c820642026d212a21412a7
zc14d63d411749b7128f185ec7b30cc6457ae471ccf52021465b657952a4c74dc8ebc5b5c7adc80
zaeec77e2cb3ab36a5af9d5dfb26aeae604385c1c7fd74c3ed17a5bde2faf53bf49502002be89cc
ze4f56b1c497d4a5448465ffc9badd174d10fd315be30ff12083f1981f261de945d911c8e0d1df6
z8bb0a3c658a19324e1d329a9bb747c17d443e30f3862554f1652b087a39cae766ea44bb181bcdd
z1d02b8a94fcf5a6e8f5017e442a9a3d8c476141170d5cc1257808ed4a571135a004bb629c44d20
za0baa82539870979f6df3892e54397b88063a90545f7ce5a30fada247b6bb210c81f2daf776e95
z62c57d78b2d532b65b417ddec6a9994ecd3334fd8b18d05b8f8423ecdf7222536f169dd1db82f2
z482bb198b06e7559179b07e79d28195629e7bda400340102e934b850c5080f6e8e6350afc1e4b5
z186f5a9acd7157606e663724e780398377ea0f03b313984a025b4979beea55b3ebccc0b046ee26
zc595d7a7decb3fe0d5ebe78880a1f44444b0290dc6d8076c1d51e0dc839451ca1061c4069078de
ze2b31a7a4b5f117f989fda740f0f4588cbbb8ed038b611e0c9bb498c1f258d81179eef8b642fa4
z8a16e449096a23f3e527267b9ac0103305fd1dced0f6bb536c6142ec03d709f2dd804908b1e1e7
z5cf6a2b1472380cac105aeeb6280830f4aeef667632bf6c4ab610e168eea41c362d505dbe08d41
z6597bf137efbcce1f1b7cfb93468d787a4b030f491b50e34bca9013893072e2eedcab66f7642f3
z4b43149a62a89dff27ad761018a45896b963e7ca757148ed6e9aecd8690413bf879278caf6799f
z9dc101215cfcdf98905a75fc3dc33bdfedaa3c91dc0185b595ac948e1fec0037453b34665d07c8
z9351752294b38159040b720be1dffd632a4d7359ee2f7407ad53a048fb62b783a01325a0370b36
ze1d5a664597a4a861da2c2e364189a2b8278a7eb34aa3835f561855db119bb3a6df372e5b8afcf
z7d560d1c09972085c720a1d9102db590befee75268ae77f7f29fc6fa24196ab762e1e6cb620388
z5664bc5e1ffbc1ada1f43f2d43c43776fa730290feadb395d779aca00cb6cff74feed91dce8677
z51d076b739ccc764ee34ef8758f68164ddc6098cc4c91e2d2b2baaa34e7e48eecf6405dd51c429
ze91974a3f2379f832bbfdb50dd4c3fc307a6f56e6116fec3ee2f70720c59410ac09d9a9b43c846
z04251cb440e519d7f80a8a9ccd451158425424e4723f572a2e556f19dd385f3768ff28db0e8074
zf13f23a6ead5d2d5c93c0e1123a573517d7714efce45df672a6d540aadb66633db7e33243af7a0
zfc0088e2f819ef8abdc1375891e9a8f03e0d02a9e7dc927fd3ae352ae6ea62e14c528dd49311aa
zc039283d55f59f0e7999c93ba8fa822f57a43e10b3b3183f31e697fe182985d2c879b07824df3c
z4c4e46032a96afb0e65ab9b01911ec42889f563fa88b1ac2b311b92f17d0facee7d0bab58c64f9
z2679b95829373b6b074fb2a18aed0073e51b70c13bb9cac152771cb93b71342b058b9fe2b0b775
z987be7328d16a09cf71671ea1f1ba11495afc2f8cd507ac53332b14c65d4c0f6a9d1fe2e5720d0
za6e01adb732f744d55d29bda0b63838b28cb7a0ee7b4c7f46286a72146029b7a3c62e9f48becc8
z61712487d9363842e1c1ebed821f33458311ed98bb56ec22880d404c6854d86b10742eaa853c87
z316eff540f75be6115b57f4790ed8ce826bcb5c5ee2fdc8aec81c9f72d530678b9d5b89a252f6d
z463755270e6789728b93382f5f1d53cc4c61a455ff4e5547f9041bc6f036dc5264bfd6e415afdc
zcc1df604c5c026914ae569bb1203384d1789f2439d7b4d2898e5e8a850a2fdcc2f54028571f371
zb4663f732a2e94269394b7bb269a24541e34010f2fe1ce657e2cc686d2f703ae7219b26baf4861
z7722f7e9690d2e62efac8ed21971e4ba18cc6bd85e1ee561f12b0394ecd059c90cf27fe8d64f80
zf5326e9cee3838df134141b63eed23009150e66e0429e569dc5db1829d4aff56735f4ef843af05
z7f62f442834af1a1f8f22c82058a3b94ca0ff4789a9d790952ce3f5c9e46e06ba73d212b41ff43
z55df1138b433e19b87f91875736d8ebebb9c2c7bdbc69487d59503bb967b529686b49dfcd0a9fc
z0ab3d428cb39e53f3d443412f64f2a059f4aaa918e0317aa9e38647c071cb552296e228f49aa46
z878941ab448480dfb06e7b2f465b95160cf5b1f5d0b2ea02342bba17d17778daa3df90c82b3c95
z9a8624da2b79a33776f156bdd300fff136543e5ec612194edd3115a22949fa60cb540ab8e6bdd9
zcdaa47a24fce970576f02c7e9e63c84ed0161f35d5c94764fa509ae071bff5c6ac74096915a598
z89c8c20fba90db9e286258fc7c7c7985ddc4182e44f45abc0f1cfc7829f16e3e437262b89f9e2b
z678b97b1b0d597bf3004648ee47f242be32438b11f143ad48cd4d02f5723972a57e1ea95a5194a
z1aa4286f3552e52bfb193a2e08cf3120f4394aa04bcc1a443b1b1a41a4c92b8b07b870ab816892
z94117f7639432150da85b2acc7500a7e81193fc55b393c52d1d6919384bfa3447dca3d92b520f5
z5b44f2fd78bf41e7128e7a84f680932748ca65fcb5f5f03ca727c5061c56e7f3bf085e8c62db0d
z98aa3c7945d4e9988e9c78bcc9d1630534c21becf1d74b4649f6760e2ba82768d4a38ae426e8c0
z58ff150a97752306dc6bf9ea19e70440e521f1b840179b91e420fb85dba5dac54b66608bd9dd0f
z6983c0c8d6731255bbe2078f5283e295e87bdcec4b33a76a1c9f67dd90eac516b03b104b8d02e4
zb8ec14564144d39e0f021a5b1cb21eb1f01e6d574fef406b98cc303f81a543423346c3ac442a75
z57b867158695a91143d72274839d4cd74245da1282870fd2599d974bdf43b18c342b3e091ed850
zb3c7c795ed1746efd03706cb7a9e749557d63a91f354e95474f28e26aefb5ead92b2a425ebc27a
zed41ee0a9ea68cf9b6b063af309df631d5b34eb55e8b3775ba72803710b3b6bf474265a4cf28e4
z1ef97d3ad16acc54152f02eb4a63dfcfc4a8ce171d5070f39d8c28a34bede4856dac40c827ed4e
zd708fda6d09023dea5104d8fa78796bfcd137b2c153706ae406425f4e14e5582d606a3ccae563b
z7057e9a162f3957df39808938ef223c22eb46d36cd4cb2d7782c94176db8eb1817d63e5430a4c9
z5b8fa1a625742d5e42e75581e2b72f1e7a7db0de9559173b31c9ed9e05129df6cdfa7cff0807dd
z86527363ebc0504cf39dbc4767909310c0211be8eb2958696d65495a6d18a1ad28b247499f63f9
z17eace339e41d84b3dd92ccd0f303e3baf2cd837611b99cb18d99696a324c9a401e13ae5471542
z021532ebd468f307876cdb9c1fc2f29573c647044420a3e34a1071061dd45bedd874f8b456cfc0
zf64ef71d7307aaab2feee9c0dd8a7843147b1690ba031abd2f35b7cf38d20b549c454b224b844f
z5f048ee6a6a426e21610fd5c0a2eb82d1538f983f9e8cfb7d2041de67695f3607d67dba8e858f9
z7168a4bdc8961ae82c1b26614a94d278847b663052ec28617c198c038e54ee7d09107d54526d7b
z4a18019d825acc1157ed1ac9a216b2f1188bd3b1be88887ef2b8c63be6178ecddbdc43f990fa2c
z3aa84d2074ad7c65071838c756255ff54778ebe7af73ac5dc97647d9451be92610e544d1e6eedd
z032f0ad096afea6fc3436d170b8199a02bc7833c55e167b2602883c4abd538b1b169a6e293b997
zda0ad472c9754ba0661c15596bdb00bb3205d326fcf47c1a7e0228cfa0bc0dab2fb42a938d0878
ze232e21137d82916d7313b074af8e5c6c79233e59270a36d114420cd3002706873db67d92b74c4
za12f1ec75a3a1275a2e10dba046ed2385ec519f5f65c8ea5dbda3ab545cd98998bc62d12dd2d18
zd27501dd1d250158b731fd7e3a1752be1c2af2d34dbb90110352cafb73f9b0e25d49fa684b9630
z7ad3de5e607b2bc8fdbdbe077f1197f8911d150d284dc2733912d7a371e76748f4e15c88fbdf59
z79e706c8ad0f24dde4c84cab265788700e651ecb786c9ba624e7bf55ccabea0104d743b82f097b
zd260d18cafedee48b8fc130b582a3fb4b8290d8fe7e01f89b50e11aec62f9be594494c0c18402d
z01aaf6504bb24c2caf70d9b177c0ed004b74817f4975248dfe6c2e5924d21f7c5999487ec99e6d
z922d459b1db933f2d1ce8c490e7857a84504b63243fa3a21a12e84f0fe053582bc1898470b096d
z0c40ffade865b9e412de36e3496ebe122292232b8adfd016f8821dc89910ea1e20940e46ccf0c8
zedf161080d63534483846608623f3dbfd31fe0632e26a2d8af993ef6f4eaa50c40d104f7f0851d
zd6d501bbd9d412459dc474e2e77a0b88a411dadfa5f9e30327588311e1e24c0fca2b3c17d6b644
z5a2425cfd702a99c0fa095fdacf0edc17f5c42cf9f1e19c84d636a01932d430762f75ee9067689
z40025865ea9c6c2ebc1f2bce3b54d5b235e1417d6731302e26229544739daee0f4a975a26d0eed
z3ddeda86e53c156e36fb46e5073f91edd4c6477165ad894f68636fe12bf73cd7812793a54a8d26
z357b9b43daeed5c923c760906d7145aee0287e3f7a770fac3aec36ac950c1429e41bfcfa5eb7d1
zf46edc7954f437d2e01f2785896691a094b7f6cc98c84ea9e304d4267d09c7b7d41bace489bf31
z268f9a55661589ee42551d7ab7b4a6d62218220a9ef6584d5706829ca07c4aba5a0fd92097a916
z736471d015361cd0e47f0b79bf25cfdfd7334de812733f7634838bdba67a61d52dd2ae9ffbc5fd
zf4bfe9195c931ccfc010e788b98ef30733ff3fdbe3b80d3ba1d399493e67c296828a779e1f5a45
zebae70807f16a6d90ac4797d030424b3158456f88c8cac0856bfccab324e66624815b9be9c40ad
z964550ecf61faa71b2ac4b2267d6b0a8df08bb1ca0491260655214b4399a1612de9a7b39348b25
z84cd09bce9bd0fd5fd877c1b87d9e0921ca55d936d0382500b3d0547e81aade137898aa354b892
z1911187bfda9976ef101d83e31571f886e8c0736f98e1464a25df0f5b964752dd9b3c65c7f241b
zbbdf187afe95e0c7d93e29596f961a4b1099f83231726a70b0fe1daf6adf3d56831b8402300316
z7462d16294ab4d449618ed9c96b9eeadfa75c3f79105e5a70f1a695825a077516aa3fd7f2ccb28
z2ca31f1483e46d0dd8e0fdcabec61d7724b3f2b082d32426066a3cf4ee8d81986249eac3f392da
z313f38d2f0c4088d9923674f3692525f291c6f7a9e2b6d2eeebf75e0c2fb5ff57deb76cbd893f5
zb6bdeb6eb147f077adac98566d73d23cf9c0fa485841de245ebb4536dc86c7c514cdd348001683
z929759772313e0fce1dc22f68d61d455365b78f8202e67f9b473a72ed4bfe5cd087429eb6874b4
ze4e82739a8ed35a7ca3753ea4bd1f67fc58503a9345f74041c06f3436c8ab55612be11fe4cfca1
z104431eb8053cc9cc798ed62476418fff65e37bd5ac3a3037bc5359704bdf8c8e7981062c5487c
z0fea481613490493f16beceff6305ff0ac2f78d9a1b6fab7024ff5e08feb7e97aa20fffef9c15d
z17928ee07d13ba18925e15cb006f10400a953ed14f99e588baf5d6227c9c8c223680b71352bb47
zb4ac6d202a274c1c398ad0675caee9e10e3735de674cac638abe2e616e3677d0c530dda8d51b96
z8018a045eb81e76ff6e565250ae7af1e98d5f78675b69cd96d7638d7621a690de545324de3f143
z6f66ec98208e2ca8cfb2e12d1f4b0ce3996a76f260174c9e7f3130ad4cff43cab1d20bde930a3b
z01565f4ebd1ea7b2551f5acdb01c246805b0a6fd11bf7d3edff6da469cb10a00824fe177aed543
za07af9c07d4e7ce35dc1de77e3b889703a55be7df25d4870029ef429643b1cbc2610690e56a527
z6042023386fcf7e55f7a2c9820759a78211b952a5eb177584dbbb0f4f3d8e6364620f757c13ea5
z1f7c6ea5bf2f97967e5e1b09cf2e835926d996c3e679e0e69de39e923ae1b51707881aaa0f6935
zca3beee8180da788a41950deceb3802daf91c6b3f8a916b3c0021c9310f184886eff1ccda38615
ze4baaa50a75b9004e6da664f58f3d9cfe70f1d332d7684c29d599ae4b92ddc9f35940d8b6dd5a9
zd90d1c71a00548f3c26c3e50cf689ced57045676efefdfdf5fc668d9a1d0eda436d83088bb5211
z4ab4d1609bdd8597c180d7fa9b9891895bfb5a24b008bdaeb0028fb1244726393c8c61123cc156
z13b4f0c2672abfd46766a7bf382664d9abb6305a0a3275440db1c8dfe29da7c157de27af0ab1eb
z900a68a318739b2c0f3aa253405b4ea70e7d2305d4cbaad8ecb7f63c559810f40e326dcf54fae2
z699596fe0d170947a1f575b76c6f982194931f349ee776d72bdcca1049d9f9564cf443f4ed1591
zbbfd56338d02bdfaa57672cf71d5891e2326899dca0364b5bb6519ba3a6746909a0bc117d51639
zcbfcf98ea6d1764617c51915040515a994bee1c9c04fbc92d516d471cc93ddbc0fd0728c4788e6
z2557539d11aaa673ca7c42b668e0c9ca614c0d1c2fc814f9b48a07f8eb255868b5d8885c889925
z227d3aa449ad8468927588f4b8aa05c934e3ff8f12afb6aae5544ed8fee1b167b1b9123e624da0
zea5ed23667fb994e0986dfe21aef01e43c534110e2ede5dd1c8b4271b613e7945be90816af3bce
z95208590a84ace1817ca0cb4c1667973a329f58983bdbb70c6c0e722f01615ee282c5f04264122
z21f3a7a360265c6a397dc01677975b436dc253b81aed44665a3ab16ab32467745eb3cd80d4a8a2
z85321597bb4e757a6488cf7a7e6fa64a1c32f31a8d3b926e5dd8145d77c9409902ca38f17d2891
z9569863f4fd9655d87d1ee3e9dc889badc496f4ab918e24fd4e37d8150c5519f217fdd7daa9c78
zc3e33acf0fdaad564964d598efc585f746c2a7186072ace9560f269a2302ba9cb5bee896f34133
z2981692ed9675f113cbbe73fbb5b6e091da3dc6ad43b29366b968c543649939d5c8e238e96a467
z0f8405e633fe4e5ebfc9e20703ab1c97be176cdf71d8ed2e57d582c8b5935685b86d116ebc2761
z6be53e5884bd044cc089f657197d063411c1c43bc718908b8e7484d8dd81b954b44f12812725f4
ze42f73d9df93591451ce4a741cb08b8ee1acbbae7aec95007fd1f49ecf13bea5d0459c32e80788
z78b7982187763568c1ea401ef7a5857e8770dc7f732fe2183ff85991f592549b5036b327ab8575
z2f189ba04936262fb13e99656bb3d73bb9dae2f4fa53c2636f34a7d677f0b7fd094d0a7bdc2042
z145d097348ce8f8bd347dfe960f76328fe96f3b2ef8c076e7bd85c61f09d8ed47c017a3b514608
z9d6678dea43016b2722f809e3385c4d94c5aad8d1407799713441aa44fba7b468b75fc3fe5ea76
z963a9a5b937044ef21fe4a98b927c2610de7acff9edf1e1a9f0884fcf5a86c941f7adf9836040a
z3e48062d0f0f60281a12f92173461d786b70d352e070c9ffab9a0d916bc9ec5ff83e67ac53b8e8
za3f4d0206c7bedf9a111b7726fc2d97264dfbba1c439f7c436db46e4a7d94a8fb1947d9ffa58d0
z4c6425a2aa79c0795c808c98ef2c6a6f2c3fb1dbbca1add2410398f44820cd2d4e8b1a419706d7
z18c09eda971442d1f8be1f5c0d83fa15ed41c765d6216fbfc0985b3f77551f166ee2159e51eb8e
z4fefed97179358991619a4f14a7ab5cf71c273f2437374218b34dbc66458586b4c1c1b8dfc0f6d
zf8c419b22f7bec8e9729767c1ebd3738b6d008c192b95b96fdc013fc0b63c8cd07e1d9fa2f4ab3
zf504b4a45000547c1daa29256df69132a6840924c54683edcb306a78bf066f2c4c56d13dc02967
z2eabf8b6ba0ddfb2471708fd464fd5d1ea9ef9dfdaa20604610369bbbf63422bc592ec3851def9
zf6f792b0813cffd8b1bd43c7f578c6de14440e60bab20cc81d54f7a2e23a4cba6b533da3a1bda9
zab39daa2f943dfbb7d36496b0a2f54adddaf534465c0ceba01382233460e2b4cd97322c76832c0
za39910ef05e335ef1479ef12fd9237faa0c2932114a98eff0d5c79bc81ae620c10de2defe0b168
z390095bfa6cd7729561bd7b5f2995275dc367c9889ac6111a205cf9fb702591c1c7ac5049d46e4
zd41a7fe13fef38a86c05924d58fef94ade37d04c94087162861c2d8bba15c3cfd3b007c4b9ad2e
z1b1e34a67aee2e7e3aab48d29106e811d827b96a932ba5311aefadebc0dcbb5c9892171714fe23
zc87ba4ce59e027e9899bdcd629cb838791814fe632b9d32c1865dd7d17c5f61410979e43837af9
z613c24d88b6ab69db344bc4baaac574ec68208283cbc74be4dad09768cd0a2f30fd7b954ff8daa
z7aa82527ef5805188cfc46ba84b7ae9ee4b3f6d51d7bb62d65aa0f8309599a238d962236121a17
z22178284b68c8db8bd03a8e9795d0fe06adb4d1cb3eadab264c599bf6e6a7cddd0fdd5c3569cac
zd23731c98f695b2c2d7fce400e05372767b64701ae4149f3152927cafb3e6106f5bba3da6b10ce
z8e0ade671bdb06726e9a8b688c3460e756aba57b09c893aed3a1adeac0a8cdeccaec928eddc160
z1a20081886b53bb6f0b83ccb10c81da750bed9a3c2d2907672b5a7b8a132db1b473d0e27f9e9a8
z84ef34dbc3d832f111b804624978ad2877c6b7b4ddfbe86c2cdd1e6cd68b13197ecce6db2adc6b
z464d9e1a231875a59f0f4714310a0cb63ac2b2b2a5201edd3daea80d1d3ed535d3b5e50061d5e2
zc2b1956fc19d6d24b70a6af4ff48b8a60bdc1c92f93063fc4cb51c04cd18346c7832a9c26238f0
zfe79c029760245d1a93cdd1c5711a2c3355ba1ba4a8d9cb6b383ce31fcf20625fca4ce6a7e7412
z1e9d12f4a0df64b542f69d1a95d81c162802cad5314d355409c8925bdd9226bbac5e9265066a5f
z3bf94f038a1be138dab6e18d5264c5df4836a9a28a646ffe3a0d09c8f27ea45fcf8b54447b50f8
z0468dfbc067584a4f5dec655b79101d31a383bbd617e8bd377c650b74431cd224d9aabe99eed4d
zf9f7b57a7e80efef6920317b15bc926241d2e13c24a4e0f3b608338af030ad9ce4c1d88744ad07
z62f199dd5b97245305ce0978b0a145d92e1eeb07e3a1a4cf58f7272f28614b17b876e742209459
z6dea59ddbfe8baf7c27a0fa92021e51a8a56fa168f372465bd453fa5d2f2bbb5dbf159e8eded18
z5e82fb7818204aa673b330d6aeceba913ba7fd5118b7a6f61fe8f8108a765d70e59820f53b5c25
zde6b96b3f27f23281e633e2b86f4f975d17fac305960478ef8dfe69e80156aa00bc063713c2ad7
z44e2486ee3ccf556178e5935100a6b3c3416e19b4695abd3d366407f8b25297d24ed1934f2d6f9
z3c500dd86028b33315749e85de7397f0f58a17478c2db0d9e1908e37cdca8a8fd2517c2ccb9eee
zbfcb7e32164167af3c2d15b38bf5f8870a46dd19d7b734bb707cedaffc8be4fd497addef3128fa
z2323a1d95d8fa90160b8cca1b60289b29b75b0cdbb45aafee7351d21a5117c46f258793320160e
zecb6f3d9a43ddb0bdf9e155fefc563b149f06f77f0646a7756c99ad437c8021f8661cb0f00aa32
z424002392eeb1472b0337aefa07f34b96ca8c8cbf368b042446b9b737c74da8fc0944c650300ff
z5da6c41f298bdc3dc2c9a4d5cb236a0e5aa5bd0a70e0d8dc3bd933eba134fb489fff006e715ba2
z0827e1bc628dd8cabd5152fc42e0afccd5ea7f1adc2efe3c37178303083f3fff6c90257a7d3de8
zc8ecf28e5704dbc3b87bb923165e9dda69d0bce97f7408ff5cd8281edce5cf73a1046a28b1280d
zb1a8384653456742f99f573c31230029a41cf8a14993b8058184b9a973abf80fce9833f2a234b5
z66acf5709167ed5a761deb914c2bca7a92a6779b60d7a3f2e960d055f1ed849b868b3d5a4a7908
z6b47c757f36a0bd8d61426a3e38c8a5a659b096fc84d75ca5a85f97ac27bb5b682bfe84d249c3c
z115a7f71da2e8f29c0a2905c4e96dca36def55cfe7468562ea1f8347e67e812601b1291f7410fe
zffa33e8ac7930db279ba8394d2d12d69e5b4f54c32127d0eed5ee72cb2481f7cebab2ae082bf72
z3e5840d1a17f15d2acff1cc63b6585782dcf51fcd27f5bbba0fb219e9a3315a793f1d7e24e8b0c
z15fbac3cc62121e6a39a3712cb204f2d0cbf641cdb7386bd9343bc1b938d66e1116c66551590ac
z70cc4919a155938d859a90089bb009ceee0f416dc92cccfb9040473de32bcd08e70f69dcc74106
z4675c4328b70d4c93333e9f665c14a51bd722c1713c43c80ed6a575515627990ff1d14cedfc0c5
zcdf552f5e5e9a0b992746329a9a51dc077231a5abf412366dd47c126ee50a859758236801a33ea
zcf94e3cc3707ff9bccf3885c0e0f35b3f5d9cc26a473d8b12f03e33a4e221affcd293cc61d30ac
z95bd788eec0e7502fd6d0089550c2731ca1c886e7a65bd6cb923c1bd7e1b03a634126e96045c35
zb790e5c1bf27837fb0a7630e920ef776bb64663a755802776ea6070ff287443e2ac22c2868b973
z62a27022666590fb18b7fea2eaeff0f84c5f47e5f8771a69a43655d5439e485cabb48ba6edcc50
zeb7919370c320e84fcdea933d060285f41824cb13a636ac2b1a3c36e9921b33c630a282f7737ec
zc05339e2d3ed92b2dcd2d665e29ffee83a4d097ebbe4e09cc065660f9c1cb4ef4e87837e02f55e
z19c4bff0699486ff7f9b62fa525943968ba1166681000a825d1464feea321ac5438e7e2173a98e
zd4122ae5b4d65a443de8289d374271763c694dcf7c20a0650b88d55ca3d688cfd5115683db621f
zd8287c5d423a66df7922d6a9e8e82aa894b7dfc9ceef94e6020240f10adabca0037d82bdd85fb6
z929f3030b4e1035d9d7eac09ebe78621e7d70f0ac3c3d08cc5962d26f150a3711f6bf5b2efd781
zdad9a925142030971752967fc5bb16c7d35579a319c32c3182c7001470f7066274ae62d37348d0
z89f3bd015636a4d0991478ce1ac0d628fc1e19075d7e91a7c19b4ebecc53e17dba46a891e911a8
z012a240108ce9c27379e2339477fa4ce04b40d0afb63021920f6b32f4cd3bc3bff89ec0495a11e
z7c811110d17dbab8da891e63f2dd73fbb1f33d00c605fa65c7905d6e4796bc25c311bb58b64414
zda9958be6ca64d519f2dd41ea30ee93937cffe8d3df4aeb63eb097aff99e88cb28b684668a3f08
zab56f501d859d16769a5b7c1adf5f7dad13bb18eac198d4b67caaf1b57c2d64f02c704d69a2ca3
z6e2f5fe13b8b6d72e26845d48ba678a98554e151a90af8eb18b153a28e0eca79b8b2d081a1543a
za02ad4d928fad15ac2ec10bedc5a22730fe42a04888b7003f36b51ac566b5b3866eb7165d9c5fb
z65a0f5ad1d9c6a66265bb10e5453a75c9bc43920ce5ac508e886d3bd523f44c094a0af03b739e1
zba27d23f6efcf7f55c03a728cb30189abb4b7b7c866941f10274cf18af47f99742f40e6e515d0c
za19bbcbf6efeb25d66102591a9ac83697493feda14fa64e8523a0d136bf0cd593423dac8176cb9
z5e3cac1d2df8efdd76f4d0c59db03e482351dfc22a248719a2adf76cff57d616a05ce9bd3d5414
z62fd0ba85c6b0282cfa2d1f43fcac66eef182bc18fbcfa75e79246891669d1d101463b54fd9f2b
z94689b7289065dee760b8d8379f07e3290a82e6fe4a78c9c1b8060479879abe56dae3a821598cc
za5f9a0d9966619e93c0026e07ace7bfcfd43ef30f68712a6107616a3ac897cfb014919cd36d2d2
zec488561ead0350030f39f904dd6460c17f6101d467eaa0ab13ea0e1b304afe437964878fe2976
z468adea1c69a2f8371173fa25d5df60c89509a7b9859fb6bbeecb08f155576fd90568de9ab9778
zc3947bcab9b1a10169dc4b7642c13d5e27dee8ad4a805cdcb0336a408ec6eea0d5e15056ac0b64
z38f303b9c0a9aebec8c3093f0aee549035a751004765a5c942c1c0ba845c8e160f9562a47f733f
z59585ad9f0fb27ecaa26290ae0da40555b6291084f5ec6e18800133bd4d051c75e9d8781b2a2fd
z868c3d1ddb9bc93f72aa0b474ba3d5aec5c05f664b87ff2cf5ab907889066333abd064d8fb5de2
zeaeb333972fbd4260a43060fb61b4acc24331cc072985cea3767c2e2eba9c4427f86c362c27188
z9d3ab30386cb915bc3ecb85f670a3c9a87eeead27c44964aee873a154653c5554e679b7ea7a8d7
z61bfafacdbfb4723244f1f1850873703f6defeeab8b17877aae3e05e9a3181742b4f10f7d51cb2
zb91296c9e631a40ba8b611f4a8600cd1815bd748cdc6690d668061a9d74a300f8f8ded5ac7469c
z7c6d719d4189e487f413eab879d9f297b15d832c0f541f71dbcd3aadf252538cc60c05109d94a9
z88e1d8815b67f14df935b44f8e199f95028f785f0758adee72cf70f5d755a63e84306a142a9c8e
zbb78e8fcbdb31a61aae67f92ed392b4eaf8021f5ff43a1d34d966b8dc93ad92d6ffe6cc2df3a21
z51297cf6d21727a5bda71f9fb393e0beecd74b64773ea0e7cab99d4478a9b8f0b522a91148613a
z19b032c31aa2692805578ab782d488289af0f18c5e8bce77879fc5d627b21f351cbae6e3cec558
z3f809525633d5ffb0ae82420b0b6fe4cfc1d11f6c0372ac868656fdcd1d4a32e01450913c309ca
ze20458b9d5bf6db35ac20ba45ab7fb79dc3c630160ad23a8d520777a17c644dd60b1eac42be8d3
z997e170e19631eb66f2f2f1c4fd1c3e24ac705d781deb554fe393b80f712c1fe8e047895f26ed7
z0b0252f20f2204c308f4016dfb73bfad03baffa4f865a916eebfb0761d69748a09ab7e32cf2536
z763904db352134dca7139b4fa54f71124e9e285516359ab6e49f5d964d4ffa6b1c16e489ec9d32
za57c7e74c5ee1e7ef0114beb8dcbead3f923f94bada2e9f04e7c2a803ae0d94e03c9df9458d9c3
zdf81748d1bff1e094618a17b894a8448ef028d7a9e9edf7d6e7979ad2bbb245ade52a648c3a12a
zb4dc2d061f0261a9138ddc311db40ad8d9aaab25caeaba8320de6f980d4bd96a7d7920250e5ecd
zb8fcb870aca912b94a282529d23fd968bde60100a5cbae9b276b87e4171b80483eb24583118560
zb00dc2a7ada141709820a1bbfc469840ca57458eb7fb4645df9087ebc85f8dcf089ac2d61664d0
z8133d60780c49d56a9161a9f1062e60568b2480c5b99bb18462f8462c0a329962f6f75470d3ea5
z0bec57b96327d264c4b5e58436bca041efd0fcf7a838622c078bba876183021eae0fc4c1b95ae1
z0bf162090e38d34fdb25958e0c0cff28f67c0651e6220d669538974d59e5c25516f2d46a4d539e
za5b8c9f555b44959a251c9b99187521ed8a0fab55e1af2b150b1e5206322767b71d6a101307459
z3cae8de118826cc1fcb4f6e5233a59150beb223c5aac828e9e7a4a9196a98a4aa802f879501819
zd82b07d81b41dc955daf666dca9d97ca40c5afe36c163baa978e2c2f36d240661f9ae2141c9ce9
zdf61b61f390a3d935a9a27305e51a40e22dadb110c498287736f44abdcc07d898ee7e535900468
z1ff9b4bdf3f9c3a49378d09baa44fca49e329b5f331638526ebe77efb3757affd4bb88146130ab
zaba3f5832657b0aea3a665e26860af0b17a8f14afd3981e9213dd34fe3b1ed15e779115a02c998
za9380f614ff55f976d2e6e318bfdb78bcfd762f905e0f0248565fc8390c71b7ee90b8c40c4aac6
z186a4d85f218f2f70a520114240776cf4f975c1a785d5f9f812ede7c010cf044534b7f4a03f735
z9542ba5689462a7fb72f70f534089a1cdfb1e9f7ce548be754638cfb92d42520466e04dc5dc094
zaddfa47ad26a7c478be85b009d92df570248715e5903de079543e328a4590eaa5512a864b58aeb
z5b3b1bf8e532d432df6719c59a00583b7eb8a1b7ac17129ae9a7b879451d3bcf4f337767460bde
z223cbb25b10affe3d0113c165a35b789750d7425d23c507b7f11e59c589a35cedbf1a7bb51d454
z36ad705a738c96164f361a22c77577fb79f3d0be054bbb40af31b6738641dcc3b54a1455d31da5
z7d09a74a627a841c3f3aab2c5efbfba8c13ae0cfa9a77b0c14b250fc5be23414e0db8012970b25
z2668eafa153803974030569c186f0de1ddb09b2edc5780bb659cefdce4b3bd50e3a6bd0f160243
z8be9e2efbca8fe4343e5f9d327fa2ce9b33c7ba3f8e31726079af63338fb9d151c665dc2701ba7
zcd3fcdb668506dd63305d1fb64245d53874536bfece08054df0353a44daf0494a7bd1e425c7b3d
z805d84532acfa531e3844e3e05755b6eb0ddc4e4e961804f93883204b2c4aa947ff692cf96d1b1
z13486173afed48364a0e4e233bd5461dfbb2787baa316951c83d0ff0f041642ea04b2929a3ee4d
zf065faff9b450349e042471a48f7f1c425e4e75b8529552a24046168780359b039a1d46397905a
z016ef608504316bab8da7e2baf8598361196ca761c7ad267ac3090fd70a507b44f2e0a73ae84ab
z886ad7be6cf59d5608d1219f04d21a63abe0b276731a054d151042ba1b0963441eef33c3a16e49
z375d2689dc8fb065f27379afe513820e101ef7b057c5b9c1a99cdc8bd1aedd5d7d0df1fadac66e
z6d3b479d066590e3763ff26f053195c0eaa9f0658859025afa17eefed670c47f2ba24c6adebae2
zab92d8e5fc3b5a0d10647fd6bbc415dd19afa7b198d3d2520dd94a3a36ad9897df4946288dd80e
z7a3038214ce664e79dee4a5e6e3f893ffbcaa39ed8e5f98071075277ee0d482534f57c3e396270
zffd67b10a82f351d904185f493b94f01a56894e313d4ee18afb708864679302dba15cf7180a857
ze796b5cc551cb1e7c68195eb3871de1d46da430219b31bd51c35165ec98147aead588a6f19de0a
z96fca09692f69ba484166ae6727a5a636ff0dfe472f0b409ded9b8d6ead72cebc012ab0d11a41a
z6b7def1c7f6493314d37a1f4537f28c0443c7cd21949c4068baf6047ee9bc93db0ea3ae489d778
zb649f61e0c117bcc27bad84f3ba532d2c87a45197fb7db10c9842e2224e216bfcdbdb24c56eba6
zc89e881c8ac731b6a97e8e7d8b1dfb8bcb4e56e937790184c9c6abd68bb9a94037fcd324845a7e
z6af5f5ac9ca081dfb2d3ffdf98012b664b9ef9bca9d05c46e47c391581c4e2fcbdac33b868057b
z9f1b28029127a7650ab5090ca18e7340926ca0cdc2dd39671423410133e8430b0b8cfa397a1f9e
ze9aa1ce7b475c6e6c5a9dcb4521ecfcf4a7d8f1adfa4ca32ac0d8ef4626a27037fc098c010376f
zbb32cf1366bd500ce530ed0500c3176e6db7836185f62c4911265eb954b614db880ffac70edede
zeefa43ff50f130bfddeaae2902bd3fb85043e9285b92f18d5a695fcf83779d1a647c20d4647c36
z6904e639a1c22c0ec967f439ac1157e64b686fd8203afcfc9c08f0031341c42822be92493742d6
zad59108c55c5febcd8c2d2e7b6c92c47bd902d97bfe20b1a372f316a97030c3c555742d68dadc2
z58d9648c291d77f2160a2e6356d6d5e7639e1f998fbc27a5d602fba9d9220d34b6a8a77db605c7
z2bfec0879b8deaf98281f52940041d61fee293583bf3d81e500f3e8a72f989488351d82319c614
zf62532fa24adc93e2cdb24412876f05fdbc74b41dded8922e5ce1ddccda400359e1b0ab320dad1
z38ce1a3a969290df8bd7e6e4aed0e76ace033df10b6ebfe3b3840c11c1b043b310808b4b22d3af
z4281e49b380c58912be37c06adcc466755a7bca5e550fad2be032c4fbc43be60b625f86a074f6a
za9c25ebb006dcff782c74d6d902828ac303c60c876d27b62629f712e3047e9576f54e2a91acad0
z90815f2d962cd76e5b7adf93ff72694208ed0704215180189ae89cb1b34fdd4b0a29a3715808a3
z9fb527f504fb64749f81658360e55369fb4d6f814feeeb6d1dcf6685c35fb0e1848bb9001fbdd6
z5889ffe00e742812a33681cd43d29861ac54471595532d54188fdd8be35b42216c67817b90d86d
zaff8b84a60312c658a097bb09a6a46f216b1bc5ad33ba241aa1854abc3e126dc90298c9b2dd3e0
z4fc84713b2db80fdc4c4772bd90cee080e441659dcf459869fc6c79bc14fed492933ef22f15cd1
z4dc751652b0ae5fde489348c894f4f99fae94b967f60a6a5cfc12c5a5b0ead6a462aed7833b321
zd6a467b149fa40cbbf4a6be3a48ad1cb519a42b0beb8ee2a208e3ab611d4f0b22d7dec74f711c9
zf3c67565fabae4fdb6feaf69d15afae0053d4173e4401a2926543801ee04828f5fb924800dc8eb
zb97064ee31bc577b9418ef30570d98ee232738799134dd209d98653035c6c604a3a063eb35f38b
z59d5aea0eedfb6a28272f4068da1ce4a60cc9674d936e4f008d7b341bd46cde5b0cac5062c9ca4
zee1168e3d38ec1cbf657e4f5764a43b0e20a1e103ac9f2ad3727b295a766c87ab5829dbbe2cb44
z5fd28beebe4651de54f76e3d150d90b1950f18008175227a7cdd1dbc62b4e167416688f275638b
zae142581fc774fbe027aac1d5fed0a3220b72b3d9c4aeffdd829d15ca3bd573e3de9ea05e801ae
zac266733d268a1ef4da1829116ff8aa5764de6b4b1d7a134b6876c36118b55122fec17b5a96e7a
z6c7045852c3ed2cb585da36a81c1ee43219ae5ab1a3c748e64a5d88c09c73cf68a87e31cc3ef85
z410e854b7575c79ffcf34fac10e9db701aaffc8b82d76ef06a1e6fc48bfe2dc79deabfb1377f6e
zc18be2f7ffe699aed14f6b57b1ca20214a4dd693cd4edf8194ebad3de4f700eef02f4999a1d190
za985e5cbec01b8923e4e78360deacddff70da3e19b24dc51fa55efc6f2c333183d9975b79b1037
z7f95c7e1ec340e3ce9f08a5e2684f7c4c259410edd13712c0dd72e7b8f2baa04c9ff88f7b37db1
z598e6e61e5a33adf223cd27da4320d18626808862a0bfe1e98c499646256ad70a9133e4e2d83f0
zdb71c3dd77e13a4c93da34422e1e97f4b4542a01d6bbd3fa56eaa912b08d4a62605f6641e54235
zb58a27098134e5f8017602dc69214e63230c16ab64bee4d65d303386880b355cec95159a848911
z764055c3b63d55e929e5e81a0f3b30dceba8bcad683cf87c2bc4653e655c0f5ebdf70f34c89bc3
zb4e0bb1afdf97a2fa9cdf28afd3f2224dae785af019f44b48ae1b0c0d36615c7ea0c288192d914
z11efcc55948e5c09faa5379ec7d7f1b504f7f4a63d9c57dfef9d7db9103e9ee9b5b56b2a7031fa
z8e766aa8d0c4890a4a94a5b97244cec638d89a2b2cf0d11c6dd825c67e6146c3121b32f5a1c1c8
z70846b7628475bf9d870870f022f4d082e5179bb5c9e9581ab02c258ef72925ad19497eb513a3f
zae45a2aa114e6bcbd07a0e40ac9cda4705a0c0fc95937e2876ca06ebe14b0dfc6597befd744619
zae7097580dc53b8cd53686f803658a5625e8534a48a287ea16f2a1f10c37f05dd5534aa3ea8ecb
z525a3ce8c8ba22d92e1aa7bd70dd2497376bf2cc0c40d388c09cc9d57cf372c451bba2c3aa3c82
z011d84b7f87523fd23d90739319de4c260dd5098311c86fb9ca206a9f8447962698e884d25f8b6
za76dcc6cbb04d3513623f114e4199771024d75a62979cef1ddc70204129aa5cff8d75df2c02398
z529473b95a1475b5bc2a0ab877f93c2e2259037cdbeec5899d07c3dd0559d6bce08342d7e9b022
zef4de4cc4ece82568bd4895f6889eb4512d0faec79e89b3578184f92f1807953b05553c3ef9681
zb034064100b97a3543545a5c8687c694ce0f8723971bef58ece4d55aff1eb7ebe70908d3c2c6c2
z53c07c88f61cdd06b1ffb1b2f9231f38ba7b45a705c0bf7f3e4537704dda84d64e363403582fa8
z9e01304493dd2f9472029774f970e8923eb87887652824b7d68efa7119f5c40762c835a115f1db
z97d8aba8b2fb03885b17d9905f1afeca6d0f8f7d117c3023ee7182ea87a720b0f0367e617586e5
za01055a3bc7e5cad1e825bb09a0d484c84f4c1bdd92041570739aa886efce697e4947dec17af6e
zcc018e807848b11626210edf8d83b72a90cd8f0ae7d36941a711d1cd4e92f833d62e50bbdf56c3
zae5cd4c2cde0cf315e9ee2ce4fedc1edacc81be424ad885c1fe1eb3860e7421e889d3be2f80493
zee292d932c6f86b0bda3dad4306c8c3c0cee7d08362a5f1d57cd1f95363536de8a8df5c405767e
z604f3984723d88f45a4314e59c9531b28c762c82a25aca91033b020ee9b89dfa6402209ce5d2bc
z24ea3c480c38a9c53c4b07ec6a1a7559f59ef51c8fa7954c3e81df5800c9c52c81c53a6d938ebd
z9bbec154e38c810dd030ba91eac3e8331635bfd36596ee367fa5fceb9d1d74937bac5e400c2d2e
z1ecae94622939bffdcd60ac5dfe5f4cd2b5376e626eafcdfe7fd9f67801e0d70dd0610d8ccf069
za7aeba30ecaee37f05f5b2e03c431facb68ba132db9682fcb500c1ce08ab25e95d3f627f912823
za87997932fcaacfdb4fb3cb0cff71ef3a8aef3cb84ad0cd1db6588f3379f8afb68b9efa2cb3bb1
z6801eeaf29a8bb41809d892587cc3e4fa897edbc9956ccda08198b426faa098a359f554b0e6072
z6458c35c757a1becaf84a70c5dcfa89a75eb463950a941c1ca13f25f01f69b95ea694f6fc69c08
z1ca813dd3ab71619aab5f8f843a2891ff47899abff1550935bfa436d549e23f013dad4c8e82765
z807f8f00bc04df0a718f0c0d36533460c3ef3738be506922e3ce54c9a6e607ed64a5bf329a7c8b
za65a4d4617c05d1fa47f0db449ae1b74cce6bbee61c7b8f289ab98b32fbcc1df1661e362ca406f
zc3e2a96c498e16d3ed436967080a38725d8421d6c6fd066ef7e4d3fa908d5a506320c88c3027d3
zdedd319ee2715ac20a6c242c85caa0a86e91b1a3df633e6791b12480406b039f32034a67d94b8e
z3d835675be2f992695cb137878d8246162d4b0269ed9f0963ecfb9f783b7a4c9ba254572dac0bc
z8e662877dc58a468c05ac690cbb26aeb3fb07727d61426005b3bffd6690688f1d58f31cc10f5e1
z9179d43d0b05b1a7c2acb5ae4ecce88222c06b0a1b3975f66b2cc34797f8016a992e7260f3cd8b
z811971b1c685fbb3af07967a51d0155a30604109b155f5e175b58fa0b145dd59926dd600b935ae
zd88df30dc5e5c9daa2b91650bc08ab627548a0fed1d2157dd51bc78225524de7b94554265d490a
z7416d787975aa86901cc3ec1942d5cb284ce6c8a25e2ad2638de2c2bb930c2bca2a0761c245d2d
z2345008417884c47fab2632a56d584863399ede5fc91c13bff0e7956ca5013e233dfad0d9ec42b
za39f047da2651556a98b46788beae54e181435d639df99836bd57b4025bbe1f1693c58038e9536
z4a426e91864b1fd9f3d6370dc3fea618d513eca147d9b2a3ea2fb756dc9af70de9a6eb5e5a7e59
z9c50c7ad0006f8a35b4a95356af7e2bda68498864cd417275ffe6487c584291c2891604d0e4176
zb97dabe47dcc2d511b88e702b1927a16c774c065f74b5421d4f84f61a64c49083f61a0fcb7e4af
zf9f7833014a5e08eeae8e1c057ceaea2046ce08353dbd763c58d33b284c6d67a879d5e42fe5a14
zcdd9cca5974c3384eaedd0fb08447a872554030333519e023cd52b13dd66d0e8dd1074f17e6050
z38071c6df873414fd0d3d53222c46bd31e5acb7f9b8f8c5500ce83e33621e79cfa5d1179bbbe6a
zdbd1b1e0cf07f15a6803d643e2504653a0b217872b47087d08235491295cf9e7e0e3bb3e850218
z20434a8621723b5cc09de35bf3770c95420a0a79f9b8999ab22f1b5883a48ab4881faf087e1cae
zfc5ed37d3b63608e1bf7ce66324e2d33374f5c594484a02a01b8ba456d620bf77c951cdd78b836
z006a07bd248b8ad04eaee9c0a65ac44a0fedb24277f9cf58e4d1d9e56638ff1eb8a27591164ff3
zfd71ff72f25d21303af27fa78ba107c94abc1c1eac1f20674ba86d52edd8189cff97286cca8e15
zfbadb9bc0fa38cc5f0551b5a7734df40a6893f9e0ec33d28a837c1f3a03ac8e350174898a1afbb
zd38589522e3fbbb634ff21c0b8d097396e0d9a834855ca9666d9a9835cbb5f2f3f56413405016f
z668b57af0e365052331bed018037eef171a357f63fc1e97f4f8aabb4a0e91586a7a48e5e711359
zfd048948779b432101c457ab7adf5d4cabc94aa90c376ca191a4484e93be19fb5a45871f0298c2
z691ace439460c0d326b15b0679998e1a95cea2d972de15f2c209b0a209c187b01b4190bebd1175
z1c849f6a3b7e89c16d6f5d011d82a9f276c1b3344147859d1c4facd18757354fb175f940ec80c4
z29ce7da1a98fac6e02173de424899175c9e8cf180ba7565aef715730e52641b9b0f75dace7b4dc
z920bea5ae0368d73504f28408edf3e3bfe9cbf40074539d10c5e3dd4a8733f097d7ab86622d26f
za768e7172204fe2d0b25906cad80db7df669e8f6a416cfb3f66c84adce14a39b6ae774b9d96287
z0f7ba3ef5b0f243ae8fee81defa3ce74900d8fcff755faf09d9b2d53a017cfb696a74bfc3c1dc1
z6f71fefafe27ce131d823061a650da7f9c834d959cae617ecaabb227c40087f2e7271cdaa7f52b
z9ccd48713009d24deb6b3d30ddb3ff31e282b47c75bbfd274a86bc59489c420da85cf6db2011b7
zaa46c6a52bf02201608e9f9a4d43a76a2ae9b222196a11fb320e61fe85560c8ebc5105a336a6c3
z58e6d30bc717bfe60e35bb474251015c3ed219378ed6f7f580007783c70d21a44034a49c2f1524
z515137deac7e0de02ef5e065d773284744940fe3cb99a8fbdf6937aac53dbd62f1a975ff9977c7
z2f8466fac5c5829dd6374e98be9a09d5011648fb5614c1af139f232bf1baee463e468eebc5186a
z6387525f3f755182f852c6e8b38542b8a399f6a738b6f0a960e0202e402dfc1a264f7d7bbdeacd
z34576e02917867e1097fa9586582ebeebc48de6701ddc15e66b607f05599b6d57850a56098349b
z1b868b18eae8c706b9bbc0cace647c6719669dadbf3b758181cddc92f8702e947219b777afcc6f
z6a8efc8b894ff96ce1cb2f73693209d716c66528688392656f86fc47177ba2778b5c7d7f596a70
zec3307f9b9134fca4c1b684f17f5983b686d68691e45442bfd56cff56d9cd0cf22c58017a4eae1
z6d30d6c2b35cc5c99bfbac98830dd0ca72a25c0bd3b26f9dc0400db504441e698ae579e3887ab4
zb0f5f1c45ab7b909ab9f1f8ae1df357f988c84a6ad1e3cc08bf3594166dbc8b1633e57e37c8f52
zf6e8da614f48ebe2e236a46b7dd43c6f99653b48b965bcc7ee0942192a628931cf72cac8bb8974
z96515e5e149e6595d44b81605450fea84cf2aff754fdce7677640761ef33a77b02428ee705054b
zc4eb87ac0feb6a33b16d2133af8bce1342d1b5ddd34e4ea0e0a96e05fa3376fef5ca4f75beed8e
z86b354884e7e511d9172f65367be11829d41a3f3a0f655a59fc2f9e6a2246aaef9f211e2333ce5
z0d45591197dfb9d0c3432998af3b6333d8fb2c553ba993a59f1dc126935041adefe44aab3aefb4
zc3094bd2408a66481aaf7c8fb7c0f193edba099bfa4baba1c0724cc31ffd42d443811c840c8326
z51d478fd3257d17770e313a8060d065c11c628a77d6f8ab5b88b30fcf14984721df6091594c487
za317c44003388e05d88fd1795f6d498d8165352ae3901916cf4774b140a4fa81b9485b7b84f12b
z69c0488aa37f7ea04bee85e72b43b8d3808dc0214489523bdd81fdddaeb721b7ad9bf6e4b64a84
z80e90b31a1dc3c81a8c747ff578ac5b2aedd0a78d29db81ff33d1bd5957579bd07790c6d51b075
z147d124b803cd32f82a8305db11aefe84c836eae18d0007f39be6310a2ec8bceda8f2c9f95d996
zc034fd5d38b7104845e743db0e21cd7286418daba975fe4994b38f1bb5d66cccb767f764cd417d
zbca6a45ab34836807c429a9d9c05e7481272678f0f6de6289e36f9ff9432c986d331322ba3b207
z07afcc8af7e8dab354f3f0a2c4180d1a3a83b3dcdc6d9dddc2b92db2f21ea0611f19811fc4591b
z5aec57c1ce24822235f26d72832fe6d86df8455501a831e0eaa55d47805b85c7a29e8454e6b582
zd6f2f38b3583d1c3e33772113358350fda6623b0e0a47ca0b49dd0101b1a30891f9f09c8973538
zf5516c378da58b9a425c88bac08d2a13efa34b9516115bc6520c999c032b61ed1d11eb5493cb0c
z1978ad6d62e30db0f281a611bfedcba7b6d1e74e504b802414e7d7db8899e0df32575dd9e0cf56
zdd3eec9d2345453810203728d240fb99bd309132405d8faac33c2f9f3dd50d7ff9af9977278350
z697a4a905bd240cc7f8f6a0542a7de3082bc45a1dd22f6d4e596647773964816118649a560cfdc
za967143cc26d192f5d8904ea55e88c1b507b7ce452fa36febdb9adad2b6febdfc084f8be00fe5f
zc9ecc0adf03c81a972e32fa74f77eeb366c3a5d61ffdc6ab82027ab28eab98fc3277aab816ea87
zb0933e27673329d99fcbc86d9c8abf57dc5c1f52e5b3d1eaa64bedd15103e5087ffac30313d60f
z98e1fd167ef581b949d4187f27c3a69ece900fbe9164b358f69655ece2456567d9a3b1b4bfb994
z7fefd5cd8ca20bfdba04a780d67d23497f35b9adcff82b5ffc7354ab4791018910d312367a4984
z3666ef4eedd7a55ba2f805916213e959c1bfbcba74ce9b57417f5c924124bc774979b673c8989d
ze943a287cb5e8642027c95b54593b9be897ac130570ec7279d1f07f0b72cab5480c2111885a51a
z1ff154828376b8289bcc74fa765bb1d8eaeb622222a682b86d14578816716b0aa34b9f4eee7965
z6d200b4c994dccbea9409a800c9163c04224d4cf01d85e74e93c5e8346536af367d2a526ee0c1a
z7018cba0b19d7c4841b6cae211733eb9b8995a828ea68771dce1278a42c17099af83ce46f8df4f
z4f0130c23a108b6a4207df65e03bfe34cd56aa3ef6334b292099fb27fd43d8c77200067f552b21
z9da7adf3609f01826003eb3e1bb692fa0670ee7bce4e6980f3cd26f6720fa842a816bedc99ee4e
z2eec5f3c6cd1afe333a08b815c25e7703f47fb939008802625a0ebbc6f7987727b8ac0effa4cd9
z0d73eb042857eebff1b1d9a0907be11217e825b18f29c71a44ccfd8046f17091e6cc1a0cce7175
z9482fc5f8dc2cf3af87b773b8a416d4904685e45132514f9ea68c554f741161c4d36f7c02195db
z1536b5101d393d0e84381c0709d491412ff0356d76aafc3096f7b91aa0a553e6c4df7a3250b2b5
z063656f6ce22b3a37044c61a44edf88aed7fdafae47b7770f85b48621a6eaae129fabb1c2aa754
ze942b3d7adb803abc2f6e10e560c069488e685f8a1b4d91de355ec0d2669f95b4a924f787ab0ce
z7aca9bac557c90804f2cd3aeb29d0b4662a194ded4002531537a09b26d3aad39089284156bc067
zcb566c26b45cbfb28751938c8b064d46d65ad48afc57bb2a45ae2958800aa6bc059eeb2197afd6
z0825def2084a46b2c0f501fccdde21162320549941e6ff27c2e74b21292ac9ea51a19af2584bd1
z5ea584024bee72124306cb08eff8c07bf292e48dacee0710c15b7fe68e60e76e621d80c6293cc7
ze90c7d7d0df1fc21a577e3b18874eca95530ced7dbbe19ea561ac0e64272abd068020241d067db
zb0d20a85f0c9fc713c21a0665a91b6647df6502be8c816909d583b7ae0268176ea997fc1ea06c1
zc63feef9c83087b81276dcbba5cb450b1f3d23d670c3cb70dd22dcfacef6775223cb620c05fb5d
z055361449400686aee53793bc1a43ff8416ab927fa62e76e9df21b1758ca836aebc5e835f58eef
z1b3c5d9b95b18cac1c450abd2d299f724b245452b079c994c96f2ed0c6f7a959b99379251f195e
z9908032ce5d772c033ed2b72f6f8548e36b48b2841bf937e63a4adcfb0fc27d1a57b03b2fdce4f
zfd55873432e49061a17ffa68afb92588f828123d5400ca7d33275ce223ad06b4e8be3feb486de2
z11facaec1bf313bf6f301e76012fa43c8ef5251addfa50db61848e8108ad9288e13ed7f3159a5b
z587594b76e913973a03ba9eb11cb05d92dc3ade3710ec4cfa0a39be8e46304a0a723f80000f7b6
z4f25375f5eceb58642637be63f905160cb230293fbcddb1c8f4fb63560c7d13b820909f2987a93
z6b52ad14b84c0efdd80b873fd0a6de1578fd74107e7553777506d90d27a4cb8cc94619623c3477
za7c6b979b71fb27f1ddc0e3b7aaaf50599d1103cfdfcd37ab3f41edcc35c83553f38096e05b179
z065ab720eb852aa572d0bd7ddd470c3f20f50f9202574afd8f58ee596f7f4ce502552c5252ab35
z2730f98aaa725b717b9ac0a392a6e27d61924397e88fe9fb09505ce731b74f7c1177fe20e41702
z0c8ede19027d67b09b3126c2532e31c5bd48b452143ceeb0065adc8ae10905c0b323b427b23137
zb301cd854f3d6ea83a232ecc3d01b9d36e124d6bd048109a8a9e4092d2bf26dadb6b208d1fa4b8
z8ee78cdb8d3d6563f3c5976c4e4a14ab86885b031731fe8de19347387048772938a656b3a29ea4
z6bc60e2ed677ab9471f838626dd333192012ae55723386111aec0ee7d52733f495c6ff2e3aeeb2
z12d34693d08ef32dcb94dc7c927353cc933501ac833cb6bf25155b4083c05a0ae29044fcef59d5
z051f7967edec8371f00481c27271a264b552ccf736abe80fc8b66bf4f5ce041a2c1c02b447d48a
z10f33e213e91ef9901f91e7c5ba0282517c7926591d03230ba1273c2e94e6c1f4bd94b0a46e7b9
z8ddeaf8d39f8cd8204e314f968e24fd8e1aa310448ef79e0be7638908e368a3644f821b8a152a9
z9c93d304220e56c05d35d201eb9198a2340ad6e7a1e144fabf8a2d97ab1836c5e11bcbb08f4420
zf6ed1ea3baf7ad70d3b410b97f8634820489f39dc7b8b4af010271aa4b7a59737f32e33bae63ab
z9444031db3a0a469e7be767ee70d099d9103e36412b40436698ac113958f8d17f936d7b1aef17f
z87e0f86a1792b9facc9fc1edd29e97029070121b9ad589d4524870661c129fccb86410c2ff9787
zf0ec587bddbf5bb674bd86d6f5de6edca8642ad0f2b744e56216753e7ccb06d315f4bdbd40aef2
ze98876c79bb2cac72a5904ce0f63c99297ca40076705c2940ef7cbe70867251f91fa29d2f16d8c
z8fff473083b8ae6390cbfec833ff74ebc86c83707589b9eb81b218b0a8da377ee1ad1ab182ab0a
zb1a520cd27dc75db43b66b419fdcc39b9f20abe5774c624de54480b8086b4d30270fb6bb1feca5
z9c8c4c25e0350466d31d99a5211590f832795d207ec9f4ab382b17ecd07f4b16b917a354f38178
z23de180f554f61d2bbb3a5aa73afc113fd72abdb4a92c28c466de58dad404643ccb18f26196a72
zd630d532f66f71fd536e8bc8196154ef394761d705ab594a7e20f07beb34b86267695ee566d555
z0c9e590af8c11df551cfbd8045a47ffb3217474fef164c5ef5d72e17ebbea1bb20b3f1264f44cd
zd3e7a1271a5591f775eba25c8a18d0786e614c1943148dca29eba8d0827fc5f99a8dc7ae13df83
z5b5c67d558680bcf06fefb8d1740a9333717512f0f6a652215fa1f59f28353369b513b492685f4
z391a91b8cd9955bde122161d06bee79f0b80188142f5a013f6009c3277dcadca73799972564183
z3f1a9ea01d724c7cda1b6ff662c406de16239d58b9e6be840ec43437f66683bd8287343b7696ae
z2c3d24d964f531bcafff1d22511bac1eb16488307a184d5e6d55129def57431feb16abb94da70e
z6b7a3fc65ce64b815d79af0493403afdd9ce3642ef91cc022d5dcc72aa4e5dfb8068cfabec27b0
z001ff718a5c567a4a7def69b05fdf5d5ade17e54b683c15399501b8608dcfc0ac4d55fd35e14bd
z8b6cdc92ca5512976494cfa0572c11e507f7039ff42a49c6514a73f513c3e2383f708ed18a433f
z68fabfdcd5709ee64a1ae1911fa39316ff18d6d7343cccfb9d8e274f94737c59a983f5cecdb64c
zc180e4503f5128af518832d16951a06a38b563b986f807d556db2d77a6b38c4638435e437bfdbc
zb15c275709fdd3b77b1f8ba8a802e093ba618daefb25797ee6453db783ff915eb26c5d629a1cd3
z9e584e0df2361a6b592f5de198dee563e984560f8f0f4274db535b1e7c7f66a19afb566ec81230
z7a7db1973a3232b7be17b70e75afbdbaf13f53f033992cb0581a2d71001b8e318f0df2b7d1cf57
z9c81b2b37433cfae03ce5005d5473e6c94c17366f10ae8dc3c519436ec15711b24b750b0bf5521
zb8ae1fef432a319547f87ff3590912d8a80a413877a719531897ac1177d4e1bc9d0cf6b5381e13
zc0e9868723ebbeff4239edd0ae901157d06d54d7ab4a2030b3b8fd4f850045e8c5d59581f90970
z426542e431223583ea83328d599212fe0955584392793314312aee510d9fe99787d81855565d75
z3d09792ed34b357edfd22bf34cb92cfab17c2145648bedb642708552c0471a1d2fe1696b23f298
z6b37228dfe2bd00c621a2019afd4902f311c42f0ac0c94c146a11b824913c3ae6e72d4e876377d
z4b8e85bad7f8001e79cde69949588548c8f1083d7b77ea0fcf88c96ec216fad7267864dc7b5622
ze9a4361ff9357257e0486325e793fbcd46d4ecba2001228ec2f11bff6855eb59d75c62a148c2ac
z7a297e48763e8de97c2c7a59656d99cc6390542aba7ce20ff642139cc585bee9be294063602f7c
z7da50a145222fa27f0e76b7477964e340b9fea3b55f9c58889480117a8f3a2e36a38e68dd2e058
z1ec89b069c4d28bd86690026b8288eb623dfcc6f9109f1671d84a401906ba6ffd9e99c33f5c63f
z81d37be5f8586cd0be592c86bea16aa3329452a2a11f654419e7fee4a03c2cdff89d425bcf5286
zf7a142cb17dae3fdb4dab65d055943362bb1bdbc88e21370ae35339f1ea81e8be3529b5c8edb0b
zf9243f136b6f4c3ec727429876bb1b3707371c7b298ed2cceabca90f38d4d6cbd2018d55a24aef
z792a83873901f8fb541241b4ec98ee780bc51b4c2c17ee11055dd13b9cc7032b217d658c544a5b
za9700caf3eaa6dac5fc8b915683d47687c0e324f4bad2e34f5ff9c557a22c9faa01008a28dbbf5
z9beddbe82c0b3eb1e6c5365aca1d06994190a58e5b86140417a889bcee22643d99cf3b1cd6db38
z23882e0c907a1026012beb8a5f9225c7c4c5cefc69659810d79e3bd33b70f122db99ec3df91b21
zf20cfe78cb815f5078a9c5528250edbb928a373afa93748393474a2f9558e322be6b9391953a52
z990b00d974c6c3936dabed3d45147047f572e8ad20f1d0ef0ba5af8334486c376ba91c1cd21049
ze309c6c564983c861f2be3e0aba6e813556f9b48d8e5bc591dcf9f37986dc0d5b7c020f262bc86
z36d5ee9046876f02834985a6c79b0e4f125e880a1533eeee21d6781d90d7ab36d7be2e2ecf2380
z05be09b7f10c03046be2fd52eb520816ae51d579968d01e75c4057a5548f73307214634a465110
z824fbc05e49cdbb54dfa87441fc919d27275c15a344d22fe4d6b641c366a184d29ab6b16b49517
z597b0d6c3b140e0c34060c40f76b85dd920ac757111bcded423298fad5c2335c2a996822194fbf
z7986675c0e9ceba45c62bf4b05fe1d36730d3c280ab340fdb91c681ce572d3fc90e3646e7dd5b2
zf4426adcd67bf7f4d94dc94458a955d51d4234691e7cc3a89718197616fab33bbd757e55a0e292
zb9007427838ee8bd5d3dc702ef7069ddbe41c3715ad7e3acee5c8271f2778b36ed135d6727a033
z58b968611c99f948edd44782084a12b65d584c3015a244e982d4a9b747bbfff925e07cefb961fb
z075b742e730890595a486c6673ab44e516f155be59a000c6310b9177e07a8f02a89f7f6b90143c
z90b4a4b158f517580d7047e1d69e5c145d06764ebda2b999efe4bbad38571e668bbc444a16e8c8
z1a4fd186aa8002b3024b6fa518c7e872233ce170c8f900d9d0ead7b83dd5663feb53492a9cd2b9
zb97265936cbc173157495da94f8da68bd9964e7b59bee07695f43939f928e08bdbd1e27261edb5
ze295bc7b58e0058338c7f439537aff7b3016009dceee15684f4fa74074bc8c97acbc50eb9852e3
z3fad996e2509740eb54c19a7a229dfd7a42a69ad5ae4077243b3e185ec02a17351db72de78b682
z01d468998f93da2869838098375bf50ad5cd4f05187054e6df673bb927765ab0af6c73fb09ebbc
z593bb6f7763d7d3ba69983798ca74f8b0bd1a302675057d519d78c0b3c77ed97227970de6c96e9
z8c492f85cca27a0f07f42d5aeaa1c76234f717dbefe3335b44bc1a193677b76cfa3f0044b28c0c
z6188635cd8ae580bd28397c3688dfcab384d375d47a9330d7bcbefc58111855655c50fa72c9515
z2ff39e5032713d654091449accf82b0aa8bbf2bbe2848a86a0106633993d9a30755ba9e00384de
zb8d068109d89473ec3eaecd92785ac3fe769f6b936ebae41eb8f7c90d9ace45c0a1e9917cbf83d
z9302580207f2bf82267b8d586994b43dc0fe55385872caee98c0a9be49af69b18816e2cb25d46e
zda895c8a8ea4ea6d521f6a420617e289e8ee8eff01c2813ccf1321962fa6da62484965726b5e44
z12ad65cdbfc2ccdbacf4c2777f949fd538d79cfe3a3e05116f740328685f5dec49a376dbe911d0
zc8fc071cd1e7bd1c822a143c4e95e05f59be0175308ffa7ed42faf8a11d122c78ccb2f93c09bd8
z9c71ea06212f7a104e6429252152c0a4970327f8858c2550ff133174e6fb001fdcd2dbf823dfee
z31e9aa6480d2b2ed665357b2949d0ac6ccb65d57e3c0626d8bec3737c43dfe64beafeef1ac61d2
z5cfdfb7f40bf3a09442d2019cc23c5ebb5039e51bcf1668e131e95fb238dce33ecfda9322cbc6a
z70142e431ba9ca3694aad2f849836de4437f9226c7b9bf33cd4057f88e20c022116ed4eb49b945
za5d8332c30eb07b4576b1d3e8a079b51f34ebaeeac951ae3c60bca59f97ca8545349dea7cb1560
zab9a967f3de23d44adefdc76bfa80d16182929210eb05997e03fd31c959cfef9be51b910318eec
z1216b0ef7da4c6253a9029fb20254f2f7049f047aec43b71e6196c44120014f84953c882f10d9c
z19528d9891c54554c0d53320fba958fa1b8b07220472cc8e57bf3dd8a6500e8a7079a5c61b2caa
za0ab587bc7d32c2503f026bc7a7a926ec9c03f1e634fd697ffd51bc7909a7e63cf8e7dd4f7acec
z43665ca9ee33efa6f97f6589625db34b50aa634f58dd5e41b9cbbfc56b347bbdffbaa9166005b8
z48d8459b925b3bc8d6d69353e78ac36ccfbb5df9acfddde76de55fa70717dbf62b83c6863f0d45
zbb1c998c2191b1baa1094709fc12485c057162be974a6dc0fc37ff0bdbd3ed7a6da344f7df627c
z0c6b517daba23f8639d2eeccc7d335843e8cc418447ca86ee9f23c5b88f17f522a8b289ebb3375
z9191c4a5b7bd7a5b2d485dd20488c5cf94de354a8b1611d352f0bf4241aca526bd70d314a79378
zf6b138ceeebb18d75c33c13f741fdd7e8b570a1dc2e06d0713a2389b44230034330a8dadef16c7
z39c456f6d8c87cf96c47229b21eca5e36acb510ecb649ca5efdf464d4d1f24b479da9878ba6260
z9458077f079a597a1ddc1d39d632e7b36945b69d5a1586d59e192d7a36697da61d7beab439e1f1
z8f7d22d4b1a6c7db963ff42d56481f5da7120c9c0957aec7768c3cfff12c7464aceb03bd8b3a51
z7061d9572548865b8999ea8bd881d9091717afbff74c02d1237412b0dcd1fe5563421bd88eaf74
z722f27f27772027c6b80a98235617de68e4f642fe642524a193b27c8204d9e4d85ee3fcbc1a5af
z27d0e3f03919d5c408fdf11efe4c3b16946a235bed75b01c926acd602f3b10b839f36475d1c710
z95ce4a29b8d6b4635b124e0c2d41b0dbe8bb77247438a00c41470168b241e1d3a959ef30b7e14b
z59f5f654d4df49f69edb0b6849df8845cd5db9fd9e300f4db94c7f50cdd6076c3beabac2662944
ze85318227b6b56a0caf790e5e08b833d36566ef10334cde9d6eee89dabcf0babb257019c616987
zc6b1c6a39f7e169240197f031f7ed81f61edce6106632469acd89ee410d3281084da5342995a9b
z9a28872b05cb4d865037faf9758f57fc2a84429e5d4939155e233d9e687676cc221ec576af77f9
zd4c7d7edadfdeb6bb78f3238ef1f1052b9dddf75a89103f732cb08faf259ed28bf85059ee9a56d
zf2b1d3453de755afea4d9cb41304b03eb8f94c7385bf58bced7ac03b474543d13087dcfdd43df8
z463f322e249f806272cb197479d0526b759a1ab4e8cbd3038920614257d3c39e1ce0038bbfb829
ze7aa912947da5b2c69ccdd1bd09ada846b4889599b22a67b4440eba7dbbbea4cb3d2d49def42e0
z6f9034a06c61cf9221fc007bd8a3e12604e14fda76270f4956a0665ec4f8eb813a305ea36e2343
z781bc4a306ceff9d6adc6222f79baa30938fe1f31386ce6f6c8738a23ae89180b67e811c75ca72
z93a6fa32d923d70ee2b210dc012568afd8cadc1d796808ea2d14a6409515f130b9e6c219d8de4e
zae04c51696011677ee2609f0bc47939b8962126ad9438090af78c45a310e17e267b7529f570074
z829c076dcc07b8f9a6a68446acf02f0e3dd2608af3ac441f2a0941f62a1185d1ace277cfba673e
z67e322105c29ff2f31ee456920ee713c4cc395e91fdfc8661ea8acc61f885a0d7c538a45ee46d2
z34eb69e5bc2abe61765aa20d063ff1f2925d24dc4b4070f541ca50badaa610b40daeb3df0fc574
zd965ff478c8b6541aea86985b93452e153025dae69a5abc29580086f04285581263c1542c7268f
z85e7fa0df750ea0ee14daa64c505196b47b758e2038928bae64962027eb729b2ec575bc5c389db
z3b09cac4c92f24cbfed5e1a7542da5a00992bdf3a392fa76cc8aba402c559ad3a27d785b46a446
zab1a7e377c8783031821fc02a995c28ddf58533aa2aa658fa7c6f2441b83642715ed1419605fa8
z0e672b58d899ec5605c55cf76e4421a3cfa0a42a2cc505fe2a09b20ffd71d652757f2d64a7e534
z50d0bcb6c55b2c739aae06745337cb56028235a479761db4c829f185d6bcb7f0562efcbfee149e
zb9f12092beca12e1ec7dc842088dc7e6a6f14f36b31a75a92d8b048d14e9bd1e7153b23af38b89
zab2766cc835e58f1c0ec00e87113bddc8c6af567ca78feaf6e81dd0d7d1aa9314f336133433dfc
z9c3e81810fba0c23eb91f14375c8776a7ad1bfe0f5ddf46953473b39c0572a7b7d0320b2034505
zc9daff3a1c6048d7599d6dd1deae6da682d231e31240d5ae2e6ef8c96eb789000c5933ae708baf
zfb5d395d5e1cdb6f8d47a0dfddc3729e3b19a66a40cd9f7bd2982237bfec5ebcffeddd630bdb47
zc4fc8cbfc37c2edcfc5be6af79d855d95d302621c1c65129190f5930d7acc5e324a753cfbb9463
z7b2005bc1e448cd68b20949de112b4d1949f66920996783377781472f2dbed3685618c314a7391
z11f58e3cfd358e57c5da94e4f6861fdb0058c1ea98f1e35c00a1de92945af5ada50780170d014a
ze74318aa1919aa4fba87df60473ac3ca1cac414b11761f2cae919ecabde7d8f7f2d5509e72185a
z1fbd5ffbb42e016fa361e4cad2cd69695f418ee2b9079d08d32717bbea0257f9cf7a208e9ea132
z9330f0fb33db8e4a82c2aa45b1750a33701bab4025da78444de8bcad35c59930fee24fd564267c
zbeb8f55160664faab9f8fd0d7644ae17019c1c40cce10abe35b5907eb7d5d6731e1d85cf809eb3
zac352df4bf045b96ac0fe7f4f613ccc00ab5b3236245fa3ca4ce40f89a59f280ced0f05aafac25
zc006417e64daf4c12e23f71d446181ac3e231e7781e468722a2fa626612d8db898eaef8a755c94
z3710cba4201e64ef8d43819a6182be865db1a1d9f8b82bcc524993f72c1ea3a659e7fddb5e6e3a
zcb94ef9f671e44707e0769693251fb4283a351cf0336ab504d82eeb1c3f39cafd01a338b5c6fca
zfa8da4a0abd859994e54a1fff7c1c60528f77378635c9e1ec7795e1602ad4e50451309cdd8dfde
zb6e323424273b4264c504765f01ab15bcd3b82d6b87fa182e6d99fe65cd163df87a268bee37670
z1c2fdac3d6f5a2c254f75f79b327238bcc2231c028bbb1ae9e9279d908a992f9f89d9f83503287
z60c5f8618ffb806cba39d7873e617af9854ff958ea34c9269f624102fe3dd8f984cc132f80f5b8
z18eb5ab4075c1333bb45a9cfff3b19945925dff4753e353dc63f73bafc4ec29b86c935ed949529
zde4230908896dea42c44fec999deeab24dd08a1388eb3a7eb95a21679eda9950fe72a88d604bf7
z769735ae74b4d2c3e6a9b7724c70f277fca394081efec4bffe4b9536df45c89015a8c933cdebdf
zfdb5b4d39a8ee1b8c2a630d1e80ed4d53b80e6f8d5ee4f3d5babeb4ca4be5d6510b282e38eea0e
zb579543c35b4e381df09f5b184ff93c83b0870b7cab7b23923f33c8bc619e7c29a01098fa71072
z206e1cbb42bdd9f78f09a3c702c58877a27edb4337a6f98f9733c508a821f6c4c63692ecf488b3
z19ba092ce04bf9047c2f7f311fff086505bc1b875a149129724aad49b16f6c39202c8b96ba55ca
z2e4dfac22fef04df5ece8bfe55b2714bc8f711cc2f6bc725a66c24f95e3a1928c580f2a5792a87
z3f9825ecd79cdb293a6a4a9ebed80148742d7916e8603cf19f2234a5a983dc1b30ec1f5b9603a0
za2898ec10110dffeb4046f5adc106819c643bef72b19258ba4d4ef4c67ac1a8b27a2657c19e101
zf7c8cbe38b9da40ecb99e0e5b31809f6a01f47025d0c48f22683d616a1c07f9dbb7ec8b3e9d529
z9f844f68490169782a1d15ca196e40c82c3de7024a9b0f582ca205c230f711b392c35eadeb79c0
z46f75e7a6c8415b345b207fff314354be20131b919c835a9270d1799f2356e4a835363bb4e1450
z5ec98d6c1fbc54c71ac36537c9739ee559659839fc866563279151c0cd75f1122b0b660c15dd89
z81a2e83e6625ecb9d354e9f556920b0ebd5cb5df7d2f5e4e75875c4ee67b518cbb69d0628f1c71
zd870c46946e36a4e57c3a84bf405e76aa830b2272f26399c9edeb29cefe7d857377bbb350b0337
zd5c644c996f3bd48481d268045350d19dfaaee5d590ea3d64108b6536ad4eb06d27702fccb5291
zff1cf91707f493a6b35f5e99de4c3d5c39c724fce75eb1561b008bf25c0800d88d9ba545cbed2e
z76ebfa154911dffebe6091037c3dbe19eff933d2463801c5f7ee6da9c140e7645526be512b400a
ze86563caa0d18ac5f2b2ababe6b86ad5e4d44f0a1dda479b51884784d66cc614c96e6cc9fc22c8
z38f60e4f7db38cb527f8909c6b3ba0e6deacef309a55171f1613063309271e824438e12535256a
z6f41ec4f16c8847eb9f96c20254467e1ce49c94f2f4642031a70d5ebe95724b496e3b0f3368e9b
z81635fb29c547d43b4cb9dbb71486582dff1fc5b6c5cf5e2bfb61220e176cbd495685e7db60ade
z0f2f19f3e3b5b0d7d7f4aaae800eca82fb24eae371c0c01415047254a09ea5f359d77af965e827
zf1281e8ad5f33fdc5b44ef5b83161b60f5b4ea1391e2ca79dcdd888c90b9d3f30b727ece310de0
z2a05dd7124b19cf40334a3d711ff1da3ba18d5acf729a2dcf9b88cfb08e8455eaa286eb9684cc6
zed76f2dab51dcc14f3eecb3e5fbaf4ac59bb15c08a14bf740833e631326742be6bbd5709fe231c
z578773daa744ab42ada5eaeb1dae925f2300ee36814417198f91d6f28359a26d08a4590669b0ea
z0f4e0a2f18eef2eb6f13d6fb824632b906da7cfa8e8e3e37ecabd40c32c3a551c1f5bb73284698
z22074a172b43c8410a494c8ab561c96cfb6d17902cd178a6c56bcbaf326c253aabd044e17b94ef
z51ae4e164fc4c9977fcfdfa9f511c650a076bcd089f67126af8bf444951251e3074c03453c0052
z3e1bd3de522fe663cb834d6e79df88468979540ae8b06e870d0569987a616cd5b068b3f3a71505
zed05ae344ce990c0446b8fa23478ad6e83d1919da8161704a991461ce67ff811d25e57fe936187
z8c29683d9e3a8390939de3e4c3ec62f41b5ae6e05e1b2429b9f8ae1f5be348da259214cdb26baa
z06e5e94baf1a0f5212acb492310071fe5919936dcd908031fca8fa6e54830f0513df9a325fd1e5
z951f0cc498af15eed8e99392535439333913deeca0995a26d9821d5060ce7443c981106f7f0a6f
z35c7db8707df4d95faf8a6a8e6c3e09ca40dd14fbc4ba614979f6e52e97f87e22a3d79cf7cd5f4
z2de2a08af013093ab5afea4d8f8056b174de72849ef2d6cd158c86d6ee4e2b149a5a07a0ca5a1e
zc46de3e10a64b76bab4092c17f41b0325be306806704c0752da633f56fc24f31b35d594874a42a
z7509c37a61ac3f625e2b915c4ab87b2fb89a4a14918e1a17e91b6d570525da8b3f3841ad66701f
z28ae42ef593506511565bdc2878b49400c18c6b6c7e168f2e640afc457882bb1b2b92fac7c97b8
z11e29729575f1a904bd42c65a236df7aec31b401900faaa77b96efdda0a073ca224bf51654022e
z82314ee110f3887e18a7e59647c8d038d5bdf08a3c5f2b17d5b1b937e1f0eb48fd44410a63caa9
z4f8ddd6fa20bb30fd45e40183007943bcb14e32afd925e3af566175859185da843e4da7bc8493e
z6b488f8285fe6f6c8a5009f7ee7f228d298a6581180fc57b03f03190954c631a98fa86b3480b12
z9ef298f4675fa3302fae8ca4cd6da548560473553681f7001154feadb96580323c533b1006b1c8
z582d6a220bc01fff5cd9e13a54b081ca17c94bb04ac586477af805fdef19e2707acdb0441cbdc9
z499281ec51b9c9e25da5b81d59b437d75681f204eac14ff2c12d223b65453ef0eb00f695ddaf33
za8702a1b79c830a24829039e21295672ca49db11d0b5b1f508e7a65cffd37f09926a945f7ae2c4
z23e85b4f85288c6d38a854de9f687a442e90143518966daf329000986e09404af4a10981f076ed
z5a67b9d1e494daec63fd54107e148c825352a0f7126bfe6053ce05f225b78d82614a3389da5160
z1cebaa2118033f866110560d8fcc7a4db141928a885e731a47971392911e7efdf619e80ceebbcb
zef1f3c8a0d8533967722d8978fa4f527ec54b83bf77b28012184bef8202d206ca975e3018e7cd0
z30b7eb864a6889b727c26833bd7fb3c69996bec8f4686509d31506c45b3cb01a20d231282f7d9f
z981876bd6e2f4321f503267b22f5d074b2238c34f5163358cce1a41f9ea227cc98575805cb8991
z9aac1643136b8bafe18b24e8f37102e10a49cd2ffe871f69c77d343421c60d88cb9b632e26734e
zf3942afef9f7429e7e1b6c2469a0b6ba270af2f914bde950fb137ef3ff22c174739e0d60941793
z8706a85dca740c5273080ce7aeb90b83354351ae0e7d9bcd7996439d2d9a8bedf0eccb80e2ce1b
zcb4b4eb0f55333c09c5ddcb6f5f9b9c91a1e55ad8755db3c9d8df814ee4bd4df495b826e109408
zdfc07cb698ea39ea7453610d1dc956bc6160fadd7a5355a90eae682695182b98eda01154931887
z13ae3fbe5a0c3c990b08752bf2b8a1d2b46d21f3644f68ba97af63eaafd16395d3ab86395d3bf5
zc265da5e111ecb18907f17beb7f4e53d40af5afc6e02f98d12416df3766f38921278f84949431a
zc74b9d64e3d3a7ccc6b3f6004cc4e0d89957f6d7324eee9e8b118faa065fa6b70df932f0327c00
zd3dd1baf7d08767b6b0f109cfcd1884897a15cbd70de4b7954cfb5ad9d10a7710ef1de77ce445a
za1ff8856a04b9fed9cfa959f4f6b68b3ad1f85520105168a323516c1e193c604f0d6584497af70
z6fb33e84eb4dec90a0e5957ff664ae406a18a8e47b19e1ae75910a615ff97a4a4c0ca8029d02d9
ze68efb6fb69166a267a148bd93517c182c18997ffe4be8d075c69b31e5fb21323f9e7d7da268a9
zbdab713452733bcca8fffa6aa7a436e67fac91c21ee47a75d79111f8e176e6c7d96c116a0ebff2
z2d916674a3c40adaed035eb233e7fc0bd8249ce26aa4fe32a477cf7d09bc9e6d68e9e448ee4530
z57d536be7971c41df2b7ad1bada76457bc664436d592660bd7fdac414859327aabbc5c29c60eab
zdc9f9906ca7d55632345aa0d311e76a90c173022c3898c105c8eaf4c98e1ced7da273e8a32f944
ze4c322134bb1d31eba53e66ab9bdecf0b170c5e4ede74263ce71c9ec51524eddb0cf2a6c9b667d
z20b70194d33a59b6e18448867b4daa3bac7a71de85e9c88255a930f2860d233ebe6f3789b1da16
za49ff0289aa9c38c76d22d12d3bfe874355ef6ab8e426d5d9e45ba66599196ddb01e6920086a03
z3547afd388f1a4eaa7eed079a30ba0d1c31b29847da746e766ab7f6cc946af9a72689ce6a51b20
z3a29abe411a8feadaebbae85ee05941b4e7822ab86041c5df8d3f94449f470fa413b18cab25bb7
zdf01664176b6a76498f25c6e1f1b5101a0a501627b98226871a4b1e03f9e7b94345dd9eab9e010
z6d8278d4f51daf06a5b04939def32213229fccf6bc60c003717959a0e9e04b99220d06c1172e8e
z5c0020dafadad7fa43584b2a270200b8b647ba616af83e700e042729d34f817bec21ed0895db3c
z541d3203251411cc64c3fd606de8724b75c9b594f47fb01c251ac888ac5816fa7d5c0eaa61a3c2
zafef7bde5a56863f55b4aa1afe12b4ad74b94064db4c68e211f303eb67b53d4d50305a3911ea0c
z5e73f860ab08a76383ee32815e25fded68049c3d0e3013e8165ca1779c4c624aabe6ec3fc62651
z2598f7e77a16fe4e3b42d2d0292dee34f9611dcae03beda8ee0b4f0a501ae55389bd3369ede14c
z0082c9c6f6ff96bf1171bab520218aeb4bf5c184eadc12cef256d3a798865330b8e14826154149
z6d0593c161fa26bc5b454c279274ceac28db0986ed6653989bdc6d59ccb9b91e9b3a41273bd98b
zc4ed63c702d5b4febf69c13f7b5ff20c192c675f807bd64f054f8a41033d99e91d6dd073aea25f
z9f03422153e45951de8a5e0877db8a196cabdd3392b9c1b544dd36e6fc6b3e5c05eaf3ca52dd68
z313022ed4066ed571b2caf91c9d284ce45519d07cd47f781910425d5828bf81a2fcecdd9f58552
z479419fa8df27da77180ded6a4aa93eacb3e5ad01e95a822435b89325b01b02d8f9a82b2dd7c2a
z650ad92fd539bc66ca90f6af9c1bd98d7222632b6ac309e1bf4f9d75e91a0f02a8f3c415ba2a3b
za6d5174df76a7e80197a52ce6b2e443cf8c65a3737ff99d75a300bd4da3ec52070f0706b23788d
zaf43d99a2b062cf678af98cab1c201227fd8bb15f98c2e5124cf6660efcf833265a2cb81577809
z650a3b13fdfc1c1bfe75234f6ee16fcec37f3f21b577e48068c13988650d6597f2a4e5c1e29a63
z4a8236c9d7f558990c0ab38e6fa7c0801a5d7308a88a084fbe25261b3b38460e2d35e66e3f98b1
zfd48c9f1d61dc9b308376b763b6ef860baa97be3476c5c92eac71d21d69e989d8d7def318efed0
z0b36c1ee92b1e5418ae93cc81896d720dc51539f36a87ccac22c17ffaaec6c2009d4643e93d98f
z0751457f434f2e1894f9e22959d40dee22242776a03466d4a4d730339862af3aec0ddd796da2ac
z8e7950004042c8e7593ba47da959689774a86a20468e7347193276b77d5a70f976f119c34d56cb
zf59b3e2b3c3b3c59530043c9b86e68ee706290496082bcec5f63730f5c000f8659f819683da47f
ze89998072c7e0dfdda26a1137541134d7def9f92b5373691a10b3fe9e1ef42cc5ad760659c0915
zd84f131c5d7031b898c1faeecd2d92e5a953acfc34dad710a6d3d70f7dec55de0d6bfd9b1b9470
z8916899c43dca469c218db82b1adc05df70bb28265fa6a33f835b2a1efc1ce5a52a20d866d5e11
zb5d85c81ef5c761b2fb9f0cf1b8ddea471c118941f49570962c055a2f39e5723a6360707fd0ba0
z974c8a66cca70aa37a0403bf4f473b6196608f3c9ada94b9c18c97c168df02aee5b34094c6edfe
zf10bf5bd540e17c7f3417e0899b126e5db6628d40d20b2d19f5fe76e1283dfc06cb994c9df7d35
zb83235364ce91fb6eba84978cae8d3606e26c1e76dab7aa31fb190f80e3f432e7aa9c33e739a09
z39e3061c7e0b9515b9f4d02d2db315f055825cc8fca31284e593fff6b6b2e5df27e58a7ae623bb
zf9c10e962dfbddfbdb1ccce5e3c9840ee20110ed3ad28aea8f3533f000a909b356a5028c9d5959
ze0d4568c9dcebba3b545cedcd84877f796b4c805d3ce9e6932078d43773ddc290dec0c4eda01b8
z3b9965b025cb553ef0b78a4f401356d9490707dc0f7093094cfdacaa43af1107b1a86545f0ca9f
z014dcf39405f706cf5f408c7cbba920f72d104a830532d8824876d8534bc36994e94736d562e13
za0b69789d17a09bb721a7b793e0d314ccbced93f970a2a0ec39961cab6555cd5d9b99c357243fc
z948d00db77ac9bf502df194db2b30b543adffef03c272c26eaa144715fd118c5438bab9dbf349c
zae60288f49368879c735a4e44cbbf8414fddd4713f7c2cae3e7bf35b73db52ffe0b34fe986b948
z0f2001bf14a6e2d7fde2a0f9c2e2f299195eac419b7deaa951d8ade845d76e77aa19c3f0e5558c
z7d02e3f989a8c506958c1961bb434a2c9ed3c637d60f2473caa761fabaedbc4094747a7d2cac64
z79b5f369222d4be0824d58bfbc5ab1587b038f1493a6690e82fa3bbcaccfb26888eed06c3969c4
zd567f77b2d09e7a03ac0a6d3b8d40dca05072600a2ff77444b4ae1585fe6b24e2333ff70e31284
zdb072f5aa9b6d7ea4f7517f4d92c0ea02ce6f0f58750619a79fc43bf4cf17915c5ca3835ee4b53
ze707be14f2145c168f0d449babbcff68b69e041b7878790243c8ffb5f2bf830c56e919d6230eb1
z27c8af673ee67f883733608bfcdaadcf75f48eeb1998aeb62996bad8bbe902d0e110dfa29200e4
z78ce3b527e7506b3ff160d2d4427c3afbe778a8adb3f761aa92f6a603cd852df14a9601cba7806
z88b836f874c7d7200028318f06ac056337aa4f9b899370dee147b8fbbc2520e16dbcdd43bbbde8
z133f97a6e9dd66b279665c21d19e1d76afa9581e3e0404f8c7929ce95dbd41b97dd34519a75400
z6b243fd405b019d6d6f1298eb34e0aa0e5ba4460e7860feae6ff4bc1c92a5387f6cdcc2f429340
z34376431ea6e5c786d949661665e4b14ee26f318594f5400dd9ee40dea828121f428208b594c39
z66a5f67175b2c990e2ba4adde23f95321e91bf135a8c5a5e55800d25336db2c5ac5f3efbad5a5f
z9fa1e4fd4f0f0329e68840aee08170306e2c5729836697b195979d564f20e9aaabccacdcc4266b
ze3d188289a3b2946d875947131f271d06262f126160628b68ebbbc2ab596a3d7107e28f1c947ef
ze3d4cf927869e22c5f0a5ac9d7fb637d36072f59cd5d2c1d0a1759b23b3d67f5e82b775a21103e
z9aa58aa2af29430108d7788d61f9765670d7790bae0d9854811fd5163be6f9a6270959b1b4d557
z32ef0f0b340c084c2f258a56bec9f496fa677b124e1decb8350d6e8b73a5280acda24ccc66d83d
z8a66aa1d27ed94e30f50385a1e567d33a626d92dda8878498c08ddae7e23a1b439215b6ec14cea
zc9bc5eceb981e059e6b3070f4706184317e5003f58e06345f283603913e1a8639333ce0078f94b
zfffbca2077fd671a19ed125d72800fe37a013d3001db8a63306d587d3e52cb8b2ab92798c75a59
z8dde83d4d41fc41cbf6c6a671006951da3b821d0cdce5b2aa56a4132b4eb9d8c78e1db483d54f7
zd221244c590f07bb173084cbc85462192c35153df29eb60fe83dac20deb0474fce61a39f347034
z1e3006ff71b0a8b15c54f84fbe888a8fbcb6d252a06d1b94c03fc5909d54c9161d9f8c39096d0f
z63f532c420c1fca63dc99fe8564674d304001af939a1e2a8f95663aeadeaae11d852e82489de65
z08d73479b6e7f47f1e3ec022dadfc7d24c41e538f2bcf07b92b234710ab7e6f44a484969704652
z302861940b4066466deea4d7153100bf0970ec64cf2e1672a1cc178d51983a02f91b4302cf52d8
z99b918ff320da6057e836c60694394732485e36b44f748e58562b7bc810bc75d285a39227ac46d
zc4f1a06f7f3b56c08b767c46bf4e80fa54ce81f8a28956522c4a1531e21c37d31739b1cc8d8198
z3d4c332005244eb325dcd8bde90eb6514adf49e0a179440747cd6412ce21c3222a9f3174cfb307
z3240e34fa35988d8a8dccb4c8742df3bf3ebd0e719b0e215d5dd72568717f9a529de29acaa29a4
z5336400f477026a9c4a9559c1e764ee46c841cb9e5991a80250b00daa4699db34bd49c0e2185b9
z905ffc7649ca7d745dcb5cd8d6489079c5ffa24e60379bf77a474471f8b9902b821261c77ad4e8
z5fafa749270cdd5a792b1f2f6a3f3a35a130e36f2f42defc5b5bf09d64f28c59b959edec0f4980
zad8c868efe6eb45d0c5cadea4092e0709788a046a6324f1263010cbd2082e0caee0fda5c927167
z603d44ab868ebd8214a98dc0a140e7b5f8186db67461a4e98fae9abdd8b932334393c1a2a53228
z729ac9800247ddf81e46579c79e14f8718a7fb0ef4810d182486f7fd6ef1b57a2aa075cb14fb6a
zc97267d0a516b2699b2300fbb6dc553c8d3bab3e92866bed2034589e72a22fc02c6b844614787d
z9cd6415c7de50229d46f0c53fac0a6bb743a8e626ecedf4b4ae81d7bc4fe5151db6330d117fc7d
zbbf53a3f8f5540b4680b0eae74bdec487e87c7e2d84ca50b9deae8181f27c843c5d6ad004a68af
zedfd90cab85dfd9d909148892912500990a06ecf408afae47145edbc8aee2f7e1eb8db175aa917
ze774da8be1b4472b89f6d20b13dc65d70d7b5cd2fcab626c9195603d97253379e5a67afa93e9be
z8d888b2895a865d64b7ff53a105ecd2e431bd4380874cb1f1ab0936492df87befb3fc85799adbe
z9fdd4502c24c7b47445260b9c2bc306d32d7c3545575e0ec8864b30c0522dc530b5b6937763689
zc4e8f90c5dc58514ef583d390c75ecb92422ca778c911741fa67c56ac4bdd8aec709422dfb48dc
z4f8644869a380bc328c3f8ca5f9f97ee8e311a37706ff7697d10dab84ec8036016633f843b33f3
zbe3403b2414f022f0c0637e520041a70c850a690d3c72c76308a7c7f36734016d9c8d7628d3fef
zdf6fb0149f97f2020b35a0114f223ea9d9abb4d66807336265cb55ccac482e34ef079d3f6933b8
z7c08722aeef12d8a670761a363a293e766a6609f98dcd1875f79ec5a0618ecf85f65c689f90b7e
z4874aba094ff57af3055614e00a9c61efd5b4385238aeb647517292d0c1605f691f02fcc29487d
z004f4bebbde2885ff0c7f4214c51a5210270efeeb0e0d1d1f39d7385f89463fdc7126329472b0b
za0fc883fe040229592bbb4b0b9a26e4af718ceeb9bf71b7a66eaab6868e7c917c522336a27b62c
zf95f4ea0f92662d09b32b30ab5fbd8368231d866c6bb38250ffd5a71c78ce9ed7f313ab3dc56a4
z9d47692910478afa64b2f87dc3c691d946a6ff759456b096a5edabc78cf25c177124937d771be7
zd6f3245ae987aa618dc6b95c4b6e0f977633ba7defa03fbd035bf31009905238b795be7afdd6c3
z1aab24ccd30434ab8f779b1642c9d1e32ff0c341406bdef06044c5e4ed16b92f6876498ee79629
za882215755f5a907c60adaaa0e2a89e7e7667b68d4d1fceef88100a36aa97d0a39ff2543247b41
z583639f60298cc528790dab9aeb0b87d44d9f5c6ad53394c538d36cf83b7791834e027c32b7b7d
zfdc9e2494e037ba11f52c0a83502e36e47168cc00438796af1fcf661ed7f9654c8b42b2f3e116b
zd10d2ef0685d8e943e572bed22cd6df434159364f3499cbc2ecb46aff6e404b813874e29988145
zc50ac51db27e19e4b9255c7dcd48519b4e98510dd638fbe9d09a152fe0500e911d15073292d557
z968744b844e36c96adc8be8d07a7f4bad778a7528d6769b2bece5011c48511f06e919dffc06db4
zf19d5425cde2306259b2059d8019719d2809847b5127d441cc23c50b37ca2fbc0f5df0b43c9c5d
z0083ab9ce95caf03b243391ecd61f84d52cfab38d349d06f5df0951158132b434fd71abacc4f74
zaa57aac25a1ec30be2a402a0e8be703c2d0127f8ea5fc85234b344d103262d479fbfb5a88f460e
z685dc174ceec704d42c92b6f9b9842044636206b17dd7bda4bc51f6a840c4c887d3bfb467a3acb
z469ec50a9ab96a531ce0016fcfdff8080d091abfada3f55b85df5c700302cb42f260ba3b0e84c9
zfebc61794b41288bfb90c97d82f3cf9a6e2b99fe5a73aebe502ae93534311b1ed0b10c8334d9cf
z5c41458ebf6c8a34965545f0c6ad9d5221aaf73bb5c2df843dd21cbef9413003b083f6e90d5101
z83ce39cd9ebe4cb1be9aa2215d74140634d8cb33287bbe1f19360e3dac411bfb220925f929ea28
z7b4acc95612f6ae75b1f71125b13946628df55bc3a7f042a874f3c2d5d5a631a6a527a45316346
z8319bd76abad840c9b0b08f62f31615256cb795617b0204ada7b01bba02d430ba21368c2368fb0
z91c872652ca93811a82679a7c9328b15d126af8dbe18da28232a2be0ba85d25f097fe01c531aa0
z27f71bb9ec94d50c0011563fc3e8260a397b25619cd37e750c4ee70e3a242cc3b1db3da5eef689
z61bd2fdb5f0f8c8c4fbfdc3fc7aadf222e59b15884fabe0a1b9fd52f91aba3170975476a1a52b8
z53dee01df7b9ca08a03a2578c1e473df4976299d28caf5d43825312a299cd7608fa8f80bc3629a
ze0c21a3e67586026cecf873811aa4df0c1d25d265f3a44e6a697a83066580333933037b3d552a7
ze7eb144f23760be3c3b5302394db94ba0967cc4bd470945bf25430032b56a69349d1da91fa4a0f
zf2c603caa6bb896211827ab6ad3548c4fedf77f4b01dbaf15eeaacd8ebff0da22a0102d64fdccc
zb2d05a76394676e48ceedbbcae5314e3e14fa5815a8544d7cb09270ed8b4001ce422700ff4cd07
zdfffc606ca2d164f112155088c8d58d7cb35b7cb5930cabbb11b4dddb0c053e78341d87b8b5197
zfd9f6fc8bac9c7ef8416bbb0479aa874b4c5d7ff00c97128af254807d5d5072993f8f1a8585bda
z895baedfcbdb1470cda8549c2987b75d860832cfe3ae8666076eb94b771060a52984d45524abf8
zcec1b59c4fbee876511a0166cd3d1063feb2dcf02927356fab49e9d584630e07204cd066ef5ff1
za1695badccbec62e316f935694bae87633aeec593bbd406a12eda720aa621c9ceab5d758c60876
z996ca95f1a89c691e834811d419d77ab57c532f7d424f8f3a8b24c655c3607359c6d842e794f20
zfff01338cc68d26cb3e6cceef0cc4e3112bb781ae1d36fb28a01e45b9fc8bad09908f3e043fac0
z6ff4a98a183775aa096284165ef00467c12ca755191ec28ac0cb8dcb35a4d8133a8e47d3b90ad8
za7431163a6918270082375c7e7b2bc0be7c0a0da675d782b998f7fde015d2411bf718ad64e3587
z5cfa5a1ddbe8ba1bdfa463e1ebbbb7cb45f980111d4c21f80556303aabbff5d1b1526ce7ed7dce
zdb4076006f293e1ce1ec6e83324c57ecda847dc1486916c4a06174dabf1b7518d0ea95c24eb7dc
z58d539a097faca6fee9f8a1e60b6e46b5aa6018ea7043b521b10a146f64bce182263b89ce7c08c
z2fbb8506407e3fac9e22ca9a6bd2adaa5cb771231f2eb9c81a7de342ad7e7638cd35e12069c6fc
z7a950542403d53a9a836327decfc6bbd9259c8f50fd776a986f8df690e73d9db4390e06d2c04e3
zd44a47376f2f2bc58912e010e9ac7b5dcee6f2147fd567f7c9334cfaaea8c32f6368d97c436d76
zb7a34efc0a4d1c7b4ed5acd4f3bb0e62b96f7b59ae544a25b63f79d91bd048b5d975f90fe5e6f5
z3519a5c6c8f29f628f34598bf3c507fae67c8a128b3e0c5d4df42df800f87491fd9eb6f7f00cfc
z5f16d051383aa66962ac0d0916087694815d39e6179c1617fb0a2825a5b5cd3d5cb5c747a90d11
z102ff1617a75fe4d98e94a2e31441c40c284245cd50fcf80bb195089e2652248b92e45de2ee6ee
z2dfb051bd9f347f9523368d2d45c53e942d139c0fc71d69dfbdc937092195d82f3278f65cc77f2
z7ca2ba5d5e7a1424740d602a6f1c2130f85558b76e461abdf4b0611c0f7f94109c57eade4f8f5a
z8cf4377756f8285c80d5c025d6929a531ea2565a03a92727c731b95fd85e06b9720c2c692fa33e
zfe6fe1b076d97215ade186880ee4b35ef69799d1148c22aa4d96e2e913bcf53ddb8c29f7519a05
z0d1767cb4e491d3f72a8d964f6cc126f0a27162df7ef3948753bdbb650d2f81e0dcd166701a0ae
zf90bfd9409cca5839d016ecc977141f44e33e74220bee6a2741b977966f6e9136328285cd72b21
z6f5193b73e49c6ffcc060a741aa74e5f6f8254f16fd4130d5d152b2393cf232b76f799443733d5
z90317c4261c7d2ea3e0bab9738122f4c6e1ecb9c5c4589067497a9693dfa30e26964e7699882a5
z2c53f7e4011ae9a60d2201efd806ebd78c6a902f1d4408673f4f52b8169d4b0ff9c1c55c398126
z5bdccd82fbbd7eed82c8158487c548303754b87f93d2077f3fca1034211858859f3de8d0d6ec59
ze33c8eecaf1efc1bbf0df6e8e16f0a8ee7c7a13481417dbde416146c8bd0f43c4244cbb8d27a5a
ze33ad13a8c1640c806b9fa5c1c23ebeb8f5a8d635e6c0cdcf1b10910a3c73c0e3ffbbdafad9b4a
z32910092d689346af1c24b055a16dfbde08082a4b05aeae7f68e266d7f86e00bc68282280c56c5
ze034b41e406cee15a4a77e9a6b30e32a06ca555fde995801174c9be6c37735cfd18fe57c37319a
zd72018a62ed9cb1ac3f7809472786a695506e6ead65caf107e0c071b26258c82630910b7404200
z4242a337b6bccd042ef2a742650b62c84647fbb3a17f77dc5b6a537d79ef7a6f721b34dca70700
z3ee9016aca4ca3bfd2e1d87b6c0e09acf3878013f127cb95f610411a8ad1edd1469b2af27d873c
z5f419c82248988e6a00aea81d21edeaad99c66a08d918c609b0de0bf6578fdde44bf5d4129e9cd
z368169c21ba18c73ebdd07df9e3e6b73af1f07c4df3678640d04885f280e3aa10faa94fd732084
zb336322105fd293ea13ebcbe7f420cc0ed9f7d7dd654771967fe6df36061bf26ca37c02db9d321
zb8ab10a7d37720083472516a56b4112150cfad95a63bef6073639926367569315667ce1a94a562
za8dfabae595449f389511394f246123d1c7009da33ab8a15032246b7f2442335469b67d90f39ba
z35daeda7e8e01ea63643ee9605c986bf02e7f42877574e213a5eebada19e578b6617bdb425a4e5
z2651a35593173fa353f9176d319a08f7d6c57521a2844f02c4a1ee5a5ade88b4feda095c26d332
zbe7199a02ce2c0db875e56db0ac4131079237151bcdfc139e37891e5839bdcdec9183890225a50
zad85ab49e7694b842c361b2c8daf27c0665c98800761986afd7fd8ebd6e84a636ca6f3373afd49
z5dc013b0dcd39b159327f57a648ba4826f955c4eaba27967a3873424caf5232e1de17dff77886e
zac1f1943e5d20b913870cf0adc95ae3ddb5e9e73b0e45d3116ff5205fcf5a6a5115120e1c8002e
z7b43fb479326d9a4f4af6e31897065ec20be08e52ffd72e06cdcab5a854cd6ef3f428f64d93296
z0c8fcf965da7e47cca4d497bcaef1de143c75a656a10fea6c332a3b13f5cb3c4fe8d7a883d7a36
zcf4256ef6eea502ae8f922f7ae7e5a3780536252c6d019131e7ebb530e8d6aed5b4f6f50214304
z0a42e6f164b5e56120f4b892e8a719f117df7ab7d021a31cfdfe4cd7c08663ace6f1a4d4beef84
z4c80b81b8db433631b2239f610978497e103ef0a2894ecd461dbbdf54df06f23d561dbc6c1f213
za98e69be91d7e41b0fdd2e4298ec75ed2e89385940aa597a6de00f938e89433e92da5696736d74
zb7606f7aecd6403b0c6a0b8e0adf4df3d6981862d0aeace8bfc4a6e1920d23023dc29dffdf1d5e
za7555f46b0223c1ee819ade7603b7d2b8fdfd2100b162b2f55b79927cdf3175e3ea8614b44ce74
zfca52f06ac2d3c8723b49838d1907fc6632cbf9e46e88bd70300881df167e458f91ca9a54972ef
z822f0051fe0bf756e89b7081c119165aaf2a6953bede93c5abba985e9ba98be552210b094bb481
z902af603471addffe3d47558cf260993d95b3acf337fa4e7d67602051011a24775f713bdc7ac3b
zcf5cde55ce6931cc5f149214116d2bfb4d6154a1d3d720771e1826021832023321f1bf6e1d5e66
zc1bb669db99102cd913bd2e265e7575c07eb90a4c528bb11b61bd6d4b2d3c99993c283d2a5a57b
z7cc4f8cf901b0e376daf28f19093933223c6c0b1812b53dc409720235f87824c61c909aaf26fcc
z5783e2d9056ac29400ba814d916ff98a7218931766c5a37e2e3a5a33cc807a81b797a52f0b9476
zc0cb0564f146b2afc77f75f82dd151d3faf13860ffd959912cedf51f6ca8e168194126a786f425
zdc2ad7ee8f570a700c7b19125c798493c7c3751e8fa3736bd08d41eed1734dc6324ccaceeea6ed
z9b5ff2ba762f4fbc7253e873782fafb6e2b974400db6f1eb20441925c9fe3829b7116be45d627f
z99f32267b9f93c994964923cfd5c0f31a1767226838cc1f4e4b78b946a7dee46770f70d6d98ae0
za6529453bbaf621837e260226604bd5efbbfd48b3caeadb6993e71af5aa10b085d98d4d0cd9286
zb51d1a7df87242c04b6926f1bccaf8bf1556057ed31e926ac002970815ebbafd2791a01c91389d
z918176b189064fc14320882058efae51a0558073c57aa04607b0c1dd5f5bdab7089b6a9441682e
z16aee42bffe66fd50a150f7f45105098505916fbccdf899614c2f6af4f88981934624bb43dd89d
zdd94f106a66302e1536168e8950078cfb35d1687c32e56571a0a44c2067c39962a88c8d63a2a2e
z0c0d128855ead39529dfc57ae00601bec67901c88382c015caac0404336a63508cc29b5d3fca05
z1fd3a0e4666bf4e900b0fd241272ab4542cdd6e4c78f2375269636caa3d7a80f330dd49fca312e
zf6192850c7bd9db05579fcd670da11591122377519877758fdb087d51342b289f087e57f9c8a7e
zc8ae8e753c51f5d45cab18c39e74e8593ee6e0743472e95721c10407b111274640da38e36bf01c
z83fd9431f3909f5c2aa86ad939ef505526e42ed500a1e80ff13fc74e9b99f9205544cf0e958e89
zbefcbcda23ea82cd76f03d031472b12d3c05e624738e762c3e66f7128c268ddef86e49b0d7201f
z24bbbbba593c065a5f1b4f2e39ddc1e84981a6139731f456f3c7e3cd845a5a9880cfdc78f45e36
z8f9fdeb5fef3b45c8e31224fc66940fdd0d81bbb4ab052d272e35a66d85b88a08823e0011c1214
z8f3e4004be411f3eda3d2e6747c2fbc221b72cf2b398c75044769fea26ea8d9afb93ee2e042c33
z31050b48ea6ce2cb22cae6fdb04f8f4c39de9519f626384b312c813049c0c93a393957d6e360a8
ze3e725ac6b64d6d0624e987b3b7fa8d201c605b34210acf299e6f26200c67693e22b3c53c7ab4e
z8211273bba3888d8e490df48fafbacbb5b0ee4163f253663289077fc71d6536852c89c39b076dd
z8d60f3d4faae1618ef9a521f07b3761e393d3d41a6f81d78899e1ae1e90042f52b1a069aebef58
z8dd93b8257d5dcecb333c578de82092d51c9b91431799c5f4239601ec9d049c2fd865ef5925c98
z3957f4f7e7e6062593ba217cb851e3df918ec0d63f25c18d76c15bbd4b11c167b49ed41c1111d0
z7efcd676e4a160176725a153bf0c453a9c9ec227ab927de8f53c81ffedc486b35f6a1d7f2f3856
zf5f519bdfb1a623a6b186d33c1112f18995d89c4d5c8820ca832d682bab1de8ea9c02c7cf1f8d0
z274cd5fc530335b4f59b2da9754e78d68c7a37acfffd2bd5ddfad76e351a382538e3f5532ecaf3
z8bad2ea99b683b370763c05506f9375cc82a892d33633bab3edce38ff4a82c6317cea36c45efb8
z99f244a25ba1dc97946a4afd07e73f19cc2ad953f7d34c6e459aa61c3adeb9bc70f1a0d813c542
zb0b06726835ceeb67ebf81af40a969963cb221104de042a9b30c3ccd1118ea92078db124f8d20f
z08f9a074c7d453a74f738bb3c107e0b35c13d3d565b4f0fc7b470cc08c194e3ea6888e38d22c23
zad4a79e32fb7b423f779328f808b0cc626a9fddc1cf662bd449fee0f13fcc0e11f517d501fb1ee
z9c9aa2d7eead77645417a77a921d634d1f293c44f37c523c0c1e19b96e45de65c6eec2377d1025
z01692d15b42baa5627da4e6e6884ebea644e619443c9b23ffd5aa39cdba73d4d0ceb9ce5ee575b
z7106ea9397d05b829b6e176dd7553be71909143fb1b803777368b280f8f0b8f0cb139435b7c814
zcf167c34550ca4d8d0b3ae77aace8d58267114e34e321460f36a29f501d4dec287cca1b3c0089d
zc22fcb14989c474a7e0e43dfbfabedc264ffdbe5d8b913859f07dc8fe81d42eb3222745888ba36
z9946b0a3efc277554a8d4e71c34f03e9eed56a508bdb9472aa67155ea0fe02583c99f0f1c4546f
z460113a3e97be35d5bece1de3f5fbf368bfb8d0a377273618b58394c55c1128a66e75735d7d6d9
z002396ce5ad85814d523d576d8515de75e36eca85eeecddb8745937de70eb527a97076c044a552
za2671dd86fff44ab48d13a908550b805c581f76e284974697d95967eb9903ac2931532673b3383
z8f999375448231a12b8d1061b4b2e82d84867aa6e1bd49317dbb7d658807d0577db2229fe968dd
za08cff9db323cd02511b6fefffc35cc54342abdc6b6f7e33d4d9f039691cec39329ae653a69668
ze2b3a91ae6a378925e24435c3ec1b2cc806f0456696d010d5cabff455397ea2e30a2bfa80bcfa9
za2f3acde567cff4337d07d1987c42cb7ff30fc6d7eb6bdfee8b81eb1e4e77a255039e1412ba774
z1599d0bebe34d4722c8720cdbee970cd6e6c79defd481f27a4434769f42c9036e1f12bfa60c94d
z29b9598f8f8c5a3c6edf2f70e7de9010dcc11f18878560510815f171f55b10bf6e44f8ecfc3fa7
zfd6a7a6fedf6aefaa12069c05ad8fcfbe3c26d8fc0eaf975bc23c9c6b15b8151ab98e2092a9d87
zb8187a5dd558f97e56cffdaaf347af394a2e54c83382abcb9a93362c98bdb23f1f4f459af6911b
z0ce5945e3ff97b197f92b480e91e73d281cc1530f6f0cc5e8d33a9609ebff266eba6456586e7b6
zd8ed5af89796a1822da9e0e04f5ec939fa93a378ce02b1dcee30fc79038253f79dac990d1bc997
z07491aa696c3fadfc178ca9412f26864208263703703f425cccb6c7255feecb5f8aef1bcace9c8
z825f839de703fed56194d6a095428f6ed3a18f09183da7472f08db9ac81b14d377ec19c9d1a5af
z48ac8204c7916e15ac089a4afcf1e3e8dbbb72f85b552f10b020311be61c6aaa5394ad7630ad20
zde6fa03a5f072ad213a04d7cf0645a46086108ac9dd1a71f1d500404d3a22016fdbc353b391cc9
zfd7fa4a4b41b3912cac1cb130cd59f18c1215c381a00160ee8caa9ae45aafab1ac87880cb73085
zb14eca3011a50575e8c93ae343770adedbc2d60c3dc6e31fac22e1e5ee12ecda78edd0a34f030d
zb6c01976155585cc9b105b16220cd1d29e8670cbd33e8e8a940fd91deb878a38ab92347e8b6cca
z116bbfa8681022b88541a818a3fbbb46cdc7cdb8ccf078579a7ef9c782acde9c02f7ff61732401
z2983fceb0858b63359154ed692e62b8c56e424f74624cb284049f1c7f366b908391b690b633fae
zb87828fb63968d4070c500ee582ddb301ffbc3a1d601ad7be0d99207bca51c1020427583d95200
z764bf2056f01510c9c8d09e1d6afa2d73d2014ec0ce036c5679c24f4de7213f2cc53c88316d06e
z4f1fe3b22a1b7cb4209d9903f5ea24be9b4578a9d6c7dc252426269a20370d61d2654053c0c439
z2045fe471ead16dfb894393703b9abe3af0677275fba2995f1620f5937e032af976b14d09d56e3
z3fd27c33fe4bcad842248ff1db2db16ea4b135b9e3f8faf53a00aa6ffa527d20560d135d25c197
z3b8db21d0f6835f4e807d34f172e98a7472bf5b76348aa8d411ce88c8f2eccc5534fa972342a47
z9f25a2076218aa7e86ba2b1f0f231e0fe9105d0d415b15cfd94cd624a28092c82164b3d5a4dce2
za1468eafbb37e2c6d98d6395235781f65b8e5e050535addfc40a29cfd92c151416b2fca9f1214f
zbc76c54d54ec77a32df71a34843dcfaf5339be2fe526603efc7c8f3afdd9cb2fad0fc96fe1783b
z76dbafc5844d0c3934142c01e605c0f3296a5acb87b7e514f9aaf05383bdace5b39b60c9754131
z02123d81001a337d73c396a4ecf1db6162a3a8323b4d1db6993199164df36fc03aca92b563f4bb
z106e2a4b43bf9fdba5d3d3cf301a654c229fc26f1699f3800a9719af690610e7b869d9ee6da7a9
z2da6c4f2f1b4e4bf061acba70b27f339266e05168e8bbadbaed30a3bf479e54d5eaa53413f4901
z6cbf8b986c474ffd4d8ff818e1138a1a6d83e2fdd77b8d5f043a3f1fd25feab2f664379ce4793f
z642d170705daf05886469cc8f896af98ec3509e1559107ef3b4c299aa01c5a572b1c7b771d3758
z8d8818e83b791faa8d2e672e29e255678501594798b52ebfadba3cb7e5dce4081d32c76f415f33
z9986eebc7c54efb76fd8dd594901dfe4f9b2a7a62fc7f4c64335eec5f4b09da4fd8f1d79dcaaf6
z26a0aca8dac2a73b1f23e34f81724b9114e318f3d19d1c154fa1fc662e401310fc2982ad7db367
zaee30870511800a604a8cb4e6b986662906d74c8105683ed29845a42a6dc7e80e22ab6682adbcd
zd4698e630510d371a0a7644361d18aa583846f38ab9caa7463794c1d07982f413cbea0a058f622
zb5a2f8554547d9461bbeefda18afb572d27ab52818d9c03da53028741f4605c964cbeca3e74c71
zcaf0cc2410dbcb35ff9ec5f98457529f9924e30809506442da1804ad4aa6be7f635d44d93c6258
zd7b5a2ba4c60b8ec03a843858eaac167cfaa51fcd31d4935ea145e4d1028b8401f68f3de9f8b7d
z4240b711eca5e3b5265ad10eaccd40347198293bfe0c14bb5b001e74e9d0af6528ecce922c84d8
z93d32ba9c7f8769233e247935347f8800d46e357e9edbae1d8ee79d2d2169d16f11e98ad495e14
ze0e213592afd973ab392a3589f32de0e7600b5835fbeb11b7a91e6270b252d09c96cd55f7229cd
z962dcee6f256caf3902789db17053992e667c1e321e2c1595a7aa39d634d492706ac92441ca6b6
z4274aa9a17d56318745c8d84cd23c25024dcbd80264e31aea2ebad9956cfdd91fabee3a301224a
z3678138c8043f505b96c2f654315e69f0fc25febeeec47284d1280fd41e40b37f0ca5cbc8d9d06
z82a792bdbd4fcf12000b797358397adc557e7065fefdca22780530d5781d917f530ee1aa9f5e28
z2f8e059758bae2f4e82f73f4f5fb6aa7bc61710a34cfddef7a381e4734b8e40ae0fde6506e96ad
z601b318936b4f32904fc67869c68e2157dbef0e28d9c45fbf5d5c4fc726930e53f41e961dff693
z9b2b3817b714d1c93da05c3e721d89a1cccaeda94ae290efaf33bf51c7c25b4046f7b48af00cc2
z26c9c3de3844138a3857373f50bfb831b3ef63bddc8aa28552ca26b2b25137f12e01784f852280
zf47d0fe84f01833636a13a0f787439fbc43fad13428063c7b017509eeebe1f4d62063d71ca36f5
zfc8688d56c381ac9e034058b848bc632d646d30bb4e293ce89f6bcc398a2db3f509d8b7c12f65e
za330807539af3d3d3c838c4cb36c1720c8ad138f106148f8069e340262ce7673c603107cdf1ed7
zc9bed328940a7d2680d2ffc100e0fcb108bf85579a5c358804cab296ad97fdf047c8c449ee4b62
z2ee2fa3497bd6e679d16716b6cee0c427b83b9378dbce6de35f42f26ffa56edbba1e22e4312d99
zb6927c9b7a27a9847e8d910e7ac6652d608db1320f452714a90fb1d0fd9925f8b00aae4da72282
z1021ae8ba10fdd254b7b0fa74b0cf91b092af0551955468c9faa5ee3e56f3c0c8906044151533a
z821f0a9e35e043b7b904fd0479047cb210923deb11d27e691d7f41baffd883650e3635f0e2060c
z08f7fab37a1160618ab3afc58412af3b42a5036c7ec9d70adddf8dc4f0a255287bbb347d67b63c
z10bb23e11ec85507d388e09eb70518189f4d6be5bf179510dbf60367890954f686bdfb31900e52
ze58dc0f3e943963d1e37c4e80d1f133330d9663f56ee78f3be633c630414b7b892cf6ef4b8658d
z2b011b7b19bba8e1941406846cbde457e4c642e65aaa9c9d20fd13871582a09320072b17aee86c
z1b3f33cc8c7caecced895ee477799899b02978a2d70126e912a703ed75271041b1ab59b9cb8b4b
zdf3ce5319f15e216d71089c26846742df40876e190e395c18d4c552088204adfbb1a19ed12bb8b
za3ae9143b232de7d6c92165216b1fcbec1e84c737a16bd01ded3a2217b73037769ec7f602619ee
zb379d34747181ae82c3b6485b2eecb87271a95149cfe90036f1bb6b67b2743b107e8c0aac9d860
z966b393085301b1f3fc001a121e5435187a7fc2128294db49ffcb0cdd32a4c092d404bfe19d646
z14fb75475d7ce85f7fa400976957d2119c5e7f370838b8820ee2e777019de1737034ad732c5344
zfcb6e1fec1ca8a1fef69c0c5abcb3ccbe7a54083a0842b948518ea08f83048462db8f58a59b588
zc2fe7f6360bde26f962f3ae8015d470842627f83e744baa3f13f7ebe15875925f34348bdeb2c90
z43e04bcbb641703bc812c9c65b80faa8e7deec35f905b93b4f8f59d67adfadbb51c03d413a6259
z8e4db2723a8b098df5d7cd4d1a8442d96b1850c8b729c59754b1dcc561bd833cd7465f5a464b2f
z1f73ed2eebdc5cc0acd3472dfaf927cca634dab7de93c0a6d64c8fbffd66c399576e615aa30806
z576a650e9641e0a3f05294fc501f2cf51b1ce6a9b62cbb19d945dd4a37dd8cddc8d2b244ace9a9
zb698d6ada34d5eaf53b549e7027e1699efd61e7bea839f091a008f925d3ab34f66527440225f6b
z7cfd8cd86193e9029441ab5dff96f46851d028e139ae04cce1a1ae58b4e703f4dfb43637e4bdad
z3da2f456def3fa9291144c25b3f97cb1128441cedc5ba338e4cfb2dda07a627644224bae5c867d
zf25c0a7e725ca0f6bbbddff848e2a04078c45d16838e77b6ca8170c3f63dd63f66ca9ce1c662ae
ze7e2a8fe49298451a39fa7df2efc48cdae1fe852a94fd8c768798f8a85f37a601c4e7a261eada2
z27badf84f53026aba11b4138233685deef09a9b5876ed647aa90eccd1788871baa0d2e7082b359
z5bc1f4226677876af199da43bc9fb601b97d73ebe044522f070d489610f75141153135b00a2c83
z607819b3302a68075d552708487a64a16031009d1465c88af7ff5532a30e71a45f8b04dc2713fa
z83f16a1709c5a09082182a5d421d2a80e0502cbf7634985ea569335552483706c53bdc033872ba
z826ecc5b568210183c7821ad8ac44306be8bd51d44809cf368937547fc68805aca4adc3019482a
z2c704bfc5cffb128c82ca74c1307598f307c44d8f6e00d122f843413e8ee4cdc4183f7f5eb7edd
zf4acd8387906a305ab73b4a5c206ae6a9e9b23026e0e5d520e8c7eb9ff0173ca563460a7dcbc78
zd00e96215dc033ddbf85bec52dbcb2eb182abb4dc90a7db163a3f6514a3bad646c5a669b4a43fb
z07bf8a0a686e34096c25b45fce6351bb91a9f01377e8d9a84106222041189c18f2a86d976ca695
z2c43012de7fbec0f18b1a1f12967ff4852fe632dc78277d4de743c9b6bd69d2ea536305d059229
z32bd7c6cb5287d5695f2924b5a31f57f30dcd9dd2d85a73e3093a78e022b74cc03324b01841747
z314fc8dd8893f6069a300ea710a25e3f1e994ef9e02cb0d0eef5e9b9607f284bd95053b7c07963
zc83aca5edea787dd7d4a41efd0ffd6dc83524b4b7200de0280d04ce407a9a4fdaca2df7f4ddb3e
z0fe1529cf18dbe49102dd2ef14b3da21228a2da0d5b02921a42b01e52c3c03f77357c0cbd7e0b9
z2ef8026c61d55c765b1b00eef14451efad4763806a198cc2ff136fd5f77042fc960972545b0996
z623eb6ba5c6620e725c09cfe0ec9caed94261a1ca780682fc159f77e3d841f037dd4c190ec2356
zff4aff3d23d5397672facc8e857e05ea4908a497f1699cd80d7c302b2bc3e27a99b1911cd94b6f
zfe41ea3ca4bb261fe3dba97460502114771105c0b796f9b56eadcb8d7286307949879cdbb60959
z21d6f9cf6f40ad9f0093ccbf81cde9832442804377f14dc6a500ae03fcd7831f1e3d51fe3695d8
z12de41b227200daa15486fc7ee1eec6d6ce09114ad9076c1577ff026befc1d7e68395f22c831a4
zdd2c384121cd319a47d778e3eb76b6a0fc430364fe59481d6c3ffdfeeae361747922b7ea45f296
zff4d3396d094f769ba5542ee6a2fbaced80ba2ff3cb032e72d2187f767cc314dcd42cf4f99a5ff
z370cde7ff3424cab9970b22da315eadb111c146ff946d0ff6119e69c55baa3b333b3d5c8dc93df
z4e7e0d9d90940003e050c0da3c95e9ab340a88d928a8abddaeb5a2d3c7d52aa0367bc12881351d
zb29a5d8171a7df5ca0b53f6d4a1765a27989faad2d576171ec94ec28322e6ed71876302e2b4e9e
zac55b77bbf4e71fa3fabd76e0f015370cfb7af24348388b96cecceb125c3583d4a9f3e0832678c
z78a46c9a5ac8e7a5e50665246a0746320a7f691063b3442c9046722292fc2cdd187e14ed49a91a
z10905a1a3908d50f456060d3e38426720b99755cfadb9ea8619017cec8c152621a0fbe512eeea1
z422da781d352c8b56ffbd2c11b27d002aa52427b91eaeb95dca95e3084224152b4d8e7abfcf422
z67a7fb99c50f25e95cdc50fbad805d76f6726f5dd4fbf684c6d9b1911dcc1976de73b993ee4ba8
z75e9bd376afe014ff6ad883b39cc43297bf7c90409dfb4e92f93c0bf3e98c8d02f1f52749f1601
z735f18461129a2ffb3809d3a3d9905c2e3d3d5182eff5b7c35aaf95a5e1a4e432728cbe9e6a072
za1811c175259bc0a8dd0193ceb145539b5a8c850c7281c3861bc6678477a2804148c64d0e30f2b
z5284b0a2337661d763836a74f789b86cc5d2e096ba43c266dff2b5e769766a1a2d3003df08545d
z15fbcf7c92cae3e2dd7fb1bd91d7a076da2a5080fad5ec4d68b0a2c8314f17e5f4ceaa5af18327
zc52356341d947dab9405adc7423389c7df5403935aa3e4e1767bb05567b2fbc598e023d8bff54a
z92a5d64fe606a499db212213b4dbc3d567e67493c0e8fd4e3ea44f29fb8bfb5e85058868637229
zea354a624f4c50d1f7af044e25962d69e21caee86dc7823d1e48e7cc124bbe8abf56548047cb38
z58741e786854fe735b345cadbe94ca69dcedc0ca33d21d9aabe5903833d4018c0dc58e7e678f8f
zb73ac33499f3a7251309b6481cf70a5e22ccc9e52ff7fb93b4b87cd9afc782f3230018c7d811ce
z75522e91156cb600be3a048a384dc2d55ab1fd412aaffb476a2be8684f197cfb9394009e7f15cd
z7f519553ce0dcb12b953d69137cd865a02abba114b32c3f4ebf5f9db9de7e7701ae6cdf7bb6d51
z23a32e6fa3f23443c29d6fc087688d4cd95fa292e7572ee44710fb7fb5fc1eb376f38aea8c7b4e
zd6d13dc6a431f888ba0e96586c5dfb97f4968314e0fbf19f55c1f245597d710df1deae3b9c9a1f
z8d1c97ab190828429cb1a60d3a486e1004826bccc90f97edd670511d786f21a2423ed4c3b078c7
z9a5465bf8e9f13119c90148523c809088ed7ceb146d6c374ba208d60e55a442e634c83269262c2
z294817dac2d2989c364fb1d6a668f3a066e5c5f0c686b33a14675391d1a42e08552b5d6ab34e62
zcdd5407afe3f48df96b56be4e49c07c374bdfe464a23db7e2056d9672114a441ffc000f2091729
zfc94be014df803775dbf1de316b01cbe5dda8e25336656ecb08ebd4745e588005046ace978698f
zc7ed82f9f7f8aefaefbe5e5a0bac6d4d398c9986379b39e1fcc0c68eda2312e614318f6f953e39
zbb68c088b6ce8c4906a57ffdacb560d4779755e7ddd9e7ee2c0be6f25210887555ea8b6be2a7e1
z1985308969ca4b0476779df23ff10f071a942bc9d3e3ff7c161ce28782eefdd6bcff535b2c720a
zc1128967102bd4407b7bc7804762267b6280ae28a98a1836462567a5bb18e5b9a6fbf78660ddbf
z3b4c0d6e54c5c0d32ce524cb269fff00cf6673c26c4992ebf21f1f831294f741ecd615778b3f05
zd7056f726f4e301f1b78603fbf77f38f78f43d87a08bf15f2cc1b3af236e59390398474cf7de10
zb101a47973b303f8c82c4eb3a2fff16347d50cdbfeb2c30171dd31924c91f4495df01f1e016230
zd6c2c960c59c39a262188f4aa9b72e9634782ec5d77675f0e3f8fefc553e1ac86ecf32b2eb4178
ze9a05a6ae2ac3e9eb172a7f90cec0e739b5d309ca90bd1a02865f3190f45a3eb5aedb99fe3b517
z7fcf8a080a2cf95da0377d5dec73a240682d35ae3117ff4e5cb420b3adaf56a0184e47310ac6eb
zfb16b2a1a2deb9f874c19dfcbb71fafbcb05ab41b6c882ab32056875281ca42093488db16066ff
zcf7fb185cbd0f2c67794556630e0d5b4df0ab43a7b1ee4b4c10a896e894a7dd660f3536486b9f4
za885b2e9f03351e7f1e7689eda4ac3886484b6ba2aa1126d1a2b1657e14685f252343bf499fbad
z2945cfdb72740475edf3c986b8ed28141787e3b0bac61d3a4c480a39168a84223a429dcdb8c64a
z3900d7fc573c82843ab2b5de65a6bbf333b10e800a905ee8955aeae73b775f021ffe505c1dca18
z1a2e3d7c85d8197e9fc12322e5d0acf00f969d87c8fd19fdb4085d85df28e4db9425460666e7c3
za9a9d49136aa3fb087a6ffbf9bbfb8a30375ed975981131f77f3a575b0253a65b55fc3b739d3df
ze2598f22abd28aa1c287c5220a5e170ec3726ab791d96a497bb16ebe063ebfa08fbb2ca2ea82bc
z7f293b36ed84115e346602d7c42e9a55357e8752ac4fed2101bea4d80f78f7df430ad5f70ebe41
zae26e11899c5e91acaf35052d2c5a4bac2b94c8130a89f6c75c6a347a11edabb263ad86fa58b07
z65b45fe9b4c71e188d11465f12783ad27bbd4fac354cc74397ca1f8024504ed7a0c3788479bb9c
z7560aa2700e4a2105b71ab626eefeee09470d014e7e21a49965ea38487d5546620aa70ec8d9c75
z69ce3f5c6c1c17cfa57b878a4a1e67e03cdbb5f26d28e4e6f41d230a65cc001136925713ca3efb
z88ae2f8c1d9af6cba5bf63f1135caa344f1f522a76a828b7ad9862dd85cad1173d12f45a200e72
zf3e6cee0811d3506151265a2133b966a1e050c5b0ab6a0301249f2be21df893b8e01fa97c73968
za974210e55d087246e8d7b2969870127fa221c57d0722107b4a103e0921d2cae9b8c42e35ce47c
z6b3bf556b4831d7a73a37c025260ff056412114db76bd1324a8205f45f70f3ba1ce1f6ccbee511
ze92e3f9f36fb616dc0e7e5ae33d3e225bc36698c2401f604b1121a607a4845b270d7673e450568
ze7c3d0a22746fa3cc78fd8804180d4f53035ca2b3e6cfdc098d1869f45feed2231d0540694e93c
za95c0711fbeccd711c78f55945df0ce79ff416d0af40f6afe235a2e2efc82030649b09c51599b7
z8b196dca9332fa202bf556ffcc17e703637d5d56ed4e9b20af1e697b84b5424aa30af5cd30b27d
z095bce09d5bc0d061bf30b6e73f2fc51ac91c2a258b5a628e51d07684418bf8ffde02b2791e6f2
z8371f44b36e5924357c8ac9e2337373e31d24c3feaf4338e73a8c061fee030776be3cbf2d0889f
zc1e4a81eb998e413af1f82eb84a2b5977981e4c29a194c30b7d26c5fa5677ea4b9c8024ce7ad19
zfd4e76c9296dccb4dff55456989426d55522762be664712704090156a35cf54e7ae611bc5f1205
z1fcd67af87a8b6fc51305834e963309010be626092dec86d67889f610e460bb22899206e920232
zf31c6a0fa6f02b237fddf762bc6b6f1f8339bf412719445ac0084311d0f2386f02ab86111a31c3
z7ed263d2b92c5494d71dc87af8d6cce920281df292478030a687a6c56edaca948776cdad3d9880
z151a6f1eca8939ae21702e30142baeefcb9a08638f24e13e352875197373a06d83ff7fe6d589ca
zae51683c1e9dd572ffd155fa14e74cda2a1865b0e897cef6d64f798203d5aa7d1d4fde231b29f3
z60211fd5849f440ac14f4b3d5c92559ff753c35c284f5bc1f6f1927adc24373112289c00ce4825
z0f802dba3f2e7666f49d8da3d53df77f4eda977aac278f5f03b9548f55493694c958ae549d5524
z092addf785ee72a4cc1e5b5ef107a96c91987de7a5a9362d5f7ab07721e32adabfecfee1db9c1c
zd9e54e1973a7d67fbe3a7ae015742a282f94a779bc5c3a95867770a58a4310065d72063a933171
zbe8e7c904a7e65cc1e187fc6346074e779d36254ac881dcbe8e3ca0aa76361e8f8c17f41d37ac2
z716af04e056a5c598e9cdf939c498bb19b8cc6042d377a774db3827e9256d637ae101fb29d5d14
z8763e55b3ae79135f94aba4809d9807377d5d0cb4e017cebc8f48d9c33a279ed2a9fc1aef01037
z89272f15767b4b452d8b401bcd3dbb97c83844d8906d91efa7d9391a6a5b7ebf13cefc40fba640
z4fafee05d40531361cc7eb04df4f5b3e413a7c25bfc12c67ae2e13855bd9faec13e6d9b45580e9
z38fc62de769e65e95312f80a03f3a7cef221e5f2140211243e06166ed9dde73e578c1888d00199
zdb618f8272c29c15f78dfe7f7da420f59e90ea535537951a44f3cf820b467c94a30856fc4d7faf
zfeff49cc184fb163b3b0e83d28d02bf35469cecfc9d11a9031ba22f6f883fa478b70f26c26de32
zd06ad6d8004852ccc6ac7bb435ef5a8dc645ed2a7c3648ff3bec7ce6b6d2a28cdb860727225c8f
z4758d09d54d6f48a0b12dda9c6f0d88acd54b9a2627a6bd5b05383e24f577d815752b16ba1fbc3
z16d9ab2afc8d680c6f2a06a7ba5d811bd8aafb4fcf2b769fc3bcfed1cdc956082d22be66b9c5b6
z9841677d8880ddfa6d8a6efe538f2087b5d53da5b389f0e8791b996b71f91a27f06ee4fae5c97d
z03d9a4b6a9b6c862e30263dc9e63363033df917f768dbc8712f881c1a8a7b503c388d0ec93d498
z9884e4a2ca3d367f07facba69bf5124f9a5ba558806837fafef888692e6cffc3a32e14a93e73ae
zf2e0414ce2b89e4b6a7e197a0f845ddd67e5ba53362d952ef698556eab9048123c2baaf540fba0
zb0bdd501fe95179bf64570210351465e9f943405e378ccb64d570b20d56d4f56442b13174d39ab
z3cc5fedeb73d882a53954dbec7ba01d9bc7a4ea0e8d47f7c10fbc1deb469fc9cf90fc5cb751359
z5de746e20c417f258b53a0e6d491dc139ac4fce0fcfa53473a638e80881d7227cb5de07da81dc7
zbc5dd6de7f39575738b12ecbf59d53d2983a7233bf3bb17b3eb72ac5bafce7298cdd73afb4af73
z50123c11f719c218ea4dfa976be3df91602bc9278c345f5c8d77e2d7d8ca834a0f940cf79cf15f
z358dddeb444b3f4daab41c046d5a3261ce97ce043d5aa8e93ca2a7c9f3e7ce3a8c41ca03f870a7
ze1db440bf047dccc1ab49aa5b329c159e3cd2f5e9a0eaad2949b688ee1c23bc512e2f72380f71f
zae4b7f87caa0a6c8aeb8d9ae4b5bb72e30409303de7ab8902bda2490c7e14c3cd061e476b6b070
z87dc9e283863349d92a387c6c1bf2c6fb5a7e87bcf3f14e04d68032b3708ba4569c4af32989f59
zc9c9049410e25762275804711cd2b819edf067b28ee8e207b5c7ec83896d3f71ff3e90227522c6
z2259f917c74a56dca72f103eed3cb2de1677e2d3f99f7a8c1c4378f65b687de26ffa51ce986789
z2d1155252974bed438df860cd923e67ee97b21dd504762d576ca65c1e2f43a43ee90e178935bdd
z6dbe48d6e8c72101c103e693a66cea62be8dedb276db0c3ad48c5825ae8117536143ece59b1bee
za43e879da63ab1db0a6846bd243796fdd506fb32aa1e946e340f6b367b28e434453caf14b2b7b0
zaee45a7a32d48e4438f765d984e3af8c5c00a61b5e4f58846f896c4e6004866b8268f973a020cd
zda0337696bbc2579c3d9ae3116a473dbf004da33fa13da1f084cc3bffbec61c6912e9fe10ce8ea
ze0a6575c96558c87b728946ce1a2f69cbb5b81904fdcfa9b8b92d74b0abd2d04d60c8f8cb7b825
z51bf72e395d2ea39b980d5614364e264aae5c87e02ba67ba0999530fabcd3a34b674ee32e7a749
zd7cafc40c2ca54451f9c2ca49c3ded0c20b5f34fce8efb5817b15e3b1c4a16e2ff5e5af94147ef
z965ed1c1b08fb0b35f40f2c901d5b9fa03819725a14c883cd446d808dd117d81428c06070988ab
zd1051156810b84a58fa41da80ef93aeba0ed76afccce3b47988c19c88d3bb118bf1179b29273db
zcd93a233b8d3f5493cade5cb1c99bb974b79f8305680b559443897bfee364b26f2e008228fe124
zc0a6604a939d6192efdca30777fd8345421b8e96f9df932359695d4222057cd1f060bf1ef4a3da
zc25fcb821c07c0d9ef333ce7c94dd653528ddc7c897b01a5c8920712ee4d546ffd4fd8d55fa807
z42c081d582f82d605dc9c6414db5c610790c5bbfcec78f735b7bed270a54d7e246a9e52ddf7d0f
z91c191bf57b6e7760083a21cb02b063733b525c35e0d8720db29ffadb61c1026415189db2bce63
z84581a7db86d926de031e2b1db575fab3b4090a5782776fe7c0cdbb56fec96e60b98b5ab0c5d05
z948e678a25fad20557ca13234b406fe0935704c533db0f3a6ecda43cef43df5e41f33457deb6e6
z0da66f004182f46e84be97e39d9149b08a1cb7044352b7bdaf7e2873d20c5ff49fd4640f4783a9
za70e4406325e7e5cba23a59f9e9887666ac75517622e8ef7c24fa6af6c7ee7526fbd8694895bc9
z438bfd429f3bb7f7a73ce9ee3d158deba227b583fbad6c802e660399882ec3e5610d871871ee8c
z1bc4d52f7b504353216b8857381f37bc501d101ff7b5e60eabf46a0340f61e07472dbf4a62c11f
zfd70dc4d9521bcab82a8ba42dd55ec9ce2ef1176fa162d0bec9323435f7ba2b70ea7c460ae3e21
z232aeef5e8a447b48ddee9caed7d97e857b4fcd9365b81a6051fd9bcfb0091f7e915d71766c986
za9aff16b91dc9abae408c31626c4f95fbded11ae489e14c7daf838e6d42bb638014f220cf5f473
z151b73f0b77da2c64b5c848ee4233bccdf69b4a84f842cf8c54972409db503e2c0ac8ee1d8da46
z991eaf6deaee4beead7fb0b9e2b0ed490452d702f728afcb905414be73cbe10fb30d9f593b3eeb
z750bd90c87baf5e87d04cb5c55e218f2854d19a5d2c04052aea4e66874daf3dc44f99d9a6c5fa9
z9599b0fe3ae4533f7568c830875256b8a3476e70dc4f48a2e66b99845ebb9eb996880429d35d68
z373f38da69bffdd9dff049d5f1343f42885c704d957da086db6e07aedd73d023815cfc2b79281a
zcb8cdbba5f2ef64a0051474e57881101c576a56083587ac4b5dce2fae811b8ff30018f60e83c57
z7beb02ce829221cc35d3b21b8687bdb4279a3d72d195eecc3e0618b7cfe3fcfb2732ebf34823c6
z9ce76526204d7162fda352c15c1b7400d74263f1741524e23b48a01017bf6d7b617a6f01e4b13c
z96358dd6d22c461ab0b4823213b71f1bcdd8cd69ebc4cfd6e11e3422c7403e8f723ab57701f9eb
zeb6f2d57d435ec3b36d78de9a0a8f8fafa582620e0668e4b21bb391598a7048625baab50bb7196
z3636ca99786f9d3923b7b17b631545f3f2e46cf1f352c4aa74ca01af945232548c8f620a9a059f
z34108781500386bc585337b2b35a83d3b922275ab5dd32ef095b7cf4f61665a58048d32c4f487a
z51d047eb632637f0e05060a4e8c0878f99ad45a6fae0fde08dd3f068d86cc97ca08ca48924ad3a
ze4e1838098fa187df56e4d7668f6b3bd9a022cbb6d6c515595821f56e673414cc244cf6bb840dd
z05f7293206423cb3d1490419b97f2e7d98e26a8ab5f04a42d68ff2f066774838257efc28a84383
z78b750477840b4ac4d9d495350fbb42d9881d9bbec87ea9cfb515c62121853529273b3bc817a96
zf5593aa408db03f1b27b6c6c7501b0fb9e26ccea520cefa098524b6d3934f85a010fbc189b9a32
ze6a6e231a615ec8360d60e22070c5ccafe2a697d6b7b6aeb8154b6dab885205f290c5b0df61bbc
z3276c72aad6de89e4b942a3f3e6b6585e150d303aaddb38b9b90401891e9c4fc6add662aa7c220
ze471203e5414f7b8b775330f44a5b9e5bf28f636776225e1de57e42dc4488e1ba11b8ba4b3ef2e
zb4c8be1a7708617572a0224c1793946b160fbc3e273e4b6fa097d78e7af1e2fbbb0bdf64484ecb
zbb07813487bff0a37946884936485f16216304497f446c166451f05f331aecbe78304dad82e220
ze4791a63994235d9401b6d58d2efead29c1547b09368e6619a0bf72774cc4857d26a40409a96dc
ze7bbb3a1957added0c6ffea6cc24b035e0fb3f053faee6341beec879cbc0164a2a9c2df6a80f4c
z1194372e0479cd1ab71ad0db06e6241f92b79f2eda13509c821a23a76221c04d00a5f3f5f0aa7e
z0d80912a43680a04c57f63ce8f1f658f69a08fd1d6b09ceecf1dd7e0862aaeae867b6f22e379ca
z776515fdc8693f5fe21c4673275980d3bf0540458b06d46ae062fe19cfb1ed4a71c69f9a98a58b
z409ea4f819eee133debf3aca1caf55b09f547bcc7d04e9d188446ce076ef93cce2487afdad7a5d
z60b0ec65425f8a53197ca7848d753d3240fed3b615c32dd29ae4687942c90c9e8025ba2ddcfafe
z772c410fd682adf96ef95c3e820804d8b8a21623006be32b5d889111978fdcfd76a218fdd5de85
z11fb338b9414f3b6c06f93ad2a0deebfe4243c317dd84db4b86df2138a69372655ddfad8b5ebcc
z066dace3e1134459e8b8560e909596101d3927e54056d2a0643751cf9a5ce8048aeaf9d89b22b1
zd003f0fb2ea288ba5839349770acf5583c3056827ae992a2e5e1cbab37878d8296431def30f49b
zeb1b1436df8a7100cf401546da9b78d9db35844c5ed33f39a4090254ca388a52c6a2a0e33aa2e7
z02f00fad93150f3fa55f7344dac173b014149c050d3b42a6906a9ae8c427a98eef437943fe730b
z7e62dbf1db1c0fa5796477b67d516e071bdc99db5af8486ef8603dea7e18fc243a8638a697d9af
z96a6b5b9d4759c75f6c55d3d58ba2575ad0686598e93b691b409f03faaf60f617d8b0adaea1aba
z4e612aa87676e85c686a15538a521b2b7dc87c0010d557104442ab4d5bd82f3961b64ee64a5c69
z06b28ba2ef9392efac05d07e5ac1158ae3bfc14864a9d2f1516c55301bc7e03af7c09f5549ed1b
zdfdf801e91430378c924352f85c7b57e2cf0b836942a9399e9dedc447ff2e8f2b7c035908b6e02
zf094dd6fb8b48ff13a6c359ae1e72c838c4fbe54ba966675e4a97d33cec2c43021bd2888fb42f1
z94c95d3282223e2cc2131fd3633b5740759c55e89395746f8028de5d8ca5c03763066881613d9c
zffb9241b7f82eb200d90b3ed8a872d7ac3f60c276495d8cdbdaf9ce35d5f596077baafbd3e4722
z2b69ae9596651e3e62fe9b2d6ebddef0aa894f1f231cd6cc63d6a10835218b919eaebb19f6f45b
z00669a44abe09770d1e403bdcae900507e8210da228022ac44cbe1a4d20a9144000ab977c1a930
zc14a20f083a8ec330efa3c627d765e3fe2de4bb907835d2eeba846973d16e07153643f2012adbe
z3f771146f38d76cd6cdd8df9e071d47097f4d1166ac3711f75c242c95ac3ac93fbc66cf91759ed
z5dd5e5dd2d5e0c82f5cfcd83c253183d175732bba0e57f1f07087943ba503073415fe1ab75ff5b
z57ec57890b9609e5015ba682651aa92c497abe4b4e5bdeea3d90b4b00fa3b50cc2e532650243d2
z3b090cbfb980fbd4cd696c62c717fbe2d872633a49c4d7e1c4c2063186597becffd702d2ea5952
z0ed4ddff0e3832e87ef0dfa0b2c0d654c10c9c8df9b949925a2b6792c0ea7f85213e996e5a6871
zcc8294cbde94b0b8a2c4678f3e872761fbde3be3251b7c9efed87221f96f84fdd9685c81a4ea76
z837c24aaa618ae1030c45a7ab365ef03abad0ae770c9b008f0d21b87bdb135c054468726113458
ze6f8f3b2ffc3b7f6f23903e4941a5b23236ef277afe69972ff222136f36839a4a1e76b55e52fb7
zcb82ec9c9c0ae2a2a9d59363aea18e13b42444b08f9e6e43072a5ad6e03f878f9210362afc5541
z542f6a856a70fef8816d505e05cc5d86dd69c3dfc4b3e4202127d1cfb73e1b408f48064a7b2bb8
z8374b1fc45a79c727252a8df22120e7a4a7325f50c5b713da14a902900ec687a285a77bd84f0f3
z1c08e30e8a0c3d983caab9bc5517edd7b89921e5c9fd31e710ade637463d01720f5ff54a7e6452
z775c32980a1202276972289e8de9957360c7b03990c91bdbc99363e55b86b721eea94a8b7c32b6
z3969836728661321c471d412e4f11c3f2dcf6f70f50ccd18c1d288ca4a300dc2fdefcb8318c325
z5a2620303b3c3be1b2e5968938d0fa338e4a039c2b54acf7f36763da5ca59494c3b437ea2afe46
z7004960adacbd316116eaf952498b8c3c43cfa90bf4961dce048ccc30aeb98a926c556a6b1dca8
z50aa76b61500622afc81459eed9d178f088f40710628c0ceaa6e622e13e24a7ef64b14f920cc76
zbb5a88871460dfe31b2564f19d8885fe378415b6cc74a2ab06bd902f4e0118b6b4346097e145d6
zad39e8d73cd4468fcebb835aed82d8a8313771b26c25655ae480df6e3de5e18c795a59b4779c80
zc393847f0a864273a532415928b37f05af1bf6fcf4fe467deb982a66514e1e5bfcb7d45489573a
z758c5474d0406bdf2931c6e85738651bc9834b75ddd14880b884fb0b344d346f7d5378036d16d2
z0629b39bc171f05465742a220891a5d278aebc092b527f862c3debf106af18b35a02382b2c647f
z58043448e2f18e069943edb199d878f790e91240d9cc159086016fa44afc57d3764c153cdaf29d
z2a868d24ed53602d726d52193f6c71b127f62fced6bef5a68d7d2c80f85364b43984adbab3f628
z7f4ca7cfb5834aa84b746a95984e10352d09ae71c78b1f3f1b548e49cb4e1165882b9f83845c60
z90d8700c11bd7d17a57b9fdced050db33b2254d40edd2bfd2cd536e1f06ce5a9086ca9541d9293
zb15b47ec4c9e69f665755aa9542ad72b805b601d78e4ff5dceb229c29f3ce5b271eb495a908c40
zd858322f3a4aa1f22b500e17c5f647c918b639fe418819f7009a898f20fecaacbc5ceed9326ae0
z43bb67a2b70b3497e8cf739c7593d15c75c57e548676aa5ad955a234d87229abb53ca8a779de91
zb0e4d50b0bfd02a9d983f8b177198c34ac3c2a57ea9712e00a4534b2a937bbc13a5461c5817c26
zdcde6e11b11041650be95723a2fd1b81f55538b883c2f74a22fb7627099e2b784c70aac59ed9c3
z62531d406a11e8a71a20a9e50db45b4375c07ffbe7d8b0ebcac043df2cb110530b3a7a96ee9cfb
zcd3f103067fe999a2498b43250b1aaf48297c5e8c18f81b651e440ea1952b4b39d3b2f73035c46
z8fffdd72b0abbb85c6480033451e2f6ebc1505d0311c0b256c99d88c90503eeb888a659b937ec0
z634a369d9d6d508f14550b898f240b106fa23f89bc7f71f5a1815bfcb760510ce4612070cd2887
z5d06022573ce3806a96bbfc7583c7f87a322d0a592d655b7724b0c83890b13d73637941b6a37c2
z088ee7d189e78725fa7b4150b5af262296eeba509f2304f320ccac4e7b33153b7d6a5a06e4285f
zb1cb18e32cc167e4568f0853f8f0cb1a255258f9640c9be4da198ee9f3b155428bc55790126ca9
z4b3e52ea2fe793284f18fd9a60bf0c75c9e7b5db019091bdefb7e9148398f486c6732fb481ec7a
ze5a6c1e99b191fac7bc5b8178a4edbd0ff8ee681a9918a01545e920af61703ab086ce6cb30eb41
z9c0ce4e720c53fb1d81159d37cc75a0be6d1837b13edfe5c5c22427e20e0f7fe8c6855385243b5
z50f25f2ad100af153d94fff017fed0110bf4f72eecc6b52a5c5ee2975d87d44e3af21b4a2685ca
z801584e6a7663683c34a941df2b1bdd3d2414e64d8d63dab9f7443d998a6c966a7d5b8c913da1a
z73f0b3f32c7d040f4791f60b1f32f20732f4417ef3874ed8c376685f1b3dc254ccd8b73b8450c5
zaa14d14a4cfe024cc83198bcd79ca194ad625b594f6c81808bd642ab570a730db7720f346165b5
z8b00d05792224484734742f7436822ac38b1b40772e75a6f5b0429e537be43b2e53f1bc696565a
z9277f0d8b0090087b869ff1ce241da7e2b7f92d69c3c74eff58c27ac79847bf3ecaba8d44d2cb0
za83b6f1edce5019d03336a1604eccfff1cf0effe3dee72ff674496ccf756628936fb80ed02b577
z3014d0bcfda4baa5500fce08009e7bfc4cb371c5762b0fe91b57aa017ee8436b5eff2896721923
zf74ef577452d4e3d2ba048c51f3d758ce011848c33046bc3f9f47bc49927d2b64758063093d7a2
zd0c835ec51f1595e5f8293a8c4caf7749f4030aec9eb2bbb4f9ed7a34cdf3d8986051a63dd046b
ze68ac5ca71d8ebe44c8dfe1c35692e27239a0a9ca26213d4688b0545fcbca9be53e1ed859ff9ff
z43cdee42826983f6bfbb1f0cb4727e8e53c5717bbeb66c186ff0d7e06099c242a082985444a0d9
za04349add3ebf108463d9245c8f0bd637e583d2e39f2eb7f317f60fd869a3f793af6167f5fece2
z7d2ca0ab362399dc9738f7087a014607cb1f10d9ce57b77f940405cd321b34da0fcff68081b083
z6577850c21fc8918e29cae34b0f2c5744504ddf1040750ad7a790a33918a63731ca2fe7d173456
z40f01682f25c0006e1415548d62090187a6eda6a182cee55261b2359e60d1b801b4e1772a48885
z3d77dc34ccbd55ea587125f60ac937921b1ac6d2effd774f2b81e7a82c64dddfba4033774af8fc
z8c0d2ae6133720acb0f614a0dcd19c37aeac0c6e545e12cb84b36e4f6266a8782124d4a9b14446
z3261bc428749fe0c4360f66d0e6f3d84e9e0077406107e80a88cbace3c0f575dca563811b4c1ef
zae9564387c097030054132d1e7b21682e95abc89da40d890f686b4ed9b87aa367472b83e1d16c1
zfc2d7244b02e46cc28890157a3ecf671131dd80fbe047b5809486976a70a85f3f031f929ab5613
z95a7974bb1d66743a4d1631642e16cf4b7861b4e10d25573728a0f794fb9a050190876a120f571
ze7c37fe843a97cfeec5ffe9ae93f3abc619330c3731c2a8196f6a73974ca8cbecfca9601ce8a19
za48a18e7d337321fbad9b8deb94848c208cb6976d40fab62312f6f36675bdf19a6cafa9cd87972
zca630e26619e35f97d22eb67a2e145a2e245b79841f0e4fd00ff86e4ef1d28fbe81743d4e0c26c
ze58d292a715069f2fc4cf432dc44c746d08d605e349b311e9a1091948271a33951a2f74f8573e2
zee997a13c9ec290f3bd6ffdfbf155d77633d56e588118cd04e1b935a4e3f832f6766b8983006d6
zef1cfb5b091fb23ccf120584f347d666e04a276979fed80e87a0be3da0c89b6099e76cc8c383ae
zc983e6e66401fe8729e55226dce54712abce61fefda1c954304e82717574aef3f73c0c06239607
z3505c918b8bbcc6d08f13da5987b1b494102b936674ac2d6c4b651fec28ea07fa9a08a4734060f
z7fb80d66e58c7d6cf75fcadc6b1d9e3c6d561d35b315a39fdb138c8b3b2787f4c0a8838cf0063a
z7b970345c65fb39979ab174b9b007aae695479c211f902d6a08a58e471867a2bb5eade4ceb299a
z6812b92d3f86ffb407d4251f19cf4aaaacbc621394f448bebcb27484050ebea839b2519673d320
zc049f088b47f861f09fe2b63fa3bdc477770eaa2500072682ae39605756c480e7cb78ccecab632
z118a4ba0b9a851257eb8ba9fb67b0b38c1b9b5b686c59565e42b611b21c895ca41f59aff78d96e
ze437b5cccb20be81cbca09bad0c3fd01c9f15f1aa3ab613fce8d569ae0e32f0c6d262b769963d2
z7861ab4630168d228c3566adcfd265d7bf94e401fdf415165689b0687c83f139e362fa76eda81b
zd27d545c4678b71afabd53032c7d9c2c6cee30f7c5eb25303deca4a127029a84e897392bae9ff8
z2668884773f07dc6179050ec1afeec3cb81530881dda4c486318c1f59bf04b77682d31b36b55b8
zcf9830194d27c05877318d8da8d0dccdf46d29b16bdce460c661508ae9a32e5b4b990935ecce19
z63fe1318667b60c072222a86836381dc7d02a94a73c86ad7515e59378e6a7f35e91cc52d214db1
za4a06faccc74c01c86ce0674af632a670ba55987fc4a517668fd4a2e7c4d453584cb824f16b496
zd3fbd48b97c990e59bcafbcb2f1078be9456e35d45909f6997a59301a144610d55e60769e932e3
ze38ee07e3b730453e8be721bc837d0c261e5b757d4c2fe424c9e344e6c76d92c9ecbeef796872a
z616fb2c519cdf7e877e6c76c812c51b3a6dc0d04917d63f484e540b9dbf536af3ac5aa2afe482f
z4a113456bdf0bc52a1ad5c901c3fa4b3cfd264fb5ac1413369d98a803c9d578868643208a20fa8
z1bc9a840d17c7da5353d25ec4acc6c13b4dc2c28af918c98cb6bd22a8c852a304569381f819fcf
za3b520e193ed1c91d1c900826ded8127aae5958be020481dbd9abf1bb461b98119e9f816615624
zfdd5314588e867b510f53ceb7e4ae6206b1518add972dee70e96c437f452f4d3bb4524a40ff2f4
z8a5bb8ac7b767fe715f7caf42058d56576f96a86d90b6fd2c9175351d5b5442f26890c17422b21
z3efb756d78a34ae33aa1c3f7a9af50dd173c9fe05efdf5c4af08c2d92bf8ba2d9e9486081a986e
z646909f0c7b7574eb47c8aef49c1ef72ac7f747b22ddf9bb5e327db0b2a66f99af23d38015445e
zeeaf78bcc584c6472fd4d8b1229e2bb9db46a8d0123901cbaf35c3f74508995e08ca4435810549
z78c58ee89ae261fceb8975413773b6ad9e3bb22ca80f9a38f45659e04b0636230ff4773bea58d2
zd269ab6394dc959dc40d9144d58495fb9b27923d6dc1e8ac32f01baf9598cd8dc580f677a08558
zaa4bfd6bcddab3a35cb5f767a5024eea7a56047f9aa975849af0a0b2246c7605907ac45710ea91
z31240f8587aa72973434f696536aa9f4bf19f6e005738db183ec6674f93c756487e6ca658c58b5
z0dc90b1331c1f019b0b8df1ad3cff0eb53bf7dfa4ab3be5443e85eec0bca8240faeff489e741be
z13f8b4f07366a9a074b54f9c7f3342995a00922aa28f417c901b685a13dd82ce168644bed8e446
zeb43e3572cb8d7346cefcb9415f9039173ef7f28f5c79e9b9937fbaa1cff174999617fd1e0cb83
zeaf772c9d598fd1ecefae77f574596dd3b4b025bc62612290c8f0b929dee4ed92240885d500aa5
z4df3cfd516c634c8a418b245de6f4b57ae922a4b90bbac2bca68579ecba958bd6557506421d657
z52538e0b07b8b2f2e1ba498a1f2976d3af5510a25d01b0ac8b6da90a7d11897f7f67d90099de8c
z532e72fde5f796c709eaa9bf3401fd93a8c04d60246c98e61aaf3520d7638dc897d0a631a7a462
zc8606b26a4ca1a75db5ec3b52f6b7baaad9db86707d64165881b69d5a092f99b83a75918ce3921
z7bd732d2bd5a50119eb4010193528089a33f61056dd1840e64f33e6e758ccb83ea731e6b6fad58
z009d823845d14db68f8a00deea99c385ce142c6cf776ddde77deb958241e6a7b88e0aa594880bd
z198db026e3715c4e2be7bdb37c2c3edfab25fe64df7e00ec494638a943a18ad54e4723b23468f8
z315c10cc70c73ee2a18d1e2768c23fe6d03f5e3f2d27384f5ea086053721618e24056c9734ede1
z6bd53b910a7b4d872178561eb8705468e96e0a99d97dac7f7d389a9731d054ba8d420342388b28
zd08fd6d475d64ee7c7600ce86dc15714573213a3def5d1b3d68ae30da93634328545136c4547f0
za67e5cfb020dc1048fedeee2d865e3273639d2de9992dda00054333f0215d9830bae21c9a2f5ea
z5637528a0dea5da70a844108b2aeef929e2b6a06e4ab17a88a753803c915f9a3fe6f30537bb38f
zd8e0f4c8b934da20b97481bedd324774a118a2551d6b8141585bf54425fdef41be1bf4249f5f19
z63129198066bb7b23d7bc2e0f875d7e7c943d924c96d8821661e4eada4246bf59ddd33265bd757
z465a2312eed19bd2aee7fb1710f56f679f0b16ed1e43a5aa802b3e85ed644846e85547ef969ee1
z5cfd7a04b677c2e8eccf5cbef8299bdcbf1ebfd1acd4ef4d1eb6ca8aefa3a18c836e6df19d1f39
zb18b51ee18024ea4348d3dcfe9e64e672fd98ffe903a4060bdb1e85d5d1ca81fceea1fe9574d8a
zdb40149ec9af997423a5b3035deadfb6aab0d89fe843f1bb1697e21c69cc2900618b10e0bb88e1
z73e11f8555d7f2b0ab6df4bf622b51e656e73528f68783e7f38aac95dd4d5d4cbbf7eb077f6f24
z3c1dcb348ce8cd0a97d145875c832dc63f5bce74ba444db708435352a541176e5e14890f060515
z32afae09a5ae2881abb0d0b62ad99063956bf78ba7e47f339a0d75be69f720cda2ccb91da27d53
z57deec6417370329493d966baa00b0f89223a70d3d71cc2587d77a748a58184f75f182b4ece3b7
z7eebbde964e78f6c4f7711f271dd52d93c9c83f98b3597e3abbdef78fa6d69895b1ef06500a9fb
z47e047c7fe8bf85ef9cfe6d5deb85cffc386a8b4469319bca7dc5edf3cb7d378d18325ee23220b
z388003b061e6b96cd4beb77b144bcf0faa6b2e053903fcf959c7d1115a335b4677fc1bb66d7319
z74ee458537375127edf16e04d4f79cae4085015ea5605fb262eb485225cdf38a5c132aa01e210d
z2d17b44ad6f681248934c461b770b6a1102be45c717f60d7c878d4b9b4eeada5aaee4d09d69cc1
ze7e67ebc17ce0cfbe61b33d0c7d090f37a7fca9ac9b694d1b50f9e551f03f73cb46b6c1b2c3948
z3131c7d7f5278df9a067cdf810a2bb0b0784157d361d3066b3376ebb015393ce4add3d181ef816
zde9f83222fed7f07a07eda78a921b66d8490bdc25d348c22a5cee619aa25bfd30a13b50da342b5
zb9346cb01e43b80c452f1ddfc0d64cef24a6d930b66ff04c8d045eef0427a49a36d377fbb2c715
z4314f8559436c0b10a2ebfda14fcd129ce2b9764dc32072c93b7158470b58e63998d4ee14e396a
z8ed6a413a4597e51ae9b9b627f251c0537e7c985d303703f361e228c471e77ee273350bf743b33
zf7da38400836c5e621d80e98e3fc5b39abc1f75e684818a1ab56391a0ae9018e70c1aa5b699609
z1d72fea26d77085d01d1c13cef072309a4452f57f7f6d145b38c3d30f2d10b89d9f79975399575
zddaba7f8089e2d851f92f0a2d9eb06a3a23214c82dec21f37896aba2782780d0401d2707b2cabd
z29b6d8a239a92311ad8ebf02e9cadf3c8ccbe0942230213f6698bac6ae31f8fc4fbe6df5dcb466
z9e60f56517354508b05915b6da3da021657a6c4da84048c3551eb6ddfe0639a49f76cf4f06c156
z2cbdccb5cb68668fba145b8e194f638060c396da2359e954d8f707c3f4b9b25678358b87d66a9a
z9bf873a52dff085e728d968a4e21112733b439ee1e8f0a99a8858e973acc0d4fcee4ad240b521a
z2e1a00356d4ca38b912f9f5adaa84f5f236eb002af83957f758b12d74c2e92d4f44d94e21766b5
z1d005602b43b2cb75bb8454146f3595f9da033360fd9e7f3e657c064ebbd96094116b300a3fcd2
z155a8739ec47fa2eb9ea580d3fa8e4d483473f6beb0ba7a99dcf854e8fa0a8bd40aa56f2fa6af6
zca24c51b2012f8a3a8fb1f6ed65589bb24cba1df7da12f2f086c031f26e0c7cbb53e460f4f5c66
zd646e9745270b8d72c7ceaa0e033367c2df2e48f313f71691985fac328f0d5112abcf09842d47d
zae992dbda26c3a99cc00811ba7d1f911c5c201c5314df06f1f2e92cd90fd0b0e8bca00c65682ea
z71a0286a2058d9adbd15f935fa07c298dd3cdd37451d67cfc08f686c18f24e656c99d5a86aceb0
z4bfc9057f98af325eb68d8613c37c4801bb0c576f2b57d3e7417fe30a14af395d77c94cb2bd8d3
z4471336744fb8935a52ceee4e8995771bc71a4c0982d733400cde39242b54487dfaa8986dc5317
zaa8a6b340326f54bcb884eeefdf402618b8d9a6c3040348d105c034f3bd2180bf4c0e2e9de5183
zdafaacf9fefb1c1f28e23d29eb8524c85c2c6b18289ad8504607f11506a7212699630b870ea1ae
z30599e612a19c1eab8331bc398a56c5f09af79cf0b705a725d83a1815efa768a4126bd10e4a417
ze7e9c70f575192365f613ae1c7f63fe89296fb18ba1fb9ec487da91f4be24dd02e3569bd604f40
zbeef4418fad558e5743194cb33d6d15f8caedf921e28c3639d5e2b0d27677f23917122011c49f4
ze722bffeba8bb772a89e4c22586e2c8c52a20084d0685ff4297ef120a97ce4f049eef4cadf3bd8
z8a0889e7105b530c16881c750401e0358aa17ecc4918ac8e55131f54f93675ae8e30b60e796455
z67e8ce81bd8bdbe9b6032268ff4b35359dc92437dfaa95d6e2b8a4b0b66cfbcd0f99bacbfdd5ae
zeb7603d71672a819a789014364b5e4836e510e1af49f1cd9d22eaf8642fdbb526edea0925ff869
z1edd22293d25ef8d265d7f69578f00a9f17a2d2ddc29cc8fb6abca49f41ae7836302c3a5d34a5b
z3a3c9af388557fdbd676c8cea2ee2b8027b8be6d2f01d90487af4402d02285d02951246c72075e
z4c5a9a1f2987d4e001806a9c37fa2fad1a35dcb3f6f8c9b27744a3a8533a4300eb3e4f3e7ef1ec
ze12172c2ad9196af59947f6ad159f98e3f099561b1eeb3c634f2836421f11b080e2fcad9e2cf8e
zfa84a6f2bc2776a64c591e5ca3c54228ef78a9fecb6a32c7744da9ae07ef30d537f02bc62f24fd
zef805309e22d31745a188591c0a34da332d4f49565517069aec9519a561420e2b95280a633bb00
za035449f48a980a084ed6502923a393a713b5c5c94816ad4dc48fc32696360b8f45b6e4570f6ad
z98cff8383969e0b07f07ec976f4775c8d4f62b8b7bc9af92ca8f6ee93358cf7c46c4d66d77995b
z1c4f57a6939afd0923f14c992158b09ba97631feb7d992b849019cbd9bead510059f0bcc794d05
z3edd94836bae434ef1cc0c82e76e192cf003640b4988c4ee781b15c7a565cfcdd3dc1191114d51
z0e19d7f957f4efc9f8ffa45c1ebec1f7a429618c97c66e8c3844b288c83efe322ff6dea8461f28
z026a82f9fceaaf403d625a682229049f39816bb31190bd9bd61a4c4ac6420d1bdc160378cae308
zdf6d48aad7976afa811ad27c876fcea583d5f136917bf519bfcc7ff328f6a7bc92881222cb533a
z9874724aee83b42371ea05c97cdb6d2f4b59c7ca80e7d1addf55dcd7bf03980d418503baad29eb
z3c01edcf1d900a88a911695fae5e474447bb57399528baac3f611ba8095967a75171506b5d22a9
za5ab4ab0f647ff86f0a78c1a8688148ef25b35c42bdfdfe72cc19f9251e92848180a65693e9962
zbd55a7d340558cb1158e98a6a33b361c0d583ad7119e3d575e4d85fe3d763afd22fea476ca0d3b
z7d375ee9fa745aff77c507c9666213af431c1acdcecbbbcbfc49355bc17c7237b7e55d48731d26
z694a4799f4ac0a73eb2e7debbd27492042a28fe4d8bbb8b7933edb2ded117086f9ec0a540f95ce
z5d3a56da1bc56a4faa275be0d4a7355bbaafb1767902eaf35664f1ac544cdfa4c12a6d487eda12
z3fb61a1a1c868cdd28fac44b893a61ca48eb1ce4507a6ec40f811b776cfa1d4bd17dd5474b7675
z09de0d0046bb087f372361a91653fb19431bd10f28f8367ce65667d59151b02211a84bf07a7d47
z62b65a0900f9d3cff589409afe5c3082807dfa15e7e58e162c5de032c5df58a1aead360d12b7b3
ze842110cb5fd6ea61fc6010ecc1e43b4d029466e1226b98f7e9a33e7e730f3f1139a76e3b6f28d
z996e7d6c2ace7de2b428428c13e3c783f18e315a8f6c3000d62409c3a132d1c1bf8836ee243b8c
zf6e0570ec9f6bfd56ff5eaeb1359a213c25d35564849758f0d05fccc6f532813fd60bbf3f998de
z2606d9c5ae021cc2d94e939d35c6982fe0779508f8f63ccee3db474768e131c852f6070f18d7d9
ze70d91fe8404dfabb08253fd49e6360eb0065f55d7c5d8e66e30f430b216b1f1f4cac22270b433
z96c2def9c8f1f1578995fc0082e4e5081610e309ec7863861a3fdb4b966303345ce1c377edefa3
z50551393aa19df2d578424b1a75b1fc4feb5e79261c683762bc5932261f78a4c2b54776f6e4b99
ze159edc77993cf6bf2b94fd8c48275b912c4148b867d7837cbfdfd095f456bf097636cf4c4b789
za3a4ddaf11a3dfe6002084d73f3899945f4aecf5e54838501579c2f14b227e3f3a4075c88ea6c6
za2996a7b353fe66f77be8455ce3cbd125ff978bf1bbde5d27f20ff75a5f7a080d1e5a743674140
z355787c1444a653536bbf7c688c9d5efd45d47273f3f95522f5a6b335ebfcd001f20af26949377
z48fe9ef8a3b97cf8b1c4a5a102f4f1899102d3bddb43fa04db16bc6df2da2e1d359470dcd25e9e
za966a651be387d14bd2de32f762fd432cdd1e903139d83d70db0d92d5d89023805811486bf3f75
z92015903c2b464d8cb9d9478dde033cf568a618ba79347f1fc35c5db10662e591973c037cc6fb1
zfae5b213824ebd1b626ef9ae57c2137dda43cb4563ea73c1e8bf6f1074926ca7b97a631d46c31c
z5bec4cedb55c05e600852b269643dcc53d9a6a40bb0ba92a2237af5116996beff67602fd5364a0
ze32e5ff988f40cb6b57c76297f45d4b05dabe6f2bbd24f25354c7f211351cf0032430328835bbe
z2f9ce2baa81ed33f223df53432a7cb1fb98dd359ba71db2fb587837c5cfcb0122eb8df11b6e718
za527ada6a56d06acca6f57c2026cfc533c590c0adbac7ecfe120b3c46a3286d5b351a613b3613e
ze601a925ff58d0ef883f032bfecaf6b656ee001192768523197f352d027747465595f88afcafa5
z8e74a4e2a3c6636030129decb4c8b25af1ceb0909d51ebd0763afeb3d1e5d01f896dd110d182f3
z9c1a1cbeddec4c412fc9fdbf230d0e7c7942812ec34197e3af756e01e12a5b8cff60f299acf0c3
z3fe8b14c261e3b7290c1caadce587649886087a3fb2ad8348f56d44c25732f16198fa7fde5ebe0
zf9dd38b13ac9edf3eaf5aff9e44b3b74573c70ae88a42985e76c41fab8d7f2701ebf6c7bc23e2e
z35c128668d605e57638bc319aeaef4a0a1890e0c1f6be37403f6618a3ab33352a13aa6754c295b
ze18f4e9087c239885f2fdcbf684e5354b18e44780e451dc971a1569cc2e15df05545fcef9326ef
z807914429c943b114226e1c057e38f44e99f432844a32fb8178e5af1f84d9d220dca2b57a6b623
zb35ac183e1847323913a83e7877396b5de780a7a9887ee03bf61a7f1a01b22d3d137c6cfb6343f
z23ae877e1d646022c998aa1a0c9c59d57ba747fa1e87ebdbf7ea4af682cea3bad0e0f681f4b155
z6674e3dae714219cabbeaae78cfa1fe436cba0c3575e9806db9a0651a406b63f411e8655d1c80f
zdcf06321a68509bcabe214dff855ec718cd2e059111775dbc472f6cac19910a70220220305847a
z879408300ff94a77d8a8fecf36f7c217c31673ec3376beae0e9707b50ec8f0f374626d9925b7f8
z6cbe6083710e1d628b69c1f98a1e6e591f11ed8fda97a48524fe5696509c0993414bef742b64d6
zbce9a6a81c2feb3f51db1a4d61b72788b995ecf3d562a0f77586b3373d43cc5af9ee3ebe28870b
z4f3110fb050e364dcb23691cf4c558b371444251357b150c1f4a9bcdf9352c7d00cdc1afcfe32b
z59d531ff5c75cfdc937702129468c6b89444882030a455704be3576a629a15e088c93921a91269
z8d08340ac081c695782254b2353f36b2aa10fb311287d786e38a8879f15c4fe0480f72d5581b09
z2af1cc983a166971e133bf96a222731fae4247132b0502a7db8f62965152ee04609f452c75178a
z8295dd446c1d547e478da53cebd92b3f679188ed240d996764c1f8c8b7c89ea2b18db6a62f42aa
z1e29cba21363994ec073e2527181ffe60a429b0a25f90448782f6bb057e7579e20d98cdb9a468f
z64fc01951c04bf6d1b90266bed3e3ec41247506f14cd4fcf8a1b84a92dba01063ecf44b17a7a8f
ze543831e4be37482b2ecba2085257421f60245b1de5dae16ebdde7b51071f9f372e98062d48dd8
zb2af95f24d5582d13567d71298202c04eb76da0dbcdc7695e4a4673d1a7c00409f5cc2bd3ab328
zc69b23b0edf4089e1ac322bfeeb9ab95c99783a019425442adbf5913187121ae793b1d173e35f7
zdb07071499626ff9c6f26beaddcbfed9b9ad1b1d8229c30419411a38fd2ffacefe4a3917c80474
z0b02a2a16705618c7aa37f381e6016879a9d92e0906d2525a7b94f1a81a6072338a491da0625ba
z39370ceb51b73cb7423f7f7ff07f9997b3f8eeaace630e73f5478b98f8b12827e4a0751b0660fa
z8ee1796b975a54474d7c5f73122212f297759ddc444c144df5d9319adba231e41df8722efcc4bf
z0f5ace4b4d685220aec82f2eb4670d73375c5a0d7678584fc5914927162df25537df3e35db634e
zb8047b144a571fa899b146fd77a497492b4c99cbbf9574cc18ee5d16ec43316b07a30381d1f5d9
z85ef15f8ebee641cd57121440d401749176489490adb8bc69147892cc751fddbbf4a2d7fe30f90
z387ab4226a140a27fd6ff710bc85e8865f431a3d049e30f20b9fc882b8a68f2e0671b248fb613f
z81436527b6448cd1b0514e94a3a86c04a7ce7ac5aaa1c3e22b159587cee44ac2e75225bf923ff0
z3a0c727ae2cb3958df364aea7b1e5f6b68f9b3719d38b097a3cb396925b9269580fab1dcf9c2be
zea8ecfdfca065b474a81d5eb1d60b9cb6e1760bc06da9ab6fb47e6f08cb8159f1069401845a249
zfe5373337e7858561059660a99002470eedbdd13d17e27f5b8a9d584e89c5e3d70a1b8df71c69b
zcec5139c710c03b187d08210e7f3accb4a534a5069ca87af65d673177cc01d25de47d90c24438f
zb11adf4b8d4ceb192985314efc47f6e0f3718fa08b6aaf37ecc8fe944c8f7615c03fb7e9a93b98
z8adc04e402c2eb372a2c2b59130b9c5a46b712269f2a191fbd4a5d768a18f20b03c145c9d4196d
z2d7084bebb51bd8343dae439d0964a47f79274acf52d6faedd000baf63f5c03542ce4c73b49c6f
z43f555f6d6aecbe8faf09de6d9703f7096240571d7275fbfc85782a9e90590cbec14d690aa8605
z7604b9bc250505e7bf680cd172c5a3498bc794c8c155b28073be8c3dce36fb5ee8b91dd3035a16
z79037cde3aa20c9400001bd6cbcba945f951678f5c7a5f471e8b7cd97a21a6560c39b12a6a0f8e
z871de8ad994a6e99774d799a7ed785a21a1b7c0ff5d69de33dc10e31bc449a9eb4b300d9e2cc0e
z149acd80005d61460932e08e77ca91d8f6984117c51691ddebbd6991f18fba212189e0ec2b6b74
z838c896f1c9c6bcacbf4aea7814d69b46ed3472fd9c5257b2608833c126cd4d5af34cb074c02aa
z4f0404c8489f92a3d7219273a1546009e3e5ebfaee76c44b74e049404ce74d5f261c8461c22c7c
z88e90bc9a5d6aea844a40ad2556ec17c1f3d2dcb45c8d5ea7fb506b41ca13955f41278c6183b6d
z3c121a7e20f67d7ae96dfdfbc0b619bc2a536428bc0836987c46fc020f2df4f97bf9e8e4dc4d46
z7123cfc48229affd88e1645ca27bf48e31cd39735ab3d17be4df4fef95ffe4a0e0367d86220591
z4e9dcdc5fcf6467cd877683da2a64b7308051f63ce9f04d631fcc42ab9b311817190a79abf692e
za7834c82dc074eb449e83515350092d995530ccef83d62c133e588c7a82b79c9a43162e7f51609
z1ab8e6f57285112949843afbb745c910a001dca1c23ffe37fdc7c01b1caee3b3247f40c38c0d5b
z6f7e50619cac7be4df521acf1818faa8e3caad06929e1a12dadbb8addfb6638525c448517d4118
ze25d254b0574ba438acdb1b1fcac6ba62287032c57f4718170436114d9c53add0e579fd0539406
z55cee8d0d30bb987f4e13c91e2098a81be1c54520dc347fe5587566b9f63ed57a37fccd58ef085
z74f2e529ca692c50ae00d825ecba49c529d8e5f1906dac558329e87cb7d1ab9a4c44290c2c311f
ze0639586addd1a58fc2711d8fdc99a5eaa5a6eadd01a0280ff7f3b6b5285317c677c05e315e87d
zd5e4a6b3ac38099e17a07cd94d5ff1c60438f7b6aa999d22c132e1ad512f171885a46df5b6ab24
zba2d6c58c070aaa7428752963157e8e8b63bf3f17c90d6588db2061de6b01ab6b692256fc518a1
z2c4ee6030564a2011af62a358b837342641dce5da5ae5c70141e6471ea6784fcbcdd3866e79a81
z5298469bbb2ab7d04a1bb78528ca1dd4672d1603e16630eb8d0e3e01495e36328a3d678ea1f62b
z707503fb04224c0b72b90edd7431b6fcbdd4b37ab7fdeaa2c0ed56c528e94b2891a96248e909ef
zc0bf940ad8115af1da3ff7409062ae6adc2def755cc2494dfde56ec269dcd8e979615c26b6b89d
z060b451e8ba485b8de9baee27a8ffe62bf9b3d352cf41dbdb47eec23cc86e8603cbf4fc05061f0
z647a4399cf9143aaa4cbe3c78fe9e3c3ac3953a0d1acdabe76c174ae618f58b5e4c0e2694370b6
z1ae97ebc02f52a7389e30a5e1eeba4120c53520720e603f89b35da9b3a66a97c11dec00e7a158f
z9ab6aa5bd06b9d47d54490a7b621759b7ce66cb07c7d0c95c3f750f5435e805fc4333f5dea686f
zeadcdd0c4dd50152d59b3eb5c92c2dc367f015a4b55443a586586d5a81af3d5bf4ea4b6c9a0197
zd6b02abac0c84d59de6ee41a99d6e96c8a467698b7ee5759e4b7a48ffcfcf10363cb97d30656b7
z74b159f388577100465b40078fa390dbebaf277eac9f8b21cef862ff1295b44e1f5d6910086628
z0d4f9a880369fff26caec430640b2403e274a18a1a880b657f2c5b0a909cb2bf53a107df82592a
zca69d826c714d9e02a0a6a8fa0ad4a90c29fe56e897de0f0d6f435298189a4dce94d2bf777c117
ze4f6bb81d1894e88dc927a3bc9c82290b8c14036a95736a636a02e212dfefbcec2dedc75482256
z21450246ad5e2e218b2f04e9f6b64220fa5832ae30bd1ea619bc3594393fd427f8ddfe8be90bda
z345a47c0c9d71bfedb60fa4eed48c32b455604dad532d05f394b713438bbd0305d8dbcc36e33f0
z653c3a85fd3dafbfcb76cbcc6d5bd9f06c8215b5172306c86794756fe8305a520d39099199386f
z4f0dcc01ff29c798a082cf7242422e24fb67843d9a25539f4e870b5670d1f7dcdfcf5f051a032b
z6b40b91f50305d2ba4b00299ae3ce7814fe129eb2eea195745a2953b543df363e34008e9abe7ef
z4ed346298589481b6385110b39cc3ed58591dad0d5793e4f430cc53e8459a2fb2bbc91b7375758
ze9415ffba9585097bac8318da21864975425d2c6172c8662c483ae15760223a3a820b6e30797b6
zdb0e3062691e3932220c0b4a9ebcdee245a836ddab26abcc7c3bda195fa2fa596674a712c8f745
z8b61c22d81f6efd4a1952b947d77ecebe2cda5d1ed2912eb6d28d9882d3e05993a776d4ae1affe
z21b707ae3f5c19d4514e6e71856b284f4ed9924ae950e367d55a0d6b5b6bd8d9a6aea738989c0d
z86ad18994121988ac807ba389df7c682001b4298f4d8b90fbab5e9f049046d17b304e3082071f3
z9997a5e90881215ac67b55ad2ed38f9179ef3697edab2373ef0b7cedf81b589a390469ce621f70
zecae022c31e7b1d7942f20e2dcf6f4a59dddf3d2ec0f438855c5b2b51bb8b44511b98234a4efac
z07e3e21cfa661b5bfc5c4c25d492114cf7d0f005aa37a0233fd4cf2418f401b3205069866fea87
z2de7ec0153cd99b543a1f6bc949953ecea121083233b0ae7e40e210688076f5d30b2d1a091d72d
z163d5ee19730fa91428639e8002bc5506881d62f76a0c06c164c017c4e2dad17ce7389bf53cfce
z8894dfa59b20ebfc0f641bcaff58db621d5aa40add97b2af25a1bd5f5eb64aba8dc074dbefb394
z828ae7eccd7efd52cfbaffcbc12809ac76a4fa2c91d48fc51d237c868001143619103648349e7e
z892b7cbd2d7c70ab6122437cb411bdfcc50500bf4f900ebc9230e44a4181193346887092e24a62
z6e592b6b98ec3093a3d50861116b4dea0fad3887a47fcd8cd3062e209377ff238012bd9358a884
zbfc71f51781a8599cf88adaa349015fb523bf60376af44b19237e1555243b5a9438267fc475e70
z3abb744443749045ea8bc3ec339df96520f8ef4ceec56c2b4bf31207360f178d41652a7df57968
zee148bfd3997625b8b3d780761c980ef855fa0c4af52ff03a4348f50175e2361b24035be39a7df
z23ed03643a91c025adcc8f6b0d7cd54bdb851a235eca9f80ed2c27dcb2668272aed574ee76dfa9
zf3ac85509c9fd47b1aa9db5b73da6420aa4de42712ad8e846bb9988bd7d01c453c4eb25aa6078f
z0f5e3fa90c94b1bf6396a03ddc017319bf9bea027015d5d31076734e0d7d149f6a54fe32e143de
z13de7a825b89f77e8fe9ba782cbcbaa0212ceb6a3a4e069079d3b00764e213087765da4edff939
zb0ed59213f11b1cfd21038410ae78b3eacc60d682db672fa5aa1c28f8340188ddbca400d84f823
z7feb3623e294c85676fd936b83c679c387891a0c2ab98592587127a35a366f234843ee60e07667
z3fe6bea26d600986470b26fda314c50b350a00c90c84ca96d30b31a19c69a83eb802f457a8e8d3
zbb819e47abb137d0b03de538f168906f8e2730f1a95fd0f75b115331e534b291c1786aa8fa3cce
z31ff42910a387ee320b37f0b730b4efb914de0f151beb3826ce3784c60774efa41f63de4d77c7f
ze352f80928e4ed8d6c0465edbca837400ced7baa771a06a8988c02721233790710ef4bbd0901cc
z54e21ea9e40364a14b0c8d97e46f3a67fdb2791e16d4e0570e46ded0d0d9724488d3ed66cf921f
zda889a437a24ff99671f62eab47b997400de2d458100c633d4b5b839a06e4084e5e6aff39e1311
z46c643356dcf76e97212a00bd854a58c9db1ab96236a186e9678f2dc26a2d3cf322a8ccdc0a76e
z895f5e91155fbae929c79ebcd99226341400c7c4612735d5362ee87be49e5edfc1eb5d51cd69c0
z1c538fd831082674f4db868ab152a78a308cd070df14f4a2e17b72a08fe1a8b99a0f362bde2e7a
zd9f2203cc7c80e86104a2a4b5ab84eb61233e098a6b4e18137689141e6a000eaffb52af52cea98
z8a74ef24418b09b49590f1f7fcb217e6c51962e59a2e900c67b1fc392d28dd97e51a1b7f702e59
z875c796643c253e8b2a920699d5c2dfbb02a3e6a96ef0758e3e8d86d944ee55fecc0a510dce816
z2dd159484f10b7b59bcdd71f1ac66b112aade553fb19956fd7e8f3839b1362473f71476037d706
z5c931327a57dc366b298099f308cd92c6c68dfc8c9008b966ff0aa32e235117af902d570a0e3b2
za5796cadbf9cb58ecd8674e217551ee23bf68a8d2f1927e72364e28cbbbec35bd1a4da67f7461f
z06cbf437999bf3d468069cd752d4829e9c8527e297e48f6fbb6256d6d614e2aa3e0b320ac66b87
zbbd1db1c589bfa0e35b81d3375429bac99e900d101bc1dfb37bc038d3c1756f2127ab5b6a10f36
z69ef889722431814aa0f8dcd28c70bdd7f4f30a6055b51a6460b57d638767d47951caa022ae64e
za7e7b17c8480bb113bd7ed213c6ce7ad5c056dc84df357f95bd531a34145568d4d205b92bcb143
zcf81470218aa1e8d9a7e9f7c9a23abf1e9ada46d24e0e38322692e543a482447d130e73d2fb38b
ze91d69447329f1c05d6ac050538df889e07b24682e903d8998d0582da9befb3cb7b94df15ada09
z0d1f6692c11b810b0924cb5d004222b6ad1216b62a06f13222cbb6bc2936e8cafc788867ffb35f
z43b492901c86e342ce89c7f10f314470fd2d5a308e53a69a373eb3ab5f57ff30c219b3d79ad7fb
z15eee013d219ad7c1f4dd6ec05f6326b8c1a3c966fb30d8be47e15628a613c480d23d8bfaf22a0
z6a947b8327fcc0a1cd574b67608a53760f084f1e0207f3a3258afc24cf2150969ddd4f125a6c35
zf9dc497cd7705da6e1fcae8e8b46c342d052f893c8dea525cc1b86deb3bd6be1839a19abcb2e04
ze2f51d5cf1f1aa1fe17b6aafa71209a5a96ddf1e48b5708ae4dcfd810bb04ba963c117e9e6c75b
z0910e98a4e67e7f4d7fd2392c6a71e17e1bbdbbc0eafdcfd729ade4ebe3f1980d0f66e083ef3c2
zd05861732fa01393d361cf2d6a996a9e6e05d2139b7d42224c1403dffce06fc269cd6b399c7e67
z7c935e799cb8ddf3bba9a363770c9c7527d27dda90891f48bd9aa858457af95ca571f9b853962d
zf18a54d98309bf72a1d667ff22bae80ffe91ac3c5ea3e1ef6b2ed45cae46b7d74e9ce95eaa035c
z875aa6ba56850e3c1f0401ce1a466fcba476c10de7b3fdd7dfdf78ba4dca75cf331c3af24c19ec
z8c1183d5ddfb0df33138bc6b71f4bbe80fe2145f23bd508be05e25e2cdc70715f150c67e5fd38f
z7068c415c9bbe398257e032810be62ba054ed300d977aac78672f566586c5aa2fb70d1fe950dbf
zb5b03b77ef2bd94167df0843485c3025621ebffc726e313f0fe14fe025f9ebc7ed4a3f0e8966df
z15ac4c14b6d6f85f0b6002e98d65c0dff193be137fa9b786b52032273960e056d1dde8883462a0
zc862e29739a4d5c3a411362679a59011ed94557cf502b3231c151e25366483b7f91aa984cd7495
z640802dc0452f8ff8a696d13f27d45245266f900aed222916596e7e1bcf165ab6dfcc5c4c46ec9
z7c74dd2e889dfeb1b272a7616b2ed40670b2e9737dc38cdc834dd612b79d97fa033b1f4c73d19e
z27e064b805a354fd8cf47b4b521b1a213584c32b14f20560a720150e60651ebc3554fc31b38173
zbd851583b6ead9b339bcdbb2b6f6a3f31dc8676657575f9be85ce82629f91595e3c023643e0037
ze938fec9a038c9b11090d8a1a44a959f9987ab283dc9fe28c48b64ad8db816f5d976693db34edb
zb75bb6984ef810cd406af5082423abbd3f7d3eed8f6fd5a7baf9ed7681f95da8919a4a61f594d8
z12e82961f0e8917bae926a118dc59bb6b0b9bef88ecc3a4438d953d1c7f38ffed456342b1ee152
z735aa0da43baa44af396fe567ec3054437caf286501eee4be8da7647a94fe205e2ec56ebb5a6b9
zb885373f0fb031ae3d23c7c032ff3cd02771df8f84adbc5bc85ebfff757686d9d7faed602dd16e
z2c5e716108251c2707f57431609e8da6ab92f0e7911727b514f12ef32e4c0429554cc81375395d
zb7834e5e8dcb2177c38e8d25d84e445e2c64deec7a9b60a0af2c82eba28f9ea4305e507b7976be
zd137008307fa8c77e82ef19a64388ecd6403eaebc55773927015230909be8993dddf8870901b96
zf37a8e8484c5ebf802b789c4929194a46fb40b1fede173703fc28bc0ad184742c9497721aaf424
ze67edb34801fb03488045eafcd2549124d04d7d142377b7669b0ec2e150c4ecfedab713c7b5b71
zd0b9797b27d49e9b999bf3e524ff472ef456e776bdcf9061c14deaf4932cceba0bb20a90a0f4d1
z904400ab553e38a3811d15b5a8560847de60c28cedb018b0fa9e39f8ff8ef957ef3f48fa67f808
z55f29edcace7adb64bb7c5a8f3efe0d33e2d5695f9ae14463f8f95663a332d3c292e1c76ad951a
z749922b46a2748e9578ae31c4f5cff47de83bf295312e2e996bfc127d14c98067503ad6dd05169
z4d668cd53f922bd14557acc0a16e4ee7a2c067a94b065afba8b6b5ffcc95fd5ceb82afe988f3f5
z8e0c5edd629d5a09d781b4753a6e5bd2395a49865ea254dc4dec2b01fa080d4be4696575bb2348
zdb77dfe634173702ec6620423e2f4665adc9018765f74673d1f96e7eb8d306f5bbc7d755196663
z8b12bb729117ab9ec370d4de63222f4b426fe75db488bc1a88613774c03e808ab93def02c4f228
z16244869693e24599ab4f0a259f4345f311174e75dbad58398a7b9ccff58ce032e8ba34f7ae0d6
z0add8b396f7b0d29ebfbfc13348e2b02a04b6ebca3beb1979d2d46bc1d066fe27e3b5de3e6be41
z70f1ad06055ea70cda85d47320338a601b2ded1b8a5d5a6c8779986e060f0c0cd5d2da66c7e75e
z9e3af5d56baa4af9d45db0b239489f166e45d659f074e3b967d5bf5aafd956f2fd29d609cc4afa
z9b267e8a2f9d05f21370c6b730955fd62d8838fc0796c0a3c0272b4b759bbc23da5966b13d0b7d
zec2e0ff3c5605c641ee7c9fde892d76cf36e9304b303aed01deac4763064325b6fa53fe3f10f32
zc7c9103824a734d0429ac701d45f7960d86780a637c89e40d31a4ab5947054111bb6a6e73d04fc
z7c3c545fec0fbd42f229440c202ce68fc433ef2e7909be52c312b24dc38576cb9d78b8652c7abd
z9c363d2a7382ba01fb6fb6dfc7958a90d5395c3fffad87ab1b4cf0f1df7b5a7321a40835508d62
zee62b4ae07e1ca4ff58759978e11da3fb1263923a8337d00729a5500614a9673d41da1cfd940b0
z8f3ba103eb82f35944db724036dcea63c9b969516d9d9f9f35d66a62f5f11cc02f536ebbfcc86b
z4c4c286f1f73bb94c8e513630865ac78f5442acd221742f3eca48c7126f4697f5998ca5b9f1867
z909e088e323bc0e9026b0b6332f37da2fe7640fbda5543c3ea46972262ccfadc1e0756a0ba6a6b
z3cf4caca249304856501f747f297fcc3d2c68b53422f575a354b2016f76e597db09e7260b754c8
zdfa330a266444ec53c9a3dd044d475c4a26ae277e5fefece65f6be8fb21051a5687f976b7e0315
z02241302e1fbb4a8b7064689aaeba10495474a3e2598dddd988f1d52808fb3705872faf4aee833
z2fb0858a4787d50b568cccaef101e1f963d4e0b065142d7b78c580015c0d9473034ee5bb4100f9
zbc77c08ce19f3982796559cda3f12d4c0f12b3984d02e72522fef5032c72ddf1070dfbe87f3f70
zc17917c1078d7e90e5838af5cf89d04314ca8a9cbcb250d8f6398129001f50dea80565e7dd239d
ze5b0eb386a4248c22e6681c60463cb8c92c58312f8a501687e01ebba68f190b54a3cafba7756a0
zb162d05667ea2acafeed77d4aeb8dfdfdc972484e7f9a5d82c142e4fcf217df82864873933e4c9
z99b1e1ea85325246836ae68670b5aed2f73e246f60c787beaaf635e84be276db84ccba67a3ded8
z05ad2e1deb351ea9f8fa35180575041e59b2d6bdf7cb189ae0b0ef9bd3bb9cfa338504508ee6e6
zf31402b58411ef4755d052e538bf4ad89f79d309ca191df04dac84e0bae53e5c588df0151eac5e
z5169191bd30697b4980da590c054ef16913c3dd78d607afdf6ef6f05dd588d9b5669acbe9a9a8d
zc7925d1e123a88102f32238f97a14eba3a38d61f72a2fe8adb51bda8eba43dd8bcc1f8d4efe6b6
z2730ffd9047c09b7daf3fdf91aa9784f8432fd0f4d88baedfffa0237615ea162a14da2df0e7b21
z84e72e152429b1d142940d343e942f6a5b63400f2845223c50567f67c899955b26f1f5b62bfdd0
zffc9bd830685cc31721645563c6e365ab9064e734fef3a298cfad3f4370eb2363811438a8eff57
z1c04dbb068397a823671077810f5763bb02c835083e074b39860f7c2c43392f0e35a26eba04750
z36d040d8d0025f612d9fe2f5554a3e401f1712cfd4799c1cb91fb6a935df0c9522ad281c258790
z416914cb1d692e5d4ba9a1962f2e8e825b0ddbaa20e047133cb95f1e898d40078f6068429f4ca1
z62c644eefd634e63568f6205eca2585120ce73608fbfac51942c98893c48be88f17be3a78da408
zc675fa3a85806b309b7a183975f90b062c09a484f5b025b0928bd60c57d126a27b2100b9bb3b1e
zc2161d8da217f2a87dbff5a3756e978ab13969cffa13e9b32a5b30845d39442a21ea4a37cf2777
z161636e9eb1ff9538186e5b35c004fbc79a65948083290c96adc29b99cbb6aa612dabf67ea8b47
z52455aff0451ce61c6089cc6d7b6e4aac206720de36671e4fd5131f681a39717e6ac954217cf61
z5942729e1e5a3ee4a0ad53854658a8c46cfb4ece24af8a6a913bff7502069ab968e47d7a01717f
z3395bc253eee38dcdc751529ed628f7445cb84850b7b53bc72fadc4f7fe0f0c85aed5531ba210b
z6f76eaba9ab15cbbfb6960823995950fee73c72a7db774c4534d9d77a4855b918397513d05ba58
z340b45d46e71e353fff9a5ad2d7d71244016acf7fbe49ce2477bc8ecd750c350254c4c050ec392
ze3662755fec94fc3d804f2fb123964177163d4e4147420793a54a59887a215dded58e52451c7cc
ze15d2aba869b6d9a114287bec55d3cefaa4f20190e088cefe770ac87af70075bfb94e818fde929
zbc8edbbd9f32516b4f35b3649f4470796b2222f76b8be826a0e3882cfdbead95e1ecbf64754ec3
z9911bd32a777ab557d31d459ee9344835a01e5205b49060e29826d25707b55050c30428e638420
z55d3583147d1956666c2fc8903f619599243ebe95006439bd70888deed7c0f05b17a96ae473d0b
z24df4e0c1fd80115696120dde24ed000f44d95cd58ce424b078646b38790c64dc1a02f4a5e9cf6
z5c4a9e817bb041dfc9e77cdc6d1770eb9cd8f1eb8578a80c0442d0f55d99f16071f6daad1b354c
zb80b1d62d2bf67b206ec075b597b32684fac3de12967222bad1e8c5eb041d666876ccb6022d4ee
zb904e49d510c4c7dc140dbf1553bcadf45d08dcec7af239b58a2a464164611747e5168a7d91234
zdc14800a1e8f158b287abf72ebed587bb2e897b4f777bfbd5d4e319fab684be09e7698ba858a04
z1e71552652458f3532ae0b6dff3d7dff5410d2d6d97d02284dbeb1868f143f85ab6073981b092e
z24136105c3f623396ed9bce0374d578128fa98bf108cd519548c6a3f99eedc138d0b3834ff5f1e
z304c96b6ef19d44fb05a113ff96a9463bf2db31273bec5f8b09e76b2510559d0b9a1829cfe56ae
z804bc9c394068033e61196bdd1daf046e54c2a8b52165221cd890cdd6e290f929fe9db8e502984
z33e95c52d389e80d502b542024b8491564e87a2f2b2192260553768bf3c275123d5c1158e97f76
z305501c29b5372b9334eead5ad63d30b02a46381c0afd08a1d3d38aa3e54946cad4e28d5f17cde
zfea5f66db68a5e486dc539af50050a232ca8b82396109198391e4ef87ee7572f63accd728e0c1d
zba532b103bf3cc92f72ff69634346a8f90fb91a7ee45367068bf7552c70558afc36e595d97d609
za131991bbed692a186c4946a874504f27782c880c05bff4612530848cd87083eadd839b3e46612
z43860d8aedbc87cb695b1606d730eb7de50df3b7cc4019f282b2d1395f96f2356e00840c3defcf
z653d9c281dbeb25b7421d28675f6843d535242e3525755f9a0525600d6edff68e148d3b9099d13
z64d9d0cee0064228731e841bd8a7e3f4eb3f7f0a976a0bb758c422b1c8d2f09d1c037dab821873
zf83e6734d2dac7684cca7d8cd48ffde23ee97c6b7cc7a69ed20a91fc3afb84a293a2117d28748c
z6624cb8075734241eb540eb96a6f7d8c9fb4b72cba759862d9920f9d4afd1db8c01654f4654666
z8c94b826de0eb27143a39a0f88d82e6e6ead17b57950ebca085d84de5d2c85709fd44b188ca837
z350da2d9031e5fd137f692cdc7009b9f77b7b5a01aca757b1ac7bebebf963956f375b8d67cb4ef
z419d13dbde33c1c970b55ac5f616492eaf7d25bf167a7bcc55a2fcf41a8ff9d438b8ed82c03785
zceb08f113915295cda5dad58f6d4e2c0b0cfafc3c9e1e35851ab53e4afe4aecbf9ef07dd940d51
z1517d36ad180ad1d637904133b76471460ae122bf531f0a5dcaf7ad1471db87cc2f180f6c9e75a
zd5001febd257934706801ba48aad0f6a99c8fb8932e890c14bdd4cb73617bbba416b4e64cc9b8e
zdff75ecfc9be568369fd764ec7a544389b443c5816f47d0446ed528872b5f91e098305c2312655
z52e4595933c6f17d08185342701721e769cae6ed7f4be4194defe6fdf665371a4901b2342038af
zd20f0c43f23098664b23633c29236c36f1cec6636cb60ba736f182e207fc903a504614b8a40287
zdb1148414179794ed071b8835180dcf916350795c955813c14ff3e88f48c2f26b203d7fdc19fe3
z99933c5dc2284428fdf601774fbefd285bb748a246a36059661600d81f4f0ee4058c3a2e8c1a4c
za8a2f7d974e01a5784704e4eaca0059ddbe0a7d9b89aedda4685a454819f27c010f6c98b71c4fa
z7ca35c9041fed58ee2d17180f27c3c41abc8078440b6734dae8589ac44f88eb42969ee85d548a6
z8525c6b015ff97959ede57acdf223e52730e1a212a1d769975254c3c1fef2c74c47680b96318f6
zf4a94cc348bc1832e4328bbc71ab02a38e1a333d48ec08d2e3eb9526983f0a64b3b9a6e374b952
z7b5715a9924970e48784d8fa22da06e7480f09b40d112206712ae1afd9a6850be2b94092524444
z77e9e06d8fc09ec0ef167418ad16628a50feae5a9286fc405eab1252120a6b34504165e86381c7
zc5cbb156aa64c39f58966be47c2cedf8f116640cd09e2f4b54b299f67520cb9274fcceee4afee5
z41a6e50f76bb1e550bce8c92ba51e27daa12f86b0ab0072caf198d1043768ed0a469edef7bcd75
z7f29f24c8a0ed983ab87f8a6061bd3d2efab166a8bdd7a60d814902cb5573f178a7e3150bf5b4c
zc0aa8fce1f2d5fe191cc2aae5d74cfe3adfe835e3ea6b839003ee498e34d9dbe281a18ac60f05e
z3fcfd025f5618189fec7e1c30c8bd7c42a6fa98ece6d0bfb8c5a86c38129e52c9730d39b9556b4
z38c4f2dd3a3dfd3da0c699ee54e0eac21e0e8107e0c112207a22e55d325b40effea6af5225d318
z6407552cc50a9abdecbb153626967df8dd74bcfabbe514ecf470aa7044bd8ff9cfd0e219800ecc
z6b38e2cb15bd871a6fdb198ae7f8d0ea48d07242a2b17f7feb2e12d8505f6956754a1fec10351f
z7a4a8b8260cb978ed3327734df339a7d8a8036d217fed456f2b7420226f496e400bb5b7e0eb840
ze4a9e6e0e396cd15bc768ccdb6ddbb9f994959bb30a461b1afef0b347e95388369dc8752ab5a88
z716d11aaf34a2ba0f48629320d3a28ff6685fbe62553864b6d437f151264d92a0a2367732af96d
z4e84216ae0bdaa067d1a49b19863a31d881bdff34971d65adc9005d6316e524a00e61888b3d9a3
ze4197362d2e9d2d60dd2d6bd8eefd07fdd5576cd0e078aac744b3178502d147a96bb4424839129
z9d49c16e428a2209d778adb720f7611aeeaad575d5fa84d22beb72fa1810f86b0db9e1e0e931e3
ze8269b36604ec53fdee0c7c17fbc611d5988a0e5cc70fe629bcff11d56a99558ebb2898a012833
z7fd766361461c8f54910447c907ad716041ea3a5a8497882dd6375f23153e86e3b388157e0135d
z8da21a7713baa7719c52bee40a009514e2851a09516b63e3daf60c0b1aade3cac31517bd12cc55
ze1d25aa79bddf5409a006655cbba0838903203dd899b7476fff3e436fbcecd99bfd2a2fa45ac89
zd2b4e7036afd7f83bf2e4d756178a859b75654805c92ea74100e6f41ce0c0c9c9223bbb1e0e3fd
z2b28a6ad7cb108d057db77f4a54cdeabd53a6599b88f356bb191e1e51e984ea5189811ca5c0f6e
z8bc995957cbd4737a1678ad20108e2981d4684e2e1eaacd2021d50cedd1a885f594c4de68f2f31
zfed0a370dee56a125530c4d4f9e325760cfc9b46a8fce5e3ba6c5f3ea2f0836431601b919f1bcc
zd37f24a0085a38eed0710fd5e9c2bec9e44de7dd961728c9b3ff2ded18c248c6b2afacafdd0133
z5668ae23bf63d3834ef0ac9d42871587de57e8373395770f78ce2eecb69bd103caa698767f2e27
zbe816aaa30080e9b723b260048d4260de230d2763e34fefee64a2a1b035c0640ca649acdcf157e
z2f7dd275659a92c171c6509fb840a5b217c4665e40c779b4bc5372089afc3ee647eae1837e1cbf
z63d72c3708910435a5d3d02924f6ec063603a5529500283a43cb0fb1c4bcc1686aaae3f44c989b
z0374403e3ef9ebd004c2b50b3d7b5ca040922894d7db86a7b916919538e581ac858d674ec119a0
zc74f6b377c0c5660aaf27a24acbb8a4048ef178b6647263e58e36df8c8c55f1a02e4032ad91e6a
z5b55c157f314764bbe6dbbcb1e559248390f61f554f31200556c5b3046a0a4194687e3f34905c3
zb3711f63a3b765d56d101bf78d018973f31f65bd3785f1fda808a348d36c8c434f28e62d7df62a
z27a7d87aea9dc2b2ae146a786c1bf1cdcce449ee3cb9be5083e3df27d19cedfc4b90952326f0d7
za64aa3522248580d4eb9ec07bd634f217428a952afef104aad12e431adb2df4566a368a7e5827e
z8a5051f0cbe7af51f2bb849aa8445ff0556e58179c3e9cdd931cca799ded3e94bdfc95d8878552
z1df7469feb3c746a23b09256be0552f14aab73c1589fa015e9220e8bfa3d13ea53d6fbf80c8ba2
zbd1c59ea9aac8ccb4750628538b59fbc8dafbac465f2e87eb5532739187c20dc779f3d32e95b31
zb2c098ed3bdad91c404bb4ca8da6649871dff0c24c548879e5d8476fd1ae53518e7380bd718241
zcabf72dcdf20c97073bb73809db26d11af7c4fefec7b3cd43b7549497aeb7d40048217721d9d56
z7a55a9b39cfb876fccec18e0b37bfa657cc260590a6c5f10dbc71ed106467e7454e1ad5c19bf8c
z6cd6162612df305aaacff1b9726a202b18450fd9680cf0ad2e03f258833017eaacf834fb0a3069
z9d3e9363d7ae7a14559560258c08aefe235c457ce662e745f58a8fe581d5f9ec8d1eca7304575c
z7d88be47858203d2ff202b05fe0ea246c59678a9cbd9edf722038e809ff27bfa4b9709b62cfffe
ze7780eb49463f0d5a13df545246d3921791504d656d17de4d83242c633d0299482f27ae854e848
z1e5c33cdfebe3ae4da3f7f56abe7b691a9c9e1bfbee3f1a040e5b9112768b6590e34dca8b2b11a
zc05bff13bba3d9389b5807637143febf7a88e44112ba6720a2e8c83b14485b99c61ca6b3ba537c
zc0b18ea547f1c798148c56cb93d1be0b90c342173770391b059f539e5effe03fea325b7c247206
zf293dd3227262826a7bf9aad90c0bc7de719f50a250bd71193823734c2f76a99840f6efae93fda
za55d073cf223c75b7229d835f845c8e00c517dd1730dbf22e2e2cca1e04eaf64be0abcdaf1a46d
z7b1ed73340006e7fd555cfa2a0c42fe4c49ce6a985caea0c45be8b024e105b7e6a8eebb13e7e98
z234b5e86f55c23f9e1bbd247569f0df50872f226a743b0823c97e4c00ca483afafac81835f326f
z17546e0ef6521293457664a461576fddfd479f7c35cfaf7463ccf583329aec9d2e1ead925fc372
zf217dec3c742111dc6c90856390866f7acc2fb2956b4773476e45494a2e8f056963cbfc4a0c0d7
z5b243886abd920125727221b26f02790ea0b8e6fcd7dd127c9354af87bf0dc4c1204201abd927a
z4357563a42d7646290e22bf7af9a7c7b5c98d319525840aa558055bb975d3331e146a2b0b24cb5
zcaa50a93ada1d362f54797f0b3b32135eb251086fd30aa7962463994b6c1847c880eb9a0e0787e
z3e1224e305ef871ae8d5ed532ee9855061488f214ba048e30e81893fc68c7151c6b5a38d63ff9f
z24a81b72f07f951a3f7209811175d2c8f5d36cf7bd70d996a82a9950746b595df967a1960f9ad3
zc10b575811a8e4abf9576371518be3915911bab835937d9411fcaf27d2d706ef885ccfeda90548
z2e0c4859d20fdcef7137f69471c512ea5c57ecff7f94f62c24b4b06850032ca5c8b5e001953f47
z223f2a39ade7dff0b8a379d2ae4103af8d74d09c8e01a56951d43739d3a62e755e67d2c5894751
ze2f084994a448f1a752a350fc2fe167d29c3145de24adfcba8c84a6990bb2a76e89e2118dbbf14
zb454442754d91e55578b82597a6459e352cee3b52bd9975d423bd966fc033ca75e43c7618a098d
z76fe7403ab62ba225e2053b80647b9a729c6ad7895e52cda06ab8a35e8216d62975994f20d4174
zf31687475ab9e1be26e47255aed3c0cbb01959f91e599090403a3eb068ddeb2569dce36d6554c8
zede38134885a294791ea04cf4f713a86e44a6efa9c5bcd64d9ac31e410bdeee3b41b4834cc9d3c
z1a6617dfd4f68a85ac1fcec9b0fd3fe335f4d76c22553fc754927ee5dc7c3891c740445f1be7a1
z2b85cf5f52ea44f6a9e72f1f5c91321909ef89fb3692d80e30af6feddfc7b7d368c357ed2bc05e
z9f26ea90603d521cfd3cd73bb615678ed3a24de6481c50be88cb7d17fafc65e5c74ac7183dd14e
z123ef43291a20ba1367903883928b96cf3b3e9846b9015d3da90887ba5eb331551f02f302e0541
za982033957d3958581b7943f12248375fd9d0b9b14a18bd15b9873552a0613c9b08f76feaecbc5
z3ccf3f4d10e4dd76275b03113c25ab489321bc1b77ceba300bdd49e3f756fbabe0ac2d4116cd9d
zd3cae20426eae8d23e82aaa5678de988e525bb50c7a12df6cf26c3664b226e95004589cebf8a14
z7c54c7acee8d13b376109cecc90c13b7221660e4fe98cde31e2ee09ff4b83e13bd474468761695
z439e08727180378232ee95a201e38f778118363296c41806fbca98125a5374c58f41a72fcba561
zabdedf1452c0f78ee8c8fba56a220d5804ad4c14bf2528e22f20d8c202cbacc75f40a6709c458d
z84391a1c88a95eb74fbe612e9e221a8d029c1f23af08c1834171361049c3a0838c905246d53f5d
z0eabac12372dd8b54aa612ff530561db24f693b461c5d8ffd74cafc65b1a1f45ab30de82dd92d4
z21bb6babb3c453ab32feff409eeabe37d0b40231f6684fa03ebf76cfcd362aaeb614211236d65f
z47d63fb9d78e1ed9ddb4623506da4ca48ae098a7aae9febaa68de51fe059404079ea27e24ae671
zb45acfa9b4965bbe43ff72255bfb43ad5c7c50bcd1b451eeb61ed5fdadfea5acba1ac5abf85c18
z287f00ef89f65dfc9ab596da229def898f9ed093218992a387796ff1a3b6290c7acce843426e7b
z046a68b28bce2cf7ad816cb7161b8a56199f0e038c401a71624a9fa6da142453416187ccf8fa9f
z2b8a9372f31c66b1075f5e040e0e0b6c26f3b8ceb836776402004261417f5a7cc5d42f3283501c
z1fe69aa43ae880ff625487ca828d7e0ec597549c6671598c6fce2ddb99ecf9264978f5d635f802
zd9aa91c357916768fd91a0c32c52e5d33a7cd893d5ff622f63843c5da11f2a6c5855ef8c19213c
z27d65d2d4c4ab2735fdd3759b50684ba47f2a06b88ba5792398c9efd5fe6b9e2394e8843fde4c1
z66a5496656cb6ef5ae7e4d4252fa2135875ba83f7b99130e675c4653b9f48ea261b082d0acf547
zeb67b04d57953efc263377ccdb018184ab252a08e8ad93b88006dd08cf68146bde9255d8f94d47
zba018ce0034944813ed3683aed698a8bb3573ee9769a54237ec9e7fea6c439d72a878d37a63507
zc8432cb174d32d734aee754b6f1966d91b9a3e83638b8de96aa8ba61a6524583a7cc2f25db883b
z55ea2c698dd972bcfd51f1d57a3fe43dc46d2af0e433ae83520cc362916d19cde05403b304de2c
zc557d1f4e8e3530c57d193fdfad7e3169cda523605797680857b5d6b5de7b4daf0736453d647b6
z9e50bb4429bdf57eff00d44283d5f9620853fac3500286ca3b4a472b2557e0ee3751b18e2a3729
zc7ce91a8a81632f7ce33fe43943a6a82d137e97cbe7e4a446aaf6cae787e0427470a2611eb163a
z6ea705db0d9928ea1a393eec92d7debf5077208f4bd3935318927919bcc202e95401ebf70a1dd1
z841e296fdd058213266455ebb1628a0d83fffa1ad67addda676f7096fcb10b652f2176cb1c8b97
z815727a9e1460624dc5cdc536359eacfdcd4ba037ffcd6cd8034357877c7b869b0c24210ce1d60
za0e24587a6d485276b50d47693a230bb070ba187b2f0a5ee2fc68f606da20efa48539b9ee56851
z98caa89b27c4680549e8b7a38f3d5dfd4587b207175217a801b4ddd0214c6ebfddec9b590db96d
z9f43a47d3f595b457a6d97a4fa2eed55a67fc4ab6ada22cc845b864803b4752b7670ad6053081e
z7e396a3ec065a93cda9cea8fd775db612826eb168bd8b058fef14964223493dbf37176d8b6f802
za26084044ac43c1c42dd4ebe600e65ca7c966da53379da3a024b6479fab3783a0059f3960cabca
z8f9974dabc76cd1549914c2c736bf29acc19c35caefda788cf9e9f134c731e76105cdececf181c
zcd81dffc462139ca534b0bcc0794c1e45d3ecfc069343283e8bbbb4b5221241026bd2291bbaf27
zd4964a49bdf1095e30510d11beb02d60b0d39b22d0f304e4b22f77557b8216ac2b90804bf03822
z630059e2c65f8372fc2f682072ac58a81c9a1b1ac6978caf1640e2d86e3388ca5d7bfe23bcf8ab
z62267b55bb679af167f1799f113ad8cb71680e157e82b23d94d1e7bae4852c899ba2e9a7339d90
z99da21e647e18d598fea4a637bd057243ca09bf7b944f327c236afeca4493bed2a36041b25f3d7
z7a35a8956169ea25789828626972ea003cf3226226705eeabe254aa78b8bb4650a1bb09ef4f902
zd10732561c6465664d28b9deabf265a135de86bf92a532b0ff794adf99042d9c4352600571c2ca
zd715d35615120469f0f836f2541cb18145d5c2c72bd3b1d35d5912c7d7f5da251f81961c2f712f
zd6d92e02cc4bf9986e851c2f814f7390bd20009b61cbc7062776b81c04d9776cbda90cc07385e3
z3ad3742a7ef2abeada1ad775ed179fcf150f19c32765544d475d6a5f6364e1a16f95271baf289a
z05c0028cfb550ad68f6f405c566bf01342b8d01dd11fa3eedfff28ff24ce8e39d83cbe9cdda167
z4563618b02f0d5bb1ffa8dfdd3e6f2bfc23ff91888a51cfe712048589631f7738af1ee2f949460
z67964ea6f545d233b16af99469263123e6d44c6661ab839998377f791eb68b67bbfcc8d9b9e817
z151de46b16d629af8d79d09a1298905fd7b3e21d1be8b5f41e617d87712958e3d67ffee90694e5
zc922702ece9350f8c252f599c89719ad47b37dce82f9af257d1e4f425754e77d2f04060d77d215
z493d6e9048ef5e5176d4a40c47bebc18698ebd238d6fe1860befe0e8cc717883868b0e6b16cc9d
z471a9a6de519fe23ae82154eaab3157f4e28ea57baa5e4db52f859a3a676fb734560872a087ef9
z5f374136ae1d92850ce856195d7412952f7c65864fbdbe2c51db480bd3438909bf979974023d1d
z6befb3db3643435fbd7202d95e52d7bcca5190094289efbcab06a413c335793f1a133f579a316f
ze5474c534f9527e84b29f5eb9b6a370a796071f25b6e7922ba53c26c6869d342bf591257005ed8
z50bd09e562fc94d5e5b33d8d597b44765bdd83b3437295b4d9feb73bfc187a5c77b2200684214e
z2310adf361cf1aaf44e39c7e434914354a08d3e4388f5edc58fcc10f3194e90ece0a46d2e69a6b
zed7df5e890eaf284fcc000f87c4e862eeba3dcc48d6f8094b6673e41a8a9419e08990b504102bb
z1403915e64833e12f157d82b8a28c43148628187f00f304be184e9fee5d8a8ed8f816c149dea4c
zf659ad2a324ecbf4b4dab9f1df3f188dcfae02ef54a3305d88ee9cedf92fc029f186cc04b490ba
z6cdbcebbc48e6226d01b21f637acadfe35f8baf7803c025af82e11189cd1272f9ef0cb7de3df85
z11dd12d9c0345b125665f8cb438ad08d72a07dc70d2bf3372843c761b97f848899e2f43ceda7e2
z253b0dce4c99340bc5dc1379b799c1a3ba1d0be295eab0ae9f4cbeb573364fe6c4b72554210bad
zf8fcaf9071a2452ecd48bbd9eade748129dd7aeb016fbd42dc0d26b36e44e729a4580ba1e31000
z0eeecab1b72cc2fd8ce0fbd48f08c015f9b4cf3807324b0bbb4952c29e2a13257441706b9c466e
zbbeff72b8e005ba0fa4754722a963e8a4597cf0b2a28614b3064076e4631663c5ab5fcf8f5f70e
zcd2d71d38c6f2dc9e57f1afde3d0fa4a38cc006e6d28618c97d41389419a68fb834e0e3fcd8e4e
z31a482c980f36b78464e847e4348f18eee01c852f422c1ef9d2c6bca054846c4292a20f4f0f026
z41c5af216984b7f67075a86a98a756415a5971a4492ae5a4ce39a1f6e3f80653d4555998fbea8f
z038855a76e00fe19f8a72cf2975cc27b9bd93615cc92847afdf4d6ca4598bd98013c5924768bc9
zb7bb4d2ba6b8025c67f662e64d11b84cd9a862421129eb8c903027871b08d5387a7dd4f513fe8d
z714166bc2fc31725ac3a3124c61816fe510d8e93aa7a482bca949d46ac0ad94040d82ebad143af
z0ae273cc2031be3d12a4685bde43eb70f5f5fb96a7c017031e863791924a3674ebdbd22821f4b0
z323dfe0df6d172e071f43a3de519e9dc32ca85911030ee92ae12e1be35f3b895fbb5f2e725bd92
zd2dc3185a71358bc0ef927f8b4c33bb832643d43d4725ae984a28ba5c51fbb54ca51a8e33c285f
z1532acbc1b0a2fb67cff16566aced8808b0d6c5d9ebde0f01ef809390e32383070f399d4061851
zbba75631d343dcb9eaa9c197d20efdaeac987292cebe2233de02579318dd361cd8b7305413ca31
ze3fedb400cca691c805e39ed85b3cd0de0aedfdfef09e2af7ce7582bbd5367e4bffb0d1dd9da60
z8db615265a7bca0df33fbf4ad98a59721d848c29a0fc14a4f4ac1d6c6705fa3e9ca1954293f6ea
z2beeb2be5e8574cf79493cdbd14a454c55f21899d47419f0f7ef7e7ca027d896d82a066f665a5b
z9e0bd1da3fc13ae9df5249637338a0ef9faa5ea28b4ddfa224db61020a4417d728efec5d925e71
z9f937de7e3cdd123b09af266da6c9ef1d708ee732e6e7f9f5f194ca445c9b8f1389724c9e6793e
za0c87f1a4a7f34053623a8daa29ed7b36546ffc884f865d9187986d765404cb90e8a14f2abf3b3
z0fa582b210e6d7809c31db8b6b2eb10af2516c34a343eec42f0f4ef96bc5ded6038424a874a6f6
z924e602647034321711af111a613999f3583a8eeb83ad43b0a9c8b6e65608560abcfba4da424db
za1877910fa55cf59fcf95eec438560ee0f6e9cacd42cba83b2384e505e9d72b145eff534571c23
ze20aeedd97e292cfc11a69b96afa69100eb7e8bbbe329aa074942b732d1cccd3e38175be2e04c3
zc0289b030ddc356af627fcb0c10eda5f13a48a1327af9f0b23264b3f877719c34b377bb2c8c9c5
z2bbe714f187f603e49844350a989e7de8068d0c0aa5071fcf7817bdfd2c20b4b0f83cc52a32450
zaec9a54e1ca84ff000edec8c46fc04631df2eb15d5d0973c625dc2a9b246e75cba0af87d9ae617
z419519d5ba5fd730764fe43dc79c1ebc476430610d41e8cae5334611c025d367b77ca8ed741d7e
z4983829bc590f9302dba54c03f60eee3895f2ba3b358fdc6178adb1de4e94050e302cd6befc9b8
z71d5a9aed959e5457675bb567411bb8178d4d45d18c5e17d2b818f53bdf4b011f1ebd2c9375c8b
z1fd1d0eb792609b12aac876d41f0b6c6f64f6273679f9829e1e66c42d1149e03b092c738289bfa
z89de667ea99194e5d2de4a13fdae26bae9bf80866ac941b39ae65551afb30358160ae7613633e5
zc4353f728da963b52076a5b541e39c70dd714773b7055f5e1485306c0fd3d0d7ce4ebb98c441a0
ze04bde3c6a55e3ea4109224802303825562021fdc1c21957af57db228662e0636c9d86a6671635
z6ad8c80db5959d58ba55d0f244e0ad1ccd408985db54478b2690adbb447f7607eb31db9e199961
z58d3c1b7ae228b8273b22b48f420c84d5ca65678d35d75893ad55d306bcc2bff6547bd0d740f5e
z0e7dbe4b636a2c27810dbafe6e99ad436b8b578375ef2e1355e8689b96aa0517425e855f488dd8
z9ec2dd03448911a5b42842a4c618c315750201aa4b7f887568396cd192ac063c0536be947678eb
zaabb4960b7c7f8cc4d676454a8bac438136ba86cae06adf1191d1943c4458b1de91292a58ace9e
zba55c2182f197a503ca3d3cbaebfa61739e3b86dfa439cf647ce97caf13bc0a88b6af2777af3c5
z55903a3a9a123a5c2f78daa118a44789ac4f66f86ab860396f57fbb460d7089e0f1ac5c8d548ff
z4f9bacf550f2d08ceb1df68f2df45ebeca3e6c6fbda68f86087234ce32ac6167771f46e1ff966f
zd03327422328b507bcb72962410f7a628a96876f86ecbe9ebda61cdad274fc33584e65cfe8c193
z77c767d57fa5e758638f55985dd5742b6f2b07f7147ecd6c020114de2d676115d7f6a88fb886ac
za8a44388cf6aa190267839a2d9d065201882fb3f71897968d1ad3f584f9769e63dd623ef329044
zec573f6edb3d4d3843e86e1b0ce97da583586d9cfd1f7e13686c7e64acb802b718cca3f00a71cb
z3141b54ec5251311b2a0fc87a5b48306287d8f78dc93beabc31d23b7d9a9e7be823fb0bb873f1d
z03936876aa1add580b832bce2a84e52adf56a26a3450f55c7f3c80ec1ff1dc11ea54958bec19da
z43350abb66c0339655e2ec958b05ae64cdd70619f0f83c5c046028948e11bbb7a2b6e2cad22f90
zb357058b3e748a19a3d30f61d7a272fd8a9d3591fef3570eda708aa2a26451199b6726c7b5eff9
z3555bc358ddc834731fa65255eda39735fd46dbc3bccb1cdd33daa3e6ef9e5ed449d1afa5f6822
za120d21b257e2f91f851c20a57cad25adfde10ce5dfd01e0112b653704a86e4e0707e82bc27ad9
z490cdafafc33bd3e63183f71a7da21d70ae048d7984faadf1dcff3f0a936b7f96cf4e9bc85add2
z7ed5ac92fa4e5f948b0a45b88b29aefbec2b1189e252b3120479909d455f45cd3a19a1191798eb
z96d31fa25854c1236aa52ae3237a4bf7dedc01b764876d8c7984a5f314a1ba6eaa64aa1b33daf0
zbb59df7d3f5ef5b5f925aec402d31d4fc03f528fed40b15b57779812af3e8b634ba26e54f2f9b5
z67512abf4d728515af98a29b9f169412eff8cf3fdf2d75317b5acbe9ff16a84e528365ac78c877
z2c68f2cfdd8d95188b88b827a1f602058b9c8df2cc38abbd00d425afdb1b1a50d77218891617da
zddb031846c7440cf70fa6c0a3aa060b330be2d50deaaadd2bced4e48302e2fafa9f682ecbceabf
zb07d3fcaef6bd3441b07b0a2aab1d734e352f8fbfaee5469ed4a6060baf6388994a4f627303856
zd2b910271e20fe13155b30429657ab2741002e35cf941c5052336320d479e978fce2f703c3d35c
zc4d2191ce8be51788df05674c23ebcc43b58865c2f9aef1923e53b916418b5a0966dd6d432b753
z6cd3ab9aff64556d6453fe1b9501fe9d288943b4d41f795ec36d5507422d25e2d51b160a405ec1
zb8ed29ac3cca866d6c75358f98fc88779a28247bf9ac6c871132277646ea11cf63425dcabc2e66
zb8ed8fb52c5693b1b9c8f05df722afa98e38cc1645fc3c993fa189ec433314de41d76306a1cdfa
z1d86b986e0a4b674c10facdd5d8465ed26b2675b6711bc064e9dfea623ad9d0d48196fd4c7a903
zae5d7e5e2d8a49d4c134e237f9b5839656f1e74b2269e364d40078b7ac738c6bbac47b969df1df
z8eb1fd8541c08f1c98939770681bf855d813c401f7779f8f6d38804984324968e82d2dc0633fd9
zce2e40bc05fb55179438ab6963aa221f9bc495fd2d60a0f3add2b5e5dcd8e36e7216a68bd0c28a
ze973b62dd61b849646f16882f1e35012aaec34a9d94508bf367cc85f1d838a4b7a03037ac5eda0
z47fd2f537093a8e743d4a0bb4ba78b7f8222e1b6f217ef5078dacfc5e64c9d187648113605972a
z2c096ed577dfc1bdc7d0df1a58ccf151eff78092e40ccb314a5febd3d6599b6ac08fb791ab7aa2
zbb36cdee67aa85ea57668d56822019a0c647a8f4a4a0c2b78ec2f9a0c9b4f6e5790d4e1ec152c1
za37b7cfa94993c770a821e176c9ebaf5ada0519b01ba2109e0ab8ca4c503b33422f6053602ecb3
z4d1cdf5bbb9dbaa0c54150e480e8eb6bedf62ae7d4322c0c0384e7964e040e43d339c3bbe2bdca
z99e48319260c6ed958264e6c86bf3e6c2a48f6ab6cf8a526051c7285206cbf4c8febbfeea1bf1f
z6c33ef5009ebeea37384f1e8ce80f2bc56156b7774c5236f7ebffb530f3480f3bd2166e43b3e1b
zdac01fa25919a0011ee06126453c84a76cf2c9f93074a7fb0fefb247eab50bbd29eef3877e1cf6
zaee21b8b0f4bea2003247f8b2f2bbbb331553fa3c20be0086bcf364c767ec2b849216faf4266cf
z336850bac2ea2348203d00d0de0e322b1cf8ce56e3514a1095a3d4cd754ba0c88141c23081149d
zdf6d7ee90c1b9bf99bf01d8fc4d156e7e58766e314e42b039d1df8c8a28d63626a40188ba334a4
z20b51b94258f18937cd5fe9959d814d699085193f5f8d269847d8f7767b4513f88a8ea0b49ece7
zd5b2a79284338e8786eb7d12466aec6c7a6eb75254c3db63c3a26c7189d18a9756e362523eb230
zaa4f3f7dcdaf7d7b1814107680b6d7bb0bd86ec15cb7de5f7fcf22d9fbdf297e77e6543971d9aa
z1187db2be0ac06ebc1c221ef3a7b76ab2fa32c08309c758f8232f6f5fecbdbe04b08ce65d03aab
z1ed28c39d2cb18432144eca90a0edf640bd5d5a4e1a800bd524187351a3f165401ce254cac6291
z36d47a82c919e81a6b5bdaa56a9ad5dad0bfcc0b58908193be1cdc8eaeb9a49026815ddf75b083
z12af0f1038add22b3fc06cd98236f4c9667d997d4fe54aed407e11055856cdadcf9aa180fde08d
z17d6b700933b4c72d1150488c1ed6ce16afa9eebc0cfc4f90b26388a39d1e4aa2cbca7d8d705b2
z03024c04baa8f0e2f4820ee5527eff00feb17d6b90fb1d2c03095e22dc5c5ae494817ad391ad5c
z9a90c86e320a6cd37cf31e64d30f7b6e88a34bc89af5c19b43df2bd9a9850ffe035aae4645c6cb
z7579a34a3c32e3b57af368962f3bc8a5aa3bc9b6c588b098f95630d98a6f017a352764fd9458b4
z7c91fc30a8c6a1c9e3ec19d2569735b42394c7d594cc92de48589f5abdc7bdc68bf7096b258fad
zff93f7fc1375477028c3c4acaea1aa78c7aee6ed275911d179eff61dd076da62c9e32b5d83fb84
z91f7d5e64dcbbedd1b05eb504a986c931d455a80d6cb0649bdd5a660f5a54f7e6cf42f19ff5e3d
z5a26301e1b178051b161991a59086395bb4f58dd14df0bc1aa43d26f02323a225767d1c23d6b1b
zd33230090842de8551ef2853ac034c2c55ee16067a5cf5d4da9a029637055c1c7c82f356f5894f
z97a3ba354e5b163d5740adbfa42f379ba0b1bf9d677694f5c00addd324f6e1ecae3b37c5294168
zf95242888cb29c1f4f7212e2996f3e699a4b835eb786896862bab23903b9e41c28ae8eeccec5fc
z190aa927b8a87223535cd631faffbe9e004a4bf0883e5ef52652124346fac93544abd65b608138
zd78b017d342dbc00cee960fd183eab58b91cfbf79d68af3110056133d57de6dae280853eb95c86
z3598dc54e3beb5c52f805a68f39dd3377c6beb96483f6734d7671b949f451ce365892fc7e9e880
zd83c897e628d4e45c350dc5470d79b17de1f8026df067c2edbbded824390f1ef4b8e8657336c3f
zd5dd5a5004600cd4693b79975473ca6549117da4656332a14f38f8a114707436db4d7e3aacac58
zc003b0e6abbed46c46ed23d361f477ae98cc306c05700c8447792f08d34f2e1593a9c7c1e0f4b4
z0e243fd4a2612a444a680ab1673adb3d7295fff83f19763aef3d431824728774ffca59820c27ab
z255aeb7d0d5267c6017cd33d3d27c64e1cb236856f9bdfa0fa3593bfc37ebbed833ba23b338da2
ze79ab7ece2b797fea61b8479ede2a01cc90f9d91cd86878f6a851392fc67af3b8c1debc023c94c
z13043752ae12dbf27f0a12419de80fcca69cf9389d03d150a2ab24f81227861fe42c602ae85ef7
z49a4c8564f5293dbb1ecfe8b04bb8679f4432724fa326691f530957b585579516bea5dec2aba21
z12d377c0f0f3c86b4f09f6391a8b55c2090bd177c0360c8b6664ecaa4fc800bf603de20ceb9735
zefcd7d9a073c247eb3790d33388bed672c6ab3b6dc1cbd9e595f45bd759ce4c887fbf768ba09e0
z336fe4fc143dfed95d3db561846a3ee3613b6c883cbf2d5ec22b150d1144e1539ef0f09d315ead
z9637a442e7c56c9aac83c0f75ac620015778b474ee742f06821d34f4afc2a72bac8ee5fe879c04
zb8f46aea5e9e07f12cab14f6c805221972d65c47d979c45bb2d13241f80937bca055ddb67fc3c5
zdcdcac589533d9419a1858f9a3bed60341978b111914f6d404ce3768764a123898b784237a5072
zf8726f2d0a8b5b7cb5e5b9eca06581317cf1b21db41a23a3014987c3aa859c44f8518cc539e43d
z3aa285e1aa9daa0ab01add641ba8fb57afe015c1008b7c4027d700bed365844fe6c2b336923388
zfb71b16105720251dae369d863255e16c96149a4c02800e046fdda389b62ae09ab298140719926
z11c053eef75ce147e14a443a470bb8d92306593d520b35bc1b9e07c7bbf8aca8098f1ae542aeb8
z2849e319d2eceef07a430fcabefeb949cab7fa28cdfbaf5b05265330a3a836c76adde81d1a7fa2
z285cdc5a9b5dc5f23c1fe63e6754a32e55e578a30857896433e0cca265f61605126a72e40cf80a
z21994672ffe2197fdaf307bd40507dec4423881590923531e5b4e6789dffb9d2f3dd19a0eb54cf
zefaecc56688c0529586348c92c61c61a30059264d1e2965bc79c17b3d12f5f5acafff1f8c42078
z59eeb63f09cdf2f0275b7215b7a7e27db36e942fad454dc1f8a1f83975914b4c904880abdbf944
zab0d52d440b62d3c498d79a81588c4e7a301f47e5ad8e7c3a5c261df3bc0701b7ccee13ca7846d
zc44e72aa008cb627a7bdcac3688994990ca8995641ce48a97095ed0fbd7d64d03162111d91ebb6
z08b61f5e9cacf1425b522e4e83cfb44ddcbc398dcf0cef4077a8a76260db67a16a0096cd11c2aa
za464158b8c8ce5d0bc539717dd73dd234a709eeb38f901d892952346e7f65e19c168e2461179e0
z7085dbe10026f1ba4bede2f0a107fafba6fc6ebf17b71ea529da43c5db807c33dde1145973d237
z48f8776d82ffa7d833b1539cc1dcfffd55bceb2f6c3849218aa5f0ec5e0cb0a90472ae9747c7c9
z88bdebaa576e1ab0cce7149340b0c65962ab4b8e4844799057559c364daa63cdf6ca51dae21d80
z4884a63eb6d60447931faf7ea1769187c9d941b8991b2e9606fd1333cd3633b4f168ff127c0f6f
zdec63a7009ef36d466321dfcf2771d9961ca470f47c33f1f290c75afa93d7a4b653ad28bb1ee69
z713cdffebc56975995a06d43a1e0d60e6a8d672691a625d7a81a310a04c9525e85c8792339ace5
zc995e191d709a85d23ead5cd3eeaa7179d937543619e49c6bd880ba092bd628950a3162609978c
zd6d7df271ba6b23db0b98c641eb5b801ea813082f321fc0a59a6bb08b15d53d4cd6fa2eac48a66
za4b7fa62c023f619ca6466631b90ca91dd335bddce163d497eae312b7d241c14f4473ab44ba37b
z28ce7b69d2c2103c7b80f5ad5e0f404b4ff7fbe954618228045afe8c8659ea3008eb7ab732b29c
zdb11725f7045f079007cf1cffabb23fac5fe7f0db0beb93f66d285bf1701801a43cafea11eb666
ze1f001378b1b31beb5beca00b26374f3374d0087c70c766d89e22a5a116b5e4e55a429bbceac98
z0bcf3831207041c2dc0464a4e6471a2dfa792a98b03f8ae3ea452fc69bab86d98afee82f416de8
z13894490fb683d5db47ec5cd66ccbaaf803096af8809890ff643dc5b9ceb1f72bd5859dade3395
zfc5ea700524eb5cc579b1b02835ad4da2b9e9fb4b5abab7c761633a80d286acb62846db428aa2f
z804a84da551bff6654c18c4eee8aa46121bb6182e9f187f1bb59e7a846897b259d701f58ebea2b
zd4987a36372702f792cf3ebb333b724c9cd0b8d310dd8d06d21c65ad5ac2e87bbd17b293e8ad3d
z9c8e1c0c417857144e161c7583348a91a1cb49b771dc32d501979309ad32eb6cc46f4b28127e0c
z85e2123d8621289ea92fbcda02baafd499c6b3b130505e277b3b7ac80d01111eb0d7eeecc65616
z1e5d530d8d1b62f52b957e5f064d0c0c073ff50597ac7edeb186387113809077ce89e439e80ff2
zb55f2a3de7717d720aacad8c5ffcadb645dcda357903a203763020ed01d2a35d24e8c81086f2c7
zd92bab74f3e6dfc370a6d6bb0f7b17570556063ab3bf5468ceb8be364b382a1aeb57595facf0e2
ze42f1d8dea6b4abacaaa4e1aa096faadde54b3a8c07f71a23ea4c663e9b0861073bd0bc9f37ff6
z7dccc14dd7ca29a3dc9a15c55eaefb50717f5334b45393d21e9f238784aaaaa0f7efe0e584fe2d
ze42def04ff8dadfe62a5d16def880eeee97e9ef741e026d82e8f42a9c01d487543d87bb37c9b86
z66d8d52f34fa08b31763cafe3fe9a15c3b6aec3fc891c0e95f0ae8304940dacf749d4ebee05031
z203e07d8c90d2262d8a899cb8a6bd1dab422e34dc09f3cc5455c698e09131e5ab1db8c17b18cdc
z8580d20490eb30da3c47a1bbdf2b53f31a5864f716921d4684e600aae7c2dcbc153ce2b13ba3bb
zf3ef0f5023b451c8825707605d69a21e726b6ca0a7efec17ca51b96a293371a1d7ae18897ad10f
z5603e5309afecd2f0eb51f2a76d77a03e758ba6553c1e9fb7dd35e63e9131b0915a0eedcafe40d
z3a23a120223a6393ec6b8c7a2a513fc05e3c0ee0790b716a84efef62c60a105b46e904063746f9
z835eeb71268344da54333cb11297f71221082def0cb0d4272f64e418d8a8af26b394a235edffea
z1fde41bb1f79a5150eb2e93a8c0907ab1cae8a4f38b5ae401de5d3e7b6db97c9b0bb026d692517
z2a7918e0062ed1c6d4eecb06b0961c58efc422b69b2b79e2f0f619a1c56d41eb58523db2be8869
z99f69d74aff85f4c8d6ea29515f7798a995ca52aeefe7945f0b72e1cd069d512beb42ffb16c829
zdcc732fa8d41f748832da29ab03544e5931de34fc0dbc53ca62739bc5c44c3a75007fafffd9a09
z3b10372eeb93a22021a345afbb61359ad52202553977fdbb229947935607c208643c63e7538739
z35e81539074db8ddefc395a19af3325e80fe79e3b185da64a4665ebd1cc8a27ac82d2715b97420
z3f67d60c438be74ded7099f555af8d378b630f6e1641104fc1a2cc2d0e1ec187558f78e7616594
zd7fafc533a81a0c05d2388117022dec5deaf9badc37587924b5a3315c3216421760f34aa60da0f
zf1efa390da06dfb9fd633a59c291a972e2f4a5efe236c81250cfaf9cee3ebc8b87f507b48405e9
z229ff35de2953f468431bb19358f4d904e485044877cf35b8b3913a7887450d6e3c14f2718f89c
z3d7b6000e21a6dfd53a8924f13f6efea90e015da2e3ea41d041a94cc772ad9a617fc2e5b2e9cac
z4a763efe1f84540000b605f706c8a86d8e176540e7ba32bab823b5f03ab81ce287c3bff1fc5fe3
z2468b9e11457ae0bfae1b62b3f906b5d4f6e72817e45a4c425bd5165a6ef7064170474746544bf
zf7028a5747943b9dd47d19734445abde7c7674203729fbc0970cc2b7924c44d1ffa83f24116cbf
z06df4b083691d8fafd09dc591885a8d87ba39bed6735899211bec40e267f0b5fc6b6ac7df30ef7
za186332d2b26aaa2323407c5a6939a6d8328987ecfb548098668c8f2adc53fb681124cd889d271
z33aa4e9382c64881ab876fafa0d81b63e0228c28a444c5e759c941ea9365755ba702f29fd7cea0
z176ac8cd5425df7118daf7bf424cc6cf8b608082b97766c0384228f91dfa099b4e3a1e04db1550
z91e7e33e33a30082b99b757039bc5ffd5614257aeffdbc3e3a029a3c4b8517f677c4a0dbed1275
zc9e0ebded8a10383818d57a5d43f92eb82a417d00e419c6f8a1ffa3dbdec1c5a67418453a2814e
zfedf7c08c266b4c3027a8834d80e9a2521397efba052fbe3bc18e84d6ed9e39cbec83a6efd5d91
zf1da73a67b59f261adb726fad99443aeaa75f688c43b4fd00dce3abf01524fbe47856433d67f4f
zb4a81b5405d37379bc3b2a01223b624bf0e71c54fc2dbfbae8a6416083a3577d8b53a510b21fea
zcf75792dc93a9b435085daf00ed567b18624f47c2acd118a5a9d9a4cff347b7d9fa07ef3df2eea
z36329fbd79a6ffbc28d70d18e95bdebef201b7043788c0c57759bee4ffe8851e9118b0f06168b4
zff28add4d9494edac0deb16bf2f3cf218ff22fbd8f909be311a4dc3da9f4dff3c97bfff65d27e0
z0fbb2aa9fd02577cfa87e1d932c4ad2ffaa28f87e91a9c477bd3c25a947c88f0e97998cce8b85d
z70dc0e1546b49399d9b375e7ac063eb3cfe25e8c5c67b884d1c4050921d2a5e23d318dcd3d0338
zba7a4aa0100a8339d6cbe0f947094ea62c71072713c0461e3e890745ecf54e9aba70f099494948
z2b6ea6ef30845f3ece30dc32697b1361aa0a45bdf8214061718d07976f3b329159c2001bb93f91
z5c5b779b6cbe1234e0b24c76b8fe482b62fbf671de6c1b0acb6fb2662b5f445f1af282c5057688
z177982cf269220f6c219fe58069d2753cc3a73c9a19bbb3b4fd9afac1ff3c2a020b570143c8705
z3195c2d36f8753ef43e15c261b0a87e7a6e5e84dfe4b19fbc128393c4db2dadbf6eda020a5de51
z83af3877fc736681d296b7f10c3c7547c620bb9ffa620f7a4d84778143f69e60fc24e337c83d3e
z5667c0fdb339835bc2ed7f6e321424c655f3aa5409bdb20123f3e983a425b4f973e22c4d55f80c
z6c2ca9088b8375fd97dbf0979d8336acaf97c3d2b87cdbfbeb118b386f852c4afb935da9462ce8
z9f068c65a65fac98a3751281b77460ab28515e5fdb212544f5f1264e34620fdfdd3cbe33268bc3
zd6bae713b1c9488cfcaa35f708a2ad58af5314c94b9491ad8e15bf0d9e8289e77c567d70d0932f
z99c42c0ce6e11dddf100c76d99357eef2b1b0991394715ed96b31a6aeb7661613ce38542650d68
zcd33b92da2982f80139e2092b293552492a7b451fa723ea2617c5353fbe7188e6e97d034c5d8a2
zecd718e4c47935e557523cf327f5e6c2a9cf01cdce4294c901a7f51737d32cd307d69d2f3d4584
z3b2ae5f2ac7cdb080cd397ba9df66b250ecf5226d02b1812f4661dc65cfda834172272ef533def
ze51eb551a30d928a8bf757c19b4a33ae1f786cf38aa075977c4e923bf9e8bb8e842291b8dea0b2
z1be88dcaa0275d982dc64761a340ac93dfe411cd1631a434bef4e8336b64ecf24ce6a2ba9272c8
z1f25d3138bfc2439aa669ee72c23a60df9d16991a3f662e7f3e0dd2407ce365d4a47ddd6dd2f93
ze78cf39ef2b0aa61cf172138f8eef3ae78fe635be4186c62031d3775826f0b38375bafed0c0684
z4c4003aef6a1f2d6eaa0d55b063673a451ef5bd0e108308a2c2484079ae681e7eed849913bda79
z6ded498d96d04513389f14d6e881a458985e6c0f04fc9ffa319c4a7f7d465bc5d48db9b6dbcf2c
zc912ee4917da114928be0f53e7d474cc8f7739d1b8a5e580a87d7e89c3a840def230393c8d8b28
z41cfa3d03c833d0f9d44179e92e1491967bf177456e5a3f95cb70323e1342f263606eb885d5e81
z761da1fc2b30a36e4dcc57e9fd8f3ba667e4b66da0d67c574f8d83fc04db93b385d8c60c5e2940
z1ccb7db65818b5dcff782789a5b89f5e33fcdf464796b051a866b485618e921784c9bc5184f2ac
z0a67fbec98d7b384eaeb335b5205fb94e5a0b6dcf9921f6af4bf3a2375f2b9bc32ba1b6c15c92b
z5c927c02aa4d18a909bc54548b1b5b56f932728c78f69ecffb46de12ddf42bfffe70b4cac7b13f
z89a19b7811bf63656802f83da7c4ea35656f639cc4a7ac85eef3c66912bb1eb80a1a383fd60313
z063b146b4a82587162ac2d71ea2664f78cf089b8737ff8d002d7632778ea100a6f2b085985105c
z7df9ca78947722f316c2380903c2dae8200a5b3f0f0be9087ea91e025f24b12e426726fcc35307
z77a84a5be308cfc5219465f9eac3226a12fb3bbcdc28d7972e5c21e8ba098aa59787a51aa55cca
z6e5d58d82ade45f7b9762571acbb1a8965357ded4981fce0c919da6bdcdd57436f44055d6f1b31
ze7b5e1cbf23a1ef4ddf357613ac04aabbd134b235d6db3c98363b1c2dd17d138f134bfb9b16838
z2c7dd86aeb0613db16918cf12614c117ab6e4cb26e479915ceb627a4d1eed80db891c7856b9dc8
zf3c6f8855595f1c74b973eea72388ac788bb1b1c6c008849d3672a654618e106b737e6b6f5c1d5
z47a2d0ad3d5b1ac7719a77d4c225f9e0e570d79c6904220cc1a9f677d812334156b75ef9c1b9ce
z6a74cf0e95492d463c5807f88fb8cdf483671f838a3cf739c43c7860507901059773b2a5249447
zf7812c2bbac8c8199bda8f1193627570cd5acb71c61c8dbb5975cf36a237f2a60b262aaf57c9ce
zbbfafc13962dbcc406c82ab9ac54034587845800d60ef70bca311ae4b4114b0eee58fcb6ab3488
z06be0fd98c9b5f7695260bedbdd31467bbdc6a964e083ebc2602b8aaeb604a6a25789462b64bda
z5b5d12a23be35fbf77c3cf2377e6077536e445ab6f3aaa25b6f55d65ea638251aea700a9213fce
z688b54d51c0c55850b529ebec237bf4ddd01e9d4e5981b6abcb32cf45c3e4aa1020e1140eaa09d
zbe427551d73347d9bb6ec8e32d9a0c06eb43e19e6ed4a550c2126754512a0e411784e30795a17e
zff755a78ce0d5128def19fd6d41a2641157520da043ca3ab78c08568a3ca359746a78498c9a5d6
zfb756927ec366da0f264a46b3545d38b78b6cc1adb113194f4b0bc7d6cb3dd1121e7d885dc2fc2
z358ce290b67762223ac4fb54e741fbfb322baffdd14e3c2e036ead56ec8a390b89447e26dc34b5
z360f1652df472ce7ac1f1364649ab6f8846eef75de3b5fa9389da0e00957d9f135c3a412d7e1c1
z6b9463103c1d6ca7c0d0ec7b2b6b942bb8c5c47407b018ef5fa70a20cfeb870fa6ce3c42416afa
z1e8a06745908430365cafcd7f5fc8a78d1fe5e9068067667521cd7d66da25558046709bd0695b7
z3bad9ace3284fd97fdd7ada0426c241da2ecd17afed72777ca18fe4e1c0eb3596627b0d9ed0b8b
z04fe172402eceacdffa7ad9f422d2023848fea570b16a80fdd767f44b0315457a39606869ee370
zd0969229c6b7574c55bf138aa2bf17ddc77d71c19358100addd3e904ac05be6e4bfb65e58fe354
zc916bad7b2085f1e7e16fc0a2f0801a2641b9c1a44244df43006893acc7fef652e62c5a8ab90c5
z3e90bce77e416c1a3f12d5a7c49edae6dd760cde1a9f43c1186c745c1adff3005057f606b5e92d
z38d5e9ca6f6145e7e0f9e0a34862a94493eab2f22246d49adeede4a5e4d9fc4c2674712aa167ca
z41086d28593fe1dfdb51c0276fe652330020999f236517f8759e3b306cc83327bb7a3a539e41e5
zfb3285f3d5607634afecf2f0bafae8dc992cdb26dbda0950cd7b2d957b813f849bc4852e10a94b
z48e3597e72238ede34ef156c859afa967b64df8796aa6f341b6877ea87e0c9b5274a7c7f385d17
zf40632d52f2e792c259917d13f6e7eeeadecd2b3cbf2a9a77328b50040e0136475ef8a2faaf999
z0dfe43f34f9acb7f25a13e57197601d8a7684ff997636468d8519e0877be12204e87d62158f48c
zc94d66efdebe1f734770afafa5c007e0c8858e4701ad93f39441b74225be4e6718df829d627124
z4c1d6aaccc74c7f84ac5995c8f1a15d139a074b10fd6183c031a26dffad80383a7a10da97a5e39
ze1d4f42482a3f70f2a8d15d990740b9e6e8a1062059df6bf21aa56f1c49242daab07ab8bca348c
zd9e9ee9f700abef6756f791ce5211ca623f79c9750ed6c5a2e3a701d34275f50785255cec45d2b
z67053e8396fcae377a7ee405498f1d108f8fc9e43c06b2ed53232b6cf7b03ad47fccf7b50c5bc0
z902067b717487f48e3a578028f2f72278e2b8e04fff18a05a32a2b37b52a364fa2f69affa4da40
zd63e3a54d7bb4342cee9f67a2db7399d259f208428e5a1afabf2a1f3bc965361c28ed59b359293
zd3061ff3aa04fb22dce3c29e83165d7416144d3680d072e53b5ee88d7757af950a93d219dd21d7
za9e371aa765f507bb9b483571ffcd4f9f7d57468f46ebe7dcbdc20f4804936a74396790bfb9e74
z05fc53689fee7e855733474a811ea283abf21c27f6141aeedca598596a4c3c2acd169096eebf55
z264945df15ab8f06115a7f6bc342c7ebeb4a02d632a90566f733c8d5f2441910fbad0d8fec46f3
zab165b0b6314408f510c54ec82f9849fd6e0a1ffdd350a5a62a5914be20e8573877e8daf5ddcb1
z300c8ba6c4fe59405f321209f699ecc1078b6b9e30dfd993011f6353ee882fc7dc6dc96b51c7fe
z911ef43f29802774f3ce39d41fcdf419c070886ec647579b50af863b598838ed0b9be3c8c0cf67
z5841e9958d1289fe7812320a796660079a54cae51ce28cf6771e76d7d00b2c2b5c7b00f63e034d
z6cc85c5881dee50ee17f610bc59961710e78474b8ef5a00f251cf45a27197fdf3ecc10ea8d493c
z6d58de05f300059e1607e940dbc4a819fb9f28ce793e15cfb09d7ea61d6c193e933c11b466da74
z59a08239c037d8d3682cff8edbb452e947b1b10309c8e71f9762e2027cdb16b397c25061abcd2f
z0517e7a0b23b188a62054fd1692d6250637b925e8e02c9d73335e814b743f0c9cb4166328db0b9
z3c716c6d8a72153ddc574b00dd922af7f927364f1c8689a9ff346290b75d5566ba64b2bb3835d1
z02f69a4a933ddeed9f4017794ab71d01bac6e5feb932609878058205813aae00af5f88c0619953
z7b87ad0568b926d8471961e9ebb173d86ea3f10798ec02c829cb41dffc66b06b81758051d38e95
z68ad2d9163ee220e4e16dcd214584f89036a390749fea4f83f4b5583c8ba2eb392bab5c6392b78
zfb7e087972dc98a128a5b31e29a590bafba06ca85c7c346ce6676768064867b122b04d06878286
zd5153a3d9ba69203813a021909f83adff8f20d59804c7ea471f306bb7822cc8f78549e79f3e33b
zec2be5501b2e5ab32018b2ae3b8108e1bad320e8140d89eaf84c31d5e2fa9f250ea3b460a4db98
z91a16d24c36ef5084e0c0e9f500ac5bc08d94e1f53baa00fbd405813966876aada3e77731fa6d0
z7cb434a00fd81d395ac25660ad3773ca77ab0187c542526d9b0b3bc20bff96863a9ceee0def796
za909e745ff6fa8da7cff37203f092b8bf336b1dc409dda51074072af07e1312a8d8717d6bf6521
zbbb3e4fcee0015c9e708404d90161e32e8e250c9615ab9ab34c1dea82751736f8067364ef0f518
zfd989c7dda9c47122330bba64d3ddfb29226c0d9f65dfed37e10cd6c4fc33071533cc316a4445b
z58efc2460d1ec10136e5d66482eed37b665afad1272125b34f584e8894f569cec072c54b4b7d57
zf4a00165fbc6b8a19e16b9d0f0edab4b923b20fc0d2d8f3d1f49d404fa151572347461217d4e27
z080588b037fd7af5071b9bf3fc909884ed5a678736f0a4f38202b7eef3cb6a8d5c105e3dc4cecc
zceaf80f35e737c396ad0a4e7b226b11dc272a831589efd1b214c5e7de16a72e439f63f598b1313
zf31b9c28baef484ded87e0c15183e2dd543980295b40ce47ff5a681be0e527f2aafc5f28836722
zac2dfe52dec2f91512b9e414377288719cdd2a5478ca4629c6ceb853991541624697b0cceaba91
zca3ee0a81a8cc55b7d9202797b3a0638a749e6283359fb76f1f4b98f1a356840a1dc6b89751d69
z7369d7a91ee17d6ceeb5ce354efe038a0993f6ded98ad4011b406a337fd2254801ba35cab7d798
z41e467330d6f7410f16efee5f862862bf7906f1c969377e9860b2e21d8f229b8774d568f3192e3
z054d884c7cba526988cd36532de59c4223c6d94e648cb3781c9112e731114e0f33bf90a220db79
z18a531c48aee496d6faed7d2179b11b936fb7c726be5ffbe71a57c5f8588c566ae7d045d9fdafd
zace00044a0a08a769ce00544d43c5ecb3f5dd94b658db41e812c088d988e4ce2534069b318917f
zc8db09505bc93d3d766de05791a01c235b684c8a0f0679e7f375a259442f2bace7a147dc30aad3
z0bcdb5a6c7794f2278a231db9305ed52f80537690e11419f209ae4b17e0ed012fffe1f3fe358b8
z368f5a5f036079fa8842b2a5ae64bca3d7f7459b252b77007eb7ef5a17536117be081423bebeab
zfc08b8d669545cb13fffb85a9c4d1c5b1374cf78c6ace9e2df3836d7284ee7d3131b23db2ade57
z0f970646678446234029bc98a8199ebcc17f1eb73c2820053eb76485089d132c21f72c44b7646a
zd9323bcd34df688eba638430fb779660a605c603ce9bb5d25d283ba0be32386a4646a41fef1ac1
zf886a44cad340ce28b083d710a8a18d0921fc363cabdcc0a4f691ccc51bdc40ee9d094a578f132
z659f43b4c8a69b6b032a2b1da93c761d676a66d7ae7a51bd968042c69ce18c6ca44a37b2c0708b
zaf18d8840dbeecb3e88d2d0be7c969699fc5663f8cea27208d1d6bccc1af4cdea601dc5f93e7b2
z7778ca9eede73b5be80bd056d03463bb90ebb0db53d513644507f78afa1e8000c5d290a7e73adf
z54cd3917296f0f451e9f2cc900ac35639fa881686e720539a7cd407a03dea76c7ea2a2f21ab563
za042040021fcc904ba5ae257d06c86c270a88cd3d2fb6d9a434f7959e3a3289deaacbe3f851486
zcaf3b9e62c0551c517381d7e95ad397309d4446ca828bb5ad18ba482a11b02c4bf99c7d42f4ce1
ze090e8950aa38b8a277db8236f3fbfdec901aa0c875b90a51e3f6f7bc9f257ca3f41c49451e507
z31f73a33f92da236a36b3b4d093088a552d298619b0539618a6096b34b11d9e3269ab987aa7b26
z7e4ec699a058baed4afd0e28608d6f87c93aa69fda9e5d2be363c7e7c190b29343575460705828
zb0ee7c6688e0cb53fd67d8377113b5e91524f9c281b86fc04d3da066292799fa525d64b70ec245
z5e0c3e9c456d8e75f6462f54bdd3cf0490960c0556d871d2145466dd661cfe99de20efd151d386
z419e6783ad90f55aaee0e883405934dc703185c3076e0b8253216eb5676a3deb6927dd04c0f670
z591a3118372cb8adbf14905e2720595735f2b9ea41c3ea2e93491ca29483e32bd6b8e24f2b26f9
zdbbbeef09b960a3aa1c80698bd86ce1ac069dacdca0eccfa2eb5420da6ac5b5726d17fd60811d2
z32b269b2d3d07ae58e067686eee1987cccfe7c16293c88365e289361b3103fcd2bcf077ab1c101
z666a1a78e57710cb8e7998f3b537da212a985dfab5bd413f0a2050f1560b2f3f3f37f384371b5f
z386fb70ef189ee5d75d08bdac31a586216fb149d71742df60544e870ec5f75fc5f9b19743d6835
zca52e7a5a7d2e9add423dd86154566e0f28f5bac1711766e56034b922d4d0f796d341b05da0583
zbd621bea5ea306bd74a338246855ef2b053c02f6aef5bf7cb846a56420c9772548151fbb6e348f
z1b6c49f5f582fb369724ae95f15a5325ec129c825ea723a290013f5d6c26c96038a478163d4469
z34f977478e06ff7d43af1fde30cdfa02dcba6b9b3ba91488fdaa97063baf5018417776e0c8d8f9
z6a7358a82081c335d8272a49caf11709fd22cab4bb3d77b9392a85baa4be90f7a4d405e1eb394d
z42f4ed21cb0eb8885c0fccd054d6dfbc899afee82082864a891c6f514b8c4a7946117c37cea937
z0caa43b26fc7f105f6b54cb1ab8a84a917de578e401e71fd8fb7da3ce891ddca336953ac0b1958
zcde5fbfaa950f5ba48a255a07fe90cc203222fd67262177087a4a174fc8f6a4b9234ba15566c4a
zb7eba6cc67fceb3929bf45b605fafff79a2bdc88af65878abbda9fa70b09a36cc8eb4a74ae979c
z2e2a3bd3bd4b5e3b1e583e192d1ebb414b671a6318d09fbd4c5eba434501f8c912353249984d5b
ze57ba7a65f4388db63802ff6af24830c9ab1476cb2a347bdca1256b46d91ecc437fd6eff3201d2
zfd18e259b86dcd39e33d8ae0d28256227511d793d8b380b668f9372ac9c6d791e8148719aeb30b
za6686157b88b362e144c3e91277ee89730b790fbfe6ec11b6aafff490c672e4d594d1ffc963c94
z8fcddff7d475257d959c3c79ce36f48c97eb058408006b1c4f0bd1ddf8008edfbe8904ae519f3e
zbefb1e8325d19f0a22cab941f1973d35a468da3c608992b9a3a996a6cd06b65735e6cce4b05a27
z355aa769ae537bc9a1c1545482ff53553c5bdef752a8db481dd7324d40a27dd36488b5855bed83
z3ac083b25cf653e2fac37f07e6a6bcc4fc83a2a80eb68d9141cebf913a7211f5cbbfa9d055dc7a
z13deb7c6b4cad49d5b440a7e9db3e9553de234fb7b3ee5b83e76cd840f96778596d84c01fc6774
z73061d88665c622256b47577532ed3adab07b627f99f1068d9acc5a49d436d316733dec684323a
z060a8592194f5c5c23a556fb79a65bc3a72e728d67aa32a4b09d3c1ece3364f84c49b7e0899828
z8a6cbe07c920045060038f62ec0f67d4657b00e089d41ef463824c72dd01a1a447b8289401e95e
z25beb610dd1c1d9c5124fbf695e7e144dc9733d6ad506a229110b874ddbc4c7817bd8384696dfc
z44d9cfede09edfd2fd1bb1ef716007347148d2c09f2c4efe9f2fdd333648322285c6dca87705db
z4d783205956aa29b6c2a8e788508aad90ec2dd02995afd3e54c8ced099db34d106832f344d7005
zf92394503cfa993840b0dce34c2febcbcebb87217df0c45a16be5e722f1e3531f5f2d655df5e26
z403784785167918f9a761248a7ace228afdb06dd02f317119b90bf02cb0b0083d5b7b763e45e44
zadaf66b3df2394f4072ef359c7895ee16e40a83dc49469bbe6d89cc24dae134a78106a04a4d987
zd28ae1c957c811aad39ee359878de0db96c0cab0581cc252202dca65cd9de2a756cb3f963300ca
zdc75959eebc97bee982214075f68d921c08389ebcb90d39c7ccb0a0e5ca79ae3ba83d431752a0b
zf67f472267a974ee6c4e573635266b831ae6bfd4990c88e8c8d6c6389fc614c1e4ddd52133d84a
z45173989cb8d9e1e02316d027e3d830474b1d5551c5bcef9cd61be17bd7cd31b09293a97d59722
z7c21c1fb67bf25deaa2d2713dd1c5ab56fd124c6067cab020d19122fd952cd10de3f92adf9f220
z05859d7c3bfdf1497aedb84893b99bd3020acb6466429337eb95e1020e982222e667f4ace301d8
za0cabb7d911e551ae03cfa124d62dc0d18de47405c28226a6442b0371ab47b708752a4038cf144
z159fc64af585a8af9568bb62ce16d239b66bc163febf4aa9cdc66301afb732a07ceeef9ac8ad92
zfdf96457a627e22eeb2bfe5ac48ae585bdfa853bcf09ca10a5117e0db0285814e5af58ba5af687
z7867a61b4c157e9515eccfb5655f95773bd71a855e7994a21c73088c6836720f986d1f039744f2
z438fb3042af0ec229325fec0ca582eccd9dd7caabd07cfa9d4c8019d230b5d0f9c6299373cef13
z266d83cd32052974cc4073961c2342b1e7e1149874aa60549753c859aaeb9c6bc8c9313e61ed6c
z8bb1c65adfb0b9eea6901cb9c3b86a11a4314b28057e31ec689bffec9d342f3c640163d1f2d62e
z58b24235ede8f50c33d1032344e45d3ae3ee872ac25ddd3860173678f9c2a0d951b47f4c064c13
z08c70165821a72b8c5a1ffa6b874a5aadcb2540c395f04da6caddb1cd9566ffa73ee82c835ff19
zbb7f1cc7c10df8184a1ad5410a4853202106e122769f9745649f5d5f246cc696be3e0215193f38
z7441288564850849d38f2fd9b152c22fac60a17087c959b2b09271545548e5bdc4232c175e1e38
za52633edabccdbf07fcbc2e082ab65dd56cc984f9a8bc0104f4d25b958324863e5b3002eb3e513
z6473e983894299e1b8aef779ce24277f62169d905eee99509bbc3ded53c1a2aa6a84bea72bbdb3
z93784f55e0215fbc7f9480e4d71593b72997b958d4a8457877e7e85454086e9f3712c3bf273ec8
z95a51238b2d58312940ad2f3cd62bb246e3543a97864d02a3ac09b25a177fa40e8678184e885fc
za8b8b34f45bc27dc426d2994e7d1153eab141eed89d3798161c8e38f46347abaa4e8762c7d3d81
zf4a5f6eeca5988ea3e3334692283c4d8d32132b90b157db761c5c33b1d41a9a8e48f5103892d26
z21715186a9736702db05ba9d2ee586a82f7e75433d5edbea8fe938769d903577f3623d77bbd110
z8fa97d54c7f0ed2173b47c59b5385bfff3b982be19d0d20985e0ecf7978ac70b5c97375fa28ef0
zb7b8ee5fcf29b475299ba9909b8ceb650c0286932f633024b10e9b620e18f6eb3fa815f2f0fb1b
z962d9b6cdd3456b5843796995d0fb07669662bcd9ff865dfc14b9b8650626cb2a81bde93f89117
ze604d6823ae9a71ee14dd41127e2fd60fed24bbee5fbe9fcbab0043bc35d803bdafa71eb66bed4
z6e67533d7bf53b45531191515e526db634be8bcdd672d86cfbf7ab092d4a8a2cc2e807168aa1ef
zb8cbf255cc63860e64fa7be10f2101a674099fd7183affb19a2c3c964677e2608c25e9353e983c
z225e9ea47f5a3799704b0e2085f91e507512c7fe33486ca6202e606a985b327bc21e4f71109fc5
z0e50ad9ef49930def9ef3ae8a2a9fbf707f7ee5ceb78bad31447bf58378a6c98f9bf0cc1de0b38
z62a687d925e665e3aa00d116d65532cd84fddaa5d5b037b77f0fbc18dd97a82725646189615d4a
z685807130e3d01508968657f18ec8e151f1a1b9e00d0b8abbbaf388113a84d470aa1b28dd70ef3
z9d603dc7721d7eb36cfc28e4a75733f58025a2016625b4d718c9533d0bdb6374aa3bbbaefb99e5
ze56bbbdfccde0f21a58a2b85e0ad7aecf7f9f05ae465aeb82fd72b47f37cde79110956194fec1b
zc42ad5ba4d3128cc3ad16d0c90916fa16dbe3a4883c7acf47db352ae0676d50bda10c5f13f5574
zb91269f62843517ea496e253c7a19572e522a092739735d6ec186423c02c17fe89ef1b8bfc1021
zb372317974ec0adb5d2bd96da91d41fa68b7bd55e55e441413ecab41a695c24581ad754131ca5e
z098304c9102f918893fe6ed6227b65f2e02cd7b9578a750b6aafc1b5c7902054d5090c766194fc
z37a19e2eda10a978d08f45c9c56206b78c7b10fcb61825f261beef2261cfc62d4afc63a056a644
zcc6e3ab7774f5d31bf0a83d4cbc172e18cfef837f1ea9b4ff99327e9b1a067a5add670aa1b5d73
zfad65f2359110e6168280f609d38d902c892466f94c6c5d2550d31e7c79f6b8bfdfb478d955f21
z87559e866eb162687cf250c5d09ba4d2997f5558dec9cbbb0186211bc21dddbe9d63673a3073cf
z839f656df40008c51b4f3ca4e48fded5a38d1a73937f6ce70765cedb3e0efe346d0cdf96f9876e
z1be9de83eacccc59fa82c91c1f447d8d925c769db40da802983d08a43054ecb2da42d52244653e
z151523e254f66a25b78c3e0f0a6a02b44862f2f5b50ec413c0007700441054077feceb3d5510fc
z96ae537f0515334c3e29c0afd46550fd0394e4a4620caff2ac5192414511e08691cc40e60fe7df
z385222dcccb95b54571f56c4dc17e58bbf5000c0c787678a42db1ca4f0ccd7cefb715e67713221
z255b6f81d1e6b8067ecc8faafbb6bba9971e313a5f53868b0f68e830441f3c73d609f392d244d2
zdf9133821aa0bf61fec4a107c255eff64de128670fa6d02196a2b9460f6afad876facce2ba67fa
zeb57052e464d4a028f6cae52cc086747172e41001758789e01a80b5817945a7fd11f2acd27e17a
z971c4734e0047110cb583e5b9af96bf32d7c5ae9469a2e9c4e3708dff720fc8a480256a1885e86
z64a515aa41239fd490f6268a9ff95c356cc75645abbfa913f45ab4cc652429b3099d4f96e9f14a
z7547ccff1932c34872a70b8eca485b9db36d1b64fbc6311242caa5333c605367f694c82917a29f
z7c77a7a39851c111442bd9d374f292ce3bc15705e2a0ba42dabdc734935e7f7e71bd2d16d75c1b
z59372877d4a588a75cc9b8f411ef09b043ba4ecf2737a36b5ca71f6ec9919de7109b9b0c105ad4
zbee90f706c26dbfa87ecd435efad9de90696423046188094d5913e7fefe66927ad854fb6a4917e
z1524b5b9bdf4b3fb810d429a0100d05becf582857ae762111c0feec6662419876d1aa7c0335fc7
z85ecc779b926ea27a46bb92a90bfe68ac254915ab3e5b4203c74999f54a7a88fd0d537fe8a9212
za75507941ab4e2dbbda10a794c9003c0e0542de5ae12ac5a00c6ecbef2fe2a16ae2428dbbc81cd
ze2d4a50777a0968d5d3474d5a9f661ec48d9760c41c2d3e7afe8dba24f360323f0ce3c2f962440
z0a724332d9d6c569536dbd2357aeff660e688a90dc84302746f711ed2614f24d534ca25bc8542c
z89f9c83c464fa34763433c9f51f910e431c26a0ffd214577537e196f6b674bfb90ac558428ab0a
zad677457dc868a9fa6ad4dc7149f118d4ee60b65958fd7c22f50ece978484d954179e0bf3e311a
zd29097c37e914898599b7e9d3b38dcde53196539780e0d88c3e664f71be2dfff60b41b96178c58
z0a7bba70c8d8bb7330f11967ecc71a1c5835c9bdd8867eaf1c5215ab6e480f38efcfdd62b6cb43
z3e203ffbe12bbe75352af38f8ffb1fcca47a3868ed0e27a2fa475131a4383dead91a32f3411065
z28adbd2c2e1639816b2214eb09fcd2fae2e2a5f41d7284d1e165594e67a0fe562d59fbc38c0488
z7ee1ed2e149d06c230577d70e51798340e25074d4278f3e0fb39a3d6b2005abd8425b9dda3aeba
zbcbbce25daa8c747eba0380d8085f474527d25a62a31befe7aabaa71fdede8e5243719d735e410
zfbfb944f7aed3d9c9432c574022a7949fd2398455e756e7cbeb0eb469b06fb2a773aaf3bea5175
z2abe878c279f4d7777f758ccc4ebca398338464f36d7bb724a5c7b2883bd10c37d71e8483ad0dc
z7f9a120d7a1cb3cc9b98236610142bf6a34c4d2dd2e5d13da1509c61190eb11d7e6f4d55bacf8e
zffd1ee5d6ce7047f5aeaed4b715d2dbabd3c515beb97f75f6e9a91174a699b4b32c0688d170ec6
zbe930d9884f5e578fb35d8f708f902cd9788489f9dd372f559995de62d3cb780f198a8d381b062
zd2cfbe484d4f1385c00cb58bde26a5ce509d3d3fcb62feec6cd2bc9a8d6815d5b002b5ed12e8cc
zc1a83d49b1d3e4202702c054a5b3d8262b13c1fdff7606e7785602284d82adb63bf6721f441f2a
zeb605ced0509f6b45e57b52f34af44312d596e30a10efd02a22ede7357c50e842234c3c90e2e0c
z9c747bc1f2a185a58655bb5fb885062dfd15ab11e50f6e5c793765b3ba6a9096cdcf9701452406
zf3d4a3d2e8cc80e21f462eb161e62373c01327390d063fea68dc0f85a01e8af3742b940676c95c
zc143cd0a9bde230594590d6d91ba2261f7f93cf6678da3a77271e8b17f7a0cc094476ec36ea3de
za9345460a1385dc8f402643c63aea80350361c8d76457c39558055b254a2fe3cc9c6a9d957bc4c
zafecbaec58e69970f4916965edeab4ff2fcd45e471f658f3e71ddca9901115c2b8205341edab96
zb41566496d0b89a068edfb52da5baff5c492e5df0746df122e6ace364e565ddf679f1a2452ffbf
zacfd8c0e57d3564d8b6793565473c8d236e84138bba4f52d36ca5211e056dac5009fbb806b817a
z70524f0ed051646b7ad2d2dcf98a53cd7a161a50395fa0f20d942a0b52d2dd1a2b6809c477d777
z5bf27c0f354091934cc1cb95de339510e5c3868c670a8f0735a097195a9e05f1bb21940118091a
za20c02a4257d4e977f01cba00da7fec5c81310acc9f7f5f5c5f45deca15600008ad4e8628b4d8c
z85a8823c1d25f40b30d2a826fe0c10fff9915c309471570555b2299421c5ac67f4e3b9e0a05432
zadfd3b7f5c435758541a9edf837a1b8572477f5ee3d74bc5be7b6042bc9e345e21c6bf03781929
z828b8a12e03a4a1166243a623336415c44538ffb7f25b60a32a85fdc3e0ce9a7334b7c79b29176
z4c406251a66b06d4e40a1e1b4922634997b0f2a65fac5795ea22b4f7a184fa864b49d37b83d0f2
z8936d2fa2e5c9ab69f47c390b39683573e5c84d1277109e11ad27e3dc5c6016e4c4c4245fffbb9
z5cf5eb7b118b39b3bc6ad5e56f1de17a68c71cddd5108ac01cb4d01a2370af1f944600515879b7
z43f9e602ae3618bed1c81b010e21628990501184637e51e13debbc93a7fcd693f35969cca26a10
z9455f6dd68a4ee60be8ee39cccbacf8937020bff1850b8cd7ed00d072ac6c2a3bc816b75d8f699
z8117d03fb4b3f6870b429d8c494efa76add0861f7926fd91633d65343ae419ebfad2f52d324552
z8b80d196dbd804b5c4488eadede49cf11f27e8e6d438c50f57f4603cc93dd2c7a42057c99a2900
z959cabc435ebffa91980087139c7264721987b580ef20ead9435b414ac69c87ca6686cfa4b749d
z6e803bacdbfb83c04ce811b45c6192d1e64bc6698b09f094490c47e6ef1bea991bace7c1986162
z3bc4404d34d950012e2c9e4a4510b067e4ac00c2246067a5a51a8403af5f843cc063039e8bb05d
za69fdbf60c680ce9156b31189cfa988fd8ecc6d974d3583704a7d37e9083d16aab10f69fffe302
z265a1ca2344d949a761394443c52546371eacd71df1a0b82cfe7001d27aa4143b6d3c4ae5d8eca
z9428bdf210d3cf2b7c64abbecd1e7d24816bae6af9dd2ab62bc9bbf334d793bca7eaddbd8b00ed
z61f363d5cd82db04f947d9d7adeae19a080d50ef48d619020b6c0828074beb8e6b60e8881d2044
zd9542ca7e8156700fed3a518b9ed32344668a23c244b0920ad8774c078de9525bb9f930b96705e
z4c63ee78f419fbf10f570c1a115e9a343331ed824d3cf7296c426c498524c479e682c6cf79f9f5
z7c024b07f63a19e312dbd96edc18a79d4183e61ce3041054c70bc0db8a8e281c25499788da94c4
z17433ae58048cc29f7a0d35f2b79a59171991a18dd15278d6edca900d15a226961c660232d24a6
z7be80bbf7ea4d6e9ea91815e357546dae648e5d2510d6edb74e4cad77d7d81c11373ca6ee6f59c
z58167e85b44d465c9c3795250cf1973656b8f0f205cecad737a1a40d85e5fa7afd959834e19fdf
z8bd22e1a73eb0bfa77e0904fd7853d03bd46ef1fcb95c32a84c2c0a7096bfe13a2cadccf21f1b4
zc54a480a750e44a61fc74642d2b55919e7fbbb2dbc45098f439cc3b408430d8374869778142ac8
z24b063b8ed918c71dc9c8073238200744f7e4f6b642bd094e88a61a7f5acfb3549365234c5aae8
zf90d5a0cea66132b44fccd77ceb9797d5f8c6e90b809701ca3c2a1606f1aaac4277903cb6bc545
zff7f8563b1b22f066749c509fd35d8572c762379ea6482b2740cb58c3cffbcc1f551439c742426
z503b1a9897d6383b8b382005df0483fa08ef5a0b41f9843714bf4735d852d97fde52d15a2ff34b
z8488f92e7e249c5f2bc97c5efabba267c3b87f1b8b0657795eb2558a1816380b4b1960d168b572
z175195028f419ba427b071c6375fe7a4693e3b542e26e6e1ab9d6f21d2aaa1abf2c5a403891d1b
zb977f33ad5ae454323e1ec4c5ea8ad110ba35d9e44782e8e2862c361234b1f46b5ebd102178451
z030bb8b84a6d2b3041c289055d30ec080117f759ff80242b61ace1fd8a3ecf5ba7fd38b7ab7be4
zdfd12f7cdd29c6cee0c9b24c48541865a187e72f5d32490cce204658105e0b1ca6144a32ca3577
z49b82e56cc33e002adf0d1e7c6394a622e061e0f1ae1199b17679843e554d3b8bee6209fba339a
zd85fe706c0b0399777769c3655aadafca8af9c23a67cddfc828f42a713da8ee90573b9898508d7
zae4319e8a052e9404012969aace95349f6c6c142f89f843b05934e04238b3926160a7973020895
z2b6bd32af71eebaa7c4592e5154faed94edb0e8c6c732484fd2d310a4c35881534de48c9e58fac
z88b3c1a57792281f0127ae09b94d35945fe4e3d793cab3ab4478961ca1ceb54dd540010f74bdbc
zbb2542ccdd675e053c0182604f3b30afbab75f83a9af46f9538296ec5045fcbeb595dd78c78303
zaf4bc36e7998401f0f0ecab081670e3934609bf7a76744bf06ddf124cc94cc4b8a543ff1a037d3
z13689b4ec7ee52e01484bf36c3eea817cde6e11489b6ce5ec3d30c450d96dd8ef60d2d719e3232
z0baa4fcd2dbd96b0c864cd4eca4c6651feb018e0f8207482a470b8e3d08236be5890e9b5b581de
z29ae746ed800dfbb0b531a30ee28fd0d1d915a6fb496339a96825aeb5f0b7e2beef06210a3e986
z3ad481986cd2c918d926e09fce9eb20aa14e5d86f3166df6a39d49aac665cc6611b8cda63d91f9
z9b71558fec2a2e1226fbd2d7cefa454c017fb470d9407993a54b800c48512f6a85c9fc7db51adb
z50a4a7e6d9f51e3774dd84ee58e68f3f6cff29be534a3e49c03090232bb858480ac98c8606c00c
z0b4ee0e4aa07ca89476487148e5e79c9d1eb2b5a054509c46032a4f15d32b8bdbf511dc643d4f6
z9c98c50fc06ef48dbe3ef063cef2b40aa499bd3a1186f116b766c785712fa84f5c5b77749fb0dc
zbea0df171b7975ecd1c5dd4fb44026c240ccf84d0f5e016029ab0317442ece16ccb8f13d3154cd
z2d928eaa28f3f5f4fd29377d6b7e02341ae56760851af72f83a186ca4539c8f56ef7cd125ee146
z13d0af285a173c5ae3809c1781aff7962f1bb7d0ad1fe23f5fb4f32eaa77168a2dfcb02f7c65d9
z76918c7141b8f30274bd18ea960228d364721c2521b92a213dfb1b8ef5d07a7d0412116b0c1a83
za6cd22be04393188345d1fd3b92bb34a4701a7b08f99b438158d6142e6d664135b0bcd185dcd17
zc2465376fba12b92062add926fc5c1f4292fc6c9fe76af3b1c748e9e18ac8e40f9964b5d007e97
z85506c19e4206c3f08ee07ec5c05fa46aefe26d659344d096c7a1fd8c18d60716f79915d6c26c7
z6cabbb73fccff50b98008e9661fa47b935eaaaf1f65d19ccfb4ebcfda801b5de49c284b8c5d533
zaf29ff4d0f11bc01e58fa446d1d88abf6b97ac1b6364323a366bde242d85695f61e3972bf3bef1
z2fdb16ae0475c82098eaca20cf10fbf97ae75164adf92419c1234ddb111a3c373361eed7a031f0
zc2895c63acaf574e46eb883067da3b95b1758a7f95626e0f01a6af1eb2a2216eec7a7e74eb7c13
zf740f252851ac02a9d1d2592d3cdaf187db445bc3caeb6a58ea9f38c6dc639b339a75ceea3abc0
z612fa3aa9f9f810ec023144e0512ee986e7e8cf10c522b7650a7e3e299fe5c0b2fe989b5b47f6e
zfe71e345eb9a365dd88f329acff13d8a928134b9af1630917a322864f7ca2c337e070dc29433fa
z78ffe947d4c5beab0e54af796361774e8c12007f7a0358d7e2b652db5ceff17b77105671e95fa3
zdbb53f4278b401ee65f61ec5db1b4de9f4092b1c3d7f81845d2f09144593e380414d2d47ab3e20
z3ecb15bb67780b287011f53a6c79977a7b0702dfd539202c10701ea4a99054b78a43ff29a34684
z02954445a82ffe8ad4e46e097dd75ff01b0e30283da5219465ea8ed238d8993d74ef396460abb3
z23560c9e11d4bb7a65e77104dafa214a394e120160ef156f47af8d5c8cc8b874ff0ece1ea069af
z6ba1c9a0ab63d9eba0e49e35d6a7a46ac41825b07440a58e796a032ce54c791c0953ad0c3cde0e
z3ccf2f0add4d4f7ad44c5645f6922dfb6b71239a964f776c33a601c39a98284dd154ba9248337a
zb46034bacbc86ef7be884df2d779b600ab50ef3a19d1b08503e4e2106ef81d0b494691055f9612
zb53d61d54816abe112813701573d63a4be0d9a05cc3b3dd3ee8c4c555460774e53e3f93d5b0a67
z1e1b8d7c9cf3760f4e6ffd164fff240f62be84442d5c4810fcaa557e73cf91be37d9540a2f685f
z41d013d3aac1cd2dbe93a548d4b648f1d54ce11b82097cb3972bf91631712db97cb010a350d0e2
z64209d98568bdea0f9bcf460d3ed7e556807f64b15e4b9a1095d7f26f0fac01bc79221846b0e59
z825850b2d2c419239ecfd88af30b2e4aa7c38c28b7e51668fbbd87a9bf8582a92890abeb312308
z2c56275cc68349034302d5206e50c8a40663ec9888423c6db182f1fbc726fcfd2172d3484acbe1
z1e3af9443cc4ae2a674648097c6ac622dbe759bc438548731503ae9e6389e0cd11373760b39948
z06b4cb715585d9a8b8f495221259aab7da584014edfba7dd98051e7c08a6a158ef2741eb68f4e6
za02d3c09f40f265a8964e21b1580d3ba60646e83ea8e4ecb11303639cd3b0f0440194260fb46b0
z101498fbb81f3c688cf22401b15769bea8056212b2468471a235065a34aff964e8a81ebed46821
zb1ab3db19826052476dfe88bbd87d321a25a67b17b37c7b95bafc35a4fc97bc1f053ae26adef15
za07937dbd7bd9fec3de23f4230466f3d2173820ec5f25c36c6264efdcea67870d18cc6f3a79354
z90102f41357e3e4ca9d61fd5ca2380cf0925a8b511c001aea5a76384520eee6fc6b61cbefcba06
z756f3351ba75b6ec85e4dcb3c0e5c7fb6e22c522e5e59749229ce0316f7f0cc50e6611250c102e
z3d8598a941d480b1f2a0ed719fcccb7870ba60aa7fa2a17e9ba11ed509d9751ea4a1605f7b6a8b
z13aca538b31abd32f2fbb3601e72a000766c8303f978a2294398bf23ce422ff2e21474070c852e
zf1eb1359df11a55c9a8b5e6f8f9a5edb2807d856b8cf93a19d8733b68c1e3e96c8b6eb60ab581f
z0803df0486a0aa8afb631889e593c77c78cdd3caff06896d72350d28b79595b02ecaa10758af81
z5c666a70646098df8620fa4c39a388af242865f0dc33108b152835e92e900993e9f1bc303849e9
z1779ee97e9e1c7a3ec83970cbc7a800f9657c833a5417bc362bf53a2313d154c76f0003b27e96e
zebba16c25bb535445eb7bd13f475e4fd3831b6d7ee3b2b6ba95b0b0d396982b00889af4e5df1e7
z6a1dbd2b8149ddebabb1945222d0ed21473d97197449556211e7c8916056041454ccfd8472eb7a
zc06f805297627672c35ecf28a0a9f764aea6ea363e1bf70264cd36a068d5ddb77f608f1c721349
zcd49b6ac2d0f404b6f4deb8529103a467cd71ae25138137c3bbb4064238838997aee3b0e09dc55
z3eb0c123db19a56707ed1c9ac5fe074fd3b3d55652ceedb879dbf4cd9471e45d75e23bb5c8fa26
ze130e0f6e2e703f200086cad776104584ad2f33ed376316a0f28ecf5e77ed1d81416693f9c93e4
zc5a4e03803ba15aa9a4694c206676d0d9263262ae97d251d1d1ddb2a671c6df91f836b6f072213
z76083b00f7d516cc4a78210b6648d98fe9056a3c7e807d33638cf43976acdd531c5677a77f42d4
zd6aac7af8b9003fa87848254a0981b1412b0fc9a0b1f8be941e1e30556eed5e1485016b6454915
z5ed152267cce1fca24f48308d9985723bb3222464b5dd8f381414fa420201917e1ec4d7bd26216
z138dc4458c7b9c227fc6445c578de6ff77338b6f63d187dcd5769506e833ba429a9f8ae3431ecc
z473b2e301a497ff27a1e2a2b5e70175e247a7ba28c0fa8e43d6e08bfee14457a85d0a7733421dc
zff7b46f131abca9225e08fae554534cebffd6c4d3b1267f9755cc975345633179022c9c909d401
z12f017f94cfd17e0c98c5c627e373fbd632c72caba492b0bafd101a9ca0c6e840ffeed3943c597
zebec628c2b08fa3ce0aa7e28a1f5898ae7eae9f08897f9841a1c5e47da3e678884c4bdd503a009
zd710c845c7758e18bba3dc3500ff7beda72026d4ad9134406f9f04bbe74f2a113b176f45815439
z3b1e511ae2789546d993611c504192a08cba6182107162a4b29e39fadaabac063d3adf2c6b2c0c
z3bc7dc4d8c197c3edef86bec4b89205414ff4733c1e0a3d2de8da3f48f04ae44d02e28c2e12efb
z144ad13e190bc66a64c51047bd77a7440652554a4e628353463f61b9f02a28691c178d3bec0cca
zdb3608a1d0cbab8bcdc088f90d2506bb204cf252950cb721c38b4d97cc1511b0c15ae1e13b79c5
ze9a377ce0e6cb06fbf7cfc5861cb6e4c3593acee9e035d7585564134ff0bf9e8da3f51c5725d11
zfe400e1aa1a8d907b4431cc33ed8f8a0ab2653dda09286ecf7d779bb81a95e68c1e7d32abeb393
z33d06c2ba9c0dada2e73c2548e6d6f4941b1fe3b9bc049dcc466ab64b8da76f514a10756002461
z733a21ee2bbf5ecacd8c38d6e142b6813f3d2037740464f7915e0c4de8ffce3bac71d955a667c6
z27e88e3341b079f1f7b422d394c8a1b25cd6e7426da74ddda4ba4784feee4980db2e34ffeafaa5
z148905024ae9dd335d6c37d635ba0b21efc3d43224f60a1f83ca353e6130929dda12ad7dfb66d7
z777d2b03b444834b0876b9fbcdc164a2431c6f6397bffb3e98e41dbe5cff321a463c63abb70f2a
zbaadd202370638be74341e543456f9ada0a84f4b4cbe83172875bde3dd168c514aa5162ab08d8e
z78ddbe3e5c19b0eeeefb36e2ad75f7b3ff4c67188b4459cced8ebb493f0c677d8b7d8c4c05cc63
za69773ffddfeeae279e2013b660729c28d867139b759091de8e83b85fde23c1b1e39f1545b4906
z6237296c6f7d53950d84b0fa155bf01609156db9b59254a3e3c6251f75c1ddbeaf4d7de41ed998
z450e68f9e2ed5e37cd7f945e62c31a792b30051613615786f3696236ba87bae962560afc2b34d8
zb799692b8b65702a11b0f2d441a0e26a221b559a6877bd1790dcb586f5e3cda333b5ba36e80545
zd6f48ccec5e8f76db6455eea014a56c015dbdb45301790f9f188ef5f8f4e48c8f6945522bc86e8
z712f2eeb3724a24125fea956d6db5b74d4810214f00dad9a8a67fab45988eb730dfc579f19e921
zf33842d9c18fdb22f55b6ddde345c40a6999fe8050429ebbc6640ed01e02a055ad3bf6b08615c3
z216ff1c0d80593d8602d25c3e603c23a50602ea54aaff146b4d39d2aacaa0babeab6697f339cbd
zd460d835e9f74497b4c5a3597c9d8c2cea558e64af5776deaf6d7d87549aba127337d9a2f2445b
zbac320f3805d331b5187e4a2e31a238dca58e3f0b77139ea0e6834c53b6e5222ef7329326d7727
z0baee8c966c0c2d15c8318be1666a17b548f27394100386634cfa7b4958cf846b9476fffe7f78d
zda4f51c7a808094fd4fa94d33f2873d3c9c9a1eb5ee3e326c58ed00630bebd734a274f27bd2cf6
z0ecfc472076bb793cac214ffaa3a5f68e5aa2bdba376faeb33904b679ee7c6c500cb3e53d87067
zeb7967d18b994f105036e7611255c1780e7e82c92433b8da355f943d7ea93b1e667d6373c1de59
z9dd0b8449f2052eac365e23feaa890c560c0e309a73bc569d73bd226810d24774a93d605967526
z440c44101ee711b6d10fe42f6387e7aa69248decd3d8efa60f9450f48232d4dcc533027f2d9098
zeb3c0573cf1ac4e4db35b0d8c4456b88425ce6b8cf7d4f2dc9d496f284519d84fd604b947c59a7
z90fa32b1c6317db48b12fb93010321db2a67a31bf9f23ab6cec35cb7e8edfbe7ef297b40d8170c
zb606453f965431b14274cdb2d25e6c7df178a732f0fa7a65f1d423f91057eb08d311fefa75e38e
z20a595eadd08f1096459eaada39d3e547c69e973e4528bb0ea58364a1efca1ab4aa26e5bee547b
z7f3ef57d9fcfdc9b013c5a4a3d51190b02ec814a46b3c78dd5363d08cf57aa952ec31757672d9d
zf8493aa9eeb7fd98189c36ad625aa06396ce85d7944b34695b9dbcb5bccf04931efafdd10f1d5f
za6a1bc8230ad10bc90469cb4fd127d6202a23023d3832f37ef3f03f01771b910c0763a7ab4ae06
z5f9e55820dbf75a656c639d5022459beaf083a7745b1c458bb0baa9e4f9f9b5a5c6aad90818c66
z83c504717d78cfb502eebd8d0ffea765d70cca1fa4d090445245ee1c63669575106098d41d689c
z991b2d3b369660f0e0f76209939655094f06dc047f67a009d8aefc5182366527ba512257c82435
zfbce0fcc7acbd459992574b0234c3ece7a228e4acd3dd5c60d61a05ce3e53fc7309047855bafb6
ze9f35374e56954d4b5168b10a56a119edf4bd73e4d9602bfb6fca2b036b385bc99d616eed9e3c1
zf25f6523162d06fe82f49355a67a8b6e61dd921b3d6053a7dc7f4a7765f6d5fea6f90cb03148bb
zc95d8de1dd7978b0ca6f031223752d65d8aa1a2d0ecdc2e6fb1e9a736307fc5c41db24401715da
z14b93b12b78267728972a90e7b4c7c71071d75e0b8d18f98b246df83223c7e6eeab80b7b697902
z34088418896d4d7ccdc9ffecb6618ee7d8616f695df682d3e265769e8921dadec619420a0ef73c
zcb6df7f612ff9bc2cb9c4a04e3d572342dbe635baa24dd161b42af8174a8ae81c99165ec9b47e2
z9a4fe3369cea9e78a062fb32e45053cccc78fbe950bfa4ec1e1f7af5d37ab4bdfe1056577e38c9
zf6a4a60839d7a674e3a8cda7089159a4cbedbd7b35c911088410e12ab3a981980d09f08ec5a77d
z52f936b90fd24f12404de6138928bc896e04e6ed78eac5fa66ae2d182448be2c07233d24d960d2
z80439b688ed6b6de897a7eda3653eff8725731060cbad6cd4d69232ab396802d78efe944a69928
zf5b707c3546b761f5a8adcdf144b968c95096466feaf053866fff8b1de277778bef6f9320109a1
z69cf56a7c843d67068a4c8996ddc57daf78d83389ef25b9c363a36acd56c143aab8d0c7a8149b5
z0c9673e98f168063ba6c0e468608f046b793e66bd8a3d75f62311c5b33f489caa69d130b23a5e7
zdf9b468c7443625b3dfeb519b8e495dd1d3d132a12256645916a94dd8fd44b954f8d5ace886e54
z870443e4a7097b1656a7c63c2dded4f11809af6dd6db9f5757d11a1d4eb0f94c8e649a79018e32
zfaedcd5360eb35002fa2d46778e77082c3994ac502ef82297e677287f6cd5b6b6da2d6f6f51bfb
za94b3801469760cec15a151345fa5293f0ba022f17c52d7bf6752bb017bc1d8dac6c23fad69359
z2c744056196fdeb43f5089ae6c394723a723327ce2800c67c5dabb706b10f60a118219a268e034
z50b20c6e86f570e4c176ee43c72e7c3882a4fd65e558d1834f26fe72591855fd03f0ee62e3c8af
zb42970a63f9c7df4b5d6b641e63cce3946d8925c3e190251bd44159e5dee1ea43acc7c51d1b141
z449f7564dec573dbbf4ca3e4a68cc354401eb6d518e303d947f9b259a74c5262e641279393d751
z8b30addfb04047e349cc2d4843123d25480a8bb471875c5a43ad717bce5254825c07d03cfc6490
zf976462dae46ac81c1a15f1321158bc0b1ed173c0a24300396530fbc1547b6b4f5f144486c035c
z6c9c7c25a05b2ddd110b3e2c984a444c7199e0907b1e44ce47d08a979ef8b82ff9f52d8df86bd5
z888c2ac86801647ef2bcc55de61f1d1f4c5e31dd1e19988e12ba8dd3246a20f47831d3efadba54
zeb797b854edbb8e744ef848e6769dde0c6f33eef3f2890c787b1fe295386b26c925cd54e2158f6
zd07084f72f7959adfd34f1bf0de1e9d31cb0bcc7d61c38b235e8dbd40ee6e3370bd533ed9b0e77
z4189ac37a6b24bba2c21614807841d4ab6792480d5d713d2716bf946611c9e9fced60847e963ff
za09e20ff9fb67eaff7e35b0011ad5fdc462cffc43108e0dcd0ca389211966967bb7d7e70ca909d
zf7511f2fd839d4ed2a8e2ed6e36a07f0cafc25b9ecc2773f5a165b0bbcae8b3d46a44b6ad7c03a
z11249524dffcf88a6929f572fa8765813b58f46c7b962fd0fb3a46a0e6796d23d1731a4ab2f8c7
zb17b28fce0346e8510d94d069662232c30ef692ca9c841bccb068b12c93202bee3505e4274f337
z953e86ab01e8671efaf7557a56faf826b89b4a44efd26491d3d2fc08e8cc2a08026be82e5674a5
za7727501829a1113e5de8b16aa76b2850450dac247a039ae7135c484c9e4f9078781a13419244f
z177d89ee9c5e523aed768672af905b0d77793fd131c19b6a4beb01148dab6aabfbbbf71646e37f
z246e49880d60c54cc1e3a0820fcdb337e602fc826b5cc7aa2b1f30d4fd7fc6998eaad15eb70a9c
z291c4d9201343c2daeba119b08b55bba3cd72cba7739cf87022a507bfe0984949c65cc92dc89f9
zb2475c730de6461e2a2b1362731f9384d11f511aa13ffa020156bedd4a41b30773bb3450b022da
z704fe14c70acb9e5f64482876b29847a10b8f407bdd8269a1775cbbf4a25f2656e2a4da5ec8231
z89df74271b306bf037a2a4142005e87616d2c6009ea13cd1bdddbea53aeaf9d2d7c50e04f67da6
z836cb46160d3a5830655bb8d4ca9be585412b15f5fe51d10981a89898d6d758e4bdd631e825104
z1fceafdf21146cfb92811515afa50bb540f4f897082e10f40048ce12ce093167c658268463582e
zb04a51df789ccb1b34ddd64bd2def964fd99938f0d3e6da992c3ec21999091be54469cf09611cd
z516b3ac84cd8fc2bfc50007bc179bd5f4932f6108777c61b3e4caaf87e49474c48449a107b8b8f
z453a520b75bffbcb326552f5f2d11ad7b826a3969e0f1d6bfc0bf137b2e56e752126bd81fa9179
z886fc2c94d6a707894f75e0ca1d17ed39b5944dcf88bc5437806a97cb7b97da803ad625d70d815
ze072ede33641f8de1ebdf859b2c04cb56470cf5423ccf71a9f4e767d554a0cc3c1b82720d468ce
z78fd95504c66f210c9c27a6e993d3b9126a0982f6eee01f92d59b3a855cffefb8ccc121739a14c
z33331c829fa34d800802d41c24fe24cd976857783204eaff08ce161f63af127acc239d514a82b0
z3b5144494814b3a579c29b284453b44d4be8925542f89e94193d92c58c2af1a3d07c106ed33591
zfd1f7bc541fd45382083ec6e7500a8a794de2ecf553a638dce33cbdee441b1d1148c087f319f2a
zdefc7133e20695252abc798c72e0bfd714e55a8aaf9e84eee8ffa3ef31e3624e12be5d715ff671
zc8922d93297f35c025a36140892db0f637af05022fec275093974fdad6f3a4645c35fb0f44116f
z39e515afcd10279d2eefa481ae0ed441d6b514b7f5e457c55bdaecaaaf2f4248e4969958e6bfd4
z351fc49bc5e7cd6e59db82d4fffbae202d5fbf9fc14504ac38f26bee844824221f932fa5579be5
z79f08424c4647d33245489d74093c16de7e11f9c02f3b3e789e64de3e344779c6a8f15f267e38b
z367f70cbedc19d5fa5d374195659cbb2539cd2bd1739a801d3320dec6a89b5d311861dc2b81e10
zf39ac7477a95417e281473be1c9a487b6cdbd4187a7cff9df1c53139173820238883558f759f99
z0a2b141ccdddfd9afd015dc0bbabe65a83d85e4c9bee28f31496561e14145cab4f144402dd0b00
z08006e3a08ed5b0c22ecbca342ad2609f2e4392c966c7356ccec436a4d7c6c9cf56a9a8f239aa6
z0cd47f9583b011f4300bd896763734ca04ecf28fbd138fe71cff5cf6d0e3ffce7fb0799aa31f9d
z25e94d42638bda7f19480065f0aca47dd876511d46e20ab2e16c6242bc3373179cab5af21ea872
z547aabbb1d58e9affb5901e2ea63ebda70f887471e615f0f9c00dfbcd38d65e1d46e008574b8c4
zc055f4432cea3a34d4022cbc5dc080b610fa451736698e5e910c5784cd49479c4115d27e1869c5
z2ce88cfe64ce595b1c4c923961664c7193b3fde0771d9087cb8a917e6f6eeb3477e2dd5216089c
zbec756aa9d3b1d148f11db0bbe6ae0188789c0ecb603601fb85b842deb4bcb979e608c43c1f886
zafbe4ec40f97d06c28c904e86107289c00060213246d02958d292cc77e3c4f8ea0fa2db269d34a
zab1f427dd19736691539009b71916de517edccd51a161d628fff5a0aeebdf84197ccf90f4d3abb
zf0edc9a15c9c66059c73582afcb9451815ec5e766800a2958b69f12b1308c7a02ba86f86268044
z0cdab3eda5e7edb01325f1ca324314e9159ff52a4e3967077f079f03cf4b122e6847b7e34370a1
z07ef30d6745f62b1eebf9bc39da444be7a30891f8f7be8c3d19b14f8047198a8eb755883257ddc
zc797efebc3a1c0af3ca492013fe7a16732a9d4647d1068c2650a5695e7f445af3021b0a9764b26
z01cd61a6a253eb86c6ce6155b0a4c2d133545b586eb43864d55191859d79a0a09e9de4a5ec425a
z2d72406ce5af24716ecc319549d434fb62b40e66fb776b8ba784183d4f00e075cd2b7fc1b6a875
z095c1813526368f0dcc8318571cd679c92a40578e84dd047b2b14f214067b75b9b48857a49e1b1
zf10fcada8d85773f59bc312b80c190575b34c4d8d10e7c330bfb1c2304947ea4528e07911f01ef
z2c57dcc74d75c5c75c3732b6f8c34ef91fffdb93b8e09bde0dd9ff391d67cf4ee688b40aa0afa4
za9c491f1d904abccea1e68497b7104f01c79c27845096bc458bce86922befc4c056a7379ef1aee
z931c4589d2831957ebc0d970e2dbfb61c97e938bbb22d311f84d343fa4a18dbdb8e27c3a968b4a
z4ce982faf7ee640d0c9548363c2945a7ffb5cdbc1366939e8fadb1bad7c6db95015f3205b732fa
z26a476fb2ab87c584f9cd586e9e93bbd87bf55307fb531e8b5175082f44cee6ebf81c66f79b6d4
z6f45d5f28da1378ba9207936d51818846ebb80342b01212e07d12689394cf6a3cbcae2b1c22f2e
zad42a8987af6ea4413ec984a6ff362973fc9a0adcef8aec5727e9f90996c46be6941edfa31deb2
ze45c3636ffad04c5ff90e7dbc8335d944caf72f1d1c8dabb1117c35abe4ce4d79a07287dbb01c5
z0a15d25122a2ec8bdf9f933ea563dbb8455033aa0b7796863f7ba7d81129e003ba84b88739b28b
z9309b3d3c400d4e5346782771ff82654fe7bedab5002054d88fd7b9568896694438d5f068b1f89
za58c93959e65ea8244935e7b8022cf989781db62e3fef495b887023768fb652b586f8498682783
z265baef3c9bae23c42ab6ffc93d9fc2f9fe4f34cf65e078cbfc0ec57d9b0affaf0631a97aad728
zc565f9582a756309c7b09bb8358f5ac74ecc16d35bbdd846df4be5d38ae9318f5fb137dade9580
z4ca83e9f83e939534d906037cbbeef2e8c8c6833192bbaaef7214d7330917313a322cee29365eb
z9acc822b084e0c679c7d894fbaadb9c08d89f79a8165cdccdccfb8ad5438edd875a8f991ebef93
zb1ef26b717b93547ca2d91e401d8512811911fcb1dbd8039cae89d896aa127c48ccfa8bbb3b312
zbee1cb0d22f5bf607d7fe911ed2c1c16732b0dd677f040081da5a81eaaa9ef75e62324eecd2c1d
z30ea6f0b97d1d586241e45b6e013823430cd8d42dd7b4fad7a50be31a036ea7e2ed56f456e63a9
z9af0193971b014f0acc067df8c61f34806b9e9c259b2d6385d90740e91d15c69e2c4ae8476ad6e
z95c89c6a0b2dd909b77ebc41e48c65681b27c96410936d91c7b1e14c6c77a31e1151636815c327
zdc3b67f8b247e21e964cbc4db447aa218972eef355105acaaec11b81ac276cf66fe84cd77df05e
zaab0237ae1f0ba7b9c050f9852bb6c214ff46b90a10b38c5c2b6ff0943927726231372cf44b3ed
zca43cb7a50c1533bd3d104ec88803ff34ed26222d7d3602f876c5470a2c46b0d6c6b9c02154562
z069acd60c2febd442f4a20b684a9b64c06387171a9a5e2da8e83ed27a2ca8167a03bd02108c70a
z48101785df9cae19c28ce436d47864f485d3e29043347bb7d341d3b61f1af020e6fd195680e0b9
z001ee8e740fe4b2006758d41fe8cd5b4f0c6b45c743b4a67d2d950689a0d76dfe2f19c412a5a75
z21a5e61de8034a13860dc304121c16195bdc2828f370bb3f84ca591a4ff47a76011df5a74b6c9c
zcf487b2b3c6cb816ef1e354951efc07005c8c26809bd95eb392250be53b94cc14e059dca13d15a
z59cdbde069891f324b39b904fdb91dbaf5213821a664fbe9af16ff317767d46375784c3d5f4aa2
z90ea380d580ba75fa7cb9371817e7ebb0a271e12095de5665bea12d41fd743c28c228a2eefe4b6
z82b53ad93c85415c410b5c2429c8197d9d4c402441f71fb6b9544178dd7923e1e8a31acaffb666
z455b7337b55b741ede04c9562632345a85b65bd9927b699d3d5a7d8f4394b4c01e4834aee6fc4c
zba26386133c85472d4bd3f1bf10c67574a88430aa307488952fd50f80030c7892f3cbf0efee052
z62a5ee07e988208a5dcf9e088b1b9a30c7d50403af4a1e8dd76970f5051d63f04d271fac9c7183
zba7fbd71f68f42f6743c29149ec4e6eee578e5de3e67a7f62ba28c472206a28adf1f9955198d64
z0947145a1be5a1ae3743997311d17836df280562c425249bb852029a05ee12b48d08473af1cf51
z359e801dc51d4406e112b4d5e7847d504e366f72a353d2b551b52a196a5a412d7da2f277ed3c5e
z44a303894f067e9ea2b409f32ff5aec1adacc70a0ad0a87160eaa84dbf636b191d7aee334d88fc
zf2886ddf78641644aa26d3b55196d4f9053590bac92630b6fb8d72edab94ca921083d1809c714f
zdbd62234ee0666975a7279e07d58c0703e839ca58c95fba792d83cc1994af1825c2c755f017ef3
z01cb1bf17f85b999dbd77b8f7a39bffc566754d4a6ee7ac3381045ea5c2f082553da4fe55ef5fe
z535dc61e6241195b14395a78afa639e5876ad11c7691197ffdcf21947650f2cbeaf87c883bc9d2
z2a733532ce770d81e7adaff73bb67c408793e1db8b75dc026b2f118c1e5d6f9e3f102a5833ae6c
zebe3510073c83521b0aba573bbb7a9671f1881e0a007a1c6f3b8e3a18a5126a0b49847088fde39
z3d7cbbf10a6a3bfcd5b6b3a0b547c9e1354a407288e17dc1f14b3ef194e6a5a6f6a8e029f2103a
z13f7be22a04428d54e5f2ad9de45b70a913a44fa1ea6d81125f7d6d4180bc2dba1d7982491ee1b
z4ef135973de7a387037fb20ed8be8cc1c4e11a6cc029e8618aa4066d0ab422372b491ecd6a7735
zbc3d5992f346fdfb4f1804128b28d7a8fe6edfb3576184263fd9716321bd6616e72bff6802f948
zb04c02ecb4bedaa3a85fc313fd0b9d1dee43170abd851a7169f8eb650fdb266f2dfbb9f6c9034e
zecc946d595e0d803e649d0fc10815fc4514f7836648b7807af3031939f8867b58c64f5c32adf87
z64426e88a44df6973d81f83e26d70c601fae516c0e9358feb2566daaf69da0b993b819d79b5170
zf4237344b5b54c4a4e089c51d3605bfdea919e1e785c48a3dc66601d9d04244487d20d8e049a55
z31895796b5d93542a6b39b59b529e365af62c916426385cf96bab787fa947ff289e0efb38fd07a
z771b18bb781314fe6ffa04e614dc7480b76086290558b361e16ee479d1def84f6d611cdbdb0378
za4e051c55d3f60b9716963fab8470ceb07eb1fc46afc81910205312059638d40c2e30d1e50d67f
z8b9af83e8c25a56bfd791bdf91bb864d9f4ca2b59cbbc777ea603347cc548809775343b514e327
z74fbe9db3ad66efa5962e483fe4c500a7583530e771fe5d87d58209bbb29b8f030603995f9fcd6
z1d71d54ca470a4fc3ba031b100bf8a77db92b8ee9dea2e18e0532badc88125019e6f6b2e5a7cfa
z136e116757edbe24d089d40cca3568f370f362f409a45eaa112bed53db0ed039754d2cf03e9d07
za47ace52d3c4ba7bdd842af8361457d4768a2f2ebdc285e3a2dfc4b8de30f50508b51d1acb562f
z1f004adc714619fdf78c2100f71f8366e031eb2548c0b3d1f86d6348259e54072248a0cf3c3fde
zde7393670376fa9b291a4737f46ae4a5195987b0aabda808fccb3af8962573737791ad7568e044
z908a4877f8379a9b3f8a7fb02c52321eaa94213f1187075be8317af167018310af9c6cb9c40163
z1b6297726c6839a92d261e2254c1ba00e857519f359dc11174bd6603fe32a0f94ed50b1f8136d9
za7d2044e20b454bb43976eab56194896177d43008455165f0465ef68397e64009d2863cb6aa69c
z120fe03f4b57c1d5f32baf092ad477f8215768f33757f908eff84881a0ec872d2575d0da725d48
z3966bdde8158f5cb3ee4428181b7dbc58b9cf00854930fa8c6d17740f26f679ba080d20d386361
z0a0e1a95f6c0ae778ee159e61008b5be84463f734fb9b55978b6be726b517e140827729b12319a
z9d4fb5ef5b7c1479583bdb44c873a00790d4ad303f15f33f86919fc7588de07f95555a983ddb0e
zf2ca02a588beaa6bc0f4bb1adb0da8a2e7538d14344b8a52355d5280fa147e3f08273ea45ab549
z8f3dca5b99798300753148a8a87049337a17a5e9acc2fb53b903bb1825375339d387373645afcc
za7fe318f6023958114caae0e4661824253140e44bdca41fc1bd1f101a87a7a4e413dcd94acf683
zc43aa0c1109186b50db8bea62d80b75ee7730182426a80116c9dfc0cd9f181f4811d6c39372e0b
z817a1572fb6572c8cf9c90a8945f6cba926ff3753f1ec3f37293e7aa332bca2278f2da3722e7ec
zad099e4a2cecafa9ac015246b3e85970bb8c9bcda177051001628edeeae37b7d8c3d9b8fc6a986
z3dde5115ce3979aff05595024977d310cc3708e32852c943c6030317dd7f6bd28b1050aa26e595
zd0bb5f8d311add6d5e0ba30f388e2839849924a2abca970b6c791a5802f76d6f3f3d1e8c2ad252
zf0a665ccbbca47c9dd0728088fd0b37d80b1b1c99685470278d0ac25ade3b66595545a285241ef
z95a959086caf04ad6af5964d1b2ffc7b96ed3bbd68c63e55f643133f3e85eef26c9c6a31ebb9cd
z8dbeca65f3d5a992e808c4db9c0fa29c9b966d6941ac6354cd41be0038c38cb8fb25a8f4edc8bb
z880d043a585d43ae95a381e4ff8abbbf47da2bf3ce60f7ae9d0b5f9f8224dd991f039e7f327268
z579fd737e217535a635e7fec297ec55f4d576bf3444c4334d597923239a601cae0d3257d01c43d
zc7878e93f3c8ca9ec0365f2a4424dd9c2ffc67e74b9a1dc9e170ff5f189ada6a2265b4aa9c3aa7
z9962582760d94932de5a2dfb680466203ea51d66898e161a498023de73b4353a9aca37f7ed9b5a
zc48bcfce085f2af54a4578cc2025c0b24258272aabab983cafe7a958aa4f033ee212c1c67e27c7
zdd24ac6f3c07ebda3d65c96f68060621e1a90c1b4621596c04417768a2cff1edb11f8594ee05ca
z67b34161479ec5d62a0c7ff5cf4af1ab64b8f5b991d0d36c950d05d26ae0b4d40920571bcb718c
z787fc301f2c27260f5809a48157f706fd1b2a14416c501b572cad48597f723e44d02a2655a40d9
z194ddc458bc2cb35772caa39b897b6f1bdfc192c397cd269a6ca24045053f99ebb594b17ec1ec0
zea1a595cd32b3beee21a8b8d8ce996a9e47832bae9b2c1594b3e5f8c413a08c9a69fb07dd05fc0
z1a035f892f4e5d9761544844cbd4aa6bff86a87100b1e2f821d4124c423ba2cdb4c19229905a2c
z3fc44612de56d4bea631c5f6d071e22dba44cf493a8ad0f1dc6360efa7b774d2abebf4cef16330
z5ab24938c85001792bd27faaf5b6d75205d040f276d333fbcbbf1bdc0b6b148e4f0d5ead004e26
zecb20a320bed81fcbf4f359c0526962e57b392cc12c026890e30f2e83b62931268c419046e8224
ze8d341e8d1e1c6a632ae60724eac947a8158c8824d3a7e5d15a4f494f6ae09cbb54a6f5f9c7c87
z4ebeed5080ed23744dabc716b9d731f5f6132e7d7c2d0caa758ae0d095ddad731154a31143c66a
z391e06ba4cac9a22ef3571875db77b8297006ecfd9126b781c1f24dcf1374ed819406854ddffb3
z686defba1402b7d649970d2abb4799df8cbb7d6aff2f8c8aa114a4063afb72458393d68003b40e
zafae966824ddf31b5811875d54d490f86a2abfd21ee4a7e72a14b34a4d6a796e33474333395b01
zd34ddea5c50ed4677ddbfee3a8bdd3d87af3e3071089efc934cfbc7ac7e09245c7b9dbc914fa5d
z6a68062feeaa598cea619b4f19c6c68652d61a881421452a4fba293c0e22e5dbe99141c9b18f02
zbe143d57f5d2c4d8ede85613380bed7938902ebe70415cd512b5c789351f4b5198e5d8c858901c
z63629ae4eb1936305e360f777d5e82bf1b4cda70cc6f034127f878447f6bc24c2d0c387f8da592
z032a1a94622a4db4253bc17ba553ab6e9949940f6806aacb4b9fa0c4faef39d9292a36bd5793b2
z7e5a2149bc2684bff9cbb01c58f57bcf79d7bbe8e3368152d95be76d97b05a673643801ab0351d
zb0b32b12fe448fc207822a704aa52ac10e92cab8eccebf2de13b80ceae16df041e701abf1ef43c
zbb8ad1504ab0e9bada5356caba6fe570bd97e82e69ea31d94cfabc80a2d1f666504eddb52bc3e2
zd108a8c83a785ea3f2b2baa60b45eada43d73d9dcffbad163969409dc3cac2db9b8e2a2047ab7d
z059afe7a392f3705d7643c9ffc9eb6caec58b162ee639a6e345c38e78a33608c2b3b5d7305fe36
z785ed3ca8485c05dbd0288659523875c671cb91d161f1ed5a01fe8560e53014ef52ba86d543707
z6e60b8e6ea268a55f109ab114c8dbe2f83bd5efdf06bad3f207f92920afdfad6c119d1c3de1fc9
zd67f4e362da22c38c164aace50883e7a3b1d5d1212078fb9697f934ab6386b60aefb9d8eb8eeee
zc6ee8c6f5d1f1a6ce6013f7d40d1183901a20b0e99157d239d34494b919677ddf8b28d623fe880
z07c1edc9c6ced05e282199c94f3fabacea0ae1d2963ff22494b4a8f57117a075ec87b446bc630e
z90fd836f622e3f214ce09ea048b034a907cc1f4fca228779774d7b9bf3a774224a40515093c47e
z4177a14beca956321d4fe92f57d6c51a17b010788f99de0453e907a7d38b66ad2c550cffffd0dd
ze74b0ab1296b4b7ea4468c1f260d6e3749d5195ca4dee32fb42963c3752856df1ca82fc3569c8e
z453319ea2aa34e0706d25df2a07be27e25881f1283de769ca9c32d0e9176f88cedb089daf63d75
zd615f95c6e3a38281de9b89c53a474cbec60a6bebdba0042e1e5215a820cd76caaa04f28bfd4ba
z702e34d707d961aedfc477ea666c7075d6a982bc3b42073defcaf7196ec83772a925b24a2d9409
z9b9a3441e4d93652f4210bdbab10c04e7ccbdb74adb7e837edaccb98ea446693fb81eb39ee066d
z30de037d08c75db795eb330b85d86dd47bd58dc214209e593b9d706eea76f0d4a564d786d424a3
z17ff03f0781a80685e505028739c27e98ec68393c9562f6eb9d73c328dfa6e200823158da18c37
z5ead3d3f4c5047f6b5fd86228a6aca5dcd91c35a0d0d94f9342ff30e4de98d50cd2aca34fb2962
zb00449f65add67d0187b35749bc8adfb5ae85a59243ce04010b245e33ae54cd7f67848e9fb0df7
z705cb3fb58cf45c15c3de2f8241dbbaa282ede19193152b3938f4bb7a526e384e5896cd317f46e
z08527375e14ccb7a9511089683f1e268384e3771ca76d85f0d7f571b0c8d9af5b07953bea19375
zfc01f4efb63acf995e9d57fa167bfb302b64c514ab8e2a1bdbd804e6850d7c4d4c38de001a0e8f
z829111cadd0177a1064c219ad0ebc475ef8990e5036a46d1655d48e3f103f9634f51cafafc1806
z2088d370a7daa543acbfde99892f5a1841a94737bd68aece9c225f840e6f7855976e57e9c962c5
z0894b07aa29cd95c139da96ec2cf6ae27de872f34771b07bffc7eb2295d25a71b9dfeedb84c231
zec0e8a6b1c8e49f3b8523a812aaefa7b3ad886d4013da880070bf151707b0019169933b6c71f21
zb26fefb8feb3bc4754a0a088e9514778fdb469a56b8d5fbeab50a163de30d2cdb3615dc4045efe
zd14a03ded052c9432888b0dd4c82656ee6e52e59956237e64454e0609ae2c7f57bedd03f6fbb02
z42e592e1ff9637b24f0f0158f9629b5bfd3b9637fd44d684d2f73ad981eee913eeb02b275ce2e8
zdc4a3e6e4a0541c8650b805fe2147935b3b6c2ba6cc0c78d4a5157c2311bf2259d5e4048aa0798
z64d09a5c92875fb5218fdfd70f4d0ab81c8f30ec4264eaaf831b8e67653561f23dec58624cd559
z34029105b393913b62b27bce29f3289f7fc80e2f217a50f90a1c09e6773b2ee00ec5800937f190
z5d666d340128410836f7927a80e4c602b8b58dbfba22cd6c75ddca8f1aecb72bc477077fc2b8aa
z7638c2adff290e6c80bd38c104c2662447c4479f3627f84975fdebce1ad304739f5ac8e2d20285
z6f6a68c7c5682631959a84a6d8e58decaf94984cd1cfefac1722ff9c2c928f9e0c68bd7d3b0310
z7a180c3d2902b8c1fa47529b8113b69459f88753e630bf19af971a53e2bcf6f485db54ebc6f49b
z84f7450704d0e49f5bc907b6933645350ccbc7d76c90dd3aff370e6dc32a424e44496df4c29c5e
z8182f0fb4639752d01359c9c17b258a0f1ed425a089de4dfe5401a73f954edce617b53c8e04163
z4fffcd769be54d60319839813a9f9c0871dbbcbfd1605120aa9435a66ec86cc4a990b144c6023c
z5abaf36347a2605402b84763801eaf701cf4a82393f366d6f7610b055a10438251e9acd8198bae
z6cc69d1ce2c41a1e5fe92d627ae87ed28cac74d0e07e4892d02e0a36ea2fd1f8a3eae0e54c5605
zbdb50f0ce2fa0ae586e0ef4d1148537d2a610bbff03560ebb4fce7e2df93bf932bc90bae3a30f0
z3cc4d133e3d36cfe56fa857b3c271a10d0f0fd1df185f092ff1d031db0a42b9279d2aff89b0e7c
zf4952a72d8079d894e4f8b6d308dc812dabebc208bbb9666a08f48bf8132b780f14dd8507f8bf1
z797d95e0c77547a8fe0e56d8aad3321c1f7b665961a4e61dfc6023c866e5f76145d12feb9944fe
z08b78933e670ac5ae59cb4d050f700ec2fd64e93df239e6350d81831535f56823d625372717984
zde14770cd9052b45bb4c3e6eddbcc729bf8b88d2aa530996d395b713f6d425d2800b03514b1c72
zda02541a327ea6664bc3f23887db842fd9a253ab328d896bcb84b1a41f529afa5f93cdffc7d624
z1559fdab7b19826e0374ea373d13a8abe457ace09a3ee24016c161507b4ba25ef226deb7be6be2
za5e72953378616d04b8bd5af8e29fc644893555fcab00aa8e7ec5dfb974c29273097474600120a
ze5dbe738cfbb40703495d128261e466e08046b882b871958e9538ca820821245cc8c4fc02412f3
z306983675e5d2dfb90ec95bc66fce1bbfbfccaaeb66827a35c68951f177b5d6e1b97154a153e0e
z07f38b53930ae477a1483af60fe929c25b311008186f11a925aafec2278cbe139898624d549094
z6cb3f2e358d02e0fd965297662f952dee40532c0fdffaae34df8ec6b6eb2a298ba2d24c4a1314b
z4820b976be24c5ca31a88cf9ff57033e20b5bab7476d5d21c4356b9fea28100ca1f933460b4f97
z01f97b5b2e3dc1cd37ede14d5369b5e50bafba9ced7ae02e9627f2197b92183d42b74231e2dcaf
zc5eecc263ec1a0aa85691f8d52ebdc607648b86a0fcae4cc26a0839a04a37dc75bd7895447eefa
zbd071a26f2d642cf86f951ff156926f4e1cf1f00a4cf3092bcf6061f83b80cc3ea59c583b2c843
zc824939ba31c3781eca5b8bd0cf1bd0183fb203cf136cf48bc312afeb23a5779e2c578e08cbf9f
z6face30f115ee7d87cf740f8f7870dd08ccb9109dafa01a0755a09708cbf5bb65f1911415f6e98
z7aa3a7f4445fbaab4ed8c01c71fe781d496585600002596dc69fc7a923c3c2f278e33677669ec1
z508d14877942cdc57b345312108bee68a5c019c81e798cbff1a2556022f21b3aeee381a98fbd31
z71dc051361c5fb4c9c34813734fd2ef716e7956cb106eb6d63023f4c3d8e346ca5f8f801308d28
z28d9eaa6b0333ccfbfcc6637e2ba1a611070bc2b5e306d5af3b6b15936b67647ae89f2c864ef3d
z803de7f0ca49d23100656ff0c91fc139b807bbad9fb5c87cf21aae0f7a9752aa4ff467de16b486
zd2d07784cf96b3e176ab0dbaa0653e1c3f3abb19759f2424f56a2c83749eccc83863fd1c8ad7d0
zf0759891dc7bf03e43973dd49609a4effe220e6151e743f8b83c2b8248a2b49fe70a7791905e34
z4ea02353b58e6cf6271fb3a21b68afa9abea43625e1c5175e587059f450752470c76bf31a30c16
z6157fcf5c2b3208749fd34e4c91b640db3312803f80321052bb181a26c5ab5728d493f004d1130
z9ae9308bbb9f3178789be76d4a764356469ed1a16484d1205d760d9bb9b52277bbd2b42c8a5f10
z183ae92834975ccb766d4d32a2c0e4254b960941eefa5edcf8b180ba938bbfdf536fecd32afbfe
zb0fc7e868207a693e901c5baa14d01efe7d432a7f9f7f795c6f83fad3515ac33ccabd8ae9c8b27
zdc276f37d3e830bf10086c67dce97fdb9f1703a087ce6cc00c77059377fad158eeb5228a30b0a2
z31c5746009757dbc541618676a64e63e0177b4d68c9c1f9ce4ef59bf259bb6393ee65f61961ba5
z887f1b6e1f08fc1b44756510369ef3c8c3f7174db63f38dafa6c92857aeed038911a69958225cb
z6aae4f50fdacfdca70fe4e379e4a5bf02d57dd37e9e53393f584929000eac54715b702597888a6
z9241f2180f2677dc86a8c65ac35add4e1e4132c16aab739ef99efbdecddaf272087c55c0163c6f
z1fd705996d61e40f6863ab1e639e539e2ac8833b756a03b83815130b396ff748e1665a8959072e
zeb81cb064f0f39024af7538f91f4cfeff680b772a7548dee3c5cc23590abd005991a20ad171d2d
z62134ce03c0718d71a4601df61db605756c4c16df0e432297ab05d44009697f0cfb76680ae465a
zd4c7e306da4f22af944e5f19699b4f627e53523d6a9153af0e5f057805a2891f190c8d3085fdc0
z4b73f47aed50e138558a62ae3377286e6e22f38e47d61eb09f04d2fd80fac1c62d8f943f3198fa
zb4071590032afcc4d2f355830dd894843eaecfd1d7a53d7dcd29a906531cab27622b553eb70f4b
z30b5c98c1994069882795d8a2c5e6b35b09a4d40dc82bb81bc0d2fab0f36f943d988d676939cc4
ze0649b7da063eb8f38d84600a8f81d9799c32134c6f758a5e9f7ea1df57b7040504a3f74211268
z3e2a7954eacc407d749a5a7c04fbc9ea0cae4e3c674b141d2355c0db8a9acab05f8668dbfedb79
zdb4ddf166581e03416305182c50c9d4b7466f688324a29e11f19e3bee368bea33db867c72e9d15
z92a9e4fa52dee0601250e7e253c9ecce89d560af464ca3052b2fdd048e3bad10d8045f915007f2
z312e88d72873efea22200618cebb14f68231a66d29cef8c375ba2c366c1e192062cbf2e6e60915
zab55d4199d8a04e4cf2eb531a00e4dd251bc09dc5360d4f2added1490649fb6c798437c3f58df7
zca34a3d632aa8037e792a7e76ed4d5f96ce0ba4447c3fe5a7f023405f7fd3b149d2327edc25b99
z677dab818f143cdc9be48674309e9a299b1d7d0bc9bda7b62d032fbdc80debc65821994639959a
z13f1fd50b8711a2086b0b8c76c20dd69cdfd4e39b23db9d224436ab7dde087e91f51f2420b46da
z6263e7c0ff666ecddccd00c4e1b47227d77b06de988a9b406475ac229151f77ad698d8602876c2
z2fa417f335b40633cc112f107711759e0ba0a65809a4a89ea6e7d69c96ce4f6708e4d9b7d0370a
zb6f3b0e28bd9366167f8b0f815e18627942fd3f796e5c36e19053ee7c57888835ef3d96f120600
z9a601660f7d7e45932222830761579edf4f7165cf2e26b5ba6704e21b3f255874627e989c187dd
zb54ff03160da1d64f20e4d78a9e78e3f944a6b31002055472549a5b09186e537a3fdc57ef563c8
z5d9875fe4e11128163562608b272335343a82101e2876a8ae76862354af445669b180cf60f19c7
ze51666efed5cb11a64854aa2bad368945f062681df6e8ac36a71a43d4be4f3eba8fe63a992ef49
z782d4f0d92600d38aeebc4b26049224d168c7161f80b9cd6080262e2a6d511c0c1d5bb26f68455
z1c65c6052cfc520fb07f677340adafdd28bd287420cd44d9150873c8c865e5a62a2ec54b6bdff1
zbd9409212a4ecdbb5e73714803719f976b5e44f9c76798daa91f0e233fd969082705da7b88b63f
z1e1b107fa4bbd7744e4571ee7d7de6fbe6ed27a593e1cd8ec0a380b6d7a574f21905c3a7a3fa9a
z49aa51dad5faae166eacdce6cb9ccf3681718878ac0c900aa03f00ce7169286447e059bc900929
z55fe8fd97fd30b774572c7371522188b08c74f3842d718294d12591334e42923fdd71b69bcff46
zeaa2774c04778d1b0a43418b511d90baae2b8d581a25dd7bbb9091bd8e28d21b1040b9db0f2267
z1368dcbcc6b3a4e64adb6f72e6d6a43c3aed93a7823252569eeb51df52e9538de8fe89d113e210
ze08d8cb9fe3a1c7aaef22d2832d310cf3a402f3b1bd99b2fec2899a319b4e7b4933530d8297c27
z4cc5139ff17508a7d9e443d2c89ae8d1436b9cb65d0bebfec169694871e249a11f6b9235c67a4a
zdad0e8c5d79415a4fd137c975a3b23f47da1d0f581f95788a42f2be9b5869957545c6f48ffef5f
zdaabdc73a0183c91883214837c9e516d5d3bd11dc458be0140d5ed8f58d44ba6b964f8ba5c11a2
z6866bd039c0b084f5a8421daa218040473046a1ed76515d5cf2bd8e2f1105cf66fa951a18e35f7
z4ec0e7e6d543ae66ab253ace33deb02ef6bc6f671fd379b0635e3bc6d0f0024607879ad175e166
zca809c9c73f62e194cb151fc1e245f8a17e5053eae20d11b9f413c748c5a8399e5f0b8f6052ce6
ze249b59f6841220b351fcabe9da4a18174a481872e547663b60823aa76bd0a9ffdfb1ced9ac058
zdf7a36d89699b1b073151b1b46b0a39e14957a26bd24d7557f2cffc7193f759e3247ae80beb618
zcc2440786aa805cb5681d131ae21875cf96457be6f74fd07722c80d334f39118b302d26a13146d
zcce9560d43e34af44cea9b2f55b0c86d710b35eec43730762177a6a43f4b64d0e16e51355fd9ee
z07f0644f62db087077e0fb7a63c4f59863ec4fe9d54cc32ab3193615a7b1e786e55c849418bf30
z5d57dfe633f8dfd06447d4dc5d49031ce2c0cfe975d059d9f4d7ef3d78f7a627e863f51ec42316
zb1f5b94509f544a0f899c71aa40bc2798d323fae59b61a0f28f6d952c0e71e2eb63fdbff6c8b57
zc124bf063773c6cb39509462587eaea4b953d67ccf5319338b48259d326bc05fec3ff2ee50ce61
zaa47b8480d057e16e0a6e493cc9f0ca89317b307de44fc44ac380e16e0838b4eb2652d5815392f
zcf975619c4dec33e2235f91290c3f4864b6d5105734c120d5a2942ae7821c02214ea6783a7b601
z02ff6b7121016e9d816d85abb2bf6cb744b4634aea3e3dff4bee55b33657855858b1e5a10dbd14
z0aa42fdddb1076150b63902e2646b2f0c9d8b07a0e47d888d773feb37db9af1f5c849d9420bbe2
z76835a752377b16bf2384d8ecdfe531310a3d991ac644ebd90cd40989fe358afa754cfeebc54be
z22b1ec3188dd76f1ffce9daa77f47d5937c88fadf88927560e12a9ef96d619e0b43c8fb68045aa
zae03d5b38df4294e1134d7f4650f0ac9d11dc1ed53d884de0e6f64207f3a52d5841f79e3b88241
z42f5227d2e4066c64aec7b29438604fcfe433101709d4612515fafc8a1aacc373a4eec2925f54c
z3186bf97df339acf4de226dce19af3ea9a02105ecb7956ec138dad914f7612b6135f1bd4fd159f
z6c72b9928f109578eb7b8d2c90c5ea4257990124a84bc0253f7e7345976d1960c6cebb60fbbb5f
z1f8d46898fbf53227661a4fa7a51cbbfe1dec9132383d43684b1dc69d525a7b603f1eb8efb2052
z192071b403fd6587658dc3e02c2c543380fd402eca385fd7df528a291d5abb3bbf8e0137487ac3
z24dd7b51a0e58d2efffdfd45b9587991d164618b464c2fd42f2f93fc86155678332b6171859d68
zc7c06884acf654960ad2ff96c25d28497e0157625d7194bbdf5fac50082ad77d9eab19a5a6d626
z74f840ccf27ab5eff200404fa06117eca4c5d4d863f98ac782a55267fd177826455c28712327a3
z63572f7be9bc121b5cbe81fcf4b9dd68b36291dc8ffc760ae173a68fc06740dae42701e83a33be
zad94e5b283344dc56c53e66829e1e39ec3b72323fa8cc49a2e13c5b97daf04ab01d87955c15908
z8d8e4457f55ccc872c4a0f87e2079b479d3f94e35a823b054cd52563df3b9315a96a82dbeba614
z8dacf12f93e92d46a2d3497018a60eff4c903aa4893a9b19a772d557916c1f6109fb5b7c69df79
z4850dcb590a90c8b8b8b0b628bb3d2e924529a8bba06bf697e95712591545ebcd8af0774988b1a
z1ce483e4d21e183d4d64e2cb39951767d87fd4590565a1d0daa6665f378265fbac177638ed6869
zbd9fda22ea1008bb56cfc6eef6dc60085b898ab013ff94b81bd9c174868f609b2aac5c3fb0844f
z552f2b1b8c3f93a8928f0c26cf12376b15a6d3b4c1da76bb2187487c178e62236732e16bdc11b6
zcfb50c1a46f47d19be965b6b7d800718fa0979190ba25c9bef933467a85550107fe97a8389def4
z9da333a72b367c0c6c35af7418cadf4b8fa535b1cfaa57b142d3ba497b4f29f9344399e97e473e
z8ea9604e370d66d284a9b1f1219ec4ef9c36ff6c94b7df8cf42a441d0726f696bf3f9393ab99e5
zbff44f9f21836f7ec44ec925ea165114f9a8986624a74db2063665d27332f00e8f05e2fb04e7e4
zda9f8caa6d2daf1bd92f364c34a27aff443da7e92cff6d615c960af2058f3f9b59bada75ffb0d6
z7c9aea620da711f6c8c8de5f41132c5f87a4aa70167f669e2361f54818446224e959caa5b77c00
z2c12f80477d3041938d8396ac132675647d02c7a1e43feb3536774439f34678b0691cb6995e349
z71a1d6752cbb9dcad647cb6fad45f2290d36ad6c69eaeafebc4747e322c6d9c12dc2daab57c9c0
z341d9ff90dff6ef5073493f925c79e3fdacf82baf969875d4cc53c24b71bfc9d5f842c162f30c6
zbad5e7175ca35c54ef8253ae9f30a01013c152e583d94016e60bea5ae3b1f8bc335b9bbec7cc05
ze5b455b156179b4fb66382e5f3644e9f6bc37168a2bc14ee63b5fe3c81286dae807ff7e345262e
z340e36c098df9868651dcb7eec3af91e1905a13841c920cc06fcb8b299a35f886f679916f47862
zf6fbc7c6c75299534a8e3da126ad725d013457475a75262165d9d330a5ba96d00692177f2e21df
z4a80bb1f9abdeb10b8a2e8dda3cec6ba35f6de31cec93b154446ff5512d759971dc6f58d0064b1
za839d89046f60a769a0a7df7bb6b8d072abf1eda8ce6260484e1dab2d9fff252d059a3b160b21f
zbb609e4d243b937eb84aab060b49605c1abf1c16fcb996d5f702f237efa7eef7df8be31961250b
zf5b7c82fdc9d1c55580adf0d11401ddbbb079c0a77e2ad42f7276cf9ef7254f6e29b95263be77c
zc43dac7397dda666b9b07822c859f4bee4d851097f735963a7ba3820521e711e90ea4f793b1fe4
z58628e5589ccd0454acb58661104cddb3ee879e94d9990b9140baeddc598c8d3411c0bc82f0e71
z111b591ae4c7ac19362f6a1b0761d4a0bc2dba602a748f85d426621c92053c33fa099db4472e91
z6246f89156af16e01f7a149c224d43d24ca6538b08250b1c040c628de0f236184950281d5c9f88
z279fd4c3ee234e91938994b1bf629b96df598e342c215642afce10604fee6f42d56a74e6309492
z95b00a26dd410ab36a7301da5039e5c09341e3fe3cbfb441a7235656b1b122acfa5a3a25063ec4
z24bc0a76a9aad8d04e75e94a4f9db093af36d4a874f1266319e2d118c51c52594ac57fc4401609
zda6713f9722a9dc8d56a941992b29bda39200df8114811be2397e1d4c6073c3be5db7a70ae7bbf
z7346e72bc4d3c8ad9014dacee567fc8bd03f38b85eb18330b754866e26fe201ead083a3c401602
zb30386ae699a67e52403336d1ddcf0f036f68b61dc6346bf1e0491a8cef05312545ac14c3dec50
zc20005baf3296933c2e81c5f772495e4934bfff84c361b85f0969bd1418d4ba2ab91205df706e8
z4a456078cfe6892d7a19d7df636a0b776a90ade0cbee0b5849357dc208524b3431056b8f453a89
zd7e14dea6b24dfaf5552a5ba82a6887cde2fb3bd8327ad3447245e1c3bada87f89ff02edd178b3
z46c7c5328677b9546e96a4a53f951c59c74ccc4d764e43ccab78bbe77bd6bd45cb97687f298829
z0f1f2453d6aac29ba01aac08be3e66c407498170a28102aab33f590e6c54210043ca76083dd05e
z47836d9944d748abbad54f09b2604f2773811a853939d9cd4b48767c56ff1f2700b12a35c9fde1
zfa69a1fa3a5619a35395ea730fdcf324c77991e2bdfd96a402ff359851c75caec518457e91f9e9
zd802ccd333024728f0cbb38d63bb7f9a7769536b012d2b2f48f7cbcf6224119eb5e4491ce7a07c
za86913d43bba582316c714a3b4cf4261cf3ac41ef9e4ec2090f95d3be31809c213c4607fff12c6
zd69858e69510ef5c8ae5de1d862efd9d767f88e1e4a1dfefd6b89df32f6b9c337478f18a0091ee
zd6c3e6a48e6808ee46796002a6385673462f4811ad2d7d1f6029eb9ac110432db23db9fdc8ee3f
z07dcae74cbe2a5558e323a95b95e20220fdaa069419de3f58a177f129997a4adcaf6c3e2581d73
zbb5dec6be7156727ff8a71e999dfec92b7184cdc52f69e1c5b7ae03720d90c9f590648ea16e8c1
z98c8852e396c5adb9a13c09f323823f5c6a5fe59b0ff7751d6a103636ceb4df0402126df003c3b
zf292b60e31041cd56fd84c649bee72ab47a5a22884d3f7c854563ca76d72adcfeb92dadac5c526
z704ccf8fe897ae45239a83afc4a2f17beb3457c2badcfd6afea789b3da9ce5c46edd731ce1b1d3
z586c9589a38a28f8388cb713ebff7356778da9a0d092c2f3e59b7074095fd8bb54f9de49449dcd
z8d8ff8062fa38ada27bd5bf286d789fbc85d4bc8bc2a67dfada8f3def9cb0bf774bef5ebac40a4
zbde0cc5fc19720a423ac8a7561ddf86d81bc7d3e11bf1f64ea3feb300351315b3480fd3f9e2f26
z366330bcb4d54d22c125a9bb476878b0dd084f27131832a2fa47368ba8379b1c010eddec9ab000
z285848b66c3b88d337417ed71892d75fc5b2bfec39bc0b362a14dc7c4a3db7bbb1b8bc4475ef8e
zdbc1ff550c524ecd6356642e0f8c70043cfd30d000a4d8da3f42c6f52ef4057cea3c40b2e845b4
z2831c4a7d95cf20f9f78c25e4fbe7535c0790559e89aca8a5b72214e9ddc51419f732a1bf71c7c
z9b020a60db009dd2c129107cd96eceeff76bcdfdfb2e5d4b9783bbcde39c2f4516db19a06e6c93
z1aaa9ec3cd7b021ca0b189175793f1222c05363776403f4ed1c9820e30d0cf1aa04826575c6952
z080fb4ebd8daa257c6eb2bab28ede7b40e383fb93b2c69dbbd860da1c98080e9aac16efe954e2e
z452ce1cb23b23766e382c70d0e625c7232bdaef8327fac427d873670954766be83438529a93e87
z736910363671031ac7db31654a17113e5557ddd46b3a91cf1b2d2640bc1e7d615ed6e68ad21400
z1d6ebc7208cbb4ddc03c7d2d6bab56f1e198cfe3213e30404f8388e738868300fae30bae625573
z9f7b8945823f1d0515b4db59b0882f5c750d0c3c515f39eab6f54d28b0cb48c073b16fe55791ea
ze250b72e04943636ebf4fa1179997b8b3165d42d6db665a05c07cb9f28960445468dd0c84c245f
z4c3a88f1b6954655c4b95f6d39d5ce0e9d56a93812be971955e3be7db2bb5037953f27daa8219e
z7b115637e4bc691c5fc64705d0d153050ad7c2351ac79ba0416ff06873a4a3bd0f7b8aba670db2
zb64ae1a8b20d8fac6e9c3a82f4e64682e7d8ac72d748688477911aa132bd04f28cd7bfc2440168
zcc568ba4ae129bf1db1c5a891c1b6593a94532745ebfdd576dfacd3c1b60abffdd38d2db4824b5
zaff2019f53fab37fdc0d003d5b5e8f95e974e944d7d1f57f1b11380c3a77c78cfac7c9f919f9c2
z8c774525372197d2a5a9125d8c640dd1411881377e8eca315ec2cf37309ef07f640b9529d3a666
z18b5dfab48aea750ae1e003aa0c1796d391f7ed311b1732931bad5a50d9832bddde2c31a4d0c22
z793c5c69510eff0a6aec954f8e8655b9c9ae81ef04fb58bf80098eeb7d0b3174ba2d13f25a3076
z4b881615ed89fdc25655ef3539e8fa13e6b879dc715d7832c2cf31eb12b424cd56bb0f03b469be
za8c72037d3911fdfc2bfb1fc586611d37d93989882b2925c69dec1a3664cf0f68e88bde5624225
z308584af13bc99aab7fd934d79aad822cb2a7a261a21e830e2e7122f450b80416678ffa42031c3
z66a528dc398b29a6a9adea87ebb20480997ac73b0455376f214f5630d1adb0aacf4784fef6f6be
zd2bfcd121714a0b90e0fcbf8d963267f23a08a9f996d197f78c60e1967218726d1bf69065b4085
z54e509af4ef2a38db74580fc24e1cc01e663f07affd589f12cf700e134920d66bf08f8b828da26
z9a6aa225042b17e079ee68bbf56565ceb39e423dd4ffc67d20d7725c7ead7cf1f23040efacb681
z2af814bb599a724fe7e48465bdce84d86c8c64ff813d117816f604ba70a4426eff499b15241ad1
z274a71a11c5f770b0f45b10dccacf6e497a16eafd9abae9748e1fcca97b9dd0696505a39d068a4
z8b12eaf4a7fe1bccb9ac548782fb62db32236240925de25e880bd7b26608ae93c1762c1bc2709b
ze7fb1e05522a53cecce2664a9569e24c554dd6ea5f167ee8dd43c722d808cd3c1230f216672d0f
z5c6e8ef5e96ea183a89c2bd62260f780347055330c1b3921746168808e572353930492f7c805e4
z277e1c0af63d405cb059906864c74cd23cca9f2eb77150b5cda1c53343d13152a587ce4fbe99b9
z36a4cf86ea06a992e4aa05ea365e4ad976b17868129871ee868dafa735d77e98ae6d08cf6ae1e7
z7931c644c734efbc584806acf159155d424a27eb8d75f1482a966be64037b3c7f7ceb89c43bdf7
zf2a3464e58fe490383c175110b73eb36c3bcb9bdfffdc207e1d515714584b513d772a986b92f0f
z743f5c208c537b6c462996af3ac023a12e923f995833c2911f2bb61b5d2c4cf80849b171c4fdf8
zd0d788a3f3d1ce43bfabee7e734fbd507a8bdba5fd9da767d74389999b6f652efa0a9daec0c157
zff31f6fb5d4b8a29ad936c84bb3df75466dc546315a7a2465fc38e452e880fb29cf1854e1b70a3
z488af84507c2d2b8ebe764c09af5a2ce3a5b4d15dcca967d6c1c883a6c113e38c82228c0df8c9f
z21d2476cdb301778eace965beee8e141867ba3d508571e8fa2e6adb205bccdeaf67c7b7df91e2d
z64d8047053780b161751ea7a862a17e519a4d907cf1bdef105c2555f7596f61267eb70bb7127c9
ze55ff5c276844e7257f80ccefe09e0a3d96d01fab0164018620d7aab43569cad1ec24e35561a00
z8ea538307b571790ad9ae1427df13d536bab9cad9a63ea9b0c4ac22ed0acf21158a1e5fb03fe81
z049a4114ef20de31e008b83837b4ed938e62ee3619ee7e59cf04dc92460f13a2f7a6a77536d340
z59b6148df584f0ec2825a24d854096ffe6552e2783e031584813280f074578b957594926a0a15f
z5e071086402a9a52bdf843a7ebaff00b98b408a447405c852fcef021c01571ace65ddcfffdaa4f
zb4339b3a2c3df4d7efeba86ae17f58947c7737005c5bb9ff62efc02783d5e6a4a9188217
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_express_pipe_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
