`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc89607e51
z10be237a0f267698e71d10abe7fe7bfcb89ad8328c1ba8a321747d68d06bc12218898a6da90abd
z0facd8cbd49e0de3f8b76f4c9f15847cc12f3859be8a421e35627d7d6a8e1fc5dc84e8c99702ca
z6e230414ab99f38a7b3566a2e20c1f814f5ad62218b46d74a3cc59c181e56c2e367d0900d06cee
zbcd2589ba8a427f586776b1c724666911f4c5155ac863fae616fe372ac43aeec37b477bab15d00
zea341c261ffd149b8cc9095891d23623fdc4ddd0905719ec3fab51d5849f3c100fd132dc4604cd
z1f80927f0b9794e4b0693a84bb6c6ef5bbe9d24e8b0b47716691923948157aa8385f7e4afd19fe
zdb0cd636f9b0cdd8964c79c694cae774bf07c8e7d3bc632194baa0674875a1954c839c418faff5
z98f407cd32f528bcde26020d24f5bdd2d632ac649d86fb96214f236c0d2b98efb8ea5c0b193839
z938dd813a6c09ac91e02ca68f8def53bd8a09ccf661a9b17389d4301ecb07c35b21328c7dc8790
zd604973c7ba7e0e9c05959a639e4c1faa7c50efb220c5f9dc251c9a30fffa21443e5074ddf904c
z2ffc9302d0278a56040a26b0eff9ada19cdda364f4acb0d8354c6720019fde9c588f4183467a3c
z8698e17de91e5fd88508e7b9f2015e959bff9e377e3a23340960580b0638e4e528cbac5128fc62
zbe7fea4a35ec4bd0f60ae5e3dd6c658568da68760bbc67d1c5b41ecfbd31c88dbb3c99c9a9f33e
zbf6c6c6a75629939027b4f0393a1fd8e7b8929b766ab393bc09ff4f120f57246c4e3be7348a4f4
zb18e32e725c4035bce607fef0b6c44b64f5eecad6b762e3e68052bd62fdbdbf7f30be7b9ee608f
z1b732e4f97255fed3a3959215793fd02854e4388dd84092875883845c204bf3be786ff76649918
z4b4b513b530c456f298fa4c6b95e540d8bdbc0bac63882a157720a1a46cb2b0d5ae18f9fb0ac59
z32adee152bee0d06bc49d386e730588da659c81ffd200f26c382dbb8a5b91a5db440203367d46c
z1ecb1a905e9973f4abc781d84ad93b728b6b5be60c206e0dc908dfc8d9ae4064d4df74b0ef81de
z997aa67a9a2103487483e4f8c4a4d180b9c94f05fe85feb00cdb360b7831345a6d765093dce0d2
z9077cdefa7cd9fdb008b2e4a880a80b868ef9160702ac363d513e44c74b4e04173651d26c77af0
zcb746fa796d8f46d63acedf4e48544279e0c2cb966134cd604bad7f133ad279619b19c7046254b
zb3127eb37b6cd2746870d20b7af359001bfdff8d05cf95911289db15d70f67dc2a390cd6c5ade3
zb75609e0643f0b5aab17787cb20270b41768e1592e8b507005b23dbb2106131bee5d32493d82f3
z88b899a79dfae5c5a8bd9e6af0fc37fa7b5f219b19f7856e4b73b0f13d855fbe207926ae066ff6
z12878936d23631fa635a22763a713c855e4c4a2ebb1278c4311dd7be5f4db595dff7c5c99eaa7f
zdc3de2c787ac5569737cbe7bd9411c0826d85067a381e361dd0a564c33625523681b6b9eb30942
z4a47a651d125f7cd3a985dee48ba771c6c3a63d3796d91493fcae030e6756894adf63222a6ba20
z36901f86bd1842ddc0366f5eeee2f4801058bd8232e3c07c248306b6b9eafaa57d74b93f74bc8d
z335f5cd83c78989fdca67dbfa63eb2323cf76f834247ed93e5e36600d7427dfc7ebd04eed9a4ae
zebe8a704ec5a509e7147a8e8eb39805d9530ce6d27f131e5216c469d9b6cdf030efac8cf27a52f
za4113666ee5e41ce9b7d80ccdb1c042b772421774edb35983c98ed34c905a51777ca15cb850e23
z3f3d487ec459a6cadfde1bb588c17e29e7a4d36d6245dfa18cf00391e34812041a4ea18f73a9cd
z7fa60095be019edb94564fe57125f7cbdf83a188c5d155db6143005cf2238a1eabce2cf929571e
zc5c340ca71d17bc8832c840a0f1dc56a0598ea1fa876faef2c2b36df424897d4a827e310254550
z50511d40e00f75e0b5d20cb26109ad4618eef25bd9782988cee9575a9f5be7c1d653519a1dc1c5
z67958de4daccd302e359e032236a6324572c6f08bbd7ad1eb659a8b311f690bf1f477743183b22
z9e994b7071b1cf0a290cc8f556b97c00d78558d5940f8946d5f6cb0538561ae83ba01fe5e6c2e4
z6029ca01c4a2d6e807d2f5feeee6f90a9c13fac446f3bc939d6f245759bc9d58abf31ce9e07401
z63be22b0195e19a115e8bcfb0ca5d930fe004df77d42d039f096ecb2cf1cfc629a1fe3d69130c3
z1a81da8ba40fca1a6f6527dcbdc89ca530deb325acd72a2500846a2e804812d0decd06d397b2a8
z4f73b657c0367e25dc6b09af77377627819348af81539d6bbfea8ff56914b36854ce9d8d05aba6
z5f9ee1daf350e4cd3c8bdfd0a194ac70d00ed5fae759979f262a3da20a575fbbbd86a834bd0133
zae81f2ea86a0ba3323d996238cc639c3c847c1c0a8eb2a2fc42ad94c8b30493328ccc40bd19c4b
zfe16fa4ebf77dbff1054b44c45b4fd798c0bc931f831e1c01978ea40c0f5fbb7aa43c9eea9589f
za35c08d3e18f662d579633b2c892165e4282df907676e7440e30e26e68f4e643eee268e5211060
z79b142ce04f18ae9290fabb368ff07d759bdb27c81cd980385b3b55d000e191c54209087835e3d
zb03a4483ed49536443ca15513b4f4b63708650212bd16636e1f13c03acdeac1563f06a6fd1a3e1
za6d14a0468e3e297722d3800be43c0fa2d4b09a06c4a6d92b46a2fe93d841efa9ff5f2bc4a0452
ze359a35bb3c78051babfd8064bea4cb381f2a39753dac172bfaa2cf188d3a521ad4abdd0703456
zf06f28b26124fe06f728901038e320f7572db037f91885817cfda35a90b98226cfa5db28b7d0ce
za89c58876670393882d7333f5cc3570a67ec6e3e119fcc3831c4647a41b285c2c000dff4ca9016
zec47c04bed0e40ac94936c84076eed827f38ada27a372dec7beef2ba127f6057651315e377ac75
zd574f64832ad5bf77604ce85071d0ac5e3a54898470c9b0a3f65a0937ebe76414fa252c85f5b94
z383a0640242c7bab83657f7271f9e12bae4bad85dd0c40f763e3adf0376d65294cf0b731a1869a
zc66f31c8ff166b7f54a9d9aba7564b4ec0a48900e487b18c85b1e59080f2a8e65700ac55c43c88
zf0ef1319bd422672a642fc6d24191fd7df80577832ca869d5e2852243c46f157fc804815b2c902
z0ddc992874df89a5e950efef7917e817bad0ecb3e5271627645a61a4e5ed31dd2bc8fedcef745b
zc9010044fb22fccab5338d539ed4290fee9a8683286bc73a27b668b5ae0886eacfe3ccef14c736
z8a4c997e78e475ab5efb04f9f60ef46d938ced5737fb01edb0912c30044cc2af1b258b95bef533
za20078e3726e52b5a34fd1d5cf645ea6a9d851263f8ff2128fae2318504e6b82532f47f7cdda89
z7557514c5c0b4df73be0af007d3a9ce67393d6d660593e578b3e4ead0048743213a7e9602daa35
z865f80cab744fd4118e4a15b5451e8a4abc72580c44bde5f50c528940a3183c3e6aa99512769fa
z416e42be4356dded5226e5b86f6d09977e49f7b95e8ec25ba51646d930d6496791771d6c30bdf8
za19e437661df500944edd605b6ee44754a869e6d09d503b91003bd58f32436ca7bbb3c819a6260
z3b6b9f47741b9ef6d76e5326ee48a610c7a01fa92d0d7db4f1215a4d3402075cec828e47133e39
zc87d8f752691b8a52c9dce28f005da1dfb45c3681f09005a1ca6f411e666757b38ab8bbaf19511
zc2c06cbcdd9edc3bccc8f989c9d8f4c6cf2ac8c2344e12fcdd5ed0725c743cb5cd745e189bf509
zbddc493f01e563000794ef54bb9bd597be615807402a1fdd85423251c2fb4c93259626d648e832
z71f9a6e41f6e1a55bae22a96bfc19d87428fedec2242cfc900aa3d8ed9ecd3ec0e4e216c30a5ff
z4d97509b8df92368c7156bf46a17d66fe01e976e4142a9cfb81481744a86e3d483327092ca0ba6
z5a6cb1a7835166134d1583a3d9223bf6cc1cf0bf5dac1d16a260f163c09e9e671490f2461fdf8d
z8c0f80255465ead3dfec52925ff9750a1eb879a3828325730af53474937d6d00de59242499b619
z7a125c8e67885bc80d4e4d8b69436828a00aed17f6e485b79f055fbe07e912cac3d5837369eb2c
zdc1b83d2d2c9e774bb54a4d58f694e2e7155349a8ca1a568ab8bf493070965d891a435eb6a1591
zc30cf268dd7c16b5090816862748044b3ef3817d492fe902433a87356635305ea9b91e0a53dcfb
z2630a5a9a992e71fbe26e07767b00e60fe63f141f4f91f4ea26aef1f7b89873a83a78177d2cdfb
za4d0f57fbed5a15b598f250652b4a7363250e74a99a048453f60825ca5e1e459c016d79f7a815f
zd0316bff82c751c925da29c4e710e4d3567dfdee3aa2ca2047cde056ff36d8fbaa1f06cee41399
z1d1980cad255f450dcdaec6dd3762d894ac3b52baff0232353e4fab9b62a5961176960e272ce4d
z04fa347ee80442d266a8477e5318c5e869fd9ff60451e847dd49ac597591ba90c3f0474828a07a
z1f8f83cbc2f604f5dea0a7b6317cf6535d6e1ba9b057898285ee030608d3ddf47c1eb477909796
z510dba8c47259160244b7f001a9a21f8d6c699f8040693582530ff8d34fb978b248dcdba463dfc
zd93f2fa6223eac068f990e36231145688a65e698905fa44af70b1b52bc71a3aa950757b069f3d6
z574fd15c3ec839e4e08621c6f98d483ef7604e3bbb9ec53ecab7bbe9e69969d3b2ff6ede408277
z443a4d8030ece25b945ed27b2b1cdee0701dc14b1537bbb813bbfba6c3f38c2a6a0565319171bf
z56039447a3659590945a0935e5a7094675fb6f7370dc6885d1bf1e212ae28050752ddb6de3b5e1
zed3b995f2ad118270247337a161dd33a718a45d589844c532ebe5a360b0e6cc4d49b4a9c3c80cd
zf52cf094c9e878ddb6f93298bcd59e4bf78367c391c8d7aa64d8be7cc53c5102f5300e232e6956
zc4b6296195567ffb9979506fd98002ba9f2e4b0cd2726fb95def98ec74c8e123ccf396b26f371e
z62e531164c61c236f1ebd8f0c7bf26eb5bdc00df80e4b8596bdf254d0bbad6c15624b5e02ce311
z656f02b731a7f62ee22e4cdf8548800edfd023fba7a9f8cbc4ab5472362d426a45cb5c9afbd3a7
z08b606887e9c8b79519818628c0b4da271144b4e9db2f0092335f3044f764a1522e52a1e97a13d
z79437a36a82f5750673279298ea3ebc485e2c39ed6ccc93001a625ac0949c2d95f78816a0921c7
zd48aedf421683ba2d8895210a5177d4954bc35d426e78ae361836e4193df56f8d2ddbe6ec6d8b0
zffa7e21c4d8c87014eccf5de10b41aef52eeef5958ad31cb66e73a28cab167fa4a1debe963d803
zcc411ca90d152f4e5ae77728deac6aad5b7896dbedd2d880487ef206cca6d23d56b1803465f151
z70051e91eb6c2c9d56130fb3c882ef092052f909771f34cb954a3c5e9805fa93b74ef003f50084
zf25cf4b39bef0f23d8b3d2a5e2baa66b04b1bea98183a0d040aa4b3a25cccf1b981672499905b3
z6d4ddc4b4ce1dab720a51c24557ef5fd354ada63a5cd63300b8827cb6a21ba311726bda69b5293
z1cfb9ea97b270c58cdc6173adca6e8013cd6120685b3320a0e66740fa99248dad4ffd052c1e7b7
zaf6f5b50e5628e32fbb663cd52fe2d6163db2e6f116b7b519a8b6e6574eb542a61385d8e06d0d8
z37662c3f5a4bf4a024fdc7bb55243ac9f285416a0b6b62678b1bdbf9b59b93bc869098fa278a09
zc17460055d8e42824b065d2654f98d38ef8d3061044207dc8af2c9addf93ca3790e978a4c90209
zcd4e232479ae53435f0e5a0eca0cdacee2caffe51bb9b5f1a89e19725a1b94f6a924e3e9952852
z32360485790a34560a1eeb1c795727fde21e348c3bf87db66da0b6fae0c49597b115164bddd27b
zf7f110639e59dd247b0f756123cea89c8b6c69c6005f39e98e3bb34fe2bf22879ff93821148f58
z50ba9a1d7f5abeee9c071e69689fcad6460aa3b768cc308f2834e2fc1a9f2d4b73899e27057da5
zabee82c0aada1c3c0aa7001ad1bf3939c145c03f35a9458aa1977e36d7b79d259fe3fd4cdbfd77
zb449105b2a71038c6d107a0add51734aee828093f5cc5fbab700668ebc01c4b69b7c3c72190c61
z0ebb8fd2de8aacbfba02afa0507dcaa6716d453b8fecc6399616298076bd4a7101417ab9710717
z7d8be9b139f169c3a8d27c04a6352f36a94c3b77ecbff4fe16b5be14d102b25bd8748d0cbd38c9
z0798271cd5711483e6e059a2c1da08c6822d72321970269bf5b22420d8f9fd15cbd3b3110eb11e
z293c39c1e62a386e5c755de82d30156ac78d898facad94fc1d99d1305d218f45552bbbc21ab03d
zd6a31e0991647a5b7bd738905c0a57713145db212478d87f01903a18a3967846e4bfe024b0e4a6
zc90f27ffb96478c3aff86722983d0f3f42e0e7fb182e3fd53b991ab371d30ac2e328fadcf9f85a
z86fb5f446628f9b1768191823181568564e248d6fa054ac461f5c86a05b41ce2a25fec37e63fba
zc6335f083b14f2953206c0e15affb4e31eb6ad04199357dd445c058a3e671b3d14ac5263797d51
z590f9a2221b0d3011c1ec4f58bc6b8795ab1688666663e39bcc286460478e16c38ecb9ecdb67b1
zde75e9d32a95b1611a3c0ed5af50060a7f0c91bd571d67966312b8b263205dade09c4cec564551
za08d1d951eabbf521bf1937afc13a506f1c249f5dc4a01850fffe18a4b7bdf3546662d00de4e3a
z42a63911a64d32588cceef720819731792b1770a098edba434a2dd597b320599aebee3ef72104b
zff019f84e0710454f5c0e53556e75125d7b5ddd04ce8f9bfba47342ff9099bdc793818c51796a1
zb56941424c0c1969ba561e9823035ce496ea36fcae532822cb7e091b25fc8c6382d231990b3a39
zf64d83e9a0b41f8f3e8d30017e2b70f4d6095a67d8f1292186b67c6ad58b7e1155b76e23b6e660
z79fb883df36ea90edb0fda0d4b8de86534179f2df9ec9948ef4eea3cf6136e7a9283b36691dc7c
z1ffc9ceecc3d3b64b5ba798a06ca0cd5c2764282b562e05e566c6ec8eb198e2fcaa516931e2bef
z669375a89dbbd2c5951021ccdceeaf3c70a23466f67b21684db91eba7f6ae19097101ff76c0afd
ze4544ff735949cc497978745ae00c889b0fefb9b96de702514afbdd3b3c34f95fee22e92f78557
zd7d14637996b688eff8dcfd510ac64f769d81eb6e1f16674b0740e85d77d0ce5bdbd726a4d8f21
z982d0ad931d38dd9ba9351691521e084a7860fc5ef59ebc08531848e3ba54a9f90e632caf7e852
z0df27bf6553d54a0b1373e910ce22900449ab055c7fd7e8c0bc769e052a1aaee0e63dbfb67ff92
z870ef39a5b889fc394550d4729b50a89ac8fcba52268f56db5d3a8f91b7a0621e6280f06c22c9e
z4f2c207685d33dd5f52d6de183ae29a3efdca086e67e6b9562bd1750cb34508234627b4766b80b
z76d9f997fcffc9120a34f1da2222aceb2dcaaa601e3b201cd89fd026d01a95a75835fe23ee9b6d
zf74979789d40f9929fc6db426b76e2f8d393b6d5d9f213b674a02e2f29e99f6da3f9aa689bc812
zacb250a9ddbb533dcc2cf4d7e10ebb60486efc83f36293bea54f8f0976988af7af323aeb965ecf
zfd4c32bba99905097ea630dbf0498fcb8987a60909f4333ed9fa7f63a86402d8a406d7818b89af
z32684172e877daac6f75c35aba04de7bb9c9c8418af9b3a4a16b51ab08951de75df40af9d687e0
z42c9f5592d3862c211b8a5847718ef6ad602450aae594f681044aed152203fa0f8316dc16ab006
z6e0c1ec9783e0a775b02fded9f4e79a6775e39c09128c846843adf0724e22af2d9b7c140202154
z0950f28ec0c4a75c3398ac88de269d8163a0ea3cd7f7db5146c1abd574d0d7daef9d5eecc93032
z4abfe288d5c3cfab3ecce524993faecd64aee66b9b91dff2d3d6a2eea4566aac0474cc30cf04d2
zc4455533b1ffd08a3282cc427e4cbc46701f94cd299ac7a0337be3fdd7ba1d04484f743cac8561
z4c381cfdf3fe1fb43fa245a08cf952cfa16691ca07e838556e680132a81894be91d2a9a979cefe
zdbf7d66c3648e210af24a1f30c8af6ab7e0ea897ee6a4d1aeedb173eb000c41ac8c4e980108771
z84b2d38c8a26d636c9fb823c427785205bedd93faeb007db0bfc75420ec7d5a513d465721c8d5c
z24f5699c8f6b0f95b47b723ad96685f775be3046e6ed5c3799da1ed7ebedc4ed6e341517fe88c4
zff31578468ffc18eb089be2a0688d7ac7fe939c678e6e930985a10d9e8af1de69666492afc0750
z8b7155f91cdc1c5774d038f1a7eb66c61af0c8c367c4356f4da78cf2ae3881049b345dfcfd6416
z48df22bdc58ab86ebc72ded3d2cabbca395a70b16499df773b96f18f4d3d7d994e639519ed84d7
z310d9a2405c9918a1c1a555eca326b2bf42e31c700678b954a030407eed54241d762f01a9bc17d
z54603235300290543cad8e895ed40fb492b7a2d516b009509b4b2cb9d76a45002efd8745c20f4e
z0ba3fdf15bf830b8a1ab43c502a79405a7f88524e529ee40b2f1035666677e37bbd4d143f09243
zaa0dc27deed1d066f675af27311be21d1dc91882597e39504a67b89e60a75a272f471cde804e06
z81a1bc2ce8178d4c7ea762d595d3bcb6b074bf7adce96a0a27cd9c7c6a2e07ede39707da367ae7
z6f8a5e84ca18c6077bbcd2e082497f5324ad401dd9e1661fcf9a8c55cd9cf27351efbd3127d721
z8738dc2d51229a3fe97afb1073fa23579ca21545ef8b8916db65a256caabac0350d1482a0f747d
za2fbe666463ff624b2507067f56ee23268aa22fe6a1528bbf99022dc3dcc3f9d512c2c528fd21d
z4677162b2e1e3de8e7bf723bfa61ccd8f64fd00aa19f65db2f8038ac85915497a830cc76f500e6
zc0c829860762a5aa97fb7200e1e6b4146684d15dacc7b68ab3eff09368de1b95cf1804b5a7e2a6
z5c5ba2f8ca204b224e8eae6866190bf819c4fcbb38f489e0e27e3f44b73a391cc4088be7bc99dd
z249d3da75083b9556cda841a61230dec5dcdde6782d84f1201581388512dea759f2c484b684712
zdfd8c63d40ebc8253c0ad346086f6b39dacb40622a9b54f1e3977cfcb4bd559c32e3b552ffbcd4
zdd98789426bb5db6e4e0aaa66a2e841cb805f8090c44d4ffb6b3cb82d8c8527d9bf06eae7059a6
z632c854869f683a65b48c809326e4b2ccbbbd01bd872c48a4ad2960aed8ff6c1c066bbba5c0c8f
z33795580626eaff84d0b4bcc72d1832fc8ec3a5b64cf3dedf8958419dffd77fe0d40e0ed0f01f0
zdef30cb97379325e00fb213d56b81a787a2361538b56fb064df2e2b49c3172378d2338cd8675b0
zac2e666a227e24b1eeabbeeb4374a06d68bd2ee618d929e7611a29f833e86863da7d327452b6fb
z6fb84ed9093cba3a89ed8c8ef88dc05759a313808852ba11199ee0b015c50e6749602d0fc642ea
z865752cc1835d383d6b651660ea4e177682334497d7d996c55691780a5d86c831d4200078c66f2
zabfd7e8b18914fe5f7b24f3d375261b5c101bfac9cb05a89abe0aa1f12e32dc3ca95488a7650b3
z2c381de77eac50cb6e9450273990c1e1707ebcd3174c3123fc6b69315171dae02396eebe50e560
z63f8f84d5db0de78995bb35aeb7c9cac27f4d9738d1cd7be2187a2b90c11c1823086fa487fc948
zcde5a4df4d85cfd76a9b7c077585786eb6b8e1f02a02755dbcebe40f448e85dd9433bbda692b09
z6a73f459b87a5ff54e7f7f76c128926c77c30b88c80e5e1519994d772803f6b99d483f1accae2e
z5a004a3cfe1d0a4d9b126c0a02b6478df752c30e33cf2de893fa9e1dfce4ca2fbec8f6c80b96e5
z0cdcd1c1f2a153689ec80e635dd65061aef09ae7fd7d28123c90d5a6a167f8afbee4b41e034103
zdd19b50f933c36eaeafc5d65928b24b2c92c44c896e6336f9fe3f9ea092107dff5049f0e4f83ee
zd7011f035753998eb739b2e7bd11e067c58e6be9a229c47b3729f5fe359b874a20d94ae1ef4c15
z79d1124eadf8a647daf0efd51ac78b386ec4709dcd45d78c538177b4ef21b2de4061096046438a
z9843b161b31083acdcfad5ac7c7c71a27ab60e80de741018ea72c77e84563ed0a1f4db65d1d248
z577373d21ef37f8c1e2bbed448b864c1d7a7879e9a0805bbc9a024415b190d6705a3c2e01699df
z6f74c50fdbca0b1347e280d319f684a2f2d408fe1b47aada7461e2ef50f87831c3fabf962cc708
ze6886f4756f94ebf68949bd014ddb12113896d6f16a95ebe03f79a70def4a4b0e0d4f3b7c3b89a
z6c8063653b78fe4d7ef30aafc5e2cc87669a7d8fa89fb107b737c992c3f8380ec705955059354b
z2eceaf4f49e9a2d8fca4a534c0029fe6b4ed3d058403b4c103b848d8b9c7daa3c16399b140d4dd
za7faf9bbc3720b3cb8fbf2bd032e7e84729a5c6b55ecbff1028d33bb58920a31e3cf01509ac17c
zfaa1a72a84813f4e9967b9837c238c522c725ebfbeb1177ecc9af43172b6aff5c2f8527a8ff733
z89bf9c9f37c6051d355ca18d17e0365327ef1ccea02616d5c41060b390b446cc6d73a846d72790
z821b733f791782e7509e1a4cd4b300149587a6b6e45f5da1587f1595654426af097dc982dd73bd
z96fef07383e197fece46f13bbb08eaf0a3eaad3ad75036f3df9cc39436e5d868eee0d270971fc0
z6bdcfefa909252da17a6834c60d5f47cd16cd584e7d16970f5fb0ccc10792cc564ed5da1d24e04
z753a4b62c83cabab1190cc10e33da577b86ccc7b5cbc2ba4d2e8a043e0f4dc3441db6b7f869760
z9fc24af4ca3be86dec7d582b78fd36f2ae0d0f7507e38c1b76a65c658fa845dd065e37a0d53c24
z16892181f7883c9220c19a7bb539a17c3fa8076005f8838049ea76c61a9186dcb298add0516b4f
z4f544297030518988fd6702419411ca92875c2213aad15a78948157ab6f7d14876799dc07c365d
z0a425d32c39acf76322599a71d35ac972816ff7ed529732ce1f358904a7c0830d173f42643ef00
zc974aa2c0e3cc1b73788acde4742ccb13ba94d44ad9cd330f39dff36f97d1a9f5d1fed77a10e4b
z351455bb05908dda0fba611838cc1b970d6d089393891710f79bef73051c153230ec64420e036d
zab8d7dc1e8e1c2156a9b22dba1268593ad5a06bc2980b6d29842a0defa28324e6b40a3f08ab25f
z8b97b1e98edeeb730492ee13eeb8ef6fa4b1fdee69e2267b120a047208a99e59449f6de389f2a6
zb8b8241fa2fe0b01c441588ba9902aa40a795fbe6c9aa97acdf761e491c99eeb98088a052a88d8
z4eeba70faff0fa26803c01beed738d06ebad8034b44ec23bce117a44ba3e91a03307c56c611ebd
z07f461ffe9a7832659d6955a601b2f2d6d9f1ddaf7198cd04bbcfc275fa55e4158fc5d41e24498
z893d11347d085ddb68f26285a963245453f03396b13400785f38a669bbfeb315a5557d0b63bc31
z77517fb470b2b3d0f7c2f6277592319d511dfc02befe4141e6a6d0c60cf833c198e909d4d96e27
z5d3c1e394167bb3689c6e116238f166229fc39a3dbbf9c6edefb7442a23de3debbb482b458fd0c
z40c856508c1923515d6baeccdde53be56db5391cfcace25753fe1b00ce05407cc213b6e80ec0d7
z5cbeb1a312b7f616c786d93df8d7100d9c8e1ebb807c1b557a2b10a1c53f8526a0a2d64da9de90
z3faf0f5191ba5919209d6f01d463fae5af47b1a16285d94dea6301ccb787dabc3ff9b0c5a583a2
zf6883cf84f3bf58c9702a381590ce193a2c94cee4de6e91a6d40cc8d85f3401ff8aa50925149f9
ze929cd27d46797797164405a11dc1391b99a4dcfe6b4728ba55be65f67e8cb74e6f79935cd2391
z960610967102b93485f3c2673bd38601e37cb234b1566605882249575c8edb2c4365425409ebe2
z6f0fc3a4948d067a9b361f4b995b1845923776621e0a87a96841244b3155561cb1f428ed5e086d
z610f21e35bc1ec25a0e9a4a0feebb6804074452958c2eaf7a36e5baa8bc3a5e097d2f3aa76bf33
zeb7689a99b0e3fecbcf3ace1f243c2fb931fb215132aae806bac17b5452a5079a6a498edd2b17c
ze01c983655e650d337e84dc9d40d148606aa9d9ed1e70e8d76d31ddd9eef967f28b66431c385a9
ze6e737cf480e4531f07549fe8433cdb0dfb6390c9ec1e9a64e6767ccc27991f5225e4f2e5d1b12
zc8271b388aec8524da7cb1279ac3351048aec350b2cb79f9148b765d9f3916015aa1c30597fa8c
za6735a218c8191f4b0abe25959db494fa9ed5046c6b36d4e89340dcd223b2381c799ad91207a92
zca44fff021fbb4a7230545d3ac79134cd3047262f13097ef9c53e887d02bf8b37ec33a80c4a025
z5561d160f173f3d3435e187c30daa34c24b9bb01315c1c08a8d86dc17bc841dbab0d2f9ed6963b
zf13ed4a556cfc7d101efb097edea25c01703188188a4632aefd65297e28c0f52df9015af675f37
z4a4f29d8c4646a6cacd8842ae66c9abbf870b3c7bc6eaff9497ff838f6dfdfda94cea0c29e9375
z87ddf977c5185cd05c588c280a3caf30766d6b60831b86afa3440020b7f22138611cb69d8e3c6e
zd7721f1f7896a73656193392bd45fb18dd3e9a6375bfbb85e87b2dbd4dc69da69068737c5c5ec2
z575f6a0b4b82e6a952b234de5736e0acea22bf5fc9206ff439f55143adf1a56d89f2629a40318a
z0b48663aad1ab541a6676db23d5c54c5e19c176dcb272ec627ae0875a02322d0bfe80e202c1ca4
z0e9c1833a44730688a21fea644a8c4f1576b288bf76c93f91671743ed4604a39f6b94b0ac6ca59
z2c42ffd0dd292083163817c0ef661ea67e148995c51a702069c8d19478f99154656f54618395cf
z229721626482fc7e33a9ab381c1f7b49ba4fc6894c96625f806a075051d58336ff81894a968a67
zcd99b0bda81ba6c42a88b558cb23b4bf167cb4a036e6c207aa50b62b5585f2c5563e8f757814b1
z69401ee24b8fe6ee196b4b6ed7de9702280051edd85450471a443f30b31189d7020a0768bcaaf3
z6c35a315b1eb3790fc25a4b3801f4a30120b1023dae41a4c62ee2840cc105548157ca52991c2a4
zabcc9c429f29d0a05a4e50857a6a074558ef741872a298fd29e7900370dc5c5683fa045e3d0056
z663ed1248e85db957b9853e8bd346a6322b887b5651fe6e29e4d15dc2be3a77f13286705f63486
z3ed0b1b09146132ee3336c03a698bc455607b56b759de695ddc6be7fbda886fc88a50b1170b136
z1a8b47496a684fb62a9f61c90bb7d201ab89f63b3e8e34c83f11f8308b9b75230fd48ddc7f8f80
zd13543dfe3cc9a7e3798fb39fcb109866a3580a33001b51850f7c0f0f9e9b4241a815f5aeb15f7
zb83722763a6f7b055225768822e6a04ea0146af721cd4169656f4093b70a6387f0706d481a39a3
zee9ab0a6826fe3e0b369005822c6f682f9c206b047e57899f7b6d4dab386516e6d08d65d9b5a62
z36b95f4b48c2d5b6b704ac96d36d5c89bfc2a454f584a1ff4fc22c98561d5020cae4f51cd78459
zb9dc73dde130df896eaece2f946c72dd8575f4ca950eac1581914acbcf833adbd101015f9e3060
zf78e555433df965eb6f920b32dbfa29dbc74870019113293a394c809c4022d4fedace259b7fee4
zea0f6307fa9ee5d2280664ea9e1da2f2fd8c3ec367141c35b9e77167fd1484433e74675ab2f498
z03c957d89ea0e900baeb8506feae6e75bfc1b65c8a823e7ad170a650c058200438e177e717b0f4
z58881f4fde464d3108b1632946fc86dc095485229e90fd7b2f8780f85039f5953bc3b3a111cc3c
zc7d43031f3ee3960f6c8655ee4ba8af0b8a38c0a6b19bde8101d2a82a556be8df1f43024551228
zee059bb453164efe0f18eae597940278ca54fe43db5c6702637c659d4feb2dc261fbb650a3c3e8
zf33f94440ec998116f1e0830848bd256e00775a22b132a015bd892d9bfef45966cd88b1541b178
zf73a3ae8ce532936cda27ba7b0226c8c607927072bf29c4bff2aadf6205364a89b33a579d666dc
z5f55a9581028d69e58e48855901e96341b47a51234bd5d96b1ae8c33b0048d4b355ea57ccd632f
ze9c099ed53d5f2bcb5bfbbd037b9308bc3004fbc407bfa6af13ef88038091f2ba990f16d903079
z8cfdcc6dfa1b938411f10427fc22b4c871f326ac2bfd7f2426857ff597ee38b86455b7977ac1bd
zd9b746b35527d4b502f001713de4edb8126453cc67585bef742145a1d2c45d5719c4a03b319847
zc6fce9de7a9b78904cf58a06735650369b1b784bac2a3260556c8b6038b10253b2a39761d8865d
z813e7c451b1b1b167577aceefcccda88b77f65c4e4936e6daa7702fbd7692f50d0fac6b82175e7
zb3fe0987ba8f63793e37e296d0cf1d1b8d6de876730e54557893a12b9af0c01803a42f94c6cfc5
z27cf6b738e035c09fd03ba1c8e457c3e6dd185bd553d19fbaa19a46dca60c81cc1438b3ee9f7f9
zb6039f0ae7ce7ff44b53bb6f276f77fcf90378d5d1eff057371b9d8519b87f9a0e822d286a61f8
z34db31f46f8ac069e510f25cd5155915be081e9633af37357d0861b33fabb39bd94dc60e014639
za81ec2d140902994d94bd71714f774b59a49b26e07e257f9b60a20d70c1132ec7c17c45bab5865
z5343ad2c704a1c8aa3dc53f9208dd5b7171ebcff388a1b1cf3a6d6e815ed27f75ccb21e4a6de42
z0928c1c4004aceda1e278a67fa8c6107af172db25b3bb2bb909c12852b2e1f45aa0a2ca2ddf51d
z0634045931f1dcc783d596f3e341297fba0d24f2018aae3d0ac698454c0ba5cad2fec356f2d030
zdef5c4f4cb672865faf5b4b6fc2ff816b69cad57edfe5e764b499ef9f1907012afba052386d0f2
z23f02cb6b0c0e4f97f643ece6154ac90ea8783fb0bc6da871e6faff17a6ff36a64ce6b4937ad5c
z74bb397f025b83abed397e82d64ed5ff1ffdbbada6b757ae2a3a9160f28f7ef4633e587383a46f
z672e95480ab7453caaa51099921adb6900e4433548e3e0c2f61ad52866d998a4184b7465db8b36
z93c7f059780b618bc428cbef3f24d2c4a6e3cedc78c7ae738ebb884b498a0be233cdc509fd8bf9
z8ded0d1155cd3da686c5c89951d375fb0125fa119e6560a9e62025e64bbef6e35a06f0f8f4c568
zd8b6762fe01438e973a0cb3462af241eb46524242a24ba9d18005ebc08abf78f414d451dcb032b
zc8f5467643f581c6373a3d81af29b48466d67bd8a695595d0222425292cacd061d57e5877f953a
zb7e5f22fee3e8701b06fa857eda062e694568043d97ddf6fbaab0687731ca6a9aefc84eced9a10
zeb9f307fffa10647ab4f150b9e208f3087b0300deae2864939d59d3354419b2b8be0091f4c1f9a
z1b0209df41881831206202c4bac3542e96dfe6e25a5afe2a79ea31ec22b62619d78fa50daeccba
z8e062da0e9efcfbe8e909671c04a0522b080e65d2deac8d9704b5895cd3135b7abad5594d47735
z0265ba07d99e8a9bc106afd701ce1ed9110b0d7f0d062783a03cb497292ddda0101d674c7abe1e
zcad67c1d42f92a3238255951ceb79abc2b5bdea6db75345ce5782edcf0e7006f520370e671eaaf
z77b1bc6fbd2de8b34f9f3d627b4c172e5448fcb8eb25c2538b2bd7a65b48b4e2be9ef38ed3415b
z7d059e94a6449d1a471bc5bd96c217f6697d5482cf3956d0d8308f529888a54a261fec12c3d526
z5314c9b63d75380086698605f63151d26b26a63b918175e964fb96792a1949b20a1922914ff1e6
zea0e3277a5e4e9bd4ea3d23b7013269ce4c0fe091e85748bb283b83a62d89045f5ee4cf8cfa197
z5c99894a425a3d47ae00d0b9059da251b0c4579042471c0a54bde7e42838bb68f5346a7a6f79c7
z955526973803971d59ea186c05fffd98d7628fffc1917e5a7158320dfe571c4cfae38359684b8c
z8d69d76a2fe91ced891747fa90e4bca52105ecadbee14bee1ee89d59c383c0ca4f3c6d46422033
zc1a8cc241cdad7ff427edc4f205ddc4d9fabe85f12e03ce36cd6be3fb8445b577a40f3e1977b2f
z080548a8a1b97a58f55dff2fddbc0aa5c15b4e4d106074d6ea5a1b8b6c6917b8f035d72d30168f
z217cb6fe7ed26fc1ee00f5733d4555b782e2d2b9c410628bc19f9eeeb3a970853508158fe307f2
z313b657de3ee8786c48ce27b721f79015a2f866c7f92851b15c7fcc65cfcfd55e955d1ed53041f
za8027784ab93f2c8c5f73c815742ff306fa5dfa4238fe3ffff94374768e72e78512d4d7f5f0280
zde686994cace3b0568bf724210dfb7cc05f7ddb5728798638ab41621953fc1d89e88819f264e62
z6e3e7d98f9c410ee6f5797f5f3da09ec40a39850d4c5776d7039e3e226c0c366c9a5a0241e1378
z81889c7462fe7a4ec8e4a63d932be143ec93409e8729100cf0b3b8a0c13a55bc47051895b841b5
zab0cbe8edf46df637ce209f4911fac4e40154ae8573c70ff09d7a1a98d671f75e69d3abc6aa432
z4d3a753100bc497cc2befe4b5d9f2d8d4157b320256094d01df768135effd0e6275cad254ee8b9
zb7bd57a038a1102b97609b65d4edd0a4ac8dbf8d6068079028da50a005913e58e957d62e8efff9
z905cbca146423e059db33944c2b71bd0afca907d82f8b4fb7f60d8f86edd8a833040ba7f483c27
ze2d6b4954e5a0a8d26f7c2fd3f6413258ba0ad029c2da17600dac28133164803e588e2664d3fcf
z6448b8d8dc2c7cbd4e4fd84650a4fb749c3cf9c62361006be28f8312bfb71b4cfed093ba54d317
za68d9fe06351097fcbf9d73acc79687577361214e8c226e19f9d32e79954bfa0d6d0a53e393f65
za1d3b3e99ed39a6fe6e9772087f1df7f76974163a1463088492ae4183156ec9617e760ef4ad1ad
zab15bceb0153b3992868428f188a06ab7393c355f313f9e2ef2a5d9aa3ca20e109871bd16fbdf0
zfd1313ca239aea175663165311d6e4660494c695aa611c267703a3d873883416a38dbddd675919
z039f5bd489be02af6e9a36de9236920e9d988eb5767ff66b5a2a803edd116ae9090487a0cd8021
z11e7b831a60d55bef0795cda3e1647823d830583e6133b0df965904fcb4504792b88f1fb1e5abc
z4c6ade3280281a63fe97b1b49a4cbb326a514f1386731c70580cc44d0a0281428698b06465cdc4
zeadb170876c6d86a957e491da868419a27a5a2eec43f3effb2733a78c0fdd83461a5ea9418d417
z873563f28d12c3ea644ebb98f627f7ebbddea44cf35eae354c7bc5b9c5fca266d5654b7c30b423
zc114131a8370bb9392102980f4a5b37baa639838ab2b58117085f0d024ed55385b5e6a65ed5a95
z0146bedccc90ba09be7ca836ea1554d897dd4d324fee0fa13ab788db41771518333c389428a0a2
zc96f9737a739f3243f1edf70c461cb266166f9372c607f893b3f18da00fca9151fea1ea6bb2ec9
zb7bc7c2b24b7d95e834395adaef43b7f5ea298dddbd696343c0f5c575c44d6b0e4d4469e3f326e
z0087bc6106b9b5c084c12ebbabe8207d7083268a990d39afe9616f7526c8937b7e7a989ac69463
zc0773ba4c9c82b2b69094a70c38a48e72df14774a78a68536eac0d82cef20fab2932621b5e98b5
zdc63c17d15a2a3c5dfdde03d9eea13b23f401e359802222410088535f7e8708ac84710e45b5a70
z7e527d8400c1d87f1a591e460459cd5a5255f3ed7d8af0fe451a9adddf2e68ea49d3e37ddc3c50
z8f360ec1d9da9d101690a668a0adea2fc3f4e7af97febf8acd5248ec905e228b9648468cdb8bd2
z9d2a5e0913de665cf0b22974033fb60b405242fe39f3032c66c3034e53ad258400ea57e713759c
z12bcb30a342db51e5f72653be13199f5e158a28b1c308f6d03bb6e603d6705ed8965b4340cbf2d
za8cf85b515784a6539bd408cfef7e9d05e57882ff523d30d03c7d744b784af3050d39791432753
zd4780f1bdd5667001f7c332db01fe45c4885bccb254f33905d304098b266497858c665cd77816b
z61a97eafa389267b49c7c2a4ecbcb63232c5cd931888450a0ffde761aeab6f9edfba98fa39b40e
z0218f0996dddbd2d27a3c2c0e0339fbd741a61ad23be4bc8dc413e5ce1c1e9af41216bea30ce2f
z1c0a8f6b25742b5123c4d6bbc6a905c78bc938144d12f7fde5c025cc17be148199f9438b30f701
z635a44c01cd41e04b3d77726c1140ed7feedcb719c3e9c30a7426066ca9b2c799ac0ceeb2d3ea0
z8209366c34a3e1e2f484686fd57f02b9f30361e24e2aa2bb4297806a6c8d68df2ff7f7552dcbc2
z41839363e63db529fd442d9dd36f223b8f20d7c7b0cbee047751637a84fb586d9930036c4fa036
zb99dbd2da56e101131d825957d9e7859ce78eff9a88b1e0bf34592026324a017e01f61b9714062
z0d88e62ee00f896c083b2d7ae7cabd47a60af45b546c809e967b5283e28a0acfdd642a9633327a
z4900f81da9d3340c087926008b25939915a8fd73f5208c5d521f326907161cc40e01d3fc1761e7
za21db5871a6e20eba4eda05489d52535539c2e8c5a22d536a91f9d3121b7e9018d8758c870310c
zb298029910bada94a8a71a3e3dbd4d6efe0a14555a88b100be45daf1b18d88e0f979bda571e5a5
zfbd2ca0f2aa3ecc0aab77409fe6e97beca645e582e7c3241acb956afa7cfc985fb58c4cdb41107
zcf54d4c1a0175e7997ca8f844c874726bc60eaf98b4003c5a9f72a8a2fbd6818ad2d41493bc7a2
zdff45f5ae516d9e4e1d5ff0d0d6434b190ea9b0fe419d2ed89343f2cff60b3df2eadaad51c3323
zcffe719dc85d9f09548bba143962ca207ec52ff6763b7b160f7ece2fadd0eabaebf805c1a26282
z96be54d4f98aadfc924b58b0b9fba3e662300d5ac071a801a1a8821470255ee91dca0d4a878797
zfc1a2c5c46e262082317bafb426c2e3341166c89d628c7b1783f0f54e8cd0273e631b9c4e88ba6
z2e12c10301630e7fae34a641558fec8426e9566be2dff23083af9283ac86c2d241d6d0da83d75b
zf3dfb9b14be7c7f81a4494fa61eb7f2259ebd6e75fe73d0faa5f14313fce0bd6b7ae09a053d9dc
za6b99bb59a60c15ea72083a6c873229f37f7634880e9714f5411c7a8cc866b5ae81be2d7ea140c
z3a0c504a6476f6cf6552efd141ed2200b7f25dd9949f1dac91e52a2c7b9df4070120b7b07a48f5
z28ebe92cbc99310f1967cf439f60c1b07b15c06132ecc21188b30693471266ad6de6ce2982d814
zd1d640a3a3b5f03e868929eefd018c7b440fa1d9a1d18b69fdd3d0d13eafd4430c30827bf6d02a
z96333ea461b4eff56528ab98876534c3fa0fce22f9b94da0eaf57b8ae7e4d37d2e5f340ff05652
z2f591958a6732a77497cc0adcec09941f1587597745e44008d3b37b79df235f38a480efaa201dd
z19dcbe836b945ec5312d3802c42641ab3e72c1a3c9eef8aa4d69f0eb5bd731f5da82aebaa6222c
z4743eeb5870962ab15de744c5f58d081d361a9e6696d0630e648b76fa0478dd0e0f06af1523127
z078328689eb1f090659dfd729b117ec4e6b0cac791873329b41ad6eb60755de1b7740f13dd580f
z12ce3a9712666076c2df99be2e64c218698189b4fb42b19515881c3d3760cd771fc5008a10c9fd
z08c67b8481c21357db84ddbfd7e2428a66472dae4ad0e2316585a8a7d63e0847c3a6c50845f357
z7981227adae17d7bec5c3241a85e152d884fe1336fe01de4da677fddf19ad9197ba910594a4b8c
zb24396f0d888e55eb10c6249357c93399fb78d5ec717ecd9e06a3c2a8562da2f4c574df467f0d6
z4b16c04146aa802f495bfa98b439b9bad5df10251e0775fbf2a5822087ceee62a0e877eeba7c73
z4afb51aa1a9c82ab00416a52d14fa88ed9a25d16b7a0bb03685d3ccd43cb84a887fea7615d4576
z3ed5a0f68f5dfe34c12317549ecc903a7e13f0788faa294c63f7d6336341ae0c52695a68f9c2eb
z10da719cdb35be3487893b986358d46fe47a87f9c3c6d49ee691a0008c1ad199b8e8bba2014f68
zface643e5643a575f34266534f69ea6ab5aaea59edd1cb6483069a0451676ccc18ce0cb8552780
z5640c30d24a9a071ff80ba3d495f4e6d163ec80f6cca08f9aeacaacdeb2643caa4625bed52c397
z2dd297b9f25bba99f9c9975dc436c336f0270ada5fca5e84dffe74900c307ab3938ec178ed5195
z22f77c1249c02622afbeca4de0717828eee8d40736916528f747cfa1c791d185312554d7528198
z31195b9910e81d0d9437c507f6cb664ab3b6e6ff82293e41c768dd7d673970d1fec115462b1624
z52292291fe9b1f04f1b1b1f50f8f9f361f272c68ee8bf0cbc76ff238a65b0e069d5535fc383334
z03a494dd87d9fc8460ddec3b18b67b9cea654526c190bb7b08681569204401b4f4f6873919f95c
z81c184b4a71caef62039ab8091d5cdaf14401c1d041d39cfede366d6e976246362d5156e9b4321
zffc6aa790d7cc432237e560b95f717a855a531d7ac49a07809466194abf8af67b0b0bfc27e98bf
zfcc22b23339247b173c1b728b0bbab922ce7ef4db146f338742448ba1cae9305052afba69cf743
z35d820250ddf1de3292543ca1c458f6cf8e0bcfa1655763474b38ecdda86a54a3382b353897c3a
zd967d557e6cebfbef8c49855d2e98e4e80886ce02afa56c44b695d60bd50f9eb547576d51d589b
z499006f9075e0a60e6408e09cdb5649a3194fed1b7ce27317ae868a4cc6f3e127098cac0b5aef2
zbf25bd2193e127292b26644e452b116d1ec258e7cdc938a4df18edbf4f78012b2be565581697fb
z21620c1f4d967a42d8ad58b8df78649a0939daec71a5a5ed76e457b698b7e965c97e3a06ab70bf
z309df32d0863e6fc910bdd24a6d25c84dbe600fceb75f29069a9022753af9e3e88098a4a0c5d64
z430cbf39a5cebf02064109a65c720f356238581ccb9f9d0759179bc373adc5327d227c813f0c23
z945899748dd8d821fe3c33068bc624fb1bd11394b35ad8e0f0fc19e130eb6d5fbf16facc55aabc
z7aef36ceffecff1f2160cba5d86c184858b3dd90a227c70072f7d5352098232ecbbd012e99f6b0
z65f362c2b5aaa6dabb2e84c4c89a5a3873ea896fe119dc67da9dd27322c3380a668547f65d76d9
z7a39fdf8bb8fc5f27ae1030abc68b2ef2649e37b60a7a854725a1c4707aad403f9e8f340088ae1
zfa35715473f0e73b72d9c58715bfb237252828584618d9b4ab3398d9571d9e6c23e0b1d9b2b456
z9a7b969b9a41cb6df7426096f0743929ade8358640184c4aea16222c22bbb09d65acd292447e09
zf84c827e9d65850fb2f095cef325fd9f8b965131713ef223306986c098e0c0eafa147c352dfae6
z323c57a1c71bf8581eafdac1cace97b67139ac94bd059435724b7ce50bab185ee9017edd1d912c
zfc2aba6c9a9b167e5dd157d18aed2efd2bae3012b75b2a565d3bdc0f775e83ae23695fb6a8efac
zd5c4b98ca5f4f9dc1ad7ced1a94e8dc8163f48317dfd252cfa6507cbb23026553f9533ede91b59
zc89d1c2b18b160bf889c5b83d51663d2fcecf3b3b1808d8107aa7d8ef27ffb7a2f9cd25a4f5db6
za45be877b71eca6ff5fb221690de2bfc00c5815e292edc11efb5f0677a412876a2a21f2142e4e7
z64fc1ff622e2d504978dbe15206a692169d28c8ad7fc2c921eba552b46524746703d2dc0fbeeb8
z3c7aa686093cd70cde004e9de4fabb19871e679edb1b9e1ca973947a33f3703e233fbd63180130
z2a797838474eb4f6905aad4ea3f0ee18f0c1b842a0051982e7756f85eda01fd469778fec93e536
z44b6d1880df89774f6d2256d72b85f372f0a789728d4453ca424ec61bbc6025c74c15984f4edb0
z87b6a6003b333ecfb9d9a4a39be4b40b903b20e0f09da2d4193e435be4c901a07932ad23b508ce
z9772f065546c22c5d994168b83d747bf614e56304c2e44968acb0c8045f688d5f6fe5661f22573
zade1e2218d1bbc62fb6084749d9697f22e06ce531b43e21dcfc818f7a20d582dfa26353894fbf0
zdc990461b6ec7cbf5c7c462627b6fb37398dca689e0535c8cfb3a94e2c97e9e1b7946a3d88a4bf
zfa45c4dfa2042daaa19af6ffe67b22fa4fff68eda2e36228ea22af83defae6be70fe0251051bf5
zd9b9d60e6e30840e2bde252df6873b730360a8753b93f32992e8b14f7aea06b439dca4697bff15
zef7334c25ee9bb4d13f92acf0a30c5f3595d81c78f4a2b97341b2016daba70007c8542353b804f
zb521310d0bbf0cf099883af5aa3b781dd2cc67d48951ceb3053c3890325c10b28993b20fa33d38
z6e5f314f7239b513ea7ea9d4b86078eac5ef7ddffbc4176247d86c68e87001af7e6c7d70e35b85
zb98b50b55bdcea2e6cb9a96dfda18ba520f27ab2f815aecb46c0e6f558e0a4cd26275f134bae43
zd53998074e6450610055304e6e0c6abc7b4a93c95171f92f103f5abcbe18814577813aacd07a21
z86d6e5bf0d8e4878b00184e4ba4e35070c14bf35301e81c327fb29b339232d9827df6be460a10a
z8d5cc97514de363f0ec5b4455da717dce0909905253a51a811d3dfa46e3a6fdc889e6d3bb55196
z3c84521ebd65c812bf72b9eac8b6e1ee21ba0335cdb1b8e917de66747e66b9c30103602be87414
z3cdada4b607cbb8c34bbff171147e7ebea6ccf4b26a4069601e0
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_assert_leader_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
