module input_register (...);
// TODO: Implement input register
endmodule