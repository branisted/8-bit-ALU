library verilog;
use verilog.vl_types.all;
entity std is
end std;
