`ifdef encrypted_0in
`protected_0in
z5e29c48b5864efae434ba8ed3b027973743e6ee284f2e9e4887338beea9244838048c3ef148ee0
zd71209dc15fdbe94e72dc2b9729ede6932df02386cfb6f6b8d16882833fb31f882f74f44ca09ce
zb21181fb150f4df095a9b152a8b7d0e6050ce1f87567dd26fa41ae90cc25916261330c143e532b
z61513d6d323a954b3a7ddd18eea81fbaeb5bcbbc1cd754c2cb582d52ed576f41c1a0f5fbe7b6a2
z82c9956c43fc3b0a2c0bd525d1467b5b98131917eeca4ad2dd2710c39c7443efe20eede7a35964
zbbc0a2d4ecbe8334e4cfeb86c593b2f278ee96fa199bc37a1281a3656ffbfd8c65232cfa9a2545
zcd26e87631d1b7fd32de9943e644fc16b2109ebaf98f06095b784d966c0f7a9f9fc2c58ff55d06
z7b7bd426862c7e7ca485ac0333b6fad42cf22e526efa1b688e9f721fc0bc8f664ac41ac716d862
z4fe59ab515360b39e0c1fc893460279f41cf0ac8d175d526acbee633a44385d0bcb13fbd5b8e1a
z23d0add266692d82fa87de0ab1854843a9d9266ff244bd30a2395d9dedf23b712ded46fcb2a92b
zbca0488549bca0cc9ed701de26b0a758d8edcd4d98fa35682d21895d5e95ad40dcb6d715deb119
z4b82fece2affd9bdf718a302ec42d14327a33a81aee03fa7472fb87f2d5c7339c2606fef317fe4
z3fb3fb3972d4ebd8a56d05d24632497bde4d22ca7f67708a54c2dc46da6f2d7d85982a33bc0357
zd8e0a0efaa37dd2dfc41b66b532860901f0c9222ad013223a778859909cc38752bfdd4d1479d68
z0ea3be643ae69fa7045028650df930772d81055c7b59a6bb54332c9be2e87a40693a533115679c
z70068ee560b5b2caa127932faf5c9775fe1b9706d6ae5033850aab8f64f49c03812fe844a31f9d
z5b7a1451b4be6b6401a832d24769d585177f104299ea8a6ce0e59c34ace77ff68c1cf91b10f250
zdb830d27ef30a1c9892e18bda8ffeadbf5aa92778c0d1bc105bc736a2b4a9b953d0c70d9172054
zd5960ff33151861d273e2539341d51a6b0b6f1c438ac1028588022de3300fbb812d952b4311e9e
zad16eb3c2ec1a7d29cb695719eddf3e11c462e30f3d76f12bbb097eee4bda2a53ab4658c41c61c
z4c5c7d232e6db59b78ddf28ea594eb2cd5b622ee6525fb7b282bcec34bf79d1765e3d283699c9e
zbf3e0ea8bad20fd2586a7bc8792982cd861ee9f47e2aaa94bebb0f02c3cfd327cf2a0d1c7208de
z11cdefeae3301b63fdf8427e6127c120ab189965a70a7663408ffbeebc731e3722627dc5134af0
z25fff0712e017bcf81ff3e96d40e90e457cedff27403865c2a641858649b9bf5e921f9a504593c
z237474dcfa2915e52defe6a6a5f04cf2e813835b5a7fe1046af147e0905a7fa375a84727276969
z7847ef42681397ab2efc1fb9e439e16527dd2eaa8dc1e9f14bed81940babdb7c2b7eaebf16f6f4
z39e82def89b0e7bafa802c0c1571a0d491958bafa2ec2bf9e9361340c6ae8ebc2b9e302b97dbf9
zc7ff3e1f55524b32ebdaa568e650f75eca6fcbaf7c2118a4b75e020de3c355d013641b58038c9b
z67abc102358a0e841e8719ead6f112c3fffbacd1ba5ff0205f4a6d35a0b66bbcb5fd4cfdba13ce
z0feb55bc1fb04e311d172367d62c9287b286f2bf5aeb4f3f43276261c0036f0f33c7ed3e0a9c5c
z86d95a1054592543e25aedf3fa554d0ae36326e6244c953c774c38c7360d738b5849d03480173e
z031329dee4c833300ed8ca4c3d1a88de702dfbccdb7f60336272ee5d25e0ea3a3d22ab8a06117c
z982eb0d18befc6c4795c46dc362e5e7948d583cbdb8e5a8fc1e66aae0ff1e53235aab7e60f638b
zc762dc27aa309a33cb499c989454a98ac20104b8a6aea7c0a40426d25afedc0d9c537c1e7dc467
z79c002452a4cc18e810fde30ee4209b407daeab5b5c025c47fc5cd99b9885b85d2624f2eca4cbe
zaaf498b098faa390bae97c3b35c188546acd8d6027a458b50c7a131d82984c50d51f4520617d12
z4f3aa9bea5fce4a525bc6ae28ca3a250332bed20bfbebc5d69818b3bf5d9ef5869b774e040ebc3
ze0a5ed34b4e3d3c670277815b5a7fc8bb0f962fabfcb3929f3c47d12022dcba0364a9710645d9c
z6b602639cdd3b8be6547249a1510100bc7d3f106130c990035f4bc3c69e85fab1c05d13f1894d1
z314b08b644925be2b3827da86ca2965cf0c668ce4e104f429698c9e4f6a576ed902215c8630688
zc75161c0735dfda28dc1f6a8de8c0a1f35468313db76840aaae2285535cbb3ec3c92a79d58c4cc
zc020397335f5c5f7004362f6efa7bb787be233daf3e04a211b6455a948e53873b3b4db446dee47
z0f7000fe671de286a7a9af12376b5c15e527f9a4937acd7bc1d5101f8c29174212686f1b1ba4d6
z7671794571aad411a0e15ec5c9f6fdf4aa88614adc74fba2201ad384b5ff9ffd9af7cdf6aff1ba
z1031ab232b2b75f60313971b31bf213eefaad8ad29b0b7e39efba7a67496d6b568fb2484c87139
zc1f20548b594a6f1a34057f1a106d93f215cf16403db20e2c94965e2ee18258d267eaf0d5a062e
z6a5487364d94012e9a4a9a716903347fc0317caa32c9dd47bd7e23f42838a2686055b6c6fc5c38
z5ed180ed44ea8eb8f611cca6c67ff41eba015cd3d42e6b51ba780e8baf880c6da4a3d5db2efd8a
z2022f775851cc04f8ff4101e4cabe4ed12d6f4b237a2bcbcb34dde99e0a4f992bbbdbf1088a64e
zca9d2cfb8e51e9716bc8fa0e6d6ea44b7a8dc9a09e5219538f124d85950d24609355e50da3c24b
z4bc1c6c3d56d613d1da6e1003588b3fa4f861afd798292db3ce7d0b29dfc01914fa477ed934c23
z697eb84b922e56960915ba82ad7c3db97f6281a3f30e378bf2feffd9d83dce046ca8f5778c7803
zd3953e31f94713d4470d50afe49a6fe511596968fc45354de3cce51b5550661207d035bac26197
z5af7def90dab3623b8268be42fd0b342de5b702f5907a17e740f454ca6519e09a7dc6e6d618450
z12d86ee7cce277c64addfe3472f9b3d1efb8e697775d244c593460efa9c1bd60d776d1ce820787
z932dba80870306a73a942d66ccc09f84cb8bff285ac8a5b88854e911781bf11250c18f62be2585
z567c82474a76529abcd4f1e156003a0287b7b2cbda1250d78958c04d0e4974dc68e8a13f5efec5
zb439b68a7251e53bfd7840784c5575c0a1f189b0d390b44741bdfac0aae9c13572ec8b0f6ed1b4
z53cd85223c6788f155ce1c610da32e753ac6e0738e4596e7bd92bc96774b9431e71d7c1672110b
zf37d81dbe1a8544921e1180d8a375872a86106df7107c8c42d2dd73788b080534b406c91f34a5a
zdf6e220a1c7780030b0acff7a104de80751bcb9dd452aa92e466c943ffc7b30b988ace8f9bc515
z5dfeaaa9763f4c82c5118310ae2e3d6f8d542eb5dbd683d2ace1a66632ea97c1a0244aa7141be4
zbaf4d44f557dd43aa3cafa61bf029802418d0a310c83acb414bfb7722056e6398c1b389030472d
z68b1639cc11bfe4d6e56ea1e71badc4f0015caed1901beae1ac3bbae3aaa4ec4b3b850d2eff69e
zf17881981aad58418dc03b6a9f301d370505ff9b5daba9a43595e467fda26f482c5c91108156db
z62a521862885806f893167cdf9a17e8ddfcea25e85f5f5bfb4d169160418beba7a9c1480293aa4
z216f4b1c72a15cd982592af43cb5ee51781dcb7186baaac4d5bb4274be6db058a215796592a328
zbeca259a8a66533b98feb0a7249bd1ce7a0c1f190642b374afa4cec21d258b39119c508e21a922
zc07f6d64d6e59b9e88701f991934e9065e049a0afe161f2f1936b46a110d48d504bbb14ef76aaf
z7d5890e80e4f19bfd8d5a94ead0afdf38243074880b849c853fb6173c237ee2ca7e0c62dc6c409
z24fc05140e2b18bf4abfb1e6ce6615202a53f9454f040d57256e29fdcc81ef125039077bfa6634
za56874956407ac5f61f6b8a4a5c05656ee3ffec11cd395d70e103ce3eee03c5b62c09cfe05b70e
z5ddbc3bd26b94bd4a03275527945e0500ea995163e488db941b4af20cfa3e7e30897318ea2bdd8
z1ac9d1b9edbb5dbf29a228627a62afa7a2229f3dcf930586653cd1c5db8b52d185ec3b93e8ff92
z7ca89c33c13236007df0eb6c34d65cd1c2e668e69b52340faae7b5997768d63f70cf869502e668
z8e280cf5e7684b06df0c063788c1ca31768adcd05e7a59f68e1745039ce59b8e6bbcc321bad40b
z51c38b9af4ae5b68b5dda1075c4ac32dd2c99b6116e6e793f16f5bf462357c2d8299bcd8ace745
z6e2f071c45a13b9835ca4f485d84bb4a43e57282a91eaf0266b468a9c99cebe67f12b648e2e229
ze6a6d18cef7c58eb00f028b4ad9bbcff8b535923cf9876fd8c58dc731d63d20742568fd543d221
zdf237c67c4af4c681e7f60b00e20cadea863eced01960ab4b02f4b66bff6d912a047b429b78c8f
z787d2acc2d317edc240159e14512b8401f05d99536047d614bf8f812353c0725a4baaec750834d
z4e0d67acd57aaff0131ee006a65f745fa2a2ef4065eaa70cbafe43ef0a64042695c40be1c91251
z8da104b418db004a637aba7119a0c346bbd54d9baaaee033211ead445bb22f61dc782d77d7cec1
z1c3769649aa72756b722d75862b0b7b2b5c1869467abc21dceb10451a654cacfd3175a9503fbf0
zac3f3cacd44d46ae23a5130227da09c9fd863e2762ecb7ed1c258fe6d867d0dc72360dfd586ffe
z81e5407ea807d4bb7afbd45e1e8b3bca8e8678fb3fdd5b2ef296d2e462f97e3f15929527529056
z86eae611f8dacc4f7a0ef6df1978966f2951d77f345158bd1002e84f5f1d1a8903cc772fa08f37
zd3ae757e47523dfc1af61e3386cbc203c10b48d9bd305a5b977e4775fb53432de30ab5c7d5ff17
zf7db65f95cb7a47c632223ff99a276f4d5988589b89fef9abfef99a5f451eece93693fe013acca
ze3c68cf8402d14c8e6cfb92d24c2f5b91dec68513e2e2efc59a719648bd34dca2c5020d90c6813
z8b63fe138353d1d52d3818a30994fd4778e518e4c4d650d15574c0c867b9f5aca41fac25d4f93e
z80f5c82e803dda17e15b847dc89a8f8cc7d7e0cb88fb27b00dc00d0a75a927a8db299b270e2413
z3067bf4ec923ed5244d5cccee0dc6ef9b3fb052768f23d0b0478471004161fba29d280dc0980b6
z32c38dea7f1432ec70310b3bb1fd54aa7af091e30872176199de818bea01c91e5bc8ef207863d8
z3777dd10c427eebeeadc8e0971068c4d7a3ea6eb60e73710a091bec8288a23ea2f5b55d29b9735
z1cbed6e161751f1881c005da2a21196c827b188f021ef7a1e043a31cda92268a7871e48eee3d7f
z84c026b12a99662295b52afd7a5d3868b74fc4a47a7d480443fbba2caba377b6fd086deb934d63
z4b7a4e3085cd4fe19ceb8abe211354f72e8d782a43a0cb0a228e68d7b023f1bfc6eb94729fb9fb
z9a04b30fdba5d39bf944e59b8720c3d9a66ad294385e6ca171aada21cd98605e5c87327281aece
ze0e90bf44f957fbabfb35d9d71c7b52438011cf794a6ac77f52537645eb2e819f0b56eeae22225
z1c263fb1bb44257e68ee6adcef3fbe98c58095e55ad2777800b9ed8a087d58e2748dcfc2759fa2
z7b001aab9b15949d9cc8eb6c24ab53c56dd48a6382fc94783f60ec0408996501df2e2acc1c13a9
z20a25a6223592cbdec9c5826662061ce634f76f8295ee63603fdd4315f41151822d52a437b2cb7
z1c865343d6ba0e5c0893c281a549ff4c38cc546f5ad1207b04fb828d4739ae1e01e80f262e6abf
z2ec331075b3bf1afa1c306453f8a5d2641ae3dc7d5e1ad28b79163346fdfde6864a7cc7ecde441
z672224d04665dc9f1a1d20b00eea9c8b3de1a41e134b52d259fd7c1f3a1af5c978a978037be234
zddf9d52001c1d757e70c25c30566facb159cec47dfbaf5bc604e328539cb2aead9d4fc9719aee1
z44f9bc3d4ae02e4296286819341b2c39d06a185f7cc8f35f74db255324f415a4902b32e0fb7174
z6d6534dc2d53a10c83ac1eaefa0942d65408c4803492a62d8ee08155ccb7ed420fb91a5c229826
zffe4599a051b8e2711339c57996faa9263769013b19e8c187d647d789fcc6ce62710e15ed5cf84
za70bf9d383002982e91af014a766957a92a459093b0b29c7af32cc3e7ad0ec08bbe51b77c19957
zc5741d15728a974bef606af39a5cb80bd8ae68c2df1cd03b86516d385277e4f554d14806822674
zb33f79e99a36bdace0996c35f11d69ccc6b85b40c59eea6ae0c187e0f068214aa37e79719660a1
z68f4d3e6c8ae45b1421c0fe9660e176a68ec8a0f41ff0889d9a784a70a7180dca3f90a4177b75e
z25f0315213a28b89f7a7153075b9ea258add137114b70f50510073ab9e7a45a3e8ac629578cad5
z1e2cff8cc6d23b517774dd5e5c07830956f47668dc5a801868d93cfa34a15f3fb326986615d275
z37eaab43c89a36b8db5ff474c4169e4b1efa4607ec2f94d86b4c324f99d736d599db4bc72abee3
zaaa7a142df53af758898ba46752dae448ce338ecedbd0357d3c2b0a647a74894524b2b3b3e9c0c
z55536e147d60311db98cb1ae20d5ef815f05b32380e7de4bf19e5f7965a65b47547ea3d7118219
z78ad73cd4fba94e4791660c388188b6db3cd040c7cf5c0d83e0cda56ba7bd1b6afcbac93a91355
zccdfb324c2b6dd03e074d7aac2af0cf5b0b90f117319590942352a53c254818760998427ec440c
zf8673a5af4a1d6538fb4161b52fed7ce6d82a78e96fd16719f2672f1cad8d5d69a18aea7f8e750
z51606ca498d1b0b46edfa469abfaabc29df8d5c561ce1f97d3d2cb4e9b910ea65976a5ed3034c0
ze59f4b8fdbecda5bce22289db4cd48544fbe525118c9b3060fbef1538d129d81d53fad39f65594
z7ba3572936f8ed1fe06a78660c87e6ced44f33ce5548e46b05e548026023dd2b3f1d0de92f4b61
zaf94aa5a964169e6d518d2108db23edaf9e213469f87bf3a60b04ac7bb551a275ae9fb97b46f76
z5034d7e7a1e6e5092b585e4d51f64c3757f7dffb296b87726134ab8b1400639185af2b312c7060
z8b86ba6e46200c69e6d28090e2667f02f4677d9458b203fe9ebebb9e289242c4716a187de41622
z44c6ca1e127b573475471e38c407b2a5b4b72f12e7d0cd7b6393c2745d7b96769c972acadcbb75
zf335602ac23fb4d5495c15c407be8832642e407e8c617d94f08875b028ad3fe43eb818150bf04a
zb50a03b742d7b5dd3163ddc70e31e4a45622c19d6b1ad39c375d1ffd1fc1366fc84fa8666c1794
z2e90bb8f3524b16c542cd7d4418d7a35709d02e8726e39ae60feea70d70cdacadcc20ad45859d7
z4a2a6f86bcafe2e47ba9f73dd3ce1e0f019449c57edfc6be3c331f40d610776bf29465d46f010d
zad0a370e48357b5e8bd7ae2f98dae7845ea373a99aba65629c7412ee01d01da65cc0bd0654fbcd
zbe195cfb7fe4a8cd01e93b362156edb90e35194592122f328a381ace43a79c6fc7825f358f8e9a
z60841c3042a768e6c0e173b421df9754c86c6a9e6317446061e67601fca6b08951d86b6672429c
z0d61a391f70861b8043db1dd0cd200d08ffad439e846fa72aef30d921e500c7f94c7aca16da35a
z80fb003eacb8ca7d687c839ee60213e20a4131653cbdc58014b3bca00b58ea2f3bf353e82943de
z0091cb46b2d9aa4bcf075a7d42033b27085ece257a881a19ce73dc5090c31333898f787e7a6778
z2c7e091fafd071071f2a39c14bf81ab4e75b44a584e97147be673c48409f6ca76d457b960f0d74
z4e0e343733d3885fa1b2e129f934815afba141384e53b343fb4172650ea2ea5fca07bb40fc2d47
z25c162b906231238d241df8d12725b6d04d1b00dc1f71b198c08ed97da61e0615b148a92e52ba4
z8ed7e0df3c1e5e4dc05ce16e27637471e840dbdcac023cedb1b408c82f7ab24e730dbf66dac930
zb7b61b006435b765884cb7271628e5af11f4d95c320d0a0b1a238d5d3615d0ea22bcd2736bb9ef
zb2e70bd892079294e43c7df1ab18c7ab91bd94bb1b9638335a0e2d1a9f5f2743b7e82da818dc74
zaec9d8fde9725cdda89121ee6d809dfcc00a15b33e38852a86eda4b4712883bb5c74de47648850
z3281b751eadac3b14419d8aeea59c389542a35150cbb0eef521935a3a5c940f74f74d8fde95e6f
zc5445660434ddbd60d03118e9065947e0f9d380113927be6c6e7e171dc9a20fa5c4e3f26992a5b
z294db9a53326a5d1f4a6dc902083b12c612879503fdf04da0513a4fb78f16b162b4f4a422aa3df
z1e2ae9a98aa6311329132b6e7b89037884244da99dbfe5842812955dd6e885f0db2785c70488d8
z87af3a17b8c4416f195db537d50d4489c6dabfe35adf072359d7766f8e2a6d45c1bf3b59260e61
z507e4d3da5849e8756ce380c8a158d53ca8c9eb094cfef963df2203605fd0b3e6e9f50c29b5ea2
z4e0af60f84aca68ef37e0ecd8ecfc77d92690c2309345da96f480af4cdfd2faeed04893c871553
z20734f75eadc97263768477b78734c35cce4d3d1eab2c8a2f0508c234f6e93f563301c33540e60
zc36a6cabd771299c51f701efe195bf03247ee6c1c0065cb414abb53081bfef075766b436b49de4
z2a8fd88fcfb682491b4db2e7f4897fca4a1f210539e999919a41b88424f2ea70f8558c3a849586
zacad59b153d156daa8cc46192175c550b19b3d190f9342ef3917174edbee629f4da941c84b4c0c
za97cfebb2cb82b0ae86ceabfb292e786af866378d8bef1d120ebec9619d78377b94f2b42fe1d6a
z1d7b64c8cf02c08ceeebd6b82db2c3d6fe3509836013527a1906a231bd954f9b0fee7eaf97c5e7
z80b1a35133728669bc91a6ed2bb6d7a6d2f73eb7924370c29ad6b9b84c3697d9c283fc2da32128
z79d9cae8008f13454e93edbe281c180bd458bce12eb51de6661398ed425e9305ebbe95bc7e679d
z47f6a3f93650bc1ab07a5fdc26af07f39cc303fb47b4be952b89ee6bd7fe6f7369d66670732745
z40dd8e17f71ade3f076f4306b2002c54d67a29ee8ce44a232332199b049d22be362a39c3b302dc
zd85460fb1b3b246fc5286f82aa274ab86db7c9b39fa7e329ab467353442bfdf2705496bd46ebe5
z64ff9a6466c8537db8ab2ef62ebb6283be43646e43b5f0013472dc62e9946383bed99ede03d45e
ze13a84b071e534dbdb6da52f8df3648a2569f6f7cc0fc483f0aa5e9aa19f33042f2322bb2b56cf
z3f7eef23fab815bba122ff4c5f83b36ab92fa1aedb0e6eaea004fca4a9ec0fee0b37b7eb4f424a
z1ccb1be21d9cdb8e14c83f40cea781c4544bd0da5979b4fc2644c2a2e2cb33add8e1ecaac51620
z6ab5070da809281dde39f06a1df1a0afad649c3769762ec5f0fb545c58455f67f264dac6e03ed3
z1e3440a3c5ad40bdeb0a349aacd09102bb34850dd10dec805ba235067db6ee8eb85b69ffba98db
zebe03c74423c477ba51b210bb60678edcfcb8cd5fd25a65df54245589614a45085dbcf3e70ce9b
zf60d24a605cf31c13130467daf82548b36b8dea0b896126689bfc191406afc55632a6eb4a64101
z4e020f58e202ac98e1e08ea590f10131825a7abd24d9b944669a6524c95fd581daf110cd0a384b
z2dce96f4b7cbab17d4cd6a2a24344255b1bc5e44e5fcb24c1b5262a83be1e065bd59f399f10ace
z325df3a56c8d8bb95b26c80f43416b231856e7485dfe4b08b305409394e6b498aa33cc56575261
z4d2b660a43eb1a962bd10e92847d20415a265f574aa722ba9599c8f4491cdd75bfe2955dbc0761
z361f8769bce4d399f0ffdc3aff3218511671f986c692fbd9b7b398cb8eaa94f31086e365013444
z356c21ab2b6f24402d7fa03d899ddeaab462214608a9faa2b3cf209c5b308ae80dc631525bb958
z0241291a84b9b0379b1484e6c194040bd94e5cc5789bea9e922f4580d4056ffcde82f4b3c8f3ea
z042e3d50b90aa15d63d88e1cc636140688fffb795f1476cb97c32f5c637df0c903c2419cd9fcac
zea6adede6f406472de075e76bb8ec1152d69f3f99a7fca236c3a3883f0697715560ed36712ad57
z67c32e8a9ef77d1b5e08df5b892414c74aa26c2a9ecb9517962129238d38abca03b944d2da6af7
zbe298164292e756f8933e80fa2aff6ee1e82692f481d23b31da5820a26cae1eb9b761c5827efb7
zed712e61774d074eb3a647ad4a43f3a8e314d60cc49625ad42c17ed14ca6e9286aadcae7363633
z0654ef15603887bb7936d07c6d13671a089f6ecb9ee3e70db63527905efe01acc314db8b3072f5
za08e09bf43c70621f05580ce4c269dde0cf62506e787bfd6233fce1bca3e1895ab78ad2e3a081f
z0aa74003680d2d175db42c4e40a63298ce63e5ca2df8c2a0548382c594c64ce6530436be527591
z50e79bced748c35f97fce22530e79dd9e5866fb7d16d2184f24f2e605672a222f319f103ac59cc
z2f660286da2375cf3340461f3ebd495c0d23c3006054e8880f8acd1a06d479643bceca39e20e8d
z71d46d72aedaa599bd3c920524c07ed31b812f60b07eac761c5212ec7891e9ad389a84ba6cee97
zd77b62c1eba3646b65f43ad51dd847c37c16b7996d11439a1c9b6c59612d58b17de98b4040c32c
za13c9d5b3158a0ea0e796cac55ef5aa14ea90a38b2d85fdeb06e70acf6d0eec906758537e7abdf
zb5cbf399051b8629a77bf795d8f5a51d14f926a071898441c5ab3f131fded891b092dc2b45b51a
z097fcc308a82907ed4c04e0e1c8a5457e817bbe510eaacdae07f7111d2e77996f1b97f8764a69b
zc19add79e150cec4bb91d14f08289f76d1d644ccf64dfd37cdbe76b78b76d1459e33346732afdb
z247ef382f3e556c2af18db7160c6501410c27480dba8cbcd3557d3ab28cb0a0430a029a761cf02
zc03174d4385534e1abd99a4b41e9d2394d1132baadc0cb751ed2c14457cb602631251c829693d9
ze762eb4c6efdd8391760822f836c3fa6a5555382e29a4aec3dc2be6bb8ac86cb2d0404124aaaa3
z133fce000852bc37aa788e236b9a4819109ca35418636e2f198b69222cd909efcead78507237f7
zb56ac115b799dcc488cc5244d9ebfff01b6fbd1836a05e11df34f11eae229b59196a077c99ada0
z255c5ceb9bdafa9b114f066e5835e73bf1930618e7496e48100f6c930509b34ffbf09c2b037188
za34a7d953e5686ccd10325d08b74500e833e6d115474f24f7b2e19d204a22cbf74a20106512ad0
z96cdf96f302924885274b001249465213f4e0ae243a93f12c84fc67be3ec6d6cb7c365e9428a9a
zde06ed2d8e2fa5f7aaad6f3c675eb85fde37ebe04e5bfc2a175ba05e6231b3e9ea1de0ceb448e8
z7fdc97693a3162923b1502885b62107e953a6c4a4e152ebf7d0e3ff4025b83e0a1107fa91ccc57
z42546795fcf27129582213cf58f53e16411d223e5e5e7574183289570e78b8acecf88d6f0f849d
z267c6c0edb9dbf1eb37504646863e74be69f294d1d3c8453c455a0e37039c543c2ea588b5453c9
zba5400592af63482691c2caebfa66a3e21130a76dbcae8cd6348cb3d0cea3217cffe2f6b3547ef
z84a0c633ce31737a7da81a24c880b0559f416b33c7c862ea1cb20842ac47e3bc686a1ea6f196b2
zd0a9d32d370f7a88edf719a2a5024af444b3f5c5745d70a4c3f3e344cd320413822c0d7f04572a
z444945b85bbd6ba2e38ccaab1037b2f7435075e5bbba694b8a1193d877e2a278b1003c266243d8
zf5753e41cb8511a32f29bfc4840b3a158ae6dd7a626463055eb31de6f8ac3a8f89326c745ca8b4
z2062d6cec2567a237851993d56f09a7018a9c66893ac0fb4da633db4ea68f90c60f8177a1f0a0e
z022d44abe4268860996e5df06f7360da08f6550c99f08bcb5a5e57f2e01ee8b9758b20ecc52c5c
z0783a0abd8e8920c896f2932407513f874728f29a3b0c82a6645b3b8e38df0b2df05df476b60d2
zb920c62c60afa364b468b8091c23bb241d90117d2b4f1072abd9de5a0a9db5fb8ff15d20bec139
za47aac1e949f9c15dff6e3df3f32d81c07b09595f5577115bc8c50296fd8a7c3b4e69d77958451
zb8cc492e6abfe8f33902fb5201a05aee7c86cbc696714dc21ca0fa024913518f49fea72b2af89e
za60c0cddbd46cc3c449073c7b236d48edbca39d4835484cf6722e07deb237a193f40ab8552c6d9
z36aee2a2a95b7ae4edf266852a93f9c0c2984272e1e9dc512449b01665bfc8a015c7ace78ca85a
z970ed43dbdf5a30c19bd3bcbc4e299d0b605b48d15a87d068a70d73f21a0420354c36f88aaf323
z20927af45fa25bfa832bcd52f6cd535fa2c121ed901afe7e6c2c16223e154f337c73b97a4530c5
z309b4b7dedb244c5b612bf201dfc7afb37b99b4985d09969e3d9e0cf4fc181349ee44163e8917c
z9aa7b3faf6c7ff8e3ad3d22892269641a9f194f4f8e9822a1e64065b5926832a2aba017778df74
zc468257b257318abcf2f41a67f7314d015b45a95cd001caf7aaae81ce467100c9f6edf313cf023
zd9ecc8952cac89258e623c75bfe373f6ec4af204080a38443aa7542664e8b85b1424ba7572f9cf
z1348a1ff26223572ec769f78584bbaaeb456769e2b1d6daef5ffe294dc5f31df0676c0dbc17f34
zdff081a2491341e3adc183162e429f0ddc16c7930d5270b28369d89a811369d76dd8a3f86fa634
ze339741e17ce0d3aa405405e1ae4d2a95837e03229402e2e045e29636fb196a2723867b06600d7
zc9ee1964cd78805f7d60168862cea7ac9705f34445274941dd0684e554956df548c72d46c99265
z94e87e93d190999e46445286cbe5ed1be0ee47e31db639c2059733ec9ca0315e8613b97a5bd6ab
z1679f8e7af138f063a96548114a91462f1f7e2a473c11b09c91d32eedecfcdb8d4f1b15fbfa25e
z5ec8b79265951a4bf11e0f3c7c0aec7f559d62a2951660a4eacf4ac5b2eeba0964251fa18e1127
z08d488296e7aa69ad234ede9bd3511b64b7875c9cb6ca42d6ac7829410fb07c60e11ad69699e0c
z3a31c8babdf8b646ce3dadd86f474f783a500e98eab48b89ce29f92b610f17bbe6d5d83c354723
ze6a00dee5e107b61a574371141ea65769417d388c0173ee05f7104fa3f11d162959ffbe2009527
z195fe537ca9310d5b1f20afd3cde332c07e8be43bf4eca9b5c32a368c3b744fd476222bf8070f2
zfeba4cb19a1d94c0076ac917f1eef7ef724235375375d9ada16345e6fa1466d6434e582baabeb0
z7ce4a7ad8ac0da1a23d64485b7e2dbb6104d69a7c57172d37af320d74659646ecdfc9f30775470
zda0ef368dcdf7fff19beb15c7a3cd3d81dabdbc6b1b03823a734d14da202b2a6db0e77b4a9af7e
z6a5e0fbf54f633f19f91be1998b7e4e55a23c8e8a085f77d5ba36a2deee6e47db6ed47e4b05ed9
zc07a1147ecbc3181dc5ce0cd58b4b66b24764d7989969f0da5aa6378a4a8fab6221ad4e195ebc7
z94c094d077145c7d132d6e2ed260fed5ab512ea92e5ba18f5f58161f4e955ff5e058cad7205656
z3308c0541b0cbaabee1ad6b0a6bf0050a1a7e148fce08c17c1d71b6b31b7f271a26772b0f2edca
z5f8f5aecd49e74172c065af86d4deec77fb33baaf58da491cd8def48a2b37285951d73f0b7951d
z8dd3979b82135d4b971502a961a86ad29929f506dcca8753c502ca952913bcf09ef0219cabd656
z07b5004e9c6657600dad6507423342de40c0f28d1df561d7189bca8077d4025cb9d17ce7b3cfcd
zed3e6439a6b836c165ca3938376dcc3258cf72dd24d8083c1c8bd9b72f6b5f60856b53e047f273
zeb2dff2ba9f703788d14e9e0c1e3290fffa8f2b96c87acc448c6de74ad6bf4f3f218875a13f296
z3602d884b70b5003765a35bc044a419277bba07cb9d5398578dcbe2a7791239173c22d49ae99ef
z6e9417de9d70db8fb5725718028ecb8fa99c7c1dff59efbe8c89d8641b60f8c21d1e61965f479a
zb9b2e9bde2ced893a291e2a3f3d27a2e1161607ccff0d05fd9c166eefcb87cfadead6db2891654
zf2e69e1e4ff81152b0223e8b39b1b0e6367084300ae45643e825740941c1bfde7a47a841574a3f
za082dc31e29593bfa477b579fbe6579d4126ed5c9e7ff0343a7a59a00afa115ed5f1e49315529c
zcc8626132bfae99e49982b4043e0e4f57e22420f5ef6fdf692b3f30fe60cf9ca7c2ce2292cf73e
zc87e306fb7a5ccc1357725231a7276f7f984e3521f40ac5abed7a649b24e66a3207fa56d401e7a
z5620b69873773e5430321595b6116710438193f662a1f6169fadd8c08de5fb430c7577b94f2716
z1d78fe22201612a69f6323088054185bbd0280a84094d0bb9770c7f040e15517dd7d299baeea43
z6911179b5ddbdb0edb49c5d12c52df718b87e18340e8d2bdb7f80a1f3fd1196a2286dd0566dd85
z68ed8fd205e5687ccbda0c8f71407b608dd7492252ebd02e4aa2a26ffe6eb9cf957b7ea1f48e34
zafe2c0c5d45395b5ad7def2561bdb07d4e8976a847259e2abde096a7bf1141fcf194c486170868
zda9d0b17c42b141bedad46501d046045f61b9971acf9904682e82edfedea198dec9e0f2a36ddf3
z78f7bd1a9ad03764e13a8c2b6e730e6a936f2a61af60cc87bee1ba86c177253d518246f4c0e72a
z30f856c72e1f8dac7fd7c82ff6382df848abc2a6d7a6febb927797f1d062dfdbb4f927d6daf9b3
z791d9a3307b8c3c9c925983f7f6dfb5b15fe43728a2ffe0a9333cbb4d0f5b8f10667ca5a5dc298
za6ae1ce54080790882a11b95249ebcfbd2b00445d8ceb7c44a37225f501768bfa61024ae60d6cf
zb1f89bd964a0f5e86e876ddc3aa4718703af928584e3b2cd1c02ad1e7aa7267147af6b327fa4d4
z74145443a1edeaa3197fa82e46f202f45a14611d065dbe6aed99948c2eb6e95afbeff86d9b4d69
z0737127220d9b6bac2cb4689b5692720866d22f5da90bcceec161892a4d28df14125948c65eb3f
z1c1633834cb9406a194190c4c6e371821885863da98ef8eba16f7691b8acdffb2a7714f6609142
z9c975d5cbe466d30a1d290a8e3c2196e11ebd4c0e6e4a76225117d75a9ad3ba326ced4700b02a7
z86fec99c8b4278f79ef3499ebc8338fda2feaf0171b41e068ab2f45ef47fccf6f2344f5ea1f46e
zfbfe2abfd72e0fd73953138753ea558095267518b7bd7343ac604379c5ca3ed20fb63f0d0bcd42
z4d35136ef1b65afd6bb2a8d3243ce1cd403de7c336d0cbb3a738b9803dd7b2c1ed4ff9a67b25d9
z6039163ff4d33412131b83bf9056b741cbe4adb2c3e04fa993398a98b7a515e68d22ab2e913b9a
z6dfdf79ace8baef61b1b5ef8136275f64046be4b96ec14e516b9c526bda8102592f5ddd9b73e82
z73547b51ccb439c48c81c3d3f491798041d6559958083a8674c051186201e797ce37ddb073c251
z0cde2bcaeee0f893093a4cda99cc7d63b2c639545dabd6afe8194c9723155782f81b98ac785034
za72bd9ec48f88cf21b569525abf7a3b120044da9bb29ac9c1ba4379f0bf6139c0c0ca46a8921a8
z76737eac220f87c1e4a20d2c73e790ddcf898983e43f6bb2b95ec3c529147530292c25ddea0699
z947f9e4968950226f074ea3d7e413f291b7255e0ab7c5b509b155314e3507f193b75e3a26b3d56
z090f04939eedbcf592632f31d85584cf92727d0882618c4de7ce57ef06b53fbb65abd764985360
zaffecf3d5716668cc8df7d9e7ee25997e1af170b05087d26dfae12aa76bfb25b9a1c95604a6dc4
zd76e0b6deaccba9fbf958295c520da82e87dfb419ec644839056ca4bc1f35ba69c90dcf47c2b5b
z037e4f49f7bed51e06f2c2f9aada055caf9b72206ea2285e6b46773732eab2f983c8940b164dcc
za0092e5d6a6f0a00d27cdbe85ec2704635a313ba5b601e58a5fa7d2321a74b4b5ba704d12054c7
z1af9f5ea3a1326f2001596d1a4fa3bed0fabcd7d63822bfa6efe59b65dea88d84146f54d0c2f19
z12430bb42245b24b505ef8a00958e6bab82413bbeae92c4e255fa556c197a9b4848490f465b7a5
z48fda5e6a94d214ab1b5d14a4f3e7e0d5db0c701661f37e2891f3cb890eda003dbd695439cd1e8
z201675580f90bd58c1e65a42c6b682ef9be3b836c33778b2a54060a312a221eda695ae613ff08b
zdb0e996d60bcef9ecf1ebddd21484fa0f21ae3a18ecd12aa43afb4f803e01e8861fd08d16e9d8d
zef39e7a585bb16d5333215b3db1d9cc6b12f33d5fc953f5c9381af61e3902a7fa72a8ec4f7307e
z4585db842e51b28f7305d7866ba135a62d23be42795095845555582c6d432d05e5803842bd6e16
z4f1503b2655a20c1952a43d25f7414f845056bdc6d5e8b35aa59d1fa10a04f3201d94bfcc0cc2d
z74088bdecc66c5f6304e917e3e0af96bd15cca59e4460b08e4007f983d715eb96becda459ed411
zac2379c0360ddcf974d70ed420765d70d4a1f30303df7f27d4de54a5c6a13bf541bc8d357f70fb
zd30b433071c585661823cfcb00024c5c38dc86178ec6da7da61bb78b2fb4d40fb9a604feb2ebc3
zd386c994499656d7b011761087cae44c13c0272c795a2d432061296f6e389f869e0103dea4901d
z5c8ed174c37f8bbaf02bc2adf43fff6e5c646c8577286f9346863c1da518f5c4354be46053309a
z15471082cfc0e5832f1a8cdadda88d2dd2d90cf1b14dbb3c3e42072b49d0dbd161eb5ba2d2984c
z106826049ed15e4a69aaffa39eee9ac775dbf0d0e87c6f69a1d63324ffbbb62f6c6011076fa9f7
z298149b902f54ceeba00075be1e4c0a12257524a9cc0efbed8f18011ff7db0cb8016207b643b80
z29c65ff484bda7cf9a25671fa49d4bcaeca6efdde902659ec7b87eeb21251966e618f3b1c1a8f2
ze0fae7160524d1f9aa47fc3b683a0bf4c6343e8a62a445effb460ebba76aff52626858bdb8766a
z6fabda3ea0e92ebb3cf0975ffb756702bec47789834397e0957a4dffd65a8a5f9b2072e4cb26bd
zcea39cdd9dbcab707dca5f78bd5e9b3268c2bd84f169b5fdad5bea252b1de73a8594cfa539b3e2
z31e83ab9c9780eecaca3048737fac316285514bb380b135b17d72a1525ee27c830d4254ef76eb6
zfee6fee4907484e7b0ea87f7590ac20ac50140d0e5d9c4bc370ba988aa4eeb1ba4485a8587a084
zf3019e540e53a2eb30f3c200e71cc7fc7973a956e6fd5bc56a6db2a702ad79e357d4e72862ee63
z259d8d5926b64b381ea3bab0695b9fa3971f0ed570795a4f9edcaa2a7a706c76aaab4c9651b2a2
z1029c8c2d2293bd380206f05d7d4137da88e83c3c84d706dc545e3ce786ecfe7ae45c4cd95312a
z26f6369038071d057e70408a657c9cfe1573b67b8098717b473a9e7b03c123e58d4c3ba32f95ff
ze911e1408b10f17eca21c313a06dba6ed74dc33bb21049d68d40e703344d77d45fe2b137da5e23
zda02f507e0d3b09de5fc2daf31d03ab1a0886ee850623ad9dd9057a9fbec170877fd38789cf413
ze6f81312039d9e5f83a41386027a9ad27ed7d0e5e24e6eacb22384ac7e7c412f56409c6d42eb7d
z201727955a9dde56ae483965359a81b5a9c9d2c3a91f45348a6e90af55385df5d59e50fe950412
z0234c972cc4cab7d48c57f5fc768e45e8e70ecb38e97ce43a4e7902065afbf379a272d354ddbd3
zca40f24c4d9c91a822b9cbf8dc614960de82f4b75a4f799fb606a12e47d77b7833e934ebaebada
z7e99f81111585aa63e69f34a2c9479490e450a4ad3e2084c6891050599b476f8966f5f7a9f46eb
zc61cb52d973d0488d0e8ee0be63c6490adc67c91a13ae9f20e152f92b955ab7fe12b662650fb88
z63953c6d361d7be9c6a04bbbf06cc6c91d55a02fc54fa1448e10ceea496c1fd3b5fdd51d4aaaa7
z2bf75c7a13be7e414d26f420c1539899849a6a136fbee8446d702be8a4451555b1b30b8ec16230
zb51a8103fed375cbb15e7efcbd233f27adb05def77d66b2b5c5458449bc67a54556762f6d06ab0
zc62a602ddb14be5aed5b6086146225bb18960e6d3779d242e377ecf23e615e5135a819204b06ce
z8f2654bb21c3d1ca4f084cd1a1a482fe67c3b18a5fa6d7d049280e1327481342072cc23c6318c2
z563b5fe073fe878fd59df9898b802d719c5edbd657d873dc7be1870894bf38845c24773c8b893e
zd1a39c81182ff30070b6bed82a03b375aae22fa01b296be602a8beda7948d081c9ae7597e30d9e
zf15aedbc96d749cf9baa061993abc3317dcbc38e04f288caf2d8810c5398e3b391e15de84c6bf6
z5d7a18ea15b0b779de5cd38040eda09da4146e88ca25847af358ccb647828ce637f5cd510c5953
zaaeccd88d349a6211f21af2a0a39b63fd235f09b34b4627f3e77d09d78f5f6fa4bc6df49344423
zbdf6dfc2a970332e7f89d40d32f3925986b91037e9c225dcd9f9720707c85bb3205013799baa7e
zb86355c173ce093543eb60c70aaef4fbca9d44c287a03ad76346e74682c6329d785bfa18f43bdb
z75d98e2f687d52cdfb5a5079a920c5131d22f5e8aaae43f97564166be11ab7da7a499d50e4ec87
zb520b2fa50e5f09594e43b5cd202d595914606c6094074edfa50e1dc63b311e0e5d803e7f3436b
zfc739a443e2e251318fc5c43d538c48dba588b1bec87fc1ce1572485b4652af2fae63a20bcd5e8
zfbce79d5de87017eac5ff8bd7210d729d2bed0f3f9f0a51d2e67e74238ad42d4ab0b59b0cbf636
zae2b9375290c14d7d9ee43cd5cb569e334d95b9300254c79a4170f56f890d640067d379ebe0865
zdf9104c031dc1a073fdf17ad4714300f4389b7c0fac961b83d206b44eb0cee2283975f7508a259
z719d9e808618a87cef90e5cc72ae81b25c9d291eeee36820a0e3a5ba765c63a0d0eb71f661c99f
z547e43848554b66a53b4153f39a9c199c745585d94581c626aee7f66ea883d09efef4f8f46958d
zaf0f9dcc1a410ba6227198ccf054f35315437469587a64ce33ae57f07267d4bc183293797aa713
zd503169620226ad39cacbb78f020442188bf1ccbe307ae7fafd3100f466bef5dda057c77af77a3
zab5602de1724d0bd6e765d27057ab1a79e102a84b2af19bf1df636d962e50e86bf6481793e34ae
z408bcbd5d28c9778afa83b04bf50a87aa73e86822cbf4c1d6fcc19e592b44d472553034302e92e
z2c7fc3f1843a6a052f72c1b190972dbf84b967d2f4c3cf876c570fdeeb373631595ae181db72f3
z3fc004328267c1ab8f2799fae8a60360857213e510955430ddfc729c1ac4156a0f567ed07dbcfa
z7737adde3258dae20a613cc05f6b1d613301df60b84392ca52177711568fcbfbb728cfba83beeb
z377f7a78bb8a5441711bc7f304d581e10e18f74eed11a803164b992cbcbdb68a4dcd3497a0ff0b
z19b651a0ae67a5ca0e171ca3450f1b525488dfcf76bc7bc0949cb238350885388a5c684980f729
z797f97e0d04efa955df4566f476be863bc0dd64bfea79b0920e2c0e180153f217f9b556b522438
zf2da196e8d0602978f0218357862ef09fc8ce5c42b67a6394c82eaf5cc1ab99050742b84402d0a
zdbb97b0b6286108e3e5f22ec81b30aef26422a19390ba50bce286afb14e2700798398678b0bb39
z1f1ae613e2dfb956791d0edef003f1ec088a38b4c0dd8342bb72565d57c9850d12be7bf0a29239
z180d0259c95a41b07241ef7af48a162d187d5d46e140776704583d4fbf541aac6135c43ae3e68d
z1da6455aa9d82be0df89b644d6e3c684ca65eece911f7972714b4a54df2c89dec066669019a837
zc242c53d45729ee8430b6ee2ca876072ec33cb33e40eb239bc415226e1e9040a493cef20d8e59d
z9d9b0ad90daab8d4d8286a7cb4a745c93021ba2d0cbba98460dc5c0925e345dd1bf36f2c21eba9
zeae3b1f5fd8cd8da74717e2b14ab35ffe0c7b916f31289a4d4940ddd0b472082a321f6ec8601b4
za09b39c36194578a18808be4ec59f62eef9838c03d534e2ed46068c9c13838bf39a46054832d60
zb91e14fb3f28b63538847c8a6b4003b82f6f2382ec4069c3cb2d5a48fe464e606591550e1d01f8
z7c9d55cedd73e853f047d3565eb1c11882ba0293221fb6b61b145852aa0479e56ade450c2eee8a
z40162f7fbe24706d5e3bf53355f87f64e1ae1ddcc81ae53405917a39b5f2e0929c7d7766e4a73b
z97c082515f297da4f6a50037cb9fce376bc2dade267ddd3448558dae904d74ddd625ed5115c63c
zab009322c05d5bed6fbcc83ba9d0328577b6901003142fa78afb29054cc9ab7d409369a6336d69
z8e233a70f9d8203a6c7c9dac35c844629df3bf42eb6edc9ae877f9f498a951f4b1a21760046c63
z07b79652a73dbc097b50376ec23259b4de0611941ee03e4145dd2e23eae157de86ea3758632b43
zfe8dfbc79f2cf1318a6be140ead42673bfb847a9973208d1d7d713490ff36ed9575ade9fcc4687
z129f45285531f1bc1e0cfc45b76eef18b49a99aa561e9d33ce6be5975e36cb898fc65d80ca4cba
zfd281be134f10492606acf4e7361454b57e530636fd54be6a364d31597cfb1d69e78713fa215e9
z86b03bf4a05ae5c68a3e6966efe687ee67feeb3246534b0c9ad01b56e824b3bdd8765d4bb4724d
z70dd27545edf1ff250d6cd6e932499ba5ff7c6bafc1a4b6eaeba8a3d5ad8110a5c78e411f55988
z007e008c0121cd4950bd025755169ac76888c6d72087c8003b4e5b394ed5733d7e30657adfc76a
za97d2a3394c3cefe69d446207bd3d62500497860b9d3471103418701805e97c4004e284acf07f8
zba51e747dc579d1f8cd761f03040c8c3540df88c2ad280c7744552149081c2c37bedf35fe0e72c
z5d8a692edcc7220503998aaedb771d2b2ff743fdd6e8316c25970ed4eedbc7d57cbcd96eabb698
zabe3a8f4a010433178b11b0bb15a1269419eba439a6d641cbd586367e77c251aadf010ffcf6b8f
z6983cbc4f42b77d81ec12f6a17deb1e4ccb3670bddaa4a86c3f76c0600916a5475bff52909f2b1
z24a76136f27ae6c0cfb3e694249ca8a6418ac67bdd4c10b524925213ce1eefe66b7a0bb7ed5d89
z6f15fbacc50bd14e9fb81cd33dbbf74f4401d975dae0c2cee778aabadfcb5405f694d6b69c47f5
z03efc9d1cb2a30d213342ececa41220c5076f440e6b7518077269eaef72ae48a338292ebbe706b
z875e2d4978b6ee6fcf6a923ffafdf8ba7b73d59d59572f1845bdc3186b5b1c9f2473859f1d76d9
z94d5777c03036908c5b3cf2301f667a56cf8bc89349647817c45a4dc932c50c6a58e8611fe6228
z651c636e6e090a0eff957dde427010e6fec71b721eacda8edfd6ae6fae23b020d44039a350e76e
z84ec76e922c0ac7f7ba7ce56ca0d2ac680009e649b16e8617f9ac7006b61db72d2b3251d10f7dd
z22185215de06066ba4a1209c2679f8bdd2624b284d9f09b5a6994587c1949820d010a092ee6796
zeec65c248decddfe219aee0cc732972a4780bcbc109890c83bde98a73b486e7d8120c4bfa6145c
z641e8b3297b04f16e3b59d53001664b0100dfa64020d83af87db63b927165530552a0f009aa99a
zd5b5f209882d7504b84acd52051cb7392d7362e1646127b60d0299da6cc28b700d235535825357
z0aafb8267a8381f43ffccdc57f1d298238a210a10c28bc93a59bea1cfb3c0d1409e2e78f101a94
zadeb15657a5635d9ebfc0ef52b294ea16f361527d6fddd54f78d9dcc70c65817172b3126cce005
z3b7dced99e4e1f7ed92935f1b58ba16ca3c0d93c489e9fb5d16d1e2dd3e3842284519b992531b8
zf26ff8e19c402092a236d459c40a487ff7a3c8e1baf8a30ac2d92c0a8e3af48e122d21ae662f7b
zc8cca7696123aff4e29bc78476e0bbd706140907e7d019075a7266a2b2f8bc0358d11c4611d24f
z17c5f883e1efbf0f22fd6910ab0e116013514db49a5b43cb35a0c44b3cf0f9fc15c0e9478c13e8
z7856f2a331beff7870adb74bde99d21ea3bbaaaf45a5981a466eb290f6afa77a0c45461d0526ca
z1683f257b99aae8bd921cd3ebd4f2662580474f2eb6fd85d74322e050b2aa5d7607afeb7d4416a
z8f47d7ff51215f117aa01d745e26cdd921c7adcb78da6da2b5c40ef991e84a01332d1bd191028f
z3fe63838729f976f5987a60bd2c99b22cd724894495316dbb0fbc49099285fb0cb5932f9f2ffb6
z1c546ce7d3f37ceca0f791f1d1ffb17d620fea6da3e42bbb000137ee69e65824be10fde6feae6d
zbeedfe7b2724477d07fdfbf30d1124e67a111fdc5556033ee4823a5b21276c252a81dc2ad3dbeb
z97ca3dccf036b2096e8b6d69e0d6d5ebd7cebdb800e8ef9a8e395f9c10eaf6613372cb90563eed
z61e5ebb4ed03177c8b0590a357fb6a7aac9498ce01228b5e1ddf66b7a5c79159805fe24ac0a2df
z9a0fd0e8f75cc0d4bd5c958d39c4810bccd6152a360fb55a71be02be55257559ac7c2882af69e1
zc7da9d2c3de80c022ab55c1bb5a52825b1964a2de6e1c6aa306b2968552ca68ba830bae7c3e5db
z6201340f6452241537dc656c1e2103fd70a973cd877ebf0f05c73d16bacbb0df7f794e11c59e7c
z869d1a623ba40f51a71841694c7eb9501751f517c4a682d9e4f92bc0d20a85dab8381fc76eefb6
zb4863987e4a22da259c9b8360c51ce1eeb8517564a432c79bd68798ac797e42689f0dc50e39898
z0506d03fb972af22daaf318232ac31f6b5ef7ebc299c73b0f80991407d4f58943b346f63215b11
z03103172f1b033ff8a9032d54fef78bef91cbcf522beb803ce050412040932db233d3ad5b908b8
z9cb1d30c48ecb525e6af784e91f0545adbac68359914845d3663d786b7ac5669ed07b877cb256c
ze5406b0f19fad3ae1bfd0b745a4c9f0874bb1044c71268d3eab2148ebacda42b0a915312353ee4
z97a73543a1f1472e05c44b90a533d633370d260dc17f3dc830403c612571ad61ba419d4e68c1b6
z83197056bf3a54156aeb4bbd0ec4de2270c3bdd910ff249035b836c49ec67171e241854ca576a2
zc4aa21d669223e2d56a1ec2ba6fb1226cd9318e732059468806d1266c9715ca7c4bd56d09010c8
z7b6161c45613f4f8b24e616e95d861f94616f3fa44568e90f09cea4ec90b125af6ec720b94dc7f
z560b914790afdf2f7b1dfa11b24b011510becb64a31b125e06ede86f13e9c646ff852276a77756
z880193b415cbbf459e51a3481ed367b3718038706de754f373996064eff3b67cacb6db3ba357ca
z7c77d66fc2e43ae3eff64f108041f5307c451e7eae0098ce45aa3b752174c4c27799c75c1c40f4
z50ded934fd92c1ae6dea4b6e0811647e1294f9ae27041436948aec3c96bbd44ad5c2f8d7fed027
zede7847f4468239240dc515d0df8d38751fefdb3d06d817f58030649498e5cada3f849359dbe21
zaccd4692c24f0b68df604db5d371ed39c8642027223c9a3ce47be4b3db09e17eb232c0c75e1b6d
z15b26dab9627d67d4b4e4ebe4b9da1ad7f30209289eadde4d08bc164f41cecf29ccc03e08e484c
z2c1632e7a1725cd72cb0d1acbe9fcc8a1b1b53e74a83d83397078380a6b396aaedf5db60ff1418
z2a91bb69078e3d599798744a57efd54566fd6da5b8833daa074027fd0297cca23cfcd2884f337f
z3a1fc0ee0496da5d50786ecae317113fa0149eb7480e9b45327f0db73955227a2e59156d7d9e95
z6cfd7074ff4dcaa398c33cf8405889e8870dce823803e4590399a7e52993ac1db740973ee987c4
zd690eb59e073747c2bc823bfb7dc929d621a6f638fe8485ad700f44ff329995f4e751a7b93d1df
z704f34d75ff51f88c0dd36ab5342ce9b4cca744e789f47077a2ce33a921ecef292013774bb6383
zfa66d497f83e09a22d0c8a831178611976e4959ce5376d78f1f23a83bbc8cdbb792f3c8c40869a
zd8eaafda0466947220c762be1c0f0387163631d08ba83c2bb799d7031a7d953f66b306b52242f1
z7c06e35159eb2d6a54de09bfbb46c6b2a71869081f5c661d0f6641c5e3fe4b81650ad5f842d297
ze23e5ea00960cd2d7a4041545260912d0d1aeb451860c2bf53a6aa0f1e1a582a63b7b5d4f066d2
zcfd47fd50bef989e95009d36a2bc9962058f7544f8e3eb8e0ee70f0c4370616dae490c4173ab9c
zdd0895d711349047cb3e6ba50230936ce5839293f02934ea0d7fd79fd13f8a2e6f504188528a6c
z72349462af5bb01740528334c197b1c32b72b64f50ce155af91dfc56fdfb7be54ce5d11d2be1f8
za28d2ef3a264f31a29063c1666a587f8a9c877e0b64050c91e3eabf58c4ffabb9335bf71c66513
z45354fb00cd490c7ffe15c7696494ff277d8820272575a279929a4ec9e0bc305ebfe73c938cea0
z33c22512ef5de14a33b2bf6db5afe43f241ca3fc2cbe329c1eb20947d9d0c25266209e48e978b8
z6a8a37c3200727d32fa733553cde1e29eff8f720771e361c37389d9bf53ae93e564e3dd7b520b6
zd251a43d661c482d7978ce052424e018d82c692b5bc91c981551ab6312898b3024782056cb2181
zb64f6aac6225d48a4b3431e82ae8678495d1c23a25e060231ff8e3b0b1f1f270eeb6860c94d079
zbc9c25ce6e979938f6950256a58ec103bc819d1fd68916c59c32d4305513730f07c55a3ea3f3c3
ze9ce7af0b022ac1c47123a528109835a79bc61f2c35f112833787220712db9ffe4713c74f27cb6
z0bc3deea902c254d39bc9f9fc656d8478adfd826bd7685f2bf56ef8450173832f51b38d153aa54
z6addd3136861d93bcf902cecfbac63b6cf1234ab9f55ae5efb533660d8806c3d000bb32fc9a28e
z85536ecda3ff9b32ca335ce8ec3dde345ee2936be2c8ef4c9699e761dc927771cb2377b33aa093
z0999cbdfeee5e11bb7960cfee0aeb099336527335acd0da91bf80565e45ffdd541f2c6811ddf49
z0ffbc1844f23ce08cb819a64a3400010568c9509f81440d1be23ef3d2373aa03899a93ad39e7f2
z6f8f27e53b7dfa2f602fbe7d596b142985cb056ff1c0d4b98efe96342eb08523ebd1bbcf4760e2
z600fb857666feea612c691a798273534e337671d6bc433d71d912d5041c7950b3867e5e816697f
z6b670d00c49d32f31ae0617b10254fbbb9c02054f0251b82bdde673b94d79b2a1049fd15fa2331
z14fda4b367dc771e756e832084f3495bda2d32e518de8d454e093ea6839d71d6cbe0377da5cf5b
z9ef0095aaa7af9267fd4185be6478d030d5e66c57b98b436a44646b2bcbb9acacee9ebc0551b45
zc691b388f5c01d0472ee7fd8d79fb83b645eac5ab897653a10e08a5570f824fc49655829f7b410
z25145f30f24abc16173e8495bc395747a505ff7c279dff6325bab4647429e38e773f66344d8dc1
z0ee844f8d849f18e4bea7d4a97499f742bcbc6d76c25dcdcd4a8468f2bc8e753395de4a071b935
zf22b0ec6d689ab8630c16f31617b652f9104fc2acd423e1f65ce5748ba6cf4b2723a29ba61226b
z258b91735827f93c932c6ff603fbbe6dd0e8dd486de8d8c5d984ad5f946330c15eb7506c7013ef
z0682a36cf18524c60c7884a10f18aa2410f2244036b48c269ef9398834e96b366a168a4c1fc761
zd0c0b24957cb71385009556ede953d049551d477548264459c8084a75bba73aea551e4bd99230e
z2255dba639e1d9faf0acc3245ea93ed60739440b52888866b7b39ae616e8569fe1f77fff948f67
z98000c7b4cd3c3d6b4f07c301dae3d22b907d984496cb65059b091aaafd6be10139bb3d45c72ee
zbd7fc7e1ae6ef90ce95bc90d20f9c82fce192c33c3e3914019b560d8c29cc344725035a432fd94
zddad754551784d37a93557b3e12915cf566577eab33d32733fd5812a80b3d4f9ef17954272bbef
z2353c492cc9ba17d524e253f9260966fffa44c1e685ff4d9aa4e421426f71b7668958ab1814c17
z9752093dc82a2392bf70fe606dc192498589f9bcdee09d0c99a8dbf94f2c23e98d515289d1c7f8
zca36111fb76f64bc607d3acde547cc0ad2d642113b1b22ec543a337bea184cb244a0bd38bbd1f7
zf0c0f49267e378888c5e940c6c6a5d0fc57f5e59eef9dcc459e58796a512e70d4dd1f73d8d2c59
z8fcff8af57ab993545e66b1199b0d027707c9625493be3be691e96dd13df6e231b9f582c8301f1
z9863e1302566fb586f10e05fd481d952719f86818a8ceb8d3a4827d246a61a944d5a191736dbbd
z8377fdee4bdc8e1a2c313e321c35ad8c283612b9dae52f296a085b2a693409e51b22e5229283cb
z8c0b5a731e7898c678e4b55aec3690a1b7be6e6e5d8d607e2be29f0acd1b3f0aa2d9250a79d732
z8e31962b2f51f4993887b0fbeeda3a501449881d10ed60eb33acb9ae7e5fb582f81e9eb382d98d
z2e3408808fce2002ecbacd863391b766fddb778d817219805a358b7bab9679187238b1c28f5b3e
z4ab5da441031933b4ceeb6f8b042cbadbc490f4f05fa87ff368ca94f27c1c88bdad280b145d7e0
z4474130fbfe0956ce38c1cf5c0eaac965238995c1a50f5c24d16ed141372cbb2b57b27ccd4b01f
z02072d5168304cfd14eaaf91855c34cff25c414b9f0dfcf49b714ec4ec9a38528ea0ec8a7c6ae4
zfbb043b2f11435778124e58dd83c619b25c02a6ba6349a844021fe91cf78920aed9b9558df7831
zf9d819adabbee4aa361907611620935c5bcaae6f526bb815dce261147c403784d0f062ade642f0
zc7116ae645ce11d71402e79195bdf2ed52fabf44011e11778cf6f34367a57a4b3296ea5c85ce3f
z6dc0cfaec6bcd2cf0b5f575690a51135ea0658fb8cc308e9c2feb5b532439e4e5406bde23af279
z37012e3fe763455df0274e70c724b7025f2f8c25efa7d033c54cf91a3c5ea267f387093a462535
z32b633be1dbcce8f9227cf74358467e4300b2deb4fcd98debb2a1f2dd208f75171885a3616c993
zb90c13bcf1d3cef34dc7f956c2b7f432e9a5705b226dd0234e8e1400e950f4b4c805ae732cc583
zeb2c0f633065b8c4b19328343f16a53e41b5fff0169bafa7b32324cf2cc77ef0fc97855ecdf3f0
z65f049ceccc250706bce23f4ba215f0b49691468553f594d48c0c7837ccde86204152fc3aba291
z29bbd34e72647d54d96f0dbb59b1c275efded2d4e97cbef02849fbd4227e93e2b14132e061591d
z97cbde9911d8260c79e386624f6c923b67d40d5bced7966c9e613e17ecb756c4190846d288f309
za775e5fd417f570b26f63cc0581670094a79bf4677d4aa79721fcfa763ea62b1d35e3040ad2904
z83b7b4ca57a0f7c1aead900756bc738eb22cf5526ab0213b946e268368cc98e3c183654d1b00b6
z54eb487a7117689153943e627b5fa775110d68a0f6b328a92918e70879a1deab34dc0369134aed
z278d8f86bc0298b60b8cc0f74f346aa12edf63e400107d2f7a8b72caed4df46d09ce01c035dfcc
za8135275433e2a0485ad5175dead3a5ff7a5976ec77a3956f94665c054121837cd7a832ae9da43
z939aa77ef06cff0bb6f3f3a876560a9d40cb3bda6f239cd7f654d593eab7f76596a8696870ec35
z8f93b369f0616a77aec7e779e93856828c3c857e7b65977920b48c98300d5f70a026678c2ab262
z35412ca650126b9386139453c1798be7304ad85b94fc520eed4403a284c56c6a15dbd1195babdc
z16a8ddab3f6903da02676aab65822abb9effd1932ecf274b64eed695a61c374861344d44f3b962
za1104099ee244a597dab22b13490e5433ded8aa2861a0c7f66d26f4a7ba0dc78e31996bdcf137a
z1e6dcb3889e9baec1600e5b440ecaee91ba0ce745815e004c8d9f95f4b2f3e7d13b6cb150231b6
zb1a9569b57b07ab791d90d6c598a42930fbe8d4779d3e925950e2f528eefe8ec6fd2f4d0029978
z652b97dcab041a36dd5f9482f69267041e4c5cdf672225988c6032d1d8b6f93401b58e719d562e
zd1afcb95763efa00250b84c5440fd5923021308f935c4a5c2c6d2f63cbad3ddf1c06ad6ef23f61
z1aab07f83f34f0523859c6b85b9964762649e6166749b8fe9f0a0587675c22618802be79e190e4
z8f580c0e0964c8971f77bc3f6d772e400dc36337d2e1a66020704957e73f685d3c551fa8597f52
z8e399a16362eb458309dc02e474de74d4182ba6db91cbdbc8c7079efa9c1b0aec605b8954cfd99
zb66039b7bcc3d4778c942b69272ea815f70930cd5c4e082a60fc9192f8875b2974d9b1afbcafea
zcc0e4d19be4fb5f87ffef5158ea8ef342cbc82c633fe6e03235893df6f9c4efae2cb41dcb84e8f
z4e8b92f68dbe31d04c7460390453c2cab44a34c5d9298e45afce52ba36a7dab6f5ef5a10793d7e
z9a0e18715facb814fffcb8dfaf587e902ecc0ea397236fb6c135f0041a629752110cedf0bfadc2
z772b66cdcddaea6b2a6e710a3bfa344c7618f222baa7ab6706e1228c9cfb1f19185277d5fcae7b
zbd5fdfac9acbccc920763522d19dd02efc94dcfd42f3dbb6ca8dce4db2402e732085273cbe914c
z0e3c21cc9312f15479ade62539416102442760d2ef674e9e96b771f849ae73085c6f75fc1f371d
zdd2712678e918d8c67b41a993a51b471d981819cc350b020e04ef8bedc9548c36f61f778171151
z000475741869b4477f416f44d866df2c58de0d41174c487ef2444eff84c5db630e66c32bdf1efb
z9c24be1e67f7fb765abdc9e9a8aa66f1852b6efca110333e79f9b27254afbfa69ed2cd53969da5
z39397e19e142beb59d16335a6291951bc7a35917107396dd7de54733e196f22482d117998c8dbf
zfefd1533e2b3de59b86f11f1158fe176be5913b3a9a38ff56cb2b5c5c70dede33aa81da2e221cc
z9ca726a02c4afee775600bfb89983823be8b6f9497f20a173065f054b93f195dc9d3d11e648e10
z3bbb120725eeeacc5d02eb201da278ca27d5a6ab3513a4fa072b5686b484568cad8aec9d5dabdf
z5a832fb39370b6a238c2027f49b50a827561d6abe8b812f043754444be0e8454332f8f560fdbf3
zcd7c0ac80401c2916e4f166c13c6a850c4f9ea59b30df14fb0202092a8644063b7f331de8ad31a
z51a9c724581f8d1b726a914044ceb991424fb59b0a8892c01413291a7c8024b809c199e127f7c1
za53943c3f067ebdbc27cab34bf96ebc9794ddf59f9df79ce851120d575030db5ce43f49229ead7
zdf22193924297cf02a779c15d0d8ca39679720fcdb13477d3f8720269f1a866ecf3b31bf3f3279
z3ad0f3a22b7b35b7353cef23d423da6300442dceaf3f7d85bb41235f9fc74151b43acab560ad2c
z49b24479dfb25a287101340e2a1151367430ac0c5804181758ac69c740c72077a0562271154ce3
z806a49e7b40012034597a78d34d59265957b8ca21fffb0feaf2173f437000458856ea9a4a5fa72
zed4453e2bf0e8895fc3c4132a1f22887caf98eecd9bbe4054282a72f1d02c29f270d362adc7886
z4b86b6bb1f58a0fdbd50e3b60e1650c5310484b229564474ee89da97bb37df01e59fffe575f41b
z9be9486990d41c3bb59cfea961ce1e3877de1c5bef17be21c413008588162d08cee90e9a6ede1d
zad2f44483d13101531d11f3319fa54e57159d60869821ae128c28ec1d7968262de2258eeac2f1d
z41a54ec274c0b989a20a529ab317b04a11db4e77728f899fbeeee32db75a99fa8c3c5d8cd79f2b
z7673e9c048986f6b6c2541b8bc4554d51bc4e860073229661a8077a6dbf82f467d951cabd18d59
ze6ea41920e3bd1be3fc2bb70d5cff756de3bef28233204b5878894e41ab1520d048da71329d527
z775d6c593c5066e357191b2ae40b7a31e17f43060198e43f501dece061320ce222ff309ac70c7b
z4d69831039041aca518dc16bb9af8c143b606d9ac66e1e58d708f1ed3858acd8440c86305a60bf
zb3ecebde2830e2e2e83208b6da54323b8ac6e23e4ab22d9b33fd4f072034888fe0ee69794bc3fb
z93000691bac09a56ad21e90904425f75c3f162dc010e6ecb6133a3ac5f539155929fb20bc7fe53
z2b5756453d1feee2dd4787c6bd131396dd34958c2f8d65162e0c3aea568f392ed8651db875eca5
za1ea1985874fea587060b95437108a2445861ada36653c9ed7fbe95ad8586cf12c67e983b3c28d
zb3b1d6d2e0ffa976153c61175bf2ddf58519557a756e34b27fef739b39e8ca82fb0b1d814fd140
z67941495edcd3c13be861d64018988cb8590bda39db6501145b7ffdbb9546456e7eebc0823962f
za3d470fd6747d42eafd8a4d51a983844f8b38b7456bd79129f3e4efa24fae3ebcfc556a9872ba6
z93d03a8cfd05628f5c15a9fb69ea93b5af8f16273cfab5dd3cfeea76b51ebde8f7563de4c6d063
z07bc1714bc439d524753a7396bffb4d5ff97345be1ec2f4211fc49d2113e4de9f8d6a56296ea38
z383a24858363c60dc512404b807ebb9e7d3de1f19fc754d158b9d70738a29fb871656a96c6b200
z3e0b7223a7976d160c49244bea169acc7d31717f250796261888fb2a3210fe8e1e3dcdff7390ce
z1c9151fcd6698f12e49b8b04193e90ffb07699115ced515e11889f69c25ccee40ded86da96042e
z648aba9f628ce4b4040d88da149d1f5fa13839d4ca77c897442b3297348ff3780a60d22c5928bf
z42678d3c4ee362ea65b34ea38d22649ce4c7ab315c40df5acddbd3d9f379ea477a39833191e45a
z6d46c259e98a649da3d12206501769d21782be74d914344541ea52436f837a877ad2f4e79e3a58
ze592f18e7f1bc90c47e3ceb55a74e360317dd036007c0bd1f1da0c439f0d87cbd5e3ad30dce0ca
ze4e233e5eee38145a6bdc1bd730f4f22bdeb00cb7f392656b24bf464c549486ecb9950fbee8fa4
z103a1089a42a9209bc789128acfd5edbdc09406e6aab57391ef1695de9e64d9089d7a57a602c89
z1d3eda1729856409460195a59a1db9bc730fc42bae1f91322b828dfe0ca1eb17b679f0618966ad
z565be39bb7a067bcb26d528dbf02712f4c8e1f56b06d7ebdb2a796b9c558955f22aaaa53ac8ebe
z2a12a3a86625f9f552dc7ff1e26ee8b47881b30565c5f91f00fa717f1a1f93601b839896bda5e1
z0df853a73eb0f48c696c30c72e3435456f76e629a48e8c3bf3aa8252c4d4b9d1ae719902c03846
z866c10799d7245500faaca8d1d007b35902d1344e0d3934ddf3afae8d451b497ecffd9223e95ca
z7ec8c7a130da11b05fd5dbae57d87ff385c9f3447c3b02f122555982c3356eba3658d3e1a10aa7
z2a4cbb51195f1336ecba49ad98fd973cd5a8caf4d207c8fdfa4bb62e186eb65fbf906f0c932b55
zac0dad5254103559de009d13dec2ea31ccd69ca162db643e6a5c21069f26fe26a54cef6bfd27d3
z15e4717f47546bcd8808a30141cf0fe223611cdfeb7ebb77e5395b40ad195af28515cda92ef7cd
zc6e2310a3f597fb91ac16ae32efe2e199673f50acecb56d79d1ad58bbd633405574edaba30a8a8
zabca0c262b48c5ee5b20d116c81e8960a5f573eb9b4f379d848a748c5354f3e5f7c74e18fa2000
z0997997d7599b9ff6e3db5eabf6b5283d8f269163bb43d9f575566a628e7a870c64a3ad7a9365d
zeace7709f7f080b70eed7b998f3c852160a2eaa2ff256c113577ea599a6ec35923df6836d319cc
zea461a647572e0ff8b9c41783e56287eaa443c7c8cff2914bc46991a44811c9e3e1fe7db713424
z09f0d7d3fb37e00a21a5b3952e9827cf095d63ce6b3a35fa3e1db05b4ee6ef8567efd9664e5fa5
zb2a6995addf9abf44823949daeba8a9f70b0e3f06a4ee0819bd86a21ae2767451e5dba3ba5b611
z97a1ddc766d64a5c0853587bba3ee9b6e0654e411121fd9265ea0bae51f7aec233861f4c0397bc
z96f8dad09b95ccb7aaf1f50f128005f12ac831ea928954f4b7fc1ae0878ab770a4b8764abe04e0
z8e04165f3bdb242df6b49c0165a8f249cb4347d75aa17b4ae301b93fe36304ef30b3e2188ea2ac
zb3097c7635080e09ba92fff5e5a655c7209f37a1a355dd6995edad9a5f12815bc2e9f4e3614a84
z1e1eb31dc1384eea57b7c9cc6481a4d112eaff5511891d0d742ce39e5dce8e0ded2fc295db62a8
zcd104292d47c101ddea74213a71f8cc1bbc42475aed6a177703618da23b12753f7cd0aefe9f275
z0dbf9d1818d5fdc7d66af5ffde6df1e23fc17d740685444bbb8f73dc2110edbea5d1347c1bc707
z643e247e9d4540bfabc6c3fdac2a1a029c99f1ea19c92171977a3aa36bb9e9f837bc7149e270cf
z79c3e50463190ace6f203957e7772840d198204f9745dd9b16f9c081afc234e7a0d4b5ee4e58d9
z3d2722433fa972f13cd2ac338b67cabbe5f5274e97a779ad4254ffefd251216b05f94ecb6e3e17
z89ceb06f3ffe277c7d6dc2eb4f439219e794f23e69ae7447581d1a1a8598c565cbfa291dd5df8f
z4d0c9362131a076257498dba8a7afeec9862ead4b1029446f8b37934a318ef8b36835e521cf342
zde8477e7c3bb8580e20ce5bfd15d80817752cc472b001b24a2f231c5c8c200e93598442b4c78ef
z57ef9acd209ef5174d5d9c4e4f944be3222c52f3867e7cc1ea08fedf303a84f460864a1a80e133
zf2c092fc7cf4afb441986fff6b0df94d7528cf00a2b454c47a849c83789d28558d6f561f5adac1
z063751a5711ae12169abcdd96ed8e7781a8df3a19f82e101480f4a0b115d64e4ced74823b28de6
z8d7dcdce5f581bb4b65f962ea1cbe0546019a41b5a4f31296e92743672621e7d9030665f715bd4
z4172b7f630c483b2410b8571beaefc62363095770c9d47e87d3fb93a27b5ea81f082fd7da9c8d0
z1b6577468f8cf9fe45b7f71d17b6db897cafe3f44dae2cc237787706f2781c86f7d76f85c996d0
zb04b4eb4a9c7b3550838e04bbf02a0add49db5a621a9d6ea02b883762e2be94a487ab8a8f24885
z4b7d7fe13f839e37c7eed21d60e6c426a5724167426b72cde13bc200073eb51322c788b7375a6e
zcf41561d50da48fbedd18dd804d2e16e343889b905798fc208fa9d9b07c59896b68909dc520fc0
ze4a5e28bf4fd11404b36199836a30a9f9e7ac496ecee2178754410b645df46db30fd21ad9a113c
z941f484b6b68d3b94d420f62948961e9aea0087b8dd9e199ac5ff0648c7c401ffe6e68a7f9655d
ze87a50139c71b45eec7d7bbb1019213f19e6e940691530f003a9ef6fb7b133735a5e744f2dfc34
zcda740fe4aabc5425159a6c84b6b4a4c86583abdffa3d1529bf761c303e9fdd50b374c6ba5ec67
za386ac1b0b8aae103bc8dd98b115d18df9e5a78c54082ef529ca36db6a155000bf492e9db1b82f
z7af521386aa49e153cdf9c47ca29494386e14ce3b0243136599a845917d326eaab716b9ad5b719
zaa0d8552ccd57436188843d5830a0d7bf812ca3d908204175cece7d5c95b3a79c543e4b2713bdf
z91ed2558f4c44e35f322341ca04cb19de94390462cd6164a26a2dabe8f201c20a3e2a3da8c6cb8
za114af657437e2dc2d2b60c7bc8bcf657eca11ca0496d52d675f30a2d3ac4209bcee70fb8556db
zdd0715a073987253cb0195187331889f0239c761cf9b379365e0e08de95b1bdd978fea0eecf7c7
zc021fb0179616ed3887ea70831feef2cb49d6b4aba4586e44bb24d3a6aaaaa75eec41bae75ba29
ze641d9dadd8fb41d1e03f4801967a0054caec05c07194548c38f2201d47af67d294c3bb505ffcc
z113dfad0db136ee1117c072189b7ba2e6e59c7f278b3f955ae90ed3a1456aa2828d8b23e392552
zf4f15e3f6cd501aa97644a458c7960ddfaaad068e03748f9ab2a651a92ec91387ea8b270fd91ba
zd67c079ae6047c45d3f8474e73f8bab28aa3c825a6360c1ac848c737f44bdef4e75bdb4c58483d
z8d499913aaaeae89da55daaf906d0c6761baa42f5172466f22df954a1237694cb5fad9696ebc92
z441164dd2883302ded89cbe18006ca1d72f7cf7cbdab6213d5079f445d3cf34d389b2aae936616
zedb8667a645286dd8a5fc5e9c93389f7914bedf8bc593f39f1a48963b4552e47548bcfcf6f6340
zcdec4ab0cbe7f1daeb62e35059f0315acb2dd8a179ad2fd46f6bf74e4df44c3e744d7ab744afb9
zcf3ade8d8e200a0da341718620919e5d144f4d0b566268e791791879827b82d25a3b26d41732db
zdb2597ffb43511a597a38cef4336de0bbf01a2259c237f8ad17cdbc3f616e43eb3be8d8afeb6d1
zd8eeeb9951945d84bfc28f9ae59a868749bcf7dad42540894ad5ea06f05dbd6deb08eb1992d621
z153e6eac0c3ff9a9d68f103e18b5bff3df3d0b2f2916c4d980c2806014d7eb1b9c6d2cacf3de00
z84396e24ad64f5e072b75effc8ba42e883c6a4e3bc9e7af30652fe6bd320072b2c99c05c3e0c4d
z70478ed7bfe1e228710a0e937821b4c4bfe77f05d8f49b2610bbfe8940d6029c88c0ba92c141bc
z11dbb6841aa5d9b8643b1e7ab8719ee7202c261ae9528dbcbb548b171db0de29a217fedbad8dbf
za45d39debc5a58cbbfc42449367538ec0a2d57a07c29bc170b0a2dbabe16a7f11fc2423f4e1af4
z69be22145eeaca2a007dabfbc015c660977ec0efd70ef49cb9ac4dcbc87d5f3a8684ebd7e2071d
zff03c3220b9c68c8fb9cbed208011bbaf4703c00f0e0fffbd306cbb2c74f990fdfd4387d5358e0
z6122d6d676a29d45b5f446d05c80817b9a43fafec016d9b83a6d938f2665fb4109ff16def46f2f
z41a129618485e08f313715adc4ff3a143b97869a07e72596cda675c46e4d3de4648f2b6abca264
zcd6e36e94101b33dcf216316e14766c17ea3ffcbcb318fd8f90608cc51c99326ec825163ba5253
zf82d8bb8eb052e6e8d44f9c7967362635172c333188f34bee004b65c8fc6d19b16e2bc52206f18
zfce299f489b78c98210c25c49695529a5f2f57eb1ee46fce31b30c79f9120634c866f80909f935
z6048cb81a65f107c3abb443b2883eadd28913c9ebfde1766e92de89ecc64613dd291fcf2fd1f44
z560d683322e6a654067413cdcc9a8836b3285e1d506dc4f36ab4eedcfa11aa68b9eeb4d0d436be
z6ee0d6f9c290550f4b6853db7bdb0e3b7cc75743d8c1041899f300551f14cdf3aca6e8bce325f5
z21c9b95d5d73484b039c7aa06e682410ceff81d956790f77a560806ac4d7005a72816c67c924dd
z3b6ac6488ad2418339929f16ef1be4e1cc21ad126feb2911c7224f0218e6fbb33f2e66cf538e84
z4994dbdbe7eb1f7bb705ce9e00478997401196bf60a5c348631a75e1ce27cea60608d53ea8b370
z8f0eead84bf980550aab08e1b4bcdc89d2e5747cdb95ef5d1a54c10c8d3aaefd1e39d13ac74f09
zb656ed03908de93f0ef0856b089388e0927a9caccce7acc2fa15e18864a092cf0147e686f24b78
z202bca6a33b2e319f513aa2b196323e40f04d4701c06e98ab085f1a7e10c48d6f4dbbdc1752934
z68fb7c654b9839c6667572ccaffa9de19acb507f6186356c119d203efb64d240964fdf9941fbc9
zf0b5d60d8c8477038e6b34b081ad081b6ecaf2e8a95116e4fc952563b0b332d7db9fd489055a4b
zae2b545f8a21138ff0ee29434c525650a7bda8ef4c9ad4598fee8b585563924cf6f7b73e9f84ba
z0cfd085e0748424d158d5fabeb2618076adf1df2a9ad2f53326233965b4b18e2920e62519fc199
zb8f9485abe4e07a6b7bedb6871e68e66075c8bfd84118468b60c09f33a0197cdc3213387d18566
z8d90b6306f37f55e6aa01353dcca05bf44e9f6131d497d3f9d13b974d6985bc5b7bae4011e590a
z5dfc49816928876d7866b78c92b3e249ea725229d02773796218701d788ccb3253397e4b21e9a9
z8aa6892e390f0e1f465c1d77dde85253f7b0c7d1bc2c801b4da4b701a79cd1ce9ffaf09d3211b3
z3b42ea13809e48125da6485ab3cf65618387c0fe37cd2258d4bc2c035fcf185935c7243844edd9
z2738a6411815940144978845099f4db50e3c6639483c3a624004d58c838e1063a3d87eeb9d17d5
z081d01a85242d1fb6364826852486c47ed5c61b4e67a58a76de9676267b310fac49b465eef44d8
zd28e811b0d97f25133862e201caf8b48516acea584bbd6161233265c446a5bef0f9ad456c10396
za7ba25b3cc608bc8952f14c02016f2d38efc8cbf4cd3a849bbd555be87166835adb707c17fdc44
z6501e99e4fe35cb74c90f323f86d08ed1b860ebbfdc96cfea475e282815e8ef548778f1925f3b6
zd9d42889de975ee8d1885bd8d73b8412cf3822b9088b55388bac5814d432fdd0dc45d51cfbfdaa
zaaa1399aae4cc0021b030abe1fc9c81566aca001dac5e692d14ae9e34062e90a5c5a9fe0847749
z73772ab70a5681e2777133a117f19ad623bd5d635029d9178065567f6bdb28ab424f81c85cf8ea
z64e1edd1173497d6effcebb8501fd8c77abc8d8e8d16f54ec7181406341b289310b76a3a5ef753
zb030dbf1eb5623107964e63989947c4c42a0b79c90dae57bad4d818555ef01266643efac631a32
zc2a8932a76254c5ae419e30736b86f709959cfb9b0aae78150884b7c8608340daee3bdd0d219c5
zdac293be54414f473336c2adf3d512b8e1a8e3b79d02b0b9d89b31bb3a39ea484ddfbabe665c98
z7b296883be81ae1dc4cfef83af1025be45c009668fc7b2945428a9ed5c1cd6009140f8b1a29b67
z60920aa13678adcb18ecba80b1335bdf104ed0a109b3e0cf75433166ec04874d28f21e2b947367
z67c21ea934e45b4b65c766d6f3a0d9583e9140f63e867463786dc6b09a684a1e779c45e5203cde
z7572f89b8f9e2ee59e89d540e083e42237278520ec544afa77f478a9d9b4c30c200b63a70c9fc4
z3aeea04cd746de113741386039f5462cbf8d08dccbe515ac8f02227880e3c2dc7d5020b0d0d259
zcb5dcff1b00b73e8562dc149edd520cc1a24600c96a0ff4f830cb9bcc5db40b287be87fe9ddc82
z6cad31acba084541a993decbe450b91403b3a7bbf695d9a32772eb2e1ae7cb6d9e827ddc1f7c90
zf878da6b16748cdae44b9203de22aa1492f4d7bcfe361e40352a9801a0564f511188cc3dfa3009
zf95813ace639e5bb8fb4cc94dec2567e737f24cb03df8976d2c4b421be0c693584aabe56d61b36
zc31ebbfad5a325f4ba399cd52dc992349f0e2b2654fd6ed14adc73864515fe481fa7a12b3a5d8a
z90ffd45809f6f1562f2a9dadf0fa831bf59fd79332fb77ae9234f9892ab77e4b016cb996d0f6d1
zb16519b1c1cc48b79cff545e6baa1bca734634b1f94fa2d1d5e74425575b5791d29feb67f72f0c
z3e03c46fa92dab78ba31185de43c92db9ad97b6648e6e5bad87e33a901b9098ba94a8361d40b21
z650215f6cf1b12f43f2087522de5b2678968bc316ee41b25d39b0d6e528b6fd9c3e6d8869a8278
zce34346986bdaf2fbb6e92cb0d8c4ca2b7e049c678ea5c48c23abde7429c31c06bb49a71a84bdf
z844905ca204431895f891320906f05d2908efeb6a13fd9e43a00482bcad6e9efb90603c7a49f79
z2179d08a5a4d877f1087fe1f335196835c58f074451e579729848d752000e13c83b5a34d1115fe
z217ac5e1926287a8765617455336f9e4ae3401532cc29231fa1f2fc39574920c43c8d5ce24ae0e
zfe1de6ef5f1e2fd2a6bd094a5fcfcbf119df7502f4ec3889b9af125df29545d5cd6e391cd50671
zf2f0c2b688428cc700f37d826e41063521045240fa4bd7ded19e82d7ad21563b87dcc857dc7a0c
z3034b9a60621890eab187c7afd500df2714395542ab95a8320920611aa71096acd912573484b93
z64721fbd813b4348c4c219de8dc447f57ac4131622b6b57d17b5959524b0da342d54665b6478ef
z25feb92d3fe5080e36658acf2d7fbee29940abea878a324fbb81ea37b51c4ca422b98895d0d5bc
z59b916025380c7c5bc58acd5b8ef473c97fa9cdb866bee6f7e1a576d65b4626a9c68cf509ea442
ze4cfe793a12fb1d35bfc664e6c7676f82659758650adb0ee1579d1e1025a825df593023495e962
zde1549f36d3f8972e9a2156d92433a8b472c9d6967205cf79fd46405bd8be5bda301d7548a122c
zc851feeb148205c864f30f6188771f69a31111ab68c437637a93c4e8e47c2d5bd4a7e7b92a0461
z067ce6828b71b0ee1eec71fa2f816f7a1717feaa439df058e8cae2f6261417fac83c51e130e8c1
zca3e9e38fb13ad841f51f6b8367091dc1afa62e1829c23c9d72d669081bd35bcd439e9fdc2b9f8
z43cd87dfe0391262b25dc289cbc12e8f4712bebb7ffa3b2df7d7aca5b7183159e593f103adacf3
zec773564df5b4d61df835b0c31190063ab609be66e6f50b7b37cae9aee32f22417e2407287e86a
z4f8750e3c122c4777aa6bea4e18034c9c891872bb45007e763fe075ff4f8f8148670818bb086aa
z9126dad1f3e85583e36196fa7d3553c8449642c1c5bf920513369d9b9d87b443a02af1897e0be9
zc298e8b471f85bc90c1c5b464ca73c4de393485f5f9e7431b7b9089cde461274f69f66c481354b
z74ca29d3f124366b003167132d488f46d32cb21739daa9518aca569f09b4ca48b2f0607b81e0ab
z0a6394b760fb0edc0740de44c7757a736461fb1ce24366b5a5c8223499d2c9b4b208ccccfaec29
ze98aa48af1f3a2d9149f60c0e11bfba8b1c6e61f14f43608c5cf9178ecd38217c41c63ee1066d0
zba9f5c0385d4f1b7c4a9777ca8d8c11b41a8fd7d050097b2dbb9f2cf8666edddf89eb28c3794ff
zbccc5b304c6dcb91eaf355aee6ee20a10359ae35ed763b8349fdb1fff5714afdc84866786303aa
zd67544cb69dd10ee9268a3c30d03804869aba956d97273f377bacf92a84cf0a7c6fb1855237590
ze746e43117d7e543f90209e3132e82ffac4ee1b6430eaf876303b219bde8039f9f989e186f16df
za8f6e1f20e417ecfd9a1c3c759de04d0d865c0a9ec81040d30ad2132b17318ed9e15746b607178
zc7ead4cc33367b0f2c4c898b310b0c6a628cdbd6313f5e178853f21d376bc2cdc792be9438d97e
zce84e8d2f9bdbd8960498dd1cc5f306120e5345c43f7152caff8548a36654bf02954c13b97ec65
z59115c89467b9d582c0713356ba07fd63647469582e4421edd80566acd3018d5a811b346e66b31
zaedb54a7afbe955612ad677ee1584a0d3cf5540d7f1c5423a63ba84fbf206f1c683edb9fa20f28
zf9548ea9414339767ab156d0a96c386bf0a51cdc6521dec609fb2be4f3f60ce68f294d814486c3
z56315a1f3fa4f3e1f02971ea44ba8da6ff017636f7331d1e5ce8235206980c2ae073b723706354
z71e72cd549b648179df2829477c56b8c6e7a284d1e751fc161987c23b63bab9060338a4cee676e
z8b5d24fb6c677c13f5c685883c2c288948c6ac08f1a5f0dfa3e4451787358568aa1cd35afdf3ae
z48ec841e0cff99a01eec9a6840419f251140fac26f1fd49e2dde9c4fae56ff64c09603574de020
zf47735db3b87c3940f15083b09ff3dd8fadab894918c08a2497101ebe5da2498344b3ea4c506ef
za62ede4e74db06d6f26d583c82aef0b1d24a02931ef3e41d832f3e376c6804821e33ec6608ad6b
zf15f47fcb45ed1fbc6bdc2a9ea0e18d64f3ad58daa5394d8a125b436717b833ba769820920dcdf
z6563b224c13e708a149a6fbf23ae1b0e1ab48c126e5813572b907ecd5c2620c29d90026382b2b7
z9adee0703d86f7afb42565eb0f9161e79629dc44a07ed41a0739f3acf36204c6a39545c3b449b5
zb08b158893188abb24886f34c156ed9b67f4101c927c9c0d9c3177eb8206032c56ffd61d691932
z43cdef1a22206fb29283699e30c7c30200b46d0d46ac1feb08836fc6360d9a31c28790f250eedb
zb39abdae3106d5bf3907c391ede3ae943a3051874bb587450b9735de042f26b32258ca0a8aba0f
z9cc32f48752fd757b0090ea898383c8108d0612c2b8fda16e13cc134ff085e96fa067c1c7ea985
z825541d7f70d4a1f7c8d5ad54460176b967cb71e790cababc0221cbf5e847859f908faa4c65798
z67dc2b3d1f6481330c6940bdc49e89b51c3162cbae1909699cb796b1b2d9341a7621eb62220428
zc531a3c53972bdfea6af39e9fba393895b2df95936b0bc5a3e28800e4ab0d5a7848e99f03319aa
zb0659c9f12087545c2042b14ff348353f7638fb435de085b14816f76d765f26d6c354be2a9370b
z56b52e230a253e3b95382f0705d0cc3ebf1c30f6fc47430b5f49521261034e4ca2d6ff78bfbedd
zff67da79f8e56558bfcda0357f5693a6de89529ca5c55404a674f9a425ed695d567b5ac00f93cf
z1d1e54dbd428a7345a82ef1beb4b95829d9f38982fd38bc944631845d9ec7878d0f076cb03a2b3
z3914967cd819848818db35cc1f49e12ace2c4c8c426467bdac150edf9533799a7b5ab50dd7f710
z531f7e8aca2c1daf9f2490d581ae46e4821710208ef984fade9b451fd08c9b3c7a6fbcf853515b
z4ebda5cb3b5990dd19717df43eb472023e014dc0be78322d5bd83b25f91ae71a88d0b368b0427f
z9f76535f2d55abc338b3a5f7361d3a4642c3536580c6b91b92245d8e10e7af4cc9cd3681796917
zd5e9d59a5ce4291501434d866dd62627e92fbdcfd3f319f270e669c57f8ba5de87ac800055e791
z6aee2b33c2db9a3251b02312346c625fd4d515cb41772f8e933f5b784a4c0322e334320b8ca8b1
z2e9d04c023397bf2962f8f01b1477f69ea616aa68400e333e39134feb01ba6426561d8da6fbbb3
zb4ed9599f958ebd553fc91f862155bed9868b786c42317d7534c16768bcddcedfb2f9576e06e73
z842fa6eadf3838ef14b72fb895fa042df23518e342a48683245f66fd8a97a6d849810f018a7588
z26471a6991803c0f06566a82bbd2453143c8f7d40b6e18abd50576adb658261202e6651f91af1b
z5545a7327e6923f52b401aa2005baba6882e370d19d50702ffb032e8c063888a866939bafd1742
zaecbf7dea1a17db1e98a25ee4302c917ad7bb08b8121173165d9bd67b9c959510fbfe44f5b6ec0
z151d52ebd21d90dcf4beb8f97ccd2a2df3dc3f5f1d95387eea33b34e0e9d42b94fc876fcee7b1b
z6baac618904f59a9b1f9ce5e284a1c147e47bddba4cd0d1a4c9537a658baefd76893fb63d757cd
z10a8c5d90cc23d29f6ad2ef040b8bc0cd42f326649d85d5bcd78a05910e36f25412f508f77f8d3
z0604541608e1cf0b64c63bacf7f4ab18742cf9a1b117a00a58e559029b81ceca64e1f4c02e89a3
z234c79e3fd037ca502013ab44b9d6bb0b3f5a245b3b0b0d8560d6aa8098618f7d5ee19207b5df6
z99eb171b396b560de93dc4c0a467e15814095e16db8867cc7c6c9eceec88ffad2b6c022176f9f0
z8d0aec13fa128e6de6adccaca02b8d0a2f8554d10d54026f3d798c3317fe89aa1285a53722a309
z7fbc0d0237c54c5f3d101e4d242a2dc4980494daee7bd19dd6250a103d42f6a079c004442a2933
z079c9e1555c6ce87e925e236e1c73aaa06c0c13b5b9c93cd6af5f1d819f3b3c183f049b25c785a
z767d267180086411aa100419c94975bb0650ab5a01ee7096a1727cc55b659ba1110cf797c664c0
ze597daea21f39faa6245d3f21175a8644e9a34001eb28b951ede5311ec4363d2f515ee0fdedc01
z1a8649717ff31b83d3c760acdd3e1c16fff18c1aedbabecd87b22a6ac1f7b59e86c0617b3ec266
z4c581c5fa8378988cac3fc3dde1ad0dee7cab2a958a01235a45e327c75003ea05d33890839cac2
zd936d1dbadccc9b0e460dd00f3291703680ea4106981a879c4f79a04175404e3d6d1a9b2ba7141
z8c86535b33e815a83dff6da12158770cd5aa132fb85273d8713c69c7fd98233bae9771a367c5da
z3692bcd2b90356bb9adfcecf260ed247a8b8e4f15c7d6a240f2b239d7f042b943b5a2f2592a463
z035716ceffac9d0c1d68c15aec34a1ff1c6d6616da1999f90556bfd76207815064192c966c0bc5
zc812ae7fc9c10509f479f60f105a144f158558099e13cc5baac93e23362481afcb209bc3dc5d46
ze84e7a8091bc639ca3f8802fc909696e226b748fa80640068e3454c4a6e55dbdf1a106b4e6713a
zfd4c38da7cda8ee70455d0ae44f2c3686972db7d9e2b4e3edeb15ea35f9b88e247443068fa087b
zb1f126a0eec165103233a0719490b655449a578d6adfd0547ec1d376528e832de58692473b1b8f
zdf18669b7ca85fae305e8a279825c29e87e0a57c3aded5c58cfa4b1b947ecdde473fb974d41998
zdb47fd397395a4bffce1d9c1723904469b1e50a0783b7acca184084349d792ef016195fbe25c6c
zec416d276803244f706264c44f4c6d9541d2ab6646aaff8ba867e21d7e98d9f3c1f923776ba40c
z43f383de924d0d97fadab7ea172cfbef89ea449cb7faf5a33f6bfd2fc1ce66bf2bc783cf3b9696
z01d0910d2c3f4788a2560ddd308d0dcaaf4c81782a8931c5ae735111bebf3a614032d1effb0bf5
z72588d8fd687874e58fbaed19ce3adba868d4faf30c3ba7cdb33b155264289b8dd3c6e8ed682a8
ze403be3d46b8cfde937b0007e3eeb909735b4561437f0528025317f5a96dc333b144ccb9324301
z469730cd6e11ccd59732472f88bf7b45be584aa2d736fa86929f45ec40ab9881059ff9d9c9396a
zdc5810b4ad8c0fb7841bee97e9cc321fbc127276b8a2f9958f115b0688686be389df52a0c35703
ze797d5294163b0e4e78e5766b677435a06c499527d502fd6dd65e039c36676d1ac07b0f393426a
ze6c566397ad34930e5b519be6ba87e2729c1bf1223f9a3ee1a32981ce20bc23b7407639b77146d
z5f7243b82ad5ac964ee62b1761609f40eb5857a1e431e8b0f3410a73b10b5317f405c2bbca6c46
z2ea7b866fc76128affde46e3c0a53b7df34b9bca43138a2d88e644921b46a2e790ba69e800ce4e
zdb49116ab7af4010dbcd25edc431d52cac556b8710962b1af2c618b49296831c47f3cedcedb638
z539faaeba757a1418d1ec83f80aebae24433c77a175223afc6223c460860c066a1e3a59e7c8215
zcc9309753571b848eec126beabb3bed140193602647f484665042ac63a8a961b1274145a29d227
z3f55fdab504e96c8e9fa800d4e3c68d313fa382b9001e2e771c7715d3cbd31f1adbf024aa27452
ze82d0adba6a26b8b6d4d39cd45d7f69ad895c6bc15203d0ee8314a98bc545122c742f8c2ef319a
z1ad3fc1a0437292474374b1977a0934d9f15cb516f3150aa1d30c11ca5c08008eddc88f3630583
zb697be47c34ac948ab53dc7fd29f85f75cfd1dadcb21c3ff826cf775e284d588d1d1640613c1be
z4913778fb3958f3f73376bd79f7437e1c97fe7a08135c62022720a444e713a2d8b8de335ec5fe7
z3490b4df9116b3707e629beec012c9045217b44b79d61923aa4682777298db4a649227b6134093
zf278441162e339adf5ae896a0e8fca62d8962c9e7f3be0379407bb7c16357094189f3150cfb6ee
zd66e5df578a573da77a5d3cd8ccc5e88cc5f896ce15e5099f06efc80435cc4fab8709805eb072e
z69699c651bee145efaa29c6d6c504753de13d6c6c9757d08d8a9bc725c7f1b46628cbfed1ea2a3
z2b3b84585d7623589cd8ee01df33a334b36cb9fa63a7c2ff1ada63989cd5edbec6a60aee7d9018
z726e6d51fdc6fa200f25569e8a3a00de9cab2664dd38a68105aca8295a05bd6beaa7a9ffbb778c
z873f87994ca6ed1dd32ef5e0af1c547ca0f31b9c38710a9c1b2deca42a004ee22bf8df6d694e9a
ze42eaee60117edf5f0943b8fc46197726dfe17575ab60cecc6335e31f0cd2afbe4b5734545f3b3
z5d271cc02b9ec08880c34afdc7683681ee1e5522c6fabc86d4ecb3bd9cc9271a60eedc3bb3850e
zbeeaf22a7cb854701d4a99329a9a9754b70dabf5230107f706955b72d594c7a570f77b563d4abb
zde2b57c8fec0214a60f81b30caf415eb121639ebb859ec3ac8a76cf9a6354d8f80a715683c5dbd
zbcff87aaa94ced91b5e71c99221eb52117b149dba4d26d449e3f83181d2748c3ad5c853e36aa9f
z87604eff37cc846db0443e61c6ac5d36cfd00718a24f468685afbf4d3fe82c7bd839f6942f5ebf
zf307da8cf5e6153c0acf57a96222a450ab71e172ef27053e5c7479417e19e3e3bf68825d5f67a9
zc9b4d9ee98d04de8d5903d083cd07fd1d565ea9b16150c5f5b6dfe3aee922843352dc57cf47b93
z3b50f4eb7af794511e7ed682695e65dabef97b7025b3d458cfd174c10e941878eaea5ccc3caa5f
z7cd80defb1530e5d66956fae19f36f6aa51768ac850a2f74df23f094abddf90346370a823d4424
zb92bc1bef9aedaec9859d15965ed41532418466feca1810a160a34005af0740aedd25306d46940
z9c9eda2f0357353f871d29be1cbe7c9ea15e5102d6418eae5997dfe9c169bde35777b6472541f0
zdcacf08555771ee9d80fb1260f019230356e9c3247c2b4a449ff6c70b6d1d4630fa6d571de1ac0
z3b73c98cfb1c8b0adb33020f93ddafce16d2dd631819887624e64a5795e03a1fb7d58591ff9df6
z2fc6167a003cd1d6782dc1d1866375d972d84028f1c02293c35d5485c18b8ef8e5539d8c0563b1
z6ea6c8a9707d96755e0b820ee6d662b26bfae80ba1eac119aaee162aa39f829f734cefa136412e
z908c85010e7675f8d6c11293512cf4b007c5eb5ec091113c02e0389b27ed0561f46e9f48d09da1
z78b187b63d2edfaee8a394494856cde1e929946cff2da693b75ef68a4a9116305be3be2dfec959
zf08d2a265ad75d77a565f313909a7317bcc4310850d10b98c04935a8e22fc08321e7789e83b68a
zde38b130f979a3066565ee01a64567bf6c84ccedf46f65836e1a84ad7eda6c9fc7224c34c6a4a4
z265df3596a9ab6585a0376045ac1a401ce1898baaab21557e9773d659cf384ad9e96be765ccf95
zec74742365120c576705384d507a113426193398872462ae50f6b23eec602b8d33c48799ec3b3d
z81e52692e25b48c907ed752b06237731c890d30ea814b4c1305ea85789d37af747c4a00a32e21b
zfc1567d2b455023926c3d6f58736c48533f8044803ba1ef9a3869ffbfd84cf49029341b5223bc6
z871aa3253be5cf3abf62da2d64fadcdc0b18ca0049aba7739af1b7e0dbd6033bb5715213e2d294
z5376e79d532fa687503766d68d5161b09b4c676878446e0d02d45c344704bc536ca384c3948b1e
zfc873913fbf504a5fc0676267fc7804b9f25d11ef359e6f0275f69b594fb745cbf9e817c18c2d3
zb455b6b4ad952980d5852651b7851b84e1bc12607e5db1276c69bfa637c9c8015ccb8b56acdb8d
z42e7427e7a0c02fa29fea33720efe1fb6283de2c268aebab495d4b2731c90145743446f4aa4b65
z572948482e027ce19d70683f127f6f63e4351092acbae7e3979a983343d0b5d7e9b3cc243590a6
zee6bfa03daed1a75d31a79ecdcb520f3722a5b0a2bf8b3a51916f5300d749f4adb382a8641e35c
z3734fdf55db29fb134ae4ca05323a50d77086d7bb00346ccb56041ad0a661a089a9d40a09ef981
z13d3adb71fbb97ffb8084323fbb251177621a720d5cce0f6641e71dd88cd1e5587a3d54703a1dd
z36b6fb974a7aed170894db27d9b6d81d4273bd68433174f85c13752fb15e5f7a03daacb4f1bce3
zb626fc3ac62dcb35542d5198172e3bd38eff13bf1dcf147e1b604a1252b9e43a6502126ebfbfb5
z77c9e387c80843eaab4e8f142f5c2090829b61df6cd46771e23a6796e6c50d703fc48956ce1297
zeb640231392c6c650815b9304b00d6a75aec40045af190f2ad6b3690997c8c4d21e4fa3a90e9a0
z6a39482f03a991d3e2a2cee6686ee8743fb740326d29c5d2f7be00c96860e99ba317fdede08a6d
z4df02417ab00df5d28494821bd81afeb464c25da21271d4ccb2efc0551c8e6c7b9c96ffaa9aa01
zd83ee27e4331fae3b3a630ca9820a643a628ec7bb203d86b244d8009ee85199197fbff764dcde7
zf4993a7ad11d66e6278d3a2a163b5767e6e81b0fcb53c821f62f129ca4dd69a13e9cdd441af91f
z33cce41fe5c57997b666f9241884aed6088bc9d9d5fec541a99ac65c4380562b93bcd10e37191f
z144049dfece40bececadc85078060de3c58fdbfab9058d4c78ca709bb5cebfcc4d26405f3d389e
za4c3eb9736b175315e6479accc04f35d446980177d8d5ca0050255eb651e6c7f1071a85f7c7fa3
z7db7a5b689a2a97c0e5dc9ac762f93ce2ad4dda86e03577f197f67e154a5b0da481ce53382b73b
zcbffe38a38e5e2372cb42576f40da84a007dc3f60d56952b172f0854a5bd71834149b1f7b44610
z6dd3d0535ad22823ec8c6afc964e1cfe66d77ca6230d5636401ea66e912c741ab65c947429c65e
z05e49784ed74bc3a49d8c0b2da4ba23971a258c0e311a9be4eb3a28adf7c373980ffd218e4664e
zf6b9bec7e1ce81d1c10da596fdb131c79585dca85eaed19d97a2062b47985fc4d327382602f3b6
zb49fe1c3c6babcbc1004f93b1c90fdf49a5ac34bdb234d38202425fb3be601ba6fff3162e9d309
z35f6c81f83d7c4604b8287194b382e5a01a8a2984a9b0451a32973a613b7605d111717a35e4c66
z05fb415324cbcbb00e65f2d9e7f31e28a325252151ed851b47da0e8bf61f1d4c94064cf8a7e943
z03a8bccb5084b289d808cd6a2ced329001f4548eb2aea3ed90e61e0371b36776ddd2892fb4b1b3
z4b528d67bfe4e86720428cc2383aededf5d052f4a633a825f7700ba705b8b0997064bd744e3ba8
z8e786c958008065de92a38a2fe080dabded46f1ec00f5cc27c703f259b0e7a91591c15e645c3d5
zcfab148af086e18658e18b184c7838c9b0334ad14fb0174835850a6c27dfd98625881a26d1ad1b
zd8fe3fd010a923b22ed146728de80c823879d46bced638af87f3b9a510e841111cc9c2cb7ae2ff
z967c81dc533e588f24c98cb49f86b6561dd4da6c0e540873152699453b7ee48e53a4b45362ee78
z4c8afe3a0b172773de60d15ad7086264afdca2670b90f083a9309de9b65119109def0af68acdb2
z4d283d15784951573de4a92c1390aefafeb469cec84d955ea21c075451258daf67fb5191f47351
z7fb6a49b05787429092de357e977ff3e778acaac1d0aadb4d8053b61a77105c442ab4d67193a9b
zd0acd3061f2df0fdae8a4a10c25c91a1f816b53a5b7b71462087c5dbdd1a0dc614b7973e26fcfd
z8afb60e177f04dabaa734b471273d748e49c760e79df49d1ae02ba96f6bc65818e3892a6b9ceb4
z2ee896163ce56a5086f481e9e14207d3cdde3f58c93ba73892f7053c1fe5d217bdf38efdc59ab4
zb141044131c8f7e467177b9665b064245a6cae57c698f131dc43e55266695fe2fbe5c08ef7672d
z9468e90d708dc3b56e1fdee0da97a2ec7bbe3c4e0da0b963b7f5c89c66176fc21b5e839ffd74db
zdffcff715520d55c586a7c666f37e9777a8ce0aeb774556fa6db121d42ec83cdadf46f33fe0419
z422a8f799dfea484cc3048c2f6c39da455b5f1ab657a82644846cfecc9ecc744269039e1f86c41
z1fa82e4f031a24962324b8b46c582e4511fe4a73b4e0658866986aca000ea5bfebb0b47e30ee32
zcd7ed3929c28e2a88d957ea930e3c9d44b364b853306f0e13bc90d7874f885ba62ee2e02fe3f5c
z84f8c70476d90cc8a1961ba8015dc7a122ce66957e7a53c3def8612c54dedb6d9aa0f452bb60bf
z0130649d32cab18c8c152882dd18f464a10be3df4de03b608256bd29150cfb8db5997691f8ef2f
zeab6523e790a6a559e45c99cb4d0a8746356ef96a427279d4c02f02a69bd863520f84347dbbe15
z99b24fd80316e947c8b2671bda642e84e3198a00f23729b48e0c8f30566648e9a418d017f5b72b
ze6191037586a9efd2110e02db2437072f93ac77562cc81efa63deec3ca579cbcc58074d7f6f0e8
z84dbf43742ef8a681d42e8832f626d532372ab813d6d65c3ff49287a2351944d293ad5e3d67a8e
zfad2dda992529a2d07922c61d98d37c5b51b6b4a650a47343baf43232446cc8872ea156bff0c07
z75e1a08a239f087719c15aa52aef1a3831057c40fe34a8cf6a124f1808f92723159e213c5e6002
z00600ae41c3e647f4b74b6be711dbe782e9960e8734a31a990b2c5211a9565a06d584de3fd3d41
z51045658e88836ab06cd3a06501c05018be58651bf399e6590ab36cf3196929af7aed660b89c2d
z8a66774157690a83c4ae15b96de425af796221efac7dc7d2207769b3fb44222c11fc48182027d4
zc801e7ee05d695e59ffd9f37946da2674d3e5a48f904aeb360e2e61778b9b71aee253526c8b1b3
z7514fae046a337e24b8264859bfca65332307e8d8620d5eeb0629d448b3144654658f10ddd67b2
zcac0aeee71575d9cc0bb75c30a895fb5f955efed7c7f5a67d58b19acd7137c135fb833553da9d9
z4298d8b22e006e1f7a26cee464dd165ab277cea68e7aff4dade13bdd726cb3a807dc479cb05127
z27b139096a7a21c3e28f57ce556bba7e087e1e611c62347789be198acc7ac852a3e5cd6ae3ab4c
z3858362e95ca58e66784097c858dd3f3f0200f1a844dfc0f25abbd52db0751ad2d0ea154db1a02
zdbe33241529fde581c4944cbef16cf0383be4ed4e017a557c9298a53192b65da6e9b60cd926834
zd0b572aacafa76d24ffcf184f48610daf13422e3c942306d91a20206412da5bfe584aa7e7ed580
z8f3463ca5779526bec2907357ab2fcd770586857a784ed31806d71370e3fb9234d18bd31348433
zea836d15c890ab5dd4d65c0e53a6b877ecf696927202c4af7e8135f02b4661c1c447468b25fe80
z90324250638053fbdbccd761680a351e4eff5adfd9e3fd6c420e193a4420b2ac515675a90ee305
zee6c8303f952f2ff9bf41d9de41f54c18dc1ee2f367d01edc05e8cee6ed5bee3b277486a3d033b
zb193357f81f9e839bf6c1695b49c8300b373dabaca8f9c12c177666f946a4dd68a14806bb9be71
zd3d50c747ea5b4712a57b154b88a9e5a0807a2f49c5c763d5b690d330834da793120030df1aefd
zf2836bfa740e6ae90be6092262282abb240c6d37fd8f074620c8faedf128c8ce0708ebed611ca2
zcf410dc699d763cdf45dd5e67a038dacc75b1859414e131e36feb5761e77380dc37969056f328b
z084974278c0a4c8233d61e31122259139b73bb1be319402b3dc9a7d84fb407ed3cd0640eb9a9ee
z05dc1847d2ee6955b71a8822c551c2628138f3ffdeb000b0cbe2021675dc6475f05bf828426f76
z0e62957593107cfa0ab103dc30c1b1f9ed3ba366aa88c24f7ae05eba8864fc3fe2a870e1a354b5
z2f94964165424b9cd324b1f265a670c66b96ed3b9f9cafe285661c4f9c567bef2b6463f2fc6d37
zc76e1ccc96716ede6bf51ec4077fe5cb44b70afaff72f8b55da11993f3527f6dd2c050ceca62a7
z257351bb6b6de9993037ff5d8ceef6b08505103466c4de076396f9bb4bc5b6c0d5268ca2a9858c
ze2088c1a89de775a91f72da22fa6ffd054864201250652db2e4aba96ea14760940dd657cc29cc2
z6485acc0a42301aeef3afa6b62e9a342c79d7711e4ace12536d481efe6c085e53945d8bacf855a
za7b28f05e2951ea033dae72597202948082877fbec4ed891add8b89a6a9b943e1e2087208cac70
z839d99f5557ebc7b92b7ed1686bcba367d8db0478cdb0143f5b7e3cda7706239642a7c57f866f6
z12c3a5581042fa3d4fcb4be43c9a22a7a08ffc8e57e5a2ea7e0ac6a4372c0d70d80bc996dba607
ze07d945dd6b47663bf9a3e219136cb043b6b3d03abdf79cfbb4bcc2419c56f642277b51d1ed170
z5d34f02ec0c465dae73fd39f9ac633b04a872b0d086bb4703094187d10aab6490cd125c2fbd895
z6aa76e53df0e226e866b080e16aa365e97ab3492380bfd30d3d333ced5b0a1dc1410e9da2026b1
z6f47af2be85bbf682474dc2e9964b513f324d20efe245f20036c17fa073efdc1434decba365f67
z75802d7cc92a0f75391a4c36e38ded1687a7b4bca65b9ff9dbad7999cb0545a1b8ee8266e5a634
z69b95073a8afac8ca90be8a1a3ec212ff542864a360bc83a7ab5161fa9c002921bbfce0cac075d
z36caacf3640b7b438bb961ae9c2bdc276a9e3a4b7fe1d68120c1867d0e76192d4e3f47ca5e87b7
zc3a98452e0f9e1d3b26586c67bb14cbaec18eeedf6372bbea899722ed3349fc9bfb6e9b6bee043
z6cbd719edeed01e55cd8dc30cc358210c80ebaa5ca6dcfd8ee0cd82804a9b9ca9d3b48edc9fd33
zcdec4a6925c93b835ad8d569af17931433db4b6cd698af84308eefbaa2369c55edbe7173212eeb
zb5bd579c3dae1a8f06721b394c6bfe49425ce57f0437d70b9b988528ad114f175d9b092b4afb25
zf4793719ad0f08cbc866fac1bbb4ceab6a95df4eb8971f13767259f9887f9b53742def15cfd9a3
z5601b9fa2d3f3e2c11756368f041ca005247dad2c54cb5f663a5c9a8a671028251ca8e5dc3aba0
zed680d2617f1807f4e874b2f69003ea05b5fdfb2bc282538770f83c9493ef2ca32a2fdd42a148f
z0ac3793d40b749f80f2f3ac415a00718d5a5cadff2c882814c1c4b35f9093c744b7acd33bb19e2
za98142af23403d03413e9b7668a729b4cfce7daf951b5926931502f3311810189add9544b28eea
ze9c5a94c49c35a668ebd47ad7b08486e44c904a61ef1de74e58c477e65fb033b8af71e962bfee2
z6d5ff4b0de3845b3009fa69644073c101c4d1b585bb05164faed4137ea3c98730999cd7315ed45
z6f1032e97d624272dc0967f39c645c7f127a17b3360b5416a8e6837633e906b63e95303796a3ce
z63cd892a0d54f0135478292e09f0fb599870c72688e02d29f4ffd2e94fa6e0521287f88fd53cf0
zf01fa987064ddfeecb6fa5d7dcb346b4a4cc38c4c16c49f5c81fa4399f9a3edb1b0e8f883b0d71
z43fb20dc443349a6fd334757be6a35a95a57808ee53d0d4f80f4b8e74c337a33db5dc142e2094e
z85b5a3bbdff8399cfe8ef2c65a01bce04d5b4dcdc2d108888c800c588f33cde53fc0b86bb7ae96
z8a00fe9dfc3cd7f1cf63ccb3999fb0992c1e089accb91f58ac8402b6e2e4d60d1d4618e6a14ac3
za897243f51c050c5d3e082a5c48f5bfaa9f01ba29087be5b9ba12ca6b48bf1678c347d8a802b73
z5a11dd03cc74d3de494410faf5bee2961b4b99849594c1252ca2d54c8a30b82ea6e5181abc969e
z9b1bd0fed3a9f6921cd4a27eed7b45e24ca9cca98c0fa3766c741d4876a800f01dec1b35fde0db
z355da8f250566b4b77580a22da3783db022debe99b9ac74be945f1b2467d2835d020059a6ba703
z742efd8855b0ca5e9feca82c526b1cf1be737b492647fadc8d97f7eee8de178aaed45e56f5371f
z50807078b135e2abe7e308b9966058551a221e5584291b62e4e146c98eb9b15e92aac67a5528a1
zba423f41fdc546bbe2bafba87caad6e22175d42ba7c27a1ce8da2367d5ef8028985c0ea3a02eca
z6e0a31835030383f8fb07d97815b63fe801d290635f88dc740236c3472a633c0811d10e9854b5c
ze46e46b1cb6a34cc32be5880545a2fc890bc20ff013c9904b0e3136c79b83ced99f28f563ee1bb
zbdecef2ffda825c992ed484ceeb2b8e15877f0f8ade6c5092143d66304da3de84a78be3a846a64
z4006deb2644368d4b6a93d3a271b7563f0f4898975551037104778138d4252b87518431e54e434
zbacfd24b139099d20bf24758dc665c47cd0ad09b013f5a3b425a92ac23a34bc4a3b1556352f3f5
zdf5c6b84074807bfc1d904c053e2f6e2c44970dbf3784720cb9e2906182c2834bab83dfe7508f1
zf276bec6907a29f0ec74abe24c73088f9ec9cd8e0d8f8b5986ef42cabcee91412573902a9575f3
za1151df6569adac9b1a38fb6c26352c79e64762102839b188828a593986f2b18d5aeb7100f8cec
z8bf60d3835367e59c8ba046d33867fbafea10cc3ebacdd6ae0a978a36394fb709296f274a1e0ce
zeafa62e7231db085db130d6a76a8033b3b47a962b5c7dedadb818cc36567e32c023d164349899d
z025a561440d9027376f6b330a63e199010e6a93821711b704c387c050a9633dfaeb630f7e8ad13
zdd20fee6fcf30c7b6cf0ef80ca52b8664a4484d9e367e12bcea5aa5f5705ecec66734c1f26f8a4
z4966b00d49c9bec0e9d68c5e9f2b060b3e3a64fda780363f2f363f9f9664bc5f073f8aeaaee40f
zabc392895cdbf028b3e4a3a9be88408574a836c6aa1ffc48f794a7985807a198fb56277737b4f8
zf34f0110559ced9166c6240d99ff8dbc9534f299ee10f2605f2bd4fff588846aca652e68a16098
ze41998729547b1c9c2f4544ea3576f31d7646c58441f58751972a0598a022f6ab5ee293823ef03
z75f9494d062c3f9ad155849c58e2d317ccfe5258ac41d3887cfc788b68bb8faa73ff1b2358a566
z8e25928435402def075948ef3d84f43bd9b6a48d28cd975780824bbc88dde6260bf40753264580
z9ade98d560bc445242352843e060a08eef3967b2297adbb545c6cb7982c1470bf07444533fbbd0
z119b625d531853f0b6bb631296504cb2dc6c6ee76800d676b9170ee611c346aae80a95a3fecf5b
zc93e0b8cffcd1532ccbe1cecd9ec48581431fd007a36ddff085082bf3fea377f2273ba81f42013
z197dc857fc16e3a8dde8fe1daba3d29bf9ff7d6587898c185db9869d0a9a301e1c17de3ce97cb9
z14c66c3b36120fc6eeffb40e8e5699b6f401b8c33a259f561b71cbfebd17f1ffb4fb5270728121
zbe618e2ecec612d749429f2c08cea3c98810c4bf055a7f8dc43c0a95a5a11adcc13661fb9985d9
z29b34bcace0b6a93210729908f10f6d305dfecc5f9ffe481206833b1c44ccf2b71ad2c49a71d15
zee12dca07d0969895abf0cc84b34cf4fc9ba8cddc5064ac929e82529c6811ca533d3d8820a964c
z58ba91ad02e502649abab36617642c460aeedf94e72cc3014999c4bd183ffaa6a8c08c32f7db42
zf134212d7d52cbf4935095f88d34ca7f1f50d7dc783d8db2f35b8c50b70f121f6f7a472a0d19de
z955d1f717876396b19a433a9062aed99271e0ddea8f28dca28c7b84ddfde89f9732b65608e2500
z7d5b89f866257fa71d6a2fd07b764946b7aa2f173c60c1705972a056edf6edecd8959070b56600
z3abc66b3a31d62d08a8cc6c332b4fa778e05e9ad6cda7123581654f44b6a3bf3d109030040e858
z1db9662b20c5f76069cc86cd1af9b7f08d8cf4f1790831732b3c0f6d3422f149868546830b824c
zc8a4caf80ae05543bbbd53ac2fff47fa449191de82c35a9673052e6a8e8bd4ab12b162c36a92be
ze3c01f4948abb97c9e2e77f0a9025110cb1a4fc5d56d1f8a2f53fb5a23c51e73b0809f6ce1e770
z440a2e7e00cf6ee0caafd03214ca3acd0ff2608d45908989ea3f31a200214b48f419e139d5fd9a
z5e6df138965d9c799b2030be4d3da3a7610caf9212347a100c13cc01d8e10fbddd03ee032e88c8
z8abef5069a633186fcb30e4160dfd70bdb264f42e587ff95fe820fb00bb40a7e583460d7ef7b9d
zfaabc10f036f24261b7bb2e046b32153554327ad07cce8e9563c61904e7354ca2036aa3b4395f1
z67149bef9c6e999333970cea4da1597212ec8509c84dbab9f7dcbea0988be68bc2b1458c30fbe7
z342955395faab5c8896d0fa2cc187423a6c498203feadf58f39ff89bbc9b2d008fdbdeb1d6a998
z964bc79dd89c3f4278eaac5e6e3183e1ab23189cdfd3b9c9962c8dddb9342900726252287c7f9d
z10b4263d7557f56e7f182cd011599609654f8f281511c3bf4b1b0bbf72c70058a11931c8993685
z8ed9b94ca0c4c05949f48536590c20a5dd32641afe22bc78846a1a56ee6b88bf67808c495149a5
za431a104451d288a8cf99323c022a63f0e27105afdcedec982276da53fa09ecfd678775b20047f
z0104ee906fd650c2323cf5b95690a23180f5ce037cff7c999ecce3b5ee6b07a582954b3e235082
zaac084b55922d39f76e78634cdbf402c7b8bdb3915679477e3d1df7a83b3c05fdd0d89778b7fbd
z1e1b80e4f5251302415e0353da4d8fc057ab0ed1207f816810153786b76636c4750330c5d21ed1
z7bcd8dc5c1af7b8d43c637f88237374b0b7e20c47c3753442ef067536ab740e150098ba6a201f3
z17eace1627b409b5df7460731e334e23fe4460cd8c600f8bb4c5faade1c92cde2dc527b5cb5233
z1d5dd1ae532a369aef437b38e1d3fca33fed6c0a5b7ab217ad0a5878eee1db5aa3eedaea965429
zd62a6b05bbbedaa3cf0342397b4778a16fbecd5b1ae419b41c25e6e1a3b5e46b3de02ac7ac8754
ze56f78b3049ccd0b8aef8e3f18a3baa7c3216764b1e1676f47ffc548c539719f70a62975d7edab
zf36c6efe02b795a045ddbd96238a939e84fbd2e822eea10412d48a9c1e1a03641a7e9c4bec3548
z2ca23aa758f6e02d56836fa30c850ccc5493aafef40d342aacc43b57bc5b7e21a75f248e11e17d
z4a148c5ddac21c797bb56a3e46a4e2ae1c5c9312862ab77c43ec932251fd7bbb5d4398a875ae5e
z25275d986e5c491745239c24f427aa4d2362b2a4a6af5a901da9234ba2aeb27a662370d6438af5
z7f6c267f875dd757b0bb9e3937df066c37ee7257ee91f79c3d9a21b938fe5c110fd68583eab298
z3f424a15f96ba5e6eaae4935675851705beb1881719568f97f3f577f12605a5181d36ce3c04255
z5dcc68c294ded8432de6de33fe091a36486e43a9f91eaf617f2ddd57f07926e3e374a2cbb8dcb1
z40cf3ecf30a265b1266db62afec7a229894d1c0df5ee3bf333a492453166a6189731092ea176c9
z7a7c9429ecdb1cbd0ebfc1772ae75c560dd1660adb308d0af9f70cca43c0558550e1b23efe7335
ze455dfd12720a51ca7a3951245c87c5535e9b9cd6c5e0afe70ebc385cbb10cdde3cebc135c567b
zd9ee03a9e9b134675857a9b262f24c82b139920f8512725815f3984cc7da9559e7eb1aea27704e
zfb943e2cb363b650e663bb6ba0e926ad1063ff8a3d6249cf762f30cef742e5474da0cfcc7b78bb
z36eca3cdabb2b91c5e0b5c6923acfe4fb882eff1e7f8a3f784d6b2b08c7d3e24b44da9e0405e13
z31a0abcc98049669496434b127526c7229bd7e5d90224a6eb0480fee0540d5a971c0cac821082b
z9545fa638f10a53be0cd633db7ca65c4f1e8aee1c3f97ac6bc4663a145050523de970f718b4908
z64e438f3a033a62c424d8fb237592920a21aa11ecea872f64d24cb03b5959d627d4b5c7249cf98
zaaad34f915cddeffc57250f157ddbe440886488956575c82ffecb743920cc74cf938ee7f9cc605
ze9f2ae2e329eb6c3966dbcf21d934e75a36de49c656a9aa8d3645ea1d6645725c4fd5c367dff98
z6d3efb00d7d10072c8a477c9e3f3384ffa19ce71c056b029716a8163d4d2e92574626990cc35b2
zfa9ad4a494e77d5afea3a601f85870eff7df10c353b1bdd4569d22621a9ab97fc67021cd3bb619
z3f28fcceca8e3db8cefabe797c6c1f879178fcfe39d5f2c1e88e56d5f9c580b11968450d26d272
z68d0a0d38ca1618ce0b9d00d5f7daf5bdb068ab974d6c730ac65ea05b61d3f71bc93fe9a17396a
z8d1aefce19cedc23c4ccf88d82164cb2f9ee18bb1af9b2b4403075c5b78a532a1cf4f0977e84a6
zab071c5a34ca00cf022b257076a0c7835ef4663409eba6d507ced40db2c65343c5f05c07b4f87d
z7c44acb64ca6b2f2926e0341e06657abcc58d7eec38de4278091d32fa694032a05af9103cda9d9
za8a141ea5307fbd09b46d1671d6be35526cc64f5c5560736791ebb1acbccab778a48b7dec59c63
zedc77d078b2a248eb21e02efc17ebd99473018db1ff8cceb162d603e4162edb08fb607c261ae23
za5b884e4113cbc1275a9136b7793437a5e6b5ba64ded9aed8af576f6177e7148147790b67f03c5
z00015d0ae1e442a92a9dc3f5dfab57e33b40f3bf18fff1d35eb697dcc9b07425e256a9e4f77496
zee12b85e610da44facf7f3c0f7c6f926813c632ade57e174371fa7e04ac7f1076aa106719ca879
ze6efc355a648eae3823e7b8dcab9e45f8ae0326d19b0f7a32dd34e81fa436187c7d6541ce62b96
zedf996902aa048a4745ec4e81823c0d778c40258cfc7e932f772b833319ee84110509df2713626
z6d3d6557166622540ac0324cf042dd4979698214893eb2544ce4c7b8c36463732e8b88da68f193
z2a30cff54f797cdc850472dacb17ce0f524e243b9c8ca8d6fdcae67b39cde2919c3cf963519bdd
zd2522e869a90fca434c06cbe8119c132a66d81e04844cc8d836579ef7f6e04b86977b52b293b5a
z053c54f15b8846bbfe2115598454176f03ffb919a5c90391e73dcd587e437ea4285e1fdddc92c9
z653b04b11b902119261cb89c0dfb23a75ef28d916f5ea777e1c3a8a69297d992e6f95f07c47102
zcef0b7eaed427dd747dd45232f14fe5d395562c30f9fb4e33d566ab2b67027613d882c6d6e3d77
z047981cf8afe57e9944ad3b56eaad59ec14d2edbb7a0398274c35cef1fdff4d58d6d540f1428c2
z2fdfd297d9350049627c0c13590eb04a748df7010e6bec602fe8ecf58aa78f3adca5e8bd1c6ce1
z0ac6b1bcc24500db87a887079604a1feaebecac28ce1502b7cebd23474b3928753c463e08ad76d
z81afd17a8467988ead7db2943f7781dc2a05d0861e6d466cc0f59bbfd8e8fd9ae021b94146d06a
zc502ba8837213dfe9910323667154248831667bd20e1b2be6e49a45f8c9ad397e1046bb07baecd
z670fd17f471aba547d181f2e948c72413ff7758d9fd70c05e894a6814ecd5c3df72662348d655e
z014ef017842642b84d98fcfe0a527d00bf7a895c8d5cfadd15677afbf4e6bb428a3b193df3a867
z9c45d652d873b02266ab19052027ee7b2d791231174697e9af7bd30f03e109e50d9cb1ae5bf369
zf1b049513253ea6200207dd9e1f97eab079ebb55bf4cc154e35367f1318af821cf5c61534133be
z1e0234101dd5a17a6d4d7742f3762a18e70f2ef25c9726e284450011f7c7bbc3994a0235df897a
z9e7825171fdd73488b7a4a5d94d43ba16508ae30e838681cc088e3452f426da60931194ded1818
za7e557f7860d865094397c2a5fefe0455d49745e5e0f41f8ee01e6083f0b677c15be8c8bb0f958
ze5679411bd12071791f635292037ee8eef00903ec9ed8fce51146db713bf2b01fac4b562ab1f69
z4b6f0a490cdaaf216ff8d91677b3292309fac566d63965a9fd517e62a5be4a856513f4650f46c4
z613fe96f33dc2af687aaea87254c3257eac2a25fcf1c1db15ae49de7c3cc3dd4623dd37d7f04b7
z6efc29547b5a8c140027cdd63723380d1ee5df63e791487ecd166eb928170e50cc2f89a889e93d
z3c74c4e7a97cdb4fcea5af90a0a49ad282fefc7548996875139d3024eddfff5ace1727c08e7ac1
zcdc571f0401947ec6911a158e95faab5b2966dcf8854fff12519563fd193115a32935a345766f8
z3eced87d9411b11829273a80a998a93a628b121c2b51a8a37816d8dec08b59e0a5400bbc2b6414
zb0747bd3119f552fa0824b948cc3796c02ef164b740f8d8b4540a6eca32b1eb18672d991124abe
z1f6c9176dd198da629dba32596d1d9115dbe74b706590431a1483b97cfac10cfe3c30ba984dee0
zd76287ba674543c3f9b78275e751c91797c26e47233a9f20169a7a592a9c589d16df5f18adfee3
zce400d2b1066145d9dc2b8d910c2c5b66d35208681c2c881c5bb21992e34187c746980a29ca48c
z434d03f9e91bd9a1d8b84c3d2a0e2c2f9dd20098803d8aa23970b8a377593c20c5b6733cf66964
z5272e8b16157d7ca34fc7699066e3a3c0ab45c136c9b9e07df0983a73300c8d7270ceabec1340b
zb1604c4f9e078d358a2f1586d5e4008b0ba2f3b9a9d8b75831953f2be2a43cb18b9d3e32e904d6
zb656bca4fb6cacac8be7ff6ade04199a524bccc540d9430f980c92b4f48affd6f8689f5ef7c6d3
z4933e12511e12a087a4e57b70d7a4c54006c9654b4a2e78fc1b485785341e20acf8fa54724c4a8
z398d670b85845807d797f6ae348f9753e01f0b688d1132d8b1bbe23a82fa1d6621adef541d0e00
z04a5aabd9a8b4c578866920ae0834bf0ee49fc95d7dc4876c6e44c6d1d1e8283dcf14e41d48c9a
z564bbfef4ab0174574c21cb124b4489e2feb908447eb7bcefe1152ca1d569595b7f6309c14ecf3
ze846af2db347976db9ff0b606f87d8afbae36339a077cfb23b467d5071b98c18bcf74519260cab
z45223455498306f247a44e056315bda7720ecbaaaa2ce80fabba615de23b8ed30006f55a19be08
zf9ed11106d976e31e8a8e9392af031c731fd46fd1f04ecbca0ff2b2e8cc560602d5bfe27d8e5f9
zeac33267e02727af73a26895ae97eafd19d3ca8192fc368030130f2381a94dbfea653139c0379c
z262708338787768f13566b6f8dee375502e453d01f3bfdc571bf1af21299761567ad0a2a5ab3c7
ze849b9e50c3a15b36bd8e75be8bca996a82f33e83b5ee85a5cdb7d0d8412eca1251209348dbc69
zb0514f4026945869a764cee7d0396780af10ae9717337f10078cdb245678ee8b92ea5b9b88ff79
z7cd6a01fb94e59f260f5aaa545d7e2c98730a18aa5a97d8061860d79f974c202054d207fc945ba
z0477846c285234b09f44c6f0269dac378f23092d5c269ffd03d65b07d6b6bf8964c293d0326e36
zb25a455e595cbfc6e8876fe63da627e58cd650755a717bf26ee7985571dc97500015c8606c4b17
z410c5b8d5c42a33f002e2af29429cc70f06a2070a7a5d5bb14fea150d27c104094c0422f074e87
ze8179582bbf4171968bc84a74ef0502a773d6d25f57bc5aac4581d01bad76ed7f917401029fa5d
z7e85948b540afcd3009087e2763ec387bbae2545047771701dffb5c60072ba0b6e422fb87e661b
za4699e81086629a2425b5abd81201bc3000b6a951c9a7b14dec4c6a9e8470c1665042511a60909
zd67a504ebbf541bae7f4dfab827f77849acefab768426973808b84e7410c481441ba39df8579d7
zcf15063dae4c1d864ca8688a3ff390206b58bbf30d3da2bb9acb47e2b71b618c4783fe8b44af00
z0444da0ca3763ef748338621a0af0e129c8f117341bd55aac2dc0e8815fd703b13c643d7defc98
z0b3a2b9375480190281a87118d46e50138fcb6776c3a10f7b953cd8846b5fb45be4535c49568a5
ze2253316ec69fbdfc8fe63e63b11e3fabea29d3cc052455e50b2ccbc2c00caa2f3f7e97fa8251d
z13135d7a55c3a169b92789fe14cd51444785258b07b501fab28d8242342b2fb1973ff01f589b9d
z60a8a272128dd43ef69fe759b7b9a273722e3efc2de150e44b9505bcd687117707b32dcec05465
ze9febe2b858bb6d02514f496f5e66a975cd97f158ec532c6e6a819067d6d4d8eb004c74a9c1482
z844408d3d7d9cbc6e7aa67defb36f383c045cec91b40c11ec39864b3cf8f6b5f9b29e587175b6d
zddff1d8c1bca9831f79962e6f4dcb856f9f018137d730a1e8100aefc3b9b18b0d17bce8f7b1d26
z9f33b51d16ecaa6a2480a14d0449849f62b0f800ea60f9fd2598665dd919f9370419013c3c1c87
z88c372d2c637eb4feded1752984293fa149959382368ce4da4a1157da5082a40233e6ae71e1e6b
z9abcdf54f39358ec6ea2abf73679b623bee1f56d8a28e5447bd81266b91cf10398bd7d7fd3bfeb
ze149841962429f072c629196e8c23f5c83955dd002b8d69aea791e411254c6c794caa25d794419
zd4052509602e0c6866cfb27e85055a0fba9dec8f9d8e2b738ea05b7896031f64017159c5dcfbb1
z461480f006f8b260d25a3796fc88d20a40d8b7637b673d2dee38aa9eac69c144e571fcde2d3f58
z8e77a01d9e25c7ee6df4eda8b251f0426b42620ecfb743c127cd3c4d116efcf04f7a660fdcb4aa
zc0ee4561b1e56c1405e15eb793125253ffc48542e6015b1615dc436c0668b4c97e4d48554430a0
z5d06174d9282d5a5131b524f1a152e7ec4b309b4b93786b2a3ed8f871314fcca8b63bac0e8c1fd
zb3dcad97541d1b9b6d1ef003ad5a88c04eb26c84c6d10597439c09d4f0895431cfb691ac7a0821
zb820d622ee050ee350d17c03594c66d2991ea32a4b59e225171204e0e4eeec86f843c132710d5d
z0ea96624174cd919ea5f67820932ad1b0c96847c58a344b020a9d2c0a9ca0abb5a71a6d33eee25
zf6a0fcac8a4cd71eeb3aa20a3f2c3e83dbe332af7193154aa95e9fc7070278185997af57d4fd77
z347a7df8d5de497d5bf14ef8353c1a90e474df9958dba76e60767d11ad971d24ed4c101689a805
ze57f0277fc6d57904c2c4311cc1e70e6d45669fae5a9de96d9254b149288efaab5660836e89798
zbb80b21bd405a7082ffd43c9d57607692b95269ad6b7e321582903f9597ef3568dd67dfa17e973
zc0c6f97ecdfad9cdbcd178353922ea8d2ba3fe5c76c46ab58c133b0b4a13e8ace0ad66e83e78f8
z8ac87c638f4ea3be7b676ea43c0b8fa26aebb41feb879f8c18fdfbd2e227f13b46b09fb4d5e938
ze5684c4286a3efb535b8fe96cb9e1421f0e2dee135f5f4605e41fab81b321ac756a316f93172c2
z60e62ad788658cc48ed9ee1359916a22b75670f9f56318e06a26a12d649b35e783bc2bcefafcf6
za0371bc9ed1b9e239194a40b3b2f4991fb97a485f767f4db6b0ee593d0cad04d51c0fcbc5f43f8
z3b72fc868b1566e9f2e4f9f717a3c91c90e09692a9fb41abfa7520cf1718e3b4d369fd4c22009e
z3914f0cd7f2fa6a3677a06a3260c47f7a613c1f7e786fe1f5d41424f8dc6e73f48e689db0eef6f
z42c82a8ac32b34cabccc10f6e586867f45b5af0e8f0f849af1f0a50981d4cd9f122427d53b0e79
z00aed4f06140eda4655025078aea39886a2006492835fc4d5daf7e4c3773e6be0e9eaa19f8144e
zd21905782351437a560eadf95db741ae07258dbc54940f74d7bd6f5ed606714870d2d406edf52a
zff1a18a736344b927c6b05c67f30eff519ff4aa8f981c7fa42f390490c6f99799a4a0040795026
z39749a3355b352e2608c643c7df7b9aafe24dccd80d115e1fcd1a698c0570e994ccd6e8a626a54
z858dc5fb11a6e2540f4e1f6d19f08b48003935d0f589e717cd6189b7d22749a361a3f6a64cde2c
zb2959362f101ff5ea8cc9c8f8129be63bffacec6f0068724c722823686f72b5630b33e891b2744
z2c44408e4bad4ca0ecac12991eec74f40a9edcdef28318d6dcd65f9f2074967949360bb8910377
z057b386daa3377281b07f3e4f2c6ee81acb97a4ce6c55553d1d969d2612eda371d405dda0ec186
zdf346059b5547d0d50a6674db92ae9599125357f477dbe3a33be9503ab63c51902597feba1e603
zb65e192dccacb015052d527deb3b49f558dcf9a338570f2ed05bac79ba7f78dbca3a16e02593ae
zee8bfd73e7f0235b71542385a4a312e1011ebeceba95c9dbf6dd09fb9aa811bedfb0732f257721
z3565598d32824091bf7dd49f2bcc0897194108f93cc8ab035482878e1cab9188fb841dee4ab82e
z9d69d3806e95fdc06b57e5c03c9a87b4196f57d79c62a345ccf69e61db4569ee23e6794b16da87
zc29de71dcd9bc976a4ec27b4164a2b18d4bfbf07eedfcd68875e53ebaf9c51d7daa26e37185173
z3b6a2314b333d2141a4e3790e19da739b9a249733b1b4058a92041d74a83b340e829008808dc7b
zd98e56d1980391fc3ce08f17481ff5c4ed8b0567d2da525d4e6dc337ee4c7b52932731291f04a8
z8da20160e9cfc53a55ab00c6963a42ee798ce2aaa995ecca52b0897e2a248cc450be17449a8ea9
z75e41e2a9e262ec2dc85732aa91cc9e170772f8223162412813b28477ef5ab3f5eb3c8ecabea59
z415608d6f7892b61dfe026290969c4facc591a9a3eb96ec2b7f37021ded0840863065c60137c14
z76033ce06102a6f61510aaeaea2c7f959aecfa686092efd28044d108107c321d3bd426dbe80188
z8dd290bf9a98232f6188af60fe87219c942c0d25f11b57e590fb0fad52a2bfcd71c0bc10c45ce4
z83c529c2e9a4a926861313a8411de5692a945ca56ab877ab4d1d4a15afff12e252481da8cf9ff8
zf7eb367dbeeba41fd2f5a35e1b5be74a414b7b9897dd3251b20c0188133ce0fcb9750914d6a802
z7638c7f864fc90e695a6db3547b3b9919aa07e6c502d1fc47b74853b266789b0459f167cd2026c
zf0151448b2cfc0e0701ee2971008287ef6f3ead9d5201f0054eb53634d4003de348b28ab4e68a9
zff7b528d19ceea07b94084c0155c001440c475b0666059a109d3ab3480683f1a8082a2b9c5002f
z4cc47c289af03ebb3bc74211f2ed26307bfdba549b71820ddcf6aa8a13bcb92f0be164eb241cf9
za3807c110540d91ebc2217775cae5d3199460bce0a34dc43f4968fe568b49837baafef9d735066
zc6a9c2eded2c055be2e380d595ffb231ad88610eb439fe34eb09b7b796662b880fd054d5e7be9a
z7a1fd9833902b0f85e5ccc458c1dba534ebf78baac0896be5d62cfd7d7eea90b65ccfea2a9ae50
z6a18a561d304314079b0307fb4ffb89b6efbe5bc29a87cc9b257d51408f488ffe35667920c7c83
z0d6b6cecc398ed90fdb7c90775b352239d4160ca0c11c14071ec7393e776695a5e500767db7cac
z1be70e3e2fab15266c530d74e6f9a8400f5dfc7d4560cf4e48eead91ec41942f4f48f520c58d55
z0a483a9a61aced0d7e0a6142e517f931e700bbb4fa12e51603a6df249522e524de6487dc8d9eec
zc0ad26851f32bb8ac013cdfd8b16496178edf95970d262a760da8eb6c371f0579cbffa7d55b815
z1f80a3e0db1362aa3ad9f0282b6c6f2756e13305a70266db94a0d8f8442df1ec2716b707dfe389
z522bb2098c41cfd6a3af830ff89e3aab1eeedb4619e4319070df9ad36df0743fef80a96e06608d
z6285b921ef43045a2904358700776a2951db0bab4bc391879061e9a94af736cd99c5ff472902eb
zd7ad28da51d5384eaf0ff5ae5f143ac5a11a40f20862b17805c466c2da8960949737815f646b5c
za5586d44be3f90505ee3962a7d9abe844936f3881dc648e9e73968e443b2cbb82919192eb49fdb
z8d1bcd4105ab428819d183a3b34372c4cb7411129a78340e762e8a28e7e798e9cf290f3881c196
za03623f8985293ef145d1a5f76c439273b0639db17c97039638329a6454b8cdfe2b3c402ff7ebd
z0027bd0ba467fbbda46a8c2652959e4447925a2ca0a00691f3421472584e04db57f430134bebbe
z172826fd2f5d8b6e178f274bfe969e9e66d1a66103241e0bea54c7b8390aee494daff6c7b6b875
z98d6f240a6282367dab0423180d1453eab096a32c920b0fa17cd8a582a64084319f70686fd9ee9
z6c22895eada6e548c7171942c02df1cfd81ddfc4dad0934301111917faf28f6d22ba85a134bd93
zdaa08381d9e10f9fe0976720f5978e94a0286f0f203599cdf845a95c5be34aaa6a3f0600b9879f
z5a5262cb1ef7d10eacb20a8aaf81d2337b312a8807fc68e7f9857186d8ed0c2a959f2e5de7bf38
zb34b1fe64518fe16130401ef4258136d70186b00cb64aaf5e4a536a95fa27731f51e57ceedfc54
z45a7cd711cdf6b167897db9009d8a95dbc25a385201d2c95dcb71ba1725acbdf884f190f7be61c
z986dd7ee590682e026c7963b2d5646dc9cfa7b68c9dd6902fea06dde61cbebdbfa0fe556052c9e
z8472c7c3bd7ca03e2a84fcb488d0aeb03728ea85a6db5b9a8859bcdde632ddecf6e9d4b7124e50
z23983ddde9e8089dd4356aa3ab63a717f861cd774575fb6d1b3f1872a91f4fe4ce04219bdd7d15
zb76cd15339a60ba0d3f9567b99069bc045d25ed1e3af5879986b77c10ce7e92cb724f2ec0ec85b
z24c647b5a9d6b0b933dd1a38cb70cf52752b6fd9114a1a1746caf8454e00b2d48b5947d6160e02
z1d1a8d4a2bbef4922532a178152aa9ea8440c13d6d714dcc763aa3fe1a034351f3a734689045e7
z6073c35da1538994b9e1039bcaf97fe847a1cce9771652b0251a4626b74beadb8167a7e8941bad
z1398d8a54f946469146b56f2d5b0bc3b74e9abe9d1c6f845f5fcc3654ec60b43b0078bf430cf98
zcdbe114e563b9cebd2e0734a6963fb4744e40e07f0a6b08ee4b8471b8d45be3a954a64d5383bd4
zeb10187783c908ee24893dcf7886d4b269f44b5c2262dd4bf56391bfceb259dd7d06a4fadff0a3
z7e84ec0f338a4e957facfc71209877daca1f088fac202d35cd4f254fd57a0103415168477980cc
z098835e490109ee820acf69b91bb4866bab338dfc4219b4dbc68ef828f5ceb978b3ff8d8a4034c
z444ea1550030eec941933bea1f3878ecf3740f64e50b8075147dd71d797c50d85526ca4abc2d26
z85b33b5ec694bfc155b1acefe78d897132e6cc87c707b5e9ac0c8c7a155a45cfeb7f52d7b3e352
z442853d16642cfb92842c9ed5d8142313f95bb7d55bf0e72fbcfcf50ad8deb31e54a7f2d08cc9c
z832468852130b5a94624cee8637fcd61e4e6460a0289d6952fdd1164eac9deeec09f8757e030e0
zbbdaf6a7ad7725ef8836b61db69b8ede7afd9e33a7c1d2c8a9da869a59ea186125a5eec8242b57
z04c2df32c2426081bd106fc28a9230cf150e9c5ac96decde040b222184a63c889b5996c70e6cc8
z2179d0a83dc7968c4b2513dc2118b498dccca8117d0de9d4eaecabf862c0944240425b2c2c5986
z4ce9e1481966d14cf3441c766ab2b93fe4da51efdabb7d0b6034267b33958ed8f4e01d09a666a2
zc571dd81b7985c2100fe0d3269abb8d60ce5b69d36a7fa4e2dfc73bc633bfcb69d16a77f1c03fb
z463ef1522f3bca1902bc5433d8198f65cde2ca68ad3b27a07d4c5daa3f8fb6d67775913eb222a4
z88235c2d166947d3ed2570edac3edabda82a535c1bc5b6a0f40c5ef04e934b5856f2fdec36881f
ze4e55fe9b032909044353b92aede0599bf0e6d6a99ee3568af207cbaa9c1d3d2c4c25c07af74b3
z43c28b1036e3f983a5a7674b9aadf400979b128a9d3b84b109bf525f3537fc417631de780bfb97
z0449a897c2060b4648048d77ea59b7d457d7df285aab204c3ff726b1f7875a918edcfb1bbf9b9a
z391803d6f82bd8c6a760c55cc040084ad80e31ec3bad8cafc7a2dee29099c08831b70d6d19f1e0
z2a077a17e7589cd654f76ec7a2da50abe67a4623a63ad4efc3aef9cdcbf00482cd906babb1e5bf
zd533b93839941860caf40c30dc4a97e6c5a607d3074609d7a13ee715307177de0ade7dc2d308de
zf971f4b749f8aa08d8953d315d517bd816bc368b755bc965e8d09a94eb46a71f77950e1fd3ebdf
z16fbe1473d58cfbd3f711a07cd4eacc01b4c4dd97da5330b5f6f013fb3a72db2a78ca0aabbed33
zcd80858e720fa51217d67675c68e8df5ebe0866163be4f0b1af5ebd5febfc2c7573a01e602ce52
zd9e8af6d6f7f90e80701f6f8b923168e98f46d69d98449cb889fac167f85153be8d32c296c2148
zfcecf479a9e7cebea39c959a522802526c1ed2493df4797f81bb2717c37c9acd35cfd9c9cf9bd2
z0d206be1607612c3be43ff39200ee75913813079e47c1d2efdbef629b41a575ee1f7e20dccba50
z31766455bb5d144161b22aac9f7dd9efc99a81de1d4db63486c67e94a51b94b3a9f2761ec615bf
z3b14f3fea9ee9d9cdf3e65c07044adf0d8dee2b3bbd92bce02ca758445cbb9effad5bee961ef76
z2575e3566b72e8cc0c4dea41d6c6ba1df0ba474bc23d3a02e1e0aa9f9374a580065f0695db8a6b
zcf560b49726c30cd59dec68f21455bc122d9da2197d46c3a43fadb837e3d1dc1971412c3248089
z0ae035ffb44af1618314a4b22c059926f14262c73aa3590601d34358097922161f3f8bcd0bfc21
z8f2ca1ba38c163b5b0dcc9d08059230be52591306446c390f41e66fc1f2d926795c447be342595
z5a3229549a503bc2ce6a180d952593413262373aaed7d9791bf243707afa6af7858b533c3d0940
z49f99115afc6d3b510775e70b8c089aa744f1d06185c0742cd8b5914e5715aa7990c9d24b28df1
z198fb82256d8fc86382242b32362b446b0b6215f9006e7f79103be9ea0ec5b53ac622eceffbc27
z0ef12d04c37aecafbefc6ad736f4f78379328d7b51278f4b1288ba3d9868d66d74530a40e6766c
z1a664278df556407255b50a7c7ff0c860f921776f0a1868df3443a780f24fa5d10143517b00020
z703e779369e6024fb0b27c14242a2c4e20ae2d1537b0cc8d5b7d7968600c7faec279ff5d9381ad
z84da7fe96b2296b068f8271d6f284599c6a4f825c81c7e63f5668cbdb2652b19e9df51f35b76a4
z01433fe82432fca2b36a4fbc374299211a6f5ca01ddef0a90a087b56fee3d312f0bec868d7b302
zcc7daeaa269a1bd05e7caba992e591df0d6e928ea3cbc99dd2337dbdee3ca7fcfd8ca1d24add56
z52250a1b6715827dbd530045aa0d3bffc256924c01202a5000bb772339f3f544b224089c5a8d16
z8f9abd65c32ce88b5c658ea9e81abb9e73a8d53a12368685c54e1460b03b5a10f767e61f3be99f
zcaab5d97b3ed346992f633ad9cdb0ab9dc80310c0705fe8bed9a6a81934e31722e35a591f98b16
zd05761868f892c5b8e2c79ea5354d3bce1925e6df540eb4c2bdcad947cac1565fb79b2fcc7c4a1
z3570ab4366d8837ac1ff309eb4a839647237a7c804534e4cf0ad97a955a1750233886b63416288
za27824bc382444596596e5f06ff9c6f92eb6283c7f5f2d1524cce1378f22c6f86ebab502c9d02e
zcb5f8eca2aa4c4d112827a9c6d95248445b4c1475a457aede5ffb44b169dce6e6f2dfd22303e11
z9b55bb6fcfc6e4cd44ec31f50e59ba786fbf70c87d0f85b8c2de2c6fe1cede40a7c0dab0171225
zf5d9c192d23660c85d89fe10992ce379c9543657a21704fcb348680a130b7a8fcea26c18df695a
z6258440ddfd4d3c8e127a9f8bc113c1378d38f59f6ee980cad551abb8343dd7d811fe6ba9e7000
z34326119bb3382e30e375364c7f54c31d8ddb42c7e9450259e09ad7ca39c8c296488e73e2506ac
z1a4973a3659e48199426486ac4db5382c480ba089104d5d1155cc16849f5f16b2c01935382624a
z7277834b6d71b6902f65d0f804bbce239a4c4c5a55816d1730c712bae6b5a09b4f138e35040c4c
z714801fb4d1ed674c7cf975972ac7fefce225fdb0d8fb436ea40f86cc600ebc058f2e646e5a90d
z1ebc175175158b471bb51dd2c711874c3e0034eda329bd75e3c5ca513cb5266057eee7dd0ac348
zfd9ae8b1996b37c4d440c71cc5d32a8111c1d5bcdc79e1bdedfb1c12782577084a0ead10923775
z0360ab9e59c36bee912e412509715c5da63a279c39d1637cf675605c8fb8b0037e77cffd754c70
z4e2fb60d500795c07a2ad108239dac3bbc49f5f11bf64e78bb0be02656e513f3d34bff5ff86ca1
z7ebbbebddde07f3623c7888604a903fa32ee732f0ffd61a56ce62b750917dd1327de920d9f512f
zbbb2faba2d099b494da8fe4069a85cd3a00f6129e9a8fba7837422aa7ddff18a35ce7e5d68cbef
z51f4e74a404e862276ce2349fff2634e9d51532c67595735dbec5fdbe494dd15ac73d43db63772
zd548479e18dbf2dab764730ffa37f924322a1798dab8a8793bd022bfc9be14baf4f26ab169b0e7
zc76c32fc0f9929223aaf1bda58ec97bac3b05035cd002e9b6000234b3e7e3d607cc7bb20f85cc4
ze32fec17a23028ae0cc25657966b6782b1a60da107316ecb7dff924b14b051cac3d427d081ade0
zbd402ec15584813661f2484793c13e4c1a954099dcd0de8e8d14448f90697c2295ce0b5b9a73b7
z1e8031dd19791f4ba7e370d5ed45113fea528d5a81cbe9ecedf60ec234486cc3adb3f8acdd9608
zefcb0054419f6e848d9753cf03dbf2e1887e2b81782fd81f7daa6c448df6df38fed41f0d430ee8
zf25d35ddfa5d23f933247e6f10699d97766cff683c3878ebbab584139f349e10e8fd00459a4caa
z3be48f48fe81bcb554566add5e2a125fad5842fc8763c4fcd247162776aa0545ce60e94472a202
ze9060098a67c9f17b3bc0b636cedea8b2c3888bbd72c23996a1b39f5d815423ab73e9df51ecef3
z9b15012d4cabc63bc36eeed631f1f400ac3182435e9c639e3ea80d226c95fe314454e2a8ce98e0
z30c81e87e4bb6c5cdba1b9434266f0b103f1e05ed3ce69f5fb8a91c589d512dc020d97453091ee
ze8755ee35ea46d496a965f5e576c453b8053df536d7c26d992ed60408e779fff6042b401625485
zdb88e19f8a67aa9672cd1cd5a9495c5358ff4087473ae641d77d804a94fd51e9d92371ba827f84
za39365e9b0fe7d2f1bd8129c0c40b083cd6b24c08c5b2d7bdafbe1a48fe281e6b4466a49f34180
zf80148f10de137f092e4c74f53e538427e258c6ac712266bc7d01dcf4b042b96c6a45be11a6335
z179209cdb9f6428299761ca0f4b94c8b461fd7862edc0f8ddf0a6a89c97c94f31d097e95a43227
z1a2dd419e273c2f0e0539496841aebb92a0784a534694260c7348b77205c2045a48d4acf1155f4
z0cf3cf1a5da98604b05e694edd60f7a1af4d292557a8c51de40904929223b81732528a7630e9a1
z250e4cb8c29f0293b2b43e7903b4fdcc63aa50892c398da9f4563360e88eb3f932f4e9dbd25702
zf2e9955fe36e012be4be445be27f8cc1e6f1e528d4a6484008f385a73c9198bd0ae8d3a303674a
z9337168ce01f64ffc82737a1b25870f2dbb821591f2937d3934da6e92956aa13d733ccbeb41a33
ze589d2c265c870452416284466dfa15c942d5fda4089cf43a29d47752c32bc378279ab736aa4c3
zfedbf4127b1e5ce4cd2e1ee2179ace2131126031ecc6fdbb95de192cf0d03bc500a9da1773904f
za730285856ffd1fa65a94c7d0d048670eb2f7a8445ccf1f66f4cd735021d305e4c9afc92f3bccd
z14a6864ef63244fd590a019a923b4220d8d32317caa1df776c452652399a0d4742bc610cd4b344
zc86a904891aa07943a371f389ecc25416fe6758ca548bea2a17e700c2f5dc369a2a039d4d82988
z9b55068509b82391919a25e4db2ad11e3c4a7672ca2921819c19b121e0cf80a56dc53dc1aadf5f
ze0ea6aed8b98f12f5a3db49d306c556525bc24dbfb73b3f273252c6b0889b949fdf916190532c8
z1a9c56e3fcfca42986680ce1f3220456797d9ceffeef32313dd02147dba011ad00a6d85ef2499b
za66616a77004c95ea36796f5911475f039e7c73a8b5c3f74a8e88340533a4725411ee0cd441013
z382dfee2adea871334d01d2798a8ed22bb729447b605fec7d14e81035277400681b37d1043ce2e
zdec577ed99bd6619c773bc1b054c538d6016a5b5b654ef7ead1dffd6942d09431c171e859a9115
z1647f43f8861ddb256127f52407cd2a38feee172af007e54fcbabbf262dc00a24ae9f10643abe4
z91402160e5b5ddf10e415273184a35a052d74e5f21953b967b698e66ab448725896a6fcabb68e5
zccb409b71b6c74cad181d0714eb1b1911221b275cf258b76829e86b7643c5c4adea5aa54f80228
z0b455b2ead8223e6934d767a7426e0256430f16704271277609226f57189a71e80f06fd4362d27
z6f0c7991553ca04cee85548a62d7ddbd3c216eb579ac508040d4cb2039eabc94cb3172702cfb72
z778c788914cff4741b478a7dadc313e3da98c81d6a35737779f2e73d191cfc3a1163347393af55
z44979faf256f81ea966f22735324e1ce347d6092a4c9ae2cc0c4ef3e35d48f7d0e630fd7c261d6
zee9c9ccd96f780d27b7529b04757dbd5b77957153e3cb2ea4c1d63a0bdd9807a4e3f34a9f10716
ze7c8740cf3f832064306ba62e7a433bd071e516037a79800f059d31de8f6d0d3d02738b187fb5d
z1ebf84eb964fbfca455cdb8ba273a3d524402c92c71d24c082ca334d541fd2ce92bb1aadb941cf
zbb9d615bd9016c6d9054247ac8558545901c44cfa98c3551fcf0a89f070a5e9e8973a84f88a6d7
zd5423b04c5ea8e2693f37c8c78a7c67a1fe936ac0d838a2f23dd55a18484aa10aeed80da1133c4
z3ee8194af8eacb49b1fe1b6f7afd4c453521d0a51e7f74210aaa76a985165c8f8e6e40e50c9f41
zff83774ebdf9242a7c4ef88337dad6ddae7c5c37bd7905415a472c6eae60c794fd6369b813d9f4
z7f41aae33f1d5730c99ac478b229c25874645ef71197a527d20fa8e61dd20fff8cd4ae4fab40ce
zde36369dcc0fd4d0ad38ec24b469c6a30886919ad01b65bbe40363c9e4c8574c408eff7b4b6d93
z640c65be1a8e0c383f88a61ecab8f5efadd79893b6e97b8038f52bdf067df0fb88385849297ab2
z1e12ea72faa28a79ab63367d9965fb24bda24c899fb714328d12916ee5cfed677347c9c62b7faa
z58b9972042f38f677769935a5f9ec4ba509ae9a68444ef705e1cec3a974fc26b2c0d500a96019b
z8fa7c917eca934cd16ac5b1c4c9206ca0c26a01c2258671b169da1fe0a7f8a1f6bdfbb5f2a1c0f
z320811e603454d6c742f920c96f18c9e68560052b6cfefcd418d171d8a5bd17feb979df6b7d425
z8e06642471431201e8c28c5b3c707f8a0e5cff30836ec4150f99fd1b4c3e2130ef4a02cfc2d792
ze32094d37eaa7183073abdc512f56d4a7a4eb4109ef3dc61d52bd4aecc01c936a24a0f040d88df
z5cb32565261cae2b3a784c84a3c529e2ec6cb8d5fddeb900783a4915639ad147666ab8c3278ff1
z400ad62a2985954279a37b3c3610b3cfd461610b1207173d3e6679c5ec96ef3d7b4ea1d9f4f8ba
z2ab6bf21c132f83a54577dc19005cbff7bb35175834fb8c447ce507d82a594a40ff30587754ffe
zc2f7f804d9dc9a0abb56d993066daf7087b9efca3e58591eb21e30dda1047788a92529c67d4046
z4727384357412a7e08dd8b4e64ff35061cb0d162b8226086d296013a3df81dc2f2c986b5639f12
zbc77ecfde0a8fcbf878bc22675fb4fe19c14632bb7c8a0b3af0cb1e877782f1a1df0ee4e759e24
zbcf9eed731bb8390a6c23dfdf2bce2593d2b47f219096730f2f0e33688e41ce198d1377a807850
z68b145b975b2a26d837c04f9a60bcf9d9efedf4ab0862d7618ef52b22a69fc534aa4cbc46d2f68
za7e6562e57a85f4277e36bf97d16b246808282a0945ef7db411f3f7f17b9c081ebb4d26d5cd657
z8c1c6fd0d00ebffa60455185d4573d8310cf71a122edd196c7cd6484cabbd0a3263c707c851cb7
z1319063b09fe252a32a5195ed0345f80d85ea84907752a73dc132c9000ad19ee74417d268b6b22
z535ff96541c6ac2ea12ef64805b59f106ed7c377ff27e8210736d3d1b8fe7d4ca16337e07198bd
z3106db916272e530deb611ab93ed67e09a23f175982f622bc25e345efe2523ce79ffba82405d82
z8bfeecfd3b160066c24352b444f450a051e1344cb1d97ce1056dd15f7a1fc6e68f42cff4516328
ze1f19aad8c7129e96fdb1618bde58365b5f9d121929560f388be05829edae0b0951679f8bdcc1f
zf2afc0a1fc562b978cb83a6084bb6002ec0f70641e1eff1382a2938ccaa8c89024fdc8f7e9473b
zd130e98db188e5d40ac3a48840db4bfeabed28111083ac487367e3f424d24843e957f2a28ab4fc
z8fe950d7cfd0e85e1eb7d2d2b976e27e40c1a867f594f29905cd5173dad3f44b3a088f81caf092
z00e4b474e5f4efa7ada1d958ba7aa5f72d5c025fb8b3a486c5a18803a23f417c537374e4ce99d2
z71b80432cf9686b3fd90ff3660d355936e9fc7368a59fe732537f78b8570b431654d203d886449
zcfeb3f72a869de4c9563194d3a2046e835a68a77cdaebe7a9751ee3754c0a83ecad4954caf6fd8
z4c432fdb4bd96e16cd7d8a08c9f5a6474294d98ade3cd59dc71de5ff121f6434ee5ef9f1eb34d6
zff21555234ef8b65af4475e28e96a5303b39245d365ffe9fc59a59f598c296662c772ddd13db42
z899961a3609998082e7374274bc72a3b332e330cf5697ee7bfc14cfc3ce5958dd345c51e90a7f0
zc884f133d9154da95e43dcb99812763c713803260dc07270a165ef37e799f8af148ebbd689bb71
za007178270c0cb8c20110f9c0cfbc6e05365e7e9fd003c96099ec4e0a10a47688de4e52b6c69f9
za5f3d1c9035e1fe45d22fd25e9a5dae18067c00fbda586245f8a7716e969d07de660ef8b541ea5
ze4c417c96f68322e39047cfa38337ae874e6b4998f519ea752c686bd1c6127307fa11a9b1bf3ce
z7b093348f991b76c3fe681166929da92239fa895eff1d122f98dc597aceac560d49dda4aaa501e
z569a57db49a0b1f6338d9ba9cbc3f1bf5a8be46848f4b9eb75
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_ocp_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
