`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da33099ba6084c0bafded292dc1
z85dd2e3925edc8b79302536c5a94d857dfab42a4b162c335c207c17b63516c48d4fb6098b4cbe1
z1bab4deb91641b63c1c6e839880afb896158ee4b6eec753c1e96af4a0277309dea144f991d1dfc
z09f66acaa3548205c8c5b56fb9262aab6d7342d4ebdbc28ebbab2ec720a3e3a6aeb6bb1179bce7
z01201d7b7bc3293cca0e580e41f9dcf625621115ecaed1676acd74dbbb4e1eb6d938bd7d0623fd
z8fdc2be2a165dcf4df0bcb9fca0fb694ac9e5ad772999f9b5d3b5d0768ae325f0a449fe4e5bff0
z75a3cc605721b7c45573e454ac78103eec590598c76c11b4018535c7b043ed21ad10a7392faf50
zea2c690a79ae2b70d7dd7ccd523109eaa19213bc5cf1a2f25c34cc93b273aebbc82493fa648fe1
z7241c2d2fffb8e97cab5f6d213ecbc3392d62423bb80e3efa0d0370b44fd88dde30a7a95860ebe
z529e24f3e8a0b84d039c65f92fcd51a2fcf1fd715a0f9422d39b372b6ea7c96c564b7fa462a756
z11d3c1b99c86def28bf847c01a6c2006be57987fff702cc0f6fea705760160bcc8f02b262cc916
zac1146bfadc54317339d191b00c388a569aa48459981cd1a41cb7f4cd63e025f816517eec55320
zf78e1e29d8efd08d023b9678283861ceed8c7412e0e3b0377cb1059ebbfc7db691415c925dbc2b
z0b5ddecd7a48ccff9f1de4496696edee1f43a0027fa2b06d60671fdf189f0bb4d5caa162b08128
z0b196e2bb737d64f22f1745cf348bde0caba59d3c7eea235427a12151b593a9b299b39f7953aa7
z028bc53cb23f68b0edc02ba16d661b6e9ae807d13d4471e3acc8481582ec0e05a40e0d5708adbe
z61df014578ca91a42d0698561a245c3aad2c90efca4beb54323f81be5015685560ed49d8ab12d4
z5ef418aed3a1c1b08e3402e0a6d58e599c6e50daa4b5b8c01164e4c47bfa3537a993e70191f056
zf43e3e6463f69b49eee83496038f76e86555a1a314a0badb9d2f579b29d76b76f86c35c6af55e8
z1957d56803083a52080e3c5f8f60beb6c2b344af7ed2401c762cf29f8c5dd6cbdba491bedfd94c
z102e63b29ebeeda75951a5a601e2eeeddc9325b6bc04f6ad9f291ed0379b754ccf004723933949
z21fc4e02ca679824052b47c1e0ff2111b6143926b1e869e1d2877cbdcde3a1f65b7c3f9247ce1c
z1499f9d298960920bda547116e5496cc8d3e9a70b23d90bb5dd341425d138cee8088db7ae90c1f
z9a1c0f924bd5a6836fc25ea79986ccdc541c78cc2c92b545bf29237c4d623b5197ddc7a97ddd9c
zd7cd45eed91a3dd226a6fbcfca8811b66b904f416505e59c4b43d6d934e1407d3ccd3125005af4
z3679d81fb3daa32f6f29edf0b6fd8ef7f5f39e1d025e8e7b1ec2799d45ef169f41fe187e4514fa
z31f4bfc56d1ab8dc1869215018bcae2188de65a41b1ef99847307e491b83189dad00e2ca1cae67
z92a4aec99ab9a7165b3ff94a7cf8e7bbaeb1aaf2f268b8432d87157df17ee427272d16576c4357
z823862d80beec19b3e38d41ba585f58316015e47b8a40579c8cceabff310168ad38247bfbb57dc
z66910687cf28af235ef93f8a14b7774ba8ebb9977c725f02d2b553ea8722503f68602a72e12d9b
z064c85edebe54582c08822fc0da8a496c7d2506f00c13a832a7a557e95f1b7574986bbff8a1aa3
z32cc62ebdf18b609e4303424aedd4d3bfa4e4409b58842712e309d38e16e0b290251b1e57299b7
z35a83aad96d952696e49063b7e2eb8ef95b78f787f910e473b056d6cee97b90822d881b35b64b0
z029b89e2dc501dbadb6a83dc9e0169534c1ba65c0c37c878469402f5eedbb0b4181844381d4589
z458689ab558ecf879c5cd7f17b170355c8f78e6b8f82a03c23d624bd5087b540eac495da3c5496
z6144333a8dbd544b13bb8e063404418316e20171d114f898c440092af6b97d576c36d56248f08e
z08e5838a9ab9be022ca712478bf4870111fd53dbc82c464bea66528b867acc3383138bbd21c642
z1eb99747608aeef5f5c5d949b9a7fb37e62de451f17c53096164a372cc42957818024658e44e9f
z3a976f777d090a71512c7982837db7e7b5c24dc930562ed10c5b1b0f803f3e5bde3651fade6089
zdafcc29cad5ba7e334c215e6ed0925e6bbe62c3b010cb8e5387f4841c99bc6c11176e90a62166c
zfe36350718108639960bfe0513b7812eca215b651a2b75734fdea4945bbb5f9f566f361677345b
zb8e25cd081abfa25d5cd5dfd134d13ad09ae597553167eaabcc501bfc199805d3335f403b2fa06
z253de82062353e75946b5eb9510d0277efadba805c257041120459249a9bf809abace2230642d7
z73a0a2c63dfb474f5b63a56f894e07db24be5dc236cb1d113a39df6b0467a1d92c5173f672bf03
zbeb46e128f36a30879d724efa7c24aecbf789a63211a174bb8f1c0c5bf087db960386081dbf1c7
zd21905a38c66d172e185f8d47c240738fbd3608659017de178384be29c38a537f826232b5111ca
zb7cc528dbaabce4fbcd3a032a83f5f310f553a941e612824fc53711a89c33cfa1ed150eb90753a
z9a8aa8e12eb301a7dd7ba3a68ab404b397af5fb46107314952ed3f9925286472d0e6acf356b759
z3f3a98667f952fc13bcb220e0c76d2327b1239c49680488d2d0b03752db1ff7d7d71e8cdeaafbc
zf717778343887d0090d80b0286fc38973dd3118b44d31e31eee4869f32566702e1f455c618d55d
z578c368ecf74934f23a8896e6113b60c02bac1702720d1d4b6798832df473ef5893ac4076f9311
z1a0fe62e8c9b9f9d7caf2ff3cca426e72d806e6a61550c531d2e85d269d11432ea83c50a6a35fd
zb3beacbb42c842a6198eb52f17d0e3a891fd75505a659cb1e4eb9b77f5efa6e91834261d26da0d
z5348416f8b974d646a8594423c8096b79b4d3e6a960638fb9ef102d9377acf0f40806fb1e92bac
zb72d29a6c92a00eafca0bc1813a939e36b442618552843efd59ca0147a3394400239e309973a0c
z83f0419abae2fcf172a603e09fcbf865a553d1173f599b399f7e846c46a8379b303f4436621c76
za2f4ed3a4de60002a3408f63b9551b940d05cd60b23587adda68b0e3b35b907c53550cfdb22163
z0c94ff138471e7f8ace59792ca07ce7da41365fb9b83987c72d78e779cf4afc705af274a3b9b88
z593727678a3d4b5e4be3c07e415e9e6b1062847a51a148fd4698d268cae310f2578bfb2c462920
z7c2a896fab58629e00bc93997936de3d24300d3f443f2d1316da1f974bc49cefdded6ee2a3b311
zf49719cbe9ca5ae1e1c6165c691c9bc508fabfd8f9f426a7aa2cff8aa212b10a314ab0498109ed
zd99ac06a8b2f1827289c5401a9d2253a2ef78fb3dbd5508fdba5d48fe00547eb06cdf91a3a426f
z1cd3fbb64949aec874e4e3b0c1e6faf29025fe51868f553fb271bb1402495785bc21d5bc4bd12f
z423912bfe587eb7670e65e1146e82f3c9e6d3e981bdb125d64f1ec8f1d75a29baef0a07a5523b5
z0c38810317c88a53a4e09042d2767f48714cb80f9be9ad4124b2ef9dde9a15f10c01b7485d3fa7
z08961a6ae4ebafabc6dc557e4f22e9fbf380add6849ca14dda8f7fbfe0b63eaeaa46a681916139
z7da176bca69d162e951a2f3bd79a144ee6e742de7fb65c7689cd1d6b01b1803bbd44dc118bfda7
z2482483272735d38e7e5a92232e9da78f07a8cdcf761ca063384296a24e6d02f6e7fe604451b48
zaff6cb358be74ab3c875bdf5a4c9aaacb3c0d37b99549bb98a4d28600b53a902e6b118892de8a8
zeccdd5657aee935851cf73884f791974c2b9382d969e83a87c8c14201270457fa9fd412f730e2e
z7b48de5a0e5623f21eb3300010e9674dd3de7b736b896358ca5fc6921bd5a3ec9d3a7061ea2481
zd8e2084bc9b2b4fd76b97aab9d6229862b8806aee14ba78868e1b5d0bea5848302d3536ed8bb9a
zf05e0edcb717510d293bc6f81ab1d18a205e6a1fbfa57c8360894f1873dc80f779765e384da6cc
zd7f495f6d8c9761ea66c17d7110c15aa1b3cbfa8d78f59c0a286b0978d24d95460bfabc4c6dd14
zf6b8316c54116d0a78c5e1d1c24844ac99aa4db2e196f55f7fbf1963d6ab1c4d035a5fc4fb79cf
z55ca7a3eff105a0e8d9de512f5a5c64d20b2b80f9da8e85e9e206d8c9cec4d3c39f5eee9e743d6
z3c61475a8eecc1bd53021b24894796f3aa2e10149b6fa962a1e2388c35f7b66dc3a1286d265c7d
zeaa862c22fff24c166b1c4bda0cb7defe7d493d953d21c68dd4687443c054df5d92cdf5a8e531f
z8f1c16e61229a029aef51492ea974bbf8557d133860f66cd438337ff395b90591b03f650eeff42
z593dce194cf281c006f77ef1ee9aae6ef26f25de17e038f1b942800f8da77580b5ddb3bf4d97dd
z0a4c9d4067fe2c3c6f95f2285361587b52c514bdca1b8c4723825d1878a6dce1e2619666226d6d
z3caefeee514a2265d003cef6720aa0355c19e5ad5e0983712c3d0bb169dba2b9fb70d99e91800b
z6d97064a109606bcca7f3e1814b679be603daabe8f2dacd996b815e4c72f6d3de7c01876e313a4
za04c327d8197c52b3d8a64832ef3f6cdf2eab8e963cb62ce61d785b5971b5a264b304907603bdc
z68fb316111e46e1f78d3e6a7d7c76bd5394cd6ac32763915a65adb8803969011e83b51b2b6059f
z2adda8969d35df8b2be16e5d172a3faed316fccbdf3505ad599582f413ae60820a666386fa1e2a
z32ae5c99656e146ef027d1ede3d48a3a02f98d8feffc6a3793ba26239f50db185ed55e6319ac6b
zdabbd68f8d4a9dc69849ecfd90d663c3f816604f20d29aaa93976665f705cec794b95bde3f04ac
z1a2297f49c9ed3e2d5d22249451171951567302f474bf902155949921232161884e879b0cf94ff
z4e3a7d1dcd7d9a5ede26f4ffa74c209e7a9df91f68d6c92be6f1b2e8b28bb22e242c13b7aa44cb
z3961e25d66c74aec73f3c7d0b34392677cbefccbc896332b691bccc66525cd711fbd327b3b2d7a
z716716b89f60a0e39da6fb61cacf7ecfd3c829464f66eccd7b04dda356163c2ea96f8741254b11
z1bf4638bd988c21cf5d8753c85bc2f91a052b7eeb29b47dbff07aefebe2acec60cac596161e8cd
zbc61f20b3185128b088584356618630888583a2a090c974b9590b3c756c1bfc1b8ad71a07a4243
z31f71a8025b88971080b93c4e9f69c9a1bbb6c2f647cc89ded2a84a7fc15a715d8ec5ae1587e75
z9806d5cb0decaae6003eab5b9d90fe7c3efeab5218728e5812658d79494c4214cd38c94ca4043f
z6fae4ba9fd84b811ff794bad94e5228256d176703589ebc84fc085c3ba84e0aa43a0a92dffef7c
zd95c10ede55fb4b43bcb7bea4a9365a994f1554d9d3dc444fcdcaf5136ee3bfe5ba8d83c76dd0b
zebd9e251941c85ba75b2848d07a98a56ed4ea853b138fcc477feaa9b6cc17e671fd5da1ca1a61a
zc9de14af41bfe2367e880a03aa2f887f93cdf39b0a91142b5f4687c6d3c873e28f5256138d36a5
z261b07cfee95d4baa1f786ae050d7819cc8d5d84d00a7291e69cc102a2337824bf35c54fc0af24
z116ae15089aadbd4cd2f5953a4873638406a56240d2e255499bf7b163cc30091a11f020e903b08
z3efda1375b726b57b33fddd60912c7f5145abe5ccc1996e56aae392c4c046ecf0c5ed255c557c2
zf7b36a59e5cf35f463ad9ceae38d22e79c0ae951bd943ab631254b9eeb858b3afdf6bb9d68cf2d
zcf50412948cc1c70c71461281ed410ba9ea0b3ae6bad77fef5cff7b5ab61a432bc37615341f0a9
zc77c6ec20f5beab0d0a5cfd77510d71a2f8296ebae39cb2c3771ea5d467bc6d1d9e88dd6c0f024
z437d32a8908efd7d69a5d203142af4cc7c76652ae60b29b55dc9351cc6f67b5009d6fe47340cd8
z9a1d6d1261590a90f4d347cd71c9ff924ae4f74fd28c40daaea0c90ced65667e4989eeeb0115c9
z5755af3426f4f8c235c6041df971a13bf8335c208e5708d1aaccf136c8ed64ac2fdf12b1a9a892
z2976f97e1722d800bff610a66d0ba9d3455ebcfefddbbb3418bd7f97862f211ce422093e620921
za87c4200c9d9f8a374d740d0d029a9af8a7da7138b5bbe49cb0ad1efd35ac738f24d1de32ab45d
zed1c71ae8c1b1e9384d3a6ebad158a53b22aced9aacbd4664b89a59b1ab6cf1da604d29851413f
zcb214922db55fcedb3337bef01fbae7a40550f36564c7d2bafbe5e3660754765af475bde5f1459
z3b36ed6e3b63bfec3b94080da712d6ea1d89bc91395c3769ab285e65a72666dfc6b26fec0288dc
zeeaadf84f914a779524a339792ee4941fe8721bf440868fe706fcae59b7dd3b3b287afe506115a
z45c52289497db0a2f26c62ba0273f0b1b82cc034aacbfc6c23337f324fd63b515d8d0ba1d21006
z47239d2f2b22ec2b8cea8a1094b268188572de5318358183c974521e5322bbfd431bd59fac98be
ze7266b90e38c2947aa178228a1d9f0459de1fee4592dbc0bfd033850dd3def9cf2d69a00698d90
za0be0650f77daed9ddcdb0c375f00f042ca371158d63e535b87ed66366695dc44ff13aafa91427
z0c340736ca136184adb1a8f93c16f59793102c3b9f783a829e0de449caa64a5a0c5ba1430534a1
z867cdfc80369bd2980776afcfff36cdfaf07a8f90a7dca888aa328ce521f65978782fcfab581e8
z10af2d5d2bfc3861b268cd0e2a5b4ef356f172500d7879e12c543a523462aa18f5f5ddc7860d99
z6d215151ba47d73ba130bf872da474aefbacc392df497dcba8f5cdfbf2798723a5e9f21f56b747
z30fb8e49d39e4d110a75ff422eeb9a46d9d5cf1724e720736a0333505b16ba18709307c4374d08
za5a912b93b616891ebc6b50d95437ce0835efd27ee3544fa37fdde6cdc929cd619a881d662e190
zd8c20d3644c350e20236802d5c428650ee9eaefc55884d0359067710e6184137d6981466dda0b2
z7a31ddc3d8299c5c14ab28ac4594e8c403be183cce6e3554330e7e2571caa13dc66981c73e1745
zcceefab2d1863182127c0bbf9778b3f6df51c1c28145798702bede5261e890f4aab7cd4e97067a
zf9022fff3566e0ab27bf561df8f441046f7b5f8d085d711de16f550a2248d52365afe22c9c21a5
z892718b2e7c933c07f2a9063026230880e06793140c81abb146a28195b1a52349456ed446a6b18
z46aa6ec31df3b7ab57331f6e3765d3097f06226d95438e9f8cb0eb655004229de82dc23a69fc47
z5669bd003052e173999687c0bd3bfff3df9e3568984088bd3205e8a03de7ef2d914c44452c7ead
zfe5b6f5b4cb36e2c13a3ff327ed0f7ce67b10d9ac2f4efd5343a7c2dc02bca3f1cd95c3d239f26
z093001e2289303776620b6bfb6530f663f0c31ddd3ee465c4ca820363b7740eb9144157aa13650
z887f2db47470b427a8181540a341c29bd15a4364e9d443ccae583f40992d0ed76b3558ab5669a0
zd042c61ab2b984b5312accd564bead9e5f1732630b19a80cf7bdc07e9761d3b1cbfa02c94f4169
z9a21528928c4f9b8b7c5608be2bdd915afe8e1005f9f5a3aead72a6a2099d9e59eac96439db96a
zed7c83784d3f383ded1bc45af35d1d5c2956188d3c7e1ab76c1503a9bbc2e1c2926a1a7d715503
zbfa13ae28bd6115bab8aa63b482727c02fa47d45f34c1f3cc6297ca861f045c99f37634b7e8129
zd6b1d086abe8f62be15521588aba3a51a51440226ed67b409ff946dbae09e9eb8920bf4a28a88e
z726ab4ed903a177cc199a72c2fc1b664a77117cff5c4b4f3abd609a28029a4ef71cf70d5fd7320
z18aa0698c7d44e54c8623b0ca3b4566c4abe2d4d4ac0db4b89bc161498495b65a65b49a33350c0
z67cd28817bce590cfd4b10db3c15a924ee815df2e33418f375c032764e3b771d8cbc3dc8fecfc9
z06080aedc1000ccd66cd676880901651d478b369a89cc7c9bfbdc526d225578008f71727599555
z8721a5b7003a4928a90c50f9297aaa07a0e7df19621240a6f4015b0f2bc323387dba535d81918b
z7a694be7ba5e3745864a56e6d206c878fa87e1fe31ba1bda141add36cfb1de6a97c5589bb9b69b
z4cf8cebb50fd502842fd190e8284124651d22f79f26b09bf23242ee629c2ac1ce1860444588da5
z9fb70734aeacfbd5432293aa8db467628282e053886f9eb75930c51d41c2a3d88476b13f00b592
zedb97c27460514de661c8c128640bf0b431e23230770a5d68f03b1d73e96d62a90fc5678b660c8
z6c25080301ab6b7098865590952678e60f0184aac187d4117d69cdb8f308051db98ed99b1afb87
ze7c74c9ad2caa0e03da84fd9ec9922838c486c3186295a86fbcfa032dcf3a2671649e3cd050d85
zf353bfa249b4b3035c5da332b6df5ad86b979ce78f46eaf94833dfad0163c8888e6adf582e4a3f
zd99fced4462ebbaaa09d71774ec76ba01911c84cac056a122fd214a39f809c7b6a4ad4cbfa8bf8
zc1cb60f3e8355b2626a748fc99bcea05ffb4b9f44fa2ebde82a95f7800f61d6c43114fb26cbce4
zf28abc8605e00876dab97aad3ce37b92af5e9fa172629b2b6c6b33cb6b7f319c3e6f020b29ead8
z5be49aec4e55f2fe4517f10b0a6ef4b48d9e3b1dedd406438c5db1766be2c8b8f3c68c6c1dc5ad
z5ba7f13ddbe599455d93d99753f9c7ee613f96bd9d185a841a554b10da828065c358418a41f826
z4eb0ae5ded0675a02fff190cae2c1fe3f5a1ac30ffb299c2d25906da521429f73007749cecfaa3
z3c3ace2a0690dcd6588733bbba664f514480f77503397a0de9e34edf700cdf2feeb7e8822ffdc2
zf39f8ca2c821bf8ff6678a17c18618402dd5658dea40389a44c997c478fcf31095195460ca7979
z0c6c5d6b21fddc08a4bcee4f31fcbc366a9188497c78cd5753ff8d7a1e6793cb35c26650b46ef2
z2ef8361d49396cc16126ad2d68a3414f145dc015bb479cf926c0c38b0a05c03a660b56ee896c72
ze24327d43f9f9111aa436643626cc5c489e91a0b49594cb9812dbbb2262fb0337e74d8918ee181
zaf2ec5ffa320dde98474f10158b512f60505de6424451b5a9eca2430cbfc97e6bf273d83d5c4b8
zce0914e6754327754c4edc9f030fbeb5797c8acb002cf484f2bc081b861494ca6735382e466523
zb53fad7b6c5e87c5417fbe3d2b3352ed088361052616ee4eaf43bbdffb2f543ee1df89caec6351
zdcee928f6b58ac1a219548feff5445313e7dfb5e43e0c91641de788fe2f75dfeb0de7b8f5f525b
z06bf60d7679f2a8a9467af23e67f2e686c4b861488b0a37c1070a7906550f84e6fc287407a5c5d
zcc5bdf39fb925d29172a392ed213c57488db3a953ff6d8e77843d474120522e48f4c9d31c03a64
z283f24c2d6b2cba5d6f0d428cf20c2e24bd53a38073df2ad41ce53a5db6bc5935feaf918ab4f59
z55b09908a831dc23c37c94994230974bac3715614ab4d87e33ed14cb1f5d702175a86d3af30140
z4b0588ac4f7f05315d4c82d8ac3972db46cdf042fdc1b58e5b10937b3f730761dd6050f8c4c510
z70809cd29c552a71e214ea79d5ba2a346e253ff78c15c351c00690aaeeefbf804ce10d964a96c2
z00313705b535c21bc6701854e5461f89234dfab9bf4685a2a3513c8ea02545703bf45ca9774750
z463eca3a41892aff44f0af9f379c670f4fd58b6524262e55fcaa5c6e61006d95e3c3d488d270db
z82e121b7af3c39907e85bf900a447be8cabfba60d9fe73223b711e1f2745e7771f4710874a408e
z4ad64afffc3b5202b7b715f10fc0eb328aa361687264a16f3770825e06ee59409d602efe05ed84
z67d01aeed67c4ea5af40ca926d51168a635e9b68f0431c31fbcea001a3dd2071966f2dd826f3d4
z7bb587a9b7f7baf3426e588a674e94a453155eae737671f28800c7815b1ab13bd63c07c5c8b846
z538d06eb4317fc1d9be2a35c52af35b8bff3ead14e64c5b934afae0622f47362072861fac573ad
zd695ba7cf7adb76551365a6c59ada1fca7825584d2f3af0efa448e93cec809a7467f4ae497c7cf
zd90a50381e3e3ca0603cc34590eca5c48fe841b418e1a7b4569496cf13a36865c8eb80ad6c84b7
z8f29b647c00dd7adb2738e6b2a70bec0314caa7a2aac7bb15cc06dae2885be73ee6e8ceb6cd4ec
zae5ae16e95a48448e9cb079340cf211f60324e9d19d13d8028e1734143e6a1e46a4dadb961d0ba
z2c40fd87390e29112c54e3fe25e62d7237f75e56f21b6c505e6a97d8f18197c358cbc14354e557
zd3239d7a56f6e82026418c109538c8bc41e1aada66ac86c7951154fb13c9a805dc39e8d52a7200
z1b302ec0f41c0a3010befff0621f9ed42a024437a0310d2817c567e6a0750f233e3f4655b1ca84
ze47fde5cf0edd26bbe160692c94a13d5452ccf5c2d6c310ba72a7ece9f8b1e3cd26337a4b1bab5
z497e45b43a855c682bb84770838ce82347e6e971ab132ddc64bcb6656bb2d65c73a170909fa4ff
z749933b3f7227f64a9cf34baf2909836de99c5a0e44b8a9ef98b3d58b2ceccad9fad7823a1c5ae
z34a188fe45287a0e23887e73c0d140b9803dc299e03b452dfbc53d5c40ebbb6f4b4f922b17e4c7
z6b1889c7d169e3dc644c12ff768009957b9a9f27fe3a79e5d61990236d49dbdfaab32a84ad436c
z0ca668e5fa8cf752a2acd8b9a58c5e10f846acba3761fd2655675d685ecc9655eee9c0f5f76d66
zc109426e6488fb375a624e2ed2da58e2d20816af91c05f9e1a388ae4df4861059c84e4d4b939f2
z8ad550318cb169f4f42077f6f209c837d5f45d0d41e418100c26f0c157191793113bd805153a10
z91a72c5dfca7e375a6321f7abcd1fdab0d1da084815ff0f8d1f95bc8bab97551f6ad4bfa60a8d8
z2c542504a9748f9921a7d07a60a8176396191e82fdc3557541efc707618ce0c34540c6641f8380
z8097e92b5961d83c94d9a478ba39917e3841396c6498210e913546d7894ffd82db87846751f60e
zc2a620e56ad4c942d7b0ab57835700bf26d0146e50a916696be77b5c2267822d285d9ec24e1db7
zcab8ac89586472422e0c09334b0bc77f938f29f8c0363d4e6ed89c9e6741cc574bfbb958e3f696
z740f30fda7f5be1a23a75d71a1086e3c57762bcac73757a34a12d2a5a059a6e2553a08d814e186
z8e7faa2ba6b5196b8c5d74cbfa388313c7d210e43cfea7afdecf540d0bc53567ea15c6e603db9a
zec58fe3b1688c9a8c39d9ce1e0f7d4a1a52a14ac309c22a7635b3fcd1429953633cd2c2b3e1633
z9137d8f2d48ff4e28c36a3978bac7ac4e4dac58cf27825fbcf57a02be038c7cebef4414fe05122
z3f81995c3eea99c7c6e3c88c287a0777ee52433b06caef7f3e178bda52eebd16c966ba46b9cd84
zf91df3392c9b50f5c8dbc9b978076dfe4feec8daf63c0f9f26ec3e7c52bae4b74c24b99b89a531
za161c6e9d1fc161bc3685b05c55c63595dba5084053679f9bed823e78fd795c506bb7385a9045b
ze2e9df48e69a49f0a204303a3ae0e80fd4e68d4349cd7613d80d801af3cf676a6f5841155e3ff2
z797b0943dd5564cf41c020e3717a9625a96b784179bb3dc30b1d356d5d6189ecbbde8e02230fb7
z80a378f816339c6e437d067848666a65212705a0875a382dfe0be7fff0a295377d276f4dbc014a
ze88b5b72d3b042334594853bf3bb292e4774673656f85ed50c7a317e621673a50210d8a3ded25a
za9e85616a5dbe5d88bdc9d36d7b2c2a24a10c0732a65c6cf42f3d52a5e1429b4324de6376c080e
z5686f01f5b8c6e68dc9b0a78203cbc23fb2e76c8690169cdab9e1bfb963e2054d30930df50f7d8
zc0bbb7bdc23941aac303e0a28914756690363c57de091142ea27d2521741bb83d68ba6474a29d6
za7fef04eb74f0869695f4992882a58b24c0fd63a84eddce6b3c1598858f353f702aec71c6a51a8
z4bde7cad24343fc43f28f6fc9f0d3b8958c478115e101972ad615a8050114f46dd73ac3c4aac5e
z8073f31c81af25ab453fbfb34aa84c26c893e27590c5acc2648e742298e50a5efbc590f86a657f
ze0eb5e5a18f597569883ffd3c3a4f2f9e284327877a45a83a093197d144efab26fc58386361188
z3860a00e378f20753f3a7b9aa54f410f85d863eb90d9b209f33bd85edead237ac2057b81395b50
za7969b08845f86c7dec1667165d13753abd99163bfb734ecece2fdc57584825533e4e0f206c128
z5b8f37fe90d69e123982f61a5b0dd8577e1fad77e32d47f1afb37db309a41bea926dc808d15a25
zab753115248ebd7f2e191ecb150880caf65d94090c4e7baabf7ab9accadc67280dfc2a27ea963d
z336cca03c34de0cdad4931807e7768058c260ae833046289b3fdcbfdcbef5952871a74e5709277
z31b8dd1cdda3dcc288d13e3693cb4c2040857dbfb27fbe16594a30b4057ee8f1289ea8ccc20922
z1d36851f7fff6e435e6dd038f93b9ad6a1c61b146ca5a61d8949a2a9a8d30f9d5df9f70bb29de9
z1e21a65579b4e7161f6f4761bed5c6a3277e19ed7e60fe336dc9180dd9206c25903f4cd1a0694a
zabf6cfe8e9ad0f348482cc9c0db508b2b5de047e857ee1dc923ddcb131c046a5c6a9f3d8788e4c
z3cddbdeb99aff43a6726103d1e31eaf33790ac482c3da32dd5c0122737fa0e4ddfe79b334940e7
za79646caefda02d2c39b25d8a388ef44d0b48f959300bac19fe1ebb0b60ff482f6b695054c4644
zc69159cd196390afc4e07a244a63ad535afbfedf64b09d34b5e06c9158fe1fe232e145caa1c400
z3164a8fe7ca3b6b94d221aa3ae6d831f422033c9e762a75fd6c39a9b6b088c6b03b6c63a868572
zaba49bcd528385ad75da2a6728b2238c3984f8c545737384d2016e9b4bd72ef03d51f79b572d48
z96728e32b5e5a78caeb9b301ce7b20bb54a0423d935fba61be63eba60037fb45f0cb2252049037
z3fe3d505be02e3468273d83fc4ac1f37d8cfdbcc8e6d014df25d2ad6f38d6ce1b3d7f568797127
z482c2df771d76eb6403e7d639871ca7be0903a9bcfb2069da6c3c042f51b2ea40f06c3096ce319
z7013d7011737e35825a68c9ab02c5e5225a02c39b0af4717fae7dc3a74fc9892ac005546f6a431
z6a0a2483c6299974fd89151074a953a96b364e1cb37e3d265c6970b33519dd753e7296853fabe6
z0896f3380a7e5fc6896904fadb27cb8d18bfac151b5eb3d9f181ff9acc9eaa8af110eb9f744dac
zb892e4bf5ee1ecae293ba8aaa3b71319e55e1012e41a5295a7a54db475e3534190699ae640f894
z188ac02fc135efd7268db463363ed802bb05e0ef6e60a271134e3ac252d8badce36f67b30bc9e2
zfd5fe1b44c026fe0579fa0a6027b6a7965f786c59eaf8acee556d47ee0c05e643fa296d4c43575
zd391cb056634a0dfa56b1459775d419a19d66eeccb35572b531fe6ed643e80b3b3f53f107e9a1e
zae3df5efdf9153f3b0d8bc6a481493cbeb08c82c3714f40764538d611c0fac30604bc6151ca1a8
zea83acd3d9e64e0ffbee02ebed0b3df9733e770fcf76395cb608c5c622cd2d01db13d72be58cb6
z0b57989be5b41c0cdb8cd62a93a7bbcd64f02cbf6319469931c7a8ac98d4cd6e7bb01f8b7c2f4a
z21d8fa6a8da15082ed8ed6e85dc7aeca7d6cf467df9d7970e4c669fda5de000d1c1c4c812c3ddf
z3aaef23c2b4606e14552412b87627d6c03ee5aa6441ece6dfdf338578e2acd7ec6b4fde3b9bfb3
z922fd98521f68e3e0ff3d0295a8b98d006f49f0916788a89dc3d44121282713b458894cf59a514
z2c99e7eb9fd41e2358adf9b960aa1c00fe186a56e5d2bb9d40f4c762c0aa76ae7d8add80bd96d1
zc604fd045f15a838babfacb2ef561dc664e0a6b67831df89f10071947771302c1283981366b5be
z07bfbaf5dfe509a09eaad287943c646ae009ca6883195addab866f6cff3c7b908fb25cb372bc38
z48d84c06727e4bcf6fcb6b14762f6d55401b40a943302eaa3088211c48736c88e9d48b3a27d643
z0415f8638bae33f0aa75ac459e4bfb671865e1685492cbce1d70470bed4bd39ab455ec80b7c4c9
z19c26b0983093832ecfe63597642c273f02366c5df77c5b02bdaa616b6779500cbc39a4cc527d6
z07f52d9ab0be53905156aadecb6583ae16be842245dceb20029ad73051392b0cf04f7eeb2a24d5
z290506c91aca59cc4ca3f870ebc976d1418e0a13aabf1345da6d0c1058502cfa2aa682ecf54d6c
z838fd18dc3b7f41b2bbca7bf77efbcbcfc74754772b30e0a8725d9a02bd431b2f9ad7112f17a3d
z162a3a706560c8f2dd9b4f4eafc19535c5c387d32e82ebbc88b82cd8c3afd18946560d734980c6
z79832c28a37daee8603451a2f32dd1be8cf4bab072e39307afaff2dde12527d43b173168f65fba
z5e8d4fb8ab8aff3a0048dfd7424a7d68c9ced67d84a48ddfc39e6822abe41b9fb6347cf909ad0c
z7b7feb4e47c69cb0d524323e2521e627c1bf25bd0cf0b17a74d049df32579ffa607c6adbb2aca7
zde5a210d0629f0ddc64d8fd854dee4de3f12483d99c28e0dc578acf4668c2b2d7408e925754d83
zcffac53aadc1fb234ce96107cbe11e210e47ada887f5a23d39b4c141ca14eb864b951443a7ec67
ze8256e2e972aee7a2a0cfcc25911c6e022b8cc0500c8caf27100ba2e110270262e199f2ce68f46
z26557ad3d65245d780cb8d0279e94ae750071cf97401ae15f735ab89ce23deba7c79c822bcb24a
zf5ec6fc13c77c2269b499fb19af367a109e56359f6c55c46756b95bc5c9a956bd706cbff887e7d
zbf534364b273a8e7f8d24d8050ae069c4c399e0dd6c3410ba4a6079185e0dec2498dd1afe88ac9
z2bbea01589e1cdf01904b1285444f7e4953b7573103ac41da0ea4b3915459e137286450bf096cb
z1823ac217b120b5fdd7e7f024b34abb2f0b142cd1d748d07d0350ca9b8c828044efed3302a41f8
zc5dcbceb48f7711ba874af5e7c1da0f7c477abb6b7965ff315a69f9684bc38462184c8a8676f7c
z0670424c3698a9fceb17dd0200384c51697f904053a9101071d35702714e0f472e9eb609d33f94
zf35ff7953daa90231ca6e4244080b12b8999234acac2cf2c01a863902413a86b6a360ea13c146f
z9ccf2dc4b947efeb4d75a1a68f4a6c43db13d36e6b55790fa88a1ee9c2256de2014358fbad97f0
zc671a0cf6618d7595f46c57131cb354a9db50a0b98fcbe57201b4a230414f3fc14de31bdad683a
zc28c8e41a6f4881c6f2de2c07b4cb9356790d69c090e1ddb48c7a21644aa991aa5f92baa8b20b1
zad61e201c989b7fb12ee585cf44c87c48b4c3a214755655a1832334b467cad39bf2e0fbb5a8935
z67a8e4c444d481aaf4236a1074760da3599ccce75541b9bf8849265a0dd1642fdac1adc6930024
z90a35e9160611981da07b613f494f9662bf8219ce9cb79cf408c27b4c332336bedc7ef637e9035
za2d75f03639c6648d98abc95de566257e6169dbf176d93a77e4a93045b65a66f060da1d2e08e61
zd4056a117da844b990b209545dd044970e1a8bdc6cbff3bfd9e7dec6b2ec7753886486429a917a
z315566b03b8c8ccd84ee511029d8908862c33603a71c93a58c884a9ff7016956998cb5fbeb6198
z87339b25335bb811afe3396d12fe53200d3c6a68f216bd87aacf27a99b3b2857a3609a576a590c
z4ab1e9199c2d15f727d7af79cf7109febda1ff16df270adc4ae963bb9b89cda1d63ca666fc97a9
z62d9733cd94c71d4aa6283166be16e1dc82d8925bf54f36028790eaa37089d6d7c43e3036c75fd
z5ffb11c3497df9f676db017e6cc4b0ac4814ac4827af20521ae036092bf7bd86347e67ea791a29
zebf5f9602fbfbc9e0478fb9707a0aed1c5a0d0df13b10003cb3661e99269226bcaca82acf0b7e1
z74b58a06c309ffdc9f964bc1adb81b61fc120a98970165b406f33e431dcedfe6e2bc245755ada4
zba343e8b3f8dcfb09515ebb47f9712fbbc70a4470de3508a6e97e079ce66255faa7f13f9ab142a
z0f998ada7a3ea353b730dd1dd62254f92237847016c159e9ed46748f6706410a28ed57984ee956
zc192c93fb901a6455705504c2cda904388bff68904d3e9e968cc30bce0c76e75e98c9d4764de10
z7466f0714dd466953bc35525a0a1ecb877d963da47ca944d80941b4ed15f05bb7d84062d212171
z73658c5060ed4681849faee8ef7c6063235e8481fca2dec79d65cdfdd3e0060b878b068e670e27
z60b519de81239f42629c35ec0a4de3928091bca882a77bfc834a0e1d2280ca3add19f5d16d5b7e
z5f681e976606ea5812566b30e8df246ece58407ff2f8cb79ab2970d0dd2dd50259a4a2ee966916
ze545dd58dcf85873ff537410193ff37ebfbfc77b899e8a0e2410d23930767bd1435858bb9f161a
z5c29e86a13c50e0524501a36f4496d5c1e72180becabc801765c3cd10478d74fea71a8ec5c9a4a
z5fe9d8d5a5be799356eb4efa09b34c0225ea74952a56999feb723db8631ef47d3d6c08e5fa31c5
zb4335d233e84571787e834b5ab2afa5ee8d5ca8bf4aeea3e02cf537a918680ce26d8c514f123a5
z8e732339837b8147d9a2d5449814c755fc1a677afacd716dca4231e68e0c6e5fe84da846290b88
z302d4ac1503eb12c6edbe4ceab4e1cca453fc54942a7dff597758b4692fb47e53ac5118ae05e15
zdf98e83f15fb6b7f9197751704c86dd4ce1a0935ae180d5b4e5d2138608f7590348ac072a65de1
z1a1d9bde801486c854f1ac59056a9fdfcab72fca089b79f1b38c1add030813c5394426c587d11c
z6f3daa34a62f7d02000b8eeb413fcf9ae871a49590084d1de4697afaec9bb89dae78d774ca0dba
z28dd225ad77a9d8567e9e031d18088ce1d0a95fa586a24fa9fdf14c72b3cc9d53cc595b681b015
zaffa5823df57d725344ecadc40be183474aeda1227f28f6571a69e46c9a66addf54d50d06d8321
z09997afa8650f4b71bb6db9a52d6785edadac241e452bd1d799f40e8652313edf7220d24bbf0c0
z279f183d2036af5b202aa2ee3069848158c9b9637ee3606cb1de5af4f4dce5404c770029b07bd6
z6cfb9cae23d47c277718bf4c7a00436bb9bf7fec3f36bbc2a6f7e8134cb15abb9863a2e0a55283
z508e8ce1643c15910c4318a5a72b2be761ce3e3f5c4665a9389b8a1be7617f01989e216c851f5b
zfa38b1d63ec3ffcbf57acb73b3b6f29d5a1e8874b0de302fff63cd16fa6c4d58323d5a60326289
z44cba94f6429fcc0534330b61064c420eb8c9542d44a21a312a3cd9849ebc1da64aa4339640c1d
zf6e09d371779987f99b94d1882b8af5720c36b6d25774766c70baa63423b560e41bedc814a417d
zbc51fb3038d5c0995051e06c43c42edf0f918cd45f8ed1ded63190e33e2ffc1b11d993ac9f26c6
z57a7daf2292f4b381eb24c4c801af7ddc0eba3a3f8448a79741b1600c7f3fa932d7256fc7ca905
z7186d418ca600bd27ddaca95d2b046a45b40640313450c9260f5f1e0ced411c7a607783edee696
z09259eb7f9313fbd09f4b6ba0d7746ad7cc8e055343d6d5381ee1bb50682dccbba77b0ca23f570
z4011baca2c3a147f09817e7d0a2647ade4530211663d3e16b93ca5ce94e8d11e32fdc8a0b0106c
zdbf9c9fa8e74860cf0823154ba7bb3dfad53877e4c0ac3f7f9697bfc67cd58f1d17b4a05f86466
z417e3204d7efd61237cbf484afdaf9c04a43fd53a7e915610e526e87f2ce62aa94cbbcf66b1e85
z8cf0adf17e47dff9606a8a44080306ac8ed36cfa20609f61c6c35b089e4960d5a434727aa0522e
z4a4177b56756db855bbb13d010061992a9f651f3031ba92fe95707fc5f9ee0d140f3e59a2e9f3f
z48f614ab002c6fd62e8a89ce936ef0455229415f59cd31b27d75a266f71488dd7f5260ded9ae85
zdd82494beab309909755f7eb04cb0a1d2eac73d15ee1954080ae7fc178aa1cd2ae1d67a9b0d7c9
zddf7a637f418a2d9c297a14fdecea85217322e7b76ebf61bc2d644d6d4524d4f4a76f4c1fd1701
zd5ac69926afaa63ca73e64614220550dfef4d03f2ac9d591afdd947079d0b0a9e912479453f12f
ze38a715784bc4d400f5de272d94c212407c7b6d848d6f50ef735330aab4f64ef47980971884b90
zf6db9d9b1dcf5d7ba7b7c34aa07735fdb118eabc1891c7780375b1dfb545dd9d1220fa4b63f642
z263bc1030bcbc07a25a6cb9f8548ecb368a761859025fe984eae78c6822cc20c74e9c7e35e425b
z38bee0681e9a3b363343f5775ddaced3aa1727179de2b0c8ed4101ce1ff1efdd8a4d275dc1ce4c
z79e0bdd74553f1ffc3fe85cba2a13accca7fdb7357bb17125ef5c9f996bc4c0ea64b985a772d05
z5ab00c9165ab4693a3845827e7f64c39c6792156aaf88fefb8af8bf50109a83133d3b4bfc768a5
z854920caab83cae34ae7310e9b8fcada1cfd37aa844cdc3731a93a612790f5f09a8f6901316fa8
z35a331380dc751fcb2a3478b80bc9d4e721c656a9d40f083c67e65fb2f07d8a39d1242202ed308
z9ba3be9685639aa599a19f44bae0162e1238c6ec7e2710a825fa9dd8f66fc34c3441de78fa6c45
z7f61c8b99db1e3256d7374ade451f21f0a9a0d3d6ce4c18468105acff4cbc34293a57949a66204
ze000a632f4a589ab15efd8edfbc4f1d36faa985a37d56335de40e1080551e6fcc8e84f910b40ec
zc9982ab69b5c3adc91124724e32d6c7c51845a99f0e89ae52f9dd80a5d03188209e9bd0ed8b754
zbc3092acfbec3d5124d7f0c29a356f3da46312c5b4b6a9af2e447f4151152ee9df96d0eefd6c39
z9801f113fd70f4f5e472e691618a91f42b09d697421cbafad6eafd875acd00060e9e6d4d2e9a78
z8209b360be35e2b25d11a41c5cbbe8bc17f9368210f427de32559325dfc0a3857603620eb47ae4
z5b157929dfbc4be2a92822c60b7ab05bf16cd126982b21f94c26d18cf77d0dcb599438a923a743
zf9c2703929040694dc13a69307ba57292acef800c4875f5b8af718c148f6617cb83cd88f2fe999
z5b332dc66949fa2c60a577764f81176898fe47108dc72b028e0b514fd809933df1edb911f63b13
z812927efb05e327f2e14ead50619f24f2cdc510855435f64dd74480882d18b9f1a2f053b34a21c
zf0a30b1f664d4c12e861a4d4282d952fa6cf76b5eff0a74f388afb5a291e28c949534199e676dc
z485230202179e953fabfb87735b4b228bbcc15038047830ba7770ce979291d59cdd4914858785d
z636013896c269c7b010a1fb34b1ac49a95f274054209b6a76e67cfd2253b17f1275beb490d5b99
za5f22f75fc30eb15cc321fa2cd436cd868e5b66f834e7c162f756b04f8a7225e57291ac3a14c2a
z9c0a01c53bf4df8d0d03e8a2eef64c1adcec698301664f8e8cf262639d8e1b3963c015477a9e90
z3cbe9633da972c97be6b123f037181aa73d4d25b507eb6880c90b202fcf4e139c8714b1d540500
z6dfabafd6a3d4ce51e5d0a2538e6318494140b0886cd5d42760361d24b86d636831694ea774d7f
z208a6a6bdbc92788c872f6441fcaa396964a0c086647896a2b97e8bcd573ba396208bb9909d864
z0ead85c4db3c19f6e0e8b2506eabef854d23d11e0f523432312514b19ed378e16595ab6ed74658
z55f0f498b0a7ec2be102b1c19247dd594433d24d974de78fe717bc9c1aeef663db85f84e3ddf95
z6e65c0005dffae30e0ae31330afae5d9868c3c671f8d29cade55f852a16dc4baa4ca5eb5d5d7d8
za3f1d34bdbd805467a46502b430e9e4544cfe5e1cafb00b3c27c15efa4e34da8b4823b30663234
zd736f31e6ae5c378941fad366b661c526831c5f5cd1633ff3922b4680724c16cea4116f12714e9
z376fe910ec9883e373169642c970bc70fd0a060e937e0d59ae230ac747b171bb9e223c04a8b67d
z26341a9d8ceb53a42ed7bff8d4682e6e87b4b128b1f7c8f375ba7381db5f3504f8180fcd1c8b2d
zef2310e3bc8d7d1a510ed55309782344e097e880c9112d554bcb74f93d07ac71c5428af301fbc5
z6f7d9b9130dcb385bec0f61736c4d004243a11d974b0b47bea6fc9a6c45d47c27c8c5b0c935766
zf16db6c071cb6198773207086d625a96a5b993e5eb9712a9b03130892a0b3fd75d5847a45018d8
z0369f59bfd87a8f00edbb209a7ce2c9666da465e3b26e4130228a651e485b0e19cd5c5a540fa30
z6b72d509cc5e43f904173e1d432cffd37b685c6aca2ace5e0f6f50ad8db4dee2211eee2f2d852c
z19faf7401b1455797547e5542ce3618cebcb7be3c169840bc4e018ef93d74884fa3f6f1dee4eca
zd86cca02bca40664ecb0e577d0320f00c9d73cdfaec521b2302c7b34bf3c8097fb970417157403
zc81b0a1b22877ad58c396dca8257b12f4dafdda9c04c930438cac37219c462a7ef326f0efd37f3
zc7e91c157decc38f7de1f1f0d3efa1e00a775f84c357a825412f1107ef2d4b81fd97dd219fb5d1
z84cc8545be9df2c2223ed81be2b9f014b36a4ead216673fa3a77c760ee236fe32fe0b39147de71
z579a0432a24785318b71740b736a468c4d8fb20fa4bce7cc952bbc1c84ec1721202e56cb295e36
z3e96bbdacf020393e0aa632c46dd2f558fc803f7e8fcaa128dbe0b8ca3b92617eb28d3b63be4f7
z42e84ed1a98a95d10f4f582dc75f7c7f06b59dafc0a495cfdbf481c142d77f26eec9d0694d7303
zc64796511c8fedd0f48e4940b1b0e515f88d2b59cccc70f2c746203ea0db834455557151e82951
z8b8de2ff4bdf398b2c8def83c4b79457a9452c4bb596732874704a066d4e3d63402d36c1594f66
z0bd68e1d3a6afd6289111c46042de3f7fa05c954b92c89ad8788368c99b5b02a6184c397d08107
z87cac3008a57e8f0850853070cd2b8c1fd52b131fd2b640e96c071526a798984303e1e5ad1a152
zd96cd733a9451e432a32769c8a8d9870c548e52dd60e85d7a18df63b0a3c5c243dd4b8096f46d9
z3e05ccc66eaf616f6ea049be47625a83fe6f288a32e518135523bac5201fcdd8d600125155b456
z18cdb3dfbee02c0e2b921fe6ef648bd50baa1e5247dd185f0ff4538dfec6f3356248001aab7f9f
z44076c1115e66a1156f8d71edcc2190451c1c13daaab2e144b30d93d818911833f0df5787b93f3
z0aa2ca1b7f6d72d9f0ee4c3e489575149a386f6992b2cf878d43305738ed19a2ad8862a2c2c1fc
ze5cde9d7518d2287d5f4b609441e13a381ae24846ab9effbf0cc70ec11fb08ea4d58659c71152c
z525ff42d1943f81f06823e9799061cb18c78a389400ef548e8830f4cd5c1648587403ddcae68f5
z750898c3c080553bdd763060c12505835f27163fb18c5b174b5158917993d6c6f5111858169574
z6b4a5d431fa9a8aaed41c34d3b89b950ab883a3b6f39397bea837c36fcb9ed773e786eb194c761
za16ba2a111387b35d5db166ed0d643b4355d70a9196985f7d16088876edf98a1752f4e5c49fff8
ze2e4303bb5739c542188f0a4223293919dfd383b5e015895e85feb62e4f6cff211deb0b646638d
zb910e74a7a43493f5d3dbe6ed24a03ceae6434730c764f7524cd65547c573744bcacf8d406a6ed
z8442776105fcd0ec5585bc6dff5b46d11aca0e5c657768d1156511de4bf2397f1df2255a067ca5
z6c855f236ccc43c736d5de70ae68122f7d88e49e74104dc00ba96901d79a78c513f58470975236
zabb4bd36a876241556e94d1ae8dcd19308034790160a04c6b99ef810eced62eba9f50418abbc69
zc1081001367c3d0e4a73f7f973a6e8ae8e0a17b9940790541438b308ecba254212292eb7bd29f6
z364885e591d464a8f5ee9fd239c51558a7439e175ed8d56e3ceda094f62a9a01548fa2e0389b88
z2ed7ba539bf1d44f8b24859c17b52bc00a5ebc63b766caca2af5aa3bcafd3853aeea971134d161
z2418fec7ad25b7dcd0a55c3602626d67089ae231a15f42494c3482ddb8cdd2bbdf8521de64bbc2
za3cd120737f31c6ee0347d89529aadb44960bcd6e503c60a9bb75e4ce188c628f0f48b3409b616
z3abca11c940ae1c7461b64189279facd14faa30cb2bf187329a04a9326489cc50aefd6e66f6720
z17b8ad471817a6217ebf9d8b2655537e1ba96b6b371a93b52560917cb2daf5eb28c4342e952055
z02e8fdfc2ea2385317a6794713814fbbf73f02ad9cad4380c622171faa68950e3108d41d066c7a
zbed8635609ba6efdfa9e9e0e586000b974f9851ab898fe11550de8d4005c25dce7b76bf806defe
za0516a822aa945d02472a16829f480ccd5f20900610f5d43e6fd11a7a0eb6ba9f24a38ec3a9e00
z90a2e633fa53267d9003a50135794427b179682dda1a50f76f4a5922b77cb8b26dbda378dc7904
z2aa55c0956f50b139de22a1c2de2e6987684d01a5b22d7ce8a015b88eabb5183547524c23bf2af
zbd8013aa39543abcef670f87ae3b709d06b17072bba395d887078e890ce88c4c71c9cc3523a934
z05cdd7cb286e9c3cba81761234c5472091c2b779868c00d29e08be7270545100ad96069ea92f13
zad608254b7c452472e93f4fab914b73643978c75a72d905b06d056f6c3ba2cffc3d36cc9086008
zfe573a034379b36ea5a862c7b3b021ebbcb98faab70b854354eb001ff76a0d5b4e88dd1aeadac6
z5a664bd2fff65436c7bd1447a960512457e145a6a0b92adbbe7bf64f59c33a38ce21887bd7445c
z68abb1dc7e3bbb87eb441b675b7cba2c06c1440abee3c97f3b213d85d42774a1a8da3c47c4fe1e
zf494e4a02ef1183907b777441a5975000cea108b93c892e20c72157c539eaa379a5c3cb0d072b0
zbc5fb79087f5e3a18b8929b8bd517e7b1e6554f0f74ad094ea3e37a7ba156b87072b113ca34778
z33cccbf61d912687edfe9728d316e01e8cdb42243af87e5290f8be457c2a00e80d623db509010f
zb17438d3ade849c9154261fc1f0596dc1c10471fd1ac0044adb8edf52dc45a3d4b972dc5fe6718
zd774c6ddc8135768aa062c796f9d69615cc8a69ea49e79e9ce34407da2d1c6836eb8eb376d74b3
z1e722acb0b2d31ca8de1d376ef96d8978815a4560f692a58c085d1d79e1a75ed2e2a5107bd0083
z2b1737db9fc2e4c16cf41eb300acea20bbb54d52addd2c1536a5c1220e50769f31dee43a2e99ea
z1a2095b25040eac44d58d19a465098bba4852e0b5c2ab4effff9217ee5192e4c70ab94ae142d52
z32f8e8ff4ed37e96ace1f6c1294ac0b901ff51107800ebb252ce95d06e4a9fbd7dd50f8e7baafc
z1b5b3b58265bc45764945142f5f014f06159483b5138d9eb9d9ae777fef9d63711d28f05381b0a
zc80eea3b0fe8540b7fa75cf3d7a942b8cb3608d61647e59948b30f2fc86a87e483c759b5168001
z0342b1c04fea6be075443ed8660acbe99b5d2748b174696bff501664b724d70c05dd5814e48646
zfc77526983c0eb435cf40f556cd81b46d42df797582ca56a9d04c732435ba5d2edd3cdf669d952
z342dbaeb347aa13f0770094e589e0b71b11140faeeed07835576ffecd01815acce97b9c2800c32
z3f8f4b4b6fc57fdd794a32408e63704d204681a1efea2e00d4d59dc7d40c156d3669bb26169b7e
z4063204e79673da1aca9af64a045539fc5bf60e0d01e777ca44b1b1ca937c3e3259cd65c9ca73e
zba6932fe59849079afb8d88ac466a46a512ab38cd9f44c6ea2a512b6857af6d4f351bcde1a2a93
z4a16275552387550d0285869181ba3608e222051bc4df9eb0f43d5e42c4e0a0d6681da35fc8ee3
z3ebc09228a6f79b6f8862771317e7dfb7ded9869050f0aa723d568bd2c75139a230e33e28cfb99
z915d30ee28308fbf2dcc7db81f430001b6a0d4191f96928583731aa75653dad2c4b20d0110077f
zeb448d9de0f895791fe1c91bfcdf7d3d417608f0be8d15367e2f1a8c4e028d4432c2c3ae4f9597
zc6086758c00e316899ed6ca9e57774258fc0499f0649fb068a07e3f8692d127324eb18b4d5feb2
z58366414042260efe3ac2b22692e52e791f8c668d8bee350aa776246982b560b9d494d93a5efe3
z7c8bfbb973f8105035544a1908daae70321c291befa9b6e66c18849237721a18850fcdb945da58
z372e9b5f3b51c4e2bc8bfcac78131b0793f6f5afd5a62051677294aada0e004ce82ebecfa354e3
z4cfda19738783a88e2bf2d97944f31cfb5b37f4bb7ea25902452f9ac1f396fe0c6b96d54966b67
z809255e6d19e3930728eed6076c64ae9bb6e5c7d64b4e0e3aa912aba7af5a599c8598244346aac
z4c25e24b7b317f2485dac6250dfb98ffebe10b9c2cb76916bf845f0787a963510c1a2c9c8fc1d0
zfa8ac57997314fe63777d917ed10ef7dff1d496b2591afb4be85204d954e22cca8cdefc02ba88f
z8a8e2817138fd96b01391d4845418be6f4eed8d53cb9b0ee7b0ca8662fb1dcf91fbd99af157573
zda780914e9c679bdbfe77ecdf0322a2a71819e3b9993d912462cae6de4e3cf3efd02fc66511299
z34af1f4397f53e1701d57dca6fb50431268fbc1de5fc5abb6506929211a6be3e05b62b14355c89
z68281e8a44ca870f6054e04808838f61ba4881e06459ccc303036e4129b8194fa686d0c367856d
z89056bd00a3d2c601ea5d1799172c91e0da91ff1300c34ed99db022ca59af6cc622b2745d6cf4b
z7d8fb59ce18918f7ec82476ccaa45650ddbcc7c76142f8794f021e054f7021b95bfe764f7c68d9
z6f188e0a64d3f16c327f724830e12ba40c255e451c1dd5333570f10963289571ee65335f18e7e0
z5339b07e470e670d161a5fc4ca08bbe84d1f8250e51a9a26570922b4ab63f68bf335f690fff378
z0b4b833cc26415f96974cd628c822cef80fd57c7ae5abcde4f461a0328149fcee106f274201255
z4619ab9bd7befb584ce96647670e1c198b2cfd047f48e093173ae1263f1c27895b9d0f6646e070
zbce8eb328a7efe96419cdd8173e90221c8b76e5f5d7f6a356b1af5b5e3500bd48f682f567f626b
z0c8ebb441cd56c5230c5d72b40b3fbc8c4e230911e1df56e083b357123cd10839686c5f0aeb4a6
z67fb3da53d4d823851851bc44c9826ad8313435a9e738c62e2617aff2ba7b9963b404e0b2ca6dc
z6a3bb5ecbf3ee44dfe0a55c09b8eedcd089bbefe03727faba861aac67f5e6a62287859ca4ad2c7
zb3bad5a9610c7856bf9f888cd2231a6c416e87e1e29e063d961fa6fc3847c92d5d099ad2fb2a64
z5d408f9f5f971805a387a9311b3cfeb6e5bead888242729da9a66d009337d0bae0f6559d50d69f
z33158b43f03aa81ecb03fdcbe675798811af32a0d77abfedef90cb3af3c89bcb4fe033e917c695
zc4fbee44c4e4c1405880a4017789bc68c9dc6dde07f5a9ac5da4d959313dbba3b5915299df514c
zcead76e4c932b6e7bdb0fbdc40cb0aa1761a5f8cd68923bebe3125f675654cf0f3d88286f368d7
zd38e890bce2dd38ce1cd7d7ac609d24d2c73e813129ecb2d660a337e3a70f36ad7c55ef78c95e5
za045e87548e655067603fa994d554994f22d4e719d3644b4d5b6498e3a32371e2ddbcce4cee674
z2cb92ac5b5ad8c05a2cbd5496c0605f1d97cbac4454e26392d1bbd2eb9d4bf37360e3f205ba5da
zb9b11fd5baf21fea1ae899004f5476f74a75e89b9f1c77cb8b3a1cb7f142b6490b9294a68a06f1
z126cc39ae4bfc1983477fc259d6bf292f658c92be6fbd679c86009f4eb633255ea744b3116656b
zb7560d66eb6ea43bcf6f8681ec753e4ec8d3e8f5edf879b7f890ed19c8fd6ce36f714b7a109ec7
z7d7ee6f83584c935fb32a0936d1b9c55f4cfff2ce1914c0cc48c917499b7b336c56d15b56bf83c
z09459297fdbccae1f998093a31be1ab4ef027703a5f926fdd58512089553f408d5cd8fe62466ea
zead6c79399f0dffbca739c11ec6058b5ef9b26b09a5f3ce8ed8aa9d4641f4ca153ab0814837bcf
ze5f7339b15148f439f19b8c529e62c3aa39e7618a7267cb4a7c59fd1502d9af2323b62a5b12e90
z9b01bb34d28e3b599a1b7921ebc69db8ccf541f9977db2f25c3892e883f81cbfd876c89fd676cb
z8075a29c7718279e3b846d8317f62b9b924cd4eeeb7dae541aab6132229aec87d24dc09cea0bfe
z2267e4f78422cdae08ca41eb73c4dc6c9a8f2ca340a48b0ef0a14e6357c3f9b3c93f700398bc8c
z1b6d67baa49c617b17273b1dbecdd34e424a6a929653794b0c94e1b0d9fa9cfce331d8dd49d65f
za4d22afab3c0e90eaa4db9113cd7ba670bbc6b78292ff72235f3e4b1ba43bfe20abc72eddaab4c
z58fcab3530f104c93085b44a718a5c0255d3fd7f1ea3ba558f1f0cb3aec678cb187523e7e54fa9
z65838232bef3888d76599693a343b9c5ac8fd7edba92ec4dc870b4e920cb8752d521267028c2b9
zd33b848b40b9227d07851f1f9713fe6845efb9439491cf14d5c1c3ed767648bfc7f103adcbeecd
z3f509fb41b3fbcff342f90efb8cdfe0a78881a2a74f5ae5296e8d40a8c4922cfa5a46479fe739a
zbe25ab0103720ce524b79eda380b469ca2468826c68a9036f0f0a2e748c5e2ee0af93f2c8943b7
zb550bb61d862450963ab6e096915282aa1f13c61f55468837f6abf242b40c20b771f82f19d7c4d
z0cc4ded53adbada8b0a02fa8f3d8a9462ee22435ea562ce5a9989323a1389b8240a5f15eb226f9
z0bd4613902021ab4e35728fb1aa518f8db6f026c0cbbeb84d3bd85b6bdb04220f6968cb28c2432
z9a406e89df53372d666bb576c2e75b4100610336f9782267694aa683abb43eb57a870dbba5d585
z91ce24ff44bb233ccda4117dcd012baecad93aa51a0e64258e2174c6df1e8bf80fc7a7ab89312b
z5dcb08ed49fab0ecd2d7873e3e009e653b6a687eed5c33d392fb265d0a30d377d292c29191d95d
zbd2c740cfb882855294550c08bfee5f6b3cfe1a0a0a3d9bd7eaf660b47eb1087721577580180de
z3b5e46db7ac530249610b410e877f3f9bf3973d6e44fa60486a8cc0323214566ff16bf7621ecec
z67b21fb2c0ce835d0dcd1db3bf8ef44c740d52f773d46284149ea1261fc2986abd2e048e51bc66
z82f7ff9d564087e38838dfd426727cd63752614c7ebe1d77842142a13464080fb199aa08da665d
z389993441d82366d300f6a4dfc61cd11645880a37fdd7b25a9d1e1fd23e1f0e0ac8c7b3b0b6a9c
zde73abf02e2c6a4a6fe19670e8a6e78eedaba7dee821d4f00b0521f82ff0125ab444c52791d1fc
z60d784bac931f7a6beb085ad6eba02b512aa7388b1a3459f066b43d4cacf180cfb5c54228fcfe3
zdfe55492a1975c6e79929a069906226111bd94c112e9f16e08069196b2fb1f776875c3fca4f632
z501b6c8f861187559fbcd2b5f089ce02ef8e068ab1518932bb2a2f5841248c3a1b05c8ae524963
ze04f27c667b5bd119af11ff984d0b958f630c3cab7659592ea646aeacb3e28c92f0f64a7c51a66
z14b0276039f21aa3d0c8fc3586582d5cc2fde75000e2497b13fc27bb212550bf448ec10ad7e5ab
z87c0cdc14e51c1b96cadd9d957f99c9ce531f10c1ce94ce5fb638e0599fe6e7ebe2f4b7d0cc9e5
z8fd52012cd69c09b75ee3aa003341b0cbed26fd7b5e5f0625eeb3337d4350d5bcc385029a1c6a1
z5de082302b55b846fbb82f7d08299fb79f54db09c60fe92481b94321b89e645d2bc00cb1e2a84d
z03487c0bd20fa95aed2ccb64420227ff000a6b918d08ea99ec7ead0be8ea4674bd1af5c6c833a9
zeac7195158bf4613776789f436598bbc3c914dbb6a7ada1ee3849af1cd105d6ff6de334227801a
z3587f63e7621e70ce28814bd1e01554575569781d80c4e4f9503798dd9e0e6ed1b93bb773c6eab
zc5c11bd046eebed6fbb58fa99df2a1ce1081af11f64142a39ec8e9dfae5bc1fe2bdcac219a84e7
z4c98db7551ed07d3f86b434949224c5fb6559326390900639c8ce83d286d561b6dcc4382fd309b
z3d7e1daa58b309dae2642812ff23fd62fb73188c6c6d088adac515cee19c594512e8539c9978aa
z9d7d2e382b03491eaa1a4a4a4e2cc877120daf65da1e81f3254173af8d91bfcc60dc667d3683f7
z40c7b5e6dabee7d7c7d6d3e0e6fc06f0712f4f02c63519505c1e697eb83d77e901de48abf23ba9
zc83d3f2e70fc75c21f809b67cf1a082899b0c7062f120334f82f6a7ed74583e8d57ed2ee4fddf9
z323de1a2601d1e091682910ea2b896590539193bbc09dc4a7c59e3c1bdf5d99e15552d2664d91e
z459d5cf6572a6796515b8e2054ccdb4fff197cf2e9bcc7bac45544a895c653a3f4f11afcc566b4
z8e0282ceadb1a5e071df0f87259d99960beb8604e4bbc9f30b88f5592ab6696479f7caef952918
z303da4b9bd356ae9144913a99585a49b77a18338ecea9c91cc286850170aaa1f0ff09b38bb4fba
zc6948aaca0d90a6020060ed86b0253c09529ab3b246747852670fbc027e2041043969fab113948
z8c0c063c90076b8310e26835d0fa95638c4fdf0b181b5ce714ed589a520f3a65a7125cf022bf83
z2ea7c55d412c045681d99f225e29e3fa3419c7e30317431aa07e41be5eafc0231b89ea9c9e9078
zdea90d8eb8b2e2d6729098319d99b7b6114edc66b8eae206329057faa8aedbe18f3d4e9b601cdf
z6c41eabe260d4e65048c5b0e0c68053bce475c4d37fb103a9a3003d615ffe62f6edfc4f86459af
z1d82ec28ba43c5f978caae407a022b216cc94a697adc98980e3656482c883d0f98e82b40619ef3
z1dc8b3978d443fc83e8c1c500d721c81effedd94f39f69b87c040dd6827d069d0f207b9d79e12a
z5ef8609536c6d09437345e5d781baf4d42a3240de3a001220c12719dfcd452f7e1632325b773e9
zb353e91a9f67e2b174c49909d9f96acfc0f5121b636f7b75c851906ca51ac6021ceccb0437dcc8
z26ea31583e7e6707dc957a62a8707853f4d91755f9e33370cdafe5eb59ccd36162be9e74ad8648
za146e47ce7c07bd42d3e41e8aaa53d04830d8bb2ca5b05a7ea9c6d0d1d335fe7437776b5462043
z556038c50626f1fd89ca0c3248244059c27fb09bdb3cbefa0e0281d84019dc02a7a7d20ad2b840
z295e3a47fc42dc0e736bd82a0d58d89237549b209b95c81a52fe383830bb76bd75a21223b6b715
z585f2d109d52880525dc5eed90a2d4ee57995840f602672e5ef5dc71b3ab17250725c52def86b5
z2fdbb3c50bf2ff5639f149839d3ae15cd804eaa8352e888abaaa11b6f3585bf408af80d1e59d13
z3bbc3903390cb22a251254f06ef9ae197c28247aad4b6c4c68cb169a50d700ea073889c24016e8
zb5944cc18e3e7aa3b852fd4aa34e192c810fcdfcf0c04ca0cd898fede3ec448d939397ae902618
z1c23a4af140aa001cdc992e8c7f4502c274f84ec1ca5b5b851182ba24414d69499ab196fff658d
z7c9d3b2ed65d08d3c83252e6de1519226ca42baf2bc3235ab9f4ed6fc468ddfc8bf52a5f25aaa8
z19c4d24c4baddfccc545c55a867ed5498f3a8c6f6d051359599d240cce68f2adb06547fa1163de
zd2af3cd969866b1ece6732fefb82bf9db1ecbd330e14784648d18ed789a8deb1801a96b58ff789
z4b64ded0005a0086625acfa8bc7baac119da68789ea58f5bcb2f596d259b54a0345556e31c0a2d
z2f4f7f584ba762c751e5abbcb2fc22e1cfbdda3ff709bd814ebb82e2bd70f27d5147c4e9d8e62d
z4c85e8d77a651ff5bb44c0c1ca1999520400b74403fa43817f8f916c0467b559a3c3645cf6dcf0
z74aa02b36746d5746c6e6bf358eb6fcc2a8ea6f5487ab1156656298326b4ef25fb6a31a74dcb48
z13951cac86698fadc79ac9e9d8312537fc61330084192f6167135d8d2c52a3b0155cb4b3f7ea53
z34b8f524c801bdeee6c8b2f67743cb11dc6d1fe0e69c18cc647706eca9bbffd12461553c9ee989
z6bb8897a5f38ac3c45758afcea9b045ff3bcd3a2dfc9754031cce2913e2977220e1c26d4c91bf7
zf2bb707839b1b2d586b68dfa6f7900df85765d182d0c069e3d5d0dd2386acec49689cd0c0388ec
zccbf0d3077edcc60df1c87ab9f09d989e366674fd74808373358d5e378851314fe08b5b24c2d6c
z6e6235be05413915ae0120c029c5d11f95a8874bcfad98c66f3e7e50dd7db870381850e45dfaad
z9a52c2157c023c2c67e78e35248f7ab22baad5e91c4b5f22a22592af0e9bafefe4bbbab60d95d1
zea9518163d7536540f2931f1d21bfa706619634fbf805cbb7b2767d7cb92b6ccb284147bad63a3
z5baf936c51878d717cf12c56fc118fe883cc07028965a2f6bfd8cc424701c5aed5ffd08472f6b9
z74db8c887beab06aa1559a0d34f17ca3dac0ceded7ff68ccfe126f36f45515ef03c6a66e745684
zbfdbbfb0863d91a02216e47e62ea63dff6bad685d9a555041c53a6b2a4445f1c7bdffb4c28fa7d
ze7f023af0dbad3e7fd34ac2bc70161dad1afc3d9b9c942896d2f41d2d2ebccb62af1535a44c8a2
z5c4d076a8da228f74ce8a31db7225f802d4600a5f66b1430be9669b8398396803e7ec2e0be06dd
z7e679addaa93781d55367ae7acdd6817e6e00b42e629b6032ba564d1166bf5fcbe03b9d1e854ad
z1b3acce261f53fa44b50426fc24e79f61ab40f8098fe010a5d00c79663ed671f2c0758daa72e9b
z5a0d3fa3d922597dff4ae61c669eacb82df54682fdfbb6c549127dfce9434fa6030c1b06db0af3
ze5583a29eb9afabbf859ac8c29bb7a657d6264d194a7566ab4732fc2c3fb9afb8e4c9ecafb8a40
z897090dddc10b554ff701addb4aa2b507af9c144edf849124bfedf753c5de419cf14bee81a7fb2
zf19869d13784d9eb5d145e81cc46bff79b9da45698b6291b30e24f81b83ee4cb2dbcad626ce8d2
z51ce469ba7dc23d119bab1e8fe245993e623e04a64d11ff7abd4fbcb20b0948840762ce924a007
zfb55add96d31f359421bf18d0c4d156d01de92d1785fb5414fde18da6779978135e042f10b654f
z36ef258adb180c333ab9cb33978622c9577f20e049bd09aff8f814345717e211b82a09f7eea048
z7c0963b605497fac6303e2973d7d65dba14e5d6679bb8076df1446221c1d134ef4ea19a545d8e5
z733a90149aba86b6cc3b51e2f49f346165940a2abe5c962b93eba3e2882bd721dfb188ed2e8098
zfbed31ae2ee6f9ac877de6c814d0be2482d1a8826253b074a2932f354d37bee84c01decf446b6f
z9f9264dce230d4b7799dc71f46fd7478855d41e84df986e0b89988d8e833fbc61cd53140dfb79b
z67b6e6c2e411d55ab49f105d294a725f340ac5445be013a7b7e067b9f0e099248f46432b9a4b57
z5a625b88bcf70cf02053dafa2ab3bc3c21c6373926e3ed1184d942e5a63d37fddd03f19f9e5179
z6ae978ad09be19ae4723cbf6cdd7c308db7eef90a6b1bccb564b9ba67c1a1bcda4dac5da0db288
zdfe1c5d7d818cbeca735aaa780cabe1e9be27f08a4cc28690656bdf001552dc291d6b342db3681
ze25c84bba1afb035c7fa8dc8948aa8cd95f19e5fe8263aa36c3d54040471b9879befc14b52b194
z1347be0dfefb545fdf4ac86a8d96901513b80f92d3c128ca816973f7de797d7e3d23a90aefa89e
zeb796db431ceb07b46c73f05656efc075a8811d003ba95bab3459cea6e7ecd033147c31d37d8e0
z7a02690eec3d734ddaa4e66410ebc682614c3aba301a5f1dd921a46b3f45a3cd2b767a1ddd87dd
zba8d1750fbc60ec459cae7f1769d9290840a0eb2e01cf9792b5dc79196daa15dfeb75e364a15bd
zb1be0e2f596ea1f870a278c8abebf9dbcd9b7ad480d32f68d3d1d5d7308772eb896a8192dfbf32
z8343680010488fca453d58ac979aa8fded13c781979e2ceb077787a2ee193a28a93aa34824eccd
z7db46797407969adba9028eed0e4ce3f309ad5e6f28229f960aae04d88d49bcaf27e3c6d9a6195
zd42d1316188b8c5053ddcf9470513558db20e703cc64e4850ca769ebce82be147e8fe633605f03
z7dc9e037e53de2114e4cca5793358b80525d602581a2fa176400965ae1a46c693f43174ac2ff20
zf8e946cb09db3a59814d1fcc66cdec3b0bbb3c27b21029bdf7e8bc9ad04558b207f5ef8ae953d5
zf22131cea80447b689037d1b7a39481de4536e81fd4b016253e867a7fe589992dc0981dada6039
z3ba29eccaf80af458418bd03b4dc3b126cf8bc9983be4c8e0754e7ab05fb4af3300716f481a899
z3da8d963f9d29eb763c703507696ef3f6cae78f5c6b5b16e109d992505679ddaacec75bc66b616
z2e907de43042392e59ec8584b29134b9667560120f9922d0d1df47da899ade831bd8a34691ead4
z460bc1c32b006ce4e948699fb19e9e368e0be184b1c630f3c059d7e38aacb2f972da8f9ff4df35
zd33cba5689797125f94dd69b75e6a6e6cd205bada5601ab60d89829a2a940895439202cf8713e6
zfa83f0d0825bfffab4c4d3719d7f7d390dd57812c8ae197bccf7679385a0a915024ab5234fa272
zc4bb96beec5d769130e630ec14389ef948647dca1fcdc9f89603e299c606e524c5d6ba3e668fe0
z736c7b3e4d5239c39abd6e6e54bcd9d62fe2431bd47f6b199a593ef7b6331631d6e74eb67332b0
ze287e696ab842b97452f7ca276d562bae0aa6162c35b07bc6acbecaef7f8ad639d8fb57c36daa9
z32287f0980fbd32ccd8b529673a8a662d0330e0838b42e720cb8f80ed459384669ef2647649185
z4118fdcfe25228ba7c69fe7f5186d19aa7400a565ecffe88536dad9f173945ff81dc40200ffd9b
z92118e52ca4b3504e1618dfbf241321a3f267b7723865c7e1d526e52547b9e17a124354d23f1dd
zb1c80b0509eed8d1e67997d7278eadd9368d816bc01df28b2a9768f68690d6d066ba6cb6620f1c
zfbd559cae66613888f6afe14b7a7cb1367261c00dc9e08dbe5c2641c108c30ba2587fed3538453
z7efd499483f85343a4023b93e2b8128c0ba5734177e0e2f04b02e6cb515f874b6fb403dfb35278
z583a173877fc96098afec5fbb4ca882ab9a9f8b16c7cdba7835fe126378836573ddcaeb33e46bc
z97f2a1f68ed12bf9ba60e986dda1158947299fb7e85dd458e993525337e7eec01d8eb726198805
zeb0700f04118347cd58cc8dd7ea0e54a5fc6d7bc5a57538587030e9b0a8c886d73ce5150c44ded
z89866b1d363b319dd1ef187917c555044b2d1764d8ee79c77d0aafc89e0a289c1fda5f6436384e
zafc63d4cc1c53081994a5b3d90e1731f4fb3fa31e5d07d977c94c4d57ef75f234cb6bdc520eb6b
zac704c6b0faef0700584f5c6d6119524ae9553ae34039d2df9bf527ea3e4b8ba0d8eae1de25e42
z31733275bcc91d07417f12dec5a9b560a497590fc586cd371d14e22e61159db4cedb9150324078
zd193abbded6d5ec77aeee34a84e51cf002a570e0bd99e202b55d4becb61f4253dcc1deff12a704
z5d4d4eda319bcb858735223b6917dd38e4a5dd0ebf975826810fa60001aec85d37ae119faf9890
z43c9780077ed3e49043561818fb285fb27738f23689d60f8e8636b1af0866be66fe96376aec5ea
z2dadac6627140833b9b59255c9b0463b5f6f8cab76b8819d825399a778568c584969eb7842743b
za91b01725922350c06deb273ec172542365a2753daa06260cdc8de06f2b937c1ede8a7624b57d2
z976f4c9e601bcc1849343f0624338adc1c2b2950e4b658242f5997b41a597dc386cb0b0368df16
z4abab57132a51c3e7f01e5ef33e6df35aeae0e6526520bfb3db82dbdeaba66edb68253c440b455
zdce0fafef15371d866fa454849953fb5c72c2968d1da35c92796d64b44c0418779b61977de7f68
z89d692079af2bfeb470fa544f9641cf671f93d98a3dfe6cbad2d2af9624df675557351b1ed56ff
zea36c9f45cf1489dd7fa56a901a7478d5a65213e477bae350f9a04bb807ed394ecc0fb8e588823
z905cc125b92d7e86c2a34142c037c951cbea6cbe03c683ae6d86fb0c98be3b5f3898be2f22474b
z3d14c5073b3695b64728e8bef23fd17f9a4525b58f5ffab26d86ab5a683040ade5ff35bc56be31
z33ada6da35c73a1e39237eacd830ff6a3f458a8789e3404a73875b2056bf652fb6ace52bd44662
z7b76d099aecaebaf35585bcce0acbd208e4366742f636e3f9cdcc0ca8be08d109379bce4042837
z0c1bd5ab7a9316deab6f04737da4ef8c6018f21f74ab11885a632cf7580dcc94fe88bfe83f2131
z21411be51e08520464aafd4473b161d2e3fb87897c7c0eb8bddb1628cde3e3902101b7ce586fc4
z2b0d9a73d0f9a358b0e920ea56e6a65138b268eb836efc4d89b58920aa798ad78ffbb478c209d3
zc8874328a17fcb064e938a84351b2cf100549c18a0039e3619b9ebb66178cbcec8900dcb20cc92
zc3985d2ce944686d2bd267575c89631df5b61a9e8269c73f490fcc4581a5daa5c252bb37b94f90
za56d6e96e70b62da05bc0ac5b1a616cf6c876709b55da7efdcd2831e5d02e6225baa5cfe1e4897
z049078418adfe3d0d5f5d7d1998439ab7c2d71a5f0f46761e25b3f1afccd61c354111b648f313b
zb48030e8517e02f2c0fa39a6f558961f5ab0964ac188ed1c4243a6aeb0a4c260aedfad4d063387
z13a8a420c60514033583df79608e160ac2db5bbab325afffa5724e961942c874b6099be47af22b
z99e465859e7a40a0000b17f305a737d1dddf2cf5992e74b44fad271249fe296bad59bc28fb5a56
z6059ad1d3c442fdc35cf34e4dea6264e62faa59eecaec85406a0d7e815bbd712b52ceb50f110c8
zffaec1829da16f529c7ef0f1f26ed84e170115e06bc70579e75a8b2020b2cdc1a06fa83cdf84ae
z5371f38135fe8fa25eeca204281c7fba262878090a7cd40b59491d6cf0f84eefe22784c1c2dbc8
z04b1796c90c5c8d17e9ea5ec2471300b3d538692a877f13996d9bf7b13d00587273627c545d58d
z7520f29af558628499a2efbf36714ffe3bc7cc4a4e9088aa05d486ca7cd1693128efbd8e69623d
z4ad0300b063e74d900b6dd14bc43007b362cf61dee077bb342b0a779e6f71b83f2a8296e6ed9bd
zafd8b592f806bfe1aaad3d1992ae22b1d42edaf612cedcc19c46eaa86f40e50f5130b2025e9f51
z37cb50bb2ed621226824694711da1429d0be15b50894f9cb7dd4c23b883dd00202e42c04aeec3e
ze23507c20a1807b4bb388d5fc873ffe1ed5b605c6e79ef68c937caab955839d92e788eb11120d4
zfa6f4405f45639d0fc52e21d2f4018cc0753639c6c316b89dab8a4fcf9ea379f15b8e410694ea7
zf300ae682b596bfc5792d2ea52486256b0bb0d715ea6936f58787d8ca36e4739f7b27e06c475b2
zd0690399cc4dc97d457a4238354b6e42c96d8aa8a36c978d240615aa6b3ec2a2f8f2e888e3eae6
z01f8bdeaf8f01c7e17c812c300dc128908a46f4974ea552dccd533d5025e289dd34f023665bc66
z06525f07caac307694eb2bb9c2b2a2f939c43b78e01244b10e597394df83aa5c265a07ed378f0a
zae15c484f6babb6a024525d0b3ce16e8aa
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_ddr2_sdram_data_checker.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
