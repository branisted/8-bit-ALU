`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026201628cee5aae21fb892db766c4
zb5b1406e11aebfd6dfacc9da5ec03b70c276807a3eb15e28ec7ab1dddec42388b9424ea285623a
z248195c9f894b36317ca6e59c86f11031163f5f5bfdba36b10b435d36514783bc1c6e60eaff7f9
za2b8eba90f8fd9a9cd7c932ce34efca1757e6b2718aa68644ba032b1bdd74efc688b935cf38d81
zb1f311df3e5b8e4d46dbf459c824f309500192485674c175e61de609f1c94488da73614dd500c3
z680b7fbf510ef6c68927870992ed3376661d943d2a929d90faac51228c485c2005ea015bbf306b
za52b2ed3688d7ece69bc3ddb93a45ccc73f6e00673486a8bcc92acb7d4412090924945c1f1562a
zc5e0949f06ac734085ed2107e4aa9e39ce4ccd2716381ae81c00f915da3dee1704ecc26765111b
z37c91301861edd467e17607d70795d4d591506508eb6e0385dbe68330b0508d49914b184eb5143
z0de35e4146b0a895227cd1cebd7fe0a0e690a65144d58346a34e920ca3dcfd3b7bae8a9a5fb43c
zbc368eb9021d06f1131291dd6d1fbd1dddaba872b9157058284d0dd16e970359482f68631a9805
z07532590445f44c042503fdbdbc91482b4eb6dac87dc601d1d5eab8b5a973c4b2858676ca6097c
z461b8368223510a4d4d8eaf6eed8ff9c34ce31863be15ecd5c71390aee0379e11ec682d501055d
z0801d515fa3a1e2df3b8ccaa85693d91100f6f329e8e63185ca8a8f41d19d17cb0236aea1bf894
zb41e86f4a1f625619a63c6f02cd0132b6fa821f8428562c0a890db7d5ac04a8cbea4374ad26af4
zcb5b63827bceadb0b83a7cc919177ad33e4551da575cda6317dc56887f652f5580d970773fee4c
zd691deb792c51933f078b10db37fe2fb4181a3b7e316c99757652c6ef2ec0de39f57e283849a70
z712b5cc5acda5c26051a7ca93b69db58bfb2cb084ced13a2a49812262313bf37e7342c66649b5a
z5c724715f0aad5f3c3a3d350caa5d58a8d9a0a096b6e4c819e1c845041364966b48feaf6dd02ec
z6ec250c8de48798a4a339d1554d5733b7b7c5ea5676fa08b2337ab4304115c3d63aa770cdbc7ff
zbdc8c09a237ff2e329c01852a311141a6f75ee1cf465825c749631815bc3cc3c805234bcc758e2
z8c5c18a385bf303af73f4445ae4f84ec9e7ecdb8b0d07befad4cc80b159ad29915927dc4d5727f
z43506d46a9e548f5a292aaf29c8c08cbbac65ebbf2510e629d3b0f3a78b705272a55d4141166f1
z9dd88f8fe0eeef5a13dd403a3ecda14ad487fb3c51c39988254d9af8ac1c4d7d89532a83186a00
z6b8b699d00b6196f2c4d58ace32e6eb284f0c68be9b7f57af4bffc92d33b0aee86d686149cc474
zb363cb97933a369f3d626682ca2f44862f6a454d108d7b32263c48d9c909bb2190ac6b063bfa6d
z60726089c68525ab2a0fa038ef11f84dfc0244e04be3beae39d5f36342a0a5e3879a83783ffbd9
zb43888c9827fcde00f23ee571aab78f4807316bb22f1ca69ecc243e96314f22e24a0026ee84571
z2b099e2b0f4aa52db7073b8db8c3a8b6a58c06f08a571230fd3bfc650c2a5d61b9b6620c141d61
z43684f4535d1798fc6e3aa269d953023f9985e0d920b5eb4b508d5b7604da6a9ebd60f6126d5db
z2587962416810661d08c9c610ce2297e51cf6195710fda7cc333be42068fa3cac26b77e58357ee
zdd933c6c2de76fb86f471ffbd6f9db98d739f26661992655bb19112cee3576fd9e6f111b2a5c11
zf6c275422967cc2de277b93feb856e54363fa389863f638560bcfb70465ab8c09a4c47d004efed
zc27fe9d129b8422e94f7b380df879ce987288fa984a9b304247b002ee87ca7568dbfed5e8bffc2
z5d64bb5fc691c23583791557d4deb0fac6634e3803678d2a09e14c5d78deda188dc82839fa896a
zcd5b9b1c22ff6641ebefd7c3e085f00daecfaf4c44bc14085574aebb543e27d82e591dc3dcbcd8
z24ff0326a55cd42039fe7a5eebcc29a4ea3317ec18dec7e483647f1eff7473f0b1e4ddaca79f7d
z8fb1bbc4f6544d6109ee461fc68d5aca553642612c174fa51c64c90bff301e8ec09023e32a854b
zf5abcd6f0612cd5c4a4f8df2bcbc7668bdc43f903d62e42ad76f4d7808be454a5719be5c24b7cd
z3d32acc874a52040143ab0d52ac0888e4cc11f35933f53b9e9cf0e6f6ab160638f14924386c6b1
z70c776a98f954f429c40911b844cf21596ba875f1333e3cfb3c26e7d444f77bb8bd13826f27e86
z48a9fad143074268f82bc7047a626b2248d81d970bb9a3659a0219130cb3527dd8fc0100b6095a
z88e7c0ce29e94464c8f356d53ce4b0509b29de20fd4f0047d65ffc1b2639787706bd505275d88e
z531e893cf0bdd3509d789e254de6242ba13ed25990dd76a86ecfce90fbb8672866bac048c4055e
z033de915fc02aaa66912cbffc9c8389b50a7535dc07a457b50060263c36a5e2517fe16cb469221
z69c54ad39694b33121c586e71d893774be2a027fc6b832a4ebfbb7ed05d0515970ab2678b5afc9
za1b7522c95be200cc077e6c3248a32071cc90ad3b2a348d041f0f559d4b49efc575ab7ceba1b3b
z22a61c3c5d3703cdd74ba8048ee8bbc25bfd7ff0dcc3e16b326db280e98f9f9229f397840055b2
z5ef04871b0a58d0f80b4442b8050b9dab6de841aba8fc16b9485538146ecb4462d1ae05a82b49d
zd0e1ace2612876234dba34fc5a66d688eab3e50c709459642bc568c249907e71fff97ef16784c4
z2eaf48ba01e41a1c5a1a3d4b9bc7328f14f1651a822a774daa4957d1515382a92b796a88c5d562
zce92840f30481a5e9bff7fbfba044ede018b470110f8ff0cbaa19a4dcab8d3310a8531687c723f
z733334aa5a8ae215ba5174fb2ed5f191ccc0acd649e61c044af9435bf08ddb9dafcf9e57847fb4
z2b5c6acfb838d3908b4e9196258aeb5f94d86d1251a7499e4b29f4090a227fd9b74fad55e975a5
z9aec8f13fa7e2911c97373dd6683c59b1fc174604136cf427c903355e545c0acb98d26b01c7016
zd3478731d2337c3261d98c8a9cc07832abe55bec6bb78bc3234718c0456548b368455f8e114c3c
z236221502e4487317cb3c6a52d44053d00afc01cce9757e53a304d9cc45395e6b3ff1ce1ebcea5
z299478f29d7d1e1e28a97691baabd73853bce2be91a337c4a9316e8730fa8be84c3e0dd157394e
z231868e4df7341f59a9b1e56788f4cd730bc3747a6a795c214966e7afc4d8d47a04f074d843854
z5ac5540d2742467b8129fb31d55e7b395bbf09171aca1d6528cae742c81f1984648aed51bec341
za5cf9fcea55e25ade739a2ed8eeb58fcdd9ed47f7792e80f0dc23c263adbe38636ca0e3daeed3f
zf11f7bfe51e328c3d335c48320abb9ed1871ab23012729546072928e5b32acdff9a75a94e7da0d
zd6175f89badacb91930a50e019c2d5036bd1f545eedeca91a3691f92bb2a9bf34bebcf7724205d
zab82a9bfec274eddb889ce295f98c7ab87077a76c989e2ba4c94a4cd94cc4bc8d771d7dd32305f
ze0ed332a9b14e0a13041b99a734416f4214fadfef8cc8a49193b6952daa6a905ec9efd6a9667b2
z04f022bdad80296b9528f36600efb6cb966015b9010ac59f6f4e20490d4a6af45e499196721f22
z8a3e0f8a2e00b2dfd63d46fb3af57b6965aa809474fad9650465df9b59697e16bffdbf0eed7910
z8a141da942f0c4943ef88b101197c51e1226325a3fbc691c93811cf762f2175935ff69d2583f1c
z01b0b00250687ba90b4961d725967e2870fc1fa2b9dd3bc2631f1e10e0cc51167a2ce106b49829
z9a8066694c7a78eb1f221bb324c53a2b711a0b21686a9b5177d02e26e1403ff44594595a03d150
zb70e82cd26f7678b0eb5b345482ece7f699852486c7222bd08c3ebe43dbe18ceefa20d0bdc4836
zbf78025bbf78aeb73ce7e4b30838fb58029a6a23b16c21e708a7148b8de292d9aacc65f866c8bb
zcd5690f458f4bd5ff6fbab3d1d646fb69b6c3a7eca6a435cfa5b1c422ca218fc02c24cd36e2e00
z5b2b2a5bb804068fd6315f11a3c3220ff62b23c3c13516f6f7995ca06af638b08e444bcb1d6f30
z4494606d045588ee924e65c246a9a1822170120abb708763c6a20e19855b71973214a88a2c45c5
z96ecbebcaf68c0e856db58c95ff2c55bae2a6eb4176d3b91553b5fc0505f1f3e6a754ad4946679
z1611698e4d964e786e76ef05def3a039eeaa88d62a8ab64908f9ce08cde21dd17e38183b3ca9ae
z42e74719529c32f6abd8179b9c0fbc2ce835f7d31bedc0649563e986c03e81d791f6c379e17c92
z267e65a071604c94c490bb652c94c3300594c5a2d812d87a5e766d354745f823c138d89cd1a672
zb88a630a0a57a3dfddc42f52caeaa4ef0186e966e7e8c9487c6d77e8aec22447f91cc3e69ee2d9
z7ab3939df27f0a022642598664d1abf755fe672f72ade963fbc85c47e909a11fa7813966d83c1b
zcafe9f62f2d9317f780516c5779759d983d67a787f240b5755e3ebbb2f91c2c7f489da7b33e324
zf43155f5f82b300659e4b0e47cffeecf385b70d78052c29ce12f78e982ebd394d88a7141ad996d
z66a65df479ed326980b8a830d3d833bd8f953dd83560eb9a316954d6a8b87857ffc931b37522a5
zdd58de9ee7b540a9bafe22abf5c43640cd2484f15c1cf378c38cd0f1b006fe24b5bf67d9703244
z74480b655e871c74354af46a45c176eb3a3f7952e58aba1b39429dea5517d70424a9f902144954
z7c00dbbaf972ba88b902c5374d0c7ce92959d3c328d175916dec602f25b05032368f00a2e92ccf
z082f532ae0b1a1bd591d230833071c46b74862b76aa1c3286c39fdcaff626f955ccb430f62c145
zefb7110542c0d685ecbd4daae77bba29fa9fba3c2d613e6ae568bfbb437ba5839e24c0df7e78ad
zd82746d832a2515c5bad4272ebd00a720998d89d74bd5c0aeca15efb7856533df65bbe5a242659
z3dbf5a2af65d1c849956c582ce735b63f8d60b828ad77aebda8ea99f3340ca682114b765b36769
z2711393dec47408d3e84081f0bebb9f25b9ebc5ea445ca836a0234c8e540a7793daa53b2941b7b
z21309658b239e562c467f1f9f447caced21c3efc5224165e4e1f442552aa16fd0fdc3506d2bd3f
z1b8863be4e41fe90df8b9b5d42a665e5cd62389d24cdc9d18a290b403185d02f763fd57c566b7b
z950c46a72d678e307fda14db881b677a08e6940da21e2221685ec97cd66962a1a9461316ff0faa
zac1ccc0a326d15bcf880249429dab65dc6d68e21116b83da47aa39276fddd5124ceb918a1a858b
z8409d99ad53b9463e690484ebcf69fbc37f28cc6867ea45cd213f16fa7c31052d8002afcf52b6f
zada0e9eb775b275e621e2e5ac4c29281ff866ea47de79f6485ee57094c644cc3c8133a50cdce9d
z823b7d2700b89f70cb74573e14a230ed0b6e6a92ea4734ee76040a99c7eb8e97c257e4345141f3
z10440c57255009a5574aaa3dd7556e1b321ffb58aa23abd4748aa2e66934f4c64b4f58b2519191
z0102535082680365b0011d3087de1a0371fe96f51c5d153c926b7720845093e833adb6faacf7cd
zf29cc235e94d82a52458814ebca79b09e86461d81af33c570cc167dc559d99776fe34749532820
z86e5e12e538c79f7dcbfe1b888d1bbae947162e4c8b0488aba08b1b1387f8169fcdf49cc063edf
z5b557f4d688c5c549f94c601bc21df7ac489767886de0ff33e53ed911732c638a3b07179ce7036
z04033f5ed93e15ea5baea3d8785e649404a31a4e6bf12d0a81957b06bb3f23a7712c2e2b5f4d3d
zd570e4f3f809efa21ef0578d2e953a0ac3000bb22b9512251caa96ea61c8bf1d9f8d71b2b8bdd2
zaf19506f61845d192aa6bb912b9d2e0b19e80c6eea5035f8f0e22c7c89925d4e598f09dd43d370
z620e0617a493b74ef4ea3a12cc07678daa638bbfbf0fd60c1ee556c26369dc07413df2ca3e3e3a
z2f883abba8c4bc3ccaf5a887ef24cf3e84b15063547b4016a3ec4d3d431c15e8bb905b0d04afd2
za69a4f3261a94bc938b0d7ccf3a97eb995bcb963b7be6d254f2983d68b2fa155fc1a91eaaa9c27
z50530fc1d083c47cb39e8c8c1bb9e82f130f577062a96bc1166ec6f7b8923b0988f68dbb2beca2
zb1953de65df5e08da807491e63d95d19ad59ec6796dd452c3c6d24924863b62391a6401f7e94e5
z9dfb03588f49950aeb5af0ef0fc81f6530e7f8d8042d248eebd6a69a1c4acca8d6ff5c3fe17d14
zf7eea7f133e5bfce598702325d118e96e3644c8c78551616576edc367cf7400cf99d3550541425
z8f801dec1032d7ab34aaf52a6d96778db45922e1e8fa255fe6b02dd263e00f15d874bb5eb25988
zf9497b01b1941681f3185c5132c7a1dc68f9d06ffac51a9bb0d0799d7e649dc81c3f5cbe387da9
z71e1b99f5a05f851ef14e9ae118b9115771ae9425eda1b95735fc5ddb5cdc9a3233d86f4b995f9
z4fd0f8f538a70c7792bacd9991c20e4ea5d385aa23250b35e92b35f8501e021754fd1475ae2171
zc43a8d90da651eea19d022a0c3dbe84c3ac12bcc4fe80e2beca02cabd54f9b89d98698f32c7714
z575d60f5ab325807b762a9a0d332a63efb9e8f58194499ff4f99509d9a85314ed5ea61a4a35d1f
z807aff1e0795641bfa5a8b19b2c8fdf456417f1c733c5d43320ccd2ed25eb1ec8f0c498044fe7e
z33d62914eb6f3fed19b0ce01cded11dd573235f7c9aafe81386aca56c80d066d7c065ee3d6f8bb
z79aaa1ef49ae4d2e0245ed7bb9849c406421bab7a3acaab71703cda1c9247d52711f884c98fe53
z3d035bc2e7a4dc59e46fd715a16b32df02d9f86498808c56771dacaeb106c1507fb3592125189a
z264a659afd43810f85de08ac8569944f2531352bcc03936e8830d135f64430985cf9c72d789da2
ze370a197de08eaef96b881bcfb1eff08bfdc606cc8df6212ea3b79662fcef4a750aaec67ce9865
zaa93d129e4c50a0c6f7ad93b23c28c113cf4023bcbc3b5b39b679cf24726d722a62dd75f89828c
zf497dd85456c7860d38eba1c2c26fde7ae383e624e9d693fa9ea8f234ed6cdbcab442ac7b196c0
z575d16ae6dd9e4cfa2a145d813e9fb70a13a4337f0db55cc6b537047d0551cab4dfa9937862188
zd67e4e93d0f0e579c1c3b33740c1721fdec07c599a06be9d6ccc0fffd28e922e70f38595d89810
zaa8c95d47fc71a73a9c159d7e42a24e926ab05e5ba274a8a5d06bc8b91341f27d64edc2893b57a
za43f93814a04afe8f157d117997866b503c5a4fe95213b9bc60647beb1ef02d9d042ca9503210c
zfff52662cc4cdd1d11084f0aced83c592c6e90c69bb6feca012395673b35ce3c1de0af0a942890
z57ad30bdedab6d0b5baea357ec78a0f56b1f9045ecc27896929b2c5acacd00e01bfd07bd75906d
zc86d2d7834a6d42cb1cbb4d36176df8aaca6a7f081cf8ed0ac1778dc5eab70cb16b4de4369acf0
zf31e3f67497ceac62e09434e3bed7e8460ddbf176b610b88ebe9bc2f75d79483bce9c31a548f1b
zc35922ca23ac064b31a15ed59eca7b48484c5c7e8aa0c429a1995175d954b38c9f15dfa4758b43
z7b83aa41b11568b94ac000a9d363c2e9fc31bf9b0af995f81cc574ed0f878a6197f832043a3cae
zdb01dc13b8533a7b82713b0dec5514e0b6defc9145ac6118ee9b7d1e6b4ac55a2e365ed8672ec1
z8b7b941235dd68df93db19509e09c8fc1752883d827c4ddf0fe0986509b4d5fc5c9501da3ccd6b
z809d73b085635a48a5dcfe3d5687cf407d2016f701b879019c42344fbb137646d23f5d682ce25c
z55860b27aff03e70bde34f79e6ef62be18fe37b4d5e480f483dc6da22229ed2593dc6d58b6fce3
z7f29e1fa91e1ad2e35d0bff0c66b96b14ef8a70e9bf234faab33307caade44638b5d9d66fa9c31
ze8ecced690a61ef45d2b4e41a0696f85c248d382ecd5bd4a6bc84445b521adf57af909ffd5c347
zbf50d1c62aaf27eeab6c974f19741c5304767a7843e0771683f13fb7dc638d01847674b6d1335d
z5aba32ca5aaaf9b32b4adf44467487371d5b94e1fed41d4a883e463610757a14c2a9cf2ef649b3
zd0ec0b90ac7522b5e0004c47cf95d4ecf12ccd3c3ef8af6cf2fc44555d8e907c6b086c01fdc7d4
zbca3b6a177de7750287b3b1229e6533635ddc3decbb855f360ece44a82b43a8f47d8e3d4ad2b0d
z0354439eb8bdd67a584cd3f32c051315abc067ebb260a7a018d98be619491d73393a202233f987
zc257b8c377412ad63cb07083c31399ec3aef7ff404ecc4470fc99ff3ad9a4e1047c8ee50ace7be
z9d0c0ad1ff87b8f265ae41153809156ce4b37b6c1b134c5a98a94ec7d856dfb0acf28037c2b56b
zb512d353b4b4329e394089942355c4313d69bc858d619dc18ceba34c85c50186733fe31ff3af78
z70fd6832e5baffbdb024a0e852964e89a9bb75a8e08fdd9e78307eee201df9b9d04d338d3af93c
zb0b2cecc183f9ca70256c6072cdae185e08c921a296fd06ba8c8e5a0b8938b1af496a90477865a
zd29a5a192f19c078008e3d3155adc50bccca6899175d2a1a1a48d29ce2553f0689fab35fb9ca30
z19606b7eea4be5339afa9e2f9345e3a5152f38014d4852ddb32ef9ce1174c7ef0fe1752fb08eff
zccec21f03ff0cf90b4a94805a0a2a1273c0390e82c20bb1f5ebf0c752642c81e43fd7cb3887784
zefd81e5f516c2432721b18695e7576a77d1c92b4420ebe8f304b48b5b6aee6fb0d14e7647908bf
z755cfa6e955c3097422c9d8f003bdb5f7628d34c4f9ed7ea56e7dc7a2395b9dfc01e4b4e1187a2
z29edd2a986811f30df1db41aaf52befd57048e3365d81cf753b6be080b6b6b7544afb68d7a3b01
z0ed0b4fb84635a30479ba7cec98769ac0cef6302976e0b0c2582bb670976e97bc44981c35c2149
z4c927cefe2948e8c31be662cea635b689cfc8dce08171b422b55e36cbf7c85d6ca810c35104e79
z17857c70a775b9aec366ba6ea49ff21dd4bfdf7011cbc9f1c5a4e4ab4e5b2d77c114a97dd212d7
z71fb8154a69d97e549c09a37365913f7bcfe3527115674fad3939cb5c642c42eadc3cdf93dd22d
z90a04eed097beeb3a96d4eb131ccbb98be0d4f5595be7631dcef1ec3f3b321c1d61d13e37431c8
z324034bbddae0a3d8cb0cf398a67d14a423ad62b66c3960cc2a22fc7cae8f8b9b23e6927aedc01
z210e15a58a2183b47499296e2882cd2272094545f8d4ea2758db3b1f2745c319d969a0a276e5c0
z863ba7ba396e1f5dc59229b131a3039ff150895abfcf833d4b30523b246d6c64e5d83bfd9b1454
z7a0659580a24fca4c0f595b78818727f687e68ba40cdc08b5e47ebe4884ff60f997a4b5153fc2d
z5ed52ba647065492d78299f38c90a5549a9b7f4bf0083283709481499b398ddabc4e073a84664d
zbd4913c57d8abb830036523d9406c9f3c86eb0c77b13226ac6b2ba6263abad4e477303bb5c680e
zeb921c540ddc5de1bd63572071d7df229efe0cfbfae11285e35c353b7313d746c7ce9e5226e74a
z1110114c7114f0ceb8253a382483246ad16035b5bb9bcb2baf59830d4ba1be2386d7ba9f4053b5
z80bc3324b8a2ff84d0a9a71597a74463a8a833158322f00b249928df749dbb23e4334b8e227464
zbaeac8ddfa92c3b0e8fcda4442001ebe138f3050dfc849704ce2b3f4c29a88378dff54def3c539
z29bc2eaf33409cce47aa08ebca3be48300c3cec0af1fa82254eacaf62b785c56c2ca62e42f8e8b
z006941d2b72a779691be7ea4d782caf6f3bebbb2e509e9c4962fb6fb404d10607f9e67f5010f55
z2b5cb6e24144e847a221d5b53ca9f7fb0d58726315088ccc827b11fa126137924a4e8a767cb585
z19c5c5f75deddd0b7ab85027007fe9299df7b66279174566c355a56db4361edb4f8433fe3b4ca5
za11e21161e2e8ee4e116be82e88a05504c01f704d24d4a50f367025e5967e0ec686bb52c9d5f8d
zcf68a7ab4a81bf8bf7f495ad3161519af5ad371087971f76118cf45a40a98bfa91fb14583b85f8
z2854a5be3bfe68fa314aaaef3e16b91a8b24e440e4df13a44e919d16adca171302235c3a252763
z3ea0c30009f1405faed1f20f4770f8f0fb4d79c36fd7d0668eccca89bdabecdb77f5ea7e86e752
z62a7c02dcdd02b22d148c31e2bd0a965e88b0d042d2dca9bccd1e0efd810ab7019a63e4fe4e4c9
zcecc637aafa682a830630f253c274786d5b87b48f5bdb817537b803e4d0e4e786816f78fdad2e1
zab75fbd79539c4066884dc598f6a4494bf982e0aa79879a46d5efee73b2f606e9ac104877b2fc1
z8f0e5f93ef10529e27522324e8edaa6d44d6244af37a563472644324a69a33f05bcb64946cbe74
z55321ff9e69dd9a6005f710de46b3423f7b247463fbaa305d252bf63012698ab4d7ff9652eb1a5
z18cdcfcbc0b433877b4c9baf8043607a36972d4914c91f9d356862d170381374e0b07ea49cac70
z802814a7a7a9d28732e74da8042d14b2c77c8d4fb1bae0658304dd59790c5ffe124c18438d1c36
z40212cbd80d2294f920a67c01b2a4efb872dad91cc425370a55a34e9bded754dcecdd110604807
za32f6a8399d3c794c23c1d08e73c4528c298aea610f3e80bdf60f386813c991f3ba8450689eb1c
z5216e5b8d621517dce5b73234cc78818c8b428fef43469e399579547c451708a1ecf92b297860b
zbc4cf53233a4ceafce588376f546edfb969c25426e66ebc54d22abd37bc2834bcbc7002878ebc6
zd1fb7c5fed4fc1a07bae63f9b2aa4ded7a8b62d198c02712117084f8d7fa1ee1735e9ad9d05a0d
zdc7178888f44cdeec325ddd5910b3f9ee97c65b5a01d73f4f389d1271c9572847ea104a375a994
zcb1512bffda9810a86e7db71b888ce3a791168b262237873b98aa7dca2dd74d996e0f4cfe3156a
z27590dc1ebb07986c4d8c3eb3d2ca82919784d7c63dd382ce0b85332a96aa0250a4b8b1b7d9f48
zcd1e0a229a673ed783553e1ae006177a4c87c752f86520bd11bbc6e2b4e28b029d33d517b8949b
z9f4460201a2de2c5e306fbff3ba12d308bdb3bb3c640766e20622247662407060f7596f403e65e
z852310743547d8d55c99e818e7fdf6882aa0b211a5df7de40d0b792b702923295c763b3c602387
z9d90b8eac25fbda906d8b72aba4a68bce1370b7623d05120c12bf24156cbf72117fa502f575973
zb09d9dcb732e8d396db727a3f4ae8799b1e475239128d6eb38c415ba86138684d56293cd77fce3
z5f3919ebeb79fe0c06d005e0b7348777ca215ea46b3a560e84e9208245479312dfab12d14daf1a
z354e86182324d205b7b1a2812a3784e71b4b52a41cf703d828fba4038e3f52fe89036587e3956d
zb101bd874e620a8e7a3f06fb25e46e3ee17f9006e9580d83bdaca1c8e8e4bf0b82fee8bf6b3144
z82264e7de31bc590bbd853eea42545b30ec8e808bd9bf100282f4b071229216d8c58f87fb9890b
ze4d706e1fb1391a0db6754eb12e93438d563ae07c778e3e0f856259f114642397487a26ccb7596
z3ce0a3b70061bca11de0012690d355d02e76e8baafb643108df1cb74c7a43e619a56238c3628fb
z75e2630b6f91d090ac30a532701b95a5210f6b8c72765029e4866d7f923b44b3beb37cf6f989a9
zc8ed9f32245e833f0e98bd7d54745cb1569a3387abf8b5f17551539d64d047db86ac05144d9600
za2c401f6fad02b70b09f8ed6d215ea9f2572bd77b041bbe9bf99767a7c0fafda30a03e34ab42a4
z7ab383f32baef9e6981ffcba5e7793c7c8535730f7c0007c2ad85e5d149fb276a9e519ce2bff5e
z2eabb0efe0a10ad7a204d9873a52fcbfddc6dfca9f9e9ebea7b6cf366896fba06ebe8eeae3ca2e
z1584acd819c2a9535cc3546750617df06d14307edf39ac55f6caf10831abe60440299125fd8868
z9c19a334209155ebabfb55a1f9d11fbe5baf4ced2e9f3b76fc31d5fc6e340e00c29bcc50838d25
zf720ae731e2ebd9c0f381e8c1a38c6241103818707a632480f87eafb2f76de9c2325fffbf75929
zc6e415343d4fe9af2e68fa934ea1bc67d12cdaa09ea274df9842fafca18c266e2a9a1c621c1b5b
z4657b99d9dc2bfa29680e313b9509c2a91ce4df5352150be320d13e7d2c4c7694eb3b3ca361fca
z44d113a9186c287eea433ce56fb221c845c417e559014163cc4f277636144a291f3e861e24a177
zfac3f4791e33813f3fdb66181c5e7015057dc292ef4a1361c3f607332c18a557d0dfc6d1137fe8
z562478282fde55d894e4d21548f6ad87863c8a6f9ddc128f7876cb30ada60e3c3ed7e8c77a4ad5
z6b68ac65ebf6c5b4cf859f56d3799797d771b2addc6c1b81d1782328b0a6667a17eb41a1536e18
z0c7552142298cdde760796cd3da0cca0abed8a99dd38cf643063012372465086fbc23ee3b07e3b
zf614f38ad2dcb490d6d70a43178812b59e2eeda6f3e1a5da13e29700157201454bc97109bef36b
z795f130ba24055ec3a59302f9e823c986e8d3d5eaef344de0b8e9347cf4fcbf9d52fc34bcd0e9a
za8e5d29e9f0dfd9e2910c16fae1ba7b3b815297a19ea261ba3a9d3000668836df021972629ad17
z454220e08ad7cba531e46a665ab4251df6572d206b46227b84c90cb51fdd94e9b1968fbb240ec9
zf4c11ad6862998403b7cbb75358a8bb943d693d89505447e0c0737d219c837cd39bfc4bc83cb98
z69bb46aad3acecc756a62208f815ccc376f03b62f84c6872ce9bd7ad7cebc97d57207941cc7e94
z647cfa5d7be548afec8391e1771aa9c29871f7f410348ecc959edce2737206d678281e2b9fc800
ze1d200219ffc14d9c101fe9e0079457cf6eb7468a6579887156de2f6fa6bc551284ba006174cbf
z832060e5d10aa44c93bd60d28c6e19162d4d98d6a316db2902e877fd741c0ff35b791ea24b4257
zcd836e8db50a19be57cb51e06806dd808b9dd407abedcdbbc4b7436310e3c7f989880c3a80dc26
z8619379d497c2ab300d565ecc9f04378a5dcf8cb7f723487a9d09ee916c471297695940a136f75
z1cf1b1b9e1cf45dc9cc0135a74b50e07e371847cb82fdd62ac4249fab569f847f8583429df0762
z5a6c1aa76489b3aea4ca4d0646cb5e5a010d771d823f363bf343e7cd7faa4e9f0a6e90d652a7d9
z7c53dd3a0780d0919f6e94c36255e4af6e1a5bb44aa7bb96fa4848740bccb1d97033d887b095f5
z5158cf60fbf9778c1363b7bc3d0708ef96de14cac830221077f725fa62f5761f59343cebcc2fca
z0b80ca5e6d6e70bd2822eab2e955fedb3737358d9c93c46aa9f2da7467b459535a78caa7544f22
z96266432897cd558303854f827236b0bd41a07790b34548e22269c5ad1618a7fb232e8878f3f16
z9770b3ce3b1060f17fa0c89c8dfacbdaf30ff6beba1989a565737fbdb709af63700661a63c5411
z62554dfcee86b3089c5c86d64bbdd68f837e1184b1ddf163bead8a29b6387e3cddd757b89b163b
z231d05075756c2197dca3b9a91b1c54ed9b346fc8ea456e83a490e09441581ae5664f0606d74ba
zd119fc2b405bfc9e4cb5d8ff151f01cfab38eeac25d48287fdc146c0b3f1393946ff5336401872
z6cd09d6de4efe1393bd78d19e071383ca62f46f1eb06664b6eeffabccc22b8587812b9def63b1a
z3062677c01d8f1acb79ff0105e176de8b8b3a40089e3ab58f3e70b9173d0dd6f0229aa6842b68c
z4c1c26374eb53858c40e09eacaf704475e21c46b93bfe15c655d84756e7d1ae4b400b7f2fb16b4
za0d90e68ad8994c0bfca4c1f53578b8b217a1bd4e59cbcca74e1e160e667214e51c9570a0ec4ed
z063704fad416eae2698f9b4e613f14e5c816accecfc776e3ddae59d0e95b9875e653f84dbc11e0
z685bd7cc78d9bc79e9f793cc3a47f4fe64c736c10d5c5f28157d4db503b6f6a8816369b378a999
z637740781f20c00e17e96a4a7ca6670dc0393b869191edc0ea6b9b997045b81fc4ea83a595a17e
z2a81e104c2879879b9d03ac98010d2a93e2b3c2976d76135a3b06b8431450531add9927e776212
z49e603d9487dbdadd6fc33bd6d69c3d23c9f1423e5553565429a62655451d739f2d0efe5465b81
z5a3d6dc12ceb746e06e95509ce4ddec336bc2cbac10d6119b287698dbb6f11c05d33ef36606aab
z8eab6eae5925e1bafcaf68ff5dca069f67328177f1b52b9d84a9e4f2e3e72481de9edd5a7157c1
zf2085c8fdfb52c27fbe2c7a525e5ff8de95f0570dbfbd5c07fe3884d343ddbd514bd46ead8b48b
zf52fc6c51e693bf2dfcfa44b520a2806a81b4ce0138b858196d761f752a85b8e11945c6f8e9541
zca5d2e1958d92913358b864f0f2d1f067e5a474de161587c8fb316e6e4f9320d746c6006a5ef0b
z9575a565b08d34813127389d0fe1f6d2209c3afc13c1c015f58fc99bf928eb784758126f7a653e
zef658b52dc65f3310373d205dfcc32b2da5aadb17a90c905a3569a02ab8e29fd478f9e3ae312a3
z7e42d0270dcc0253ce6b3c204332496f11b69162a3b1c24bf0ae599a3f2fb13c417c1efa6c73ed
z0f568e00770f0c1b7bfbf62b17304b3f889a51c58cfd2d1cb323d44bbecb540995250c5b55855f
z419955d3ad87952fe1627d38ea7a1e3335b63c83714d9d6e7369e5d25035df2e57451063fd10ab
ze537cedd532a0a31b3f64478f074c5e12252514a857d45ecf984168cbbbe05350abbb031aaa447
z3e6607632313e14b7d9b6bcd0c415bd9563e89b33b2bfea84efc8c648f4b9bd46076270851a651
zef51329ef7d8fbba8d6356a0dc513419127456ab80d54cc0d1c879d974d7cbc77b390949fbcf78
z9efca94a3f9f22d9216c95ec9fefe4b563c8535b16840b995df2928b94e0f9b38f088bc046a6a6
za1ff7326d22a04e4d11c720c462a87779ad1de0f00c5dc09ccef40baf6d58fe93ece9c1e70f693
zaa74c0ee2263c4993027d8a148298dc6b3c95342797e53b93fde55cb9f7ab6e893fb2ad02b0698
ze390ad56c84e6e0cc0c45c521c02747c7b382b6db29eeda6b9b37ae914b94a36485b7aebd6d4c6
z889ba3f26bf31ff44fdad1ef9d46d954680d970a1d11aaca8731988a95b52d16db3ce761c169bb
z285965cc43f2c9c142671be6ec098c7641ebba1b4145c026dddef61f247e14e533f9dbda6a862b
za48971a7a78aad17c6b46ee1d50b17c19f5429205bf1623d3d3420a9b35a0730357fc4c20fc360
zfe0e90a2f46025ca18f291d3688b458fa2738093b4febd5b67c1393e4ea959cb93c1bb9144ef5e
z6fd73d3f8c7c0d301a7bb72d11b9dbaf4fa3d0d4e3a9a1010a3635a20f27931fef61c12fb8b968
zba29844940b49c39176feedc3e45dc4533d7bbb9eedc5c201f9571386c2589376c848cb9b47248
z79c4a71237e804bcf744f3f9de8ea258791913914d25acbb774cd35f7302accf44d821857bb345
z032bf81588d537a9176a8a9bde2128c1ca32eb90c66ee1c4f7136f02cfe3244c190b30c015f0f4
zcf512f41dafe1c8b787da35add80b3b654030f96935202d47ca31f58c544fe72125104fafc6590
za31d7baae17b64180ea65a52731cde96988f834d6dcd862b9a1812358615cc448c16564641e4be
z0d94f52c05bd9a3ea8b630b875675d65d925d23f86ee33dcd48c52f9d7e7874ee5496748761738
z01b97f9b9f00d908a6ad295ba0d928332238677c4e9a4f027b9837846a0775de7d00767ce834c1
ze1859f73baf8bb98d530a160b9ac8f69bcfd74c6e47c15667f05f80c122832a70efd129656f2ba
za12e67172022bb35b496c240fefb286f5f2d9427f732b2473f19eff3ce11f0cacd4422ebaebe42
z80c8fc4e94f034fb2598f077341ee68872aa6f1455513421b43bea2f8812411fd1aa0a83d43f7a
z0e60d3510e27a20c3ed50b7ebe066c66cc3e93a855a2cf04597574c28496f0ebd6da2c1cb13fec
zad211746042caf390343c22c77c26052ccaa9831c6061185bfb8175c17b66d7149099130d0479f
zf1967a82202b18bdc576608fd80cc8c110d7f6c66028f9d437871f174437f23be6e69b6549549d
zcb422b159fee86171c409c54c49d4e2f917054a6321c311f500f1b7e1a2e39fa6a4d38e75cb8b9
z8fad731d9e0b335df35e2b45dbb49abefaae8ede833b7ce0bb2c98ccd9269b6d29325892586368
z6e38460fd95807d6f03806b898dfde5d7a7d1cdbc875a1d58545b73963120738edf3cc8eba0096
z700965282b362920e401c60a5e98523b4a792ddce15720cf69932af99563f3a25ea2539a260022
z0d81c3c4a99a29f29ae6d4c4834df71a448ca58d8b72287235dfc5aca17dfd3e58c9afe2785c53
zb66f4819c1994b8ec00493f02d57ab0bd9404ab058dbf77f5189b51a22da6646baced51bb9813d
z037749e714daa9f75ef3f5e9705fd01c85541b9357012e5f67b3493a52c5c6a6c977313ee5b5d8
z0dadf54008de6790623c2e85fbdeddf5e3734feb17ddf3bea337cb4a85c39849b401ff9dd965b9
z07f7d81fe04594fa149f1b6e6f0f236ecdccc853aaa88b6223796d30dfd7248a318641b6c19f85
z3f93a301f9efe9c1f16bb2da72954592f3e02d3b37fcd9b1c4f2162dda362999db7592b880ffad
z9668c658ded38082cbeeae0c64fda3a2569d5dbb6e81c637519877c5e26f04d123e73c4e09fb8d
z6e8f79cd9f409a2e5610c2a94030628b789a123bdccfc1c5577013fd004e5b13eca43a332f6ddc
z682ff33d48e9acacbc1621b16ae3d5cb1aeb433cfdcf6c457836597eb62d49354d0fe763a86578
z093dbe2f2e36adb0dae81047e1f79a036539bd3af9dd4bfc0db8d2193c29b55d6db6ee6e056327
z82f0ce29637d84d3f72136703dfaacf51040f17e31a5115389ec4e25b0a5bb916a379f4eaa2994
z24a47e66f94155e970d5d5c9b84eda53cebeb1bb6c1ec9f2d683e17843ea99baa438580566a49a
zec1188bea55d557b6759c3bb811186d688619896287b4331f4f151a0f5cb9439acf84b4e57fef9
zc51047b172593e5bfcf019c1b609e2e1a9f30eff4df6b0d804b34d8687cb1248f5bb3d290adb92
z6ffe88650969e24feb6a7f58bee42472aadc961b81aa547e1698e640e08db8c4b5affbefd27ee3
z74beed6e7804f2dfdfb3cacb5921491c13688f1695be2a948fb2975e19bbe40b85328e287dc86f
zea667eb12b975c050c8b549e555aee38afd5f1066cd8d7e8f6bfcd9208f36c47984654e23d616c
z0ffb89dfca9bc23acbd597674ed78e8d8da0f80e252369ce2985377ecc8ed0c8d724f00f122e95
ze66484686bc1f826bffc2b55807d85373fa2d0d80182466e5be3a113d3e8793a822d485e633bc0
z01095966695db552e6689b3b8a18372272d6ab2bcbaaf2c8d18221222fd42036c4e23390514bcf
z13a1ffa05922bb92905f9f891550ff91185383fcd680452bc677d691fa779c1a8d37570518bf5d
zb0646315bba11b46dcad254018b7551a1f117c1851887de2dc0079680ab45aaa14b580cb478921
zdda660c5bca590653f8cbfb8ab07f5654dfd8f89654799e8efa988174197c390fe181ae002caf2
zfbf3ef2709ce617730a70fb07771d92055a71c255ce1b2066bd22c0b8d1832a52705631154cd1b
z4da76294613117333674fe23e048964a50ccd26857cfbe22c5c93429723214fed92b7a3c4d57aa
z93e8e0d6acbe3c0193b0ba491c57327f113b1009cb430519f56db5b37a04d069816c92c122a5d8
za6df0958498cc4a945ffed6ea68e2490628e16d0f94b8f49e978b989225785f216288cea8101e5
z63933882e54db8e6052c9a3c4e696799daeb853acea0069ffd8ca2b1abdfc715716b6d539bd7b2
z2d96d43c8ef3b507bb4b3ea714510621565a6afae7a5e0590dc180e4bea6d4d57c668d0627db6a
z91abed79bb80be1ffb9680acb2a2945cee5a07278dfbe8e6fa065c6da7cfa4af6b8e11244bf50b
z2ae58e12e3d31659466d3554270b3bb5b5cfdf243fbe7522a6ec18bec8dac6e5699c20d1c65c4d
z7b15b2a8bdf82b1fac80724fc90b8e739999b301f530e857ad66ee76603880443c02cd31d577d7
z739722155957c98434fff9323718ef0c83cb705a5d2abdece3879c214965ea88dbfa50a1f95294
zb3363148ae94544b5b514a4e51a4fbc979ae3382c05049959386ed63062083aa91c9d2edf1b24f
zacd49fc32e0848cada010305b01fd699fdd4bb8b579b6ebd92ef0cc0a5d724f50df9ccd79b54e0
z5eca63babcc98293d5daef6e6d229dd8aa7c70be7470fc480ed5e9e5ad69ec2d13c7f1a38d552d
zd81490df245aa7381150a74570c5a0b9ce88da66f5d0e8069bbf02d2cef6b5700b96782ae56fcf
zcb70d99a952adeaa7f04a6fefe120432bfb2d84f4d73ae6f20daa2da2f1ddc1a59fcb62eb468b4
z709c1abae4ba1f4cc88a0518ee0b7781cf80afc75c52f54bb044c84982fa3d647bb5947446564e
z5df6150de1089468312c7ea4c83dfe4c7733465df791c6907c74bb394358468f4f7167412133e6
z857494aa34cc6c820777de7143458c6b8b7eaff39e797e9e55ec6ff827464659476d3e8e711935
zb332ce6cab94d3709271662fa085f095828b468381a72f9e8bff5669641c4c5981217959ef79a6
zbbd4779a01c7287ce26805e6d39237c74e9cf650e07fc23e93c889d38d464f55eac55d0abf383e
zca80b1da2ec5e876a7d85edd65bc68d76d68c73e8f16a4890c2d95ae92dbdc011189ac7a4f6259
z45b86c5c9e80e73481ce683252f48e9b437111b58c60e40ffd7f5e970ce3c6275d31ef040b911c
z84f1a81b2771d23e18f7f60fa5f6d8d62332b73ddfde31ed81674f56c19f3f31b354e06febf5a1
zfd86d004f9d96498954190e15aba50d2865f1bd937bea81428f54d266554794a4e586bd0b5dac0
zf480b8758dd0b35f03daf2e4e0801c38aa0c4cd8ad71b95976b3625648989a6c4cc28e16283d70
z67e2df0656a5cf5e0c39992db14e161afc89ad385057baa713aa92aa6f9be6217501b3f72a2c9d
z9ea4737021d38b5b3b94afce2aa8ccaa919b5ea48fb1316baa56ff3ff4bb8071dc0a89e17b0d2a
zbbd14233402ff137083db88a72f913e70a1af0f7b6db53e820208ff21833cef1f648aa875d18ef
zf83258792798489bde4dd3aea168ce20bd58ad9cafb06b03b0488bbdf2c8a32fdb1978a454c1de
z944d5312cb0e66509e56641e8506f10dedf7869bb8298af886ebc16e5ae3c096597b8cd4c9866b
z96bb98d98e2feebcfb12f5539d1ebcd492431dab6d480428b1456521db8f8541574cb7fc485c54
zbe4c3f34e6deb18fa90e9741dc4d10b8f410d16b955d6223d58569826ad2f2021a3cdcd2166e37
z263287b27d5ee485ff310deef9e3fbccd92e0aa30bb4ec8632cf3776c16e71bb4ff8ccf0458efa
z6de432aa4e3b54e305ea3c1be505562f8e591d439087c5f549068c30caa011a505d116b8047b4f
z89cc189ab908bd8b5a9de1fab8ebff004b21680023c96f9fbdc60deff399d4c89009dc9f399617
zb35dd33a97fcaa9be3ad5fc33384fa3ced8fa40be1702f8f2fc952b82a93d7cc6620c904fe5f0c
z1c7d7bdc1048c16439682bc7adae4ff1a652cd7b939b7308316a87cbaf4d7bc3c0798ca423af86
ze584fc43db0b18a23a0a332cd8ce84304ecca7c0c92639f5c15688e7d436a0b26760e4b3d23f1c
zf1a4515e1eba367e32096da8ab6f503117bee414c76520b2afa9ca8696c9ada83089885fae7196
z95e287081cef82925918d172b24fe63f3ace7963f22006e0ef563195607eaa4831d4e809695aef
z1fa6dca3b94b12532ee2908c6924a539e9151554cf8a4f82179dfb3c12a9ee981c81f3a793c5db
z2b92f1a21e54d19fe42415632b9de56ca86495e03a55c12cc08cdfa0cadc26b4d1bb09243226b9
zf4c04dc3bca70b23f4f164b1e3ba712cc04703fc81aaf1effa57983b8b6074433958baba6da58b
z8c8b5a085671b5c1012fb961425ef4debb3e2a3e16db77cb4e806da87f8bb0aaee5e8d08f0964d
zd0b2f1209b5eb061f61b8d8c961414cdcdc3673dcfe380f7a9b00ae249444ea619e06e3558b964
z70cdd965a17a48d8de919030143ddb2732228a7d4009806f155b4b7a1851404a334abfe8d2eeb5
zcbb00da69efe0197cd9b565523f745100f7c7c17fae0ea88cc92ab8bce20b737096eaa70114973
zefc84ec7fd4e428c9d8641e06c9a8eef7ee6314deb2ac722b574c6c16fb26afb139758e66056dc
ze6ed27ce88a482fd872b524256ff63545950c5d37bee2e1ae15bab91cdccf5cbb63792ec824b36
z1bdb00e5eb1f654f4b4419817cd47972c724bb34edfd942fe4a139c3ead1a2ef574ccf51c757e1
zd1be4f4808e26ab0a42673ef0c76489b13e89374ede7ef6633e5e9b8838693b195165e2d8e8578
z3f73f7eec46489a7eaa2f1c07f24556321d2fc06997fd8da4f85126b490a71e43372fcf99cc4c4
zac2cbfc72d05fd73711a27854fb5b7566dbd0a906f8ab8e8a78bd187f278ce1b4ab84d945e6c2c
z80fba794f3ecc33401842d2e756356c1bd3ff037341e13f5a0ecb0d1aa997d4a640ab8809dc4fa
zc61c9a4bc6b4207a9cbf23cd1db53620ac0d1d0425ece63d8b1d3777650d80011dc2a5e212ae40
z287033387f5a3d2cffcada86178e161145484ff4485e0aa190a5c3326f128382bc86390da1e028
z964becbdb163a1359e708e58b52957e333d28ab19401daead65b97fdb20ba1caa325af1ec22f2f
z7d9cb50dec15c665ade4c65da02a9d879d08f635ca6a921df36132bb36c681e6c525aa7df1f33e
zd9e1d15dd6add75dc13c50d233fb6e018f9846f5e4c55b039fbb7688a13d1bb08e353e1d8d1656
z46ed08290f1b583d6ed5a68b2912f707b8bedff2a37bea8e97a009b536aaa812ffff3968e1f8ee
z25cce080f1f9978aa00db267f54726cbea211097163c6af9bf419f1d83b752c3fd6bd7f9b3e914
z2d8c40f6755cf8c3bf70caabc7deb1b9c10f00f9fd558be218883b23d081fb0de9b1f12e2e8137
zb0049e481a9cf6090b03f9c5b9f3fc38c402c9911260d653278b94aa086d3d76977f7da3b55697
zf814181ac15535158bbd4ebc2478b5fdb59319c2041289d9125044d4b28b3109560e271a5b188a
z9204c3b3ba3f7b33bcc749e6f277e41aa4338398f1ca8ca19f3782121bb0e198d8555c618b4c20
z0c00d0d16c3b1f81d2b1e832ca6dc881a98ed6721ef6dd52b7f7df87c524eb8a20983e6b65cb7c
z07f65e59215185520a7538612867f202751a32fa01d5603aaaf8f06bfef14e080ec34e1afc9d8f
z92727dd3d8faa9ed50149a8c253877d21606be08dad03cb5b359fd9925648d0be0e6f5f2aba049
zaacc4ee8c53fe0e150b7d0db6150110fbf9e72c3e764a32ecd2ccff46a42174337632fa61ccf7f
z68ffa621bd4d2f874126d28eb3abee9f62fe52b2bc262d110ec23784e38ce18b9d97596877a79a
zfc858d89baa187805390a1d00e492bb6260acd4034edb947b9aa428043b8a537c4a9db94d0e4aa
z57a5c3925337a1bf951fdeee4ece0cb82623c128b4add443ec16e3f2b219ce71a144e10f5d3b08
z17ed3e7d79b2705f7b916f998525b0b9ef1422b013fa98c5d61fb9f700c7b1d903338e6ec71884
z5f93029515ef1474ec095067f10a0a9e39d4a528bbee3b8251134c8a53e872ecb0ea7ca317fc3a
z7e139020f3ebad862c90d8137a4d801ebf0d04ba6e057699c3b2d096821ae614d530009d26cdff
z7a054cf112a4f8f0a98c0beb224ffeb6c05a6f8b1e7437631b54e05964f5608ed11034a2573b09
z8202c2574286096002c47587d818ff78c19c471bc8ad225921a3978c61b9bfaa25c97ce07b30dd
z1cd4d5d251a42cb9cf96c7fc086c4f0d25c138fa6687277dc4438923280d1bcfc998e903069d50
z89eb09596584cc5534777efaebf12063cb5453c83e03feb638325e872df23cd81a85d26af3083d
za5f4297da2494b0530bfd5d287099f13a504d931b252f927c6d94dccd77cc6be9a0dabfcebd6d8
z231ff513f1946d1185edccbc072d36ad792df0ed928757e66ad3fbc2390ae8d980ba4dc713ada4
z03fe4316b8b57ebf51eec6bccf2b0cc1ae03a49f7d154f3eb90c313c12f75fd2f2017fc015ed4e
z98426dbdefaddc83bfaa5e46a39f82c439ca9d3923cba5e75c89a9375c7881369c4c0614d80e30
zb1ef74dd6a3db7087972e4475d0a0d7d6882adfa8f882be596acfbcc24a00efb91ec66b36612c5
zfd07774f24b71094b03d00b42409552382c9e3b811af2ee5dadb23f424766f035278b9b98ca4fe
za11b320777dbfd68611e457d47bfbb72231d04687ccc67eb9194ded6688e40202444f86143f303
zc7d264870ebfe1e7eb252b7ec7f56ddb641b1d4c83ff7905ff06a60aea4b9575915efcba2d23f3
z20c603e0fd8e650a92977053d8c348a549533985c979c433dbf0da92506703414ea79e61924261
zb144fe6c67b706312df462e6550988e2565b5860378a5194781a65853deda886d990c97471498b
z68a96bc7041f3bcf67c7bbd3bee5bf56b6aec29c9832971db6990ccc5bface4151eb056fe424d6
z2145ecea762f638b8b5e32d656cfe9bac210107544aa5552b9ae6b61bac5208c1ebb677f5513e6
zbcfa6565f1e7c616d8195fc2965235f6239e442990f53b3b59c045c2fbfb1dc0434186112a9c24
zdd2bab4f4e6f50b982d3d1d67829566535448acd6aaa4be7d3b854019d13bce1760d6864ebb91e
za6d1a3d383ab422230ef6927c3d0cd4170951995a50e104ca5f4490988337092a4f2933dc1d0fd
z910c29556936f86f062ac0b5e537af26d0d6140af1efd7f651157b3b4e37d46c6c4107242ee15b
z53bc2a2e10ec28ac8097cdd570f3e392cf99229a5e4fd7ea702a09b78d6a0d6e6119466c3dbbe2
z6cc768ab987d49bdd3eaa067ab6093566a8d03647bfa93bdc5f3b178186212cabff64754565203
zdf90b899dd659e99e492833ff6fc3b6edb02c6059d8772d59874cdd4e9c0a3698fb78ee6db69d2
zf3104f3728476bdfb4ec41a69db66756e71cd95b6fc6d685b689e30a193076870d04df9e65e523
za1c4eb3e57d10e6a249520e6abb2b5b97f4c2875e8f5950982262ebbbdc7dde4c9582872656dd7
zbbe9807f8342ed14743c93cab9d85006d358d005e736edea9461d67578b90d3b74d56bddd5965f
z95d3295f5e17b5e6985758db8b4755c8a802e16506634fede7b6d8a2bf9e136efa713ecc6b6be7
z63dc4eb1bb7d6f9e43c7602aa48ca19a516b07617b14f3f8f93e3f6b21b2ef1746fa18cb30a66a
z32b43c49e3c51c7b4f9a2c3f92811f4d9cfd4e72acec0b331778a8cf4f75cd52fb76521d816a13
z8aaf6ea0fffccbba28e13c5cea18fd1b96dedb8951cfe1cbb4b84057c257c19eea6448e21e9346
z857716cb026cfdeee088991c9d58a61662fbecbb0f87add63c8140623798d651864d077108be07
zeb05b651980ca3108ac39866c21f9ecf7554a40fa11f1665d982adf38975b801022c46ef0b9358
z2b6bf460a3c27c489679528d76c0836f39ac4e1ab16ea8f83127a7158f8db277ff28c74e234d62
zb52bea51c691dce9da4c5565018135886cf156b2de568d8bd92fe2b56327c2c8390defe02b9977
zb26e2605fb0d6d0084733b31ecb032fdaa504376c5496af8238d38789c80c6c0126259ddfa48f6
zade6bfc0890b47c3bec9e4bfedfe1346333140df14b1504d01bee232be087260ae5c0affc94890
zede02fd5e5fa6c78f15a69f2fbe40ea0ff1de55640f8652347cf930e5c25d943db14d7f7073a90
z8d373862bc8d46fd3882c9d3153eedac0ccc9d308705357243c56b70f0d12e036c39f775c94d24
z639c3519fe57eec67a26ab61268e7500b32eaa5ccdf6d89e72d37a0ca56383f4d3faad9db0652d
z119ddeb8f5b7337c3b5f061f8b7c0b5aec33c8a1b7a32bc2636905fd8bdfb7db3b7a29cba2b0ee
zed8b314482b89923715b1466dda8fbeb81d84dc60279db2f84635f2c9e801d2e4b605a528cf4ad
z13c777cd3da9164057a874c679d94a947253e3af2ecc2c26a9bd7b743c7d11437e938b6225907d
zcf33f4bbf769d1147557ff36ff1ecac571d4fc8154d2042416b4fdbee5e800ca670ddd2415161d
z9ba8255eb61b532540554a9686bacdf0f6afbf314355e0d98765095d535693ab8502baaebc3972
z79c693cbf3b6ab6c3d641c3d1e747a8b1ea523583179fe48479710a0c060df813059415302b985
zde41c5830b6ce4e09b5b9cda9d3e20f4015e30006ecf53f31743738a704bd49608cfef3c3b4736
z3a9c2fde1581f4349e6f87af6d587ab090018cce2d9284a2429753454946918451ecea91d7cece
zc2a2c3e81f9a56b9fe549cfec709856c7f804bd94e69cadcaa5403f39d330a88b81f1045d80bee
z507a051706508fb3a5ba95d66721f5de3c79de24c5f15be68c4ab042058079956153e7847e90f5
zfc546db8cf3f18246477865b045e39c7174a2529cb3ff731e7d9a85992930beb81cb64e4535320
z8c22f75fa0bf16b470ab5d970060e57753454ecb02a16809823be85d2ee74c7e939a959bc4b094
z4d1b734602acbddbfc30178b88196ffde3cd177ff505fb70bc54088c2356a6fc5b9aebf1a3154e
zbd648ffc95c2fc1b5aa75a3262db1f33215bb601cb98ab377dc5a5ea6d0a4218d036f3d33f69ff
zc4ee245965c40304e3cc763d51fdcc48bd3afc7f998980495417bd1ebda5b04d13d80b45f36140
zde9ffd4aaa6f2b660249bf3137de402f432a381dd6395e3641d0a692f3e03d094c1c9de5fdd7e6
z9517140e764a537e59ca81d7aaf2deb484a787a96ed67e2abb927962dfe9dc718ea33c365a8bdd
z33cf03fb08d92a7720077d05d64256bfb2c532c8dfa9a33121aa618319b1414b08f025f15301c9
zde2051410ff7feec0158055e8711692d00c716087bd87fef2447c755f574dd6bfd698614c75645
z6a04f8ccf75d342be3f338cb24eeab5d10a12fa4d0a0fb8dd939b1ffb45480e4739b258e02550a
z91eeb150d0a80509b919e72c022005698f66632ed1a5084c0396d088cda816aa52dbff3b8b2c70
z8dc4f2f19e3c32b151ca8c6e3f8afb6de874160cb2a1f165919edcce4eb4b459f097f2f400027b
z57b6b1a9c9eef5ca02d7ea2fd9c1e3aa919a9a4d56ab57f654680e4a581bf04bcbdda7c5feacf9
z984e2c55740bfc814a9c79e24e97a59f684be7565662b0a635dd5c285794acbaf302f45556067e
zf15d3d6dcc1407112fb220bfbae81a29a12326aa1b34a2a7e050c94b7ca412f5e7f67ad44fb9fc
z6888df02dee2c8120f5aeaa245a613ea7c8182fa46e2120f306e8b6d6e24a88454d464efcb0688
zcdbf0b5e3bd8edf9e087d9159373214643c78eeab8f7301a81bd6a2d6ad4132c23397aa3df710c
z1183313cdf4253851f92cc6e40f83338c9dc7b80bc6e76e64abcd40193997392616bae3aebf1b1
z51313f52fc1ec3eeadf995ea4ab82588de82559540c358e49cadfc42db26fb48a89a7e96f93705
z9bab94b49377e2c359031667f63043a7abce9e20c49a73913da779e6ed46b66ead8d9b40678894
z492999ef1397379387f217ac9d8cbab8456fd2074ce3b2ec1547df63c7e5a6cd39f2225a66ecb4
zee18dee456370a32cbc1911e4530e2cf90667b7cf067d4c8379cf3a299257113f7eeb5c31a1047
z907b677b5f7daece984fb81b775f779d7546862da240e240a5bb5ea81d51a17aae4ad5bc43c115
z939081fed97fde4ddadc9a2af7083f7537625635e946d5c9528361c2c1d4ff5150dc5687810c2a
z071aa1568bd83de62f06a5efde0fdd161edfd397aa0d3e5407599cedcc160c9a621b42bc895878
z0706c121879981067fc50f3ed5ffcb3ec56c4757d38abcbb88a0b1ed500fb5586710d2827c93b6
z4243292a9c027f8ee7bb2f5fcf2894a8413534ffbc0b00bb511e3a94d6c0308607af88fef6f770
z2dd46f5138915409dc8959c9eec5a6e603823800bcd0461cc89e6090f9eb362ddc98caaee86a14
z2ee91f1320174d2246255c2227e074772aa8dfa9888c493f76d17c24f7dae0948ebf2415dbb8b6
z283dbfa64a0d3785fed575fb502bfea7a2faee64f422e5e580377038d24f1bd074d85b3040378c
z5a4b549a26a22d82852375f907b30333259da738aff47f483a885b8cc2a392d7c77724f3db8e98
zb3620178abcde18c86b2322701088797bfe1242b619d4cf82528214d5fde9eee4fd81209649daf
z4e4483b09722caf423b5a14e7a6f2136ca9d60b22d20f946d8c3832f45b0197d80c9d8038ea90b
zd3628c396ea9c2dcf7cbdea10dc2acf49d7137b2981dcfb269f9e502044421995044ee8536c1ae
z834fd6d6e05b0a404a197b442c01384605d59d7ab1506c301835c929a0e190d3860798e0258f8c
z5d74c0bc202b9b0504b5438556855f0880316bd01eaabb21bfa0bf140bc14ecf3b101140fe95df
z98de9aadc164e1024b6660bafa1d19f77872bd8c9cf9dbe83c41fd3c71451b3d7463d62e24dfa1
zcbb30dc4b0ee344f0de88707ec1fe6cbb7c6c6aa3a22e3e9d46423c5d99876df5944449a20946d
z8fa8c2028471ea022dd53b66314d5d2fc2db73c240f5aedc89c9bbe24ef71f064e52f82ff026d4
z2957f64a2954f9ab40afcc005fab21da865fb82e784bbcfa25582a9ab0f24109f546532d878f2e
z2f6d7bbff61fccd3b6e91b3acb2e0b68d6fd18ed754c2452ea6f9c7fdbe424e0379171a1ac6162
z86955dfb063d84cb272d44716c9b5a97590152c48b3aaf37a110b11171bfcac052a3a8f4dbb12e
z52539a7112a177353db5dc63b09b7a79142bd3128e8cffe4adfb72f8073add7d42fa5f1039cc36
z8c344971f55140b9012628631dd337e03f8e059540d00932c93f003486a75332ac1ac84233d86a
z935a51d4277dde1cb4ef046e06bc011deb49d8e66616a098f6a1a764249bdeb2c968026792ab9c
zc2bd232f09301811cb04458ceb1fc4cf225f69d46ef06d2ad8bd8d8163e8ac42b7ecf665df42f3
zd5a9fce32430048bfccf6438181e4c25a3f80923c0f113338295da05cc2f5c6dfdcd15376a4382
ze855c3507ccea9af005997622d39c1a5d8434f3c4fc078796d9388a92c5c6d6eccb0c180554724
z6bce00a7bdf9a38a0b4ee1cde9057aa9a4f6c20cf6798bc41c87a702ef61fc5ba3f3887d4516bd
zb948585a0a4a741076d35c54edc39f90b0b8384b0060fe5c5bb43def95c5afd799ca5fb56042db
z85160676386dbef07889ebd4ec6323e410f027e50480cfe796fb090d4be72146c4ef31d29f76ef
zd7e54b75beefeef53f91192080e2b79d8451c358543777d7f0c1abe8117d7ce7bde762f8bedfab
z7ec24f7652b9de51f1aa55f910e4824aa0d4b528cdf0b9e18bdae1ff45fea892092aaaaf157c8d
zc822963cb51ba443a6b0a845251df0fe58a5762ab39004e56a81e74184207fe2e38baa9d7abc69
z8b8c5df4dab23db74a3421504d3f8457c4b44cfb97e807fa8bf855e4021a0f5eeeb20705dbfd05
z78d481eb1284689ab3e0e2394668825fe561ea0510d65520df94cc1349562619807c90cd0d6613
z7335fbef343c629820d4ae35920381e9d89878748d6d0939f955b1d87cf1fc815066f7ade25435
z893c3ad87ea61d0268a4ef38794e3540a62059c5bccaf6892057cc4a9bac130b784866a129bfd6
zc9410d41fbb60317f09869abe2e4aa54364b47e16ad4eb21d2a85353059dff68536f49e74650ad
zdfced662cac7069d74874554d543539cc523f2c97c5efcdd803a229aa7f4c47b4d5adeea2d5fd6
z674e1017faf3352af4fde051bf7cea15d39f32380db0fa0f51971d2943374fe44dd92ee3d4e3a6
zaa0302b604cd97f542db5d6775001563c546ce2f2a003ff3208531b531e0791e4f5b09c111d101
za0841be0815586d5a21831ece80d4f64df03bbb27e7439e784684b0dcbe8087372fa4af40c2a88
ze49c234a30889b7e0c99a038c67eb36186506b9974f12e63437e5cc92ba8558d0c66e43067cebb
z748cd28a586e11f20128111c2ff4cb669c53e073e5f1ddfda6baa2c025560c7393c4d62583ca2e
z8b5a8cf3934aa303ac00265342f4df3fdba5155fd1da277fca57f918c500daa502c1789bd6e1dd
zed2078693ea93b6c2548df5e87fec2837275b2d73c84671b9c6238e81f1a0431434461e5026c90
z93d65fa3d704a505e2cbfb7aa388ecde118c5d1e938b410d43ff068366aa974cb8e33a7afbdf9a
zb85afe93b0a488088e34bebbfebea35d359440f53a40b3308c89c7e301d0264cbb5723687a604b
z211915826e12a9ab73f4494278b02860b2df0cef59ebc586f490af183167fa0c1bc2418e294461
zce26919f67728cdb20446d3d3352381a8b380ff6fd4bcb10cad84147247eb18396620ec71876f5
z7218c76fdbde614ba21050de931698df08434b6636726ddf748b87ca6323346c47fc5511d18e63
z3d4dfc022a7183e839ef9c0bec476904ede9d077fe233e72b8f0497ef9b11c413673c499863889
zc2dda02a98bc11d2f11a47e07377510e76fa9a30c2b2c6614605e5a2edc5d47b789d311c2c9281
zf26df86f3f21fbd8174b657824cf6fd9f9f5d827b7456553dd3f919fd26030f74970ef926680c7
zb3d038f0c97f32c63a753beed4d0b051d0462c846831c4db1fcea7ec721ae632dd9508ebc03097
z33f42e1a60618a9e284533b61de654e7de9870073e56b4a35ae2e5c233ffee984fb9c37ae45bd2
z3feca75917ee07cc53c4933b5a3d793dbba7eb18c5d990ab7d0677ec5dea81113027b5913d7c0b
z14b81f776a6d8523314d8635e6d6734cb1cb91aadf27f10dfaccce09dec5045ccf0a49b67b58ce
z48d735fe98e7ae142caedb7857c1103d28c532e54227a35b566df6e13773992c4cc1256d7c0f5a
z6ea6de914b272e8b4f786f4b22dc0314963dc66b3d021aa665c4bb19c0609b25061bf5171be3b0
ze37076c34fa74c0bf42f4912a14a4e1ad5f5f7d6f8acc16a3f7bf3e252759de6c84bfdd5d24146
zaeab10ed21075fd87f493bde50c6c01536566f07c453dd2544d9f2fa1bd4c63c6e9d887cd3e91f
z0bff01ca51df7406679bcbfebd1995043f236843732e26ea96d55cbb5f76d42a47a5664476454e
za5a2a4280a6a15a66b0bcdc1572ebc1664ca0c482aa102939245edee16531e1635d71b96b27d5e
z919ac5e8256b867dbc17a8c16f5c27c3eb291b24762b3d1ebb9d719de719624e251484f226a8ea
z4495eb00de7a4191a6cd12fc12cbb64d7f4f5b48239b8ccf6b3120e9b8c2d5934267f92ef1a00d
z7218ebafdc33ec131b505fab6fbd90943aeb96f580730537b28452bbddf078811d92a6e9d03991
z4b0573b53584972c5afa1471bc3dbd623f5c0284a34e8c8b55b978dca66ecd588294a1eb964821
z36872e9db49c9b778dcb0615632fa08b874a43ff5b3562ce8f727cef43837bef5d4065ac7faf08
z18856381f5c8d8bc85bac506e1d4de5600061e646d27ed7d2ff283c4745d5642fcb21e981fac9f
z7b2393fceb5c0cb4444b893eb8a78edbc0cea6c0d7aeb0da6cc86f631a749d360af36e653a86bb
zc9e3c3ba5c7721363a155fc4f82e7cfd439a67b4b759631be85c3156fab9844408f3b332a72991
zddb37e6aaf57e50fe6503dc4b689cfde78ca5c1cb5bf3b98646bfd9c9f00feb45d5bbefb6e35d2
z01a883c467601d76dd24f02624589cfa8032f9112f4ce24d412908c82516d7bdac1a857ba41a9f
zb6171b504151bfed09e2a4073aa575ca32edd2f612a2c097456bbee248cc6018f3618a17bee90f
z46c1f6a9885a522d2c83cba66c6a439bf28969d8dc18ab4468d4e19a09bdcc3bfc41db90343db5
z1293c86869d00036d8a066db40dc81e3b2a8ea64bd03db159dd5bb1db5e162189c829cabcfcc96
z947e6b48c1d1ae4b3f06f3cf5b79afeb7f69e9d0e81ef5a7eefbd82acc92749cbdc745a119871c
zfe063ec8fedf13e75824439f84aa65ac2d3194a0f4a5dd33a4e56acfce6c545a91e85b56b0e268
z5463a0177d4eda9148f279d26b75cf96a94a5e1ac40792e28c815cff6e6993bbe9e2f5fd46aa40
z5cfb3313075961b6958d5ff544188d0cf3ee4e0e955f5a677a39111e91b5160ae7583a1d5ee19f
z65f79f208fb86b7e9439eb454ad26422ddb302fecf3e953275d55f14fbf53a4ebb0cc0c1fcd643
z05866a0c6db877f5aae1d4ba9febbbc4cf176185081981dd57af55b5e9514d49c2f082815ea395
zd51c1f5815956e9bd4f8d9ae782132e289c84533a7e0c6f37aa9170abeab76435f70fe885eaf95
z9218246a237c4e185e8fe2fb7b7284e25d4de2390a6c94c967866108fc2a25982aac481500c311
z81bfbb817128005416c7b7d7e0b77bcb499d810c11e5fd8c9f3f19091f43400552196eb2ba3192
zdd2d620b0f04694ab80df9f68a41abc136f15cf0d92abb7e94153c3784998f7fc7318122e34365
z80dd764353ccf3d26a7c523faeacd094c3aeda2a0bbeb11259927a9463d69e679cda3857b6469b
z3b65a17522fd08463a467abcda35337c9085a9894133c9d3652b3c0e1df75d0955400ab52050d7
zdb3ff6edb8fbbe94a51573eb90351a96164c5618260588d9c288f456b4626a577bb9061058f7f0
z1d373fd26739e32e774f3fd13aa404107abef5a9482ff4d9ca34ff3f0f26c0d81d9fddd0ca6fc5
z0f052c26bd18b083a11dbdb2492f8f1b39e5ad45cf30c670e5eb4a0e2ff499a69f40848664fc33
zb720d21390b618b2faa0deb3f7ec6ffae58f96d72929bf05438d7992fc1e27b98a3e8c1a824620
zf6bac41a5039a5c8a95b7dd63a393ffd65adff63d3d192dab0b8bdcc5a0e974b3d06f899aadd76
z682e44ae83484325e69503732de6734d686bd33eb33d24ea6cf9d926d5e2f9a31a360c47d172b1
z223af6f31b4183251032e13116b8a314e2cfe2b4563afe45ab403cafefec4b636a6706f1f1c0e9
z723514dd49e02196d744b5c96e79706a7d99e66f54dedca767ae167f466ea1eebe2fe985ccba03
zaf95c393323d121d577c42745e5307925d07a312550648d2f4343997f9caaccb2b96172b2650e0
z0b39035aa67f4ee93c950ed12c9d21c2eeab2c862da222ee0296bbc03c78e9fc5610a0653438d6
ze906acbc5e1f525b702943a6050af6a0a72d44fb5e02ab2397cc3e2f2408dc3d3d2d290394b8b6
z4f678994e4a8b32f1e14387c3efd59ef16a0be53cac10854df8fc36014859854e04a5ab1924ef0
z5932711be6f87a7117165491a18ab74fbecb9fb2bf6d1bb5c5f335807a079aadee47f443ab2b0d
z6877da03cd02028680b19054a8f296e80c114aa2b58cc4bd60c037d38f815c19ce4cf8244c35cf
zf194b6a0819b340ef9e326f1ef4e215a5311c3b8505780b2bfc6352b2db8c47183f328a991c515
z50770ea24726b98d5031eea92e31f151c56ff52233af645787444009204da9ea58fa545520ebf6
z0fd8cc4a35882280c1de931d655ddedd606c3ba42652c4343e1d1c72a03621bc141d1522d2f5b6
z6b29ff3e16319f4e9559707cf2c2854648dedfaf9ee28b5959cbb59d40ecc0aab73befde613f53
z9f34d83c014fa0a4354a71075dfc90353948be3382097a4a1b83039db1bacbde262bb5c3513dcc
z98785fb7c5fc7563d1d97d1a56ed14684005fa307195958ccb2f5884b0070b85b435b5a56be8cd
z8d1423b8cf54604f8457d84ff1585b72aaf4ff2330dbec16dca5db95677350302a8782fafccb87
z2e58405613f37a57bf65d23f68ef83aafa348e2c7d5786403ba45b93888ae08c177fe1f859fdb2
z61a7ab8e80249d84da7ea6346b5d7bf202a5377121c75340ecfff72ca6c0b14ed61075ae5ebd93
zee367cc6c22eab1fc4545bcdb3035afec90924634e107bbaa7e4419b7d22f50c859b934fcdfc80
z611a37f9e5942c64007ad1100e181f158827739cad860817bb1038a26b98311ebcdcc0b04dc9f6
z406606cf6dec3fbea7728afa80057e723bf2ca0170eb979b6bf14f1b00df61dc87f593ab28c392
z76fb9d6e448368a6083e66a31b4a6e3233bde75ed1d9e3161d9b50c59c1aedda019d445b48282b
z4092f9f44ced400b072eaf6d410994f137560327b66e3ae3a1711d8621a537b6e19f65fd01d220
z1ce78aaba09fb78e2a786ce23cfc62736a3052820a6dd71eb4884abd41386635ff6938bfbce7c6
z2cb6d29f31386ec84ae6538e55e91e906710b814d87ca22c753bcf64639728ad8622aef227a582
z417907ad4c18d0fd4d184b9682aaca6fdc5529d4114904c5a20d070fd6969c3110b67fa61787bd
z4cfdeaf52fb67bdd00dbcbae125ac5d101e992ae1297e175f0c2210e1c7f31a781407fb98d3863
z3199f1a2f197ad2dcad9b7c7b752912634546d60054ff8e7d4a836dcea9837e3ee59698d54d994
z95cc629e1a215f436e4bac661bebdf43b19701df8a5bcc6fbbbb13e8018cb8e6cb98ca582dcec3
zb05a5b8d48312d0a2b544e6d34c4ff89f343b44b52d436f0edef305ee61081bf78d69ce5477822
zad1d3c085cfbc591fb5b47b55a005ab9402a75adda07a96cf89c78264eae855a1adf623d334675
z63255c81db5a32fbccda0eb3699b1f2229f9952ecac74640a6e8c3e1ab82f29d22242d092bd060
zc375836471554ec8554f512b9fe655facac236b227641678d626b7e18ed427d17f11b7df992db9
z29589aeb3d2248094242ec0ccf0415bb4b5f4837bf5fda82058a4fa5466e234806d6f49c10cf59
z5a49dc59c22cb5dc0bca61ac642462fd7ade61836891fd23f37b1b77b7f22ac692eed599364e3f
ze654512653f8f64067bd7d42520f9a00dacff21db6f9dbecb9aabdaa44ea0a4bff897b641d610d
z1c042bab7238ed2a75f9f8191ef88d2f501da9cd315152a982b9d800866fce599269f5ec1b0b34
z788269e9eb526dfd0a1f39ed8a96ae8915ec90e744a54760fb150a2c5c7bb0c0c665244f77d887
zf426252fde72143b650acc52984e82f75d4c8f6eda0f33b2a452b2cba150cc10cabda88f403296
za0055dc0e8c0cb33f4cd9179a285afc789b43d808eb40b4d8b473a82c17b38f3d4c3f25659ebe0
z5a2e6e7beb595fb93549e1e2649d8b2bda22b7e2872ce681bc66396680da5a5e57f0467874fdee
z96c6b3c707d63557e796ee404e5955ebcca80c15db3482ad46d2ca4d8484d25bf85cd3ae4f48a2
z19cb97a170eda8e646299d8f025e4f3d4935c4c7d1c26765e887ebf02701d99dd2142c9f0372fb
z9dbb27691b50ad75e52b82f2c2e293adc3b47dfb5523b34ac3f1025d65eafadaad0f0f81fb4501
z66d9ab9e1c4190e091bb61bc476eddb3364f41a2210ea6244f8e1ab78d43a078bbd5d7935fa428
z860504463900e64ddfede5eb9ea3dca248a0374e50372f547a3e41b2240fa452b65aee10c635bd
z2a3cecb31c198b73472c8e686665539c60e01a54a8408fc1d46b11f2ee7a385cfa31419bab7a78
z5c8ef3f52a4662fb1ff8c46649c13c589da17c0cfa0cebf7695d5e2ab303b7abc2ff6352ce0558
z354092f6b831a2eeb658ee9170f085df898e2e60141887334f60378c8df6d8213e82d75ff2b27c
z7edd08dc4c9046fa9f8015633266d252a098176a5192988239a5a43146e7da574f6038f82caf52
z61d7ba797172ef7fda24bf150916ae3b9ce1b5a4dddf50ff80888a2d99ae502b158c6933218065
z7d23c528fa4ea1f675b0f3040145353b8094ad0a85db7655b5204aa122307cc5f2c216d6831bdd
z4a5f7e4b49cc537f4544cdfd89b1df99a708b96171a0cacf87254b3adae45ae757dc593b596f5e
z23f8e3ef0c83bcda47d27549482fc2c5128676e6f3a97e7bafa0c8d8c46685e44b35aa68b98e3f
zf3267edec2bb6dfa5c789885ca62144d16533e014a2cadeb0db10ced0e2b5b62a8d3e6258c9daa
z8f0e708a0da01fae37b8b21de77b7ce1e2830ddca9d8b6621eed14a96dfae767c7378398ce26a4
z399a95deba30b90d36ac0cc0ae39085257d2eaa954d14daebf973d6efe8793c28bdf538d8d0886
z3b82d831d9930c750cc3cabf533403a38708826f8122fbaa763b0c8937c8d324f6641041cecae3
z63f4d9bf534e24120bbcb9081b4627bef985b459ee6dd1683513d203c9fd5381c82a29e52bcf8f
z5d2a7b03bea7f4f490a19274b1da5676ed4e172c144b69f68a1d464b0cb992dfe3020d0b6f54d2
zc72928fa2dc8dced973b8bb3306afa9cf14919d62093e328c36a0a5b4a49f9d193c09dd97a84f6
za35a41b4c75b5350f3f607319ba3ce89eb7e680d9b150196ff450b31fa3195254da87cf0c54a80
z85a3643824adbdbd5a65100128b155a4598b232971e32d9d33adc56c6f2429ea461e47b9cbc756
z133e5d426c7a74da067a7f9f815197844573c1b6a421ab68de587a19eb8e9b603e86706fc51ca1
ze4b2750f9ab9ee772276e36139575080cf96f14b8502c3885db25e5f12bab94f4cf2cfc106cf47
za5abe5245690a5029b2c4cbec0d3d8410183ddc4096021aba60ea4af5e64afbab5d8358c1bd5a1
z2647f90dfb36670221b16cc3e30fb33738ad9cbe664004dec7c36b9efe2439eea0eb32525b4e9d
z2cbd7bc132ff17f2ae2e60e8854df4e2751f53357899c94a4ce4c5decbec96e37870b1006a4cd8
z4b2c71bfd3227cc9fa95b1096d801dbb005e3c43af4ea52fadcbca5bbd6de48f85c5cff345c7df
z5059bd392c9b0a7fe4ee0ca7feeacef0e284a5f079701d6b50a4c328dddca5e460142746bced23
z37d856ae72fdca5f3afb7911273cdf00658c736d76a872f793c927747048d6869b3153bcaa22b2
zc40773637441991ab29a5beebdce2310711d0126186733d0cf237a1756785739ac0bb308c6c738
z80e1952b264a67f07500d2ef12a974cd7a75fda5d997fb38ce7591e1ba492429cfedd8f3a12219
z5dbb2a434f61398493f1c4a135c6bf1dfccf78b65dd9bb71ae8ba8e782d0407804e6ad406c15c4
z8abe8a8ccbb8ce40068a09d94aec80c2fe5b704efe791a665e634aaa2e1f22a5a3b91b2cff56f5
za1ab30c2d4af21d26e4d84e5b1baaf59d37607e30269700a1354e5bdfc714ebd9847d0bb5fbb00
z3b2eeb0b471a04618d6d22232d7ca64f508d4168b85256e34eb11f3df973328ea8c58f29e727a9
z80721562f313ff5fb8a77b56ca65089a3afd6f38c1f289152bfca21f85ac1a30a807b91e6689b8
z3e4667d2e2da49c6f842a4396155490bda4a9f2fcc295406827d5cdb401900642d3a0b2f556a14
z87a989fb69dab440d873fd2038d6ec4b20ab6ebd743d1a85a860aa69639fbfef4576bed33429c5
z3e85796b14c474af335f9ed9ba5795f6483aa642c30a5dca4bfbac9b06a44fd9f1f9e19e85fcfb
z69cb14c792b8da4968a18ccf45d8d1cfb8bef5964a65a51636eb75cb09167c7423bf2bccb7c30a
zd319ff9f02a15ab263b5fd8d119447cadce6bd0c3cb4bff6cedcefb8a0eaa726c29e4b25bcd95e
z06a76e9ffb355d64c23483e6dfcf42bc14fd7c8ec3d03bb6bc5702556999797e64f25a60c39c25
z9b60157ef072859352f17a3f244a9e08eae820828c1ef8e46d126c0aec1aa546f3786a8c632369
zce55b2e8be2284f82e8a6d48ea143d413ae41afbc45864d87abcfffd03eb5793838155765fc7dd
z7b5c846cf23cdfa7d834474d7ff723e81e140fd0b4998086503f3fac79407afb69370147aa4182
zc845c65695d0ab6d76f61c1b1e74ca460a26afdf262aafa56a85e3832eb3b451eb892ebe0fee98
z7db739919c4442a6743df7686583ac8641bdeb0f81ccf11bb2f01db0ce36f580a65f2150c6a246
z030efcb8eed0e58ae8717548b205eaa318b19dfa5cb5c19fe14ceb42fdb0286e5849aabddf0d87
zeae6b5bbf6a3b65116d26e02535de55fde3e4146fe2cf8369b92a10764eebf15eb5811ac555320
z3f861edefac1fe5d21d813ddee26a6a21af2abec070f655d5de280032e3350bea2f68d493b42a3
z6f4d9ec78f170a0e7cbe9d367264058c8bd30261583582d720d52c6592ce6591f6714ae9b8ba3a
zcc8436c7d4445f4ab535240c68e15dbc5121ed97a79363eea70a47f8d5e1597438ac91fc1d7f96
zada6307a3f245a42d9e72006f1089a2d79fb869f80ef5973e1a6b4646942cdfc1058c66a72cfe1
z45dc2c64d88d2ddd5c94704680882b3ce85801568483b4d86e53ae54a3e391756a60f4dccc423a
z6661b9def10bb4b170681b01a39f70c71d87b9253b230ae6f3a750707b775fa4ee30d2ad8b90c0
zbbc3569d9c3084d108f67a325ee40f9f02764cdc98db417563a1f8f75ccc931d1541d14cb247ee
zfb925eaaa42950c419fcb89870a14a21a41c5626061dd8540d2e274c5c6958fa037ca788a4a1b5
ze4c74744c0edbea8a6b2dc013683dd07d0cf9519e6009b32e1ba96f7c278dc8cf60c42e78d3c3f
z34fbc81842f8f3f11c87b50d3370a677872d05b4c542633f662b3695532e2e397b8d830d234ab0
ze187570002ed8790799e6054f8f61d6b770df5eb8dc65228f9841fc71777a8fc37409e79bc8cb4
z838d174658faed1bf37c4cc2b44c91e13f0eca99d9b8419660c89195816fd625cfe13117b3a1b7
z7f9dc27f4bd9367f0dafb7a62bce6600165705da089b8ff004569f1989fc92c3f53c34dc118a65
z0026310ec8d35624460612033acb4f91aa0c7a04270b11ddeaecee8d50deb1f03a9924dfed5e28
z9890dae17cfdd037f9cb49e4718a744b2ebd9e91520fee79448cc941bb543324bd065733bbb224
z999344bb540980fbea508d7e7b5c50813d428491093d07feded5dfdd9dbf7aeb8d7d77cf28cce0
zf146c7010a3bb5ea7625a98cf366c9413f519c5ec6fda849ee1065e10a301941f84c63cc877056
zfbd304184846aa8e50115e9386594a70c6001787f4fbd588dce8811d619a5cbf2ddee903c851c1
z1f76ccd78b612fd4fc0088ded1847123c60e36f562306777dad947a3573a0734228d066da17de2
zeb52a321106ffee19207f60ba53235068e0f92d62c13144b85afa527145dba88d7213fabf5fa5c
z979982b7a91950c58eead469ce926702f2abbfd04a40bd48109bafa6c9d105ebf23759f42d8040
z822744fc2d6379aa9d226499912436b759743a91557acda91ccfcdb86a12eb8521734e6856214d
z17abc1d9618f76c3415a84130fd88e3ea4c15d20f3b5579defedcdff398315aea07220d8e4572d
z40ad0fb241e4a44af04f1091f60072d6302decc89f28c388744009f0ed0ab573a1972d2070590d
z7032b45eb122e3c352906543919d16a327d45d779dc90509dd6d79bbe678c5e5993d90ba179071
za96ffbe41b6e17001fae753e28b393e1a39b4eea715ded0cbd88337688b230cc68874fa783480d
zcd0e7ba6c282ba2ff7c65a9dc295667b6ece7eebe347a233865672ad550b9809482c5e931f1f12
z52e9b451aee49e80e9f5932cbbd46f05a68460e7b9bbac928356d30a139f8567edcfbf17dfdf36
za6047d5a904b46441597d4d9ab533d41db9fd2b384cfd438d75782fe02ed41e599973c08e98e1c
zff24308b86a272ce41173f4c081e1ea2ffa012b61d73583172d8438125016753f7663d7c4cd138
z4ee6ce9ff412f7a33cee8f06e5e7167a51e6599d2345ade0b0adbb69b8f8e2d4cd4f5f83737e68
z8ea4f9600d2231d19c91b4bb00b7f8454881bac11162177ad7492f5311224c8726d9d056fc6316
z2afb077db986d61a8298a0f34049bcb4d9e7bfb233b33e5c8a74f2eb6dd868d226f76e516a48ca
z81f5b31fcc1648a73ac1f5697c560fd7988a7a8daf4888c9e416e5da9f475c6e1324fb50138a0e
z2e4cf10116f2359cf7b6dfedc7f167ab847b17eddd15c081132003f8bcf28e97f70a1185fee0b0
zba10547cc826baa9d5e628385655856bb4344bee5b968f74667d102cdb0c72e8565370a4084cff
z30eef19f47beb93e812890fcafc8d2acb323cd5a7a8da4823e769c07276644caad7fa532414d04
z393deb4dd6c3630b0b7e4414fa90171db94a6d9a973389c7e4be7229cfbfab0e34a5fd6431acf7
z4a62b6fc51b3e2287e31f70ff11fd3617e46b8fa7b58817959d53e741cb3cf93f5ce2bad2c0f75
z8d298e6c14fdaf9c8c3fbe20afb229d9b84800cf5168960131852cf8f8b33eb1f026be9243cf3f
z7a9776d901f5be5e4852a91bab84e2d02c538f53c7a1967635c9cd3c1ba09e9bf1e30f41500120
zf01efb005a8f0998d81d4aebefc7e0a20823ec13afdbdd080f380d0a5a514e81468f47cc497900
z97af0ab56d32807f821d2a39cb0624bc7533d0118413ea416889a96c9b253e1859902e5e1eb17d
z9ebf31ec0f0864d4ba5412b7b9233377da1ccf3411950cd34e5c74c7587b466c62eaa1addafee0
zcc0587d417d428b10de519bcbd7186047e0ff96f473dd911ecd69c718b59244a815c6746963b50
z5d6c3ffd9de5131fa20cb9c84f99471229ce4c7ddb41ef9d980f5171ad2233edbfd9deeb630d17
z9835349895647238449a270e10c1603c64cd214ab9b2dcaa4bfbcd752b3ed677e2411f56dc8c3f
z57081b8a91fc92d0e226ccf30f8aae60760937bbb2c9f414efe1f0e980c8c4a3d6cd01ad7bdef8
z30df159df87c56a2198abe03e88a671406302646daaea68f422d759c8b885881d8ced22bf5dca4
zec701ed05ee9595b063d1cc444a6f6eb7e252379b8c05921076aa9ed69f9188c00505b6f16eee9
z0b01c6044132592d5f2639a00611eca0a7ae6b9606df7fcb07cc54f94f59b27e8c094ea37672a4
z388e5995a07e608ec064ba8be3ee428c2fb6a12e8b83755da3c569175dfb196b9a70036158a01a
z1832313076a129aacb5616994111f6b319e1288720d1f74e055fc30ebcd565e74e818a972c1e3a
za018780a5fcb9eecc067b96df5191fd4a348be17b9b96bf6c0af5876f30b0e3a84d90157a86542
z6fc2c40b88916be1c06f022f265c6c6a0981f873a27939cf5b3272d57d6c0ec07aae2ca61a270f
z8a5fa98ae2a7953514562b6056cdb98076b2139792f78dac853510af5b9b58703324850408ff07
z9a14aa32dd7afb6fbbb9110ac983939b9adc9ca2467908b15b665bc342ab0047f3f36f764a2d72
z4d7753edd15b20fb685740c3cde1b17679a026fea1b05c8252e7bd516afec97339c6561dc88e43
z332639e7e25b95a6bcd0265efa8ec152be2d23e374ba2e176d1a8603d4e643ee15bcc7127509fa
z593ba209ddd528599845ca04ec4e5829a503fcd2b6f32c47e4354fb6818e99b0d5c35ae04c15e4
z8862d17a72ab7653a0609b08d837b9a6a3569f6cdcdcb190b21e0d3390636e7c55fe7901877e4d
zc7ef19f2321f20fd6af3306b5aca14ceea2e098aff8e983fdd6dad03313e5e0f397a9e6d694707
zeb80158e744b0cf95c94f280e543584ea3a9ffb24c6116f357965293c7e1db0eac76792ee31a25
za682f2c3717ac86271183b7a8d26dd6a41f2a72c46f521032e51dce93f0ac006e3d5b94b9621a5
zb8f211997d7d1b79771ec0fbb40cf06f9bbf2ffbbd0a3b40994f6f7d065c420d824ce92d7eb6b7
z06494d95f57c2a68661dc4dd90e882b67bfb3235acb9525c6ec5444bcebe314d21f2c5e474b9a0
z70da5c70644980ba54861f776f84a196d710c3e053b821e7925256870a7f0134e83da841ff0230
z18cb2643c65d1f755b79d4c470866c37283f537ea73746ee46e41e41aa842e855c63182c34c006
z47f13df6f6127d04b87f56dc4e87f7907856bf2d1c34ca2d5a046552390f51aa3b2d309096dd52
zcd3c15422da3f0962951d434be7a7fba4cbef9f6b16ce69c8480d9a90e1520e33af4b533023899
z88f6fe81ff6dc11163576dfe397942238f1d58c8eed4e0a72d6ab83ec823b85d94b231b5b2b7b9
z2bc318c70d1fec22480882ab34e984220e631c30c9d032ced651ba8e0aae9c9aed1176833edeec
za4df40d7ef4ed704570ea73444cfedeb60a36c7717a514395f78d292a56691c0984be1a13f5770
z6e22c1bb2b1c188f2633d7c5648621b9b9321dba0caf941ddc86d9085d120e9df07a3d0d906e05
z907b6f52a5fdd8a270c51bb85111babf1dbd5af2d0bb5673a383f15868e44efca6dec34f29afcb
z29ca34dfb3ba06c9037e88908a36d1fef44f726cd8f8331ab056ace7a267d4d85628eed2ac0f12
zf3d4a37465cf85f4e2447af0db28bf6623110907b7bce4dcbb729a6e5ce6f976c918aa1db6e831
z1b644ba821b554194f957e01d06a155b2e90ece1e174dd5fa24f4cca5fafafa177d8cd3dbefff6
z816af892bc66bd8f4332aa795cd0e7b8fad94eec47079db7a3cd4438a677f079bab316b119b79e
z145901e56f30c159fb0a04377615a5b8403b1af91069ced795d91a6b0e0eeacfdf5769ff26b7a6
zd69fd598b6f4761df0fb2a47ff8d3693ca074e473a3a03e353736f49c6a2e7cf08f38b608c138d
zbe93d8b5566e45b79374e2a72d0370e1b0b16e6775361db91fb5f12a580652881d008b31ce39ae
zbd25966dc608fbfb5c83839e685df4b08b895798c341522e52f3a325880ed5d13ca00e57bc13c2
zd8c90de63cb3770056f579da10d8c86a04355dc2482b86b8ee01787b8356a009bad1729ce427c4
zcb155405ca628ee501a464a9ecb6d9ca8e90e71ba16169a07a58ecea1636c53d4b7e5919efbd6f
z5c5646d89fe90c31291ac3644baedfb7bd6252707395608b0f5fcadc00d2cc24d282af20de886b
z1455ca2b9af6a964c9c6e5824c79ed1d3875bbe695e738a8cfdb783ba1ae6d241db3ee56de5dea
zea4c7e562de7587fc2ae2ddfa29e65e5c8cc70d000bede5993a95420a1afb66276d212e39cf470
zcb8d9c52e9be54ed254511ad9026ec25798b429f9db40d1ca9549494c3347e34359871503716b9
z99179220398915ea6541fa389ac647297050e2a73a3c5afa7f798615d372cd16a7989d031af2fd
z495a392a6aed6e5b5a6f419e300fd5380ae836e0aa0bf4f0feef318bc29e698a552977284c2cd0
zdd5b124748b708a075a8395314aaf69c6868048cc1448aba2a6761ea368d07820f743cfdd67886
zabc8205737050bf6e823a47a8ba8697c552690826b41be24cd9a5f24f56fab8eaddaecdcfa6186
z7dac7c5e80abbfd8dcf67e1912cbc48e0fb0dab64931270bef8bd67dd4727ed054375d9941bb26
z8cd883538a3e6e13438c69b450253e62570c2df4221af2e4fd46885b91bc83eae596433e626434
zc732fcd99b1104098be2eac4af054df1c4b705dffdee23272dcf1da3cd76c42060506ce9102c14
z18947f325fa19a61675c45e8bbbebd4c9f3b8f36dc1bc7d53fc5de52948dc367fb4ff753535544
z3b0c4924f8b153182574985a10d0131886ad5b997c650285728060d8d1c10b2aec2172063bfbb7
z642fe83e987196cd9252fdc7a11c370eb98c0009442edb26482b57b2ceefef506d97416877d519
zba6de55d0561806c44974eb8917c45b68017e7e35f88b35e8593d0f4c4295e0e6ba1093bc6d868
z42b7c70b7ed28d83ac7197be4457691be51447a1786d9d3fa99629609f44845228338e85369005
z0fc56f79c6e6ed60d211492f92014b3d3720708d6951510804eac9c5a8a6de054b1c45a25d3a6f
z04f20fc7086b711a9c00882930ef253d464a72ddd4a763d826967ba4e61cff03c670705e86aaa3
z4eca64edb2f607f55c8ac070b5404c06cc0b6e57ee61a521270f91733def1411d76b48d332830d
z771bcbad99746781d998159e19ccb88c5c998d2074d983b4940b272356aa7305aa4bbf75eed6f4
z29181744988e5c41a8f92e37d6f13894348d34f5a90458c2c4e56eeb7bf11bea3d2091cbdba6bd
zf13107f5cbf6d7613f84384893c2eb8acbddafe0d9f04172164dc83f8d3f0e4a3e51c6337cc2ef
z29a7ecfe3ff420f18cb764207d5e49c54b30fe3293388d15a0da5617bcf769352ea31e25c712fa
z6bce69cfb779537abd4b5ac2273b78a4d512bba723a18b99ed7afcab4cd2267d5b3b89c128417d
zfe6478857b78cf720d48b0d2033527b8602adbbbfdd6b48a6d9581bb79ff8c006ceea68ce4d498
z509d17dbdd03c12e2d557bb264b346804cf2880a5d35d68b84917aae2b17a9180990eb149e97eb
zbf3ce6f7ae44746aebb2552bacdbac4e4e2b8cebe1e283faae0b765fc2bfd96fa44de5204753c2
ze8f883eff5cee87b148199d1f74e9524717b108093549bb0562841e848f011067fd6a8f3a95c4d
z79ed38ec7c1fc7092c2aa10b90eef26d6a56888ae8749478235113f4ffa4b0f5c82e6ea2fd53f2
zb14f7dc01ec55eeffe29d7ebc5ab7556530a9a3760f098cb4f4494f9b21cc4547e1bfd268d8e92
z557c62f0b0857723635a772d0e5f916ba6ce3c0d2a5b05dffcd8e3edacf7de458fb3ce17f29ca7
z9d29cea610d7e313d1457e969f7c0f5141c34a7abe503e006ca0e4782fdc371b4526f4175496bf
zce86950f3775726a3755d3baa80b9428705f6151f6359745e07636867ca6a721f5321e6bdd037b
z02234b9407056deea66769fc8b8b954c5548388b5d68bd16f0486a726c9cad8c0ca71241d4d7e4
z33114d9bea794c1773833134f53853146b59c1129791f63256aff061d6a00c5170d8bf2352f496
z2176c0dd113eb7f8250dd4635121a174f19cb9df6278b20ff87c03877fb7df660bf6b4952815a9
z8821885ac15c473d4a480111692e1be68dc9536c53b4d05b74dbc1970411cd4670565c89ac3c54
za846262c76c930d4db7990fe6f8c1918526280fe05d81e57ce5ccb28e07a95374d10e31e62b038
z20678dbabe2b1d5f420af5056fa4c2a488316338ef2648df77a3758327959eaea85f8b260a17ce
za5c281086107c0efc5fa60d43e4ff8c730a6066cf56acd3c7877f4a6e5829e0631f7f5247c7907
z9bd4754ab57047e76e28f236af929a858437593c0a79dc28b87d5673fa63ee79c8394458a12f65
ze4b0fb45f2e22064797e2eb11b9593071638e3a8fbae06df1c0e93debf3fc661acaf232288266d
z40b5a012380c5efca57f2ce41a2cbe99ba1987846d4a45c2c2fe28bb11020787478df25fddf762
z58b847a295b4bae04c0706e74e7a4b636ae2026db1751a0e2ce35c8cddbca02745f54889582249
z9533a6c02f9594931224f69ea7dc4fc56313ff2ffd76af35878fd1e2405a6a331a8a343a51d2ea
z1b75adc073d3153c1cd4b45289e00952c544624298798aa5d372fe93f7aec3d170ea535f55d84e
z182df9886872f9b79a300d236f76fb1a014f9ff95353a41f26430a30edf7b197c3f2bbd828930e
z045b12866454aef72b892f337d463bac732e0d868b8462fe9f6726d4784aab477ea95bada4381d
z45b69a90ecda4da80773c7f8ff55743bcfd7ee0ab57c9bdb63cbfc0612fd6e39c01dfa396de79f
zc9d307ce47276ae128d2ea367acbcd44f510d67bef58d7fe49cadac85473f212485d6f5d47600f
zc4512f998ce65a6cc76848017383ff56f2d34da23f92a4a7e076124d62ff52748d2e46a51c1fb5
z39e10977ec39470ff52f840d5aff41b82fec9ce6be65507afed37638f0a64bb1d904e570f90fe9
zffdec6821738b30e7fb873542b0ef4c807e20fb2167115c65a28c9e26f3aeaa83983920ac463be
z6dd2683b3ab47ece4511a0b32145c0fdb64b1171e71d5cef1eaa0a8cba6ea0ca7ed1dd94eccdf3
zc3af99527b5a1fc8c3959cbce6740c8d307dc743de232c1f148d042416b6c0ca7d0a6daf407431
zfc23d4f02acb6ed8beb5d3ba032a71c321fc4ccbf95e1109ca55941c1ae9df19a366f677e35424
za5d71a1236153d236257555dd808cc00a3c94dd80476f174ba0d745e4da295fe6d94b0fd0d0d45
ze2266b64c3f2b129286c243f777c3a4f9ab47df6407f9c7ae3026866f9359badad33c9769a38ac
z78a71581c3e682b0f57af6bdc7cd340f24feb28a7e264a43e0b079906af627c45738478a491be9
za6caaa5625d4d1d90ef239cbe17ce45a91b47b777e46ebbada5d4550bde40bdc780d0d54aec269
zac2de96684feeb4b2514418354e6e1bc90efc7061e4333418e5d57a726564367ec2bc7241e25da
z3bece58d7ccbc468c303284c01b1d327e4106bb1214f6004bc38736c85d4127614d902f4c23077
z37a6a2b60278cc615ff2ce71a7ea85a500a781f11448f018b43d0521f0a343df61b1f46eab0d74
z1dcc74824b29e954c9384cad32326d07d85ccf325bcd717c660b876d867a319ef07415cbeea6d1
zda1f765ae18119802e67ce93838973e57162a70a98e5b4fd90309ce54d8860901d3d57ef052227
z159c50343f0010b9e5816bba6f6810e8ae7c6d6cc2d6134e1944fbacb8e296c4fca4684b27d90b
zd9a7dda8556bfd37ae043f7e6a6d74a2f8adb9d66dcb8de7bb373e41ceeb8acecc678d50389e83
z41f40b25e661d906e5558d49fa361a23a7eb95dca2a9c93a7b01ba8780fd1ee408631436234786
z89ffd671261a1a8f0572b4a84fd5fb5fa4987ab75fad7c99157e462c7e1d211dd0baced706e26b
z44aae5f1a238113ca8e28f08e453b314549330816011b5a3ab2b5ffefa6c4690757da62d952595
zffffee185003f35b968ec80bdf125584a66edd3aa9bd8e4b5ae1c24e225c64f3e3140e0dc31b26
z669855987613d6b1760d416e2e5bd96d427717972ed864d20929b823103ba73e8ba734b93ae674
z0257b185846cf4652f35da0bc0aba53ce51b5919bb60e1bafb2897ec47e38a31913d8f627cea3a
zb9cf40fac44d7cfb779ea1f9c7ab2ed261e518d493dcbc331c993337b91c3e9e47982f58a7b94b
zc213cbade372895bf8e5be162100e9cb1894d75c6ba361d2df67f19bf686952b49d4b63c109083
z34d283aa3d9b9c27de669104aac350a3bee8fe2d38368a4e6d0f3df7c9add920ce3e8baa6706d7
z80149e7cd3166c8b94454bf92c35d57759bb3c20954376ecad9995bc7e15f1cc0b7f5abd92aea3
zb26ea3f939cfe15839bd2bd830c0cb28a0d5e0a91993bc9112931dc1baa2324c4e452c8f825978
z1dd75744b1875649a056dcb3ba5dbd2279cf316e5fa3c2d275eda28d9ae1b959b8fbb3f6694635
z3415280c8dd03b8138b3911f0c2885f03e53089a76ba1938927ae0eb40d4a73f4be26b20db9ea8
zcf7d9d51a25020c4468c6b2f142b45f6730bfb233dac564e3c587ca4eaf3e0ae0f6380920f8804
z7294443d87bd023f05422c1da6b059d278e900e776ea730b29d32b66f8c638d2d29d365151cd15
zd019582a6f20b7a74c8beb411710d99b87b35434d72c8cc6cf93b759b644aecef57aa48dd82455
z59ccb7b31b0341e15dec27d0ff48acb38bac2e5b47377bd7d53865b4984d53512be3c3e4d8e073
z8544b81ec21285e71587c8b878ebd9f930fb33831a4ae6e426efd050dd425b2de813765555c9b1
z3110a2a337bd277eaa1c0a125b37baec1f0697b45c853e1f2eeddc840c2e3ff8a21e337e4e5683
z5d246a85769b44a3062c476742441e1655aa026107dd7bc33c407e541e39fd0826073fb15bc226
z3a3d3c1a7fc3d114bf50d7c365e7c8e073681e1ab3c93b868e29fc1db4bf9b3c8739072a57bea6
z87f235a04bc7923d7f661cfc03b61aff90823ba6093d1ffcad59432ddf82ebc5f25b55001b7134
z930ec24ecd7602a3cf38d4b6072ff3dd4164bb54f948c553251caf0a6c0c13570e55ed1c3eb68f
za69aeba01e3d95d08354bd868c5d46e82d934fb4853b870f38c9607f8d3bbb3107201c987b1ed7
zec5e9a00653c4792b4708616756daf772bbbaa81b9a48e5b8c3c7eb2a3ba557cc6a44c4768855c
ze3b738373926ba29a67ced2587a2308e7a88629cfd3f9869a0322a50b1bce64313bcb9801e92e6
z89b86e0fdbb8452b688f1bdee409b9c168f4a4f9c837c20560913bceb9ceedb22ae863570e42dc
z2418a87ddf8b8f34d2e0abe890b2a13f454b95dec6ba749b7e3bbffce93e9129f6d74b7d4fbcb9
zf88298f950cbc37ab9e09ccb5be235ca393b9b9c921ad50bbbea9d37011448c00e2be19314d9c5
z645361f3d6fa93a0345b2a5be2d0e638c47e76b3274f00bcce1e17c3ecde8eaac000917f607dcb
z40d33159951f3c2df9086970f1ed64903ed6481a9ad2dbdb0c5d384f6c7b6825491046b39c2d05
z907f4a961efaba3f6e341e3601fee97251be431173bda1db216de0606d713591140885d6d87df1
zc59786bc26c271c5f11c3d9f78e41a1f0dc4a080ffbc427ca7d0bc601346651021c13937302d6d
z403bdb0baa0e81a50e2442f17d96bc2cf9b84f9eb9d8c0531ffb31702d7b704d8434f3b09b0c4a
z38fa7520fabe3121da2cb1f5d5b88bc62520d1aec837d4a856a592df9580e4509bb8ca09187dc8
zb2572cb048600e8c60802fb0498961328e93f30bef514dc0d5fee8801135f160f3aca19cb48e8c
z727b8b57900ce29dd55d716d0a32fcffc484fabdfbc8a5431becbf131e80764cb87c914a2e45a0
z84e9c9e0472b331a3c81b7b24f518588e39211a7a4a1495b55051eaa3c674d365c0d5f3bc295a0
z648c0bcd53184d526ff5766aa57821b5a615bdc29d2a02ae6de89d85c7101fef187880d333779d
zf8ec653580aa344adde963d1198ab856c0dd0882617b799ad175935c65704be3632a30c45ace40
z8f4510f40f30410e21a5561f10c02ce2a4880cc810038c67f4863dd84ab00f778483fcec55e2b4
z4a6c20738ccd92253885d39329a2065cff6819b67b327b15ffdf04c8c13ec4b7c3bcc4b7abf3d3
za7f0375f8f4f223724b175cbec4409410baaf948b5f0a37bd457682fc7b0dc64a7d055a61fe8dc
ze516fd974e94bfba218853563df2bd0312bfcbc5ead0b690fe1fadcfe14ee51a53c3ec241cce17
z422a98c0ea4c3cfae95957bb4d928be8117bfb36b32d149ff561cd0eb35af2d359806c9987753c
zfd088977ae54a69325b88852c569ef8d1866aedf8869cfffdbf78c3f8e90bd3a25d05f0c3e86c8
z59527bbd7ff86356352d160cd7579405352af9eea4d14e8fa735c24bbdbc3d5879ebd763bd8790
z29f8fa9d72b1aade3d6d03e042061cd318b5ed60c80ad206e023d4f20a157aea54c11b2022eaed
z58d6ebd4399c3a98e91fa713566485d526b31d212ba7c6c20e9b4e5d74d0a7406a24134e1c551e
z45b93436f77d98bc0fb70e8eae37c0bbddbcdf30b0b136aa87dea2b96a05d9041ca12ef706e69e
z03bb43cf98848d9ccae99f588084a898455de3983e59d0bc287c4e4617edaacc2679574c1fe156
zcc4d8d57c96820448f6e81783bd2565fe2cf2714d3a7f72f205d4f627bc4093890fa8f6f8f2483
z37b1605cd1f27dffcda009bc3ff01407c89e758ea8286d13b73becb78c5b860f9358f8fe0cf6cd
z4395f76b2af9ca107b257e8b181b906521dbf3c6c3e48df222962d8cff5cd55e9f6bfb0cc57283
z4fa7ef06f5061f6d1aebfe1db095872efd226f789c012b7cdd658d202c41a4aa7983ce7a0570ab
z2f0b0feecb71e0fb7b5485320819ecab705c1e8586d4ebbf92e0b76a1b70896873395b9990ff51
z605262b5e62c18a070c0a47f6db4b2baf0b151b8f652f774e7d9fe673d1c2b33fbca4794fb321d
z8e82bdf04a512ec97cc7e82640d662203c3907debfadbf5f69725628d30eae6fe0ebc5e72899fa
zd797cd601ce2c1ae060c3b91ff003642ab2aa86cf7f51d82c9a4694e026dde9a8bee63bada8a39
zd36da2afdd67f39650d5222aa39ae786fb68424a5fcf205555ed94d9fa539f205102f0514d2d36
z110287380b0934163e3cb177d15058cf3a9e93c68508e9eefcd41b9642edb7a5eb289fc0e6e215
z2bd2e615d14813b3e6798dfb37d0cce927f7fac08e94e2c1703d97c38da92137656fe2e8b54e79
z70f312991b7a58878091680cd345aad432fc4fab251e7d079433c1c0e14cc7fea372adb620f65b
zb5fbde722c5e069a0ee0c9b82f231b8ba02a80aa1ad9300e439e08961118dadc732af3ddff835e
z5f9a241ba16ceecf0fbd88c2686b9b8a56ee72caf27467745af0c50d372654f4ac9498e8d4d006
z487c88eaa07ad412e238fd93571aba3b0f22e72840d4358b76eb3ea1d47c7b87d68f00015b79f8
z96b0b3f7f52cdad8b9b4277a5636c0b7bb5284f7cb9796bfb55c210b65cb3b9cce5f3bd5f0e3ec
z2168f0107ef74e270633e8720275f5f1972234f6c9b59a7608f50f46ceae0c088d6781ad72e3f2
zf97c724ea84eea1af39b16667da749f0e8269b07b51cef8db672d22709615c3dc2d4737ed04864
zf3b242af4705923fd1a21d16a4ff560363477e1088a1dc60d9e605024623a4b30d15253fd7cb68
z70650751288318d8533ad1f980649d53bd1d732caa32de10be5a7383242b10522b3b0e7bde836c
zded49198a0638c6d4301083acdc182b820b7af6454c3a2f3f34baa663fcd66c061ee61e3017898
z2c008a8ec265aeeb5a321ba9db81f1dfb3ec4e7cf50f108db3b37e631ce1c53f00e336c20fa5d8
z2ba2829fa860fd22c06db0bbe6b9f1fc14d51fe8a2c64c7305d62babcd2ed687d12aa40fd3be7c
z9b84442a9090c26150f691859cbf50d747eb9a8d9cd8f4d2a10b83875e2ebea8c23edf0d21517b
z11be8dad0c90fc39158a9e433a906b178719afd95eaa53a872d543276a13947f4a7377487ecf06
z09412a1752f09a86d7825f6fbaf55b0c92faf690c6b7ff11db66edcd946a671f56ad3699992a9f
z8a4a376ca11388bb08036b107cdea2e6d09e9f022a40112f07daec01d3193a147484e356ebfc3f
zec77e1313dfb5cd3c6cd99a539c538280f78e88398922070a7f78f70d8876ef403fc8451807cf3
z2b532b138f483d9b71c3b38372f5ecddf4e64206d4c4630dccf3b9b991a1cfa66e9874fe214828
zb7b29a44ad270d995f4db78103a274d75a6656c235f625c393e9adc476a9e1c5d52eaca4a91246
za822d247c38bece10aaac39963afd162478face52ba87ee34def9484f10c6ff7c73896f46a55b2
z4a336829bc9b2b483351c3194051cf35badb2a1e844497bf551a2801d025f001ede2642b03e7f3
zbc8b7abf9e9f9781f945909626d97f839b9517388b94f4a817e6f0c24c9d3602dfa10410421924
z103583feccf6d4ef06a2d8f69384517abf4f89851c65f7d51b6286430b822bd350b3d0c38f7c85
z5d6eb1e4692736bc19f132292070e6fc51a7e59f9ba9d4e6ef0db4052f65c6afb8381995f13c0e
z36a6ba2b76487776a9bc21f259b4db1cdafb7b10769ed83511f7713f2c9416536ff67cbb0bdd9f
z4544da333f33feb0c1c7417a943c0f3e4cc7c6ad1bb8bfa7ee9f5bbd55c682bc1f7f213538efa7
z560f312c108c29f93fd3375aa778647c9827212b2cede3bb30c69a57347aeeb4a5febf110cf6cf
zb74cf16f4a7a83dbe4e1d70e633fd992ef506c43e61d9907479eeaff53811b66414631bd749b34
zae8fbd6368d3fc5b2cbda7aad5a90067dd0b7dfce4c1c3ee2cd170d56b741c5db51dbc5835a557
z25a64575c28092f4241d2eac2e104bcb3b7b0864d088e647ca77dd58072e96845b6267204b22b6
z02dd7ba7f2b7674165f43a23c9ac4775400ec480f6fb45c93e67919cb8f049d5c383146db63bd1
za91f30dbcc678b70f0a07977ab369fffd701d3b7b304ce763310832d60ab24f32108dc6f19ef8b
zc000cdf7a91323297c63695a9f1f1f7ef045ddbdc2af1625c7a950d4a8951fe6540ed3ad5fe37c
ze2828a19f6064fe4eec4303d4aec5b0082eba899d4fe80bead43495b40e7b4208643c2e1c178a7
z448a615fc45a5dba4f87a50791eba50e03c434d19844ebcfc6f9b99d5e4526e3803cf3f614d410
z0adb25b88918525251b1af96b10296adaae2b279b12cc54ddfad60f71bff680a7d6f9ad0e77220
za3c9492c16a61d71842aabfcb9eb7c3f5eeef72105c83ab35c217243202f7ed123af7b865d589a
z1018f9f14374f7d18cdd68413f97cae576002ed63c3968aeb7ddf6520e86340c2143163e90594d
z65c69e85a42542b425c5c86c2132494c3a342559aabbaad1e9642f8b61b692326732ee24577edf
zf5df73ec375da2a4efe71b0270fc0dd9da6e77602560fa0de7e5dd9bc3790c15a7897cdca60daa
z70051354ce6d7b3051bbffe7a81a0ecc1c3fc39f51b51493804dcfe2594d386d6c8be906906c4c
z5208dcc717deaebe853e2e9dbf0e7447a6f5d1dd52a8445b7d3a9cf120d02f18a6945e2bbf782a
z20443f8b5a8b9fa05e81c7781bfef3e1eec3b911d668134b9e574c882d88837270145f7c2f009c
zced2adfec987f64346a89d212be39b5864a4e7f76557a9fe663a9ce88dcafaf2db1e22b79c5a47
z6d6dbb40bde569f633315a0224579c5e6b50f519b1e4aecf82ad916240ccd67183483f346e9066
z5599e0aa7b6c9a837753ba1b0431b337117e5d728589c7b212fbd8fec0ba8d289d619a8592ded4
ze36cb69746d9de20c1c38ebb127057683ac1fcb541b29c7483c14911fbe71dcb8e262dd4db1dac
z4d7ada7485ff3aea9795fd55d32423df510e550e786fec6b530cfd1c8226277bbd2deb94ae5727
z4194e0b2495ae36189472228b47d479af342098442af21fc0d3e7cd18a7702e36d06be40d9d55f
z1e442c56270d0b2ea65b4e7dcafd0fd7ff0ebd5060c9a576771848eda57d33c9d2dea8e4d7cd32
za7985b297193c65faf31013c727617718fdb17b149f13b0761efb288c376e17afa4f0cbb46e222
zc8bc26eb845bda696bd9434ec0286e3378d4d8627b1f3dd906d6c88c52add77a690bb7f7bedb98
z1120aa4ed3df4659aaf53b21d6e95839b518fa9b27668bb73dc736296a28f21b2b937e1b1661a4
z4204f1d259d0fd251a524834bfa12443641e2955195b313c97aaccc92f0960d9b611d288f25dc4
z98db5b88cc6a6715a8c2201a2b536c95b641a417bdd99add13b7c186b79e23dac3e824c9e5ec50
zb4f4dc254cf2c1276b19cb6c9c88766d2078075891e78906d9d414480f332607cd9e875c1f683e
ze41189aa93a663eeb6408602c3bb33a26527b2edc903ecc721ef2c08fd93b26ca9d44ea435ec7f
z6c16d612a00d19d9cd7242a49af7ea589ef6b7cd603e98e3e8eb5d46bd04b73d7e90dd015a7727
zbf8f9fa066134865deb5db22f6e75cd9a6b8144a30cc6b4a6f1dbd12e97f59c94d277a78542c8f
z358e79c0fde8971c18d085dc99960fb0df624e4efac04f09bbba34c837717ed4423cbf2dc0a016
z1ade1fefac02034704fead04d8b7899b3f7347c9d35f75f974d9115664a98691e55e4df15f70cd
z1bbde1e1606dfc52699a7f89b133f5bc5c4533903baf8dfece5d5bf8de134dcd54d41672d6f8c3
zfd84a5c40804f73dd539082a1289ab67c70f81a2fb908209860fa32c270e50f7d23b71901c0cf4
zf159722fbc22bf397fbe477d9469eaefab752ed7583179169431440f807adfb3b04363764e8df0
zded2b998033663fddd910a614dfe249a0b8574922a6e90566ece35e24c5543303f17f580d9f82f
zb3a7eb9fb1ad42f3c5f1632577e893100d4275868ef18046503893d20b816f7852fff854d5aed1
ze9bfb6fda1d660c4d0df8efcdc8e1056d7521fb3887a68951eddf19b62990779d23c5b151a6798
zc77dfa500b33e03429a5226dee8ea8377254f18923c2609c389062de907760eb4d4d4751386132
z5fe365381b28528c0f7b8c64e237d607eb17c6994f7ba0ac68ee3e5200ec3842e886452b313a9a
z7c03c047e5284cc7110b23f3f6242dac1377c1c1488d55338a094fb3b7bdb52389e969bd7fc0cf
zf5584968915e803179262335090e1fa96f06765401cb202af5de89fcd23f1c0966e760c06e5ac9
zaef35e32e2234bdcadaa2c938d35ebe52f43572f8365ce8a6c1ef8466dc128b95cdead4b10a6e5
z48e43af93138d5d7d33979935d81d82f6caba0b67f6a1c080ce9efe374d9f86bc6a92572ac836d
z7192793307b3a236b26584fceac2aec099b7a3678b7891f311615ee859dfab4fcc03fed9db1e22
zd8cbc1ba3800b3710df1a7efa5febabaf0c45b6505b622266afcc4d8c51f444401edc774151913
z4fb692fc6a05a7d0e7f46ce5aba0292dd3
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_sas_receiver.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
