`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bcdbfdb1f2
zeefd6bb31746e3ce8f77c3840cb2256360194c3d47ae2dbab74c0906f37aa384cf2472667f53d5
zdeda35e5e25a0da86d76dd5ba9c3e8f1a51e0c7985a38da19a268fc0b58a1952ff828cfd84626f
zdd24efec82c8a9c8e659e5f9641ee91585223c6778ea5487d3771b6be3023f1cd7666ab4846f62
z177887a462ad5ae73ef8b11330acd6c73645d39b006f27bc8c1f4555c34c35674b569bfa76cfe9
z8559c530f1494896efb511b503f1625d48c1cce5c00e506edbca8b28c578f5c39a0654879870be
z641740a0d39faa9854e6b629dafed2dcab821738d3f824282ccb8e3f8ef7c114ba2d906468aa20
z9e2c87b0df5f26fad95ab7f4a2b83e1319ed820ccea3ba58bbda8b8c26b5505ec5f285bcef9f51
z2cc7a9749dca125700ab7674f26103b389eac129d3638da61441cee1d479ea984cb522e7696afc
z00f37abada99a27ed5c5e62280880f17bfc41a18b0803de6742ff445d6800c1d33ff0283d8c7b8
zce756253b21b2aa046ccb7aa9ed83301577776282ecb48d6c55f39e6eec4a2dbaf723d45b31ebc
z16a23735aa0f6d2a55ce5cb3773885c36c1030b98ea75a5772071a672823cd76b5916f76028041
ze4e4e127290572e481c7e1df25f5bd40984699d73eea1114cf30936d8ecba534090ca92fcd42e8
z11a513c65614c939b3653d1ad59395aab2ecdec54eadcf4c9162a1d173df54994d87940b952e3d
za4a0064eaf649ab6fec770dc482c3fc6d742bef87322f7d0f5ad65858ce24a33f9107673b3716c
z7f4abababea22e9861b656372e91effaed0847eccfcfe85ecca0c7e5c8c7bfec4d89c4d1322774
z3fa15607983b8cfcf277485a3bf161d6032edaf6015202e9919bf726989bd4c6bdd9797e30cac6
z2b9e4108b4702ec8fca98e9cdce351a6b7f7bd9e52a858a9d657df6029a972336ed1beaebdce17
z3f80d108d859e2155fbb5fdfe389e539103f54ca99a173eba64c8ac8b627e0bfb347de7abb9ba9
z98a017c318dd8820a90805fa7b3572134d91cfca3cd89f3e47a0ae5bcb3ea928d3e9de257a7ecf
za6856636e3fdfcc490ba52bc96b1718220ca185dd412eba3cf87cf72cc8579213505062b761414
za15f743e0d5604adc8c9154656b57bc9fdf3f71bf3b06ebfdeef07510cf0040fa8b17c9f174c22
z8d4cb9923e65f81f8535173223c252756b4fafe2997090871d9c9652ea6573ef8c460da60a5eed
zeef0c31b2dc5ea5e177985766ff1fd1e43b13dc8fc0aa908d118893d5f34e0ea6980b5b15c552d
z19dc115e4e7b2c46260b64579cb474624c4b99d20d74d8e7e817a7d424920093ac47f5a21b8b41
z5ef1b524d726125700473534c5591dbd12375c3935a7f04e48dee7136b9b75ea8ae11bca0b52e7
z3648447a14c32e18a557c0411704f3330c2b873e31b1d1353b7b4851ec9d3091db9f1696ed3be2
zba2957e14b28d8679a19fd52894e3bd000e6396c0d742156a567f65653e1b109a18fc44cb50424
z73a209075160deb195bda4b0221ac8a459ad775c14852ca6e4b5374e85beaa9968a1499fc0aaa1
z6207d1677cb191c3f8acc3f950e9d2b97d9e7352a2581b2868d0b15b125942f098d0397ef0bb27
z0f120ccc1545550c10ad53ab40b0bc84f2a5b502353600acec414de00c8f7d5e2a66e9f20af218
ze5fb7df6873bfb6b2bac4690c872ead04594da868f516d229f5864dc4068fb477345c655b05ea4
z9ba89e389ac6122e8ed999a9828dcabaecb3270e8e5ee195bbe37b5239bf546be9dd3baf948491
z88d1690f974b3c8ccc22a3e3a387823fc7b839881c1d0f3e70849f1366918832da8c664fe84c76
z04c00292f7e6ec44ef267646416bf76add61c2bcfdb4fca66c90d13d05123695fc9316ffd96319
z3d078ec3fa2ab885dd6aee0a6f410e398b003653a9a6c3ffcdafbc663982495946bea0ec959d47
zef8221caf5edd9bb6414a27efae36ff2340fdbd8671c47d274d7b778a0f2d641cf668402eab36a
zf8a0fe758fb7f5a1d17a837fcc20b734afe792b11a1576b97de38b81e80f2bd7aa4e7854c00730
z3eba2d5b76ed3a98454ee4f98d1494e73cec9874f67101d7c247165f159a0bdace7f9560558b8c
z074fb17bacd44b9debaf7d326faa6ded719a0bc041c1ee3dc980923a89efc016fdbd418d2459da
zd955e676917d2d16b33c21bbd91a5c3f43cbe6d2ea63a48a7c02d46c3ceea875c1112568519546
z28d8f8092e2380708f7fdb5e1d4fc695a067f90e65be026f79aa9e383fc9eefdfffc73d89c5ff1
z1e8efbb03b1f20613164ff5135600a45ba595154a773821941fe237663e7034ede1070d5e84057
z0f9fe44d07446fe3920a4e96b8943ce318c2214d80d7554d879acf988e62ae270dda2115a73bed
z9538635b2968ed75d645ac2b728da29224929f74b86e10a3162d7037ff1216f56d4b66c5274fc9
z02d7da22557b4edfd4e7eed12a362ed3f53708e073e289dc8f8028c8c25d42a99aea8c796c3d38
z28a81221ef421b37b7bb3a9fe0f90c9c3c3fbfd74c32eff9919c9db5b12039574afdfc462ea854
zad6ad917f1bac20a3aebf8d4295aeb0a0ac4f9160d77d85ce722541c67dad4cfefcc21c1085a25
z2719ec51ec957b889720084618d8e5b468326f1e7b88957cd8a069315b1b939de438bb6fdaf740
zd1b891dbec678803925e3942df863fe3bb8b2dc3d92e253902444f8786d24ff558f52f10cdc143
z0689caa11b4caebfdbac676606f22a2bc2eb57edb2e0ded24fb6d701bb9e2b989344a0a4c1101c
z3203cc511e87082f034e42f0b608f80153fec343c1f62f242d3966b4d686ccb682e1187036d8e8
zfb7e9069a247def8efda25ed134048214972b83188a7c4d32f29645f066fef814d5c6ed96069a1
zdf66a469d3fbf2aeb835a9c14802b4ee5b7229c650093ee5d2fde00608babeb4d0d9d73d1d85c8
z4f2134cb6a4fb6cb0ab216bc75f9c410a50f77a8cf6eb5a383132ba48839680caab73f98b3d7c7
z3742f9618e6757513dc65fb09315a201f478b356a94ef1abcd93e279c7c11d953bc10cbacb8baf
zf1cdbf70d7f873996c1fd5929bd3f0d9a81992db615cc032df1441f5c232e13af47a0f5e8cf557
z393f6ace54838f988ff5ad1cd190910b7fee04bf44b66e497a2240457e01ef159bbd8910625606
z5e1138f8e04d51cb619865a241a431798857eec923e785cfef0cfa339b272e069ed173851322a9
zb5547cd3ad07e27259ad798e8e980d16ac1e1af9d2a15b870ae795c0c5b5f2ba1f97109e695087
z47dfd4d75663f6057ed56310ea313f295fb9066a4e2eb8f7fd1d005ba356b7121cb225723237db
zf66258e4e7c213fd484afab585f18d88815d4fc28558712cab9f691b9f57eded417e46531353bc
z5070da9d8a40d5476ecf61ee70281b1915a56932d98cebf9ad9c8f0c83c85320b62732ea9fe606
z447656102134a924a83b134f36fd755af2926170af2b8ca9e5c8fd496698cac6e63da5b9ff0793
z38af003da5b32df4de53af25fd8773247bbb381b563f6bd4adf4f20b6456ec37e5db75d4c82f90
z3db747e7c25fc7b4feea2d2e45e80f365a3d4107544f8bfe2866e5f733c103309c398c5969fdf0
ze0683d13e03b39791a49c162f2915e73deb6f1dc1723d38e11ce87e1d677afc1f76666615d0117
zbe6bf16b6007b1cecbc66034858a45b5d941c0b9f5ffa881271e15ec1afca94be1df6dded401d4
z33038f6a6a94ece99728855681da6d7243bebc8e16161a93404ba7cea4dd1a447f747724b650d4
z6d32b441690023a11556f1d972e856dc74e2b5594b2894d6e6c4472d82568e5a11cd429d30c6d5
z77e3c2a1eebe47fedb9cb5f1aa4903cd111085c5a228dacddf37b692df935e1ad8fd32155d6ec0
z8ef8774f23c357b2dc18f6bf3cb006ba3debd2703d2598def31fba11be0d8a8d1212d53e1f9bf2
z9ee27d9e20e1a6b2eef391252c08d6fb7e54cd7886e1ff1b439d82d0ba32329ff6eb9c73e1fde3
z2e8dd2cefd275a0478698ae3535992251da93f07434f1c4c6a3b1acb6c9878ee2594b80a4ef360
z85da1a28e232a421f4e032f941ad09a5baad25e223639dca533f60fef27f67d3ad23c9bf434e5f
z40a701176df31307c45568dba1bc10a413ffa9afa30c5d7fbd44bd642b7095886707e29c980705
z7341d76e02dc3b721ebb007a7e8178dc8aeaf084e6b42890e0a66869dad94135ec7036daf6afbd
z413fe50b30c05091a1516a74817b5571e6ded0eccb92203253070f6afc18c5c997d6a409e4d7b5
z22d4db78c38844f1d2936507b2b7d9e8c8eae9f30cc40ac3ca23383027298c29acdb03d4db27a2
zfae385db4c833dfa5ad5e298ebad0df49727ea4e0746bb948dda2a97c3d304ada45bb43666fd8d
zf9c839f336cb76d479e260d9724c8fb44cd3a1882fc68615e5bb2710d8713aa75fc07f907fcbf3
zedb9a1b7b43a6c480efa9d732ea8a96b7f1e168c76e498f47a3ff81d1287fddc5120a6dd8d0075
za312d2ae3e23f4f1626d70c38cdb62946004458ededb7b691da15887c44f3d2c13e4c355ef8625
zde376e5812d7e9a6ca91727c15aaee83a33f00ed50eeb5fa14a57abe8db2c000de8ba30e17e4c6
ze44871b6f1d2253cdc5d1d40a19c2db882408cc9d1c5e7a8f393bae54bbc7821aa482e83c1f783
zdb248ab30d704f27500447ec07cb4f6d793e04f36dbfa5636b7d25df6944c51c0d99bdf9fb1482
z7d1b01583accff53a40af1927d60a6ccb45c2d08937a0b811f0c795bbd12c931f1aaf569c3a552
z687481820cc04e924c24e9303122718300abf144970fe847d08dfc57fa35fdb7a666e9377a6aef
z1fa56908c3331131fe5b710840df710c5850ef47ac77f2496f5a6d4da1ccae88957335eb08bd32
z04a58a328b19ccdd0906feeac771cbbc15b9a66ae4607a0f9863ded9dcfd932f9b98ba1133c757
z3c498cfa62f3776bea9133072277b1ab577417e761b0ecc264f7779078f47ca5e2c2e3d8555740
z3ef66151975136c394b96d5e59d2fa0a0da3cfe9791da64341adda9d1d38df521ef169310ae88c
z3b441dd17a7c34c92be55caeb9aca2df0b3191633233cb4e28ec6237ca6cd70ac388db546ce790
zdc9120d76089b8da9263d2685b35488b9cf3d927110c5663e51602d671a86ac9ac402aaeee8f83
z3e0dc6a5ae9ae46b5d434bfc04b6c8189eaf0d046a44826e9944586e47a38abfc960b68d4f1e98
ze426db857605914ad7f05b39f4d0f6849abb03d7d71dfafa63a4bca1b895ca57ba8abb9eb798ff
zee0943cc2b0d0af67d365627a737bf3137ec82d3e876b1b36daa95f753b9e7c64d77a295b42e5c
za07ad774188bce56793d058e0e0cfc16ccc880594755d6b78007f1f7c291dfea6c046de5668fdb
za79a4c69c4aefee0d5435654b20b74c04a9792f7f30d5a8c6036c4c464c91688155a154245dc59
z4c58d4c654c5ab6a3a5a9f787d97a1daf72bb3f3298cb3d1116c00181ac3eaa693b77bfc4d4efa
z795f17130e1c66d0b546e8ce1ff47a2e07f5bb69f0ad29a1b8af5b186bc8c45253a333d7294cc0
z290f8de43604fc2eb3c6e838b731e28c50ef89a3168b451b5f657026dcce6a4c9c48aecf6158d6
z957cb0a75b15449c8b76c2698deeff5719d72f10d399ab08c5150f0527a5400de4a2ee5c4a8c63
z772602f5bedbdb9cf26cd0978b515bbf93c2b197fe01b0bd9c21f52193f0880d72c3aded4f0492
z931dc8b300264b6f465d657de96f4c774f54e4ac2c994676e9c3cfaebc86f2c4c1b3695ddc2ec9
z4cbbaf94045799b84aecdf1356af04a9266c3de8d59d166aa528bc94be159a83a118e41a61684b
z873a9696965650d5b3d6f80a5fc2f2eab310c6538c1a00d10ef37a79c315e7b6fd9ae5112c9d6e
z75037e18d5aa669d11d464012db4165238e6b11650a4d6b1da09b8ac809fb792bf9b1965a46e41
z4c8ea86816adcbc5ead1ed7c089eb0d2c861514ac4703bd48046740d9dd736e4f7c793851af909
z8180134df29116ec3685ae97d09445b889b4aefcf5101859e472113c5c780a1e08bf5c9b5e21d3
z7d75ad334cc4d86c254223601f4d77c3751485c3707b19b5bdb9214d7db30fd66d01d403144544
zec48253eef316c2170ea5ac25c1a2a98312640a075b758e6245c7dbb1c19c44aab6372d6cbe4b5
z9458f1a6cfe4c708df2a8a65dfebe8091fcbd22863078379dedf1f8886950bc2e3c9ea681ea003
zd0e03ae2b49300bd25d81a6561c95189b98f63a742ac66122fd56ee1180d2e9ae818602905665e
z9e0a772b3895ae15b735c90af0b7799b406fdd05de06f78e0056308b6afe5f50234d9085218f92
z2edf0165ab63a900894ee867d2cd1f30b67998d96d30cd1698700728411dd8f10573a7d2fdc262
z553a8dbb1ce9ea4dee019f16513c8159f3d0483cfbc7fe4c2f76a0ba0d70fd4a3d47d86167500c
z1b59c78775ac914b9ccdab01a40393dc485e4f1869203bff3c29fd3b8f37c06127b51fa054559e
z5356bc032d14a65f13c3780e4711254146ff44ef32f05dbee92a0d5e2b2abaf8618c1d5e828b74
zfeb657df43593b405948a5bcc40ef847fa2526a8772cc3042975d1a854343dee10bd25ea0b8709
zd4631eafc816396acc4397fd24b795aa5b237d95525700222166d92fa239bdb0557dc9cc37af3a
zcb95de31ec12db012b3a2fe6c22ca4e5ca5fd7684b06c2c35fcfb6d709c69f2b0fa6075653d01e
zd9d29c82eecb29124b1f99bdaf997614a02a6500335bf10b2713ea647255186ab2facbb2c9b4c1
zd256130d2d40e43203d4867975a94cfee52498e2791d3900d1065a6de1a3452810345e55962390
za3ae183d3012b4fd8bbbcaffe1c313dae39efa92ff7211b8507e959122e14b129b86d1aec67f1e
z58c925997bb6248ffedc54a314b67a1550adf7efe4448f2f606065802128c6022c5186f7467f7a
z14603f7727e773f941b82cfeddee89008160ef8a7b453621d99e80baa2ff3193d46b2da524b3f0
z2b3933376693e6f8c00aab81e643a764428a9fec0bd203ebe729443c4036bb3024b3b0dd9b7549
z58feb0a4feb00b1d5d675b5d2a215660b60ca4e9bb7eae1283a4d6cd7e49f19e8a458c4382933d
z569fb51ec4527bc4ab4895c9e4eda055fe5409a6e5d16616084e36b49d43572657cb637d7030e3
z53d5962bd9b24382772e2072c71fba3e58d74b867aa7a87fad6cbae98e840abd13e3369b9a3a21
z32b05f9069c79b0a8e6bfe6ad8dc9af155e40912f2e6085600a7d74de76cafbf5b2b58bbaf3509
zc4910fcff06f22aa93f3571a9f982440d607f9f7e9d2a829de135037ff5634af2a1510c44d9b50
zd8b8fd669e6d16618551d952f0601d6e3e04b99dbb9e2d1c1a0570779cdb90a7a8c28c9e05d43f
z4594436f0db740eedcd64ae10e5208176467cd222416e02fb5f5fd6c097a8cce4b2a4e5f3e6eaa
z8b3a73d90932f981ff0739aeaccc9715fe1d91502e9a9e3962571f8cb7fcf5756979f11c82c243
za9c4905e6a13f64ef9e2c19210becc0b1a4c80d3f28a0465bb7813076a64dbc61cedbd4314818e
z91c497f6b53aeabc9db3d961658b66158aa8618971e106291d0475e58c92e9484975fca992c2c0
z877a812b4a55a078709ad7c6fd119d438be131441a40d052f2dbb39b22bef514035db049074749
zc0c267dd9ea94b7e4d8bf03529775df2ae6e5a8befa64ac2ffc905f749e0176a41b5004af3f147
z7c338174b87d6959abff5aad83280676a0f9917a28e2848a270bc33b877354297d4d9ebc198a66
zc35a6a68c361f9356ed7490230f8c5b4627222764b2ff11c69a2839f4db4deeb210bbabc7e73d9
z525e4cebfa32dc66a0eaa4aefb90c7d2acd52c8786532ba05d2346b96d1e75840d7af81a36705e
ze368f22a30c70e27950428745622ef86216fb97b3e3287d74fc3ad9c68e3ff06fa5f028c43e72b
z7bdc05a82e7ee7b259aef6badd7813d466e91f674dab4772e2399db993b1d1f0910f9e82ee3040
z88b5664f71f9a37ca2a39eaae23fc294ea40e3bb9aa587bbb6e9ef4160828577f06d3a68e79ace
z844cb36693dd674fd87be3b17c46fa71fca7b0cf458d15c4e22316cf7f7e1999cb7e8cae7bc4c6
z4a5e708a822146b122d6d0e23fd349b430fbd1b86f72c8b33d6d8546f304c7e859f69a4d027b68
z5859bbbfc5863b0e4eeb3007983892b675ea557029db63b3e7684a47016770e732ea5592e8cd19
z905a05e6139d57a038e17d620d72f6ea0be31a07be119c9bcf185bd418c7df640763c12a56fcf9
z2259e40e1ac7c5309899041058be7e9bd05177c4bafffc8764156fbecc3ddaf3fb6fd4afe14af0
z251efc0ddb2a08b17f694fa6fb33f8f2e1f796dbb74d578a10a5e19f8bda26e0891a0939e44fbd
z68d0202bed622bfb706c329888fb07162d94e7676dbd056f2b6021a2076a11eb07d092c34cd066
z8d97e645a53ed779c763f16e08d14db2a68ebdf7bb5103b7aff55e7322650916f82a4146b0dd84
z1da9db3d1a7f5a380624f5923495ffdaf525c10eb463a5973a9d35b14e5509a343aac8957ea31d
z70b9f7926d3f7a5cd845255c358786d09bc261fe408c3e4fc1497f347575541593c7880a0d1a92
zc7bf997ce08f6e7979afde2241072bab4bb023b8a504df424936c32828a5e6332f9c7ec00b78e1
z6f4e726927bef86743044162a6c036171e78d402e92de954462db5220948317be802e2a809ea53
zbb0363110b5bba92054e9e120fa2182980d60b2aaab6eb8f103916eb9adc180e14d0b7d76bc99f
z7b8966d01e8ec959773e5917d911847a5d0208399a0751b6c6318cdc94e23cea2038ce2b8c9bb5
z0826df68e0a50ff3ed9b8f4fa53b7db785e5ce3be4f87c2bf2b3a11696463aaa34b1909b884289
z6006ef0fd515e09e0387205ef6dea86129527d391cb9fc18702498ea14b5de68e4ba0c1f4c46f6
z2d7621c72eac64cebbb753856288b224434500b05f2ac8aa4a28054b375a2dfd4c8fbe288d71e5
zf5780f4f9e396efaa4fff38adf46f5617aa7a56ab15c8f89f6cee2babcdbda8bf35b473184dc2d
z4994c0474ff8e42858b4c7475378516feab1d487b7a997e3a508b032badeb7d0aacb37233071ff
zea510c760c4bc873a59480930f5b1da0ee914744b56d06a986c912ef4fa32085a2253220a7ea9b
z52bcae957d39f480f0fb597c86e684b9acdd589c4c29c8dffaf4ac838f94f1f0ed521363303593
zd78a963cad5ce07028d7c68e5be01cb5ff350993bf61b2398e5928494c1d03b78f7141a7ba8efd
ze061eb3d4da7732ac89c82227efbdbc5b3baf708b28ceba46a7fc4bef88febeadf7b4fe4dd4d87
ze7e65b9e0a021e9bc16623bc6c5bb37cf32c86c173c757a4b278a7d4165807af0b36993f3944ce
z8af54fec40388ebb9888f410862a0d508f984029c71ae515f87b47c885728aeef54372729b5c7f
za4a499adbfb77ca58b1dd8b0317b82585ac5f156887860b70d053bc0d27471ed1df067371c57c8
z8f57bf41a42a0c44b02e920c9303b59c7060b16309b654c6f80cbe9a30a421c08df814c7d8fc89
z685c06ec61bb001cc5f29bd38abe561b40867938b22c3366877d894ffb495498c158573ecf76b7
z6694bfaf20497dfbcc59f20b9ad3f1546c588237611f71b7b0a882724386d49e25ab6210f049bb
z4409f33191032d4502a13caf27f2a627e32a8ad690c4271b98ad3e963ab5b9ee5be45f67b1d443
zdbab8f0044d9584acdad8a35e2dbcd294c18c7f8d90a8055e4eec8dce5013422a024c861f916ae
z7aa29dea041a509c304f2928037e4f6c140b7d1eec7bc3a13fc7371358fa3257146602ccb30239
z97cc3de7d30020372fb1449ba9bad6789a82bffd91f8e831b5a8e334e943a0222afd8fd5067e85
z842904db51fadd904e3a4e35384492cd4a4b825e18f9e0632f22c84c4db93449ba38feae71603f
z02bbf5d5cc639ecf14da15fac1e72e49ac1e532964060d5f0bc704070e5a4c021cda4f3cc5bf22
z847443641b4301e812bb1af74d02530c3dfb3d01516340bcab983ae339fa34caf4b87cbc967956
z368e2284b45ec92403bbef793510e3bcef546c6465fe95cb5511540534e826d8f4a5783e4a28b1
z686088dd9a480a7544f986e4f1b572dbc5566a1765a30f4e2e14fa8c7323813985cce2b43236df
z0b840124247204f1944e44c8b8c16cddb137704b74de2c7449ca70a22d7a059f21758474505781
zd5b0c406135eccc816ca943403cbcde70ea98244c8a46dda5f54d059a8fc0e14e09e6d4b9b6829
z3ea5ffda607192972fb77707baa97dc72509676e2db7d6481608299a7b72590958c780fee29ecf
zb570052cd2afffb334b86af897d90a214c328034a6a3fe7c1e2ccb2b450b3fea2f52db466b27c3
z47a70c01ac1306d70356cab9799310be43dc66cb994850fddae4697548962400992e9e69fe64b4
z94490ee56e87f0c783552d4d67bf7c02f080f276ba2bbf41c01d16957b64c3bf4ec395cd419099
zf31a9c46875f94a9ff74bf74216f40a41d5165b137920d36e6da1b102ef04db9a0d55012f12d13
zefe81da7de410bd9fceae40cc985925ca504bccff5d98a713655c6628f11354c8e2c18370615f3
z979c3804ed928f884cfe5f961fd2290b589d457c91c02f5c9faf79fd049ced0368d6ea3d13dbf5
zfdb8dfd9a9b95ea681a073f8715379143d19bae5c5856d0bf6ba1bdb496db396c71a19372c19c7
z59a9e77e1650c577e5211b447376a0dd8c9a889bfaa9fb96142f71c7e808cc9ff7286abb61a31e
z54fbfe4e38fff7c5e13d006063308216aad56f43cd50164dd1298ca0529a2696244303094f5395
z513fea9ac9854d6196cd6d5929dc2c145f17ed3eb1d0cec771b0f2fea39abcfdc3d8fce28fd351
z14c1082655f6929e8ee0e2a89e0860deffaa354d4ccc07186685a57ec3f36c0e1fd1c0b21e2cc0
z21cacbce4be1e6387b5766f885343ceec80d29f6cb45ff9b34c2d88e3622a3db8c17e86bd75f5a
z75e1640cc945491a2cefb6fb79da48dcd79c0be473adee5a25ad7baaf88a89d7328b04ff3940b7
ze241a741839c37c295f03316cb21248f9fe54cfab7096c54d92c298df68f8e6044b23d9a7694d4
zf4b0c12ade41bb9c8fcb926f0c2357579088449993c5e2246a2c971ff553d7393fb6c7a4ffbe49
z1feabf9dc07e8627940bbdaf3b5c480df0bb6e44b5e47da880a83a3f5464d0b9335d832809dd42
z7213480a619b4995d83917c2ce309d2cd88f8c481cba727394c50a2e3e590629f22e359dd33c
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gray_code_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
