`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026201628cee5aae21fb892db766c4
zb5b1406e11aebfd6dfacc9da5ec03b70c276807a3eb15e28ec7ab1dddec42388b9424ea285623a
z248195c9f894b36317ca6e59c86f11031163f5f5bfdba36b10b435d36514783bc1c6e60eaff7f9
za2b8eba90f8fd9a9cd7c932ce34efca1757e6b2718aa68644ba032b1bdd74efc688b935cf38d81
zb1f311df3e5b8e4d46dbf459c824f309500192485674c175e61de609f1c94488da73614dd500c3
z680b7fbf510ef6c68927870992ed3376661d943d2a929d90faac51228c485c2005ea015bbf306b
za52b2ed3688d7ece69bc3ddb93a45ccc73f6e00673486a8bcc92acb7d4412090924945c1f1562a
zc5e0949f06ac734085ed2107e4aa9e39ce4ccd2716381ae81c00f915da3dee1704ecc26765111b
z37c91301861edd467e17bb93d5e374e1e91c3d7ba3c326b7180905901191f995e97041dfe92a43
zac13264e5f9c269b6e7a2b22e5cc8b0ec5aa75177e1c8a2d5c5456d5269c1ef0d82494bce3da12
z4598593f8470c230d8cb82868e2e8926b86041df29c6f868fafd01b20d15e9158055c9eca0eb1f
zbb75e94bdfb4e336e8888b859ddc98e14841807274add30af47330407dc3fe4317c3617f953577
zd4f5e2050846fa11e22136fe1d04da49bfccac468a90087d714c5853724d5847e1f7891ad9c470
z73306d6006d0e807052eed0126c794c03087ec8ceaf31379819d317f9fd5324fc9ab389e92c9f5
zf87f11ffd3a7c0bad30910b0a9ea77952d05e3fba0d239dde3f9125ef3aaead1e1207717047c73
zb189fa783b565c0b5b80a8e5c3281139cbce0dfdfe225634179911f45e0cde88f30c27de391149
z382b51a0eae4d2c9b552620c88057ab506bf655c16dbabccdb73d222fb33195ad5d88137daeded
ze8768562c518640df73740465574dc1be86f73f1a2e6f160ac27789bd73ab387a4a5b882e9f759
zbc93c683fc934b63308dc97e65d7f7ee1bab65c25a19e9fa02b58d7835ae7aeb9892e4b26c83fa
z73e703e4bcd2932b6335711c60c644067a80c1373acdfd557f5c4d7aeac35376b50d7cc7760000
z277d4c95254538a49d0a0193114173cac900f719d72a525d502081d48dc1a45e746f84cb105f90
z15243878b73f263b5bf8f99cd4ec9beffb8d6ca482cf34cb2973ccaaf48a8de293d1b90067eec6
zb3e01475ca6181ba24703d6c258dca0d02c27ee41fbedbfb872623127357871bb2f76c1685aca3
z21a994e9cda3d9fa168c9a8c8a5ba4d222b524f39dac5536175a52dd9bb39804b9ac9d01a1945e
z84968012c845b1b17b3fd9a5c29ae2fda32804fbdfea3d591e49c6dc85dbc08482c0de762ec0c2
z3770ef8456ed8e9360322c138b7c16b6bef579120f5579af9d9f0bb480851bcad1d3ea56d3ac4f
zdb0839f0f9c8add210dd8159a07ec872f6a3d147c9ed38a44036feaa7b60283de37f9ca55473e2
z1fe7563c44c629c45e7146203e4ee49f3727840a892eaf06052bb0dd8012b433e63c08e039876e
z547e83304337e7338c83b8269815fd849a40d76bcec23ae95a999955dff37b8ec732f0426b7328
z1877ea3dd6e65c800978bec72c6fba80cc38eb825642c0189de6753d901bd956f73c747a045ec0
zdb4dcd02173825918a713b15e52f119b4e703e1e0939b2c92999bd586e1b575ac9f15f7a20941d
z382e2a651549341320a905e069ec4c1a7e34cc42adf94c13b6e8cfbd09c151dc17c71a2bbc1b8e
z3da9c978575354d12b7204fa84b1c9e955035e3e0008909e71b9e0819b99f3f84da020a40724a9
zd6d693ff47b9788bcd572798a51e971c29cb1c06158e79458fe75b1bff8ee3171e43a532df85b2
zb1c394e4fba23814ce9fdb7215e3558d565a0f735796c42d6d785c025cfdafde08f6a74126afd8
z5b14f588c736289b89c6d8d8a569620252e5a15b9937c0f5d551be1fb4603da06c3ddb9ec2a288
z8776ac714077a2b538c5e8817f6d0ecda1c50098cd92fa447fd7a6ca21bb21edd7779a944c2255
zb9aa0a0691b3eba3d5ac285d1f05c2d1eb0950ee373a41da8c383f3ed7c5f9b79f7f50a4d2b2dc
z61a96ccd71d190c795c6cec0c82d3b3463cbd4502c97bc684e4cda8edf46e6385b46c98a9d1e47
zb8c9d5dc23d07e4a89a8da20d33325415fb955c02c68c707b20175a3de7bdc4bba98eaf8e92ce4
z622b9e988fa86df0b4271000dabd7ffb5d93fb054a3a9d0da423a732ade23946b67ab9cb7c3fc4
z8f372db0c216edd2c92214505247b618d782a11391344444dcac0dff373888e740c10c92bd2fa3
z138c1dddb68e94f8a4f6b5d935e3411fe0fd87cfab7a9e874105f00432571243373a7f6a60c258
z3a4d10d3c86cbaeb7d3fc140a397c82d198f3f1c7bd3d50725b03013d6dfcfa42f1d7c0f723b2b
zc1156ad386602987ce92cc972f8ff54a6002d193e3cad2a170f38e7fa92a05859da8069394b73a
za25e0a82702c25e39ed85c953f0cd974b92d0353b4f741c70a7576dfc74f425b9eaf1896428af4
z8bf7fb036b849e1df40df87eeed399b8acc2e25a5497f1619db8d44b1476a12e9d198ba0633d9f
z9c4802e280d4e17589b7dc0b1a569fa473b0e6152444b1fd16d6033200c3a6c199e89a3e02f19f
zed1d222ed9211af7bd6608aa2c580db91b6187115411c51664e3d74b8464526fdcedb5207909dd
z8bea745c55448f1bc5cac233390ecb360a86f9c61d99696c184c1a7769555d47f5f5b26951aada
ze66b64fcbd63f20281c05685303af571b62958322b07dfebc1fdcf3086de54e32dca3f19a3a891
z744ba8733485cddb7d646d89be572bf589cf53ccc4d4819d3b634d888ec73247ea20b3eab19f24
z3ec344a9906fe7457e770be9b6db53035a089b222b74e1d33bea9f00e4f17e891ca7262b2aab37
z0b284dce7a5e9d78ec86cbfa65a1917ccd5f07dd5b1d70e6dd3a87d379798026d6ae0ecdc6c22b
z4adf08974fcaadfd06c3104261bbdf9dd04479fd77705442919c832d4ca14ecf05f041cc24c473
z94b98dfb097c901dfbb8d3db11694fd87bd8c7376196a34a37b770d45055d120089591fb31ced5
z3f8d5b8b73c30f93dc0307886114a1d18d906248681af92b2c8893b9d4cff18c599fbf537de0f0
z7bd9c615e89a0b6cce74ba3033aa6c869e42f68da0a6efc280cb32a71134ff6b04c5bf2a409f1a
z6640f3be739063c781d90aa7d450e25db93a1108321a0a9e489abdd185ba9536e1fcde2e832413
za757007b4874b6e9f7a2db70d273e7622e0c23c7607a06210d688ce3d154abbd74f7165e612a3c
zfa674678599b8d5255cbc7a9c9bacf49f48c7c767fae7a8b7c17ed771d2f5b0439f543ad4fef01
z1604832647316755c3df2b691e352959f583419b6c95e21450a5375f2489f07f1e56546c57ba39
z331ce38469ef6873fc8843a2cc73d667599b178cfe771a76d6e37cf682ca4539e84103d19d6e80
zfb566e3f4f10bcdaec2de7a954a47ba7325cd666b44f19a3717be6852e3301643c1913e9c97a28
ze939ae53e15de156e06a2f3043d172bee1a0f4ba78afa886e1928571e5ef7170e78fbeba51d6b8
zf746d37dcabf9334a73286bc702e2e229762c4d5109563097f674a2c2a1978dd8bc3f9b958b89f
za1b1c9c19ea757dc55bd6be61dd3653c9ad6c15bcf324dabff8aa29a7986f7014c4756c085bf95
z0be80de7612c29a3fd708d8330471163c2b994e0a29acf3d71215a6579700823a6309541178b4d
zc127f64aa33d613cda08bd24ee2e865cde2e2691e6da62d988330eadd8f7c47912badc7ffb4380
z064b358e5faa8e238d18a213eb1f9e221ad23d6c602e8e1aebb54ab071beb6cacd24ca857d55c2
z335693a00746eb1cbcb5fef877e42e848735eeee053d534292d8c67c4615e03af28031904a205a
z1f48d1ee425c11a09c3470c62ba01695595f84b776dbdcb0bc612ff2469b3a318708a63986e437
z56bff9a03e3c79d23cbd16bcd31f71de4255ff11b5ef8a0504da05cbe8bb355c91c81f885b6071
z50b3a608884040a59822ce3b78b6d909787e00f78311c7c0d0cdf178d6360981b38406b26b7f18
z8dd0a22d8bc7b6b5a1c80aeb8d477077527ee117d045c33f9e917fa616ae7597efa0f216e4f1ee
z540faf3a559e5fa7980b167df79c6c3e48e97b091babc29c181f2548adac64c71245bf0863c9ab
zc951d8e7f2ece582a8826b5e86ac8ca6c8828a71dc277503a46b18ef1a50d8de728b55da0476fc
z434f73c66ad80c2dc9749570a1e40dec851494552317fcb9c0f71c2e25172702390e97d4ceba8f
z1e0f4264237c9a9373d6b595a4279145f63a3913c77a2300c2377b288bde2aef896cd384bf37f4
z4fc810155a22440fbe4079a61e89bb79606ec8bb5044cca468091bc543471b5e1ee418e1766303
z52df7198712606ad06226c6b23ad15781448b478602d32606cf6acdf71f88616b0970183462e7a
zbb76c858b26dead071ab4eaf508d1f3b2a94e0e238e4de22fe700c62c37106553d261ea6c93a94
z44e81dfffc936fc3b586d1428da5215bd1ccbff1ec2b18c526f3b553a1cef6aa35eb35fc9097cf
z79a6d582d2f31408a6d452570632b639c1ff6cb76a2a818673b039a8a4e6fb362afd36a6adc607
z82b2e20cf07e175abcf4f32287013e395e23bb76a22a3ab82a22eed05590ce92009c317593a882
z5df86744da261064557113bf2dae0c542b30382122d72b10e55c894220b4d55aec4032fe42f411
z2ae27b433a81568ae60568b2d59885f591261a077e02b04aa9ee9bae69aba5582e138bd7de78e6
zf24affaf48953447879805a21d56866bfcfc7b8c1f594fa7f0a2097c096f00b84bda7f5b3e4e9d
z5c680919a3872b2f39a2da91f47b2877380d0029d0258f1c9be88bf11513e85f012a4e3afa1d93
zca77acd1069b2a1d6678bfc046ff3cbd92a124173c6062f82925a81a09a44fb0a930e96986656c
z5976fc4495c0c1aedac7d275a146382977a7646776d7995d84e53431e5a37fe6747f7812053d09
z4ce8ea221bdeb79dbb5d199e597b9d2575aa5cc6c2bdcc9333705512fb9159745c05a91072c65e
zf8773ab32b6c076f577de196535ce70069bd26d2b5a5d338619f31f84c975e0dcf88cd63711b9a
z58a36aed061f603564377c19965f5d5fbe1f928aebd1557cf389704668210bfa24945a78727aea
z47ccf8433ca681eb347af8392f887db4ca80a51124a8824aafca9b86fd4a5dabc5449136e079c7
zb0ed2d4510f50322a00791a026bced84ff4c2ef52b1be66624eb47e3c859def1216933a7d1c422
z8ff6f6c6c1a121935332b324d57836ef84a18e3008ea014438dc9be20d3f5326a56a2067d17f0a
z5e909503b82a0bdab5d5ab528017325939efec4965828051ae9b4b2015120ca79ad5327c890c7d
z9dd9ca02f71dcdef1d54404eecf63190a0ee829c5c56776f78a7ed79d9ca80dbe759eaeb0d4f87
z063e3bcdae67cb4192eee86d595e04a7fe76f7a69f17d2c72ba8bb15140020a63da34a59b0db73
z7b74f4d0b685fcb6f7cc61d455ab2a6d481ef8f23c9f9345de99f33da08b7558868bf2c970e4a5
z1e555403b67f10dad8ca40ff8a0a87ccfa9bdc6c91f9fea75251db258f57f33e6bdee4530d0756
ze3cfdb52f5dc0cb69bcadce1df909572b5b7d29f7ddacae2a6f927fc8dfc1d3e99dbece3cb4a2a
zc1d4266c720afd158cfe553ae4acd64e3946930d47765eaa2cdf0f7c7cb2dede9628049ea19c86
z887da56733c595284b6442a78e2230e80ff382c9e480106de1a5fcc55e8f5794d99090166fdbd0
zd51cf50c1665d97fb1c5ef07b509b7339a38b2ba31fb25e81f586cd9c2b24f186d27ea6d40b5db
z95c55c9fe3d46df8a430c50f7d05a7b76a05a353720977bcb0a2ebf023fbd58f1f50580b816ed0
z53df264cac03007f947eb905594693eecd8c22da008cfcd3c60790ccaf77abe365bc7c40267d45
z99e5bd70b0a565b4d1253df81f8787ee4065c579d6ea993d50c156ab4aba55d7c33443eb5769bc
z66088a91d92c7aee93d262fb15a6f429983623bc9e04215d6ecf9ab180318d92dcc87fc00e23d8
z03ebb234e7d5e457da64e4bf3f79c050e6f2c767b547c9bc84020a55af0064048c5ca759a323ce
z8c0b24e2b109e7208e65d7640a1472d5aa435e75920bfb3104c124d9b0b2b39b500eac93b4e57a
zca6405cd4e5e1c516bda661943a389826f9ade3dafdd3e06f77881dcbb7c3182455ebe09648850
zb0976ff2b779c4a5eae6bd2e2b596612ab8d29913f106331637f4d8369dd6ad37a0abeff368fc4
z45ac37775f77c70ef3c82b32d696184a592caebb30dfb7203e31fc41bea773aa61b823754d2abf
za1d962765a8d55458a42ff7990022e12cdf1fc0c89c1ed90381e25be59686c405ebef7d4fd1cde
za548a8a74e93146765d1f10845bfdbac543288f4dcdf016cdb8d6fbb4e98c350be17dd71676fd6
zee8369038013be198751c3b976248f582e4e83b8b0c2818b8f6e4518729f37317de041d3a19b1b
z55e856f47a3f5b4ab6ca10c0634df9718aacd1a21cd15fa66f76c92741f9bdbb12ba44900af201
z5b85447c5ee3919a0e0a36fe8946998a680dfc0a93a7bfcf51a7c672a43b8348921c118f4c7d8d
z8787a57c83448b2bb8f2e1b082e88149a1bfb8fb7142437bbc476e54d90b18c6f4cdb236345704
z52faa891287321e79afcc0429d4da597bebae6d6fd08e843f5ae39bc87ca555e132da3a1268b69
z835ab6f52e76cddca5abb9fcd1a1fe884caa369f879ec55e8f919158e9f879c30777ab5cf3d735
za2656285ea7d67b28b58011949f636c88be20265518bee129919343b14926260f8ac9514e79b65
zec750efb97371366a530e37c928a817162aa0b545aa277c6e0d8bccebc5dda5e69e4af351876da
z382db304e33c21fe7f4194ff595e993a3642176846a7b4c166f6a77d2742caf9fc8a2b557cf19a
z189347ff83c2e2ffb3c9da1a1f1beab15452654076ac9601703ac86c85a06082a0773e04d69663
z0eac05aadfdb29e38cafefd6fa7bfd464a7692c406533fb122f429e3f1280707153da1b34bbee3
z3da390c36787f2bbbceaae4a71942b4d79dc789909f07c4915aebba36c1e213ae6de575a56d18e
zd8504068f8512064e26a2bbe632a85204fa570bddcec930d65f4e163d060beca5da60536ee2ae8
zc8e7f87196aab27336c487c24ecb5d69119e0608ea6e87dc00e8c0bcd205bac61f004d864de9a0
z4e5c65672395304f4e2a2253a0d9c956f851030c2981e62a2f3775b791559f8fd9274353c24719
z9970e76e8fe50875f38930678bf41806eb393aa0c94ec2f8a2feef1c97e7eb71a124935e3c1e98
z873ccc1762d80adf124342de3a1563dc1c2e927d2ca9172768fc99bb7602614fdf076685ab0a98
zf847f12a1c4be65ca7fb58d68977298f0a41d94166a60bdf543679e8e9d2621c8ae2725f2b1713
zb8253168edc6774ce9381e3fb8518317f204b8313951ad62e43ec238c5f4e1a7e3da5d678c3a34
zc600ba7b823ebd7e8897bd8811a0857cec482ae195978756647a4a5ad7bd3e19a348469307f1a4
zeb1a1e2422065222cda637343b4f11e80365e53aea506df5c315b9b8c3e189509bc5143368e16d
ze40eed5650b9b0f2dc44890e151a9be338abd2238cdea5a4f98f66ce0fda5d1be9a52a2108b517
z019a3061c3cef8ecb4c69c0288a16f32dde6ae985eb99d41492baa0e90411cef3d701fc91ae4e4
z8cba44e972f27c12444d143a4cd752aafe80c6bdc719100c10e7b67d4c27333dc70adb9e9fd801
zddf8e60ff29e7a6d6dad441e301111b5916211acfacde0ec6f4081e3a8c3a19d01cf6b78903944
z3cf235a4c13ff15879460c840222a834f0205b47155e44351bf86b79fa57a0aba15c9c52564cde
zf0faa9e90404ff5b40bdcd18939158d9fe07e067be452eb202914be7cd67bfb8550a744c7c36dd
zd490bbd73f6b56270f2b742e62b810b125d56beba625bc13e9a2923974b2df465fcfa5ebb6737e
z0937a472cb06b467d7814e4185f984724cac4939bfe7d53f22efe2204c4294166613595a324776
z82d7027a3cb64c652de923d175bedbc4cf1c23442c0311aa9747a6cb02ba1203003351edc756aa
z1330f917ebe71e64a10fb27785607046a7e280a65170c17e2a276c093666e53e9ddac46aba28da
z56cdc5523fe870fe876f25bde64d4311ffc7afb750eda7d196edd071c8e2c699e47af7000022df
z5e96dcf06691acf407fe46537a62f49990a677a33c2053730cc5462715403441c533d62df042ee
z2b2100a96e457012dc5efe6a58fa74dfcca34ac26f2193ba9882375c7b19a0b0aa0c8605c9b282
za13f455d240d58c4a4b0b78264b47a3ea600654223609790759063bf2c3737bdac9886642a07d6
z11086b4ac2bc9d3d74a8433de869d3efb41af7c87e10297faebe7b9999d456db3bf58d1998604f
zaea7a69f7f4daa0820f2d437188ac7bd737d74a4cfcc006a2c8a1afcfe6dff5f164efa5f7058af
z1e8c7297f9f255b4c9cb8f19ba62f12c8455f02f2d823be009e4dfeefd00541c06a160f1e90048
zc5ca341d4803dfaaad0dd2f71b7d28b5026bfa6b516a3489b0f38a24c2be6bbd845b210faffd7f
z9a215bf1ee05163f6e9b5e94af1e85fc6f4f063dae28c514546f5bcd31c19463d69570e80cab72
zeaab3043bb453f8c3d272998a0d4fe6cb6f767a15e20174f46a458f05830290b9d4d72a90b6d52
z8f1a3fd1ea3e49751e6c3854c371b437bbf5610dccb15aa050242b513a32ea243058c2b5427030
zbdd67df6c259d435c8caf8de79c1fab2e81bc3107f5f73bdd73c9856f9490bf205fab7f8ef620f
zddab7e17f312dd2d1e01dacd849fc36d31a6529e944b37e552b6d4eae7213637d625b91dd0a805
zda1625e2187fc3aa968ca232b12657c45e9f4b0f457658801ed801ae9f16cdcbae06f3044b9593
z4cda8948403c49befd18f4c2fcb5effff1eb8e6909bb76285e6d74f75d6500e8ee6851c183a087
z5ced93aed1336cf72e522dde3842f8ed3ad10901e3a2b070f12271c7f3c38a4e3a06d3cc85f7fa
z481c31d104d74fbc9295407fc0e01335ea6f6c5bf75dda5f6ba1c4b28b9f59c6811ffe472744a5
z89873c1a62a49f54c3003b4aaa58bb8af4abe3a81d86c8bdf333f78e5ecbf1f37b81c93c844dbc
z484d3a30444004fd40d462af5ca6933d06aead72f88218191206202742f3e1168905e265746668
z4c783f66afd19d054c870386a980a73caaab497f74f1fee8bb02b32c67db77cf9e87e83404e556
zdce1621d61c374c1a7439e09ae3331bc8692b72c994221d702d351368faf2b635eb302182a3c3c
z035104601b1951a0d4ba7be0d4a281cbba5b5ebe055e6a7f4e98849733a32bd1d56f1fbe2c326c
z068e244f9b2feba850f399b484b0c305483ce5fd04e10117cce92dac7f766972255fd55ceb5d26
z1242ef57e9a2b28eb754bfa4961252ebaeb0f6a78a0b3b28db9c70fa2a7739ed6dd17c6f78db22
zf3b48a40a2d6717bafc62ce54344ff40246972618d8769a0bb8f7ae28ed6b2f9bacb6188cf14ef
zc08e4dd1ed0df982373204a9556bb2f68b50bc80665cb61b0b905185af8d739ae800e5bec74e10
z8d2dc96f0a4fc0eeec6e397c2f87d1bfd5910221bfb7810d8a6b8cb19d99fc5ca38112d77f1e9e
z7d1c57791a3ab00088effab272853f05f27a967f0e88e86c169e983756c0debcbfee07a0073a14
z1d2ba0c4694ffdbb798da4a69a5cdfb454c9d99c0d57b46fdab6cff6617ae19a6b75a564e8671b
z7a8be484fda6835acc39478420b2b37ec08255b2070df625671dc002581b7558dd61b6bdaea297
z5c91b0f19512f22e3465eb6d9d86eb8cb8b67e4e00e34b033817fecb9d89f3ceb8e146bcd88221
z058e1d332e994129979026df37761f45a60d37b9395874e47acb8060457b2c708d6b3ff0b3fb62
z3028682f26a6dc780773e38c6ae437d77915cda977fc3484e070ed9ac3c47e8369667658868304
z89def2b8a90b196701445a244ba4e05ebe6ebb7f0d756e56b075f302e4259c6359a85d5f5f5de6
z004e67aa88f61e3aefb88c6235a69eb9b7cb84c070a9e2642975fc8fa89d6dc56acb8838217c92
z5b28dde3139501ddf674145042d8626ed582f0f637b04aed3da157f63780007966d5a9c4bd0f39
z621e35c8c6db9131947342354d418e2964d67a03390edc20279661b44e84ab96510cddc8da9279
z533e66eb35e33e983a929ee8f4a8783c885397fe16d4bcd360ed3ba8b1753566217d42d407bff5
z06ba774bb179629c672e1b29a8d9419c1d28e18438fa2fdd8d1f7caf78aa27054c1d7325ca1fb3
z93426e51dde45d35b230e14ff1b6383c7f877cc0bcbee26224127b3cec7b56a6ca7184c79889e8
zb5c3a08bff04257faef6f2856ecc568ec473091c30b038428fbf154425087e325d8f086f867da5
z799afeb95a7deac98798899476664a58cad3e389831fcf6b7a7ffa92128d0c07ac153de0bedf8b
z390d5195d13287781087f5620809f08ca7f4d945fd8705c7f0d91848df3455812a3b29f3533a05
z460f34d5900a52696ea131d79a9406af32dfc90a9c12d346497e15ecf688b66eb3c465689a7329
zbc571781f95cd610e78c9be6ad7c5fad1c1752dff46e00998f4d5868f2f8e033f2149a564144fa
z585703a445c480e4593a28dd5e44240d9f7b1088dff67a2d16c1be4ebafb9a8e3938327d743e58
z0d84f53290861c0127577a1c89f4e7efc39acc9c9607398f489e53dd0050ed963e9f00c66fc6b7
zc6b3e64d76c41f947e6f1ca962fd0c255b89f0011295a51ce46be83156369b4324a806fa21848c
zaae7064cfcf1b0a432c0a3312dd5f2005c08af40821b2d09aa7329fcbf7bf558e5dd433ea9a6e5
z6ac959d5aff83868eebd295709b915e95d067e6281ce8aa6806cbd39a61286b9be67670db83ff2
zb03ca374ff9fea5f11aae67055c27ae55db36a7ffec4b5e97cb42324e98f9885dca5b81f28c007
z2f41f23db2ecf7f7a3417c22cdc8debe729aa96da6fc84dba6560ccc584b712be7ef6e7256f17c
z6397084fb9c1ce78441a0ad21c9d65a2c9fccd3ac66e896ccf35354c17e4da8de8f46817c7125e
z8b4014de8e51a2e402869b1ac5e20163cc490ffc414ec33b7059db96c3f2bba01f1a87537b1bca
z37c4bf20084a2610f97c4453809074358da30e1b27b52a6cc0532b58e624554bb430ab4133cad4
zb663bfe38a312b6778be4be67ce30998ed80e45519d193fd031134528e0cce0b671c9648029d4b
zdfada532fa4fccfefb7cd2145b13f86273fb7a7553f34987e1cfaad1a76e416038cb44f52d75b8
z23601a7d2464b11eb7e125c1ce7b103c469f16f86b4ea091b8f1931bdbd52a15985829d7dcc013
zdada128c756316af431df933bc1e09b41be7039d095e764270f43b9f9ed9d4510015cbb9ba4349
z172defc36faeeebf7ab9c9d8e422664b0b69e08ca02454fc0facba7c5f5e1ea68c37f01d55d2ff
z292b387de302ccf1cc9b7e819517cd9b57dd16ac9fdcd9d6d6ab5a25bf88b07cd937a46d8566be
za100fa82bb42c1c61e4d97a30a5270060ec758f7ecb8c72d84a2ac1aa52e733904c5307bb6b79c
z27dd795526f05d074b55ede60d9aac1fc0e71156734a3e065ed8b8352856a30cdda72a67a8d19f
z537435696be68f2cb4d11d05d544df0946486e11c9ee08f3f1240cc05cee77f379581e02c15e51
z0b49df11966d1261c6ff942c6fe3d58eb58f365a059c8263a05f7b7414925d80d2d0cbab5265f8
z38296fe4031a7b0ce867ceed842e02ecd248505e5ab3e3e6a6773e3da52d048f9a1583d90d2e13
z361287250156ca03d0cfb73fb49f0136115a5a37c52f6de728aef197f71bbd9aaba92515e4e708
z63dfe507deedd5580e013ace36afc25eed362e6dd513d3d16544fa2252ba90ed944191e8e28267
zda4aeefb1164667100f41f3d2bb16e41864dbbe8f48d22481f58e3ef36462dd437781248833615
z3b136b058c9bfecb4a4e55fd020a9e9a08827f7f2b61487fb289e22efb558cdef787d84fcf4bac
z2c8dcecf0137dc01586af5686d0f7c8ea5b51a061ec8826ee147e08061b78e2a551e63e3036b9a
z6eb0ba0aff1800b19b254cf8e517d6ee446fd32d9a4c690a999303763c6500f9a7dff6aa43f1d4
z54926b57b7946aeae9d3dbdf11b773961c0dc8016b493936bf93f9e642baf7653d708833aaf833
z1c489d8793559d1875f23741e3ca5302ec4ec1c68389de3da596a268c09aa8cb316b52301eeeab
za9dfebbda54144aabc8c1470b836ab6de0a8b0f270c9c449b050619c8d4f7bcaeedd87e6718a35
z5b0dd70e55d2e72422eaf25b3b6685c7adfce964c559f568e612d94c595a55557187485f1890ba
za8127acc47cad55a1b661da58334317411b490700ec5afe7f00acaaa98adf4ce0bbca63a09b298
z7b61fc730662c406e41766de9bbc2cfeee6f45f9e067f417e50a9937ee1eab2c0ab6a00a3b21c9
z115029ea6a03c72c636a6aec22a9277008d2bace082f2cf08b5e0a851c00fb332912ecf9ae6aa3
z71875be5bcde6deaadb862b5e7f72d70ed3e7b6d5f49b15e686e019947ad033aff3d22b7714e43
zb83393946bb8a4c127640e464d6af07127d39f1e28071015fce5b88f8b8a1d1c8e57cfd8838ba3
zb552fedc2f3e9d8a9d176215011bd8c51353e95e26417b30ded8df5812c19e43ab4726e92f0d01
z89237e6f115068d4116d2a5a25244deb77e1031df3e64218d5e913769819d45047c16d1cdd7fd6
zb8b9f07476669436d21d61a790f4fe916cbbe2112154196d322fc107bad01f9b4160824a7813aa
z6abf5c52618ba69250cf6d2ab4b6db82f91ff0e749ccf22206fcf51329db279a2cfe66e40daa42
zf68f7449aa0e1ce26eef29a0046cca77253bd7904792884fe593a8af5ba1b27b5227b2131a7a65
z5aa29d339789621abff16793dd2f08770547e723726233e86d101c6891a5a3152718dc726f93a1
z2583fee1e89db02aefe5e74e867661825d2579d64886a6c7b4263ec2485adf32eb0aa90b59ab8d
zb947efeee10717a8756c61e0a503bcb9be58df6541cff899ec1f216339b7d97970838b65824d1b
z9c9cd4fb405b57f5251431f3e7c742c95dc285193f56f90ea5e90a44f53207d83635e9d49163d7
z83e0e6f430a4914b7d3000294d3019a4d4d2d130ffd690ba651eccf7110a07b1c5860260915528
zecbe60e5a77d2db3a54c4893323de981744a4fb1c97ca25271a95ace8004b06d7d9bec76469efe
z026ba83d75aa3a4f011a06628873fa0b6a0f3ee4ed2f4542128f84a87d12f286cebc0359032d3c
z1c06fdd11540cfd28b593ec9b9ecf58e42f688eedbd1242b6663291ffc92de6b90d560941f9df7
zc7d5d451f70679977f80dd90c4cde8f1692641ee504967d35625cc41d2e49b63e48db339e571ec
zbb0b2c23419e43e595136cf02e4d2b4ff0c292edfc158a1523e9c7463c2fe4be8190eaaca78a61
z23a5c142ccb96e9202f3d608138f1a8d452ae9e1b062a2041813e8f17369f721c85fd84124798c
z11c19a3f0e8501572813793443c012b97bccc6a9a9b301e5b2e136951f2e92f1fd803259fcf28f
z7cad6db123fe5676cf8d86a09971574c08256a2eebc9faf262549de3569ac9cf1deb799c5dac57
z7cf92bbb043e666d3bdfe635af3c41e8370833cf7eb206828f5be4005537982f1da6cdf72ca7d0
z6ba9354401c1b639e964f4b53a44aa76cf6ab27a6bf1c3ab0f4eb1f24b6e62360a41ac91ae7888
zadc3a9fa74db92f8db188d9f97a0449dbcc3cf83d09d554694f51eb0defd0137a587050ca1b557
z0e7bf6bf6a38eea220bc33ba55728ebd11a6517eb8bb9e1c6cda675666b6a24fb1e6754386c74a
z56129f920109ea1b7c544c6134ef667ddb6c38478c164d0e546f5b583f21e308eb4baf2fb68bc6
z5fc99c995689dce9fd40e33225055f2baddd70bbfb1f7d520f20c3996d69f9315f78ec2de10fba
z537906ef057cbe25540f1858e7f3ed1ee14e3fb4f719fb2b6a35657bbb5aff35b2e2788f2a0919
z4c0a4d345c9403d01379c3490fba545d48af8c91d50c1c6e02b0f1692868a8e8ea08a6831d5d93
z4b63c82b0aefa58b94ad40d1afecf5f2a0a39c7b03f03dff32407047f3905b688014a0511f6605
z054f3a8927fe12cbdfb2dffe5f304b560518e85617d132fb3ef2a1e842ee90a92981e3b368fc2b
zf85f860e2af8afab4eac767b52a75c08e78718296408409927f09e8663c5407a75bba3b3629365
z920a477a1907f4a4dacdfb4480449b2a1d85a3d4304676b8448c64f073b8e0d54f01a5248153b3
z7f4897c347175ecb409ab18704eb837edf5c14c64cf4a34adc6dfca1a70b7024ab0384d18f842e
z03eec3888b1e2e33c8045ec5559b7adbf75c02911cd3398b1188b2f1836f6a9074a7f5f727a219
z432560fcc0cdb783f8f71e6e56ab15d3c07abaacf795267c843f52dcee0c76e07d21e40da28cf6
zad082042868f82803e9123b4a5a63790115ffcad5fe5559302d3d0fd6311a4117d614eecec8498
z6ff608e7834e17d2a2fda41b1a6dcf6182c2641eda4922a9bff8f308e8ee873e7852dc6d07cb99
zf61e1f5435c2b7a43ce88d8fca25a8a89ed64bca39a1b938366b4a625bf9de410cee641bde3564
z968180dcbda0816687cbe7ee4bfdc5908a9b64459f9b3fe0e01ac5a6f993be1b718a1d53058eca
z7dc1a2707c7e6018355f05396b2dff7040e462096a4c9ff8245538b389744c2c7ab7404ae4656a
z629dd115d0012a048bc063f26ab36097d2b5992b23d06c2d3605122f3b0cdd939fe286ec41001a
z745a6730297b0692b729fe2742c1a07df736155596815ecc546b001f9c6090ccdf9352ecf2c66f
zead730f7e08aa2c2012aec2d275695e2e4faf5554991e51aae9da2c0fe59c21c2ad2534b0c1875
z64aefb67edb916704885edaf69443253c367646271089a67b3f61c4a4911547f4a7d4a9217288d
zf0d8b88f2d6e0bf242dad7ee87ccd38e165223f7ff111c1c9ee2e246c7702f1a5fe5ddd0c1d566
za3c805723e94a618e032a9c64a07476eee6a236337257b91f3501294623d5721eee27747254bcf
z964f3908089435fd30f1d32eea743634fbc2152b0e14229c4e41bb60dd11c3f9183d947fc1be92
zb33cda5f64f4383aca6994b55acf0a84e8045f0307e5a38b2b557b1614f3c95697511cd10c2404
z6e6934cc64216966c33bf1712383c1a99e85ab83fdbecca08289e624f70ffa7ab819cbe94b4a2a
zf74d9afa3c689ece3e767974e70189727c8587ad785c47d2b69e21abbf1a7847cb27a4be6e6b94
za691ac38dc652ccadbbed6ae608acd428ab381a878963aaa83994172d171c6187e7d99d2e432d1
za4fa454ac474215b068b1b697496d438e1591d1e64417a31dbeaecde20a74401da2166762c8bc3
z301db0a2fd174067da2c5b0c5eed92ca89a541664c0d61d3d3b37f28e74f9a0cc2cd81c575cf6b
z1586a799cc586110b0989e21d64f83698d01dd5a11dea2c1133b7b5e9ea8e98d17ad7b9d1864e5
zdd3544fe36c506a381ff61087df50e6eb2f7f5aa8aaaa97324f145393894faa6f5093bf88a35fa
zbe71fe27c06a1448597508982dbf50127a8d53bb20ebf372ebab4bec97e916888d69bbfaac4462
zb8d616ce424c4b2d8fb17b8f6e4504daa21ebdade28bdb84d80d71a2b8619e78e7d04c850c6362
ze4e0b6944be4366041b09e28e7288ba38772f5e2978b8bf4e9b4246846af6bfe1eb5a523220e19
z3021e51e56f1feed9ecde2289e4c8329dd105e3d2bcccc1e8f2b4ebe813c77ab6009e515f1ca18
z643ca5302e0056ec21a207b115e39a0ddd1e4a04bec5bf3d12d4354b8a5607dd16f461cb731208
z1aee154c8a6ea42daefca7f5c4f236d5a140aaf97a881d4a38190a5e4670d02b1f99506756c65a
z09795de9288f74a8ef893375209ef70517b2322148bda4e0149ebf6ac4feffa5397b58c4249cf7
za19601ef004370dd8074933b1cbf529820890ce307600b40c0916dcdddd51655adbed1e6a540c9
z9e5ab725712f61d5032f44b49c3c16804641d607f379045609dea1cd53f8814dc89397659279e4
z95116f961b3f68cf5cb88c32303027469b319e3e015c1c1b2e81d46468c9aed7bcada13e4aa674
z4e2543264e567f9d39de04124a7acc115521e0ad158e322c24f41ed3d635160a4ac9720248bf29
zf8769bae472e25c41c8b6b6cb538cc16fc87b11ac5a6859711d90f6e586a001113ff4d611dbbca
z70d24de3f2baa656295d2b7b7ae1fe2fbb68a41f811839b2b16a122e3c5e7a7e7598cf0b716b4d
z7aca437c189fb99196c041511bfc3862ec5e109ee152d1c6c1c6aa87c697e7f68e3bce60c21190
z026e93a06f614d63bcb010d29894726720427144aba1a15bd8e81670e013cc539ed7bdec6747ef
z9b11d04e2bff8e492289f4cfde7b584d1cd8a58413318414c021e3f0edc464e0e11d7fb8bc6ab9
za6bdfebb532ac3bf7b74b249acadf278227a884b42a0d7cc8d679c0b3bb6fb5fc9ab3080090e46
z14183472eb9a2152c22ca50bc3aa8b096d8da0eb5f5ab4e9f852c52fec4507090f41136bcf0e29
z7c9ea4c57b2683a43faa852e9a2d2d36894323ff77d0e7737c3af7a588159b20306f2d1d2a17bf
zc15fb3441488cc911eae36371134c111b0174585ab33900a14f996db570595bec3a29499e743d5
z7900e017be0d182efb959d5e14a58ef585345985f59ece4f05bf150a4749bdbe470b87502151fe
z4d7785903dd692447708fe795eec524917e8f4ce03e5d5618406693dfe0db18582d8b272e36268
zec86f9d2386455c16668733bcc9c8e2aa84cc87ff45d9e4a611e0f0097dc3bc8f31e1da820ec42
z16770af55ab78548a61fd028d37bbac940fa8ffa1aa730243bfe744bf0319ba51a833acdf9f534
z775fd8b1a4e079b251831ea1b5f5a2f513127e37f9adb6b92f1ad8961f1bb56dd8560ea1f04cab
z3fdbbf9a706531b9d8fd79ab66a385303cf28cc0f3ec6cb85d0a4e4168c146f1735812f706fc3e
z06d4699e4ca7ebfc37edd3526841d7bcdf36e7aba0bc2670277efad4eb4ccbd99627fef9c929c9
zb6c5d8dd242d47b588c6970390848434f8a451b8a71066335ecd2880bd781e3396e1dd956aa20b
z0c4e0df7933918466441c2aeaccdb70dea70332e44ce13bad634c734fd4907730c6566b6a28f8f
zffcdd8ed7cc0894db80955f1f4f47e8ea198e0248fe0cd5a732bd01c5c1563832827cad5914b5c
za50d8ee0377c13be1d256ec405e06e8dffe3d51e0d3b4f2226931749fc1d2cfcaa90d1462f9673
z8ab70f540993536e594e16be3d8799f2197c400c762e418c376478ff6ae821f21623c318ac3b29
zbad55348caf1d819cfef9977f8b21c1760efae76cf80e05b7e74deb9ba22dd2226837898d15b73
ze4ebcc62dfaeb06bc02786cd467f335080412dc9384deffb7d28ff718817195ca7f98dd3e62499
zaaf298a7d982835107bce0806d410633ade392507868922d7f8149b6bef25b085dbeda5d8fa789
za5ca0e453c7638f78a1e27c216d931127e06dbac8b3610a80c17cf0a786002eee84bfc98a5a222
za88fd7bc9fe033e825b697df292b2a124572b055969f3f19f7987d93db4609f3dd7483df73c61d
z22d9f3e44501541396eea358aecad3d29fec9a2fd794d68fc7f58b12faeba34ffd7bc2fdd7b3cc
z5bdac4a7431c114527e267726a0987a5fb353a5b359b3c9804c42d4258a378d676a98179ff640b
z772c84c78a2b9f7065cbe1ce7880cd0e1e684072cc24c81ee57f0b9e6017781c0fd972b80b91a8
z3d448dcbc837f2b6029f73a6ce069a7e61ae51301027ae0033fb4034e5c77886e658a4d994debe
z3ba10dbe2d196865c279feb2d492cdd5284ab719e7fa22054c3ca205044e72195bfb2311244de1
zab020c7816c5411c9873041529df964c7a8476f45bc758fccd853f5071d4d831e93341c362816d
z3dc76041894adb1bf8c598476c1d28f910ea546681bbf03b0541eeef601219321aa7adb35a361e
zb2f19f44ce9e5e6746e456b009186d7c2191fc6bdfc0f0919b78770b237345c94c09f62a1d08f3
zb4cc86f923e2e0cd45071fbde9807e238ec9ef7fea784c4384e1fffde370d72a36b3c463a3e82a
z145a97ed6bd4aeb8f767a58d64deb84bcd58240179f21fdce3c58b0c057b7241c11768b799f0c4
zebc94184952796a39f897decd34fae7b9446b9517ad28ab4f22e1b0e4f89470f4d1cd8176d85e4
z5de2b308317b6bcb57d8f05a5639d388f577285bc608ddedfa72ba8355434e2ed927fd04d63904
z84f04cebcb7a2a7f067c8b24025bb9d2e1294d7a2c47dd4fd61f216005d614fb8f9ff66f435c92
z38c34e5e7ebf3220403e056c186d7ce71c2133d779e5548f02496e13dbee03a88dabe896fba57e
z84d890fc10d2c7e260506d5dee5e879dc3a27f2fa5522eb947f25618d909aa1d2164fe510b2c12
zdd32d6ba6dd417fd228007be71f92cc69596c73be872e0faf1517c5f2004ec249624982583fef1
z9f9810b1493c7364bbadd5de4abc41f25e21c47e47aec75c3ea226ac77acddb35d11a8145e30bc
z64772cb5e84cee9e8ca2d232b3ca29cf314736e9da5222d4d23b67b847b835bcde966a098e6318
z1c29ff185e8606588e7c7776041417aa4817376acf9b53ed1b122ee4b0828ca4875c649bb3b410
zab61b97b4abe20439b3073bec80694c269dceb92d0aa37ce080735fca38468a2260f6211a55612
zca26038c4db267cef593f442576a6a2db5232c14407ce6bc1f1682734a98415707da95521cddac
z506fe70ca24833f05c57bd9cf144eb8b5571e5f29a1b170a8a62a4a1e12d62c6a5bf8afb4e5349
z09714566be619c2335b792a8b38ecd682b4248d83bafee8b0cf3592021a67034f175f967f1afaf
zf695d59afab683378f0b005adf1a12cd033c04102d71c076e9943e41eb3790fe6385f35ff52199
z623be893391a2604d090d93d450e26cae3fcbd6fc7ca170c0d7274aec0d82827450cb202a0a414
z2bc0442854af7a9831c03e7a51b6b5d1d8b4de096813f4b7f610476d89c758567302e4fff98599
zf5f5aad9fe58907015ec3024f7a347ddb192c551517d2d4cce7157d90378759566ca1cf042ad1f
z452cb49b1da4ae468814066efecf8f261f31bc2f3e720341ec4da24ba6ccb3354eb1f484de14f3
z54c83514d12a5ab05d21e5fed985608bcf458e672bbc0a8b4948667c7aaa90fdd7260e81f8a6a9
zc57936e95e49cae105d6eb64e5cc79934ab695b9108cb436d424eb328e6e71e09fd47585169e6c
zbca607eb58adc3682de421b7b495779b91da030cd42641155aff0cd71b7b17507fd85b272fcbe9
zf531630084d92139033377f9ee76a64bb4c3abb55d9b4a274431304644ba2eb5077a594268e5bf
z060fb3942a1a48cc8906e7c40b396579943c1125e4ce13f9d00ba3c65c13ad1058118e825bd3cc
zd489c1b64d0015fa8b808f8db69e1a1f623fa940ba75d92071c72f928a7c90aaf2e85d09bb28e1
zfdf156b46b471ef31566f2db19cf881088f25d538ccd99b30bc0f57c7698c33a41c3732864b90e
z2e615c89c06861783342e7c5fd35622da2f2762bc3b10ef76f6533d2a28fa97bf0f3b597e99dbd
z1fe2fc36411da5c85f4461a85ebd759f3589f2d00d3eddbdfb47a100f829618383ecddffe69992
z96c7b94c3830ecfbcb52d6f73089556e33b0aef9f8e0be5e2b4c53702d4e7617f08faade2ccfd1
zda37537816ebb6d0172df806364eba337bb3590eaecf336b7abbbe639f0c778d19529b90f4adb1
z9d2c1d7f862f2ec7a19dc1a5cfd366f1888800ee7476e7d09aff5f9bbd3f2fcbb163ed8b4feb41
zb8d289552fb3d172781d79f20a4edcc9283156f7ee79e057f1c24426b5201c2e9f105ed85bd44a
za40bac8765481763b588fef99f876a0c88b4e93f47f3613be075a6cab77c4a16400d547c9cf5d1
zcd03521c2988a214dd5df90aff87e1c80da0b8f3535a073dcc9a42632b74c7c6ea84cd2e878449
za384d5c64e2e1b62b206802d69201ff4c8224d8a509d7355d1edc4d6ea89c064c72d576a397508
z15448ed46b9780a7a07f120cafe2ea607e84238cf83c243cdebbce15d8c044634463ba65cff70a
z4343640acdc236066a486b20dae6cb8430dfc84c210039ab15033ed8e58979d89063f6af410572
z1a34314702e8c853c1049f2917bac7c8f265dfabd2b6029161654c0624191d19af2d5d8596e32b
z1b32f164ba84e40d3f6902deaed8360c2178119e9ce608f8aff39e4935c4c4fa9da731368b5cc2
zd0e978bd781dc6be8268b546205fb8e482d327a274c32021c310dbbcf1dca1ee02fdf3dd9198a5
za67f847e3328581f05b8207659e2aa560c46c14e46befd0ff520d52ffb50da10e816899d745c73
z9c6cb12e4687d4ee0b931e32aea2790f7dd2a8a3135d7c58badd248d271e969fa8a5ba87b2ace4
zb7a3950d28e5732e9d4e489b79b2af32ee740cfc6f2f064ae3d25d4cba2607a64db534d5c2f036
zf7af75eaa0457ba2bafd5623447aab4ebe4d70d30d576e39e8f90867aa7a49f094092a1be78953
z2a6c9c7984db784e437eede3d1743f7f66063066c7f219960935167c1c93ca34ee9f85e56cf5f8
z23fad43e9acaa59bf9cc97baa709090a63d7480056d9221d4d8ed9c4ef93f4d41d73d434fd3149
z8c810c70f7cad9aaba747d22cb2168feb2a172224b3491659d15c0ff22aee17f2c3edf40efa699
z0f00571901bc99241715ce66123f428673f9a2fcc86be1aeb35d534bbf5a917bb76ee6eae5f897
ze4f79abee690e3d0aa39430cf3503f852c5b623980ecabac8a022876de26c13f7d7011b8196b0d
z89e059eb31bdcc5aabf464ea82dc4c02515c933c0be75c6a04d7573d1f18eedd0249802d52aa53
z35302a7cdf2a734a4e593a7b27f39e1e597dd4fd34107136b4109e50254196daf9a1838cec12d7
z50bb757185c3229ca1ba0cfd568aa3bb3604dde3987d579add775b30652a4313c4287f5c5c2f27
z97b56c00f9f03ffe73be3f7c2d107e6c6f37e725c4de20e2d143d659aebfe87e8c697fc6fdea53
z0dd84b34af7ae144f2c060a9e90041bdde1d90a48038f5862652c95dfd279c191b084705a27ce7
z5c2fb23bd4f0d5311e0911f5fa31c58c8011ef3a306459e7b686b16d33e5e00d696e8f7214eba2
z33db7ace61bccb1033cefbc99cf451a9862f66785a63860f1c75098ada59c9ad49a2b4474eef48
z74472d51235545558436920fa4efa371ab5fb778616d58c32143b4c6a54f973bc40a917dfbc758
zc55c024b476dec12e427184f327246c13d76daaa6729f0ef69f2f3e105b652ff4aa3059a428890
zf43f0d9a73a9ce3e54e220d9b7e2dc4474da792b7dec6ab44564d1addbcf8d220c3e56273b7528
z2a056144b4f1885b9d1b39498a1ba7b05186636fca925a741c3c6ba5a3b8ff165bb5b45c3c8820
z98b118a340999680862dc5feb53fa35e6e93de7d594b0ac84bf9e7ecde3d8e781affcc303b89c3
z6abba6d5506a78be941be64eade73bc277a69e7256c1925479429bdf3687a72f875bf3e0d25b57
z0bdea62325acb05e91221d2261f170f8ef01ca595a3a46e8b455f65babc0997e4c9d993ea575cb
z9ca6f544993548e779be2844d0cd68ab9fe52f3064cf5e974a9060039be254b9187d99487544fe
zf74197f38e4c567f8d18a3728e4605952446694d14ad5c94440d8dc5300b43cf936d5929499e3e
z2c64f632c47d2da24f3ecbf23dff1e2f5274013be148e25a5d01a193f9112d556900d8df7f64ae
zba931b4c777b3a87218b40ec27efc10dd20d19712c688d00bb27233b79d4f0d8637592f4e1abd7
z6d259c7546c9009cc6d901748f826217e4d81f8e3781f4b17ee004d292ccb3a1f39efd2a2df836
z877f297824a20c1e848c3bf73ec98f3e8058dd58379ecddecf8c9c4f8bd50dd6bb8c5262826ecd
z3390d8c035cab65de2e8109c2aa0305fc61b5692148148aeb3f34712134a1db51dee9798dc2730
z7153241efecfa90e08efe07d215a9fd88ef7d44adf833ea315ec65c04bc3e3645b6adaff7cb357
z35d7d1b886b808f81317c9bde1617ac23ad5446fc3a4e3d51d5cccead1b9dd24f1c2c026c47142
zbb388035cd48e9749e9d6dd7c452583551e104de5be91795d6811785a9cea8220e7b8efc887729
z475fcd3cd36012d6965314535dd142c1a8b9ed70c76f84ee59682819a567b332886d154b8990de
zcc0829a5f3abb325eca02ca5f8893390ff44077577519cb55094e53e65b5ddca49d5425ebc24cc
zd39c0a330e84595475689e6c3850702d32360ebff7333239a5a77720feafc81b8262f81b2b91d9
z4b5e731e41933f66cbaa6f8a63933a632898a99636e2090a49357559ff86511a4a5f6772135baf
zd8e5808854717067bbad6218608374d80f99b2ddc23bd358ed9b6ad710484d47e9eab34e9c44d2
z90e6f5cc02ae1592c19556a27abb3581eeba3703cef3c38edf86e4801ab9d9fdf3e3cf773ef2f2
z95b9ab28811b6da02b4a46d60c5897dccab87d262df22b61561e620861e130777d3f9ca3ab1410
z29a7d770f5d2ac6d7b62d02c0461f020b58945c75a03094033d4a9cba9841446b9c1c5855115e5
z8aacdd86126ba3c1a525960b9bfcebb08b5da022c3b9378d0229a4c39c13bb93dabc4041e986e4
zb8176c57a0ed9332f8fac4e96ec91905e5430c55dae368ca9a0d638774841ee20f2c50eff9be8b
zea40da41bafefc59c12128bbf7b25f17c5f85612d4f954d90a8cb79ca551846947c33380faf03c
z51b3f63a63c64e271cbfaaac48a978c4b359c23106f9ebd68ffd47b3166bbbad099a08c586b5eb
z04913ff9e57d8bb69d8fc299e94af683b9627df57f2a0da32c83a71d2067db333fc7ecf67c7b41
z95bd88fe750a769af8575fc5fea70665ea145a0375bc947a3b0c7e1d4784ac2ff2cd886b9f52a6
zc1bb86557548d383890005fd2f2ad98c8004d0d3de612d7ce90c2c59a843b295587636c17a3b6d
z13d2e7da5979d6e9d1cb6ada6c010c915889a6acaf65b9944bd00bd66eae1900712aee4691440f
z5143e8e99e1f4231b391072f5a98a62cad24a1dacae8dc5c8bf1836d0991d92ce3df4ea7b7b9dd
z7d4dbef0f146be93f162565d3773c1a9109f843d57c8648aab992858c73a2c11c7fcb1ae9412da
zb7c4210de14b66217dde1ed1eb9eb5f93ebd2ede783ce02dfa51bf3d78a3771b74e0c3c7b1b1f3
z3da2f6a1b449cb6a5256e63081cfb7b4193497c80e5abef349a55fbdbc1ea454e1a10b2257ed43
zbc00f40f68b13e5b0f9f2bedefa8a9184078a7c9afbcb4adc9b62b1f84d5508b9c37f44e11398a
z4a5a8faa5d5b3e9d4d0cfb29225f608495132e3da4be3314aa64c121c97cccde28069e11b3bea9
z269d47c589f35b01f0266144b3178313267dad624433ea5664af85d6cdfa3eb281e96e12a566ea
z07e13baa73718526cae753434836d7a732139d4fd65f4aeb280de2229ec73121711b6fd446e14c
z19bf6aabdfb8c151f1e4aa840dc87ee64856bd6f02110f751c7faa91117236bc3b56cf963eb144
z7990b7a5128e8f580df6dba2e6b761bf475e8efa575e3cc81c093f5bf00d71659e0a6fd79b2553
z5df5cbea3a918c4c1d875fac55cea2109c5d2519d7a160444dfbe985338a94b65f84f893241853
z32b46d816fae4f914eed849c6969eab078ad3fd534a09b2091800cb9d1fed32f40b7b65503bd4c
z215504c124a067efe47b18666c4b9504be5580d7e53986c3674c353c23d5ab4c06cd0e28ddf41e
z11db948de7e96195c463e06d9964e2325dcb42517e7fe15e5dc375954737dc9e6c20a8cfa7e4f4
z13c5db804e4c6f05c52b6dc0ba735228c8c88e9f051cf852278b9a060a58775c5d8d9ed2ff378a
z972a9db06e72a8c76519c77391210b62b071ba48faad0a9d6da04be22704aa0dddccd1d647b131
zf3c76eb47063471e7d1b92887abed186727569535d250d5c4f5531e2ec3819dc39192f61dde68e
zbaed6dc3e9f5fac085661115bcdf63447dfc5c501d529eb29f30374f474ee8fdd4d736b1c5d4e9
zd173409dd3e946badbef202b07f193f6de2ab17f5fb2d7043a5573a2df2a8c8c726f1af7c4cf4a
z755d4e54e31115151cb0c3b7d23b8b25a50771f09227caead2b1b226f01da4159b0a95dc83073a
z327be85fdd8997ca4f19b5e69b48c003fc380c300a3916218ee616d72ae7df3f22210c8b76dee4
z4233c79ac2663a36e6b599217441732470a969860c2129483166c47692a111a834071180b60b9c
za376cb047cf22b9ea5d83e89edc3a2f85a423ec96df098c05d2d0efb02338f05c1b36fb378f10e
z636401df7e1bb64cc907b565c14d3b605e73aa667e449071b70f25d5451253f6234ba56bc03c93
z72feacac664ca7d57df7a6fb18dc02c88136279766195aff3f869f6947f2c20b32dbc97ccef385
z7709d9e9714bdf2d51e9f57876bdaa379b034b7d806128f847cb81dfd3455a7ee9e49a78dc88ab
zeb9dcad3cdcba1b767baadca40e97a2cf3cece950ebc802efad4ccfc29989e2e1f9e4dc6d150b0
z79d6e4009628f347eeda6b5604fbe995d69e573e10946d20457333accc835f08f4eb4c16ab810c
z200f7d6366fff96d3dea7ac3394f737f5181419874ed39edc575cceeb914e224ec25490fbbf864
z5e631776464f5d7ca1af2d148066de72f8be1a8ca48e170f26b4a7df82e3283ee4e6e99e4c9a2a
z72c0b4a514a930cf71c5ab6baf053dfdd07eacb581b56973dfe8735c8651255e4c19fb39d62520
ze71c0ff2a1dd911e867e30e21e315ba75bbd39859d47014edc644975b62e2d56d4bd673ebd0445
z4e90941605eb8abead07f115bc34183bc558260e4dcb8bee35d110317e161dc6f5d7b27cb88e21
z39febd4ec546f2cd64dc08638c38332446db85f89c8a05b7686e4187d5a7fbcab6e018d6d4990a
z63d7a6f57e9d3b288a7392faddd630ad7c07a25169653a834df6d6a0caaf74dced6bf27bcde5ab
zce03269962a2d1f2a59245ca6b96350d5e77f89cdd40b785df872dd7976c4eae2b8d9bad5495fe
z270c4f08ec68e8d77b54ca9fca69ea2f5e3acad867723ce732c2d9512d41f526328ddae7c2592e
z8cac1964d3baaca353fbe8d168ca29f2d9d74827d7f8ae19ebef0a3dd7cb5ec845d6a503d13871
z5a1f8a84f43e1d940514604493925dc3748d3b928b3f7d4fc5f28b5ccaa7fda7aee0326fa3babc
za2e28c3491401e3691d74861fb8861174cca8d461969dfe889320ca642bbbac4bc6c0dd2a36d5c
z8b0c48017c3bdf889d3c01aff835db3bc26de30bb6427727702edd4b0c95167f52e22caa60693e
z48f80aa62d77f003ac4f937d766713362b3cf71fe7ae62550f08cde635d295f5c00fbec2beab49
z094d899e32bed0250f13b76140daa60a531cd1756c87c3caaf1542609a180105fcc78893a16b2a
z0bca9ea15431825a7d4b88ac370fb319d92d16eaeeac7ddb1392101774e915a9fd23dfa5240128
z2a2337449b2c65b4af8bd95ce3c519c56069d6d461496751b8078bc8916c4262212d84893d1294
z58a406ba406a7399382cf43f48c920d36774e3d782869bdf8ad8cb821f65ecacfa33e77aa75893
z269f68507212790f839255b133e6d4c5da618b5e1a00c708da863cd3b3191646b942ab52379aa9
za9c6b4ce0dcda8a091b8a1abd08b06dae27faaa89c1555efd02a6d876921aa23c2db7af7e951c0
zfce0304564b4f6f163137c1c78edc46b471a4cb4cac3ee94d3f0e151e76b8fa2aeb07162714e81
z39430bd609845022634d0763c4cf966dddff8f323abb46b0fefc7c9bd2a5c982b465cbf5523b6e
z352c22104e0ab509c9172c09eda974ddc711d8c6bf11e75421d6dd6cb3427ea178725c152e5f8d
zbd4f38322eb13cd266e36ed5e62e0703baa6517d1663ad640cf08202e469882dc5c5ebf130dd98
zc6d701627ee018e28c654c8f820fac26333ea1b8fa33f4dc537474b0e38dafb2fd4eaeea696425
ze363186ac2049ab555120a1e8ed68685328dbc70c1145a07ab27f3ab817d473a1fb1959d21f6b8
z1d7549915c9862833dbaaa54060e3aa1bfd2b17278c6c8e0e406100a41d88c64ee020ca1112ded
zdee85c57a06082f9c4321b28416c08e4fd8f3638b7f00fb58af1a1462471f160123d66dde83972
zed5240100203aba346452d60ac5105a7c459ba919b08a1fad896427996b38ea46ba5c7807ca510
zbc8c88939181829fb1a0a32db0056f1be33831749e88dff26a8ea337c9667c0bf5076ab84e4214
ze4a458a806303be19f2f1621d5cdd2c0be2f528d2524216bb313110bf21342238053548ba72b8f
zd4ffa161ece2fd0547efd11d95cf6072b3671909381d68a797632d70c2f8c2cd9d1f951e2fc0ac
zda3470a5b6fcdd55948ee4247719855a3e47b8f44ff5560742c6f5ae1ffd2148a9506a56a83901
zb898bd9c2cd7cb77177a4ccef914c85670461234b03b2cee5f81d304e436ffcd567c6dbe65cff9
zce8a55bada18933c6d6f79d421d178eecbf4f4f3034f11f5efe5f553f0b78f218de9cf84e6dfd9
zaacf3030a4b279d1b0b11a7ded41f892c3125824212ddb752c2049ae09137bb3e1c93fc9e3478c
zb300d9de950adcd64adf546c4ca91d82a016b13c9143fd1e6d0e162e5ddb96b34f9c2db04d0012
z551784098682ead6454012d700531c4fe3ef468d12ee230bc47e09177b3d8b8bf1c46a8a787443
za4eab09b3a8b63c346b267489fa5d0b202b61d1559dff06d0e258e90857d765117e48763791de1
zb55627a3ccac361104bab639c28fc8cb4179e8f212d9fecc18722fbe898c38e2ef678ae85520ef
z80317b683442839dd3751f9c0a601220d27a53a969d695e8797c92ccb0fd4938af3a4b0d859487
ze4c35b26e3c7f8d34971f99d0870ab5c2229b13396857e26a719f625eea7f588031c65ec7c9731
zfff8122575237c9a0f2155db9f08558494f2c4ee8400eeb081c84cfada18a5e792fe83451ca276
z466952cc0f79fb9bf1922dbad002a27cc6522a59143481487c5e150dce08911903d77b042f7723
z0c0f5dcdbf15da1ea3a3c6ddb2b11f8fb2a2717094afbe883f1604214989913a9e0855a27612b3
ze79a72a21085401f2317326db74c3b947a082825a53a08e6f86a9901f96b882ef751fb36bacb7f
z0be277da4b5ee9efbb0bf73baaf26c0af9f5d7aec88471c3af05b5a6ef0599de511a84260a3b31
z3f81d2eda91babb18c9302da603b0143e2f9237c4723192b299a03ef419174d33847f40b26e0be
z73b6823f89253c17a9967d152c02b413cb2094300cfe536d81309221c63fd8ec7c8843f0031357
z304e0b6e2e6478fd59e048a416ea4a2837a6f67be9d5d38f48755763e210c4b34f831c275773fe
zf905673a40b1aa847f65ad626e0c312d2c6f2d154cb07f0989c60d5df53c2f16beea3254c48260
z0b0bd2949f2a393f2e564820a8733a933b644abc84b6f804949435764b8e90380ecfca25b48b2c
ze80d33cf0c512fbf0335139366ac3deb6db89240409ca348aa56024f526f27b455af7204aa97f9
z4344233fb851cd4fbf351961e07c6ed3abe340e89cdda959c58a4e389aaea4d005fe6dd46ed9e2
zfe29b2687c0ffae1c197d6b4e75c5147bc257d4c33da07f1fe33124ee8652ce6ad9ee338f0eecf
z4f2194beef9234aa7480c64f7fb6038376941a3f4102e8a45f9472222d7bb62e6f9246dbcbad0e
za2ed12dfc8ff130c3fcb85a5dab2513641054bda8aa6a73a5f636a796c4fa11024c2b547c44a17
z444baf308aaf750f88eb54005338147acf257b2184bc93184301509e538dfd89ba8ab84c180eab
zdfdc2693a87d6a733b0fa65a21f5e89387f6033ca5852768fe3be268fe95fcf95fccce401a4a72
z1d7e0ac27ba933ad679894d2722d3f5cc4b12d52dbedd6577cbfbbbfdfc503efed7aa743a27053
z87024a7628980032cec1e47c5830a5b1aa645e143e5a64d9b5edc44283b28bf0db337925bb4708
zf7a5c84929f1996702ab0c6cb969ea29a52c08559b8438f275f14375c1a171836a6ec95a783ccd
z1718413342b63029aefd54a34a73f9ad1d07f06ee33f1b0c3efbf68b163220124d3a3525f1174e
z442f4cb946709d995a6493163c08439221a47de6b9b26631aaf505ba377622faf687e335b73631
z100d5850318e7205b045ea10b7d15276238731755469cf99bda1c879a1c91bb9096c711e7f01b1
z4bd546e43236d4a3233438b9656fbd11ab20b339430ae37583378ec433bf539d46cd71c9da5963
z28654bc85f3e2f6f46fc7d091261d8cc1aa6e908ce106d710465039c15d2ff06b84c9eab97fe88
z612caa64b256ad1db44293a4ea03617e601c3068eaaacf984d2004f9249d548f0eb4b72ce12f0a
z6f0424f7bd69a1bf6dca8bcf505bd65ed1049c857e5c300667f511881fb70c0e05c8f3f145b703
zb39a083035e19ccb130cf5f9fc3d439ccc86eb949f0cf362f54ff572cefb574d8412f9847e6627
z1e36e3a7c952bf323233034ba3148c2284010a23ac128fcd4896f88885319cb29cfd648bf9a659
z42b0a67bb005d8819a3fbc933c6ad06d5a6fceec37914007cf18c272c079a58bbb43d7cc016113
z331dcf5e7593edbd40bb79d2258fcaf52b33aa2feb3003019aad1157f3bba4d7474438498bb2c7
z1d841f351d40df188b945bc40f7339a5c4bd04a21e6714529ad5e84fee438ec252ba33aca0956d
z3313eb8c6449d849a784729f8e79abb21e6dfc8a196d9a20e9f7b6fa832781e2950b6f705b4ebe
z3825320e55c8b6ae6d322f0f95c18facbeab437b98d9265fa050bdca8d92167731588b2b43f5df
zced4a037194bcc120d68ec84699cac49b9c3aeebb5803d53ea28cf4b9c51dd266fa5b435e23498
z7904de70a677d56531aeb6c4f1dd076114c82a57aea03de7d1e8e061931c6dceff05617401474d
z7db59a5909524c84efa37e39be4ccb05df4c079caf8735fe6241085d60e7a2fd929336c4554ae2
z847cb770c37f473a40f291c156190cbb1318f21aa28f9337b7fb8c37dea11221dbe02502339e6b
zcf67dd0c8cef4b3d25efa4086efd5748d226cd2fda7c4763740a138793ff97152a9dd4d5806c09
z2a6a542caa58a2477d0b3fd358f43d85e06355544392aa3e6738bc2db83de76ca0c4eb67aa8ea4
z513d8987e09bb5d53b3e7d26cf931f30b2bd4b2dcc41ae3c0a1b0fc2fd066edb017e48d9463c32
z8bae0931f6d5b8abc92a987f2f2694f3c595733e538d4112aac86326a6e3cb8cd9a2475751431c
zf05ebadbdc3095291300d64aaa6da63b0948a7af3595d732fce39cb4c448acee4907e8adc2d3df
z437690d2d92acc24ff28e8f76103bfd26ea0693b5e3918513e6638322c397c4af711537d571d01
zc13c1c54b46fdd1f0218312f9971aa2b0250bb98577c74fb0ab586bd96250ac2041d6fbf400eb7
ze400dd86e3a8b74ab5f74398180e3130da33594d2597e938267ed547420b4471c81afdf6d141de
z05f647802a480de9a4de33079d0442d02553db0961edff7013492312775fc17d29c897ee85a949
z5ae4738b43aa51770a1f93af741deebe3d45000fc3b37d4482a2e0cbe76d008e4b1d96fe0016fd
z6205f17c7c4df15e59190c153e70b5f22261edf678b3af7915152a8794eb6f8fd8262dba0fd5f7
z3c5cd98a53a443797c04213e5fbf37360d5f0702d2b6970e6d2cae2e49e8f34fd8567285ced957
zd1aeaf68525d28dfc799328b60d7cd69d6075b3cd8e375a5a709766cf94d59d2f84eacaca04503
z26ea976a2712e87fbc333d47dbf0972182d1750142f3db108241af833a727c9c146ca286e7bef8
zd8b1b3b0f269efc74b821945f702cb845bef99a278a94f3c83ae167dada2a6ef27263d04ac33ba
z9e75ef2dce121cb4e16d638c45e60c7e3faf5dddc88e5e34fd7036ab66ff765a252bc931a8e9f0
z1eb2f9396245c9ecf0cdf5024283e173949473aea6dbbec05faa491373d442cbf3c024172d0a83
za7945858f5a38350f48c0c674e3f35d33269121488334657ba17fcb9eb9ad404a0623e3ada20e0
z5800e14038d39b08ec9759f4d25f0c3a0e524958ac84d5747f8b44402a42276eebcc61f3b9c8c8
z313da66b2947ece83f096032bbd8ec04f236e03a7a62a224558104fed80b55503cfb4f4e98a3ed
z733edb1882b79ac1b00cd26442652b323b6b54d7a815d167579c73b0097c61be1aa2c803a65e67
z5157dc3105bff9450afd959732b8a2b7a38725cfe344f9c3f91947d322849bd573a4bcda748d7e
ze155b7e592a5a1aa5669fb2187fe0e529468602b35f4288d3b4abef1bdf55ec7dd6de6af10dbb3
z9c6ab855d89c2ddb7a6ab1430e65e43adc1aaa1fc5898c7be418e2da09095ed430b2338a02650a
z6c8bf3b60a8e1681877b6437abd2dad6cf4534bd85f60d96bf3c7f833eab4d24c94687f84c0727
zefb99d765470cfef540f99c0de36279927f03f859af8b5349b70049966e74c3caa0470380540dc
zcbe008c7dc535369dca9925361413e6157a62e8d1a1c6540636d96ecb23e73539ce9f2eb544c63
z0017b6bcf26940aa978c1361813b53c2d29ce89020a9ec4e27bbc95e26ce5531196243e72b5cde
z49c44ab6fccd4ab48b55deb77d7e591ba6842aef11a170622c78de1466b52a92a2615f1bec7197
z6aa5b5e5dfc1738112b2220f09239f1e58423f33f4412eba9fad0b12ca4ffe11355c0e2cb1fef8
z2505cf6cf0f269f7840e558836d24aea5d508d7de4ac979b2a93db120dbdecc0bcee9e8ac9cbd9
z94937d08b2fc652ab33d4c5b076688363d4fd8f88fd42fa465df4836d147280ef749833cc0a479
z9aba83095328e0f90117d95d759d4cddba0132e24305485bc1a7922cddd8a8d72711a92f4b0beb
z555c82b508a9b66248a2c7cbbef0318a97670e8dc230fe2ce273e7444a192e19736293abda004e
z8eaf28e300feaddfa7da393c4b79bd759611897490109bf4df3ccd1538dccbdb17644836f82b8e
ze49dafa43d442099b3c0138ba42a0750f29545ecc4e29b06411f20d8b7f15490e0166da3cc182b
zcc56965f0fa6b4aca3cb9b537829cb55fa17f598f8c66944f6ab47ccb19c09fc64ca359cabdba9
z18b7b075c1283c86a2e5628ad420382fb47a2c3d23fcb21b707a48ce923fa482e103fd5a54fa45
zd6dcd8c3b7cf9b086b29fdf51dbcd812cd17733400f9897a670a60e2b22b31b939b2ed4d39183f
z5bec9fa6f61e135aa98934209221149bd5ab147a1ee697bab74b4c449b5eb1dcded64a2b4d3faa
z191b967aceefd03c92d15b2b1d3acb4d8b27dea0b985a3559df01bb935752dbee428e96a9f40bd
z7e472c13165e9ae49e11263cf7999d3554debbefc516c05691db5d6b352dc66e869ac1eda566b6
zbaf3f6acbbe75be57df08edb9c407c45a851a9c9301b2c8931296ac6b49807c3e7078fcb1dda38
zf9fad254c876887cd2cdd005cab66df339dc35fdfc3efb11969f3c786316ba2579a41ec445dc9f
z878b14a685c441411eb986c151e8ab67d67f72037f77a64bef526f7c78fb31442ebe3da41325b5
z35864a8062dc0efb9de78176d61ed2cf780b14ffdf3382df67329faeef6f93f8a0949b67f8a42a
z46ae8a8337b871d414b5e2e9f42fde2d19929629101f6fe1edeabae6b7d14dd9b9ad0e191986dc
z5a1b5f98c48b8f185409b3db81710ea7de8f75699a81ccef0cacdf8be0098903050b6b9f87c003
z01d3d21c73e0f504cd3fc2855903c57836c220312fe7aa6e45d04407317b9821fa6115e983b8a2
z536b748f324c9d24ef5ab77f9503dd300eb17a9975d954c5460c3bba9deacc5f8277eb687edf90
z37860c130f9d31d42b6ad2d9117157a832c184f3eda8ad1ac58db974ba6f8250b9cf2d2f4683b2
z8a03dcd7c8bb1988600a3b88ab95476c543255468d743961a9729d15cfe7ceaf95dac26a274115
z2ed004f75fe4d8d37c24af1b9f1c3151e2fd6a5b612a28f518253b678e633e4f18a161ba13a60c
zd8528d8f1ee3fac5e0814ad5aa697eb494c75a3211ec3b3c4d584f2dbfbd499ffb45386a43f689
z6a0d375a5cdfc81b48039e9911b995fc85d3d4fd7adc6dd3d4deebe599c6995a955752423a8c4c
z79c88c14c16951cba7654c10fbcc7ab109d34ff189ad6f664a17210e666b1e1a7ae0a178f1667b
zbb700449cd4902d7a1d764999420b21248e9f2f14d585d5242ee3692d3cd553be2a7384a51f031
z54886ffc3f1cac92cec4554b83753ff3b9a7dacc6ab2fc1eaf4a9c20e46e9f0f51812bb324fc32
z4f98b7db7928952a208df5b764f7902728ce86bc93d6ae7a44c92dab0a4c0bbae6dd6c31386b6f
zb01c8a6275c807ff934a4378422e043820c75f2ee5a5cfa0af747065f11f1c7e321e7b7daa70a9
zb9b27ab743b91a4b7e3cba1665747ce50a4184d65df8b416680db1fd275eb6acb21fd99e8e0895
z9d049457d154dfe58346a68cee1d7434fef04f5a659a11e3d10454b0e1733b0b5eec6a8d4cb0f1
zfd57c2c65193ecccc37b6f3f65118b502f36cf76d4545b5d6e78a4dfee0d387c0e24fa37fb7e76
z8b25f0135a6b03265a99fa4a6ca7f6bce735abc0976b755ecb3ce742183fb7a44dfb0a8900c74a
z64293018a6ca3a49d44de95131b595e0fe7c795c1a6a0ecd28632e1a27b9383419fb7ba9f03dc2
z16778ffd1da65750ddd93cc7f57c8b5163a4d366e741555d904e91ce81c420cb539bea19c0e198
z4123f5ea5be91075e3fa0a0e88b7e9dd84679a8633d3685b56b3642287b3a114a587d5ec1bd50c
z72ce86b3e0006b9fcf37e35d691fa5511a4e6bb61ef5d0175b55ae3beb66dc6ed3a4d928f7c6b6
z11206a197043496d9b0d371e8e71d0b378b0303ce57b83132e77ef2744ba6eb265cd14dfc0b909
z918b200740b25d3160a06bb68de65dc9f653632294e632b94782fe232dd784a2b0bce6d27c959d
z86ed835bfa8209b3987de97b1a8abc6aba78e0f63bb36ebadd9fa02d42aca966359e6f0dabecf3
zf5aad0dea7de37221cb6f5ee8604d889bf23bca65e7e71d2d693d4d6df36d15d601c9362898b30
z1f0bf4fbadde08e62923821384a515125f8d17fccc9ab03c1f32655648b414233941cadba91d74
ze436abee50525141fdde6b3c4e003236931b58959fb1f1c2c8e45488bfb68c9a122dacba7cf6b8
z7cce770a09b02fa3a72f5212f1b98d2e3480006095ea44c15aeb5d204af96ef746531f3afa14a0
z831dcae7e896ff2d4c01750deb09453d8f9ee6c441c7ddbe2a9a7de1cd33baff5c3ce55f8af0dc
z662753f82c9fc3baeb6d9ac3315a620031bc267edd56d7b709583b004f08a2afc47c1e24e941db
z3aae5750e5eff6b66d66d271152031ba6ca6584acdd6505ce39c8d9e8acec7dad84e6e5140932c
zc3cecf0de151ceab5b32843b9ce2c5e8b54bac58d7ae05e2344417af8522e741545f0e1b79dcec
z06f8f35b378623d2c6bedcbe737846bd9424bf5cb0bd7e181ade8c33925a0310d1ba747059f233
z5300d6fbb0632c07ab0e208e638aac7f2538baf32a835a348b3658075d022815d562b46adce3cc
zc3baa55ea36a03b0cc82cc9482d5384329ba8e31db8d2da3953ac4a4bb9c53d29806d58d3b0b73
zc871fbc1651cf8ca7f89ba838987307c095c8a7d74a207d1ef9aa9ff842e3c3ca9901ec42f70d5
ze6b6f0038ad5ff07702096e63f5bba977d29c7e1c3ab915c9ff534f2b5fdcbde9c9d50820d6694
zda16e27af02d69332a4f936738f67c197890b5bc913f7270bf5207fe55e9e9b33433e4334df042
z4f7698806aeded6af04bff6e88d0e4f14454d8de8e9298a99e9f772bec05de09fdf06beda66aee
z284aa1565f300415ef1d6b88337fb667758894b7edf74d0d961ffb3bbf2c6f3f0b0633a282c6d3
zde8ed5bc6df7ddbec949547953abe16a3cb1d70931b392c714808ab6171b2fba8ff0c228f7a634
zdba959b8de71f4afc15e36e60dcc938492e59a9a59c6d8cec05e5ae4571f77c8061a28e9fb0fb9
z6165c191d72435b4922f7ed636f11606614f7306d27de227ae0704339b8d146bd1a1e6266f7d76
z05b3796da70a5839109c6ed688cca799eece5be62af87c1f7e064c49500b1c7e004e18664a26e2
zc56e75150b053dbadd2a53d45c0f5fd5e6e3e83548cbda54e4e89834f13f7438e150ee0b4bc669
z576f214844849b03870c7100567381fd0efa01654291906fbb88ba36f4a75e8188ffce7855b6c6
z11f00371b56ddf4d6c128619f687a96882f193c991b6239bf556b888b5905b2dc9327972c2257c
zbe16870e7185b0453bea2a0980bb789570c31bbe0b21a2998b70cd14c0c6fbd9f5ca382aa18697
z138a9ed371b3599326b71b34e2b986d04f51024fcc44e627071213094d9bd6f74327d9e05c4fa6
z851ab86b0216af453dc8bed2c698ef0891548b9bef6165422241240edd6b4a110ca6512b02a0b7
z0a05e654fba5d94a10710f50bbd21c31e4777680477ae741343b4220c6418064c4741c80bea661
z7c06c75932552c42659f1aa66c6a526705eac4c01f0ce966b2883aa7f278bff79697e048545241
ze236ea19f947dc4deb0742a2e8c8e8507cd0a5150979e5841ac66aa0e51c48b7c60941c56cb36c
zf2c97f3f2a028d8c8b133f5ec8a1b2d49c459a0956315a7c8bab304ae15914fe6a9b6bbeb5bc44
z765ddbcc56181160739b987bb7469be00138314f214e553fc2c7f5038c0484ecc64df2535d6215
zb4eb83f6e8771837675d2c5a9a2012ee439cd71f95afbe762d1e5857db6e1f6df6493201ff71f1
z0eaf32dec3fe54047068619592b20abf94006ef986a2de5c752ccb1a7e3df1af4645a02a9c1363
zc63a00e63db392a7c06c72a211c1089d0001fa78497b7e426eb495b72d9226ab376cb23f0031e8
z348480e12cd03a444a3e6b68a0b91577208e9c44d764b5609b476a08c89b0ccc8d7c1110e00d2e
zfdc7c8174d92d74cf5988e4242eecb2abfdcfe6dc4b57f6f9bed368fcbf36803fd0eb75a60fa3d
z36e675b70377c16b2ff265c8afd18133e8f141e96e419d503d77d21e67e7bbc3b648ead004ee3e
za84bdc74c2907c554ad028e84d52e458e247cad07a0dab93e0599264a4ee0c3b919fa23883145b
zc31fdb3a8527bb6386884fe7fb16b19853127169c0b92af541d3b10922bf8b2263f459627c0ed2
zec8c9f79884de02efdd8b5802293db1d14ca9329692440f18909c54df2eac46588708689273937
z303eb38302e1c114547247c348fa310d9aad6c52533bd8c9a67f53238b55a5426f18848b08f863
z30a5e6fcf9a5552b5dca9e461987d001bcd9365d55f0cfe16184a187267fce4b83556df96d2d73
zc422ac5b3f0e9d1a83173a9b4be8b031ab0932858ba525e4e3f74594d5dea512230684131c35ea
z7d5037eb4ac279d1d6302716fdccadbdaa23695b1eac4280a14786349a912f54a3481cf9e86653
z2a9d2f6d5b7c8a39719964c902adfe3392ad5cd5b913682ae1f40eb48e0af920258279e49c5a8b
z6cf2fe08b4d52d9ed32ba359c78e7a30381f6ebf4a47e402c51cb65b3695ebae00c8690c2a2f13
z5baa19fe0c2c40fe7e75b2d626896d000149fc679ed6d25434a9cce6529fa8987130dcb405869c
zb3cf29aa983833130f643e3b8fab588cbb758280a06729e7dc0513895d12577e51485f5accc667
zcefa93e27a92ea38f17d7ce09cf297b02cb0e00c06593701e8b76dcc1581c942fa722598dffbf3
za650338f184e6ac829b4b58092ed7ab773744c3961819719d7003beb0b8b529360bdcec4ae4508
z5793e30fe8575301f4db84732d989331fbb91944dc65ab0fe275bf909a05a2a67daa4832a5896d
z022dfdab49d3844eb20befec662724d68930b2411a8e216a5bf7f58647b49eeca2b3459eb9e2e4
z3528f80a6b7e0be1f67688906e7ac11d7f0e2758fae12d6bae7bf3c8e9c8829036eae3acfb6769
zd5c8036fa9702120e4b4a7442c687465847ebe82ea41a2e95da36ed7f9e197f7d61983d7738e85
z091a7c9366066bd8608791690f1e90545861661d5318de2c19121237b683e6c3d659ad5a964716
zf85875bc84844ed50380e57bf7c4be7167287ab6931fe71dcde1910af633adbfe7a8f20b190945
z5da67026053f65094632fb6b9fe1052cde6f161ad53b8eb9e47fc15fa686ada579f8caef0732a5
z078b3b42fccb374acded93772d6a6884236e833add84350957b3035d444f85d67500b586fa122d
z6bac63d7c0e8549538f4a836717520d50f943302b6a268f787e657cd0ce8ce1ea02b3b2c941749
z38d0fa9d04794dcefb0ad7d9e43566c86b4e1e6ceb4b41eae763cabf65bca05f117f183482ba5a
za193a964d7209a9356ab8c01589ed8c0baa9f96683001c69e83a6a1d5bbf9c2ce8e5713ff1a5e2
z4f053b5ed34d0f9f89e96e6563b9256e4aca4c745b93909e9212e5cea465ba59c22fd2af58416f
z9d173789e4a59714a6182067a02842318d9bc5ba7894e9d6474357e45f6c19cf6380cf84a155f6
zf43579d60885fc24b51fbba98ad7a1b4c86227d3dc427791d7bf8e986c69d59ed8719adde6531d
ze1e23db53c2108b9d224718effde7e335f4c887032189c2ae08c2f3e45b44147b1caddd19c1590
zbbb8d037be16daed3e1692a1e5d98896ebcc733aa8aab4696cc14ea032d394684733361e4483d0
z80e7c112c67e0901bb30a346b692cb30a6ca3950c8f8ac655c0591b7573a6c744101373016ac70
ze404a765d6d7b01742d88c37e42d2917c2ac8b6d7dc1a0a74ff44cfcef63d2a7685b61a0ef7234
zfa5484e667d933acf9849c693d1e9f089aa4be2c41c74d76cb61cdb195b818d5db096d61f213af
z219e9730dd23d3d93c5ec7dc6e2ba826ad497422b77f16908d2614e4c84121642d827a4b9f93d1
ze3bb06216bb85dfa8895a5e74dfc20f816ab0deac9b806ab135188e72bbf51b0cb6b36b30b1155
zc5ea70e063f08a57bb1e31c9e73e6f0b28310f9b83b7304913c1d8cff97315fae43a96994cb913
z972e9fb925f9e1e4b12710e6f324b18ffa3c77135a863f4b7e1f7aa5a25715e478098360423609
z2eda9b6a2c1164e20790b6cd89883643fe2b4758d74613911003a68eb63bebd44a537d771b73cd
zb18045830116df1c88d0ee18dd2b9012e0bf3c076af7bd9996e1c01f7ba6378cf7d5ee2d9c8f87
z19a1438a128f42caadc3c2dfb9fade73ef5f612f6a092549b89387a7d9a254d3c351101c118f58
zd1bb32a709a5ba4c37af9829c4d0cea7a6d98dd926eb996cc91906f7ed99e53907829606e2c872
zd705070195e1592ce94ad35b43563ba292f6ab930b512f71451ae806cdca4c2cfc066fa9723703
zbeeb294f1c0511bbfc8c65b2f07dd884d2c408f75072c2d6ac11e65cf892c06f5335283a877132
z7665f90203c69dfeface29c64c71b014c71075dd070cd67845c6620cd27eb665220edd1befcb64
z499f913cded38e2e9cd9d018cee716eabadcb881123b43d09fa9f787eb8c834a7181c12b678be3
zd97da710887f37b13dd1c6db42f25593c5aa5e4406fe2ff802e105f8d30f5f892a483c12281726
za7daa8e7bc41198f6b8de15c5103cc9ebce94a5a9fa2102d120f96d069005b1472fe01ce39b150
z5c1c5e742a9a5acc4643a82f8c159a4bdd31b0be3a3576dab91da03939208494713f62ff3df472
z741fd8e916ad775046470d21cb34abfc48bdb2e211f1dc502264707bb94834d574483cbeca190c
z8c84f4bd1f16c488e403975ae02b3f94fbb4c451b60ee37d90d02c7bc3bec7f14cb59af8960c57
ze031fe46c27306c6f6f02ccdc7ff00c85641067b5bae6eda0d5cdc93ef984ff27d598682f35b23
zd5b9ae35e207caebc72aabe594b1b253044ceaff8bf966408c9388f80fdc4ade1994fd55c00e69
z3acafb7ba77ea513706dce62f73758dfe7a6db0c5d3ab8e16d5873a228c0ff4e58d50e5d023fe1
zd1bd1518bf43b40f6e4b7a73c05db35dd59531d81ae1d8c96fb80576d85c8922e63a3bfa328b63
z920bd1e3fa1fca7c5509383feef119b72731bd71100b08fea230c1d6ce180e5fa3719358ff202c
z1148ca0a419ee9b87474eec31a2d191543cef4c0595121d3f80436cc1171d5980f9a010954317c
ze89715b9a549c0350bc9676e98951741fcb6b15852099f040cc24009ec9df401fa90de831b8272
ze0eefde34d66a8604b0bc9b2f8868a7022e1ddcc546fb7d85af1fe998ef310a28586d409312d9a
zb9efe7431871d7bfdb4e20821da7cbc5aba0c72745a82bc375a68d39f70e64f70c07ba633730d4
z78fae11d1f2a78ceb37c80da2408c7f7b6a23af36d4f3d42e8ac391aa41666e16609121a10ac22
zbc3a13f3c2b910ba5aa1577382a9ef2da9c1adcd11d612aa389816934194765e194d1cd39c2917
z863b56a55dd8916f3369d0167cb8e61133fca66839e7daa33105f0feadd892330d725455625da0
zf7c0467622cae9e371cdc0916d866288b368009ad01ed2dfc51f7dee4a1bc8f43e250c633067ab
z28a3f405bb8dd7f287ec4351e4d77e2a3812e5f0821492899af04d991d385ba9ae7cb83a61a812
z19273286e2d820e6e5042a09113199186eecd0a5b24429a4bdfb645ece2071b85eb80b1e50772c
z343094d5dae24e303ec0c2da1b02f56cf2d8f520597b5f55c0147e6673e74a466655b4c130b88c
z3842665664701ad4c4e898ed882a473d039fd9d9a2e3e48b0b3831caa2b66fd895255f6c0543fc
z1915f25d4327f01020295bd665ea7f1164726dde52ec70ee5fe8161f0d3d18dc58536226f8723d
zff27a6509a6621b9a7984fd4f0c23372673527770322d06c1b799da81e84e02a8244dd9fe24db2
za0893b89c8eef2ba0b7574ebe88885a5ac7948f06edbeadd86dfe1635eb4e8fe4b5242457be085
zaebee75396b5975cbad4893a6f9b3a00b106193b20e40d3dfa22cf44cbe98e3a4ca5facf3b7290
zdeeea5beb8de433f24ec688d9438cc78e23c0e6cd5a50ede73fdbd92fc348268ff9b0e00e7aee6
z4b99097fb552676499f7424ac579e2e394c764bf930ff540560e2bb4306a2d430f8f9b65f2853e
z7c7f41a598c9327f38289f5572d347752f9b5ae5f686267d2e55923cf2a1de6d2b7a540337730f
z9dd0446ecb09d78f00c486afce3d9f3497d7cb538050746f73630d4c086858012cbc88d9c579e7
zf05724b96dab25bc678d4950689f2ea915f6d424042e91b62fc4255a7c314d28babe217e49a64e
z343879ce768b617abfb1224c8b4ddde97c3324394cbfc0360d2edc6a0e06ff396d9cae7712195c
z672c506875ea443435b524e26af6acbd5cadaa4cc74d533031ad305fc310fb139a7ddf4350cf48
z8e1894ee9a418533e9dc7e2f10855854651fac8917e4514ecd40279b8982f5a3b44f9e733c289d
zb9cd77973d67b464a86f44c0dfb79346b1fc9fd42d37c059339fc6cb93823b250d9cabdb38fd2f
z831780e45d9ec65f0fcb99bbe41986e604fca3d22f17de294d5c8cdea10734cf09dc825605e6a2
za9e8d0defed0fb81aacb6fe1775db1a915a07bd72c7223040c88f53e7117ab02d558fdcb9eef6b
zc1b0e1fe189afc86fea65622a358cdf8aa3864d6e85249fe4dedd6e4b43685b4f6f403af107752
z7787588292e469bf25657cf58daaa9f28daf9264e83020552492015a4b6a5ca990db574b45b2ce
z60912b490c32ddea89d2d50184b87723d3a355bd76d9fc0daa457fe8c848411e6dedf107ed06c0
z97910acce6f24a54aa0335ca1fd511cec5ec1aa6ae35d1a33075e9bf8aafb8bd51287955335542
z3daeea064013c0722435e7d0da92d12be82f461f137e3ac8c10e87c80ac1fcb5d0bb2484194001
zb1b5931e9f6dcc362869d0294c7248bbe03831c52b2aedda3a73bab9dee1e245589a6e763335b1
zeca32ab2c1801ef5fa76dde6a69ae46e1bc674d526cfb21bd54a68e2f56076b18cdb29de9d7d02
zd76d64753539119edcf61f401781e102b877ac9cd07324b7a02c62ecae0214077107fefc501136
zc84ad80acdb347275bb829a447a9ab1918de4ddacee3397423be67ce8aa0ac65e26be936358acd
zf69da1a381446eabc9041d3f1f5213860a083cec60451dfdbca2ceb5d625595322c4ebc27d86b5
z616147d9d084cfe304bda4393fd3da276c5ef329eb86a6681601862981acfa7be0a4ebe1985c74
zced7eeb805f784e5fa2c68e13545dac443a170f48858aafd0f4798c6d146425fc79285d50a8f1f
zcdfe16b522d01d30b21fb0ade261ee907b7d51b306bce33d19c6e830766f6273837f57019b6e27
zef98ab25ce8ea18601bbc72e8d6fe1ec7785e31e85d86f45cd6a4f340d769191a122e6c7fbfd7b
z2ed1d2b3731d94c80986202fee65b85cc49ac7d6ea1c4d384ccd810a5cbe2440a6e718ccc03eee
z66cf50b9b3de22d40be5f5968424a07e904886905d6ba2ab6c66449eb422f8b8fe6dc829d4e33f
zc81f43ade3bb786ef645be8e936c67f30b9867bf23c1172c04b682c594ec4948a4f55e13c887da
z015f0e8af1b82e4e23dff85076f3989955c113cf4aaab4d651d8dfd62d7498a0bcfc81b61557eb
z763f2e8e164c83f5f654eef70df076e8ab9d2801ae17a9761d6fd7bd2fda28d1787bedafe2626a
z5842fd3b0325bb142a6923b1b8a862914d184028fe2b30affa01887c600c908686ef2b286a30f3
z8a9ef60e5ae957ba8bd5dc245e8d64499ae35f7405b714b472462527280f91c60800b84313226f
zfce017612099fe1e9d19c19545fd8cb00e743c66fdfefc7567b3af555515aa13759d40002f364e
z99c193117e26b800c4c07547c0f4c879b8c6496002f00d4d8e8b9fdf2b3155833b2390e8eb8424
zc7f4e08fc93dc2d19f32ff8551d9712f3dc496d4fce3383f7c7b4341c13251d58b04b40e8176a9
zbd0f2f5b8e407fcbe907b9e26f30eff0e9f7c4e34a3622e5060e068e2497ad5d0bf71dee194445
za29bfd500561a083bccd1a4f0cde20ee054ad6176a4751b9bd1dd65a04a0ad29b9a31c1e9a2b29
zb0473b0d0e4ca056a2f8195d2dbda1c0588893c2da3f671d5984050be32f2332be394eac919bee
z89fac1b74e96b19251c8d84ffa45b27eb4a55a4dfe43b4bdbaa1c63eaff77d20e8ede449364305
zc0dcc16354c3b898503945f13f7a320b2cf78b4e6ec686e9ff020b12b7a1831aa33da09ee9f62c
z8bc1c67cf53161182917726693c76e842de193b30a89b62a4b3ed5febed46916604cd645678111
zd4672d85058b575ca54211b123a79a70ef20e119129f60af2f3102565841d42259bb58bd3ff7e0
z048a04543893c94185f593c5d38f99428ebd1e200e255df4aebdeb47f31cdb745dc8aff08b671e
z3af0b27284c64df32d779185285bc030b716864c23ff44584f6a43ad03c2ff173f22174457e443
zf0b51ba7577f257d057c68a56da221e206ab8977d85efca70c2a8ac00e53b224950ff4b5acce4d
zc76da1fa116211af882993ac48412bd418a56130e5a7a9c8a2ca6e99722089b881f2ff79340e98
z98bd1881030a378ec7925faeac39df248816b42549f59aa7c413abce665554c773682a421047c4
z0db1642eda5c90255d9610f981091fb3ee41c99443b583fdfa1c4235932099c47e5b921aa3eca6
za3c85533d931f158e7b8492e87e562e9bd78e245a6ffac2ab6b1c430bffaf3a6a172783dd1e0e9
zf32ec00089dc67ada6bb509b35702a8c8426387b2163a933af1dec540ca8e4743814c1e281bae8
z014db75b52ab507a24b72acf16eb980d962c5e2a22825074d5512580c760746d6a4f9dff6d4d8b
z517344a71e25e00ad05d33c689d572442f6f07d48edd87a09c2be41a3cd9a92af0008fea2fec64
zcabe4cc45205b5afe88f2951cc9b0e23705cb1687c1b5bbff06b81e24c6d635de1e5bf05182a98
zabb9023c0a38edc977986726220229002c05ad7e473aa96b0b289f6fb8f14b41c1a050a17df95d
z5917be480647d0c0a7c38ff1822d58ba4a6393166ca0f9f6ca4cbd8da27c2bfd676d8bda64087a
z7cdccc1f24a60d972c8506991aa360b1845c2ed9bef13ee66739032cfa4d75ec414cc45b3d4e81
z8ef0fc9bf8d35a8f4cc2fc303a372af49000aae1a71aa89ada8e45adbda6d7d6bd2b21c2813a6a
zcf1f73d0cb70e90ea8c1f0ae6a3c5445f155bf87bfd8f06b32891091fbe8a3a646ef21dce0d888
z5e88b07ccea9797d3093fd95d882940cf615421733a4ca5e0f54537824288425457977cc266e6a
z2bf6dec34fba4907c6e988e2092e81c683dd9823b54546fd92bb7a0e65024a7232cb54d6d13ed4
z9f29c3c0a910336942938ad791a45c0834197fa2f7bb6f86eaea519a8c060f872c164a8496093a
z5907377dd0efc54c62f0d5539af1de805939f14ab4653939c3cbffeef8fddba26479c1b504d3d7
zef4b5df84078216e6c6fdcd2cfac2186f354a4bdc593935f9d480a0b50b39af765d637610540f1
zcc873647bd9cb46bdf9d4dfbae3f39de825b146a1adf83f859413771f9d67bba4cec156f7fae8f
z8859cad3b7bbd766e18b8c359ba03bac3058ad52cd8ba3a9f1695ee1c96850628623ad5819d699
z4254ae9b9dee0413441769e822c8d592bbcd2c61e27a510a5b6f6d1ad4b124e6034c64ed736bc6
z734a587e753901bba389114e6f8535a1b935e3e55e6b63883f9b11d55490aae06b7b6f9130f27b
z5c3321aba6325ce3ac8b582d52e45e8452bd452cee7deccfc68ed3632a5439aa305e6e0c8fa22c
z820d21f18c250a5fc47d199c4bc0fa112def45500e1f860cc637d0703d16ceaee6f511e6484868
zed8fcba39e1492f845b1d5c37d3a0caad3205742fd61116cd057192403eb7df356420ffaf4f7bf
ze19492001640bf0f15f02cb9285e35dbe1542448df1225858e5c4d307702acd64ebf487aac9a3f
z5bcd9e96bec3cb1a42f8dc60bf6a1fc91eab9f49772a03126c9b85721769e3f86060e0f00a08f4
za5db4a13f43ab88d43f457b5867dc42860b23bf58d4f197786ba7bf7e25c224d360aaaff49fc90
z271131cc1774bdf0e1a1045193ceefa24fafb3213d9c32aebba799ab2a9df755077a95b92c87d7
z8b3a273f37fb0e3b28a7d39ae84b50625cfd891ef10b3a0264ee0f637624110a32488c64cff4bb
zfe70abcec74d5a31c8fdcd51bb27d5e5a03ffe43049170b4c5f051494f12e1b75ccfe3a145a620
z7871967f0ed997a03bf8c1cc0045023011968d883dbb09b4badc2e9e3658528295559b89b0e2e1
z3246718d28496a1328b41ce57febedef0f19145713e883d07f2733808f3bb288822e8cf4929ffe
z51eb18c54e32a6bf6aaaa2cd01beeaf56c3f7277b2cbd6427cf0d91bd803f288ec99fb9b8a5ef6
zf8dfb64f219d951e502fae9037a7dc40b48f338694d443576d4649ee08fa0112d2c2cdd79e0dca
z5b6a448707f5671fb50eaeec45f5a7428f4b3a9e0c736e0015090c0f63a7d3216bd64314aa5933
z0a510355f75a422b125ef85714d5ce048b3e27429a3e3ce11a90419a3481dd24cc6a435489ed29
za6b66751ee8f3f7a2c79f836439c5a4d9e17a76cb0f932e8da355347c3dd1522367b86f7ec8b1f
zb8a234776b0c4ab1afa3b9610e8f37c4cad8656c38cf3f3c0d27793935728c378b0413dad02c9f
zcda15d833381f70757e6af334183b10f3dd55279e31fc81e47f6e4c464146d9c0abc9d968c7c1e
zefca998baa62120cdf8981d9d791ab14d4909c838d7ade7a01b873214ffc8bf902959be718bf1b
z91147d2b98f64c4dfc270f916b0c71fd2c3dfe1dbfdc3f46f4b2f13c9357f5618b84cb012c5537
zce23af6ab02bcd70dc85fd00e1bbc50250e6d6322ae28f20d5c24e3a09e18418e8b6a73a3a040b
z66d7e40cd70b343d6abc3e150d78888883e218f145bb6bd45114c6acacf0ffaf8b88e5252372ba
z17bdfc576a9b5350919b692e60df2d02f0f38cecee38701597c0fcc4612af77f9c2c0bb908282e
zf9e08d5a5a0693d4bd31d55d672b8ffafdf292abd2641f256cd74d52ba1aca99ea6dfb4d8fdc25
zf3c92dcf38c4f32bb9df963d4d920d56e7f60d445a1dd536f784be31976f36b2bce3b82fc56498
z084edbbf4390f67bf2cbe0b10bdad21961f01411fe0789e1a3f225e3a033b7641e041a0fd4e706
zc85508d7f9528bd7d50a8288ab0d6f7d1d3e77a361850d465d9683414ff547fa84138d5bc6b91a
z3d145b34450ce98350fe5de5f32f011c63084fd2331469b7c7c4ddc0a0d0bdefaf500e3c94b30b
zc515354929ae3eb47c2235ed83edd760ee42507a1a5e300ea0b9bb6936726943307714163cbdb3
z1079556c07a62d614a61e534bf646f49dfc51c99befee7e4d4ed0f465c38ebf547375e6886585d
z577cede56c821ee65cd9d03c1cba11e01d413eb6092a36a8bb7f42e1bf22b9fb1a15719327ecac
zd82967873948e543be59176315cb0c006824163dba2900fbf2e9ee824abdb2e7ec68c71b553242
z98521a020a46dec4a26652e483226abb019849df5c58a5397489a1ca8b2821f51ceb9b53030f3c
z59ad694577a819210f1abf339e6f11ceec6538e304fd71c99b73a5a1bb6f6f5bcfe41e6eb48f94
zd14f9d6b867d0d5c7a45789793afa97c0ff145ae49af90e286f1a246bc1ffd725c4e098af735f1
zf8635a670c26c34f291d7f0391feaef237f0d7f2729a3be2a5c299fa175566ea5e34b7c4bd286d
zee4e9e9648a5d3ad2f1cf8d8e1dbe7ff95adbb395287b637f84f9800eae31b4838894dbaa6acf2
zadb695735bc6ef950b466bec06025fb42a886da90f9f2feaf163f26d87eddc230bd11039c291fe
zf588d87da62030d993d8dfc981efbd8bb6c4a4e110114961e7ad9e6a97a07c99b2011bf30aa686
z0a998b22a10c8dd9e8a8a0abde352c8a8272aef680b08e8f40e95de425c1cfed96997e3abba9bc
z406ddf4a2ba67719266b566f2b8ec954d57ea20ff9611614930bf980495a9f8125478562a96829
zdf6580a019e84acd5766aa4063dd50ca6c56e23924ed9f53296e795664310b83cb6fcf22bebc5e
z99476a8533eb8ea9d464aa3120705f7753949339a3faf6d34da6ed01aa9754781eb15e6042fcdb
zab739b6dda52ace5c9b765b989733c9ecbf30211315f5a2c847392610197de1d5b1db3987aab65
z1f52ece1d7eb9940ba832147ee3f9d9a2f770f87a74dee99afc11c18e08af2af4c294e4965aba9
z89bf07867daaa9268c8d389010d066e3a77a782dfe0ed98ad6b8129f653ae4d1ce542d1eaa1ec0
zd207db4b08b152cd3ebdc9d04259dcd2973e03e7d2d7dcacfdea7f81b8033586b43b5f94ec973b
z85619d2bf41dbb53ee8fe6d768f9c39ea83eccd8f1a7aa5fe5f47aa25d5b7f7b61a745d9561e4a
ze1f6518266314772336328550dbfe7572a2b274e4f75bd92cc7d8e1d089023e19b3533ddfd1209
z85f2d452cfceedbd8b6fe20e2d6fccffb0013c5eef34d870c2d25ab4bb6e7639cbdbc2039d5653
zeb066878c39af002749872b58c1cb8cd72ce339725cc3a7271df6e03bea0570128afc6c06b5508
z3029621fd672170b1f3b053d9ada3ceb22a2059f3641a9db95fdc16947d0c8a7b1e4c1a27387bc
z13e38992145867ea9b043151bac1feebd52344e1189cc00b82edbcc3b7a85f0f47f89243668e17
ze597167fc7b7890bc0f48f5e26395523ee8fa2de053f915781bbd1ba96c71538a8d8cd07ae0415
z18e5d69b1e89380a3a545a0246366e6935485a006a0d90dde122d58b2f3012c49297a4247d3a4f
z5eb4d6c290faa2ae27564fbd4a9de4b574c056d011ca26c40af4750c4393e469f8406db527306c
z6237f55681d631f858d28c0af728fbbd7a5746d0d7b772d303a80b7b74182f760783008831c999
z0821eb5d0433a3c4686d7b684e0f827c004cde5a52be7d42bdd0a0ef6c93217e6fddeff998994f
z6ffdcfde87f17838050b2de678666f6954aa8dcb4354168d5b996f9d10a52c05f829791f7f8943
z89b1dd328d1ce62dff009ee2f5d45958e0bd86feaa00189419259a69ae5a285d2d38c4dd16945e
z70ad8ad4b72894a6c5653adf17fa410761375aecfac6d79cf790d43e674c1bd3775163732a070c
ze4730305a6e4e468bc7b05e22786f19198f45e62dcc4ca3c0116f941c6298e15cdaa7a0d4d3d3a
z9f16f5f2551778a4f17deb5b996ff90ecc2ca22c5642efca7781d4c9707eea1de40e9cc0e1ab80
z772e551a9e311841503192874f23917b439e6be2792bcf12b8dd57f1e822cb12aa0f76fedd0814
z7b32883e6db71e198318f73e8568dc6a6d2e121b1e076a6da2da20ff14c941ab2a1496fa5d721a
z54d20905d36771f3d264a9ba025a9693e84f0aa088c283ab598ed829166d4f7e4e800025876227
z2436f3c94e64290e0ab9c126594599ed208da29077a0ccb1370894020c2bd0d3bee2629e57889c
z1a3cf76e0b405e3ab6105fa5f607e0e9472c6a4a5d0cd5ec22e98f2a4180c35da2917b4bda46b1
z5c8584eeb2bdc1410a1160c00b0d6dad279dadb2d87f5cec6c6949b1d0b8aa489252d0a0f6c001
zc2e54cecb2f4b0ad541926446efd1d856ca823460e9bd00c8b86186560b9c951e519919f2f8fe8
z8009b5da3fce67011336ac7a671b144a73bf9997eafc25515325542a8a8ec2f8ec70abb4aa488b
z7604ea026e9389c1f81adad972d10f26228efa60ff3a9606e346ce5c384ce1ef3aa8ca22a71418
zd387e479ebb7c2b26695b8bdcd28d25ab459a44d0be5457f4e00c85c103ff4d7eccedfe303cf92
z9914ce1dfe19475dc4da40082ef5e991442f210a5adfca778ef55e717f749dea9ba4e324f4f0ee
za03ff804706e4106f8cfe256806a67f4bc05cad3089430fac7c330af9b07c82665169c94648874
z9408f41e3ced76ddc66b2bc71727f3dd99801a931639dd934f69bb703daf005b5ec0f658058d06
z567a74f4555eba88668c7655b708c3c2ef6a0732fd900019f7acef6a162be0c5102c52acc1c585
z164d99f9eda7390945901ea70289b679e9ad4f1c0656758c9873efcac2a31a9d3eba4bb9e4811d
z6f0d9f36bc7061690ae6213f99f3601f78c96298f3e4dd4fe3d5b27a7cfee70705c109b14af78d
z44982db90699f1cf5caf81ffa4e67d8ecebb2ee12fb575e81581bf25e4473aaeaf3f1baddc84f6
z0cd376e76797fe634ac2dcc345e593879e4d42c32c91a890b6c4294a4c6003623afc9c9823ffce
ze2b9fba2bca975301c044a6f9febb4f6e444a2f2ba3d6b1ebd1d771d0902774dab00329a89efc5
z98a64bef97b4f0f2cf3fc5d97d2bd5eaa4b215f8cce28653c5d1202c7409e8dea7acb69a9f895e
zd69be65c948ee814058123f86890a57cd49139a004c78b33c2a5a9df9788f3ae3d3718d9c53676
zbcf9c48144a6e8be5655bbe8a3603155fe878f0c60239f67a72447ca072c8a08fe4f10864368ac
z28ae67885290cf75a78b5cb35119e9d16725a3574f726bd03244533fcbe907d2cb42e281ab7f3d
z32aa97417c3b4ad65cd1470c61ce74876675ccee867fbc7ea3f765441032197fffd6321fd79047
ze2f172d29bb61df09dafef510f94458b6a3e322e72a576f26c5997976cd0fddf62c786dd3733e6
z44de3554045b7f5cdf5144cbeaa1b222b0495d0c5612a326593996d0353a4ac153358aaac61a35
z8ea3ff5923cc58d1d93209e638b172180c609df65ee1df61944aee2643d44f37bb787415a08a27
z8dd452d50894d1889a8c3cc7dcc180c56ed31d0a0f798db13452e4927b1f8eccae6a2fefaf763f
za396f865fca4a2af6539a7e982a92e703c0bbc1d5f77d8006e91b9f08e7b59254185e6d83459a3
zc43495642d4bec62252ab19ac21c0ce97371520f43b7e8f606b77b65ee627ebbb90b7ccd0eaf22
z9bee13e8a108429ffe73b7f77a56d01fc1261a61d95918c9256ac66d447fe7427f641459d07a07
z6fa00103c5c007d82b508211c6f6ee925813c5a3c1f4b62b67250448170d5788c7fa673cbc26b7
zee078368ce7943906795e328fb82544115a5c449fdd3ecf5ae4ee92c92cdbcb25c2c220b3bde89
z15852b9992e4e9e96372f8f7a4eec64182ee31b67c3492e0650b82de51c241f41a21d6e96c3e72
z8ed0f82d2ea46dec2433e73c5b0a7dbf80137b432361dfad1266b2d104dc4c0be7cc1a33493aac
zd858a3ff1bef5bf29cac3cb338cdae680831f104ef776be2049b7cf9634a167950c3c02732414d
z3425655f0ef190a39387e16600010f4a21d087d527470bf78ea5eddb2ceac2ca7c16e5f1949788
za17de3819905dd422a936d18b7e2b8fbdffd38cec1d4bfb688ee74cd5f29d153c201e2d9b12f74
z48da9fba98daf37c6bd032dcb4f6673a6c70ba3ff5be7792d0539346cea7c79aeddbf7d793aad1
z56d0d24e23775c4fbf0300d12ce643031c1d03e38fc7851e6df402469fe19141932a204ef0e595
z2d7970ce8ea7623eca47aa05537da146e99e7e1f2a634311c424237f26447b5eaa077f24994b5d
zf48300da7853655a34dcd38c284e385d3bf8ac744caaa5f0da55bb854bebb498c0cde574aa0ab7
z808884f8a1008075e80f1708df459ac6be00cfa51ee4a0bd4500dc2a323fe28f49ea0071e7f10c
zb52fedc8ea5ea8d20848b600be31fd9d0abca37521b9d7910a1687b84dde722c49ce3529dcc028
z644e48f63d9454d21f450d934e0a7f82e5a9c98a428bfc385f8ea1af4ee97575e71ba7f4aea1c8
zb6888d4bc4f4ebb0b0590d8feaa8fa80d3524a1a2bc80623e712d28a22f328d31ba526d9c0594d
z4074cb28970f48f53d58b8a70bc9fd4c622d8f36640a06139f02c8e4eff72a647ac2309180617b
z6277fc271329add5c2325414adebf96553fe7e3a1db102a2ab3b0bb57c1f1a5f0a4a7d4c65a455
zba792371c4923472b14b26b92943155fe136770a317ecc46a5a1b30dcebd612a4c3e30551709e4
z71b32fbf6ef2888104df55c245cc824f9b39bfe73356096835cc2af65f8b35f405f5f26baf0103
z6821dcec553c01a1ae739db34f768f5e2e8b1f973e833ea1941f869828631c896aec08d7195af8
za2591cd2e29ebe370b3e7a2aece4e9c4406b842a32e8225420b58560ed219f9c094e72a0cb5a44
z4ad842ad4e55a47dfe13f2524ccf7cf7184f27c2fcd8331eb706880f71d9188244123409e1d15b
zbf98ae471f273c2c3ef18155fc65dd46069e4a1807e5d4cc743aff5059497fe585d83fa8525386
z5b9b9c1f549a48957ac34d2e7f5deaebe7287157308a83306a250d74d30975a9ee3e352a1abe26
zc2a467eb1f552de5db2fa28bb37073dfe5f5b77b762eeb54136fda998c7cab9df8b1bd0441b52e
z4e0836e7c6945503f33fdeeee018de6b880cb7c30d47fcffe10dc0a545174c5ec6f81421ca31a3
z936eb0571d5f5ee86fd3c2581ae61054cad27cc2b1bacefc357bdce773a28b234db444df522391
z599bc53c559120854ff144428729b4a15f48927e6f085738d3e1e6932724ae2c27d996414dd35f
z5eed199a090ddd5ef381e3eb3b81211c2705bd6645c5733c2f214cb6746207d5e66989000b3627
z534b84fc388edfb961edf1f53512ebbdfa7bb1fcefd6059b4a79fb9bc5e531f4ac2b5a24f864df
z1f3bec29bf811cfe4634636ecec7646e04cbc57be9eaa9ca4c88b283f76e87dea7422eb96656f5
zfe12211f71a059d41849f192c5693cc26548ec7d64eba826df80a7aab540a06cab9dae68708a94
z2178946f80ef528bfcada82b8cbae11b4896e5ca0d14ed71b7e8d55e5fd3d402b406109a34adf1
zbd4ffa9a4827f8c6eece0d1093a7b5286804e506c623f51e27dd815843df3d06c831a33c8fca89
z46761733cf90b783e1a4461f113ef2738909da60b8c3001b9c56995293b8c885d7b1c02e52f39b
z5bf36b67165058e72817cc7efc9b4d8853129b38f24e86c32ec88f58200e6ad20b1900dde7b969
z593773f1977a8dcb5d391ce40ff5759cf3d11b5cc270c512111fb3a9aee937fa6be0c3702e0a5e
za9457e2e01eb23f9713b7ce7dec92d425030d323ce90a739b0bcfa55b81d47af54ec1715d7871b
zb537bc48ca8624828e1e9390724d88a4610802951f74d94978969df330e65ffed2d0951615dac0
z9e185fa81d292b5ae207251570434f8f3cbb309f4acd6513c79c45386b1111e9571a20bfb1d0b8
z3ac12175ae258b44d5ff65ed924a3500df0d829f8fa141077428651fecfb2b6d9a3c55137570fe
z3aad32e5afcc11a9b94ab95f31bb8787b3556872db8207cbcb52a593020d631e5ae5a24ddf5f1e
z8773ff5f35c0384e4e41bd8cd63661d95b623d43f852fcf43433f23bf42e1e9bfc712e807ad82c
z94280606e6b3dfd132da433f80e2b088576ff6a48e7ea30b001b6ffd31ee21838832d40e9b110f
z33c94dc2b58b053bc65956089910fa3a806b97c646fb26884bd8add6a260c16495927f8cb7d198
zddb9f3c56bdc63e9f017d1b17f939ab4a07637011843f8739c0245722ce5f9bd39b3cb4e7d26eb
zdd5f0276119a71b6fd4dd5054619e7cf21be62f248e2931e59f4dc1d660b75a71c806c40878469
z13691267c04802751379996faae1647919284aaa77766f2b240ba9983e58a4dfa3038356732f88
z7a7294dc46be235ce1a12d192ef3a01d7c9d50433623c0c39d3c90e9fc389db9c9d1586a4aa7ad
z13c3308e328b92cacfc130aa132a30a7e7b961c0c02a2dde5101473fbd27cb18b1a376986fec58
zb16020f9f0315afc9649695d38b3f9f1affa4c7425e410182899d4bce49068563b1368d8789715
z0f9b83c923e3e10cbdc5f7c20311a84649bc4fb8791d8fdff5db05ceff191d0a6fbfb1e2c0f60d
z152968d6304880d07fbb71fb32a5b3d688d2c3224fc5fc5c0cf62517c1c1b5e18ed2c9f26a3e5b
z9097b881d51d49f4dafdbb40ad7e0bd009fe3859a8a3e1f6b6e95dd46070f2a028099f42311f80
z20fca04d0146d5cdd5f11ed08a002371351868f362cfdac9b10a214a0599ff5e317888aaa13d1e
z200c18223976946a3e7c8a3029c1f86f43d790501ca74bddf0f04984e1c7c343f96e8372fbaa7f
z79f7f147bcc13f56e8211d2b68c4e95a1e999103959c9f12a7c1e42eb591732b17df732a9435d1
ze6a5e8267d64d28a33140bb72f1a9672f30aa93484d41d7989c3c84f0000a8f8584dfe7b4a800b
z9483a9a09cda5877c7060977586743407db9f1c3cd0698c0d61ffd197ac10a8796b02e2a6bda62
z29b3ebe229a0a9aac1ae906a9d86aacf0bb67b8addaacb7af53b1aaf6c2f56a0f2cf4599419108
z488df839222ed75ebbc5f3e16fc74155c29561492cb36f5285a3408125a8ac52ad6f214e041ffc
z737cece09d17b2da280aaacaa39896afd5a5843e1f1cb3f4bcc9e8325c573b79e804dd0b61a8bf
z27c8a4f37b9b9647a14612381d17f6574a27c812cd517edaada517ebedb508b27155b670142cd3
z9bf695d15bdc5452ac9a2f9148cb2c3115b5c869545d9aca0b6a4b465ff89cbb0eb3895da9b376
z32cfde1b724d269d9599d3d120a3e41b54352c633305aef1c9e08c466033ce5c8039025b12c989
z60c27471d37d7a4eebcd17e0d5894ae44d0426c0659228488c48fc3aa2943079d664f53b9838c5
z1fa5051d9e386ec0cdf0f1f9ae0fce98f043dd5699b08fd2598840f1fc4f8058ba90d64eccb2e6
za04a62d24f8494e6dc2eabad83f74da15318b90a6dcc2c685e3cf88348174231c104769fbf0852
za396d276ab07a0fa6188aa782a5b01da13ca95875bbd9273b7c4a25a52283c56a61380b5a58ed6
zad15d02327608376da9aca7009cce31dbe131fc889e34c53f8e7a0027016843cd1a66b88bcf376
zef53529bd27900a7c4a983362a385862d92ff47043019dc5041658ec0c9ef6de9ce791667f8351
z99590463f5c5ebc2420fdc33acb1e2bf039872755cb298867fe9065b4e37f3181ef832f4d699a5
za9bbbe0e53f4d4198f3dc58a308e90796510d0acbe16f7d05489ce94610f07e61ff0f5f6378dc0
z7a1a1c2b1e774dca6fad864d4c569a71976928af53d7e87178271aab937018dde25a91736b3550
zc013e6ae77f18e9170a88dc1a889e495d75d0a876aa8747eecded03c6e985dafc3a64d508e9bdf
z20917ed138cf0e5f04027a6f592120ebaed529cf48410fb30b8d8a59f6456847867a2d78c50bed
zc41d11deabf36542c21162749023fa33ce1f1c69889cd499dd2d1fd8c4c0e769af12e0addb5492
zd422664f689bbe3b254dd8a23847a033f09f51522c042236aba773ca4f4a7ae913561beef75aaa
z07fbdaab1efc375e0ed3b5e7e778a5189405d14987a304093b256d85c12cf6295ab3b8fccf53ae
zb6398e0fa7ea2ddfa635f2fd32c2e6eb764f62af9dbfa20f46645ef3f2accf4ee2fddf3ac04b12
zfe25b8cfb6b46c05b4b23eb4d2835d02280b10bc7255b04550613888650a34e3d6c5cad9d1bb85
z0d686f44eba314fb6f5891af6d5777893ff52e95f1fc6df783a29a9b541c434fb1d11779f6bfab
ze917236019c0f029b244d484209e61426c5445bc0ef2a1f57daf8d5eae6f1402ebed5a3225706d
zb030bc269d194c3bcf5acef358cc4d6d858190c7eb09ff02430474daa4bbc185f63ef09413f1e1
z058f429b64c1ef5936aff3ed744f042bb173b9198a00d9b144a679d46f813e3765bfd648188185
zf31acffb3e1ea2a3316cdb3103119063db86d675bfbd44edec893fd672ffcb004bf94676b36925
z527e005b6e1b56a1da86898f364c22ab999c3641cfb918616e5f8ab610e9d892b939f7330634f8
z9d8e540a2094fa9bb24a1d8476a5b7d03bdaea4834e8bbe51b744b4fe82f615fef74b3c51ecb29
z1ea5236b93e8b49c92700500bb10f6e7439cb80644869e230cbd6bcb3fd3145a1f764a51dab907
z56ca93e62028551f05cfd9be85db47e0d4a9efe7dcba87324b54b46e1ef6bcb754cf08add181c4
z75449b8a93a2e628a53b780052189e1227ab6ab153cbad897c1c49b85e873e72909478f667516f
z4e4e8d40e484b103d9a7c0f486f6e7858153ccd53c2740f00b47664bf74d25da5932792fead9d9
z3ed50e61f4e83202f03c97b1d7abb24f7f9835836a17a9d8a9e2c70e70d20b4a31ebc083a4deee
z649c3d6a21ab4ba991ed47f704babe7d13337eeeae355625f9e71df06a6d579d15bb53fd8d9ae2
z355cb574aecf374c1285e2e9963ffc34fd9d9aa45cb563a2eeb28cb1cf2020746d0508087b4d0f
zfc1caf35355b31a6f6a881598de61608c2c2b2be60c5eef562263bacaac833ad2ecf336fcb26c3
z7b793ea1e247cba802882e6fb5f78795f98092c5f97d75489d08b11307942017a50906650271ac
z48cef63654f45ccf68494cdde1e1ebc2fb951f0a6a22c57724559ecbf0a15970802f08ea00ec16
zd9f7c9ec50daf6d14c0b754b9eff6ed033b302e15c21cdd8d03f1b3e2e280dcd11213e539b8c4a
z8f762e87a05b224caba7006260bd2fe40f41419ae5b61629dbc8ff52d380c5dacdd77a87aee13f
z1f734d55ff09f6488a05b713c4b8c221cd1f37f57faea1b37106e99fc071705e79e8597240f21b
z3044aeae2ee62710ea4cc54ac883402e181fd630ece8e29d909830639023374e1944a54d1d7abf
z43a1e393e03129d8a1ee09245de397e11e190cdc89bcca2843f2b3f97a8460e58e6f35342e5bd3
zbadc87b7a31f13c9044ac3ba2a46345b07de5b22e535215bf81a9c04f5a5e920338e656a4bcdd6
z56975f21902c35a8a3c6d583e5d234a3d10cfda67526f8b0fba32836b9f17fd631f7cbd13f0525
z7063783b9381cef2376e76f187ca8f695b233ff049ebffbe88d570daa94fadaa80ce0bb50f6b57
ze2c025a6d47542ac9b8a949f1c2243e8ffd8171848176ca28cf46fb63dc0a30d7c6a11b138a889
zdd065dd98a34f7f9a5e13f39ddcd4a9a49b1388e149f160aa5f63f188ae7f3d18a3323dd6de8a8
za713c7bc5bfc78d06a60eb81e4a05f47db4c8e68537f5fdce9242be54b740aa697fa587626fb48
z81fb8f20e268321a95632de43ba6ff82cfb9209971ff82c51da007b11011a2345278f3b311342e
z8ea947d8bbbcb644d40b12035a54ee7296e377e1a9def0b9eabfbc5b8ad0b63a15edfab612eba1
z7d253c2e1a579af950e92528d1137e2f63a82ee888955558e789372859c9bb28d5ef75e0794723
zd1f3e78828493170f6e267d7b5b726fb56b38ac7d4b8c8d21db0f5be73699a7b68e5586f6a9ce2
zca3bc85a25ec9f21a1a6af7886087e828610814310488407dceee0dda1e15885a79a71569757dd
z7361c560ab801d5b3fbd20613cd44f06b4ae656cad0d3be1d4734532d017f35d4c1bd42fffd0c9
z45d8eb578c09385e78fd350260f0f5a4f0221720e144677760c6e03eb00c7bcec98e00c817c80b
z56db5ebf9a324270d2899016278d60e3858cbd1873b4b0f65c623849bc45fb25e10971ea9c4d47
z6459426fa9a8631b0568ebf5aa4bc9a59505c94c92c231fcc16d92212bc8ec402023cb5bc15679
z291e429a5c16bd95ea0b6304e89fbfc15e198a0a99b73759a8eae581812eeac11cc2fc9b340c46
z44462eacc37fc3176f47cc79cb9045404eff2b63bdcb6754defc0273a0ed1738876581d3bb4317
z43fa554eeed27c73b79cd606ce923763ff3879836fa20cfb5610fa137a08bed8b35c696ab78ef0
zf1a4247cf13fb15d66f76f20249df8ce16b8c4633235112e97a2f42c2cc6e693738e73ffaf0f15
z2e4cc39a56040dcddfc94be5bb845f19e8792639a98e501c71da2f87e5c33467c4062139e2d1b3
z68dd817a91b906ee9fc52f39d25342f08a9512157f42ed58fa257533e5a6ed675110913f64abac
zf4ed1e8381d7dcbca2b4d77bc735a1d57d14276ffe48183f77a6d84fae3ae25388de94a03c129f
z6d70f4d41e93105b86b84546eaa1a890501c785825af29e1707d3bde722d79a76af5b00f58f7b7
z14840c44ac2ab18925acd7d071ad3f35ff86458575115cea9ddecd4a1eb77890d0fb4542503ae5
z72ce116efb02e5ab77acbce07825c667415d5dd5cf74330eb35e2531d8fc138de57ba6b54b8816
z5ef2e2292fa0d804fae6ad1bf1ee7bff0a5824a0e95d1c75503863ea817d0e9567ba02f30e8927
z5e05e347f857abba1aa73ed700315d0b7a62ae8d35bf5e853e8a97c7f79c944d091b74183ff996
za5d424f7ecaaf8e35e67ecfe248ae4e79b2c9991b7797108ec9523ea475a2ff801ef82ab2c5d8c
z86b8f2ea11cf49460c76d2789d72110ba1f9b3babc5ed9d669b33689ff9200ff3b5f68f635ff41
zcc1e2d111ebf962de72c892a9eb8577012bc725e000fc819c1f8693fbc861be7782f8f1c679778
z09bbb0a040b4b8f7864524728d7e9f24d57e32f2945ef37532521beb0aba70326b7b60554ab0aa
zcea400ab4a9b81cbaaed61dc14d380fcf0cc952df28f7d0d7511334d5f135ff8f313c9777ba89b
z4f9dd54c9f688dae4c3533e373c1de7b5906b688602d8de56a319f515566ad57da1738cb7b37c2
zcb3159b5724f4b096f967725a912671e4288804de12a2eacc827824617744a25418d069d6a5349
z1512e0c29c7c5a74c21ddbc40c8ca59848eda0e6e2087c6a41df1fcb6380c0f063ef7a4a18b9d5
z7f6e1a501efdd3f23983e093191e953fd0d4238762dee9bfddbef50f040e0f2b676397e6de29f7
z3d3699a4f31d8663435857a2515f4a290ba95915aefc16823df38e2f25a8b06527d61594b209eb
zc99c8c7177839c8c4b5a9f7ef78d9eebc92770609a50b1bb7aa3ee986332a3d368aeeafc709520
za72a82f19aeba47cbdbb70356f6ed4688c9265e90e2efa10e368c8aba8f2465a616a16b6b26b5f
z1a94b085d66e39f5c4b0befb9bd8f07c57094e6981c7dd57a2e9bdb13cdf73d266f57197c273b9
z640b4e46fc4258e1fbae9258f2933f5bcf45f1853e23c2afc85cf0d7cc6f44f7003dc1e4bec02e
z333d709789c42d7b4951f362117bc7e32af10cdb7b65fa474de43ab96ccdf9def4a9b8d3dd8d34
z7d563f683f94c0f12b4a84465d14d7df767f7b071e1967a5724e5cef744979743f59d384996606
zd42941db0aff672c8c8862cb5803140bb2d3c7573688c9bdb2ab23a29b1aace2e9c99a938a00cb
zf55325d963b31041c8ecd3b6d75deb4dc735734a05366fc35a793b7b7dea7e4bdc9b1710752e5a
zbb561252075ed30693a2f7bd9f4610bb575d6bee02abfeafce1d049a3f430fb15b31e57852ef3c
z14e457f4c1987e142f9d91e926e919785cd9c08980a1579a75dee12c59bfb0ec848e55e0886da1
zdc77e93d93128e5401e0de8a62d2fadf45613ef0c6ba4a93bc5c9b030f5f7554863d20d99d18bc
z7356b5648a9844df9eae13e97ee10569db1e021d8d76758d9664be0892d2ef08cd08debe6712e8
z20b880f76d24afaabd4befe97d603c2bece67fcac0392ffbf7790ec529de553ce92f2b0cfb3d64
z55d5597c8d1e2abdf7d34627e6a064a827f81f202126a5c8c330d4dc4470f8042be59d90a94153
z1d721a8a5aaa1a94121c242e29663ced361010cd932febcc8add119b47e9559aeac4c3ac374b21
za163a5fe514d464e0b1d013f613ebb262517659e6b00bdf94db98871b85442efff7aa8f157ec06
z89ddfe22a530891dec791d18d47737bf43d4c797d481e174a0c27415b3b13cd4fc30fccc31d526
z8cbf6fa68b895ffeec36da908850bb04f8db084734f9a343ca253d509e712cead71298312bb574
z89520cf6d5e648f185d4dd636f4a828d6a969a0a6ae9b93ce6a71211bbaee5025ebfcc8fa4176f
zd9a8463d0ebde9785a8fca599e35610d40e42e5a1b2af2961d47e14e3098c09eb835076b282f0d
ze5e9791fb2a1a2169fd781fe503d1af7e7065f0f0b17850024425f34edd255848ca451f9f8e3b3
zd37ebc99aa880ded6b2696dec49d373c0fb50531ca83177a88f74454fb4db1e6cd26ca77939ca6
z6ca377fc77064453b49e59361b63d924c7e297a293d81305b9caa3aeba5060ede74310f3300b0c
z6140211bec3312a32d5e28e50fc1aed529b32ec3cc60feca32c97c0252db1d94e65319d7d9bc60
ze0cf22f0813a95f7a91b7d8d00e08ef1c32274ba099671a0f8ae9c6f8bae2f66d563136eedc05a
z3495ec53fd4493bb9cd55843f633ee431c12e72d36af4c783ffe2d9284d3aab42f5674d2192d02
zd6c32ae21c828d3c4ef39b7cbf058ab5dd35b4756ee8e3448230d258e7796de84d1c2f0b84f79b
z6a106a37511b504e1c07d8d706d8d39bc14e173f4bb796dfbc48047e7410ab737f86aa5e702831
z9fe1275ddf9b288910eb6576efe0d6ac2e4ee044176d4403c5f51f1b6945340b7c9dbd37c9299a
ze8025c77c964e318d2a84bf4071db377a0cabe7cf59cc751cdb0b5477bc80f7cd10f77faf46f52
z1e84fe612e6aefb0d1721ad251e28bd044b996e5079b4a2994fd1817f2c36f54daabef44e8b31d
z0550e5e875e1086659f1fe5ca5faffc748d9d1f305f0d72a42bf810d1f7bd18aba12ebd60e94ad
z578a8ab47927e166f626beb6ae232c7fea7c70b35a89c79372628d73e3ea4097fca08106bd7f5d
zff07e0952e230ddb9e4b1509ed9d72e048c13f56dbb1a7d491d44eaf1b7bfe78cd00fec14677d7
zc810b87147d09b972f3d5cfbfaeddf126c0f8bbcfd54b8a14bde8b8798949ddbc413d059fdb068
z3c6259ee33e0bc7b401986005db9f65231fff4c2448c8f35338d14d199d6d82455b486a4c8124b
z2edeea41ca58cb15cd337cdbf1d3e29e78a00990a7c2f9950997501deaf32febd9f4192785160b
z44f3ebf979149b61c9fc787b34e9e9d6d51b1c3e35771402076c32e4d8b37b8740d8203d7ddc49
z9e0403f55e4922debfc7c5427b92b6066d90b0eb6d7797f9a9d50c9d41e489377817db95c3b0db
z757069d88bd38b00d5ab56c27cfa4c9e3fba45a86d435a826fd4475e666de6f2dbb1805094a06d
z9c3320f535f910cc55e61405856a0b60c3ca3a70fd21d15e3fad6af6f7c11a995b2a6a9761d17a
zfff306f35ed4486bbf865843521cd792002209788fff379fec13d335d166e8f4fdb662409f209f
za40d14266c22619a2bfcf4bd2f250d63015660b99e7dc6c2346d645df4b8876441c2e43b4e7bdc
z2d9e93672968e955f1623ee35641fe226376ea898cf4bd7f2500a50e628b3455d163d9afb983e0
zd8f7fb369a68d9baf4b335bc1f2f4d752850cf4c57a47c1a29aad395e56d7ffc956b064d621b36
z867b72a14b6bd7b0f34881e6028af22fafe76671705331dc4d0c50ee542d1990501df08b569705
zef41da32c4011ad58c328eb7acb06075a1c7dd82211b0c98b41fbb3d82db88c531565a5d97253e
zb547b7d1a906355f3bb629902267fbca7d8da4f71fd713394481c07833a2c771faec06a6f5d7fd
z8d7418f76369effe6a1353425bcb00fc570a8d550a0d61934e634b9a18e12f7785fb92b3065789
z6901ec64f63f8e4ff5f73a984f89f31b72486e0cf38809a9680d8cd09c55cc1dff9fc4f2e528e1
zbd1012529a44b3f655d0fc4e5a5dd9377e22666c618a30d4b7686d8b57dd0ed3a77be37d39a7e9
zbbd45865165723275402fea3ea9f7ffa76a180086faf55bd40a6d53ae156e484b8ecec0fc35bd3
z4ba88ad2178d01dbdbde0bf47372d339400967cc1d1ab943383e404d82a54093a00677121156a6
zfa4a9fe85dac775c09f226105c85e24d9ba9d480cd3b3d09c14651e06ba67832b63eaf1c81178e
zef2b5f92d4d3b7f488c044f7a2e354830d53ad03a800d291b7c092b3daaae2d122b25c56fe1abd
z039964806afcc5bfd9b556f00ba23a03f7a73fd6b2725f9927679c577859e739a5d732d2cc2df3
zf74dce256e77ddac8e224f565a6b5e7451642a7e2f32e67303dcd7e3966d8f5ab2dfac43e212c0
z9a2f12978718c79f7340a98d496fe05b2186061f4b2069db4283f8d0a42a3ac25a80a9d4e3b557
zffd394ee6f388124ff391ce4b38080e2124d92c2c21c104242fbeaab44eba1cbba94de08de3e90
z402125767ab38b94af97e897773b3604e96be0daeef9f5092f84f48aafd6a4d0bf5e7db7d9ea91
z4ccd69c47e81c7efc3f319d59b47c6cfcc3ed7921fbdc58c527a511dc0f0a836110793877f48fe
z96c174908a7d7817d769c9c4aadf062a5b324ca5cd11a8b0742c58809e91e201a23cf75b0b5895
zae3698596ac4edd9547e17d41431a7026d3740c17e39fab5114af9e8139ea938ff558c755fbc6c
zc3b85c31cd8bc2200c119d6a40c43303b366a6416b2a57136d1ea5e6ed6e69c0e436221d375bef
ze4e8394e88bdbe269645b96a3e6c79cb0942ccefaed15ea241951b646b85875b60e09411bede2d
ze367f400debe660511d79dccde82072d12138c5da12586988de8f464e6d24f2f033932ec9d3a63
z4df39ae3a5b9d2aff9b4153f8059db97de2381fdc494b8de261be0fbf435b43967130d23d9dfee
z9d3209a38f6a4e75272cac1337d758af20d24c03d92c33ed9bb25c44412c6968f33a11a86a7971
z5173406a42fe9629301483e285f60258bef0763dc08eb3eb5ef44341d6c5239fd9ecdee713851b
z3e76a818a7740cfff21d657d9ec7c186eaa617b9065aea7f362525e1006bee1613b19f7822ece5
zf1e5423b9d99c17816b3491c430dbd33b6b47ec80e8669a336169aca8dd19718157108e28eeaef
za79ee255926f69fbc3919c071f1fdd9b35680f2c76f5fd2e9668cdcd9cd3889eff85c7ad4321b4
z78f3fce449c78d1bab5b145fce22ce828c33f2a80407f37e610c6484d1d7f69b61fa4bd5c00e33
zb903f5bd81616ec725080493c3c3fda5c8d7b7f54e60cee42f77fb75b0db3c115514593bb15989
ze81934394222c3e0f84a5bfaf8b7d4012fb29f7fbacb174ba74eeb52b327b692f66c6554929251
z68983a332b5b826f28fc104254c54a170cff82195fa9e7567ecfe074289d45633ea99053b78ef7
zcec05fb612c89927c839c7231a96565b2f86d8133d19359c50441d28e9ec9f0534406ff04411e4
zca5dcba28de41b02f323fb8c289e67eb520a4ff09d98c649165e541593fa42d820032e8e30a118
zf70d7766664a7694633b09d3c541350f124244591573e13f56d6c3c6a1428759fd51735211e656
zd72683b1d4a32e25c80186bb227f3e2f35a96c66b08ef1be8e0483413de8d3e690b8034c07efdc
z7577e322a3d2dfd0ea264202cdc63bb0c98cee7ae3d34b7d0946a183a50cbf908bb12d12c962fa
z0a342819b8408d28d72806f19909f3a8fcf6959f4676973d4f0882cb6b746cdfb7affd6cfa30f9
z64670f9ad3d102e45216078ac7ccfafce756760f2bf2bf7a26606890c78ca452accea4573b935a
z02e10275f442e6f79332d48b92f954d9513b38ed7c54353f6c7bd385efd17c9ea840da2183173a
z3782db2d844dd6ce5f66ace40e486eb74cd1e02a5d8c58cadf518910b8670f3d430ff442d0b707
zae9741c048b8309b452eed86450557f0a3597f457bcd4a8f80dcec5a01daa481fde249d920c87b
z7fb44850457a0ded6927304f3730f1f2d66ceded344d964b95d0c4e0f2d1d708bb4ef5bbecf039
z8e990aef8602ae5c3c49c46299b3986faae00f2c05608e8d233a5d6dbe773cdb19b43ba82b943b
z50b7a7ab1b6856b54a83a9167bc49b4cf9702a462144b380075bbdd94c391d892942a467d66d29
zb47c1768a7f87243fc4dd480a58a465b3d2e398ede28a71f48a7d08d22c61d63d669bbb54bd8bd
z557b1ad701e3f7e5f7991dcd3a47c8f5fc0a1e59d0c6018e2607cb8135c8c2d512c354c315b31c
zc121affa0943e7681925fb7b7495074a9ff3ce4bd732f0a2aacfbf448170efdb5624fafa9d3ea2
z7848ff0b1c099ed2766985f831794f7ae09c46a61955aa47b27d3cfd02ef24c9fce89c90aa2d0b
ze20e92e889109620b0f62705055a92c52fa8296641168ac1a55daec8c2fb11fa9c97f8e9def023
z7612259be363286364ac1de70c7c818b8eb8454e3f87ce14c0a34d258d9daf1b6541671cd97bf9
z978fcfe35b74112398be5efbd0e587e3c25413a44e47ad6dfa4f8b915ec4747cef8c3e2c545462
z4f266dd6889d2d8e758dd010d69a77c433d9ea6956759967f4815b65e9bdce4ce4b82f77770efc
z2207b757b7f0bd3e6d153ff88db196dcebf573200f58311c1d615a40e88b323d84bf71024a5dc2
zfbe2b133a50fcf62a03b6179341391255a439ca9b4d682bd2ae1abef99c826cc6701f847028290
z7bcb0ff1fa1dd361c6d1d4930eb2e108135cd9ad601f3b6f0baa7ca73ba623b8edbc0455885e79
z0c5cde9637c00e421bad765f4216ae033f0a19cb1885a10a7bf0643b56bd2b640ee90357c5b132
zefcd59302b020f3c076c7af7acc4757f994bbc745c27092ed4b335883d7734fca9689cad43bab2
z57568e0cf268e1c7987b9fd9bcbf139fb9745a9edeeff2b763892e5e7faef704a94c3c8239b29b
z04d573856aa6acb3eb2b46377adf9957d0a7d0b71c6b4ab90172c7701748de40ac08afa8d7302e
zaa7d69abba4030a7da7885d7a5f462600915fada9e3fc96d5cd0c9547c0f7d5dfb776dc0b71f03
z3aaf95cefaba6bfb8e8f1567d8380c0fe335379cee175aa72dcc050e13fe66ddd9c6f7ce76ec32
z46089baa4b24301cb2a82cb96acdfba0b8914a375d3d66ab691d21b1da8bed35438bf5ad63da45
z5014fd4f2b6bbbfc20e0999d99e12728eb319eb187200ff4e16d7b787746e60d5d4db308c7e979
z984cde57e92e71f21021fa30b2b79e88ba5530aabfab66dc714f813d56260204b3bea6744e6001
ze01393923b3f74e5eec0233be9b09fb95ab6bba712aac4e03d1afc273d137acbc1c4391333f9fc
z4956a0ec147c4126cd972d82f028b54812a197ffdfc30ceb3e7eae67f4d8b636b44618919d2026
z38b87754946903929d5708182b62db9c7ca74c583cf80aa7370f1acfbb21ecc11af59ba85d7275
zd51314e3b9d3b6bf9aacba77691e10eebb1991adc6675601f9cf8ba7ef8a7dc9adb73353f8fb85
z8011de07313ea10476bc8f3e029ac8121b5fae0ee0f99145972e8a5df6ecbc85ba73eaa1eba3c1
z6603ede6296b9dcf43283b5017d72048b6118d3c2402c2e3e8567129dab2cbf357b4b6d34ca8be
z516a16d6ac614bf70f6caec75a8156846bd1f9190e104957cb370e44e787ce2771fa2f28bf08ed
z56369af016d4742415d8f105d29636117f0bebe8111136371378c15d62a5d78d346a0613d3a884
z50b0fb62772252249cebb47ba8bb4b66936c1a6d4cac93e35a50aef394c731b8976dd94eee3a31
z0e9fffbbbe3f38a3ecfe815f2749dd269e57028a1101857612e41933b1be0957fa7138bab7eb0e
zfd2b8a5a9bf3103ee56d803119d467294b2bfc1aee70357bc2562f4ee4b34df74917399dafe3e0
z810bff906b68de8c0ac5a34812c7de3c8c7c7fb4ea22f7f7a40fe254b75adbb9f8f09c283f4d55
zbe42ebf106a86219fcac1176f4b446e566b286b91aa0a674ecf6cc3456e8f31c5dc80f6a5576cf
z1645af855d3f5ed367ff7207213b709bdc52315c8cc39e9a4a6f6e7ea6ff812f95bd9f25263dde
z78524519292b5a5f4ebf6748529d43a9c1627949bd1dacba5d1f4b9f795c7fe4144b074f957111
z9c8524b43308826b7aaf2dc3b32a4dda41faf2c8166b781d0b158c819682fcceb7644466ae2d4c
z891d1cd6c2d4f6eab4b34633bd8375bda406523dc3644a6d5363161c690472abb1383999da8279
z69913cfff38c79ac3372f122be1bea0e1fcf768691655dc037764f88c075790490ed679a41a5d4
z57c3728dbc0b3fcc3ca9b266abcd2f7c3efc4dd8d1505552803b15bb745cf15502188d6c5a2560
z781684cb11424dd117fc96736c04b915633dd802e2cf0eddeb909fd4273cd993a49034fb9632e7
zadd4b8379116ce56a89dad2df4d36b2f9251279f6eb05b41b29ee98fb1f1c6cb18c72c97066ebd
z9484f61d1ac21a7d69b2cf8489d2c1fd2e25cc0003b90bcb9510e5532a30ce1c7d9b436cb1587e
z413dec4c4b7b50556020c694cbcba1db17d17b9cab71ab5bd251b0aee0700307050571bd9d283d
z267390eb2e86300b1df9eba2f570d28a4aa0fc3b6c4ceaf2dc99df45b571a1b2e828f114ccb240
z2c9494b4f83c7a8acd631145a19f4c811f388b0a2e64f12eaf89e6fbfc00c6807f16d6b5cf2474
zb62f7afd40240113b595a037c57ddbccbe526d1ed9acba685c1f05d53289087e37a8e1fc4a0ae1
zf4375ea61c8ca85fc643e3e72804b33e8dc1bc4561053be43453a1c27f1e1d4a72a1b0616c9696
z927f6b62671cc5a108268cda40e8490f7fff38c1d0a78e9111ac6ea63fc626e74dcf1dd3b73c2f
zc3cf3c4e6185e2ef218b8d9f0aae738fec720b40241d5dc552fb0bf88708f02d22f2a4a58d97e3
zfff7a1cbaf3f147d4f43bb48ffce60441461b1f12786e24dff45e5b1179f310b0436b68d6f9312
z19324813ea7327801e2e2e66b75ee6768f7f0d0ff498b9301f92e3bb594ce43d307d3da059a7f7
ze48e3d379d2425ee233d952b7a32a97d63863a0ace4e60ec7f8a566b62cb3e2b168f222dcdc813
zebecbd2bb686b3274a80bb9cb7e01668c22ed460faabe01192f485420add8d484f2d2f5b8940dd
z6965d19d58fa20f3bd0e5a861f11c4461be66c847475bb2fc60245514319856a2985b17665b208
zdb0e9c02d249040480e1bd5f1a5e9818029077a2371803b797ebcf47fb5fd4c8892e84ac50d596
z9ca0237a009d26488a0712d48d31fcfeecdcebcd5d7b9d74ea437b33c90b0d52b2955c136723a0
z19124ab72f0ce4039568f386ca45ed7a5e0b6524a0307b10e5f25a1cc96de23671b950e26599a4
zd6f6674f0b67e863d4416e0d16903a2e5b30aa8333904ea75afa30c54b9c809ab34344fbb210d6
z295a1c0ff6f06c0ffa03453d096686cd42ea8157f67c3379e5f19cdd1e36146c235dfed3a0afb6
z1c247f08b85eb5b484a79d4f82a25496db0d7bf9539e438fd0757853f4149b96d02a315debcf2b
z2c4601b65bc478de4befdb96d7e860bd458fb567df04aed4c4adff1efef8741355249519cf0841
z4247f07bdeff2a6019a5c530b3ac2b83b5bb3fe7dcb563cac6654055a1959dd1d151853ce13cb5
z568819d817798a60ba080423bf1ac30635af159c9020bd30db2999b73ec3e496aa40a9c5247185
z06feab952a962015c73a71cd451783bd3b18f6ceea0e20c7d7bea8d75293c9f1fad39323e00201
zd5a54bda4b5c034d52982c5b2eebf17e8ff3461a6c76b33e4994deeab739577301ad59fec7e836
zb2c0f2a52e791ff67cee2c1c43b08f30b03a47a8371bd5209bb2c61d1328fa1fb7f308e8e97976
zba7a6b43fd3459b05348b73a4bbacc36391f8e066fe388e77be69657508f1703a56b91bd636e1e
zba6af176b433097c6d117a5c78aabc6f755c9af2b16a6d3a6e784551bee5972557950d2dfbf145
z5417024d079304bf8c8db65ddb0e6dddabcbd1d78cbfa152f5e703990b4d304868a08c4fafbb2c
z2c43ede100e7e97b1347a9f46f8795a2b852cfaf3f25c20abbf56a7132ab634e845b3efa0919f0
z7070db5bb785939279bca8cb05903354c6fb18802e570743a9aa1228413334525f50b1e709fea1
z2d054921da8dfb10bb61abb06b9c2d54ef4898cde1b250b4cc29f99a1e0ca1b639ba48dfe50e78
zd94a0ab8c73ef528cf433cf97f84fba6be5c3149bc986b9dcccd15f2535f2f124b2c8e181d6b4d
z93a7409f019dc35bfbe73975a85d3f43a94c4df3f6852540e78af7d074656fd589b05a038af7e7
z1aec590d8f3735c6344fd183be7e4cabd4edd31b5067322de1f5a0c46c1fc7ae925265472aeb4f
z68bb7f642a385ab038ca152fa93a8b13ed2354a5c2df1afdda044ce705d9022ba34b9f7ab5cffc
zc6493215c0133b31338a727855dd0ab8d11afaf0561288dd9c99ad873d4f340d46623925d01755
zf8622b8443dac8af71cee824930fd73224dc1735e8fd68a6aac28859de690a7253fdf2101f9e62
z4aff2db6ac9d4fa746df2de99ad7bcdc084fc46659805c62959f508c89b68e6fabef920e30196f
zcca29da00f584127b401d5a7bc3ba0c521a6d77f896251a57b6493c6d96336df7b86e2bf3421f2
zb87d00a970a06a0d8076593809ed1c79f3ded43b0f36e730e7e2b8ee9b320bc94e5dd8bc5f751e
zf760569074eb77f214a5255491533c0145e667bda5dc78a0c1914b1f9969fd1c24e3ab7c5d4308
zee8d73bd511380f285fe5e74d6ab5a4477fb9d05bffd45778af56ace6e6fb425f808a6e8e12978
zcae53d9fc973df5047fbfa4d38c803b6530e44da5aac15a3f39a3bdca1d59a8e3c41046bf1183b
zaab6b18c9fe4df4662c4aeda7904245ac183c2f8a72ebe44cda00c0af1943a6505966ae7076c68
z6ce8f593a74b2d362d4dfa26278b761aca46d6e78544ab55f68e64782b94e819e4db4b94bd4b50
zbc2d91e11c650adbe2d2c5b6ad719728027918332fb756b870f98fcc3db191d260732d62c517e3
zac21c562097584ac688815a387b167d9c21f5475a73f0a539ad618b59be38cbdddaa95fa049c6b
zf1ab091824248fa18357f7d12cd61c2b01bc0293c96e9fc48df042e3d77b3efc61c3bfbbfb5c0f
zb70a203cb41b98f4cf0c47a93b1eff913367f2e5967094c4ac41a4969d02dc6442a93dbc75c8f7
z4b091e06fa9d6ab56ec4fd45128963d0a6c253eab1ba214492746a9cd1e5a8f888dfb6ef575e08
zda41299a5180c4e73e7a21b9e4d188601cbe206144ef1b4e20338a25ca4c7cb3e0982749e64b59
z69e25640fbae81d035c4551c22ac720a4a03ea4cd589cf9f1076ea29b70c08eb87bce2ab193b64
za435e888abfa8d460c21d0ede95d22481e1ad69f5e8e362e4a52d4ef89a02cbe7fa6211ca4615c
zff8bb3efb21cb0522d31fd7c9c2668177d7778ea3ff0131063f68bf77154b96640d02ca9f5dca7
z1b46f6467a4c5faa02efe7d72219eb47c4ed40a0cb5354ab7c1a522cfabd9cac6fbf1813fd938a
z2c0eb0940f7cd829bce8df5745c275c9e811f4329e6ab83f8cbfbc0efcf1ef7fee326963358343
ze0094db75ff6c6e0d86602859101525b1d0ba199bc9f8a28c01ba765adaa778d72eeb5724a4f78
zb7206e4ff39ab5c23753d33c9acebd8e8dc360c13121db7080fc7d5aa85dedb01bb511e0f62a6e
z835d7434b0a60178cca54c875f59fd3b585e5bce30baccf3e00185c51832db95f9d231bd96cdcb
z6452fb395acc1a7d30e941b876ef5401eca29c51ff4fb3f5116a233b50ae0dcbf6047d00fac088
z39284e74d6fa2f5a1e6b6f6d1a9d641e7626376c5f67940abe1577b5efabeed5b2c8201390cb46
z2314acacdb87e9ec3ed21cf035865be94fff4425e35a7c27d7d34731ddb154ab4cef21017e884b
z7e3a0b19b426bc96428520a9a0fe5712c14df33d791237d130d7e37828a2abe4b1271fe5e9789e
z72c68c94f61e1e9eb3272deb466f76ef4ee4d0de9f726d3bf6d9b0508dafc630e0ef4039723c67
z16e437f63040dde660156ca9c8558f92c901132f5699b83087c2d51105aaabc19b66f21b542925
z12937fd78725f861ed3c15a8af8ed042546d5ecc254b14d68e7252459b2cdef7cb192fe0e6829d
z74ab31b1e5e776546b393284a4fa7b4a356f0014e8214eac31c9b1e08c51b60b2d0bbbc1558770
z4fc235900a8ee580a3799433ff55dded727574747ab432362ebd3e769e5f021b5c4a88b5329764
zc108f969ded59674190d3877d8f9005f1622a4d1dcfcd2b66e04c909ef11cc1ab083b4fdfa4a7a
zf83839e9c5c7586c97d6e096b0127ab7fc935c3be16fb60c5793f5c1eecc532dbc4ef21702c084
z2fe658d8752bd2f46816fd661bae8a7226802addc99e8b65dda3c1580a89bdfbf75feb4a9b637e
z0bc990399732985b8bc079ccf96e59d54d1000f7e7fe4085e7c51ada900c18b6cd03dfa0f1d6af
zb1726d560895071c70dd7b2ef1c75465000739010df8eac35249f96302f98b410cc2b51b3782cc
zbc5bfeee26d4c6b81047c7ccaa710633ac7908852fa9c3c62f91f44720da285f12ee1855b57351
z1199fbc76165ce2d132ef46dc4728582eff796fa20699ffed8a2cb66f6c0681f344382a517d8dd
z2ca89e950aaea43d79e9b230e2121dc400284858fc919d1ae551c8cd8893446caf4e1db7bf71d3
z11c9fa983684664d82d8756ee0c9906eb8fc1b744b5c0c217da6e8419b8676fa518acf11ec0e00
z1e541b9795c82ee265830d5f18e9d198fde92c8ca72e206b5c695bae9a3653706c914c662e4501
zba0be5ecf49d2b4a7fdb4d9e24ebdc7a82e0c8f8dc25083ede02718d5b67e17e32b7a600af4e2d
z95428b0a8fc242e4673829a4b353d33ea7fc1666a9d166d055cd680cc760abbcd75b64d3fd1843
zda021ac9f7e12381c5c2b498413396f9e2496243aac48ecc002c428fb5b32ba21695e0639c5ae5
z2a11420993b13fa8fd88bccac41da017a0125ba7ade0b8b42f8715a89fe789964cd1b4ccf6bfa7
z05154cd9cc926df09344077a75ab941307a1b67122e630c2658570a481b5edf2797b9f4fb411a7
zf4c951aea1d4e2bf8c296821fc390510d43b50db61270d6472f1f65bb42676894e0bdcc7114d57
z65bbe3135034d11d3799e31a41195a4c0d9e7e4cc8023cb2c632eb4f013170d92b52c75f67af82
z8613a93530cb91f23784d2770d4de888cb6cf5b40cdb2858604bdb16856593bdab2e81a1536199
z865053c37f74d56b13dfcecbdb30e566256a6cff718cd85526bd416e1df7548d9f7787baf548b9
z5f4a27fb8f3ca37157d67cf8711f6a8dc85affa68b7a0905af8e72984d4ba46865af50cca41036
z3ef07048fb310f5c67c2fe4a0522219ca737c9040d085c74ad6ab30959e440de95f2ebce3fd670
z04faf0a3b207162dbdc35eaf2d4e07fad0365d4319eba3f062079ce44f6c3df1bb786bb71b3810
z4c96735110f23377a9121d80d4ba44c3bf76910d51f318ab0013bc233c14b4d0a2ced4f3aba2a4
zb3b9bbcb9bd3e338060e2a488e8b22c8eb0a130839eea5ee246ebe70c778be46d3ce16dc08a8f9
zbfa9d6be9cc1672861375b5623df3cdc7be26587eacdf25917125fdc360b867a47e9142e8e7fb2
zf891f768ccc3e2b1838821cc98edb5698928ada9cc9402eaf33bf1e848050a5b7cc577d18c347e
z06ec58f15613e01a18a63ec2dc8845479335ed735f550d79bb865811e17a36128f6e0cb15ad5d6
z34e242a0e9d031a000dab44bd355a0f2771c05b0167bc9c4a5c068c7edf28191cee0001b18ee13
z945363fa2290902b76e0a922ad0c5ffec3c76a54dd40feb5693c7f9bebe12a0d3cee4a526e17d6
zb45b0be397e35a39f389ce81600385ef676c81e43ad7e20ad5f19c36fadde60268d4e7c7cdb1e5
z15f46bf708dee3c7ac90add0f1530275171a1750f05d5dae80498e99436aaba675a6b3237ae1a4
ze1f2d26dbdd8c76237c73b3397e5dd4b8e54095eaf98631ec589e320c03795aee9dda9e5ae0f4d
z0a4fa7ce9c752503ebb1bb8a4d6af9fa9417aaf4a8de5fa984bef4798cc85ecae3265dcf597eb8
zc9c9eba602d1a7b214e2384c155ae67f3829d4801b74ba53c97ac6fb5fcfbc6507b6579ff5e185
z298c74643f98325c5642e6e25010162d92c5dd40056766497d5aeb6e5b89e1adcf6e8a6eab8d85
zbf5d0f624794efcec7593adfdfc0d28df7b5e1ed02d32531c3553e30e17d53fee7133bdaa2a55a
z96d6eb0c901280b772e1d7d1b85698e40a7ea173ee84a75aa3675bd68a62737f8a6265792157c1
z3c735c95a132a7a6f255509c0b4f21fbe8127945fe5956df47be2bb2e322bd48ffdcb2643b7145
zd5d14e73af47d2ada4211fe1fd4975646d35d1820ee14c808572c4d394e286aa81d52b78c3f654
z378898d6e26a080f6085a92aabb11587d057d6fb0b48c951f7d711b251a5a2eab61e7203461d61
zbec971f15076362d9ece2ae5ad84671d7fc8e7c19fc5e596f0c8150e6f035913478f00db83d968
z8b514f7259f79b082bc3f1a1b016db05ae26aceceb48c101b92f7ed645e50b93ca48b935fb4617
zf057d21ba2c81952d1f158c046a3ab2f2eb140d9453f9157059f3fabd21b1f1f58e4c4c831be05
z3c6e692c66c527a8d1fa04685893c18210480afd146b1c619721bf712b7d0dc40d64adcec05a72
z5163b2ff81d0666e239ffc60e6791c3da7ba4fb4ef05361547c18c3a9019fcda160941721cb474
z4a07b3f3ce9a86bb7693b326d3460f8444f87b9f476719e7e9e3af8a789c25400ea9007538ff12
zd56e8cbce45958244793cf0e8c49a485c8a6e594f7f018e1583158067d1ce6792cd3034111a878
z38fdac7b6e60265c079b3bdf7a8bf9b1eeed235141221722c3c2216bd7a4083cc6967d235c00c5
z0665077ed7a52847a2213f6cf11a6acc64665a87d318813def7585217894df6c48362789383738
zef99fa6a808aadc6bc44a7c998b18739fc8e66738f540cdb2c48dd954ce9632efa5383f897689a
zb547d8ad8d705b40f1e08ca05a1768053808bab471191a87ee8dcb9bd401b9fd6a951fb70dd778
zf61dfa78745207aec44c12da7ca99abe3f47a4e96508a68a1768306408af0557df886c983ccd3c
z0b193844d1a6ff37f9e6db322ca5c4dbf76a45e43e847972b965c4f378b29af49e62b2c97028f1
zece62b63dedc24377e890bae52e27ae3c4242241a6b980f26ac9c1d310a019e760d5df5d6a23d6
z79ad6a31a4dddc877ffde0a99e39ee6adacb698d9f1643b595718e635f6d63ad53d710199ef01a
z441a375abaa8829ca0838a76d066f6b4e766b88b9cbae83d102238748a421e9a0e96ec323da08a
zf5ad4ac532fcf729b0a6e8894e5562cb5ff2f4c77884b13b33d7816d310f60fbd111a60c80a7bd
zdda82d66489550560a4e72bb836860aa7c7c817c99bc8d64b01a09f6e536334ff6f3a4a5878447
z57462c1066dea30b60e94feab2be280d749283171958f8447437728325b92f6c3b0cc186d9a25e
z9ccd4b7340d08e515678618195826e8934fe82ed6be35c505b505456b7c560e596782fc5274b7e
za0e2ecd5c5a584b97257b41306b43312dd159712d567c5490f349b6ceb03e351b3888a162673d2
z8b1e8e2a5443ef2249d5fabec20942553dfe3e949e476a3dfc73d177bd213841e2a4469c5860df
z5c26fa58d51ed26223715329dd57acfcfac94154c2f693b9cfb769a68eec120cfc6491fe22ed47
zf394e0a590a69ff9c9108ea231257d42a0950461dad9e238f2537feb28fdb6b01a8658a03a8127
z3daa9317512ab1628202012608dd7c00ea014ad4d89cf11ec8cbc18196645c95bdbef6bc2d034b
z1b0b93e34d11295e97427509f1869aa9fd507ef49dda2e969247928af703559a3ccb013e8ebb1b
z3ad261e8dcb84f5eeac324395770aa3d6489141e0f9a48fefd5841c7e175504d50c72951532ec4
z4acbe0642cd822d33705bc00ac823b82f03b8e9a14f51958fadc3fcacdbacbdadb03b57e55894e
ze1ceda9511dad812249b145b48a903f2d2e6376f26e050152f9ca60c8ef151a9967db46c1399ac
zafea53baf7f13243edc9eda5035e7a9be5031543f0982848835a185e625a28d241a8607b95759a
z922a80dff560ff659570d7ca80c4d67183c5e2865dcf720218bcc809fdc4b362580f6b6f27ebb8
z4029503299602640dcb805be70d480be07c486035eaf2c6aad8ac9f65ec813608a62e7b3b782ca
z8ca9c0c1140da143cd4b5450b7ef2d9150727ecec2747ba1de75b5f905ac902c2b5f7fa4a173ff
zd2ea3ea8d58eb9efe858b7cff05f411229778291e0c97b0962edac00ba21c601d7b87ff9bfc1f2
zd2c867734e8ba43cec34222af1caaf9d9a82761739a3c2111d8bff222a2fa0ef585a83c3b25339
z1f212d3176848f83e46042f690c6817b51b8873de751754a7ff981100cbf89a717efa0f45c9f54
z9428e1476d8ae5f9f11da95867c17cfe2a0a37687054460c0d88d604924774361ccbf678279e1a
z994944739bed47fb0c372c7b06fca54204c7d423b801bb772c05a51d69f6c0117a916ffff4ff64
z7e58f97864d3d7afa3e9633a8a8ae1cc074d1dcba785f687add8b1e96a8a552af4c57962545d83
z3d679afd9989852d57534086d5a3ccc4e8ae22a554df31595c87180c1f8d23e32caf88a636a18d
zbdda4ecea2f6ec02ce81e294b13a321162d399507661743d1c48ee3e8dc717f5a39e5d919a98cc
zca2b7ec88ff6a9593a64b53fd0e1be1465f9809c01a6f7f54cf9b814cf11ebd6fae10504f01808
zd9946d300625cca48ed801ac079ab579e78f9493a6c11285fac64e4daaa58c1e16908ea124d847
zb5d670e7023fd94ef83aff36a7862047ae00d9242dfdb9fa461fad2e7b83f27f010da7b9a85564
zf021974ffcb30988b8351a0792270a3dd9fba07164fd0169488136f6dd49b2a177174b295cc7b0
z0fe220cd92fd07177bf6c4ebf32e0c952c687e8d3cba9e279828b8a9e2751c4634c6b4449fe231
zdd56cbe8c81dffef98ab00e61c7070003b8d7ca085256f25ea47ce29ff3744026f735de7eebce6
z39378a6a4480a2d88b365aedf8afbe30c9e7f2280b16b94a4dabdb6b1b79923dfa8926f82aa50a
z39f51b31f646dc6668386bb15c3f5c20ae398576b32354f3f332fbb9e6ab3f45a20536c10a6800
zbf6388065ad1f6acb7806ac428ce0ee79e2133d931975bfaee254856c88f6ae943370877b36796
z9002e89a0360831c0027b91507295af0d9d356f9475f957690eae6fb4159e733abacf2efc512a1
zb73d138524faa062cff9d9f20d9404a61c79714bdc092a7e2c9ea70b39da1afe7fa30a860a536c
zc84b438288f755b574899cec345b7476abba09dbfe6be5f4cc3420a09b7f205579eea6b0d53502
z856fa6d321ea660769deaf4334bd0301fbc43d3d945be140a8b53ede154600b50e559b5192b2bb
z2a0c2e3149507a500b3bb66e00223922bb3a2fbf8d6b2398e97ccdaaa91c7f59e37dcab84df0b9
z35c444d056c0bc04c4e1e7c21ab1cee13bbecf9a379fc47d368407bdb46bb7a74cf5febd75406e
zabfbb84ecfb627eeb9e71c55f975b3951cdebc2a13b36f793681090c49c4cfde58d103a790e211
z4bf6525d0f3425e64b6172217b9a9df76be9844ead25a7504a2cc855a3cea5e08b718eea6250d7
z1fa90ae24f4801ef3fc63fcd3b350151455e8bc42e34c0552eaa72db4400d70b77b11e9fe63bdb
z67089985d4a3cc245c11113de5eedf03e4e32506a22123180c9b6d762efabf5d16fccd7662f7d8
zeb8da730ac531a870d86d834d67dd39f65b5fc8daabe0198b59fc4f807009c644937d02a41f1cc
z758d7099d17aa13191c6adecbbcda42fa5c80b7c56252c55e84792741c413892fb835b5ab66b61
zf92d47985fe2ca5972ac69c004b8aa2c53703b673e10bf34b9d83b2702369de4c0f0c380679323
z553bb24b6da8611168a5088e64a2800ce037c9d5d7dae41520235e70853ccd41b85d8ac8c66c5a
zb974c0340e8ee0a87e8e263d711c835ee0214c45267ab41978f78ac2531358d7eba40574c35720
zd438474287c4889b7b36c88a08d39f935c237482dd971f6aa3f1efdba7cfa21c840d51b755e623
z4e2570571a5aa5a8b358b5951ad4eba5ce6300c5ecbd6089f37d09fcd2bd931fd45cafdff5379f
z7505e9b1d9786d40d5d2cfafd94affb5b9b7a04f5c6402741a74bace881e874f82cf64271af65e
z906c55b8ce64f3f74f0b6d281dd51155c71609e42bad26391c5954811164f288a4e1d4614c844d
z357be7bd451e6bd3a854692c3c61f4e7164e041bc923d8512d94f3cf1b7e9a765bd65cd245013a
z30f20e4266273532bd905dd075e840ee2e510efc71c7c7bcdc7d11c52ffc1ce96a213044ffe062
z7d353adc9c25926b38cb869e86254fe42557adfa03dc0295c763fe37741b0e4f67124f868c6424
z58640de87689c322ffcddbee741f5d2fe32d412b43dc2d5563848a7be48c55fc7c745220a94fe1
z3cfd2a47df4e76a43fc32b0a4c90dcc3e2144d386d90e6be9f101273a96554c7bcff4489bceca5
z21e4bef97366e1d6827d92799b39362bf8ac855bbb1aa71c49714d9de43f0c66f89fa5385b98ee
z16c71083784f6e9a06eed0078d9b9721755fc5af0291e653e698ac8815e2af22de6fb35f2595cf
zd602f3ddef7cc6498aeaddbba19f90ef93bb70ec5222244c6dc524f7b0fa99c97908e95f7b2dce
zb35eae2b96fad36902576215e2b9541ea8d231d2f1190b04afb7445c4d0067cf1eab41b453ea56
za36647539be3876ade7825e32d8b2d5a0fa1461bdb1818eed0c8614184b61f09f6d9e762b66688
z67c5ef0c900ef3351b9dcc655ee358150ad652e81e0ba9ff91d83cf4c1218e4558f16882ca0a26
z142ea3763c9872b58cb5ef51e805cd8daf072c9fde957d9c853613087ba9c4b31c00c36dcdc1fc
z6c8e7d7391cb4db037bdc65b7052afdef26e801c4f41cabc5142df2f49e462ffeea48d8864d7b8
z61904bc364a598a5bd8eafee9011f6cb4653df6a86462313af2bf7a6126f9f691e0fd2f45d20ec
z64b86bca380eb4e393950765df55d1e7fc9c3bfc780e9dfcb35e73cd1832664eff36ec58c039a9
z83b716fa6c6996671be3635c851ce5466e38f2de2df40f4be0563082f339a861d8645450e9949a
z131ae519bdcc917b72c2b10a2a207b87b8495cdf0d970372b14b3ee102bfc23b1e29f058a0e1ea
zc21a7804c4f992f29765ae8820ad2343434e0978fd773829179fe3e576a7c7293bde2c3b85f25b
ze5fda89e6710d99acbad3ffb12bc4cd2a2c2e45d8d985af40a343f19f1d16640da4d3a165d3735
z2d1877eaf9a6c091e0f8fdc8d367fd47cc2c288e0eb607965936d4e205b2da90bc65dd23497492
zb2b8dc0b281480a67c52ab85ce45744e60c866f40f79b27d3168ed139c91f23f3290b44fa4e9de
z43b5776b0994f71f275e9bd0582d8c97bad1db2789e727240646ec76931e1a62ab157b74f8a285
z189e9d4dd12a14e7b62d4cedb91cf683300e187dc432cca5f4383fb32b71fdec00fddc02e21093
z390de56136d2cb4dedaa4407d668d5f6cc8406e40c966bb1f7de74e3ce1b6cd85bc5bac6510040
z4eff7848f1d0998844bbe719398486ab250f7f284407f4df76861d612d11166f5c4b68750a4e73
zab3b6faa85e3ad769aeb64c30f788ca49c3263bd9fc5194759d9c7ec7b37cd9a6cf8a7b4cae5dc
ze2fc273574b32f60e4c7dd3d77d75f1a392cabcb2dd58da472b6668967c4dfd634819ec4c9572a
zdb24c8e72252f4b413ed1e81883ec4f3fa9c42e7d5e9b7dff7e07e99add24ff13dcc011b29c1e8
zc5c9fee4b53ca5d17dcbbf5237152a48c5bc6e4e5cd1add1dd269b9dfe7d6fae6d6453bf9f10de
zca5d8ea10ac0d50c16d23f44dcad4218d5e0ba19cd58481d7b43ef5e7128207b5fabdfea132669
z5784eae8e9d1273424c9b4a6dfb2413e8cd8e5167f240423328ca83e2aa7cff6e3a66e7bab2a37
zb4e8f3e9debd90bdb2e2cf898e81e9b0809ed267c4b740ffb99211b3ffa937252793294f84964b
z2490e8a1adfac9b9809ad1582ca91b72f17ea8ae42edd163b876f4b0ec0e8523a919bf8ce669d7
zcc493b8cbc559061519d10a4dc4d0f4504b8c4be4979ae3444ce8fde4fe43dc63ef60cce74e8b1
za484707ba954664ff9cd0abd7c78b817fa62c00e20729ddb6235931b4c4170ae1d20140a141012
z1dbf1dcc41dac3ba278375fc8e3d41ad64f9ce5caca45542a45e64b1ae3990dad800aae2575413
zb648d272b39e80615d1a696460e8bf3a15e63180643d3118b8445695707c9ca34fe2c20fd0ff48
z13c597bdfa69c7c5e352f8636b381bb119bab3fe251cbc54d2d6d6f81c4cf21eac7c4943c225f6
za71d710bbefee6725b948fd11ad907ebfb119a6911904448e6a2a7f69644bb84748ff9f748649b
z87b7e111df72cd06576f07a875fba1255c0d0557a280e43433a427e73165b62569bf9fc99ac17a
zb953cc4dc0769a9fa4a71c463211cd264d93deb9b3f0bc32a45b7c8291708bc2ec90285c95c844
z47060f5a9bae709c830e8816075bec1a631ccdeff6c982f1d5a7d037e6496a9ab3d527f06a2aae
zba935f892282337ff6eba4281738f096ed7529fe6841318376f0232fb92fa66efe28b4567ee9b0
zd886c2d8b1317fcf073d29087f3eed28b1e5b5990ffb0954b6528612da26924a162d016c5547ce
z454e194ce70367e616e03fb0a35501bd1c213a718bd932b508052690bb92edf1cab8cbcb5ddc42
z17587cefa8b983d54c9a9d8b007d9780cbdde8a0d04fe4093630da16d43b69faa2c328c6cb50a3
z21ba6b1be80a035237a2199dde643ad70117e0e264976e97a025927befd1b93186c9df73f7ec21
zb0aa1b77f3bc857917af30f1b6a5d2090666e58404b4d0fd0503c6bbacddb913528bb93293cf77
zdf57911a6ad6223a4af134027ac453b006082016e407d71646f0d470a3a002447d94d388c24e84
zd848e06e452798cf206050897cb1146de86105f0e97cb84b44289ad212b4b8991b699500e86856
z0936fcd919899480bae46b34ea6621b37e1df2b07c4e3a8c3f7f069c0d3f3481f616c2c38083ee
zcd39eeb81f6b9d6d3dae26cd42f22f9a424362581ebbae86a31a5e99ad7135cf634f93bea95924
z78bcae26aea808a4d570f588eaff6412c4309490b098cf807796dcbc8e6d5a16fe5544e5aba7ff
zef0a8b9b2927c03bd2bd170d4ae140e46c4def6793fcafa0ce1cf6e35908f60ae6be82733363ab
z2841cb5c93a72bcd3210ae715d5c032b32972860b208979ad2a36a2ecacf147f82b9d2b93e7c40
z34cf5592a4d8554603c910148acd4940c396406d9d59d21d8fab61b0f0197be60e19d8bb0a5fd4
z8311297101e0b46ac5305d46da11f69f3e40ca27995110b5adec5616a8c17f029e1dbb561b0ed0
z6faf92dcddd73f8e55e8c6fc5f57d470146e9ca6e776f5627a1c4626c5252983e1de89b67c00fd
zab06cca28a6def7e4655ad5042702ebf8a90a3f0ea8f827e5512cb62db01a717614551fc81fe0e
zb465ac6fe2a5af1d52651e38f106b15dde72939bf75c6e68d2a6f6c810889d42b469f0897bdbac
ze93ee87d1cd63e9e885be2a0a8b435f08f4479bd4ea9007e6e76e22d48aa8c894ee4707cae2421
z06c2b87f21ae7378a1814e29e55e56bc33ecf41889c7e895615014bc1cce6b3a62121ddae2a855
z7843c5d4728a0d772cb323a32162384629893aa90ca9738dd2d4d91b72b86ea31a3f340232b4e8
z2c5f28462f52f39537fb5e560f59bad184346dee81e440abb1597cfa0eb518358e88a49032557d
z5ca19007e45c8fd8685f9e96e8a22ad6dc08aa12538abe2a719672addd488c41027a5757ca6e35
ze9b490af75ec2b066a52ec5229fc08b22396be9409e2919d84f57b69eade662d6763dfbd225002
z3b838a97a9b2ace5b596a4b1ecbc47336823354ae7161376356d43f01c8b939217c7b204767ba1
z3dfa4b12830ceed62e9b1acb87db8add4594f469f9b50ed7e1c7c47ac00e77463ae19caa3f26d5
zef480300c6ebf7b464e5d70a2e9557a440c3d5b8d9c4b464e8f07f651fbff8994dfb60c4fad031
z28d879994372f5c672c05cdf072661a6bc6aa4d5c83d2260bdf8d8390dca8fba1d048c28db9458
z805721bf2e5b1d43dc2a3f5ad3548d1f339eb060d29415660922055b139a462a1bf0dedaabc5c2
z9b46f5a5c5c04a7436c991032bda73f293448b52da24c17a0a27aac8dc5a86cbf2ce2b74e6962a
zdb4c46e77a004125e10a08280a25fa497a88b404bd40e3861c4ee20869754999e168113da91f73
zb6a3934530c6f6f93370848a3fa131480c9d32fe2680fe2f53a5f6c7698fa2c65e794b6996bacd
za708b8cb414acd3a0d821cc945f677fc3a658f08d0381d8e370f21ac116e9d89537247328d9f60
zc06ab2ef609bada97a090e0da066a7506d903582bbe114bdcb81ba6078bf328067727d40452a8d
zfd882c3e4623377e15f3034fee49df2cec55a172ae1ae474590933ec437fe9bf2e7b71e221d67f
zef8a2ca791f05d31ca73e091aca2a120c0c5848b79db99aae069372ee43ae9cb00861324fe8288
z94e6736ab8b5db0e1cbf70a0558793c073ed73d61776cbdcb3f9074d16d1595dfa5e798b89f70b
zf6be661fa327465a2b41695f437201e41eb1628bba1a38801de9edc5389c6387b1a3b844e67600
z653fa50e47b0b9b6e87e6dfe3112e8db981c0226de30d3ab41ebd8ca3c74d70d71fe02d1425740
zebf9ad87538b45ea0019f36fafdc7d4314e8037e9b7ecefdb4b4f8809dbf0c1cee71d514b60da0
zdddcbcaf3ca44ef8a3e3e2899441bec822e254304af47009814c3bf94699fbea10350d3f78dcc3
z9b46adda852319c18a776d27864deb11b95ed8e002a43f3ff74ead8903ecaa35ff896d91822df3
z4c89924214658ad10828d173ac94f766668362a56b2ba1b4a3ae88908315656056bfd831be30da
zd4826bdc8942348a3869c731c002ec70b1f6e9611d918dedbbe78d8095d61acb8c90195f2bf616
z2b0ebc2d88ff71e94cb39e82fbb39cf2f51f89b9fedda34769e587d35cc84e108cf473d6cb2028
za38a20bb3b9e59e8e5a8a1bb46fe2dd7b87343bac59d5a8f2efeb9330cb38f96f89d21763a995d
z88cda91ed03e67740f7611be2d89d1fe05e1bbc044f4f23caafcdd0b25ca748d7561aba715bda1
z2ec650017cc6172caccaa7c6f1edbd3ac16bce8d64e292d7bec344f4f3c39e23931dc90209024f
z6d1866f9aeb6b78ed99e5f495228475699e85090c75bb87bd2cb8c15a4c66d6ef784894dd14306
zb06e409059bbbe1ef25979b65b5bd188083a4f9d87d28ad155edb695ee00dbf1e869dcbcc7ae8f
z96d9f27cfcdfd45a72637f1e5c416726603bb6218f1230601193d6bbb1cd4d510ac772fca8d807
z9ee5b8e96914be54bed62bb5c23ed24a12139f884b3373eeb80aabfdea33731b9663a230c3a111
z2a8c8a58bb7eac62f15dc9a0b7a8693701667f3445d23f5c8191631c53605bb0b5f2f7f74062a9
zdbfad5835f27e63d234a054e26f693a50a4522433d88c8d9848de3fedcebfc1802e0dda2fd05df
zd9b720faaa1d157138a235ad0309fd7715c80821b13f533b4ce48b585cf0b9c9e943653747d6c5
z2ba47de3153a7a59ca722586c1c7310fca781cf26761a82ed9edf85bb41abd958dd0289b976ac8
z415569840cbc73d6901abe48d828d9824fe81f902f9027221ce32277f9c260bbec2883181c84d9
zd9d66da9bc93c0dd31d4c6a4179910bf3b9810fae20b528a057472ed3ed6c12b9db4fd81ec64a8
zce30367493d32becbd2338065e93f663288503b6e19b384c7e5f3f7998dda818e7ea3013e906ad
z147f2a8dbf28125131de02d6b0134c0b2eca8e7617736d3c53163bacb38ae4e2a732dc3f2c2e77
zaaec94364590335db9167273ad86fdf07d4d80c8aeeab203cca4cad8c6b55fad6197d320f1bea4
zfdaf372287d627462aa89cc703c33e0e10146ca11906b26b9e7559669134f9056d6933a15ed06f
z59924f1fb0186e614ecac5ab5ff4211c68acbe358945f339731d4f25e36e75b8162cbee54d4415
z8ae0123f3b01825babc5519beed3495738c31b947c394d0369e184212b17947d5010e72a2ba6b8
zc26adeed1b808900e6cadf494239f2460db56ddf8e91ad47e4d899066715ac5d33a268f07c741b
z07b5358fb705fdc848bad2b5b9539482dec79deb898c5e83092b188281af7936b2903976e09f56
z889f7eae76801967ddd4ebc1fa162659e96caff0574777a997e337a95832fed192a14a3a6b53cb
zab13e4c81b77fbff73bf500aa16be57593ad4ca4de789ca76679ba2d28a609f7468dcf6f38f8fc
zf2caf411d14902535723e14c0a63d50b6449eaa905a8437b1576f5ea11ce23600613c7bc890c6f
z2af318357c312f310d133dcff61b5ea26821a1dbec69416db85cc1a21a63832c6e8b6e376ccc43
z1b225af0e6445f0413716fc7251f75589663ab98cf1decf757009126c32999afc418b15a53c0f0
zde2c0cc54e0631cf74fe80728f52feefd7a84765e0a6e9ca9586160c76ab05274a7148655ea380
z35997a7849c3c882d463f5573711ce6cbf7cad7f75267099cd132f2244e7a59a1f2b73f4c5e3c9
z1e956f2a9e424258a544a505f252f50c51448bccda718c6474d68480c2b3c756947bb11e5299cb
z961c38b6e2ed35992d138fa80298ad7f5b87a06a9ce31c84e75022586769155fefffb22b16bdab
zbebe9e13d7d8c88958d5401b5d231dd2ae4acf327d3d6d6cc98da90c0f25c43709931dfae7c8fd
z417ac72dd04dd40b29a68ee905631a94ac9de93c588bd8151cf4cf49ad790e67fab4b52d422cae
z3ed0878931e4fb52b29d1234c1714d233f0e465f3105c426c97e31a47436861ddb8258b34160b2
z4489161622263890521408c4da1b2f0f998737b43a18d336e7f71ed128d4617d202b71e76b3000
z55ec88e418e1c3797b378c8b262f05ccb0e1d5c7d3fd47c202a5520e3cbee57ed5f3dbec712f02
ze29a08ad87fc6b98581a4a0de6f2afde3c626d71ab7b0fdf7bf6935ea159070328c0697a1ff572
zf798f693e92009e267e0e8e8cea053d1d7248e00653d06ec7d46c8d6b798eb35819f3489738666
z61422a271222721a868599eb3941ddcfd25a557c8888f2ef1b13ad531475f6cb113978bba2574f
z18f4daa54097111ead19026f4f9219f36371c9c2e5f9c8682f3ca997b78e65d84d9d021ab426dc
zf516f415098d8703d15257d6cf5e4ebececbc9d2fd11dedd49264a091cfa6a5caaf9f6d912ac4d
z2b8981e8b59b85d334513b002822d6482c4d3a64872d9bd90141f4e6887ecaad4b8f9bd662bd6e
z00a6770944541a94bd61c5a9d1f1a4e79d9d843c32cf88e5da04966d6e251fd10595eb517d86b7
z158180e3196946e0333cb300b1f80935842e76873a6b3c24220afd6c502c4fdb8ca07f30c87955
ze3888f9750458b28bdb9ba33ed905982826b1fccdd33bc45ebe26c4b4dee84773181748257a7af
zc4b7ec8b1681c163cc6ea1a7fa5320692f3fbabacf1402ffeb277a309ef2f610df61cb780417a3
z4ff7ed506701fc7b02bf17fe62db4a5188ccb2fe303e1561d400d59c3b5b031f07942b8f932a8f
zc68b24ae258f5d2507f8acc54a2fe3523e1ee46a97ee770d935ef4ec7ff9ede8685bdeee946632
z911caaa9cc0c193522bb67d69d44f7ac50810a1520c015a4ba84dccce9ca180944056a2b2c7c43
z29dacb5a7664416692cefeab2a2a74761954807c827a539aac04e9046168f6c437ff957b486c8c
zc0ae6d36fd7633927f5787260eae27d3bf3f0487830a24d5a8a365b2c57fe8764e37df5a0fc5cb
z8ccee2d2eef3f2ab9a7362b720d807e5a2579b7f2277d93379e15cc57976ae78ab98260e4276a4
zf5d3ce155844b3f61fa6d3930c33c99f653571b6092316d72bfcbd3e3a09f4eec7e4a31546cabd
zb118e51e0db997668ec69c5a11ac989f4a60bce5aa344b2ae1205a679334a5e09dc384c167995f
zefcf8ead5e89545466eb68ad783e16f85494d9ecb2a610aba2ce1feee947fc71b9b320bda2d46d
z1dddd7276f4ff51dfdecf57dfd33916cfceeac00be9ced7be35cd1460b54fe25063b161fd2a171
z19e52285e25bc5676afe73c3742a0183b7138ae7e9b3f86ef1149d5e01ccdebd267c9eeb3742fd
z5352c3126cdbd2a5444a7e51779beed07a27085eca3245c4a4d7c0ad2ab6f21aa8d77abe2c3152
z27a4c67cfcfd058f80234a44b83f8cd56221d0f7c5c359cd851a2dd0106f8c3dee1790e85e4775
z536082ae651a6225a1ab7bab95b16c0467300349cfb68030a8677006a10e06de8d78580878486b
zb8c181d5a400ece6ea3b1f83d4cd4103d0626a771ab046de5c85a113bb53831dac2bfe690d17d0
z707a29ce4863adf04ed46bea21e3cc159bc9292687c8744597998a0601f3904733cd1c52d3685a
z0710bb6b92c1c993ef0fd8fdec54f7660d43799285f8c824d499d8be6fdcbcfde85c96a8247258
zc022919a07588641d7b22c2ace5fa6331a12601fd96e913fad2690af7cd2065b6a8a347ad48159
zc515bf050fc1f37fb7997281ca0d67a157a9186342dd5c6104ce2cecea7289f4227bd6c126ce79
z08d66832637672bfba3deaf8c44ed71322d51308048b219f48f787dd7843b97dfdb1f03e8194b3
z8d2d59df3e578c2fca0377727565baea0e6f488d19e302e0d2a499bc0506ded0ba101e12da269f
zabf054d7ff1b0e9fb7ad9efe061a7b23990a957d16240611c86777c8d3bdd4927b92efd15d7837
z96264ef9c1af73dccf313ecc6cadab6547c17e1c1b5d8f177ccf33501ad69d8018679e5a9f2ab8
z347b8d1b7fae5f0e80aa0e93629a2deb1b8fdb094802b35c934ddfca76f5576504c80e2ca4cfac
zf0234acb49469ac75f779933d41b5fe6f10e1f1e67f3d1a2c7f202db39a7bb7dcdb873ce3282c5
z05caf7581226ef938c1b81bd57b799eb3717b44aa7c65b5a094467328e17a49582894f8911ca2b
z4bbe2007dda027d506bf55f56d2bffdeb3e29b01f3d1f5c8a67cd10d9a89a52f238355b4728549
z292715fc25dc4ed0713e72b0422569ee9f8fd24e2a3e06638da30e299755d43680c38b9430fa7c
z2230f02d8a19a981c775e01558ec5a53325d820babb84b9bf8e05da1789a632021eaad697bf0e5
zfd692775c832ed1eb4b02a394fc14384f9caa49ec826ed4074cbde6dae1bb2b32f6354ec53a76d
z3adde1c26405bc9508ff8dbb85864050042ebf6d3cda772786d60ba77038466c373028a6746264
zf42e64c961758f3c09a065989aa816f073a457221121956f804ef1b37eedcfa1c35f22f91b1499
z5ac0eee150ef9298b775d1d6e10c53330d1d4fbc8ad04ef3ba6f89a180eafb541f20f7b08e14d8
zab77320657c7358d2fa58f795e07e8f65dd7ff5eb194131d273bfd4ba6878e8f380ba957e85e35
z6fe86007b43634373620a6805c1255e837d231238e057f891536dd8af5c3b3f19823d8b3e6e990
z5d50ef3a93623481214b63844d0c18e6ae413fb9c101767dc5e6d8c1195d708e19a99a9c820af8
z4532b5850d7fb0745ce3ae4f495ac4de7d0c468f73196f2b2237f2a51234d3381574abb88228fc
z73f686de6e97d8b92ed39b79dc0576550dd4e8b55d78819ee7238f44715cbef2e7ee7bd1f801ba
z985672a9b03829ff3015511f106be5db9ea5b23550fb1b72961e66b2779c56fa7f2c0aff0877c8
zfcba2fa49c2eea4673f620d3e1ed7a4c271f5cd3dbb4de8744e8cf56109162c1ac2898c1cac66b
z6bd73d1d30da1ae406a51303be5f6a8b027ad3bc32b68daa239a16a557f6ac7ed45e4699b818ab
z8eeda51ad3f10b7a1806662a7e5325ef9f8d0d105ccb475b77bfc976c6b6421a0b1eb47f45cb79
z99b2aa258d03a1b3a4e2344d98d9b8aaabfb5eafdc06e9112cb52d5f10351e191b2e71efa003f0
z4ff5b528dda02c2904f44d1555e40a42b58d96dea2594c35781a49d7e3b5e8ee6aa1e3bb4be87a
z798556896a4740d8de897b183c438e32902e8964d6d9a2eb8ec3bb7650719fe6de101ffa3b7b52
zf13997f0abeda54b1f13556fbdc8233987509d30dd2b69463e38cbb1aea47153c3b5bd329990f6
z0dd068806ab99bc43aeaad1d2317bea86f665c1de20429e1850e3578b2facaaf5990fea9de8d33
z7688bccbcf7ee241ecf9e6ac2f47c97c71a077c6e7193faf9680771c4506ad12fa86233f15f53a
zd72185d3e5336034c90e4a42653bf77c016a17c5c51c018e19bf0a97b73f8b6c0620f4a9a3ea44
z6e1bc688c95eb93aca548f02c3793dbe00f3cf7ca3477f12fe637134035bcaf1b37c8f0347d160
z7a5a1565574748f4e79cb41e6be3ea3d549ef94452d9917c2e1c5b141e5b033f53fdfe5b430426
z10b176cb43355b9d7f89e0b181cb22156beedea87c876daf3328b44af6374ef452be46ec92e16a
z6ed34e332602924e49cf1ecf5b24ab09cabe00c9862008c6a9494a65cb3c079c48cd48f51b16ed
z9a171532a5d88dd82da593467b5dc68c07404cc48ce2f6bb17c138c61742d8e64408b3ad3c9d55
zcbd66a6a2ea896c1ca76f1702a5e620454db3aa735d68e11fdfa680c9b68a791fc4ae2328a30e9
z88b44a3c4302da67a87f46973b59f134f98f0c9a3411433859223d6b3f931874a6ef26050dff78
zbfeadaa02514a1bbc428ab2778d1e1df752953dae448b7c2d5b173ccac08bf9e81c83420d1cd0d
z38de9326d3d5efe6d4df7d9fcf856f993fc16ca42fbf4fb2cc16091db8359a06ea6beee3776a17
z241a3d11a43b8a1da0af1ae3bfb1ee4c30e3f726bdc321b34ea158c209adf58d54fbc62f5baf87
z99026e85fcc14e9122759c66fd162adc76de52a715b9a9f2ee68c446a4e88e35d37bcd6ffbd0e8
z05c82f9b401417c60c70236dd4a832c6e5c71fd1e8ac8968f4ae5dd32fabed98641b7f76c17c27
zd46d6915f9ae169844bd18f0143a9dca65762d163d022c15619a872928b64c5016d89875c2b247
z4607201b4a7a2105171c8e87d0778fc368f10757fddcd58e15fab01160b35c1c2f26b7cd3e373c
zf9f4425867076eccd01882ad525bd8c35c6bf394c3d8768f408ebef13a7c26541bf2a839c3a13e
zf5d5a3a8eed1782d28d236fb0382fb48177dfda5bf5be5a598023fdd2c4c23dce536d6d2052e80
zc82ffd5d961771d0df25f17c29dba1ec2dccdae127cba69e773d54a727e815b95d47f325d10322
z75212637f0516a8ee429b182ed73ff452a55438be1be076042f473be48181c0fb79ad1519dd41b
za506b4723bc4a63d20a59ea9fa1c6696428d0fc6399962896a38335865832acb2c59f3313ef9f1
ze08eb51fbf53ac37e281176a88826174f1dd990a819d6cd99cb7edcad3cb8cb3ef51e1a8f8761b
z5d6e12be260b0dabe1c43643e332fa43aee609875feb19d9176606b7694be654f3ca8d0508e9a5
z3030ae268d503d40f6a457f19690921615eca4688ce4a9771a3b300750649a5aafa6a9966c4684
z393c924399706a01e6e61d79ac3a5aa5933ca74ff40f6025f2f910795110a5a102b1d72d747a8a
ze1dd33431fa38aa172ac31939041f733386184fdddb7dcc260e903ce1443ea6daf8f8016f98573
z87f47ee40ca4454d6967a9aff5bd992df04ff4e780b325bfaf152326ec0ff6347c911a5b9248ad
z084ba73ff393f1245fac8206725d304c362e68681e20e7017ae7e1d63d13fc2c53c72f30bf8e62
z9aad48dd54b631f7f1b58725d27775686a195047616358b29168f6be6a15298015fa4b71436c33
zefc7f247748ac1b18b57b8d6ed68de881fe17227ca80e00732edfd4bb3bf62cf619a058440251b
z8db2a73da2b30085f46cf6cd1a37b5e6310dda494aa04ce886476d57f9c5d3bc943abbed53674c
zb056c912c07a1b7568cebc4b23ffff8f91b78dc3cc3a3b15643bdf593d5d45ef65549d72e1f1b6
z9f136b1656238d43ffe5436254128faf4766f47f32bf2b993e0f1865bdf8c14477c04b6d50fd8d
zb741b98709314ff67d05f9d0370b1e5ab849602aaac0b77f1ef8d1ebbb4523ef734516f933d1df
z2344447fee7db40d1fa22c861ba7d1e34b96816e4923f37b2599e034e761edd60ed9818feba3e4
zda9dccb77bbb8402837bebed476729c516ef0032b50ce68e5b065b64a69d2f5874cf4722745977
z2925b8f2700df9e6cd6ddb291ee8472f4deb7763d432d0b036783a860ffd7fec90e68c6669232d
z224a5e16e230bca2af337b300e21d64cb6cc829c5847a968ae872767ab5ab10b5f5d5a7833c7de
z9d280c4691aec9aa297be9ea736ab48af7a416be6a186e47bb18d07f96e8b43bffc4fe54e86ab2
z812b63140035853991daee74aa686843e921a5073f9a698a02ce6f83bfafb7918161bdc147552a
zb05d2381c49a3be05423d27c1d42b3d602e1388b7dd99b221cf3eec8d4871a8c486aabf4f86635
zd02576be2441b6a0c863ca5c522a6b42c0913c38e4e8f463f06f988f3de2e60e5794f55d4c9a42
z2c82c3b2a4c5f65e2087591c90f523ae827e0c04d8276fbe4bb327ab916ec53a873e9de8eb47c2
za965a5f7178d166db11d46026811afa3298eb91182985ed8015c69dcb9666c8a2864975e7d5273
z6f41d542c9c4d72abedfd0f2512616a6ced282ce7fc0d6a470bb7f1ee5b5e8a40bc12eed04a2ba
z3be50e7172c6b4024fc35372693b54ba2b815fd9697b92b113e57ddab8bfb139b58ae046e50755
zbf6f3b100aa5fa9b78ab3dab85cbf3cac5bf18adca6d366da48d0d802bb61fd4a14d60d56b6bd2
z0aabc53d84973b283f3010779ae440440c3bef259f16eb7f453bd79dd2b335ea9257ce3b9054ef
zefd8427d08621e73c0b86ab9a94d044727c2432f00a7d5555c668adb7d15e1af434b0fa5858937
z05f5cd3bb3c6d4a1751426ca92b9da0e70d039cea3969c28a3bf7f11ebfcdf78bf9ac3fafaf9da
z6d3d8fcd8797703f13f60b09cf2bb09ffd553e6f7b6620cf3d38cc633be0e6505b99364c8d29f9
zf191c64a5ac6080391fb0e7d6841d8322f53a869af9e91dc765b7b65a84e64c5b78d183c2b5c80
zdf07c3006a7bddbd29c2bc634e688d0265124a54236bc8a89a37bd2dbb6379f7c5f750d422cb5a
z889c2291f728375e87e83067f620444c0e7ef94c6310838eec0c0318ea2e9a20e67f17f0a8040b
z3739c62c28e837d8f1ee3ee9dd899d6d3cd71ee3462e17fc2ec341dac29c79673690335c0d1092
z1b4909e4b33d9012e10fc8818145bf904607e1c6de6860145d2e1dff61ea22bc665fd7a8635552
z22b52837743c30584171c99b276456e8498219ccacf3c99b8feaf68f53f02c5d8539b19298440a
z36a4873c15d830dfff64a4296f4000c787eadc5fb49ba00764f67b53da1e9e857d67d0a2f45040
z32cb7dbfc5e517165b192a991b743c4fff9321e2084c39482dc514afc9eb9c13a6c621a56ecc9c
zcfa3da83640895d35513ec2d8d04b546824b034a3f1b4a9943245f8fb796bd6c148d3cea1048f4
z69fdfac23d436c8e2fd0ad4af08edd9e073f41a43f62c85c8e6217af01baac1cf785e7d187243d
z1db890b66238c53dfb2574679931d695c6a18e34cb00fe1ce7e5508857113f88ac65da73ad5e9d
z110bf5d323c161a2d3ecb6b975e7d698e20e705396bae8dfa4312fe31fc11d240ea4762342ab16
z2f8088e5c8859e50ffaffbcb2cc5b6c5448ea4d0f68ae36571d3793f34c25c2d1697be82651c50
z3d4bb3a65767ad2853d6b925192e0230586c441331a4a3b32256b2b9a329d09e9e5ed785e5e378
z228baede2dae1de76780fe34394c8882ab4e472b823634a3b88f292efc5339bef93c7bfe539f07
z677e7cb42dff91f8bf73fcac5ed2c16e4dd765be3aa01db227b1fa71d4e0c67495a8849f2c619a
z4a64f57abc38a34f34177624025c4fbef4d12022246e5ed97302738c0da08bb5acf511f0d9f87e
z6b04916e7573df1b704ab7388c41e1fcf7065717a5c84826963e67dd7db92f0183f63a8b9eed53
z6a745e7240bb1c9328154557e2f6d5e4793533a009a6b563a739c3dce95cd7c6132b7d820ead25
za17c756e8de33208fbcaa211f8528e3441265f9b389c148808c322211b21bd8a9a7fb1c57c21e1
zf80b1857714d29f0e8bedb86ee2c82c54ccfd73a7731344017876841fdeee8059e871713e601e8
z441434d8c1acb92bde0933c3f6515d07761045a8b6dc58632d82346f560edb05898639c71fd1ef
z51b0aaadb999a1628d292684f6cbf7740869a0faa6968eb120c86c30871f8cd00d04630c87ed93
zcbeda8d16e5e04d9b2e9b3a1530b49fba092148abb19d6add11864c02827e225a3bf7d4bff4ba2
z9a821f3b90bd9235befe0652bdfea93c154827052f26c559321e23d5b91733e5e966862ea75a41
ze20305303fd83e1579d40e76c7caa6790bbdf1a4eb74fd679c3ab2e655c0fde3983e98f9d08a09
zb564d5e5b73b8e531d29da344224d933ac42fed58a5a98c851722b2525be33351554ca3192f18a
z306bf1c1cdb6bf473a2785c0e6d24625602b49a12b1e9e91b15ecf823469125f9b41257b49d739
zf2f5ecb7e109cbefb9178c0cf52f067f77a725d7585cc65f334deadfaa7fd57c0a545e9be836a3
zb45dff3a4a6a2ffc568b3961b6b5feab281774c75d858a18060a9eab035d0086702686b21b5004
z0afba99e7d5ea516ee5102af61d983495d2a7cd80b0599dfa6d0a773baf468bcdcee5519e00376
ze64732518ed4fcaa3ab0354f352678f308497d742a19ed7d332a05f7c68b4761d70716e3ebcb18
z3d3d927ee4c514327d42c668a0b6479835600b3b37124ccdeae60eb8090b956e80dd89dabce151
zbb4627784f25977a64f6f098db61eae53f4c7e1017eb8d1453d214b00ccdf89d48089ea121fe00
z11433ccb965831006f70b6d4b68b016a5bb2e79d304fbdd91cc0a9be373f2093f168e20f3eeb37
zb7edb2df0df5ac18046976cddbcf91effbdefb93d31a8f4d2185371fd2d2bca3d861f4cd5a0bd4
z3cc1fd2965ac620b5d4f67110edf3b62b7e2b56f7b08d7d38e67639967c6761fb82eacb04d2fcb
za557fcc2a8eea7ffb97b59eb951cb7bdeb842a5495678e977f8b2fd81eec72b86f39b0a03cb054
z154afae65990575b468c654251b42d1065d0741398c665f293b04b12ff80d16dfaa5be0e62922c
z53d70b6160bff7d6e3cdfa574d329f7f6b2dae9d020877a2a31828f4f19c56779b39ea63042845
zee8b9972c51eb97d451755e37f7a229e8a99ddbdcf488c8891fd52cbc87b0162518a82f9912632
z6953bb72eab09dfe148cddb3f4f5f68993499a33e61cfdf763d4468430e5b3375c50874c9f21cb
zc569bb74cb63bb39b96f110cebb22865c80083c1810f1a002e0e3c1bab83e9d4b50d8da57ba3a5
z50dad3b4999849edfa9a7a4cdd47d5d1ad7ed7d995d29e8483e2e31b5a4795236e03c0de38bc00
z9f87ba092d7f873d0cff88441d5e7170c99c897bd59e8b090c3d1cde4d8efadf9abad4f707c5ce
zcfb3ded4aa6a2bc191f9ec9a5910ce913700d11d92c2a4a70b6970b889fb77a00c90be49c4dc5b
ze89e84585928150a410a9f8e2994d0d799d2e2ba5255954a62b48e539c102ab0a15ff5d7b2c838
z32132921e969d36829ff49334194c6a9f7a1dac5cf05ea0759a26bc3334b9aa451cca3f7fac51e
ze505408abde40874d2976c19b7ddcd7ed6f72020069ad2d6a5e2b150e5b012996b0236ff8b7ea4
z3ab1625928866fbd86b8509f5ecbe61ee81cc853311438221c7b0d32a9a8f42008cce9e982dc09
zb8fc9ea88e748af4bea001371fea9c353d765cd746ab0b2108b6011b25a61fbb323224ebfb5be3
z459c6df38cc8bd9c7c79199626b921fbe04091c1e0d002e1c70a0b3dbb426569fda5752811e696
zf53385ff42c6ee20d5496ebb89be605aac1062b4853e54701be859aa46bee59664d7c694933c2a
zc3b18415091a67f55e8442cdcd368160b6409b8630f5fad92119329ed45276e2e0db73ee1de355
z608c5a5b162ddd7ce77051ecd84ca44c3ed2d807d1ca848a350694e6234dc85524a1cc36866d32
z1b397077044a5a862fc5335d53cf6f6ab813c3bba811e7bcaae412cc06a5a4b467449d8452baad
zaf40cb2173020826b16800bbde463068a2bfa91b8ccde4bc6cda11741fbd6f66d9a95ffe396176
zc1a0b30a07d0d9a17f5bcea9dbdce1dcaa24aa09e38de8946b68071cd60856f7b0ce135d26e8a2
z73b4998f1228bce35522c24b4062972efbb2fb4860707f2a796d8d08479a72e01ed5224c431cc5
z61e49c9f9d230827b6ec8b37f285233777ae58f1d22617d55090ecbad4a60b36535ee7dd7064ed
z38fd37c72271ab677e99ed784e33c3a5d3b615b195c4bbb2a6a8be93ddc0145d254c0505160ef6
z7decba86279c77f913bed9173e4b89bd58dd0a62e73e96bfa78998460d20351ffc567cd183104f
zd3483bbca7498a38e1bd693e985de27de115e656c2b58729c0a38f4b093995cc0de91cf6bc5c28
z2674653366f7789e02e5b3353f23d2dcbe85df8927272dcd222381bf9b78d6eed914c746e50a9d
z1075597212224719ce7d07652070cc6b6629d75e826a7a5a1a0a44c1925498457864dd85694ca5
z473e4bd15aa47aae75e1809b8491fcdb93c707cc13d9b450014ea55d724ee718f65f527b04aaa6
z756be72472fcd87e94d88badcd8f8992df50cc87e66b51e46c3c57d83e1a71192eb3990c7610c5
z8de8fa351643d3be21ad97f9d52099eebf49664fcc5319bf1a240a441c5e170f248c05f5b32cc5
ze97641b9b0dea873ffdb75e79aea2775a41ac0265479d9a9cb1fc12d7a34a1697630135a9fc193
za5ea00297fa623a98e93d4b67c6b84a0503cba4ea14bf9d1205051b76a3bf1576de2f4d3b1b692
z20316dd697f4630bb27ff515d916bd4a2129b3de9738cef30baa12912a2546e0379f15b7b87272
z0a29c2910688de6e347c58d59263d62229ea22da2a5f2d6e57a51229b5ca3a15006f1912bf8488
z7bc3024ec2f4e22688d08cdf9932f9114ca1613d6a951e49d0a18d63bc8f00d78bcb88c8bbecdc
z2361f19e6efd93ac6a208ab326f048739ad5d848c6fa11485b8ce3d6a8c8425ef80342b5c59ffb
ze4eb6428acaa8c6daaed6c16f88f9adc8ae85e9e82d4f1607c24293e2ddae88aa10106f77c4e98
z50b11a7d119758692c644a00b3fdb39b1ba5721c98eedf8707f67f3c72d4e3167a7c86ffb1a1da
z4463ead83e4e49b15a25e7744e6994344cb493d6cd29997bac6f5f8d50bd3c1d088833811fa887
z8ce37c247f4afd83ea3d59b4df7b680658b367929b250b89aa72bc11223185c0adc0e7b5373dae
z920b1afbbbee2689b0210a5016bb9d24dd093738e0f8172b35213dd13f0b8bbacb0b3e971f2e3d
ze274c5b9f03254f078d5e98d0ae26cfa4fa49dd642590d6904936c0f4a29901513d657af645852
za43af507103c787278c3d87abfc4e40bf0a9e10123ad088c54ec2ce2aac4470577fc4d8d436119
zb0258e02c61c77273e7391a08ef2bfdf02431e2f4a97438ee8e722b65942f0c7cd6671d4f8459b
zcb53041a683dacd77ced30a3974e0683609c1ba6503981331a6c349462b8242cc822a2f048d748
z322cb16d58efa9b8c071bf7bbddef7390c0673cf9a0bbf60bc7668cb926c090998df087b062be8
z79bff6b80d4a845ea7f7e654db768f9a0b5d33020289f3cbd5e53ada9287becf38e8797da43dc3
zcde7a02a78cc464dca6cfdd48661d25ddcf4c57f160095b8a281888b6bc7ff7f33fde075a9ffb4
z20bc119ffc840f7f2789ab4de74b7f1461f48616473af8b561ae0a5b8857786f2d4ab8562558b3
z7cb6f4bd5db28da6eb1370b86b86b14c3202a8f50712ed9364e03e6331f38ec1d5e0fa84c47b5a
z87daca0058d4cd38aad79d6218c12ca08c08b661408578a2e4117fb1584d51b9f18b8aed725466
zc7ccefdefee8ef9baaa5b908eab600d362dd6715601064857da2aeb61743a8982ad51c491813e5
z6f62244af21ead52320124cfcdbc8404d0318223fcef05d9b50b9bc79b4701079edf7902f96d24
z6e5547754c2383c946c014cf5862e771b6a5b19f5f700d0d0908f286663c7212af28dc209f8336
z87945ff9dcf0a1e5074d8dd0de7e6c27ddb2e8fcdca61b9b870ef39ad0eecb46067ea5d0f02dad
zfad1c524a3f902cf8c375624ba8554e3215265b2205e6c3352cbaac137ae872b050e375ca75b34
z599965ffa51a8ef91a1b9fea19f1a82dd88f8344032cd8ec557f0ac689fc09128fb080d3cc605d
z22946da31aeabea0294622b165ac5ddbf71a827dd7c7099dd63ec38cb1484d995e9e455567e2d9
zb3ffbffa68c062ae2ab84160e80c9263efefea03fedd7aecf978cbc68637794f3e2e870988ef13
z5f5a2dc60a2e6421fe407c72521a4f50cc1a25f70cd42321a6ecab35dbf957749a8008610f7b1c
zc05db3721bbe655a0b9e89e3cd2c23861505b6b22a4558aa62722c6bb6ec9f43affb33aa567026
z3fcb646067642b38f20a6601e364168981199125eafcda31947491e3b1375092e889059074a43e
z26c0e35c3fc9f9c812cbcf7f4c6468471228df350427cfabcc36c7b4309f1510fe249ad31a6ef8
z749f76406135d357185db1e1d01f414d89525d98069d6ec4fa839acf27e54bea541510f886fdf9
ze6218537b0ca41d7b73cefeb784661aac8e5256742a1a0a8273ea82a0ff1751cb074fa877b200e
z5b8710159255b68f8b38dfd95bf28cf980e9b63dc502379862abb32672779dea9c8d28d946d4f9
z55135ff68a640eb17fac38a24ea53c856fecf3153d5a3409f07d815bdf6ba310d8e20b47c81353
zcacff87c4d423db2b4fc353d82cf2c889b67c4ca648537f93b0895b662eff19219488efe2f5ff3
z3b5d5c27a141703467dcae614f0fafd26fee263008719970555df1532db4ab98b4f9703afd89a8
zbff392639c03f22fb758228363eaeef972ac70c3c21615ade3a2d8880368cf1f36d40316028217
z53c0fa031786d0985dbd40ca664d27fa237277a7948649adbaaf003e8c8daece710ef890b46de4
z195baa639830e909814e4b0ad372e56a88292624a5a30124e9bf148dd890bec9f19ad94e93ae34
z77d61ff65f40230c1e870c624bb108452cf6e10dcc52b6a2e5c10e3b6c48baaac4e8c3051d7184
zdc2ce6478aa60905e08e0e07389a669ceb68c4e8c8454314711e0a1e2a99f2c0999a0bda0ebcee
z4fb2cb1745915c0917ecb0822dea1f5dcfa310bba4ab7e28780aa7b3b73abfede97abf5eac9aac
z4008879da86ef143124390799aea553617a844ca64d785feddf73f54fa42233d1246610bc62182
z86c1ea81727d03122606ebfab7aafb8f7062cd47be3b6ace9c13b586cd391c3b0315318805b128
z696c5f25c85fd68e7faad66d8c321f82133ab7bf6ff2327ba5b42d357d87bba3ef5de0caa831c8
z3ed8611e74d94639bc5375f02226c52d4120a912e6a334399cfdc906778f204fccc566a190da34
zd86aa071f6267c96bf8037b1435c7d581868f7b27b85166e02fe9a4b9da45d7ae10d209f4b8236
za6075237120d380769e5c0570abe3e04a14fdd8c9ff6a5c48ea5d1e019e73a1d7aca4a2101267d
z7df9f1639f2f31d01df5d373ada71c3bed0613ea5839e895f23a7a4091b9c198550edc78a41e5e
z7c63ae0a48570906fe93e9d40e8dcc4ca5babcaf26c3f1989e1fd7c3b8f9f9baee3ec4a1089a18
z945d8b49629526894f9537401aa46b658563ef2249c3f2b8ecd7da88d10ab5bf49e4df1f5ad252
zd2cbb9b50feae7936a47318e14d59be8379beac01eee85909f142f886af3dd26b2db6c9018cee8
z23b2803fa17e1f5981abf5259ee04ed4da28b42023b019624a29fa55a37282434093b0b53b7813
z8d2fb9be00d76ec3661b079bb004bd257f0eeb4071e27272d639b8858dc6b0a8bf546d922f0d66
z7764e096eca114aaea557a0aaf76b2ee98d596e0eeca7fcda5639f83299da66798879acac05efb
z0419b5b3fdc204af3dbe7dbf3763839544241f56dd3b3436dcb84c8a8fbe50a47733ae57e344f5
z48e37821436cb9c149bd220a7c562f96c43f9b6f3773735af1240b22ea5a420c7596218f2021c7
zae83816e9fbcbb339e1fc84aa12930a02859e5c2815621553cc1bde14982a45227d3859960a1a1
zbd366d54cb181c0255d27e3be33adf1b7bdb9056098132eaafa7632d65be32b8e5c6c6d1d4801a
z744de95213d583e43dc1efc0aa355ea573f6806ba00b7efdee2ec5fb8fdf60438d9bd923a4d243
z4b1f455399680bfb63c31f8314b8140d27536d804591b362bd547d6d11dcdd4e8d2227d33e9c16
z4f29c394196f27f8a08536cc0f829197193375dc37f393e0563429f7a62dff87e61fa846c274fa
z14c1bacf508a88940bd24c1db0f00716af8dc26d6ae81169a05654aff9f86db8f1becd2460d8e4
z251d9ee06a09c8a64c067ae4d6cac7197a4928433647060598573fa02c760a6dc00045ef3862ef
zc89f42da31220c3e8a3d57e3204696627640b4c455ca685d4e10d2d9942f205f0cfe14a031c59b
z351338dd49a4e72bbc6fcb4698f8dd90cefa638a88f9a96be4b75f9c80cdc357086a9db89e400d
zbb90c21156f4e3103d20a9a7fa77aba9f5f4e292932e646eab670b2c90f4ec1111bebd78b0ccf0
za0da4f4073e8cd61f9c6623d61d4da1e1158e63a3ab6a58e7c240a4357f1afb664eafe8769278d
ze56d02ee8b0640a6a2e141863d7338ea373adc097e93e5438e6b135a644ee5394dc4e482445520
ze85d6f077e2de66c7a9cca27e626c739374b1dca07fc79e98e698f2edfe293d986e0be8c803f18
z4e7acb16c5a2665f6b223624ba8bb6676be3668d669f7d0ebb591f51af2c65ff7ab00cece42811
zf67939e1e69f6ef1048c1b5ab58bdc5a3f61529b2be681fde4cbd4a0602609594a93c20ebb4b87
za35ce7258d5a2d750e9738eefb98844771616149ef564c42e9836bd4f12235dfa5cc48b6140c04
z5b8c71c7cf7292a010fc806703fb5288eb8094ea98d10ed42bf7c80fd3d0c2c5c18cb083f7a39c
z4d27159f63a00f84562836a4a8a2ced254b490649d49d028835bdd9ce0e7228c67226e96200992
z49dec8fd48499bf4b03b9f3be77ae17b16d23ddefdb91625ad1fbbea38a301a63193c798d147c2
z7b0d46e6a230ee5fae3edbfbaa31e4d49dbbee525797abac6897d574f34f6c2a946c87dfc975fa
z15889eba6c550b44f43a0ad14e3a15bb159c48dd8c85519c855af3769c848df2104a8debb52528
z9a1ce8a105cce506c04d80e79afef2a07c66f0bf52826991421ae04cc5beb0eda7d1490726910f
z938bd4b08a6f7010b81ba29ecf3a49c59b18d30888c8af8fa4551e2f496d0abed7f2384a5a572b
zebc114644a08ff84eff23f208de5c3e432e4ea7d1eade3144aa6843a3bdf70ed119af1677cb131
z8a6cb4ab929582fb2f506733198db8b2e37c3e0a6a3f94a09ca69628e70eb861b5d5a4c74c6f8a
z2a26361841017af38a829475826c3f3947f706b8428af27d651cc208cf6effa4be00b62d51e0e6
z0e03009a85038ea9e93b3984f70ae46c932d5ddb84a3256c96b2735921c85b2563fb6fa7256cd4
z2ae08de24de4c1208fb77f48585943601bba4cc53b7f3a4531141127b315a08672df40244c510b
z331da96fe15fb739ba73f9bdb67be5462b13b95ddac4f8901612a5fcdbf0d86e78df7f61402b6f
zba158772915fd6502b258d79879a861fffb77467e5f0a4df912c41a84496bc0b7c4c123903f99e
z9253149f5d3b5db692a1a49f2a2a4efbe98c9ee0831db29d28cb5b2c6b06266065b66b65a484ab
z8fce69705c45aa38c4571467f9afd7e25d3de4737a6a5c2e8629679ce132c9c0d10dd71b97d9f8
z51c6d7cf7d6c125f3a430b1a120647b2e1376e9684d2f8d4146e38e8bc440a8f583876f6ccf640
z9f273cade1c0f4981477130d5ce661571010b8c1dcdffb17c049989014aecefb56d906cbd32e32
z858845816a10467f95ae8450fdd566097c92329def4f115ee30d5c8d2fe143f0f7ee49ab69b260
z361a98cee690f12c1989abfa37a429cf67e7d6665ea87963efde89cb1bf65cbe1902e5fb9eb890
z9cb99a3c8fa1cfd728e8e5fadd31f4ced7600ef482c19045a8ea37d5741ed2f6688e21f2f1e08a
z6791ba128468062daf3f2803b1ce05692eebc38942eef6de94ab33ad39ca1b344d0e2477a6dabd
z09e16b02fe450df3c8c8ec801cdb18e4de180c1378840397d79a4254aabce3e8bc9587e829b39d
z85c5d08e7f6f9b7ac6cd3a7ef81ef41073793294e2f1ab490342e0efeff19907cdaa6b816e1b1f
z5d9639f09a4aa32296f7e79c50c0f2cf6f80fe48b477c513abd2335417afdb1e0adef900877285
z314946faa6fcec43bc96d9abcaa9ac9639c1c74913e0391f78394277dd272329da8edc3e537819
zcf3a494eca6cb9c7f9cd0045b8d7d8fe0321b1fd889aa033abc48aabfab407930db28316d865af
z2280671cb366dcd21a5cdfdeea1b3f91691364f070af66d1781cdef1d5621f81f4bb1a998e1efc
z0c13191bf17c7848ba56f1312a0ede91494a7b390775757800f6ec4459102b1e9399df2a210966
z6dfb69ee93a5e0dd724c279fd1fa364d26b3790b7431dcf0d98c984cf96ca07b4594346e557ffb
z83cf79498be1bb7fcd4b6377278b252110aec907b83b70d74af330ccbc4fe6f615fb1d270179dc
z64327a4ce99adaf8f59669508737c67aa25cbe8201920f92facc4dfe52f1199263555168e704e9
zb3e1e036345232db2867ee94208b89460927b8f7c4aeb031ce5c98fda1b2f94afab9f78bc8083f
z60900d5a7d7233b73149acf7ae697cb91af6b7840ae2eff15f30a21f8939d0e40054b91c08a411
zec9db93d0865838f3af38b9b9bd4367efb43c5efa9af8cbf03f973343f2288932189540e56d708
zf5152443b9d22eca7de76d0752359b291dcecd9e0141f0857524952f11cf6939d842e4bb7a4d9f
zb94d4915342c7f54a4d15fc34b47acaeb5492eacbcdfe267c1c1c3c81473bf81cc91f935d860e7
zb97a9df12f2507a0a0db69e0d5ae91765c8fc5a5d7e92ae740853c1768ee6d8bb725d8407f3330
z32cfbc8e0d9f17b37fafb33969eb80b3cd7342cf61719fd96c1288d4911a15bdc75c7364bb24fa
z7d178a7b0e696c0efc1a26a413313b8a1599ec768ee99b709e8f13400ba7f55224f3d8c09da133
z1019c7093433a87453b35c787471c11cc848091a3a541e8356cedc63bb7657d4f51be1cd951815
z6011b01a5dc2e582c74790720362904ffa5a66304be42a0515b89c9d43df320fa7974195f3e49c
z721d4372f3c1c2171514d55faf72fb4a8c62a2b0e01375d15365add9c68ea6b72838a73539d5a2
za50ec2b885c9f5433f2a03845b4f2a379807099fe2efe6b2ed084709dba88e550bd294a5032bf7
zaf8fcb02867d8acd0c6ce06ad5a2178e236504d52079d93937ec7eda1d742d2c90e950f2da7efe
zc49f2e4fa8d60652be25c064772866d6af07cec1d37688a097d4522f7de5c4a6efd6f90649503d
ze5e4d2a5f45e2492ea851e73a773bb9f160412402d9672edd024e5620a3c5267acbd4f4614edb8
z0117bfbf9893428c0e32201bb9c79d3060709ac43ca514eb0f4d356352b1be6cc7f8bd800da4a3
z9a30ae1600ee5fc2b5d5974cc343441427628bca80cdbdb42b1120a217d17f17322e24bd90447a
ze879d6e7fc3b4660d175ad35c1d9994187139d4ed1c2e640e15e4e05873c7eaa1e6a700db8b224
zcdb6b0398dcb96a0f7a4ea665c5827706f7e060356e47bac8247d0d14d4a1aa9db9f9571f27d9b
zc537c96aaa180e7e190b2ee9bb45b8f4a08133f94866b9db4122e0585b8232d10717a2fe66c143
z7826ca80b18b64f805a851439f17b63ed098fbf62c0a8d49981717df5b9cb44bf17b52332ae941
z7c297658b9756a2b602ca0bcb814a0a1c41fe3b1e4ce8af5cfcbcddc72af656b0153067cbf87b9
za956045fcf7aaaf2acc54072dd9d996de2fbb745c66d3c244ea85d3b702260a1921f37971b51d7
z47466c66d417bb3ccafce73aee80592f91fd9dd835010eb38a3cd51766d7c914dd81137f783947
z80588ef963c22471df8c647c77f02684e3656d537e3cdd7612b8134f8a20663fa65c10727b9436
z3f5cf48788c6e76c506798d943b3bece2d8080cfc7f27080a828622f84eda65af2aefdab054eeb
zf2eb404c2952ddfe6314bec375a132a58744aaa96bc8da489e4812831d05ecfe43d9d150d75983
z9e6fd6d5c9eb955805b815b34fe4b07ecd6b5fb98e7b38442e24e073df5084c948b85bf68779d4
zc3733efdf8f2762da3c60f28c923eaf0290636f09882c14c5ca8143573ad949ddf882d2cb3a2f2
z0417fe48611e090426853280a4b5ffba279eec4a8e3244af722d8914d72d90c25022d053d98947
za92ba7d35edfb0f6e575a0c15c56be7157e3bcea0b63d560cf9b2bf5de5a1073dcd3a76a006958
z1f2035ca6f99b3397e04a0c46fc6722c8f80225be4da3950ea0fc3837dbd48739e42fb295e2f87
zcc0d71dd46898fa2430a79af90591ff94366ad69d6c43ef519a9ee0750d5e9c9a0f49acbf94ae3
zb322a06a4555f93ce578ed31546cfc8d9415bacb0b4446ad23eb4b3ef908553d51d15326fa71f5
z053c18fb069a2850a63217c5d49ad8aa8256afe0906f39efbda17a07920777b560548ca6064c2c
z6518473d6698f19840e1a75f7cb830136c4c5d603d9ea9dd4ae3f9267f33f3fbe2320329fa803f
z9443803e8904b3dfe962c90d31934b996248618a2236b41879db58927b54df317b5a3bb0c8a2cb
zbab39a86ecb750fb3bc708e544693cd40d636098e5c7410fa4b661c8b3fbe9664e76182c196134
z4e3bbe4e76d33ffbe25590359714394c59479266a8954271f39d1594a61aacbadd2e1e8d5ba640
z48b7b3df0982b2f0bff53bd129edd9e5df90b7721d266c77051346cbe1d6ee64a55ce848f5cf0e
ze4bdb0eaa24d0dc1b54e813dc65d9d6ad53e5aac79ab6115d53b8fba01aca7cfa2670723006982
z8e5b8f5778c8e4824c65ec92e03cafa1b82794214bb6ee70974a982c8a8e2397a95617b9ed2aac
z1423688e523cc8c46bb13bd8f918b09e5470f2927c4c5cce65321403d6db737acb0e03a3d2de78
z10c3e3e70f8183ba14478e68bc26ad5c3647c70d2f8fa9421c129364ebbed650cb97ee76ceaf41
z8fae127a94eabf2c9ed935433ac5573acc7acde35871a4e131c2a0acd39b7f39c65fb7e667038e
z386a9fb844971fc7c57eaf45386df5280c527354b4c5cf29e63d56861a6faafad306afdbcdf261
z5e8cf5e1adc622a78c06bf617bc3bbc455c346dae1e2b3b4010216d197a297b747ae5fb2db5fbb
zad29bd75850018a94506f196a2a9e9d50888a53616bd973704aecf149b6b5d6b66e6267d28ec59
z58945b1532ef687c8260809d1be5d5fff6db0ff77ed75819fe5728cb7e98403ef981c770ae32ab
zdb33279f2d37e1dd7ec47b0e744aaa537ee8ff50ab324dc3a1da555ba2400f11156d37dd6a28b8
zdf5fa14ffb5c5319db6898b192ab0fc433cbbd13efc1b59a00229691ec7ea7d5a19b5b9fd3c626
z03b4a379a090f77c4b5f9b6c4f185f747c2d97315f5a1847e2f349a65fe323b339aa9cbd5dd8e4
z6c4745e2238e2059977338b8a4ef23e0911e23d6e3ea9251c849e57e2efa3db4ecb3826c16f910
z92cd9ce63823bac634664aba07d2ba1dbf28785560237b2e11f421d78b79a00677cc868561b4b0
z31a6e2f353beff15b54df4eb4ab9b5ac94c5f1bb0dbd9da006232190b246cc0749bccbe1c7a719
zcf7d5ef7d8e55246ae00e5290d8b8f75a019886c7182e6e55fca403d6e05249527826ef13bd2dc
z0ef809ad9984af0eac9396e5b86985dd6546ca79467ffd01b62c84d9ab8afc88d454efd3827203
zeddbf0c4fa82a0bb7e7d38103fa84896bb7f8abe3b7b160ccca60c63e29350e47dd0a62e890f72
zc608f84f4eb017ab2e3900c5b2191200c3796a4e9ec8428319cd591a297a4e5b17cac8720b8643
zd9dde6c70b2b99ae26758d51709deb5b8cb9373ac48d06c5addf226f60e2a9ab84ab6da2f68380
z14bfea531bc04913144cd9f9e96d5e904d350d0b84360ab1f66e7e51b97bd379096bc2f1148ebe
z3463eb42d9e4d6503c37a912a73fd502e119b4087964152e72cda8ef1a3fc0648ff3a3a39d633c
zfd753844d76da1bfc15017b4f090acbaa01fd408c0fcb5dd43fdf6b1c9e31f2a306f2463d6b43d
zc6dd0092fe0c07837f0cfce79f3c1b064b4841ffb43b890227085be045564e1eb95d299a52c71b
z103e911cc1fa5085cd34b4dc7ed7c8e07fff8b35d208ba6eddd013153ffa1836a690874a28eec5
zd999a0b86253322bd7517bb470fde179aa0c2b924ead0729d30b4c487dab8faa8db451e5ef27ec
zcbc10013f0422b488601a4c45c3d0cc4102390cf74838d036a065ed06b1afae3ab0d3f82c3b699
z96057c96a22126f46430dc91500efd15d8d45167bb214f26ab142c311fe347d17441b5e0cddf4d
zc74df60c45661a3735291a85d0ae57c037d4a2202807e99a5722aafd9bdafef4960a44b38bb1ad
zef7a06810195ea3c6845a6344ed705ca2dc3eefde55f86e306b2654bf57e832fb9abee1c5f2429
z0ffe09911eb541119a8300292f4a9592314f75d19c00b751b9200a53b097a03e49e75d6bfb4241
z645fe29a1a92c4b61f90fe635f3afaa197f720ff59b0a9fe467feb7465be6f2c228080ce0a60dc
z51b2b15fb5425bd42ba7fe974a79abf6a765c44b175051e515146c40b6f35f861dff5385ab222d
zc8bc93ce2e1b9c914cf3d217de8e2febc5fd6a471de7b05dc2e8b7411515a3640a09b516d1a226
z7d709a36d5a949668f2d307979afb3ec88b0d65d2811840b85e1b961afc9d9bfff011503f1fc25
z60235a2d373da8b77ab02ff89ead39c7d431dc54aaadf5d5a554c5264a8ab7b8b266b6155d9ce6
z7f3b77d3e11661e8f175709cf133bb43a0ec86615359a756a887596b5a2d028973f80a2810a6e8
z70c716212224b86c740ac3a7a4f1cad653d33114d02762087b7b7a27b54ad933bf481d5854f34e
zb15d903437eb5285f97a8a6f8adf9f08e642a543cf46e776f83fe942e97a8b983e3e33cba5b4fa
z41ce5961337b7e6cb99166a4325df0df38b0509b16b372a6b3788c0c99bcb34563b5329fc64c3a
zc92e31cb3ed94e3320d737b75027a35331f7df4e8899da3ee7f157dcf07c6fa7ab946f3a4659a9
zedec9a557acacd511c8890601914e0984e673ce27bef441defab43c7196bd26bffdecc8bed886c
zf915b37c6675344be5ae1faf0727eb909b4721425ce0b83eefc27a3148a1907da6209df83a7982
z0bcc62696ed427e7ed19475b6f8a6ed46a96183f5b6d68794708f75d18feb21a9ef7e0e5d9e506
zabe6fbd6e1b94359c908d55371928d2361b0bf397c6f4aa4aca978788622a5ab9ada43617b1ffe
ze39f25333f5e53906c246189c60d3cf499d97be7967d2ee0f75cf88457bcb03d5dc4bcaad9f28b
zc52fcc45e4c1087e7b4c6815d5c99c92056817a3221ea17cf9e28eab53db717c69f801de8a048a
zd9e06d8e7f1703d6a94e6074a94dad22063efd24bed5e23a377ec2ddd5df187a61f8ea9d88388c
z3c4594c345652744aa8ade6f4b1aaf76569e62f061124a6e385d5660ebfe72ecad54bad3b415e7
zd88cf2d5a5c41c82fa98f17599172454554228e4ded1a443fa6104ee6e8ae783f86fc2fd946bd7
z0c043514ea1415b44d151d1e92d514c5b8bd6c6625c3510d448ce151d0d34d4959a86388b9fd15
z38848469127078b14f1c230ddcc7e0bc4a38fe5e71c2f3e0dfa34fe1f6c2473d4e7e5e6745f8e6
z7edbbd5bed952f97715ababc90c941896604dd6406e87c7604ee499aecdbd1aa5fef31572c0280
zf58f276fe1977021ecd9e7a096a2b1299bb45d55f204f165f8d5cb08c6f4b8f8b98ab3f29eca38
z1c1b1a94c036d7a2d382311411dea5b47a3180749a049bb740d23027ca3a2edae055b79ce49056
zfcb5c5e468da134f18c34acad05a39a249a53826e628277671dc62e9e51c54db005c8c9d40dc59
z6645e9c9672da0a1abd66db00c935ed2d84551da4d7b9768047f8fa9f171adbb7b9edaf8e2062f
z09e9c311582f929ffcff1ebb56378be1ce486d5dda9d2e63c1d35eaad8550ba3f4ba83224113dd
z95bead3e8f0c9dbe1c1ff786655a0faf2730840146afba43189ddbeef07c6e0f955bad76dac458
z2cdcdaaa1fa081e265f50929834ebabb9d185f887153bb57f3ed1d1b27de1fdb2a73b23bbaefe0
z787eea8c032862f97b33f90f744d39e79bb8218d654548991456df6f9e90c1f7a2f486c12ecc6e
z9d26306da0a03ccc370ba9f98f4195c5687e38677b8453f5e87adfd22a3ae091fcb517df7c121a
zf159c8457b127a76a5a49ca3c19c70239a42938b67ea2d7e914759f07f652296934e5ec12c6bd1
zdb8e890db3c6539c5252786f88b115669c4caeac0573e38e0c4530efd0ac8054667fa477f734b6
z86ce355fde445a3da0a38542a8b3f37e32a05c2f492d1cd75e4a465dc2a19fd4faf11b08fffe71
z1de9ae90fa1068e21261d8cccdf585453298c46124a39114b506529e63b07b64f82ae59fb73a65
z33bae637707edfe96ad06c56b17992861fd8ae74a5cf06de9d12a0eb84c9af238e2d347b5f748f
z70a3ab5bf3fb27bcd35d556c2be952eb7f7c969e42f0b040deeeed8cc16fb72fe34b465367bb80
za9f32d8c9874512df2f67fced2b6b921442641313a692a1169c1449d29c1acda0735e0604b0073
z1d5ff165c7b74c9a38c236b93d07048c8ff09236a1221c2dff348a366cbcfcfafa597b891d6ea0
z013bb71d8ea6e8864c288b1ede51a832e1cff54c5fb321cc9839900f3077bc6b9ceadc533cce85
zf5ddeb13dc1ab2c764905ab7a97e1886dc73c27db2e571ad7027b35c069f16c87b96c10dfc6115
z6a7c97276281f67c5776ecd5f68761ec673db5b8d8f3393bf3411c65855b444792155c82009bfb
z05f4f50d7bc8b37490029643036bbea4f9b87a4823454ec9f9e269485862b61b2bca086c38f2df
zb7a0ef08f30d97d08f0c41467b0fc370e7846cc690b45d5a8b691849c3d815487489c58d5ce239
zd4141ad3ab4c55240b12370a573166ebf360cd916ba3a93874524fb4ea87ae793fb421b799f0ca
zcdea19bc9085203d74258abe6617d6a3062cc1f5869302f2472497181dbeec8ae79567a4a6d5f0
z9ce0289062a4a6bc703cd5dae30cd12db01bb346a5ef997b33559d322896d7a1501608fb5f621c
ze1f6405c949e5f0e8a6020a11588dc14603d6a5d3067dbefbc881982eb6d08960d64d7cce63c61
za89f6341d340771d6aeccd80f8c29a3b7a3d16579d900c1e6f28f44d713e68281aff15b37550f9
z9da9e221871ded7be57d810c16226515db154a782bd573da3b9e5e4a6cb6ed156260c0cfb09dc0
z0c44556d1d2712625edbd7df2e4899a567cd6d5ab51e37974ba25d78d4b9bd8db9048a4e8a1f69
z59a8f03e1115bcc242129f7d92873d3344f939dbc49f21123a88aa9f43e6ba2b1ac519f925b209
z72168c3467b9dcd763224067f7f9ef11c76f5d27d49b3bef9b757ce1303ad7656b18fa356fa11a
z03df0b58f17bb5ff06146746c6200153610a641f288d621a9c61c0da2ebaef8f7e53c757712427
z3f50502c8e068625fc0593505c5aa647a02250b6299246edbcaa9e173c83c058586b7fc6484a76
zc8a8cc990cee5c6f0a7089acc32c07675ce94f30d99eddffd9cbd3a4e82cda28655ac5636d5ceb
z5e5ce8c2b68d408cd4351f7fa8c59152fce6a2867389c6883f48f8bb957d2c4e0b2b858dd246be
zabb0393c44fb7e4e37240be337a1f0a1c8e901cec3d3f2e3308249a5f7c69ac1cfc02099e1d6a9
ze2794ee03059851a662c066d11ecd6c49f73c15b5cb970570878eb6c1fca76c0aab32203105db4
zf4d4a8ee527c811fabca421bd46fbe5de522750a8b7e75d728c71867653fd67a2a1bc24148a941
zb2d1029fd70c59eb8052e1b8571c5a33cb39fa47c1686fadd9fafd8b26f16a075ca584042efafd
z484383a30c0b71a46875abb3c4905566169d0ca36496473eacb84fee30a946a12eb4f215fd36ac
z92b0bdadc75c965a6ea93a1273f5171c36b165b687f4d5e6d489127f0501dad45d8494e3c345e9
zc34f8a25c1cd534419e2dc7df5dd36136a6f9b2bb5879556fa312e306c444e6bdbf92d4f3c0bf8
z0ac03e0d27391b2edae73a1c547e56533b93e927d3e74051904e3483f769df8429655840af1485
z2c36eb0d4a67976648e30d53de2cbb7773a1d45a4f61b4040e84ebb27c2364ba173e8f1e1bd039
z07dd6397eb2f43b9fd0e07da37a13d7295237a9de7773f17df48e0af8929f076e4efb93eb254a0
zf4c2da029703575b560a28632073d149256aeb1db4a8ee387a558a652cbf365aaab9ca3745bae4
za855d1adb63961d392439e0b2ac7549398d34cc0e613e9425e5f9d5c4b6f19169a3a22b0a6609a
zec4399c6152cb1f28e76152f441c923f88abe9f6eb3a2869314a7f1b0fb2cff3cb2949c1c54bc2
zd3c6b1d9bf3a9a299dda3328fffa57b89b8715e2ad7717b285ca6abd9552606288070402a4da58
zb3c8c25a8f722dd9b47f30295c56d353d989eadddc1fa76deb30753b86f92096c3e74224b86e78
zbcab01e77ecb1f4b715a3be91e56bf9026bc5a02cb41b48bcddf2b0ef951580d8b4ac9cefe30f2
ze645cc4b1d1bbf08672137a5bfb8c036a782ae5699075925686c49ccdc429bb3e8185758ad5846
z0d98f796dce27cdbfc86a8288208675a47b3d506e2b80e4b72da1b3f2a0b08de8866e7caac9ae7
zcf93f3f9470bb17e9da8aac63636da8d3650bddb1b2a1a78ff22d9bf23f6886491f2f23b6422ef
z71c47aa1b4a091d2e8a0db0d2e3cd8f2d0d95a2bdd6a9ed0cb8493f05d1e7eaf0ca3357d026417
z9387f0c10a6ad97ca8be6202b772d7c1bc0de6790b7bcca34ebe1042d4042f1500b9b7e4cab9d4
z497f186fddc499250f614051bdc9a264ebc5336f00dbb364c84cc2015188b7c9cad2705618905f
z74f7fe7c6c0d32f13e84a118f3321c200158d650eefc56ac142cf1aa2b7d033d8d548d44273b77
zac185a4c66db9afa305aca8e709cf8587d8151302e444878031eaa5cff14ae96d3cf5b2e650606
z61c6a1dfea47a2ba4898c27e9d13f72a2cad89295b71399a072848c104409e6be816351029a245
z7c6665cd480ce6ce7666c0b2b5a2faa2b37efaf836a7700f3f9fa4765968de0d65fcf029dd2321
z0d4351a77ddaefcf8c54f197865b0b07e86260969e264c24741b1df6374d8254ca01d2fe56c616
z2afbc4add4e22bba370fcc4e7a19e1fbd2b3bb3b6c3e626ca726c357a0a8a44eb076a29cdcebd7
z0e91f510b000f0f86db7b1b319dc432a629e4dbd503f49c7ba4a2cc38977271cfd60dc47352d3d
z6d436f9079c4fb39b406dadc39e48a8485fb436665a1f60026da3ade04e509c2c195d6ac6f7870
zdc50bb8789f66b075b818f901abc9d1e38c818d8e783d10e4a35072a647e71ef66637f2cc01b23
z4c8af11253f1d6b3bfab0c1ecf0d911f5eb7050abc2a445a46c44ba436cca04eeed19e7d3fe959
z9153ce0f4f1f4e21cca88927855975a315c1ce8dbde00d2062b252cd8e00c0aaff3d044fa367e9
z22bde2f0df850f38fc5c6d210baee4facac022ece0499f780549de6aad865b0c2fe28ebe42696b
zf121f03dd5e2128d59e4b793d59c65f7fbe660eccf6af8d390308bac21e7cc910b3f7764f5ebc9
ze997199a60943ae83be04655ce5a9f9adce93a5bcbcf6373ce2b09bc4ce58d77a552abb53171fe
z0cbb30583cf36a657f1b5456a1177508d858b8bdb800b7ca6eea218e173a4c15b829285d8e6c38
zf3c080b974072105a130d1d74e82fc1608d0a38aec0160e0f092bad67b65274dc356a9235ad4fd
z1be0b8358a753ffcfe87a00a601f787fd35a97552b244a69622e11135452bac5cde86849c7182e
z501b5dc83b22c1343a506e9399165455e31b9275b64f50aaaab6d77089d3c83f67608862074121
z45d9c336a8ebce11153c089d2e66c010a7f1728ab9fa6a154f7c90516ec5c3721f670c10275b5c
z4ff7dfaedd717b47baf322eb949dfcd20483d15f5a32dbdd0a18fb7b1539653572997a236b7eda
z8a48b1e8d72a15866d216b84b4e4d1a6c824d99d03e6b9fd53af5d81af4a30431cf42e0a6d690d
z8f6af989caf3364813cff06b90cb639c38ec182eb389f3c1424109115be51256a45d64e8699ae6
z3242c007c63a27c337e0d48037f06fd68e441cbe52b7dbbcfb1ce4d060698a5e02842cb087d54c
z5b55dbdcd19bdc7f41661ac68d6fda918d545c4dfb2410e565507d73247fb6f1bcaaf03080c64a
z85d199b7f1d27ca24582196c692cbe90225f33bad26bbbb94bd291acdc77a2cbdeda3a3c7f5419
zb34edd639d93689fe3893cfb9c7e7fbd20288f15b55a1f275ffea67c0d0884ba640abb63362452
zd9cf28faeac422995f0ad602d9d4da07ec098999d52b8c169e473ce4f614d60dcf7d9830ecd440
zce6e6320ec57d1875713d0ae8875d6cde73098d45689c7e299568b5ddc578c0157729c3b66629c
z3049b7570970b4301c9eb25238130da9b938ee20dfe7e9d7c91a0360adf92952c406318b64a943
zce01df15c55b053b6d45c1147fc190ce490e96a432447d6d84c8498aa90be9e2f10bd0ec9708f1
z792241617cc70f64f0054bca21b6d4cb891b698d99f307e150a1c673c752948175b89ffd477cc5
zba04cf72eebf4e0668f924bcfeacbf46637de20179bf5698e0d9572da1bfb6799668bd89d310c4
zc2e91c3bde8dceebb2ba28120258b7171c9764199299486e8c30079d6bae2e475491633371c7dc
zd12f3be252da457806e21a0d99525f5dd08a75f57ed8d2b9c254a520f474cd2e279c81ebf22a8d
ze1e1816159d7b342d0a7228b5241003e6f7156cc28f0305821645a7c826cd69109cd35bf43a94b
zf536a50d599090c05d6dd2b6469a6b006ce246eb27b968e43c3d1c638ef1566264a62282285689
z04bf114e80093ddea4e9470577a040e3bada6efd3ec8b1e3bf1c13b653a9b359ec3572f4b9d988
z422badd84ab33218a0d0a603aa165e8073baaa4f5acd0a0426a143c6fd602fb6605d047972436b
zeaa6fce587ae74385b18eb22c448bcfa6852fa253b69896241618cd503e6496973358fd5691d43
zd9b4c002d6a758e98f43648b37c221a38fe7536086f72751f929bd08539b5c400b056be0abe0c2
z76a64f950b3cb68c984aab52ee77c944ed035a75afc3a0d3f55aaa022bb0426851b8520b303c7e
z38e4d9672e6eed58e10b3af6714f129938e67d99965105a582137d9d368b42ee6a54fda723fcbf
z2757056bfccd7d93d0727c30482a2adb9560b6ce9a1687dee866b8f8b0994827f74a4a45a1d27a
z8fb4e7c4a7654201486f7df5cb57df5b9640c75384137fbc322c1dc31c09ba08354f22ba5e2bea
z01df66359099c29229db31f9ed68ae63d20965156d288179f0641ae9bc85a5c76b0eb5b174a55a
ze94338ac4ca4356edc7b99bb00e49524ebb5c01a5172875da9ed9f872cfec0e1e1b9657daf5091
z0eb0173ba619fb069068528add032ca7c0dfeac58dbe11dafe9223c386d5503dc813e9c0f52d14
z59d2d4d51d69da569f0ffe05944cfc56a89512986bda2542af2fb63bf93d921c4e3c88ea310a61
z287a8d50f27ef1696078c13b3b81a9c39bc623a2d96f92dc334ee0545441cb98f50b1e4fe2d854
z7fe1c52c55f406930b90574a41840a492110528b6bcaeccf06d020026c103118f6de08736e4c03
zd50eda23ae929760c93580da8d8b05c38d7f5a3aabe338cd1b02f7d654a03be662e24f1e8cceec
z327b24bf107283b3596b9ecfcbc02a8d424e3b646d1439dfc2d91fafb00f775cbf3abd0644e0c2
z67d3c5be29f5dd673e3b9827d901e3c72318129cab2d3b6def29c120cff95351162031cb120266
zb87b5895db73ff3e91f6d3e3e0f8bbc6a99db7d1f255b780e9f4e9265977ce5f9c94afdfca4ce4
z4a3daa0363a0c54a4e4b7a83a8f8fc222e9ac596d58e1bf3de26d480384e95ea1e095b110e22ef
z0da21dd14aa14cbdc8db40451417971360578b78fc2c02f0a2973b0233b5d435d588bfa00259ec
z063a2560631105786ef8e0cb7318c5799e8e3a36e5dac19c0cbda4ee394515247d3564a79576b8
z7ad33fd757f52f524a4e8af00fb2969f87101c3f1a6452b85d6d41a00bfe41a78bc4e0761fb2b3
zdfb5a289c24778155ea5153acc9c3c81a3b846d85deb5288495fd9e0893d4290dbeb845ecc4176
za47515071341562fe97c0a096098d48441868fc6c7e54724583aac0abd59a19e667d3311f3524f
zf6d929a6c17b337547bd76e9846720894a4f820bcb2c8aef1e991929bf5671ae6ad8b2610ba324
z8d076be60720504ef604cafde89031edc12b262063925c9b5dfe9e7ce55f4cad41c6ccfb11fb75
z601c74ec7ef274b481d1973df58392d66423d997c3eeda566739c20b1a2f93a8bd3ce7152140c0
z4eba5dd8947eb05bd69563ac9865e6240491d985b319cbac3eb39b467f168e70f2155e05aa0ef9
z58b69506fe066118382aa828f16c4c118b3bcf4c31f8d350ea01d85e5f846f7a1a96229bfb56dc
z4b91615ac417f69bb1f1ae516af69e9b5f376b1c9b90f2cb2adfc2f1e6340543eb9379b90dc38f
z07e1bc5892591b447d95b07947ba255d5234dc050d5bb91f8bfa0aaee8630a60cacf838d6a1c9c
z0dd375670e58867f86c1c085f4b55fcd743b85626e77de69f38b6000b11620c0ab140b8a53bc88
z3a3fcc1a47346524c93200446f589476fb27747123fdbde8f6ff1717c813692410b5893b391893
z5900885d670b3b9a072fd9b92cd4f7b240da428ca51cd04a51a39b107bb053c591ebd548f91441
z00b73b7e58aa3cffb0a76497f572ecca63a1c079cc0ffe52d08704a02bb0f4d7af745cac6e0d99
zb6da98c78ef34622a442137a22829145be54b1d22472ddd9d245473cce36b6e50e4ab0dd17a648
z0fddbca33375d401f7fe185aa69ea4d4987ee63782dd476028c5f362e7d95abe5b284769121520
z60cc252e459c5f85fcce9befce6d5cf5ebb95b5325602990197a194fd65c2a323fefd0913b891e
zbbf548bd239a2f866d56eec3e94f028542642520492f3e4b84948858ae446c96d22c407c230f1f
zd1e8051e03881891019505ac3a714d8e29bdbbe1654b5eb71ea9651ecf65276bcde4e3b7f7faba
zbd9058061b527f6d5a35b3ca53671bed66bf6df25bbcaef96d4a6232431de1eb99b41a6850da00
zf35d8e6ea2e5ef4606858e4333f5f953fea46b03ec2bf482a00568740eb654b28b2b9aa25129af
z61852bff122e928ab715c46f8d7d4d46047898d550ea91d805797181d6ca4bfd636f210bea8a83
z3bd5aee69bc51300bc1ac0ef26be79322d19b5ec092c760478242e14712909f5c8edadcc4b545d
z14620baa559d82060467f412333476070ced1160617e3b30e53e0c5031f3448b9e8c4962e274da
ze8152e07f357ca5af38b5c26d7bbbe2dbbe622695537d0ddf895eaa9cef4e0d169c0e74fdb6429
z0f1f3edaa1966b466f1fba72f68ec340c860a415b8c65acfd27644923b58983e6cbb555faabc58
zcb68885fe1b7540d958d6e105eeb48e81f36ee5337c8b334dcbd74dedcb0bfd3c46b4c9b1a0bce
z6dc563f47b017d6e48528d7747a1ed3548cc3484fe3bc3d53ad8cd62043f075f6c4ea2ec935823
zf5c9bb6be162dddb2a3123cd89a90018684a0c8cad39e69c5f49c4fcb1a93a37708ae36d5a3c07
z878fa4077cf78c30bd8235e6db19d0b170f8120ae6ab895557400a0465220a2b6de738211895fe
z797489c7e9d2dcb85c09c526aba463adc07dafca97561b26217890903a52c3963216186169f2f4
z78acb3213dc573d1ad0ec81516cbf645fc3ee61aea99a6cb6084241931ba6f9252ede3ceab4c5f
z78698bee284fe16c57fa86e526d52c451f4a8f5930300b62f2129a271a41d73c79c93b071a027a
z5de078167d758515097471c16fb8882abbfe138e3fb5b8f2c4b8628e9d1aa999806a249f5fe6e3
z8936f14a6afba3da4d6d43d37d363ceb33664585723fc367466238c8fdcb2b299150c778754995
z7572baac4befb993a1e0fafff980fe85eb1fa907561587a94d53dd7fae36884838d4abf30a649c
zd0b5d72fd4dd6922c4343ac350e7b23aa0656e76ad577449ab5d064f0ea7809e82c234e434b786
z942c11d2ec5c881fd749cb4260f28767a7595f01045b53b5f9f982b7e470d2f9b2eecc86956e9e
z0dcfea8948efc140ed7d989c1b221619dae5c4c044dc12eef11e52246af903ff1293b4fbf60062
zba4a2b639d972a541cc2f55e4c8f7793d466f525417c3b40159ec2d7c5972528a782e87cded24b
z483f9ea87627233ebbbadda69e0b9488cf72919fe882d0d9aaf94ac51336d2562190a6f0b907ab
zcb2587f23cd169873995da44dc8c36d5cc213fb51804ec5c73f62f078f5fe02ef7562c74341ea6
zce5688e7023cb63daa4be3c949f8dc2e14fe235ece45de1ab144cebc1951e29204436cbaed5384
z5d3e42fe47782d538dd281733c0cdcae0ce7a862f619eb4d2d52b377ea4ef0c43cd17ecac85f4a
zfcb7196e2dea5fdae898ddd2db8c9bc1f6610398d865565fb74ac36ab1b9fe57fc741090f18df2
za7ab30fb070d288a387476233b8d45e48d28669edd7ab65bce11b0a03202fc1406abc98311de81
z220e1760cc50f6ad563a1b2170c271dae4667243d69a8cbb86bea40b7a39ee319374d477d9d6d3
z4072bfe9fbac4eb249cbaa6d4d1f665046168987480f300bd1cdcf542cd73ffef2eb19dcd0b7e1
z00c2e4606383de40724baf099df46e8ce747e6e27cd07ced34d7243ef27a0949bdbd0100ddba44
z7e1c4735e2743fe5d9700230a08b24ec118c05d119de793257972f0375ec2a9e54569800223f0f
z026844626010f17d214e964fa14485bc0893c06ed4fd3603c39953595a4fdf9af44a6b8c4eff10
z95a3d1a1e4e5d7e5e8fddce59b384b73162747b3c7c794a6065bfcfdc2012fa82cac8a6419cf3e
za24ffcec01014f9793c1b0fca695fa043df521a54254f6dca430fea3040ef4c512064c81e52dcc
zcabe56e92111ad3fcd61ff675b820e0bf0c635cf0f5f1c4f54a3cb3190abcb1c549eb6ae5d050e
z74d97c9ccdd9e78634f0c62039b4194b51e3ac272134b8c4e33596ee7aeda90a7e7276bcefcde7
z645e359b49d1c68ccf4f3337c8067ca0e306aa38d2eff4bdb78bdf5b030de66f7e4ab9ea259d93
zab848096318112d9b19a67b01072a10a2bb2380eeebd31d7b67a34ab37991dae457d7239a7a6d1
zd42044c9ad3ea06b56c017ddce0f7052cd2c8e3699966e9c9f18986409f98acd1c2ed4fb6def4f
zfbc62c2bda6b9c6b3e4a14ecabd02a43d2089f18837496b66e79b8dda702a3a29ff0b235397220
zed722f1b7cb51734e69eb996d36709801a5db70716691901f99886b1a6a81f55908de80c6a053f
z9d4c84ba72f1b817ff3a6b35e1aa227913437518e7df42b10ca4191e0a5648240b4959824cde4d
zf95f25cafb8424435068d7e5ccbe3b1f8699ce4a98588934779576d75fc5c0a11d39e6a3664deb
zc3d9a682255eaae2e659bc9eb899eef67891ac87621d33b5135fd1efa4b8fc389e744b55d9b188
z58f8017036fc2ca4ff9ea40a0196ca99084d335b37b107b2da90f8f45282e18e0d6c2604c16b52
zd0a678b802da7423e7f4cc8e240add9a4dc6ec19dedbc51a21cee94751f8a56a2eaa5c4c904cc7
zb70d11ba6a65334e5b4f63cd21c3dc8f1dfe54732792324ff8bfdce6a47f81371ebfad55caeda8
z92b23a3a87388775b2cec1abb01d1a0ccdc5163a408e0890e112ccdbea58f11ddd83a4fd488dce
z970a45c5ca876398c6e9ad045c400128a157c3289e9a5070f0bbab132c2532a4232ed73f42ddb3
z27fe0fb2a8b5a643ea2b6dfc7e1f1fdc860c749254fe7f73e7946384bbe794dfce1c133d9344b9
zcfd7a3ee5b6733b8154a375dbda32d7a1956107fbd991273971075b0a5f74867c3a364ac1c1ee3
z35804fd6e67f3b56d3e6da4c6aa946af0bacff99cdd98ac540a4738217b50f02b9387b4fcf7dcb
z51a7870a91e46bdb7db8a39068f2d1594e9cd351735a1cf5a6861c92242420e3b3664e29306dc9
z8018764bcad47d7468dce6138946b46edcdf40951a2adc2a75b33d4004059e20f06b7de59de7cc
ze05f13eb49feba0591ae8c34e1d286dc8d4a0b7503e4c5859961186c4811b95271395248d96d02
z48121f8b1eeaebc3c038f051d51eaac5e55c9ecf31ba9e9ab915b1ca046f33f8fc01e16e8eb4fc
z469837cd5bc45bb0a29d512753b9611463f7c39de48d2fad8fb5b182e9c5c0186f0f0052d108cb
zf8afcc1dd84b460886f048e5c726f92df1b76ea251793ef1dbf80b30865c48626ddc8a8a966c1a
zdf8abceb96c0e59bcf1a4dce7e52b54fd8e3b679762ed75313aa0cf3ca845512847ca1e1cbdf37
zfa4d421b9c62a1af7d29db8a2e8791804acc1c762e0adb0d15c35ec77fa6b9c808ab6aa5667830
zfa2a7e9ae8916b8534b7f2bde46743f2d198d779c19a81be49c3df444bba9c3edfb8a03c0913e4
z5551495ed90dc59beaa3311b7f285e8ea9876895e51951f64215686ab24aa1841e5eee65bd7fdf
z0d840ccb7d984485d1928ea714dca2f1c54ea6fa54b987bfda642b47cd9f9af5a1fcb1679072d4
z55ba59b18642946725e05025a3780a3941a0819e6aef16016b85b0c3b27218a85d981dbd1db5e1
z9ff958d2efa6cc59a7a26e645d0fbcabddae1a0ebe0f22c2dae4e339367e27786a60f946fb58af
z47d785ef506aecdcfac7d67f64e3bb5c7b34b7d7b32602b5a67302c642d0d103494aa4212d579b
z5c632788dfb2f2381a086c005408815c79289b2c1041ac82f35bcb8fd227ec1cfa67259dce34e6
zcb9b47d7e8fb7d4fd9433776943ba6e48895af5439606e04cf1b6585aed06ad744275229a63530
z4af2db5bb67d0919ab75b3df1731d288db3e733849d657d06221f6bd714926775fad822cd6557a
zafcf4ebf38047bd4734dbd805a5f5314b6b34e1da06bba98fad4aa08001fbbbdb4518d56474a11
z0dac35365a3ac81d121b4715f77ed38e0596fdddd51accf0c7041b0cadec736cc45c0294451785
za9f36c34540cf0c4c7830cba7800bd668a86d5f4709ecb8dde49a8b6fbdffcece38270bbf267fe
z7a7a9b3d7f118eed485d41747b3a25a92bd0c994782029620379d8f0ea278badcb8f68e9a16f19
z99ed8d55fc15e5e2cbf12f2104a56276fb604079cfb25e4ccb5f95e9b75eb38bffd159be6fec68
z23b494527ca86efeaedc90f62955cdc3110a01f1665a0d1289a779b3ff6311f9d98bfbaca09784
zc98aa1d9268b9f46e9fe1cc8167ce876f8616e615806edc2d151f72d916fa07bc63e449ccb7011
z7a0742181eae1b8f8abeafa293b9383502ada82a7f9750a87cc8d42af9416252061433c6dd6ba0
zd00d11a43d583a40f1c9496ae6df70a31a0b9a037d951ea45297c4b2ef98849a5ccf0c6ef24dca
z01d2e4ba5d82345ad07feb8dbd7c1a7842915f13c497c825927a27c4fc1e46937d718b4bf6c6cb
z9d405b0703d81ea67fff08abbaf9efb9c71ca19f9a6900a7d5770d3082bfe21bbcc274c39feeed
zec01bdd772020d38b3cb0cf06b220ccaec346884cda1113d73d879d63ed552bae5bb3e2ac85116
z5b6a026f33c89097f0d7d5e6d145d858f42f84f571789a21d63bf420bdc74eedb0b9ec7f5490c7
z8f0a68b1c1dd91438405bf2e1809b21d55cdd018c760bdcb100fd5cbbf1e80919f730ffd747efd
z48e713d7a94ae24b98cbb70555f14acc60093b80e2213cc764e551a6c0b780fda4690a78e917a9
z88330481fa8fa81065c5cd4f7b5d7f4d83e2195da9e1017f308c3f34b8bd296ea51b6f15aaa668
zf9b76a0a576a23ddedee02852227fc8cda6e393b041bee1046b3ffc58e3003572e9e14800ae1a6
zefd7c6d52b62c162301542676af9c2d3f3ec07bc10f141b3343e3fa04c91d3bf4c37a859cda6b9
z22e1690644a7175d6ba9ce49d70ed6d594791034d5b1b8628e55d58a2ab20742a1f650a5e6dc2b
z8e5d2c33086d95d56b662156189d214c617a88c1ec3710926b04e53d7bf0ed585eab39fe7268d4
z5b914c540b9495e6d4fafe5e58e2ce30cc84b103be029113f4586711984f9c1804dfb084a7caa0
z06e7df4ac6f3d2d65c81557b78ec5870e08709d07afc510e4a82316bace50de25f99ce5eec46cb
ze5cf5799c459f9a9e167089714bc7bcfcf4a88386baac9709f60648716b0dd2dd9a4cb92909940
z7f2b609090a3c40309ae38992a17cb2630efdaa9aa28430630410da390d5db8464efd56d7fdb76
zb03f06e575d553adb325ae49622bb47a632737c83a5e81f50f877faff4256a94cedc91c3ae3f56
za4185bda8e8f4c04889bffcc0f4b9ad9e5d51b73751d68036531804d33f0c94557ed63171101cd
z47e6c3beb715a602dfe257aada707084b41c7e5d14b2b668a00b175403b415b283e0666bd0f0f1
z6a83c25f126910c41c8392f2a62bf2e409615db9fce3794fa05aebe0ee4f150f030985addca609
z66e5ccb040d66eb4ca18e35e73a41619b8d9ac165331cab7bcc0686df4dbcd4f0a0a3eca1abb9c
zec6ecc0ff34b6eff2afc44c601e858b172ed58c685a79dd1c94bfbdc3ff460ab9d607788df317e
z1cfc0a42df0f9272d3dd73b60a696cc41344e6354747fe0d8ec081ce7d8ab49301efb334cb7e85
zffc6f4c094257eee830a2e354833b34e4e8b658ce1c996fa5eef0495b109da7e72bcdc2b428eaf
zfbd412741475bc2004c56d559d345106b9524a05928b83609985d576e3fb8dda5d14fa30c586c7
z4a2d1f67264765c9e264ea1c065f9f875891860d60cc7ae6f2f34239a74246ad47b2e77adb819a
z5e5c569d5f893f22fe2090f8c7b64aa1438fbc51ac7464f6ebd86e7c38d054d21c0146d89b1b31
z6624805e2f5b54ecc3a127973fee7cb9f167db7e03eed0ddc4bb0e7c8ecfea873452e70fe39534
z9874bdf031df01f7764a3bbcc1a4247b0405d7ace4febc18b2f12c279a5e2597b11d4001cbc745
zd8b4e528b856dbdd5dbfbd3292a3b56127fecec85519a4faac15c3b94f201537d9f76daa9ecd22
z957a85ee53c86350a474b36532081d2d099436bb3c347d36fd80df62b3f0882683d53a01b30b9f
z68d8f383a70f011a8cc2b48b9244a069227ee0e42da7f7d8c71227de8a69e9fc79fdfa3b925329
z9a75fd8cb26fb69bd60c882b212ff6d14c1e664dcdfb38b29bf16bd623e786867d63ce816fb79c
zdd8f88efab01f2397f93fe813de93cc684af7f49fbc36104d817fbfa7ea23a9ff6bdb3377b985d
z98ad4799b0b943efdf1b84ca8b24ad170a09fa2fcf705df4020a487deb88cb28333088f4f590e8
zebd9979da5b2ce50bc041b994652dee0b3ddd66e9ca82c91b8872779d18349b51b5bf9260c8a63
z19ed26b4fd7f77c6fc91f7c0c8944ef3432768f02dc9c5c7ffa231118205c730fa9de02085e1ae
zd8b738c27ae56c2184dc9c3fa3793b26fc12bb2f0667ca53a542254adfd83be31ea08a1328af0e
z06f1ee36bac500a2bac75c8aab079986a0b2a4207de4f3dba5fe7b3b266d6442cfa796e3edec2b
zf3c9c038fd1a51cbde5fe6ce2b65dde58d6aa1079b25942c0efd82088ead3f1f0119fd49f5e2a9
z230f7c2cd5ce67a26596bcb9cf825c2fae1102ab3fa60006104fc551ffbf0a6a0b456d08dab886
zcbf1e65fd0ae6b40e5efbfbc6e23e96dd3f2fc8666345dd2e712a9945796fa57b24ac8272037a0
z919fc07dae131b40c24620218ff207854f84470e06adfae732fde440c3b3f2c9a13d26ee2608d3
z73f8cc14f8d42070af8122bd75b8864c0b4dfd04f29ade91869b1a030edbbd4e07ea62cf2c6d1a
zfe539581e900d7e7bf1ace21d2052fa79aec9ec1343fdfcc614ada56dfe511b34ab588df9fde91
z692e11d333b037a0cb8848fd4ce8aac10ee2c69e23d11e4d49c95bbf029654419da32f349d760d
zf67bd82ff49658d74f9b36a595fba4992cf9fc5605b5d203074e90f0f0f9da6bad64039066939d
z24f93684c2b6a04f054f06911ca55e5853aba5df5fea630dfa52eeea6d4ee7cb78b23becfdf460
z0d719cbd5bde6297f083667cf21bbb159990ff349ce0f5f892c5832f8930dd3ce733c8d335d679
za3be1a757b0d0a610d0efdde01b14b5ddab216cb4c1e8b2732b59ec10de5a0f2fc58d119377984
zbbddb1c1f4aa8b7fe62b29aaf599a30ed486c8726fe513120bc140f343a93540f12df6048fd61a
z23c0af9350ac8d64778cd5ff581993e5789226f5a22889632c27af6b531b8d22dabb14b7384450
zb92a459afc766cde4f0312846694cb6d0b7b93e0b802b5fe4894b9dbd07600a21fd9cff4755d1f
z3535f6366942c26d5fa4c6793606ea2c7cfe7a863f4f47b82e12f7608cc33d78c3293d34fc01d7
z12565c6425431e5080832832ffbcce48cad121c81d01d8b4ca535800d9abdb63e7a2b2083d9867
z0b76b821051246d64a6c416ea62f364333c0e1255f9c0146e93fbaf4c2c32d7566a5efbc723501
z6fb2c197bd2a04d9eed9a4e2dee5cd46d71bb20450ac346fdb92a29a3e24a7f3e989c9db2d6907
z135d809a26d115ebdaf3dc6875924aae36a105c8dc1262b0474453bdcdcfdb896c93b18fa871eb
z5ff8c29789c7d862a68a9b97480532435425e81d4e0e10285b80d637701fb61fea1c92fdb5ce5b
z5583121d6b10e0dd4b7083395ef849e7df4b37986c87199822307a57bfc6b955004dc9978cdb77
z27894df06d6a817d3a3f25528a667aeb4cfd4ede6a1f1b4a3a45916979ca0709900f6e8554cdde
z87cf6b7cac6aa246a28bfd9b46390d44996db64a3df284f66a454171636149ace22e0e242c6bcd
z12c32cba807c4cf4f42d674230d5135af64a1d728fb082a4b79d53a0b84aa56385f91b3ecbf851
z787ba6256eaa0583d3b7f2da4b9af4351b084632fb42eebc06636f3e955f6a43591f6796defc50
z152a56ae66fa41e2359c47e571323155054be0f702122f09a160b931ffda7d5fca1fa9ff136aa3
z2fbc1172b316b164384c87d3f885327f208ec8cbd0e4ad3378d3a87afd91494defba19931438c6
z16cc70e997b4f11db5161c7af0ee3867c82535257a228b8bf10100ebed5dc2465eac83ea1819e8
z4866b73aa6399d30eb9020597259ae0a7857e65b832bfb1cb9bdbf8b2207fa608ca1530e87c5db
z5d8559b368877647c572c751319ed92c70da6a58fe9aecbf38c02f8382bca596a61e9cf236a3b3
ze4ae66738c07f18030add19954980538bfbcf02311d9d44d94c953b66e9eeac083d5ce70faa9b2
z9b5b2bcf5b25eaffe1b946e3177cccd35509a689c3c9179dd02a115e454add9ad2d67b946e7b73
z5fa5be0f01f0d92eb67632210ba95cdab9316f3f46918a34cd59e4ab43af9b184d400c5e13c5c0
z735688e14f7d1357e63c65c6666f8e7cc13d7ee7dbd87628ee65ad59527650b925ba177a82184e
zd9a2c430e9cf912be6e3cb9734029d792d66977518df67af2f8033f9f7df6ed87c91eeb122ad04
z7760be438c153a40516923afc622130939e6eb1790cd71bafd131f357106af851fd273248411dd
z8d7b194368c28ec93c968a18773627a969182fc899c278d5c25623f946c7172992ea22dc58d84f
zbeac0a6ab990d5bbdf98a8e8f19f9e3e492fcb12592f216c47e8112eaaafdd456efebc6b3284ce
z89d55df73356bd9242f9e9732a53fac94cd0a9c5365ae58e2823965525318e27913f755acae323
z08ebe6163734daf07c10731a1e13015f7f21e5dd3a114c7bf772dc6c3e653d8c5ce4c451d22889
z9ddf9ba7d638137a558577e1bf3b6394e4d131103993deb0fca3d5d53c973f5ab5530edbed670f
z447d84288e182519eaa5f4c057057ee91a48397dd15971b748d84efa02e2a8399e067692ff5b6f
z9284d9b8b0bee790700346a251b1d7d6b3ddf169f95d90e0867cd28dcc301b13c2b7321123fc77
zf1cff60fd2adabc7c382d886886ccc7c75207290cf20f3b7d4706ddbcef62db0cee66ab55f1db7
zaeaca93233fb684e781294e46ad2802faac12476af40055fe752398e7ea6f29040ee543088f926
zb7728ad2ee38449ad4f7e2ed5242eac610b8ae5c1cc3243ecb5dd8bed022724007f2e932079b16
z8dcf4b5f67e762069b526aac04be9e78b93bad8a2d551c85180218dbb62fdc1962f077e5cb29d6
z2622a52d0650b179ad653e15cf0fa543aa8785ad032f1abb4114e7f5b78686b9ba094dab2035c3
z1690d4f8058a06b3dd5b6a5267e8adeeb7c236dc2cb820ce54a06d616686a4cd31b806d431d9a4
z7414fc86e443ec5e3caeb401fb7b31c6a475e9b8e75665c0196d6db831a07528f2d3990916dc4d
z1f0a60c3e4b04f705da0e814e805fedb626e163d74e9d64108860d07ab10f595dd06025160e107
z211d765a15c373cdf28b8a66e5f4e205c8f33dd03cf4c49d4dcb72f15b97a89b6bb3773a9b612a
zb8f16c3cb5e147024a7b1f86831098873bb09cea929770719551d6a1a01584da2bc1bf5209d053
zf8de521e01133772e911e8496ab80c15e7d686a4c10fccd82107253dad5e258be50d90ea23c16e
zb1357b80fb78f3e4e2afaff8dee80cb8aa37c584aea8f7ff6cd2b38f9dc3cb485ef251b1832f9a
zfec82e6efab833acc379a5a436a570856d7318241142bbf75e0b197490e0c0d6ebb228c517fd38
zba48c45f44718b9b65a4dd8024db71f64da90a76dddc8def036819a5a4feed3d52727100b84dae
z8dbfc89d3922f770b459a0f5b251d88b8d81e7c12ab2bda3f8b0fd674676631ecd440fecf978c0
z637705c7aef4c2905d19a5743a0681986dbe1ea39e9ab31bffd2fdf34873b4ca51e24ffc71697a
z6038eca336cd80ff767dddaa243cadb6c72fedb10c380fc93506a432c15537f4451d76d62b6f17
z5fcbb2cdd181782d17b9a3aaa45f02ff27b732e999065519162033c4143bf292730b0d5ef4b4f8
z710aba9cf1daa0c22e305317420e9397c117191356408f85697f245d0eb84519d06310fb3d5a28
zbd8a750961d1f1c6e82d33a226b7d3da674e272745ec78eaadbaddbcb0bd13a864dba004371a17
z959c7c06832d38bc3e07973be2b0cd6314f151866917e369dbfaf6ba49fc79fd5f6c2aa7a459a7
zde2c3a3eae747743b55ff32fdbbe0e83bf9e16f3d877494dc7389a5dacfa3822e5ba8e1cec97e9
z4720aa00b7aded1823bead333c8bddd08a281dc5fc2a552fe29a1e10a53a77c9de83ffc33442d3
z6ea8faf39e8d58969be8864479bcb2f32f0462b5abef0c9896200d88e060166bb3dc576fdfe91e
zb1f9f2d31883e3bcad89ea32ce1b79b36c76e0741658c1b9dfdb749c003eace0273de3a4fd9856
z71d9029db15b611101583809ae937c5324fe94bf486f7fddf3a6738e1ee87b47621a93be236f20
z0f1b612e43ee8a13002f0e66bb3ea4dcf20e466fadf588c0204a981b3a2230066b0cfed2b940d9
zb441a3dec2c500999ff7a6a7c379c584b97b80ceb0c023945145162a04bb74793b2caa09ebf633
za337de753e5f41bbccfeab76c883b83fd1e26100baf387e1efe4e03ebd91fe83fee8151647a692
zc4d7f2da411913e1a679fe61a03cfdc45e2f45b29110b770c9472251a9821cbe3ab7d61adc132d
za54b30cc7b6573df760269f93cc7b5e2decdf5a1a6415506ba2cd7d552b666f760b58ead99b8bd
z1f9422d784cf9510890b76283fa79c50cea07c056b79fc17a82a7aa0c8f9e307664a118502b159
z9201039717a09a626d68c335bee72c74f74352378594b0ad5a9efd2157c6e61c35c661a53cb0f1
z0f73c56388436581e6bcb61b12ed6704876e255c019bee7a6f6a1356fc3790991e525f720082b4
z81019d886ada3708284b9464efc15af081043fc483a6ada78f9a97eeacbd4c048ae758bb914161
ze1479fa7514ccead3d033189694b60559454e814f7ae9b64a0f704b9dade4808f33493c12b507b
zeb0da7cbdbcf68e4ec4654c0de11d156ff508e7c5de0515a3a77fd8570057f8a15607b3a9b2bc0
zce0f4daf472fecb21d1dc0b93fda386b80c1cdddd51b12b190c4e2a5b682462d3701607792aa30
za9efffe63e2cf7e87d2064836807edb06e43ded5d5b80a18501348f2b7625917da06fac7654449
z51f59c3bfdcaf9cfdbb7a43c5118c8a4245b3f0856f28911f3dce44bf7b38360c5833723042477
z5969e89ccd3ea9e85b1225a5b0e569e386a14ec5a3b53e0f9918de734cfa8fe4f9df4402947f5b
zfb713cca1118a5c792a39611efc52dbb6b4f72ee1a94df4d113f0f9bdfa32069fee80d7a811839
z8023e3363534e1ad8bb35a49ab58d87a26845cdf7957f46d61e5926ba6e23915b73c7c92bcb11d
z413747e6f8b78507315f4ab5e606cd7a27ff2798b605bae68d267cf38da36242d30b9a98751471
z52369a0ec5c289c4e0d292449d2a3852efe299cbf20e1aeceeb1f6c7debf35898285e63235b530
za64bd14266d0bd4be60c08d28db5fe92ee6c3707b70eb967c313327c6c72dbee46f366b37d5c33
za42b45d83dfecaeb82d8817cd35acb7f803f3a3486214a41b94f53f6b8a30b35cb695d4929a535
z50242f1e267ffd371810108765833556932af5d2c273bf5c13756695bf37113414a3c8c232c8d6
zb4a65ccfb4cc9e88b9d1801a0310ef8a5514aef32b2f18457e7c091608d5ab212db0722387866f
z0c8095eb23e836f95fe7e54c454e374054eacb0d240683c82e3618200acd31e2ea10da91796501
zaebba4e6dc13bf962f0ddc328e34894cfffffe5b00b6af95f749d78e65058953ff2879294c076c
zed4d58411f73e606d4687e23de0742be840c1254b7cb325846927ff9a4b477270071b2aec8a57d
zf69ffb6b899914a1ebddd8263e16dcafd9581fc040d7fe520af76d664f2c5508466dd17966d347
z1b7ee0dcea25c88015b99e8d84536738330ecfa3efe58173ff9cf68546989e457fef25e862a02f
z5d818ee3c2229912d98d12892d250036043be306592deeea65b7e50b756533a91d57606a89f711
zcad0365948a1752d7f3c2f0ef1ec250949fc2b003c168b87d2787b684f985226d428c32039b9b5
z66dd0fc7751746a750ac04bd9cd64963a139f8d3834d2ab81431f8c09637408b783a5b3f8209ea
zcd9327c83c1663251446503f5b0e41c2297b7a830e8195a8c1631e014064415949ca4ae1a804f7
z305cc3005ef91abc6f4b5f1318de9a9654593b64164c255bd28c1e16857cb56b39190ffe2be504
zc42eed43a2712d4582cef9d7aeff70e4b4ac59043e9f44219f16d985f1385345292ea445ab8bdb
zc78aec3385c08f231fe0c96320b51eb686bfb0adaf36b4e9334cd8bd02aae2518a192906cd8e81
z5938933323b3d082f564529c005f24bd33c17523fec331ea0004347e8553019fdf7afe58e83763
z338fcc86a0c51ea5f34cf4a1d50d5d34583c38f9706b3e1acd3cc919227665b670ebc33bc99ab9
zd773303a77adee6513944bcfcf1ee36435534e246bbb18effc39d2df5077fb50f197420483bd7e
z451fbb7cda533302adffeeff539d9e7b8e229c96be16dd98fd89973cea75d0322308d5c48570db
z9bc09216bfdff1e239cec4aafeda49bc6f456342d9fc4544fbf1c38259123ae3aa594b8f01ce2f
zaed9d63b6646e71671de92fdacc8434aaf8444ee014e0f213fa72a7feb4ebf5367263a0af799c1
za1015912d13d680c96e2e6c69383994b4578fda5aa96e46471735a8b566be281347af32f0515a9
z10e11fe9b5a538f4f44d2e9e86812850c6173e1521fac6434d6a434209914630571f466fbd5278
z5a7ffd212326f01f1a7a8946014dbb19b7d85befcf0cc3c51820362ffd5e86c18c8b61d1004e10
z2d07f41b901c4c8e8a5605f747de77d28c10967d0f05407b96a9b9a68220176199d336e0cb3976
z8ee13847ef21b8743f7850ca434b460bc59cfb4fdd3ee96ee38ce45953c83a35185b1ac32b5234
za93bff56ccbfd6b5ca0fad29dab1e74f6ef7d18231cfdaa56786d6013aa5a69331a209c9f13b0b
z2aa921e41f62bddfa3c23899eb1eb2e97268d561c59a97ea1cfff3cb6c09025a682c40e3a32c42
z0bff4892911147f7fe811db8ceb611fdce5bb556235f7ca34b248d60e2ffcfbc149868028b704e
z24eda86e1fec5df783e6a8ae2db54ffb59a5ae46e3a6229295f5edf9e359af83dcf45d7ec3ab16
z01bede7ecdb4e8d4f39dce0413d9e03ff483cc550e5fa68ceaaf915653afb01b02e0cc0dff6e66
z1d5f81100fb6f48b59e9c55b57a0195a9651f8927d4a1f4f7ae64a10da6069c761a6eb3720a7e1
z11860fe50763f81e25e9c68d8b9089a1dd9df85df7aca9d50c8a326680fa2bf2891c247e570414
zcc08d468a3259db9b945dff42e6b048ea25ffbf0a69e22296adaf3ea5bf90f4b39eede4fc600bf
zef5cafc14f9bbbd683daeecc728f56d1b9a02589a491656f6ed3c41c3fd3694b498b6fa1fbc59d
z4e80e4a6ecd5f83c359320ff9e8533d5da26437707a1e716efd60971a0739cd8caa5359458ea79
zad8652e8ab92c61bec578c5a1f02ac656fcdf7d4320076d47cfae670a7592c0e1b4fbadc405653
z6522cb6567cf1d5f54d463663beafe3a49cdd304b399e54b0240bd7beb9551bb746d08a22be858
z6acdeea7b1285cc80f38cfa77ce00598bfaf5b7dda6295fcc8169a91da378f3c91ae53b5f0daca
z841ab730981c2df9a01c2e00ef531297aa1137ae3bf70fd215f297f646c614974cddd9f3ceb91a
zd436fe1814c2aa2d0de08800b4465d6cec27e1bfbb3ddc9c4302730f0c05f5b4b46124820cbbf7
z3f2ee09f9d1f00e0f44c1fae972c7ca8f2910b483da284c83c2295f3ff6216ea2adb64152263d7
zf722462322b61b8c1447f5c8f96c96cf0e36828279a5c335cb2612647229823b4ed32a309ae18c
zbad756b503fb1d6b1c3d67278029a758da23da1231bef83c6015c7efdcbb66462b96f280d08c00
z75c4d52d615ecc530b5d186cfc160db1db747a2567e050acdc95aba91196da4399453df5fdaa86
z4f553d0d5ae038b0c2a38e831b4e105758a8ccf7df6edcc434164ce2e696089390308e09a8d8ca
z88a50c63ca25251de90a183d11cf46ff59d3eff9a5db8ff8256f97bfc90bdfccdbc02edf7ab746
zb9b2207a5aea8c79629752ac7af9dc9e824028f7b6c56ca72f01064ded1f80218f213288541226
z5147b0fa448fc807627538390260f5ca976ee296da4da05b9c6d900b13681bd0d4468e8257af90
z42d71cf6a4d633d03a039c70282620a14cd7018627f3a8356c94dc15de173e48496242c8c456e5
zb45e152f3db2ff428ef79228b4f3adf6110259e18cc677466d99f09fa67a55a9921aee4c1eab97
z36c9735c49b488694edbd9c90d4a7d6bcfce8e0aa3074c82380c3a1fdc55e0717de31af5a5bbb2
zaecd51c9a682221d2693830f3be7e8da2916e83822ed0e0175340f68161c783906ad645bafc97a
ze73cff1105b5985906a4a306c2971132f50df5777287786ed2bd132e936d66e89b4cfc92f1db22
zd71fe8ac4478c2c06f735fd19376b5d47c52d548b7ee06b4e97c98ec0054f3bd48c5405b6fde8e
z2c5e4cefe95e41741054f1c15056b4c3bc9e3a3a8e7f38c924e3a36dec538785f474536fc32fec
z599047a468d986bec4b4b19aee0e241ac936a7a13602776b40a705a2b1b71df87bbdc20e73a57d
z6310dfb169b17e8450ab5503f0d0cd65297c5cb0216310ee66d639fa0541040c58aaf0fcce7ff4
z524b3d8e10b5ac0a6056d13916117ea070a56f1e568e84c1930cf6374d34173b33a683fdde933b
z4d5a9dc4f6e52e98fec74c084d4bb18bf7a7897bf5508f7fadcbce8fe3382cb038f62230db9699
z450b3620d086bfa4d7d9acd87907d841ac43376dd458a1f68fdee349e0263dbf526c1fa6ad2d4d
z9392183937cc52c636529e108433be76dc70ae777470a071e22f3f0700d5448409d9e3a86a24fa
z339f51c3c850e2e29c089ad194baa6600e31e12a01b23ca1480314ad875a1994885b3c9392879d
z92a7339cd04392d3d3641f747613d7525184250d30864edbbe0fa63305a487c2377ef1747634b4
z2bbc644c63705ae589bfb364a4366edbe3dfb421f82254adb8cf4d2e2f4f3eb87e881579303e27
z7204e895cbe59528f08459df59e7f6828a9bf361c135fa5b0c232a334df80ac03565bb3c9dd0b6
za3712c09649486054f484e0fddd58fe5f41b0e0cf51788edbb8c236e1a5e93fd7df379264e28d9
z313a4d2de09b242d4ea73942f0db9b7733fd0a92bce6b83e517f453c4f90bd786d4f52dd8518c7
z6b085f5933e5313c2a413ced4f3f9b0782aee6235ccd4b5762d28ce7a58289b10e23523aef838c
z38c4ab1140bb0d182f8ec64fe81a1903c999bcb5c2fbe9915c9d91f1f508d200ffd810a12ff2c7
zba99db493809928b171fdf2467f2da2f2983a63075d743423a5fab5486e8a4883090feb7715891
zf39230a311d6fb196d37ecb63861d05928548f280f37a59f75ad1148ff84cecf65640376b71adf
z6e999a862e92cb8070223f7c641c69f058f20430ed54b1aa4c5ebe15f3c1eea99aa4ed77330718
zff0842918ec984389e8d942d6ee2c0de17e4b8e85b64edcea6cf594228c8a416ef7e30ea0bd4f0
zfe68434ecfb3b1b0e8988e51aebbafa0e21a5c79ac406baf93c9e45545c48f1ee73bc94cee6bfe
za6195b8672938351b843ca817fff25e55dbcf0d10e0f835843bdcd4df8b3ef6bcfab1c5f7c8d76
z940c96113e380e8d9784d88c48c5ab8a30731d40d152d7c1a34deb69c893dbca929d07837a1340
zb838859a8655d7e84d1a238c62373304fc677074a0f305d83998bb70331714f5a8fa3501626f08
z0564154940ec266adf63a54c8bc15b63498ed7b84e20441ff61498a6ed778c7ee7135b35ea5917
zc3f9c1605610f62a7d95e9aca40cd7773a0c016ea086d80fcd6774d4247245a93b0b8b9c2a3744
z7f9e828d47ca7e8db18e3890db3146291f797d83259267c585c31b8dd8fd36d962fb008bc82eb7
z05562ee8a651abb349b558c3baa53d4fdfb0f54704b52d7c38a3b8e10ceabb2d238077cd7ba5b2
zc1c510c63d2de1c820b3998b589d9fc1165a109df27d101623c695bf4204c853ec362c4bd1da78
z270f1a887b74e1d50f8af61ea4534571449a9a8cdc00aed141f75d3682d0912448460e1ff5cae2
z66896514e2190e5f1f01fba97d6733f1eea425a8545857fd42edf2f9ddfe102634de03433ba408
z1f5c48de6cab5546d076dd6dccee4197ad3b3f67e5fe72ece1dedc5f9d01b9844f79f99cc13595
zdab39016dadca5a000b26312362791841a65d30b9fb8d887efc1ea08ede248d991da77452c8ff8
z6dee0de880324b404ad43d8f666fa889442607af063dd0732290c99c1cc914a87bdcb724842f35
z44ea714ce95b255fa2c330048f23d4eef3e8ccc23c9db75074100e651fb0bd1876bc59d4645101
z7d2680ba3a9cfde1c088f74dc6a8ee057478cd43ece4c358dd6090eb7fe763b78faf4768500cb8
z414aa44645376ce578e4cf594ef905750440d9bb8f6af117b3a85e8611c24860532d417377a245
zb3ebdac2ebbbcdd676f78c906d7f25089a5f1e77217a3b4a65e88840bbb2faa6d7f9bcc34cb175
z0aa23008d125a664979aa969809028b3dcd2de83e27fa389bb74a0dd60c3a5419d75bf9571d5f6
z37f528e3117477865452acf9507e0451991202aab60b8d2d637043e7d1e590e87d63a8079bf301
zb9d2a2f59663ed63ce708a68b994f094b4834519fa0814d230836deebbc95d40e73c8a82728d5b
z70283afdef27fb74bc713e091a9ff5d7c6eab5d1cd975e16d77e6fe28c1abfac1e2cf97e7150e0
z23855c6d04b1f983e4e68f75b19d353905821f29907ce23f14c1341b71314e67d2f1f8a51a2e4a
z12a113985c656397a84b9bce898552b6f1269a4a24cec94aea609804c783380c35acde3177ea6b
z38c69ef03e10909e3c1c4eddfbd5e532d66cec369f36ff55a23942b428d861b7a438e44e2820a9
z27ece3fbaaf233a4ebda7df0f63b5b720dd75b91b9c6c4d66f31a0fb8c99d1b0a2300d1f845ff1
z30e8ebb5a575422daf25c98d10a5caafb53de0cb0a2ddd91550eb6871b70cf079c4161bdecf4b5
za16d5d2780cba58ab065e2694e21f3a80ed7bb0a63fdb86b9214ba170753ec3e19869a3da50007
zfd78132ee47c882730f9ef04fe59f791c3e32790795f3e928374bd36b13557d0607a3f2effba13
z34fa9901b2dfea4a805b53c3cf5acb31ac4bb8916b544c651f88fcf98aadd71868709a880b57b6
zd3ef590f1012be3a6afd3fe92b1d78f25a20dd621f10501861b7ed8b891e4588a88d352d21e127
z7593a653c70782b580bdc44a01aa8ae4c8f18dbe1bcb84fdee895c31c086c9924fc9e7dae6ce20
z8d38a842cc6ccfbdcfa360a842322f4eb9a5b2cdf09d550532349d74f0a7e88dc75fa470ae2940
z8c197267877ed7ce98e1abb516a06afe6e34f87f7f53c729f484360f0c1ed0cd7720e7cb4b6234
zcc2e196dd37da0241603ab214af2ce8d425e02ee162543e8e836e4a9bf2947ecedb8ae2f1a07af
z36ff243bd422bc10fe4c8d2f794ba6770afbe6acbe1fe1682eda8651b280483ee23108a1d41ffe
zd3aedf96a9236cdbe0abcc8cc2b0cdb1d9bfa01b9f57b8221d7d6a6f7c934a1b941c475786e594
z0ac8dedf117a172352d04eca4d0a81eac5a152795c0a2cf0334aef86cb8d32f1ad91e49837cf70
z7837a7c48d3fad1731f5c98d1098e6376b91b6bc877fc7b65e12c764c9d0d2af9aca3bab197d9d
zfb749e8aded07fa44ee5b9d6e37f9e7f1c545af294abb17bbd6bfa890b59353a9f6ff77f51fe79
za749da1bd9a2122623adb54b9193feefe2531503d6b2404f1140ae8db174749e9ce3888ab075f7
z03c37792dffb31e40d082f7cb8d3760bc09cef09a054b04ce65173f1f91e0f17b2f72707077a90
z443ecae4f10118cbb573d4fe569461f81059472c2190d9ddf83a2f5cae06c613fb3f2b81ea1219
z3e75fc034c0b3458aad0ffccede5b0947c8f19678562e9c7cd21e97e48445da1867cec0d452c32
z5ff17f2ef8c118844a6a327794d21703f6038d7b4bf91f0480ba2f3a9cdbda10acdcc0dd123815
zf9fcc8e5be72fe385e9c22f1534ccef8425c98d1c9fb756e382675fc03c62f5cbc5914056acb00
z1c9de09aecffb3bf5c489153e53d9500301ad92d63856e2b899133c615d1f5c86d7b3262bda7bd
z2f704a87841d58cf2b24605c957b5d39414abd2408bcd55d7b3d4a73d729ba3dc3c1ae2faf7349
zd272848098f40c731863b51bf380932b61690a63601223f0fd18667a7f257f5caf529d0a321e56
zc84f62564deb36b9cdd2cc73c28b44842ffd054c757904a3b63284e44e9d21253b889795c9a657
z9797eae63e7ae81077451abd02bebc15215f247bfa01c43a368427bc6b0b36790f26401ab62cab
z19b92066a0f1f7b776cb5eaa57949315ece7cf6d4a73d0453e0b72893d14c891f4d3e7d4f6fabb
z70f55d0319a6963d6f119ba372c2e6ff7c7a364bcb7e3592260c0354940ed75865147da4757efd
z6caf5d0283558865e71df65e2fcab168f12ccf5ce07b2b53a86b112a9d0b63b898164be50f5440
z93aaacefca519cdccdbe826b2d1f1660d8635faa18907cf6a154080b23ec2f02a34b7818d022ad
zaa1bcaa4067b67a985bf11ad5186f1d932eb18ab38a2a8415b03825ad79896b699f26b50f28b56
zd4c7698d0751efa9d5d26a75bc4d3074c56f5c43b2928e6005615253e561f78c24e725c400b2b5
zf423d0068081b78016e7afd113417f43e2f46a1bc6d6827be1e23fa7751a6aa730144748c8be3c
za3f47596b2795c30b8321449cd29e8b916e5cf0ccc94875781076ba1d64e816a9fe577fce60acb
z6a575c6e253dc7312e0a5b4f2be6d76892d70a2efa40c98550f7a2f5c7cbd048fa3174254d3430
z0343dd37f097599115ae066fb01ec45b2b722df8f6e59832934424287c9316f9a3c49fd1675adf
za40e4e3d12a9626afbf404380cf8af2bc340b5916cae3c9ac6ec90e75ebc9985d4c08192731273
z8f5b793a0b9be9c5fc9b96eb98e00eb00cf673d8240fcb4beedb9541bd7b1ab2210ec87ba1e7fa
z3d3e0a6f41a3d5ae22d99c7dfc118b28642984984f9c2e966aa90525aaaeac6fa7f02df1f1ff64
za965490b63e0cf0cd707536f470d04f8fbc819aa6f8d6e56281e676b764bf71051d81d6eafbca4
zc2416b9b3f7afb94f712e80642e02be428a54da258b1a943fe3139170ab614ceea7cc67703311c
z9acb0c7852c715acad72d8617e1a22164063ac1a49122c5d3aa3d0ec60f99cee8fd20bdf100c47
z84f3f1d9194f320d1b7d636f7d70f792fe704461585144ecef98c2aa90e506df25d88855610573
zbc449de03e3960873bfbe644d2aa4e1d62bf8d06176048e5f57b176e9306d393b422058940406a
z58db0b62ed60ce61ccc2b3ccc068ebeffc845869696d3d52c5c1f3bd5c7a0e251efd0c02833291
z995f107ce70d6569dcbbdf3477f99edae23896923539c9a29fc1f1d4e7e1a704d53ecbd0076748
z0bc9509442bf7457b763a5241f4391a42a9fce14261357b4e0aa0f12769c33d7ac8dd7e33657e7
z8d04ed40f9f5a832c4a55db3f7ff6a9120536c547b486ad98be233ad477c506d8fca23b21b20bf
z2d7345c7c05d304889c509f82593be6ef83397f01f1e3d8c471cb582924e890d305b4b845dc9f4
z208d155a68d770fa5c8f242401348a010b7147e148ad7d64c97d3c1751f4e05945db2ba886e4b6
z9fbd916fa4802f81e6f962013ce5fa95560cef6203f4d32e1a9688abde1bf1a71e6c28f0b59e26
z1703fc75d9b02d5586acf3c55643d87dba0f703984acbffd25eee45c4669dcb2afa31c880f4c67
z288b1f367d646acb7bdfd6036d3beeb9906c728ca143cf553db34c09ed1602d30e1b8cce579e83
zff3973e3ba23ad04d966fdfd5f9793aa62b3b75e9c3f0ee526218c91fc720046a2d6ffb586e035
z84bd19d426c3b3ff5242e7c895678c467f4a460db7922b3ee7b27832255140784c1072c084f6be
z810a05bd07d5abef8550cda710841fe3e10297d5f8d58ad85b95f36f8b59d7bdbdd068cf205f5d
zb6f909bab8372ea7cd0c8f0004813b9c97fe3c88bdaebfca63e681b72ee9fe0bcbc7fb222e4696
z0f5c29fe0f7cf2ea32582dc1fa0ffc9a446636e43159bd9e87f6b9fbbaaf0a5d11057cdada438d
za5058cb19cf68a4dd5a2bcdb278fd71fc7430ebf3b9986abc69401fdce44cc1f00d81e8fa36d5b
z50fe4adfeff853c2aca67711b64bbbe747d1450fbc3fc53cce291e9b1f5ba13058a9691a2080fe
z46a5d3e4925b3316867c6cc4dd636f7d647449850d56e4ee6665b8ffd83828e9ff7f6dd9b7bec9
z26878e62e8c9e549846abfe725a3f3d9a96686bd6d7dda744c322cc9c13886ceb247c39dd82119
z2109bbe5245f0f2b718a404674a4b23e3ead0f54c291fdacbd58cca028cfa1dfa624f350881327
z68d115fb0bc2e801a57090094dc44cfd0b74dbc406406ed78f27663ba0e723e66925cc4c5a6797
zedf34261dc03c5f56c8bc33fefa903fde4188df0ef8206c8dfb063539c84a9cb6f357fbb412307
zdd72760a005baddda604c7032dc9fd986b71cb48f967e6b2f3b4372d7d28a629771a4789f7cbd3
z0896433a00c90b72f1226d882d250a13d49edf2df128ac11e6230d6507646030c9f5c6c1e40186
z595be51cfaa91b64f4941fcce4524a0529e98ca87c5419d96ff0abbb3ff2cb7f31889b8adab65c
z2723e313d75c210ab45e79904a96cb99aa76a2356f506d2312055b9d969109883ebaad64766b4c
z94576afc2c4852c645d2021a74603e108ba4378b7c7da4cd10cbc07d66939fef68482512b267ee
z5e83489e7e8ad4a284214ef7aa9a2620220d9baabc73cabbe57b9cd60fc1c950f1e7105746bbb2
z7d3e7f796c84b696bb7a946e53000d96527fe57b020f4dcb8b417abd66111e081292a70970332b
zd38ae9e197f0276a95412c0caeca7e21602870f163b06a73520700ac557e8f0faac399598d7397
z38560bcb81d75d9d296e26d49ed7dfc4e63c95830d06cffd2b3bba2a2eca5cc4ef38cdc14fd26a
zf3c2bf600ec96de1fcf7eb59133493eabba27c2af8feab066ab641403fc3e95495efa0faee42e9
z218458b84480ba2e12d80c2e37f10901803b199eebeaee610ead726ec78b04619ddab2bc7c145b
z930441e2ce2b9cffa99dd03e30e4deca32f1d4a3d7d2f8eb1afd65fc887b1d9db904e2aa1ef686
z9919507f6812d8812a3b6399f8df843f0044273bb33806886222ef13b9373e63bde34bfaa552ef
z641598d80fe5c3a951ba437e00a4d8bc9a7879db52139ccb72338aa80fa0a4580f37159b9df8d1
z5c33224560b2ece57f577bcebe8d0677b609215d35c0f5eefe5597e2a060410446f0e126a2660a
z060fdf24ac6aa245ed18c4dd966ec95255cd3cd36c189f1b6a5665a5ee13d47e1dc1a287a46a2e
z64b5d321ccf3666b70ba2382343cffe8bffd6b5f1599a8f2543c7e393e6fdaf9bb561e95dd1363
zf1db74fd79d5ce42bafd8d3039bf73af13df1631fee1143312410cec62d0faa128233a6dff4e7b
zd6e42d53ad9a82e82646ff308cf7858d337738d166a61dac5b4cc886fb627b2c4f28aa80934dd6
z2c667700518307737de926459c6e0b4a93430660cf2232d319238c64787880ee4c02ddd54d76c1
zbf1418f33ae391ffcc569465eb071d24c5c7e45cbd50b88ac750008074d9cc0b1af56c97a4da82
zac0415cfcc790afe921cd22e88dd3f4d63a26b204e892b47c486dd34f983342d8549b0c60d104d
z77658d9abf88a44c6d90cf810678799607484b4d3e91e5c01d81a5b1c0e253a2b19b0f5420502f
zcfb894847199b812a56d81ff1c5ad04b40342e3c814f64d0b64a04efdc08933b40b82e618ba75d
z9d80aa2f4d9bb85f880e2b92964c0d1c3269e6cee8986175f18b2d95cf04dbe0b31958fdfaaa7b
z272c3167ab006b89be3131a3b51577a4b0f648131f6ad186300d0cc610b22c8f54cc12a0cb2a98
za0256e7089285929e4336e3ca2eba937b052b6346e3940127f7c04f24a8b3c878c07c6eeaef7e7
zff49909d2183fdbd3966a7c2608bab973df79dd836a0f864889255ac58ebfe29246714b4ed0b44
z20f7f4424dbab2834d450fc4856f95d7c70388364aff12be36727f31ad29f41e9c912242a7f8d0
z9b64e22738c16889a2cd65f5446d9e286b99743e0f982523edd5f8fb036d14737ef453f7fb3c03
z229dc7c39180d99bdd52ca5ee94a3e289501097d597627eec413bb78b4839923d51c0a09e13e64
z9c012d3d7a64d1db7feedad3a1e6c6588b36e75f980df578089a1ff24a90d97319c8f6baa74405
zc0d80ceef205340b8f805cebeea828d068bcef92a47e9d45b579073a892284cc8009188d970ac9
z0f4c58e830818e06ecea650f5443c622b52e66b614ae4c3b1dd8e2a936368e8d0e590ac82226d0
z6db15c8e0c677bda57972b7e796da8369acd64cb74ae2fecc49c8b820d7e7904a8c84bba1d634b
zd6a5caba2dc6d23a39c3c2fba983a454e06c2fef36cf1ecf500b7ef6b24948808c7fd1060b56fe
zca9dea8d4a8c1f72d77e48f9362cbc0515d33c82a0e6a4ea3154e47f4992700912f5ff96abe11f
ze6c2c4fd75a669d88a483a5611c70a9eb3b73224200462058b1fece284ce00b538135cd9957608
z72caffa8b9eb8f7e394f77727cc538dc401ce3fd5a14ddcaab643885d6300294379805a71e6347
z52e7de5dcc93ac8bbf1d16c0c3c9e8f0a7d554c5607800a5271add604b7fe98ac03d90358a1ce4
z9ab7d934e29d8e1c0a3175657ca1270bd595a6956019d9524969a6bb6874afa4e57dd5ed8a5148
z4336068b0ac7d669c3b03649adfb309b5fca994e616ac4d71934fc578dedc6f346600b9e361a0f
z0a8567785202fc7f769aefbc5f161bf22c0ae620fff06a0bc501a12ec3572949b360c5a26ec017
z369b954d5cde39edd60a702dff61db146e5d8f5526166525b6e7d4893d0113e99cab1ec75853fa
z57b6b84800223a069aea986bdc735c2a27d8d3939bc9b58593a0b8d472de064c663419f94443d8
zc32c6e4cdc6fa056fd40140a9536b5479d00061623af653ca123f03bb9ba31e270b82bc6d8d2e3
z460d55e92118bfa8460c9c922e0c134ec535f9dbb954fac5958ef633f058fc3a29831881069c75
z5f7428367d38796179645e9d558d9e11014c14206eee71258d736ab687bd7657d0499546ab1852
z795da55a822f08ea01f45588f9638ff42581c98b7f20928338d4566e7cc635ed124164db29138a
z0fc4ed3beea94a33f9f22b0768e4dc90df9ae01a564e6b68ed84bcc31d108b8750375babbc641d
zd20a96f22201f6850443dca521d62762f3f3b70e0886bb99e91dc73fc0893d5c30847b88b35ee4
z09a1cd56a833db983c731cfb235714f70de44daadf5111f7a6dcc960859681490981ce1b1c524c
z0cbcaf2ace74cf20bbe51bea92d42804e67c660d87259a28209cf83c4e608470541a8b31f52382
z0a11315493052d9a34819877a15d20027d7d81f607e4cd1435f19ed6a2f15da21ede4bd9c28b17
z3d0f0452b0185bfe646f322a53903f80a3f74b9cd1024b2db9bfffb620bc904c7c2a3b2106f2ea
zc6358475ff4e5477bfb08b8a5e06e3f69431c1dc5d5a29a3987eaa76a891cb327db56e635f3502
z3107ba0fa9eb0b93d9860ecd30f237029e31d6c74443231a01b5b08d674969222ec713a7f40719
z630aefc5a432d6009e88f7701e23ba7ab707feb2cc6a4f98295002487210c11496d673408f0d0c
z37e1223cb3ca26ef1353a75931207f2b09c9a78410cd517b048f862e95b501960aeddd946a670c
z93f95ea05f9be8df859555959e1d25a8140f9ca683fdcf654ae8bf4d7bca8de645f5ff1137ab78
z31db9c3fdd7410b14de83137d8b35719e9153652bd69d2b5c03e72b4a21afeb44f9112ce9d7d45
z614206d8a696a7575779e349e5e59fb4d10dfa341021c794f3765f8d80dcaba68396d5dab013dc
z56c6ee82d7b61da21cb16b9bcf1cf668450b68eb2e388a951f1dbf47f90dc0596959407784c5ec
zdbce5289f109c4c8763f8c409676f4636e3051d5c6c6c88048c952bb7744b85b4694bc4d6be273
za24e87837d89992b31317b27e1a4e3e84def88f033ffb19f99cd41c5f35081b26eee3a776e6ec5
z8e9ea67c55e8c54863621cf541cea20f9bd72bdf0f535627b4df9776e2db7abc807fd62a6d0362
z84cbeb4d1383bd91ae9a017706d387aaa11da83aafd19ffd7d9a43ff2435d937b3b482a30d328f
z6933213390b4440b63d0539785434f4a8de62773e7b649e563f605ee32e3f6f86ae883433fd19b
zdf3ffdb1ffc48ea12622b50170465940fadf7f106b75aae1d1747264426406975f760a19c7ee97
z1a11df4395dcd647def098f7f78f0b83dcd6360e55f02cc33a1e50466eae076d496fbfc8fcf32b
za1697b05a7c1a98cf3093f714b1b425604182aea37d0a8392b3a20fe20b757a13f3e23bef35bf1
zb91994dcd5d5eab942b5ece395db991584c5ce04394201be6d4439eb3f3472a3aec6bf69e03044
z123d58d09383db2d1c8e32281a627f6dda0e16e2e74db85e747cf3987b57f0f5285e140470bd6c
z5b682473bbff35678412a2acf26f0620a5293af24cc776d51205291148784b3b89b76879ef230c
z65b469641b7edfe02f95e7b212d75fe6813716942646410442c3ac21649db5f60c337cc7f286c9
z8d565cdbf5dd7e9ba3848711ec823b293286c0dffd0fe0cf9dcea42cf6276c00e2f1dc67bc8d04
zb504077af260e9c74193f8440b2a8075d4452c02db0bc6e447e7652a8096331f0f6def0520f1fa
zf93d2e12116ad32bc671eeec1293ef20ae03c0f9f67b8b725519adbdf7f612b69335bb305b7b69
zb23bba4ffaeffbae96f69cbbf4fe3529dd091ea2c6b81bc00dd9eae1f3ddf7a477ee5f6cda6c55
zae958377bfce713dc1a8b7ac28565e5ea6f140e2bcae13bdc5a0585a25ad0149c6bfeb05a5a84d
zc5598aca94b298af86455edc17fab20fe1da931459e488086cb94ca89260b0d3177b44526625d3
z81b70d48ef21a0e312c89153e2588f5f5a5f5f867567d31fb5929e80eb27ca70bf2b75e9489cc8
z02133f365d3541052b7cdaf72536303c61e8b83e75c1d94871bf5cef07c7e02fc3fb1f24b2e529
zcab256e6f953629bb3954b40fae372ebca97d117e0ac986e90cbb94be61a24baa1426e57ed671a
z886ab19d5537ae54ae4ede990a7dde4cb22ab16bf18beeac18c15dbdca4531a5ad7f49899a198c
zed69d0d7362d0459804c23061412be1d1b60302f1d33858bd05fcb0ba7c074411480b9ddbff628
z1d4ed0adf096840c9b935e0fc2053d7d9f39e61b00ac13701f7cab8eccfa4c8d3b890e13ffd6e8
z3f2ae41c94c6f1f483bed3b4cf05f6b328037a09a2f568a13e5fdf8a1bef3572dc4399c939c610
zd4424a2e4e187097e97d8aa94b91086267dce946ab20a227238a571a872ff8573dd5802dba6421
z9d1ebf1c4589e37726c17f6a1db4b59a09c80773c66672a365f0b86f7c09136afcc22c5b88f50f
z4186f9cc01fd28accf54dd5202bb8bc022a514acbfe59360b3e887b3e31c1d5904f8feddef322c
z42148569d1133167cef8fa10fd97ee203f3fcc55fd650894b0b61b8521875ee5e3edbbda15b6a4
z0a61f5dd6720e77a17ba63de07187d0acd0bbad9c2815cdf8928194fbd7c2c0fbad68526e08aac
z7fbeb5c3ed7198b7c36ca85e0f71cefc7103fe677f24424e287da073ebdfcd060912f8048deb63
z2f2687b44317fde23de495cbf55b009e1dcf7360d54582f39edf41b18908d3c4263f9e14ceb7ad
z80576db17f936d5571250001afdc8ec7b40b2f3129f7435c3408df4c00cbe707f39ec86f4d292b
z8e836cd62908d3d8a008148f09459f7213cda65ce3237734f5fd06174b8260add3251bb3ed8b65
z72e9c47e915cf9d48cfc36736d86bdeec72ba4b1a75b7efa83a8a4e77f8dd983df1f162612de35
zae6acb6323f190d9178b5f7b17129fc39bf168d7f17ee5777c9c277beadd2f6dd8c69e7e2454e3
z4c20da8d521aa351c5ff835eefc0d650e2b6667820f148bfc4657f0a6d4513e07cafc0ead77218
z18a5701db67bf5bde89b86a82f537e395263cb214154172f161d2c6d84f41a3a4ce9d8f6906b9f
z05a695cb20217ca1f142890ca0153f98efee4e455bb5e65ee17dfd4c42969cb31cae276093b30b
z86148b7dfd4f6c924b674135f005bf41f7e4407a3c45551cb7a49b90525bc538246b379a366e12
z6c5d37f29c526519713dd0f0d857c33ed39f589c7458987f0e2dc04a1f63a7e3f5e72b507db038
zfe1a83a75615a2666ff8c6ae2ec48ea8ad4bff674d0c892e697feb5fb2b67523ea16979f1aed67
zffcbafbdbe9e53cdcdf72be14ce850d87b3256b81cb125a2d57bca23a43a2da4e503a0228b2f59
zc4feb2e29da9e8f249bd9e1de0502628594b8703f8a68dd9002460299d5609fb23db804f1036cc
z8b8d6faeba0624f981782f902eaad5e89978766a94868f18a6c71e50e55dda50f532e2ddac0aa6
zd613f12bb87537075c893cbf522da8276d8aec540333a638d61f59063e615d6b93599763698e6c
z86f14694358595190f9e13d91e1baeebbc6283bae80eaf3f3f9590bf7fcb4a479ecb87f287cc0f
zc94cf7bd6ec58a05e36e2ca7a338e3e051fcdfd6b3e1043a7d132df3866c9aa2bda3121f068302
z4e1a61492ee3134ef194595d7cb4aacead1cb4914a0d1d70083398ff8966e2f8b757502257d9f5
zb8ebe136e5ccd60ac78be63ab690d8da9565d059497575c869967ca3586766617dd8b5f9c6effe
z4e86d485258c5499894a255046a0d140522dc294c82e81df6fa8e063e59a78c5398b43f658d0c2
zb9ec3b7dd993c0a71c01edd9fe3d795539666a7887a206a10a7b493e4c23d295e802dd54bbb635
zbe9f6ba3e73487a6f04b7a9280d4108595a681f6f8ad2ea48f8e7e3ebdb05f50f4e4eb93851d25
ze913c41dc685006242b8ea72a00d1983e412d84c95cc83fdf8e5880274e109df9b6c2a64b70fe8
z73e787a6585f172ee649de384364ec8d7497feb7606dc9e82f981f2659ab5407f814e938c8effa
z04e11503e0aaf13763350e6015243909cd7afcf42b7c970dd72c3013d4ab8ac38c335d7785a655
zc74a229d5c289df7375b3d20f243ddb337275ab4c3859448f88219defc493e3010796d4b8c1639
z15749b2ac9c5f8629979bef5027d5dc6a270e8556967cfdca263b5783c55032cc8ac3700c5e808
zb09304e05151ed72f70b27319850ae4936abb39e62f2a01ddd9eb8ea837876a09f0f43fffbdfef
z457f1adec1c767906183dace4140011d9a83ef5b99a2522bccc4e3da3406a4c556dd735f7e82b9
zbba70f7afb563fcb42ba3f66bf3a7e535a19cf69699db5b1b5319470c54a5314c538859ce75f40
za7ec256e9b9d4387842e2fe8bf450fb05b2ced33c90549b243bfc4830b7272b6be7ba688b7544c
zca049983fb9cab52be15a75d0cbb09eddd41017c80f1320817f4f42671478037dfdecab15cf52f
z37f8079aa6b4a14cdc0b302b087230f2bd13a3f50165c959039d525168e00d589b91b2096580ca
z5f45eb6b7c447f8774ea00081255d2a6ec56fd1e56affc43afffff76625412fa66b39ce8c1adae
z2f9eea8e340856cdfab74e8240b0a36fd58c643f7966cb72492b15e4cb3b65ce0c94783ce23caa
z413228a37f7124ac69873a908a2a93fcf135174d4b889c9787f7a1ebc653806e09e1739170e905
z1c7e5d2e2bd03542700affaaf50a92500c5ffc9fa1d4d531afb8e2ba74406bb2b66d8109d73abe
z9c3965850ccc2eaf1e35f1113ae92eeb9210c5a4edbf6005fcc9f9b60172cd762e041dd11c3a16
z6683931603c38a8b2455ba1397c9d5aa24a40c7830cecdd03c640d3b210d3bba42f783f880efb2
zb9b32507f879b6cab352d1ab93973e1a068ef65c2660fcf2a88dd926999e3a5e7b0f44c89e814c
z2d744508378fd9c7a2b8d092689c01d78e953d6d2e492608ab58a5893f425b3fd930a9d9d85c2b
zc30652aa94eb8863a81bb3fe8e8b63ea298de7e731a9bee86d695a408eeefefe24fe3fc05445ad
zd5c1cf77e82732abb4ca59a8f2397ca73d623d46661c7e187891da1a17c380529069e8d842fa9e
ze797de8b575465c62ebfdf2c4150b0950734ceb1034b292c6462ca1f3b77992d540186dbd25b57
z0375677b99befe04a9786b04507566de016b9c381e666d27e9f590bf7cfc1d1fe9f9a79139a1e8
z5c5f56dfac15ec52b1032cb140e98a05ebf86feec95b71306c374ebd012f1fb3180cc47f611420
za7676c28aaaf6b75457c78ed881dbca97589c4c88983a89b349bae1a35305e81714946cddc2db4
zf3359fa0b0360eb1a1ac8f8a19616a92ca77fa2f557c9cda26114b2e3264a3045522bdd1737795
z6e258f3664b90b8abfd5c74a77cba860d755ae44c5622fee77052da4fb267be3845c827d0d9eb2
z57defdba0d6c98d4cb914c19be7ec979b93d8c09ec64ec7f91f5ec3ecdcec5d3fe7ec7633ca4c6
z825c3f29281f437422cbfe1f971c4cb27c2670c31efe8ab970fed32865daa116003fedcbf9edca
z5b3f4ceed574a598f5527b7f06b29ac09058c495c94b470810b613bb4a24d4e1e5a4662170b20e
z19c660f1952ffbeaa06712e866fd7f1aadd5caad8395a24266bc7bd09ea5a0b1ff96776216065c
za38d943b5ddd1d74c6dbd31e04d2ac9d29575b9dd8cba6e1ebf1c8f5df374744f7939465007265
z38fb227226a82f27d106a02024ad030333edb03f33c217a6ec6b56308ec03dd56154554b885b40
z9ed19f48f700f43ca55a6d3bd8ed5682a8cee61ef684988e2d7f5a599035ae5a051f1bf669c37c
zd7c1188443090e1551c7877a01e499ccc6362add09d15f1c2faeace7e8dca94d34ace68f1f601d
z4c89042ecb468b3577404d63a70aea95720485dbb3a833cb74bcaaa8b561ec60d521648ad8117f
z3cd034e7ede8e0e3008b06b8d00f658b9e1fd63eb86b7bdf9e9e3eeee40fe2debf455872b9829f
z605c3ace8ad55cabb82b05489218ffbc2d715e53fec96460b2434ca3f53f531fa0c79b39d0c6e0
z5499db09277f60812f7d75ac27d593d8dfb6f44880caf31a6009c9b8b2762ca408798eeab2fde7
z43e4ad63029c18a9c2be96e41b615a6f6d18f55ed984d5cc11c10cd65b062bacf7f5e639313ef0
zf3421fe63528b050945953fdf035154c8c4a308a5aeb9bb35902c676367cdcf1cae4f25ffd557e
zf7b057a4dae15fdccea0640c3db47033f4b12aa6485695c1fc707d7449bf0ba41fd08661522013
z3c6b771d01f65c2f42391be30e22ad9e9c0373e8f170e4454ac125ddb0a150006faf6dfed60916
zb77bf9820730e82833a282d87af760b3b7be720b18df6b0e9a84ccc1371e5212722b4ead7bb03b
zeada3379747f9d2253e5721555e1d7d3be1f44b72e6731c21ca7e9ec91470ad393b1b0bce8bc70
zdfd75744e495f2b4081ae79b2d8b6d5db2e32ea35e91efee14f6c5dea60992f3c8348713455d5c
z3e55020dfb583316db5c828040f422310c0622736853b3f9160bc6b4190299c5492dfc882b147a
zd44759541a67c01d9f6f9c093d7f33c87ce15a0d44f9cd97d0075e8cfde57e7a0200bd41db8435
zedf6dfecf11216d087e039e6c5da9fc808485b7bf3b29b08b29e37752e7256249b0125709a73ef
z42863f64d3cce90028afef95e3b1db1ed6e5161661e533f038d4d03aa117a87f946072aee88cd1
z498f16456317ed558537fca6e5d7da08530c1f74bc90c5c681639325fa8b92e716dd990ab4c6e4
z373e33bc1c20782c636f6727a5853188e466fe954359297306790e8286166fecfb79edfe0a3bfe
z9d4bd51c60cb234305724ea126b39944fd425c49b2e15be0843b9dd8b675a150237f5b66990e20
z46af4e843658b000483922d284f5c7ac37c331333be93ef55c505bae8462992d28961699bdfbec
zce03fd8fa2b3304fe63f5d0d95d64e49b2b7076d8171d51b9fe255007ca68f71e9c8ff03a3d261
z8d9847debf2151a4fc772ceaf26d28831b3d7cc74c523f57079aa8f326f795bff8a1aa597e86ba
z18e940769b08270a01cb7461c46f28e4f33e606a8948a4ef0d47b1d1cf4848821cc9446d8383d8
z5229434fb21039415b49c0ed5be06d644859410ccc3ed019323381f8cff8b735c2689ca361a02f
ze71fad52fbe5a0dcba998edf68e8ac4354d490ee0397728cb58549b271654270b2e66ee446dd91
z952a3329a3647d7a182c42beca9e69065bdab633d4012f931a08d8417b848cd0e9d44314051432
zedb42996eefaa2e6d8e5076fd171559880c5d422e07fdadfe687e648af6937646b61c3c800bb62
z8f6b6ed63db5d70fb31c42694cf38124110226601b29c2e20fcb3bdc84247dc673ee3518485cd4
z15182659d92aa67d744108d1bc7391d3f204c33b89fd866bd08d41fb13120084dff679b37b24e9
z3c006cb2bafeff4c0f07ce7531c667414c316f790611dc088987692c8e8b96f9620f3a124286d9
zef65da55bfa0fb9acd0bce04800428477a332ff6061fa3e19decf652a51cbe414ba00cd772ce74
zcf1ff28097a5814684e2595ce06a637e00a5edcb240b0a30fd916403c6c90e19c2280fdc6cfad5
zc4e7b2652f156530a9b8a75b9d36bea8d35f57fac9dfe0e3e73928210a5cdac5d28d7c7e09a298
z14dcb8213b23a5b90133d39338c94cecf32de91c2b9999198603fd4574ac9625dbff0d44230420
z5321ae9ca34dc2319cb11cb96e52ac2b4823181c5cab68955d30263aba9b26128996ebeee33af7
z3083cb225bbbcfe3cd9237739505858aa469e62e90fe489f30aabb1b521dc7558b72eb82657caf
ze37cc80b28fbe50f1474fcc3b6d04d1cd9151afe18812961d06957aefd01d367678d734443aeff
za1eba6e58cc11c5352defa58ed6c1d20ab40c5d0e3e76aabb01e7969b704f6bf3b332b1106cc22
z070d9745fba34a223b58eb27132b770ab58d8dee123e0b85b5bbd4b0dfed044b589eae22c70bfc
z8ab529b8affe77c55b8d6c45a7afee36b65346676922aa10305babe03ef1b0f0787db3211a1538
zd52d5ca740f4a5d76b5f03f1b3e65bdf6a485aecd326bdd1de3c9a6dc2bda3fad118b6a2c2e4d1
zd78930e0b34be249545758cc55c2c66fe032240f23e665ca4033118ae797394c9d64cb290acb6f
zb56716eba747cd664177c0e8f27474bdd37f46ae500db981ba8a250741a128955f08915363cd6b
z2a2c1c3f32673b79550f1dc80911cc2857ac9c5ff1e7a066f6b0ee8c9112e07c21b694a12737c3
z2fb359d07ba8790f1a78a5fd3bb61d5c94efd4fe2cc0c615c03ff5e132396cb88bb32204de93ef
z3af5ec069c13cf492bd98d67358b1bc51bc892b57bf0ac0f2f90fe331ceb10e37fead8e6890752
z84c5c168d4551d8f88219f93ed72afb90b9939bd6f5da34482b71c1fdcfff0e30124e5fa6af9b1
z94cc8ca648c9f30e1821ff3476b4c0a17e338c6c136de67152ab6c6617b12602c0a78c0565fa75
z625e77a45bf1b6a6508aed606b35ece7c1ba296121d662e326c05554091ee69ae286cf144ba8a5
zb27ec9ddf67cdfeafafeaf8e069f1b56cf1d2f7cdca335c473a3d658157ff61a1a1050e8da9cf4
z0afbf2263c1ef7535a83e71a2388b1529bec4b7ff4949423f5723f03b8c907c5459a3fb1de4e93
zefce13ba48e107617c30e9f7f87f41506a436b6bbc8aa32e2fd038b69715cbebac0d1100e57343
z4009cca86802f1b4cb3837ce767d6fb694a369a4f016362916745a9fa54c4489b9753c0a3de92d
zf91fc0cd1ec39334e222b8fda871b18266bb0673a44d1b8fc78210a03cc17d3fadcf32cf5ba4d8
z92ac8beee84e726589f7c9a35accc6a344a7b1abc8c8a5fe2b3df58a27d1cf74c2c4345cc5346c
z48888500507e19b06225f614e8094a8e019e5cf4a481487fb7ed2bbb06595838a97b5492bb97e2
z8471e5c4a195095de79d6d7bc28ee02977714d298757a0b94b7061611790e7654b05ddf7c59b29
z89891ff68eacfa85fbd215eab362380e0fc7ea16903ed62aa3f9849139bc21c94308457aa54d66
zcfd647a720f3fecbba2a568f5ddff3278a764185aae73faab7d9f72f638f355fe33aac0b5e123d
za493738b5837021ef54911a4a546b11877c8a68751262822084535ec52a23092142ea93cb35e4f
z0e225c40fad5e6480909c6addd19897931ed4f7edf4b5559edc5c42cc5210ea84a54f79582c3ab
z63407d7d8a4825e185c9a12f3f6ab7420d674b08896df81acb3596723681060d9b44b9b2eed967
z89c66aa1745e52d665db3ee55e4d5844a351e983675ada33084eeafe377e1a6000edd503826158
z2fbc4fae081645a9357f093ee2bc25b35324fccb1aaabb4040f47104640b9eebb163377d6d3535
za98f87f3141a8fe92da95650734040d90a72eccfe4a0b5fd03860cdb653ead6151b0eef3a58712
z1823aec60741eea19a875da1000a8d0c62c911a961afd615347cb341c2f156ca31edaa3bddf2a9
z252a7a4cecf8d35b89f77a82fcfc4e27ee1e5dd2c0bc74d77e62ecd13b7186a4f83bece3d35491
z14115730f2eb5103ff7e0a56c51c8a3fd3b5913d997ea816da220dd4f04e718d198e4f75626d0b
z3f1223bf5a6b6eb034579820aed90b3d749d65afa18a2263295b199837ede5349abdcde15d2174
z2bc12efda4e7ed9dca73316df4f122ed86f927fb2b59fd6c0c768f30b63fb5845188939b5578b8
z94c92a9d4454cc3669f9cc416d3bc25f776f7152608127fac2515385dfb996fd51e2137940031f
z9c623a2e04fa7b9b949b2ffb3c3e71843a84089ea0212078452884f3d5382fe4dc5d5f6479f6ed
z5d6efbe524d860ef5e4aed1b5c8563daacf87537b56a787ad281842dcc2a77875444e37ba279fe
z6ee306e6ee1f196dc6354260296d2f5f5cdee7d2534d430015281e184393c537c403b60c1e2788
zc45e8731c737fd9bb91e737189cdccfdaec0793617ff570a49c28eec0422e8d05a18dad2004442
z8545ad37e7c486c8033b6a382e09f28f2025184712c0ea9496fd28bba494622de6fd6aad54ddb9
zd7322b0c2d5a001972e14ae90ea94017bb1221ec2a479db9ed83e08e80cad61f69928781771d3a
zcd0defbbd957051ee0246432b6376d4026136bfc2eff185eb477709a6006847abd443b003316c2
zac8d4bf250e4d9a1017df71b3414435963778358582437882e45bb8dfbeffa49006064e599a76a
zfa02dfa3052c4a37302cf616751842c0c5b75ca0446c17bf4f811cc4cdb818b4019de58290daab
z42a1e8acfa2ed7f80f1f0f9171e79c254a53af44b90458d824ac2e32c74bb8a19cdb72f2a30c68
z7b4dcdb3b523fbf48994bf896b418d659848fcb781efd528fa713b6741ede0bd39cc4816d7b498
z5fba54cc8fe71acece325723e19435a774323ee503f8f9ecd0f30925504a3b38d5365ddb22738d
z7311639977718e595e0bc5e606e49f1582481f002d2961fffd023aef54000a1b1f3de3fbbec65f
z2efe7732157c666f6c25c0f5ae600078b1a311daae1cb982df6cb9cc76f4663e077b777fe94343
zffbfb7ffe98a11152d4e9364b4aa0da69068effb22436e7f0aae8acc40a6e25bdb725859163af6
zbc7f365738dd6537df184092dbece0221e0698063ef63e3618a10b428d9f5b9f4e6b21d691e54c
z7af1ae8a3c3b785bf0d14b623d22fa8581fea4b8b8dd0f2b22089f9bf26a2b9a3230268d6f8d12
z06baca98c38d28a5fb8d654de7a3b9d856803ccd75e96b63821d7ba462b078aebf8ab319a6837c
z901fbc9be36f9f67218db950710eaceda8c416d032650d57a36b287d9c2a6b5b11eb72f44b64b8
z8b44cfcf8869592e19a367c851984299341390da45b29a3f30c477fbb107a29c91bbcea2b32ab3
zaf5ac158db161d2694a977a048ac04e26534ff514090bcb93a5d45a6bb7389ab144dda2b5df6ae
z10659aefbdca3093c7193c3dced3999f840bb7b80224c94d21bc5937aa50d56c1269e8880b75f3
z120fd58bddf488a421be638e835c1029759d73df10e035c3485c4670709f5d7711375b2005e0f4
z9cd57079f1ef50a35c7fe68c2721fc081b70556f5b61e69fca10519c8a230e8c744159f98881ed
z70170b40eb3bd5b2722b5c76e41d7081348327e3714bbbff7951fbe0467f8f058c7f4b46621c1f
zf963c1c61cd5c5360c4c20726ffd829c14a1576f8f37b38a4cf0e6fdc9278ce849877e47ac190f
z953b924f76e02a58e16a927d5ce89fa5faaa63196cf21439c8e0a1a43df934fba2acd749d1fd2d
zb65e9589ec2bd786089fd296484861afc44c3ee5f6bbb049fd438811ea2fd5f7357fbb3bcdd10c
zaf3b2e2260f1c035261d1eff61e519defb4ead6ff09ecd57f8b320459433d5c939424f28241b70
zddb1bba270a318fcc6e1c2ddb846cef4f2a700f5c7ee5efbbcc01b781afd075c03d1b32b8cb925
zd380d653af6c14fba40a923c8502a0d2b1af15a8b4d3a6c40e74b8986b9b8d6b53bfd8c2d49cb9
z5622ecdc11ed98c247ba612ee4c4df9b7c28e3babdbe56bcd01d0096bde8668fa1261664dee96f
z600ce8f0583fccbb7bd04b0c7cf60dab65649d678b9dadd817dedd225cec6b233e731c71ca4e97
z48a6830a150070f09ba44c0cdefb30c5542dd142a5862c17bb6d5a50be846f39127b68c9538b9a
z4ee35950eca00cb16a89b67469b837f64508ab8620bed340bb468163a0596ef4f1671d5bf02498
z5297ed5c664ee0f35f6b2a1c71936fd920b2a9da8393e73d3590bc12fdf68113694c83481a1d17
zb53076222e895ade3d1c78309aaf44b92fd521e5445653afef1b95bf65ee713c4ef2887d2f1442
ze1ba9155e384b4328eabf08eeeba5ef830e923ded426021fa08b577cf1d53b5518f5f71e045885
z33215a4aba089aec065039d5248e4f13db672d8830cae3ca0c1b3c3c0807feb899e1c5f86bc143
z709cc2a92a451bb016289ba5b0dba6bfc77becfa8b0400d6f4e287ff643a763bb101a96a90af7d
z27358a38a6545310b3cb38e60c4698ba661bfe3b78d4ad4327869bce9ffcbbf8d4aae36def9164
z082e601c10019a04e17f8083c2121fe2d9d4f56c21f9c1312d90f2a33a5f28a1d3c8751c4b8bab
zb993d45806fc08138217f31e579f5ab6fa6a5c0158f3bd98a2191e22f4d5e5632fb288b2564d34
zcdc997d3dd8dc8acb152787b1669fd17e72498963884797d4d9cd989737f6a9a211132dd048719
z9330927cc9508a746293f4f06d376c70b6a17ffd5e01ede348ebe299e18bf3d7589705db0bde06
z725fcf1eaa73a814b23df1acfa109cd33d91842aa28b4a6d6943b94326481875fea297b719b6ae
z7fb5f7744dda70603f3290de028563fcf1663eaab4ef71041b9a58cd5346b0b061e43a2da2d5bd
za0bc15eb4e2568fa551dcc7d34a4a551250b3ab29df28c2e4dc306330c2fa21a860d50a388dcda
z64bf04e6099a9b3efc9cfa6c5ba73291343535182945fae6c43a2ed173ba169af36c35cd9edb75
zde86a66e523c473a8cf872f32cc12dfdfb2fa224f40b84ffae6df888377cd8071d06235045f4c5
z5e548213416a95427cce1a55dd02b8f492af6165af69385fb4db1e074196c644774510eed240ca
z8f6aa46fb50108d0c3f4bef28a8378eeeb847f0ede02356d79026600cd4b78b85a49c428eaef7b
z40f35896ee5e0ff6f08a0e886613f1d89971a292850070951d2d1fcb1c54631c360f0ea4a25b95
z00a41d33bc301dcc464e102617b3c658342cf7efcc9236b196e6c95cf7528b9293c8fd0d3fca49
z5ae21585e8fcccebb36a1e21d4a9821afd2ed2579288a099ddf985c4b5a516970e891e3eaba9bd
zeb09e3429771058629e32811f860e50b624886f96e6e689ec07ceb454dbc22257b9a70a14e79f4
z35363442e5ce14bf932ba019feae162e758eb7f368cb3145dd6ee57d309418431c92e4439c9a8e
z5783b1736459d531e32aab740cb927d4653573efd1910783ffebeb33a2912bbad6ea7aef32e1e5
z06453ce536fd259edf862ec36460c4b8e91b858c7c61196b17041269557ac7e2ed3589cdbb188d
z11d4dd9f49e94d8dfe8cec03b80680d8a866d3e75e2ad8f6083459b97da644cc0d2afc7c38c00b
zb578aadcb3e06dbd952ef16cccceb5f2311349972073cd4a35f692fe716eea0cecae5d38543639
z669161f8ba55569cd139c767fa627f61df3910da6f61d6e3ec7b87db37e07fbc415248b8402f1f
zc5a2428ff8539d299bfb4d4802a755b39774f9870f4d5ef23e7bc303b73013b490705e6045abe2
z0959feff8da42999a8fdbbe255b76d4b5b7b99b91b7369edf807da4f796d40b561dd0a03c085fb
zc0a2275085a8f4e9e391af799299a854c17b35c14bdf1e6aa08fc14a7da9867bf163ed111b894b
z027512e835781c0a36510ed6f74fd3f85d433cc5090c489e1f338996e4b00739011529a79e8a3a
zb32b8d9a748aedc6bac8e588a7abbd6d1cfa576742f74df0432f5e426ad18e9c14116329a78294
zdf48b43d97047c2e9f729730ec40e66462e4adc5fa93fba4e4c320452c0f6dcab70185f2afdd21
z15cb0f65ec74e5a872c7db315159ff05e44a57a2ece09f6484135e3e8d9fe24c5f42451ce3b3d5
z14655aab828b7de13693671eb4c80c09170bf68ec56811861f5332f8ccf064e155161fdecc5193
zf3511842540a6854c6c557020ec19ea4cfc0d832b0eca6e18a588648cb2dd652cbd1cd34335534
z7a6a149d8ad8c68a63ee9811e4a4dbe92e50ea58b69ff2a77699261556ad377459da4e1b5cb1bd
z7a7abe2899e28c225bec5960e34a52bc0bef7ac21619e0cc671c31983649ed532666a8db5e288e
zc735f867624eb4b90028e55af4f412f19225d3dad7963780121019b28ae5cd25db3488cd47ad84
zde0882368e7d3f41ce8e152ddc3f79bbb21ec8143e24391b1eac6a8a78231063451dd0e40c7fdd
zbf17bddd4c26846198ca7bb2b8efe28bf7183c6aaece01970c4248b27178d1be0b8203300d116e
z7df5e6517ed51e48394c7b4ce5b1612f16d6c9045fbc6636370ff7a96b6c15f8e266c504b97915
z9b8904f75f4f821ee7eedca2147ce3be35c2024180c440aec039958bc9f33b2d83b5a198bd9342
z35477ca372abbf74774fc41660209b244737f414dd7be21ebd3de51d9e67f6a1902a9e7aeab039
zd5f23e8e1acd54f5046afece63c4a1533ae157a56dce505e3dccd86c22585bc3ca91a34aac0874
z76557180a34660413b4949b01b39aff8a699fadec147c9966878ca8b916f4cc641419468a30d90
ze4c4de62bd0bb3b65146aa0b01898d16dd92c28c08e3da2d57c2c887d73f4a31b79aea14c738d3
z04770303912b0933f1298a00d307d674d604e057c986bcea1ddd410e104ea64600a37823f3a57c
zbd89b7316405078da06591835c2ce3a690d41ab79031f0f22e0ca35db383e32bf3f67173c0145f
zb64f362f342edebe4686995aa8fe93ff435688ead581bd028227b1685ea714cb4a2503bedfb513
zf1ebb0129000720ac2070af2319f46b6e45e814a707c43df9f46530e363a9d57ab89f08cdcb53c
z68afc0afde1bcbecf8a393ab235f2f937fde4ffb24bf48bbb0fd232016ce4c3b9e1c78f52695c2
z6dad436a66478ee2f5342c8b33ecbcdf86265093fe45eab6a6af51be2896b41b8bd3c5802020cc
zdec862f83c86c2393cbda29e0ac052cea54e95396e18746f9a0b866f13a7f467643596152bd273
z204abb8994a2d2ad06a4ba970d4d00bfd14ed4d859a1c37d16cea54311b36770417058c680acad
z18d2646104390f098e1534ff72e97c4fe9e6dba832f344bf27624cc581f2ea6f9ce5cf7c6f185a
z40445749a2ce98d235e2596be8e5c3ac13851563853b9fa26e30cd717f86cdf0ccaf71047eb495
zf0811913d9e360911f97dd643dc3eeea85fd059caebaf7c6750260a09efd88de943475d3d1b3ce
z06918c7bb9ae78a4c2b963a3c147427e1372cb60fd1e912b30c50f920d4ac1f2149f3885443005
z375ff026abc813179ad536a98f67ad6230dc3426e9bddd113e913ebeb57943e0658910ae7479e7
za4c4fb4c5a95009930f2667bc743232e6838924e173e6ced458e637795cfbec6a55dd66d48b3f8
zee104d0066d5ec1f4fe8b13be567afd82e1d35f1c1963802d2e16b0aef8340ea097e6e0df9d6a1
z504e833c6aa3eb8d1bdbb6cfd7de8274fe39ba0ee7f0995acb49b7fa8c7dd7a9fd3f5907291afa
z0be738a0e90e5395311ae063c002c91a8459ed7ead7d882b35fddbe0fe02d388e32a82245b30b9
ze95853c6fe502efcfd63912c09b29c97e3593247cc62e7b90969b5d02464d72f5cffb6ff771474
zcc9cfecd7c9ab428ec4a51d0c5562f256f0f4dfd6ad9706bb0a159b76e676fa78f25d798a8bc1a
z7761671e98f8ed369021a7ed15a0a868fe379d856179eff6c7ddd2bb8e50190480e766ca8c1008
z07cbd96f5388986155fce887fa2a0b22f623c6bbdf02ebfa93ac5880b7a6d1b384e7aa3aab9fd2
z486944e396c72033bb4fd3795bf63552e69fa4bbf0b4f213f433a79a0c3374639ad1bdfb3babd4
z3659fd2d6244f7297f42204d81d765987afc889bbf0d37323d4010b17f0cf7fe0869c753ae387d
z2efda9bdd9364f7441e72c7aa593424a670c4a1f674c1f8ce8e91083bc01a71f495361a7e9a4c0
z13572a6db1b2bdc257d89d965b90b70348dd02f62e61879ceed4870e7532ff4e85e3bf518cdd89
zd174b8120697c5889f4aa84934f6acdd743c9178aaf44102d1efab60d199dab84ba086b41cba94
z4b718c8263aca471d68e1bccf2e09172f0027a037dfd300dcb3b2632f89e7001f4bcf03f733dc7
z5d7d77e77b78c263f1c743817a51c6f36f560c9c941236042d2e3ec265797f0345226e44359941
z8b7f6733a9430788b48a0be28abb20be54fb42f7118c26c27411a31d1ed68839b8bad145dbbec6
zc7045bd3bb234b2fbeccaf5ef32d95798eb3f0ca4fcc57656aec8d7afef69c9c230152c24d3c46
z75ca3d784a5ebdd5e6a7e0182438a4816d10c82833855f8dfbf5c98fd888393ddf2ab4a6f1375d
z5a9fa8a6a90f35cbbf828d382aad55688b133be22ffb5855244ff856df3099bdf06b732576cf24
z9a93f50f5f5db3a94af6fc7b73b632c789a84bfe5e40728ee40035fe6bb8540b473a1987d310fe
z985aeefcfd386d6f1df2cd95a3cb106b006e893b71c201ddd0f9899674b21ca1be02bebf2efd96
z7906c679ac76cf662a9877ce8e1af818d511ae074e7471142f6190d0a87dcb3eb4552422e5de54
zb8b7c83f38deb4fe05c22aaf392bd78f22cb515d8ed51a4a139af97055d9ca7417d937e7597a3b
zf5d22161bed89d22cb2584a8d646470dc940c30709ece35e2cf103d4b73b4ecf2a4dc26052414b
zca1bf6c63bcc104a290e0cee8779925099cdf4ff40c5187ca2d565268d41b7c4d8b31ba9415173
ze4a6ffe74901de74c2865c9fc084d292bbc78e7f029f98cd0265d174f408423157cf459db8b309
z628e5bce4d2d9dd5b08cf2dd414eb059a77c67c32c4ee0ff0e123ef6f340bed78990427351489a
zaba87afd92cf2f2d798ada3e6c65f3b527a15ad4616e875c5158c880b13fb6823c42ef79476fa5
z9eb3d0fb07980be39b80ed2523397d8f0fc279ea21f819531acf07c7dd61139f71c811acff0267
zb14888031a17b5127f949b58438d1102d12c4ea99c6e3edc8020709a4afa47317638a7dd61a15c
zb1c83d6e1eaa9a00aa9c2cbb88812bde4828b91892aca5cc31437d4a646d03b5571c663105d9b6
zf4f7024be3154edd9684241736b427afd986e4aaadd4eb80ef3d29b967db8fbc94d757d43bbcd4
z2f783d345f10995b43038f35f30be325bbfe0828cbf69db672a4f29e1110b8fba61d017a521746
ze7c3abd2d1ee127e456b58c21470cd629a09579d93c81f30259e3d44f468d1bd087af7b2649976
z8e2b4cb34906f2a7de1398722b630e4ddf8f2808b94ebcb376d7ba1b10e04c0347222177eabd9f
z7c07b55946bbf50c5098ad1355680ae4f0fd44a17015cc2faf06a8495e407ce524969aca179719
z6114fd703d6e3d965381f359aa0ae83e905455562843a786c7234149b1aab613da23755670b726
ze8ae9ce764897d3ef82f26b80424dda68a99e45047738613f24d9aa9fbb07db4784010faf887e3
z793f65080b812c0994160bf277c500bb5aca366860b30a3a6fbea6dd7050e72d2fd42349032a87
zcfc5c0786b819ffb2f65dd567979e6f98635c3d51f9d93ac683472a132b4ad8fbfb1c292ad9e2a
z14fb89ae113cb5893d56d05a7ec1591f97fcda3f4223248305628fad53ee563e1721a967d21e1a
z50ad71352d9d0f46a7c3ffcae9b98b8dd9f587cfd73968f947cb36db10373cff8de040cc3bca70
z3b4811d3be176190552755ea9296ed361322218bb531ebafb003439f9b764a772557e507757785
z6200952cafe3aa859ce2a0a0b9d6b2c5e6f9aae36e7d84130976dba0ad87921957a4aee39c282b
z3b412dd0070f8f4e01b5164236974e4e563d6d1fd21bca49ed2a3d142ae56aff54a25255ef98b2
zecde7ddd333ec760fb36541ac04276257722cb152771df4c55b7afc52566110bdff7dcd2646466
zae035dba853d6cfda8084092ce6f96841f9c9d037e7e2fb61eee9ff8b29a6c5084e51edc848ee1
z494e643b0b6e798d4f5acbe169f882a133108540490df85013c6668cec250b148f90ff863c7c66
z3ccc0df71485fde1e540e745cb75f15200fd40860f860d0252668c8c0948b2ebf2ee1b35e0b748
z4deae99d91dc1e49a4824b82e16596574e8d44e26b8284b0cbf752ac2064cc6898d1fc6ec312d0
z788f178fa520f9ea0d6d3eecc5017ea16eac7d0abc44ceb15b208214a6ee031b8743416df9e801
z207703b7badc1f6f98aaffaa5b7c1ab10b44b2c1939cdc80799b712e48eb48565eb12a6e84e3d2
z6a09be04620be9b30bf4910c71ba7012adca0697cbe0215d6a0edd0690fc6125dd858f82398a71
z7140a2b6050bf38b9337a2bd4b477c53c66f586a8b803614a8fa64d6ca7af7b0fad2bdd5dd6459
za3becf3547497a31fc3ca1963d5cd4501b87603091d4fa94f3a37f47064237e60ef651d1284cab
zef635cf430fd1c6720709741923d270ca5a27b775d0f44c6b4610614c1669a5233eafd1860c64d
zb165a0ecca5011879393bd4bdb667891e0415c6fdbc50e4f771b562720a403e078974c34bbc8ad
zb9f39f98468f02fe0f66eafa270058e85546decfa2cb6447eea1921bcf2171c0ad73e99136dc6b
zec8ee04460f3c782eb21d64fe4c2adb16959d76faf6d23d6774711f33dc17e13937624b354c7d4
z4f4c0ac2d7265eafeb5afd41d1a7748c3079cec5d006d9de2f51f967e2e00c990e557eff153770
zc605244642447a4e1f248a9325495365299b63249d5bedbdcf1ddb3e8a517e67fda1c2d1df6e3e
z9fb230aa7d9535d11f81ad707b88bad9527157a89b9940d283cce7bea18ba81d619891f3127a1d
z78eb7b41cd8dbb379acb8e06a2c521af4d0e4f126c08ba0a2a3678ba94c24fdb2f8ec1b2e3bef5
z0936b3743de63cfdd78b552a9820b7a35860c4dc2888646dd8ea96a7a7a42a5a92a5adc6ffaa26
z2392c2ad2e4666b3ccb13f54d951b982dff6fe24d59419bc91121c183fd63504361c156ec2e1bd
z8d8076b6c4b69fb8dd54bd79205745db3d139adaeec533bfaef367bc877d903c4d28510a41ed0b
z63741e486278a69175aa5a5a7917ae91671c38801df35c8a9ddb748166fe5990ad211165812738
z31aa50a081cb1b46d72cc4bb209a3f1006846142292ac6255f6828027e23712bf8e252e8cd79e8
z0f766b96a39bdc9571e5bac32a9cf523a792eb76b1528a4d64ddd00e9e9e057320516cf2665c0d
zbbb436434d645e1639f5fb5b0d8f73385cd0c9bca260c4218b23e8e873dad176bdaca55c331819
zaa0127526c35cb34a7317f8a5ef34aaecbb270c89ba1a2e3c7846386a31b33dacefef0959d8445
z6819ca98164cebd75b2469ccd2c185e3472d759e2b560d53b0c4c355b1337f6df3a3dbc7f44f33
z0da3ee7ab84a8286ad11dad22ed5b510fed1527877be6241b24616d88c9b3d86cd0dbe344c6c9b
z376a3033e8af7f1305151c809222e12fedf48f8f3d3e69cfb997758a5d074d6ab631492b230828
zf472e47e618bf0e6dcb3279b05fa6c59697ea8aa281f8ec285ca49ffdcaec59a34ee3d93f08493
z24736d91cd6420d19db8ad96d275960ab366bca6a38d2e7e5c5ba67b5073d39d0cd27ba0272b02
z540e0f1c5de283315623c6a5533537c5bed1b6f9e0f9bddf99af4f1bcccb80d0196d5f0921e42f
zaeab7c4aea84fd239ce09129b30b0d4992b325dae690b340b9b3aeda3280696cf28d2d87fcf872
zeae41a69be9c53b4080f81209ff92dbb5fecc0b20ef850f84f517fed864ec8f6d7832d474318be
ze30a0d470c3455a5ec153814284580dc4b313259cf16217a40ce9199306fad4d014cf834a1c4f2
zb845d535bbf5dbaffa7f38f72a3cfcb741acfd2403cee524b91b7c81377030cdae462c38cc957e
z9c4dec17fe46d332503716d9294dd1645ac0f56785f3ebe4ab08fda333abeaca6a3d55ca06f7c7
za9aff52e8e141173fd03599fe862afcb9e9e1de0d2718913d6508f98b3290fde3ef5f9e000b434
z7842b33eb3206170d553599c842c20d86328ca6303063ff0661469c9bb3247492946cc66347e17
zca882f36564544512e02e3aa207ca65b3fafe1d29f9013f85503fe6e5ce4b09fa8055dc1096449
z7abf33580a2ec124bd9f52ce9902949e849be6a5a2b1969db6ebba7cd5e59efcbe5bf8bb9e8188
z0292855c42befb169bc234ff32abdf9917905a5799d5ad24e7f35bfb0a51a0b3333afd061d696f
z96862dafbf21eda0583e254831373dac76583689d9b70b78cc56022f8eb320159c10f5c1e4ccad
z9151fc41dc3e36adcee71b3d37348c6fa0229520e1499883c3031f347b0292a6f02ec8b2b649dc
zd4b5bbb9fc9494024dafd85437bdfb20784757f4a1e85d5648ceb1b58438c6bcc3c33a45a58658
zbec12a2f2c8e64a6d6472d8c095dcb07e8bf0780d9fd246b4b5c188ccbb5ea785132c6d8ca9116
zcefc2a7b9f1cedc239020fe29657a67d09b63c64c4cebf9218045c7e288e8a40121eb634bba0fe
z9a016de504c36dd98c1486b55aeed0914647e65dfdc6acb2fdd7d435f365a97af08515ed3da953
za436038d7f3de4882186e1ec52030607ea8ef07196683ad0653364ccba90c025e7e9acc0b47021
ze11fcfe013b19ba988bfacdd44d32a90e44fc7c7075fa471bab0a6383cb5b17938ee1b15762e46
z3aae3e549feb509123057a26da6471b72e8ef2ae9e79e6d3faadd3290f59d4fda67c03ab9ec4b4
z083abd0319e1437b68a917a2cf5e220bd2a58cf573b57b88f007a344dda7dccab0bbdf86c7aad2
z3829cb383c329cd1ecbf443dada59d8b31388e72b2b877a557f5dd655014894e2f3489e109ccfd
zaa0b77c9609f1cd7e0d8231851f350ce08043ea734790e1f0a88966f0a14e38c46bb81079ae1f8
zee43ae78dee7ac2b51c77da83b7483712551e12af4e9404dd327bcac4bd18ec2238dcdd7a232d2
z31ab6582816d1c28cd8a104d420cb4278ef0545e86d3d12123208e23d1f097c4d1ddac45c02f19
zf2a2246452f380721ffaaf4438343743ceb90eb4b9a6a903edc72fa1f4fe3f7f02651b591db965
za4c8ea7310e5a6651aa07b9da55ca5854433b0ae42307a7a456deaa55acc3db9053453926af0e0
z2865deeae69531aee297995195fc5118157cd58b9d443111cb69dfdb136ee859b2b8e5fac6c94d
z785c153939ab6a5e28a16aaea2fb528f0c3d86c2d119afda6200747b90cb3b9ecd7d9f2b819934
zcfd183d0c365094fdffad5eeb874bd050cd4dbe23c88ecd0c14b3bf23e4890d636936fb4429fcc
z693a65e41d45f4dacb89c32b8fc6a781e16ab817b4a457e884783695ea0131803691f21825a8c1
zbb73af8bec638877a1ee1cf980a378a79fad6f296e7d40af62566179cb26fc7085b26cb937b936
z23c5a80e2aae02bcb3109d8157678b9f1550360dace9346a3666ee8cd7c1b913a0538b7679b92c
z962362c203e35c0439629f170aef89a6b249f3400beb64feced5c1d35dd71c81822b44d0135935
zb8719faaba21ab2aeb097d0219f7a4e76785ca65e008ca7d6b0b1fb77ccd50881036a52f3f29ee
za3aedfc0a7cbd053d00ebb6fb35e6cb5b127a957e09b6ed36c4163b72890a29dcb7cc0a5fd94eb
z38c9451e4180e9f4028cad3e645618631d35d246e172c85199933e419ee5b304619a805be122d5
z6f52869f0bf6e1707a28ae00dc40f3a29829249fefbe93c5269f5e2c345f85307232087d3a20f7
z741d6c85541ffde3c87fbf15c5007cf8ee3f06416a7124651bf312434dcdac13592e977741af65
zd43543871511012faafb7cbe42b2dd92de209551c0f842720c9db05dbeedb94c854319584a5466
z54cdcc8d9ead254bd6b70ca6b92dffea8583dc880eaa675a6629255f15fed3a74da26304cd3acb
ze7fb3cd609bbcb13b552d65f11fdbe7222f444575881d4439178456e7eb60777a5c74c8436af6a
ze2d782ac0fae3c93b976744e1485353a36b278654907402e21f2963369875fd379629895146f56
z788d9bf524eb35eeb03540ed09aa5e44f960c9e1e60cd431f161baa9ff0396d7bfc3e262da575f
z4ebd9e16a2a42e716ade6c87eb0725933d87a6e714b1025bda3cd53cacecb8cecd431e70121d76
z0cdd1ab1b58f686a5895e5f0df274eeb13d9f471ddd1cae475b5cd55851285e4afb32014b7266a
z54c59e0bc2f429a92ab5902ada53b3b85fbce423cb1f68349090b81bd218c3c9157855c7c0bb22
z7fca93d0967eb5fbee0f93523315cf16c5e676c647e0716d84d00095253d3090da7e26aa88e52b
zfdf40e073a5fc21c1bbd4ef345ee2b3ce639b79a65557a9736bdc988e74cfd23b843d5cb78a8fe
z73baa82beb4b0c0edbbdd9b9726ae502c68092c4c4a876b508d3af107b054a66ffed816da211cc
z049f08bbc256d8c07c1e66378e72224d91f895fd6dde75e6e84217568de536181fe9caa10ca924
zd90f7a657bcd311b833a9b4d013c789c5b1d8da7a81be119beadce0a509bd0f6f585f073b90804
z2ab4e96a8f7e28ba0e86fb74690106a9f692701073276b7ad579ab8f65fef1d430a5f4049e4698
z030bf4be466e2724c5aa29a22e16e0c4e9553c3b2de08c6cc246a6b855f50b8cb3101c0198c8ad
z0fa02b5624d7894095fc6aabd08cfc9dc937c99e7248ae64c19d71e4d169bd182f821251934ad4
z416d934dc0fcd0533823e0744dc3a088923190fb1069ebb214523d990c225deabe21c7bd6b7885
z38fe8ce2b543b5782e59e9929d88f0f251ec18f509cdc95afe4f819a899955e08863e2282e2897
za52775fe46f05a42e983f8d44c26959f3246417e79b43af5641a63c9aa343a9b638d96af9654eb
zf2a6ce9d50b6c83a17ef37e0e9854751cba195e72efe7ede675f602a364e758e322b70ce6c651b
z3e47cc08d2c18e2968f6a9c9ddb102f7ea4ec0f57e88014c572b0246905795dafabcad9b53e833
z007093c67e958fefecb3d459d88b3df740345109a7492357379ececbcd32c60aa532f374642e33
z0ea6cc7a751eb262be4eb60c5991f8578197b946af8458f7903d34c22a584a9fa20646e105a7e3
z0d38eaa43e23ad14b07ff576a2461a6a642f9b6e09fe33c06fe74e1ea023af89e57c6e9b82aedc
z92d6df8c9ba3f80110420ca4847db2afa8d20175d7d049d8dfd1d57c10e52f391a8d6b42e9330e
zd929b4d4cea20e82e9658c7a5ff9b571039cfbefa4464984441641fb4d4d668a4c5b29cb01ec9d
zddba0e6f6ed9ef71d3c4c94e618f8d9ba1c7fa3227f94e6845ebeb6536c89fe1e409e46d981fe7
zc7c9a3c9be08321d7ed44d615d92482ab3febcc8f6ee73f9131ecbfea4c77e848cf332f5c94320
zfb4933408b79b19ad07f9dd65c166918f9ef2f68d38858438059f6726b4368b89e4812e9a9d739
zd3259df925762ef44a46d60012026274e8c2abe369e691e911dcddf292a5c78f1d10881c9ab73a
z07312db7846e524f96284b9405ab143b91b24bf0341d190f56ced689319acf955a3c933e0fa5ab
zf21911a24d079a9b4b73ebff677424b05f0823270c298b99b9f543bd878e04041bc9c8db10a57a
z2f29500a6085eb0c1735593e4776d0e974f4135208e4eb61cd7b04f03e4deaaa9aa03ca500d155
z4228f769a871935b575502b220b88a065f391b6a537e15c61e5b288b947446daabeab9585719dc
zb2177209903d67779b2291488e73a15f290aed3fa9d3351ecf28301bcebaf2fe2602d548a6d753
z985332589f2a8ce8bfd51bc29c2b17838d4db086835e4c16f2cf3d496a976da7028e007cd45728
z51694eb535f7eedcc1d93c9fd2d3b580ea5edbf00086b861f35d1ce6103db73494315e4403ea6d
z67ab46c7259610770e96c7d3c133d71aba0ce2c05fe78cf81b029906a8d4aa74cd87d87212a266
z517f295068c65ed7ccab313e979eea8a442cd99dd68fe2d0f50ff6dd5f7967bf65df48fa61b093
zcc62cb622c48375269c51a1a22976f44a74c8d3e30e48043246a8a5f895697d9ce6b5c522b5c59
z782cd3d27a2c6ce1797a38d6d8dbea086cac181bd3fa3ca3c28e82aca86b8b01cef724ec927282
z2d33db237218437c94d1bbfedea18c35b337af3b4c9bcdfd4b9a82123d9d9e08444113d7daa67f
z195efac042c939bbd270932547202ac024e95bb05d72356d2e6683bb9b380bb9819a25391b1d81
ze6f55c49f1e402ed6ff58ac0239fba42109844b74e838441b01775d367c7fa1fb9b09a90601997
zee08470fd4ff3afb2785c6829371d19680b31b385149cbaefc80f45d4e12c4206a53564747026c
za3d8e0be62b3d0bedde9014330b203375f2e52131bd502a0317049bc01107bc4e39e7cf3aac56d
zd0fbe72d3bb1484d019ce67c35be48e5b4421bb5b1090004a6dad3c3614d147286670ae27c59fe
z31a5301603a9e12c209b89399379b2ebe518f96fd7f8510b84c57457e64e0ad2bd57fa7025496b
z3e339b05a70b96c84b67c3f51a50d3692fe4970fb3a9e1e6b76b65f5b66434450888c9851d6081
z161d743b7ffc048251f8231f96c098180c22ebb5bf5c1bbec1285484a85a7f948d95bda1b9f096
z9252d0c6797eacb9c9d9b59271f0303075da3f2822ab94121f6ac2336d8f029f6c91e4acc370c3
zd0af7701515165a6b6192e5b346e7f3ed9ef35dd204fa463d7287d282b3969105c56da3d5c95dc
z527d43ae1f71a7b359f59bb5bdd8ca05f86d6e756ea90b61a5f03442eebae9d25764b9811f968a
ze4b9ce0427962e6b69f62626d1226fdc1e1d9d3ef470a880ca55fed97cbab07c6caa03471e3d87
z956ee92510cf53c5e911398b56df8f3fdebf879959a8e7a1cdb3dbe11133e50f0d3fe28832119b
z1122757ee37a7bf477af7910072fc0d36557bb4e168a688c6044c667f7c1f3f065c1f51dc4d6dc
z190a2786812f0a5c9bf93a96146ebbfa47e7067828915be34b20781a65b1a208a46fa0edd6369a
zc0b5d71e17976136da006ba3be734748a79cccd2176f14aea1e50afb7404bab34ee2a78077f6e3
z15e8e90a5e8c7d5d45f914c5e76942ab2b4e9437a0b622dce52f66fc670c531c2b41d56a243fc4
zcee676b24d0479d7e253c8567a6366cc96e39d5e9f73065ba3273fd670629e1f69afdd5cc096b6
zc7352dabef35c61ce6fd2fb0598703a9eba13069fa3ae228b8c1d87f1a9b83fc82cf281998f9b2
zef5623e3d8b88d68e3108258bb76e0e91fb30cfe4be00a8be2848777ce83ae5268518c02497b78
z61c365aff5d4fc689e504da36eccab9d02efe0e32cf43d72e1930bd511ae565aef797893be35b9
z2ea9643c2ec4bfa9d77147a388467fbe19ca6abbf34dd8018042d4a9b778812ddff5dbb084ab12
z26975dc6146d169cc7e1bb13c4e015045c251b588d9b8adb5a959c6187fc08054b95012d811e2a
zff922fb33e98f0b8ff2b29298e3470af5acf157b986de513710ff079e318276de2f5a592f14997
z624a0ce30b0d512e529c89e97d10162941678cc72673c157cd3718ce951c56fc86c195273a2d84
zaa125ea7200eae4331a951282fcbdc919cb754e7cfa4cb273d82a8cabfe45ce8a73e04da47b98b
z2265165af63459da7dbb881cdab2869a197d677868e08aa935db8069ed675a4f469832e85355ae
zf6c82be93f56f4836a2ed0b09fe5da0e643e0ea36de9afc43504f080059543313918817ff9b49f
zbfdf59edca9dad95eeecc61bdd10cbf8724a0d455735cc815a64720325b7c807d0ee910ceb484c
z281b94b64cfde5b74ef8fa6d22e4bf1cef294fc65c0478436026149bdc38cded4e5b70c33997c9
z91083a6d38bf41f9de626f9ff5feff1f74f4d9ca4501e608e5dfbb7ae6a35954cb23776210f772
zdfaab9b2e79f67ef8c497ed6f2350cd9ce029c9a854de2d04ef83ddd616ad42fcb33d47c0c0601
z297277eb613c632acb7896966882c3b77a2f1507c81f00a0c5a7bcec72f44be13bb0f88944e216
zd7ce761e1e1da6a92ff2379e4cca7dd7d35381e7e5d0f46d6a52c86526849e95194b1899d00f16
z8e330788985f4e8a83003f96dbb3983ae241b59fbe55119dac815cfc099a63ea32e1f92047407b
z8d728b0ec102517395043bbc23eb2ce857120dbdbb15e1409808caa48d56a776ac1b4fc0a1b287
ze58ffc476d4b4baf1f48ea0ee4ba7f3b2b4aee322c14e575163df4b3a396894b7a332f2122d86a
z00f9c06571f15435141d1bc408fbfd2b95026f994b93633ad53cc41d4037148eaef4ea94dd10dc
z14e7295a4c1a542ff3a288b7efe2b0a193856de812717412736faa33ee564bbd6e34ea3d756ecc
z6d1f2cf33479903ce0e6869ff57db4b92a95598bab6093be2fc1deb2fd8c8dd3681a3f82a5f284
z012e60ed6fa10b3ca00334a7aa77c2c7337e3a213b58027b13d4bcda637f3024c6344dd07c2c86
zc13ea53ebb6a47792e6876c353a8d409f8d3f021505e32f1822da2e49b9487312af3abc544115d
zcadeb6663ab4ed19e05699bdfaf45324c529eb82130668341f7e28c15f81fe9bfade0f31578ac5
ze12c44a18ed07a867d7d88cfa45a7ae3620dcbea138f5819502df92f95973da8201b92e6ab3c92
zbc2e98f050f234b635830a287d8b9b3f1c7fbd13c2c2dd6ed53dc9093f7e37d9df927b0fe1a19e
zca5d71b7c212230ae0a24e9fbab784c4d60b13371530ac45393ae90ef8078da33f09c3bea9c145
zeb59575bc342294735d1bdac813546f1c7dfb71fb36829e5cb4e77b212d679e7e7a5e95f8c4175
zb91ff625ee4d85565485689ff47f609ae50d8691bf6da79af7de376f24a9c0ab31a207d68d1061
z59cb1245d37a4fe0f6b533f07bc0bf9ab68700c239bb5700346053d740458bc8dba5b49b90ccdc
z559ff88fb1f255bf287993b10cd6beee870ce1884e5f7da712ad45f013c68a587e3605bbb605b5
z072d610e3845082b93d1cacb92b3ec641db7f92f8b5bfc4cd8874b6017bd80eefe182f615eaf40
zdf4cfe794789dddda8a4848ab74ffa2ff8fd7460953ecc3745636650ad42a25be13d893221e7ef
zd3122700c5895257b16c0c8cba622455227f9c4f9480b0bfcc0db5eadee04abe9d81db5d8f589f
z99f3879e4bc35905d0ef8b04ff176d20a675b91feb2dcf30c7749fb92f69af656bd3926e3d9775
z09cd9f4412a3772db116702e27fdaa9f1ec5e861d2542bb885b9cb3650c3a7880b30f29a5e7020
z163647f6e54f313fc233f84f2880c3df37e6dc728a43936065f3846017604cb9338e4d65e9dc61
z5a49236c2f15658c25aeed68ebee0f94fdaf1a1e3d11fdd617e86b94b63bf32c56cceeb6c762f3
z056aeca89a27df4f6d5b92811cb2ecbbd08ba7d49e832e838d6bc32e92e05c626222344e738498
z74c73f06df35dec720231f400cbde2865eca4bd2830c26b0308916254c9b862d7f5d9f9a6bb2e4
z50e17dc6fd25a98943eea994e8ae618d80cbade8e2ac180e3de4e56aa6b191fc119df494f01582
ze09c7535aad1715c64d72e6bdd0ce4078ebbe52acfec7f9cacd84eaf79a9bca6e354a44d095ad1
z5fbbdc2f650d8d6867b5b9a0fb21e6e7d34c3d9792d150d7ba5367cec0270f752e024521724cf8
z283ae1694d12a1b9e8a42d2815023f500679a8d45215b7ab8c5939d2d4a91c6ebedaf5cc3caa4a
z48d04151b79e5ac506a0b27487a9e233369a83f23aa4033b377d379dce0f2be3ffaebdf970add4
z33fb9cba5b7560c4c6097ac086282eed4de1140c12d3b5e19ea51d8f6c70a881f0bbf1afd33ac1
zd5eec3a63b7bcb5f7d4cc9ffeb051397016183759171a157199726c548748d4cea17bd57e337ff
z69faa728b4ab7b17fd74fa331efe81165130225482a65223590468cbe6b52e607e90be7a3aeb7f
zd61afa20206e5a29918643abf82cb876e4b6efebdd60bc7dbfb2521da85e557931739809a590b9
zf5367b98bff59736a82b56a574d0bf580c65df8c3b54cc2d5eea7e73366de65ac3be05f2ba7b37
zb736461650d2da3ce49ed4814bf7fa6cc6a025b9f7d9a52fab113c664b079edf5165f9a64051b2
z5e211bc0425304eba04b2d1b19677bec1aa7045f3948ab9ca43b12e13675b1306bf007c3a502b1
zd83de2d233274637914b85467568451d4c348f30b14880c99030b5c7ad1f0c5fac58489a9a38f6
z845f20708eb2f7158a49f1c5990fe5b57395f31f8fadcc0bba01a21a2997bf7b34705e4edb07ff
zea5a2f4f1e5e88b8bda61b1efa06eda3ecb264779dbe472f635af8211d69bf9c14235c4864780d
zb3d83ef0f6cf1f7b86b19972227364cdda22fa99ff6351d978f9f531fd21d28bddd335fedd322b
zd2c5ac9d1bdc4c041a777eacd6d0b7978d9f61023095400b86cb842373f87ec55bbc4be725d268
zea18fcc897c323a98d821230bb7bcbda28e857e818b64b1a77c434d500b856c630d349fb5830a3
za12a44e07cade64929111b3d416f6d3c16120e43e9e377334473a3738b212aa5d7f944bbbed94e
z5b918cd151c37ec250901c6fec8b1697c0527936c1813aeb3b8b47ca6080ff09653e2d51d70756
zdc082c472fec5110b0ba056648e378aa6739ae6e4b6b35d88886c2cfe6529ede32590d32f3c58f
z7b2e39b1ced4e64eab995894087d5260698faa0bec6331beedf485b4eaae8d9af08d413f7066f3
z9eb738580dff8711af75f4cd27b79d8fc974c5785be26069964b312dc5a01f81c6ff5fd1f2d582
z5e124e4338b933aa15edfe78a7476858b5de6d5319f37c986ae6cb4230192986ebe380f2fdff42
ze735d683de8e0ba2fd7f182d97873eae501fdc1ae0c9aac40e921902b1cdd859fca6441337d342
z0fd648cbb8d215bc9d4bd9b79820b2f0dd61bd7418c579251dad8670b636219496f30071f30b64
z3d3068a78daee506e7cb18fd93d083ba8007df43df7b4f555d25b5a0b1b808f405d59577c2b8f1
z5b8de31150bf347f44805f8b71b9404636d73ae8bd5bc7b7aeedd75af3dff6b6732f4211ea9bb5
z5360f70592546ba9bf56ed4ad1a74dbc8eb9e169d858e49fd748e3ae47cc7c4261d810932831a9
z28f89ebfb22a340a7f8962b544a70aaf0f444d193d6a4b295e4949e7ecb7fc161e425db91de739
zea0c76ac15e29261b6227e9946d932439aba3fb24c2913ae42c197e615dbd761454655a48eed94
zc28ae58d4dd79821046fe4f98fb6b4c3dc50fa814862fd08eabdf473ec038898713531ddd9f063
zcb597660a59af1d8eb57656656375ca49ed9d15e77a8c61b3a7991e4e7946fa6c124667b4b061a
z9d94b22df0f1910b577b5fa3c5e1f53ce64ff7f76b64e06511a4f52c0a3d0f228f135194a2bdbe
zc75a3c9d0f1339bda7e85e2ce56202bf49cee91cec93a35944c49811c4d6affbe979f523693c81
z6c91b83a3fc6395f0869eebbf545a030b5c79cbc57b0a433bb192ba59a63768c2cf5dc17b19b3b
z589da0a07a4a34e4aca450a86d27621c7eca17fe974137e6dfac3b22c798c3cca1891a305c03f5
z02b5cf7c5bc34da48ae41b0691ddc579743b6ae2914357a6e10dd781d653f0b6d1f09bd9614f4a
zc25734e533f91b2a759bf32e1b969f9d351a4ca74103b5d5729367647c01a1a29bc0dda1207578
z1b4f0b966cae5c68b1e6e7b065e9684d3b7f1e8b0a920cdfe13e71106333cc3648e808bcdc1948
zc8d367debdabf96f6df4f5c11bd58820d290c1ff11e58b1782ba7f8250e284fef5f6ac20fc0b1c
zf129bbd91da9b5ec9326ddf7717f45470d99d24d5d21634c46e24be05743786ba44e9f08fff58f
z1aad7fd6ccc1ec2df1c201b9568acc7b297359c54ca4633d6717a69eacdc0003ba5b040801ef97
zd94b9d0dff185901cff9cdaa389dd7109a16315c391171661ed814f0f92593b0ac0e2883292f73
z61576d0cbcd6fda0d154bc919a533929577c5505c067c3201d6d772b46adb232a26222b2038506
zea34116751c93e7374705903c0d15c20e7ca81a08a763cc7cd7cff12573089a0981869d7607f34
ze032d024dac5f968ea7889bc54eaaa4ae717e8507d08cb324e411e014fc19dfd5f6a705c34674e
z50df2b0069abe507b5ee2234fbf2214cbb8e0305ee5e3166b7c7ebe4f24241048b0362e646d01f
z90c6e4402d168511b6701bab9ac67bae3afdab7ec5ab825bbf8058669899ce2ec399bb27993ed5
z395ef83c77d82a11e5fa9d3abba1d9a0d4dd440a3f137ce155e61b28df5d8c48b118c512f061a9
zb00d395467203726ad0bf7d69d68bf569c149ceb1a12f8dc56146a6bed5c4efe041ebda869b51f
z496bbfd7e0c9374fb9e6904a286e497acbf2472ccb46f243f41f666c17a73f9b11da088450ca03
z6992dba1c171093e04fbbaf9c5da9ea810d5a7fa578bf937e767cb120d969828f47340d59ed573
zfd195a478a99e396b17889c29ebd9f044b75380f783bbbafae7168ada976adee62d68e429a7b6a
zeb8f69f7df9d03307aab3f008c59a765caea7aab60f8c726df1d76684d3bb0e35adc8c25513ee1
z0eea7ed7b592cbeee4a64257d08e7f6cdc364ecd7e196413b8377d00dcdde49bdb59c4c36bd9c5
z8b1bf82830d1158e3311341e2aa2f161ff6b88956248a12d2f3f729aca3dab507e8f2a20dfa24c
z8614016cc4df05240aa3893ad0972a09715a7455d7334914c9da6285e64343838e7f05140b8b03
z45b7a4029db14b0aef9b8662aa4e7a99c918c4928a5203e910c6be7c752282deb8b3ef30d20ff3
zb93c733f376742b0dbc8786d23de591f2158f5331cf9699a9a70c10f2828cfafb12dea45d9fc6a
zf867c9ddc0215931ce86860c7531a8db26690cf8239b134b3cd66642b9dd02963fe72554ab8834
za71313888fa826a92b7eded810f11c62b0402f3017f70e825e43744ed51eb9c1f9db5d71a57f14
z71c51c33817f0dd63fd5f54bcb6f20a3c279e7f26778dde995b51127b4773d11b7648e7978f881
z69c64fa18ad0cfee9e2c133d1afeeccd516a4c5aa63e47ec3e928331317ce7d860085b5e3c6f91
z68adb7d7fec8e4fd0caea20c65d522e0bcd1aee93494b9da127461a5e48027a0609a4488487b65
zef36f5e37e1aa43dd1b73de073f11556adb017d58afa96902eb7beb76c8763cd79930bb6cb6044
z7a2eddfc7d834672792b56a4b30abdf64ff6af9b934a2839ac7bc55c5b416e759084bc7faa8c44
ze99f96f1c4f29abec06e90b198d9918593462cfbb70708746cbd844b1d76c862604648aa0f1669
zee4acfa1a9375bf8b1272c632a7c14b8ec03cdc61b3d9de5f95e562d4fa9125db62c61284c20a1
z62508ea30d896ce539304c77ca4eba2eb0b4ba50df6e2c3937f03d1f776cb5c1e39b9a89bdb80b
z9fd24219365768dcbea85042d83d1cd8e23451c69c4f4723745eb102d5d3b20d5dd654408e21b3
zebe65c9389c2beea523c6db1742e1f4c5d368a282eb10d28be9070d38e813e0a65d057eaa37d5f
z6204f4193e029e5b7ce04212c99ebf39bb621477e89fc5376f381a1ca303984070ae3097b9638c
zce41e8ffbd7e037fa8194f6c2258e638a1f097392894ebe727fc520d45e988fb4bacfb8b876512
z3ecb84c9c5d9ebe7a0f7ed2221b3670ef1c04e07e781c4545cbf845817c8609a512fe84166b4f0
z184f8ca0e22a1071eefc538f977301335d4ffe7828d1b477c293f2a644e8d58d54a1fdb61bdd06
z3ab149ce5d9b72cb5a350beaeb43cb2bb463086e25603798a3f5e7b3e29b90a2b1d9a25ba206b0
zf966e5e6c734cf931a76c69d78d1058e09c4a9d78daebba773fde69c12d1a0d330c29624437b1b
z8bd1f1538db2f8705159e5a72efe8ba6e2c9ee7d861cb4baac71c013c0d4962f0f1b0cd643746c
za0f84617a321329fe8c4f91ddc0ce05d688f81746fe3da4f4df519d6781fc807fb78349981fc60
z2371c0ba11313bca09a1213889b11bfbc2e3a9790257fe77357061902d72a82ba858ba23630281
za7addbe59dd8310cfb2caabe63d5013f8e2ee41b87c6cde4bb37e4099ac9201c8827db2bea3ea6
zf2da564bfcf5399a4a899713da75313ee6b785504a84ff89caf3162c7403deb667efdcdd2b299c
zce41af016a01e35db20539ab5f77e9af5f2f3dc7144535e0e749db73505cfba461aa1fae5fe402
zbf300d3e050624f09998981e210cd366a3ffe0b7362201df5d843566163182efeb8aa6f426dd4f
zac26378d90a61b36989cee32cd3c6a2d02c06b5f5dc754eb147e540781cf979160301ca268475d
za0894b0814103ee6a843bbbe24f33d67613b714f662b11d02dc91c1c7823edc0999a607db9acf0
z05b8fb75421e2f9e8cf9fe5a7eb6fc8fdf07ba210158b39eb0242181c0a85079821d5abfa5bff2
z2e04af445fd7e942a5ac938d1aab8683b3c9dfa349482a74baddea1d27b5f61adff8ed99134477
zbda854b67a2f9d77dbffedf7bf6d9725e49806d89c1fa527d4bf67ba0326cf95a3347cd51f7dd9
zd9d4f33e40ae22b4bc72ced1aa645708bb711cb293fefb0b3c6d856f827585aa18e108057b0b57
z9a5b80488444b0a0e0bf9ec0d32aba120ecdf726a33e591ff8e12f5565161b324350fd1ce429ff
z84c2ec31141c766362793c37ea1933e960fcc800bfbd10f26e68b1c669552a201264ea14fda055
z898d48955c45c883064c612a2a0220d8b623d9a0fa022777e2a9c1b7fb36df0204fd7d319e78a8
zbeac1eeb638a736a5bc4ca62fae5965319e513636525ec9b1556831abeed487ef5fac7c0d2663f
z3a213f07fff5970a021c4c124fad418d1b33ef6040aac6bd9e444058c60a4f2ea207431378fdf1
ze82b46c2456a27b2a398c4f55bc62ee76b24fb266707107c6dafddb414bd3f4e5f21e3f4ac308f
z666433df75fc5de6f3db39fee91b391cd73e0e3c6f9647a71bd8e86101487fe9448be042195f89
z8ed9c91c2429414eb47fc070ffa7f7a5df2dcbe99b82987d9ed28661590cf16325f0bf68666a88
z4ffa2407f0ff4d24b34773809555c46f94cc96bae59f4c6b140a70627d805b08e0553c9b19f0ad
zd171aa1c69c6f07d2703779b76ef0d467d676bffbf3937585c09589ce5bfbdd950453f63413aa8
z1773ab83b07f842309943bc7bfeda1a6b78c10be9ba24fc7dd9de1f3c677fe8a47dd81e38d0b8b
z21da158e90602585cd2a5b80c51076dea9090fa725a5abd92ac7cb2afc0935276a7161896e32a4
zc0683aa68b84bcec1868e399cbf365a128ba3d9198b182053229654aca1ecd8d249436a60dc501
zf6d6e09916961ad8741e4b78635fdc590782906b1537cc16c28e0c0243e300f7cdbc82f1b25c8f
ze053e70d7b60fb460d2a55581913e04d31abbfddbb80d78fc507a7bdc5edeb403ca0f55e134b78
zc7f8ec0ec3fb0c3a597c8878f1843b4967f71f61ce643c9c57843064ac2e9f533508574f53bb91
z702e49f5dc19c8f0c22a47de8960b1129b17a2e21b72d99464f0faf12f71e75fb38af8b38eb6eb
z34f53853c7cde61f2d99116bc511b66adb96873b4c5131ed596faabfed9a6d12688d444893f163
zc97ea0c2af6cfea912b415f5a2dd5e9dc7cf9060459fe0d0707b6800e680e76d97cdcd36299a66
zcffbd91f8233b87792c3cd2b7fed13c7fd815f4b9bb5bedfc2a2916afb0b9a35d8215963d6c1fb
z2e8204c912b67b689a901422a1f29dc7a7c2b8511868cd9782c45d329f641d0c176c7741780c8f
z5359b8876af3ac05d9dea4299592097fc12fff0863f3b3e82721fb7fb46f2958552ed45edf714b
z66c057e9ffc6459a832f0854a1026b7cd1d19a66a0104c729c8a9a2afd6a4cda5a8f7c95abbd9f
z69d2086bde958d4f092b6f29369e5b2f9bbb1c9807c65dc72b04b909fb75491621afd9698217c1
za0daecc50b5da08ac60551c1f70a5102792c76302447ee40571e62c41db7525cf527cf8d34ee1b
z1ae6459e753a7b4e3e11c24c048306323acd2bc6f18e5ef7bedaa54c013ee36c0537efbbc260a1
z694dbc28ae7c4c1f6f23a1ea78c3b9cd507c8b83b018051252958f53768735f80626ea2b91fefb
z0189fce76ee0203c40c55083a7514f98c333888427feb9bb22b9d924761167b607bb11f0916339
zb2c3c359ce289c4b356303eaafac427c4d9940749c6bb02856cb6476215e2bb9e065b27212f4ce
z10cc89f624eed0f43f640e781897be8fc234c284341106b11eebd1ba95dd05aa7172c7df9367ab
za29caf1d986f149b46d18fe5b3a80589544bfd788aa8f8a2e563e9f5457d2f10eaa9faf30a12a7
zd63daeeede2accd8c00dc0c53cfa1832119dc08d0d4bc404db54b37bce45171020dd8919f793a6
z2a21cebcd5540f01c6e9f049b6f519a01b26e989a7af2e3a2e5d703e01b5515e720decd2132dba
ze467af12bb3df66c5bfa45ac35a563b1394420700c2465377ab86e14c9c4e685d44a821581803b
z4140290f6aae59dfb12cfd55a89a72f0ac6d25638c2b56d4ce4af61a998054654470e348bb93b3
z8592391d3d783dff6bfeaf87d5a0e5b6e1449b52a65063d98a72a481646c037ce24844beeead93
z572177066719c137c1fc9abe2ef45c877f534191d7bbb5d90826f850c4f28a3d44134a538cb5ef
zb30f607714176b4e34fb2b1d4a72559818c26c65211749080ffda1ce059a58936c4d0aacf77eea
z5dc86e87381dd4f320c04834577494d76daa38f85b9a278b2e3eb60d3cfd10cc710c6b5a4ae90f
z83673c6bd96905ea5c3c49f0e506f75927b0fbecea7b4c92a2a5bff4d8f405cab6ff27f538aaba
z1610eca54dc3011c892f9f0429251173c0f51119dd8f234c6dc334f720705bab2d6d6c473be090
z099046d1002477ec11e73832ab6ca002e0c552564deef0feea0c8d135d28467e05d0c98545889f
z70b0356f603da6da171887eb801d88ba5bb6bbc28373f931d0598873c0ea46e0d79b854ac621a0
zdcf8782e67f4d5033f1e2fac6e79e47096a65e4fb85317ae0aa94c698fbfcf10ad8c2452d513a3
z2459be2bab0b9b32f03392d6d705ff3a387b10be898cd36dac3b8be28515691825acb3453d402f
ze9111fe38f9506919cf018515ed5c767c7ce2b37e1f67c79651be8e44bd115e41b16a0a20af8db
z87f8028ee4cd06d24d09aafa5585de6dd45676b6da7ecc75d0673d9cf771591b88d95a9931cd9f
z8bbaa1a1c9a162465eb8c28c42073295e346480f703b2eb6d84a6fbb03438995e7ef010500cf91
z0b8bd607e17336c7ce17823fbd34ff7ff6b86a8d575dd5dea5d230a5f0f2d4d74309f92d431f22
ze94b836dada933b1790af7ae5f8185286df5f6bd3292cdcf0eeef208c9db727de2a9addd1f772d
z350bb5e38ff2761651db40b73d190236699d3ffcd53f39a54acd8d8eed1fa04f48500d7860f32d
z109d344073babd355f24a69852a7f74fb43cbbb721a04614448208a9a7e85b523d82a0a4a4cf4c
z4c8d9ecf6b3422ad6998bf4500a75c2122df12d3738995a20360330e13767b9a2d6f907573d826
z7d72eed16cd31fe004a4404f10469cbea6903bfb46b6103bbd626395a7d531f7d266d9a0ec4ff8
zace2d19c224e92c9523b93a304cb2ff241799b9431fda2c5a5cad844283e137557fa77aacee811
zb0dc9633241f7245a85fa0a0925575a75de03b88c74878525a2623c4294051fffbe489d4f49f2f
z274a529bbbf5aa163467490216533dea24f2584ff101366b87cafffbc88327d3dad6ae5beef006
z01f0145bd7abb1820c9c13558ce7013eb6cc9a0a65756cb142957c13446228d62c98ddf24b497f
z17b3e49bdade1530bacc5a59b80a5beffaf1f581b6a6fdddd224050a25a200121435e9d29150f1
z1ff2f9679cc3a30fed97bff3b19ae9f4e7f4cd824dfde09e6f382e3309a53d8fbe8a0a3ea6a5dc
z00ba3bcd204863591182ee5f770efc20f7441bc86fb7c1dcdb327907e354114e650e932d76e66c
zfefb72c408c5093afa714858dd4fbb32afa2c099f17654ce71ad26fa1a7ea7e078575d98bd30f3
zb3835038e46b766657de7f99ecaf2c4b3a3de012b1171d6d436e3e151d3d7dc794301b119085a6
zbc737a6e325f6370cee2d07b4b6a0d848d500b4f306162d4cd07dfdcf7b5e4a07d3f5aad6b8baa
z74ea45d1f5c92a9901e172e939dacfe76b66ba2f584844c3f61d9e4850d46a40ba2dbd54d8865e
z3d94512045270367a02ad2266eb958004f98394848009a65e105b7e0efaa65d88bc46b79c75b7b
zc96049a43a99994a4c933af5f2de823a126526823cd1745acd7b1e8ae70e8206f6cecd45500d2f
ze1e285420c28d84e50dbb20bc44da3651b0158bf0505da509b10f9a9f71d590a0414cbfa4509ea
z67b05bf386b8a54142810d56ac1de7e47407b859d2b0c77f32d4b4366ab42c160c16849deea7b7
zd731ebf18d1a609f7121b79f83910420bd3920c39ba67b28bd10965075b2e404366876c4d52706
z6c1a12f0abead43af8ed6ed8aeed0330e8d42e6a1b16c6072a022ce492673d1ce1a12c8a46e8a2
z080308a8e5e7c402a81014c00d5e8f1a72b51dac40ffd18aa41224679e4be614f63f5e2323f9a3
z774a6744e98209ec98495e89fb00c7b3061176b985d37d9692e6d16e63d7e4edae7c777c2a5299
za69793b158fee5f50e5234c74c1b9179a28f0e053e0097d2e8a16408b54c95243325b675153642
zd2b9a27abee22018eecbd41588264aa1c6549473396edbbc1cfed0f0d60a808d4eee0d021891eb
zfb823cee71920fe93028fe1dc1ab950498fd4a8eed1d970b56c197def48572592b6b01ac1e4580
zb72e682719dda0126468579ebeb2df1a8325b06375cae206ae775d99ff4e0d9de6e7a0c67ebc82
ze8b7b415a491d79370893cddea240a2a6f31b298cc1808f72a940d60bb51ff8bdf6fc0f25d000f
z361e325fe46703ea2a63b1fe82608f5369766ff5ef9f46c05cc27fb681bc618467cf5f3257ff1c
z886121b917f8182ac64c3450dc51c35c997843880e7d7beadb73574d10ceaaba8f1d9ff057886f
z549a9dd77e59134997c8ce17450506c1a84dc30c4360843f80687a9a77491cfcca34d1465dd016
z1b76f778b1b31ca3fc357050bd0c7ed4162b06e8bbcf3d923585beff52aeaf915f97fd1ce1cb93
z986850883985532ff2b6f15bff458bf355cfd78f20ee3c03396618bbfa47656215be36542ca58a
z3e4105d1fec30e71044f4c41fd51aece2fb97b2802d91022292664631becf32b10736f5519c787
z6f64e7e00ffb2dbd6f9c9acd4e8cfadb4e304639844ba957d175d3ac34c8783da43cba899b8dab
z388bf1170f5c6d98de844edbb90ff737907cca38d6c10e93cc97dfdbd6792331ec640926385b21
za49824c0d10ddac4ede1a3b3f764a3b644b9f6a0c60c2442fdca89d79b164a5d7a8572c75ac7bf
z98fb27e5563939dbc98bba1c1567a29dbe566c1a90214b7103eed11b4d068d0d15c8878dcebbb7
z8af1dde13c6fc50b6f16d864ff4fa3499542603e1d0067f12b8b230863d553893bf82369969c59
z95a335735026e8bccce9ea38f322fd122d41c1e091177baf5c7e52b0226d93047c77d59e8edf88
z73b77c97b48ce3985c518d2398ba6724ab8a65d0465cc240809ddaf001e6aa0ee59276c12f4303
z4332e578ebe191c3b7b3ca43775bc25cddc50de1f0b36c567cc95f61399ae8a89246f4fe9b12fe
z26e72a78a2761ee14a9570155ce5ac3c897dd0315d74f217abca84ba2f81c5585511530c398c9c
z4d5add27fdb380f723548c1000872f8ad9dbc6731de802f08a10669dab75e6e70c0d31bdc33059
z9fed04c41b3dcef9e0c2f020e153441762e5639b7f2de7fc69181d9f8036b0e74cd93eb1d52528
zb02f86887dd73674b73837c78d12248eea1bf3f216e62fdef2d9a4bb0f34d71e2807a50083cb77
z19d5fdbd0fa28eb107f2ee0bc9cc5f88764b63f49f4e3d8d772fb6b8c22715ffead335ecc25cae
z918ce62d16a22bb3470a9cc39310431e8eafdc84c3e341a78f30c985d6c4c53167e74438ea70c9
zd555bb4d21992fca6cb024797e531c088cda27522adcacb25326b50e3b7f04aa820c589ea41967
z50cedccdf2001d585674f8419c960364565510b94e638d566a10b17a869138b120c3d9dce91d77
z8da423636fd0b3c51ab37f401d4816259dbc3b553471f2e0c17c64f59e6b8728d84d04d4658ac6
zb1599d1f0e124d1e07c5448877c35628b83734c5c1f14b461065e99c6c4a9d15f6e53a0410ab94
zbc109ce06071d9c09c19f50da89443e9fcafa460604ae419190623f890549eae8a5f90b53cf008
zacaf2e0b543494a00fa7c728521f0890a58187c9a2a8060125042f0493e16968142f8ede89db51
z9e2475cb37716f1df1ac99b4c8d1709bfea199043cc6ac5f454929765fcb17a783377f4c660b87
z65602a4590997236f58240cb3056c8fa70545a5ab0e3b5acfdb40294ac36d2865ffb5571a8a975
zec94298f1dee922cf9def443e5ed3e00020a01d38ff66fe77ff3d60573092a4bbd3f52194eb5bc
z8834ed706297f20fe556f6f8da72e8e72d6e86e26316be5ac80b926ed41467314370e530b3442c
z689ac68a6249445cad6c957c47e1ddb1584b75e489947e5a193eaef0f0b9e281b298bb5c349274
ze0ba1d27c2d9234d84c42ddd0ec7803bf3a696af2d13a5ae801280a0d866b595f8039e94824984
zc40273e6e03c6bdc5c91af8297b331beb5f35c42d77ca614caf81557ffb1c3943a6aea3bbef70e
za0ece5b2c9b1cdc2fcd6ad660bfeb58af13b0fd3d6b302f5d389191bb7b8c554c239a582095cbd
z3547a60eddc43acd441f521ad34fb0825f7891627fb7c2f52bfea30a9df287fb0adc5f7bd3efe7
zef70063f410f127dc10c88440e5a0e3bd6aef9d6867b9bad5f6e7e04a7fd1e1ef6fa1fcfedbd21
z5093dd4ec3ba244f2a43592b8de5dee8042cd8a64b8887d23b4410084c1bf12a60eb0320305746
z601c721b26781830f9b96468745f9dd656354e616db2b5819187a7d0980d4be12dad5771f37d6b
z9266d334caad6ee63cbaf52b4d8ed7bc92ed59ebcb262707f016e05e1e9516a7e31c8c25e3a6b3
zc7ef5c9dedd131853baf8d91bbc0bf66fc32b566932b50fe4445d0e524b15e72dac1b99b4fc030
zea42213a06431626deabba172aa9465b1617bfe07b817014a4706a0c02e27728e17fb68ae9f537
z81759a4535b743f5d4c22f3ba4c355a80bf19f893b2016441a210d59db47d72fa0e16a8f4b4be6
zefd5c0ddc1ba53826a651248438019420037e2ea44f7abe8a5a72245348491e424ebb106fb66f3
zf99799b3f083af0054b4c90c4ef646e08f8083964079f101fa620593eaa503be59b8f5f77e9ce9
z6ff3b48444e24d2f33f7bc4aa3e78f4b2cb1af3f1dc04e80620ca0d2c86da33d3406fd93c56924
z6dd032e6fa788f8c4e78fb9a3c0e5b250ba787c4b511771f30db5baf57c5e08d71ad79f554a038
z219eafc9039f80c451c88fb85ebda9cf6a7cdb609ff5b909989fb6171c5d76a7d9949e4a691103
zf8deb6e1ec139fac4d6791dcd017ea59b06673e40bb87d8380783dd0a7ecb8d3966cf0fd24f658
z397627e44e9239a18069ebd215bc952d5c7ef1efb03453363a0468797051522317e62f12431787
z5c503ed4457e5fca6451df699ecfec27546a5ea44643bf693114b462629ff49368da01ba249ac1
zd6b6f446c3aa82e2ae8d2ee40ab5e0d083237340721067a248f8a5a07ed2253c9900a55b18bd5d
z6999219c6b88ce2aec3bdc9802b202b0eb3c633ba680fa4a7c0dde0c399ed7b2569b22b26d6277
z67988e01f3b818454ef7e7955639d8d2c137d2cac2605e2f325d6ce155baa8849e2d95cc612a78
z843abdce03713968f4c6d72e57ce47d00c0c3a3886ff27c7fd6bb963221d514d002202f4838cc2
z5dccd929045c3c5da17bda896218ad1f8ab28d02fd67c98cb0853c15b755dbc33cea6ba9f84f78
z36e877fb0d67d38348311c65b45d0e432065fa25b832a8292391eb78110b0cc4de1a3d6ebf2958
z764aeaf9a9ade7994b249653095ac3a72d575f9da6c653429239ec78d787236c9f382ab95617ea
z3cc5b3e35c47350c404f42120b8397c6a1fe57c47cebfebf61a4feaca8d259b5e0ac4679fa4f91
z0729808a68316a46a96eb7d26f62724a16f0ed5ce8bfa91a7bdd7832af4d4620add9c43aa582c3
z050b2f08265da5358e3e08fb08eff101d51d985ca732cd3a94012b96ce750bfc32dc32b9255512
zc03323561cc8fbc5bdafcee55df51ae37ebfbf5f72127f3a65a5fd1fb17e09f3df59de60e9e54d
za30e21c06d7188afcc5b30c8ba3793f15ec5f689a8a67236abb570f6d94ab4d3da5362121d0f05
z5896f9a314ca03c190cd660c3b3be844c3d7823f106efe47900c8cf2126245337debee019e1b05
z91206ccc24aa7d2c3141566764bd581c98c147fc644e0f6c272a814673fad92d7ba44c2c146094
z14fda1c28fd5519a406784a19498406283fc255870424ec5d2be35ebcecbc115bd7eb83cba40fb
zb8f0356cb0d561fe467e75e188bc3c5a8fcf681c00983b72f8d5f0702f8895bc95fc21920b177c
z0968958840e5ee925dcc54e8fbbe4fc133e9607580658f231ab201b62a61200a984f08459c2765
z87fc2bfd5c51667ac55e0df2004a5a2a8eff0c132d54f9141f2b881315c22ff48bd435a8a17bdd
ze2376d7b61970a5afef93c1a0736becbca4d359988b63af7d48691cfebd5c48b996138ccab0622
ze36c4cb8df35bdaa2af66af9e19b8f823d34c3a0ff36e7acc65026f5a71a2d687fc172b8b1ed01
zc8b2c7524fcac3e2ce3cdcba386699741486ce34d856ec8bf41a5e0d3ba471970d00dc91e86a9f
ze1b0a55803917c28e9f7abf361d7df9ede9537d2259a58b1191680cafb649b2492f2296f6dad48
z9550693ebefd5fd090bc9786561d44772d3b7e44e20369c7a6d73a7658ea9f91a66c51822f119b
z26ce9fb15938b4de9f932eeabb930f17f5687936931492c1896b0c63def807990a61dffb40afaf
z76b2592668ce218e12c7b73e610f8150e865a572396a7e87fc5ed42500e69e291b58ac1975b3fc
zf51c208b780fafb481369fda76ddc66beb936276b5123704a8bf835fcd02c80868dd29bbf93812
z63b483b8157eac5981f0a84a074646776d872d3117ba516e146eeb81551d613ebff76a534b3acd
z744c872ac0e7d12b1961be6aa854f2f5a3da5ac2554e3d2839ec80487c1a61d357a627dacf2a36
z2f20c6cf09a68073817e3a2ded70e055fe94e70ff4662a20fe22474c31394a2c5f80bc2320a5b2
z7d7377e3b1f4210d84e1fc5d50d9551ab6564f3d7e1ac5c0002185aa5c05d30a53c10b4485d83a
z4df7d75f09c516c6fcd8a669d8ca9e02ef414b74eb3d3dd40727f07029342cca68b62007eac223
z4cd0035bb8bc43aea6d9f509d6ecfbeb9d6284f7c9f295762811eb403440f4bdcfe302af332fa2
z54d1332a0bd443c32cfad7f49deb58c60372090e90ba6d247e99f538876b1d0b0bdbc141afa3b8
z609a8759110bd2eaba3f51a5080c32060d8a4db27d5794ba5d5ff2a501c2aea1e8d5320bb3bae3
zab9a14d4e8610665bed1c3352c13dbd82cfda6237f61f9420b82549e65212d6f5dd32776eb2eb5
z58bb18e3f460de5649e75bed5512acf535cc86641e954ef7b5a15ecb7d4e6d5753a1f414e0053c
zb24db6d9faceb2b930b4d464d6dfbd3349009914b315f32717aa2ebb264e2f017d2dc90f6fd4a8
z836a61c296291d9342c2f332020aa86926afcd857e9df11080fd5663819f318e419d6b29c56462
zdf0a324463428b9c416d1423d3c33a32108577ae995d21b4c798fbb1bad30ab53ba0c5ff401593
z5992b90dd06f97e19b5d7b67631062e59ac20047b1c6049e85ebfa7f17e50e7033cb4d19e80040
zcf05c9fdb182351014809643ae87f68f5dcaa65d9510ca2bf9daff993c2187668819c671e79024
z65d5026d4ef30b5d63a477374718c061f2f86dc775933e348ce047b11b42596172252ffa00ee45
z54a4ff4404d8049dcd05f1ba3f9522622dd31c5731b7325d52f9197847de2bb4f4009772b6aab8
z435d5472f5a806edd75493e44619e64097e5feff6ba2272ffffb6466c0bdc5f8e75f3485929842
z7af94eebb49f61f22f94e05871e35fbff6acf9c8b187dc54bb2265daa94336d06f0e681d057871
z5a90c2cd164478181ffb59033e7afb1832e32a20601faebd28fe39313f1428c71db44a7ac3bb6a
z6652bfc36ec63c4f67d2c529478243b4b7967828752e47b1f331405444c1329ebb1462f18b26c6
zad4e4a46aeee0fce61a96a3e1bbe1fc0ef3ef550061034594995ed2f033e5254ff0ef8ebcf813f
za8c15138b495a671f44169999f276eeb94bb2b25b5a9ebe554d06b7709f84ee3fb085c6bd14a0a
z63ada130a12c1a0596cdde2f701768ca570088d6ad9c963dc9bd5fe76f9aa26a8cc6036d6a2c41
z61d62e133c4a8cece93a231ebbf288a5231b827090a65bb0b4e2a8f983a125849dd15f137d51e7
zfe94e87eeb17e7b83a3cd5f852fd4c6707c56dcea789e849ba924e4313cb39e7b8f1458bd59a9f
z03b6a2e7806cefdb529d46526efbc921509cb51d9267b2dbf6fcbefa851136eb3f6355cadd1a5a
zcabf5f59f6be4fa5af895f1c70020cc5b84c87a989ee4cb8aab2c6e1a9c74f79e778f293510a59
zfd055d62a2ccd0855b48ddc8fd50585096c55185557791f72f93a3238e76d268a508a72970e74a
z96086c5d77e27944f3d5a5a24c71063011681625aa5a505e4aeef3c55293d3110853c8eeaceaa1
z7b483aaa8cd27405a54ad941e06542f28a31047dbd5d2ab31cd28e4eaa3bfdc5e4c1d14cc8b9de
z40fbc48123720ce32a6fea84f90b72987a705c7b7056caff7bc794a37cec81579db6631ec5e0be
z1ff97357223dea1df81186abf48351b6fc028c1df2e2e453fb259179bef64e5c70c8eb3857df54
z796f11194de52fb88485eb65212c3353818208a4c18f0cf19918d51cd29d2bd28a01ece9afa0cc
z697decb456a42983258b65e2202c0bc6119325c7848e16d0cc74878d57dcffb8109977811c0998
z6d751df6fd6602ddfbe3c88b40f4df19e8bcc024de29bcd256099190ece55c6302e95c0d37e2a2
zd00c86e990be760841ab01600971a6b09197dfce8366aefd858692857bbe40a555ec7f0d39ea4a
zb3da43871ca41a3b986af27c1bb70ea21b1e3ff21a5106f93ab31573814e2cade4270cc47a8a9e
zb5ce439c696bbf7fa94f024eefbf264d04f86bd1a22724f39d6d0c90de2c3954bcd681b81aa051
z06a3a899ff0a7b69bd94da537cdafd3e66b3af0e59948d4188402a49f1c226df7dde4aab14f38a
z43a5e1384f3448a59c94a4ee6f6cd912bbb0778efb35a22f20015bb72b3854f3fb6445d8bb8379
z6e086ea8368d533360ab1a27409d02ba10da90d3ba7556e17c9196053d87a4c25cc8da33a42c3d
z7ffe63acf5e6263c567e70675cfe851497afe778fbc7cece9766175c9aefc0b11e0d6e75e2d031
z3bafa8aeb4f319b9056a5e9a4e0ddf59855099e777efd6eb8840c09378d769972dd128d71c4378
zbc2ffed8943538cf09d3615b9ac877bdc899e60fa2e042353f38ca54e628fbda6e001772612d6e
zd4d7fd20033888fc29f2c88bc2a1829a6509fca145f2e0a41d86f8b471485843c569d8992bab3f
z0f68b2ca874fbfbe219a6bd14910ab0232c9df61766ee48fbe7b376a6061df15ad63870a16dd59
zb40ccaf4d2015dbbb82ca1ede4433d995797ad64fd6d3c6a6d2fe9b84e44242b80433fea826986
zebbf910869ccb4a232a1af098b834aabea08271652c90c60fa1239b9ad3c7b966c349bc9ca628b
z4e65367fa0f1624802fd368cece0c6ee3e4977cb914748285f468d324146d93f9c17fa9342a8af
z1060507daaa8fd9cdca1da28ba7d47ddfde1f59de4e90e1e40f1e762908666569b16d1cd48a76f
z49b2d6e74d1a57eca5a70cd26d150ec04315efa2cfb39a98fe7bfccbb43a76ad9116f64fdcec10
z09d85038b99399226b17e30d8f18e99612cedb7ecb7d88e4934323e1739bcbaa3a3f2cad30c9e9
z3787bde11c6491929ca2facff971aea4fd14b55c17bf077077337eac730f97423f81fdeaeecc45
z114b465d6c4acb0919699099fad01fe3632363a024063ef54ec0d12af8736b3b656a805f16a480
za853dc4257d5851dd5d42ddf3e6718a19ad69e0a81e77beba331c8b8f5bc994692ebd236bb0bd2
z2b99056b18ad4cdfa461a209d861829e99e0048c2f94bda08d7480c0ed2d0bb1dce0e91145b6b9
z5cd7c86e4b9067434d285161250243a5091bf3ddcc32afa579eb782ce07007b16c80cb42e511c9
z39874f817ac5067a544bb19925b7cae1ba933057b7f1c06e9854406bb096ff34d06d6ee7e3a015
z0f7014ee46b8bce3218b439d436b33216b18711845283975182fdeb20978b8b36941b0d6ca4476
z39526d98aebc400d3337a73dd23921086ef7961de6761b67a09505136f021d5275d9a9f85871f0
zee045effc0e965678044a35a531d965b2ee4a9482687d6c6c875256977662dd8bc3f9ef8986507
za5c22ab7e3183bbe9e0a7530f8f469faa17bd2112c31488b7ec7e21d2729ac62e251577316bd4c
z6753a1ab6a4eff7e9b2acaa87b043f269ffbfe6a6d17436d948df115b42039e76c2bf0efddf98b
z823d9906e4b51adc2d8e7dd05c5dddaab81c0707e8e72fc42f03bb69205bbd1a171f7fc95ee240
z80e19149c8146a06457c84468ad4cc62315d13d1d7109650792777bfc7a61353850b8326e4d763
z055f2d65cbcc3222a7b3eaf84b5c01186a7007bbdd76f4c3ec6ce06e0ba0d1bd5ff6283343c4e2
zf100cb6a125023e55a25ee4696d88475896648678fdb93b3a2927b66e0b9f04d938055b1b39446
z7c33b305f909d2784bbd47d63d568715669f9849b366f3b4203941dedd759cb4d12b8211308235
zc2f85c3bb65f2f19e6fb930d50fb7428223f99b0256b18144130b70dcf774f8e9eaf2cdd382da9
z4497463c77a07d4860f5ffd75d8f3de5d1c115b2e27c449ee526e02be71a4aa4299fa33a25fedf
z1721756d7a526acf4f681d3ff8d6261213bd2af8bbe7555dd83d08f8af3fd99f604677ffdba0ea
z156eb3fd5bebf77dd517f6e6c2cc5488375293469f629c855e0145c88b41a9fcb46faa19ebf573
zf34af39a50bb5f0df0ca8e11f71c6c61917d4e7154599ee8b413863df5e2969b0c3fdadb9b8355
zc6a5a1f5b3849b46b5785716ffcb54738d9010c41ac9b3320bd688e87a9b5fec27caad548f8c01
z084f75cbb21b9d5cfbedd3606ffd501181624f5b8baac26851a31b1acd6ca12c672ee2eaf887ab
zb2c6ef2979a726eee209d35e27ac0efc4e536d6dbfd21397bdee66d161e04596eb48dc92075388
z0a13984bc574bbfc3f4078dd4ad6b7e8ead2d776cf13338334a05cb4e33093ec0f3e9cce2f9b75
zb7a38cb3ac8e1c93a5af6fb896cd3e4a347aab676f76591e1f3860cb1d004fde5c197f5dda4b91
z82e0c259a1e74ffffd8c95485c50bbaf840f8df323e3502a66c42acc4c6abf16990cdbc365dff5
z9cff79b2ad1ce3e0422a1958b378379fbb4b3851a80b6af06a7bddd5e67663efa18dbe8fcef4b8
z071a41db3eaa677e9bada544636c8994478a5ac12cece72869b151cfa89582bca39750293ae849
z524eb3cb83824d7828770da2e4ff30c9822eb7f7237467bd4a222b5026f20839d6a9e76f4d7ba3
z53ac97488e8bff30fdbfa5a9b266acaef790ad31c442dce685dbe5a7d29f8cd227b1aa0bcd3ce0
z82cd7617586759b2921d3180adfce248ee0b9f59afc4804d7a30ae3ebfba90fd2a4798c5c61dca
z3d99e3d11d78684edba7f382e46bd484d973eb62a049dc805612bb9ccccceee5bafbcafbad3bd0
z23b34fa346ab4b958b58ff2244f5720343a01d0dab6ffc7a190e75d1d0b301a91e78046f9a0f77
z57a02ce4885cb377184642b0d91143707259a0bad34430b726e5a92c3782ceb88064ea58829193
z27e9d84d732e188e8906be8a5b3c3af65c5e6971c77c86c7df8b921ec2bb11071bd6df964bbffd
z3bdc9bdeeb756534f34e94556c0f6350bfef0c78bddcb38e19d8431a3f069c149b0ce29ee606e1
zbb1f986f4ff096cea8dc5be653b06946c9f05633aa4d52ab8f5dd69de91aefc2c4b55553f4420e
z211870bdf904cc813d39312a206d4f3cc02fcb63db4b43988360ec93f191ec72ccbc5fc90dd79b
z92c59e03ee541f175f2eb3b8466f0fd39810c90d6d6644f9168298f7c4e0281328b989cd8963d2
zf37f846d6a7e377257e9525663ea12dcfb78b3feb97e47da0f47a5212dcdf455a9a9045fa17f5a
zd99869fec2936327a2370bed1e32faccf174516874814adbd07939726207cb0e99e5fd2bbac380
zc6c1ed1f71ec3f08cc0ffd3fe4aba3730cae46d594a0b8d2054e91f037cb11d72df4bf362b72b7
zb38da2cf8f731d26d9203c90e2c5f693b23135e520584a5be341e92f6790c472fb8846ae445d65
zb891053725e16c6aea3d5ba3d91deeaa86b7eaf1e295b2ce9d2b61ceed251b55fd51685d2838c0
z1abb5ef3cd450e4bdec743be252dd96400324203f5c076ef059a71710344e1000cd7c9136c9d2b
zd3ac57127a506e0ccf71571efe4dc36043afffea2ca0a769ae999b094dd058c93b4fa0679bb377
z5ae2c83a4100d4d3be9b6d590264ba07823f4babd3d22e88935a54ff476eee58df21544eb64546
zefdbb4424f5614d586690208fa4af68c9547837a05b4e66f5101bbc04a2acd988c8e002b91cbf3
zad76a3070e71261f2d0ebb2d626eadac0da28a4bb2a7d06d9aacacda0bd3a8824ab36091abd971
z2f68639d70d286a16a42e4e1e46aa1f61bf62f9685ab926c5a8c5e5dceaceeda42b82680453c79
z3d0e15734d9082088786641b8edc081a0b5eda7292630b31b7e581151f8e57dd66daa5d3915dd6
z06bcc5e21e3c118e2391bc6ceb45159d5a37ea8af973e5c76b60ca85989380334d5bda82b3dbfa
z33b0c17dcc99b03ba4d58b91447880f3590e78e360776fe4fe329bece0a57936e2ee2b2f5513b6
z82bf7b3c3d074445c96f623dea176e376965cc12ff77c4ede7e514e1ecedc11f63b166005801af
z2c999b54fd648bfa4803f3f84e9a88ebe74ea745d8f21254c9e77663b34e82ccd9934457cd2055
zc48e515bf2f6c27331927e565bdcfbadb46511bc4c60d6617fabf84dbfcbc13f5e67a1ae1c0537
z11331e06d90bfcf9cc4a767ff2435b497963d5134f1753bbd72af5ca2aaaf1f002591fd75b3e73
ze24b53e426e84caf4c1bd3c63538a1a87e58706b3f0d9a89d9e9a6d515344e8db07c67c98b778d
zcf95b83a58cfd7e52cb5df7249972e12527770780fb1209f87089460c3d06c4382a43ab39659a5
z6b000f40658fbfe0ca430f1181e7783c9a31e41720bab7baf72f9327f079ea78ab33b2170832ab
z046391e58587a45bdc3d46864e433365782a6d47cdede1b047e84ccb9fced2a4869315bf7cf334
zb819a5c96a7685ea05ab9c89a1d1fa92ae6d851da80dd93be73b7733afaeb8d1123addaa251a5a
z3114c23a4c9777d353f8b98fa4797ddf0204b5e9b5ad67845207ec1b1b09afb40fde9dcea6edc2
zdf43125219bc4add6c1ae17a887a7248be7fba9963b576833a25c3b08931c7026b4eb22e361152
zd2e621339bba8317bb2b7b8f2f0ccd0d764830cf13f4b3478a806c3d773b546730652494b20457
zd8349a529a72072fc1b623a75e55fbb1c01151591661673b2cf56221372d4aebc38b0563910069
ze34d44b968668d9df9d500096df1f15e7887bc532217d2b00a054f8776e471cbec059dcca283a6
z6a6c0268249dbcaf7c0b6d0d9f54ec77925b05ad65ae15c1b9c500a511ef202c9636b4f82e3ec3
z635724aab17d9238bfa74efa30ebab0d2e99e734b46a85ce897fbfd5b7bcddf2f5acfe3523225e
z2b53b899442b370956b906d47c01e35c768a32b548ddd6e9c28064511732bde5f9c9ec6774bddf
z558e7da254b256a8c91e802f884f37a6fc2a90a49f1aff3f78819fc641121fc5c1369e54d31d0e
z66681467ed6d52352a89b2cc7d0d46ee6f7e642796b5ba47791d9ea156a90ba96574a801709054
zb6a7fde9db884c471cebea0308fe8e67536c3ce0be5b2c4806bbea82ca750b32198d13b3d42a4e
z9ddd131a111405ca1ad0b97db6e04af2cac2837f78052cee7da557cd401580d795be750ddc0981
zf26617e159169c1301ade77ae77844b81ce88141e7b4aedd0446d54fae23e4d09f4e289c08b1b6
zbc4aac3ad5990d501bc04d5b418b11b793ba30a96a65bba97715bfb0a53bffdcf7c4ab482349f5
z6a7afaee273f4dfc2b720433c9732d4c1fbc528be3f3984eb3b8b0f2aad4ab80e1913a01d90344
z3fead97ec598b0da8125d9948dfe4ba2c51221706a7ffb9bef926f5dcfa8af92897e05335b76c6
zdf3a5782b8569f46f9c436ee3cd8d6bae64bfa05c7e6eed5075bbab23191b8930c01311c950601
zf699f2ccd71dd88e90cc220ed4403f5003a4338e027a54b4f386fd23425ab8dc8ec23958b68b11
z2488c179be216e4aa6d8a49fd145ee874f7da8635bcb9e12983da4b4ec466e50a81186bee45b2b
ze1bbc62ee6c856ac3a6c85c9b5f3b77fe6cd9be91e463af9dd3dfadb7f4e269f7c806cca4a8bbf
zc427275f5e2bf1ac36b3bdae570ffeaa1b44f620732b18ecff225c307617708641b90c4e8de843
zcc21dfe695938647c115103e7254fa98715f9e0e0722c9254be96877689fa5a6cb1e9162816f31
z559bccc1021425790d55f37453a457968d833956cafe71e5e5af0698f49b3abdd8db56b9b1c196
z2d48bccd670481e2046da6dced7879d2a24c6fb049b21224489a3c40a87600e3faf40a619007dd
z209a27b5ee214bf83d7fbd1d4132e855f3694c9afc570a58c0e284b5d7b17b651f1bd24a4d5e7d
z1bdd2c239e222631c74ed47f4888fa237b5b8a89c1af960ec3c8849cfaa2c9c6d27dcabdc32a37
zdc5d76e6e612316dea571b0a88d160e5831e38c9864c0ee464d0f2c64e5962734ccb9e2ed6b782
z76494e1a41a91d1d898fa1ba9dbe117b69b32bb63dc7a0e1d2aaf0b26a509a3a2c73cdc4fcdf32
zb951e6593859d7f79158acc1433ae781bec6bb3e0fbd5ae6c45f8c4633e4d89da58ac28e69c093
z71e4daf986a9d30b64404bdae60fe4c508c5a47e41a6b4391bfc3cd29dee6ab48aadd2b0c1018f
z76e0f354415e952fd0d3dc6b22ac02dce602d3503a5604a9463120f71ffc365fac478516dba3da
z9cf5f38fec1688bd871ff6191f978d08c3edf0a28c442dbaf2336ff173114dbdf6f20c63823838
zb97a6320a259d54627d73ebc1797dd49386970ff3a713f8ce4d798384da50c3858f9522a6deea5
zff72a20f926098827ec3f8e285cb8303385f0da6e6b53812fc102d3ea88f9ad1b787e6c30a38a0
z39f6b234ed0b79a939b544172370041783f3013657ceb4839dfdf1a151a4c36a63e38620ed299e
zeaea6de9d6f6c7c2da4c03324fc109f6a759b0b8763f20c1b5bacd32798e4ef3df7e708ae3326a
za2893b24043bb1cd0d70f70319d660e6fed31c3fbd378aa17e6b3d5037382246a7244fad2f2b5b
zbef59e2848fa801cd94e7c8409e6759f3fa6a5b0b2af01e11b8459ea7284a41f27d3555e5637c4
z85bbcbcdac57112f1274ff060c91497f8b1150f08c1d1bed0885b6afe0611812b257c46616e33d
z51e7013f64dd66e14515d069023504e974ba9032c0efca5a99e1bef268f8b8ede4d343565fcfbe
zade1798a591945d5a13d2d761cef6f248bf90b9448498c370db04d3a8947df588ecb2f5bc89d17
zd3ab04204aeb821a7e4c2ce111b5809938d518b5caf5ec04c481bd5a6918c5132a3376e61a41f5
z729224b3865f6b221a107dd59dcd30ddf1e215d1e84bf1822de7c65a9430b426059b378686d7bc
z0f49bb014ab28c4d7ca57387ea219c146bc3d99c60bcb3ec54b580aebb07bda80b22faa3a1635b
zf987625857ad659ae4d4db986fea2375a6900807e944db80b500fe741c74feb3cf1f88af150255
z161416e16ce97f320cd6258de800a31d2920533b32cb065d171252042fb19d9e8ac036fe4deb62
zfae5c801f7f7267a77756bb7efc14e5fbd0a4bbef86cf6cc722f736ec2928aa0266e58d7318a47
za2d135c68cca9b3cb91f6a0b223c47a0cefcd2c5871a4d97aabeb3a4ee496bdb6e82d0f32868b0
z26daa5aba1eb23b4ca639ea4601b6fa8dd5b789a2c03d68edc89112b192957de4674af8ef1ec0f
zeffbc075bae1667b932f1b054ac7220bb5ec5f94561d178c4a54b52c0e35f6479c413dd43383d1
z671a7b9b465ba48dbdb9f2a5915dd9fb14f6bad16bc330ab859d3b4f8f51037ed73fd0716454f9
zd9034bb2379a8e3a4f21ebc65f550b53a1b715e5e0974d3b404432013950e1da39a3be27232b7b
z418094b1bfa3df2ba9ab45996d876e4efbf35e44e54b5b8db580c1edc582a2416cb3b9185db9f9
z73e107c51cdf1f8689e9d59fbed0b238a46a30626004d0e3e4be492151a5da0b76894b01a6f032
z95ded7b9cc305504ef144adee419e4e75dc1aa02055cfae2ab09faa60e7299ca0f31c77f85be78
z2a8ec0b1de5caf11fb841a53fb964e4c7d87e8668608cf915ee874d3cc8aecaa3405e6946f4547
zbeba8dd22c9f9247b204f8211ced3d8b45d1646b4717385ad9c5eaec7c5423bc1e5490550cc940
ze62affa735013ed3d004eb9339c4589a8b5ffb8d187c67912062ce2d0ca6a025158fb28d30288b
z122ae756a1c85f261959e07f43ba2dd9eeaa17dfda57c1be184aa992354c31d2422c6fe215a7f8
z6a05ae2012f7f857fdf92ec4e9ec0108d7603c7a164e02442f22ca56c9be64c319f95b04b379c2
z6483f69ac7d80af44fc0a6cb029a9568656cc237525c23be3d3e44752126d1e789d213aae57118
z3ff9e46c70ae3f874a3f40fd52cddb878df353d1de12474965c369296f9ddc9a688527a27b6422
z0c0d1f2a5d9f5152b33291259b0981c65cf6cd227a5918ea135c0f9bafe3b8ed61cbc88880814d
z906c8b40353b577898473d9c6bd8aa0dab512b261648505a5eceffc4e077707c0016ba036cf693
z69fa8d96ba5c52d30c1f2547e9caef955716615694fdee6b8ec9cf62981e616d010d1ff808ad3e
z805902962b1b4f94f920eafdccad5ac1ffabbe773063ffbe9a8e8d2bee5f89b5cd60e1b88076d7
z73d9d600a1df29765662ffe4c23d55978bc8a95f55fcdf596e51bae636d59c4817154bacc9eabc
zfbad71d203ebc0ee787b65ba61a04e8b9b527e029876dd9f26cb56308545d53488788f5d331a9a
zc5a7d8c022a3c50db5cc2be6b87e99c049f3c8dcb4f2d04c3fe003eda226186779a5737592782a
zfe3a5cb8d4c7e63a4d58ab27b77504865b76206ac4ed71bc1cbf9f14c232e9cafe5682ed1709a6
z8812224215065059ee3ae20fe659e10a9aee665e774d04e2795b3d819c1fa91edb2ba8c47f937e
zdb1c5853a32d83f4e18dea2211e01f5eca3e7c599990c590cee514294e4056cabb1d083547017e
z047d604b9e5a520b2c47ee7bd06342939d7a602066f9dfa65015201f1d2e5881ec6e12fbc79aa2
z81f4cae1a5d1edf6429774bacc23cafd912cb7c162788dd7a494d8dc1d03db318d072aa20ba60b
z05c11e1d7634fb0743e93fc8ce00b32526c269dcb7101a14f04e3fda41ffc2e7c8285ede0393f8
zbfd4bca5b30c6d69adb9a7c8cf8a589a72fab3e1b071f09bdf491d8c763a786470053b8356f3ba
z9e67de23629bf4890c7274d9cb0056241657317294188b4acf4c300ed8443036a3eee215108457
z0c49a8c5413ca49fc5c2a296cc69d1120538bd7d19b8d0e544f99aeed3e29b7f75fb3bc123c5ff
zbab3a0055ffbf7a90edd8026a4a1dc4dea14d443320eeaaac4bda94897aaa26ee899d08f632a60
z3e88a988fad82917b05c4fc36183165595c002b61ed926d7e2fe3438590d43d5fa6299b9948acd
z374f921541cf24f91a8c76d502568ba139481efaa48b644484e524d46bdb94b92af1ab8a230ea8
z106808289ab188901f7a6151a4b1096a4a766ae46caf2d58c62e7bfc3228e47f78794e8581bab6
zb6665afe815d50ad13173785f503b19964f844de8259166b0ec75ce36c95204c9b030593b89fe7
za54bbc837233532bf8078929721a97ec7533172a0f5eeed1bdf529f3cf0ec9f7d6287eca5c9e0c
z1fc448b9da7dcf48693d207f9955bfe5f27c14a1a0fb36752dd3df35c23d2903b81daf97d690ca
zf83d6c32ada90bd2f32eb9880155aa1886ee5dd56aadccb098d2453b08e5b12d358c5f31cc9760
z0b21bfbf5368ab7808341416c06246b39333ce5689982a97ea01a18bd5acd9cadc5e6902d6421f
z2e5d535e1638a74a1e26c84780dca27a577aa6acfc0c9402b554e88dc02ee9a762d462082af451
zf4fcb2130658d50dacb22cd41f13c6f4008228b8e2acb0123f7f5d5f997f85d29ae30a539a274a
z8936c3a0ef0bfbdf18d78e95ee7d4360cd7e45f9954fedeaee346b8e0f852270daa3a3fae63b1c
z1faf607c9fc29251713f67d84a7bdf56e62a765fa6a07d46f86015f140261d4f3228e73e13027b
z19fd02adc5f2cdf312473a062fc68691ca87ce3f0fddc1663f14090c228548558cbccd7f8878ee
z5759ea0be79d5fd569f72d96761f106074c9120fc9ccf9e87bfbbc53f669eade5100ef21ae9cb1
z46bd11a3860cf4adb7e6bab02c67dfd2755ee5949b68b3c97fa4fa2f185e9bd7c6153f51813d16
zf030d44149bc8d3a43737c42e99e41eea52021c343d83cd59e1bd7361bac2bb018d534eea8090b
z8ac084d32d1749c695ba525aadd77a09dc44a33a0b86faee7e60902a6089ba812be5c9cc5f68b8
z997e381db8efc2c0a35c6a4fb5111d6af0d4f9064a8b46c62fa6770e27db6d2b55dbfec6306443
z0dfd521212a9ba517ce5be136bf334855e188de758327122ecbbf08ed43f64fba58548f2418945
z9ab0656ab79c834b6b71f72cf6a7f077d439443e6d42e0fafb4e21b8fbd0ada5abf0d6f59c7dc4
zb3390c27bbe39f9c7ce7598aa0ff8e2ff8c5f49305afaefb095b72fb41d95a735bf2378144469e
z955ad5bfb0b6016a3f13309703ab19011174eb1e01d0ff985ff8177c6b2a81fd81be3d8ebc494e
z0e4fbcd57776d190c3c53fc812eb02e59d0b583d4283a5e2602283a7d474466f364f49f97e74fc
zcd5ed2da43d540c865046663be5b2a0ba509e67e9770d1cf90cf494ae5f599b50a686794295113
z0392b7ddc804834d7a36a0cc33ae4a140f12134d5e5d8251b5cc7912a9c03d7a782b7d3669a166
zda46d7a652f37d3ace42517c8ebe07a571eeeb415d0fecd94d55cd2f6d37a3fefc353e05dac13e
zfce0f7497aa2c12b1510b1efa2d0b78cd7954935f8f79bec0ccde23f3314ebdd6f3170686ce99a
z277eabf47b7938901db205fb39ed3f2bb6258e92d72b62fe4d7bbc71d058e8ab14ebc967f176fb
z9e9872b849c1985102a0e36d8dceb11a156d2b18e51711c52a874e181a3e9c0746dd17a25fc37b
z94496cc4397a7d814ee53a0d266bf456461c27906d432d804fe608751a6892002dc22ddb62793d
z9f80e3d3680c401643c4b58db7df69606048079159c4e252cd2a2c403d4f4d1b2ce2a3daf75941
zba93ab063ec202b823c820a484b6376efae67a704b9e0e2c04b5c7eb9731fe89e0e3614647178b
ze9ed96485c14581058bf79370b8171c2be53a11b847e1817f801ef867c603964c64be8213f7139
zc776d32f40b66ad9c7d2969e2a563c16b411ef94eff620754831eedef47eec6af95786bcc52864
z4628b43cd279c9b6d2eacf117f4bffe89ddfcb9d35b45b31d1256767501f5ac3ef42d176a4f068
z67d651b6df39510677c4f7c64b42b3ada0dfad951c176e1b7bbee78d4b21b0ed64ba97657bccb4
z5541b503df29f3853922ce6525d6ea8704c5fc31070c03680343b345d1dfd30776d836774972cb
zec6ee2bf011553bc7c1a32f0e76311e004d0c12d19d273724ae3b651d99c3687c54467f1ba7307
z6ff09ba666e980f7ba5972bf1c46c88144f51fa05267489a41634d91951c619778ae84685274f1
z8e16b9881c1383e4c5c3d7a3dfbcb41006157f3ff6ebd6ebc648dac160d28b1c375bd9f402a93c
zd640c2552a2b2d837ab7bccc5cfc7781f195f6d1e7fd93ff8066d91550f31cddfd0cf27d6cac22
z53821a234793de5e34d52a13d21a09321742d027567b4fcebc414b4f320bc5058eda6040858257
z6922963b3204d78e2b9afb0b29a0f8d16c5cab6ae5a3cf8cbefe03829a6b86831e1ac3deef9362
z97f0be2a1b0161b279148ba920653186f96b3fd80c84c0b7e740a8b7449ec57b51344c1100649a
z7b5c622b92b6ec6d2dd86b8104eaffdc0cbb157c2f2cf7fa97da4fc917cd54d123c9a35df232bc
z0860f87d1e0b2bde5ecffc2bfe0e7efbadc5ad364880b9e4382abffd8e245cc69335279977f72b
z72b06830d9e2c6ec5e91651c115418f065dd6159b53d654fa2cb55bf2b0fa189f3a7494b9edcd4
z1ddc25cef30c9a738aa019184c554cf53e8a2859dac1b3647c2489610e4e5eb6b2d5353c7fb034
zf052e408e210e991464b9078201f6b8f264c8fd9f56e43c2f684e2548ad31f94e76de3ca6bed62
z3b8fca1f8dbac0fbe3b86fc5ebc27562ac6461adc78a2140c89a0f7f149712525f8fc92a128a65
z704dc1ff56b2e7881173ffc8d3f03afc8f57f007c587c2ea1992197f19eb4b0ccfeacc7c1bd69f
z9f3f9843b098e04b9d58167590c7aca61f36779aa044632fe50b882fc3df199f19555a31f3804a
z6bc5d1449f96e7d5b02d259ba823d90733686db9b22571896b73a1c07c66caaf1bb63414f5bd00
z59bbef6416ee845bd75021acc6b7b46b5770806ed47a370400531b5e85ffbc56b4b86912e9e1b9
z6c9ff049733ca62d08fce061247e480df5aafb2b10ebde1e7d40519cb1d554909776db7996eb65
z044fe98faf37d3d73b4e3de4552aa67e7ddfc19fddb0cca57d6a7af5f8dab3d187670ebb3dca30
z6cc2f0ae1318d6d0dc2f3c8f49fb69cdb8b9495cbb17d4c1c0fcd9a516ef24041ff19bd28c1547
z7aecc1466fedfe106fc226f5aa1160abc80090a09a89a8c406d9dae4428e303b2e6d49683dbc84
ze50b49a91f88012adf971676c7313faad0bdaf9daa1220af8f5a9f82c976cb45d700bcb50798b4
zfb71a36036c188ee5cdb4e830b467047feccd0695e93b0057237de34fb173c73ccad829ed4d763
z17e6175c962130b0d087bb5de42a1723da37b505df07d0ca4b1f8404105d5285cf821391e1864c
zea6e82df1f8ba016aa71662c3b95d6d95da34c9fd08196bee97880f9590146a212649d24ed9939
z09120606c34f878e3a12931948c340528c4c82eb23b3561dd45a1ffe9e458afc7f46d76a288490
zaf71e30bec59e8c9d7698c2ce8acaa307486fefa4df1707617700af2c788ec8f2065cc9eb93ebd
z45b1674048c6e98fd5da94259e58236ab63a8284f87682c7e48f07d5ff7c880c0683b0a9378d98
z26720ccc1aa207a735d15d29f5ab31ff18e01ba6ce173b98cc1ba3579babd1fa7928d72663c1e6
zde2caf22147ec71516c6f794c5b9787f0b5e1e5ea2cf6dc9c9805aad5fdbb680ac539acf6c0972
z4d772bb5b32b35468156552cf95a45462bad3dbf6b107459b5a91fdd741676277359b30f85a3da
zb70e620e82ab6dc9b3a4a1b18674eff47827054f93de7906f08e758a636e7d955e2a425b1e0490
z90b5590e919d8cd0edf29eacd0a58cf696676ae8498428eaf5e80cbf7f9c4fc24dd1b5bdf36495
zfe4f75b1df2d4ea3e11043914c9c7f0bd96420a8f2883dca88786cabf9c47dccceced2d46eea1e
z6c02c0ceb6937a309410a97527fc9326e6869fadca4188ffc5efe8f98697b850be1c6846f16c82
za3ec892ff832135adf3624c2d424d318ae29f9fd0b1144e658cecd58b10bfa2d74618df53c1669
ze8343e3c55fa0d3fba37a5a4c7f1c5f52a79c665e0b84781b875bc47070bc3d475392c86d65b4e
za7615e63fcb4be8c3616195530ae6a04cdbe3afdfee21f7e0f0b46ef45215df88f1c4777ecdf8f
z365f0b50d8514d17e66cb6cb8bf899f4a2c97543c3c8162b8f9fd2ad346d014528fd1782e9ec01
zdf4c1cf9752107b82f7104a0b4c7e08a9931c695e7213045da1682a859af12d75fcce57d7a9759
z541e06a3f6581f191fb5671956f898d956a19246f8281dc31643b2fe532f4da68abdca0436c945
ze007931cfafcbc31f74e9d7e9080627e3fa1e1b6bfa1086d68720dfeeb4dba919c2bb3cade22be
ze8077ccb28f17ca53aa85471848d42d5095e65b4043f592f0a77c73fc2ab78c280425acfc2152f
z2f48ebc8c065c2e29d3c198db5f33161203a3d4ee3d42ab89d7d584bc682aaf77882e165660f40
zbe38d443825350249acacf42adc4afcedf2dc388cecb2d5bd99e6c2d1b843c3b6405310b0c346c
z803e291f2e333b16305b53dad12e45ff5d55932b385c15f154cfafae47f2c899f1e50b95ac9034
z815042de2443ac9fb908e3753d83ec7d474e8ec3169189768ab653dbb3a41a4351021956bf7f92
z437a208d571302a54106598c0b5395bcbae8c69ed594713ffa8097318059f14e6da356be20febf
z1796de928b901384047b1f14ee4cd6c5f5ea482f05a6ad5a0032c02893d2c625b855509eec98eb
z560f2e76c9a5c61d946cc602852afebb52238ed34367916ee94c3f28a71a9877ca47f9b1cd24d0
zfaa82c13a039d52ff1d124e474fc7b25af6e5ec0ead1daa9471ae4212260cd2e72de67965fdbec
zdf5fc0ef940446a138f51f929841bdc692fd1cc4f50109928c6409d067e91fcce94dc966df1155
z442b72f149cd73df75e4aa03e5009f6e260d170574f89570171989ef73182c6939aeb43f73acef
ze6959aac40232705a3b9518cf1c74760030cd74687e48530522d17800f43b6e8fa038ee5e495de
z5af7d8008298f87a679811fa12aa1673c31af9b362814f9a57a1a95e58cf6c04d08e75c438fff0
zb8011cafea318071a35f52b08b1bd4d5f4e54136835b274268bbb975d1efeb4ce33188fdf5c8af
zc545a52dd95bf67f4115bfd7d28d91a67cde67bff4075f07e128b60ed115a0f9fa89af4878f639
z1f29f441da24a92db084db6730f8287e90992d6ef035a1183049012b379fa445965a9f51157cac
z0fc08efc4705c391a8dc4d10bb99927b3b1faf7ce257cc065eec9b4f3fd55e069585044b27a97b
zce8fa5d7f2bc16c2d98c99ad4e2d96770cea27816026c2ae0a3f85726855214edf526c97e67040
zfa42abde613d4c724aa8d2049f0d2459d517915dd90a6c5674a8b44d145fd6964173686ee9c2ec
za1bdf0bbb88bed82ebdcad5768b11e77961dbb4abf02349cc9c117af5c505f67d9a89c646ee179
z8ed6c87c67dcd3d5c1406cbb4d7ea4039f888d948210e8475f6ddedc25d052de635e5103b21bda
z29d2bf99860f50cbcd5a1a118a424acfa27af44484814b84ddd55d790a30722ff2b8912f3906eb
z0216acff65cadc9508cf793eb9e3daab04866881b01c803ef517683c093d8a8f92fd5105899cf2
ze0573320b23b84bc888015f4d1897681924fc3d2b4471d87f545b75520e79bb0cd27ac1ce3fe41
zed982572fd77b96b1c8374d838ab31a40313192444d03ac0137db9a19c5a25e5735e5486783221
z5b821d440ef217585d41f70e7d26c7cf8676e0a807ba9cddcf3ea943d6ad5b2479fd1cc3cc86ab
z8853928122a6f02effca92babe546a2e46263439f3bed5f50db5c0f030ae4eab290d107dd5ca00
zc327e585de6eb3705b02545781764ac7c15cc832fde14fc465ccdd708d1a6cf0195846a600650f
zbff718fc30f161a54f9b550eb4994c949eb60bbacf5bc54417d0c500c25d5c95bef3dc2e29ff26
z8bf1994fc040ecfa4be9547026f097b0ad481907f9be55d7f9dbe273549b7346be247756c27239
z77421a73e1fbd88fca126d254c270dccebabc9c3985ba35db4e8294f366391cae5d404e94e39e8
z60d50aa66d2f10d41f7974b9effe3b5d173e0c0f5cc868d93dcf613b0c30875b704f7a10be304f
zba026c75097688d75e03b841ab1a1182e9a784ddc82646a714bd4b175fca29a893f3f1ee3523c3
z4c10f2f8f3d29812f6c54dbfdad4987a7f36ae206da2a1bafcec2cedade0a1c616d0bfb59ed34d
za389988f00c5ce3a8ce0c8b3ea0ec6955423f73d15acaa0cb591eb9448a8b934ae418d39c73693
z48a7f8bc5de1c67ef000c1c472ce45075931b357def7aa1c4417c97bed199f3c669cba2bfc6505
z497e14ad2e61d5488e173a10d1becdc59c4e28428fa52d7b9439d529febaba78f1afb917dbf7e1
z09555d776733f5ac2479b081eb0c3bb8560e37a2e0f6ba330dea703028bbcc52b4beb6b0513779
zaca55f7630f330fb53285dd143ca463f78f1905cd6161303fa4336b47c4bff46cfdd07fcbdba23
zde8d49a8f47f671b2097739a0edbf334042631c17b272a2388c045b000000ec3d273b8a26eeea1
zd4f0870b18f642ad32a2bdf016ff38be50e2ae4bd491c1f336e25af12971bd7735f984cb424162
z7844b9666270fc157232f01bba97d055c0d7cf6f917fe870a8a4d09b628981a5ae999b42705f8c
z3b61dcb408b7f363a5822543e19a1b087d8968f2d9686236a958487ae9dd6cce5770d329e3e668
z6d3ef7e50c55f6534f28314678d7ecf68d076930bc6457915aae652645810875ade0599697fe8b
zfd36dda5b04ee5b5010f21dc641ab5c64d4dbd4312dce8a682b1ff880b829d81e935f266ba1c0f
ze254540851e6e24ee36729f791b08c765d9534233a6a79f6099bc0c031378be388b15eaea7c6bd
z925c4d01bed7ee94c169827c9884ebf4b1069c465fc8695628c6b4448a62a8dc2a95002439b5a9
ze4242cf39ea594e59894d7046a1c4928ba71531cb582856ac06a80747f0975ac75adb73a56b6dc
zf256f0e0dab4c10e7619340e2d5afb3797909a8197b003f7ea180549e8a155488469a3f924bfa4
z8154be12625fd8ea59b85753a826726a5b6825b5fe52036057b5b35c3603e86a1d75060f1d41a9
z27eb024dae85cad3a1e7e1b743824e9d7cdd656245ee4280e4b49fc95b0681541bd4b68a1f1081
z62e7f1de63261bcb66981358fc401d1cef55e5b15a9b60285cef33ed04e03adcee41241b597105
zac53dca88312cb0bb1ed2a0b53f6f690a9af658a4d5789a690ccb8a44d25eb100b4824eb14c037
zb3249b779dfadc04a8a475cb92a4ffa3419c46c8c797e263960a7468ef547b71d94f0949769a7d
z37a6a755ada2982578c6cee32faf1c6a8646e4f3a98f1802b02244e826a518efd154b0dbbc52f6
zf8ea0393f745548d4ce0de48e7cff599bc76e49a025d14b9a85576fdea19bd8304d4a07402c2df
zcfad399ff79a91d6b4081a6ea0c00865e9aa8a80b14ea4832fc3c5413faf061a52777321477a70
z3fb886385a49602683278a71fb7a779a4572c15dae3641018459c9936d78ecb253ff8343a22043
z8975118d2bb6c962582f7b29ab86ae03e9f79111e9284a55b9ba369afeb7f3d29e8b845e670beb
z9b286a64cbb15202bf38007110d47d6a01ab6ed985d8a303c8d9e1d1609bdf4a6410391f4656fd
zfc9493089143e4555b0644ec616d61becbc25a118a33ef5a3e222870732e068d07e8da534cc6f8
z57f3567a8a1a80afded5000e0f008ed8f0a1b7f70de436a8aa4648bc722d9fa25898f6334c0d61
z22203cdb515423995c213eb32eaed2b253d8110e445a1dd86570008995e2b899deb5f34e15eab2
zcce0f16df3beac021c0a729a7e2e64895554f794d12a5c5c6faf481bbff398abb09394472508ac
ze469399a83f53650e0cc30436d9771c5dba671bd4e8e65f4fd32a749e55874f9db20ef1b596974
z7217dd72276f287b9bf2a55093c3bbbf0ce57d22785dafa97794ce009a7256d1049be5a380230c
z9a5bdd4493b4a427e0fb50ced2f3b924fd228595ad63798fcabb91da946ecb763e9a202febe108
z4658feac35ad21694ebf7cd4e8321b662fa450a9c96cbff8030ea0a478e9fbb854100bd48a3fca
z86110f455e07444daaa525558b7aadb849cf4cd542c952e3700418c7e31dac352c5b6142881e03
z5a1c83d099fb97f6fbaa989f1b970cf7b730d45404dcc3b6c94b8137838e90e98aea69198dcd98
zafe07ec380de40873dceab5f113596ad1739ea5c737573144cf44cbcbfa0cadf0cecf352c3bf0a
z3fe46b48a60f339ff372933fa9a015f10cdfd7b10e08502c92faf83f26cbf74f40dc009696d6f0
z5ecad8e055e81312efe65f418d0b7a945d60c3ca1629feddd71a279c97785fc84ae2d9a7f95af8
zbd1319c4d49523727ba7dbb64a6761f5e2fbffb394bf7624477e674466a59586aa1f86e062d5b8
z0420b3eb79024372327600cf3683a60bfa7eafef493fef008cd72d0eff155522a91548aa5a24ad
z59611c5678875eb21a35857e71886e5e33f93b8b867218db3a17b58b738e86e8b7c0a66b240798
z20ed6c940386ae2cdb4609b114e72481325a9f6af483094f06b0da5ee43b14f792cafc134dc7da
z42d87bad2ba3a703e7eb1f52abb9fd47c9d29efa08ec38ef7c6042dccb495d4b501cf9a2c6a641
z3edb843759d7b113ff23ba1dc5c137e7235ac70af9903e4a223bcc8fdb19cb4132e5ff79661a9f
z4867007beed8a9579eedd8b9cdb8f0e9ca88bc1bd6d9ef3fc21b9a072bb49a44c13eb1c3e54c94
zcdb124d15d27de547136a6b22e235b0721262272144a0768bfb8a01d92f9b0f8792223ee61d437
zccaaa7b7fb77da464dfe2c5e75a37b6c562360a78e843ff6d29207fdfb0d163bfcca3eabc93260
z25b8175cbbd216bcded29be07190745d9b7693ed2df196a58a2268bec77d903993f7c8b4dec44b
z649608734628e1621c892b5d3ef76059e8f8182cdc41ef91855cdb8a64fcf3d7032722f5aa8b80
z3bafe2ad17fc2e64079122c7e80a61b2561d4a3289cf1874b18aa1bb1df992e71fac0f18d7cf05
zfc7e79b26c78e230a9297e43f9be4508a35bf795a48b1fd80b30e71b85c3ba487057959cc14214
z4e996f74df711a594d5f0d75b2f0ece7f49b7d5e7b7e37b7a65191611989b05a66b1e9b28a32a5
z50137016111f9b6ff31565fcef4cd9528951f64c2d81fc63ed03ee9a178223ec55c8afc42c820a
z8e8f844e53e12aceba60e7021f613542d8a0d0e9501de6757b6e67d415a28b0481180edd181c61
z02dc6d5d82f58afdf13817d3688989885b1644c9a888fa9161fd1d6a9debb969d4e56cd1a6ac81
z8d223506feb2d25774a2aacaaa061af16b2a6e7d4b5b9fe6050f0a8da00aef7d1e7c09615889aa
za23f50a44cfbe0d09e54ebac7f3d5e45fa2317c8de59beae56260c804d95d9e77e3273a4fb5adb
z3b4236a2d074771d039ae191c09cb5e7d3dcf60c6d4200a0b2b07b78a4aee6830a139ad6ebb42a
z3c776aad170025763039a7363ca3f4e470a2b034172e480265cffddd4b261daa314952c189aec4
z3ba0cbf5362f082313312454b15acd8190d16da4b5ff161cc1ba7965cff03aef79fb77bbfff0cc
zd59dce9a046335ee877c92348f01a110bf0bbffd229b0313e57c4d90de0eff5dfa68a98770837d
z1ee2e424af385fbe149fe1b4dc2a67e36fcab93d55f465207dabdd7687e0f6808121306f4a8dbc
z9c5f117ae5c997acfbbc87b944e1c7c7acf7b0ce6c9bf980931ba3d1e5119a5ef05aa67bd52d51
zb8400428b58b6676900f2f950169e096a155dcbf841f076dbdf902b6b9a4fe0d2e96850e14e8e9
z96b9cf9e0e796c312fd80b876a2093b1341bd2536f042c0888159bda46ad44b1fe4734e5c63411
z5a369e938bf57e8e746bbfb6201aa604a440773bf87e7dad2e2871ecfc68ffe9d963e744b5e9a3
z249d590dfbb496e97c4600e94b2e9c5a62d6258324d12f3ffbf1da50265d570b96ff4a69a91f5b
z383ef22ed8de8dc6d06e150e00e476cef0ac565511a1a88fc3e3365b07988bda03e1ff45ea7d60
z41ce1c1c92c172c94e5c7e32d8b7b5dd61e9db0616fba20c2c8e25ff3cfaa0c869d18ba4efed20
z5d5eade2066af909b62057a78a2ded43558601962c468b1933245f163bfe2250aca26c5673ebd3
z4a28c1a0b46f4439371201d97b6b4b39269c9d2a32dc3391703abaa5a1d70ca5a158c4ce96dd29
z52b573d828c1fababed7be149b30a270ec1c03731979be2f3db1b9fef9bdf6adba5e8b804496db
z88693061e6238dc60681a914a60592eadb09c31d04efb5d9cbfb0589bdb50ec7d0afacc3173056
z93658194bb2ede6208341a2b34e0e111aaa6e568733b3c0bec45efcb534a0d1cad1df580dda220
z931ebac8c05a763c97be3588ae9159e1c9da2df3e30d8ba3cee19227d13a11bb4105c19674793f
z49d297493cdbe743f63ffb968183f9ea5bf8fa864f294a3e37f15ce17f9bd9c78524c800ee1d4a
z99ff06cc29b1498bca916f4a22703aaa5b39e52413bba7bc009efae8504bd7718615ea0f5fc2ff
ze41f34b26e0f89aa870251c099a8207a9ad9e92f8c54a2ebae1dce5e60a5fed8c368499e79212e
zbfe89a97e58e9828e1e3869612ecd860118f161b7f2b1a3f90398e6e06305b2d0653d151243ec9
zd7cde8b3ddb92f9f7a6186342247eba0f409f38983233027738cde5a3c7852db8b4505315873f1
z79f4d390b2cf467ac626bfb762426e7403d428ed5799bf3d071ecfe0eb46fad49fc3524c3512b3
zb11bab1fb11c3f5fc5846e8672a0e284a1ef54b1bb449de5a06a3130b89557d8cebe6d6d283340
z49659b427732e414c357150b56f5a0824db5a9dc3b9f7b4b6e254877f4e29436bef22c783aab9f
z2bf3e3a10dd53f828bbb6600377161b2e9afa6cff68b31a9bd8307ecb879f925b997f1e66e350f
zc32a62bad64ce4f2951eec2ea780b3bff921ed3e588b89f6eeb3a33db7c55a4b070cc21f8ca538
z5b95d496f4042c2ebab032dd113c7f1876570596aaf6d2387342da7dcba06a684a3d911cefce1d
z6c5bd2e8daee7e5a3aae620027376bc32e43f3e99a9e4f8d9096ce2b9ea14b58e5cfbb7379d155
zd9c0ff9acd9713963e4c4e94c62a9605ad7704fb39748483b240361b14389b3a7670672cf9c0c4
z64cae53274c470066ab9655815fe2a25f64fcc8a1bd5d09a5e8f2647cde3e374fed017586726d9
za99c0b08298439c81cbd1ecf6904394eb757ece1a08f16e9361e6d85595f80cd69399aebdff2f4
zf0664b2779a875597f41ad709eae6888c2f2624f95537ccf1c2e984d629dcf5527c87cad04e37a
za7759ffcadb8d692d0eada7e9d1a1c42ff16c71c78341ef0a6211c96e6556c27fa04e8c6ce953a
zf2d68c915e00ed973062d4ec5d5a2e30876cbd4887afdd8a13c81fea2a8e4bac2e3ff65efbffa5
z684f838403c79188cda565e452807937078cfeec86c54fe96e697a4f57075025d83ec6eeeb9eab
zb934633ec755ad0f9e38e0edfe10754dda2bd9c83bced034d5a8e2e5e9d04c6fb63eba0ca01029
z1a6c9516974aa00bff863e108267b7c0efe579c0db54533d31524c1b4bc6e41da91bd71e15c955
zbb3c7552cb3d144db81f88cc5ffe881dc03ba5ed210284e0323338503ab5e9686f68a4bed82e15
zf38bcc27bdc66259e07d011a7294a7ab8ff7d7e505e9bef3ce0e34a2f40c56c68cef22fb68d1cd
zfe268c7a745f27de08f6af3b18c3d76ea0cac64ec4cd85a913f5c504901f104a8c22c800818b4f
z647dfdfa6c5bc1fb4bc16200e0b72298c64cf2c53b0361cc1598290681871631bc6c7346d73b15
z586d6e62d230f6adec4f057ebfce4b2d3fe2585708936bf4ef1e41bc8e822d85d1b06a9a24d9e1
z1ff50f684baee6c2f1fce4f985afb85f3b9bea0e786cfbcadfb4fca3649dcba491e85ae1843a43
z4cfc9da7cce566172b46d476e3857c52945b1ab1c17ba7a21c5667991ae9cc5b5103c114aa5720
z7423bd8f5ff22481795767b3b13da4dc32474fd5a87322e7f39c09fa4cbf12762420718af72ed7
zc5d042ad79e2ad1fb1f95a4d1b50c5de3476090d125434dcdaeacd82ddb3edda383f52f738ba5b
zd75c97b02880b6fad105569b61ea9ee740dfa42e42a0265cf9e49c9a4b943013c275fefcbc2bb0
zb9d13d431d59d4855405e14aad641d12bff2182ce9373eb3d6f1f8e92b8f99e96bc2813759c2a8
z55118ca1ed7fe193250ca87e6963eb2b278a589fb0dba0245aef73deb5bd358c2eb7d5e00f8bb1
zbe71b3ee96d2c7daad74266f43b4e054254d25930224314f0b88f4a1ebd4463ce51b9c57b88a0f
z2499d9e0ad25113b02c0922a16e6f2048cc6ffba17a9710e5ef1d536220f1817131c08b8fd36b1
zb96e9182164acc77f7e1041c35fe14aa82d0b6a5125ee0c71f3e45ff383b8e9c944020cd9714e4
zda31889f9648bdac19e462682c3f95ee82b439c4fb032c324dee6e1ca74fe37039ef97d71d6492
z4913631d306e2951f7fba161d4396950f8adfc144eff2b2e840b5ca7d179a2ca5f3624145c16a6
z1ae4b6f398e6e6edac6a912cc1ce3e39cf726591dcdb9c9505d50c8ac1b0e452cfc35400ee0c91
z72fd78984ff6eb1a20149e230fc40c9ae78aa2ae9e7f0a5999345dd29577fd8db75252ab5e3159
z67a93ffa3755b7f30de0089647591f226b85c57baddd907c90b27bf8c360e3e03ef7983d391b21
z6ac2b5ea6836907fe20eac6059e61d6291a837906b7c8470ca94e76f19380ef31bf2f979ec5b2c
z5fb78a290c325903e76d47e91e39c4684e07107ec2876206be40db85b6da56626d99d8f11f2410
zb0b5fdfed9fb4b8790bb42cadf76bc789ad117e04a98c437f767a7a69e71beb48f43b8955707fa
z1e7efd3074eb1534b3140760b3cabbc6a403d51d64e049a9e0b3ec4c7b3ab6849efdd05cc4f5f5
z252551a9873ada99b761db5491682118f7d7fa368984b9a21c48142ae3ff9eacad4659fc82da07
z625cf173118efcb31928f3b8530f0394a7896e7b6ba1fa22cd08b2de1456783ce11615731a0900
zcec969d7a139de27b3324956f20ee05c7dd0bd47b6141cc004ae83a242519820ee1933f789328f
za1624ef3b99676f441da3dea935a545314df732e076db5f768db25ecb5f1778178346735bb3918
zca88e2687cb78a8c12e508b6efc6d169361e01b058ee13a07ae263038e9396e14bc62f08be7299
z3ad8a31b04796686605643c73e06e89531b63f6275228be8097b87d5f862b73b0046385226cea2
z2c66e4201d2092878e2f64f658b51ecd4efa30adb38a9c5d7db93d69760e5f9a6d0e7bcd3a85f8
zd24883cb15971bf272f959bce7cff7c4db5d4b6dc7ad320629b020f06862df545f9dd1850ec69d
ze9f876a1a53109cf4ae77bfaf941d82f7cd5017d0f30608330995e1e2a5f2d3aa27c9abbf5033b
zd6b8647911facc886721575c512369aa1f4fdc48d17f577b35581dc9d79dea0a7fea3d97db8134
z19122ec41db55bf4ddd498cf24b14257a33660539e74a370ca52ec570f4f837e5a76e81f1e389c
z0a8701e47462890d2131a0e49f69fb32013841af1d2cecdac3e771c29f4cf9006ccd3091926d4a
z3a65556859a5034f428d964cc13db355e6792adf8c4adae463be7c3549a16eb804285fe7ead2dd
z835688485a6c893e307dce0ce47d8ab55b37257c4b77f15892886ab036ac08fc00e10052b509e1
z1a8eba1eea33e30de7c4e939a8ca2bd123ca6fc2e0f11a5d0139cd94bf04b722d3a964f939156d
z049e74382d699556b0950d3635a2a4ab8e4d9c007c6f1018ec0f1752495504bd61bb057298ea49
z1b98181072846a34e53f29473faa9a59b8583b25aa2e73f90a60a76645733ab55a2f0364eec34d
z596ad92c86c6793d2445b6f316489c0b413d621bab0d8e55034346702d7b35fc7643c93c05e893
z9acbbfbbf89560662bbaf3b42fba8310bc031c35fedbbfe22c5a818b52bdd36cf24dce119eac57
zf5f3344760cf9df0887df382c74bb77b6f683d7375b6c0a5292e664b5e4a37be6c737f08f9f966
zcef470663885f9de5be3a81ba11ef0dee90a403789e736eefdeb1c00f26e919c0c898c05db75e5
z09ae3f3619c0d4992c2ad7fdc8647b60e1d5ed057d185736c403628e0e706dd17b6c90f9f5806d
zc31ed7b81d91da39181ec9eb34f1eb55f3ed1bc371e2c6d86ed1a12fc87298a04d517c4dd5fa70
z34ed22b686a0e8629690c41c32bd7978cac39561140f7a00de98fb6d064e62a6ca6bbaba80971d
z97253898a734fa66383f97cf586ecb902ddec2806434c629546075c3ec154328609b108634f936
zb0ee8ff7410f134e13a531915de2e7e653dd53fde5932ed9c7f39ce7b4ebfcfa5edd66c920e45d
zff594c14c8a57eaa294e785087506e9d18562da1134bfccb78263551b0528b5940b00c1649e458
z1b3ab53ab16d5f29296c940b0288c944088ca4c213a6acfd3ec88d9852436ea0bd1c2b22bc1bb4
z5ffbdf54b6a8161db28a0a542779f0b3f2b447ac3ed075189001db0fe7c3659d66fcec2af36a50
z4aadcb5fd53f0224da5171189925829705e5353039b173108f01626cb33f7a080830c3976090ad
zeb7e749eedf1bdaf291e8174ba84b81b29d23a7ae7d37a3ffb74ede0aeb35904f6075801857316
z7196a83d00f1e2d7838324a6f83bba5ee4a283a9922e172ebf13589ac797d4729aaa785207293b
za81e1fcdea7e06a0a5d9b9c37247b3166520996a3abcf5c67b7313e1a68f1eceec91a5c21efd05
zee249a01a6790698470e15120774b96ef86b7ea6c466321848ceba0c0e0e107c28cf763d6910fe
z1f9f472b22a50c26c7d69483075aebe88d53b741a569ef99ccf4e95fc6bd98810e25c8f746da4e
z1fec9f183d5c3020e5a0d6ddf4e5bcbc2fc430d78c26bbfac0e0e3d331de7bb9f8d7e7772445ab
z8478985f288c7c9e2b64553aaaf032319e839fdb9608c1da1c19609d1b1808f11aa9db919dd053
z43363252c814014b4cf0807c5668b4da70cab53a463de17310c9010d2d187441523d8a5a49574a
z6fc85b66da9495264c7e0579ce7ffcc63b9ceb587021a7cb7a3ca033dedc83b666682b86e63dc8
z4bb44f60176998e3374c2a7e1d7f6a0ee7adf6ba81f374ca24f99840d5aa6e2fee30b37d1d4f5f
ze00efb24251a6709168fe520d0093f748a500928a42a4d1f4854f789d14a2e8ffb5d541afa307d
z6d5b764d87d49a07ad9af0ce5d576acd84d408acf0b623ddbdf97513c40d7404b8b0b4de9e74ca
z9a0a03637536abb254fa6dd2bcc2638ce27af3456c88e33e267d3ee0cf61b9d371971a0d5ff1fb
z7506cb7d57514684bcee67e34cd56f521b8d146a2deb70fdafbcd8ef0f423513d513ce66e661fd
z5e7a0754ff626c0563236a9e912cd04ffaeb0fd4fc61d8e50407ec59e363125f26cbdfb6f56e0f
z2d49668815fadef097057b87748a9896f84279df914c0a1a1228173654259a58a02e2005c94d61
zd80796f08d38c77d1c469ad44c8574f4060d49470859240559f6a274e6ac5fbbc85f1b2f5d88ea
z5bc2aa0d3aa483ac8e8ca2ebbf80d6a63ccde16ec16386ab4a34b044f6b025e58a418e3cf27075
zf032d9139b4ec772dd592f0b4bffe509644c63aaf0615f316ce5571e4c972cdd9099bbaa4c4fe2
z96540c5312a5201d0819b5cf0e7f85dfa626dee28666e1834407764cac5c887f993181b6a138a3
zd42c33c41996e9a3b0792b00655ea9d3a7e2ea070ca8a9910acc3f9c2b5f3c6a127568e1fe6496
za2c664dbe569d17bd974131d7fee037f0f608f6af6aafd8c56cf9c1b9191082b8f7535cb583451
zf3161faa6c86d3fb33b71b823c7c33b3ca0b26163964d489dadafc3c59542a2fccc8d389e1d871
z690d3d2d8af3ebb1162a8025094e30ff0bc54f9ebbf9f365bb8124107a4c09509264cb2a524d16
zd1d256d6c84afe3501968532f665f614710867dc7a3352b8133726b8b62e587bba6771997afdb8
z591a85d5331b56d234e995c373bc644f6333c3715e262342be4020fd72539afaf40acbf94174d9
zc9e90654c1608f4af33cbb45028812d64f4b57d812343f08dd46f926baaadc62f43a5825757ccd
z08743f0bbe227d5b0ae0cefcfd010b7ee6cfce2f7b28f58b2363978046c6be44d005be9c0b204c
z7c80e0a7c95094ef1ce3027139e4b1379c29be8d675b17b78ad34b0fc0c90eaf73ddccd0a292ff
z1f4344a2b7807e85a4554669a397b710a8f0223365023cb0bed70be54608fb99a4f99e015d102e
z8691d7ff0edc9bdccaabe88a9fe04cd471a4d786e8c448107beee08eba5a7ceb7f1f0b02742d72
z4396a9bf5ce3208937b6d8f59c06c483e3950416072579335daecda76bb386c0d8183a8ed17e3e
z088f6feaf2bf24502339d1d7a5eabe66c127d8090b02fa987eb95868a26ee93041a8a5535741d0
zd38837acad77a43d6307957a37853898ffcd0d748af0ca2e9ecf6d7a02a30c73838e37748ebc10
zd048c229746a8373de806377f381849f3c7a63b704086dc951514acd848315fb7e64821e231f7d
zeba95022673c28c875088f8c5cf4a7bafac67470660e0633057c0e625a48ab515e0d072ee84e85
zd7eab9a81ed7ae88057c7d25bc414ae522ec44941b1e62a42426ed7500b622c3c181ff3c70844f
z048bcb20fc52abfb9843bb1de1c5a99eabaec13e031f3b04224d8a9f5fa9d53a300aee42d5f8b4
z0c3bda879ee2b3c77c4d613cdbaaa294b035608defba164116e06bb7cde18c1446c56a2959252d
z43f15b5ec68ec0cafaddf59bf772536d76224a7e3c8d03a0a66e889d2fc0593d6cecc4051102f5
z153c12b335ffecdf82c32ec5fe43b652ec6e1ca2f3414611db4de26e6e92e3676e8eda89c53c6b
z0da0dec0971f52d6a5d6c4c8f44705b3500de1b320ffe8015c7aac1c7f60d241e09221ef22aa2f
z6a4b45082b2b85121ae3a511ac27317410a3d3c4bda709639b7802a034b6853580a05e4b8f9b0b
z5b508d15684dbf055c2166b2da999844d2b1526f40e4f871bb601bf35a23939c76bafdcc453098
z2949bb78f8f89fd72c500c77b3a7f079bbf171f4775c5efcdf4e85747bdd0d7a8636f22d73b88a
z77b567bbaec91882cc22a9f737f6b875d67b2b01cecd79ce658e5de8f2b5bce9efb4ff96305a4c
z315a7eddd64604352b67d753e863e7f580f1579e04a22fb46b45aa5090df8619b159774dbddf33
ze11d277117c4f1b2030a4a647666ca5e16d6bc51f77b05b95882e44476174f112c58afe0c1b908
z94fa37d440af5ebdde3859524ded96e168d2cd58ed506315929ec840a0bda2b0d1f0008a65fd2b
zaedecb3e44b148c1a546311a7f068799bb229b3f7c5eccfe40156fa5c0d9c48c6ff297638eb4cd
zd7ef6b6962404399036392cf43c4fd419c532243fc68e8cc5a0db459eb5415a4153e583b500f47
z4f53ec2dce7a632f1c5e6e0aac22d2e95f337ba1eb33af107ef6904ed96838ef67a0c43be85493
z6805020765816770a0fe41a387bd60e09f5209baafad59d3a12ebb73277a4541e274e0c80db04e
z1eac6cea28628e3ad2664fa6fa83a2840c8f339bf71222819635fc78e59218a4548a26486ebfd2
z92e35be1285b4e33558c76a781dda4c2f3346988a7122ef2597b414e86e9f95a864aee3db3b588
zb4c050c961b6e210c1d1e7d5d77989fa969d0af730b02d94f54b80c388899fff31493f6850df92
zdd42ec70f09cce956dcfc7d137f862ea87b020f8600012541b3e1c6e551972aa18d4322a668484
zdafdc54da1618025bac84927f57d401e0e9d3f35d5ccc1058d806d7d5a5d365993823f6ce77199
z0027d92a0cd6becdc1a60e637846fd986b9119a28617105de36aae557b8323c204a5a6f017e9a3
z7b1a7c4dc9d4b320461967bcd02c81aa46ece9bdb0478d2234589ee535f4d7ca34683047681f26
zd62c710e0b390596d368fc2d51b6cd0a8b2e56509e0189409038f12edba1ebcf193de6b1dac944
z6bdc8922e9b7447c7d828b3492c314c4f6191db06cb10058f4ed91aeb13503472ec277f8dd0460
z889ebc77ca27cc6f762da05a05a0772cec4733e25c964e83fd40455c401e7e2a0ea79f72b7e0c9
zd9680af65c1bfa71cf72f2039a2198d12f5ab6763e2f52694b1d1cfd3e2439eaa01e30b5a1a78a
zea048858d39fa7a900442ea482ccbfe4124292b6e6a44d8194a337cd55d2c9c949e22c995b308d
z77f66de547bb72ae56a013d9f373e3ff5ab9473d78fd0645bd8c6ae1e417f11dcf686c45562844
z79dd6947ccbc569cb506acc5147e3a3acb7a4b9decd50746f8562885c6fdf84894b47e272c9274
zb3df3bb0a91d03f5dd1c15d17a5162d2e42b16a9b8dfdb8f449e36fc954dab12272b0c22dd982b
z3a3b846361263809ef88c1f4d63c2ed54b24f61d9133e65e4ad851bc6ccbbef9604b2502d71f09
z52dcfb7987aca488c01832d401e52e42f7e483796788fa3abd06611a002e8fef6f668b88d23d2e
z784cf5db0a557357f301bae178c191a17a7d6d1a0cb147cf7349ffaf527c9c1dfaf812380a5eae
zf1c5975a70f70594e9746c22276fe96118a483f3bd4dc2081fbade6f5e01b7d4da7ecb4fe87206
z20cb50f1e26afb52edd7cc706b2c61692c044f1f2cb9d79f580f7a5e219c611a4674c675554476
z9fb146297a7621759d09cfe19546c874eed6c9245a845f80ae2eff3627efe7da6589ae59697067
zd697f2854797ea98a59d63a0f42ae3d85cdccbdd25d040fc57e620c64ac226de47caae547b8c28
z1f592a8a3576ec818e61c730efd4eafc39e0754cf6a10db775a0952d2bb915ee2a9300c8a887d6
z90944faae2cc2608b19c820624336e7f97598e9a10e8d3e7b439607966db954f128a56662f51db
z7d29b203017858bc70d2a5c88c8616317b7c1a48adff2cb9de63afe30491f18fbd04b8cc6bfe20
zac1ae8a6eae11ec3cfa5534e459f450a74986212b2f02549bf4c451b9004892e72aeccb262040f
z1b4559173aa7af2b904e9ea5ef02793f9d6d12838cbcd3cc3145514b0c837db657ccd7e62530fc
zec3e65ab3947ac7a1ef3ad081a50d0e4c6f8cbafaf396c63b7030bab32e50348084bf4c605c214
zd7d49b97ac76895710d4c94f885a89d440679a09ee862242858c32b9044be67b88cd57f71f375c
z3af4d2cc3c003858e843b92bda313e6e0d31e482c10deb6b16f1a02207a9b26493f90c6327d984
ze16b4d5fd4b852ca7d9ac91ff19fde4c508e44fb48a322c05b93059814c0c42f942d65aab6d293
z7e57c34b65439744f05cb2abd07aeec4e6b7fef529c4032d560cb92b2beb20e452772e3feee327
zd7fdb228aef085f97649060fce479b5e16c04ecde9f29fdfb4634cab426193f9d22177f06bfd8d
zc9fbb0e2d10268c04b9e5292a18abdea76948606dee918df2e94995f86a34a85a4172eff9b9834
z2623d6680049859807e7880e6da8f5514a2dcf264085d7029f0a2340eb0ab5bfa254102a5b286b
ze60e2d9f0f052e98ee88c9df98e1ceb02d3e9a38284c35810a1bd06ae958c9de4e5237407d97ad
z0d362278c52a2b5f1594fbd543d0b5a796311e425d00e530e106599a0493e67a50c9fb6ca7d6aa
zb5de2e3fd4d6877739eae7675fe5f8c2497ea1ebf83621b06ac7a0f2244b188b97f3830c6da15d
zfe36ba5526295bfbc5e7553bc4efa6fb701f5de0cf5f9a06d920685f073841a191f65bea0ba674
z63de22aa8694c5692c5c7d0afb50a6833b5bc98952db069f963d19c4a064d8680e77b464d03cd8
zb36df4cda771a17a9b2dac03fb062981c135bc5dedaa0ff3533efb7a997cd14de4e06fd0b920ba
zbf5a6e0f8f25715e01576929d86ce1e395acda4c275b47fd8537a48bddc32dbd6dbb451697dec9
zdc3964409176dddeb6f59dffb67d155b1ae5423d8945bfc655087357b6b1b791a169307b151762
z65ac36911a5c5d5edd280cb5867b02cd2a439dd8df62543b5f6556f8f66b0e41d37c31528fb9ba
z9143f8cf6ac211b2c52bae485b07d81a530934b891375a0640e3aebaecd69db199b11ccbeeb8b7
z1170a179729831db2e6999697010f9441add974bcc7298d21cf38a19325c544947739063a4319a
z12ab55f58f8686182dc1049571fdd7c8552a4ca73758d878d0c6c183fd052cc822a495940c0d78
z8a791cfdf5f3ed2a415f0690611b7339d9cf6e641d0261c5bf563faff1b38cae9f1d43789edb18
z1dea11c5d1f4205703fab4b31fb4c001fefa8af59bb2de538ead86343361689d4c06404c5a6c80
z094abbd2a8e76108e199c7b7aa07e668d60413ef76d658016b2618a1855a92cf34da0fbfbd2730
z056eec448650198111c2c189000ee899d124680f8906dd55ab9dc2b0658208f9f3a084e0355cdb
z068c0727593a1c7a2b247266f11d7244b0b04509894db4a8970562ad6cb40675c2881534c3f906
z020d246f8d996c38368a9f92763b464f20861165453000f2a37bf374852a4e219650127926a3aa
zf7b4d4acce1756b79226546e8537fc9cb26f7f04edb6079a1679ffd2f3f1dd160c6bf5c3676d50
z8efff4bc46944955e14adab0480f6245ea1f89c8c6b6841839b59e8bfa812ab3bd88d7824d7113
zc05897f16977f438d347f521fa32dcfbf9ab206013e51d6f9753f713e73a03a385a027629dd428
ze6dff691346b40e5098a7314d2e24ae701070ef6ff7c8ef37bdb5595a3132b5c12bed3841a05a3
z16b4f456ec52c2bc63a4569965b289a797078084a6147ba4c7198ac526938208696eeeb78c86cd
z7a42d9a2a0f589e4b09a6db5a2d44642e26e9a28313608a156347fe0c4145b90a563447fedff4e
zcdb95b6fbf5f18a6ecb0450a00abb6360233d087903f6f91de121cfa2508ffdcd5b2cc5763a1d6
zf952e9ff42b139e3c78bb37c67be92517317c0ad8daf9d5bb2e7e948107796b33cc29e2897fefa
ze9bf4b201a5f67dfc94675489897f86496721940879b24be1b8e10185c47535b4b928c41c9c41d
z88e59c6e60ca7339d796a3bc0d92e008093a26936306cade8c6c1e3d6f043b1765da65feb040eb
zf16a6769118c6d2d396fb5516989d1428c9d5badf5c71f25452ec0ac59614ed2b2f8a9cb97a005
ze019b1caaffa40df4ba8f03e64019ba08a7c3b15c1a9d0bfecc660189a20b7a2e658d655834243
zdf398b901a1ed3f35b5fe308a0e90e4c95095b1ed30ff5e986480e3dc18b2554284b31150ac647
zbae1a501ded5a83804bdcecd307427f3831ee6640bbcb18b81031a12015a345d89324c9503c154
z9d2e0e7ef253181f59442a582b9aeeb5ebe68a4b9e130e100d15ea105b197f3ecd2c225a82ec61
z34b3bad6795a96dcce823f2c01b84102ea1b7dba2a302adeaa8821bde207425b5219f7c6005e1f
z88420c0838459a3894a3217d6c96bece52917c7566f961a61cf5ef15b4d8a2600d60fbd4d010dd
ze50fb0670bf1bccec50233e005f1a66f92e82315f2d76be45161771a46f65ad1c3e7a1f230c96a
z6056e45dfb8dd05b70e9d0d760e8b9f8d73221f3d46540a372a4aa2db6c418504eb39e1b02da7d
z271760f0eb6cfe89ac9aebd209202bf9882f74bd04b1f3baf6ea820086f49b86d5e18328922b5f
z1537f9b76a0a05e542d98ff957bb4449882efd69e79eb465e182aad782baa08bcd1e07fd0e6807
za5c0753fbd4e614d0bd27d118fe27cf0ea40148d5ca9da31ef2ed4658d0de724c8e4675a084f59
z30a087ae4ec28c7db34f57137db7364dcd703493e9139b645369f07e810bc684c11ca872fc4d7f
z3a00e111ca5b78e1bdd0f4f924ab8747342befc6eddccfd40f83aa596a726b1a2bbd0b7b1bc84f
z15c93fd18a651c8ee31b3f0a568d706cd6cc66bb466cf0b42cba6afcd37cac620f1a338014ecf5
z953a6c329869ada21bd651973b5e1096fae184d8d6c36a78b1e08a24b3ea915c88d30e34ac735d
zd168a19eefe788deb1a247fe121aad873fb9b50aba7753c4301bbb491f2062bfa7ec8a1eea86dd
z7bdf029ffd42a5704c2b51afc4c66c3e04ca3d9b9878083dd815633e49ca1bfad7598b621728fe
zd32a6e8d2f05012f2e1571f5a9664315ef4a68676c4b706cb3b361da62f566e2fc66f2cde1b42c
z56d01f59498588fad6fba2192c3c1808002d6858f344f5e61bf07c144419bac94ac48fe729936a
z53661859be7fa8eb3f6c529c0c8be0c060f257b4c8aa0345ffd430e54ea20841fb85d59f7f90e3
z224ddaed979c87bc0b6bd7e4f8108ca4f2386152a4cb12535980f8e446dc496472d721d46e1153
z43d66b1f3fd3ee443821bd850a0970e5fcee2e61c9c93e9e15fd89e625981d78dfb0b6869a63c0
z1db9a9ed5498d7a09971753457c3fcaa2cbca6d235cdb5d6ee6486dc1714a047794361b7875ccb
zb27a95a1e6c43cfbac06d27a612c283e4bcbd0375506124dbb0b01a8c0ede450f8c529471ed8fb
zcf7ee50772effae9d6b0748fab8d813ef4aa4560c81f15884a70da13daa1f3d06f30dce1385102
z011f4a32cd2856c683b21c0993f4eb4aaea0c0266634e5154c65a20ed76b0c82a7fb882edecdb3
z514dfdda8a3a0bc100b890f0dc9aa488e47573f766d37324a213a4838e8b21fa396f180318fbdb
z9b438ef957756c25b457b490519977c8cee198f8822a63b3abe2c1e51470f3dd45f7827052e68a
z22a2ad4253b7e67d45ea40a436060ed5e89714df37feee66946854ba6764f1e965ce42804c9ffa
z5d7f70115df458cfc159494d55238c3096c3bb11a50934948e0582843a6a6736ea677d79ebe588
zd89e79b39ff9b9a3e368a97e48840dbe9ff244e2959b53af5dfa92d8aa572ee7f0d2a45821a066
zc8ded614a62c797e0854304954e97fa11396b31df2948dd357df8cab76de027f1c9e4c989d6476
z64423b32e3d16eaba2b9e341c62d3be07f6e38dc9b0b76255da7698165e165bd8ae0037aa5f9fd
z6d1019847469c8c4a7bb3a3794dab6ddb6ce33d8c932a61c77fa28a864f626a954423fdebd14df
zc403105c8f8957439e496c5e0b793cc4c5efefb99e391222bfef9e95a5bea377f7fb9b1302f57e
zef08a2c13783fa95b3c5034d0adc028739bb058c1720c9020b73c05431bd490e584213650c448c
z55241b4f694d8163433704e8889f44cd8eb315b407f5e9ac1773374b874bf78ab14a05b0ce1da9
z51ad508ad6998d631fb39062522523057917d17f7718659f8774351845f881d5139d9566329e4a
z7a7418f1f0ed17a36edf9553bed254f9d5128c8c69f86b1a885630267930d1046ea313aee28602
z9e9bf264d0a8ccae1b4275b31adcaf73512dfc909ad51206b8ab04e032b266357c1b433d1c91a7
z55ecde7c4cadcdcefdc80fddc53f07172d22287fd800c33a49c417f003f2ea6d1af06a717a6b37
zedeed3452e4d401861804a8321eb928ea25005537a5aae2e755fbd7b804a7192fa31e2d7e0c8c9
z2e24b1ec65438854e50d1d56c6514c1f957e97487b5240a17a4f1c39ea82d25dd0bca164169045
z1a470ad0c65ccb026b37b2850e5a494fa3398aa276d898ee89db3f88a32e283fd907019ec556de
z928959a3442560ab7f9217ca7b84f0795cd03b7c11cabafe31c3874002bc2a5c0113eb50c27610
zb0c4a715d089de0f62a4c8cefc36a8460d3b3371067c358e66917ac72270202e54304ac840084e
z166f3676c05785a69b1e0a6bfb58a40640fc340ac513e1ab9c24acfc6282f51ad1963da2dcc612
z50e5b9f1b91669918b5f705b0371da9d05a94b9042cc324df6fa85674d8256d067af01783467a6
z8a103b8782940f5ac6dbc9fce5a46573d1aee350f5531e98695686c355bf73c547c3ccb64d1b05
zb85dcf92ec82f3fd31270a7585ec4b22cf825582dcdbc9e159a0e1e56dc86e194433755b11997c
zaa4027af4ec03fe3d1ecd201785fca3a8dedaf01794b2d7f3b026cdd10afaa2e0c769e3208eaeb
zb292470b645aa9ebbaccf50e94a3edf64066f8d3300efb2fe98e97ef7350d8b7015a012a41c29a
z98d3166352de8c3155885a5be87c3263493a361a5826fe2de6dabc8eb91c4447cfaaea4abfe928
za7a1b90e6f2f553130d55d888f48b06c22a911d3c08b74d6d765a5a11b362d2fcca41ccd06b143
zce7e03f3cda38a8cba965d426494933707805130b828fc9022907801581e3432a903dccb92e4ea
z19a06a1cfe42d21ee7e6bfbac0ca153f2b146173c1e22ca04a5e235e5bda736e52db6df14cd369
zcc6ff1ebd22e8d06acfcd78a48428b16f3a7cc314953b3c83497ca7289f416406bed1d4a6ec8a5
z1e5635b276c2840d572a5a33a7aecaae847baa765d796c006ae533dec0731358187d2293dd00c5
z385df7decf9f6b32f36d29b2910a44723d3dcc4622e5f78a83569ec88819f190dd84869bc2d7d9
z00d9a2ae968ca4401bcadb142d349904337029eaef69f59ad6fd77f95878ad791abd05890f6063
zc72f314e6d0abef0c0db432ad85a47d1c6f680a48b7d1b5dcc2253f36ee10bb07327622211daf7
z8ec680b11020a797c9f3ba8cf5e79ab4712dafbeb37018939c2e535056a8344021df6fd5077780
z31c9e5b5be12cbc5ed4b303f6a14198d9746473b7f4b8f34947546b368e134506c51f91b4d99b8
zd495ebdd046469be2f4d856ecff45462d43bffdf17e84c73cfcb39ec61716e10e21876244b5dbf
zb0053f51c015935700ab3eff1962d8bccf0d744318db1f96858b539ec682988bc6aa0c45669a45
z1e6a2fdf432a97656ee0b086058781e8afc3261e30d563e23949f9bd29163113428daa5b28ee40
z5047a30aa3695d8462c3270f00e9f45b383f1458e78133f142ca5359f8c75e25fe909ea2961380
ze4f22a04ce4a8fbbc97087cdbf42a90d8addff1b736049eb41acd04f29ddb85d2ed12151acf5ce
z942fde7cbf5b3f838d7fa46a7ea7e456c690ffaf6e702f1bbdb54d53791cff3f023a1958e2d8f6
zf57e536b015467c990d4c2ec5d030af70c9f8b99549efa3d4ede5b73038c6baa1c7e6e58dd1c3c
z2eee10cb3b451e397a3dfaebc5ecbbacf15a0b6b4c418e79ef07214e3a20c5dd65fb61099137a6
zc66d0515f3017964861769cd9a991c550c80ce2ae5d73476cea2ab410d12f8fe000d52bbba86b3
zd282b0d52784455f8860659e481740831417b43380d7659c5b975953fbe39b49962a379a4b6b12
zfe24d925596861b2ed2838ee971366cada5a6857e8379ec0d833775feb456427f62f06732a09fa
zfcae1ae3b2bea8245f6ee82503759df7fbe4bf8c574d36e4e73bcff96b3571d856aca0771ac677
zd2d5143b43bb93fed80520eeb0decc370c01cecc8fb0d78d8079d324e088370e482d7f54e84f16
za8626ad75193cfd410ba90a33b16c5e7ffa909d1e211cd9473653ad2fde8ae0ab47968f89c67df
z9efa08632ef99b5848e08218a2f353dad2e8f6f9a5009d484082707d189e95ba3db06e1bfab13a
z7c2a74b24ab6a72fe3e11cf1d19cc5952141e38a0f8fc884ccaea55321c9b7cbd4965decb89457
z7df4c3532b9c6486af1ba4793de7b9b791bafcf712240b98b5d46ea452f6d1f07e7463e8147bf0
zcd425b7f64c2ef8a3012fd4777623e5e3bcec7cb010614b76353729a4f063df7e2fb55ca8f8879
z59a71d2f83082afe4e6716452f5d2bdd218b739ecaa94d09c542738591a7dfb5c3a73165c5b4a1
za09904d92162b0841a655a25d45c214ecc1e11273eb926b2dc9bc1c0b7d77a86eb8560a708da5c
z0d0a1d23a731bf4c33ed071983cb4f9cbb8af7ee5a26ce9e1e431c43c4974b3f757a22bb43cddb
z710ed215a520fff05a14ba05229a5459acf6925ebbb8d67d2cb3b533123f1cc0784a1795c77b36
z5cf18254450514d2067eb2cf926326e0d26c828f4654cac3216bfb2fbb706557e5f07c41a61d34
z7c8b8f3415152153cc60fc42ba4c9eb53b684dfe6e9234a3b421180522e02ce1ad2104a5a8c95e
zad598c1a93ef73a407c0e9632dac25b07a0e5a02fc3b836f9ac723bd510d7a01351ef6a3a259aa
z3b7dd2384e0ca4f889cd20813c3fd2a1b954c18ba88c9fd459fb691c129f66bf86632a322fa552
zcdd847ead686c8e7f71ae67aa9c429ddd0cbaaddd31b700cee01f6cf0f872dc761ba51a389c0ca
ze09e6f236364fe82cd4b610337cec442014fea8c13e7e48b40442ee97b1465e5fb6fe36adf6e8e
z608c5784a52f9302deee485a3b7df4651c16b358da006469f5cd1a3d289f73b1b7e6ad0ee04b20
za76a360c757b32842f0cfcada0605161fae1fa33fe62b290da18b8911e113452f9a378a0e01055
zafb6559c896b23f032d81b10d76fbcd2216dbd9fa64200e87019c01616fdb6c116d2126a148af3
zc229736c6912783f4faaf4c27ad51626cd03e9c6ead8dd0210f5c80c3c0ea3dee6a42486d8d34a
z7410124414a2beb5c507d020c5106a5f01f397474a9229b7a82401aa7db2f2ef1fea7b5c583c0f
za2a4c03723bf836f88bd0efdc4d03b003bd3ee13a5b3c478559cedd36a7ac96d024fa64c30869c
zf2eed04dee15d3563245c61294c3de1405fce1bf746cc90fa2e45700982853e5dedb2689668364
z22e1c160751065d646cebff1a84591fbb61550056a900ee02d337d327ed092b672372408b31191
ze7e2efa285c26b160b24e8a5ae89d9cb2cec19e1cc96ef5ac2bb6dc6d65975fc53ae5684567a73
z06ca19c76c43debb915348b087c75ec3ab8adb023cbdd4b735f4a0b6efc2978c788acc3ffc4f3c
z1cbb04cd31484c1136fed3c497d7f180e71be6c8ce71fba97696fdd3c82ce0798ba36758012d5d
z5b611df7753c7a4f3807c33b1be7c33ee6e1df679b6cd9af3644f082fb02f3545cb53f3934650e
z8d1b5002bfce726bdac8720b19e4e7a1b0e3415ed87f5b3666b373ec98ce55657ab6d3641a07f1
z1b3aa1852b409047500b7f0f7faa43a512ea836f3e693355685f05240670e09073d0d5a0cc9176
zcc4811c1e0611ef897d44d0da8a321f84af4a0bf0dbb46450f7f3b0b0da8d70fd4d58a7593661e
zeda56a357c2e08ec85df1c96d9f17970a7fd4c8ce1f98cc6177decbbc9bb4eefccacb0044dde2d
z8d0d5008e1fcc247f2db79320632547c2912353d0f5ef0df28097ffbcbcb4981abae0703ce6629
z2b516de1b1e9f51c90e5767717f455f06cac90d796baa7352674820ae75e795ba557eba1dc9b52
z86461d45ff496ca7e06eabd8f4f16fee49e26a2f7fdae650a3cc23150bbb67d1e4c9eedfadef8f
z016c175c3005b6b3551b08fd350d35729d9396405658ae9b215933c82834f76012157e4e45c2f8
z2b4eed61e9cc5d7d55a1179a38fa7dda9103c635dc6d4753a655eced9a67d2e4b7e55133c3eaf0
z4dc42a5603a660b5f169c7323fed9ed1fdd6aca76ca56f1d6abcd27f3655fd7c8122e5d5a6e88b
zcc00dbc36a97c68f2baa2b967be8f7adfa1578520f73f8066bb77508c6eeb5774fc812b632035c
z78a68ce1639cee26d28e4bd2e22f09ca29aa362d87be5182778f36ed092bac09da588c2e0ca320
zca49b0269a84cb209fcb13229d5d4bb5caba661b186428e9d202337917a4aa422c4f52c688f4d6
zbb69801f49fb912e4a1d79638a273b41534e4abda1e9fc69c933f28379f68128fab9fc6c41b78d
ze0f0e96b3883db6fd004fb243c729829b9eaa2c6b6cfc8dda1f4edf29ac5d1bb4b3b1d9a1ad146
zddec6798ecc5e6230f3ecbe5a02efbccc40d16655bea8957218aea6cf0639a1491b43e77d22e95
zed4f94d55fd58ae87dd4afb9ddcdece4015dcf88055c07d99e40df85d8267250ad35ef7ce6c4bb
za9e3a3247e50bbed2b9b83041cbcb1c3652ff01fb64d966808745fe2e26427763c621ad660b56a
z49466cfb2349138273322a95b4640db0beb7a1fd9ec0940ff0853ec32f3f190eedf793a2d05899
z0ed15f93694fbc1b0721ff529f51b63c59ef74ac36aead35d5711fdc9482833845a3ca702007c5
z0c079cfce4c20faad28419282a6c077e9dc9ad3b26f2533659fa48e8fc01552e67e38783a40e9c
zb367ee2a54df7222aec136f1f2f07e529e8f58ddebc5ad47df7b0647e07c97d4fbfdbcb70fb8b0
z8081265f8c1762dcc5a2e89a5902ec76a3e3c9514f0cafed74988b92ff25e17f01c7c6d3b1113a
zdfb837be48f5439f8c1f3453f3353b0a1e68b27d2a62557c59b5f10e3562cefd882a3c817c2a95
z12898b905ce86f7e8ee2e1b448037c0752b5a4b1d5e759a383551e2307af960caec593ed76c603
z86312db96ba3da9f44e1724b182585ce6ee3792e5dd0e0d43a091d10f2edfeafe88539f1d08d3b
z8a370de401b4f9b26b89bf213143d23d6d1615af3d725a0a720cc8d537a126e03b6e7bc15c9582
zbba34069c9f1b922db07a31354746d8fc0fb19738b2267fa6d0f7a0d51f02f96e9d6879e64599c
z35d2e7b93c67a95f22f480f40c4cb76046c1193e79339027366943a4286228caa6c3dbaea4bd22
z367086a66f99cdf6b3f2e9c78eb1af7d40e1ddb1c69a7f40ce871df1a070aef78f9d8b035757af
zb692aa114d48230ccc3e0f7d4bc463c72e270f92631a8f2eeed1d41334e590e6ed1a35d2bcdeb9
ze05e13c94ef81139c1d83417724379f64b4a5576a05e19aebbd5704cabde8677e2f2ff280d959c
z471eed2b524b68c9c23434c835ac97da02606f3d2390e054b5b191c83691ac881dbc1a0b12bf52
z2d24a777ee9cf2dfbb13027cebe96120fc3e061a7c35b1221b4069c8c67c5ef6900d68b59de74a
z99115b71ddc59c926fe121602f2bdf556134550df8703e4e6590d75832b3196774636b698cfc9d
zd07a445ba1835dd992811a7dfb6e6b2a646cd2e9775ba429d42091f45aa82606e7eba8121bb712
z1fd708eb26e6b572321d1c5b0e2923822e899cfcb05fe39b6f431178e7f4a796283e2e709800ab
z26ea636b38e6d984cb886300c9c10534c15a052bda10605543b206fed9034de5b1ec3c081d15f5
zeeae8736d07c3e74cf512b0173d45dcde933824ecc7c044c383441271e0d99b974ffd93d581550
zd3b724cda0487ed7f1df9ab47692426bf6bf7a7f2cd31f44c2cc131a4068b48620b6af7d7ab1c0
z34a37408b8ab9be5ab68647b198599472e73da90558b25545148c37c447cb9d46818ceb3ad370f
z8207a0869529eee05c8d9795c544dc74217bef3f0df6417517ffd3c297977d3c5bad43972493cd
z062b033690f962c769e289470c23e14ace757e1064476ccef4969dcfb30becc76c91c4f7f18a86
za3c46b1afea161441364786949f299431b5195edbfb847fda5987fb00314718e5718377ec3484d
z44a1ef77568b9384559e038921ea4a0196581ed6345469d9ffffecb713f631c8057e8f933c8e2e
z81a3ada3f129bc9a58c0b1c639aae1ded4268327bb9b13af7d048ed99a8d8b96c6c9932e8f977f
zb0208267980a25ed456ef4cceb1cb6955952c84ada3006eee74f249d8c56b57cf4f61b6f7208cb
z560452521d2113a76a8a847245c5d9d56dce1546cb0d1572e9a678cea4d485f48a9a141ca1d81d
z922c041770754e7a01ff55c842aacf3aa979b3eb1e9a189e9530c66257e46eb153f93813e52e03
z87019816c0860423bb38d5f7c78599d99b0de69e173c12569ec9cf0069d2526e18662a5445751e
z980b2084164bada0aa1f3d9514ba699391f592a0d43c8654c70e95209b1dfcfd5e1efa694dec47
z9036c23c1f5f2d95139bae3ec952e57e96ecf3b68e14baa9272bdd50ac7a4d21fd486c835ce137
z44aff9e13a676c7676e81bc8ecd02fecc99c8c7c5a7ba1219fcaac5b9bc77b91e30eaafede20b3
z6b1799d437135cd003960904ad8d5b4e1cd7e9f63fa5973d8ca16e8f764bb8559d9fca2d43a799
z53ae40954e0fea5c89ef60d1c1eda15c1d9cdddb32fe3920a0d89e041049fd5f7cf2cd21c50073
z58319726246530878752cf3de67585fc49ad3c94a350997c4658a2ff718a949bda380dc0610c1a
z771d3e4b9e7b2724aac494649401dad0176a07253130a2fde4b0e6c82f00bb9c65e58982095399
za9ab59ac8413747ca4b672c7cca0bb73e2bf0499b77b96ce552c607ab243d97fba10436e564306
z377a5be5c41df9beb1f27a52ede1d6c5558fdd118cbbfd249e705805f02e01e40b7863e0482f00
ze3fa4a2c9d58edd424960110e9a802f24210c186bc045591669332f7420e5a1fca2230f92cb3c0
zd4175cc727bdf7a1effc8d24098fac3e225705618e5fe73c651438d6306da35d2ac46b118654e9
ze2d771218c16fefa4268998a96b4e04c21e45e9087f3f79adb2e6bcdd266fd91b1ac16646bccf8
z65f4c1f8dee013ed69fc9e98d4abfc0bcc98a2bf2211da0e7cdc0e4241f1a102ba2e8116dc2f90
ze3cefc696a38f01d55e6674832771d7c21a76374345948be958fba6a5c92df21087e1347c3f0d9
z9e90a904c6204fc784012e782d4a5e7b9b5bf8d3591456b303f0049ce013da4b136a59fd0eed3d
zada499fe9e6d12d1a60c8c1805b18a55f79975856bd6415ee1ca0e1557ad2ca5879216af637575
zda71622d341ad355415dbb3c7fe7f4bee71a4e7bd679e66eddbcfeaef3b10cdb51087bed5548e2
z3a8c0c06213be751da0d33c43b03e28cee50758a109d72d70804cc1a475277a7db87a2b21965f6
z0bb84cb178dd5490f558702c4124b982ba455d7a052415a718a3ab8c710c4ecc403b64d505c672
zbcc70058ac671e75e2cb982473a498034f2fb775bc4b3ef087961a3ac707d41c8eb03da08eb1fa
z64f976246aecd8942ff1da164f7c2e78eb5d7d2d7a51624dccf29acc77356fcc31b63222982fe1
z81ea41c9ab0ad340745ee38a13f7ef22fa5c5805d7e158e11a612fa37b98ad4c29fe8b9d4fe057
z8c141da62d826314781792389f99ec0fc3dc634bd4c2a436974b9bf25961365f9122b2d29b7c56
z77b952003b7c5644e09911c85f092828906bd9152cfb092f0b08f498458e4b96bbf1cdf0193f25
z7edf3c3869c29c4c90471838508181bcf7954fedff6b47e6ae4a4ebca7cc91b4402aae90da75d6
zf8800496cd4653a820f1031d0d350e9be6cbe692211646e8c0720cda753f68069908bbd90dac84
z57628030a037539f43926dbe94f692f170f24a6652a665979a6a0fb23765464ea7d5fc8455d6e5
zc3b78293764511045e92a5b5172e507c146bedfc52830299f4ee7d882a661b69381f8db7f8b5cf
z12ff303e4028959e99a9dbae57ab8ff6989055c85bb1c505aefdd1f8f9018b5e1bf193dd2ccd26
zc93c0813ff7ab678b401db37acc4d1621dee97cd7ca3007d0a752767964e7d500c5978e6c520d1
z2c6db1ff01b606aa81acba639364ce35250a6cfc4a55f67f2d0d66ec1676d6d9bad19e182fad2f
zd11cca57d894442895dc292d1fce9248f9eae136ab9a7dc27bad1fb5fc9b8b1f9e57aae0e3f1f6
za413b962cb15597577ffa141a183f3e4f5ba580c918751f0db96f4c7fb745a4b58b0240d062d40
z6bee318fe946edc4d47ccfe58c1ab62b009aa52e49a6bca1380f8516bb217a5a8470cde2201a81
zbf5d05fa2f817bf86ab5ffb76cd427250a16d0e7a074ca751669f11debb00469a6eaa8b5ee9143
z879e0a0a26ecf0b6647274d4c4fd9e663a06867460287ebac55b21a3debb13e8397cd9bba1a8af
za260d4465dd3ad100a3f8d965c345636bab64e06fc808ed54fe8f63a9423c31aba139be8b7bcf1
za52f062f2a754e40a72141ff4658b831dc57f34961359d80577c66235e80e95961fe27dab42b47
z9025121089ae4743a7b5bfdc6c86d587dee34813d7c3597566be925045ef61f7123432914ff24b
za5f747aca5923d054d03e0e0e1283d21a526caf8293dfc0871dca63cb8367fd4bfb60e3053a0a0
z9c51c6e139f17259eaf321bd38af17097deed6e475de42cd169ff9238684ceab142d4c7cfc6da5
z31979e28dd7e8145e4d6f8f3ea87f802bab0c3a6e5080780a319dead22ebb89b4765e1fbce11a0
ze07dad77d2cc4301fcbac2ce688eca6993eb79266526fa807ea8a1644054d16736264910a46efb
z0f563a52bf65dabf432970daff0633761eca84b1e9e682a9327050055ae47a867dfcb2f60750e5
zf7eaf730e4dd61091bb642ac03e3cd1a8a315fd22d15c3e2f9622a782d2272d1644b6d481f7cf0
z5f6a2fe3d778d5eda32b5b94f71da471574f0f9bcb95109551243e33f290d67c630f45bc7be9d2
z3ddbf3af909990a0fa81260c042a3449c9563c41c1fc4db2dc703ae09db20bc38eaa69cd0ca1b2
z11b214add7e1e7c575147b0c9fe25419f946e65ea9dff60675e80ee277dadbab6ab8431f56812c
z8dba3cfc43148627032216f77afa31c887571f8bec2832902800a54f5fe2b88036c353d2971f9c
zb1425b411fa3417def37578e6d126759653dbb7be0576d2b0bafd63f3805a0b7158fc4ff22f24b
z0732938926c9859c592622cfec02314c26dd9f32386fe25ecf96a959d37be6c7d4fba87af2e316
ze2d0e8b398a5843d6bb1b00dfe90ece744b9f4770c863f81d280755cac595a53a1e3c299af84c4
z69d57c17a8438b76664089219bd3e62c27ed214dfd47dfad0c017b4eb38130fbc72cc51776ef32
zfb0033ef063acc967c190191cfb2f01e44e487e8a251e906b02e091cac9456a92e9f08b63d89a2
zc8b5ff0ee178f58a3aa5921b5b93b040722c78e1411ce896cccd5141ecb4ba775815981f91a40a
zb60f75a5c72e284e79798651106ecda4ad11145a88a2f2942413558dd14dcfef619b137703383f
zaa6ed0962154cd849033ea381e39b1dbcfa22d600588fe6d1d4af431d70e9eb736bf04f668436a
z20cc7e111ca96626bdc117e10b9ec1260231a1e9c8058fb892a97bcf147afc36b2038c8c7714b2
zd5f210d28c2ef3e4c2b4dfb731a1e1a32a2c8ed6ea2c6c73ef39d12a8c08d292bfb00b117ad5a3
zb683791284d5eaa106fc2087dc4d347c49b0847504ec807b9f96aeccc9cf66fa85e48a805e15e1
z7398c4886442ca544bc3afe326709aa214a64555650a9fbd562a544a00f5c51bb04188bab7c2c5
z78d23703bd91fa95ed8380b29548697e8ee346ef7c397913940d51505040202af883d5c450df88
z61d162f024ff6e9d02a25388c330b37aff08a79d859fec965dedc49818636b0bc2386ecaaf616e
z558a68f9897d4d70e0145c242ad97f73bada0c3ef47ccb5583c093e1e5921fd4ea97682d537092
z97e5f3d07dd6c00ab18f88493706de3544395874c2d8b67d3753c3e11e439ffe92a3666ff84f8e
zbac9a934ba15e92da711be9494b2733283133cb63bdd2425748a3560687f9dfffffdfd1ae27c5b
z3a78d4b7b1e1c74f88daf8ad8af69259182d8a50c90e51fca2cb4ed1865cfcb4fb446c61fbc343
z9e8c8b825cdcc96c375cdd9f99e23c4410dd433f02773cc9e09eb37062668d911bed5dda422224
zf1d2000ff8492f9f1a4f79faf693b576977cbe91eb161a1b8f3bd05b668bf0c59482e33412c954
z7ffc2bc1947bf76528d8b75595120f0650b689faea337d7ef92c3d8594bb646866bb97e3d23fba
zabe5865313d26a0a7c872f0a077382722ba4d40a6c1072d4819e3b63f726766f3ef9db16d9f3a4
z1cb159611e6fd953bd2e7d5eabf5b9c0daaa941156581cd5973829a505ae9c77c0b5124928654c
zda4a4505f7059e64d26bc700f8cff56db045d411f394f9ca98d5741bc4b5522c11c4d461fa42ba
z7bf9d0a1c8c7b07a0485f90bd05c010255992bb9e15e092edab82049b4c809a7893d980ee3de66
z7daaf2e92c9d6dd46dd04660d11b00e3d14bb39d5a3798b40648adcdbd2539934ee2989aa73b41
ze935702c7a0602325e355fc116d6a60b34d969f6b12ca63e5d8939d70c204cebf499a0b3e7c9e7
z16cf77d9dc12770aa8331bea22115a64469bbf63d01a3fd4b79e0183db31d25963e5ea888640cc
zc946233684ba96d8162d6f65bdd945f56b7e1181d7c4fee1c58f08cc5047915e6d6f25ec0677ae
z7db851a3b4def62ed8dee1c97bb947e81fef6786967619a8fa943942761c898de584847f373175
z1ef7590b9fdb3da87921a6a759482eca157276f4beec71480d915ffcb577476dcce8ac53369177
zeab8908cb0c827d4bf89482a17756d9658d374d1a63816bc5c2d959a8607a1c84b06dd0ba6475a
zd75f576da9d1a806e9700fea7bd92725176ff155d6a178644c01e518748a4628a6df4dbf580883
z7d8fd3e1c472debf919dd119cc9f8171ea0456da0620bfc74afb6c628f5b6addb9a0aa6fc9b8a9
zb96517af396322feb32d3413e49afaab50b9d1d5664f72dc9bb890ccf90567a7741eb20b5940af
z771264f07912cb6cb0fa328d34709272a54ec84f0b1365b739954ef672d3f14d6bccd984f98be4
z3df581be600cbd4d78cd783c2f23d8ef740dd53d836833714a1a23238aa5ac45b78fbe44b4072e
z1b68918180d8640c2c5d26af293a0538309a28643424b8e9e344fd526af54d6f8a85730a0c8aa0
z5fe4e4a1a92890f157fb10d6484de7ce5cf46342247bc0ff36d908c29aec64e7520f9fa8621659
z2d710f214418173fd6e1f1eabd6ee9db6359ce724e1ee2476e7fe622748d925044c088d28aa68f
z7595301859ab20ae5fa4cdb6ced04791262caea1feeb74b9e871a525affa3afaa04d6498b31292
z2b2d5533cdd7c2bbe827dc073a6281109ccfdd2274f07251f18255aeda045f7a82c31cb485d70c
z654daa1642ede3c0dde1f1265cc051708c66c6238ca79d7c1320400085cc0ca0e723d501deddbf
z32c08857f315f28012ade5e860a5eeccdbfba98fcc9e974418b645d412a6954c6693d793912fa6
z591a6bc173b486d5323f4daadd34a5f0f2f306c700ac7017d20275c1e516df4148cbaf711db491
z3e2213955ed8a4c600514ba5d5cfe35a48e43a19c910e267b7a5d264d0ea5d4c37efa90674c755
za74b15acc164e462e60c5087a722609b4eaac972f53bfe2d5271d899baece0473c824e04e9d142
zbae523aade339df4b235f688b1c3adac0dfe0be80695e8e17fe70b1725390615baf54ab8b3aa05
zab2011794a02916bfce4593da1af7c647d017aa78f1af9c75d215091490a5bf63db2d4676513d6
ze8b5f578dd184f40b4db269b3839bb4a5b5b947b24fb79e22af006c70d4a84eb5b9373c60fa9bc
z1312d2f658cb30e71c1fe67c821e15986f7f6c5c8bd3796895ffc331b94c8d3be5a704e63f32ba
z8cf1c59feb34f212ca0a25dfa6a2ca0cc6edc4134faee0702377b5e8f5709795ace45fec812d4e
z07e493277367a02c88ca32331661d4b43519b6edf252d5a1be43f35bc8e959cef38e9ba10fea4b
z8478016c2deb3b69e58a5a84a4a1d318486f78019a594487188bb8efa036e23c92643879c6c5a0
zd84ef83624b8dda9183093fd2db2f86616e3f83c0efe4de5d407e3262f6f57ca2e47958b4fabe8
zdd6e791fbbef5cb09960746ded295f1e0f688b4981ed8a6263c5ae054051bdf50ce53f0178d432
z8243b9b8c03ba7630862c46ec9260076d3374e210a1a6d6d387409210d91449498a1d0ae4ef861
z0a3df5368b5e5ca3ec9273120e687aaa2977b67fe6ebe293529449534338367ef43450ba4c9952
ze17937b4e1a9627f68acf93d92b3a0d04c63d1897f1881c32898f162a04d365efbe7685551c335
z4086a7c5fb248247becafb6c32afb4d161be92693fa049dca982e0991aa43fc73a82ece03a59ee
zfc0134e9809ca5b0537bcc0ca48134889d1fd17c245749ed020fde6df6c5d1809d0d8185b7c68e
zd99c0f49fec7432f3476d28d82fe42d1301842713265b7568528524205b07de135dd2dfc7765c9
z104d019bd58131a0da65c70abc05c6f15f7ed54a84d30e10891a5239e6ecd2c8676f59cf3e7425
ze3344b4419d18e72fe4548ba0a091ec5b8098372346d58956f5730a65de0c1d5ebec580ec1deec
zf7a106ce4a8de6126900f83ada244e673c116084371ffd03d7e19b55acd5ee71f1e38fe7749c2b
zb9d2d07ebec7a6ae25985bf624e97d3b952146838f3cb70218d66fdbbc74242d97610c951b5c5e
z6171c4140b66b7844f52a5dbb4b985f0de9e459c3db1d14c6e98a46fd2cc0fa33d68c3b35de1a2
zb7d433017ca6d854f4aae1706074329ae2ad287e03448fa190de6be89140e95c653ec4756835db
z0bebfa1d24a785e5ae2537c1a7c044ddd5740136d801002329d1a727fdc8221d6ee5b44f431bd7
ze8f5cf93a12f7525613647f3fe4e480a134f564f28e5b486bf6c13297e5ce567c5d40d709081d6
z0c94d8bb8c8fbe58512a27bc5d67bca0ee860e5973ca2b2f5614aec50d6127c6c30dc3545accbe
z44a064421955e7fe7ba3d6cd926d8b19d0e8def310dbca76a32fd9f8d21a9299059335fe16e858
z8a329aceb053594a3bd7cebd1a787d856ff10fc53de3cb0b93d7fe58992864e22c9dc936a60717
z339bec5482f1175a140ee6b3e1853e3beb6b02030d13fccff85e2e5c21b63d1c8ced413b0fdd21
z7438d93931d359f698685c822670b426bf3f9d462bd537668c3bf838088581b1a3a824c83f993f
z5adf2f42570b645924506cf1e9c9cc2f2c78618b9bca7efa146ab5dc8be2624ce63b4973393ade
z9b12aebd1dba252d6eda7a205c7d5546ff34ceff083213a4041026b97858c1031c11164533438b
za4e4614ea3b85bbf964265588b62170fd140aa4b5f154b3dcca4728bb06002d87949486f7e8287
zc20a7dc149064c1d2dee82c67e1fc8b0d8c63eb69759e99bd3d50aa2f5ddf5988433ef7dc1f0f1
za34e725c106f416c2033499e11ace7c363e0b1a9acf4614b59b62472f07978ea56a49cf3a6e668
z70d8ec3591c96a3ed39a168c7de0a3926cf0fc4c56adcd1980c1b8486bfbbbe0a2e2eff6f7c981
z599841ab5819d861068a229584074f330f0414968cb949a42e6fc0fc7bdaaa9386b3b062cb3166
zc75693f40cbdd017583a658f71594a5a5de251391963ed281be723050210f7697d11f58a67e222
zcfddd52cbdeaae227df69dff66b992fdec48a3c9445129189120b4d65f48d56695c9e0171e13ea
z9a9a829bdbf0db9601b4c91c0b14fb4ee2514f50637bdecbde1977d6978c03aea0e37a2344fc4f
zd0af6d7f1c8d8673ed9a979959e300caad9beafee45c2ffd25d6c863f54dcb6b1807d0440c4258
zeb0f00148b6697e43107427b47d6ef05004fde1e83ab84e7ab07f4db34878d6077bae434bea08c
zf532d4cb0a8306698b93ff7f5849907469f38f09b4b1b1eb104dd179bb582e73c83aa4d7951ec5
z4274b98441ea581e93f9976ade65532713ebf10d432989da0967672252801471a00f14429dbe7e
zce906fefd830b1e0883b3415adc6a04e4d8fff305014bda4d5910c48ab74c19306880d98557a55
z2b48aab8466645c485805c05748ee7e3f05065d0bd7fa2447b59d23cf5ef488cfd8690275d074c
z7f166441277d0d3c0e4def42f12383080f107b2cc6598e8119ebde16728202a656151b58c1df7a
zf2249c154d7026292e8840456a8af99441a72e3d736260c652ccbb4df37ac0f1ea55bb55698655
z14c1d8f1163117f79c72ccecc0f4631bbfb89bd32162d6352cb68a0949c6ed1940742e7d38f497
z9b5dd370c65f35c88f09176f7b5f451c9d3a3de350ab23b42f22568ca08f5b76aee138165b4eb1
zaff7da3b6576172f9fe026fa33418c2242f7613987592999eedba140f8fb5340a4d746ef75f0ad
zb6ab219dfbf701f58b03fed303b418b078e711bdc7c8364678c6a910224b4df597275b35095495
z14ef06bbda164e4ae02ed11156276ebef97a7cc3867576fc35b9f59d181a81427c1c20dfb0520b
z1794156cd37a896e5d44462515e9e1105b14590d5443ebe7868ee038156484dc41adabc48e8414
z129cae313d4dbc33c43278d0fff57c8f526194ea00dc9656b5275564c8e165a7f06c0fd92975c1
z819ca6bc65771d40eba407159c0346875100df4ce5fc1af4439d990b0a15e0cd9a270cf674c354
za67ed457f54c17525d9184ddfafbe7b698d552464d34334aca881bf216c2b9d75184e222c3967f
z137e1af8933d07deb494f1ab9418a4b2ee3df3de2e2675cdbed230db70bd1ef326c0d746f53cd5
z8d2ebb5b836857bd8fdb84665269b9687304cb8d2fa851ca7249946e09d43570c689b72803abe7
z1e59c1523479b7c62d693a68248476dc5015afcb1d637788d28fd1b7b2991d7c447f292f8d60fe
zb6f381f802b7bec260d4ca473bce3d1612a0c271a895c991d3b7b4bcf45779215c4fdd2e5b50b7
z78792a261efa0b090d97c3eddcd37f7db3a4e364c270e39559d9a24673febf7e027b747abefd5c
z86f158fb03028ac36d9084bc36b6fb58a231dd090689c82a429077c1a6a52a1442b9ab84ab5ce2
z3f280aca1cf6268185810d413403f208bc20440f27a7a4990469e66eb78f6db57830ba3525d8a1
za3ea95e36bfc30f35ac6282ff122b86a304971ea4eea8ead416f883edfb89b67c6975a5b58cc6f
za5486fecd4fa701b4701f8c8d04846469d80048c480977bb1c2fc709d786e6cd1120d018fd2982
zd42ede12be09684eda07bc398ce136e96241fcc20d4a974ea154d21f1ac7505c5711c38b7d6458
zcb8cff00bb8ebb146c2157fa3624e8f0e2c29e0bc9ffbc25d71c8cfdf35de687b0e28e19b78cfc
zf7d0ed2241e247e7d3601c666e0e7181cacf5b4548fb7daed8f032329cf31bd70e5c038ee62c3d
z3ef91d3e355a5c1f3fa5be44740eb98845c4163033e95e924061f118ae7fca53ef87af167df55c
z6f941daf5bf414770ed37f13378ecdd3b9c458c24aac5a4f888e11b927aadd97d6f2fb37d29495
z7ea963d11df035a64413cdc582273e3a007b878466110cd07a1126e23c39d2755004babbe89c18
z5f05c05c307260014587f7639a85852fe524c283f5c88055d82c4961bb341b4f25991e3ce152fa
zff379aa203ebe5444eda2098c1a201e5670294442a01a4f0394d8d7a34dc3701e30fd12ef26b46
z5b5e2ba007322b4333f76846b57aba9b5072ab332e3d4947e9c2da7c007077d8aee3086972a144
z2e6f63e4dd2c4f66953720aee439b77530581191835cbe376c5ff168f8b6c799d52a8d532ceff4
z175641e22c94d0bdb9cc2fb84239f5ba9fc9e5927414c2128e845fd163a6609a92257596bd2e58
z8c4f20d617850f99f73a0c200d110919f98d5bd9e19d728450c6b49fee6b7d0d9326e516f03ca0
z63f2eaeb8ffaad97c2954cb1bc9da5381e7da0e5e208a00981c40a5f1d2d39575e8ec28048719d
z27d23a7b4916c1e890f032cdaaaf0b31aa12cb9cc91c13992f5b61a71084fad2d8f63f1590fbaa
z5ac3b63410e56fdb07c404f9b64e6bb1d6e11c00d1d49f0ec61b7a146a7dcbc03c47775dee23fd
zf91485f80e8b5c1b62695ca82fc8ba117c65d421929608dd400338d7d2a440f994f9f038d22599
zbb96b2fe70c323b8c2803395ee634938aad849edfa5785edf58798ac63e777098d2ef0c76ebb91
z960549fb313cde773aec6139f4f33eb57528bc27bdc34396939e4ca74998c8eb1a3d7d35dd7444
z70cd23b895d62e4b0566c41c5e39bdc5e1eaca3b2579b812011be7d138248ee6a573b0c63c4d7e
ze623a5c751ae8aef6f6a6292356d516ffba17858dcf1b113e5f475574107c193b23d97243be8e0
z89cfbb496f777a9791be4f3e94ee1c9688be73c0d6b5df6d5f0aa8a5e1ebaa46690686e6449427
z4edfe8a08d850b04116731d8713544b047248645b84c263e26b24b6ba59dee20d3e611c01b7d87
zc5d23a3207e76b18bf93eaaf28d205a3e168d4df890b693fc6b1a7bbbd71a016c8e8e498c7a23f
zd216194cac0d82264073f0340d09955137d202083f1f59357f7cebf0a9afc4863b83910ea37bdd
z17820ab3b29f13ebb187bbe5e13cd1a0fbe10a7d34f56d0150beb634336ae3b99987fcf9a63729
z803135867f977429c30bae656538d8534a929cba0a1155d55a29ba59e4decf9ab2995933a74734
z4202dbdfba32248a7d5fdcf08df17c7b23ce1a38d36b44c79260482b4a5481bf304d1a0dfd9c43
z3cbb97c554e87fe27547cb1c91682942417a3d263840dc1b690ec766d2df6b3ae0cdd18d5c3554
z581adeec9a4ca439fc69a3cba3300b1bb8ae648ff9cfa24f9403a004302cf1e3d1c2ce33dfbc45
z54f4a8bf910c1a5a7825e152f33c7826637a81ee33d90dcfe0757b09b29658e6c4c107a2cff157
z7c5f80a0b9708a295506b91d360b994ed21136bee0ac38f0ae4fbc2af2d5963532ece286023319
ze93d7e12ec92b93ac9f4bd0b3f698c47b08e2004abe6d84c30015a20bcd6b90b5ffcea1e446744
zbddd604bd6464b8cd1e1607f2439d8f79c9e45a7bef79a6b4b5cc3df39caacede92e05765d7806
z1d63455273ecfdd804731845b864b7c6f5d268c7c076e042f87e4f9a243d5545b5ebd201f8f025
z919ae38a656dbe8ee422c1ee2076a2f8817e2acdeb37e442ed2bfeae06097a59317e5bff816cc7
z7a3812b8f3bf62c3feb52225960282d908d6a9d9958094e8bdb52e6895022dcea146fd7e13583f
z82498d2764e806e9bf451d9d2a86c7f0dcbe5036e93a515c19e4f5f20391fb944865b799d79e5e
zf0b21a6a4a9cb6409b9cca2bab432dc30583cbf5bd268a8ea94c3b52d134155221752e55300269
zbab6778c1f0a47e2cb656b9e5dfc6c78b3730767f1ccbea3f858c22f457587ba5f34e3940f4cdd
z9acc845a58e956c769cd3795f3ce26cc7e187e1b01f097bc12bfd5e5f379b78b0c8ccb9d108ada
zb8ccc8914822921ca60f9b340dcaabbcca152139fccd97a8e8068e67844ca9000162862a0545d8
zcab63bdf0075bdad12c3c3ba310065fd5686ac929bbdff22992c09332ad88089cd59a329ae4e83
zce87192c27c14fcbd99cb6f57f0697bb74974f7911ccc2570bb7f79f92ad6885b2b6876c589947
z14bf3112eb7a2b0493d10fde77a7268d82a0ba56507f5711f5746a2637b443002c125417d28691
z6796ff0ba835079de8f985b4ea0d90b24b54f4f249693c8a8f46eec599492ee75381d2cbd8e45b
zc593bf4a945f75bc409f18ca2a9838465f58aff5e85d41c6a5a14909a0b4f041922fd602268b2c
z937f9990f06e023dfdc4baf62e5342c38a724a2dbaed78a7a9cfe3260d217b8c5c43581fc03df8
ze1602a761b3c01ce52d226fa0e6818a56c9cd4ceaa1eb16be27dc747d063fa1f1f7384e5d412c1
z1509857100777ff398c31e59c1d01a1024b878cb8b3ae4197f98b95ad1d002bc743a9c79cf1acd
za53290c125dbced880c0cdbc30654a00b3295e261022a9b3410932af8eba5bd25a939ce2a60582
z40002eb1deda2ef48a53b12a8243ff14718792bd9bc7297f2cf317d88a9f3c1ba053aadf1c6e4a
z7594bfd7fe7eccdff569c63ed5b9f30eebdc52b162a29b34d92a5b6849c2a093c6350a6c396bf7
z91831292fb1202092c45af686c3d54b692144286835cfc33660bf6d9ff1f1830695789ad2d5f1d
ze5f10adc40c733e86f6c0efdbc5432a1024b2f4db89194ef52ccdbe691f467cb436d56518347f1
za00fc92df2aed2b025e3d35ddbf87a0a01f38813176c9da1588224e6e5ef2342b9a52259e133ad
z95c0bd1391c67cee753a239e8cf1467117f46a5dcebcd35f556784ebbfc0dae8e21fbf475f55cd
z08986f3ab6793e709c79a0109c47706552db1e41089d83df4795409e920d3bbd478e36593957c6
zb42ac72ae05ce3f4b522c93274e9ebf1233c35946348fe47e639a43ba3780900828f159964d547
zda2174ddfea4f733160d9223090fafbad6e0368500979d1c1b12dba108d4454ea919181e5b1f7d
z530cbaefd9561a0f814cea6b9e2b394202459774b4c35f24cfab37ab3143d767822ee803f2db0e
zeff83f482acb041c90e9a0a71b1558d50d3d6906a8d83a72efb7522e4a491fc6a7e8838e2a35c0
z07460b9004bf00c3a578292aa1fcc7b987be1769de6a51fb37b45e56f767e56fcd8819cd9d3af5
z44a1e26bab2073d4ab8be27ec3c74bc4f6b61660dd084e23330397e38141739e0ea331bd243f01
z8e4a971c664bc23d3d5d107be6906e4a6884056275e556cacda0d4ab18a3455cdc91f81d8307d2
zf11a845c6e09eab9e9a0789716640de39521efbf0aa990aa82dc3c2fdfb913640dfd4f94fe09e7
z4bfdd3929eb93b09f084ef4b5a2556334896335eefd1f1efb2a36c7201fc74103ad5521a95f5b3
z144140be75432eafa3e5d24b8f56ef42c6de48e6a18c40796bbae0ef0b07c8075cf730487b0040
z7d285582d35dc02d28a8cadeee8c750a9dfafbf62218dcc549fe8ead05d173e9e95edae17c6eb1
z10a284003bf52e9c757d9bf87d68a49087ac6a888a9d3dae0e76ad5b04dba11d2204b878e96a8f
ze5a074b6941f7452e153d48db09bb4719858214ff9e2e616b99b6d67950bd4c41297c0959e8e66
za1f05c54d990db26fe2287f247d5986554e08400c70161ae68ba4631903bf13e0154fb4f0435cd
zaa714caad6997445af0ed364180b59433faa8178da3f10115e2d894da190ee0cac0021638eb08a
z426a8490044b10c6d425a868d3f64445a8a38c33207ace1552d38a7cf22b33e046c7818e5b7d77
zd06d1edb21c8a99b1a043638d2601318115e91b6974de7a7df631c0bca2c970c6dba0697f81729
z02247ae880104556837d3a775700090257effd5c45921af539fda6d2758bc4c9a41bd0c7f57f85
ze8f7b38f8c1a6521bb12366b316139d6a0b1c3243b3503579585117a12dbc3f02bdc8e3cc04628
zfe83e8778421980db106ed33f8700ae1d56ca033103e696d5cda396ee9e562c49c540588744d0c
z3e683075d704cb4c0ed0f3b079aea5491dbd83859b7edcafda122ac506e50fb92091a8b148d95a
z94c53ab3c0039c174ed1c7bc121495716da2906acca93bf8be3467c633d61611caa21086ab74d2
z43a75f04a02b1e7b9dd824698172869cec83f95d2bf67c6212d7bdda2ba2d1ecaeed8297826edf
z6aa3c54d4d5b7eda32bce7ae330611fcfd328e852f9715520c31c10fdfae3a6a61d0ab1c5a7b07
z2b4fb19046d35fb4ea152faad1513f5c177377ad4ff82194dcda6785890e8495c721d74d39ea7f
z718e910d8e04c4a64f4002dfc732ca77b3e30d1c9e89e9b8e78931dc5b72a14684cec48b6033c9
z0f9ee945832c12a209f345e7f18ed2e6d397c761f4f51e57d17b44ba366c50e5b38c84440200f2
z6e792e78b76f26bf0059255b82ae481e414ccd1698b92c186bbc2150a67adf2ceadb7e249f02f8
zdc99a8847b735e4caf22180d165a6fa5396edeb9bff9631a982c6a5ba1c99d15e983d7a3ce1cbc
z0f320435b37322474ea1ef28f23be8ddd15fc75c693b33812561d5671175c8e0c9399290d38a76
zc6a8e94b6fd4ba56323442b8e112d9e03e28537f049a042ca2e29d8ce5a5b469ca8d6c5a9c2a0c
z7f33aebb522f8315822d1125c1ede6b2ec6e87e31561e8b893ec2d988feb05fa1f9823b523b1de
zc4ff797cd069be3da49c84dbb0f91bee9834c941f9962ba7a6291a57e119ca1200aff6717050ab
zdfc3a58f819d32d538f6a4ca23b15cbd9e0b383fb02a9276b935fadbd12a839a0dd17c9f2896e5
zc98f9296bb1689768205f71e409914805fdbbc2cfcfcf7455471e113e1b62607ffe34cf88727fb
zd0037d1306964d46ef257e2a5b4f6ad563da5ed6b314b4dce8afdb16f9804d37f38c63d075b735
z1d964a95335f484bf61a6f7c51dbfd62079e58d23ec27f423e3f38cfe8cea72c9bebaaf47e1be8
z579a000b87c8e2568a06254646929f8917c04f6c236c35f03aa6706e0e19884a560d3dcae39b0c
z4044468d7f97249aad9bf97a52e11c6ea48aaeee009d2bfb507b6d61342941dd829fc6b6e94894
z839cc8d9ecfa1c791bc2b7a2bad1e05df7844963830bb9328f401fd94226dde499338ea4475451
z989493f926dc9572a82482d713caa2e05f974b2c299b78c7440a5c3e71c516abab8ee63d9c6bff
z8fd9ad0a855c3ccbf4f1cc6f5cc8080d0df0886f08697e1d4b01c8e532a9f29a7febf79f9c95a5
zbb8c04c14400900db16e066bc4352e2ea9e59ed274ec8ceee0e0a5e119441d5e43e53d872f5f32
z9b7911a1ee71dee9380728c20c72c452febb676621d9a8df83aeb0be0151345f37475b188acc49
zcbe3160a3a7f63c64daea7a1e46fc5432e9c29ef03b85720e6406eba8416e60a1f2a9821ada516
zd910f6d40a1b7a34d3220462e9b52e9927d97b6c9430435c7114f79025f921bb4332b447b56a51
zaeb83f4a9b388e24c9eb72d86d4e437a3a19587141f0e040db8208d616665f8e645934d4ed552d
z5694ee097883e7f269e595486bc3b883ead68c3183727b2c7ebbfdc19598b73b4a65da5a7e9bc1
zf6966a53de5b5ebc9acaed8310ee7f7649e31d706bdba44dae0e93890379404b3e136a08c2b3b2
z9d1420ac7e2fff72c5c0924d7985fb6ec85fdea143c91ed4b0c07160f5e2dd63ea4503bc57cfe3
z3e19c7da58fa98102eb293342ffc8bd3b674a3c37117e4e1efcd7d689a37b6fb7aeb876ac1db2b
zb7cbaa9d4885204307c01dc1e54e19b07cd9a7a5748867574ad8fc2021bb3e0575ca7676449bc6
z5d0c712eab7d106ce55784f14b7e1a28360bac0deb591df9539e1844692e15da239e00417d428a
zd5bde0ac15d2cad9aae6aa0e0c61189b979cb9b195fa22b390c5ae15b583d067966f9b77fb2cfb
z75dcfc5ca64e599f55b3143e73efc996c821c61b963c72898ff111b79848109fb08c58ecb5fe27
zf1c4ea0f00dcd23bffde8ccb6db976d08edacb63729575ac3ed64b3a5be514d69b4a0a12cfa16f
z7d65d4260bc02753091d0a31021d07d1c7c0bafe7ceba3c0dfee85cbbf957adf04ad24cf61717f
z7cea26ecb4a2943a71d6e03f70e205a24ea870640388efe00d8469ebfaeea7c7cef3392801cee3
z8d4074604de046b082f30873ce17bfe0f0163f6a65f70f14ef4a1f78feefd2ce2215b030536cec
z9d414efb0bfeb232626930b0bc199b5aacb8915a4468835990d045e1b4934658c24e55853ee1d7
zb118c24120db2a731c6cfedb5752617471f7a4936a82ae31e0325158c9ddb55164de7e1e42c5f2
ze2e6f9df70aa048196198981f8fe26d92bb6a6242d93eef03598e7c2c90bfdf0e025ee0fd82476
za411010b9fa51af3cbb83fd916fe15e491fe163181440465ea2d71b8772b22c732649e48a1cdf5
z99d20771f227541c23cbd73d66622a79b5654289d0e380aa9a97c5166c01c6f32ec567c7e3aecd
zce2eb5d6a4be92b7b95ecee88c8371ebe2f50ddfd8b735ca1eaa43f3ad7bc04fe8aaaf854e0343
z75b788a46f20e1d47df3856526963aec8ef26318a416e27cc727d31ab14c250c9dfdbfb078dbbb
za9559bc217f71531ec134e44a0044daae701cf133bed493953b0be155e0f013607151a090d0044
zfc7a16347ff53eddb3e5e85224473403d31882f0320c73f53aa4e2cde3af77564304aeeb588c30
zaaa54b81b4d784c3e7d19d174da595a184055f1a02983116f611d36f698cad8261a71a42042e56
z31d9a945c4a1e73b52770d393d93796dc2ed3a84fddf8ac82223dadfcf45a12277095af50727f7
zed73eaad78e71233c6080b60414847509070dfc1eab6e9883007b5de0b379377ce617180a50234
z71c3572f4d784aafcd984d3e16f5aad0d5677d64348156bf0c273977bcaa8ad7b6b7134e5945e7
zd4834942861c91aca538701293715276356bc3db6de556d942d4d117652915d336cfefadd0fd72
zbc5cd2904030c99d3291e812566bb02a36818f436882803281522fe6bdf3214b20a49cec1af7d1
z4436761f8180e1e9cfd89161115ba1bd0b601ba56996b5af492637dc71979ed97e6b57f101be99
za56a35fb20d17aedcd2fb29d80b512e3ea572aa1aa2fd011076fafcd407f77e798fdaf826d391c
zfa3d5791afd2a5f40c2c1bdf079e77169c06e7db744db4799376ebe796a80a27853e568b2a8aff
zc709460e7781681fe0023ce402f900a6055988e0d2d9851d45f5f747ef364798a9262155698c74
z1c2222929deb77065f448fc45bdb739d4c56475752461011cc764a49c346022908d9d5d9a302a4
z8cface5dde3cc8e3fafdc581e9b248bcd5b8a8f380a232dec0e725c31fac9be62d5550366f7cf2
zaa67502e9c88c3f4bb8f1a319b3fee62742fba36fe3172f26c5b32b728406a89e4dca8a9e8876a
zabc74a6947884df865dee6230940ce2767d94a86097cf1901e2bc33af244bf45dc0793989ebcf6
z8c4ce3eb2eeb7a88f0cf1934305622da27517daeafdc6e8a1ae8ec2bf77533f059cb130401036f
zd4adfc25468ea586d6f3232e8542c4c869f3097ce80f94ca5bea1a44556758ac0acb312c6f2b3f
zfc1db5b8d66f0f6d06f05113f98a1bd2762b72c399e360511bb937e5327105a86dfc361f682e97
za1bb96ba7934e3834a2e0ddfbf526b13bff22fe89b2d730b491035d6fab1653a559588c9a4a49b
z23aeca3471ecb58291abe3e4d4d8597536a65efd10481d8092a5179a94a49dfcc7c35e78846d6c
z9b5c80649a198081c1e5e0490c0aa724bd76baeae41ff75092df107b7ca000fc6f2d5cef126889
ze2e805671a5dab5403712d99b40cf0e7ec5a434c3e9f822e91bd2ca7ab827e042bba60acf7a36e
z8da58115a2e823025a50628bc8f8af41dd43d31980c3051cbf6c54b2d418870fb21740184d6584
zd974f247d83f4c73573752fb558d3b79716018f25ac8557fe3e3eb9a1803df975499315bb58a34
zbc705bad586988803fcf116df0d329ca436f24461c6d66e4ad023f6932a667e4366a86ba322ee6
z789c24813a3e4ed16469c035c13bb193e86b8c5073cce6214f22102ee09cbce77d4f61ed83cf7b
z8b9be84418ac664fd70d62f79e32d27fae4a0485dd46f081312128f50e06c41efe58f2a9284dff
z6f7e993283598b9ddefc3a6559b98360995f334bd4fceb936cc9950b0e957d6fa40d3734d938e5
zd6e4d0861fe2fe6506163647eb594889ea7c138936f443cef06b6edcee26598ba201f27341cd5b
ze1ed59716805ce19dd5ea4b101b0d496369e25440a7ec9924841d04701d521020ab07df4f7726a
zcde33178aac0775007011d1bc87a528cecb0f0b4e363241dcfd1fa615fc0b7b519a9e537a67edd
z2af03a8ba6a6a4142e1fce53cec63f97641d079486431c509ccaaa5f15a0423f811c6342e6756e
z0afd344f1991b8fc351c3ef6942a1aae6e80431b9f1265e56e2ac5a8f4dae84b4f69e938b60cd2
z5c152f10ffceb55a640f7b5ee9766eae97be929b514d7cc3873c00332bc5ef7c45e4a47d001347
z8a09504f1530f05e9e4349200fd964840b9249f5651de2d415360c3437eeaf5127cc7129070f75
zc4bea6b0d807a61cc7ac8a2c8e623b7f2222bbdc99c34b05d86be0881acae33cab41001ecb213f
z87fb8c0cf677fd69c383b8adde3bc3d35e2fdd374ffaf865ca76fa36cfab2d6dbf5b09d30a57bb
zbdb54c398183345e3457cb688781f70bb64c56753bf07faaa024263ada94476832f80e1fcf7313
z54c6c6767540bf44abc4d11dfa2163417fdb311cec4b53f7d9ca28764a3cc4b7526d49bd22aaef
zd7d245d414ddd84b2886244513cdd969c5ce246b48fa0273850ef9407b6a5f825daa2809d691b9
z77ddf78cf0a0e69c52039ea896c25c5a4abe7efda1fd0f9a9699fb21bb6cfcb88e0c43da7860c5
z4f058328c3a4ce5cb3b80d67f26bd81c00d1c039a6203614a0062ea81fdd84f06adf90820536b9
z1cbac9b8addc21f52a6e8f59e4bdeddd204caa06da65d9b1fe47558d0365b9dcd9cd67072c8c5e
z059442105e1c7d12cd74e9388d77cecc70a69980c6d72e93311ace2da6e8453f4962fee39bbb66
z88f5fe6fd3676adc4a178b622fac6ac1b0c50c665a4b6d5f62a181df30bfa5306c051e865a0fc7
z49a98b719088c5852e07843b7a0fa7599735a595ec75a3bc88ab76a210301328b116bb1742a62b
zb3d6311519f737f6a004b26f12eb83adb95c2322767e56aedc467b8a9159f7cf20d514abaae5ba
zbf8ac2820e4d8c17678eb32b7cbd44b2b037adcbfc22fe0232d0d6d34dcd7b4494c4c1bf5bcaec
ze8c944986dbcf2c3fd256c3f47487ae3ad02ad232af222c728f0da53109bb65ba0c8d5356ef59b
z420a4ba16a8773bafd9ebde1bbf801f953da81bc9295818b15d9ae6474255753fbeee1b4e22fae
z69c018c1c5d731c4fbc0e1d612cab24d538a27a692c20da25da01f2e12824a4872a8d7d081db31
z1a119037b31473d6de7cce9b09ec0cae213c0bfee5a75bcbdf174c7cdd6803bc05c0cf49c2672f
z08e5e99593ea0b16efb89fc27f5c43b003d30f4dd6aeb9070f1f195d0452d865bc0a3b3db61056
ze7706a14de895e103ec850810e458aa243c2330e6f93cc512669e253f29000c6eb7271a2380d37
z4d3e9eb54cce482829d90450a94fd6f12361b9e0c62c30ae461f290a85202c466cc95211370ecf
zb8f19851ca7376f24c0b9c8a74cafac1e9c63ab606f866fe119338cb9ff07589cf39e5c1a65e44
z2934895cd81821209406af16b0e0da9e9f2eac00187a50f4b066365d744b09d98e8b439b9625ef
za009a87e1434c817e93b41b5defabebdb7b170b477dac4e9854595599b36c9863216be19e40495
zd786a1caa77e581b7df5f404408c8e4be87cbe874b0f7124a3c2e3c15d7747bdd4d3071b45b7a8
z727d19323fe0394fc484c1e5f41b8838b2e4604609f2164a1cdd1599e560f81e5214165c836b4b
z43ab32f3ac0140b09740395996b4a0cce43a60449ee42e168086f1ab9cd88a920b759853ed172b
zf2a3d17f1f674ae56059f063c1b70f9da9908d6dd34bc7e4d89b06443b5109b6d5f0cc74ca7170
z6f8c26bebb30a3fa0da8bd5e087094b69538c82fefc696821f57cd45ef8bb4e83a64ed45a529b7
ze9676948cfdb7681a637695d279d3f087f0372fd1911da83a04674f8344835d3a313808e05bbac
zc3c6816f08bc98a18037cebb9f39a6a4714db4af91c284c3cabf064977dc6ebd722cd7a72029af
z2f3dd92a59794c11f8a37352eb96adcd3091a81d55d8d2f32a7ae436c7e4e96f9861524a62284a
z8e446e2a661ea2cc8e34575e03e376b09ca83cd6cf452fa289291a28bb97ffc77698b1d5faaacb
z2ca46bd83c5d7cbc221c87654d04ef45a07644d141017e8db53dd77b66f4d7f393d7ab7f448081
z2f63408886b8dbc4eb07ac4f1173b4be6eb57af85b85aa9c09e46d0575bba9cbf4facc93466390
zde7b8984c6cb213bdc5b14cee65ba6d03cfd8053c0af12a47f2f33a3c45cc08eb3767288290c0c
z4480023935f6d7afc338a8e40ffcced1b67f4cf699e6359c1128c52fb16806909ec1d4f7690779
z0f364109a65f6747fbbe774d07e32537c86c8642be3233af90331266232da3b28970695a10b591
zc239c3dbc96a3828ed46e487e4a3d7fb898c9e53ad604814a524b0eb0becac2a5a2370ddbc048f
z5a325a74ecea99cf0064fadd3ff337d90497e438fd030c0f3d18deddbb68df38e18fef4b5c7e48
zf70c32389f4c07e15f123f0c462e048aae12038fda2c3c4e6879082994e03a98eb7e233e1358d7
z28cbedc49f737a313ad95be69d775394c323298f1266f1dd581713bfc7bf12aea535a3734944b3
z6f7501cca661701d0eb5a5eea9e70972356599f4bf4f91a90d288ba69bb70f356579b1e5d8a0d6
zf78df44602fe196a1eb1dcf160a756bcd5ba62e4993a865ef34df03b6c9b38e270703f093212ff
z9e0c585a3f0a99cd60ab452614867f0f4c32609926e3ec972d82704c4c7ce7f6842b189832421f
zbd4d7abfed0ebe13b93c83c16e13732e406037a9a7fcf0e06a80ed6aa0917eb0fe6374c5637242
za99fbb995fe76efdfe4ab166305ef6857cc6cc9f331e51b5d0d4616e2cde307dd65cf975f53cb9
zdebf443cbd017a076585ced29e22372425ab0431447993b2fdb576847524bd8b4f06583050ac2b
zc7821fdc7a3f9c19abfec1116a3cb35eef9b97bce3be78f5eea5e65167b4c863bb651ead9c9dbf
z53c7ceea51077003aca7238753c95f1145510bd215208ffd3736f479539d46866b0b2c800a0a5b
z9654b20886d9a3fbc40d665f2276ef362bfcfc49e55cde079efff7113acebac27ab6e524721ea4
z41ce335d4e9b3779c491d1c2282f1f0ced5c9c0f4ae48c3ac78a4d71d88058610e1f61fa7a246c
za8f8424567dcf2a8b490fde570a8bf82bf98c8281b0bda47183fcf7c0b4e71550b65281db280f6
z389dd50e58fea7f96de57538efce55de5c26aa1fd3974fe18e5e2530cd206bf148123d62ef0fde
z6ce487dd00f7959071a5cc6aafb05502aeadd42d6083398d80b6eeee5ad9eda2be9c74b1e9c371
zc09d94f4ba5ccd9c67c9619e8025ab1e3981c6cffda212c138e0898ad06e8027caf3687ae1cd8b
z4fc09c45049c6dcf8adc796da8fb7c0c9113c20f38377d2bebf11928ad039b91ab46b5cb891d15
z67568686c5778e2df35bdd0557f86d2ae39e1c1e9774e0d1f6cb20101e5cee861e4f7e16277708
z1d3f2dcbb6d5d4e740a89c7cec0a839e2bc6e9124b4a956a7214f39b01b1d4ecf95b3ee4b34aaf
z4b414e5ddb5e0fc18145b2eca54b1d1e31df2f8b4232a3a351c65c9c7894e39f2da3d9c81372cb
za089bd186c655a5d04c25d3bcb2fb2c289aff01fdb1866e3fdb14d5e9881c5fcf5e94bf2e15fe9
ze0bc4cd17fbdc9e8ae3854edf98b5633f74ca2872899dc5d6d0efc05b1b5caed0a50bbcc42f7dd
z59ac67728afd9d31434830aca73bb8a00a1269b6c5222115fa4a31c835aaf198f4ba141460e91f
z8e4917d6e4bb353c1c429403b22a9dbcc8d939470bad88d3f837baa4cac84d5b08399ec13dcc22
z467e6d7b278624a31739837f43b0ad0914b32c303bdac18ed4e7d187c553f5ac0296d73e96aa30
z952068208364cab4fa18954616eebac9901def90ebb763daecee2cc0fb613fcbcc24cc7a0348c2
z0d2379dea4cbcc941d5a509b6964acea5334d361076bdf60c23c49da14b669561170c28fae679b
zf7811ae248d010f99282afe0bef969aeb4dcd0d53162cb9719bf90331ca4ecdd7c1b3e3110d2e9
zd5ab72b0d5ce9f4479e85435f4690db4d2d6dfcacbfb5664a6fdc38cd65bdd10759348234f22ae
z25e1385e9afbfc55eb5e91cd6cccb92927ed4193f2b1731bf4f01ca338efd2ec03f92440d9c5c5
z83321bfe60f38b015b9b6212d77cc7eda523944523a47a7196b88003362afd0c51cd1d502ab122
zca73ce28aab8e2608b1d93a866a2b9b324133a4fa75acbebfdd7b728febb264532c7a4783f9cc3
z442ace56b9dda632f4a0726ff49fb31c4a11f97e4fc15be51274f818462cac6526ffc5b7046045
z5e23eb2593fa6b29dca2eec6437ef33d95059d09933f53c6dae081755e18ccd4517b6b238e4216
z4956ec76f76f4c248f596356ec789d39f0ccaa56be49c4f22aacf9a73aa5a842723bf9a891b330
za7907e71dbe003ce84c708804a18bed0fa6e679f481d67a18c4d69cf5a131942ed2aa48228a03d
z2faffa8c289c0c90782c608e5d5c7eb04c0eaa9f3d6b854d5499857888bb160565616af23985da
zb284b0a742729610bad8fa0363f2b0b9ac7fe01bcb2b96fbc83d2015067cf972279f7c89a83ae5
z34b6ddfb27fb7dd40efa7af146ba722b15c677621c96d951da2a41f1eb568acdd506446014fd7d
z2b743105bcdc5462bcec04d3100e873b96d196af54e4c84a6db558f77539df45a56ba2a09ff035
zaace86d74324e564dccf25e792c02028066be09b05a857672f4fe9126a33d2ee43f5ec8e1d11a5
zdcafb0d34676b2ca6fd2f85780ce4d0f28e4a1dfb1172f0e47a6deabbc4323095e9066e7d1bbdc
zfe1a14c837ec247518b35df6006f5e1771b9544e471ce10dc40618955cae839dd5338b0069149f
z3e73fa6eb9c08a823ea164158957a28325ee5a8ebc2599b99c3169902703227141da05ce700e04
z04601370c3b839081cc5a82b94e670ca6fa75a1f0ed2ed117ab071a7872a5cf94729ceeec22b99
z09f5bd593c2ad84ffc74abd5ef87c7b40c965872b83edaad7a7fb8402a965f7c0465196dbd933b
zd6b16a283f7a85a6453ae36342b6ea6894430ee2ea2600c82c76093b5545c7599720412df29fb8
zbf831a8cf8fe131c137a47c2bab280051e65a11e949a5e0b2d3cf8ca0b74b19df326a04c1043ec
z6340af236b1b967acc92f709ebb823596447f6164c72950f0d73dd71430c31f46ac27d5bc5a2ad
zc6543643dcdb81ed151b03a327a466fcde150d70ffd9fcb4ff89b25e55b6e4d4b561a102db619c
zcf7196b1669ffe50ce058c59285f4459a6098e593eb3e8e09261955b0d41b067ec7c28c4b82979
z1d920e7a9b01aea9496a529512248bb12357e4055a0249b0343bd27fe048d9ba7b173aa304ae23
z1557930e5daf21eea8d0ee7dea6ce59ba40f7d44bbb901281144b9e938b3d1a93486f56a82cbf6
zf2e47968ff863d92b1d0ef838aa312412369231e8ca7c090d1dfee140e19ce2fa8a5a4fa5f9960
z5e16d4eec1275a36667a56aa769e4d3d2fde8a45017baa550371cd79a1d83e4b70b6b48ab9d782
z215eae7b52ee7a523bf51b274855ab088d547dc8b38d2b18da69e1acedda618de29fa0ecaffa37
z8577f1eb41a554388e536032b556e20a195badc771b17c3be24c6eb2aaa546662eafc4039c47e3
z97ab1704a0d4d3b169a8024f3a7e14c5bdbd0cd8524a92da829e2cf603f333d699da700248815a
zff3f6efc65026ff66a7729636ee7d42203065e2fd6cd233fc0fe728c4b1ac9c76c03d06875e5c9
z2e2a479716f9cc1f8ecf928a89348908696ea16087f2e42842c050f241f2ea8d52eed6480d67cd
zb62ed860b49a898b11b4b434547909d0eeaf98e9572e878a97274750d6f525b7c4e3a3f0dc3009
za39b29d22003540d9c7e3005158b2cab8929b5a6c8cff5fc92cc0ff80d31eaccf0da915e31f76f
zef4d6c0138f0ce9e378464a1789c0ad731f2942562c66e195ad97d95b1e3b2f0791edc6567ac3a
zc446a0f6a95bbe26bc3057daae122d98e1112e6d44ac5f171d8d72fb3e1ba5a9f98afa991c0c4b
z32e3405558ec9a0d2edaa20b713d0f236398cb356a4761043ae16cf7f477c2a5c92d1e31ab8e71
z70223a07dd8711b2a09185604178f8c4d26d6e848babac08553039606eb5404cfc5b5b36fc649e
z7b3b2e0709b813e6385db5624f9061ef1a64aed1d8f8d1c6094aa7a7a6eb2e0ca360f2569b9bec
zdba6629d959b77ea0d827d1e1fd18d059181eea58d259ea869219aeb7aaad0bf8e273734f0881e
z65eb0e4746b795b8a8c39b5d6cf87139928706468298307a10b30c0dd5829582ee6bec80df8d0d
z59c6456fa1861051e4016678009bd5cd453b389ea5fbd507b7cebb820ee919b0eb436c28470a33
ze12a5e829369092fc4d8639c5cd831053cea4b16fa0a4d2cd31a72d4897169a471499d4dab3eba
z96a5bae5ff6916811a8864e329cda80098e057c517b2c04781b1a1551fc82301f9b7bf53824468
zfe3d4ac8dcfd97c75c5f4eef458ac10fd04ea0b09e38e7565b536cc009db19adbac0f632a5639e
zcf0c9b406d28cf91486f125ea3ab0475c41893f0ca09e526e9703f8eec1f2f006f8b3865410128
zc25d04de609be51c73b03e7eaa1e58af431dc82f4e7e6dcb75c1e22f42475e004ba40833ab3641
ze045199ecf0e05bd4eca459c30ee2b9a225c7d75ab96a7e2a1c5a55573d5884a283b9383316aa5
zd9d8bdefbc80d846af6bfe08a68dbe293af72e99e5479e632730bec2589cb119ad4e4baf41f7bf
zd75064278c8f67c2b73657734dfd2c4a064095a18e2d28e80206325524727f90f273f3c4f2a891
z2abfd87532b2501432204e29e20d20867479169d80af0852b3bbffabca7e2e49260763db0870d6
z2ac4931b1d6463136f428a9bcf2582cee6eadef5a108eee522a850060561f348aaaca6d777fab0
z01504c5da4fe836bac769bbb86cf81b0fda08eef6136cd5ef7b1a431ab18d837c7c8bdda459275
z573f334c89d042a5cc59ef308e5778f2e6127fdb2289e4222d3b890bba48b119dffadf61fe94ae
z7c4c8d6f660a09d27c1f77fdcf69395af6d7c0e7902c65c51e3ee49b38dfb24a75c63b043263ad
z08e7c5e410bc09aaf3e1a8664779c556ea189f39e8a23bb02dc3a41be15d702965d3c25377ba58
zc74844da31c2177e0ca44ace250f7a94154776b5163d117a8c49af0980e1c758fc60e99c19a383
z30f22e70aea9ff279141f8ebffaf621bd94b393191b799ce0c55f7cf100e5fb6818f992ac8d997
za7215bcfcf23666edd7b0a5814542004ed274172ab451a7732cb87f8d6b60488e506a84c450488
zed5b3dde35f70539d5f6bd9e96ff55d5311f7ae4aae9850ff14196f25217f842562f7bd90c4035
z6ae871fab61f77cd8ec452b40b51c44118b3d7f9d935f6542306d06ff2688df9d8cc050942a770
z02f2012a10402314a90ce5494140c2ad2b0ad176fa5e07990121438d6918336c1176e1e6c00dea
z7b6482c78167bd54935fa04bd2fac5154df06a6dfc6674dc304611692fa3078b8b5a50dc4dbb02
z03848557547464c14da7c8aa1b0abbab4f585565ce2f8cf973c2a66585507e093b8a88d1e38796
z4121ea96a696b587785877439f9172c38b0cf64f4ea855675f7ddc65e435bd0f5e7f1a6131eae2
zb46d06db493959597b91d305ef06e6caf1f53302bedcca52fe762a4664f1a4e0c7b1b7e3c0e5e1
z775cd37192f291e4a683b50ba0c1dfd84a3a1d499e9c2a71a908d440576669c3fc4b2654b8da70
z4cd21a45abf6eadd9a9d52e5e9ab30d951ca1682ee395ee6ac4d935e48841a40e56311e852c622
zf2a9a81429187a4cb37ba02571bbda15b87af00d458225052b0c5a1235c2c9210000a70fda5bd3
ze0c0271a12fde452fde958fd1c8daaf27671766e31a2fcb316f96cb73bedaae575b0c267064d0b
z32c704bbc814515afae864e0aa7016079090ad8bb943643ff2b10ca5fcf5eb82ab97906da8706e
za88d25a65851acd4614f8dc8986a29de520614e735bf48d1d1f07afde01e3099c171bc4e141d82
z3e109f104522b3b696874319aaf5e45abbafe3b5ffec52455619cf8740435b7f70d5d63ab5569b
z44a046cd655ae68acc930b61db2872156de6c8ee325e49a3fc7f1b5b2b676881ee498c861bc7cb
z54618b8bbb9fc6179029a40ea11e7471e8f56b90fae681ff09e90b3e4a12d04cde26adf9db3eed
z8961b082c795081ea49d17cf2fa0f6950ef41d416b4f27ab593af258d9eac74a60a1560430c21e
z0bcf5b96f1467eac9834d7c31e5e780eb5e1c28b755ac8c9773ea5c46529cf590e8c8d4d3a115a
zbc7efe692e067b6ac705cca1b4239eb538d4a2052b4e433f4b72707a5e51944f57eb4522bc0afa
z0dd7e8833ef9927d79e2512891ec8e921bb4f3118bcdc6b36a95847345e13d8da2353c1bd51159
z7aea30173bbcb8924d1b4ea0201e814c684b7aa04f1a91a8d2f10df47473631b199168c222dfae
zaab80805f031fab34e48d0f7bc3b8eb33ebcfd14fbf5ddc35733a1e02cff6bd771f34301e09348
zbc02e5dd161a3d76d867e3afd59e668949ccb813c5df56563aac0b3eaa1c6d9bee06320bfc11ac
z7833c7042df30900c8f8d3cc87c7bad08d43ed3fc7dfa7790e94e13d7ed08d8d0f41b75df9d5ca
z3f384e55ddee9f4c3977e16d9059018762bddc3baa8b1afa257c9c2508a1545b458f35c4fb8f41
ze097bbe139a75978c9a51cfa43a8f68f2abdb7289f172ed6cec375f41cb27f0c4a0ad902289321
z4112ddf8f60480e92b31ba21ea1766fbbdc490ade36e2d0d8744df252159dbe4440b5747fdda1d
ze9f2e19441ce3d4b0d42fc22296e5abf5e19193e0e965bfda5ed2782da40c56f70bf0e3967b7d8
zb4be1e897f39a363d412ba06d947b856cb795024926fa021121ac0ddee4b5b66a06be8ea011ecd
z61493ef677639af41e36e923a5af82231401fe9851887df7fcb7d007193c9ed6569737a03b3736
zfcc8fe5fb71ad52b33f0a372133b959f7e4cc4819a96104a8d1203aa334c009a5c90ce537e6e05
ze7cb6865baf25f43bbdbe1b1a85af0675b25092b1401845e357a71627e4c053235d98ca94b56b0
z3bec7ea140031f9b710de850b83223adef81bfb8b35d8c35b6dd81a6b671b60419ff15c04a7e79
ze4075581b2a740ff3f3909fd88721b62474c585363a4496a615f7edc14b683d9f89e7f5878575c
z2ac01e741a82de5ecd7889a6de76e74092a1375fd93c1b0f1b3f95e5bc3b767b3372509d15dbde
z28144cbde0ff3afaea947cdb8b59ad859abf5abe4d8931cb39c20d49a4c495a98a938e06a808d7
zaa13a21e92dd7e982fc5a02828cc48a8c01ae8b822fd012535fe91337defdfc7600cebc474815f
z0a35e491ef6bc4a95020704778618057a78d1c16e0467f0dc8148797e2861e9efaa0ad21fc221b
z9f7877fe0ba4a008308f011557d48f1d97cc7b9fac80c05d652594f28c413f805ff0a846cc0dcb
z9806daa15a357c6e358d24daa12072a894e7dfae4f5f0d816bda0a58e1f774f0f103e81276d29d
zb621074fbbae008f25383218fb18cb305bab78702a0ba3e4253286b2923c56dba4bdf7fada5985
z2c862847a6f1469d55d321a54dc3f8fe9bbe954e88f13d3791ab324a8720c46bdcef05908bad8e
zea5cbe74dbd5cc05a8fa26e8ddadd653e121688ba395ebd9a94f340526ee55e4bb7e2be1182583
z16ecde2ab0d2da4a8dd5688bd6bb4bcfa01ae5ccff3b3be2eb0ac081a4225e74df50459006dd17
z4a0288e04b82377836fadc98f47f0aaad99f54dd8fc5fcbd2e40bbdd87a145250bb81a00bca159
z484ed41344942e51525979dd5b940bf5d9eb59b922b85fb043136b8b6d1c346b8b74bc69f2e95e
z2a2ab3cfc9006a20bc38979ae75cc9cd27db817f2ea1917b09fe9ba89cddaeef9c82bba9661326
zb4ccc8cb433f26893878593b321d8951e2522991a12d997b64c4ce7907d57df8d0fd3f3e70b2ce
z5702f931f860d2d8ebef8573e4fe84a22e7c4a5a4ec2c6c4d68b34c1787fa39af578e6fd1344c7
z843b9d62da1286e04935f578f3692af9faff45c1c27fd8ac8823efd1b46aec23efeebbd34d0455
z4c7abda29ad0cd01b0852f640699144c834284c185178c47d824d87c9fb2669ff6945514398e94
z6cf5e8c2723a5fdab6d6b31e6acfb6d7d722402e511e77c1b226d4c819c0cf40703f9bbbb81538
z06958c206a59b95d7cb80a779116372b58612bf23f10dfb3f6358b203a3115c58d2d5f100b15d4
zfbb579f21dfd5e539afce02b8275852e62f53289d03a2c0bca3a3e6678ce32af7d6369a04ca1fc
z8b5869671c310de75edbe04c9227f0fa9fac5c1554bd0cd21731f3d497e8d88fadcec5b0b85b27
z8aa3c7836a8dddf446b375ff4f5c0bbb538d202b0ebddd081786323997c2957fd3560f644a24c1
za5106b0d813971e70abac1b30e56bfd76551da449f5182dc588b94837d05bd20f10d6546d7399b
ze9b9f5595af68fe2bf452c3c17a51f3dfb44ff649b186a41846b4fb82b81ee8effa1693a246780
z4b2781eba14da4916c4d6f2aa41cc62ead3467eefb7f9a1ceabfc887eaa342360371914f3624d7
zb4df4a592d0b2f62e117e8479c416464e8f542009a3f883a1796c15a22cb83d7da0e5e1a55d7a0
zd6e6f9c5496875e112a49f8516507533c5751052259aa1defce33b90e0cb7936cf1038e1fcf01e
zae322179bb2ee785d68fb033420b75685d947d8d6fff382aa208ea72c6977bacd5302d6098b795
z01a211ffdc1e9eab14ea09b69b47bdeab283e9fe06884ce01be3b51804b1ab4701698296425488
zc4fad8b91723f3aa4646a43652f166de23d9a766e7c20f6d41e03304d97e9e5356c8e8b1591c7d
zed91f27af84730e386d51e2d36f3001f99d36ed4060f84926973f18682094a94783f0c45ee3e0f
z10168f857ebb580c32e7c77878d3e4a97146e3b42251fe791ba4c3bc032eb797414a5eab0806a1
zd2ab9022236f8c960f20860d8c3d8b26c502eac19270f3cfc25a94fa2bbe949361bc375d18dd52
zeb726b789c18b3eb37070db43c609257a46381d15dd4aff246e67cd3f62e5ad9555298a3011d48
z618d72ecc71635b1e45c90c6071a547569d6f83458cdea25e3d548583923d99806bd4ca11f00c0
zb6ee608d84aeb66b7e21dfac7b80ba809171746d16fbad1bef93c854df982c2b26c509d6e1c8cc
z25facdfc56c9d9d7b40c7355028d0347c3ac8ab47b00c10e86f4b8085a5ffeff47ff7a8c71c1ed
z78cbdc3ef5e433a101cf5e75654382ea5a9dc817bc1881f96ed9572aab682923ac86a0601de24d
zc66fd71ce45d057e61b209cfd7e465239261cfd8bf80861bfb20b808780dbfff5cb01c5628fa1f
zec4a398187647fde6eaacd1365877a71b0f0caa2d2e6ae826702171bf8fbf8e93ef4e169e48e86
z365e73a3dd2e0a2c77a457631e46924c02b49f35eb4efdef55074eab16f6a8025829b20dc354c7
z4cecd4e5835bfb2ee8d59acfd0f8ea2a0c9010d8b9e86b7d412f14fa3bd615b0c8e8093e8069b5
z8995df01efa7945d24fbea6c69fd6f2581298fca2fbfe6e4d8b5295b50476fbad1088201e1b1e0
z6d69a3ba016e1e3d01ac0af6d8de13aeb71e732ced18d4ecd8f5003ebca8d286850e4904c0c08a
zb5096ff114a5db2b7d199bb15e55c4166fd3461070ad55e2bfabc3f62dbdba0c8ad01b900aa1b8
z4e181ccbf78c8336f44ceef2945f5d93303690195774bb5f4bf8dff372192c0fdd53ba4259c821
z277740d03f58067a489e79e3d6c5db035c2c8dc88d27e2f2a57a12859b2dfb35546cea3d998bb7
z0ac19e3f9ab8056c6da6d684bf88e8bee258d037dd654578d27ca6c6daaebf3f03e0d019d85783
z1c6eb1d314975c31c192e712c69434d7f306eb5dc47bf66f6b8d7fb244214c124b5765e8d2998d
za20ad13eedd17e45f0667c250b3e2184b5b3d5b6dd4b5b9f520daf5727867cb8030b64ccabe45f
zd78fe22df98cfd86e069e9f7749b37d0f06b8fccce7ce7342ba2a2f34c64a1321efd759b07ea2f
za2b4d8a4c69bfe00b64c49dad0c795d57a2229f04e30f7e8c6b8e7178a90c24b2f87615de71bc5
z96ca1f1f3f4281ce370c6e8afde6323ce2f6e745599366000b1f07ab983c703d2a2cf56934ccdb
z0c5103cbc5726cb524aaafddec165a7b8a4c3bd76948734c606d9c6c196080b0d469a3c3fd6068
zf3eef80d2f20934ee5277e9485520f1d7aba7ad75f44760367bc157cdc8f23e9c034a6a29e03a6
z5cf79bd7ffe6f35ee9d38c6b86a4b8fbe63068752d82393f1807b735aae3305e93861553b6d619
zde96f20b9ad2c705216b8216db0c7049244c2ceefb13571e6c8e8e350bc1789ec93fd48385ec6c
z893e32c14f78d5eebcdc2dd84009dd93ecf1211fc6349281042204d20ccec3c1c2aa18ee6d10d7
z532986e1528e10ce6af0856ac996543dc41ce682df59feab88ce882534dc09a2321927d9670ddc
zc48ab1c01cb2ba9666e036152357ad1ccf9b03b60be4d5afaa7a6f517b90e5be7e8d78d9b60742
zf40e4d462bbafdac859b65a9fd29cd58325a37263e7dd417af5d618afc23e617a98dc28317cbf5
z8d995f7fa7c0f45d8419a44ec8304b6b3580c952747f505a5ffe6b456b1f858fc3d9aff6efb01a
z97cc06e47194aa493425135a572c92303172b067839bd9806069b7700cfa9d03105764f9f0dbcd
zb7a09fa15c66be72e9d34fa955c9765a7a077344a9904ea2614699f1de1162f55f1d1bde3b5aa6
z59925ac72c08508401490b42205e55251dc3d1b8b3d0cccb13fc5773281f53ae2f95e061429b09
z53f09e97f5e9dc35eff9f6e72ffc64e5057136c6e35765c074aaa0bfc42382e189cb3966638748
z0c1c6e1a0a57d7c002d56c00b8fcc958a07b24ce5d2e67c062dc40277bbd83628447b558dd4e06
zd1a306d096cd5d4665348443e805eeca7ef317391e1ae602030e74acf70601dabccdfd61951c8b
zbd88d050f14810651c0e02b64d52dcae0d151702dfad7f51774c14c9a8f2bd9822dd8c495d54f2
zaf886a6ea93bbac6794bd1850b5e97cb2371eb44a8310b7fc351eb229bb08581b2dc6e4b96472b
z206c2a22c9f46b3b7a49f25c1fa24fb7683e7e3614faf261d62c76b9c17c84ca94acd7119b36d5
zcdf05b528a4e1b80f8297c7c01642832ca4a80ccc3ba5cca8c696690c8d71e246459071f41c9d6
zb36d42d3c613c576ffcf8c9d736c1b53785b2bca5ed24d0eacdd6abf38a7d451d4f9479203bf32
zcd2f703e9d13efceeec4ce648a13e93f09136c1a597183a311735b37aaebd92501fde9a08190c4
z4d64432aa8380aacaf8cbec98a05334528df765ff996bf53eb2957eff013e7c402ff308619f9d4
zbd8fda829b7cd92fcd54995b2bb69142ae3967eff09425ba87c002d7f2debc7ca735c1566c229e
ze348433e4066e3af6b3ecc21c7c412e7e90e81fef44ddd815c651cddf00a1384f60639aa18c940
z26c15fc6baec3bef8d92302ce46acf2d35c7dec075c03b0d03b44f262bd5f2a5b6fcd50b9354c7
z141564c8989bfdd3148b9cff8e562924f7be7f1de272f077bbc5b03dc4c945f7463721ad5cb30c
z5e2c2db8ddcf0ad5e929c759c7c6ca7dac546545a020b838d882c5e07103181b70e4c9bb764167
zfffdd9533c5a03f76c66c82825eb0d6c5e5fb179d0d1f99c71ce89335d77b8180c5d2447472699
zcaa3d68a48720a93333b648fe23eeeeec88a1a8ff93ed9b428c25701f90e41f70760391c9f8956
z1b839b332a135b772ea012bcf37f7c57e9869c113ab8c649cbbd2eb86815df44c365791f1bc739
z37a57307d2c6b8fc391bf497e519f954f5cd4c5aaccb4b56eb1a0195fffbce9b2de878eeb3b13b
za9a16566bd8c3e7d764a08444a8243bbc37da53fd2a7d3c63d9c8c8f65f6483995b15a81048b78
zd2a8ee0d7f91fd94c6edf0a71604c64a6af2772c1f9e32340ba64937a75e25c4857dfb650326a3
zf4597e71f7d560aa998dc107547ece6417e2430fe06d9555ff91b451ab9c73802c1895dd3e3514
zfeb2c9b5210672caab44f402e029b16e1b71456fcd57931c32bf6be735148216a2269a95a4d72f
z7764f66429122102dd8556c027cb9e925af80a372ae32179ccd81ff54f823f2508b355a4949532
zb7649a6cce052c8b7f533577f081f6fab66aa3bb34a31dd0403f07cd0ee277724f6576dc3182d2
zeb10185f6262c54c4dec16c91ac88a9a09eac42952cc269b6dbafa6c9b77d9e62aed08d871ff75
z7d55915a75f7e467e25251fae2ad56601b687d870771f7e9b56a2117968f0e14052e7e4a3dd992
zb0bc7ed91488e40400350e9a9752272f059e83b510a3aeca9edd400cefaff33ad67a236b9f4d93
zcb0d97178ab9c69b929e68de87936f7921222366a245508a06bd1c39706894f0f96b4bd60ab7e6
z5e53082cda7a029a11b4c00fb4b5186d302e92ddd9129690d2c7f6caced87a1000ad26504b65c3
z847fbb9b937eea6f00d954c4c38d69ea265001b7abfc827ae7f840be1965bdc21fb7ea8d958e2d
zc83e09fe070ff9328972dd41eb7042d130217e2504a9cf7a6fffbef1116f7bb45c4fd67a4f259e
zb2cc701b0b8d38618c7939ee301f039c6ab9a92881b0f60ee5f7a7f14a18adc14ebb2d570566b6
z50d844290fa18a3984516396262d28c542093171fca53dc7b906cd24e78e4fef02191029255acc
z16b13cfefba82598a7798ec865d38bfe97df24350d9f3ae39de55eaf25d065764b9f6436cbfa55
z59b4bee17fb55d85114a952e4efd812ff5de632426604e7ec50c762fa07a55cf606eb3a14beab7
ze6199e89d749b0d8617b47be98415b540c7da34bdadb0517599f5ab425185160b294d96962be91
z71d9f784ce9f2e852a7e06a20a149c7c3c3cc8ad4b2fbb057f000afd32b7f87e2ab37f8c9ebc10
z28ea85268c23ec1c8e6f207d33fa0946c82b0208ad5e234ed947eb7a0e32ad21e9987839c998ca
z5f5a9851abbbb2f74ee82ddea0af79f790c9e5f50b5aa0f6507cc918d23ee1f25979e69dc63c47
z473e83413c62265583acb955d164ef49867eb8f8d5c15f9085ecf1a125efa391c600e7d7fa80f1
z1120a967e2dba85543b57c34276aa127925c5edce8b84437a71ba1aae61830604b29aa4d4177ba
z6277fc151dd4bf90fe0f4698ff74b2619b5cf7b54e8cfc92d55906c5c8914161f89f122a46b826
zcd1a75b535f367d169bb45d456292893c02656a8f76faa8567a25185341a70ffd7a148774c573c
z2221f9baa2c8c16ed59b69a8c76137ff21ff5564358993569da66fd285c5984f8a36a78b2127f1
z94e0ae16b8b04e6a005962cc697f23ac754950174ec42ef0dc0f49f63d7a38fce2f8adcfd6f791
zf7bbbd9ca5b8ef1d2245f0bfadb3c39f7748f4436a3c19aa6a9525a25692dd1c56ac9cd5a38f7a
z40a47c6dd5dc127eb17e1736e9ba9dc5c0d7ee502eadf2517be8e9b4622f5e4b8da602e3d35ee1
z17cd63d3a39ffe32f91c675beb8b4621531467fb976b3629b865e90388d2f28202cf69b351ddb9
z7d7003a673fa2b2e629b9dd7a2a625951956869eb0f57db98bc88e9abcc496ff42cf89bbedd81c
zd992e10b9840693bda575c0f2f5a608929f1532f4067c52db52602c941f5b0341f22a5bd141863
zbbfff5b763e9d93131748c283d4206a1d0cc58d8126dde8866b6386e8309606dbbd1b404162947
z539a4f9081dd58babf2c8bd6695a68ddf85cbf202a918ed13839c58a20ce5fb71a8271aabcf00f
z6b09d8a9d1a9c0e13671bfd38e44264d3585661cac3ed2ab396af4b76f0d36fe230f226fd438dc
z195e830c0e10443cc15f875d5651c79f4a98d0041a20ca01f5bda07ed9b0baf87bce6f495b58c9
z905fa9aed245b00ee461c77391dc232eb56df62c9f24f786aff96508fb404d311e689d4386235b
z992ea0d2be11be6079e5b3c08db1e996d24cafb4a33d2bf739f90b9f960a9b3eecec4e80d9ad0d
z43d5f67180d9d4a1f3b14838651eadeea217212f45f71de12cbe7087c6f8ccfe17f90410b87800
z4c1b1e87799f63f5cb8cfdea820122163b5a90427293a000a24144f2497442d532ed874ace5e50
z8b9a7c418e4271ad6403c4674623a1332fb990f4cdea333baa52c3200325e31b71f354ec17acea
za8eefb67aee48ee1910f8f2ed083d242c95e96b28a0daa7eca460ac0dd448fbb2767e911311320
zbf83a3b015f38635ca10b1733d17b8d36af52f1f18cdbfd6bd422610f9bdcdd51d05f2242ed3f7
z855ddf5c5b81a94d03dd9f1ceae3ea0e02bd094f3a9aecb6c5c28371eb39faf6288d87f2262638
z12c201ba182e1ce604da30e97771be5d20f90dba23fa4b20d4219e822cda1be340f77197114a26
z522cdad9e71c61affc4647e018253aee1b3ec189fe559ae0f71af9b06adb5f7d9b7b5df55fdd4b
z3e57579f1e40655ebc88733a8900b10259400f9fc592ea189475a0ae03d6ffdd72c2d4ed6dc920
ze23a3c680a1d57ac8f564f4f8edd715ac97b24a470d57354b64e62fcb55e95496e5ac6023d5fa5
z57e75effe816c7e569e234c5aaba82b380da86b63e4e018aecb7435e0760493573176a3c2c5311
z4ddb7e2776c01de606464121da07da945107618a87fa16585e57b3224eec88eb62bd311aac64b3
z245b83f2cbf468cb9e6abe996dc22d6d18ad60a2451971617f9242a8b9e868964be0c830efb73d
ze7ce1392806d308beaef885cfc65d10e15b84bdf51355d5587ea8a19a80e7d90a9115eea13c0f2
z40dc8e0e73023b87d2ad7c433cdeba3c6501a3bfe7e2467d0c4abd3fb0fc3db4a6fd64cb92f138
z11b0d6daa7a3b2da1079e887b4d9d7bb686d9a23a4d674b43b464fec616661920c112339884a7f
z13e963de15b02f41c0b553d91812e7342a14b657a0a46e33c8d85f8b6d7e4bb05dbd81ecfe2c3e
z4de15801f44ab285022536eb1870c36cdd97b9b739e5a00afb14ce1f8c5422b9177d9ec85b571b
zdd3a6e5c50f89791b1ecf76b93b2e4bd4345c5120b9285081168f066b790d13f5f4c763b7853bb
z94029033b688f4f560e1f80abc38d17c6a2298502c45792fc20dfb9ffb846505a9a04f147b54c9
zc84910ed6b5b1efb99e587b398afea2434c6894b33780df669a5c69ee953b093338154b853f4fb
z457f232afdcdb5980defa51fe3fca523216dbc3ef115869a351cd8c2f479e2d9ced310765e6697
zaa807d323027dddff82c8df50e958a3f6d11a9e89d33eebae99606b5169e5c50f31bc3e81668e6
z82387b9261428b9c759956b4e0b70048ebf4e7d5cb474bf82ebf1559afdb5023c5ba2bc974ea71
z96c2e69382a12c6f766030cc2c38742692b9a532a2dcf334878ba2725edf282d08edd084826827
z7af8af40d96f3a2ea6cdbd9d7b789c7cfb547595d75262dd465493ecbdcf735dc8311d65dd5bb9
z5301b4425cf8885013d0fff202276a13bf0b81360de8fb6e462444ab20e52cadd2c9bb8328b8ca
z62853d5890db762570809bb0ff05e5b0f3b9ceb42053bc75fccd258bc95593d01b9eb831cd350e
z2c0c3ce797422f557bd2b2f40289cc7ae0988810b26dec1048d53dd00c96e2fb40a0b41ad861e2
zfcb52ca6c7dc344f72b514568372174a98380addd65ea0db78c2851a13f4e5a3015cf04b24eb2b
z4b476ec6131760de51e1dab3d45e86175e5efea8e9ad712ecede10e27df38396dc8d2d304f9805
z0371ec8c8a44314cb9916c1e523a066d1b7027b1b3ede58fe546f3cce4ad7e73141e4e75cc8df5
zce372dc8d3a171ee8b1c8b8ecea47763ed685d5d562283f78e4cf4f9379eb0fbbb22dba3790d3e
z7aefe797b7be391f240b5c01409bc858e88a91ab5ea1fae1c10bdd610c286e4d7e65ec35c05be1
z058fdd2732e133c9513395e07a2b173badc572246f7b19baec236a717d3a33935365919721976b
z23c85ed9984b72dd2415a60c7a96878d7762ac35ea51fb75f608b7090238b121c33bd416b67b7d
zc615dd0541d1ee55b08b08fcecc9b8d332faa7b0a56b97e498e5c673974eb74f633d5f67020cab
z2fcd98c63decfd4f69b4e925a7794ec457e758d125703e42dd651c2dfba3a07d98e101719d789c
z85a305491b73b813c789a4ed79e2f32c49f5c68ce8f119295127d6232c10595ce89bc518e60035
zb5936264143c1dbf954d05d94de22604f070806cca8cf04e6d4bc0a8f69a6aaa094a463b3c8254
z76ba7fa043f967c30ae0d22688db732c26fd01a5bc40467f834b23ed3be49e0f8fe0bf7a287aef
z856df84c7dcb0c547d50b0b5acbd5fe378c80db4d79e3ed35a23d175030b5032b8720de1d98c5c
z1f76c9f939efc62e1243ebbea78d010c5ace4dfd85e4bdece69496136a769b1c055e42f29fe5b7
z98f795bf93a524d376bd0ac6894cfa8f0f094934e55662c98fbfbf4c4fead884888b1ccf9d43a9
z958ba2be9860fb0b356391f49c78ad0e67fab68107e1942443647a76d3055db77dcd64e15dd4fd
zfb0a09b13f036b3fc1493841969c06066f011df3607a956b96540af3b4c1b02f2193333997427a
zdfa8738548cd79895ff72f9c16c037992a331b88d294df3f7172c24aeb2c1a2d9f6f37d16e7a58
z664f984ceedf91a5c138b745e184171f0f0603ab38f0515d7875b72544c9600557c54e729fddac
zad2050c9cac90c8f3f6c8af427ed7a3b8abf1be33bd2fa5f12501af14178754feeb52f6545c340
z8a262a14905af48037b97853b0c4187af179e2b7267a344b95576550751139db3b059cc1e6a7e5
z33f8483559f0a042a561e7ee05c35efdf862b8ee51a89dd53d4e84a81c446fffb0d8c55591ca18
z95a19cad7c2d73e958ade780e748d468d566996c11c0dce0f74c54eb4f450bc5d15069c558cfd1
zc7668dc927c1d5c95e2a5ad6a0a395316851a941f3686516b66cba692324d0d0936b2e787a224f
zea07d0fef66a32103aefe2395ae4b359e206ca97961f21ad9aadd3687b58549d6f3d6108dc2dac
z5fe6b2dcc7ab2103fa46e9ce03bdb8e04c2d8d58c7f5cd2379f744a7bc374fa195c8dc155047a7
z4773055f87ce45892ee3c2f950f9a48f1fa3ebf5101b71b8284feee30fac470352b0b5efde2bf9
ze3648509fd1e1e7826c0f3db2e092285c775bf3d41eedbbacdc36dcf0cbac64e0916e2c91bf15b
z434868829b510e1be4399378fe270caed49b1833e01feef78b752d43c72a5d679561b57da1d80b
zef989b7f441aa036ae70af71950eaa1934bb2248476d95d4c0b56e7ce1d32c3da6a497b7d946a8
z72c629428b750286868b06598551ca43e586a58ef091537c69ebb4660dc0647facda74bd53a4ca
z67301ecd57a1704cc66b6b33dd7e530f7e5b68e2fb66b90c89f87d2c03f47158b403054bb614c1
z0510b76c10d76ca2d0dd172aede253c59f6a8144792b24c82d7abc27b678fea7a50fd68c77c9bb
zd622246dca53fb32e999b432fcac6ea85664d8c69b9adeefebaf59824fa467ccaf9ef535dfc6dd
z14d8f96d55cc09acf3fcb58de18029c9637e363e078530461cccf52e59f90fbe433205bb9d05ad
z801d9a22e0055b20cc7e1aa57dd8eba67d37eb2f5d8714f8e2f989ba286653d460667d6a845bf0
z951e29373a5eec61c6c43a1b2c169a5e8c0a43bf04d0d5a10948223de8af2d64553561e8be969c
zbacdc8e390af779eb52d414df26e2d9a8a30d6e172d703f4d9ff8bea02f5cf898475f3d4ba432c
z0a45fd477f8c736c8e589f4174a17d075032fd0e122058ad3e57cad64e8e1940a8663c079854f2
z29bfa430c30e435085d5ce1c460f0988ef96f4e17e4fb5bccb1bae4f05c2d3323b0a9ed61986e5
z49741b3d41f677762d190eb461610b65d782fa51e082d6370f732e1284bc0db0d86293f4abd5de
za5aacf1ca2674b04d9a5af16631828121316a2993c5f4d15a3f444e00078182ae79e6fccf70605
z9a1090cf6ac3919993e534d8a15cb460ab9e47acd9a56131093983941b67f2e2d05e7a02a94669
z689e3ab0b8ae010e3fa6b832f21000c8533c4fc4f3278505c7d54258f428823909e87a924127d4
z36ee8053e125320c59e408326f2a0c8143ec6a4dabfbfd6de7435064671aa558d1eaaa773b71fa
z2c16d52732b3d13a9339b651bf509efb17571ad50eada2d909f461c41eff9a1d2b6244940a1e80
z9e582494f39aabd265021bfc7370a4ea3f009105f2ae55bf9f1533359171df093d8eee91ec9430
zc84085e743d8aa32d935961f74c1551129a2bd032170ec68d71fb6625197ee8466d281e294d475
z0d3976378e1e50129d1c3eebaf46cffa0d0d91a01a391848ce68f3c5342e9863f1c48ead773b09
z5b0cdb2101ff94f25d26ac388e1c5cd50890031cafcf560e0a3b508fb80e786c0066737f8297ff
za89252ac236345f7e13dfb4a88c2d72bc0481dc23269208880b3fb5eef6401ab1fbbabf7aaca72
zaa04f45b01a3488b38a273ffa5226d632ce9a1adc981548c11d0dc15e0d40e869c382dd31a9e75
z2af05a4ed738fdad929e772ef358b044ce4c99fe4095ac55e9e06051edabdd8daccc1dcffb0007
zd274b81763e5a8783646547bc2b73f55e9b301ae7406aedd3898cafee9d073b3da7d16469ac326
z0a72106f62ed208f7f06f013759baf3e9b940220629c4ad5fdfad4e436042c0d770b3b382b9a04
z2a7216463dac1a829b1aef7424e2d25878d2ea3cd1265c2bcc555bcc9d908001c78dc198bd36f3
z134f8fea92c92d979dd699da02780f88e5cc99fa55f807ef90f043745b88ae56a9f5f06f8b19b8
z06c187c2019a66902f05dd54ced26f58b739fa1e13c853e9703c8a0a8f911874611366a7001e18
z02ed4e16fbe7686bc07a4d8062f92cf65ca02d9599d40643a969d3aee1c6b8b3b47a0f365c3c19
z7a7b690b404c9889038690721df01fb5827842ee39968173e2f33a229a04b5cdf12ff751391ebf
zcfdad0aece35745d56e47266fcda0b1f98831858dc4422d6d5332fab0821a3b904088bc94062ee
z24bd1d7a0f77af49c4e03e9479981c4bbd134243fb845579375f08e57adabbe7b63a3942aceae9
za7ed35b086f8d49fef3066ae9cf7f7a7e4f74870eca6bf27cb165b605b0cc87e6add5d9211cbb2
ze67e78a2943728536c63cfa34f00ca9524d45177326736a4cee17764c6cdb2a4351d10aca2f06c
z9f234ac13463dc7af0272d9fce176fad14e32b50b6d5ad6a098b7d95d8b5c5b6a70c62af248deb
z7646602073ade7c11ec414b400780cc0127823429f6bc408348f91d2d13debfc43850b0875772a
zb6e17c085f13ec03c5ddd88010eb9bbd0eaa22b7561b2277711f5be0a37c06123f4cb194646eb9
z34a87aa1f3885f29a5471b48380166333c247b7c34dd91964471340e169827bbdc7b192a5eeaae
z439688ffbf3544dbf7357c15251fc48e364569e9b20b3af411cb150df33558f509c1573c5a79d3
zb8bfb2ba852dccb406fb3fc8ca809712b0b338970cad9e5cff61de9d3c09409b8c30c0813ed357
z941d63ec7f27ce48356aef07e43f60a630893877d92abf1780d6d0aea31ba6804a13a743af1649
z5f378fad4d1657f3917f9598c6d9079427076103f3f7e55250bbf511e3135db003d75d573b42f1
z129f0c5917ee95356402e423d4934ed5e88ff04f1b1bb309e2a49638f37c29006bf23ae64865aa
z5d8742beab7d9fdfa0da8a63ab554f5795953a05ec6b652f2921d5a1d8e29baa256e96a03afa0f
z7327c080752ce741368404ee060f95347f6b1ce52d30055f0a4f5844eb61ae4a88cf9f6e0eac64
z7d448c5cb94d32da57238b38cfcf026b66e16ec70483280b7ba3516307389f6e655854236f5df8
z0d389281d91abbc9ae9e280eedf2423bf355edc22805b8858e789e7d8f8a32621144afff19ace6
z6e92781dfd6264006986eb63dd54ea0e9895db8545432765398117eb78c578c071c3a81ee92591
z328348994a47cb523e1670363644c6874e0aba98d04130bed6873b0a493688b1c01ec35c9dc56c
z764469674d13c70d85991888bc30cfd1d2d4c2922a792895fbad134b6570c773d325312dc05a8e
z603f0b637f264cad8bcb3037edd2832eb031f465636c170ff4d46ac1a311af4c9f8e3a669aa28f
z4c89898a942a532460d005c760f762fe85bc259641bad6d5ef5218cebefe46eec5a2f20c6e7d64
z6e2785a27f526bd53fc80100a560e407d372c9248875f628ccd88a8628563625a82cb53647d30d
zbd2407d24bba763e7c99514f92d5d9cb27ece955e7ef25cf3321a77f183256a754f7ec269b05be
z39fdcad5c1c0d4315fddbfe3c464fa02671310d50992c1d626d698273a0c385ded995b1820feaf
z4cf5a618e0728c3e17a34154ed5c9a8fc4767894f4ea0136c819fa52a6bb1a5074949d6c775590
z428619efc2c1640e5302176b02cd1c027515c79a7f5a64a0fb8a9756685cdfd8c23907c14a9927
z8ab11a8e5c3bf92395a4e18ccff04c03a960cd9eea94b3a75fcbc3987e03bcfba9d1f2a5c5b24e
ze621d740acb947184a58dac0ed1de3feafffefcfd29473f3b34ff6b754044ead9c9172e5a28ab3
z6ce2dc7bdc623838225acf57d913f8a2fa45ace2c5db5d81a22f0351df6f8d57d4452f0f1755a9
ze4a64f683752b422a895769e89693ba032ff619dcdf87a35c64445b32d6ab0ccede23160003f1b
zdeae7a28b9d116916d95b2b09a4820ebf877cb147038d91b174404f29462a0f12867c2ed415c6b
z0f4680fd5e98551d681900d1c0d862480f2ef0ef1a1bc7ccdb2913de5f31789e3557b838151d75
z8d03ff69fbe608a29a6a975925e4ff0f77f98e9591acbafacfa60a0fd09071400a083ad9a60160
zb7b5d42ea879ecf101c9c2fd3ca1ee99cc3411b60bb0b5800fc90177817e441d797075753f8ddc
z4c6ab0cfaf465cd51566a740fd026928e75c17354f32cd95644c919cb97d65dc96c5405f10b52c
ze4b09741fd9e5ff3a712f4c01c82a371274472631486d9b08418e60b9e1c72038a07d575ed1cb5
z0e605a6042627432643a59f35980973431e1058c04fdf728006a5a66a418d8d73d26a31a11b23b
z85d70b89d734eafcf08e11bb6bd23568273f0f4d3e4d31b6f2d43b6741c44b2c38a17ff79e5577
z0cd0d98657835945a0d950ec875fc1fd2632f4714ccc6afbcd664cbad89955e54015648acfa407
zb0e0c302ddad818c5ba0fe2a2a9db2821479a328466c19a2f641bf74c8dc47a391ad0b685eba39
z027b62cfb028a472ee01dd59fafca35f57f5660541fef3f60efd4bca18b90143793a5c48f3bfa8
z2291bc54ed2217e652c52a8cb229f6bf236fa8113638345dfbf13cfe4e94de27a33ea4782d26fb
z14b393df6e211527fb50a48a7f6f72d3c26da483ae5ef8be13e770b5665c96f3a101cf7104350d
ze5e0d68b45a0b2a9cfe96359e84731162f858506b2b2aa2adab44cad9910f916fb754ede07b212
zb42fa3d9c5f5035273ba827030a9e5cce1470189c146813b0a81b7ffd883924102628d0c94f576
z053e95d0af539cb532026586c64762a7d1149436543b11d5097953fe54e23c961a93a52fb971e6
z2d6dfb4313b3f35960d36ebfbbcf0691eb31cdccea596a567ce4c44833f6a8b02aae521a985edd
z711f2b444206d146fa8a019e921dec127ec729a9c37976b02efa1048c3f845aee20e31a78674f7
z5366c97c2162c3cca3e1418f8a1e12d53420c1b9ae797ac9ef65509707850494c876a01a737b8d
z6de787e7438c03a082a9403dcc1d1d7853459f34e61ff408dbaf7b083fd00fa32c617061c57f95
z464462f6480d2d9ba9c5cd8054545b9a5509e52ca4d5787b6f7c0d82c36871e38f68080417766a
z4300641710130454caf8609e7fc756bb75a4ec76083cf140de31af0e86d2814072ffeafecee902
zbd88afbac45dcd7acd1a7b7d5fc8228b422fadd082e7886d5aed48ed65dc97d26a43e4d994c1fa
z314e45ec7dbe06a87bd79db4675f7f7dbd348a2709858350f3a51d6292fe24bf80d91d72c1b069
zfcfb1571c322a21f1fabcaba379d2e8e1c5a70f164fc4f444e8eaa9e538df5e871d9856f3c3648
zafd5af1cf6e7a30856f1ea6343ada5b85523327943fd3b018fc6f1daef35b5402bb1e9e0f93efd
z34f385ef41950c6e7f975c3045c9b8dda2c1d7e769509ccca6342142d9251493af308c93730471
zc6d3f87d46c261466dea10fa59fd683e0c8e06ec6ce872cb5088b79c55f2ae63231caacd1657fb
z5956eed4a57b48fd27aa92db6f0e4891bdd25d19e79c48f5a2edce50b1c8b6b89af27e90b8bdb7
z4a1efa8f7bd4aec861f4209ec39beaf7bc3c0d42888ee268682aecec873eb1a973e73aa0eae653
z1e0296c594f0ca89e95470ef8cc02dad64c595fae324f9c37305d1607333aa1857bc7b110ce4c4
z0d2d94e4ac9775170f5a8349f75ab1c4a8ccf9f1f78d1c3ee06c4abe31bef144880177dc5bbe78
z857d50e91a016413afcbdd207d453f259250b9b31badaa783b7573121a19237c2acdcbaa65c1fb
z007f5e68eaf6b2bc19154807bd9f7370f8842fa827676b8a3f7b16f9c86822148f408db6175f0e
z0717fc2ac349006f62b230a229516e2d9002df4c25b817bdc69acbda0a86d173d26ca5729bd7ec
z1dea6c9fee89f900257c671b75e0ef00bee191f2866e5b833167002666b103cc9302c8d08dd1dc
ze4490de8b3e12ef05b7ba883f17cb30beab77e4e5bbe73998404807c290eba1b95d0174665145d
z5e1ff7fba1f290937a0cb57577ce820be89c126a41ac3bebf20696e55bedaadbf25c0912808903
zcaf57889b2520277724ba078c3ed4444a35ef5f49f41dfb949ca5d661d775c4ad682a5fbfd25fe
zd96d8a9bd3d0ded4a408cc39bd14fe080742542a67b73f4859a0b19e17dd441805fe4ffdc6885d
z45ffd3fc1db55b62331eeee67319fb4353a1cc1f9ba1dcfed0796a8edb8c4ffadd1a2dd43fdfe4
ze4cc6b69eb5f47225cf6536a88360de730856a67daed19a21aabebe0e759880badf365fe41b5ea
zd3277bc71b368bd390fc35ce9bf056315d3a29ae9226c64dbece57637620167dfa8c663718b912
z050d4602c580e1b1dc80b6fef67224ff6dc9bd2d1207ed92bbce28574cb1a4896d922feff6c3c9
z5844d24b4a0d69a0c0c0b2cccd032b33b13a471d4ff59ad07c239a045153bbceb2a9a31fe81cf7
z7737dc6a512c127258e08108ef8ffc674b060aaa93cce32719eddbcb4205ea55e6e4afb39972ac
ze32461e695245c2de0980a2bd5df4704a6fc002551aad255e3b00a79d7cc808435906b7bf5f12f
z9661c3259cc2ae1b085e3205597167df2865e45381a5d0032f60137f2d8162958ee0740d0dd1b5
z7ff555871812425ced8f714c5e8b59c9895f4a59cac3f88906229e177e73178514bd72abc7eef8
zc18aaf27be7684445c0a9ae7d9dbb2881f743d8ed9c9d8dfe74ad075e6ea64ed954d2677c59b44
z242878e54a51c739dc881fbfe8b13ed23d065587415b5c7eef00d5a4c853de36883d5c59f24b90
z11a1ab357e971335cfc849d94b169520afc5f651595342b3b0ab5970391f34004c96c969050bc5
z1d367ff70eb5e5dcb2bab8afabf0119bfe6dfdd5c2b64a8c17dadd4b9ad5658995b6011f819529
z29832454a82c4d6d8b6b93b494503266475428cb48806cf6a3dc779e7f9fb95265d761a46b7d39
z41fd84d60ef75de179cc5a24decf52c26faf99399469915c6735662b5d36a792e5dc74b6432bb3
z7a16f45e808ce1fa872e89b88902f49f81bc67964d01f99dc605d1d34a8d4310b0153fd15f0713
zfd72c188eda488cc70d546ac07097de25ad61f5ab440f0fad040193120c819df9478a2c6db247f
z80a298015c707d637c080dd5acbb7b14d93e9d9a3bd8b77b3de599f1ee459a6bd5f1709524e22f
z2859c37be0fb0a7ec35d32e41dc611cc558e34c7d9894d664a95979a651be834c0d2f24c752c91
z83468f799a79105cc6fe41cbbcd58d86666ea38bd2e25e52c74c6dbf1e0b769ecb21f37e3b93bb
z180ff967d740dbcb740b115ee49c6e3fa74f00c6c4d72c2f0a4d63182b6a41e0966420c8b97198
zb4894913b3155e90785dd7ddc032ea9297d02cd5dffde1cec9e80ece59ef981639b2d4c0e4741f
z0858d3009f95aa5fae374ca768905655561de35aabd8306db574de3e68ef4ff7cd24c9adea5140
z951f3b47c4c9e2e406e93cc8d40a1f0102ab877196c5723c611842fd84832efd7008eee32e56b2
ze84d621076d17d88abaf6c74ec70dd1ef277fc0a46b0cf77fc3eb693aae02b089f8b0c9a139445
z44e454e58b68cf557990b8a091f642bafa2a145efc2392a0813e816f9e6200e17ff74f42117453
z6fc0b608ed295162cf40b855a05339f4bed47027eb11aea9735a27688f0b5b682a08203d1e79a7
z1c538439c319f9e6cfe60d38e7a091c013edc23f08d46df9f1953a2f6715615e9a4b5f33476ad6
ze46d5dee9d15bfd7fc245152b4aa70eb4ef90c09972774601d33c4700c6b781a5c0e0477c0a823
zf0f4627644bde36d77f00f34acd6403b0521c205180a8a715fe5c752ee88f2d2c2effb263e91e2
z5ef8aae7e7a1bfcc8c1b02fee1261fc370819c6ee184a738d7d1b291520ead424bf1f534abb643
zbb45c85e9a81f9e7f5518bfd0644df7bcd7bd12fe7f57b476800e96fdf21e64b81b03e92fe5254
z0c5bd9604a375e0fb468d37cdb938845271f2596f26ef9f9b588aaa1406eda03c4707fdd4bc932
z7cb233db694266ae3e916790e7a2ad802f97aea8776b83973c6e27b418ec21658d25ef6908e6e0
z639a88d38f8974cefbe80c7ffe68904660180300adcb4ccc8f5a389eb1151e88e86018c0dcd348
ze6e0d484216113f70e966f80da03b03003aed858cbe922b1aa0c62d58e43c2e419b481f3ebf58e
zad50f7617e168d66073ef1bd9f994f0a85875dc713275be4a4a967dd0625adbeec48243f02c83b
z549c2518d45dc2932882038641b83370f6ee6536248b129f1e04fef5912b218cd12d976e9ef0f2
z443495bdbfe9d202f65eba47b7e0d34d3a53ba3573898ed69971bb3e40f21feb08f6e8393912f2
zc728b8e4a74fd8af6135a3b0d4a9526301512c700b69e092d4a8259364d3c63a110294f1e78fcb
zf074c3d1aeb220432029626cf6752e93e38073a66dce974191d1e50e7dcdbd9b5850d28d2f4e78
zd8dc76dac4e78694b6cc3d90303d773c0c20fafa5f706cc2f2929cdca26d9ea8218880aa4abb11
z66ad8a6cf84e836239f0680bfb26fc65802ad7b809eac9e279fc85fd398987e3ab7b22abba6b11
z6898a3421a5b4222d39928c32c71c002bb86d7afe62b169de2b360ad3945671c1dce3747882edd
z0a8af1038dc0387b62c61c89dabc93f3402f5bce26dcb164f2cc3ed19790a44a17193655888bcc
z7e350724f1fa14ec431f0be88551c355b8a5b973a102aba62d604d12a678c4c422554657b9b02d
zf2cf631041d4c3a50449a8a74fdab41f5c3297e81c020ae7cbe976a3804e3b516af7ae01eef6ee
z89a65c9a67da2828c1b71c75ce927aa77f06cf3b78b6fd61570550b8e4894ce418d522634648ed
zc34b0b0379644be84fafd240cd02a9fe54415a7f390bd13a8c197b11ddf64ccea8fd7cb35585dd
zce75431869f3306720154885c2079f2a1bc0df983ab79dd19b0f07cb0eaf7db8f20756727d7370
ze453e35af493471f77375a7a0212a509133a8d849b88bbc84b3f5748f4aab96f0b21173dcfef5e
zd3115be7b5cdd5d8e54f35fe3cb97d5a9e7349f4a11f634907d96ed23ce0dfb5d2619ececc0762
z56765bf70c3f6bffcbbce3381db203009d9acf4c704f3f5cc22a68288385164cee4ee1f303f43f
z9f2c51bcef6bf3572b78fb37eae26c6f517127a917cfd4389c0ffddd09f63a36737856b416d08b
za796c8ad10e659a8c242d9511ba6f2f1cd02447374e5676d5af361f2b36f06b75e5d2ef3ac39a2
z604904391734e5a092d980f9868bb6b6dde8950f144e4a6efa2c82caddf07bd7dce7b27bbcd746
z6436377b635682a5db0cb15694d3259fc48292f0a1c60646c9e0389dbaa43f3a4d1aaec916ea46
z11b4bb66f52ab124472ffeb941a71e9ce5453ec947ede46573479640e8a46798e598c4b18d8fd3
z08ece01d2eddab150efc12ddd6b385631e770fb72e6eaf1bef7f879fce0eb331f81106515b2f5f
z43e761fea1838043cd43d4ec0220bc1db1e7f0a512c42a7629fb2d8c3cbe2df425f71ea24e4aa2
z1148c2b5d82a021d132f9c22020d5335ae8b96b353f12972f6b6513dcce1d0bc628009755c4322
z7dc8f73a5421f924a2c2f2dd1708272e9e7a0a33ed10016a0517699a7973869c67e3118da2ba7a
zecc892372e8fd688f2bc8c0ae6d857a0d8569236823597b808503ae229173b5f6ad9cd8168c393
zc8cf562ff754caffedc8266402d29f9974007e4f693f5807c4b95edecc28f052411487f9820901
zadb7f4aa52443f941a4ade79c2cb2ed03aa1208b35cf26628f05bb3d2f0056e56ef0baac0d5fe8
zcd37a346e9e05df242d77f850651a0985d4ff248730d12f1b4e4a6907810f87189bece7a6a0c00
zd18e88e441328752f5530684368dde6d3c0802bc057ee4736f4ee7c4933b6f5e89505d13575672
z9f7407d276d56f3d2cfeb20df34940c035494aa39874f99db346591ec4a21a956d5f03c2e42031
z0dc55162021f7c865b29fed07aec3d4aa7c1a4dbf62fda8c648f387c5c4dae3a0564b53e1a4b8e
z1ea85b75b4650c4d570266d75d05498c94b03668dfafbb1f7e5fa28c7081637979bfaf391aa6ba
z7c1283dccdf5383afe15fb14d93abb4f98aa3949669f056787c1d0dbc6ab94ccc36d751dd20bff
z39a3711ca0fa36689c87952bb833a67f80cf950b63e389ef87ddd71ba1a243a4e7cdfa47faa330
z1df7bf7dc60da26bc94262e51c7f4c40fa8c36f7d36208dd6e92711cb5554a4ad5f378e67a5b26
zb33313b5c3afb59a8923cfd0d6dd89f31b3b38ff508011b29ecff576d7b6b16fac307924740770
z92202583084e57073bf5b12a78bc97cb01a301b8f9ae1c0c7c060cb190781a319a85773c41ec56
zd7f547e5006ff1ab0ff1653cee4fa98d25f8c6d63af40806332758ef65e9ea3139d6bb987f3f28
ze77ef55441e69dc76f7b3ec0c410ce1aa7ca0db2310bada9ada47e094f4aeea71b7cf1fc7752ef
z1715d6956cf13c14f3d44ccb252c4467e6f55a39d6638cd38cb6eba16c16115edcc9268f0dfdba
z9ccb396b1a080c2071860c6cc7d7e260901450a6096686404dbc0cc40d5c9e875aa25c6f11a1f3
z9cd07f253b39ff2c00986380c0582d421b5179d9e75bf396a9cad6e433862a1683a8acaac7aa11
z1d7830f1ab16153155b1182d8f905cc9ebcfabfd0841407fe6c47d9f22ba3581d3838d98385efd
z61aadc62365d844fb41af31c312589428dbdbeff975b74fe2b235421702b2674c57604a7eb2968
z311f5557afbb9313d2f20d1105d1a1c7b2c09b00522648a059528c0175ed74cf2519ef285dfce4
z4d7fc400d1cb829321e3c74e86e70e24fb41fcf2c0e227d108465cf299af86b6618e7967fd12a7
zdea2f3dfa90c0175726a618f55f8c523519aa1b6bc07bd3611f988a43c31b02f9f65d8190cd1c6
z9d4e8d5dc8a0cb39deefa6dd258e4590d843f9773db9635a9febe103f50be643120eac44978559
z11c46d76e9dadac57827c6469f99b07cde79cf344c3848b3825b4483b590fbe849cd1e6cd93ba9
z37710c886d645e78bd2a99a2c46cbcc1b94b9f4d28e366948441d2ed268f119b914785e14feaed
z6b52da537206bf3fe5ccaa70d1fc377995fc16df8f7cabb0f470437ff6198a2d1058781f848f82
zec16e1e459d8523fe0f92057b46c2e3f5b4060299f6e47446f7ffea0be687ffdd923d16ed7b8fb
zaa873d2f7ab928687830f839e47cc119fc149854a74e1d99cfb0874846f8e8c100199a0c41d60e
zaf0d2610da987bfc50bece21fa60f33f22a50ba228a8746455c06aa8b14d52b46ed09cfd8b22fe
z6252b797b9cd37849d2c73f10ea3246325ff82c7297162b2fa97aaa6a5e96ef24a5696c416b2a6
z5fe9925cb06e635037ba94259e9373bfc0cd86f0b73a282763e3ca3010530d4e18bced9b4eeeba
zaaaddd84a20e53aa2fc077fd8e12a04be00dd6661fc3abbc1f844057dbacc7cc478521be221ff0
z97b9cc36cdbc0e32d34c209d5180a14edb6e12c8fff4860fcf679fe932a4bae488edde584daa36
zdf256525f913f09095bc2e915c861d88725a8dfb74239b877ad8662a1a4d97beb03ec04a31922e
zdb515c0be0639b59aeb75a2be89fe5999727eccb87af23672a7f55f0a0cb25eab17507b8c73723
z90fac9cc3c54d577b99f57a6321c852c7054a9beea70d042eb80a512bc6e09b6c36455144fea0b
z2f90f4051a00fe6d976e52847b6d500d25903d0f1ffea25e78e1f9226a907cfd1229c731628ca1
z5bf4e83ac96691009ea2adf9592f83465fee86b305784e35c0ec9db395b93ed51c610d8fe75e3a
za53ff090d69f895689651b32b17140200fed1a16c0ccfb50c1c1f93d0c709c8624465f5b8326c2
z91578fac27d0b5e3fcd76e5afdb3da855b1f8d66df264d18696ec8b3c1764f252566cea7de78fb
zfb5b5a5f5203ea8ec787a51008fe63bb4427399d48946639da091600737a4a02eda6ef4ed08717
z3d970d0661ff230ee6740244a7b0cbd1f86cf8f1d37119ab692b3e1f66e4c20b5d81b334248668
z69ae7b81bc06cd9299ba34edf50caebf244d0e290d63d7ed3fbc460b499a01b5e980c8180f9dc7
zaecab53239711e6edbf1863213ddff4b89b2d6f4a626b2b35be0b5a45f06415938dcc79f7aab88
z08419e7b81d2a392d56dc7d39798c7c57fc5436a42e497257c864e11937344d40fd79764a96198
zf2027cc53f3ea72d8f155f4b1e0a410b0b91c63296a1fd98fffa1677424d83616411e5588441eb
zb2027e320382c11691ee398691a3d759ec04120b531153e28f77b7136a4d52559540292a11650f
za187718d952a876c97e19be4f4a903e6a7ffd498b04cec1dadb84aa27cb8b455d7a7cf30b2c3aa
zd4e321887b88288754768eb3488c9e77c3742b92f9eafa7e83a5bfd24a8b8e83cf893341de6b36
z607050c47dbf666c00d64c39d3d15fa2e8020537be5584ef98bc4cb201d0bae9f4d9a0cb83027d
z5c598e1834e0d0d6d3b9a2633e62a559f6a2ca695ca96aaea1c7fd14854de6d9c59a5d6e9e5cbc
z6cb77537fec37c9db20fdcdd1dd792d2f0245bef739eb8216e05b0b493f6b72195fc197cd790e8
zc9af890ed4757e9f060dc9b52dbdd0c126ba2499f2ea43d7865c29ef53e94aacc4d5cbe91cb764
zdf9c084749eec69a2cc84a3f0fbac7957c4b9ea4c1bbb37f5fde8b7bd54884d6e856e5789389cd
zafc7072da9b1de4377fe5c513a790cc6a3355dd5b07f8c0c6bc472af42aadf7da0a948b1ad087b
z12c97754744b96d47ca142a35a3afc62729fdf22b1005b0caf377b54cd11e3590329f8b2a8eca5
z95c1044630bdc9099736bc3731ab4dc5c3edde9dff05d31c948ee84e2b31b7dc00d41232a3de29
z7812d478f4c42beeb6681933c44fded1db1a11bf447fbb0f745e3e40a0763ddfcf398ae751d66b
z9f3718f91cce05f5058544de225961885ff899c675ef9f97f3168ca7d20bf1af1021690dd8ebba
z600d50521372a28597b0091d306092e10636e2aa6c48fc225b0d5f6b07981f9d310f35e5b00767
z051405f15958135548021c076a7dc5c2726f0d2104036ec60aa4082dbd520fd6a7cd146394ff02
z4cb13fa9fe4bd646ccd4d2dbed038689e2e73e40b71b0782a73a8ecbce5d635bb15f9476578bf9
z643762a8aeffd44c0674e3d1126037c6a30b6c63be787a9a0931bcc720da83911e2efe9525a1e4
z29a1ef5f1bc50cdc12f1e879331b051fb37737a3098a4e0e01cc9ee0ef900cccb27aafa229ed0d
z3d195b6df713f571f8f1b188f8be0cb94fde9f23b176c7beec03ae48470e3ea3ce20cf7f926658
z39704141690cdccaa232e07c0db38a2f5e53fdb20b638d997e34a74643e4f2f7d15e34475d85c2
z7901e3a202d62891ffc092942256c91be446f45f315ddbf0045f3e81ebd939ddaa86dfed573eb7
zb515eee28305f7ee7f4b3d1c9ec9e49e3eb70568c24a6bceec2034b29b69fa536595dbf179eb92
zb1dfa784124ee672144c7375b06d29139ef619f7cd777fcd722588f288a81fbcddb1033961d1ee
z2d87a89e84aa677eea24fb4c1cb13f8f6783c842bf0b8e930c052aa9827b2f1f47103b2452ad62
z31f790a89ee55f947f0cd1274986399e7f840c509ac41b1e520d15f916d04aca9e682176378559
z7907a92546c0db3076b0a9b502b0742c57194985ead258dde005de5e5cb3a0a383bbe180bc5edf
zad29dec951b3da350e836c2668af4c7c9a007286803caf31e185bbe50334ea7bd1640ad71c947a
z65cc2c15de9a50985cb839611584913a1bd2b12e92acab1614c329057aab91f32b1844b3488b96
z70cbf04d0bfd77caac99633542320e887858ece75017ab39666fd6355aa31da59c51e7556ccee2
z5eddd2ff899d9c7fa0471b4a2532d0c6d86f15544424c2682e2281d6ff9a0bb94195f7b8a8aeb4
zadb782a54b6e01d64c7ecbe59f31ff9e24d249989b2d4beb73880f02d6f49c88e5220dc5cf0527
z8731a3ad0d85fdbcbc7d76322c3c55a9a05ff477db53e72dde4626af7016410369b5b8ea6c3f04
z87b7baf849cccacdd26945be71f86a330f9f2f819eb802cf0d3b98884ef323863715d658228845
z5724da082c56f27fecc71715726c411ccf03c5f2985254df5cf8bb80fdc188ebd4ac4c91e0a0fb
zb3e3300a625777f34b1fcfd0993263d5700579873e7cac2d7ec1c470363604df9d5c041d3b0bdb
z81135a1087877df6e627d9844cffc63b558582e035e8981e8f7cd54352c0136eeb79cdba25725a
z523535895073374859773d60287196d64198ea80a47d031680b96927462d7a6b6ec36512e6909e
zba210aad3ba97d39dd61e0adefa3238098730381be242e45d690ce59f1ebe885edab0bc9cb3691
zb206648b2f32243d0b1740afcd98a41c2c1ef604ed4fd1949207bd91d461cb0e6d6b2a715646a6
z7e22adab6d6009547794a188bcf1be69787358ffc250f1fdf0958bb8892c88c9c4611caf5a1566
z9b8b3628f734ff1b0e377750454b6c8e350953e1b47d7b345b8e4ccdaf5b8f9cad416b33bb5799
zb0593826dfb8efed97261acd10853df35f76fd773747a96760bc89e550daf72cbf951810b35f46
zbb56682e4ef99ca77c2646c0670f8a941b0ba8fad8517fc3d1c7a0a75c8339f6220d6c15604301
z3802174b3b5cc9a3c47a3aa0bc41d6a56467beae8dbb7a7ced316b4cf270dc4d4267ec400c361c
z1f5255bb8c8159eda200e4b4e94f72e6a1c413e8ac4a0e65fea2d93c89f60336a2975d36d475a4
zb8362c8afb42dfeb7bee7836fd2365e0b33a871f871cf25539e961c6bcf2e7d30a2096b8533028
z096b147a0b49f861dafd001a5eedc0135c859e1ab5db809fb31fb0cf7c47e3e09c375986988f01
zbe33f4ff88ca18762466365f7e27fc81e764e64fab691d2a9362a81a55ed382e95edf217fe676f
z3addb2f1b3b2057e2404baa822d975fcd20c98669ee57b8825cf065e6356dbe21e238084f08662
z28b0b9ba4a85d88f8f3e3030d7b34d44422e7fa493997e9250b67e2e5cd5eaff675f0ec72c7628
z257be4121625caf90143addf19c13a9ca031b4e593a68779d38b17ec6a194a3df1c16d46c9c654
z50dd3f996d3986767223e382db748b70d54b75f7c3baabcbe268676dfe8f9c1b9c93589ac1fbcb
zedc61fe42efa7253594b343383516686b0c0f37905babf4ca83db25d7a53be5c1764cc37efce7a
z028f78fcbcc81df62f91f17cc3ae1e2313f14160154152086c568f4f5fbd9bc14354114967e2a8
z306e2151270858acd9c7958a7ad834f337d4a76a7fecb3d82bdb9f282b95fcd0d028748880c590
z4fa16baccbc17b6619a465ad824cf0043677a96a859a58556bfe356c1e3753f5149a236bceabd9
ze70c214963346240421d0beb1f4a5e7630a699020f9e3dff1bb4c076cd39baf919d40d6f1d42b3
ze6486c996001560d9e2a6138ddaef38dd9ca959208c7a4992f52a6dd56f80e52cf4486977c2a04
zbb0fc47b2cdbe07b5509200626cd206972a48d7ada4de141787b35cc5d118e5b278ec8757206c1
z541efd6765b662b809495c81f06b5fe947df0b42c52b0de2b8f5770cac3d8c7e6013eca2a25360
ze742990b3edfe69c316118a18c528d223c88f0811b8dea9c976e77f385f97e5e88ca603dca184e
z9bf7e131e92eed076280a0f1b3f0629353be10a30c1d3f14f8c2398e85ce77aca3b0b5f78416bf
z9456890c5d0fc0282d1e4ea09d17208cc8feefc78c7f42afebccad03c2fcfffc79f2caf8da8c92
z7f782defa093bb6dfc2bc8b50925dc3be824fd23bdaaf8be12ffcf9c7a040890ef64fe268bd68f
z1ab5b536ca3514a53eb022fa8aeed7900a59c3a1e2b721f3ecb605ec01705d64ff9bce7466deb5
zfb7ec1d9613bff5e67e54ab660c98d06353eb62539422c25737c16f7bc569ef71203c3bb48a172
z941512a804238b5dd3ac2fd2d0904be2cc8ddae0f826a41d6de952cf46492c4b2c15c4296c1181
z93f874c1d4c6ac621a8e45fd2aebab1ff7449c8f73da2533cd17bc08ce67c560815eaccd167a4b
zed2235171495243e465525d67f041c1138f606b565c15961bf1427fab8f7cabb15750c27e13ac1
ze5e57c17922ec85786c2d5a7dce8736e08a88f0aff8802eaecf8d335c72b66619f8d4a7fc7cf6c
z13bbdc6eba23266f5b6eb919d8ad9469530aa8b9616bf21826d711d650e6063c2ffd77fd155900
z076ac412d96e79f570820f94ecf995bbfd948d0d98acf4e67aa98f159fc64f4e0f42f2723e1a68
z1e8594ac4fda310305de3a7625e87da51e03d933622afa4072be97a5f8fdbb3ee0277bbac1e83f
ze1e8e6babb5c2b87750a765459408260b992d861ccd4c16167ddee7ce7b0dd57f23e03bdc4b1eb
za4cf3790af2b697a24bbc90823b4d4858e61a346dac39bf738a9d0c58266306dcd2001f0536d75
zc2380ef9e8168ec57bc0668711e8ef91203959f44de3a5a8909505d6d09a4307f2fea0a4e24f5e
z460fa1d52230722ef46c03962879dd8c49251d6e8523b04925895d3563d272db6be3d390374488
z86974c308555cb1ce9af15f17857abb62e5746d60d47b3ddd9f425539a7ddfa28c54962976b986
z677e6728221dd635f04f6a10a1b89a5671050396514db6a68b635b97d134c298d7664b39369014
z21066f29f4e3581c13de7fb405a07c65b386b84309ba688d9ed8c251b8c254bba65546a6ce8bd0
z2d5b25016585d5f7aa90e0cf604407a5b4bf83f234be0f235677fe31cd825b6083b6000d697c9f
z39d8d1e68417ecba825c8efc46d1d782fbaf508aad39ae113658ad4c42b744c98844a6564719f2
z8be82186939d24ca86ad66cf8cdacaa7124105615f55f4128c532affa0cd7f37d064030fc84a4c
za48235db656ffc54f9df30cb123436bbcf98640358752427cc1ddbeb14c99dd23d73ae008f3d7e
z5b56f2d2c6a14b80231d7c33b9b24150ba50d624d06bf273b7ac370e872f408fb44b0acff07922
z83435a1c24beb2815457050f01191eca1cd35d1d561ec1626322e4156784a26106ebd811e0ab98
z59311eab0fe92d059eeed6e7d35cbed6f2f80e47dc8a3ec5d04d0d3571b70493d66c85ec5e5991
zf93582905eeca49232f64d98e91f0aea5c9aa7ac2d3908207d8c53a6f4de6af0aac134faddc1cb
z579ae12df9090def15e8f2eac2940c2b2ac0cb40e219cbe620e0883a5ab11c3f2047af1cf91125
zbef1a9c4bdc5398fd3e72385e08f1113c7ac6b1064539cb545d38ff9668459b21caf47a2cbc71d
ze91461c08130753d9127e3140d8a26eb73888b2b0e80b12f35d716f6b7383e4a790464fe514c98
zf3a17112dacfe9e731014973abc1bb435bac2a77f9555547d78084011087dd0feaa8cf8b0184c7
z408d9d2cc9561933d873aea7a24eceb76ae08b0f396aba5dff02bd9cde914a16bc91bee3382f60
ze9cc89ca61a7c123a721800a4050ba2cffdacf4a335a0f801533c8db345bb808dc46b559549c7a
z3859ed32478e3a54429f5d4fdbd1c795202ec6abddbe2575e24c1dc9a107af8c123c19874ba4c4
z0194c505b115acd2046184db44609f99820a3c269a5c8c9bd5b65b94c9a2c801613005e7a60de5
z04c274af0092e123a383621bbcdf046781ed90e3b1bb41004ba2dca8690fd6fbd1899b10bac94b
z7df44b6825eaa28d0e1358f8cea6e6d75438fc550597fc59313b92871fdeeb7386a00aa086889a
z1ee650a8694341d3c6a882dabdaa5004470147ca50779896c183812c7846d813efb12f6bf03286
zbda9b889b5e95e7dbf07d5e973c9f600109171fe3ce00d8a4378fa3353c8842bc4993004929420
z4f890103c3bfcb508257b316fb96f3d6c5ecaa2455ee1ec049c9fade20049e6b3fb94aa1cfe9df
zd5ad9009c0ef3434c37d2e59755f6752658f2bed43febb33d8c7ce1d2dee4ba0484bada2fe446d
z67c8156cc5ddbc1a5eef84c3329f64113741e46e8d86d6d2210d67b3120eed375313cdbda14860
z19c517282ab7ca4055225075bb5d0331da935daaaca11c9f835beaf2c327850ebfdd5a4eebc9fe
z33ecb598b5bacf569c1d25a033fbee70aa703e065a26d37eec86defa3d233a1cb3c7542ef53007
zca2377bd98965a662aa561b283af433828060226e3670e3b44116a77cce27c524c91698a277665
z9f66a093bd230a635eab2548b1e7d62f53aeb1f3e38f519f2fd7caafcdf36ad936a84ce9f534f8
z3a8971606a169e2db836c322694de0d98504329ce669b9eb477d7afc219d14f9a5a32394cf105f
zf705b65758cdc283a087898e4314236858dee27a3fdef59a55916578cbc1bfa1defff3ddb9235e
z4bf82ea86b95511b1303c98060f2191e3be2c790feaeaa52677f228b4c47eeec43b51acde0fe6e
za42fa5e7f1566eb7da16db9850a60e09a58a86a93647fe4a65843e1356779821ebe13fdd4c7f50
z51a2e055523faad5c5e895ce0a0486b9a42ed0d997465c0502096c88156933be4a0482eaa17d5f
z25a6481dc41572d397068aaba9733ac841b941f677fa0d25b84aa334730994eb3f0d0bc848fc69
z71b952701499f658a469299d06c1a15ff0fe8ea7c48e3041972ed538f4d25246ef219687aaa9d2
z660cd2d4b4625c0fd498c3753d23d01d66500cb6c4e6d0144c6ba6d03dfa6532223e172022eb7b
zf6868f573a576abad0c84b48e672efcdc838e9f015d9a92f4f465ab374be4d737267124f27d759
zb40e75976ebe8fcb63bd1854020fe0de7866fc0aa2219f0fc00888a22e0140ff8921d6031a9a6b
z00816d4a468058958e20e5da24834304c147f0d0550eb9819449ae1674d1318b924877341817f5
z6af0f10ab7c737300d7cf16af37256d72d26eec0eb0bb281ab807a2b2ebe5344264bfee2185d79
zaba66bc0e031bef985a855b6b2613037fe5f7082e3488e59a524147803ce5ac570f77386dc6d53
z02369e902c80deeed91d02537aad159fbb0e0e214f40d7bd23a1bd03a1ebbfec3a8470150ef8b7
z0192d5395ed0ef8d8e8a809c6b4becc16edd406c1ce999a96cfced1c302bae2a51ae76cda90bb3
z557285d8764c0c04a7a55a48fdcb4c5cb0c04ad4f6454f1847b927fc44011a73b0aab3b90baeaf
za176898e5c00f4a5979e4957ea2a46f28fd475ecb07ae7194cd9949e72ba1570f9a956bc718581
ze4d015f58d0e576edb1c77b152ce33ecbcff125079a590af51736b91a8b02b18d61fc759bd6472
zbcb1a09a4fc7084becf77f8dae542ab0accb8b13eaf46d054c5a12554222ab6c951790d85bb853
z024cdd94e7a7458f75233bdfa21046fb2c43fc2c97e74f8c1b80fad6b3135caa6220c9f336ccba
zeb5ecae8c6557aa53573df80213176b359ae050dcbcccf17f22122194b1b4759b3a85658b01742
zaa4c7dc76623d0300449272295681495a4e669d1e77c8ed2d697164946dcb686e472622c02f6dc
z51415271176b0e239be4532f1de3b2bc937c3fcf11e91cfa9a36d50d5749c3cc1b208ca5d5e310
z09dbe890a20978aa52afa769a1dc7c263ffa3b5574df34ae9a580cbad58f474e4444f569612713
za16bda690bf325e906e8bc493e016589ccaf3123f3b74e044678cdf8ace12f45d59c2f03e600de
z2900c41699943400f56d37bf543d95e97436793b652a698fe91df4451d96b2237c97d21c39d268
zd2825ae4db18be9fbc99f2ebe9aa9c7143bf9663692a8b7f2247c8081257c8ece927fd7e1fb6b5
zcdd3ed13f8fc38e891454d8655a573f89c3b4afe968e70f7a2ce249fd1f7defc415be135d0a4b9
z6c64cc0b0bcfb0a65dbec6462140f1dcaccc1befb28d8a256a3d599a604c8f084180401c2dd93c
z49cc77e1da89d26849e9050c2e81e67943e0cf49d449009fd3433fc4560987af0f8a6708eb1230
z518a48c5ba59bed93a394d3b58c66b2f8525a3cc1416c77973abe09011c18f1f0b5f4c7441bdfa
ze66a7dacbee53fb6ec87206a8e9dfd204ae2c88f1f07d89624215e986ace48456f918ecbdff5f4
zc5ea224536fd51af58733e7c75828776a04e789d32a545adc02e0ffb6c54a3436155c543b29975
zd15ec9d3c6b6351b39dcc7627dff3337c30515f846bb26fa0d8a18699115b1b043c77c643f7317
z142de9250067e95fc3f69513787cb751363b5abcfc04a35570cd851b8fec3ae4ed9ce5b5f90d09
ze5740226afb927a7f6ca9a6feef8c9ba75720dcea5b4a6b3c44f12faff2a7534f2616525f9665b
zb235d37cb794effc2bb147c128bc005f14ba756338c4dfcbb288673d075cdf29ae870e740eb0de
zec08d8d0c825242d5bdd508e163cf2de5615d9cf8f2b450e8b4401c0d2ed4992bcbadca7170285
z7c57c8927aa7f090a4a6ed101cfeb121753646d8a271429fe672c5308dc787829c7001f379756b
z7d030fae191602f8c8a1f721f429729ed12fbdc38e36715ae2899dad5ea06e0f8a6f40f058158d
z1bf43c3c68b1f2978f037d53873d85ac00235e318ff242ca531123112105c6ffd0f20bf5a0cec0
zc46cf5cadda0f8841eb1be808d7bed2b960a57c4e33fe664285123c0322d0a8b96bfd556a8c574
z4e492508f06f98dcff60cd67dc43c3ab433ad0dd862f7d86efc6cad16c6231d1e51c0b343603a2
z75acd0487fb2decd89472b5177fcb48e0d192998d9113799b0d25fa8580d5a84c1511504337f52
z8473c7519baa712bdfd8b1b86d55a621b5536267bfc2526eaacd286137a0f984b629bd52a631b8
z7dc9a17041b59117476ba9ccd46bef92bcca9b91f23120a4aa0c81c2d0695c2e20c0bfa4fa6815
z67adc82dbbbb97a8070dc13c060c4edbe05c15243e9fc4744be6b3b27cf7bfedd6605a67bee170
z8abd2c170a543f81a1df2f3a6ffac18c9e3ba65065dc0d51b7c33e5a5999fac685dea82eee947e
za45c749dd28e6c24d1bed51926abcf35eb03d4d402c2a4ffeb041fb7d4c7aca6c901bc95ff0298
zf6f76f2ec7386ee4c54a498887655d52afc4e2112876c08044b20f37a3c7640c42bd0404d12405
zb658081bcf998322cca515e5a669d23d2ed26f35153e0342a00c220c7eb0d4b40c349d3d558fe9
zbd39cd93a9465a87f129f414b7a7849fae45c27790423a902071c2f4eb0b399dd1b41805cedf2d
zc6c293a6c60440349c274c3f4a5a0068baede0fa98e7478c1869b470265a18e51703cec7734982
z7d883aa7a4c30f8c27739a2588b2def4d4de2f16ac485f6c0d8ad9e7340324dd05e9bfa1eb07e3
z711f197823da2fcb4e01dda89455f7c60cc02ea2b31d369b36f058f5e8e485c5b4e08df4cf6eb0
z0fd9b319af0692ef33591ebc92456c5e9bd09f01ca844ba8eb7ddda3a1aed4b0c8d735839417a9
z1018ca38f2b488fd88187cf39d9ff829c9304c848cbc618dfc2e7888ad126b87585ecabd1b4702
z84de69684e5e16d71b8049af697b5cfe89338b950f240a512759b30b83adfe4b56fc6496f5faa5
z0015790755d1c9af252b00c88d206fb078cf64d824f9afbbf2a41971e1b275023827586b229b2e
z0c401a7274a0bcdc3d18a3a1522becd3caa67cba617cdb097eaad3f64c51a5b6da8f983f0fed78
zc90d50c06223abc5aed9a0b10926078e1c0671d0e12af28b1569899040a6a162d598adb923a923
z7ec78b66db0a082c84084be7bac0da78876b12124695f28ed930665f8c609d85bb239639046972
z2c4faa255b6d9e5531d40f3cf1e41aecba1754f3bdc08222dad71259be8a7265d01c8372ca863e
z3547bb10b337f91628dcdf37ebdd60fe31daf7cd7cc6a23d5e7399081d3046c695d9e11ee7f2ff
z449e17bd9cff0daae5b7d4b815b36e05d07f423dd6cde5075974937b0c5d732aa9e468820d9660
z49d8d1bd130899fd19136dd8130377ed3ad2bb8c49afdd0eff574ef6a86a2e2ba8c47cff4dd849
z9dd875bfab77d77a5b3980c85b35c1c5eee6e979e09af4b7511571def5974743725a7540d2ae36
za4f70de47644910ecf931ea992ac36b305f88af4fec88164282315b8af4b42b00c433d531ec00c
z2adeef168b7acb6da1df9f7552d5c34fb66264cd013bbfe3acfd8b090b6068865224c79e2241b9
zf58cf75e6bec2bca8aedb3f969a41ca224db484fd8c2eb6e86508109eec7105279a2d828789e64
z0f269ead1f38dadbbda1c4421f96364ce2b91abddf77a197cfc1ece8631d899a28a1f4519787fa
z067cfa4b55bab56a5aad6b49434e4a27941352a396a80ccf6b7a7ea411d862f5b6f91b6f67368e
z869d1e036f535ff016ea3d533da0b22bea111e5037a61ae1f490011ecc994e414ce19b07513f0e
z04aac4d8591be50d94edda9bc0de07aeae1db3059d07cc3784decec50e4e36f9fec9d83e22cebf
za6c99a2a156fb473ba49cb4a40c4ade76bdb8882734d8a9c2f99d5cbe1f5699b2075114b5f1c0a
zc23c2746c6ef2366f23e76c6ea2149732e57507e9c776da8996a2dce1ef42ccde9183f4c1836cf
zf9226041dc720229bc263b5e5947c16f89110846561f0ed664a9c5f7a560f9edb55d40d8116516
zae44d7d412fd2785dc63ac2218818c805715458aee7b5411b1663c4ce43b36ddc58d2b2fbfad8e
z9eb1904d18adcc3c199eb10d7b265c38bbc81a3c89e5f1f7bba9dd04138a49cb74b75591475a6b
z428e08ae4847c2e707a6e15282d039cb05818c71305da873f23efe7499c82ed973f56496641ba5
z3d3c3d1a954c02858380ad8966092dfe06c117fd8c5679b8d5f1f9d5e9b4b09c28dc8f41225892
ze7b98d774b6dcbff9a1003f12a645ff6c99373fe71275a272610fccfe5948ac544b0e084ef4ce0
zf04ed8bcd5b04374443c2293ed2ab94a8f7aca146cd42da0ef6e041e55667c22396f8101fe1f4e
z4d11fc457e7692adae533be4cd88f191e12a609a466e617732da96f2b4e1c75a715329e2b48cae
z356c834d8ed03933f0c6572ba10c041dedbafa82ff9c368f93d19e18077d94db3bd8377372ab6d
z954c980ff3b6b99b581d73979de7f06c32e4a1379f7858ec41d969affbdcf471a9ea2021ec3ddd
z0a6206c29fe7ff40b64ee03602b25de4e3cc611929fccb99aa211960f9665a8d733d3f54e8f429
zeae1d35381c35a4929ea2c28c4263b12fef6535bd51b284f0a53829d621915a24c618dc9917734
z5d66d3d7cd97bb97a7c425bec786c058aad7668fc0bdebcde5ca1ad239d5e91c171014d9f142b9
z076679c254abf337c37d977bbdaff320cf2d35d22dab88ab999d241718c4c70fbaade28952ab53
zdebbd3632c09c9df0930c2707c65c58f5cf3eeaaf0cadbd90311aae528358b7c19641687ccd2ab
z05684799856745ecb6efc170e15da6ca746e30e409fba8152497c1d5a6fe98851670aa364daab2
z3020096004433b39cbd59e106a1fd92039b34ab3e797568bfb47ccc30c1b0b21dc798a975cddb2
zda5d4576d52615127d64aa57aff6a3fc18ec99094ce0cdfeef8b3750428065bd3e57f6c6d44b39
z451fb016788168fd97fb244747af5b1a8fefc784192b1a9292f93ebd3a9883420c209c9ef18af7
z8bda872b98d51366f5502698504f88e8e73004e784f37b64ca106d7f82aeaaa45d69522e80916d
z7193a5446b9a3a13aeae55214f31b25773d020d5642eb03ea42db838d9ab27dc9a5ae4e0fe1d84
ze144a7f8dfe88b54e3e0b009d650cbb323285936ccbacf5cb172cd387d12243c95023a88021937
z665eb37b6257487cd0a6357817adf1275d2fa8e2a8c12bf7b1430e9d8246ca3c49821507f52016
zad5e1f4c4ccc5f69fd6eacd77ba1e750a7ec3e2a274a99d9dabac7c81f1fbfaafeaaaf71a43903
z570c4ccfaecb5b0aa56fba7aa7236175b1a8aa74a4bab79b8dd2c2e2404bae7727c791b4658e24
z955733a3e30d50c31c5de5ff61e80d2b649a820149fea96b79256fc15c26f83cd32f9d4c04df60
z45ffae10c1ae6887c5960af4b1c0fe3559af644554d1e66521ecbc4cf519fb5f5160681569c46d
z818b683221998a4fc9bd6f27df568f007cd8260805f7977220f51004b16b121bb4a71ed2881d24
zf269a96b500a7e6513dd219d64ff68ce63fb90117db4e5d58ddd21c65fbb167c9062b2d7f5efd1
z34bb390807db1eda8bee077d2af8bba887aeb704486e2663ccb672a8c75d3a0e2ec87d781fa3dd
za13293cdebdeeebdc39affbe5822d7f85d5e6857cacb34737f6bdad68db2e9f37829f7e2c3396d
zcd088e02bbac14dd00b157ee601bd93cf550967192574dad7ea85b5d761d84699837c577eff3f4
z191a306ed880b79e5644f449e0efb141fa7bd283744f01220fb501728659155cb88ce8711be539
zef97ee09dc9e14b72e502a1c38c680dd81f02d5a4eeea6a618897af1fb7ef5541898cbdb8c5154
zf393a84b73b625b7561ee68f386f4478cd181e503f05412ae763bc5d639d2d6894391e765e949d
z6fde4ec933c006df58800c7e69e0f2354fb8e8068f6a41d0db3ba5027aac26d4ddd805eaccf94e
zc0fc173e80f644c579a94d6c33f0a706b05b4dd1c7ea052d4e05729c24b684b6eeb02591d891b9
z8db84cb7c708f8e0a56e8096a6f00d522a3f89e862f0c055ddb26b94466c9848fbd08b4b7cbf73
zf07f78a1a69b48bab32eeb23ff951edf7b87b3dd48873b9cd072e933c2bfc365566204ad1e970e
za5c30fb3cf71822f9690881504d166325d57d5a8cdcbd9f40ba86b883ecf1302ae58bcf610e75b
z61a3ab891ef52871f3b8803f9f18764cbcc2662e8a08a5c48ef7102b7224f8409d8f481851b072
z0bc7ed58175a8ce601e73889cbc3950b22ad79c347786110d5afb1c3a390f03b52408cddc6cf4a
zf1daac5c25429c9fea5a037198327628da1dc2af5bf6ec1a1b50f322f814038eb551ab8e0a5ef9
z0f4d6e13b81712265b350bde7a2e19d0ed3c8ae6b0d0be08ff99bcf53ad57e0636feca8f017348
zaffde549a588777b1de6a20923101d00707e99daa83f49b0be0903e47385508691ce1a0017a13a
zcd74154f00264d1d9f8d3f76d33b42fc1400081eda774694dae63b961db6749258d8ab43e1b456
zd8d19ca1f7efa7e0349978fe5c124af93ea4547aaeefed874d3126f80eeec25e3b9209cfbe4dea
z466a566be896cbe6667f8cb3e0cca28b451c1f0f8d0aee6eb48caf53c0735fde3dd48f4b8da689
z94855c123d5b9fe8fbba944593bf3d770ea5894d37c3e21093c8f588734512f890af6b5c25d721
z59b5c96fec5687afa4710080d69f370049cc0ad71d2811f115818edb14d454b9c32704abc7839c
zb897bad6a7243759f580312d74ab2015bd964d1b3f3960a22cdcccedb54a72ff8a21d34b0f2626
z835defe1efbdccc274feb418aaa7ddc06c991bac9ed458a3a3ce38f6db62be71bc9574a65632a2
z925516dc7b060ea847e49829903a284dc20436994cfa359118c4fad4685e23bd2dbd37ce03e6fc
z53187cfde2188df58ebce2c4986c5db957c2e52610bf5fba82045f259a90f797a8351d7156b913
z2f1d8eca57d15d44c68ba2eb203377b28dcda888c9ef114bcbf38d045601cf1b8ed7a9996f97a7
z7cb79832ba1124b4e046b61eaf81d82f6730edfc461a470d222976b03acb6cc16e5e134115b4b1
zd8b7a6183ff6f3936f9af1ddee2393d86404d7644b5fbc04bd64e981293e010d54a31ad7f722be
z0918df8f148ed8a1d5c06e2c193d35e242582db9c82b28e22d44fae77b6a09de787a1e99889771
z10944363313ebb7be520b5072a6c08b9a815e3a556d5881351183863c47de1297018134ffd7847
z756cce3eb115793b6317b4d13f659fdc0b5d073c103cc8ffd3fa3c574f56b9045dfff1a014d001
z80f726c214c05830bc9f643c16c7819abccab885c088343ffe45b7d7f819e3647ac8dcdd995715
zcfad6075319288b7d973da6ffc920d62b1e832e7b6b8766c1558bd6c8de38f46389e569c9c424f
zf3deef1de0a18ae2d5048e240fb9e79ac43a704c923e521c8f633fe54977ef347c928591f098d6
zd4feea3dc40ed93b048f8ddac58b4a50c836642a5d379607c7f93a130705496abe3b92a5b94746
z8ca26c84e58a0237797f4d749f28ed3dbb0264408d3e47578c01a3748f7497b526395acb868e6a
zb4217dda34b51362cab59106d5061ee12b88de0c09a2f92f006e9d135c999658df075055179d5c
z12644974254fdc555dfef7f480e0adb9ad313a8b2c5036a9abcc1777eb587f591c0db32733c10b
z21204bbb83313b399b02aa0cc71c6d4e497629368bd446d596145600af7e221a391576fbd1666a
z089dec663981c953175d2c29b5c2a316bebf41ea7e1178166869362787e1028982fb8f4917532f
zd6c0d495305c5820a27aa89a9cd8b579d80005fa355f77fcf5228d06ffb98fdf3e5a6e8da4cc9c
z5c4670ace881ecc840e5d4ec7844db00342557a6826b61cb00e2b13077686e534b99ae5b5f1af0
za51d07fc9a5be2664baaf6cbced13b4439f77d1322e9b9293e0c201f8063fcd65fd50484adfe2d
zef5c32f003cafd99ab7af6ec7eb177efe2d0c999efe2afc2fc170a917a4f1c1c8ff0120ac460c8
z0d47993be6497bacaddd264b0594e982536256ab79c2d1a21b8e4397766d3b106bc46d69c3038d
z50c4ca093f7e44d16e1310ab644cdcdd99ffa3877e6bf9e89cea28783735da57a2d1da817b5612
z5b835db909ae1be6f293767ac5c74f5ee982609a572ad29ec82610cb5fef86c0e7715371a80edd
z22aa4b369ba57762b8e3cb7b0883d16ad425bc229c836f736a5e9e4aaa6e3880d07b4b87fb6ee5
z8e7787f626997be8079cdcde1e7dc755037077e5e348bf5f0c16a973d1b34f9941b782e38be96f
z2ce1a5e255c88352469abe4c392c00c2cf463eaac998e4d52ce2e86dd3807d712f85d1a66e18e1
zc394deca90d1c5272e1aa73a61db1db056e6bd2b7f01c751b1f3966cc4e5c66a17c4db79291111
zb7c6e6811b88e890c34de1ab390c0cb0074c96b850e2d8030ef9ba6446cf81602e6f5ac6eaa03c
z4547986d59e57048712e4fa1a94c1aac870b2cd2eea9eac823d01590ac5b0f27a8c49412892f50
z16cea6c5a0308b86140e1896133cc3fe7588cb35e0706fc24e3f1e4fc7111b5436e87db63112df
z5b8c1c553ff7bac10bfd33850676d9d9d02dc1750f3482f4b58146ad1681d70fde629440847f26
z50d0364cc1fe93fc61800ba163543c1086722f198b863b86fffc6abe5b09eb1878fa5189513777
z29ca6f0d9f8f8c56dcb622942afba804e2c75ce898e3cfc0f62aefced20d4ce608d1fd4abe5e03
za7b6bf7e5055594cf523661665163cb0cdb1809f4a796b469d03e0720abde8600643112bee8f89
z384c458522e34ea2d23572dd86eac82220b69835da24f9e1738c3d16ac19a7754b75335d81988c
ze98f6e1da131dfdfa65619dc0994edbbcf51176fd533d45da45b44e37f8995d9327c490f112aa4
zcca20b1562b1ba24e9d8c9d1b4d33094dc99b38677f170f9f781a296a402c0180fc2b127012a0b
z3611d715bb8e42943ee3b716bd0e6a56fa722765e6369c6763ff7c5e030a3d550aae02ee2dbd8d
z1fa99862644a3358e59c44511f4bb771617b4fc252b377a4f09c806147ec643de8479d191ce953
z2f9a9a07f9d2d6f5e2bd03de096d17a830e6eb02ff3b4b44606b7af956b4b07da7f1a4e47f8aa4
z021cf75b890956ed1e265b8d0e288fc4639d6f37fac77842e92dae2a2fc8dc2c0d4e99516b7e39
z631ffde9c03182cf04b43959fa7d0cf1c4014a5b1c6a2e06a975de254c9cab7474352557862719
zc4e2e0fc5cce141955980678cf31530d55f3b65b1d8c9983b9e8e41952851c9ff52e85f0379838
z4967fcb5d83820abc0cbe038414143282516794da37757821d7d9c9a1e7ad828554f4d29666a63
z4c460d3e87081f24b6129ce678f870362f0450f838419afe5307b821660b0eb232e7009a755ecd
z8f491c23e8f74bcb1191d391d79173536caf102bcbf09743903c6ae47a51beb2304f480bcda6a4
z02222c1d2b678a451bf0622788ebb44a07bec0ee72a54a5ce075cea31b8b2bbaad94dd6904286a
ze2d3f07b49760e5a96509741608a262c41f38a9bb9b4a7348a0d7719633dc116bd937157faebfe
z50b38d349274226899f133a53661593317c7107dfda9589976fe5e73d58262095a94aa183d5a57
z61ab3602b82539355ac63212a445a74b7b4eb82ff1c001ea162f7076144ad122bb368895b74d15
zbd1a5799e87a3303a8ce313ee92c28dcf10a6054e9f1b66a069c40234c0ee2d726296452d44030
z74e9f730a6dc8a2f6357810442146c5bbbda7c0d80a9316f6f80c5a6934f034a209e3f4ef9d807
z56a1b09f95cc80a00458b27628975e353c208954b6102eb2cbaf77c9e8535c63a508736cbbff3f
zc2ce5b674a4716eb497b1d721aaafa088f6ad9e76e146e7d37f77fe087ee8f587b16aacb21b642
zee03bb4d9c1a2e4286a032bc8505a90ec181a0cfa49c98b51460cf744c3140ce623d162b726cb8
z32abc88e12c8c311f5aba5f267bc509a17b16c55896bca00dfab938a20da4b70c1003fb94eb692
z4584407254ebb3998fd9b4565a271410f02908af3dcc2757b3c636e9195cd87185d85a801152a8
z316ef67d98324f21ab5840c4e12c3ff6715a1af15458857d0b65e928e28f71b90e138919b2cc43
z2ee1124a85d7b1824565f2fa8d62eb35add39a6955a768a79281d36ebb0171d1b223ed9e539ebc
z6a2965c7c87c5256ba5208a252965bb08b43bfd038d86c2aeffecbb26b8af85bc911495eaf4b6e
ze58d8c5317a9fd5aef9807cd2611041fd5d9f231b65c301c9e1e5736ea49101f09fb49315e60cb
za5c47ab5dba7e3b2ce9e017de1259d17b90c779c77b24b288f257e348e558f5225a1c1c550eb0b
z09542619f83f85b7baa50d0b9a2d7a92c75a9a5cc535ebf46158466c3457a12bb88e33701375b9
z0e2c34eb46e3dbe92ff267326bb87db44bbbece06abd5c6270236d6a8608d594009549e50b73b6
z668cb00234ea0b96d8d60393331a2c8be9fd83f5be6c4b94431058fea93deb5b0ebff6bc0e316b
zbc33ea1cf1f38f59c0549a62f4db937e218a04093900b4aaef0167510ee488e15d39ffe3add13d
zbc4a2d13746ed1928660501dfd98ef96673cdd084097738740c9835dddf29d213f0520b450bc5f
zea50c76ce7e9c0aaa53cd9aef62e76c8c52eb83842148ee21ab8956fb9c1c9470829b9023d6ece
zf151a63e65b6bf55cb5ac7e6a395844960b44d57a3f4d8d8f87f637cb1d03e758f472f8eb6e300
z72730eb04cb053bd68e07388bc016083a83673d4b09734be4d2794e93a3ec268a6e8eea4d2a3d9
zba74051271d7f077851ad186cacf6bbf2a7a785326f560e7682262862e4a1389af52ab1559e5f0
z5f9a686f74019ea6923d426c052301a3d23a10d2f20615000a1e24b526a4416be2f2479833f4d8
ze47e8ab9596da0ebd8088d2b1b02e441df253d58fd4ae78a3e792b9b608b9f0c28f9cd9140da4a
z236210dff3bab9cca6deb2cec6b3144fb981c12b1de1b2c31f7522d2861a6b90605170425c9332
z5007255567534e7b049dedc1675cc0989600dfc6ac3befe52c58311fa1e97de2c22608772cb6c9
z8cd1b9120faf22f49014d82d1911d9d39ea698fcb9e17d8d820c4dec5e844c76c666791bb717f2
z5e2d86158a9503bbc0bf57ba88f35cca88a0958caaad69b5226cb417580c1a4e026c590af28516
z460675d31c37a52144e7226a4cdd28d36464aaa401edea8d66fd7e0421d4d175f6a82d0c15df43
z3a227185925a2b64dc048bc81a6dc4fccef0d99935e08222401ab8c708e5cc9a995ab988c70e92
z8c078a2ce911a3afb62dd8becad4e86763e48b1f6aba3969183157dff7eb7c30aaa643b2dbbfa8
zfb13d6806e03f92f55fe1c6af479e3e899887b3e2a756b500b96dd965d56e2a85d63cc34c71db6
zd6b0a8e1d8f5dfc3e85c5613b0cb3540d5f40444ebec1016f8ccc74de70a81f984030558d336cf
zd4de95ac446d504072cffcb21b0aa3c6df64d600b45cd3963998b48120e1f60ce8459d2c0172ac
zaebae5d56841544a0a3ecd1f7ffeb9f51347f09cfbe86dd186527be6fc0547ad00537217f2c28f
z1edee26c1c3b027b2b45e278c1557126957cfc3a190db6206bddf9243827c1e7cfa2cb055525b1
z7749daa5457232c4eaf0ca68b4fbdaa9c83a8b59b11e8d636ed6273611835509a04587656f4afb
zdad6f647702af4f053547d92c91e38f255cdaf0d3e0676cafb2ed9a1d8bb15dbcd96f0e12c11b3
za24d11797bddc6330d7544443490c63d1ff331006c4c3ee03973bb011a8d67d545d4b2c098e31b
z551d58f418e363258a4a78591b12645cdb66bbbd5e986150db0746ac226ef407a0cbda63d7d3bf
z1d647a7cc2650dc936ce83ecfa5153138b9388add095dcb38edf39053704768fb5c08f03a1eea8
z3d1fb03e1bc0afe9d773478e288008612686bff374fe7b0c74e169056b65236d0907476ea32c20
z98ea4d2fefbe5f9852691f867479c6f81b14953fde23c6387676e4da2c71025ac9ebd880197fc5
zaf2ccc6be24f7caf880595fc10848802f7864712c91ac03805e55cc7788c5c9f99ea6ba1004286
z9469b67030282d054be16b6455ba35a0f68c098c6b3a9eab1744405eb14c7eb8acdd53755165a3
z736113bd434598a0df4861a5793640032ac2cc265e0b9421f31d1f0afe422868bbae82a399d1d8
z76de3527c443a1012136621d95e50324eea37cc939c6b6e9a4ae0bdef584fa5424e6ca83aaad49
z4a7089917fb45b671da39c5726884ee22110fb4ad1be690fe6386a48438ee1ec44ce1149f0131b
z3afbcc2aefc415fcaf533725cf8e819b2ee8a749c2538d4a3423ca3e48fff257f37188995f5d17
z7a5e680c1db4b9fc298002e0c16578804178f42a7a648ccf5331cd86feb3023e261f29cb9e1115
z19265fb70d3ca7edf0f4e7caaba2dad427a4451b3eb07897fb776ee966c987bdece385a376de2a
zc929644a8fa51e91d5cf2aab79f01f0493856e6281baf9708b6f9b3ff274a27a6f2e734e6baa97
zc5a74cb4b8e56d85b5dac43b2f4a9e187d0c5c0229508236fb7bc4e2a4096756bd6717a0610861
z048d370b98372f27bea8eafeb867c57b6e893cb7606e31f1aaff3c2734eef4eb634ade1494daee
z968ccbdd60052bf0119ae45d83281c29b4b0f8cc953b7c3c4bbeed9e64919c8d5616b73f6999ff
z348a8e9c747dcb224a6b90b704abd2551cad4dd50d0773e8a386f7ec056cdf39a653fe6e16e450
z7db23b9c750952020ca541bc29a8ec9347d91d7e7620198c454d466a155cf7ab0700674537cb74
zb33a54b360fae61afa293cf278ac15b22fa9ff4c59fb70438f10da79cf762dc2616261a10cfade
zdb3b2003dab0752fc12c792f7b516d07231352cbae8f4fb9ebc436082f20b64c826e3f615cbc2e
z5511565786822694759e675a26803e40a3d827e1f3ccc7faabc24bf018e1030c96c65fb48eb8f8
z78899b128e50e69a91cb94e0059d6ab3bfbee9fcbebc5d5053dbc95b61f24295ea49928bc8fb46
zedb754d7b324c411627ba3bc62e2c3c99874152875b99f3c22c5a7f36a432e71328390da057de3
zc330df69f5e493bbe7ba31389d75cf262645e7e6ab8267d3750293390ec6cdae6ff1d5465341f0
z53dda289551107f280793cb1fa77afe47c35c94c25bdae3e736d243c52bba25c536a06b5842be6
zb56060da2f0d4a8dfe70fc3388e46ceb0d16f4c81f465b97f1e38183cfa8f6a9f9285c96c4a308
z2f050278d186d74de6cbccdd7ece573e5bf5d479b12296468070d12da3f5934bfda369237b0d6b
z78b8bb73906f52d81ad347bef01e189a40ef116082aebe1dc518aa57d8b1b94948db5c96944317
zf1ed6231d3e149fbff726cdd962e02bd99f926f4675e7abf88ce27461c44fefe18ee70b992be8d
zf5f33d9906e2e7c9c1b00ceaecc288b181e5028c55e8f2f72dd421530ce78edd8a6e944cb8ce73
z9859639333a3458a3f66441ac27ef0f3166bffd06d00a5babcb17a7f94cda76b3065af52890b6a
z90b935e7b650c3eba9a10470861fc6c77b75547bdf423d3cafd9881b251751483006cfe2f00829
z48f38d3f8e6ed079fc2f33e1d4ef6f5571ffa8e17a1700cfa0049bf6d17eeb3e0a340addb6d88f
zd0257779d129ebbc83b3afd5e2cf0d16110fe157d0e4b5201da55b325bc1b30d058281f11602c2
zbda1f896696f3fcc7e5a2820055cf1ee2d74f3af0c7b3db9db81cc518b494d16f9a04f0bcb1496
z92b57fa1c89c9a2a9706e4dafbe743757da73c31d21829097ed38af6c5b5e884a7abf9d18c57e6
zfffc6a94994e88be9b487f6a7cab6e0e7ccb0e822640e3d78eb9d93d03a06b2cdfa2c00540d538
z1453c2f1c5757c646a6be1d0645bdaffacc1f4f4d14ad6fbf5e78c723ce4579f36f51b0c9d7f58
z8857ff1cc308bc3d93c197e2a8c6d09740f0b5c3c163c04032e3be3fa5598019394b186a7fea93
z805648d3456ea16fb400b4a76290467287a0f0c5b9d8052436e974a879f0c84202f9cf820468f2
z1e1ec5e08caa33622c0db5fb0b47c3ff5afde39925cda6817a9e1f2fce61c3022600f4f7897ac6
z6fb2f6d315583da4141b5861094132e7a2a02d1a3bbaacda720702f0d830d91693600f0a4e250c
z8c44a621f40c8044df7192dc44fd8c0f1304a288c3e04f04c953632da5a3cff8d4da4aff45b224
z375f2193c66204c8c7884d8cfd69dc4fe2dddabbf330ffe460e9ad1f12571a19ee3842ca503183
z8fd1c75d05febc4ff395ae9693f19a82ecb0abd009233cc25a611c69f3b8bd44adefb8bbe09fc3
za3a24694180c1f9eb6b5935b8cc69d9ea2be1bf32e422d543dcab0b85e4f2ba476f0460dee8cf4
zfed0e10324f887f8064a6a68398f96937d89e7186fdf47e72b2a8a5b069f393dabff712ce69656
zd7f0d6238f12cde7151322488495189724cbee411f14272f19d317fe91a5e24e346d22b2e5eafd
zf97ec316305e3bad66107818e4c265c3fb5b02874de5f42b4c0e12bbc86fc6cd8c198a957f8f80
z85202d98b256351d05c59a893c6ec5fad8fdf98b9daa5f3f8dd8de176e634423c1a77d50f3b472
z3f23899f940e6c9dc849e780302255b0e0272e0b155707c78419478f909d6b730dab60d9384066
ze4bfa047df29c38e2395a7f1a5f1219384f5e635c2869ab973f4a50be68f1896bc85daa10f930e
z8c26ab910a744935841401d5e13b68d509ce1e3d372d252d68da137ee7f0df3111cbc2663efec1
z9ecc2ce317b6c412178916aef22fd32f8dca7f881f2f43ff540168f4a6db33162c2f062fc6fc56
zfc275eaf165fd01cbbd529ded91f972cbc0ddebb6237b7a74b273a2d2443f2e87c694c5d793eb6
z10a591cf6af19cd574dde0705b00cd1def1c97a12e736af550fdb01d9e2dead64dcde58213a437
z24fac2a82771191b1b9508dcec87df7111035a0196351010cf517daf44d51775688bc6420f2fd7
z7ae8bc2154c3ab5cf48bddedf8f3c4e9bf706c44ba11463639d832dd5549fa8420274a4f6a5fa5
z41fdeeeb03db216abc7167a8412f54896514602cec2495ae14933f5d9342413fe0ec06104eeaf3
z116a6164581fc4d5ca55b1a13cb3e8766a9f8f162d466385900e435f623bc77e9e6cd8ecc656e2
z6766fa4619abfc2de379089acf4f1354c152d6074269c1746c3888c775639cb4fed6cf8bdf3ed0
zd7dc3b90b6a20e24d9d32143463376aa7d22fc4cd3e74fd4abba408705fe62f82b00b9c191c217
z61bbdaccbf74e8ac0fe978791edc9022a78482f8c1b9e0306783c6a8dd5b1bd279ed5ee5f8041a
z24dce79a131a22b9eea3b16939f51038940beb332ed10dff9fcf9fd6795d5483f34c011db6bf5d
zf22b5a3987178fdd7d2cc28d17ef3a59d7534d00ad19fc7b5194486073dff2ab2ff15418b5a4ce
z95b74c2aaaf157aff468e5c19237e660ad7d0cb94b07faf37bff4111de52298483964a0af2cb02
z781f6a04f48540a5c4f5356c508d348e4e42a57dc9344124245fec70c590ff15a61f3a2eb978d8
z444f961a8472fb2ebef281eb128422c505aa822980f4e64c8b50c03f9546f2a0af5c4af4c34581
z07fa3210b65944d085c2c80830a0c0dc8a8e177dcc6041f00e0c67adf499171f0123f66c3f3dd1
z703f72e5d8e79e91f527208ce44e8f9f889cf4ea9cf21ee155c7defaf4cc094228b315212c34ca
zeee93ac519cb0ee4d5d480c0cab2f61b8b9e3f6134d14f6b1ccb1a85986c9a16a512818c21f5ec
zd7ca46caa1d12ed4b9f8b0484218643f69937bc9be1424fa4a26019e2e3d93a37de43711f70c62
za1eedc1e27a80b5753c82474602490407e6367e9fdf3b520315d6043116f47ae90cf15e3fc4562
zb4b6dabbd1cb507d7135db4de0ab1a8248c79847b3cc786d70591f338232f26e2e60720ffc6c47
zfc29538c1440cb9b394206f31aec523341813616c2aa035479861e85482882c8b27c8d7340fa72
zc0c7f2e5836df2a99463ee1ecf6bd3e9918605b2e37f6ea2d39f96c487e24b0efb48828edd6325
z85ba0d248643a17c787d02043ae01e207aa9a0bcee7f275b0120ea9af84e28276d9033671fc697
zcfb095b6e9138d87ddbb634939ecf121b29023572221638a4d9f42602355cfce52058ceccbcaeb
z6efed1d8d48917d459109c6b5a54855bc0657fcf3c26d72d7dd19247c6b159d4fa0202f0f8c597
za32267ef1c183ef3bde2e62743b617ac6ca61476306a4dba25862c7f5685af01f24ca60fe99a54
z54204824d25087cc8435cf990df8a51dcd90de964fbdfece287714862f7c868e7cb610eeaa8d44
z00c568b73b5d46f0e8da2ae313415bb7e2f2377b507b25576ba04095d51ae06ddd0741ac0c8b32
z379c9461e7aeb4ec3efe09955b0a8fbc3841f6f87c5016d80005fa98d833ae214fe876da427a7c
z2ee633b0c0b11efdd3972931c93cd41f76c4af15131df81a872c90b097182896eb2b958b630b57
ze307ffe62386ddeaf77a7a781bc20ccf7128250697b79786bc49d2d7ee12f2fdc2e47aee3b2d99
z328b83c4e20a9befda7d9bc1ef48ddd0f84df7abe927c961360a9d3504a770815580b83c8939d1
z4374f82fd2c3f04ed7f61685fbe58feabbc2d35ef146e621ec17cad93f7d71dce6d38aa36921a7
z3bae5dbb98ca0d7cc6c9576da9d30fef45ccc61c061d50b5bb0abc7f595363e8f5cf9ca00f0b1f
z2335acb3b84b614b4964e2dac2a8aba0dc0e6ebe0403a37f3767812e03c43c3afd18c179e6f638
z7fd397cc0f74efeec6b1ce9b24a6266389a297e9480d8d0a161d3181dfbd17edd35ee3ecddf3ed
z126401715d3a870a1a4bb062ed162fabb4b47e12bb2d7f37adebd0d51e59b1c08abe7e5bcd8116
z565b2abd0384b7bebbacdffea73c71e381f06b1679d510adeb017141993b37bf1ea6677fa78c14
ze1431e79534f574f0201ade237752640a3f258da356486f90acdc3b1b5a773b4d2456bc650caa9
z36b04f18f73c99c121bcfffd8476d6cd25f998d48b449fb763243e1907ee255239b49797a01e96
zebef75609bb2927fd2c052d4c6fd02cb47d70c100de1df4b8f10014d6f40bf1d13ff7f976b7a46
z59e92da33ec648531cc28d766d773e4b76ba27f49e5aae5b708bcbd29614dd35a48d47a5af91f7
z3a5fb411cbaa8d80ce4063e1e61f1218c43f3d021d29b9fd9e439866e2d241ed028689c95b64e5
zc19c1a3c20a3a8065584b47816094fe4cd43c85ac27823b61c6213d8c27546ffa10ad653e32744
z2cbfc99e4d53300ed6aadb33487238252ed1ef9d11cde199d93c67e962fc851e7782790c5b872f
z6462f4d338c5b0ce2235aaa6fbc257a1f44b16eb860e50a344173b9f808e015d9aee6687d34f6f
z2d1bbc8f2edb5db268900fefd488accdacc66e18d6520849dcb332c449e472b2a57b1101010bda
zcf1441c55134671de824dc2278f9402db75a8fd7314197de8e3986c076c85244351560266ff0f6
z8117b4f77c8003dbf42463047e494a0e6c695d400ce74a5992b7d9b29b890a181f134b9f62789e
z59d02b8534f3d76e3be769e6565a4226886558539b0522ed9132f116ac09958f2609abbe8de1fb
zb565a677b4cd18a230851f3233b025d53201ca35e659dbd83c1c81c7b7d410d1ac572a1e47748a
z946ca8859600e3464138b2518c1cecf73a1855b6fbbfb8349ca3af38b19e6e0859c24c9409ceff
zfa93fdb53eb8caeb313024670671582dfb61b24ded99a775ac73f22f12ae60655bdb7aa770d51d
z2bcc94a8e932455188d13561eadebf660d8a5f8faca38a536df5d1911b38c2562b6b7b989e5399
zcd7b08d8522a59641e6efb1e0e506afc96e5e007ca3dc361dbaee432c00569956deabae713dae0
zef8653712bd1c7aa8e719e0423f2cb2fbef0ee007a56159cb82713619cf4b9e53f6e4ae1f7e8c9
z1a6e6be42510ffb2c37e4a09720f3f508232958b96b46928548847ddea0329acd206064f7c5f4f
z4bd2d4927f906a760b2ce6e79c7238fc724740f8af3b395657a39a8b8c1b076cb5f681bd2c4981
z2a76369b6fbb1fa4b9f12046f80e3ede8e65557051713d04789bb27fbb36cfa303f444ed3d7e30
z5f702655f119425dddaca8e73612c05b5098d0dadb949ec6bbedaa430b58b1fad23f0db0aa78cf
z6000834ae5258a36ea8c5805d0c121f2d5e15476f1a8adcf04d53845e4079ce599392a4c679e43
z16d1070c59c23328cc0c54cf639999564fd8151d813db48b76c8e63e429ed6eb81b0d1dee5a044
z6045fff85e2089c929a1f30a0b68ea7b05ae6b308d39864daf547a69b5ad9f8cc9f1d15807158c
z33e9e8116f14980e8bfc9e0702961fa4ed111b732efe1cceccad76691984ae5b08b1e1552c140b
z750717623283ef7762fe965e223fcaae198983cc5af9ad1972c705a5e373a174fcb2d80089c89b
zd4a3961d5bbaf41c39f9fe101858d7cbaf970b63d71a991d06ab6fdf211c98d9d2e667046aec01
zf3cee91db3c3d41e918728f4196a70febd751448cdfc00ae30f9332c668237935b9b1cca4d2d9c
z6a15859e59420568835a68a47d869458c1db1b923ff3bd92b440a7feb25257aed1a43010571c39
z3be4d0fe9ee0609f102e0f9cc85948758243b538150df276f82c852de160693606a2da4f6c41b1
z06ff4dcab73393c571d725cc1718150cfb63002ac76fdb1aa6ffa959f9b0d4b7fd13369ebcc70d
z485042f05eeaf1a0e06b365433016eac7d4901c3755a19728a0aa617f1a91f43250a7f63d7c37a
zbf7e1acd3a6e41f0d555b9f362888c1233158d874b39105b05c0130aa4dfef6b80817626f9cf6c
z1c7f8adae619a337136deef42b423a8b9345ad8df5546ebd53c93415147ba4354ddd5eb4974e58
zaade80fd06f2734223e7ef1b970243dcd5e2eff24c41b2ddf49a00ac5afb65bded260252f3849b
z76748fdaa2a6d1d41e9d61560b3fc6f7b4609e7a32f16d0d979c9a2ae19de106895b56589199c2
z8a514fbf5c5a91ef900d3d82b787357615e57e2587d4dc2adc0519f7ef9dfcd673b568c07dd8f0
z958348c71c466485cb5104fc34492eb16a679ae1f8e86fa03af4e03b8ac803b15c67758f32bc3c
z1b668d17382d0a0a1d82df9094a9ec09b88ccc66113b088b68cfc0d468b77bdd6b8673c85b098b
z8720765b1064dc0eee616e73fa5320e0646ee60805591529b1293688220258c1b733461b8f984a
z9b2885e8f1313fc12f6037489bfc7a5c6b10216b318d71c17cf6ff7c44948e586146da7658086e
z5519433c6889231747094952599e783081a26f5fc9cb53cd354b25bc6c58cf6ad459775d96e37d
z4dde0969d150686b2418196ec899cb7be50fb8c429ea7645aa501237804f45223d86d984a09aac
z4ff5f33cc476c1e970f719778fb0ffadc9081bd24df533ba72189f404fa5747306c84806f71306
z131b3ac9406d17aaf14c542327c32e9ce7dedc4391eba401cd7b2e48283172af4c2a8aac62a8c9
z52b3c25dfd1aeb0019ad5025c7d9acafdf5d4ca3fc51805f994bc556cd1dd40eacdaabe163adf9
zd17e33032e78e5c19f4a37ff8729d56a75be867e927f1bc3af467b8611ad28d4fcc1d2a66ff939
zef9ef6aea4b3d64dd4dde9fb878e304f65bf899046261b60eed0f7d8c1abb6e1352318febda6cc
z1da1a75eed46c38a8381c8708f7224d093cf6021b803626591f13eb405073630663db8de1dd534
zd33ff1c64f92fb6b8e3c065e206ab856ac7bb713ab8c9d242116800ed7e61459419dfc0e7fb07d
z2449188f08cdee03e661cdc08cc424fdeb6b2cdd72919decf87828e67d3945eee06aa15ece808d
z82c4fd748422257df7176338e16b6fa3b3a200fdcd99e564f1d7aff73d67939d57f19fa3606d1e
z5b1196ff862672b2ba3e7ed69ffe3f63d5541623d2ebdf435188c34358188c3275d71e1559294a
zbe38b6ad0141e445efbf13aaf17123b277c8d288b97130672b70c6ec8a0fa5f763ef6f9b4ace2d
z1929b072646f21ba57120a6c759e16bd0ff61f4ff6efc82470af43be940c09dd0b40490dfa0bf6
z0f90f38755af2ef3821d456f86803eade51982770d3e18bea52875408e0152fcd13a430f2eb3e5
z93ac442893f1440e122588e3c698eb232c949a7b593616074f7854b9a021295980c5de05fb749d
z33e0a52c146d6e75420c2b7988526873a0f2b138a7b2742e187040b88c17dccf0c4ed00ce589aa
z2ae92f602a2ef45bdb84b2a2f49d0ed720a6ffba1423533351283ba7cb3fe5eb6fb024aae529ca
zce9028c3e8de31809cac9a128d8ce9fc23cf918b88306f239a295c564bb9dc2b94a841454b6cbf
z58b1f60f54615d4e06951051d7caa2d6f0167cd14deb046f092e39c4fa6bea2b0cbb4919769661
zfd9baf2e5650aa9373c96fd6e1783e1f5350385edf6988040d133ffcdb9b19f53fff05072eb5c4
z2e9e3d299013e56a2227a29eaebe92636f69259acc71877882f29a9773e5f7f908667052c0201e
z13a4e32b3dc873a09ad12a05428242ee2dbf0017d146c90e5416a22b330004130831980fb382d4
zdc6cb99e32d6fae179bd3393e154979e6799ddbe4e548bb33768e80d37dcd43a4c300e0510b272
zff8a97d58710b08c667833c6500e0243f6d5252b0cf17f174b4450341e99027a351c014aea3298
z1e64f76f4659969ed975c2a94ef0e69cad7141a188e03ca145db88c819455abfc771998ff4edc4
z908f2571003f866e1accc74b61db30307e3eb3d1ab6d5bc512e086139efc94016993353b069120
z367efcc44ad66d2e125e304d8d84e7856bd9950764513dd9b6e231e43bbf679e6c52f0c06c4c0c
z4f422bb510fcbb4bde16f3a9bb3a96f05837fb08e2f30782cffb133e75dd31cd317efe6299a374
zda0a45bb48ad4507b317d88e9cfe9c6a74d305118e46aafad7da439904608804ac49cd2c148003
zc2db2788a7f605959922e7bfd57c6ccdedb59de00f683e416f5b629ca4134b2dbda0e452e05ed6
z4b8a4c80574cbab26ee3ee7440f1dd8ea6637feb7bb5e389f1833471d12112029466c171b74cfc
z9c5e4c42f299c669064aefd9eae7d19fe68381ccbc95d19e0907ffb576144171f32cf4eef73f49
zb7a1fc71f3d4602c063cf586f179f84290c7ed560a445aa38d0ebf5bc1b6814dc863500ea14607
z95ee51258fe1d75b406c8512eee2a485df035e8d0776ad99be4eda4b8cf5f21a7846c29c0f7b60
z4ff76344b1c9e932858072fdc383dcf85c4292adb4d61ddf6dc4285ce4f6694e0a8fe83fd0be4d
zea77dd3d08d1a57aa99da4c511419f5fab90c760801449c912a6f1dec0c3533953489c48753031
z3880e2d6632ce63f2399495215692afbd7365b7fef5225d114d532046d4063288b1835bb12bd5b
z351e8df2599179e33f1ed736121f470e4707ae8696823be9bae145caa15dadc6724c23482e4641
z97ddd29dde09c2829baa679c282efc07a9b988a493da6236af1a17ef4f14322592e7ef33136143
z1b8f10fdac93416e927c3e112c285ed677254672e6cd80e33351d1ed974158434f66eb1c826b7c
z78472405c641804c5712d83fb7ad26b845528b903f7c6ed112083bc48c32790f7a9305c5915535
z09c9b70403b72f79cf4a0796af7d2b21dc027ce6bf1536529d67e416a4a7519058ba2c1ada0510
z89327dbb6c8d180a802150999ac2c7ae8720d8ff4ff032c5c082ad28359258ee110a4c20d134a4
z1f3bddc9a07e86c44b1083ae15ad018851ef6ac7647cca585289196fc92bc1ff289946ae3fcdb3
zd2523e66b7714db4f57a19fe925912eaa2efd095e71828df4766d107042f571efe6c57228c4473
z210b0e618e4644151a69578036330b72fe46607440a1f219543a338d45a4f2cee2f4a8ea504a48
z16320954bd0a4ecab56a4d970929287a4c189676f3cc31bfc9f70d4665f7a04c2f3688d0ab6708
z936d4d1c6eec2d0f4d7c2fd549c2502b32dc09144b7268a41e78872996af22fbb6f2c8c705663e
zb4a9c4f0433681c74f57209947c19f034a01ae83dec55ed1375c9a6e1340570fb77c5a5bcc7a32
z517dedded6b62c35588442d378f96ed4a0440eab0c0fb56e8add65e430fca2fb66db66921c6c2b
zff89b4e5de24630034d5b5d19fa9ae3697c90b2bbad9c436ce5df91e730c5120ac8db00ff4608d
z03519c2bbbc01a494b0c5290d119607f28a1904601a88295ac7a2c6efecdb13f9c650eadb1b1a0
zcdaf50b6817072c365598d017057ed5e6de0328e4407b4c5102a94b659807bcdba77e25ae1c260
z8bb4b7388d6a4cddac3e0b68cd3268d34e528957ba897f2e4abd8e60d6d5f437ccf3f982710019
zf15d734f00c32ce72d553e1d054cd1616b0117522e35547448c2e7f43ca59a7b6ecffb5c8622b2
zc390bb34033fa215ee415c93bc10f1964e9ca522e82e80236be60fdd47c2473767b76b0aa9ea60
z5c031dde8523b89b35c1eb9c829e1e29b4a961cd13950eb8274fbf213788fb123464d1bac709ae
z62cf68a6530f355635f4793e26d2de6758aba3c8c4dfd9128e3e876f76d29c1c11931a4433df77
zd330108bd2c31a39a136d2ca02debfc6e996ebd2018966946df0b1feea9ae28830e372cc5ac043
z47cc52564e3490407cf6f73c137d9065f0cb62f2f7ecac2d7e616024af043e56fb1dacd45e3560
zf2ca4552b5eedc5dc22c4e557bcdd40ea6182ab321d6b18bb6af6753c69825f42c8889bcde9fab
z04d89522ad894fbded4aefd8b8e3a42163a72742191141f8f450fee3b7597c1697d722762eee51
z4f7bda53d63954e703190a08a678bef9236f75cf8ae10a542d95ab68b298c97dbbe75d0aeac93d
zee931fea07a358852549679f0dc141c7e6acbbee300b3d4e361cc80f642ff8043eebef38166fae
z3084ff5d00a4c649f92a84cf74714db11b284f37dc6510e24cc394d20cc705e29550522aee6fb4
z97225bf08f2354dd21ac9e3c3cd99601da028f7b497629f36217e64eb913b3affa387b5ba8df8d
zcc879a553bc8d41ec82eed7a98a358dfc3c677319ac24281d58741fdefb397b2016233886efeb7
zcc32c0f0236ea4ba1e06f025fe32e872603498c7a94e170cbd0462b2da6910f10650deae90f90d
zff10109c2d5bace2025557c28cad077f97242ce0fe6f8484fd3e43da8c45d1714d9d7a08fe14c0
z0741271e14387912bd80d214ace81663b65aaa87af8e2e1c38d093ef216cf0db1869ab14b47773
z40f98eca1090336e482cd87772d4b8a4b2c288f4a53787015f06ec55c83003ebad092eb09e3393
z62f4321783cc62abc3d66c76fe2308319e124d12b0c527d6f587af3a87aba6a80472bb9b10cc66
zbd6365a31bc2ae2b0e373fcbc21257369e689ee33faf72c709532a2783d01aa682f480fbfca628
zefab9ec3398152dea2336fc464eba76649f69c3806ea25f38db38f76acf4feec2995ca107fbc27
zaf72b7a4ae1ea0ac7ec362799511e61d471d4457875882029a8352489cc7bff5e4e5646a6d4e00
z4ac348099aea623072846e24eecf18c52edee88c1f1cf1bfb6def7bb87fd0021c48d71bc39c08c
za9e492e58525afe01a0fc97a9857b8185a354b53eac8241d1c86b8807c5e5a35c445b838b80f29
z9081abd11f5f65a0cfd6ba0963389cf2cfa533c0fd360f78638e6569412de4b77cec33053e02b2
z5f411a9996e8f4dd36dd6001503d17f6d626eb4af29e6750c84d9f675d50229e26a4b642fd3ffa
z2daa128baac55f4ddc2465d200ad18bdc61a56ed555e927061ec09d1a6d64191e7d723b6857478
z0e581da9d61c44a50990202e196a56d9551367456436fba82c88c93d4946b4f0852aa1e4e06319
z89767dce5dd6929b90508e14d9379a2fd757c081b5f3f452fc24674bf476d9e17f361c63a2a754
z0886185d3ea4b6175c82ee75e13b60c9c84963889f094aff7ec43d5aa39ad5dfbeef2deab9b523
z25cce23c5e80716b0cd5ba2224365986c207b2c2164b53ec67edb65d990dc460946f9cbb651858
z8af0f73596800c5d0066e026ff93b43249d3bd24bcd28067fa9152db9a7b8b46ef0d65a4285520
z5801f6510e2236e2b0dbac39e76c0cbcbf98e9c02a75cf8d87a24cf1fd351b21f2d5a94d989384
z3847414c20dd0ee970df4d539c1e2598b7cd1fddee676f91fb3b26a0fd9f44e0d2215774f279d8
zb957fc888fd731886fa6a683a8571c0d7dff5dcecfd76f01162b3016795a02a5e83f7b2a3031c0
z2c98acd2f60078f02baf496700b3884c5c5142ad2b39a8a033bf03a90c5b57cd3ef796792eedaf
zf9e17671b7f1c70d37440a110e23da9620f285f74713ba7ed5fa6c6b3c808c843b80b6e8dbc987
z73ffd6d725c39bd865e6df7086f63364ff49a77cf17a798ff59b38ba580e3f15047fcbcaad5e84
z67644383ae5c6d0dd18c03c2fbf398b26fc5991aa17bc5a71f76a6119dca4d7beabc110e6669bf
zd9f3a42b0f0d4090a6facfab93773318283cffba74e5cfba6df0c9af901a34c307129d599f6b82
z6c2f6d7ffbbd480caaff2dc70e3577487f01a936a640bac2c68de9e65629ffb0c70a9a5d911632
zc35298cc77bb48fe4bf8f5bd4b1a3ecbb557f0cbc3536bf3a3ebcb6a8c9639fbbb101aac4288d8
zc55b782689a7b13d22e0decae6e35a4cd6341db83cd7b7375a8fe90b587444a73f7cf992302a9b
zc1d681f677b3ab430b7c95ce0f3dc9f7b7dcdd452fa41004dfbda96f4b9d0e4e520ec2705c9362
z283440692c3766996f1157827b93c1750862a4b471364c4875e548a8af78c6d61a65290ead8cfe
z7fd8810b4cccd510309d8035ba244f6fceeb6b3509888d668d2c1bfb6cfd716f29d1e4a63a0cd3
z70c27970ffdb5f7da9c468e8716a2a243a4d529f835b095940270e7886e64f123a47e17bdf8887
ze25fc36b550f843c97e1e5d7ad558b3aa3ab7a99df62a815bcd7068b5b6e3caaa0ec3964447ebe
zbc2d8c0bbd62f392f6e42fd66e86a1e14de1af080ae803104a88ff5349fca3d5697bd1a6fc4104
zca4ed376ecddd220f6b4a0b28548ed2f71ee35fc0954a44fcadd235109b37682450ad56a083096
zae0d2d2fef297d559315cd69a5caa1d61a2277c448897f34920a606e317cbb040498f02f05cf01
zf423ba270ed16599791246e1a1171f8690add2e036aae7eac1d0dcf7c8d17c6255623fbf0a6083
z098ff2fb1436bade3b7fa881f99949c477547d51d8b7db543844391cff2d223fcf97d712044348
z403d36db860175f7f94724f57d7affcf52b78cd3f3f32253b0d86b011a6d270159b87cf7e7bf1f
z6b6ba162f22dce5ab61c5c6f51540929454e1c027595657367be0d8ce5e561429560b7a77acf4a
z5e33146d857326c4feb0caa088619578377f1c5c300586d5f8a676c851ed4b90d88e50824076f8
z43be82fba1844d37df2ccdc3c6f87615fbd1ab60e2e30c1d43ac8d8903c7048ff898752aa38c50
z4d4bb5a5486bcc7b0be186056fc1fc661f00850757992fb2f2f330e39943ce6be32f71d80144cc
z18e530e76d33224bdca981719d33b708253a69a5b5a50fd1d8903058c5fd34e5eba20ccbe3a144
z39376e978ef55d92e88aab7e8dadb69c737b57dcb985d550b68f26ccf1e501a81313d7319cf66e
zc5a5363795cd5efb7d770131001d37f5a517fb56e776b7fa4c35f45336e0c54ebddef483f212ec
z0bce65c4fe102643ac4ec19575155f36eeace3ed371a63fbe09f0ba8c34bbade76dd3c3a027acf
z147851618c205d571062ba2aa02a3f9bb705b41c039733394d07758b49186ad61a41698b8366ef
ze69a1639a2f0d74381e424107d21a130b84df83d8e1fd7283b5bf3f7c8eef9a7ae45ee1ab64f1c
z61c6e75fa86e50c5486792beca10b68785777c4004dd23deb82dabc4b559b28130980ae3a26c52
z96d33046ba9fe989e958f361ed7d7b2201cd4464187aeb87ea05daef85750f5df1a19eac05e823
z6c64a66a6c4402fe67f9fa5705ae5eaeeeda07ccd14f27a14882ce55e1255352596626858c10d2
zc6ba8143e27522b2d15ddd2d9727332650190b615ba2d58038e6065c9d23e1295eb80843b9c944
za6a95e2ccb56c698c6ab910bc63789bd81987aa526bb03ba73f516f9e448ad63a0dee102ba6f85
z8710d834fc3505a7d9eab3c9af25f2ce8822118db8451028b6c6156909d6da1e7b36e33e4bbe5e
z0e08ea43950561b37ea630fa221cbf9ac8d1631d7faf86a5638fb60a0200a676e7e3983f75df1d
zba697cea746f41550791657e973c554ef43c6393440fbc90900ffa15cc4f4e12e6c671cc37e84a
z2eec0f6d6dc404a17551a8b46d098c6dfe48b4ef88ddea2b15c913b21ab814bb382122dc0fd89f
z593b96e16e2bbebabe9338705c4bb2336b9d458dfbf90dff08746b62370016da70050c0bdd1380
ze2acad4948025bafddb9a1ced4628da48d22875f39ffd8e8c863a8d9956405e131448016de33cc
z8fd6cdd135603bb79afe67b5c2f417cf8f25b0183e2cd2ae3c41e649e2610227fa7fe8da863fcc
z533bf91d0623f7343b20b97f476624b35846d00d80ec36eb6e1621f2eb6aef8db452e41ccddb38
z8067ec2f2b5c2b4dcd19556c52a94df5d679be3f4f7f106dc4671140249d226261a1097d764034
z6872a0aab2baa7e5d0a80413e6c0e40378c2b00b08fffee4d926f218320040870586ad9c0adcf7
z563ecba858302b91ea1ba624712f3529c62e7078dda2181b4c3243f41f7a83354aaf0c604d62de
zc0c117f97dd37d615d0f15bb1ff2c7534d4f74e3e773affd8f46c76c728bc1f091b29c85bc4c97
z649822ce05bd48479bf6f2bcb5b5cb70b3c02e54805fb34e05daa89cc65989049e20fa7141541c
z92b79b94f12c17eff91b7b91e63747a51d97f4f409b3239fff7fdf07a275d85ef0f8a8500b0e36
z52d13be9fa875c8a9b56749f76b629c5155303c597261256a175505737eedb9318b40eb0fdf3a8
zbe8fb8340663a2e46967aa1e5a2aeaf5a3d6378da84f81b90b8bbea9d9e782289d5b36b1f8aaf2
z4ed1582f2530907493e07265327f4c0431f5a8caab7b523580c3369bf1786f9fa9a6e52ed12403
z9d977d0cd92684f05f11dcc982ad9740c9502b1a19f1e6047dd6abded055b5fb68a8b87acd190b
z25851956d7e0d7ae146d4e1e0ba559758e34f90d772fd2131299068344c6aaed19ca7d5fc28548
z8fead369f33f3cc09bcc9dbdd20c9f7886b06d9e0b49ffa11806d9bd42446659f5ada4e74eb33a
z4656652a51812992d90f7ebd57d8e51613d441af9357c638a401bb8d8476ab4b30e0dc48a513f8
z544c6be5976cd4e4f812320a42e10ad14ccf5fb224f984b9221379ee2054b87eb7b815e5914bd4
z2444529afb4a87314943e83ba5def581e98a35e4c5eec009c9a3be4d42b709f81aa4663af8f019
z73bbc7b3b3d8ff59849ad6e4fdb7d65cce16730dd3b2aa04b9fc2fcf6dcdded1853783decad0b2
z2761963a22bb386cff775b49d44a2b140bde184c5e931011c487053b313a74ef1bac5d3341deb1
z8a16e0d9befeea7b9efd0974c119f7620871d742adc476c1185fb252f0ca6b6c67a9b186da16ed
ze570ad61f49301b1b9d8123787e8b2f882496543fa21b7b287fa55ec4e3c843eb5fb0af0fe2f24
zd71b4c40ed4bf79d7d35025df1e790213ee521547173f72396a682ae4d44890d7d71a67def18f8
ze32f7e551ff9688d6f9710848918655b7d94b0ba57053a6da1208b0d2ad7d3ab17941c870707f9
z7beb54a8499284e33679d57dcc4e4ccd8ef5e35ff02524cabaaab142d7f4a8e7727098812e46a2
z2dbe7ed7b2f44a0a6d1ae8b6d39d873cb380305003c5d757d5883ad7d21caf958e55b8dd1344e5
zb1a8042e9311737f4ba503a9f8ecd2c6fa9e8aa17febc147606d7c89d444c3317293943e35b273
z4dd3a3116b17cdcb758cb0fb174e13b411e1794c86ac21fc5192ccb7ef69a8391fe95814d219a2
za15a05972de7cfd1509daf97653ece62c5d6b829f87f48fd61d1dbe6c71f1b51b83a6866121677
za67647edd3f61dfd03230ede326209078358d9460faad2f3f604a4f3ad72072d36b76ee2323c00
zbdd2cbc15fbacace9935e6847622355bac315eda2a6d32a532cf9d7db3937b143b09b046ca1273
ze52a1d0de010d3ce45f31d3a23cfb2c62c5db7d298f63d50ef1c6f3ecf5a901aa92706a18d9e45
z470c23ae2d23e5b6a20276fb07741ce256ddb5094570271ad827794d60beed2f49cbed4c608764
z50cab704670702bd6046e0e9ddfa0ceeee2c126ac675a7c4055c4d81b71b03a13c88bd5f568049
zc6e0b6d7924d886454ca86fb7ec322525451562c2719b4c645e9234d7793e8b01c1380919a89ca
z26cb03253be3bfb4aca1be412569fd080031f377b7d35fd03e6408b9bc37a74850db6f5eaf673f
za19a6350526e9286621d6e2e58234f4f22b69d1b40076b2cf6f6bfd9bb7ddedd30167ca42f7b57
z4689c642abdd5e2c0bcc2225e0381143cac76256903aa7b0aa2107f1b266db6fe820744b846781
zb0b38e69609188df2097e356dbbc1f073a442aaf0c95766fec5881f83baa5cda6991907ec6ea22
zcae4d0cde7fbea527bc0388db64615c7e42d490046844a38e4dceef77f96a1d6012d3ab5e6b417
z57d04b33fff325152810e422214135e652623ce14a102bcbebc2974228d8af10c25b8f205c04eb
ze499a6954913081b1caff968d11144f1eed89fd7eeb74e21c009ed0562c3868ca293c1772d3f6d
zdbc4715745e5416c3356b6ce5bac6310205d60005d58d8a4b2c1e81895d18f9fa2a0ca2b0b3f98
z2f23658aaa7fb19e3e116e05f33ee137eb55282a7818766254404294256e093050ed245377c06c
z32c7f03e01e68eb6064f8275513bf7aa95fda6cdb820040eb54af55470f74aae7150071b6190d3
zb8503b20b48bcb391683261b329e04882622abe8323aebad5733a405cb2d28c0209a7449ff3af0
zd5f2be083f303b453c6b278d439f398460c841a795bea14797439acb0efae31bb12c62ac10ce63
za824c8f6c34adfb82919f04652889feec03fa77aa5f6374c4e0d68fb0e0b0921424c84812d290a
z2114a6aa3420f48dc54357d00dad6d768ddbc4b3482b2d0cc2fb676f1863fd7b28481f82d9b5f6
ze8c03b775b02c9ee9f33f31ab21a5e48ae4b72cd4d9061cc96957fbbfd0f96953f6e0962024680
z95f3e585656ca45c99c2e3145cfbf3fcddba358584bacf415daa379c47ebdaa0447f96e051f71e
z9512ea02e2359fa79ddf863be957beda18c5c938dcac8caa90df9fab3779c331fe9fbc4f8dab46
z7d882b68b17762f9606003fe4568958fc390345d763b25d2b2ed3d8d100e50f2ec158dd2186baf
z58f3f3398cb36eb3128f6c9aff02bf1c2e8cf5af30c8ca6b02c6277416737d5539a5418f60a2ed
z98a1c168f49b2fea276e56258f8c3c63e9098362bc56828cae5abe611d50ddfbade0c330321cca
z0bfdd2ce69adfa6ee2567e76330b77f6eab8926ca0935421c7e933cca3f0bc4fe8ea8633720804
z5844baa8608867d1b0a7117c634af84f1867df0c91d8918f23d5ab6ce6131ab2241fc63da2ed99
z12ea96cf0348e19603009db0b2210f35de4fd69c2ef0cf64c361ca387ef43a2ad67da48348abbe
z0cb5dcdf55bfdf39ef5fcca4b6ddad7f54241f18a642561f7279c671472b01c5210b62ef30f198
z00a26f0bcc6b8413a63b2bd4e63057afadc3afce7fdc51becc405b95ed396044183fe2e4c475e1
z87dd8a950d87f34b5f1cd86d58bb9f687cad935cd82e09bada5f319eace1651126c658f50fcb04
zb0343d3de1157ecc308a91c6dfc89d4dadae52e8d5633e11355c5674c77f7b2d2597550d89284e
z824345f69661244fc96b627fe75e2dc497e8ed84e115060b87b17358e73a3be34e2b4574c2acf7
z1323150d64c2e82f9ad7943ab1f7f07198b8fe7708f90371d14bc57a101fe6c573536878712433
z1cecbfa83eb8600986f5f14a5fd928a516cea642d332001717c1fb19a7950ade9ec83dfc804619
zefd1f78a035500ddf87f96f8bd339eaf8cedac27e96c1e97c3292dd21dbcd4fbd6809e31ffe9d8
zc049c858fa47dae7c13d9e806c258e49e2208638ae87169a6ace40754407a00e611b8bdbe943ce
z189815ed6354e83e3fa75fa8cfa279d930c7074f0fc92f05f45ee6c7fea123769f3315655db4cf
zb8531b6c0aecae1413f68004c1ca47505bf40f5f1bdf033758c8b90c7a6b6866d520e8a8f238bf
zbbd803e965277b1b849af273f6d8bbf5124b469bd222942a74b9334fc057749895f381675107b2
zda32e235cc29e562485bc3de28707a624810bd3e1298216e1845cb7783c42d5dca8adc3143eadd
z5d4ea37ab88cf3f2a07e4d482bb91640a926b315ebb742690d62e228efbef625e25104d3c9c711
zbbaf79663389ad07151ff145451ca88e807bb3dcdcc903ec5fef915ad8c7f65b6825db7c8a4bc8
z782db738c39c5c9deaa8c80cb34e4ba5c7a88a79285bb2dfc9100f9a71967c0194693ad85b5d12
z69e6cd54b9eccb9d9511d1a35926c36f825694b6907338d53d2c084defb9a708a56e8c53d0a722
z0c01362ea14e02fb80c47d618d3633535cbc1926ab6f1daea0e64979651687a9d69e2ef18a8ba0
z928751503baf0788f3a12a2aca070d8c5208f47aca3702fc5a192d9879d32fc839809a5768c0e2
z5370cd161298a0824fbe1531a83b7cddf241504e1cddf708dfb72a15302afad942ea198b62c2bd
z1113a8432160eb7fed2e057a7a68a04c42b50c86fcb097b088d1dab4a51eb4cf8eba96c623ddd4
ze5f1e423d6bcb9b593ff049e85d437f50dd1c61043ae4124a88732e9abfd58d27314f12477b2fd
z8fcd904d1bb3fb8f2ff61f836c3854c5f556b23e42f65b3bf2a040116567cf22c9cfc484c9ae0d
z3e438a44f36db3116a27e724bdde0385440d795cfda39f82fd9570dd2be62e18ab0999a86c2d6f
zf718a4a5a7eb2280183a49683532228ee76159f84e3a5a20216fe9ae376337c3c2685af0227724
ze451b27479d0f38650fa18be430dc7d09c9714a3bab56f62bab00b9dbd4cf249b9a6bcf4b7337c
z43e8b6c54ca854aa8d0c2d1a0d2b4ff35ab3bfbae1fa044dab62e3f2221c71f82522043c527182
z4caac33ed8d0d864b26063734ebc2e79a778c79c7bc4fdb2804b720420c38aff7fb2288bc468ee
z096dd0ae6dcaca5c7ac784bb549396afc88c4b892476e18dd00b24ff8254e4c9b010a8c4e47ffc
z4ec75da70f41ceddff2b51158a874dc73e9761add171a11ee4061fa1285944d46e71b638e706b3
z4b0724d15db04e13724e4b3bf11700292dc62ebfc8f0d569ae031f8eb6b478668f03ff70b8cb6a
z2669be25563a93efb6181e9ad496d6ea028f0b16a5422024fc61f94cf66f03c4eeec46cfd6c8d1
za4e558ee33cc97e0574f13a1435b5a686526303903d921901581153aa08d618d6af3ca9f184219
z88740a8fd6861c734c0ab9cae7d2bd1f9ee12e8e5b8337f9a0735c99be30c0c653782750d398ef
z6a0158c5fa52e7ec4e48009d2e19a43e522719165a2d1e9a8e4e5015abfa0e0c93fa29d77ab7d0
zea2f4c00990bddbd919edac8af28c5a5b3a8267680a5243292d562776124e975848c63510c7e2d
z00e274a872e5d0f046d1c898f13ee75cd7b0b00a1ae539e9c5d773fbb95ba1409c670b7e22e0c6
zf1596e2ea1f484fc571f169ea2c18b342f83719365ad3a1c6dde5c67d0276ab0bfa763b32962ac
z7f11f794e398ca2bc8b924173232a7c46c92c89dec7733ca6fc3aca0bd3e90f92bfacb523ccbb9
z412f5487f285f5b6d0e556befa08877d31fbfa9c0a56dd4fae5d866eb2020d254f362e57e87463
z9b396eade5e95fccd12334edfd6c1e7a9647c8939010e7fd49282c19d8fe813f65f12aee144d8e
z68129d752845f581b0424bdba270bb9f1531514ddc748d95fb8863da84628b7292984af7e43dda
zd78b3e7faff09151431fa1df3e59af25ff647f4312ee329e6fe31fe98cb73cd9c1e7945a87af1f
z337c055cdb67c6f5029c54165a5b3ea89c1bc1895e7ebd30e37cd81f5c9d4cf05370a56422e5a8
z0e9d2cadfc3093c3ffad97719ab2795af7d1030be63a8dcee4ce690aa15edc306a123051f1f68d
z4b3b1b52ef4af9c41dd98ac00edc7cf0cd296179fe99703239bddf9731e044b962c09f0fdfb83e
z649fb04f776e71fc8499599a980a5f7dcff6a3dc06b91b2a3af2c2e79501e1da27ba32fee2616a
z91e0ded474c8612853b369c26b00113a72ada00181ff374974d0baa4b2325d97eaa1bb528fed7f
z374d691141f8c395437315911c140f103d99160d18d43d4cff2e1635c31f1689df3753da9462f8
zc3c9497082f1e4f444d855757f4a4ef6ec33d63ca3eec2454cc14602150ce8bb24802e1b83f533
z34be7ea9636e370f357d895f43d76b7b9377cc0d023f895af60444ebd11b6f2c23fc8cc1db0954
zf35539b3f81b3658aec7cd414b8d02874fef408472f49b6967c01e0803aa2f24570f41598a9624
zcab5f655360c15b556c99a23d061b896d7e9eebd1c5a2357ac3bc97b29173a5dc2b767c55e1bad
z52bf33549d40101c36f9a22c7f45d34d96c3a751788975e82835440a2cab45727cac2666b7ca3e
z1fbb9204fabfd44caaed8a9e192841fa5988a2a28936bbefeaf6f10cfb6f59cc7103c29b71ed14
zbcbf36ddb9d9f60405af122c54be516b5f92cd0a806d38be108874383a71f3a3206aba307a3fcb
z50cedd048a91579642b34797fd351e1cf4b3a6b0875ed0af0025405328cb0741fe302ec9af6f51
z53148e2831a06f874a50cb318a947ecdda15de8d09832a2478304c2d30e64f82b31e4fff0ce2de
za9766b5d3f53b51c94bd6ef44d749b9f7f291f89341921c09eab75f755627faac6d255ec95b7ac
z802194db813557a545e8ecbd133ad725899b016c1e0201a8f393547203714e1f50692cf34ef782
z12a8ee3b5c941b9eb0f3c87efe9020252935a89521548709f44d7ae8609c2cd2c79898e6fd4f48
z03e364bcf6e780843c7910c99d7dbc943e1a4b0dcb582c0514b071cf792b818cdff8539a9fdcbf
z10bc82ae5fd8c20100d10358ab5c47dd6c4fafb858c7d02638e6052025901de9639db54544f177
ze090c20db84497175bea16235f24b2561fe0eac4d15969cc232addc5c0a1c3ff61bce72aa27747
z87abab265d9e5a66e3611524395e0040e15c9244ee08daf6b274580c4a20309088c4c2669ae951
z63411e2e7b08d40f8e157834e2952d96d3ff76911b0f0f6ac137f42eeb5d1a95aedb6f276dd1fa
zdf25b08452a9fd39f2fddc20d9f44edb7893f3469a4bb853d6bfabd75474264da068dae6efe90b
z967d4ae4ca7bcc6e929ba3179dccc49a1bac95342cafac827b6a31232fa5bfb862ea4bb38f7789
z490795eb028e57523a603bc55610e87af477e4a92f7aa2552d9768fd01162b68c69d83b9123ab7
zd1fe8e37fb6a3591db79a3edb22231fcd93ed3d770c04319653f30f3decd7b47a94a8b7f9de9be
za8ac6e55e4ada2854614779b42e3c2971e30e760eff3a17ced82810ebbdeece1000314621bc6d2
zea1f843dde8a11118833fb1a639f6f9d664482e31eb0064899464b1577e26ad5147f797dd4d3fb
z587529b4e97e517d7ec1e8c391116cb9d299846ff592bd5a6562017fe43ca255da25328579f32f
z725d0b0ff24ee3b78a6c567da8628d584c46c8c8276d5cc7ef870674dd36bb7fc46fae74280902
zda1d78a71ebe5a5e408b33c8e00e4478014dae0b22f077197c09a86841a55e3309738e3b5f1b8b
z82957c00d7d4dab6e642ef9e71860c02f05688101ab5e5c52141f7160e82f72cac767e62b6a303
z6107d68172b4bc341d1b71e9c12a699d7d7dbfdf7679e2a091ca48f09d301cd141bbe263eaf267
zf0b8be251616dda9047ea67c963ad553a2917f5832d75c74b7742187e0f06a02e8aff731eeb0fd
z05c72c61fc15dbc4dfc11d51f683a947a4c8b4db8ee8cc29ba5c00522c19c069e29e08133929d6
z869d3334f308bb3af0333c5e01ecfd4306d2cc236cf9a12fb993162f68810db52b6539aa817eed
z0cdb15050a6c6e56a859a35b95ff20511cd0958eef3b7084d8908f3f96aa2b3e0f5cc19d700549
z76cb961fc0245efba48c388a20a1f707be9a69df1f89c49ee9c4281cc7aef4123de384a9b2a633
z0012ee216a301a2e7e53c6bb64c4725218a410713625607d5938a22db54831211df556a6da28f9
z2ac6c866b8ab07c03f4b599497ca0f273898d8118d135b71f442670072ad6106df65f89fc8c5c8
zac63e941c04b7299eff311cdd5a683cbac22459b8fc409127aba15f3be35f480fbcd21d7a7fbd0
z87a39ae49a4eee465bc544384cd33b5ef371f0ebf33e3edcf5216e036e83df88e324d3db8c6523
z4bd4fb162f59a51965c5e422efb005095bdae4623a5a1abd8317b71f676ab20eb4dcab787f9904
z3cb424577ebadeb1aae077111eb95b79e43538cd42f87f7624c2093c9fc9e0dbb165d9897e0e28
z24adef3672733fc6487669eddcdb3259e8aafe835842b3aab7c95dd98189658ab85587b065f61c
z01ce533e84fd25a42104dd5bf0e94cde211936b41931e663d81ba80a6578e2ecffe6db8af061d5
z91d4b11f24ca99e60e0dcdc335f88568264f8cad2e1b9b5276e76506387a26453de698d488929f
z161509337b7259eb0b0ac3057087243efb32edd9337b91027b96b0bcf6ed6491cefacb12eb717a
z67b63f801459eb312ee12c71f84172caed816e4a74da19ba0b915a694b21135a81f2d9f5e7a633
z5c5c42e8688f467647f59379cd81415951f65d21db9d2aab7c2791e7a1c2958f1ba65ac3036598
z95bca06f4ed9e3b584ace4be71a0a216b1cd0f2e5231f942c5b4ffdeaac43eb077195008812ffb
zdee0c4b99c6f4ad040ca9a9adbd182cfe01f41f53658540531004b78ad62a7fc84920a2f175462
z93d8993c5fddb2b1157a1b40c4056e8e4d24577f5cb1fddae91169d6a4c09188b15fda7e717918
z8d7f6fcf4f61bd6f53991bf9af01b6151d8cf9f8fc2e167c8f7b38e11a34b14c83f8ac0217650e
z2b2924d8b6be15cbae243f03c6a808cdab1462f5d322fe2b6b5cf652c11431d18e7a62f20f5b9e
z9c798f5040a0d29a4e80d457dcddfb496e5cc5c57a0a1c81f5c66b4cde099e47e9f56852cb2200
z630569af3fc1ca604cad233d4a5ac07fa0b9321b94796e2083641ae5513d8c239440a673c38b08
z53ef37b7601691aaee53f8c9c6ecf56d6e597c032b410da2c6b6e7c4bb0e601b385e2d04b43f8d
z888f28a9264713be15ff2e57ea57649bf45ea90a3dabd9cc2e6943e074a5deda28566832f467c7
z79065356ebb8e7fbcd52258884029de478dd8f03ef53f9c830ed0cf608a93bf933cc8c966e9b5d
z07a518a54f4f88f66745b78b2f4f5dfe461907a3e372093edac72a007458f4a17752b252975e80
zd8d498f3facd884482452efea64f593d8b07b33e8145b9014d5ba8e619da84cb2f545c4ab3a8d2
z59393884022ed4be7bf23e3aaba6cc380474320b6cb9d636fc6498978f1593617394964e46e4c4
z038b7d0af44e11a104ac6a93f9fb98caf0404a630003c33161de07fe647888c3e80b2e5e7764ad
z72c730d75fee1602265e26467fb55af739f96aad4e3e0cc9f966b958923de3bf4b23f4631de470
z953780c0ce6e6e3c2cf26713301f3482a46c0c93e1e6f354663fc0ab6d6d2bdf63f45175f3a228
z99395012d9dff82a79d6640580138c64ddfbc401a88d72c440c21883980532b809bc6d486d7fe0
zb7f1922222ae53d3bbf5b3bca8fb7c7930a82fd725dc135862f523f2b58223d2539c31037be13d
z2f01c7fc8c027613b26228cab2787cd9d771f9415ef2f01879c157f8833984f950dcf230bc3ba0
ze9ce6a4fac8d4b09d179ad4949078860a81b942554844472c4cd8fc63458067403e5b94701898d
z5ace02b8c4f93c4b180b3b0f7cc7d6256dc9eb2560f83e355e6eee22cde79c2eb713fce463656c
z0b8a6cf2028a05af7f203b10c8d3de670fcd67fdab4d18877d96d47f51ed76d63dd6c27dce89d6
zc2f98ed0d5c8b9e7d69537a79c3a3f81e89dca6dc87072babc56ff407e657a7143111827ff7c26
zabf0a1d0a11253c0ab32d0f07a44e7ae3667f96b2d51b98a5bc39ae3c8cec7f0059bbfed0d67e3
z407ffc2bc0120c23a10a983ba21aca0dcab43d394eb6b5e20831a2edbc8e23afb6f458f11983f9
ze4cea7e4e31c276b1cd73f77354a20ba0f97b08c3450aecc8b96a4aa8e7b04fb770210bd59eec8
z805b98ce5a92e3a548f1f99d72034bbd58b681ef96b68275f33d75cc5d14e46c827f940a1a44e3
z01418704591a037da3a6d0eadd6aeb20502028d83ae95896fa27c58c2b2d30334c2f122bf3f6bc
z8791e0cc065cec263c30503f3fa14859b84db4ca9ca647e0339130ad44d0019654cd87674348dd
zb6f60ef23592d2e800c9c10f9f3eb243de510201d5054ed9a27c30ffd2fe32b019d015cd572e6e
z69801d28c9f429846ea4b0f4830f0f792d062cb178e100a395b05a72d8843b7d0ac41e50354562
zaa1b7561c166db08bcb750dd2596eaa6f2ec3146cd1743053f129221a6d164f10e08189d2d5f82
z810ab9842d29235c31fd357694b3e6bcd9f90f4fc84750b6fedf91066fd1a52b937335d319f82d
z479e18e3b478612bc6c548ac9d504d804362f5cd4fb0a9ef62a4a6e5ef735eb7de6d8e719050c5
z8d0a375f62cb3a931083fb16c8a2200dfc2d250d6dbc94ee0d4cfffd1bba0845ffe705cac532d2
z941f500ef9881ee69d99f1c3e4fc75b55af1c386fab78d03916c136181ab168e5ef0854114f035
zfd2b76e49110acd0dfddb52ca034b287cb24e53851c0437840eb37204644be1cceafd50d37780e
z7c54ac8668cf13edea3ca03b4dc503bffec6cd1ff3ee60f89522d3d130a054e292fa4c3057ed5a
z90695c2dd7658584fc5189c34e00dc5d5c5f3071e047b29e0cbd493affe3b21d73c6b742308e49
zb3267826985fa2468e2e0a2bb6537892316f6efe46a58d26fecf29e467c435c9f31fb3ddd596fc
zb542f99a0caad605887e6d41d9b52b32ccd47f5d0418e6f6c446a538691d6388b29750d77716c7
zb3ce6bc1ed7d6c5ee186958571e6be87fcc5c1ca45100a033293ef4915fc0aa37c403ea93afaf4
z6511dc997426831aff481f47190f6eb4a43a504c2ada743a991209bc2aad339d4a488936c49257
za5cc1d78bc4ffc52cfcd6ee6bb0186f09013968f9ad10c2bf4bc5a31e29fcb89ee1457dbfccb45
zde55278d3a83e0ae12cebece21b245c1794205d543a52f73e91104148cb70d21647a02fd5cec35
z67b1f6134b8b4913e23feb4fe0b1f59323051fa67288e9bb15922556087f9245bfe9dcd0ad4c2f
z9493dfd46b55c7d7b7a7ffa1ce3757a31ec0bd9e1070c9c03dfa62380d81b5713ecd96d4fcb754
z3886289e1a98ad567cc90697194f801f967961ee9632bac1b3227c901441b5ff2d1f90da9f8f0a
z2ad37c12f309a890eda3bf960f250a7b60cd689bcc796f6752aea33058c0c77e00753dc021fcdc
z46ade5545262e7dbc488a0c6ba47497c84eca854ae93d056e8ede733590e755514e0d6457c1210
z2b45600f67a0f7cf9357481e7e409045eb4817f43ac439ba79c9416d2dbf0a4d3eb9861c1158e4
z4809785f7c2d4cf03e1f0a1c2f422fd4f4e7c35da5fccfb17216758cd0fd82ffb11b7dd9b0d710
z889324c89c6b9319a210df3282b1845e86bc37e6fec4457c1facb43ae7ed7dd64465f57b61fee8
zebf5f27e4096abdd5399399625f8c66420f388d3452cbd9975a821a9821663d3eb4f35a40c5065
zc919eccf7e60eae632ebb739cf50f2791b7ac158ec1f737076927ec8f2f6a3846807cde75c82df
z1c873213269cb4c67b569c83fa4f46c04419c4d5c106194f31f24926c8a798ad9aff06e53c37b5
z1682e21c029d485ec24346957c10cda3e4f6171c9a6f5313038bc60ebead386821a655716cabb0
z7e359a5c9644c44216d8725711260c7878fe04e89e36c19156a47e8e8653729bd372820b644ace
z74dd1af96a3b1d91814647526268ae7e1c69a99b6ee2bca1a79bdef1c2c61155def3bdab4106d3
z30553ec4c7b7c67fe07accf50ccdbf468c2dd7214b488452e77e32d876222feda3bc657f0b6c58
zc420696716d6184a889bb5be29e4839ecb6110a1a466bb9e1033f862a36c9503155eaee9444ebf
z96c128d617e366c827b4611e0215e86121179f697aac76afc142889acff7089c33e36dbe061c78
z02b6cab5b9ea2de4e16e2b93427bb14990473b523efb2075a2367769c2b75feb134227c1c66176
z4eba939df68aef133036d27ebbb0975cf87929d4b79d967db52ea50adf3390f4bb1d4a3c4b3f0c
zcfe97ba4f5214829bd9c6ee9eb99a77d780bfadee7b4ebb23ee0d67942d2809c5255d8996a9d2f
z0d62b542b2c167f7d04c6b52d004e01f3fb1f9e9f4dad5c99de69fe4dafcc72fb6fa5ffe00d2ba
z04ea64f8988896d798ff11d9f0c762f300c81dc680363efa86d8c11c4505163a1de217b4358236
zc381e1819257a79df4a0bf4af453aa929ed3428b4478b2824b40b09b3bb12f35186f2ee4efbacd
z362bd8bbe6c2671b18252143b35c7c61175ffbb79995fb691df7697c671c8f07aede60235d1333
zb04924b16b420295215706cb250c33076f6ed416b85ff621a84a54ffe66cedd752f5b7c0327c9e
z8df2c11a3fd423ad9a6845fbcb6fb08f0a028488dc7cbc278c5428ba35d567b6112a28597b0695
zcecd5a50b609feb5424b383c6fe026d8424eb9bbc5bfcd1dfa800f53aa1ecff2bf11018253cc3a
z7d4cea73afc2215dcd8529044d4772969e983568aa26963116de3ee4eeac63b5629bc56455c6c4
z293fcbbff8e6fd97e4e6e7161446c1886cdf70dbe89daa95370dba28505529a0cf3fe3b94a7e36
z3bf0c2d8ab8fa101fb1e277791f84e6f85711662b1d7361d23bcbfbc1f6cca162010a380f26453
ze9a8a43ea2545459652b28cdf09e0d6ee5aeb971f1262aba161aed9fb3e8cd170e3d3e4f7113c6
z5a4073f9724afc5c655d65ca44a21d539c7fe0a8445c9b843024823ccdc86264753a4f060037ab
z7231386cf7af071ed7737d6ff59f1b86032d73d95c1900be14154b2d02ad4e4eb377990da1da96
z0f7ae853887c3ef037c1ec51b5c0a675e134857daea320897c7c29b888fd23ae3a68692aab5e00
zbe24ff3995c5ae7daef0e74613a1059e002fa0d71e3812ef35a3f55197d3b6e132cfe86c273d25
zbcbfe7dcd7486340fe34ccf1611c70a8ecc119e5d226dcb9eceb7b663c4c55c4889460f52250bf
z2edae55834a0bb652e5e5ac1be02fdc03416765f49a2f818bb0f2a61a7c04fd68c5971175ec3d9
z3f621bcd5252b70d628c2d3f63a618c31f04994a40e0581a5630f991059b96c109f1b2543d47ca
z44e8fb217d0c0f0faa45a8831f52f742330c6ce0981a1e0cf0c4060618ea07dc33bb971201b415
z9503c947b6c21bf41024377995feef8acafcc9b99c64bf0e89982edf2f8d434ae18f36fc5a78cd
z73311726a57ccf6f52a502dbdb1eccd12b2bcb73f2d621a40911ec595b38cc1c6b0a5b9f8ded5e
zd799cec9aab0c88b2062860025d6250f32758b5e958700b6778c1bf347e7ccd0c23efcb981ffff
zcb59c84510630660963af74d9846cebcec11075dccbb24e85d3b395eb4a70502963f5fbf1318a5
z4266a39b559ab2b780f433e72bfb7d6922e8b8c5595d850f57d243822d94c6f229766d2ebe436f
z37b058cdc49d92205ac0ec83f817bf8b1a296b98f3bfafc2bb2d73edf09bc78a910ade453a9b16
z005b47a8e7c1dedfd7e58749a1a28a5855e6447464d63469ae1dc8298b18c7eb10d6b6700a5f59
z03d6ed56954ab67b7f0e6a55de538a1992381be325205352e238f35011eb2443c5548139d99cf4
z8256ce71b4530a2dc9714422677089c3f32242df8a5ab5749179c73d6fce4a35c3e7b6e9b17076
z215a53e47984e6a12001d4bc66568c352d46397a70d854538384bf49a7cdf3854563947f4efe69
z55f0019389a63264b328fc56f10c15518e34509c398f00bfb10b8ec0970a3dc760d9110972cac5
z1b258b2a0f74af1ad921bae92fee13fbba8187cd2ed02e7884d975eef7a7da3a2d4b9924e87f41
z94845526be73ee4375727f12c2834640373cb13717dfed03b92a3f51688e9206a0dc82c52677b0
z3ce524061d9743e71e08ed9be333504449b8ab888b292808488bb6c34693382a7e679f4e70685e
zff8c9139decd26ee283448627cc7c0da9a9dea3eeeb01767c0b791cc3db63faf3d0bced390e345
z767399c59022e9508e22b0e4dbddf9caaa7494221b2a3371a1d03b2bd36e131b434639f303ab66
z4bf8383b04e9e81b576dc5fa40d91449e0197206d1770b6d99d476ce04ef070f32335cdd3711e2
z451380af2c8974d658d7f3761536a5a298b766d845931dd06828ff7c6073fb7580c6aa4d71ef8d
z7302ebfe57ca67ad44b1d785e0813a11f4399819d5b4602002529be5528e40977a640e8fcdb6b0
ze2ba51ea380ca325d8d8fb5deb1024d27bd2e6a3d29843b39423c779f336cb4c3d787411a0fa6a
z27f5c7e031e43b0329a2ecd7e07d574dd9185b464e12eb1e26ab4c1ca7ba895896f437c026712c
z8470d460769429b35fcf80ba90b9b3a70522708623daaf94e8ee92d7c16d4690f061936704ba99
z3c9d97557026173bb3da424626a726468af892e9d71bd0536d4a4f1780b78c8022812ebf76ef1a
z84d9ddcb0d3864b5047f5d5e55c1e8604896aa60ea3f579ac731d81be0c292c2cd88106a2a01a6
z604d002fa6e12f3b56d73c527a8263f1337f242f167454ba1e0ac3eaae633213dc4be4fac5dd76
z3f18ca546158c6c3f55ac3e479365f02152ffb649cb54dfb6dc2de3c3fc41e353fa2c2c6b41bb9
zaa39de0c25575a720da301a6caa4c8bfca0e17ab3d06c98a5a250d5298777e27f1a8dd4a3bf93f
z73f0ad00afe47b5c7459da4194488f7d4a65ba59c3b09861461ea895025a505bb079265919fb0e
z3546a3144861dea72a2588608aa3b4bb2412806f3e8c04fc672aa78051569b8e4a0b8a4eec1339
z7e6cd8790f173dcb143851dc16c6cac20d2f3d1e3572fee7ba5a348ad3cedfbb74dc892cdf14a5
z215a55fae726ee08df86422aabe5d7bccac30728708185c6945e3df4cc48415919dc3bfb5ad8ac
z260c024ed4b9325ca251f403e65df7f088f3232c29ad93963ed9df2900e9047e8c9f3b71382d70
z8c45152814b76cb34825636a99e3b3823a7380888d1a09d8c76662eaec03c1e4be0f90a239cc1f
z404abed559b9f942171827901590086df648ad336c3b7eaf6822e2307635be97ff150e4b2f043c
zb4b669e31ca0e675afb27c0f13b01490af69cf0329e31001b242d101eecfa0ef18a89169b29fea
z9ee4a2ddb0668382157de8f71aaa6dcdc9df85d8d1c06859e2effc48c0f454ccb71e209fa184b5
z6d7813296490ebd22838ef397ddcb040ae23c9aca19eadd4b697821e353a3921f3c1dac455e3b2
z6f474d7af5ee4d86f1fa94b9735937cb13b6ec9723c30791efe0f0b5b02cedef7e80494c446796
z37f9ec995e23d14c2763801cc732c59978a487efdb9f467587c21bfa897817dd4b96c65596de2b
z232a966c2443f89f6bc8a443773319eac3621912ec0661eac1e0db67afdf9c9b999309192a8c41
z0885923f62b073cdc21f89a050baab832e3a007854ac57b1fa278904c3e9d39abb71ed1c176a62
z6f21eb1dd1623b4ba4456bc165e50301d37a1f91bf7c4e293ebab4e6b17e46457df487c31ff0e4
z9c9be1e56b60bcd43f6d04658309b17a445a2db697640f69afe0dfc6ba4c36f1ec2c1540fbb8db
zdb674a4f29ebb0102eff8ab866912671331233653102e4c3f25bb3622e8abe1bdc39da008bb7c1
z9a429fca09251171d908e4318d1e85746ea2e631e21ea8c18e846e4f6f794e1c0aaaeb4d2640e9
z427be400455cfe4c5ac602ca5dc5b176c7e3f062f73f44dd33db74d8a53f641358de7b5333655b
z0f4c98a1bd728cfa71abc0cdda2de9d89be4e84f60611d455036390ca3307c64ed9a28a4aa2a64
z048df6f893bad9173a7b7114b7b68d12530360bfb1c455fb9d8d0fd21951ce45ab2487f5db53a4
ze6ebe8763fd65d40dde81a48ff5fc02c5a4bb7d1c0d05fb213898c213b4cbac9140d147e96f773
za67cc753f53089fa88e6fd94529916cb18c90a738db980cbf18360ee2dfd00b7e5c112d0328e71
za1f1a343b9955b65b2511d759a0f04e8e7843dbc50734c092083a316aad644fb9732fd2972bea5
za5bb1d28daa3f552c4360fbbf29daca75cf79a76550313a3188f8ac31c0134b4d937fbc7ff459d
z75c6311492b6710b2eac19d9d71390e12b1989a767f6b8aeb931971287e8a96cd5d6571e02b0ae
z370c66ddf52504973906001832122b38323220003876ceaaa4b88aa0fca20d093c89fc721d48c8
z63c84ba565bc4812600dc0bd839a844f4119da45391c6ff840cf53bfa729fed3eed853bb7e3d0b
z1af4a34fc7716dcb029d03b172d8ee1836736fb654801c729afdd2d717527a79e6c16fa362c292
zc838699bc51e489afce2b22fca60a33e9db59ab4658f07514806868f0b850b69cf414f5dace311
z597a6dfd287f6158bc2b57d9f1992fba832216da6b5150c549635da53a038126ed8445672c1243
z9ea5b2181933d13392c181fea2ecddcd18ac27d77cd37f3d212cbf7fb7be37c81ef7668faf50b6
z4d0c5af6f293586d4f819d5ad1a559c377a059c5e3a988d67e6caf3915fd759e72e9abd916fd84
z26fa434d42eae8aa58c8ef83b8592dcb84707c0bb4d75df25a77b5812cd5e0c3a17c5d42598657
zd466f7f1fbb5a19d084b060455de741a647ce71c884db63bc3dbb8f1a09d105ce5e0eaf327bb24
z88a3c42909a32bdb1ce889d2734aee1bfd093b8858114d3297f2bd4b30d9aae81c9def2f9bdf9d
z1bf5f559c08b8ea5bd32ffb14dd08e673bd5f04f02482d33c37a2ce9c80f3c60dd5d7976695753
zbcab3893d25256b12c109945a575de1e21d60a0535eceb05f9794278bf6b01d82ff3b02f79f19a
z4d3b0b96235ffbc9890d758481668c4afcb58c75c74adea9082e39549492eb784cd2fa3acd436f
zca89d6960435266abb38c038722f16c919dd02e6427c51e0d32815d9f05bff4ea69b8ac6f27dcc
z610e2682670c3ef04960b205b340700436d6bae420c7e6aa153892a7f835178f30e48a2839606f
z7be2657c094614d1fec0c64d25813026963b56d40c50899cb87389aa02b90def04ae397fadd616
z6d557c784c16c0ad7f83118c4a7a5926873adf71f98cbedaf6516ea8403db4c73d6494dae4b128
z1b3e3f0192a04d55b25cf5f7463190b686381a53bf460e576e706605120981e5732222e19347e7
zb60c020b2459ca73340ca3a6b5b52a1daa3f5c9147b988df77dc402f4f8e9d080697e222bca4e8
z7f569119175dec08965f5a0c9980bb09e9b4743b161d7eb1c9cee16e569cc1dcadc9a8b3abdb89
z977c180d084fc9d25d25ff1616d3312b8029d96d3880f8fa8a761b890ec7ac0638ee17ce0c7111
z458260172ec7ae00be9160c36beef375ec865f600e031c968784ce722718e680ea4e62424e4ff7
z4ed13022b1dfc34745cd52c92dd5ad57b18e204c499a381408248aaeb3f3abbee4d8bc76b839d0
z508647bf9970b58fd81722006318e1d24f730c6c88a895ebb76adacf6cb1706a9039b7027e07ed
z06bf97e57fa060824935b55920a8c089a6713b7b8ac24cb6a639e3a2c9156fc421e14e1ff1a530
zfef286beb2827c154d9d6efe1e7d76678d586cc8d915d606aaa2d5f72590a97622003c241c5d87
zd94076b208e7d8aa500484a0d7868a1e5d125c77c095a7e950128b40ce90a235c1fc76e76cd396
zd33ce7d4dbc86c5c7d32f42a1106d59374d202dc5e0c97b24ba4d4d4f09495cb9b3595c000b245
z63810e7b4a1ed7b16f56f93035083557ac113d56322821124a055f532a8fc77975ef648a6ade42
z11211c5412d17dcf78275f1a87fbcf1ac3aaef3551402ffc3733310ae861b631d322463c2929ce
za81787e810696503eff3fd6f7a83df74fba7552e0f7f5ad04ed23d346f3b01f0aaae7165cc58b8
z72cda85abcb79c0fadbeb4246738d946a5b863ead6b3dcc69b6a91c9933f4cd524fb56c9e15ac5
za1e21778387fc30a5ce8c203f3db5ebf19aff2057c56145ddb523a044d8512aed4049f84adb738
ze2af10f886fceaecb97032bf88a3aa81f0592dacb4c9ab9d707bd77f3ed2c79ccb8925749b6014
z58883100077132c8854a699ce4740b0e3237ac11c6382a5937489ed8112078098d5ca4b85377fd
z24878037afca9f639ab5efc6e2c1457868bf059cbb925afb4415a3e2ea3a73a4fe221ec90eec98
zd44ac33465c69faae86e5bd6e97fee2790c38742ce5a501b841444f42db5115d2945a8b5101987
za004e9762bc84edd0e603c5305ab3dff4a27fadc69870296f2bfab188cf8bce11ff281fda5682f
z6632875a6d2dca8e5c22181a40ddab27b0db78bfce31e3b974ad694abe6203223a3e0896432ff9
za8de56c4a79f365ef0cfea3e850fbbcf821790f439e85f688ab47afe4eb42a3c511cba4535af28
zd3a5275ab67a6029dee93b6c2817e0bcb50b39527dd9554960dc4602790c9fbe632bd7c9f3d9a3
z9278ee90d1b0fa106c37a8d3126f8e980d806e16ce52b69c2bc94adba8ff6e739ca04fa780e136
z2a5629019b46ff0f896b171d5ffb7a6e8b433e412d29cb074b3c5da9151dd4800792f52d1dccdc
z039d9cff4f07a6f0184c728c6e840944da5ac6f6eabb94c9226bd553370741986f1a82cd0c6aac
zdf2504135564a55bd54c84d5f827db83ccdadee2d2904882134430cfb5ab707e11edc5efb5b965
zb453f848f69c5b729adae866f785be7eda5a199f3a18c6ee567662e574ae7e15c3b32cbc0739e3
z939d5cecd3331c6534e1580a8b6268f3c4782c71070cf57f67136167368d0f37623ff9c3c85355
z6b03ae52c694dd237608aa6a7d75bfc1db813a0340cc314228525dac912812beff1d6ee79299fc
z1cf2ff5c71e8638f0d8f13c196e3dc9e2f4bc62dbea447b941b78144ba4165fe1ae7430edc14a4
z20d97bedbc718783afbecb716d3254541e62e8ff46e52209af5446e52dfdb80c543e772c00b549
zacae2e5f6972dd7959ad32baad65bb3364812065b3cb7e2acad6c2ec39b02d6ead2ea43560df36
z824fe42e10b96ab22c061c9fadee44a0243443d02dc42e4dc5bd1c48f88cf515c9e6b9f0c62156
zcc7209378a4c994fd6857994ac2e1b22d0b57659a1726d48ca7f75cc9a026733f7b52f0758a840
z8015834a12d09b137970203059685b2cf2f0b1e0504208bacec1a6f0728ee05b3ff03bfd05d1ce
z81ee00dc8c678bb27915982fc8232bbc203fb02be15a89ebc9043c902ec080e2e03bbeb1ae318f
zfd73f5d5fe1df51e7e1d259366e2baefc91287e278c2e3f6ce8ef25aacf666f95fff2520331e67
z639305cffd3750aa8526eb28f2c0363d3a82c572f5b64303d472e815992b13a38b56e3ce07d929
z3d990878754876e7b2fc62c5da6a2d99f5c2d818463d8801a5e097c0b77a57a3f8946348f30ede
z5713693720af6e2d0af787c330e69a2f7e809208d1d94ee17efa49d5b49482ce36e05078d74a34
zf4d64d9ec5cfc6bc0eee14fef45e2c071ba1abb7941b17c00e7d5b23fabf714269f61419267353
z2dd2e0b81bb192f535c123554feedcd3ae254699fc999db0c293e675e70c6f8e049932a4098baf
z7a4cf4bb505b67c6763cb0446417038f1ac700dc577cbde76b9919ae15175ef46e0aa511269eae
z47e2b313ef13444e79a207e3dfbd70d6f0bb1b267d82f5ed6a7cc4f0ccd52e3ec8a1619af3da70
z27260f741d5de033092c78296faae714a391f0ebff4f36a93fb16091015c2b096505e5ad5c873b
z1f4daf9d556ec198a31212dd15bfd86883bc9a12a5fc3e37db0e921e409680de0876bacc3fa579
zcc71f183314e86adafa354a4d323f5fc671a733728d46c9f8e8c2f31b928a5d95818ce3558aed3
zd44734b23350c619699ea02db63316d47852d62d4a031d0cd463a4d2c80fb70d73697e5c73ba79
z4a28ef77d4e6656ca4dd5ef596cc02b36215698fa47a47f708947a640bad80fca9a4bcd7e1a55f
z4295c1874bd7cccb45ad2438f8beb726dd6bbd0ca28f8a6da95ca645c3ccd06e499bb9d976124a
z16935cfef094471addc8b354003372ed3b264d254e77dc7d311e367dbd3607af16db03f3b67c1d
z18e1c1af63f1d72cba45f5adf1db6692ac4ca5af115121bb40d0156aa586388058bdbe48b12cbc
z388d2399227c4c89d2446d8539fda93b6f4d0ffa8d7a5f0a85c47b90f495c9e189b7279091b5f2
zea395abd1b7e0631bae0a0c7f720064b28d8a7b7e18243207a6d5e2549caa9899b281b816d6dd4
zcd10dc12f20c8f7b9e80008c5c90fd5a520b4d519a28daafb41032f785bcc77b38dd18ca88be2e
zfea437d88050eb1745f1a81bebb34c1051f97382c7842647038ecd6293e8bc085b46f5f972d2af
zce8633a23720e938d27b8be1dad6ae1e075e373a68c49a3aca01f619ed72c37e121d6b917876f6
z3db3d5048af4001982cee2223b361d6645aab5a50e02d64c774548f6c4e59737ed317849c96cde
z0ec26894eab58849b7574b1bdcb1bfaed48a59d303d7225ee373350fcfb2e1389b31c090de3d1a
zbf2d7483160576795ee61f74856f159c3bf7e7b81bac8e6da6c2aafeb5cc14d9ba6d315f63defb
z6f4bf16ba11a288b13bf6518ef6f7bf069d69aa7f46647e88e09193b8b11d10f34a7a14363ef04
z8e3dee70b5798dc06f33320f2f5429a61ee9f1cf53732f9dc7645d77b710b3df0f337da97fe451
z33f85493f0389e2812252adc4f238be0096888660d728f12dfe3ac3bb6fc1526e128573e642ba6
za90b8b9e5dbd4e37613c6c2415645c73427463759910029dd05c3db70e96e992096472f1582b2a
z66617d57c65f95b544c110fc91c95f71d83ff872a4ad2388a193467aa28c5ae08821a5fb90cb89
zb041f811839589e50b0c29459e00d5813d624d1b90b383b9287e09d18eee8375f26f9e1e14576a
z1ab288f6c39002b41e12babcca11ce58fdbcd711cf744645a63c79ca8479c06437fa689f6825f9
z3ef68ae1877767ca63394d7ebf7abab9e583a4caca9c649284556d1b04022af0e233f49f61a5f6
zd905bb3ce14ed032197579682db405833efc1d2913aab414eceebfdbe5dd58699cc8046a2c9303
z1f5b59a19b3f0a614b717e34cdb087f04a5494724bfff7b1d6ead4b4943429283d8f7569e70da7
z191ac62a4f73f5124d4a51a7c1f24f3eafa1deb0b0b6dfec4106a47b56628ba363be7cc62407e8
zc1d12ad1606d5a2219256e45ea1f528fc31050811605d3bf91221f918cb18a956e3c64f4864b5c
z0ba5a6c9114b6609320bba0d497e3d73b6d341e7cbcbd9944f2a48c7849c02f3b7ac6a1b2b187e
zcb5e7240941989ba9d62575048931244abc13f95a58dde449a5a3f1835e75d6873f5525dd7b875
z2a375cc2464a97b51695cfb6c6e2ef46bc55ae9c0467731b65a6659f8b04b61e707087cd01bba3
z6137ea35cbae77d6ece3949821dd2e450e83985bb35ec48801edfaaaae18d60dd5cd3d81f23c78
z2b14b628ad472d2bccdf83d951890d890c519be67913806f6c4ad575b516a3daf36bfb2ed5b031
zbb376c5f13fb97b225d60c4bde1b2781fe5bec808298ae9125ad31bd52315db74fb8b10caec2e6
zd973b3e96f69f57208b4171feb8d2dd7d4ea1478585cdaa073b9ea501051f84bb4b8087628e5e7
zee563a5160845c8fa23e44b683fb45f0fc9b2d2a224c12ce39cd78ce7bd375693f33b43579cc12
zc0bb48150d1182ce4095b7ee6ae496ab60e32106a002beb83cb62cc284a1e92b0ee0cfcffd4163
z0ec621f9c089ed97af7f23b0c0a34fbcec0ea5317f2a22c5b95f7ca40fae9fb8e2236664fd322c
z44c41df0aed2bffb3554806f6ed814c8c3645eb3f95ed53fe81fb0d53c0ca822cf833ce0a3fbd8
z7ed686c250dd0cbbbadd5a59862a6f4a78f4c0249da685e2d3aa04250aadfca5e2a3e624bb59c3
z65f7e2da16c728411a0050de0d1986d4eb980036b7b8e9364f5b4664ff0965b176669331e3ac73
zd80faad1609dc3c0cc4970dd95a2048094c72abf70fefd36f8bd5696d1a006f15c8dde8f7740fe
zbe066c6bdb667559655939f53dc0065e882c9e7bd8caf0bf268f458911c2a1a84f5e56ec44a9d1
z6443a57e1be7789947661be53f97c9f5eb0d1ab70f41b5c71a19296f1199475d73e19f4fc3a210
zc1580e99c5a25679519ad2c61550704810b5694874ca70761708483d4175565da193a789e9f2d2
zd7757cfeb02f8047e11e74e6de616d685258b4b9c3f9645f6cd91971eceb6283e2146273f78814
z9a822901f3b9ba28adc7b2354b0eb0723d8fdb2796e883cebc5a9984ec7eed3bae43be821e601d
z9b3c6cdf5462477fd07de494e6e3a4a011acf1886cc59cd0eb908e5c91879992ff24defb3b39c8
z10665053cca84e0445e4a3a171e187d37df6839e4ec1060f122d73631d66118e2084386493305c
zb80525f7c4c1c99948d80311fd38aa8883ab503ab0af8fe99da5a07849b272e6142c2e22fc40f3
zbf55ae64109f966cd94290c1616c52230fad47cbfe2fc788f38477b7efcbe46648efa7e24ad4d9
z9144142af1c48e21a802cb91710afbddc4b9dedd422d35ef9b4b7932d71f9ebd92b3be545d27bc
zee32fe87f03380a2f5bf13461a2fdcf601ed4f1459343cb2ba78cce5b8ebc948cb433e7812fa88
z6e33f1270c378a6062b0ca046c4a2efb365c37ef07d17ca5249344ff8fb0ee69c1e8f4dda079df
z7771b33a175329b34e331f7ad679516fca59928c34628f7ec76c0e48869536ca657aac8ba50123
z76a1ad9b000da5680c70e47bef3ccdd1a1eccc5e32b8ced80e9815621c83a02152980aeaaa7db5
zdda07a12e2b29ac47b248f9e29d050a68a010c060b40fdd4b1b8312948559c2eec0df23f209dcd
z25a6ee49d57a96e0d88f07ec944d2aa6336ff661f3e55bf41b625d439aec4678b24b1ab813089a
z10dcca95d460bc78bf74c0390c2c06ca8f5f5c544b8817a09aa291372b20ceb033fe301d82d626
z1d353ecb356055666d6a4ddd1a4c0483d9e9ff95c1a218abc9df2b298613ed8fe537d65c43885f
z792572dd451097ba5120e9c5387d272090e909488a00409c9378b0a465d7a01c8edc9e17054e21
z31adf11a3d436f5fe066dc30e108ffa33dafba936d22f8f97a69d524717655c901c534dad41eea
zb93c91f6fbe22b84add547c53943dde6a39c861d3b1cee7c995d62d5ddf2acf3ceff5a6957e0db
zcd28c286fbb72bc346c3979f617ad18250779c907c6f7abb1197aebe617a2553cea76c77d01ab8
z3554252b2db1e4ce6f3e39b11775d970ea6942b3723ce4515eee16d0b79834bd0b6ffcf1a1372e
zca8d620cda8aa66c9f7c43a0e3282738286272586f06ab3d69ba833d7aa92127ddb4da18a46071
zbc4b2d0eb5776a856a0d45c39f7eec40f38f6765e56d9a3c44d82bd7d81e149c0d90155ef994e9
z26373f4e79d7ea8e1ecf737db133e052a7665e518f79b2ea7e3b6b8fb64aa70099fe98ced4eaee
z64327ea223587ca0ce445828a5bff963ccc9e68fe4079f0227f774bd3b0404b7326cc9d1daa782
z0cee798df5b5f2965db76dca1de69087dbcfc97fa125532eb26e08d4b2befa9a09c1b5821bcf5a
zde8af8e43a1028d7cee03a00a5a891277cc93c2d0223d23a05b906b7689b4b4937fc894d842af0
z184e9a293409830ce2fdf85139cdca8d8e4131b23d823ed42fd675fd6ee01505937598ab4dd438
zce8981bac9ea2b2b5e3d4cf42f0c483e0f1d8f5e21a367f5219b8ff4280be81deae50a920537d8
z74afedf870a01547a8de95e5d579777be3c0567b569427515e1a8024f34eee246f99402f4a4f07
z4e8d1cea1289a041b579052c9617906db593059a152e34469a2ec4783cef7453a8c782a4706029
z01eae1eca7a654359b54d469b31380de96ff14876471c0b3cc3e4516fee22f3eff4b011cbd28b7
z513258cf2d54622551e65fc8aa5778086e2c62d16003d3ef465c8a1b3ebbf6a4cc821d235748a1
ze64555656a146c3455b00c04d7da09f39da450cd70d42fe11d0a0d1c1bdfe2b97dea04a369e6ef
zf42f2136ccf267b32689205c7785e9ffe239ac4b8fed8bb94fb9181e7480089e964e9dc730f6db
zc98720b3900e3ed1057894e627ba0a818a3a92c5f03abf712a185606daadf9ff544b6017b17a40
z97642152ef627a67e78abbbff9f1f00b5942c4377ee4f4b8298e94c9d39a0c08739da2bc1179a5
zac016b5afc3b139225b8688d27c6d072b94a06c450f36416795dde07aae547ae2bc4d87d8d951d
zde40f548bfb10841344bf91e82d1e59149256b734edc30c195d5f4d60cf60b07272c8e2d026740
zddfd749251fc087bac6b385009f761ed2914f3c2ad13b125feda4232d59c14a9a1b0d9c0beea66
zfa2d508ce9011f3201c21cbf81dfe626e3f01a50decd4ebfc4ca6ff2f4c55a3bd408324ced7d1b
z1298b76f25163acacf55ffe23782504446cbc328d72af56753c773f209ecf87db5296fd0b37ecc
zc5cc8499d0a979fa351ad0df51edc5d43c1aecfd14afa84d1f3e46af631054f0277b57bfcf4ed0
z0f73d560871b056dd34f9ba7f11e8ea411355deafad759deb4873dfcf3539cf7df3f383d2715b5
z85974ab6cf7ff31678e197ff353a49fa8fd203d81f3a53a403ee2e7d4f75d16c9ccfb6b7671015
z7b7b15e3087179eda6caafeeb22c745f1d345c5d800209168c09a93848b7fc43bbea117766eaa5
za5d29ba36217c4c31abd766d28a9b893961c69c463144a9dc5d77f2d40c1c500fa31b779a8b82c
zf84e178285061b88214d3b4972a02e9738436b1b716304111712ca50c3b271e72efa66d80c2997
z89be54c48b238f76cec02082bbc37326894e6c11bc0db948127f6f6abe7b8be3e76f1716f4372c
z17c2b9c10b47e53eb88d6801dfa87e86173eb810dc5904f6dd29b4d1363799204e01ded95084cb
zee6ac9f6ba53163229df0f704285c4568e4695baa52c3ebb50f112c15dafa4357fb82205eb20fb
z403f86006a2b7c984467d918714536924c58652bf04287cdb1320ed0bc6ceb747092cab26cd64b
z7db8f1e2e3ea9ef6de71752dd7530dc1e4c6a845cbec4b23064f2e26ad8108128f446731e67c61
ze9a095b8a3ac3eddcaf0f2e4c93458d9d1846ea4b52d2dee23486a6dde6b68ad0aa31be918771a
z161f7a53c7ef02e130f26050772efe0169d512e394c2f7414dc29caf29a56bf5e45604be9bd311
z8d506b3d5b044e9e20604805167c8b6350208176de303e314a9f00de9e206d82ce9cef97ca05b2
zaa4fd882ed40e39394f97812fd635971cfba2c5306cc2e8dbbbf7af7c5274c30dd68a96098dad3
z0113ff0a3db2c415747967f54181b6ca93fa1c42fc63b5c9492de9012c95a61d50e702c9b36230
zc182054bc39b12569375f317ee33afec4a35ccc058da9e677cbc190295b28c403eaa50372eaed4
zeaab82a12c80cf20209139a7eeabcb52f347cd419241d7035d5a7a0f4ac4c9558ac73952abd2b0
zf7db915b80964b5be918a56b454985abba7e1fbe92875a15b023914fd15b949e304ce49659f68c
z5675d0bdac7b4155cfa7dfe890e7dea7f2d6a01fd9b0cc9874ca049994b4ce5098134bb079cdde
zd85844f3effb186f0f549024b113f69792a0b8b1b4d1cab7c9171c3632fe84e192b59f11666fd0
z0fb5ed7c7dd972076e260c0819f585157b6b8e0f22059287aba6f86a7261d8b579cd5740ffe53d
zd96671813fc2a37f575bfd583af6deb34f1f819b373b8d2b17a36cb35ea8d7282617a7a0673c58
zcd967d0093d2139f19d52abc8bfcf49a0a0276e3b65e0b34acee427ecdbecb757d492660696ae1
zf4ea27e5aa667698f453746466bc0174a8520cc4f9524692c667deff193e792de0686e9d6cae74
zaad6062094070b0b1995dcf71199b6ccfce56ec7765cf5bba3e4004ee789395836b41c620d196a
z93744ecb4a20f3203acb20ac144985e10cf207623e770052e7fe50776b61f3561649f482ee4967
z1d8456ea567f82c115bdcbe3e570f5a9b340afe9dccaef6752c6237f34179e9c425168bbabeeab
zce8ac06bc27807cc9c24d084953065285a0ece3da56ea2bea4312d0bb4bfe8f7d882a5a95f520d
z90fd064a1bba0c5cf5c0ab53b8fdd98629f7a617365a006f6aebce1effbba8ba8833144710ee5c
z8f5341f4a36bee622e7b6417ec40141dced91399e46dad4e2cfdb84e3ef192a47a329e73bdcfae
z0c118b514f1eaa4d1c7a2ee3613dcec5393d826ca4c3dafb7f0d04832875c9d0fb5ed052555373
z3dec4134e9f20bf4d0e1a6f2e70de92bd5246c555dde8d793d3b73d420517bad3103c648c25386
zd265d5d3e6279906bc1e661696cde0e42eba7912856802146c98bfc5957a1bc9bc75d04e0aedd9
zcf2c57a988280ec5932ad7efe1e2df90b08689d686cd3e8d88a549203b5714ec1261bc7f4954e4
z9d6784d246bf3081706b3ef7bb6d0b2115b298852b8932e44146c5e01270384a3611a17dcd002e
z6f1149ae4b2bb2e053df622828e3e621f2eefc82219ea310252f5d9a2e452f82c889345ee99cb7
z94d9d59762848d320a2172a41507151bfd0be49e19ad3f596d36e694288a4b59e57e0872fb18a6
z852dfa0211e81b716c943109cee0d861bd773d33f8c754f4ee17b1dd401a3578b2c626d67749b7
z11f5da6f1159464580266fcdbfcf4fd30e23d9dadbb1d78f761db5f220b032934d1ba1da45e0af
z0f1e8f156ed1fcd228101df322a6f4e6d25d33fb7b8e7964d48cfaf360886c21673bcf9b42e1ad
z6898a66f4a1c45766b99a7caba4ce1b9c9f55f88cbc05a2666aea0f9133f1ee0914eda6a63e782
z8905d139f6b34b37950c38c8129663bee3379be01de99d25d41a033f9bcb4bcc9e67d5b276197e
z5af040ba44dfe494e98392aa523add789e60f2b5c947c40c814fde2452f1a3237917e6718f019b
zbe31ef1d437f2134f77314e4c92f6a0134665eeb03a2baf9375b0c73b774d5cc814a538fe1458a
zd14196577b4a75a02969944c1a5007d373bb78e5968161c0cf043d40eaf94a65c54d24b8a8bc52
zcda24a4986d93342af62282e04c166bcf9376ffbe2222b900b9b6428f3e21aeb9201d993ce0e2e
z4f7a5a0fe2b9998059f763c054abe2969a5769939dcd49f5dee91dc4426c1c6c6188b59c133ce3
z808b53158a2936d02b5324c5724059016a778dccec36fc0932e05a91f7aa624fb9598a832aa6ea
z392dbf23bd71605b01624d5dc4a74602a3acabedd73050c42dc8a490bbcffe65c21aa58750077f
zc05805490bb9adaf355c04de3baba96aaab6891bec195a732b7d0ee38f954fb0d05d571e559d4d
zb7b565a534bc1ae5ac2219bfad7cf00d0b31e77c6488ffdb9ee43d567e1f6d26ff6d355a2e394a
zb32e4df1a1f93b90db3a0eff3327107ad9d7551c414bafc54e2ce6c4097f67fe438dae62f0232f
zc9bc5cccb374d1eb36e3c77cbdbdd8662b97b2fd44b7dcdb6825002c2315274864412b084e8b3c
z913c7ccb2d7f93af1add70a9e6bfa95b709e7f6f6dd421b5fff42f83081d94340c4c1c1dfef76c
z5176563c9150b555e9b36e26d0b566eed93bd1ff97075ec317a23095572c5b767cc2b2ad2ab5e5
z5e81c21df89ab402644dac552a9d4f5e592786dbc1a4a95ace42164c9e08c3d18d43e09f096b99
z53f7504197dc8a4e7fd4286da0d039fee01fd1e1285b142108f8be0506e771dbd0019c23574b8f
z603356926207ef07f4eb49f6e7ae2c14dc20e39f396c87874253f4fe2f6331094cbd7ec4ffa9c5
zdbfc02a6c1ebd134b8bdad0e97426c4f4f33ce7e0357dfc1d7346d663bf4fb981e5c9fb00d809d
z3e13abf5d20b072a7d50571005514c1ad7f4e2d2224a652d894cc361ad0bc4d0987e41d7b9bbc4
z5a733c85a8abefcc696fb0b3c2e8da68c4f91aa509a9fd76da8b8c7810023a39fa258a6947aa8e
za5d5207c22fa3da11ecb2abca9617fe03db065a260fe90a352ebafcb9cbfabcff3eee1184bc424
z3ffb55ad862c610e3725de0b000df295bb68bd846392b4670098ca5c025e7ce9a051a17b90dfb0
z223f870cef90f58bfd475f16b2f14e56138d75a4d77462f6d63be455751faef89653f445081754
zbe233fa862aba0e6a272e8f0c5fc51f8eb8ec0bb0c8926dc49addeb7f0fad8aaaf4a4c6dc58bb1
z4f1e7340197c040471e262284c542645d9b289097a895023a45a51dd151badb34ada388f33c9fa
z56b15fcf648123587d3d02e48d623d309281eae27da6879b0cf68d34672948812b6414685818b0
z07d83e8df942de87e5cb48b78d8fcb2c112c13a846359b8efd26837899189ae4d372ecda15bbc4
zf1929ff0ce7f3481e8d504c69b2001743b8013d864beb14c7ac38c2df060d305502b80ad50d57b
z94c4c77843461706fb2b293b64b8f4c220d880a6b83777083d8cca21f86e33c17f72b6bc8f796f
z4425e262503852c3584eb4323a0fdb06507338325660dea8f1edf630a9f2a77ea547e03daac428
zcb5519faf6df5cd79850a5d600d0443aa9f4a497928f93c2c8f1ab19fcb84fd8315f437bc9fbbb
z131655fe5301c1409179d9456ec40f179332b92a28b6826304301c8b2aaccce9323b390c6eea4a
zd18709ef0bea24a180f5f80d1c258db5f047c0e3009c985e2af113e402415722db57cb27c33120
z38fcb94382746478ad22c4512c20e02b959cc50b3703d7f3405943ffea4cab9f2a1303d5184d9b
zddfd58ed0e70f03c1774d94165868b82b8902997ce9d5cdcedcd5a4541772e62b239930abc651d
z85a51802ff11c6ba679e2ec1fa10b2946b425de3b3863a555b8af192d153fc5365e29ca130963f
z6ce85128a7afa0b0545f050b1014816177bb35b037755bd374f122583ea6da29ce0dd7106430a2
z96b467edfffbde8a091201817633a26f600e53f2b9981c406bc288e24d9a8b2a7c21e701819ad7
zfb113ff8cbcc1b6f26fb5ac3e59c99a849652b11d15f60c498395620eccc5ed8bd76ee326804d1
z5707a1c90ff65f4ae546bf3f658f2858db1c8955b0b2a2fe25eb219c900833761e3c75ba65c597
z4ac380c32c7872faf1a2ec02cfd5c17bb572147929f04b4b277f21ba07157c2dd46b70852ba199
za059834e84b2c591fda71ed2e4327a8246977a44274c6d5b04c79a9014b9358b92ed1ac75a2031
z97fdcf4cd6430a9bd1bab5234c7b80b6f29c49877c3c0c8250eb334de0a041609c61d57d898f4d
z2c631f47439412e777ffb1d5e4487c12cf49716a720adf3a827bcaba3bca4158d9eb8c6a2434f3
zfeb7bbd556b6617a329bdf253872a02a4c15d86a111cbc7a1391ba1552f4c1c4d7479b4626d2c7
z36ad11595dbada8eb7e959f1b8657f15f2aad64f4b99d2dcc2b73b5d30963cd6bfd577b0c53d25
z030cacfde0f7f2e8f74b87210e949211191bfeb92a6f575e37478b3ece340a39dba31628d4012d
z73453d244412c787a737d37d17f20af0f51b5c419372891492c98ee7f6d066a78c57c677e575f8
zd8f059955c8cdc3f5fc80736fe1d21a1b71b6ab2241359f0c5a9a6245c1794d3218c1e3c28ae5b
z85130df9d01abae28908f48d868ff31142cfddebd206389ac6c3624cd877acaaa14dd0f3bba0ab
z14eeaf77d89827bcafc56cc51d96a0f21cbba62cda1ece55ce8b7eee2a5af65ef6c2a12cf33674
zcee3fa802be901ff3b48c5eb38a4ef80dd325bc88c1c94cdd9b937b27203498ee648e0a6ac0282
zf3fd406b8ac6b6692e246017957bdae749392120a673a5ceec0fe4914fcce7c4b8bcb7e0323337
z5e6286265a2be57f5aa8eaf8523b6653907bd69f36354fa8831085f9a044825d7aac27b25585c4
z690c677e9eb5a9e0bc6a647aa5805b0978e7eee6867e4dadae84be6105847ad379fd355bb78bbd
z1fbdd6cc4db0c6832c8824d0148df858e0c2b48d374120c1be0ca237a28a0fe8ffd2fcff800e64
z27d42fafab91f077b2a0903bc115bb84a5c27f0adf5874dd9db42ffbb9ec92ed8d80ee9e25035d
z1911ca0666248e1bacfed363e828d835596bce67b6ec35e8319f9bb0d1d1fdeb62b2921fba9c7d
z66ccff562ce3962b302c56535f80d70a45870b8fcfeadaa34c7e1bfc0cadf3534881458a3a9424
z93c8bca39a578c3215a1f7b57f47069219e83916cb6196ad4e56c73f6b75e9d47ad077f892585a
z776bb395e9e78532ab140412058edfa1bbe8fa33e38ed24b7468f8fc4ae8a280b786ee6d250944
z0c7bd609501f4596806ed89010acd59301f584fc6151b86dd357e8ab3bb7943c279bf7927e9c6d
zd1c74d6bc2f051e1245bda01986c5400e2abc3b71d238e12d2fc934ae9e2df6262d008e299e5ae
z84681189a3a99199567a6a37cd34f5473001fa67ea4428561f509f7ee56a257289ec884fab0a5e
z037f3b77b4b6cadc3b18b1eefdf3493c436789c2bb421ffdf872e351364b0b8766bb29a58280b4
zef614f3cce8784762ade431db1e7404da0565c190eb0fa801944fe690d3bf18fb26480709b6bad
zc416c3e70ea47eba33dcfb4b4bdaa50a639119640724ff82b1cbb9fb3f97aa538cec6035740f8e
zaa0cc74d79681bb0b2027e5952118d60c17dda6c9beb7b419dd465f7e4e21749d1f9b348dfe752
z6668ab9967877e7f1ed6c7745e27119f6f1e640596c160655f93cf7163451505dd3804591114f6
zf8ac6a8748e8fdedfff6f54359fd91a6fa171d08e7b98ad6be04708767154fdcefd88bfb5ee812
z1e29d593d546c9fc0720c5811f926164e0ca264ab080a91af9330a18e19bcf42032308a1ca11cb
z36ef5ad7374ec043482904aeb5da2cb0b751215b4f5bb78f427fc0e06daae6c456fe55f859b7ce
za383260428b2ebbe825b654b9f45cb585f179a28ab37d8aeaa37512308849e24cd8e25d4380e17
z40f6c820f975caaab642d979d5cbd7ede81625d5c635a84b65bd9e1ab4112b10c023c9513a3870
z46cf5debc8a0edaa0d96c2ef7f832536faf2e11bdccd7e8c8ec751a9306ebc7a7b2405c8b4adca
z4f4b06d505a748b27c69ddb6a40f9c44e5ec11b77a8c50e93fcee6b1df6cbde3e4f810bae882f5
za43cd4d0e8951c92186dea4a3b42874d8a6487b79845442d56f239271e6ecc8c52a33db6045e79
z221bacd92b42b3f0360944356a9c734a6408fde2796affa0803ecb19b8a8e3c42b615317f685f6
z2562c95a40a9608ef242af92f95213f26d9885c2b35ec1d6482463f6ef89c8331ad6516acd21b8
z0ad8c5b6015340ab30deec7c466529cc797a78dbeba2e17c7a3fe7078c0ce784676ca9a8490d4b
z681d55c85fcc14ea3e1459096a9acd4ea482033455dfa7c442a97982ffb95770359745079c5379
z3c48d554a3179d0fcb8902700a1e2a4d259d7c8f0dbb5b8f716e4c91f345f9db0758afceedace7
z7f5d56b4bb9805f442e6eacc44d70dc353b6902418602d301c51e23bc69cb3aaecd74765c196f9
zc4790b56dc139239625d7c88a0561e8ede5c65754dc5edbece1df1d4a00caa92ae79d205f64769
zeabd735c1f4ac984679da41ceada0e054b71624c4ffc53030b0f9d581548134cd7369beb7454e0
z5036a6d3ec2d551cb0bb98eb35d39fc3e6e94324e5975c0d7f8d9d1e4914a838948fa47c90e8ea
z416e7c5d1c6e1387bcb9dafef5cd98b135a4ae34af00cd1a2ef8da3bc094bba381c83f04c4cfa8
z8707417174789c3fdda3e04e9a62ef976af01e10c583b067a98584e4d57e03b1eca4ddacc08f2f
z09eaffd39ccdc97658f5f54a6f753af37268bb68755c203462a8bf67799f5faae4d055e39ea7af
z6b055d8d00f0ac5bca1efb96b69517eda48b9f9e24421edefd3d06083231c9579956cfae12ce5f
z39e98ba63698d369a62a7a98b6162d67064f1f9e1e0a80cb4354dab5d22678cb90f0b75c2fa0e9
zaaa591a7f07bafc2b3029b5861b8565dec38a6bf4af1845c021daf0230e178565a59d858614109
z41ceec2cfead59f4ebfeb0959610e38bfedf59362b5da914e89dc8ebb2b0654ca8fe87aa779913
z7c35bb7665f308deeaad67128f0f07feeb32cb068b1c5a5caa4761f301248973598d887f6211af
z19cea2ffa331393e5b76e2cf3090037cd8ae220658cb6d6793356bceba2134c45a2b2a1e19e90e
z6f723696e4345b218f68c6792c78208a880b23912dd6734c2698e49f6f924b4849b46186911037
z0c8bb993057e864994479e5eb94bfd3d6674c224a99d4e9b5eecbc7f212b6f5ec8cf18beb5162c
zadbb727fdde61d937be2c006bf1a87febcd2358763e9bd0d1cfa4afb0fb6c464093807fb54329b
zbaf22ab6f0642b76cbc17cfea789c325d79cae15adae0c642b665f6b8e4306079111c012845769
z9b606669f2903a4bd5139cb95e8e25c068af679ef7e6b63aef9e99c867ee259373dc6fe0ba452a
zb134b6071f0123f573b54c7e143adf820aacc6b2faedca80679ddedabef165a4b454bb078ac12a
z55b3808eff8d4b01164ee54672314b6fb69f07a669cc3531c6e40db24f89bcd37d8f62f148aa44
z1ed81faf74b3741ca02052b00b05564bb4c4e99b2e6d91c3b519b3b69a71dca419f9bbfeadcea3
z20528c588b4a8a3030d79a9325d2598b24b031463b2219a5b90d5357e9d7b4a11fb7b9406d0600
z87710f2d4105bf2158c1eb8da339eadfb7360610f7544750e8b292b07cb3638617cd56b7910d75
z63fd970978fdc7b6eb755bc825e43a4135ce5db3a892bdca2cc76b42c840d1f7a1f892ec8777e3
z3b21191c085cfc9e993be67c79b4b75f93f411acf47d4b5d32b4a4d5752ca307f0e4a6165f9bff
zedace2f47088a3a890afa57c1e9418e40a5aba4463ddc148fd27b4fed094916ba60101ec5f5f52
z670c3cad33b1ed3180cfa78739792ddbf24b839e711539c550cf8b4dbde44af953b53a86345d2f
z80c461210196741ff8ca6548baa26a7c0605ec414b58bfce5421e74bedc11a109ef78ef50c163d
z4dd5a67b15a7531f83588d2e213f3d619d55c11ca7494f9a321de6514a32efdbd020692cf9a959
z28373d0d60de90d4757658375a96837fbf4ea4d4c0f214d0c414b4cbccfc42bf9d6f2b83533c95
ze68921dd4e225a89705fee9ff36a4dd77fe2bbfb1c4d91f70bfa461ee9234a083cb2fb3b9de737
z81800b35e7d00f64d9c12d44551f0665ac20d5274f6cb8e168ae22c59aa435d23bcbc2e397ca25
z80aa16ff89babd5ec927318ff844fdc049c6430dbc838c947eff6904764afd9727f9067ffa28e1
z3e68a39e4fb54c0f9571f92e793ce67e2a19dd4a4acef9088c10137523bdc133149e85b50b1db9
zccbb23ba3544392e0aab74f1712822c5e2b6465f1be05c607c2e03a3258cf75ddec5cd3747623c
z5f96104a3f30e2a3904881765cc249727ed44c1fe248b2f9644da163d699a108bb172b90c9d26e
zdcfd8f0f2059273670ac7b510a341dfb98440077ec05a634d1451597951a09cf8d9e7b1f3eb46b
zc45cbf787b9eb13ec14039fd18d9409f2e5067c9615419c609fd36d8973ec2351960ff515ab172
z064693968915187290f3d0b241873c1f6baecd92e61dccd7ff51580cf6478fd19a3e7cd7c5715b
zb7a4737695ffd59c3f8341f38ef8508cc76fcc2914cf838d886ea0475e30f51f2f81b53d27a3c5
zd68c4c5ee650952f5f823762eafdc6ac49b5b658ec2e7bf14aee7fc3b5d79b0d3b612184def58d
z32dc82036dc522de929b331771d74ecea5a8cb836fb75bceafad96363491181bd9393f11b26d04
z0be33dd227666dbff2075ca58349d3834b74d70294b9a98d8c534d8b5943b7adf7a45d773fe1af
z115b2f52c5eb3f647e4f1f0ff89a1142eeba7a17d0bdb341665cf375e4b836fbc842ad5c836178
z38fac4263085b50f490b1f621291575f677d9f4f2a3934698a4d52b603125d7a411e6a381a5b5e
z147bf6bc680b5d7958668f36723f5dd6e4b34217ce85ce6725b3048aabe9c6731b617cb7292c3a
zcf1ccfe60f683ef069ca1867cde8a57de4b285a70731dde1da130f9f1fcd70089bdfae3d379a04
z80097e60a14489291040344b838e7e60a277eeddeade4c4beedcac66b1a1519bcdf734bcc7692e
zb36efae1307cb954b8d999e631c30bcba0df575b71459181fe3c0840176e2e70d892b4913365ab
z0ccfb5afd1be0d797cf5c8e48c0ae91eae57d8fd8d66d3b576bb515f8c7da397d54e761f04f936
zae66b76a754cc78b671fcf7db2d3eed8f148b446807f85d1b8cc997710c90a2bc1cc163b880ad1
zb51a6233e5e76e75afeda34a402b149dce1673e8f474b6ea55dc907554921cb2fefdadc0aaf53a
zdd015582d83e4447ca89c28dee8a76d0d3154e64cd794da875c5fe8d12eb1aeb4e41eff39f4144
zbb9f6dbca9ed3d3dba8c6f8420dc316ebfd206c45e222762e4d88bd855d2ae6b856c0a8f582a54
z414679108996afa68a113a403b396528f4964a3c672bcb5db809f0db409515ac2db91e7c26f501
za95bfc753587c148dc4bfb825dc74057d213649572cb9893e6ee4883b546020b9a8fca2d7abe4a
z114b40fb3a7341ad874c750e55f8115d3b82e33ccd8cad03a66aca8ddadfa3b9a099ddf4014a3d
z22f12fd81d48aff720c2d3261868448761ba0ab81c5882d229f62c99d355d602ffe253b64d5cc2
z7aae04648cea5ef9aac55860374079f97e5589f4bad8af1d518909d5040348163e9dd015dca6e8
zd9a1a456c4b653fe8713b88fbf0d2cac32c8bea1f30a9f40ceafab825532aef6dee0bf6a8673da
za275f39408947366816829c41432d2bc9a5dd57e1bf98847038cec1db904ea9b470dd9bc07c7bc
zfe5fd1123f79657a42dee57a6dff39e5d3f42b1b7df1a9dc7d3c6a654a3ff3010fa2c9664f627c
z228a800b96b425a4a04f91b60f7e604017f7b05478c5ccf9bbc98396649410cfab99eb5ea5174d
ze040a3d6bb3d509256088be8b47e94fd5e150960e423f95bcaf792624039c5ae2719c0dc7112d0
z471a56f7361f9f83f0178f057aa1b0ea70624c2b00dc358a2c26005ac9fe3bc19d1dcc0a5fb2e9
ze84c54dbc2e726c398abbaeafafbc8c0b4f93a8dbe21d725cab63999074a5abe428415ade76ab0
z3fe08a8d28b674de5a7b27f0c41f7f0ff6baf40a9a36250783812bfa8d9e00b39ee81a32512c38
z3bb0f96cb640a98e9d8590a4107c6e58469a0790bb129a906d716565132ddd5d62280fd9c6726c
z87ce78eb0a831679b75ed7fe2141a4aa0f909bfa8e049f0fbd8f4de0ad04b8d74291dbc6432d0d
z7b16ef96e68d06072383adfe08c34c6e4a75f28146fc70d4241ab73b21cf6f13b3fdc560b51b5d
z322d9d6109d661865a7fa4a78c15484f7518c9ef6fa850efa387fecf3b2b0c7228de27a1875064
zce9aedd60d1229757e036f6deedb5636d3b37f499adb8dcfd844b82739a677177bc4633fb7bb50
z9864532cea2d99031cdea3d7c99f69243cb7fca70fb91ff4bd4e082a01e3ae68432695be689082
ze63c1dad020c126f04ae2531a747532e8d3b9f99b47a86b04b7271723591751dbc372142dca46d
z7d0dce1ca362266b0ca4fbaea74a84bb0284415004788e94aeffdf9973bc7f9b64ab44cf2e45f6
zcaf7687f738c163de172c512aff104d47d425110e980e1c8d11d4fb283f3335f0009ed5ee5e31e
za4889903c09fea12d7c5e80966d0008bf8f4b594fa18f925b5ce8a28361ca2fbb060c1ff68337f
z2aa514d9b19fa01c91058a8b60cf038bcca5050196ac2fbddacdd7246ec78caa11168c08c361fa
za6724c6bf55fa173fa1223ff2fa5174554ef38e3ddb133d843f7c37917ea9383aa9c2592a7202b
z4b34041591eb38931c90bcf155cf7c3dbcfdd9a5f0a7d46612b38f60a05da4a952d869239dd9f4
zcfd04bbfdd95d23ea480d8cf4c10205738dd52d008a696679a9850fa037bbc21ca517ba4913f24
z1f047998a765320238f8745779d5dd9e216b18a26fb61adb9d7dc0f478b51c253d19097cae3979
z78c7d98732800a021065a67ef7e86be7cb0cd094b305eaae011d3ee4888e93f2d36a533a49005f
za0aacff1f2024a839f2a767b09a9f071b880e34a84ebca3db507a426c1c56a33c390fd94cfeea0
z3f7545ec704d9d09e67a950712d03f5a7884044cfbf87813fb3283e0806b796e0ecb67b5a47c22
z82092811b07a3e917ae854f374cb5664c97cda0710dd965f83245eaf11fcf3f0683dfafe9c9d02
z292c6930db0886b34b1756cc6c9e94b8349a23c940cc18247b040da18ed94ae1c2b78632ecf73b
z8c92b95d233be28d6ca8fdbd4b22a5e7245e7a2999da00a42ccfc7a3037c8d8c67d018eb6cbec1
z335e8173c5a789146da1c77874b275c618cad2bf5bdced4af7d10ec718e2e1975f8a2f71f07b99
z48706a7dd88579683869daa2799c86df5597d4073a9da8b808e70e4e018484725bc92d757b98c8
z15516b38b6b3df1acdfa7ea63893eabab763d2b8a78706ff88586cd4ce22b7da9dda5952b16db0
z0a2cd47378f41086c56a8c5557b28b71e6c09609953e88df1ba347878a4b6292e46bc080b652c4
za6c22f82416a42561b3b5d83fb5c7a4aadb48540bd4a6aa3e6e2aac60764b53561d4eca4ae8044
zf356cd589d88d62153239de1bbb4d151abd95427e3c5e16c02ef0528a2b8192f5cc5d2ed7ac33b
z2a59a35b7f94d44ed961b0c836448bac1fc4d797ead72dadf9efe03cbf1ab02e28e0e15e9e7e10
zd716d1aded909c4b170a52ba733c1e00fd4f294ee581bd95849edcc8e3a03f238c1a2208c7b94e
z27181163a3d8d165aafd05f90386bd65f3c93a18298ec325c6ad99e39d0de27b2ba47547958d31
z8b048a9fd49cf64cb14839bffb40a6231c3c0985d25936ac6b52a49ae92c8d47829bf579760547
z56862fea719face3f1f48d4287d8749163194c23c170513c8149a2bb5bd6c5ed18bac5369ae064
z7378ef1e61351eaed3c70f46e90f595b6e49de5d731f3d390ac3b1469c6b38dad763a99e4ac3a5
zaab24969562c04c207df284e3c181aeaaa9fe82e51da655900485cc7888784a9e665154ed77fbc
z0d48ac51b090016078d5a20b5b4756e98c8a0fa92b397020700da1c9e61be62e581c7a41efb1b2
z420d460a2f4d0a2d8c130017a62272690f3ac886d5d6b359d1446aeffd92b8d63b528d5be29275
z3775d4cc81a496fb4e0042b79a9770abe160b4f96d9170e7ad2c558095d0c17d0db3ab904dd29d
zfdb53062f76375fbdda064e5bacb24461511c54d3fb04772838db048a288e37a3bc86b6234a68f
z09366a9cb7dd6a2ba8e6b7fef0ab5a32d8e0132c26ac8ec05756ac2ad00bdedf3995ef615a13a4
zc42830345d66ab2729e8476681654d6afc3dd0064eef02238d969f634dc39f77445f9e38dd12a9
z8b219af715099a1474152fd84b2d78d88bd985a3a5ca1a79b105570b411f881e3b1b88a1aaf041
zd2188f50fdc8828640777a2a3656ae654240a9179dd7f27dac81f5bdc5f3c94dc456ce1dad4d71
zac6aaae04a4ea79f8df650d3f6ee8cf1f39e58cace83eba63af51bb417f09e2ee4acd37e7ce894
zb726a37431019c6722bc7f6e5c3c3fada5cf36b5bb5a1091d14af03f8c54e26061738702c14e16
z60c3d54557220a912b1eb57082f4db99c89dfba70777517618f9f48cf0a715b03480c109a59b6c
zb537121c8b227e4d1741f7f5e96b8378ea5a42d8ef6364a7facfe30202f36e63d9527a8de78a99
z79387e4916e93dcec0ac9476f0aeb42c3211904cf90d6f2c09ee41264a8b0428f0bd46defd0288
z73eb1765fcb09d0c95350fb510d3c871bcc6295c6dbfd7314f1752c338cc26435d2d2d0bcb2fa7
zc244cbdac3ee8c79b946f9c9d4a9a2efc83de9b6d2b058748f1bc4f85a56fc65e931540ae49cf5
z2974b0ef454ae41f0d36c5cce8491392c815a75dd3a3e4c1b0f1599f427d6763909d4337de2afd
zfbd960d9a1294ad4dd1c3808d24412233cb75f698fccdfdce85cebc95f999928e14e3303f14844
zdfdc202f548d3986e82ad2ee4572fa33c3cf63fa63d049652e9b4252bd66767846b8d03425fe3a
zdad559dc04b36c831f67a18789b00055b34a885e2fc08109a938f5928b2390c53a9cb15d97b26f
z091f519ac35ecde849b9d176abf9eec2ae03e15d729d26a9b418eba8109f660e5909b74a7fb721
z3be980a81b932c8f2a996604242a021b39b2c1c546180e771ccef9519aa48f135531f0b7367eb2
zd12158ea0d5ab59760983335b0f1327526354d5c6c9cd674f3b78160b1c90b989df2f795da1e24
z7304f1109a84ba80f6ec748ec551b710a05b372b8115ebb5638742adead84729440220f2f67656
z11beb5c5330583cd64c499e8bd9f617db5514e65bd9bf372e3e3b7fabbcb5dd640ab4cd58f7c46
zdb425d2881fd03b63991398fdf866c4a7ce4c6ae36618312ea331c67945f2e2b68cd549530d249
zd888cf7d50404a49b0e3427381f6a8ceb30128c6b322bc1411cb61e3025d4653e0a91732d205dc
z183146a855d5215f72cea01915ca02a1aca5a832f358f81b98ab4911ff163851f3a1dec371489f
zbc7dea56af0f2931c6feac648319279a72a8c5f24497b7ffa3ba687f809a7615cc975f69b96207
zd6dcf0cee46d81dafe416aec84c6543e06356e32788a5d6b502cc1a24b2f6695c7f6317563de42
z413099a9b677ea82b68872ad6e35ef3c469a20b23b97ef181e53ca9c8fcc4c00b8801a80e12d51
z9979424d0f4a5605fb091266bae08df4cfefd5bf0c3cc9dce1e653147dcbcff3eb401d9b601b04
zedd1dc8bc3e2c12e9a5243be971a6d2128cd3fd1dcf84b3b22dfcfce23b1810a4c0da7d748907d
z9ee593c45c5727931e9b3ed4d5fc46fe9a9ed9b090229f61006818c1306ea755484b5623c00d1b
zcf6d2e510dbf4461001a74f1b5b72119aa773005c089b0c636d9a39c886974b2ffc5bf4a067c34
z2e4622c2f0db438d77ead029f87dc2dc741b9dfd40fe322f16b0c740681d06a910196b97402ae7
z615542079b2f32cbb5843c2d77908d6ab84d8da0576f21a75a4e10896ea5a5e56fc11b4917089b
zd73457a5775b84758b920d1ccba295560af6a820507f13459c8acf785afd20a6e8f536b9398701
z2a7f6949bbb538b70d3c371f2aa94e6a3ebcd8dc37c17bce12c491a8a50bb8d01f1e2ab4295ddf
z25a2953101bb2fef767a7f940bb09073063cc9aad12979bf19e972b834a2bc60c63441378cbc3f
zb3bee2a847a3677677442d462677d109fe91b3e4e2bc40c0ad42c4a6dd0ca08e357c5bed72e5af
zf6ae368a39860ba521afa998caad25d42f523d4fb92beb152bf8969727eb4f0c0e3a7fa8abe1e4
ze70e7680d50aa83d0ef33c6649783df098e1169d9769b492fec52e79defcc6fdb3df669cb7f9e1
z2acbbcc9340c644b49f396cc9647c868513d9272a4aaae092be98c09e5cc6dd36f75ec65ae51f8
z0ccb92856ed9f13228cef610cd3e573cf41747769aa944d8879c07057f257e14c7d29ed04d2c1a
zc52aa70b1a541f3aa2273db065aa6f05842b3ed5186e316514fd3e1cacf9c20374f91843967ad8
z574014987eb4fa4024a18abcf388998c361a2dda0c4b984b65fc65bb8e4ccee3a5935ee2132db4
z56656db7f371085e8db7ae5b91871478f58665c3663a1e782d8d61261f60fdd93ad4d9a5634c0b
zc38c143bd802bba4c5d93247c7fc4564f889ca3cd3cd5e29bcb8e201cf8182061d75df8d345eec
z62149449f6e3bcac6d9b3e16edcfd008d310115014ad9c65e6ecd5b61c88bcea0d31d8e2e04438
z363411a519702b97f0fb024be3a9225df1bf7d774fad3ecf4861d9b6741bd52beba6795b864888
ze60b033d7a4a73abdea20baac9cd260a7d0eaf673a6c124e713d80d488655dfe238cd65ad6b21d
z83e6d29707ed69a5068d00d4008e3590997f4b0369e683cb43352c69d14b15c4356493609b1834
z86633ac0f1d01e93f3d084d3552681d3cbf5718984791007966609393db63bb5715635634681aa
z0b2b9ba41a992418d2373704ea9c10afce8ccbca926626fc060f452d937907928be0918882fa53
zd058ba0276619fd03ccf15c246b9b84afa3b6be82b5a4f1101e3a27ed1813e8ff2b7df521630a7
z057bd7dba3336d72f5cf94eea8de326a78b4971acae4651324a64d2497030b76fcee8525a5a1f4
ze3a1e1f3b2415d9ee789711c56117e71bf125f80477bd0b44c209f9b5c952b2e686d03a327d46a
z6a662101b6f504e35f5a87bd98acadf87f30a274fee3e864422d550b3cf3caf14e4f6f9b0a405d
zde844ae49854e8fb2e284d44245ce69aa995d103cf6ab39e7048f011e54c4efcaeddc47c4460b0
z26d019cedff7414e8ae55e78874f488edce0cc4ef9b6b1db2f000f38f2629bdd88f66d0fcb3de2
ze163d0fee10df69a89d1ae5ab68c47355804b51f628b37ec7984ef65c75d87c8eac464ad4a6ac7
zc5dbbae47db4361026700aa4cc88ca3b8f4566b51721ba8d4ff4a70ddcc974cf8c9acf326f6f9c
z8e71f3337b09fb8f79e226d4e17631fe74383b27d410db5c1614a7c0e9b768db86184b0d35f71e
zfa0d73d96a3ff20aa7abe29936086cf8c086360d0f281afad12c4f1fb843a125226200703879a1
ze4ba1b2a6753c7c4a9a41934f6a1005bf45078fc04c2057740404c9145d3472a150bb2a86fa2bf
z4d355916c38bf90f1333b2e240e30a1fe8fd2a4bb0d6adec9543fe0f31828682fab42d5842a2a1
zdbba32de7d512c2f4a03c6fa64fb526ab5bbc13f8a23c15b41198c373d9cf0d7db886917e0e1ac
z646eb89564c3e072f871623f32aa6d2a5f07b5bd3d68bc9fc6ba319ca1f21c024247477e72c09c
zbe45449e559bb11cf453664303fa0a235a88666b3922bebe362ddb9347605b3913f141b8df51ba
z44ada59e3c861714995d3e61bb27b9d2a11e7f1e98d99029f084cf5629547a63b508e89bddc364
z58f573176c1a5876bcbc599ae5b1bc95e4ce7a11c8217390427d1db75230154f9c1a39e0cef906
z50d5dd29d80cc4523f1f6a1f442055265cda5f5641428e80e77b0b6e8f3b587f1765f02f313e8b
z07076929f410eb613d164823dc85a8469061c44c7f5eee71abc1ccac259bfa0a8efd12d6adb13a
z10e82d68b24870878db48e9adebfd91c1f22bf4c7d090d46378de49014be572a2db93db6ca4646
z8851d6b58255ef7c0efff0408dc2bee97e85c8445e5d30fab0cf0ba4ad60adad5fb97afc2d1412
z7e1a6940981e156fd63ce094a0be8414480a3cfcef66c87ed7b89c9971e57cb331f1ef01a80dc8
z093cae6a2603a7bf1dd43b276349c478c67b14b463e758ad813d256fcbfce3be408bb1e4ab2b01
z67a2324c34c2999b30b52532941a8ff466046a252c8ffed9f1a70cdc7d105bd7d7325d7590cce2
zf14bb572a7541bd0294743bef490032e51711dd163f4108c3bcac9fd42287d4bf05c79f61eb082
zcac025ca460cd6bac17b095cb0acb35a0b33bbd89f03dd6a184d815ceb548543f7777de787c995
z35931c69b57c0a544269884a946f05767ffb879f026791d237a9bd7913e7486733d1237d5de9bb
z1c1ba39a088c1c38a1bcbd1d722f97ea0ce2677a9fe80f9273020d88603ac90b930a06cc95b251
z4b3fb760e976a93b15a0f35bf2466f66e0207dc283240e75b09cf78bae0cc6b5db283a4aee79a1
z06f00b4adb4aec6dd33c1ad3e78c07d53d7c9c16634fc4b104fde40d68378c4d6bf3271b8974ac
z46797c2306b4fa2344a95fda7fd0d6754e29a3a89892a44c019325f82a15be66b9f8c8d794be5a
zda246410592832f887d43cedb8f2d850f62f81ab6316b8187630ef7545d09527ca4ad6c0d90f2f
z6419417292b011daa9a5d117832f6d30e32fad92f35dac5cc8d0c086b8f6205974508e258c7311
z57a9c2d297b5a53871ef927d26eaafa0deba27f095205941c59c8b2acfa41723db992e5bc406e5
za9e713d36f9987a4ae01bb2a49ad47abd6d4130b99c76f21429a791d28bc2f22ac2e8c6416f3e3
z517742c3fe3460de5f8e2db075cfd8c607a85044a581feb4001b4f78609ce123f3fc7617097674
ze7c6a6f365059fa07fa2ce472eea76ff995819b57a3ac60174757aa7004a0edc0dbfad189e555f
z98c6d9a1393887dd928939f625ca960a9a828d5ae0bf71842d987614801123cc27193f6f6e3333
z1cf2c541b6375e7b42a618f8ba940cd9a32bee981484c8dc78aeb3bd5a7a1372b5223a3eabc26a
z77b58a1a2931437f9bb10c9528d801335fbaff0c844cab62e9b049a79e87f1c65d18ecb5570629
za436881a35030098fa967d420b095dfa742f8c9c208453525e60c3b0730fd74a192987898ab470
z52decd87f347d90554684ea804e1f12b063d0aa0f55e4a74a9648c8e0c5bb27a7f1b933445b4b8
zadfbeb0300f6523af38624d9414ceba03630216d4a01a8996485e31c278474117ae01d6b428d16
z246674cd6927929af41a448ec40f865c74e91967a3f58c8e694396e9ba94ff09414a608be23dc2
z18824531470b40e0ad4e42189b82ca132b03ad0ce96c5ee9ae1476a4883e1f239e947469e7b58c
z2e0eb7f7e8f71d2fccf193919da0d0f087258c7c8199e1c97cdf37a68548e9dee7a00e86288a38
za08e33c41fb49528b8e3d2170317fb1504aa98af0420d5328a94a905f00962c67845014c36538d
ze9cddebbc04aae9b31b2b63002a90b2a29055e99ed2a8581db8b4bd46c94cad4e38421180bd0d7
zda8d81fdfcb30049915b0bcaad46e89d092d2f1c5f27f1f171daecea5d6f403db7d5f8987798a3
z873ede235a849aa2b7505fa91d07305f502e17b9e838a651a2b6df786e2e017890a76208aaa9a0
z032eec44d5b4a6cac35a9d5b4cb7d5c87cf46bceb93c612e2828f6f766e17006a34811889affc8
zeedd9ca766ce12ab9977ea3ddbeeca7aad22549da9b84ad79695b43ed239cd649b909b2ca2f291
zb7658e62e341f4e01ccc3ba4dd593e93d844e7b27120dcc1611b3a43236003937abb9c04ea07a1
zd9fe07604737e7c0a996587faf3d05e5533bce6fff21485426c4cf992c28aec248e97224c39f93
z561c084dc299b01284291cc98d11a64f47890ef4964935e24d79ca17869688abd80d92bff688f7
z5ee938d39a8320347de8c02879c0ebc26e02c8f6031ad6d7c6aebe62f517365886fd3ba9dd76da
zc6f7246bb5e6b4adb3d125c47a9e284395adfb322a45541eb41d565915ee23b4c552815692d82c
zc8d9b54ffd6d20cfb393e2aee9b86ed7174df7ef236534b3e8a713f0a6c421a286b0d170b3bc9c
z7c85745e12b5de3d29417da42ea3521f9156ea3280f90c05707fcfae21b8f9a709dd9dde59730a
z99893c88dc2452442450534cf45548d2c8c0600479a1bfd547a4451f6491fad4770468f96532ea
z8070a94fc6186ee830f3528f82a7da358f8318cdc878c65001018adc07f1ac8aa5c7fdf8c758aa
zf2235bb1c13ca18a5912ef48b0717e26fdde1cb594eca467abe2e71fbf8ea56ff0c7538c9f40b5
z8b41c27f689d3cee404ba18b6d613dfba2de8fd1bb33c415d48cf6af0c873f4fb4c55666d8f9f1
zf194775bd3eabde668d34ab77813bfcff9758653384ce22ee15eb56f029b264fee28a566e545a5
ze35c3f7371dc01c9690022de74adb0ffb238e7e46bea1c095d8fd6570f6a080068fa283ab11dff
zee75fa64b409ebd7c6a6d576e6e13fec788f43aa136710800f8c5ff60c5b5b3ba5a63dc002f229
zf40ee8a78d1c1569f35cbf8baadf63e6528a613322f3331e28ff04c456b637f1cf1641200654ee
z4343027503252ee8f1abe15cabe89e4b1a2b94429bf88dc36eafce9001440b853e1dca5a1f4488
z5e611a40c7947a807a0af32b033733d0660fd522e6b6bc87b05f423dd2f02e071614f769fd18e9
z1fea26d85dd91748c37f9b6dfd3f22eb6b16bab7a5f44bc95f167da16dc9004dca363d17bede88
z570ff9efa9ef97f88fbec90743608f0a7975a133da3ba229ff4bae00b89ae433080ac4d26b0033
zaff2bfde313b4eee21e627499b4b3a6c3ac641ab21ba9d1504c8f2981061bc8d55d037ede24f95
zf0ba2c7723e322abb55d09cc3575afb2b1e0fdfd9a04b6760d62f4f96686490c8d7f022cb4c15d
zb20b8e00422d7f9d96a13acf7f51be2b42e43a779d7bebc6e7b8be32971dadc2a4c3a52d7c20f2
z3845c5eee43fdbe7ddef6da6212bc50aa71a7f3073b2b13ef57c54045473853cceb5e0e4ed9db5
zdf8e614bcf0aa09bbcdcb135712b29491a942adb946e52accbb9e1d39e419946d89984af746df9
z2a10689cfb5632cb2adb803b7e7077e827cd9fbeff27b37af3f341159380033076928390c0ed0c
zeb05a4e6b3592a5db3de161f850d2fea4101e93637750a9d9ca6d4c01589af665d96ed4d4e06ab
z0d9d74c0c3edcc2444fc71551af7a08856924aa91c492aba040768aadd58d9aa2986aec6ca5345
z59c9794dd1dc5ec1b45ffcde82bca1eb24d1de88a20b112de5984ba01daca3c3f31a08e330e020
zf9cf1b36a8a0ad0be7933b5f52b9a4015402a35407b61ba25f76868eec5ae3d4fe61ad53d3fd08
ze4bb3ff339fbd58d06ada62549c08e7d3888540e37104f8e7f6b3975a9146ea127658aa884ea5d
zee32560a522ebb7c182c21b181248acd6ceb6a4e8708a2066bb90fa5c83201065f9f5923081c50
zc8d36b7ea11f3f6e4c27d57b9dde5122481d35e756f4acbf17b58df13995f3dbb09a04b9b66934
zb9a30a8baf69d5a5d48bad0bbae57f9860ce3a63c566ac08eb2a728f044de3d4e02cb943fdb00d
z9bbab852efad0ef796eebbf01bde61df0ba8f67b581babc949d2aca58e9b94a90aa45ba007054e
z93c31ff2523476910fb6e98a96b44df8c81f5d57ca22283cb697aafe1e36687fe2c0b6840848e6
z05cec4fbf011b07d0a8739fc7c5ab53b138ac0eb4323dc9caf38bf73ed429213af2d47ae679edd
zeba59cd831dabe284f76b975bfa0264f7e97a64f74b5bf4a2ab883fdea989cc9998b7f33d61d02
z5bb527d310e789337e78936b54cdcb41a677eb82307702dc1841c3e0e2f499d92a2174859bab35
z5ad37a0995307ec9492ef05819803be7ac73ee15f56a14d0d54be31a62e552c1ec86b395bec191
z916b75f8663c9bf52d109ba103a85f180c6fbc26c0f4ca836f0cb1718cc4d1fc622f63408aa474
zdb8f7dd445fcc1b6c5227c5330ae3790dbeca78d358cfb61d9984ea55331f6fb685a4a7770609a
z4b517d953c5c67b735bbff4654c980441120344bcd06292a60d03d4dedeface4b547d68733df5c
zcd81b5fa7476a085824624db1afb9bf2c1d563dafb5f15c206925b9ec29deec87380102f99d03e
zcf2a8045ed7afee24a978880f80cfbb2eee672a97030a82e2dd5419b34c84d2afb8e46a2eae855
z53f94640c35eb912244f626021342edad893bd1d7bb49dc11013a3b493592ab59d2f7fb124ef08
z0ecbebcae89e9808a63e76288d4766dda3b1a18d793a18d16db6662d4eec9f455bea5ef7ab33f0
z69f5a99f83de51c6cdcce3744a8ae35b4f6710e39766e6af742aca43141a682fc696e9ae0276b6
z735305f51df0c2d0c5789e20c1f8f6daeebcfa58062c86c0b373e4f49b45ba14815df9d2ad8ff5
ze4e46ccc22d978862aedd424a735e172812861538315da775bb827d326f71f09232098f8d6a41e
zb2034fd4b19c84e479205f8bc5c297613f939bb63c478852a415deb728cfba89cbb5a3d0c91820
zfca32701555430c7e5d720c682b7b0c34fb180fb90ab0d7f8f9cb69e697552dc62700dfdbf50f2
z8872ca4e653d269b277b421c28dfdf8e702f93880e4a5aced52c4b3fb16ac972ceb5b09aefb42e
za7f5406c99d4976d0d739e0383a818e5c0c61520f2a2aabe3725977b19d141badffb20f080abf9
z2e8a1085c11a522d7515e2cea45f54d77297370fd081dab293421c6fad53cddd1ea04480a60bd9
z8fa3e523824c63c30cb52ecf52f91f001865cbcf00c024ae23fac5b37e68252c1bed1be8ed05c8
zff07bbefa2f573c1e5256827d71cd57e1e59bd21018f2b96caf0a8517dd571d6ab4de3a7bb5d27
zdd6fe53002dfced5057e078175a9487b9738d2bb069085d79da25c47430a915aeee97de5d288c0
zb0f1d66a05a6527ad8e7dbb8566604ab0913aa88f17a558df78e955372761fbb4a4c020cc67db5
za6e3f6541a65a819d6105d8eae886b8079a62400298e0c5a1b287df7dbdabcfdab1b4d99fbdd87
z7d64dc8d94801b2aae31657246db104a285118d211efb5a6b51eef55f27b2c6f05c23d3a210d82
z30c87d898af9d2334ae0ec3a272f6516c8b6aab418079f837d7a1ee1721f19cb80fb02ef187391
z60a4dde1374e3940dc6771debc73cd184a5bebc5a9d953b605d7f190e1e5c4c28a59d9adeab803
z093b9bcb3b59fe26389536db227844a481a9a2a24625e56e3ab3fcb84d4ce018a03e36ab0d1d04
z6fa8fe7cabfd4ce44e7c9e24ef76db09c90f413d9187d86773d20e6aee299a11da7b205980e889
z8845ece05f48a95f6a8b056272f01406741a3ceb31654b1152b8b55b025d74265d82a79ee66f01
zb8d93823617938e3b225d72c3ee25bcb74546d441a023baa2a2f062e5c2fec43a6a8bbd2409c91
z2ceb33ba1fa98662db29ea3d817aa356bc1d48b0776f50fddbf75161e6742d8059ad59a1b16eca
z4282c774667d63ca099a0a8fb60344e1d49711f0201fc233e7c26cfad1555ac7ea02768631ee47
z8b9194bdd48a39db2c5900349c3776c9bc2ecd1dcae956b440ad544d395b257ae19a29c136f4a8
zafbe3b48bd38f5b85a4f83c3e0551ede91a6c9eefe51e747650e334aaa9acdea41210d9ed2c2ca
zffe51b2f75084c6379aaa90d22d1cd7087706983108778f8b207319fb9f1b105ae5c4e5d7ad64a
z7ca246310ee4df2ea67a389a96b519633e3195c0264a07d47bdf98784f0560f3edc54ed1224dfc
z58b80ff07a38645b2d2acd6b1a18f4036057e0df64efe717fd08fd278027c5b099a158d75785ce
z1291c41941b18baa7834ad6bfb7d4b89da53c1dcfbb509b36414e494812cbfdc31084ec5c21d47
zb476ed3c66233a1efcd62476f42e576f416bafa70090def0929bff904f1e3297e6c7a784b1bade
z9336cecaaedea2312b2f458a836bcc784a6536df4d88cccb8fb5dd0f51248f9310e7895cde8380
zfab5a6ddbda0e81c509ca235ef804aa301b46d924e6134df3371edad4d545c15a7ecd143ae24e6
zd27a49d6513b89989c5a3209816dfd11bf8f2226ba1f64b518e087e5a4a25f640c6d39a4068f6f
zb7df709296495c65ae9c4b26f036eb34aa805ee3314e9c199aa20bd2f2c28378ef510c14f0ec7f
z1c593778b47893a6ba845cd5673c7ddf9d19788e449568cb84a417fb27f152a8e624a228eb9058
z1cd0d908195a06fc1abf9906a92d25a2713521e1320d1f5649c6c27deacae62019cdc505b4c969
zdf1f7eb2515843fb78516d122f5383e40dc4bbcfb99253db39a413bf60e2a99d26b6d0fe524888
zc6a29a3cf542e55254e1e5dd11e81d0c5469b26709a3061785f113abfb1a89425ef04968ec8fa1
zbb475edbe67a5155d8dd8e76f610554608057c1ad3f74eedd3e73533e83081d3d3715d283c577e
z881c723d699bcbafd504671afb1728ab8c4d1d768ecef71ded91956f62560fab41dae05467dcb5
z4b41484e92e7699db146180d23b7623bce8192887daa5f53024c24177819be5093be1c83650d05
z970e74c7e89fb6c0c6d5280a19edcd3109b6d8dc28492c161a048a10762a182d2f6d4e8604a775
z0177a9207e9c87ae7959f74b9eebe8e16f9b702e805d740c5c0ba7ae7e56e2aee5bd28933d2ede
z9d0667075f4722d3565c4116f5c23d166c7562345703872ff02faced648c025e052617320aa98e
z81eeb12d37dbb0d2b7b505b1aa4045fe0cd04f6e16406751ead344222f27defcab7f8e8d8d18a1
z919a1e5fb05711acf5ffb5a84004f32a531cbf47b963245db19e4a5084a1f83e0d05a25b4d5711
za0c034d42088a3bb82739f59949dc0ed48942a67bd8cfb249655fe71c92b43e49ab49e9e124a12
zdf8b46061c2c19406b52291a4aefd5d38920903df3adeb509d41e037ea9a35ad5062b881b3361f
z0cfdc2b47548b6b378232700b716c81e9d79cc4c8355d92169d2034007a24f72823d99c817e8bb
zb330765f5737d3f9fe654ba7879f922f85c181610f248563e3c1863dcd207b4c5e47b599730748
z9697c561001d9dc96265cd2fb4b68828df65808f7e3ef122865951d1f292ed2fc27175613e0a8c
z28012e7f34df1adf547f9f35b8dfd91f551175ebf6163b6fe68c3e85f4edca3ec39b57ad2819df
z5c280794606c7d1b7a64e5089a208f6c4db6ba1573b0898b48738951e70f532c0125a9529c33fe
z228a4173b071e485eec8afe7d1c8770edf7700b3c26474ec0f7584f2f8c6abf3a01c4efa7b131a
z24b0d3970b8ab5509fc441b06076d3359f080026edac9de3f47fe4e12b69d6ea7ab89928c2b400
zdf80fe1c96abf33ab6e8eaa9139fdc068b8799c679fb88fb845ece46718ce97339cf259b77770b
z88c24adbecb61f367e62de4e67197c73f24ee872c1077726fba8b18038d66061f03c426e8483fa
z665643b33c230be0dac269804e98532bb70e7de89c9a5a5fc8a029774a95d56c9c2ad18342da55
zfde873278472e3000ead97c83ddb8c5d05a5b80c5861def65c08262d0fa674863defdd7d416306
zdd1b7d12ca1628113f9c8e047c7c2be3c70952543066f3854b09d49707217265e2b8d7a84c3e23
ze1d7f7fafeb04651d5c0e2421121a1a3a948878e0461bcee753f27766f1366ca8dd15f4c585f07
zfdfcb688a7f1a5f77118c329ed0341b9598e476fdc53b905d99eb3f2aba49d90390aca38c1e188
zbc75e25d89f808f48a94ab918f381a24e0c527d550a5b92f7cd284d0bc01bdd09f76da6eba3c52
z98633bc979f7b0565408e3aa89d72ffe1a2ba329b903f0e7ea0ecaf5b99f00f37b9308f9b412a2
z512b65eaea4ae96c3d0be189e6e7a45b4dae873d73c5d969be6d94afd8d29bae68e7e0c84d81d2
zd2883661c90f0536facfe80313df962f32d90fb881c6cd6af071967bf6e987a3fd581ac5b3deae
zfd21475efa40787f13c976db1f5d6c4fbeaf139d3e10823022a460a2259f2de957eea81bbc29ab
z697fb95e45515598a248de7d3a91d1154b2c4cdbccc0ba10e1c4056754ced9ae6d1d957efba7c1
zc84d2c8831e6c32a03006045f65646ea54faca2ed0ae9af095de64889e5f978c3b546f86b931e7
z7718c9f8b635eece4a6f94c1aa0ec3d3f2f12f5d01fefd6c9a559026e1e4cbb9c4f0ca480dc3f9
zed1865cb7a0ab1c165576c1924dc78c4cadf910560aee1b5f464f5f9868d54cd87e4521e44dd7c
z511eab6ace05744a9a7267150c876869c9d61767c047c2dd54daa27b733fc6202e5b635b43ef8a
z5e370800412b2da9a810813e56d6c112c221459e647b82f65a8370509961c1deb5370584c0887f
z93e25575746f8e73a5d26492bca8aeaefa659c8f148cf676f453a955a6caa8fc121d49d6b83b57
zdb794fb4fec319f76c605a088f02d12ec328d1bf2181755fc8a869fb30e290d2f2480bef3ba448
z300a13969f45d1e50a15b4b5f85b3223e5bb5470ce05924f669027215aa78cebc9bfd3f0c6653b
z6f5b0b64633d755ac8d97b932d510e7306975e57adc34413828ffffdd50f9987174b5d12a0f62c
zb1c32b88c082d32b86daba4558a3d3793ae6009c1d78b0872bc757267e7b5903db344d51a854df
z7bd4acc0739193d5479879ea5289af4a093cb6eb81dada44a4f45a46d51b62833edb4f6c86d273
z8a4c843616266457f1c518b4c83cff1cdb99e3a747555337bf5f948c6301b51c55773390e777c5
z342f1579fd999cecfa78391551abfd1561e2b3bc30cf82c004c0c27ac57c4a5ba3177820e343ba
z572f00a98e67f086187c26b49d3c7f4158a2b2929abdc0bc965f072233ea605a27c14b36d8c5c6
z5625e8079ee1fb8bc1fa96eea479b92854fbbf45ebce9bc81796b6b57fe80c24b9a423189f7542
zf55e313549addffa42fa0920a886cb911ef11acfddaf0c7d43b093dd822b677e25b2bb52a63f73
z278f72066eb847cc85d6c549bb9ccaf9247d242c4f307a2f45da1d84b64f1446c20b772ed61840
z51ef7642d5df565a27c76d662c1d0561de481ec0ab941a83b6fdc595e4f438d7764ab95bf0dd02
z6002d82a3dced86e0772797fed676d90f7a2f9202e71bc902908d5c798f3b5993b1097fba87c01
z8618408445b01b2f0a156fd78734ef4958e3ded6fa55b08a9fb44cfac5648721760da821b3c441
z9b9cb2e613aecc11dc512ac06e2e9dc6862b231721957cb10f54d88675d1e39d424c97d81a3444
zdd03eac4825ddbca8a6bfc72c762da7ac995acd1a2f1cef729b01d9dc9cadb0a22ee6c6a9b118a
z577b88bbf341398a2a3badafa5d8996d320cff28dad87164d1d02e3089c31b66151324955f1812
z184b1ea4c836919b4017d0d4a879091036ffba15fa23298d507c1b209f58ad7797fdcee6354a2f
za0db37a33b09a262c975ee9dc9a1191f511f7967bf1ba590a4f34dabf79fcffccea7d6c763e7f0
z36987f392521d9cb37d8c6eca8a0f7249b88a7323f34f6b49bd6044033b1bb2770a778802aebf9
z533bbda06920b605c234e1a198d1996731f92a4d9ca45c219823ef9b3d55bf45d943593470f14d
z24b41ef933b554727fef6bff2f712df3de949180536cc34a37496a5fe3a4b2ffb17f62226e1575
zd693da6f32d4d326bde28b6a0117302723b1f049721dbdefdf0207cd8fb306b4354e5799affef9
z7b844dc46d1a5d45842776c0b7599de42f8461270803bfcbfb46d88d46432ceb8f0c72283b66e9
zf19356dc7e9e6a3af42abe00a4fe252ebbc7c0b8df5161cd9ebab698a89a5100788dc1837baceb
z2dd71c0f48bf71b2016e8b7abe3ed952ed3198dae6efc8f1129d2eda9f7dcc46b91ce5784228bc
z48ca514f6aa6064d9eefc44193bd4c91746dff636a616cd68d737be27a8be8ae48c7820f6c9463
z1a38f63bd97515042a41df616ba0a1bca7da17d2100b76b92dfab4de52a3ee3d7c021c516073d3
zc58a598bfffaf17daeffedc7fb889d7a7588fcb0078a045209a3557e5be4e4e2994f96a88d4b4c
zb31c7ef5bc366872f8da43785a8707b28fd9c554c806e8468ec8116b33f0936047e8101369cc7a
z244f61b593437d5576d5261ae46f8398f70edf6ba7bdbcd9dd23ca2065562f458a3779fecd24df
zc4661eb32ec07c13b89ecfea01ae135d187a41de169a0f9c05780ebafa96b0ca4d731956439283
zbbf2de8dc3b8fcdb5848faec898a76d148ca5ecd2981f4dd69f1d9f69eb1345e8e8b7c1f10be15
z2586a3f22eff012a841511ccbf5b74dab6ed8ebee8e6a6b683ef405628d0589a15690590eceb30
z0cbd83395222a9d75a32d6a786486773425d55e4ae18380bf171fd2a42bfd219e4544c7aade9bb
z6c84245094d5f40e5ddd2b948bd4413c68b35a3e9bd64fba3cdbd7364b61c58dba7c620d88b161
z3980c2c1576edbae529acd016c74cea6392382b2fb418be7304fba97b3a4a907498553b1f17873
ze4d43635942ea3396ebf55bc40c9b0310f5a9b11a3c5b477e94759e811e29d95e4fce1a04a4e63
z2c38d83b2ad34b35721b91076755b65bd29df4493beccc9127ec11e537b9ed3ea0a20576fc3256
zd8da44ab83e9313e2bfb6f1f59d29c68002fbb58de39fac6d580926a9135793f43110f94bd344e
z64e6642b59661f97d64a3f5d4cf41f2a33ad52d29e7239aa37fadead0f11d0cc83c789d13b5341
z740aac30d8b759845128b124dc7a11a9b0205ab7f0fc6b6a159806fea3d23b70627e108fb5bc2a
zc341c1953c3623901a09c94dd85133bdff045031bd637a121705f176ee3c6efa8a3a820b76e61c
z4f867f464fb8c9f9e9d0d87e8dd7c1427f7793dd4577d7cb2257b0ee40a29d3bb6fe332ab0e309
z0455f2ff2c78b6b428c04c681b90d40ecd7a80b3626e7e6fee957075cad7181ed79817a8d10de9
zdf1f5a8978b402fadcbfce330640498f97a7e82a0608cbd262df2d444686aa6c63abb4a4ce6f97
z90e282e073f934547abee0168bbd1b63bc2c83e20c4d72441aac2c7782b5f18625d86c9ef708e0
z1871a8f303fb7073c9e5bdc7f4b4492be78a610c94ccd9b20171b95ba5201753bfb71671b52b73
za0dae5616867bb23b1d0a3c68c25be4fc0c2c888deca528f71eda6d8a98330b6aad941bc3d2b0e
zca160a96fde7827d79916c0837a6f68a2077952e67103844f8c1d9336da1735ddeb07127bb3829
z00b0bea55c0c80a99ee934ea5bf0e5d5b3e26533dbde7793ba83f78fd91df651243b724f11b185
zbaf2477f9996527196df347bf8c9fb30fd9a0a2870022b1c2c08bab4e4380265c4822c02de7bcc
za802b0ec185dcab987bce2f60552ac666ae2306ed686c174e96f4221853e1335cc7bedbb504f77
z4ee0d5546b2096821d0c0a32ac1ed67fbd13c21f67dafd6685538c0d785d583eb105f933580c42
zfbaef7de2bb535e3c33b7f36a9a7d1c54f39062ab4b95a2855d7eccab3a0acd65be1a5a75cd405
z70b91689cca9490cc452fe101e67542acd2f5fec2fca1b95a252da36573efa40a2e5f1f70da5dc
zc3b253f2016d55ee1b8435b0414847ca4131a3a8983bab9c9ec1230a470925bfb82ad37818c29f
zb1dcc78a64d7f10c03d4f0be515282d2fa6d2cdec104206471cb953f47f7a317ab5e7283e6b768
z0bcaba0c85dfd2ba4d8a1668f74dd2d0bd0b900cd6bf669324e553b4870e59a4b5a21936364b2a
zb4430e0847c915f01d37cc4ef52df9116c6168b1e6b911c8ad1df467ca78e3593d783fad740874
z15fb8ba56f6255369bab57f7edd01e533e0d39871b4cdabd1d2c0a36776d3b6990884204ac6042
zdfd64d322fa94f9ae94e203f61a55ae487c1915e18a1df696874f01f94a8a5b726f057fa1b9083
zcf0911ae486bcc6999abdb1c01535e01d4cb26572e93b45b1a33f24f1cc005c3ecc5bd27f71f2c
z7812f95c6425fba9b47f96d5e69d843ecfc8d0038bdfb7a197083182d78c76464fe9adc64e1698
z01b84585f00d3f2460160115d9db1ecb66c0edf5eea9bf2f2f014e74880e2733e321a155751508
z166a601d0649d57e68453d8df291d9f446f939191812b6c73cfb11adfa9662478d78aade77651a
z28b4817a2a0e00b433a28d04ef96b8e5c02ee62d726987abd9f76b19dafe4cdfbc91df19338f23
z84cee8f80235c2d67b1e5ba36241094db343cde6a70b3918a9eb540a58b31f338c48c0e5731cf9
z796cc2a43f70b73e57ba786a77a5b10d5b00cda8f335246dce2e4ee5523fe128fb88277e7d1256
ze0ce73dfcba7f6f43571fe1aaf936cc06ef0d0cb754a19b02d066204fa169f561718b127ca6b0f
zd9d8d811314e2ee5b5c3636d2546ad404c54e4ada969f9eb0173b48a8a61e73f166ab41abd5549
zd653aff623e2501137ba944b172f123b118be357bcf57b695d8e417e2cc6576d550e3878974a70
z67cece2549079550f9b56945431aac0e3548e3f889db288e2a6ef09d17661ebe53196f58369ad0
z4da6e297eb79f554c9440f64d1a76cd5145906e6ebc60093af9686421075bcb9f3c9ef830a2063
z4a6b06337e6516171561e463e5d82ffa058ccc11c8e6854f9a8f319df36683db0be4ef674ab7bf
zdf8d64de686a4776b69b379af5f7deb8fdc87c2f13632e8a5b66990320468af4770ce7c6c3eaa5
z74d58d65f91b82b194ed5b91ccbbb543936b60d5cfc0ebd1d6fdec461dfa5756f964a27aef141e
z4d57cc1b4853482800bdffed9f71fc8db7a46744f6132433405b570af6cf93f7c1bbd273220861
z49932ee58bfc5166b582a05713da25f13d78bb5a084b67c472fcd646316385e20cbee9932ba07f
zb57904153ee31f341bdc5c3ead878b7197372a560a69222a98c9eb1e2395a573eb8ddeab5fb73a
zb25155987f236f2b433cccce5a090da0d56cfab643f1033eca7d176167cc4037fca96c11e9f7f9
z8dd50d240c88f427e000cb7ed1efdd2d89524305805bfde80e3a42750b36b552db5332e0c56afe
zefdc98ca50f1e60d311f703b6e13d4b6714edb49d91bd48633ff3838dacb5686fb2d031176acb4
z9a6571e857527e9e05ead56d77d56c0cc38c92f926e90daeb705d9782d2153fdad771f8a606454
z1bde5317dae2c3879c53b5fc65976c3b0d346e206c5e1df8d2617d81a4699b7c189b0da7e903a5
z020c546479ec7d67e261b15739dba22eed7320cc333a519f05e46c95935c8662d7d9f97d2247c8
z75ca8f07d9c01e2aadce83478dfa5797898402207d53748fe5c3d44d6524664bfb18fe77fefd76
z90de33d8ee03fd1cba9f60bbd114fcf84d3c196d903ece31043703765aea49286ac368e23ea458
zdb81e4ac98bc39bdc7c4f5e73b65127009790f015751a09969fbaf0995120ddb89dce2ba81f65e
zfd1f6a311c82bc24b84defb670d96f52eb2896fa9c6f645eda60ec70e83b4fdeca7a7bbabd619e
z92004b57c189097f4001a2f1346d58e8de0e477f60c63343c27a96ea3a3efac95a3d1c3359e500
z4010e625fb4f3f9fbf2243a490a6356b31635608a194ccea3a34d71d6d5491192d7ed1aa3247b6
zed958e3ef926cf637dc1d20aa7feeedeb1b2ea6080fdc1e61b6490f7b3aa677c332982f88676c1
z16a8a3390d37d622bee26dc955a1cce59a08e46f4d48dc6d30a8c00eace73376878008ec0d831e
z18ae3664450ee2479178b7d61830d35205d7e4e2e130b8a8c907480155dbe68e255acffcd144c8
z03024257ae86bba454a98f0671d1c1fa682d02978983327e46f612e4619f681f4c019e72121495
z30e984d8efc7de5f7e1fa2a95d41aba5dee4e46bf10118dffbe393300bece4648c56071de3a4cb
z2b31e520cbc91a6a57fe31beb7919b5620c1358e1c641529b2c4ff01ecf2d6256c3e9bb7f39fde
z42ba45e64d074889748037ecfa3d5e3172418dd70cfa0193c3aa308b2f785756341c7af9fb12eb
z61bcb7a367d1358cb1be95cefb5a410c9380a5aa2ca4f50f2b6d3620323e3180b1a750f0db4130
z32d21e2e8e932b24b61f35c0a75dd3a548e0d5048fe2fc13a4e4b26419233ba981a7432fea4266
z1cbabc157cdb270faa72299bb6aa375859f51270380204bb955e0ae6320f4f8f91c04ec17d7eed
zea48d64873380e29b177e97d600cd99b436a5b10ef65dfb4fa00dd24027e1cb6eb11dcd5f2266e
za205df7ae6da20e62b4e683cbdd81fc4e33b9f2e4a5277cc0bfa92e433bf1a65b0435630efd0eb
z209c2b308ff33c1dad275257e36444a85d461a5bf5ee882b120a246f75baef870309e6fab6942f
zc4b9163c8ff63e9f14537716fe9a20de37678eeaf90a413431f3c8c7bc84097973c79ec354c4f4
z7df983073ef856f6696eac27d3e65e3f1c59245612d1547eb3f3418c29a435298adfbed1480878
z4117da8af7269d83a0fde092e2e4c97d531d89c83c410fa319523ffabdbdae549c73ed75f309b0
z9e9c9871dbf99a3d72fcbb7821ce519e889fe942dbf77c3a6ccef71735c8f177b563dae6209510
z3b69e2152f224fb9cd242135ece58aab024b4501cafbd2213bc6be268469c434ed2fa555b21532
zdcacada38a57522850dcfb74755a1c6fe933bd549e197697d9c57df5081118d779c7c2d949c2a2
z42eddb29c61939ee6d613b6e44320ff1adaafeeb0564bceb84f57b68f54055fcc8e79a00b72850
zf38e6dd0f8c8f567264e92176ce0bbb8ade760a0c5ae1a4cd2420b2f1ab5a24c7de2b369d027e8
zac9b8e8a29afa021646f29dace20455e7e1d2d28b1d6f05da3a16d9c92525432aa8e4c3a8cc7e3
z7e934e597f04bd4c92e4d2c163d2a0b7c0884e62f7abd820b6b589c24e100f3ad9cd61539511ce
zec5439eb5c6686aa1dd74168ed16e0ad9ced919d2b4944cfed8392da074136ba19d533f8d5535f
z2516ff0a601e739c59925dc355fc2eab9ab85a80fe24d86ef645f0cec6d7f57c7775f6cd63518e
zebfcbaa7a8e3b443bef69facc664dd51098fda3f967addc36308176e360a937760b7d9673f8db1
z1a3c81a37876dc6867a2566b0cfae16329084ff4c62ae7fb43e0efec299b671c49afac187fe0f2
z2beb8cbf35b0301c6c4d3cbd43186f1fbb4dad2c4ecc6abb86b8098d9fdfe6ac98953e55d7b49d
zf6fb4c5892a93cc26869970930ce169475b1889cd66263ab101de13087cbf090918cb9e3ab32e0
z4d594d8425ccfd02fa0ed4cc413f14563babb8857273f68ad69f9cc8e5d645c45d44f22f3379d0
zb566c24e7b0ec55c5f10063174ad6eb84dd861153bc652ffc3b1750223a0b45179052173e84ca3
z77edbf8a2f695b0e85593185e5e0ce6fd846bb89c222318adfd19b3ec5a13084b22adfa869b4a8
z42d7008e07b5720f87b9090825645e4452d813bd5d137460ae0a9405b290de5ccd4ed3944e000a
z685ded3cdb97a83f65d7eb80485110bb573ae9e9ec36d13392b2f74322bac1d547211e2e573e3a
z6477e1089846f2d24b9f382f37c95a43a0662bb9641e63216ba82fef6755b9013ddf0e1a177c9e
zb1bebdf584350790c91f1d3572d4d664a390148a8493385f5986cec2261bee6fe7f97d76c4a107
z24392000084d006a36a7b871dd353c9ae13194a9bf8bde71f58dac2c9a1cedddc5d3275a96fc10
zab0dfa64dc660b6e29619c00b003c3ad93eed36e038663e258f0c51a2c20625693ef5b92241dc4
z6789c327e26b26141ff3604a8d8749c6217890c21e009f0e0919a6c50045ada7062c993b159d73
z6ac24219c3927997e9620fe04fdc8da703d511a2d9a8f3213a6abb24b57e54fb427e8f14f9f39b
zacf288ee432be5883e644eedfe1baf8a7857caa9b8aaddef0dafeadef00a8e64071d925b604be8
z5b9b335cff1237e96f4913141f3ad6eec722e3687d23fd5d2499dbecd84cd93308052ce2342857
z122618560789a9b89bfbe2f830e824505f01ce6a0f57dfa989a78e509b196543d8780a33acb53f
zad81085252ead496f1bf155754b096f0b23b64558a5057a6d61af4eec812539f63a6273c0dc3bb
z11fe44fb013bcb75414c2a3571754e517603278d5cad652b128d56006aaffadd89d2b8c6d21d3d
z7dbb48925a889343c1005b796bb09026530d2a58ca97ca8876ec7b8d0563299e73522cf1bd35aa
z13e6b72830f4a3e64fdf1621818c960716f22894e3904cc199e77735031352cc6781e76ac1fbfd
zdf8154dc5a040ec7e582bf10cb94801f98a4dfd6a51d0219f6ccc8c743c8f704e2c0c583e4c764
zd5bcf8db0299dc4e575aa10598d4e6e49711d9a1df88a88a4d9d02c97aa65aed6fa04e407249d4
z6da16f49d03df36e5905e2a861fbcba45f356e8e5614dc6c980947ef55e8c1ed67d71dc9ffba44
z872c61443268b51334c17cd6930d369cf2497cf9bf3e5f3465199f6d8bc426bd3bf16176f65aec
z63663ca7d2bdef847a838e2a5836a487308720c8f4674fd5f1d5106dc253d9f7f1d3ac9f2a8b22
z8ddd26f69a9dd27559ade80467febf763f55de1a9c9e75d62f64e9cde534a0c89414f2237d3d83
zef68a6536441f2634bac7c2a3131fcba5e1e9988245d75521c60ee5a8302032f21afe92cfcea5a
zbb3a7e7fc7b509d8d9133df20c13253852ebe70880c2f189cfef2192ab707f369fa76ecd872526
z0e0f14a297441514e0d6826bba12ea1af8a242b2e7eafb8fcdb3525f370701ace288c99b15e245
z155a255daec346e6c8fa15e7c194c14a83ccdd05669ff56c46621d7a1151886898a9b4f47facd8
zdfc7d23df35114949a26fe53def25e797a0f050aa15dd8fa484c73ce5b69a9e2665905daa7cebe
z64a08a49d35395ee4352b54e2dca42855f73228cbe78f6c7ee83bca37c0038bbea08ac045e9ae5
z6385c1b4c903e374e514ef9db12fedc725a7d68a04c0d88bb800ca75847ddab8ba3054c596057f
zad6ebe6197b437abbc2682ae4398c96c510d0ca16ab3395d51df064d96b7f6bf815ff1b08d9fee
zd8cd93593c0c7df1124439584935e34ddc5658bac637bab2c86d5f8ff570a25fae2966b7ac6db9
z2bbaa163a059dac8e526a206aa8afdab0cabb68abb7dbd6574c4eab2a04a85bb39a42deed50dc8
zbe5ca57dfc66075b8c72d90b2e578a3ab2bd49c5a6fa43702ee5a3aeddee67b00855799cbadbde
z4bad5b8c87ac08a27266482e0605eab4a2dc2bd5fe1c7fca0b37fcf61bd00dd781f2e7cf0e144f
ze77b3781b15a0592767b16286f4be30868b2cd1d369522d9513ab5712d008790f400878cacad86
zfbe5138c29c48a41f285bf6ca07de75c758897b2af484baaa832ce91ac4d71d05cf5efd3c0d1dd
z092e359738b1e04f4118309884e226e37734fcdb0fd201cd2473b0a55e787b3a1126e49326dabd
z1487388f85f23d34bfd2bf9a6b0cba67e7146790e3f90a37675baab662eebb9fd99c014b2f2ac1
zc784c8291a1f5db2d2e389fe46a7e00ca7c4907d4abc47b257e66352d2d43270299552cc74908b
z40430f35e722b5c3552595cafb737ed50a3794a7cc4220370ef7576c7b3afff59f37090278c2cd
z8fc5785b3ffb1c0dcc79c6b2042490b5ed9afdc3b9dcb7d936fd39dbf170c100963af539487115
z062dbc8e2504d556fa29f9f561b5ba95cb452dc06c849eae7d87181dbe8463409c47857b583788
z998ecef17b78a1abac0f599badeeb1a358b260c5bff99b50514b6a02dc89e85851e9b71fce16e6
zbbf8d42874b9556774ad25eea5b42133e236575b39d7d1d011a086b7b52e05a22dabbcfd8d3072
z4af5654cf7cbf3afe45bcf315c09fe2010d627e26d6736dd5e1378d4d8fab43a6836f728d6c953
z5b536f06cfbd44225c9e7ce872b7a2bbd930bda2b146db3f258157b3dc3275e8e9acaec6af36e2
z0c487d508a9cc5ea7a5c95b6649a29f7297e409422e5ebc57275863be50fef5cc121153281b7c2
z582df485250e81fb68582692d98b18391769673baad6dc7b065137155ba0f5d7bab6f7e66ac40e
z79ebb49b4ce8bf135f3a562b4ea48e362a86b20621a1bb67f45b910ccd55c54e35bb5464c0aba8
zfaabef4c14dad8c90e9f591f3a43f43b9f905197952abb1d89075925536fd17d9009facf584f4a
z44970f3475ad7c270fa8be52a8604c15d9be931c0e8d296bdce57aaeb971560afa706198c11175
z85a8958dcf23896b4c4342008908dcb33e2c0f917f92900d145631eee4ebc781ad65b27031b6fd
z75cba0f5a4cb8e7e21989a4858daa1598bf392d09f4705c8151a1dd1e1c24b7d4c314250c3c718
ze7d9c26ce9c90f9be532d74b87463628baa3a1769431c533486e7ff584e2f2d0806fc11b3e99f5
z9cb25c3910b829e8024f506fa826de65b1ad3d2997f7f61b919f7bffb2e231226a3439cdae0b35
z44686159692c13601268fd6129ede6b759b2ac40184986d9ce8d89b0fc4179343aa3f252345b65
zc7c7543ae92a6ed44fb3e690522ac7b169c3d439a6fba14e93952eaa880b471218a46ab592cdcb
z1af02353a680ddcae597b82f495bd6dc0d830bd255a7cf5830ff1aa7db21169393876dad89f3d8
z2d848a69273bdddcd9bc4e4c0d66143363f568a55dc6f061339ffd46171dba1efcb35d5ee3c415
z06f5c7883dad0b24e6edc7727200cd7e51a4ea11b543079db204ee9c844b63a884fe1591462b4f
z9160ea01736c455d2456d1a462f7ad58d7f05a04390f1d005473e7168f477359743fe2088d9ddd
zc4a613adf8ff734aed8c038e15cc96fdacb068a4e4b21c0e6c5e765362ac2ad327c27f3b70885d
ze60623725af841c4ebffbb0b20f70d18a9f8a0831cca2c5b988eac9af0aaff152841e883c7ef5d
z4c6f2ce69dbd40dfd3c06fc541e8662a380cdd35fd2bb7889fe3711308757c97bf16d9186ca8f7
z204c57409932ee580d01b16cc88d95fbeca05919324b1ddb7b16a442a7823ad158c6ee5c186ce2
ze7198695895839e2bde39e95d7e5e8f12cd9b6efc892b48ff73bbb4c3c3cedca2cc8bccb5f1777
z59de2a43d6c2d0c922f0824b270ff358cf0125e5a55ec0435f6bc72c476e0ae8d3d4aac128b86f
zeea302ee1813a570da7a6caa5128e27f2b1902f01bc1579e8ed3d449670998c62d84343978143d
zb8bf839be5a1dceb23d2a427b53869790e6e72ca9e67d7136c7f455236295859b9442502d97c92
zff11ee2ab82ee09774f58accbd22ad514cf4b205417131884c1852c5d626a0780f1dd81d6796eb
zf76fa5f2b9738828961d3922d37eb36180c0ea500a00e8ecebc553500ea54ca9fa5b35de87d6a3
z863a5324b9679bc0925adc2f4092f48d5714bd08021f665f14bad3deba022dc48cf1e0143ad615
ze1fc50c0bb074e375321187322a5b2d4f6ea24b9db1308f94c3718eae36dcc12b95e186f12a22c
ze75fd5a096d14589d9f8e481743b52aee709c6ce9ba77efdde6e74aea0a76f9618656a430cf0e7
z72bb40ffcab1b11df9ba0c22b7d79315ba88276d798d9c867a54d4487684c83411a0eadbc4e34e
zc05b0e3317716f09183776e5c73ea0ba51f0fbd65d4b077c9bfd4a2edc58a4bc8cc56e253b8ae4
zac34e6a54f94cde1c0f3c4590c04bca05c201a47db67ada3a6b4b261748a7a6983c929284c86ad
zf573be7f4d5823558e61a48931a67910d7569b9e109387d658b214aea4df2ec8376182bc087ba4
z89d3e9851fdd24e239db7929337fe8b6f7a1ba7d9bf1841c6648a22d777c9cff64a686ee5a4f95
ze08abde615d3e6e2eeef5a4f3bd214bf884edba76a46f8dc714642661520777b4724f8866dc6eb
z0413307a8c46194ae7d15d379365498c294b3c7a1e65a0706931fa26b64a0f75bc545a07a12af3
ze68367cb1ce74f8f3e75dd88702cc49fe5df781bef25ab9b48a08571c2018ff723395b54017707
z1de970fbe4f6092561cd4a20b4f166d435c4319d4c2356ebfd74a49a8c8b1329b2c22fb5f30a9c
z57deba2207c268755ddf5934a71e3e491cdb9b385e351594f698f91216dbc21617fa2efeeeaad2
z1060ae7009957345ee8646c971eb6da29373cdb2d22d7cbbcef96ea83b7aea81780ceb2bd6151f
z4e97fe149621a0110f0173d724ebcd741326d6657276d6d6302068a10ef8ce1c3b395a69b8632e
z7504de2d25500de5010f27b4c02a6ac7db2ef17a326ce906038caf82d3995e061ad18a2bb31a49
zf5ea786514024fc1ae5c6b88570ae156a0c8b008de25ea9ea5b73305e987e87906e9ac9683f02d
z64e88373f4c041ea40a2b8a3ecf3df7c14121fbb2389800b1a1bbf55b4365403bf6e9f7fa92dd2
z6edce4c656d648da20ca00f7daa2c894a3e29da3217f4406fb26654e21af1a008e299191a84629
z67f3ed03903be64ecbf06cbcae856d4c166a342a355d9081100a9b53c82e8aedac39ec3e1bdbe3
z612e88f2af7ca33436637987559b8e4574f53f3886b8a182bd4ecde3af07bafe0ca85f89cc1cd8
z5f07e984a8dacd975e7ebafb6adae19afa6fe3a1f516134b20d47f5ffb9b4fafbc78f735d88b9b
zf5fe38dfc0c96111a97ffde761c9fff8d6e93c403af0fc503d334891e836421ac9b0b8abf73de6
z7dbc73628120aae6cb04bff094cd99b986561c52c7229f323bfa3afa2d2458a0fcd4a81623b931
z9128e3bc9a793f6e7df264280eec325f9ce6267692c48cb8a7e29e940d85ef99ad7b0646804bc3
z6b6e56f7a0460e9a3d1c268725c5c3abd1272e113eca17c4bb9355235248ed40d9d5f6cea19892
z21b6ef0f14977cf802000af60b6129f08bf217111aa928447b18287cf34f7e81e772eded9918d6
zf46e7569df8e9133dd3a18d9e8602a26c103ef18286b6f02b2a8f79a8b1840234d95eee7fdf4e7
z9e75c11af46a206fdcebbc7ffb9ae106133376b38ed567f3945e8dbf25377aa93bb9aa7d76abe9
z96fe047cfb726c8bb250024d43f02f8eaca08ef240e7993916bf659b0a13ca8bf68b4dbb6aaf8e
z3769714881c127efe95056e1e4b8146272cd779d05e4a072f9a5a81c8a5a6ceb4d84947c9a6b10
zc12072014b4cf4acb8c982f092ec3c5a5b28aa3a79d0994b46ce72876f023efc2e27ac665dfe68
z895fa95516f32d2a55f6d7b9f2021694291d29dcf558889fb3981ca3be7456dadabd9104981f47
zfea6f8750904d7d37929582f613edbcf84895b68d46adde93f6c5373842a3a8f617008b3996f64
z487cd3af3cf8cb44f46d8bca1bdc2d056db83003546011edd3cc9976186b2ace5ffc5d47283988
z08a0ec2a3073f6667dac3155d3802c598c0f65ad5261fb266f3f004cf02bb275d5eb241c6bcb5e
ze85e0f41810b4b4494763fc1431ed569f261d2d751820a7477dc22eb3e37ad072e7d691795a027
zf149d36e7e469acf993f4a3714f2c0212a92412b806a10926507d15b76224eafc7c9f052f1829e
z10e680efca5483654e1cf2798b3df7b926325db057920300fd6a0c28ee07d1015bef6eb0416adf
z9d11730576fe559497a7156e726ecff055b6401e489d93af3051eb70fe5b9cfbb1bf2c8da5b982
zf9a8d2c79edd4a03bb034b8e88e3cd17144d82d65b38362e47de664f1261e4cbc14134fa0572e2
z0cb04d3b96896dae192308a0effd92340d2d20877c7ec3a4cadb27a2bfd2d22577c526633c8d4c
z04754a661fee5ee88e2da4238998781a85abfe9a820a044d168e3226c9e97923ebc082256d2884
z001b17c1df3be48b8293b853e89611b722b027d0a8195ae2d5a5801ec76bfacb375630a70f855e
z39e15f42865152694d4ad6cc6155c8e77936a5975e03c384525d9b7718c777de6074f888d1d4fe
zae4d39b424aabf22c1e8c8f3943b1dc34bf6666e9443e3db4c65fb98fba6be1a8eef26a32cb59e
zaed2f832aad71ed7a7d6b67b297e53af93ea2546cad9506283da424f4ce352afbd7d61c8d0efa5
z6d98a337b24ceec25cafbcf6f81989618cb326b2f776f69d9c638db435bbc099939756b82f97f5
z9ec168fa126fae9a395cad7bc3067547d31848ac02c41565274742abc226c68cfeac61d9db6d5d
zd44c504070a50c2746a09334b670223cbc38cb1ec98e31d30ccd0d15111cf79faa60ddc5bb11e9
z31cce130b4026023a1affb467fff5118ef731c267fffa9fc0debd5f446858b5f73d83b0cba4425
z59786cf6e8e9f5b42dc18cb5e11e694e5250be144227c35b4544aa5db8422ae223672749ffe017
zd69f4beb20f44542049ada463c3ec6ba39e8fa323ec01d2245ac788eb43ee9a13e28ff95a7b48f
z7be72fb3a805f1d73637111e429765b2e99562d257438c29b527da29f49aafcb4311945867f69b
z813087691f068f4c8ebf556a18f29880f721153ee15b0e5cedc3ba9954bc5b792213aca8e4cae7
zc450822fc93dc00883061d568b694af3ac41964b6f171ed8fd6c0165db9752decafd5ea6ee4dc7
ze14b16d1b410c92714babe80a4acf819b3caddeeb00077913b2a7ec530c252b9ca0bfbd39cd802
z622d8e7e579cfaecd2c08b9d76c92c96e41de05c42ad5224f09d4541415795d46821a7e78f7e0b
zd04943dfba671bfff9446d45bbf5f263e805d1c6c49aa56c5de4cc28aa6797b43e311d9d988e27
zcc1f838df96f00df4a7a532e3ed1f7934ee232da201ea18ce96aff3caf7e4e39a29f69ced2c526
zc9b5660216846ff3c549b9ebea8701c784af5fb5336db62570d8d17ae74c32cc5a16b9129e60e5
z3db7a8c50f941ec95249838d27840205c5455eccbaf0ea1148d65541e0c88d2e5858bae0c2addc
za69c854ab9b1fe8e3db94d491b2ef433a11d8e3c1e8200224247d9e865885d58c3eaa55384afcf
zf2529c2688db71ff431116010164a335c6dee84cc8ad2f543369cf8725da2c19f0d415f442c28a
z1909b9d97e91a743c81a52537107a33bd8692bd18a3fae57f9d426af2d0b335c4da14d19f5b4f5
z1ac079cc2cac201125dd649ff7494a7b93d955b4f6fee3efba662ec2b9f59747e7fa5c63863b93
z46a2ce24d70fb1a257af3b1154911d603504fe9a4af6a484a7aee823703e66561494a43e04eebd
ze038f85db2a90686d933bd5cc99cd63b3a411dfcc62e4dc898faf89f66a13b2561f94c01e6d8cb
z35a40009c8cb27ebfadc65e28ecd3d7e42661d041f50c8ec31efca7c88bd70ea89c7fa68706c4a
zf50cfdbe37df57566a3f662b146c4666e099c9417d2c6c73eff8bf4063e24430b1d3daff31eb99
z11356da277744fc8f9049037d4f0673a552a0b5870bcf2399e57e073a43e1fecc7112ad14cb401
z6596bc8d80581132ed8a795318297a679ef6527aa9592ab71db9e071626edc6f02890bef26066a
z280c94e4b205075c8ec88ce1c1408525c55a0383cc61dca556bf841168976960ca866cc3c28019
zeba8d9b9fd08c008e5d6e67fda247d115ac1470d9e5ad5975aa952d1ca745cc7e9d7e9e2a0d892
z119332a5ff21dca180e607b9a14f16ab8a1122cf27a7f7c7b7ff81ceacbb7b7b9bfd7578200292
z8350dd9324c76e583553d524b5480c90a020b4c8bc4666906b7f75c19971071f7a2b2697375bd9
z5c04d4f28bf439b4851c165a1c11bec3e9727dd9556c36d863664a8b0bc9088e95e15315e806f4
z3537c549716f02a9b896e34591a9ae6c2f1fec6310259b658977440427426176aea13afad2c723
zf22c0f625a468fa204206f70f8babb20c75752d29fc130604b5e789c2d59310ae44afc19819ade
z9aa12f57be4239433658b42fd269457ef2c502e023a69f07a516ea457529199b71e6dd0acec1a9
z393d7935fc08f3ac273b3df279c659198f17280060eb2e680919e74bcba906c5a800f72e920ec3
z75bf27757f796ed3615294786d9b84e9bd6566d2afecd1b13436817eafe87d2131170e24f71408
z9024dc156fdca8ac81ae38c61fdd9f8634e6c24755fc660938dad08a7bc700c807ada0a4e5a9a6
z82644ef9432d71088a1b3485af8c169238e336f83c7b80c3842660282985fe2270111e1d1df4f1
z0bcb018e56ab6bf3f2566fc9bae78d4dc86729fc7b2d391f1918785eeac10697cf5176390734ec
zec31788d89f12495d5e98012a6e2a58cd42896b0c1d5edc86598c6d9400aecc92c7f8749c8c46c
z99695185caec87803ea391cba7c9a5f47f93e4bdb24524fadf15fd6d00237386caf170f98d92f2
zeace29023708e998df2b1ef533a4c405615cd060d7e251940b6b3ea0f096b24cd34f9b4f5bfd5e
zab9f7f310cd04f2bcd5c09dedca1cd141cdcc1be722318bcc98fe45e7f98fe9116d2a8cd49bd16
z8cf0c08b0ca81954b145766c02c41357272b966883fc28d54e7f9bef6c0de5edd661a688544940
z7fb9a2254665682ad65d9b2a2190141e79d8436f19764ef823a4deb4248cbc5ae3617f1ee9f13f
z09de0cba2c5646e4dd6962065904f92b582c509f85c25d6be1348a04e6147064a1bf8aa3af477d
z8b38014cc693e2789604377b386958e5a874c0b701a4d4e386b3aa6abe20051569e25c5aa6d307
z4550b88069b2f19fd0c104223103e181b5bb84f767d0aa7369bd45e132222b4082295f6730c1c4
z39a9ed33d295856b0d866e1bc969c5b7e3ca28cc5b319db01a64403cb02a3258bb25105aebb1a3
zfc811b0b81fa5ca6b9c5745b080ea392ca8b6319fe9fde9538aded297626c91e284b1e7d72c45d
z57926e1cb88ac2bfd926904204eaee4fa2202258a70adebda080435b930a2e5a81350c4a151a9f
zbb0341f8148c490a10da72cf7e5b45048dc6b7cec9b37643915fdbc36ebb0d4989ddb06dc1bab6
z2ce1b966257a098d618746df315f39d3afd52a903f9b33c601f901ecbe82df80d9cbae5fd1fa49
z08a2f0eb9098e9a767e4a8c65d6fdd4ef818aa7f28c588e1a9845f0571095b55a7becfa9ee8570
z6949afd4c4a38685452cb17a7c5af4ea5fecc0b02c8bbc9192268fbec2bdaa2b2c8af3bdb7f6b8
zdd707192aac2dafeed3a48eee8d89f2ad03ebfb81881ba63526fc5f5cd8383a4ba719234314a54
z9177142c9e50b47b408c178afe92ed9db65ae94f632bff10af079f8200019a548625cda70930b0
z68e9dc2c85973f06a69955ffd04603433b2d1c95231d81698f00c91109a2b8d3db4eee5be46fb8
z6e95f3a500e0de2adacfc60978686d4a879a139ab1d534f548d3c0b847818ce62f4029c159f146
zcf900ae3dd6c34baad8dc787aa2e198a746567711f78ef044c8a30ea507f2944efffbefa43be05
zd68e71d3eea5ee1d117cf659b2b30d7c0c5949f03421c8d983215fbcbc53ae0040f38f73443bd1
z9d30b388691887389a6f0b6ff123fb2c94b4f27db0c9b24dabafd61ac3248b2a0f40245dc1bf96
z88e3a8f0874845a9f986dbd3e97145a89b0fd2ae0e7936e31c247d2f3809771aee3e700c2d97ae
zca7f8f313a6b947e70954951893da5836f9d3787d5748b32d1e3227419b8f65f9e18794f0e2afb
z40927f1be04151740766484b62ad37988c7ea4349977c7a87a68af51b38b1e72b667f8023eb6d9
z51b92c5cdac03e9cdf54fad418d75d4bdddab53d43342563c6a9d357852643c4de4c5c1b2af013
z8f7ac6dbb7e43408fbbe70ae00d74e73236d2174d015d444655e1ce525eda529d9543b89c9bcfb
zf5a147cace9ed0eb3146b3654790d8527ca3255bb66869437f5ef375981bb714cf3c269b3c40b7
zbe6d88e263a0f8827cd076c6a4600694c5c01c7667c9b692b51ba504554c81b6be5e117a3b6e2d
zed751dccf45e2464f598b82522396cf3f64a1ff7fc31a9526a04e88a007e1d5e6fca10b87a6c4a
z85c9058fe8a78303b0ddebf7a284baa8ca209b7fe5d40da5a348f445414a1ac2573a75525a8136
z7485909912173b57ea3eb6d2b75a4fde93dae7b9eeb7e873988facaf9bfe87010c692449e05283
z40d2f29bcf1885d63d458f23721fe15f1eaf780eef72b3e3dd9dd1c75f8d09a0dee63df70a1028
z76c7c415ffa224e6e11ef155db8e720ef4c860781505e4974d3cb5ce48ff827ef4fdc86872dd4f
z928daa97ed4852d53a16cf6b95501f940ddbbf36a7ad237b7a393d5d497f0d92fbe5e749067418
z1254feb6b190e3c29cd0c1e82a8acd8fefb27df4baaff3eaa4be81801b74810dfe6604a430648b
z1102f90a593ca2506f727bfc767c0a0bdad9dee633f74bb65b170d358af153f70e577c5cb999ea
ze999492fc2c555bbe774c5c07f0d7a6b52dbf9b9e3a2628ba36e3471d97481aa40ff976653f390
za2c855f2ea60b6e7bf7afb5594e8e7eda5c2b88da71e8609bd0bcbc32f09ddaf6fc9b85803b40d
z34cc46e2a104d19ce875d1d970a92bb5254e0b32d190ed8167f84bf042e2bc32e3281b34ab5d15
zb941efe89e09e30d41e158d82b838b79f51d6e580aa6e6f6514d6165e17ab4d7e2d3d2c371b436
z4b99c842f179b8f0f1e9148330f92b5cfe91e9e673bf8aa07b1800965a5d7426c03ae4b69bb009
z841bed6f9ddb773208094f54f325bdb5f4e2da8f267403bcefc33178f690ecb4195721060ecf54
zb8dfb66d4f236767698c691bc7cb37e1f5912088c2bb908ae68ee1dd31b990be8774ad49f57c2c
z2dc4c67e06e0090a06bea4ddf8b675a49d9e161132c2ffdce64b784c46667882ef49ac06784853
za215c214617d7b1d8f0f4a0be877eb8245b68edd6c262c2e8fed63f128678512742f654fe0de8e
z26187fc9a0c879257eccbe16906a0855fd833de0c648a13f7e72f67e1a7062b1174331818abd5a
zd93c3823f72bf54cec8947cdbc36d01c2a0963c9bb9519d3a6e4426a4c4a07bd070c209c4ca285
za24499d468d2a56318ed9a434d2ddfc776518c5212944898b0f65515b278a4151318ecbd5914f7
z2a35b51741c8f9c812ceb534ebee5725ae90f2318b0fc5f7701d7a78d893068b251f5bc15676e8
za7ec5be912ab0f0eb4154930ff8e5cb30303803396d2b2f381470bc47972e3dad49fec3882babb
z67f4891de783a8452e3a6364cf83293ed5e5edc613603a77f000a239c1fd810273e9916410d591
zd53b49310842b1524f6e2247f7335391cc47629a1f561187e4dd74a11ab32aa063369ee4fa2068
z787c60274c120fff7ae40cb63654e083abb69275095afd7a9feca028e567ddff83b3a22d1d8103
z27235e6dd7b9810e7b7bd965d55cdb727e22b1285709fc821a58ff78a213da456edd69f86e8f4e
z6c5ee2a802d367bba6509d99897db60796f0bdf3e7bd1c07a65928dce15ee2bb0c1854517c639e
z49297dfa7231ad44ac4288e7dde5f63d373681811f54706003690204b95474eb1ab2edc30cd0ab
z98d9111895833e755036d1593d57bb57e1b6d972092b4c4dd1e62e6d5c3f9c58e4d67249a9b569
z39d7f4639af1ce5bc9ff93ba02dc68a281242cc8baac22bfdade8721d4d0a32c06d59370fd279c
z5e0c8766e8f5ce09c296bb1687e1aeb4d6e0145fad10acd31a9ae5abad128ced9dca7361f59eb5
za1650ad1cd7cf866642ae1b7447852f9bfb77105b17f263552b034e6c0439e78de930d3c45632e
z7c6803a26533c07920bb9e16b0da714ba46af065c43dcd05370ade0e01973c4545df752f5e150b
z6a18910bea90b80a380805cbc6f72a6b54096c8a6cc7dd303c92fe7c14c5e5787a6b97671f2f6f
z989c6ed25f26ed2daba95efc8d2d9fbdebb1b5fc0b87fd6e171522256689d77cde6c9c6bd94952
z6fb72025ec8d651f34de2834f1ba1155f0705d5d650bffe77a1b6e9ad77bb1c9d466974982c224
z52b4ada8b9c63bd487c509338ccd9d39c43792fd4a46fe19b2a3ee30c61f3e033165d23a03c65c
z88ffcd1dc64938e43a29100bc2143bd7ad294564ebebba5342e1e77c5db2090fe675afa8ffdf52
z92b3c27d718b98d2e67e2e9c66e22ac57072a2e132db82d5746a3da64950271606e1f62716c3c8
za292eaeea1850ea12801f5b100dfbc3a333847e087012bacf00087c42162b15c57328a980cc64c
ze8949e1ed7fb56eba5fabeccfadc20ea2464076abd4828a883a9eaf58780c7e66f863fda1b84be
z0d7daadfe99a4b266787cd5b0af87204442a2abbcae19d5aba545133e62b5a2ed45608e577935a
z10d4df7c44ed41b1afc5a87f696730cab6cb9d25550b511b01657c935c7294dc925313618a69bf
zcf53bf0b11ca4fff35b606ba52d18614bf70ca7b81931c5eaf0bcd11cd3af67fcdc6d6cacfeab6
z780b48cdce61af6a2fb3c8582f6f53b484d2b4dc07a7b10fff1705f3d24a9256cd64004f575765
z82930d0aaa11e2b8f2351bec18819bd356ba6febdc7629f148504ec8ece94db4b0d71cebdd7789
z67aaad5c23c5162f66ae111f6b9a2a8db561ac0c4ee97ae111884bc2daa7c0ce6d88dbe1441d24
zf88b1ef0333a1f66164669705fa023e5a1179f0d355c59c2b38416d9e2e109e781c096faa287c5
z000f49b0652d27da2bf791cb3b8cda8b5f79334cef416c78f4f17334a736854de2c55034a92169
z8c00a891af42971cb71fb38ee4d0d7504b75ec297de61acec42a293cac455713dd26a0dc578070
z9340324628d52b4a6458bedc2218752c2262e86c936557e4e94004c6ea8f556cf8c6dee2d9ee1a
z84b5446d3fd8c26391428f917f9f680bab39266b82534c447c91798429e8705365e935fcf78b6b
z558a323f4031d73b9a8cf0ebdcb95c24c6c03e2756d66216d8743e98838e6393d5608941177083
zddbf09e3be42f1f7c01e25fb2e959e51c26d2a73b70f6618214d4cf86c8690d657d7d04d6a307a
z884dac3fe0ebcf6661fbceafd45a06a1362ecfe9948c07ec0b99b0e23d654d24b6a816b37c7277
zdd4e3aef4c51f56d1d4f3c45104ab79969f847181741b044f81fee531217bd7db6ad1b32cf6d0a
z1d73cbf1a2c5ff7ea1836da445c90b74d8580e731bdffa7baa32da53c2d705ca809bf86439eb00
z63e8d679eff2bb2177d2ba0375a942304363646e295f0a4069e30535df01bbee0ca5a56afce31e
z2be1503cb1a58258c50dd05bdddf0eb7b2ed108075f2742abe17128c8e2e8a6a17b9e4d14b1c02
z0e0d8cc69c13076b47e8e4b261a75e453f588c93ea3bd31788554a18ff1b62d3af1428a005e9af
z5aefa98075302fbd300a2c656ac03694c9300e4e306e48208c5d926e0ba70fbe78deade846ea0e
z4ce855e113acd83dc0e773a71e122e99b7b79cc620220da63603dd5520eb4d9ad50d58d7d45a82
z25f274a236176d7c6e83d0523c396a9c4f088bfd3f3c397bc61269e89f4897f8bdc6ab78ea7705
zbff96dd3a632186ce1c7ca301fbbaf404f74b1356656106319e0797e353cc2333e26e9b299ad8c
z886627acff0851241cfec4056381f95bef462add49fa64ea5a1848d600e3833bc8a013bc821fdc
zb600b37c05515d72da0a43417940738bef83cfcf703106c21b06d0127e51f1f7d55e6811f1edad
ze6fa720824124fccd0af19f5aa4d2c2144c181aeace6e9aab55591b3d0a41bb7628868ae38f1d2
z5e3695d6f3e3df1a9e0715d2cf35c9397f9a7662eac64a5ad882ffcaf9c7d290caf97666ee8843
z946eda0429defdd7a187c4f0c0e544b4dcb8e5bf6882097e128d8a9b8d31934eb0f1c8852b6a87
z298e3470bfc0a9e26b2c8c37613dbc03fd2d45f9965c770911bded225f0acaba16cb82fcb089e6
z3c88ce7ac485507d263f9fe53b8f9b70bc8c16a12ea08c51c69e2933b89af0341f4cdf9767280e
z581c3222a1a1461ec311054f201d764098ede7683886d88870cf9aa3467bc555c2ad7d538c08a9
z307876bb5622278ebd208a491427c983603523826a2f78182ae2dddc1aa64a43a25f630712c249
z9fe59c8247edbc6e0560210ac75bc720408cd1fbfb4d1d3d6de67a3e2a76171ab7acd5cff1bcc9
z3b69ed2d8aed0bf9a3fc9e57143f33fd61353cc7c6eaa2aed487cfa4b532923436d89f0a224390
zcd0b558330f47d899ff0e84ca38b47400296bd974b73dcd04fdda94fa1352ba79f906c1e89d9ef
zb6b3d92ea2eda257dbab4d78598a49192b06e23feb4b4589af7eca5fb291fafb09089b85fe2ca4
zb9f1f9b9446b250330d37de1fef1e2eb7bb85be11df61ec7c72442cfe47821d4a608e79a17f6a4
z0fb354d61665e1b185ccc12374a0ee4269f38410552b202826d613f25923da4392368440eda062
z03a00a92082aa3ff4c1630ad74cf4833dd393d845224ff32176c1bef7e47548f5c153975067125
z44e5b4f3669d8eef2849d25d1181eedee91bb5b98faf3fd64d066d86a876041801196ffbb73f35
z0beb4767d496a11d0d34c7525ab4788b58af2df6c60a2370f7ebf0930043ca799fb1d7e6d4f1a1
zb53fce52828f75261360c52f116071d6a10ee93ac5cd3210860b0203222abca27de9e5a44ef4f2
z9a09388f1cca70927b7ea5524343299551efe21a05dae60226ca98d02b45f02247a0b9ad14e37f
zff341528ed362fd02bee2930c53d1ae9b5b0fa9ef633eecec97697e30137d9e53ae627fd5c1565
zf0d8c362f038cfbffcfe88ed93154bcd8afc7f85ec5f4cb0769a7348685ea439da694ff54f5cfb
z2177080b8694ec7d982a9f6b0d8ecc48ffd8bfa5f19e4059b0919f0ce73c0186aad151f8144b5b
z10bfe656b8e6460c71365ad655212638132a934d10b42488fb83d7ec4216a729680912108e59c3
z26f2d6084f3acca7d04c72412493712cb26000866f7fae6b154eb0fa3a7c59fb18c123037e8481
zdcfe929823bf3a9bcd1e7a038937b3acdc6895d6bc52348ddc4178cd6028007bd2d6b57e1b8c9e
z345c5a4c051596507c8f855240e92f6081b1f06c2611c49b97f53c566d5ffdafc726891d46048f
z86256ed58706a885ed0f5c335c77d473ac678d13a20941f896bf732e4ef6a497c1043e4542d7e5
z2150d067e43f0781dc43f11fd3b8d9c667c74f2545f85d1d5b472365bf392899317f12a7aa4623
z664b91b01efd06b031f34888a2dcbedbdc4928ce6eec64a8e02ba798aee61f95dddbb553c0fcef
z5ff429efb73158e297f6155955d3ed7acc3c693f791d03cf71f6335cb356eda4375827ae869040
z44c34acc1aca7d1c6079ff1910d53fa9aa63710d39173f55737c630feb1ec6e9943769100ae1db
z6e6509bae549931cb76109b640bfa9e341cdeee993e5e50a7e7508c3df8a5ce75359168fa231dd
zffbea956b0ad9ba96e23c2610947c556a977b84f4b9845c24fdb51d75b5dab4cf6cfc840dcc3d2
z169deb05efc7c9ff7775712c208d2c340ee148d20a4bfc1d0d1fb92a52613cb0bd618c31ae351a
zeadadc0756e9a05cc93c89dbd8d9d82f503e140a79dbb7f050cbdd515cad21caac513745ebe433
z2d52487e6c91cbe85468da1f1e5aaa9523540e2fb808e6a0bab4c5aeb7cd92b6aea3d6c559e9a6
z2c333a563a26a0a6ae402af31a34946526f4982bbd4c1c95b28ee7745c421c7c3b512fe4b30c28
z33384c9eb4be8b9525a5077401a63e9270c6cd171a185916c1e21731b5f36fe936b26adfc9e304
z15321e721e5d44cbf210861250c75d52a637f545b6fc655e5b28ed0396e87c84ecaa9cf61b3264
z9171739b1e66e00a2eaea85e9fe12643a8274482a15786cb780e6d899443c9818efba6a2fdfba7
z8a8f5879359cd102142706517a14e738c5e234c8f24415bd487b06d85de85dfa60634890520d0c
zbbfa5584385d66f4b622415b637730801ce3d410e3cdb50777a589e6648ca6a622063c21a8eef2
z726d4573c2c5a8900ffdc16b0c6f570d5f13478dff1622d0b8a18f9dd85e7735d6adc0884bb777
z8db171b87068224afb8e75ba7ff5c96d9f437b8e8464d271f902c72298af2c66914082167118e5
z2471e9fc0f5ba506bbb8b025e19fbcd45b39053198d7c43ba756910ff8331a634ffcdf853af8d5
zaf29741bf8171ee04009fe92c0f417585fc938122c30a8d18c554fb8402bc9846e5ab02c8b58d4
ze7c450b81bcc92bc61ca98d42dd6a0e86911768f19e526e22187750c2c6f218388d99eb372d98d
za493156ee7a435cfaa9c02690f3b5998310f18429a70d5b715360b2daeb54b4405a3df1f75b8fb
zccdf87a55d2a9090dec715e80622be938e9fb185cd912b69f48d3f1f39c5724e7f302936a5699d
z216154ed0bd838303b23c82886d43cfb3a96988150dcbc69de6f030c3c83c7cfec44fde6cb5a1c
z650c210a110d21a77fbce95d06259968e8060d637590b9956c1cc5879158e31de04374553da7bd
z09f8891639fadb9d5a7fe1c2118002b33ab47da1b6d2720a952f6a211587b3b38ae1d454863f78
z802d1d9e2e8c1ea7058c2d211e44bbb211341456348727e0395f89887c447bcac459707d0cd79f
z4040d692136ac184b4321567c3bd1c563f0404f2286a217c50d6967bf1ce697e29ce51bb8189bb
z9ec6721f6ced8fe27384a500cc19146303354703c2f3a0e4aec619061c82d308b2ae9ff7ea35a3
zbc177a7d0bc54f91f722f901c13711b0e80a472303f82dbc4f5f56b178c2e0d0ee5f60a1038c07
zeb728db01d5bf81e26041967caf3c1a10a829d72b1c12e099be2f6999aa017f14053ea984a4583
z03059ba3c043873f56e4b9a7f7d3e7536854175ff8b735196afa8622e67ec84608dcae77643574
z6fe0ac5bf1f2995ffe649bc172a592d2f55dc55cf6bcd1aa84776dc59b53c164667f8f4d2f64a9
z5d53ace065b4c85ae3e4bd8a006e93daadc2c751d2e53396c760d85acd674765d3dcc12bfb08f2
zf0a9413d9240d65eefc334f7d02c15eeb64c2c06204fcb10ed204eec94e30b81cee658522e1a44
zcd664306993849a15295430ac44f29775b59d199147086e14b6a07d5087f0e1c8dd70d5028f0e4
z0c9f168311979ca7c9636457142448a7ccb6a5e4478cf8fb471a1c48bf719c0e3da2b192faa9b3
z495387eb7dfc064157e89ed1e35a391dbd154140ad164c061a367100255477454a4571ec15209f
z4091b366b60cc2cf517e49ad3eec5d2032e72ba78e731aa10fa898fba186185143e6f3150a5219
z244f49060d5116f096b2242039791ba6f039c6e9af2a24031d8070cdb8091080478d3fa2f9dafa
zdf6b753dcfbe591f555596c11aaf9677ff43b911fda6af615e27604898084a9c670f7a94efa27b
z612e262b3da3001c8a077b0be6a0e66b7e61a7b03922916c4ca6ecc67216fec80896604cf4dcf0
z096ab1a202d45ac3bf035d2ada9299c44765f5eba7186e1cdf757938b50a4ddd6ba54a8a5e4cd7
z1e280c2b1cb524ba2f8740cd04a9144fa42ef0de0bcd5c94914ff166cd006a77ca547337e0367e
z1770eea3b11322057fd318e26534eeaa5bbe2a4d71045d46e46856ba38246d19e71d32fad02763
z7f070b4d2b9bef7d1c7c17dd08d3de984ff3b8be3a7b95dc39298d10278c62f79cb777a51d1fcf
z09fa44009ce2a3a379ab6d1d8e53064c84da6fc59865685521aec4e605796e30854db38636b185
zdd6fee6b13c336615d549668f4e9f8b6e2830853259e3c8be6f4da2f70e6838702a8722053bfbe
z9390e63f0c88559c661a49fb7e423f0bf2cac892a55f74c345754710318546724cc3b4b1d10847
z2abb77bc33f251c76441aa2fa0c37117e73ab5a4cb1f18ee2ef463b4dcdc6b6ab1aa63f97daada
z561102463e05250f5c2f960dc5072883ab84dc4bdde786bce2c6c199743bb7c6c2ae34e3d7e6ba
zfeb912d70def3681589134c7f0d7670708e9684718fc770c988d3bbc9a3b4a21a707001b6c8835
z7a9dcdc163bb8f32b77315d7d440c029dca691308515ae45ad7c72aa74d1b5586b8855b291e4a3
z10b644402c415c8f7c513b09b2e277d25f062dd7fae1658952d6d21bc3b46464424d39604c7e0a
zafbf76ee84749f840f74061ced33607f4c5029d6d085ceffa01f8f445775f80dd2519ee3c766a3
z3e0c71f1ea340c3ef7dd6704fe35e5a40704054471622c779b77d93039b635a14c9c6347a1ee3e
z6b6ff5d5bef097b69bbe74242641bb66c871c26e0ea03b4e55b4bd71697237834a9b01267fbfd0
z931888a441eec6d9d4d48e9d14d7784bb1d71fb240dbe39a567ea07a66c6059c9a78b93fcf5a5e
zfe64048488031ba6dc8214ae74103d5109c83dc15b253cc0c52063e6bcd6dcf041d5a49dfe6d2a
z243de269d69c173b1cbab15fa073861c007bc4c07af7b5398f780cecd10465053cfb881c4161fb
z7888c44b2a04203074257eea605df82b2b2ec9efcdff3e87095486195940463857087caba976d2
z879cbb30b7c3605112e436e46b04310a35535322adad51284c3d723b0b5f4271372b04e330a97f
z281c3dd85e57155e7690dff5ceceec288ff38efd47ea7ddbb99cea902c7be48845b718e3a794cf
zd4cf96121c741c74176c3509f9bb313b841270202dfb18e879ac762addd07b12d7cf5944b6e211
z05b3a230b78086084e8949f3756d6df02e1932d5d36943c01223aec7a9c1afb7e4d3962766aa40
z750d380ea035348e17311dabd5dd4602400e35c38915ccd042808df4be116751479c11e9af74e3
zc04860cf3fe80037855e0ed7be3b5b57a299a7e2693d09968876c3b1066ee9c7f5f7885adfab4c
z7421afe2bfbacb3b8eeda77fe8b7738ecdfe8c8231928ce939d580d257af55d6e570f5ad8ca9be
za63d77df923a0d3146bc49e9e46db7d80a7dcf02d5d004f83b958809e2538c4d2b41098edb67db
z9cc291783b5f7878ceeac55593814fe40e62ac1bdb06bf357b64728567cfd66aad9eedcdfba0c2
zf23af711ecb66f47e6a67e210e06a5f385768ce7be5ad0a3017b1dcb6018675d9ac36ea935e4e7
zbfc3a5f2a91b0562cfb87fc807be5e692a83979adc5f92514cb5445b7c80f4330c661d2892eb11
zf07a83b362637575ef4617378cf58a4db6f54377e4befefed126c0e214187111bd364d912ec332
z90970f820333334043980cb2daab9fd1b7e553fcfe297365de75eb24b8658b4c1312a9a18f5f19
z1f210e31fc52c007b5f105548f20ebdcf2afe9068750e7fca6e0a0e17a7cd8346162dfe5127f58
z66f630edaacf04f1785e83cf8bc634a48be71b07756ec0bfdba6b760dfc83be101dd481a3ed3b5
z0f81577ec4862f05d7bb3950a096b704c8a932ca0cdd476804a1bf5b9f68e62e9cecd499e007da
z0b1eb8e4b657f8a32faa2cbb1516e42525396af12a3b98f27f9d721aafa4235f92988df903d598
zf8d75156576e5f694ebcc377628f22506301c946b54c30d6aa0e23b3f52c3043e29aa1fe5ff5a4
zd3e990b27c0d61c62e0d1ae6d762d550c4b6a29cd905ac75e38dc3df4b1580709805fac43802a5
z8b21ea570c9a6a42a4e1ae86a15e17b077ed722c35ffeb5056dd8fd1d649120f06d7e484a510fd
zdcd5eea7222018f27c058852f42f268044b95b754206c487f919daa8e2f1f297d91ec43ee02543
z0328236120cf62c34e5c91ab17ea3f0dc0c07bfbd76a821ba973124bbb29ab2aa12ed773c64fd1
z357a38d383e3e444cb3d873c4ef12da4853e2c52c01ba5cdcb1b5d8ef011f9b836982c3899a26b
z9cff07fe5b4ee283a663db43e3903c30d63d7c055b9405b7dab0401a8a48c7df646521d153a6bd
z10785fdd73cdbeca65aff513231c0607d926f12dd739591e67cf5ce219cf0a75dfa01aaead9b26
z063596c3201b49d23cc4e6596342218a8202766b6437d207f464ae894010dcf62d0499b5aabb21
z210ae0c54912d0038cb70d3405cba270aad4860c54ed580bba35079a01baefd3f1ef73e80e59d4
zb3456bb278ab4eaa0486c9873a11107f9157384e09c71e95cd6afaa2c94923e6b5f9ac2ee181c7
zd33c3905b42f8eca900bc634ef8b451ff72dc54bb3a94fa5ce5f6830567b01912cc72a1dd1de16
z09f6352472bb4ff47abf2aa6fa16d5fb1d745cc853be60df0b1980bd13829501a11e07c56dccc0
z8dbe6cd2a71facc3471ba443c6f87be9f069f4097dec30391df273aeb5181ae1596c3b08d558ac
zdc4890b10c34ffe7ad9fe213b37635b2b50543acca911cf140939811b46538f958244124405c04
z7d66d2024b2ade171cfccff8fb86d1037945c358341c77ba275a2e5f76bec1cf202047a20bfe99
z5a660622bdddaaf0d665477e0506aea1b59d3bd38d22134eccacf19200d671b929b8a718115261
z37ab31dedc0c03a79c0b7b4b1b9405243b322ede34b8995b17b3af19abcebf172de00dc082d752
z965bf4477544c5a0cc196c166f05a72d086b762c772cf02912769ea68bede7bd9d17f2a8f0cec7
zc067d0776f600d89b3c678f534fdb9fe579cb7a128c14ff0657ea6028c05691438a72a2c16d4c6
z30d3e2e818df6b03d36de12f9846730b7f9863430fd75b59b60e56541cb6351c576794ea52ba65
zb1aeea37925360dd8d724056aed7cba9af871e4a6a140136e693c4e5793ef5cd753c0a2e68ad05
zd6d20c2d9e29e88a7748054cc7bacf20d523cc64a7fda1e2b64f2ae8ff31edfd9dc2da94c60c37
z256d5305903289d7452b557bee7a5a5fad443d082e2b275314ea9029ef850247c1ac325632392c
z61ad971df6c8a11de8ea2a8a99151411ab5a8e096c4d122ea5aac70d15a6eed19051f17059f91a
zd120627132ce67d073ccdeffaa22db19cad86a5b52251f8fbb0951a10c185795a1cbb7719b23f1
z8fdf423cc74f5f39e08820671478e72f93f47c3343bbd7d03dabfab8adc15743857c466d251af5
zf058bd87ef2f7d89e35e03609a2fab75c0298e853177a61ec77fc6444229ea046f83f7dddcdf25
z1f39d51bbda245977f382f81ac5894fafaf92811ed9710983f1c45fbadf2a79da9b02c94df0ae9
z9511340dc8b351a0c727f208515fe9d4c08d8c13b785324a7bae73146bc3a1e19260b39add12be
z2af66c1042f6ed3fe86e76fb3efb463c581e3efe6496e646523604c460a3f8776f3437edff0833
z968ea9f4098b553dfc66f37e3bccc33a4d21ee7496152fb8d6c6a2a3fbe3811724fadd1af13b97
z30cd281277e60fda66e3231a88b8b4a8a000e8b0b49ecb77bc15b781a91f35a9c5c4876b7d0314
zc106d4a8fff9d8b4ca047e8a73e7fdb06e0c70961d35ff14a4b7ecd408dec6c97e565d351f01b9
z55312566ffee8380a53ad0a747d3090594cae522dc57d96b6998710fa54cfd5aaad08b65dede8c
z7ef02323115a3d9602062a4693eadb9b1e9d8e5cd53f017551d7ede9671b61744169ad68c2fe2c
z38a085397c062d6ad29003bb96442d675d7bffe6ab48f87f341437700501323c0bb37b1437e096
za7a1b76cc9ec80459835bfd55d832ad64a82ec2740271ab84ba1931cf9d3385567981afe5b4184
z63497805d122c31529aff1a402b4b661103e402142facc51a40b30ba8ea6d7340b71a8d5439a50
z369b45427dcb78a6d6c8e19802b484d1d934b63bcaa20ed8baa1bea0dd8be30951ffdf14af7b78
z527c6b5bdb9daf3fb8d0641683480ede3a227c6f08498c3617fdced39bb9f7a667e5dd2b89e82f
za50a5fe3b08b50cd197cc1b5ae2c4216ae2324dde375dac1dead33d1bab37bb1f2d2eaadcb0370
z3dffc32916453466662e478bdcdef6d08a866716f834f3d9f18ee1a648b484910b1e9d0748e1e6
zd4a2acc05209b804e0ceb8ad7afe2f74b3ba0b82da32f53f2bc2631c22f678f30e1e8d1583ac70
z17282f557e1ed2e1952e9878093739511c7d7091fbb95790241faa673ee7f2c3b7f2117cfadb02
zbb996a904fce9d16537fe7ef2c7f99f75f2c0f91e5ff17e382d70becccdf20800b9995086720d0
ze007777f386571f0ef1ee236c847f7d3fc3fb9541488367a522db5325c0f8a7cbdb841fc473ec0
zaaa87085f11c9ecdd7b4be988368430350ccc5935ef1d6936e0b446a3bb36e2ad9982c06423de9
zaa5a02b1514b42c4a19a22fcb34b6e2706604c218082ca7a4653db7c03812781864abe92e7ccf1
ze613e27f64ebe8a686a1bae0bd7dcd1c417320ba06145eede22f8a59ce41d16959abe9d47ebec6
ze7ec005d17877ecb358481038509ad299e2dc9f1694a9b014a7dcd837638ef8742aca4204255c6
z87e2ee03d90cf677e678f296bf98d8b51036c447b468fa79959c7d5054478fbcfa46c6babbffe4
z244b4d30abe904cc8644c917721c2b99338a12bc7d24f57d2df9ef8b390760d892d93e3869f517
z98b2f52625bc7d3e6dffb7e751d45ddf4efbf28f336110445e35dae6569cd82031fb0ff89e8252
z996f8d639c792bb630b2dca99039faa851dff840511d4a9cb59e9cf919afaa6858d6e408193b7e
zab6229e69e1962b54f088d9ed148e50054c8feefaedefe805745e26a49ac509bfd193882378aa0
zd4aa3994c34aeeb7cfae0d888b77326da277cbf9d399f9424fe23bd9723066b32f529de0cd95ca
z3ce591b55455cead2d5eef6f83b6b553ff1c0fe5538aed2c65c73b3fe2d429e5623589eb93ffb7
zb225bca7e1f3a5a0fc5c758f4abcfefd2607785b60ffc1c90ddec7b425a4f748a92a714da4a268
ze7db264ae78074f79d25141695bd7adbb820ea964e34025c02aef535c0ae954aa98af3315c28ce
z8183aae74ac60aeac2d9db1d1867ea6df38c5e2fcf96aab8ae7e861347f85271621b7ae03c373a
z5b0fc29a5c153594a0ab189f76d8905f19fce77206b6c65ac465daca4d67d309ed16a074395792
z569c1e78865022a600b16dd96c391c4ad07f2d31749ebcbfdc1f5c08f1f23fbffbc50f19fe970d
z7fe907c646721d1d40fd540825483e5128ab7a29ec8a98e80e3e34100bd0c62dca2e9e33d17988
z785f46c2fd052732e272263957262c049370ad67840d40ad0fd897a94ddd2c9a59538e0144a7f2
z96f84c5e81c865b9c715b284febfb3de38246970ad036ca0cc1572db2a83eb0fec81d6e0299bde
zffd67675e6257a2b04f446d66bff5fb443a29ce6b599ff861575c0e4852b2710d1fac5f69a6187
z33d5e54d3a33de71a20bc232194ff9e74e75c176d46220541ea98ca2221e125834cc19af9f36b2
z0a75e5fdf2a9575b0318e7d4265ef207c83413f9a369c5379e625dc54d98c7ac92be40db3968af
ze4d79a9b91446093932b9d6350db3c2465c86f720a320d8a33cc0caa3f13263764e4d1792e5d80
zb1c27dc2866f937a6f946a07644198a4a37fe99a47fd0aad78ced7dd8899bd1012bd99c6f14b74
ze30ce09ee2e4c567860653254b0c732115a30770ccfd160950d156e872975aa7b77061391c0418
z689a6670665ae0c4768dfb1f42f0f794a6162d961f1312a706587a3e1287a476937701baed5efe
z7927cb9a4daea2a9863a635fef1e0c83568836ef26eb9f74ca39216829db9a26636c240e3791bf
z2d2b8a26e7b36851f50d95ea27ed5dfed9b748f711fcee16c32e1c4f0c0269fa778bf494f00195
z12bfb18fc104ccd0593165b63a246eefd484df2e9427f97c03c8599418ca5f47c1761b49177467
ze89d939fcb8e6d0181eae919ab3e357031067191de449956748890e4caf0a5bb60c0de1c89efa7
z04b9a0449eea4b7071572cd44a947e814895c2905c5a776499e9ee67c57fa962e64f5973c56847
zadfc1ed0a050557c26fff149a48c8c3a8636ce9e51ab3512c994b2497cb4b1db20b8914f60655e
zb6996d549423f86792540f58e9894ddb4c47f2d56776fa021efc441e0a196a194e4df384f4333b
ze2d3abfd5b3c1b12a56bb7a4f52622c304f4f2367e720983f080e5f6d213c7ba494d5ab5f907da
z2ccde891b5a713b0fff249f079d9cd97de0faf22bd876129ede3178b1725e99b1ab793c6a86ac1
ze7f89997af314d445d593c2aa136cfe91d614d10f80093d6583c415c137ca6853504f9187b62fb
z9cab1e250070556979067d7e9c24e8db4d7248701b92b0e566e822460e14e0e3aa47acea0a98f4
z12c45100f47024f74034566ed954188eff2b4a927ade06693d9ae0fc107fda1f18b91a7aa6de7d
zef6f77117dc3e6c8507a03747d53aafd9a783ec3dd762504d2660506ce0cc7131302c115e94567
zc05a3cefee199893c3b1ce78316ba9b8fe292282dfacf40cb74e5f7044356dafcaa77bb8a08a39
zd14a023c7892124edd556a1bd09c3cff7b0612fc1a09a40c1cbf40aab4a9768a31b8597cd045f6
ze971d542259e6f1a906fadc807ac69d5676a04cf739448b52bae16be26043607cd64486a9ae9ab
zfec942fb515b9832c5cc8433bbfc72044b78b39f14a7afbe104271cfcb93bcb3be2b134f5f6523
zfd278cd6b34a7e8cbbe09f7e4ab85c541c45557674da1e39a779babb36d36d1321b95149ae52c2
zbf9d918083a03bdda14ceb113ae13e32fe61f543d321f40bd4c827e5e47261e53e19133409fe9f
z57e7e3bc50fa82a34013e9272da50150bde2ce49dffb420064c4426c13dfc2a40959e9a5fdf2fe
z5b254bdb92af3d8a85451efb611edf8707a697b9a9237a38955541748c8fe12a198d5c78393fdd
z1666b8e96bf868721307d0ed6af0d2c33b455325c24105261f65365fa30e0c27cdb04d06231670
zfa267e3519af5a6ce8425785689ce4db9f77f7148ba27254cdcba6118abbbb2cf2545e6ff36711
zffb20c6899b40bf0e09115d65e9fb99222c119582aab1770ad4f45269783e3b3ac6656f471ca5e
zd56978766000e14351e3c93b134448ff5f4b97943d13ff424ed98de39ba3e8861e3fbc5bd51117
zd127d3f9be32d52c37b28c6d69684562491dcbfb5fc3e1d1f76d353d3d50c9b84cf7aa492d9733
z5bab4feccc665f646ad51cfd884b4697f261553a80f1849b518d680d87de980cff0fb25bb79c75
zb1bbc4ae05ddb4c539dae39631396883b817ec863727fd04ea119fae3ba642c745d04e8acaad20
z52728a737af5bdee218b485ab12c22109c983a4f506af91ce13278aa6c750862243e1d51466e0e
z5858851c30505d79cf889fed930b6d4c3a5dc269aa9ce7f7555ca53d2b599f31d31bb4c8eeba85
zabc39fd12a11da8f0c2e56e1cc1338b54c47632ea7ba29642287ba745e38db09f977dda6343818
z39f81da928f09f5354cb1380c7de42732e0aa37c5ef650a11c1d54094002b494445510daa8a2d4
zc7bb5c1d47d50e016ab94c0886dc08318c1c184fa2217f26a11ccf2fd3d207c5434238e2dd2b72
zad1f5fcc28267bf9eabb16ea1a0ce11777afc3f16d7e0f340e0bb7f7756e6a4b50e3db2363dca0
zf2fff6c55af2c0d90bde1b761318212daf16004f2d95ba52a17ab81287b0cf8c3dae7bdac5bee0
z96340581f04a751625d98a151401c5c24ba1abdd8f4f3e7850e2fd5fcc24106664cbe7e4998765
z0f7bacc22013aba4c47d6143f6993085408181b30347573c2c99e110a53e43da353d41e694dfb8
zdd1b3e248b7cdab06c33c66d01acc98140604111038fa51a3b9dc0f306b72dbb48064aa764bce1
zf84d47c8e15426aec3ad50b5b360eafd5cb328fd6e0e56390a08933eb6f4879b1bd6c43bb4292f
z416bc418cd684d228db7acd3c76af2e8a9e50beb97cbd70296fa77dd120bc3e67edbe5b69170e1
z26491430523388993d64accff3b5ef2e17a7da6c7cffaa81d13f935d115bcfb2fefe9a37f2f896
zac460ad7e8ef85a1b17e39b6b1fa425f25aa03d30f7d3e17e1ecf49abca8884b789d99a6e0f592
zc7adad3fbbd1f2c965395cb920773798ada2081b363fc494252f75626e906961bf7576822f9d2a
z6f34a2d8dad684036d339ad22522e087987ad686db6706462358ff13a0603600bee3bef1bfe3ad
ze88a171903216307fecdcd3b56d58aa4ac3ec1fd51a8cb54e013c5fbf42855b960a9f1acbf00c6
zf77889d33f3c9445c35bd0e892fcf5ddeada7e2147e4ab2f62df2b6d503f52b63714fb3fc52f3b
zd592b85bb3836ca281b5afa7a164bdcac193d8674f8f00338b46ad55e227fe7ae52c530933a185
zae6e176d73ba121517fd9a7608e8be7e8fd19ed714a1064a6640a330a5dc56bbcf1473446bcc84
zbb394b7ebf7fdc9438841b4bdf83a110fbd5c5352ac2aa20f22e3a2930379cd27ee8b0768dd80c
z48d7d9842598d1811c6faf41812067a1e3457cc65cb03d9a19daf2033e4f431d6369ad645a3b8b
z4de42f2d6754c53fc025eb175bae4d1f74a607da5fa9f191910d6441b236c391b72746cb298d16
z9f5ca178d6efa4e342eece958fa4c949a32e8879bb57d58b8b4ce2d76cc0ad5ad6346f94863178
z559723a461f60bb00c8c5e14e2e585e0caeaf780e86429c4ca73fc81d4508f72a040d149667033
zfd0fa0090c9afdd5f9b5e0cabdb70855e9b9d640b42214d3f69ba8cdff32fcc8b05b9bde4d5b36
zb9e7e8dd27adf646445ff7de162b91d5d686c6086240bfb8621eb72ed438be410b0cc3732f11fd
z80c2065fd1de36e7d805774c4e4745f8161936d7e27f54d33c229eba6ed24d77d55bc23d15ac65
ze4168302e4425731a9c57616b6d92075f1dea95e3c8c6a3fa868f911dcbf8e628904df32800266
z1ee8ca005b61c60f856f6562b0c766e2c2a4dd4e754c5a9b0f4a08df33e5e95600857f8c4a5a92
zc61cfda6f3528840b3c825465d5278e3858fba153f4fc40e5d013580501bd8ac215ae1f8f1685d
zb1b0426123d0e0764322f30009a1e21e5c3e2274697ca274619373e9cd73cf10ba64d88cfc9514
z0b9da9f48afbd2d9a04ad65a68a2ac8692417dc55fbdcee5c91c3d5b95b9ca1c91a0dd78ad78a0
z862158b1965a036be4dd59a483ec4c7643a27ee6bd96e431b0f8abbc654cff4e196fe66d55f2bd
z0722a65788097ad8b129579c2e69afcbfa429f229fb03e29b50e70cd60379cb36174e51c1481cc
zeac07a0bbba486273f1a03fb020a911b969e0020bcb2aef2cbb3dc4879575fba1cf14f928b00dd
z691430e6c7ff6c80a8f7f3fbf527b69caa23f571ce6dd0cdc6966adf9a0b68e53e9906fab76afe
zc73cfce22b71bccea88767405fa0053654519859ca343586a40978061db501cb792a7b15d8e380
z2562de3146dc2713dc9967356bd992d8692db31bea6ff8c077f885283d8237ee480bfaaf55e66a
zf24b72a0a1ad74bbc7c580d7d7000ed86daf6d688b5441fbd47e9e170b26c826f76897d232a4a2
z7d3edd720d5704ecf00931d5dc2fbf5ebc89ad5bad596ca39039974c1fad579309056bf07678bc
zf81b7ebe079ab212226a31d956bf0b18261accf2f798645fa62a2a2efd4c5617124c323f5a9013
z18b9dfd7daf6e61c4710ccae6c19b09401c06b969214f4638179ba0a44050ba820d6efadf2810b
zee0d4038dfde92834fb9eddb8361e8e771df18a8e34d206c15ee98c9d576bb0c1a9b7ec62fa950
z5e18873ea7f745f75e1c86393f6594a630861ca8883ec600b78662f688f37e824eb6dfa6885cd2
z0b57c49e25ff84e9f32f8af0696c25cbd948ff8b697d3b0a36c9d2a61554a106cc0413123da033
z630d95d1fc2c892ccfd75285d523375bba2b07e92e6f2f29e8d0cba52b20ca0e488ed2a4f25ea8
zeee3500a631df461ed8456efa836e0a1b73d2fc594df4cd35a6fdf865e05b8d67d9cf603f918de
z7c6da263803d7141135eaf7e4f7a2fcce852c94204e47a06fb0d3d5a8bf0a4f8a4cab41a612ce1
z5d702d06e59cb90e995cee20dbeb5e9b4d33f3e8e556fcb83b33c0250c04c61719c16fa0bb031f
z4a5309bc3048008f31770bfac588ee0c2a34e57260a87fc7c765f2336cf545b7b8b07bf29ed666
z9c3578d89c2ebe0abd06b5bed0bbc385ffa76d16e7860311e88c9cd33bbec92d2ad5a6058300fe
z05a5e44de22ddd3141d683bd9a37a2c96a18efe00e7ed6b73e79f68beeaa809c6f64b1e53c9593
zc715653f128646088f866a1f119ba79e0fe404c1bb3fbafd432a778927a3c2346d217e9840fa2b
z80495f75b4dfe2d10bf0ddd0e96e3d85a0354b4ac67ea344a5d9a2b8e4ab7b1c26482e9f21fa75
z388a3a062aaae0b26415190e7c1b0213c737208b79ab63749107af8c4616e1033ee8b59fbcfe41
za59d91915662615f8d06b499540d67753d547397fa3bc5cdbab750e9d3e5b2c65c740ee0caf36c
zc2b6e8acfaf2717f7ae60181d0e514308551a10422bb57cb87f1c6ce8873f63cae06cbb0e76399
ze4be9d8cd7c5c5546909c912de6d2b337e513f04805efd8decc70c89dde1bb3f61b9e31048cb79
z775c35a9c5826e7fdc1e1df13bbb4161dd7d107723988a1b5f273db34448f89977b6c3a7de729e
ze0769ecebf410ba333624bffdb9e026eeb339881786e566c36613429958f8a6b6681b662b126a7
z0ad09b0dfe2111aedce78b2dd6b29f0f9e203ef26983adcafaeed5d77eebd09d14f01a5a05b114
z5141fc2f559d1b277a4aecc3ecabf81de3feb77d616cca35f33c5aee9252d689a4d4919e9a9c9f
z876ecf0dc5cbececc5068d5fe4601523ffabd860ffd75efe7711d53380689ae1acdbdd503d0e8f
z070d4f7a49ddbf92a7ceb7d610abf8a303e09ea42583361be00c44282662b076fb8fc85fe95120
zb7955ba2ab0f75e883ea6fb807554a432d897d8a2fd9f1432734fe77f432daa094d46657cd1168
zedf4421ce926d1284fa18eb2c33018f0eaa345da2fbd4db3101c791b464ea477b64ab546c9dcc7
zfbc95ff326a68b6848a36d1ac54b189c0dfb1a46e3cf565285ebf8df389faebaccdffc61cbf4ea
z0f2536f4f55fb312289efe75715a7dcda523fd45936c401caf6b97c0430ea03294755d3ed45d45
z8dd617e9fd7dbe931d1b3fd0204cd8d7be4b61c2cf398d0e9e1dfb7dc785eb1f08a632ae9bd9c5
z9f20533222e0b6b69b3e97d7a8f3ea9fb7ae72317d3a67986af6d0622c65fd97b78ad118510050
zc5eb0922a00e1aae9fe59ab194d496ad2f2fd43b8ee951eb3a8025995d510d6846812e054eb448
z374f3d38249bcc7ac197e4a44da23e8d115473e0d97e214c63ea2a9f5350c4cd6efb8bfbb982a7
z2dd1a29f1c22eca2b884c60a89402047035c17bad373f9b3afbfd046500c81dba37e2bc5a5adf9
z5a0ebdd861b2639b0d6d5a180efeec6d57e0516957f0e0f2e2eb2efe43ccf9a82dbadf007d3a9d
ze0b08db01b5b72f2d7d84739379de77657f8caa1f503fd7b54a992ed4f5bac59b7ade10ef5567e
z19107bc012582a5ccf734e6f415cd65e367515b149862a29886958dc5bad9aa525ce352ead2dca
z2c4fd1963aeaac92a2940de0fa7d0029fa428639c47ba5d6705b87fb4bbcf8ad7ed11ec4d7529f
z092f1a30aab0f335f5fc6cd3a9edddbe63e27e15dd3a488270721f268cc118fc3f6289a04933dc
zd16c2e11888a7b8b7d17f5e903c2fe148bbe99bd7251905975985b7f73f9a69645834b0dfb9e9f
z1244742428acfdf1f519c507550fdfd1e54d1515a258629ec43a97fc5ea0aebc064f1ed9b625d1
zb3122a0aba0069ca2c00205c86d2b801cae3f86b4bc48ba9272adce44a35d6581ff03c7608deb1
z2846fa6b45ea11dec673331d6c4113f65b887c09bad5553a501c4bf69a17efe4b2b329b8c16721
z768a85d9b2be1038369db26f88e3857b49bf2f3476899d19a01857ea1ce579dd250f443a564738
zd8460de4490917f32668f2dea2bfd5ac9622133b89f71b986dfbb9ba295a004adcc3886cec83b3
zb3c97a4038baebdeaa65b0f4d2a9d57ad4086afc831934cb20e156a4f860306105cfd58b34a8a6
zfeee3d782f19d858141cfa24aa11930132d36954218027e41e5109e66c16471adc630c3a050f6b
z1b7051f17b63514d191cb5d42c8a6fb6ba3cbeca4c202098baae0587b5b03e279d5e600602128e
ze67114acca342c284a14b1d85303a450d9a3f00c53e9bdf4dce31306e5ebebf44e7d31bec5d80c
z9a6897c92efd833c3c47173bef348a23c4645bafa94b090cbc2b9fe7341a70c210f5486d4ecbb0
zcca37730532fb2944eb14a0eb57352ac52c670dae79d8c05193710db673f4fe1dfc39bafa2f6fb
z1c63b7c80d40b8651398d8441cfb15222081693690b617b8b8e98e1b121ff7141f54a41a97491c
z349b7d52ebe87a11cf2a2209ac8285045cd271b0de87c5e70ca18ecfa51ba39ff5f80cbbde7248
z7e2216b97ff35947d8095d9421f43e51ccd66ee6ded9c418b3d4ee4b78fce353623d0fa45fb22c
zd47d64413d1f9865a92325a7d420eda02aea2c1a6c4216e5365c79efb4faeeb4679da3f073cae2
zb0ca90260d83f796a3247f27d8160bfbb38676c5e0e1363e675e366ebb214d6ff1a26a9bf7652e
z6aeda3edb607bfb7b65e9e6fce48bc8be3da155debede052c878ae4fb7e6f486fbaa09c2f97d86
z6608fe6530798a254b21f5ead51443c9bd71994ce14bb70437d84c60b90b6dee33b4c6f303bc84
z729c95780b2b044a570e1d4deb4888ef463b33f4450dec09644e1a1e0ce7a0f3b5cf13d05b2b9e
z618920dac189e44f4b33f4d0a479d894b27a9540c8d0830ffdebff20039953d5e378257d5bebbf
z923c9bfb639a0d17bbd4d77495e14653e9f2c1ac02167d4b527f00c86804ca3aced7afb2c0e60c
z76bcfd93de2cd38777fcb98adcdd9513b22a7516aade57a7ed6fe0e579f40c5dad86183e72aac0
z58ede0b01b8bb63bab2120797e85c7f90611c2be2bb285aa43b67613de0f1297b1d8bb4c1f62ae
zff61f680f2a27f2f1e09c98a89b6ff739baaf918daef2dda60062abbeca628fe722bcd2f42c65a
z3be623f1c74d0b1d3cc3009299f62caba625d3a9092c7201745bc4900e9eaacc0c849bfe34cc69
ze8a3f473bac881ac1ff3304c25209849b2b98ee92ca1c0f1263091bb3850c43af5dbfcca5a25d4
zac9a261627d9f88dd014de7f5c6a91eecc4c00c5f1625363eb779f7b85af708149696b8cf518e8
zb6fdfdd312781ad4ef7f8c8e384b35b228c2cda6a1277395eba117a303d595b0f631ef00f2555a
z7006a760682553b6f40a50a543aaaed115e5bb61c381899946ba057dd36d35998a6011253095e4
z575c7e02605c4134b7ff38984699522e500dcc29713c582cdfca3b3b9a07ebbf018de49f72ef42
z3f49949e66e91960de1a5aba70e35fc04c1c2bad45bba02c5ad65f716031165324bec809e6fe28
z8a4809b1c1132a41db1a931b106752cc95ff6a3c0c244fd471aeff8755a2deefc5a654fa9b604b
z62f29deed3b21de96f5c416113a09ef83c04f788a082bebecd4032dcc02f5b22a2f4bb743df4b6
za21d6fbe80a68ff2db04d7ec00b1d6103ad29e50713c78a9b6cef3202f9f28eabf63415093cc5b
z486dd5b06af80b1bb8890396b6a2e61bb98396830be7a11e9b51d2b826fb86d35bcfdabfbaf544
z706616900e2578d4686e70ce1fd9bcab46da7763493ea5587886903a539315c51fc43d013d0730
z4e054ec8d701a077ea65e04f789b44a0d2b7d8016d779ba5bb6e918cee30bc2b56a6eb3f55ff0f
z1cb58a199b75ae0198317ec368a42e680cf4d504a0fb1db5648ea15d3354cfc925bfdc5e462d3e
z6ef13d5362f98dfc2ee61a874d6dc4a9d1f4b8845f912b15c79b2c06fa7d87304e088fd7b0458b
z66e78c7f893ce916bfa53f352295daaa2241ea3da38e7c793bad39d40c8558d3728fe4bb854403
z331ded7061200a15216fc8d7f0546372efeadb825f4599b6d9494434af508c3c1a7b345c32107d
zb654be976cc50cd9645baf973cd25d653b6447a1ecff7ae1bb124f0fa8b745d71e35bcf447fdf5
zabf3144c4e98148dd6505c8bcfb291133eb1c19b0fc52e19e8bad36e6388a57039878a3d6e54ca
z3e12f6d0e2f1b55a071805a2b556696c294070621ab1bd0918c0eddc1f4d2daed72b8ff7dffa79
zc3b36c06749c6e25f9017ba1288b5873c2ebfb9c72358d97e56baf97ed381730851945ddd8aa5d
zc94166f3fc62735f422f1f22570754ff12cc85d2349c90536a261e51e50a2c126f42bc8cc07188
z6160304fed183f4ebc50285b1eb69094804aaf4425c67b89d31429d0a19c52e77744d28ae3e4bb
z572de0404ec224c487ef0ab419a891845e4314cb6d86bec2d673b93a7a1d59a5811e37a00935a8
z367204632d0f6a8b0c095a5e24a1cb554c441fa817c92a938ba0b8d40b35cfc982827f6843c29f
zc75a33efe7d3f008433201b71080f58160143f824d5227dd163af6ba9c5be8dee78b996b5363bb
zd6beced16cdce568dd0e3d542542dadd0cbf466f72ffd0d8d1a36910a4b0d3c35acd121921c544
z4fda1ad3b9dec64ec91ae1152a4bb7cd06e3e0fd0a62a79e529ec0bffd03cccc2802468da33258
z7d0a8b70ec28d2727df74aab447e2fda5ff7301908d66b21a5c43a388251f59d9ac43a9c48d742
z84743bbfa056e08e60e75aa6703ef508b2d737bdbaba629cfbab55a1d32cb945ff45f75342ee4f
zfb73f808dc091c5033fa99a0eb241a88b73cbb5ab61dd385287745229d938ff8d797acbe57a938
z871f9e43c8f72f34fee77ed222f96acabeb45adcee376a311f3c18ef6103bca79509ba82e732f6
z99f865b5765c44a4f070277be9a7814f5984462ff436613c7af8a14245ced13c9238847ff7c586
z50e9c9e02c46c7d865f6b9118825a3d0725be317fb521fa95bcf0f5eeecd2f7652e419a67972f2
zc92709c5f07fc19f45051212d6189d57b549be46a38e9bd92731315d4d8f44d9bd7f294b3d2c89
z19c42589b8dcce16094026ea767ad6ff3a6b605a609834f96f25bbb428f310da9e6cd43dd79ddf
z081c7e6189c249abc47b2d1dad7bce3afcf51c12cf5044ca946c6a767a5659e983c46a9153a47a
z22f5c50d60c27a0ef8cf488365e57f1b1aa486ce3c60de0afbb73adfadafa4077666faf8619258
z4fb0d1dd31dd62726fc5fd2d1f54817ad5900a31c1ae4f9be23e9086a3f7d1a458da0b1e54fb11
z91400611c2c1629b7bf69bd95042a0bcebe640684d68dc793cab820ccb87fb9b00ebbdc39fb379
z071a03493187a4a2cefc63f334eb5c91637c4e2192d629946ab14ca39543780d324e5fcd30da6a
zd3ff0746712d9dc5bb1ae2374bab69fd5e0bff535d597ddaca294b5785c4b6fc404a3047e46d2e
z5203dee3da8644f255cad5a6dd9252470e14c9c8044518311164701b3c018e50b4cb9647183daf
z08fd2da0cfaef4d9a3f690ec78121d6bc51aac80d2a100c82102f2d1e9d40377b43fafe77120d2
z7c2697b14ac4118671f174399fd90b878c5dee0c086e1c2510c8ba81801809e7b2339336fc3621
z095a391dd5649b9ba617c67acefaa756d3ba6c8cd2d75d5a9ef0a2d701da5d6b8153079909f96a
z15b92dd3a97aebddcc1bade2bf3c3c98a07c7b1a81afd1322b460389937329cd15fd134628b343
z521c86d875459064f94dd2881882567fd50948e125d8803bce4acc02a3b816d971c70ee6ea26f7
zf4652bff666d875252729b38c76e2687b7a63db57071c955ad6ba583a5855fee67268630a2d66c
z623cbb3fd10698a52a77dfd9a1072e6c8f0c433dfd725eece5acf14c0bfc4c0cccfcef052f32d6
zc4deebf330142cb0ecb7dfa595b4a97b31a925fb509dcb60d12d4e45b0aaddca7d2090c9fcce95
ze45e54f1aedd9c9f57d9c58591e8fc5497b318fcc67dd8f6d5d11ab2a3307c84ab84224975c446
z5ed524942fc3d9442562029ba36be435e8faa3f8a98b332620317cec16bd9aba99cb8345a8a1d3
zb1218bbb745bc23c10f52d0b25c41e5737b539382e74cad54d20affd99d05951aeae5a65f11fdf
z2caf6e8c3bb432d8f422fdd83b12bd3449dbd4b08bdbf78599844037d30f6bb4ca273debad6240
z5e0c66b639a3245214d6324e2b956b1849755c4333d973d2108136700523ab13915a13f2770fcd
zcf47b23d035d091d1d49dab2193e67e9c151baa8d21423787c059adba6cdd9ff8389bffc9a8701
z386a5b9e2db8d7a0b70f01730a0da24408c0b966bb67093edf951919224ff581d8515090d26a76
zbeb4305625539c6ff3bfaabceccdb191806d1719900830eceb2249eb824ffb72fcc99b30aa133e
zfd3cc91df523883080c2ca7a1fc4787eb969dec37bbdd7d6cd76a91ce0446fa224eebd2f5177c8
zbab473e687f6076105c4c99d4279f8216ecaf54bab4e7821a710758878e13836d5f7c16be8c717
ze288f8b1dddad5ec71f9cf5cb037af78d05d7c1c5787f1cd62375ce40c38c1bf52aa5093b78b5a
zed17c0d03b32f8775dd53961c1fa4e4223b0527a5806d16810778b9cf8f389e4fd87f328415f42
z7d5e2505baa841157e089eb8e23071710b44f80d38fefac0abfd905c083e2e6ee02066c47ff59b
zfa8b380f7ccef7cfed4371c5f89e66e2f3e6731953b7354a6c0caf926b78010fb83e5635fbfb9f
zce6807d4852b72de56b4294ebf26164d9f497fb3d29a665cec9a80442309f7d196afbdf169b606
ze621e8b01c51fb5357713f30b4295647f262e820cca6411c6eff3022a2473cb3a5169583175c09
z9d6944fbecdf26e752f28b6b9a1d4e780f7d509b716b6264257a8260f539bbfe72527a1cf5489d
z7412160aa64735f483db67d4df483ae3d361506784662f29b086c56b2a222d7d1e490bae831c64
z56ae5438ee3b5add65673668664e790213dd64bd867dec1524587a4dbd0d01fba343fee7091a78
z74526e07a95d32fa9e18c5cb190c9eed28d48599c6670f4bc6a9036df335984121649f7b6c5247
z92c3d74c643bc77f48b1e75f4adbd11aef1ba067abfda16c9e3012bc9d07eebf8207bcab913f3b
zf97c932f1aa9cc49cbd5e75b45fa0a56775b721d3359a737d49dc14cbcb4934cb44f1bbcabd54c
z1aa43097f052eaac68c80cd0e7c8878a910311ceb15cd16d35904ac62aef81d526bdf7738b29db
zd6ee0135a7a32a3a2623f0e151c7a0fa8871ce2677ade445cf808569585dafd3f8c5eb49427f3d
zc1b621073f461966e712fb143ff76ba6e0cd1c9e6710c10437cfc26b521c1ccb5b6cdf1cf98076
z4349d6f1fbc6384968c1028a097a27e8a048d2734024320b40a99c6bc4e32176557f2fa782ec27
z03bcfea09756e7382f4264ea3f3159e7a8da633c95b87de9dff4f874290c35edcc9887cfa50a5a
za7aba1d2937e4a3335e315c8b125e2c452c475f346bd7610a62cb5a09b0b301caec69c00bdb523
ze28cc6d0679c55d0ea19966ad821d0525b28e784c75644c5b694e54055da45d57a3049d8762507
z280bd2ef402f5661cd69eaea65e248234f85f9ecaff03da3d201f800e53c7ae5eaac59bec83a43
zf41321f643476bc23a4edb4a310f11d88db3cd84a6102e15467cd7e0667acf50b2faa51483c777
z72e737efc6f464b3dbf969bdc31cc267c3d7b753f7d3bfd2b634ac445b09f57679d29658a54f7a
z15f20fa86390e53037b16f8f264dcc624c249d757ba890ab43594a3511b3a46a7ffefd8f9dd736
zb0f0bfb45c1cdf6035eeb8969e16341399cd58f05989b1df8e115dc13f59d2184e5fedb7acb49c
zcd05ab125badea7232e52dc2941ecadc8fb1962100414a331f68e41ecd8431519c98eaf5358109
zbf23feace308c0a4b86f6169e8c78e7ae9702b9bf30e2d38dff35136433523499087d503ce098f
zcd7d111040022845a8ab7bb212bb7dc714b0f90fd1e43cf4f57f2430c059830960a050908609b1
za4b28db33709c78a80729a4bed2b2514cf9230be4d91924b0df30b30e3b18de2fc744cfd23edb2
z32b84b996f8b81510449f3db11931b8ecf7cc22c39935a9eb8e8657a0edbdaaa2006eb67b7640c
z21287755698b23f910eda48b83a4f68246c977368694dc5d3aa26adecd7d8a4475f87623ecfc95
z8f8c9764359ad88687846c06eb742fcd14d90ba7413eb1e7ad4722da3bddacb8c5ed2a3b22a818
z3bc8433e7e6d41ef27e4ad5a0b8f64bc600490fd2a8c4429ccb0944dc041c5b86368f9900640ea
z6c6466841f66bfb319840506c0b3f3d6d03ad997af5ebc24aeab27163f6faf51b7a74bb7412883
z55a8bc4b40fc767372ac80f38c74e0af7f130359ffaab176039ce6483284f8d6013a540bf44a22
zd8dcf8aa4e5f3852de4d4b38d12e81daf4320f89a73aacbe0a4c4b37fbfd31984095ca69cfdcf8
zdda04bfde2192e5415a6b6a2a1b3e246294e506ae9eb47e7ec4863f61eb34eaaed66542b80382f
z5e23de7e0b8e0ceb41dd4e0516d5440a98ab36b64fdb6fe6d76903008a36d5f7b3a64847cc45a1
z35387e737a42417522bf1f1427ee784e8727ff2b7cbd19458a4e3e72781e436fd5ba6528bd1714
z8c1ac87969720f81b9702831b8a31d6259d3ed7afd3b8c6ac0384523332bba10db9357d1a4e834
z3cf1d4a9b158b6f44b9093e090f0e0fa84a451a1ac25c5dbba7772dbf6a6579b1c4d3409f38bc0
z7f5b4f24da802813d8a14f20c0b6142ec03c79dde95657ff3dff287c52f182c330cdc09437e0f6
z90e8ae3351b6fb36e7b333e9579df63361f69c6f726781f6a4f807132ad82c7334ab35121c694e
z5a0fb76665dfeba9033086882ad2ffcf7ba679861fe00cb44f51db56e13d5502a29e321a160865
z323a8428acc9c4841537cdb0765f1d855df256765a724561b53bc5ce4ab405fa7421e5b6bc8426
z66f4d31076350f3f7c92dc739178e26c5b9700c761d3b4ce1641a124a4e80c4b0da41fe2fa22d6
zcc131c9679678e856640bfcc111e8cbcee112c4551e01c17f86647d62a27886bca12e196e4f4e4
z62c2988f65ad8cc27660ad52ad49da9a3c494b45ea00c33f861d38980160c4e0cd0211bc2902c6
z2e034216e492be142f1eff8f0298f58c4e9138eb6b1e1d49a35a218feb035b27327ce79fc980f2
z534f3b09e3fd31cf9c97b43117888e7e64033a12988c94deb6606b6251751e085f04e8897d0335
z2dfa143149f365b07cb78b4359271ca86d4d1a24ca7e67dc920c45384254a715c10e6247b6fb28
z3d3e6570097c02bb0dcd917f53106c4dc68229b11847c0e976364f544bcc9486e33036341e1a06
z806c61b8ecd2738fbc8e83d7ea2f7b1f54a07db9e768206f3bc3f7d63699ef5a772d89bb3abd1a
z26c8ab96f4721b81ea30c73b451a82548b46057589536a95c15f1617d3d82562a0e761f9818043
z427a2627f39fb5547b98e019d5345d00a32874977aea79366d5819a7d81789f5ceda0faecb232f
ze8b95be96beb68328aac9da0c412db8111417b6e2cdd8b63ec63a8c4ca499312f05116443143ad
z06b37d60c5e60a90bc534d4f501d7603082085e58bc6739599cd36a1d695bcf19f6358aa020558
z09737dccd29dd0014f203a4f822890c82cd3b5e714d177fa9de554505bed8c3f865485aa8001f0
z90ca0c6ee5fc70323faed16f9400598677894359257d665add26b30f90e2efb94b9ce38ec57d24
zee57350892b8cc3cc0cf208f8132c972193a6e35ee6b2e1f8d6782df073646ae762afce8abb058
zd7009f87764ca1d32074dd4160b0f29c8db05549dcf68c138e2b21a6b7a9301347205e233c7b84
z85eb7caf1e152c40973e18727b6778a35deadfcd9c4a5e88065a41afee81f8310136812d7ee052
z9fd995aa6402047f10edb1e93328ec47e39a0ca77f2c42dbdec2a8dcdd7b3051b8dcf431289b41
zba8f59b6273bb7172d34c4b7a07e3727feb1271abb0a02d6f3ec6f2319946a103a40dffde8c6b0
zcd660b36925ed95959387d0d6e0bbf97f5e3a64ac8fd21d6512742b7c083697a937126e78208d4
z1798bdb21b61bd2a1c4a370b05a01a2ad98e56d75e10bf5d2a55e98aef756c90c0cbc62c3b75e0
zfe5921d917e7331873084ff5d2adc26d44c17f800c62b6c701883289a7752ca0b1d7fc843700d5
z691e0fc3f8458d8134e78e6f0127cb39ed397ef1d56703c86a09fed836f75427e0c7a0bc4dd0a4
z80273cbdfc2ac1c060a72ebe6e8795312d16b4332edbc91619159276db807a0b741940d49d8f38
z046db6254424467483e262b725ba793297f4ed7eecd3a98217bb6b335756a5d6a4adba060832d7
zb963436bbdd761b762ad28418d81c3ed999f0ba9905b301272e209da28f57f6e2b9c9a90c3248e
zf466a1cf23c47fc4aea7f6185cc597d0b707de6a9fa568d95b73959fa7e8ba3e1d489d6e03c4fb
z0d93b9597be5f49e025275b6280590f103cbc50d219bfa1bc4b1009e4bee3efec35291bc4a8d39
z01c48025745f2dd6242074b4c0bc84556ad71101c233922d86d2b442df99ba6d4cb18d76551e2d
zb2485a6ba585066a99eed1668e39c98f69b4332255bd496a7dbde5df88ec6125c192c5fcbaefd9
z9a4d52dda4844cb2811b609cbdc4084ed5bcc7780c5b955e9c5972bdf3ec42a64bb2e0f4afda82
ze9f3237ab6d2fe6f4b2c62fec3133dd1710793ff766c26639a0b8f2aaaa646d4d87057f24f44c9
zdcdb8e61fd70832da93e5a08628d4cd0383cd044b9d359bbf6ba5828bbc08f53063f9cdd9374ce
zc9cb1ede229f631735b6b3cc4343a76901364dd36d610d86508b429e0c6a7834648b769ac10942
z7abdd64d806a1850b6c449adc0528080905b06c5675aef4c634906cf777604b2888a7e8ee470a2
z02584512f98253691f80f19a4611e957eafae5f4c0b7f71ecf641feed7fe99da80633a986679e0
z1179e8a3c5fdf8af06336992cda9ecd0e78046c7e9ed802cd1b145bc0cb6c48c36f5e59c63a0d6
z1db052285a92c03b49c254d4d88eb64407947ad9c393ec559eafb093eff6955f8322bde576c7f9
zd04a187d7dc8c534e86e5fc4e12fd7348599d2eaf6434d73133d9a7c94da98f440016a7c659e94
z804dd5993b8585719f1df42c4b3317e55530f29e72a8c1b0059c8ebc35f1de6983a2209f445ffc
z402286e4e22fa972d571ebc345fc4f39e1d0463418525612dc3caab2fc891ef18041b976064fa7
z2505da711991e7e6847da84df9b359daeafe13be4608aed6b4801c2614702c3cf28040e4aa8e96
z49a7d60da7fb9c1d82bfdfe2477e548d7c0ea400639fd1f4f336d861f8d3fce052987657616640
zfc6af5324d18113e05d2237a777c652b622a08ca1c12db23af258554f9679b214241d6075e75e4
z08d277bb82debd1350372de661c6a4078ad1cca784cf78b2acef3b0b9cb567934d36f285dc80c8
zc2dc3fa8a437f2124a3f5a7922b2c3f5d3a305e596a553bb81ec79ce93174368c4bdabd10395b7
z39966265d3698f9476d72818c088085407d41d737a2c6321e49f3b3a06cbf8b996090994435629
z22ac882b301f8689de2c6544afe29b41b425f580e052548eade9e6bb83206a4165df6bde9dc83f
zd0ecc24776f846fc94a8e4c60d714e0b59aac525a84b202c1955cc67273130ebdffa46728d7411
z2002b098d743a0305432f4c27f0b44e1f1d72cea3fab6768e80ad126d0f32d067cfeb1cfd8f5f1
z234b0e0dbd5d52caccc844af5fb69212aa47f528128fb204a29bcfe5de3c838d74e4c379af752c
zbff1660b357fab52883b541bbc86c4e5093ca88cdb86d6ac05b74668f685f6ec958f3e0ea5828b
z0901f56369f229e048b5bd5d93c89743e5824556bd0840b9bd1f6010e720785427d3b4127c355c
z597a3f382e6bc8d06d0bac54870b81ce4be765228bebe29708bb0ff3d0565eb8234040b33ca95f
zdb2296f66f162d101a093bfdb8870f03b5d5e7d1d32e3e3a3021b51d61b006e4b8544bb54c6108
zd461a6b87531d6c9ad31b996f2b5ab8c00fa2665757408a29e623a8a0cf67b9b5c582d60bad01e
z434940d6c123d40bd5eee5b42df11415c3d430affae9ccc12501a00e452ef990ef4aa8a0cc295d
zdfe2d8daf863bfb07b96eb2d9e062f75dfa7c1fda0a8444ea7850fa0dc9f5017a7c9703bce5bba
z89e1ea2ed1298d0e37c51504f58cf637728455a6349ffa7d5a7e161e0d0356b784f7fec4735807
z541b07a6e21b24d09919733008c6fc801425e048d0aee62fb9514928ade84006d6da28ea1d31e7
z75b27018dac1f362f2866479051cf13533d1727f6a66540a6af654650dd4091ad923741508a152
z9a1575d495b509295f7eb733dfaa50c8f535bf6e86be8016e3db9f0819736e51b662bc82e41c5f
zba17a7dd97e4851be6400e73d2df48631133478a448d45c048922fec0475edcd1654c8b5d1cabc
z5cc33c9c729da565c3b5824c0f29effaeba2b9732aa82cceda893189b43c3e08da4359c0f99841
z6227ba6cf6d25eecaf62f6d714676dea85efb92132294ece3ffab65b62b6d5e63f97ed7bc1f7c4
z63392f73d97def12a68f7f6a10ed30479486d348fdab487640aad3848ff95ff9e15cc62e3f61fe
z2643f1cbe57427dd084854f866c7abc27164380515012a686644829fefc36bac8bd2acf0839a3f
zdc661c0d02b3e0d1e4af634ad3a2d4435d3aaa59272e02e99eee0c2bb3eca9f4a8dadf8b3414aa
z403101bfeb3f3916425efd1da08193ab5e57a6be693388ee25d77902bfa5f570f9efc548671cb4
zaffa4cf3297f073a2b5014dc5df9f403d5b50429ee2a25fb2528e014be1340165551c2cff9283e
z06761a6b5d99dacad76d55407a7b2e9b6ad6bae5d5f926ec35295a6d8506466c87d4d3e8f2723b
z3d13ffbb95eb6d3ef58fc50cf5f4fb476cea1c7ffee344afadd651672552d5a42e74be8de868b3
z7fa8973246139584a54508bc963d5b54e30cbf0bc0e8012c04804eeb08ff7d7a51342627fe644f
z45716797f336e8298be46b91c84efe138f4f81912231d5087cdcab3ee6440b50180579e792e3d4
zdba809211a7169516e36e17f87beac8bf7df1ff8dcbc93eaee684a0355f3f4da9642c6bb956233
z2f56e906164ceb1cd66439cda212f3a3d8a3d36fbbc68f17ba239fde2987a0e3c50ee148c5f1aa
z31004790ef26b25325fa3c32767f1c165f6571e1d2508b15c7f3cd9a2a489820632f7675c77651
z7ab1fc1774a21fc6464f8987b07d10d1de7b340055ab49a29221cc841229c8649da004c9b3db39
zcb9b1158c3b1e90f358df81efe4cec9be78785b272e12cbc06ca6c0e6e22ecc43d3d140eedaf01
z7378e62427e2379ec21a7e11b5a2a2ecb93d098be6410e5664ddd5ba9636154578065f8d4e945f
z3e5e65168a8f7b920eadaf80eedfd8afd73e3d3f0b8bcda0c86ad1615bd833e313055af7eb0aac
z925b4e80737f880f144f2ea92d7a0055a324d6d1a8f6ba5df7d23a9b1d9907330e2eddf5b9e209
z5991795beb55c138a47b168503c40805ac3007a99da7e52a0c971f5442b5024a4d40a25ad35501
z374c8b774f8abc01d77c2e7d13f5fba913b62aa3ccdf6d08537c95eee4120409c9d4003ebbe6ee
ze16113505f05d05179bac64226a89ca51d73481de0d6ce4341f95bfcb156689cb6b72cac321456
z3e65c3c8e95527c00acc210655d8f7a3ae6e92ede12048f3940b7018f561317a534e4b3d5ea5bd
z2a1f099570ae28bc878d8142bb4339617682d15465f8ba9b6e4f9fd26494422550c781cb4be829
z3ef4594b693fbee26d6bb376bbf6880e3f3da2531dd269d10f32905da4ac755a19c018f7bdd6ce
z6a0f84cc3a84fec1979340ed5da1c9f04c0d195df610ef03be5ad6bb7edfc98c5e6dca1da8312d
z7524f8e319c1fada149dff74ec52d924ef4dd4439590d82f44fd450e1af61aaa96ca75df38d100
zd973c33308dcf0332b4ac14d80e23d28f3dbaba141f5ab288c758a516479bf4803d6aebae29afc
z33d8c16396d7edd73de3a4f966a2916b463509e56f1c71049dfe4cccd159dd9428c05fad56efd3
za9e97925fe06b4be6423ba3cd84d102bcfe3fede49fb256988775429d95be9c6b90e7e89d924d6
zd33efcd963a114a2a4c1f09cf099012b50276d34ed431ac2621ce688f72e107420bd5e72615175
z4c0e0a2cedae010bee789fd6fe3d83bc53ffc21a8f7c10b7351e4d344030e66c1123a2e270f7ae
z0ab9d6e098d0877941c44d6e855796996dc2882c3710e89088431cd7d2033c73904289859ba398
za5f2fbe68c4d71550b662b17825bad1fe7982561d36aee84e9310cc18ec1eead22229d872bc5bc
z2cf7b935ac2f7008f1c437c25be902db8b57f93f04e6ee1a34a5dfa1930d47ecaa8db106a925ca
z1bb88e734ee29e5842b04d19453219d5132ee3e7ba9189c99bb8bfd5280d7221c940dd636262ee
z64a545b1ed14671b0710fe416c985f33173e403e352892096b1f05dcf4905cf38996d39476a34d
z773a18862585248e483afc277711d587b88b0cb45f43b3e76d3913105edae29cce916b6970158b
z3af4a2ef48fa3b6b20915bdb2470f05d2882d4df72dbe8edbf14f98fa6398936e7ffd19cd705ea
za9b2cde0cbf7f8be9c63e33941ec597f1f72c1a2798428982682dd3874f11ac348080189e5e409
z411bb94f1a97d8e59de51ea6b7fa8e4956ee934c517a3acc81505e64edddabccd877e462007608
zb129bdda222f5949be7f5c2ca7ff3a001eeed4ea3b1b3d94707f5dcd859c5c917de7cdb6b66f77
za2570c8f1c4df06830958c2b96ade6f8ac7f1f951e401b09f46904b5df45adc6036be6a5446ed7
z3ac60e975c7f93d7e76481e014df6eecb960d61924f45e535318a2d40cd1cca1665dde535739cc
zd130897f8537f9f3f91a42848ba019b0734649d0952b8a0f787136b92f9b28510f64ba4a78fec3
zddf3d4fa61bd05d33ed8c7126521fb2f0568494313f24e4a4ce4bd9978db5c472931b5f9fbdd6a
zaaa5f3550b7aece835082d2cd803923b88984bf13dac1cbc6de6672dc83cb5a793a7ba8adfa78d
z34d85616e7b409d68b88c5f71dc91d6732e64cde375a5e092f00d1940535ddcf803710b3b67ede
z6897ae2dd3f1ae41d2a7f2e5c98d241f31b03a932b7506a41dc74f4be0ca25d5616f11ae25c949
zebe21f689270a839b708358c4b236f499fc6dd31891573c95483bd9349cf391b001c37f38182b7
z84f5ac5e87e87f747eec88a5096ff6183fbd31b0cf8618a2dc2b3e9a1e434a41a8e51afcf4ed99
zbf87158bdac02205242901e6a99a9da1a1307a868d4fbe91ebca4b1d1cbabd75eaf529d62d09ca
z43a03509e8527276913528143325d3a71e9ab7287bdf8073ea274a42a854fb2e13e644364489c1
z7766bc8f148e0d3d43dbdb4ab22f2e974528cb78a4ff65d25072963b668852fa693911b8b76949
z6201214a651f5a7a5926f5112124e80bfd179f46aa80b27939dc5e2eea8107fea574b9530301f1
z433b7b6b557a2f1f2671bcaf58945af9daa56c2c720bc500e3fe972185b2455fce04dab5f50586
z253dd7786aafe7117b51a1b9fd1dddc52b4257e1c7ceeb117979684393b140f546d34ae9b337ea
za52245bf1a49bd90a99713b9345c958ffd8a0255547d4bb9b7faaec4549f84248d20530b51cd34
z010c6226cf57ef74ad9c374da77e0f1a7c500f1576baecf1363c7a120b086f32e3c498b348b2ed
z7089bbcc812b464868ea0fb2745c01f6e62aac158b72c0052b2087b85192c758c3a8f3dd1b7779
zde1b3fadd7677ac09b27f4184f68babbacf21de51cd56039cf89cd348942eea41bb20ccf4ca6f4
z9ee528319b9fe920b97c77489c73aef7f23dff3d8b763937f4077205834b710686f4483f29e3b6
zf2a8fc1ed46ff3f654f987c7f8d9b82c59474f99a5176b9cc19894aa1ea2a88ad26a30a5f6f180
zc847498a6538ec69d46e3c093d6b8a06c4d56830755e5206f279f64752ad856b24d93b33503548
z9d6ba9b22239eabe95a45f0006e8f0cce553e1fecd213629672379c687bad1a6cb4f2620278a75
za30da93a1ec6277a5bd9211e96f5c161d8ebf2fedc4a0ad23d9507a93ac7f849106ffb11e51c8b
z6c55b3971ef0b02b4157ef0db82c09cb7d66f23e88f856fe69a18c5b194890f578199e880810e1
z0327f9a07a8ac5475456392de36a9588afce55622de6c17aef413eb846b0b438b29fecae84a9e6
zc05423f2b6fe4e601fa98733abee42068a6a4344d5760081c40aef567615f026a4e7ad5cb8f479
z0e039a262c7be357eb885bd662f562a18f320671acac08aae27756c174f9ee44214d656e1f604a
z13d548e48499e55fcab61a1db9efbfeb5da425940012c950e0fc5f658c30072009f6ff877b0e75
z712ea7cb4d3aae1af6603dae8fa44f39ee829a6f852a554e10d4726411e3f862e885e47e62df2e
z04f757c0ad1a09b2a07344fca1ff771c4430cb0cedc4a44932bd18eb83c5e4f36de150abd62d23
z6bba7324c32fb420dab9ea29cf7ea7796a2b89a7ae8af95d523bc0e6bcd95757d06b37d98f7ce5
z282c777a029a9927ac6f6eaf7eabe55245910e56d01934c59d0c3c9002c397e0085752274a0898
z445975e8a84a53004dc046de5103b3b03565d15aca8932b2c9d30fd113ac1d4b072b9baa6f1df4
zc0d1593d99f1c123cc3fd672c8e1c367779504715be64332980e13fe11895cd08c88c0cf73658b
zec0ef797bbb8701544aa5805400da15aecd6f27bf58f7d4b543de5d4fd8f1ab9ff68a5747c6b46
zb12c692ff459ea24ebb57ba45042156cfb1d98ee25ea83c80ad6640e9ca8c46040375fad1207ea
zd1b0675e83bf27a352120799b400924992e1d2f36b3fbbd394b53492f236fb19a2b35a567ded87
zf5638abbaa841fd5febcaf6beab6d06f445e0f774e651f9d495f8b8ae6b562049fe107bdfd8973
zc94b2883c0298ae58b9fbf1db8f427c93d1d373d9d1d7ed16d9e34c0066360538365ab254ab55c
zc3680f4874aff79b7a74e7142f82b3ec45d1ad3b56f351f12d650359198c3ffddaabe4e4597640
z7cd408f2c7fff23d112ff63e4a7bffa05e952f34bee84e6f5a4d4460cd84a9a969efb81a9fd4cb
z6aec140fb603b9eb06fba53e5ad566bdb3b0492739743447a3863828e49ce3016e980068f4c5ae
zab035d97dd6dde7aeaa9a69fd8a6b490db802cc5e586ef3518f7c20d76e74bbf56b7f02cf5d0be
z7a9a372110930fc6abe1073327909f44ee923fa779d91c689f33d7e61fce738f49ff799b4e2a00
za7d7cc6184aef8bda23d40e65875ee7ddaa9c404043b96405b2bfe13453619842e21b5750751d1
zf8d7be49bc14d77dfe5ee9146df514436cfa2107e2639193b0cd1c595ded77634b3127ba742a1d
zca73aa4381c17ce22d9ad139c4e2b691d41957610c0a87cd9ce1cebe75e04eaabd49457d081cae
z99a4aaf2f79fe334fc92c62fef5c95397df041b77c34ea0e2ce70d055eac9cf0d2d6fef0f5cb8f
z551123f9e9003be2252b7e991a853dbe993aed7e8e1d7ac4061f6fe051825c57315088ccfebe00
z9972571d67574881b532cdc670248b9a8dde94864a49dda5b811559c37dd7b5b4d1b52f85181fd
z07f09c7c00834015119bbb883ce2e50f84dfc33bec883da2c5e13bc0f3c8f82ea6904a63b558b3
za7df3613abfae96134e160c014c730fe5a2e4387dda7c9ae81a45d8088a9cb1d479b5f40b49a39
z481bdb0c0a679c0b9748fea5379d272c86abf6cc3dd36123112cc5f8400781295150698657473c
z2b1ad4e51519184d78e5d30b59d93e6112190d15d1a241c6b8f7be4f3aeea709377cbd00541e06
z12a5ccea2b2788c54d984ba3b101b9c4155d88d9d869d45f2585c59b92b327e2ac6eebc375fcca
zce8638f9b4fe1bc58ff3d0ff759ee0360b2767b57b0091a72916cdec1bfa25dc07e2129a48a7c7
zf7adc974927e178d9b0a023b7687d46513a1710e3e02ea3902847f8d225aa48b0360a5c219a3ed
z0061ae45209926818d9c3d24eabc0ca051fb45a4f0c8c82d33d623bbca9aa37b628e369cb939cb
z45d1014bccf490d4dc8590739e2c6b4d1e44ef29784b55d4741b48023cdaed6c3c83a05ae1606f
z88fe67e9971839da811f85f5550b912ed53575fb32462d3cbf9d34f46df26e7df36f1fcd71e4df
z6dbb10f7cbf70997bfd99bc5c5b3084416c35afb46540d7e99e575ae1edee8ef278dbc47fb8861
zb21110411e031ce59c57f6feabd126aaef061901e5c5c69f746240df75dd2ad448ac3493b34b2b
z4248b6edc1d4c1b283d2c086dad76ae6a7fbd0737d1ed128a79f976cf4c7bb404fe3e847ed16f6
zed37d7f61b7f0d7860320d64a22a8e2e85eaafee227c521da058f30eba10312c8a0058a6d0981a
z0055d7d3ce07d943a7f248d57060d57b0b8659d6943851a32ec2cd5489446dc74506e881ea09c8
zcca114aa977a15c499a1e3fb74e710a495c1ff2d1bba1d8749ea53d533eab31a469211e024917e
zd29555aaed9cb60c56fa7c9283f8101a27889ebe217f3d4cd1cddb937c0c4bc0d1351e55ae9d5a
z00d509a8520788b2497ed346501293d6af9a36ce23a31b581b3a64b8435a4498ed5e35f6b3a51a
z72466939e9a2e90c106e9b2a7ba5d154e3d351138924411f48d86f22aedac6e6875f319689f306
z394dcde216f847c8140ebd362a6541d87e8318b78ac2eb8e28601fc9fddad95387ffc5ad4362b5
z8667b7eec8085ca2032b021ec5f228a8c165035c8630b3c456c073484ad199db41b7b8570a694a
z99475ef16da94456fbbf8b2c64de0faa5c73c275ee3f96ad3fbad65c47fde71e182aabb2ae2621
zf1ede678eb6ab899db72f2214543768ad4607a09a95b61750092223aed667e86abdda216d0eace
zb9b44e8a1266b5e2449f4920f22ead2eb10786dcf8901eb0dbe04290b2a32100fee5822b281bb5
z9f8e580b04b0bf59c1088f283034ce6f6005242f26b9c58270f322c98e55df566f86e1ab780853
z8ce44e1942da8ec24a75dc1278db42921d7cf821d9a5e10455c37fa5ffafe6c6b51003ded18bf0
z62d1d00fe911a130d88c6c046d5cea86cbb2182caf64593bfc44291b9ab4f91524ee91a05061ba
z9055c1f8157a54518141f9a0313d99f7c065438515848702d782c63cdd764885030befeb9366ef
zfd7c635ed427a3b174c7b8043d4626121a4f3a400aa13ca20a3d5da2997e17ed38f24ef1f03178
z836618c75d405c1a97c654f7fd4d494e58e8db55e4ea8fb0c06f21cc25b99c86fe47d600cc591f
zd5bfe724f76ab2ac95c088132fa650fd002e5408f59cbdc5060458765d53067f0ccfbe6396a262
z8609a03c3b0eceed2d9dee432195dbb26e187c3776560c10838ea9d83713af3873e6e3f8335af0
z5b698bf6f8ba660c0f96159668db28a2caa9d0bc8edf091a5ad33f022fc26543f1fd382a3386d2
ze4d578197acf81a35552db2e78eacd4274317dc7297ff4358d4d5a9d4c811a30a000cec9011983
zf244e0238a070503eb6d1ba5b00f2a73a1ecf4356e6a79e4e4b5fc3f5339e385a10786f85c469c
zd1da88df56ef5c6f3b0e460602015f3547a5671b8f0205aa451ee05f823a076f2cdda1fb9d3655
zec88beaabd180e61a03d5142b09cb362a01e6dfcc4a92d111063a422d3ca925b7da76ed99d1fcd
ze7a592c8fb35ea928012006c7a8dfd1f840a8d6c2fe2799b0aab8d72d4374c9ef02170bd578157
z9edb7195a8d7ba004fb923463361ac2aa54ef3bb00440932fa3e04c4ab58f5c15d673bf5118e0d
zb6d2a3fed6aded3e4c955b816f65dd593f2a55eea503e361cfafea965ca8a54e1e4531f24d8fc6
z94bdca3b0bd362aa77383bf97fd2c4abaea17ef6805ce99d2037c0ab85ff37ea7c3ac8995268d6
z3b485bfac1a65f105d7bfe9fa8add812870383f97f0eb66e7eb9eb22d004419e46b4b537b64d8e
zac4e2931923814fd08370c4acf43b441a2f34cfbeeb3fefeb6fab03b9a745fb534816a03cff8fa
zf3edf381efb956250bcbff24a56dc86630809764389271022eddf190c18c284ffd3262ff65f73b
z61f11f3f3c16726e22a71eff0fe7eb4e6d3b96b68560559f228db442a9938954ea715a396814ab
z4ee23ddb081b9e3bb1f227f0f22b465b5781386ff85ff40ae8eaea3bc0632aeca91c4fa39a0f7c
z2b4143ec7784cb0c1aab9a471b9351ffd300deff19959c97a5c8cd856f455e038c7dad45002dd6
zdc8297c92a9ddaa91c000722c444c7221f3e720510833788c2911813c238d3cbf01a29ffdb325f
zadc0d27f2fd2b29a036e5c6ecee0a75f752facc2e096bea82b8733928a4626fa2018198e78bf71
z87dd414386bd2ef130a5d56aa8ab34ae2e75f731699b8e9b832efa3a753721dc480e66b2a01bea
z21a5ed33d8e27c1070bdb7581882947a2b0c56130ef1316c4c8c58f5e371ffd9dc43ae3b054b35
z9493b56ac07f5f9a17e4c8e076c189c1f30de6c85d5a9206a0f849c1c32045f0d49692988ec8cf
z84d891c387d1cde0275558f18b237c33cda82a3b5f91e078725d08760c1a1dc882b3b3d7d19f44
z8c52ce741525130e6ff9ee8ba36436758b0ed910fd359275409acdb2f6e1dc02241f2006fd3241
z7da6a1c295d9112dd1fd38ad2fed84d0cbd6d9844305740e51ca9a8852ce408c45b47199af7aa8
z102da5b5f303a18335efa54faea3d7109e1f77bc438d6e24d9659a2aa68e163e462fb71057aeb5
z8fb26e975b7eccaf5305d2a0132ac78bf61848036208da27ef6a59c95c07c6ad49832a3fd7e7fd
z3012dd87cb8adb604be9d877ea1fac88109e47ffa2697e68da32549c0a2ae12ee1ccd12dcbcb3b
z1e1b41bde9f4544f0da18bc22dddf77add0a19eae4770cb4b6a3ee666fd8c5219fbc451b429999
zb31b5a850afcdddb7ecd3d71a4668ba7d956e4c59e8e9a8d3ece49577c6c785c7ccbb0f54ff1b1
z1b14b7dacc323033ff8e83c388ed4ad22112ababcf4daf9f65d4b4c3c4d296d71a9ba1ce525f00
zb949b02012f38350d4d92cee9d5ccc6a59ad05bd7ad56fd6f211082f8acfae2409e7fa006db12e
z32407e82d574805805f00fa7cbf7ba24be604767446a868a33ec9d73d9ae189e8ab027b669606e
zc9c8c89bdb5c5617b429e39ab2e21f6e00f0a6096f841cf9df413d8a31fc731c537e7debf28f24
zb20b910c20853f0ca08b772f8b26605a9251bf2864cbfcad9f60c804e68a1f74cc6074c1626eb8
z21d11a1a11543111cb8560221f2662a71d39de47151a7e8dcd7b2647bdf002c58ff62df523e6e1
z1f01eef3d3bbf6e437a1f062d2118b0f7e60ed1c27d3f32042d25de3c9560a9cf94cf61d8d712c
z15d364075d33ab5f914e35e07ab075a6306943ce95403d3a45f7b6c6a30f6760e5212495365c18
zf636121f7659c24aed92694e07307eb6b6c5b5870832440cdc6297aeb8e5e8f451c9be4ba77f17
z88b2b5e14dd6e80b6e72671040cceb19ad3bec706528212f19a958c10bc1b2fb6fc2f1e0eab828
zf3acbeaa0d0216c5d05152b489ac0783dd55a4793b63beff8765490e86488913cf253a0f6b3486
za418b22767813c99d2bd86a461e058dddfe4056b65634e5ef62e44059a912958893d26952f9f08
zcbb75ac709effd3b807f1e72bc06d1ec359eaa5654590ec8dbd8f46cfba12dd1d6a4cd24446ea2
zce861c2fb516205436819c42b1c0dffd0b6beadee279663509be28d867d6722cc5b225bc1987da
z08887a696aa4f597991a285687f58a6f578a396be0581c99bd0e3c5d37fde22dff1455f5861f11
z55e7995c56a1dc6f88bf9f034efeb5508add4c97e08254f6a45bb2bd1d28e1cd0f2da68c3007e2
zeb197e9d3c9e5597a66288a39acab85e7fa99dfa41fd05214e9433a34790b1d02ddd5b010b59ff
z109d83d25665bcc3bf05364f552c824534600da5c7a0540dbbf59ca9424f726833fad773142135
z4f6f131142626531a4b0992e6bf681550fcc2d15fb8b97b25d5c57de4684176c3e0a0c566914fc
z1290828778b5b06b4d77b7b0b82451fb5d4b30c307b9abe7b86b7a89d049fd399c8afdaa83b1ab
z7d8482cd5c6c2e7fd2d78ffe75039c27a64d1d7bc31d63646b0447b17a1a2383ad36bccc70d187
zfd30a43ebac6e494268f59994b6a43426035ee133980f2aafcf2bfb7721d426b71f366676b80bd
z2ba2e531cafb2d6116bac08c01495e0b88eede79c1ed9a4767290f9d39ee1c39c741115d30ea83
z1b8d076d40644b7c75341af1c4bf8f1273f327c694ddd6a0bbd00aff8665f539746087410c94ae
z28e77829db2fe54e0ab3df5c86c4b347890c489f4d04da9f14a9f83e1a429713e724b8b5ce5abd
z409e0817dff11d4b0f0b8d0db91fb187399473cead0178fd21db8c76d5e0e465745062d562d412
zc3974fdf4bb860af76ae99fdd9642767733bed297b53297c7bd18abf48c3501997a7bfb39888aa
z8e35ef66f8ed30e54f927875ef425532add318db2337b76755c3b38df0a60f934e74cdc0884a18
z9361ceef47a975d4f4cab5e2bb8554ac9a8bf30587ec31dbc08c164dae40799e0298dc8e9970ab
z3a66ff6fa03130fe24b6c064f7067aabe0024052fc88a803695058123c324e3ebf6aa8e7d8f901
z7531da7d27940188d9e5d5f02f899d1467f6c90a88b7c25ab39850a8de6905fe94826353088432
ze4afa81e9508964cc9c5e7f9275a11d67ca2c1df0c2b695b97c2c750e6076b38e0514159506ab6
za16ae8a995ddb8c27ef725165626b1b10b48211ed5f4fdaaedcd2624e3acc9e5c7b83c0f774337
z22a04f1cdea8d28f12cf40192f281d2b5acf4deb0ebd0cc141c24d6d6ea142ba517efd70ef7274
z3c82feb7f3638d03cd5fcd24362425beffa80597552231b4c99ed16ee441d2826792c57dc7bc0a
z214f94afd71d7a140c6fa536ea5f248936ceac4e018cd43ef9e551fc3a62b89c2a20ccb6141a09
z271724015b221fe196d148363e06064d2b3ca91ff30f10a7d3d2435046dbbdba88c00ba32aa876
z80d01ca4a81e50a3cd789e444fc5458d3d4793fdefc3f72f9b6b47d5db5f57301086dbcd3b80c8
z6703cd9d277485af522d7b60856fafa9d6fb0895117d8ac592e998fb983abbbb593863f12b8526
z44add833e0d203e6f921d57d76d46fcd6b3d7297b8f26e08225a7a31992e713aa759195d753d14
z92550c22fdcea5dd2ba46259a04d433ad77e63fa437068eaeebc65fdfda5e8660589bd86177487
z50d552aed82f2d07475642df89de8557bb26cd96dd3bc2bf074f31a876b8601ec7d9f070e3ec35
ze7a0d1c6f4e6963f6745fda8c2b0d755fe70f826bd5b9bcd8631c1c1274898df7cf100656ecff3
z5d65e54bba1cd05b4e9efbc33366c5ac710ebfdad58643a7f76e4ac56c88a94bd03a2c70a532e3
z7334e5f1d8363b784ef50f1bdd367268c1c7a54319373113e99f88ca5aeab293ce90cb06be9f3b
z0ede7df4d372f32afbd1e9f4136a5a9c3e2e33b1d5df432a89b68439f82013f882202cbe0a51bf
ze22ff9d14f0ced8da10ee0b1f5eae16005aec65a47af8c3fa15e73ec162492daa9cbfff472625b
z29afad1e825777ff40ab31b50b1b423e82cb687c751f2d400284fbbeb8433139e61dcd50dcbf4a
z7242fe75bf8215fcb5b2173f3b0b58e03d0742a7e4b0ca105ad0952580c2b4eb588341eae5ec04
z987089b08ecb3ff6980013bea02d471c45f1c62c0a0b21784cfad9bd995c469d0ccfe3359419fc
z2f951ff9117bd1ab51d45c2872bdf2c57f699c6c197b2f4499998ced8edbd2360bff1a85c3c297
zfd074fe79351225a13d0ab3af416c0b061265879cae7616cd6d1e84f4eb9323ce38b3e7d716fe1
zd11ff4e03b3259ed1d5115e8ad20c6f20d9d46378445cbf942e584aae19235bddafb79ef172c90
z1878796398d69ba94e3b325f225b32cb920c6669a17509839ce4809f587037511fbe06eb9a8f59
z223f2258435157f1655bcb80284558549d563563a041b2616688a9da301e6da6a3ac36963e313e
zccee247c129e7c3c53defb66eaec09430acb60f9cd9b16ccc269570ae95a659877769df896e1e7
zd5c251ff8f349d661ab8706e71d718b563cb22e7005fbe61198ae943febb361c36fa244d053ac1
zd01729e6bd0bef57b9aa8a13f605d6ac5e67001bd57013a6ce315049a13fd3760a5e75f4fbdd2c
z4ec861fde213dec27eca87fe216ae9a56711188773db407a23190d6b48ae16341bef3e67aec9c7
zd014be58a2dab02fbbd7f6f4dae7d2ec8545280f7214dde6c081fee9045e7748501695e498cf20
z585adb5a410a3c0563f463982e8d531f15fed9c3a50ff526f0debe93f84ede44a9a15b8be024ce
zbf36e6bb303077aaa7ba761940c30d6fdc4247479e6661b3961ec0a907da2f9005cfd4c4812d1e
zf4327ef1696eae4f62474bfee06a44d0fc8794446d9368b034b48d8e9c15e79183bc93c45cd87b
zed5606046f95878ea46f072150f6a3f1fe9f05fec1a7e615d16cc61ce33be0904e54dbcddd2953
z6174a5a132eacbca1a7fb744ae03268da863fffe26133be9e858d46a75aac543330b49f5dc539e
zebb6e50a06f6f1451464af60ef67efd16bf95d8f363b0067c92a1d47fe1b3fc7933b48e53f6371
zc642b661e6629b34cc1d160ded7f61976e6cb908458f6b8e311f1bbc917884be370156c599a45d
z2b546fe66d9a3ec0b5de1eb01c27b5ae3ed5cfc39f94ace89bdeadca7c64d80d034ca7644b5471
zd9c609fee76eee63d60a0875961e273bf65f19436ca70f62021d7bd2f30fd306d5934548d2823f
za39daf5bb8dbb313ab2be8d657a556c302517f814db4278415ba49c3f693ad4282c2b2c29f8199
z05cfae05e8c86346551b561894cc7111e672ecbe2e80392a222cd200505fffc48ab0b9dd01c4c6
zaccefcbf596bc35c9e20f850ea0edeaf89a77509d2a508919fc642fb02d9331b98a4b7c4d1a5b6
z307691ec924944ff0967d7bb31d5f7b06b7b04276c7958f8b4162a4fb36df84cd0e5b78e2c1ee9
z81771238c22371291111512e3ede207f6e7ad2309ccedc4dec7266e1eb439e1e7f1129867a73cb
z1323fb386fce050f83bde79bf6917bbb771b606d2dae9edb6262cb4cf6ad9311e451d6f8dab3ae
ze172cec6c81589278d068d7fdcb797d4323712b31fd173e56211bc12b7e16dc89cc1978683869d
zde8c8a3b3e741768194f494a76c88e6a9fbe1ece565193c250c60679de53541a6fa337f4337c1c
z5616b8dd37ac821b8b68d9c75acbee635c3b3bb55628e259cbfa488a88d4a7e1e97df6582427e9
zd4202a8a497ddbfa9d36df1d72f0e66681ae9f968ed6bb398148c2b412b61f6c1cd72ed24098bc
z4e472cfb3972bdb96c4b0cc31256b3a3c088532e100f950a47fa6eb8bb154379b688767be2c69f
z85fb777f807ad837b73324a96b1ab118b0b6385650d102817eccd75b4ed7a1c250c451dda0bbca
zac5dd3f17fef80ce54657bbd1b1f1575cbb2ee781755c83bb8c4cd743360570bec41f5c36a6e4a
z27a0562fbda357a9568671235b3e44eef01a800175f1fd23c16f28aa21b4fde9a921b39e1056a0
z570dac498dc8a4456c1eb506f6c85630aa769cebdd0c10c48b340853b7f301a49bc5a3f8975065
z9a49a06f0ad42547b8b3a0bf60842194dde070da133dc105b9aa72689e23d441c3d618c91ae7ba
z0b00c46708f01e8c24c7770a3e19c6501c41c372455874ddc75c8a807585b59512e236067385f2
ze4f3279ae5f2607b702f833e61aebe19e4d26c76fffc0478244fe163eb45b854e02da8e0d88e29
z01f22ca6dea5faed619621aa665c04f7014b49dffb8a1484046a8fb7d4ca25cc278538b840f35c
z0dc4036dfaa712d714cd3296c2fbeb9d54ee2fa94719857164a7cd15c26c11871e879e0ede98e2
z8d9219f617c36d774a41da4ec25dd8ba0c550048e41d20f477e99db0b46adf8e3dae9ac2bfc68d
z6cba0657fc255a39ec03e931cdde4d6f01e25ed2dc4338f9bf5f66d8bfd0bceb91e13066a956a2
z80e5bacc5605ab3ebbb4ac636f3285e71cd0bce24cec7cb577149431b6593f9a13332b7281d774
z27dcc6e29910cf7ae6a490c584d6871d5be77bd16650c1ac6fe37a13034e402d89c866710ba313
z12a29872829e16723b06ad2038a09fee3d7195a0901ccf1dbcf834a993d8ec8cbcef701c20bf6d
z32730456ff75427f58a6bd5017f480e31ec0001b83ba2c071b5696208ce6b9d93a97f75eb3f36a
z4cab340ee6cf58688125ccca3628b1d6770602c2521b027359d92deff710b6480cc408533a8380
zab0b070da81cb28aa1a38d03b46a43b65da0b526da486a39537d2725c814623bcf91d0eb3efb83
z5173ab47f57bbc247e698d1c55171ad2a2775bd4fa54aaf8e741651d4d9cdfd3c2831c8cbf05ea
z722453787fd8a85f7b0833fbf1943e56caafa03ac5720ae27cb38692d4c08e548476029d893e91
z2fced47456d34fec2af7bf0206ec6832b2a67c0b91b4ccf354c0b4cd4d460d1776ed9258b94b4d
zb3e514155468424e027a3d768e4b96c4c1469a466aef76f7087d0d91986cb23f1efbf274cec7ea
zb0edd56d238b2745987a38fe77c0ccb5736637d87cf3511e8bf838bf43cd0d05fdb646e2bf98fc
zfa78c1f2b6a6fc0a3d614567776612ff580a5576dfb58d398705d0175fe1e01e52637c593def70
zf7dab7667c2ef229c3ffb28899e65b3f73a6a0c3f8ae8ba2dadd294fcdd141ec8182b2df440d98
z643cd576ef12a6299a0a100b77b82d4673e55c3a36f83fdb8368d6603118083cb058b8d602238c
z9df1273ef5a351df12193e4886eb9a64da39c4d60c2fea4bb5a3df80fa125f8189b40a52915db1
zc45015b9ee1fc114dc5abe77d06ede69d39712a140f7548cc0b87c00cb72a85ea15fda3d6acdde
zc6d721e7e7ce5ff085d9e03eb5d7903f4f1076aff0ead97bca7c1ab24c42338c29cdc2a21e53e9
z555212a761308e9a0abe2aeff72fbeb6c1421bf74c56f9a240b39ce54978a10e70cd84eecbb86f
z4b1f84d9575dbcb5a578f394891763917db3cfa1e0618f975e1708a812bd763622321d45d02ede
zf2c563dd842a5fd8b6283186dc2d434df080afe602b6d690cb30d8c840e9f2c7ee3a47743d4137
z451db84cf9c0b0a13221cd6dfc53f9fa5b2ef6b7c7028706afec143755ea9d16ebd589cb21918c
z942abca64ab46ae58365e8968f5262ac5351a23543ffc4263c488980701fd194be6f8f95d87761
zc6ce9b87aa9aac7245fdb2e66f0bb5bdf8f33560a94e4df0c09542abcd5fe58f053d675e47f4b8
zcbe0d6bef5d0e56d4c1c5fe2edbe1e86bd5ff481786ac6fd524bb9b1fe08979cc95e6ec272b458
z7c172daf9302a58aa71e3628562bc79909f65b5526d4144c2a7f9ebd488357b7059d2f36ed96dc
z16910a7b14ec7b445475afd7679245e13e9db386a62d1bf244701ac5316f9ef7fbfed6ebfc5273
zb79dae95349317cccb1f4951bdb9d046e999957ed3e7e51066e946a63181a276f469a4ffc4c3bb
ze10d7138c5afe5b010b8d483ec406d533a73307b43779db52d5acbb6be8abc09631ee96d1c143d
zf3ff27a83c9c3946cc80093f44a1bba2779945d827848457f8a02e752948ed4053c796f0b026d0
z9ce2c993d2a6f0ae7d32df6c1308522d1e6c8ab9c51eb57e8e28fe8175a20b486bae152996c9ba
zc061163ea2bdb63ad2277ebf7bb437e082605bf8f30b6dfbc2932269351b824ca6961bec7fc0df
z919e283ae8017dcef9b45196f704f07a8ef11d0ef165d37431e454e896ff228c1a2d7d1dac9c9d
ze73d62c959f74f76d97455df24ed5c680cd850b3bc17bc38ea197e6667ce232867219331d47a06
z1ef2f3b08d031d4f0f2053913127a6a9ea998790ef86212585d97be7d67681a519be3ee5aa9abe
zc4f8fff5abfa0e1de565ef73aa404133cbde13a0eeba973f7191a318eb7db81819e6f51ce4420f
z91d0a787ea70c719fb757b90442f184db49f54d912260e5b8bf53aa2a887b37b600252df7bc14c
z1600778e83330a29b5a07212bf730b03ce7eb2e096596493cc0bfa017c3e4bccf75baeb1ab3c49
ze9766e40df94c601663ad985c3db79b5e8cc844acdea722aa2ef60658458e5e3d8b8833a2af56b
z1a38e9d0f90cfc201624db0df080a249dc0a7192ca75fe7f77ac4bc9d002c7bc97ee7a39abf678
zdecd0ad1619fcaff053a37048418e5b7d7e8f4f521f498fdd5417147dfac3a72c8253189658fa9
z87f29322587e8023823a161b5db7636164243c0b99659164cf840a30850a86b15a1b17a366ccb6
zba7261e3c71971ec0613080e33e7ef5570dd34f736d4f648ace8236b894c9e6459f4bfd2c7ecbc
z26c3b8b6795970f14c98a46d21c9e9fd727825ff01562164e2631c7a82f88fb2eb789edcd51b12
z5a5793e6e784b573ecbc20defc85d9b02ebb3e4ec502ff9ead7968ef393c1a8f72489bbeb5edab
zc6885d131387ca7d82d6a28d1c6a16027898a5efc2e4a3cc271240422a637a1cf6d8253c724934
zc5a567225dd33ff30641ace76270acec8403271a2eaaa6d97ec9fa2c0fdb9698895b64d15e8100
z86522f036e8dbaf9edf3077c41c84086c5684bb3475c433a6cd4f102afc37d86fdf46e21c29c26
zc27e69f79307fa21d56f000a43dc1f19334633c4b6e87fef76db3bd7a400bfe705a50176fb3304
ze6d5034495b3989c66ac44681af18eb8e3353afb0ac19fc56544777143089d3f3fa0ca3edb04ac
z8ed58aa5121c91880e046138977fd4c3fbe7384546d6c002a41e5f62618bd21d147bb1038817a8
z25c8e4f2e47f41da5198f304e87696591f62ae29bf879157818ea907c3f21f9e66e68b56261c5b
z89a7c0b11d7c145b1c06d278725c4df1b5dcc08a3f3c1f33a996160f73b55b183f5f5f47e33f61
z8fc08f70007bc894b221c36b9617bbb7daac38e91f2cf2caf10f40cf925de7d9683b32ac79e081
z7b27d2276e48ca69c6d2ab5d08ea8ff5a7f2d402c5e76b240a1961e2fe695ed9287dcaee4d6213
zffd0ae91ca1f3415484572d9595c66e7fd3ab66aefc5c802136c6ab3f1ff6c0a7497528a68127b
zed9f19a2680918024546d0400ceadacf683cd5082ec8de98b340d9ba6107528a1addcb94ab673f
z99042f5774b234f62e4f4a0394d7a9d0e2c9f59737d93851e52fdf76b4a2e91f1b4cafe44ee978
ze98204c982adb7509d45b9dd9eaaed4adc146fd38a909d8a44120e4d625e6ece59158ee0e074ef
z0ed8cd30b7f1f718c6bde9ed632ce1d324a5a9132022a78f1d5ef69b8f15e72b6f8c114599405e
z5bf8230da81d421ddec54b8b05613ccdf3e6c647a2ab4e251bbace57067af04470711d3a4b6811
z5e1d2daea64d13ab73f64a2e50fc99ecb63ee6b01bde1370ab3b1ff2982fbf85e1d24654cd75a1
z4a8186827ac735f71885ba5bfae4914734d2fd6810062e8b1ffe2c59bbf2e905bb6ccb13061e86
z105a4a8357d35cb4f253e58ebb1927382972510b9bd825454d0db212b45042b9dc63997f824c9d
zf6f292253227ecfae80552fdf0dbbade7f71589ed53a57ab3e2b050bc01779b12a210d69a66db2
zb34794b95b55914a7a62c05e104b591579e6353da45275e10df440d263f9f7b4ba32d638572dc6
z86104e9cce9c69be3caf01f4d0d7c0b7be7f4b49855c2b17bc7cc52cba99170874f373a526fad7
z53d1d86e330ef97c1eeb5cfc3f5afa4eeb5f7596aee0d8cd1ffea18ea01880fa56a8565286a24d
z4e34ca254e432752d34dbaacdd1c8b053d2029dc522371559be4d8bfc195efc14bb20067ba3dbe
zc44ae155beebb8b35568402b43bcecd3993ea0679c3209d92bf8c310447475063f7d40b4cde1e3
z3eea6c7f571da73bde9b63acdc7416e5c954ce7ff8b03c57c5fafacf5ec31820b0152ed56e959d
zb15667484554f92562efbe2ef3967ad18ac6db45744b4895a5395c35515b4348c3d03bacc313a1
z7dbb5ae2cb0f1d78a963e199ae82e3ff7b83ac6ddfa7117d9d6bb533072de776f6ba5627a4d989
z47f53c8c166bc2cfc68ff5bc7acdc19c96bcc7f1e6478e02392e89df2c74f154f9921bd9477094
zbdaf254e7e81db8b1294f0f5c68a1324ef5dc57104e1fbe2db13a0faaa0d594030da83ec5586b0
z1b0b0e0a926a28cddcd76b90f22f90bbee7d62283a0b048242a7372951a2ff4ff20cd5b56b0caa
z81d864027de55256c922bbaf2dac2f54ce707ba15b31d0527358ef496d64c075f15454a38a1b5e
zae4bdae2eedd1bbd350643223cad2a10680cb9cef6b0b01ef97f75e2112ced2015fdbd8ad59dfe
zb3b1ff6c7eb210b656ec76c011ae7be04ebbaf77b5eae8102b52e53edaa99f7e5f15c07834ffd1
za724b272040942065096a04d953e2a3c246571adcc59cc6268710102fa7fabbd61440316791fc8
z854fea8d2b99c1c0ea1e2c8c10509f5a515fb636c8c449bc7a9d67b4489c4dd5b1f51273f91db3
z24f612a98eec3e3cd9dbe3832a1ebf2370f98223ce15130c6b0dae18ae4c8713349f57066e5404
zde13347cc60ffe63ce4b4434860e7655f2475be73f4da1ecc3cd90b51c9f52140243bc5f990751
z9b43c69aa2871daacfc2988a88a8818eb64880990ce2223152dd022d2dd61ace499b5716a52b28
z4d5b799cbaaa02cc9d1f256a42ae4d580326418b14c32dc521b641287eb589266860295ba18a11
zf4c49ce1d16c1b90611e80e1adfd437da986eb09b5ac194b40ddc5593af453ab8cd2bd3e26298b
z0eea61bce348f416be78250c14980c1d59bd9967aa3dd7e71c13e898d68b30173755896f139fdc
z714d5176168ae590d84e5be77ca905165e6a8fdb8a56fa6cdcb08eb58464bb2c425d66b52fdb51
zc71e5a88a39b8f02ab2c0b56eebc5d455a5657203b51c7343b0545319fed72661489693992ce7c
z1df4135de5ee0ee3fb23676961c4a1d498533edf51946403430ef3ee10d1484888b431c54d4e38
za09a069ee0098f63e2b6033d9832f8288fdb7a5ff6af9a924bface68637213b37d9f9285e5f00f
z6ca072014f6835787cf0aaceb0af5dd2a95738dba104136d214cd92dfa6562a5e056401f60f201
zd7a0cb07475bc8e672a32c729970179114d09932bebf7b45694b271ea9f1ce892c98aebac29492
z99eb4e38bc2ab1fbdf9d57967308fbde91e1dd3ce5e0b67832af4dde8832ad718f65ae4808e73d
z71e147afc32167284118c91d99f49d43b538605af7a256e6e862722c9a53c6184a12ab8c1902e2
z926da34467426ad12195468113821b04cae68b214f87dab288b8af11ff1283fb88659bac03814a
zab10f872d0ae3ff2cbc0369340c35bb4e57f799d8efabf35c380e5dfa5fc35f2d5a274e94b4818
z50c463eb3f3623b52150724ec59eb8702171ed80679588dedacef87da6700848180e112d0287dd
z881ca6fb44db144dd166451f494181ac1a76fa76fdb87d02cdce5ae81a34b6b1180a7e09c89917
z0f34333da446629082728f70b2dd70a9858f25294d37f7393d6756ad1b90d3fde1f83922d92541
z316884ac2dd6202b4d7e8dfe366ab2d3f6a91be600b49a823c62ddd5861fd998859520746f334a
zd06e04f36cb198dded8954c6d450c305ab271b0cf7e8c48bc6c5503bc554e8d75165a07edcf37b
z224d42f19c522b10b9d744dd1e5d3b8cfe2931faa359b8c6f8be5b3432c31e3beda4dac624c29a
zfccd72913990269938febffdd6602771a6b7277d954a53d9d4d67243f4ae1f8745c5407b2f7159
zeb0fac18d5f8e440f8616d8b020272ade4bd672add1b5011266275437cff43b37e41fd45befeff
zc8c7d1dd2bc52a2562a768e877f42412060a81c79b21adddac29bb0ca0a95242c93a16571d6d24
za41c46312bddbcb9004ef53ba70ed6e46603ea0123644e6ba01db3b4ed1cd58286cd0cac79c3c5
z124e228dde9dde009bfef29d74ea9c89873cafb5a584da1371745e61d2975373cf6d430a8db0cd
za89818aba3915680910c40b78063e0f8a33b30cf3f3ad3e6191613ab88bb62f17ff675a30dec85
zf3b66bfaca2f3a47f159a25972bccd0e558400f80fafc43d01d3f031c07bfce45832b6f08cf126
z1dec6849d5475366d908262a2050fa7546155c892d9f836e26bf689840a55b361a312ee104efa4
ze59ee8e7c8a7bbb80f3c3f4c04acc5d00684a10c4dfef78334bc9c162ca9f30e94f25a8b301836
z3abae17de6426fa3518e8c6d13ce2aa9277787bb3b4f21d54a2d733067de6c9682c66d9d3c40b6
z965fa5bb51b6ec6bdbc118ef6233c4249d2622e56703225cfc5f88ad424a2f909018daec458db2
zf85178d7d4fff5fbbd8dcb93567858ed83d34584fb4d08823bed7f56994cfadac8fcab045427f9
zae8d14a9752083162c59ec30ba6722c96dbca3a4dd275dfa5d9c094fc1a47eaca10a501926354d
zb7ec2719e884cc198d7df52ba797f2b16603ee079ef8d9883d12774ee920e094f0a52e477b38b8
z4dec842c7e6237182e46eec75481498de563df7fa667a204ef32d56926478fd960cc5dcac768b6
zbe3950cdff834324509e4548aea601358dc78ea3d56dcf2db9b5ae36c87592e8e8decb28af3cfd
z3e9aae4513787997e6dd3b6cda7cd154d1d7e89e1e50c045e6b5eb299af599b72545004d44f272
zd4cea9c41d8e36182a0fe518d52ffdf1ecc05805be5b82852b3fb6ff13fe20b5d386dcf1f6ff15
zb8dcf4999f3650becccce246e39e7ff150605b1d484cdbe67e50bff6c709e92606551a9da23887
zbc84e8053af7f527c1a58cde236f9688731f2ed814d4e90c973e8e5810b284595c9f11bd407c44
z36627f9859922ced8958228d3fe29246af120f9677fda101cd906a7db8f09e2b5bf1469c4a9f8c
zded4973f9bd94214cbbf2734a3f2c680a37b97096da9e63ed76989304f7c2c4bbefcc72d638119
zb7e55171911ef878641fe189bc3f904715586aa42c8a18bed5faea1bc4f59fdc0e2a725cfad390
z94a67c6c650970e74fcc974a3c379dd79d9da34c2c3c8b6007b833e0a2eda5eae90eeeb3e20735
z3d2ee2cb56e5d124300fcdd86d477cfa059fcebbe6de6b0d8d7aef778b5c3104530e0bc6843e41
z5cb7d4084cbe0d0142bd881b3aab90079d35cf643f5cde477977923e413f1640e4615a011332c1
z1698b1f3d69a41b4714bcfdbeec0984087cdf464ee4896473cee1decce0fcb8a494da9d6f1eba7
z3a9284f1861e295b638273f1d835308bafa6e4d696f73f86d42f141ea009ec1abb40eb75765e5e
z07c8a524b8e8af3f63cce3a4a0d2dc0191ecda1b2237d6a6fa0966cb4bd4045b5b79c5238b70da
z9d70fe67b0a3366b6e753066a416c773de98ae2151e2e74e6d53cae57da0da56ad0ca74c25d6c8
z30bfc2d299e6f9d21b53d4f5910a8cb12121574cb85d4565ac9be833aac623e1ad238e8c9d1199
z5509267005121365b5223f0797832308c40ce2cfdd6bb4eff0dd990c72160c12423987dc7788e5
z8f07a53f422c6e3b1af7aa0e83a6e678f3a7d5514006cd898ea6fb9eb573db016329fd060d3b2f
zbf8edc8a3048aa43da42f9d5cdc8878eac21e7c161893693bb940bff85871e6eec8a06c1583612
z679aa2ac1f09f2590129343fb2eeaa33f4c2d29e3c312ff2e84d414ee3da446950042d901f87fa
z74593ec0baee873463322a17d0118ebdf8cc1b57d626310b417074f42feb7c0478c254a1cdb83d
zcab2d74eceb3dd54ad95e0e1685f5669dad9596cec4663fd83bda7b9dd1c89d802eec284f5ff30
z3295baccd2e3a3eba2a24b6810a64edeec00a3ad728802e418f91ce9031f39d1e4a93ef42c4ceb
z21d8a7c7c41b4fe97cf0bca81af0b18cde50bfce5b8acca96c184ed5998ed432ece060c00a15d0
ze1c77a78325d9c56b5c8fb03c0451bb98f874685c13e5bba3a5c3df92118bda319eb55314fd87f
z5ec0a032128e698ce89edaaff77dffeeeae940dcce99bed6073813227d1d430f512ecc287bb92f
za051f71710b15ad6799039b5200a33c22fb3134a74a24052fe3b3baf78a652de781d502e9b0849
z458ebe76982e4e03b9dda00802b69ccae0e8a5f9cfd98eeb03dc174fde757af258425b36e89f72
z60bb619e31275ed9f014bcab944ef084b89b0f542f8e08c8202d197776ca4a6080e94128fd2acd
z56db4ae6ea022c26622f4f8a523f8a45926ac090a9c4307db770e661b2e36c83d04df2753c2c18
za86db92dfc0fb44d76bb963b6a7be17b96725d23129f694e1ca0d79a9f07cca7988a0ce9d6b283
z8ff15c01d2f7ff238fefd36f917fcccca92cdd1db91a70c2e9847035669cc32d0e0644f8889ab0
z20f9584b00ab0d1a31be8d5495072d5fdcf91ea07f5ce7a6809466265ce4bf40c737d5fdb2a91a
z14940d898c0ce1d29fb9e4a9e36852bf9dc591bf9efb9b923ac3d6fc0271cfc6b79a54b2491142
z98cd422ba3dfd73dea3affad1408e177f2786b35f4c962baf6c876c8625939ebf0d0922389f24e
z296ab3d7df4c1f6f644c80bdedde914a2dda8f0e59e00c552c26dd0afeb642a1063716094996ae
z1f8150b7ad0f29ad36ff33e4db2d21d5845b31a004314f5d4e40067688a8381c4b761f9f5ad840
z6db89c3974f5d866ac8d738abbfe20eedfa473098208e64d26f856728d541608220618df1aa1d9
zd5586e40bce7298f7e3c52c372f6a8fa61c9d5858db6eb572946163f0904fa854698abb4911d1b
z2cb87b25b3ef0431d56f67472b5523a1eb1e8895f14cbbe5445a6c97e621d03293a209a898213b
z5140574c8293c9240ce2eff79bc406b3985c08399a287c8cd655a637e944ce12e6743447ce6874
zffd30a6c5d6d5415359da5886b5b3d415045144675fcce96a5832aee0ff762d2746fca1c63cf0b
z0071454df468029113c6d3e9208ea56b2a7ceb628ac52fe21a1b1af807cc0efb1daf527a90e8e3
z0f1c37248f0db3bc0498a583a4d6b7c4bc618d9485d171deb740a47f4b5b35cb6e7d3cba0a4cde
zeeabeb71176ec6324fb29ca3f4d7464eccf7c1b8e3e139e836dff89c36e68a3fcced27c62148b5
z358f0968711746e94d2e4fcb0de6d781e92f37dd4ddced0ac9d2c596117983c6763c38a1614351
z415e1a0e3607c268a3b8e66625db532adfc9376e1d32870223178db6bfbdd3574a8619b76347a6
z31492a3206742a0a99499c0017815d82ad1194dcbac5ed0932c5407d8b1439ba6868c5442ae91a
z2aede24c50a36975c56c329bd97b0438ca44375637ac26ee9b52e586730675e0e6478023567f59
z028c5c1cb322af9c544de8741ce75594eab34a953f73f01bc297884d69c99fabbc3003730d9fa3
z49a79bdc25f93f73e649203df32d4db078d2c7528b4b88ccc38d360213a3b5effe959da9ae015b
zeee911774d7de04607ceef08b62b58503576b0e8d8f4d8af15cad5fb14a7c1986c110e976f090e
z15f6c22ad3c54a65813e590ea75fc1638f921ba1829d04c75b1f3e0a4d3bcb94bcce7db21a24b8
zcffeda75eda01cb3921db02703a05dc83b5acbf30ef28a4e20c1b6962275d1a2c678e5e69ff31a
zbc4ccbdf89362b07bbb2d05d565d012b8e373312c6cc89734d2fc1dc4585dd5fece71d56868d19
z4f33edd72edb1ef0593a1ad5c22f2178d02d9f946572415fb4c77063df302e2590b7986759c6c5
z8a7f61e7443256aae517d2698c7113926ebff27f31b94673c370ba791e696f7dd48abd1d4328b9
z1357d6bfa6dc5d3925ef0da52930b576634d032c585a6ce9ba0eaca9505f8bef93c4de053b6bf6
z2be0ec885ed2309a6f3933495b26e9dc3a4a5d50ea6ab19ba0624dad039e180355e9a0c33974eb
zc69625d6fd1ee474e7e83788dd1cea7847fffb5a0ba7aacb9df84f525df0da3efe85722d41e5c9
z68c5182895c53d3f30b211d6d70e0369f40d4ef9f19f394209cb631c5274a3a44923ba9cd1fb1f
zfc441458dd1ad6e781cfc6a834c82dcb8cc3c6b1de8e1be69a85a90977b86233e49e8e56895ab5
z7b5de164edd1074c16af180ae2ee78b2027a72ad31f99156970a36598cd6a0cbea97e87bd47f94
zbf0cc7d7fa2d12930e63d0181090eb0c254455421c05334fb3ac934ffb1a22bdde51e3eb9ba679
zb82778335363adb2270bac5c9d96432eb1e16953b2488a4cd704b76857396a1fb6608a4ee257c4
z2cab69c9061a1ba09a9258335cd43687aa8e9633c90a7f2becb17e2321ad62a603e69281b2ef78
zcdb81a61a82f57e6771b18396738b3b5f2b0fea25eaba908a106086a46fe16f4d645d9ad092bc5
zc285358e44b155aab6bc11295d0a1a5c9b3b70a6733403d27f7d59604990e0c8fb70b3e90865fc
zf9e2ad245f9f70788f4ccdae3a5edf5efd2851d3a7476f6fba1bf9703ab90c0687629592cc6b9a
ze1c600480da6531d79d4f3d7721c5c420b2d83ea8378d1e2de9336c04e2e60d919c4573cd0334c
za7f29f71be03bdfee169f5047aa509aecb32d4c99b08f84a58e2328322ec63b0f1331440f86f33
z21f5729cc3296c8480af085a1961ff1d60814ad58b015cc873f176ab8ba7f34cd51b612fe0ac2e
z20d54265bea21431d9bb7498dd067ca9822a8e57e1b1e0c5af307b520d0945d589cc23ca223382
zfa61294ddd2d91a74fb5a253c542783ac581c6b2e3fe188d02865189a134369ff98f64e1e29ea6
z6e5696b25ebae929ab9141e3834dc50207add78d7d7870fbf75e62f3a3ca96bc1c3b62cd5bf13a
zd51ff675fe536ec9cc62f4721421afe9dcdeededdefcdca5b5ef1ddb74c80c78ff153d00be3e5f
zb44594ea41d5a08eb00717af9da7c5d9628c0eea187c9c343161f321a20e40f2e3eabc9baf1fdd
z6025fb82e9a495302083ce6f8c8b72e6c6df20d4b72f5f6ae6b3ac627435862b203699c4f3f1da
zbce374bd8dbd36a168d5e34647e62aee070ace206458358a3d551e218126d12afc59f52a0caac9
zcb708faeeda1c7f8519d1d91e801bbf65d608a23a49ed73a63a2d61a0583ad9049d45abd1b92fc
z4a3f059cd04f458525eef063d92a38c62bc4ec308f1ff54e9da5ce29021269cad69f3b88d28536
zb5cb072d431f68800da767e9e0cea693768b460626bc6243921223b8edfc17251069c095f233ad
zecd080f9a72581d44d26c69b8f4148b54a12bfdc5ebc3635399120d373e0abf4bb0219cea14722
zc8bfc59966b0c4901bc68a82df840d017f9241c32045b38579653cf5f5f917867b7d348d96efca
zec2eac4a80b302ff5a590d96a9607d7c093a224b48e4c63f8979c78095ec300bc31c64090d5fbd
z78d81477a7ec5c2bab1f71dfaaee76e023ee1c693ccadbade493c71be4ac8117094ca4b4819217
zc157c0c394ea2ce8cb790a8d65ea0287e938938d86ce991bb721bacd1c50475bea5df125eaa653
z4a84425b7841ac92c95644c7861612048e45ea969c8a414775533af5b27fe91c3fdd8388d1051c
z7edef27784a4dc6e7642b1a8a64f0b58d511d44e1355d14397f20ec895c4c5412091ed1fb8fc82
z296b4ac7c8571ed0417e40247e814e9104674395772fdbcd4d37b9017ae297771fdc14233eef3d
z983b2ea3d947ba0dc99d3aeef89c44698005a2355901aadd13d14fdf3a2ec1e944c089f79a2e0c
z1fadfa7f11238496c7551d54412aba76861955ebf4377e46ffd5489aeb61d23c69148a94cb03ad
z2cc4dc32ac87d282808639846a3531f9929f3caa295e4fca453d1dff587431e82571d378860c13
zf920a697b96ae8a6f2d172161177782080d4b5796a9fd3c45b00a05b2269faed19f567704525cd
zbd03acccde314813a5286041224add71fcebae80ca9aa03aa6a21d94d312a36573fed44ab3d210
z49d0bef2cba80c62bad43cbbfcdac33b85c04a8b40f80174c25f3f06528cd5a0009544905204e7
z52e8c0bb9c027111121d86c20e1bd9ef07e7641c96fd093d3063180a94be83756c8940c7c3e6a7
z010403c8e41aeb6f353cd729bcf357dfc61f33e936f894dfd5a378a896f1e976651e0cec56f1f2
z192b8e079d43af31348dbff2c190e02cc46e78f646d9357694b1e5eb215cb076356ea142768ee1
zc83e2c300402498fa8119f0f3d9efef07abb47c85c1f72e851fab2ae3cd86b95b450351707c15f
z04a00106790213e9e2aba31a7882f94a456ecd53296fa124c64aa581bd6d53d5d02598993fb5d1
z9af65ef62a98270fb896d0181b88f050617067353a5873eeca51abb7f3c585b1ff31bf8963d895
za686fea6533f5a424f6ddc6ef798aeac3686ced17b0ca98960c051be069828fc4a6749ab357648
z2055d7d936e0af3adbdf57c5184826165f02846793d58dd6cf31f6a34aa007b282c81593e365e7
z5c537c2764ea679707c094b88284653f76cfa8ca852817979b29ab0a5e85edb83bc36e5294453c
ze091b91ca9cc5e5a8d0cd36e58b5dac015dc5f57f2fcc71b217b326174b34c28aa96ff4d7612b7
z1a040866ee16c4f4c449265d69b76b5f65dcf9cf2af7bb9e92bda3367cb7c0bcce88a004b381ea
zf9dd0a0f0e3bb377d45ada4254e6c810b74262ec990c69c0a593d4ce465826f6ecda68ad9bc459
z507edf693f0f68362fd51253d48bb07f0d4cbda4d0d81b783a6c23a96e7654774470fab1aa7f64
z7fa5344f4c4c80c938496493f92726cdba8fe6f018f52ac33732d4ca49920fcd5899d2dc247343
z2356b6226b9ad8e4a4f986d4bfe1f90852991adf3f82439f83956f87a205cfe9535748191708cc
z55d8d7448d5fad63150b4e7c37ebe2c4e0cce024b7e22bf91e3acf0ababe106429d43d9a278bd3
za66931a97d4ee8b650f64b7966fe9ea2c12605af050b06e976318eee70eb6f4bec1f6e4298e389
z19b47076497779a07ee102f2d530f806cdf163908b48aa7babed9732a919e4e88b28f3abaa1883
zd06504e9564ea563f262d85101d69c687e34c8540811b86318834c7b6d5a2d788fe5703484d0b2
z90bee10194f62ef017c4a282ecbc12a1541ac2b4587c2072b18f95d63e0c559b20a6206293cc59
zbbdadafed080b26662937abbe1070994478861ca8312470bfa697589713a44645dd3310c456a6c
z6576be66c1925393083e118f1d9f5c4456ede2bbcb510534f5a55addf188dfb82443e775a249a9
zcd1d3c63b329c2d0ece11a09789ec017ee4cc9c74e61390cd1eda191ae8034c214d84c307bf134
z150239748e070eed02cf04af52ccc52754f559b9480214da2120a55732307fd52f1dbcf05340f0
ze9f89dcded8de9be2854e7aef0eded5d02fffaab92e22bfe1bc031b436c71859652c32241dd263
z77fa11ec02eb9bbc6f4e3445f45b48e7ce59ac708a32235fe31ef83fce6f3694ca29b05eb6df0d
z552e2ea4c3286785df1777af70f35017c9091f458ceadd2d79e149d65a6cc4bf51f0f4e2c81806
z3ab0c5f33ef536c836cb890db93e39d4115ff72b68bbfcd30a547053c398453876e4df64b3cb2a
z6e906b30f7c41d56491f287b48bd085ddb43827aed14ae4f77627adb9c10daef7c4996d759611c
z76c659f032e011a1f0e30c56bbeb1844d387d262c7aa06e4f544d12ba82a22b04fd0d2c041e3c7
zb45200293e339e29b58b3ee4a52b2f69a959fe43efd636c6cd27f30a6d0a929f1411d7b440d462
zaae80d5e4a73210a6c25f6ea6220a274b207c5105d5646e16614dea9c20ecadf427864ff2044dd
zb8e04be06288a4884de724916dd10702a010e705d14aac1e8ab518c3a81f83cf83445a065d1d06
z54b0c635573b437184791d2f5b5d7bf0a7216ba36e966b9217ed4bb7095230e4acb28e2def6fd5
z330b7f088345b9afb4999e7f5f2dae4b44b5ab0c0b487cf5e87d896dc0233251fc4e5beb2692bc
z6d98817fc5112352d00acf4fb1a82e2a7bb49f3a11af963ece5f4fce5fb4a77ebc36e4a4227fd3
z0e351dce35547143dc3b78724b070dec970257ce3820fbdf5d0eb68b5bda39df58943688cc302b
z54a59b6082c556730d7271f5ed05fe82e83804b1feba87725efe2149f30213a652b487b8169c4c
zfe450ef8af5dc0947286890e80e3b0e858acc356ec87b1272e505c66f95b10a38c91a777c6d31a
z03e445e3ec48ba2c217748ab22124e2857e3f0ec119d4fff53994d921b0075e4796bbb3e7b7c9b
z9d23b168bd6e1aa6af59cdfa0d8f83d3dbbfb2bf915a4cc21c9ad0dd463f3e530e40715f66b480
z6bc12575c7e71e4061b9f60fb15ddd3d35dad0ecbb37cb54221db9225631275c0f7c09c75b57cf
zda7c9f758ca0a57ed3beec24d6e11a24e9a0cad16d22c5a04f4cec70c193cf64ae145a2485e637
zb27020e2fbe3f49d1ead2cd48882f0c61ca6eee548e8256bd72dc8b09a49f9825bcebb23decd03
za7e0b508a115fcb891709ab738783b3e2e7a9592259ee5199634ba86d5cfa76698c692c4089502
z3ae03d35d834f40ec1c1be424471cb3a576f72eb006be28413c131c9c5d43b6e1b0ba254f47e4b
z00b849d4933a3d28796b8c68cd47b3f5b54963e5e22615b938e3c73c62106c9868147fdc63b85b
z81881eb0ab914ec2718109a08c95d8133d23dba135ba94b1d2b036e86cd290de489696aa5801d3
ze174df446270595747fb981a83acb16531f01225c88cb2005f7815c40678d54baa87e66d2346f2
zfdb695506a22d6946a371b20e31596a33d64b5a823e6d3a60b8c5fa35379ac0a1af1ec47daa8fd
z138b84380de6fe8b0781f4fca6902dbede0e3386f09944fdb642f7ca8da705e04d32e518f4e633
zb7d7fa187cd91a2697efbe15a45db9eab9f72fa725bd0190bd1337180e01c5e981dea4ea18bbdb
zf1c4a59f1b25d2a5623ac40d0e42e9a0f80eceea1f271082fef48b96a4c5bfcb725392f2a9e841
za81c36e1ed474e16570a81f46305dc4ffe941023e34163c4190680b8abdec64291c36baf45b261
z1e7c5afa32ae0ce5bd225480a75b88a05b12aae289e926039b46cc76cc5a7996bafd30a3212fed
zf2ec6403c2ca722da79a7d455b1e203bc06f64879af047491af32d5f51f26af149842aaae404e8
z84857effc7b3f53484b373934924afd9d6e6eedf2a253b6ae4af2bf185f6d063f40a8bf784d109
zf6792c8099edac4c2ea2222d039550ca9bf43150acd45420fd1b539be9d1a43b7f6f0f5427c553
z7e1cb30ab31dd9b8b3c9a7ba38339010ba7950c9a09fac03e23cd0003a7751b9317d2aaf57ed02
zb8d256a86030ad1b1fcb3231624805f3a7889634562996d2bb0c4377f4051281e715f189f21c8a
zf50b4b93f717709472e15e5790f926c6adecc026cd58515a456952458667a17767cb906c3d7682
z893592f92e7e9b10a08aa32b56cea7ec1e5a8860638b314765f3a054081eee4557263722b32f40
zb5594f087a1054e4c399930bbd81f76a14f31dbc84539579bd15ed648c6508a985e38288650d9b
z48a263d5e0087b8fe98331979c4e6ebcb66cc57f6c868d18807c736f4eeec6f0c17d4f3a35835d
zb1071dfc5f97e0d2f77187a2c72466f2c3821db733f4bc0663388a967584aeb2b983a6e548b01d
z43c575190f16d1803fe5d9ef17625036deed56f9af1abc0542b719e178a6e752e3f944f254a20c
z7e76f870da6fa5d4787e69bbbdf945d3479ed810ace824d877fe2b4b2e1e7185a8e7d2bd4496db
z27934bc2670b6be6f8221559ea9d2e2dc369b9a07a73f451b3fdebe15600ccfaf5179e9c0de77c
zfd6455df87e8d78c143f91e9fcfcf957cfea4f285433107815a45355a9417739e1d2243aa4579d
zc6e013d46c3170a0474fb701d16c1e10bea408973eb992eb9a62ec254b0863f224f709910146cc
zf0d27393d947cf6f0d274c51e664eb6f3045224eac845ee4ac044d995ac3497e5d6f39e3db84ce
za659002ae35e473597192cb1fdcea6ba6f8fc5c65caef663db554d3fbe755d0e80df32d22a0482
zb8560e98228141f7aafbf3e6e20696c008e2df746a7b5f3afa3d33372f40a1ef9e5235d56d86d3
zb062f3a9ead4cf2160274443b4026eab9a5d489863d26d78bc1fcf006c5870df7bf6a8114d46db
z311f80725a06b98935084dc0bd65b36e07beeda67285e75d0d95ab4093d32588296f2d07c8ba8c
z1fb8fbb430fd9858371e051e003f46be7bc62a41ad7a8888b49b63b1eb79f288ccc1fd3b7b2378
z4d9455f590e8dc0bcee36197c4141404c5d0d93d233376c75b39251dc61468011d9626696eea5a
z1dd4f8601ad0e8ae974be86a1abae023325aea463870f28f685ed0fecca00dc53c861dd2374ace
zeec3ba5a37b97ce528f0fdb25b8fd1dfa93c32e0c77bb7e611ad7b68ea2383076a156efeb81c5c
zb5d5a58d82dec42fb2a01348687164ae28c6f130e04166cf544f5e26a03402653e0f80aa47565b
z97d3936d4a5c15ebc4066217f1ba957412cd0c208fc8e9835f2da6b5d347e96ecf2edb0e63e555
z98c29a223d461172e0a5d3cc65d5c4dd1304eeb84dff99912c538ea84519710bd19c6dfd406357
z1f764299afb5b466d73bd1b01802f6782d881fddb6262405e3259d6f749d5c918ddc8f98e7bf8c
zab8eaf5bd2da322e8d23d454ce3b037ebfde22ce586d38708c7db16e23d3eb5153c10d37e8d037
z6ba7580999541fd72ff1d71b0b056d66a73becc6e1089a78df62891d5e7f5966ff9a99dd8d910e
z0b20659c0376487b1c27150f46eb3c6605a7da8af01abeb609b6e1ef96c8f86a2fb8930c2c11ff
z547cd30d2b87df6f556522a11b0490bcfe6c39d2ed1f74f4d3defef4041708d62102541691b42e
ze1b6f9df85b5c9c046334e33f9cc49cd9c7af39826be4aeacc948717318281a1084672e2d0a470
z740dcfb429611bf0d16e92bc741942935bf8779636a19dec49651ae0ca84be293874eaf2737a60
z329001dcd0b75540ec73a56b0df8162f8ac94e416a5dc88c94e90af2663c877f1dce20e9c6790d
zf33d475f34ce03bed735129f8772179e26f5987f287fee36c31b9160d01b356dda5117cbf4d5bd
zc0351fe54d7b6004c9dd129140e65816c3e8ac309521072e5348a8875e45a7d6fabcb9cee1791a
z9de7f6f643ebe29ac74cfd4efe5d61e430621f8d1d08514eaf5e52129b662e0a522e07332cc183
z17c2d5cfbf021f389f09c1b07fd6e8f0be44cd26d7eff4b7db79e563ad3bf8c7619e33ae0cd17a
z4712fb8b9d91dcf07e680d13c3e86eb84a9a0f8369e100c3cc1d194672621c2065a4b1a4f10d5b
ze8f64b3045c2551854c5584547a08ce71dbfd71b873973aa59a5dfe6e9f25213ed18b86aede4b0
z134b48ba51ea06f5710d60a7037ece5e97cc2cc675706dad12569725ec44b6b3121ca1996b9237
z40e6ae680da87050b29b4462dfde516452a43cd15d4d1d33bdf118ecb24ab3908356b300ca21cd
z344566eeacd48cd0644f74300c6df9bc701b7347007112c4d5c6a18727110d9926a9455224e6b9
z862954342f331e73850fba3c102a7a1ed5c978276ae3237a9ff0df243b613acf326194c6ab37fb
z1a35c7046613cf88edf85e8d439ee3814bdd2fb73a5a740f8fafc75c68842a5e0b5e5b50ec559a
z0a97d5b7c446d2e3fad2b066c1a20a39c05ce73d12795d8b14bc4f3796ba60869049507ef8c153
z4813ca0f081314ebd99a72c545c6dc4e4147bb34d469edf8ced18b2f3d3348962cc1b4cf59495a
z84603f702c0b65074ff122ef73e8493284df139810803058c30695507631f5752c0f955d4a2030
z26ade7d2d3f52de02cd463f3d284a6f9856d61333b5144606887226b5c41de1f6b6d64b09241cd
zc7c1e8c1e0b214a64daebe0dbce8f20e2cf5319278edda878bac5018901c85577855fd1f409981
zac9ea24e70559f00558530d538f22d56fc2893ebd1766f66bb84574dfef31b76537a02608ef3b0
z187c3d6ef283acd0ca1bfb1daa3c284e687dcd6660b001f1c219af59b794c10b3f5ca334ed1463
z58b950ecf812fa9fb99971dceeb96707738f971a475be70687bf7651829e09af4f842eae7a66ac
zf7c0f1dce748708469dad205de40408bb76de30fab6b77762a213eb252b349459a3d42f39ab963
z7e21c41fade68b31c037f24859a917e2bb08e35f1f198ba473302b04093f1076f19f51eca8f7e1
z82a0ae5e2c92324e8b9966819e6054d1b01b08e4edc7c56c050940a0b02b6840d7b2c3bed1ab00
z539f04d1dbdea36bc01b20ccd66f92ff25c825c8d30c3b5bdbfa50d07ee94ec81bf7f0e4b53140
zbc7041805cff10b8f0683154ba28232486eef2e6f8061e1a73633d8c04a15bcf546a8bc255f9a9
z9fcb505ec3fd5362cce8c4c225b6229d8e9d52004eaab003c2bd393c0f26d7c6a5178b8897f26f
zf2929acfcf3985ace2179bbc22a0f39ccb54bf021544106ea1521562a90064d0aa2ecb2ae2c8d2
z7d7dfe33d0bd9703b15f770503ef352e22456ce40f84091d6c5a39f2ccbc1b6bac0f0e94b5d84d
z1e46499acbe7ff4f7514e19545ef47e0f9c3d51cba30a0c4712b4691a70e0628d51ac3788aba50
zaeb8668ff5433aaae3eb9337b2397c907057d7b82d3774cf7375ec303274f92ffe4e4f6604e419
z7382b3f76bb18e1c028d80f8958a4684808a5532ccdb213bee3e4de8028b92e070e604be4efea7
z7cab5f8efe02b32c07b8644a165d939ed31d92b3fcb15ef5ab406b38112123e12ecc1804c35adb
ze6251e3b2787094237f4208e9a01a435906ff69505a15eb6aa33a4069bf751a443a7909544fb64
zf2417ccb7b5c0e0b70a222272d39ed80f8786503242694c85c500db20fbc907bd436b078e99e79
z11bc79be273f382a723109ad06862a7d247edb33c83e0120ebff9561806409910fe7a421eb8e9c
z092b1b21c7645583066a503f7799e1f1e668fa3e27d7ae915eb37fca903820011167fec18062c3
z04c17ac01cd1295de579f792586126de48397d1f854fc9efa21d5890898386747afdd4f453aa32
zc62af72bed4a0078be2f75c8b867b9c5e2d763ae43e501c9d9137e4218b7cdbe7837064c3b8dd6
z8d157d005e6d0e4ff5ad684a9d7e2c43e7c32389a272c865ed6bc1526052fe6665ac0594331b6c
zfa33cbc540f88a097c2ae6569406e23bc3a99dc17807ff36b92527029f14e7ce991a0dae3c3f24
z9bb62102fa5d8df4e4be4f33c139e991ea3517c5de80ae3934f3824604a5ac507780baa42bc482
z7bcdf2c6a7165efa50a965faae97a51747cd33908f35db009ed31980977147df3436ba7f9d40b9
z5904afb54269d5747ab6956a37c386b245c8b3148eea5043ec0590c1582a4f08a4ddd0240b7c75
zc8e00f013660bf182deaa86492ae7f6a3885fd1560e4bc6cec3d662baf401474bc27b5d0ccc5a4
za5c1e454bc0a31aa8fedf110339f90cb4c8a66725173496f86843901a1de828ab58c0c25feaee8
zc8dfaf9372277ca45a5e5467556f5cf8d047a88c820f24e9df2789b87e200739e0db143869e06f
zff730f4dcdfe584f21e207cd25ba9a26dfbdd7956f959f0e60ba13c687706826b6a6217f167043
zec1b3571b2a75111c2a6ae767ee7860fbaa9f466391983da33edffe1cdd63dbe97909b9f33457a
z04bcf31a9211d4f0b166575bbfd6a1566b3b1de2d68ba35c2cba1481cb40ba96db17d24252617d
zc65819d0fad87d4ff1bb6db62d550918eb747f618afdfabf54597dd47461127a81b01357b70748
za02dc04ca30c5ca416ee63a5cd8660502bc4f1d4e585f13df4e62faf567022757c9e634f614e43
z05ea00d41199034f8ba9745e0c132c7b694357e0b484b913dd06b454ed4f801878d56309f8e030
z1da83d7bd61699bc2d774852f5ce3c301c3a0d6d64862c4d17801a10012fc67ab4ecfe57e709db
zdb5a7162416b21d22bfd1878bda33637b66956382e66349b0b6886bae19174cd09af71b3a72ea2
z015796dd400ae762a4af22c0a2b2c52a9723c3fd06636593f4c2f97b4345596d2e295b6d27473d
zd90378356a5edd11c165fd2fb389de86a83a21a452a25c37d837793e6b9bcb048874429d91a93d
z526d5ab89e9f1dd7d2a5e67f6fa3526354e91eabba7cd8cc05c8c8cd3f49a55b5bd6416e3df802
z2549fe27203535b9657201c0e4cd15edc56f3237843e862e84aad1c53fa35c67bae1b833b03e2a
zcad2ce79ffad87790e6c981c365a59d4b77a4a0fbf0a23108326d75a8d0c20ac08850e84b550d4
zaccc04d12e4fe885a1a2fc70289b8308b6172135c12f4e6b43c159776e300d7466323d383bd73c
z5c1a193c00d420576b4a61018feceb3a0970179013eb626e071bb2908c560f7c642d0446ce226b
z45ce1ba04db5278d5495cf41921ebab6fa082101a532ee62540f5f3cdd12414fa1e97934c9281f
z7644f746d4a5828d3318928b33385f5f07ee213a746f24085332dcf87879c501c16bb1db5d15cd
zda9293494af46c62ff7849a0b499270939a1044de99bfd21953ded480720b8d6ad013c1e445ced
z6ff62b512cdb55c13a0ada09c847eea646e7272eb9577acc11d981bc99e79275f67e47bc6bcc04
zef24bc0a652dd5399c233c4a57338752b836edee192796319f3d1fff8b85144b959d43455c8fe1
zd0c9c1e54c5ce9a0689331aeb7acee510befca100c60651dc44870541b6b5162cbe52381c21eba
z87c88ec4f4882c06c1d576b0da1a707085795d38eb017017ad9e89491e73a41d7e1b99a947a6c7
z4fafc799582de9619af3010f04ba261258659ebf489edd9f5d3bd6ffa4c1a0846c9523209aee8f
z72fa5890f42aee15226b05d7e83be9513f2b56898896047f35a25caa8d7c81b92ec9900a1d595a
ze7b27c136755a638bd8fe096ef6ca665f0c54cb012fdbb7ec2bd3f50f53576eb16ca41df8eb011
zb21b8429c274162fd185bfba99c922bd17c8d00521376b391119efca31196fe385ac5f4dfb140a
z41928b06a830d52d982efad2786b9d122c51323c6ddf54b4f8f220c7a69bc2b870b98491881a9d
z6116bd547743f538d6128c9a2ef8f5625ba5a21abdcd3226539556bb7a9bc200afdad49324c86b
z148a077e42085df087cfbd78d5656ee9e04a3169021ca6c879658094a87ba16fa457a97559aa9e
z97112fadaaf1cbaa48c6b17e4176a4f64bd72e773a4f4bffdf4f27bc0f7cf60eeac74bc90cefca
z56facba974f47f761f71549fccb626edadccd9866b25eb24eb27d81e24161f2819fd31a8d817f7
z56669c15581ebc045323e00588c28fe182ced67f13c46c083c079a571e40c5c6531cd846a9c3ed
za854b846d9dbf9749479dfb0eeadbf23a9adfcd406bea38261cffa5928f542c37e1e1ddda69aba
za3026ecaa4adb930e965c19e85432408b43eb9079bbb8f3f7822a619a73fc8de9bf750e8a9b693
zc32714633eebef29f7a91fcdc3aaefcee0a67de5ff6a2cd312b273b4d8f372197e27ab68e019b6
z601cc7c30ac1423f6216a5d9cbb875aec8f6e3bc831202e255e5d1900ee2531b7e357954ce753b
z4c1b2f08f2e684ed78147a94f25bc63ab04647cb1e643d2460ff732d81b908c40b0631ad1082fc
z686a53d8ea94421b0671ab2e272e766eb91f041c9ef9b46edd62d5792f4081a6fc70e125f3251b
zad8f8dabda5e5d883b3a8ca35f76251a9be52ef2b66fa8ab58d3329eed9a375d07b6f950097a75
zb4cd0b838f516a79d95eb9da962c90ece9e46a6e1c82013ed668f005eb0c6504750ac9297928f9
z41afe3f78d5ed3005782988342aeb9a3255f1afb72b0ebad5cd49702fb072fc44aeaf77df7897b
z4e47f6efc7e06574c5fa2c55e7095aad8fcde04a6532d1ab3852414179605b96ae1c9d272ce0ce
z160c3352f647ebcc11d46dac1f7ded8310f1f047b0a50e2e3a6b921b76df7183a40cd1339cb26f
z150d962c552eb724110dae7e33242eefe69fc36372099fe2a674709bc46dd1d3f900d69067ee78
z8466345c7b23621f3f7ccfdd6f3ac0a9595ce4d03d16c49e6b68f0909a2e96debc528045ddd033
zd5cb267c5401f761b2b2eff96b18ad4078211556a0191f391066f566884b10052593926732c62b
zfff821214f5cdfbd8b3b77883a8ca1a4f40b9b18b24645ee255a0cb3c37d8f3b6da691ad539884
z723819c760cf5df145a5cd0598d6e0aff6df2424b669ea1e11e9da04d5e829bc6ffbd7f71bce1f
z1a48da18d448253ee05d30ee7ca4b52b5ebdd3c2a5a7a8528208339f2f89d7dd009e716ac35322
z24bb90e4f371b44e6655234654b69140790a1fa880548c6413d776b91264e337b1409cc6c42c5b
z24fb186ade749e9872e0f80d30a722fb580ed2a2adeb103a767a41dbd6206b18c2fb1a0f220e98
z4876eb537a16b5618a1e247ef7b047ac2fdd5116a29acbb2f8f509bc287f94834387f432f1ddcd
z7e0cf42ff847c8fb0dfaaa0e17368b5a60b12c417711dc536b0edecdc1d9e259cd2c06d5a0f6db
zf60b79de5f39cae518714daffadd63d79fa9ffa2f6da077dfa742600a0026f15e3018b26600de8
z533b67e1b50afd3fd66dc0b96429b5cda9ed28ebc9c82fcb7f8a43d405146a3b712f84b6512759
ze334335645f432f6c2dbf6d19ddd89dcb3f79d76cf697c4bd90c625d4ac53dfc1ad804bafc116e
z4bfcca82b9cfc6150bf8cb3c6d763092d89699514abadf701f1f182ecedb0b0c46b897d023c8e2
z0f718d182f0798b2e28f07c3f00383b158070adce45f33af0ea00720fd36f29b7ebced10f6ef3a
z787b58c4752eb975027037c533e8fc1df8efb6d8343ea8b7f412d272d13fa37fea9b7067395e12
za0a8cb4884a42c93b1d89404383e89a150a979d0f578086ef452dbc79652c889ac3459e15e6d4f
z1b928879a8a6e820079a6e66f19d93b1c9d2e86b13fc017db16583258775d80ef76d320b41f7ce
z5fdb73ed410b2c7df51bcbe1a68a76d7a836fd990efb7f504dbe21d76a25ccee47bb0369a31e44
zf058f630caae2f430ccf1d9e56df9478beaa75a991c3b4dd6e595f78aa232d9868a6a8e449ec1f
z3d11fe7e0aeafe13c8b96f3b189c555958ef02f9eada0f895a9b95186bc3beddead48f85e0fec9
za558526a753b2d87abd94e6bf140e6711e61a340ef6377dc38d7ab057dec2b8a448812aaf03067
zc2f6de5a2541663c54115b458e9c2558ee7c01c518782ccd2aba74763a20ebef9daad122bb22be
z877ba2a0fe572c7236872ca80de82db98c3674767db1fe52a05e7a7be1d001f586baa7df90645e
z043bc8db9c0b7641b35f7b5e40252331d65456708f85346b21900ad07d03ef1b56a9e395f52afb
zc7689eaaee00a01a8471cdd3b72e5897b1dbf06237cbe6080a21b030fbaf883f892fdf08d84c89
z51e75ac462a21db98f266b23a77d197ea0afd254e2ff86afa3da4f24dbaade34d2576613a27db2
zfbbfbef07097c9da03eab6d62638e0dc002e23148b0c051240b7200fdd6f1dc06675a06c0209d7
z253e6ca8d000b16810a6c2136d933fa3699a663c65d634b9e81111a4b258744cbd5ff15f8505bc
z3e700115629a27b9bc0bb3418d996bca9b0e80bdfbb2a82da0d416d0670e41c5d72903602ea46f
z1e8c01c0efb3937adc8ce9eee0f2df1f0142224f9d69fb7d785968973092311bdbdb7472a795e6
ze1e420175676c2cf7f41d82534c480c4caf7b3b44437088a0be3f930807a31a1ed59dd64bec729
z3cc47bc1e0031e6a44228917c0f32cc1e9ff38687d76d61c2de54366f9c154626e54f0ec995a51
z6c45016ffc6cfb47cd2592eb1fc03404c5a1896ea7001c94db0022ef5e66859d37f8540e9e01e8
zb8f24459b012c36f692ef40f1354a8c341fc9d9c05b40b4b6419791c7af1d700529d0aff2b9e63
z00a628d6e8b4d82dbe6cce7898a9089475b8862d89f659aacf730a5bcf764ce53cab1f67e79c0e
z2c6b9c02936a766d56e662d1c29ba83fcc1ec066b5102baafa7117d4588ad4e39415cd87a74b05
zd68b3bd293e5cb5a38c9a3925137e739bb5f39b1f865071d39b439468d605f29e544898a0f69af
z77d61dabfa2ebd0027b048bf0ec4c91a05fdfe0dd86cd92cf8fd3645e6f154c2e1bdb0c6d056fd
z459ce6ae95a4a6fca4ee7580cd57b1ba71ab2f820ec8aca5062b81ef7f635c3440c562243b695a
zfd2cd0794289d0f45e2821b9ae711b75fc947309e5784cdabdf343a5994b457fd02bbcdfb14e4d
z032f659c57c96b9a8827d3377e6077f21b3876215e2a99ccc0881a55a15f95c132739d41b12892
zca335b229a526e0d582062cf4013118605d8602751690fd9e351dd3289b1d027d7887e77d260b7
zcec7e2287dfdd426b095767fedf49b212f82c3817f3d22d9c31870e026a2c8aa6e094d11674f83
z9a4856100f611f69911faa6274135dc1927987d1efcbf0de368946d40a567cb329a41c6f4824ce
zdf7410aa0662884f05c8dd7be508ac1f602546cd1865af2d17e981ff8aa5714c77504a6c102245
z92895f0300d5c04afbf40a89e62f532a4ef681ad88231b745309eb66476440052b0e0681525f12
zfa78e00e1100b24b4a4ca356f5755a838b0c9e80f4bbe79ecfbdea642c8a83fe2c6d4b3528aad7
z0716c1e650081e0f60cce96245e6e178a4380b52254f04cc29e2551d0b7484319a649b044f3c37
z6ad02fb89557e2dd05b071c1b96ff656327a24ea96c267c84994f38671ec8daf64d8142164f475
z29ccf65afb3d77693010956c8e1e3c49896297c1908091071ca2cd37c32ebe83f836dc2aa2b8e9
z12c12cd0fbae2ed0b3732733b05fd3ceed5ab65645df50e77ec0831dd78e41d41097a990742748
ze2d827dcdae3271a27f65b6582080d5b868f26eb9d57b0c66f02d50353206659ec1bcce84206ed
zc04752a8d24ff6f12d99c178bc6cacbb7a1eb3243861d7b23006f717a6bc3d71619ff4cf6e73cb
z84c154238155ce1ef7a0073311c59374d688e5da13291c56d1e9bbdb04807d461e5803b50c46c5
zca74d2e02c773192acf8455d731102ac361fe5317a8c43bf133974b07eb8108eeebae937976247
z969f1b0e19cd777fd1ac01878be5831cce635ee8dbcb8b2216f5b508804ff005ca62cbae1b60b9
z149a58aa01dd0178f299553f5cf612191280684982da32e1970a85a26bc4f3caefd5ddcc72690a
z9ad1315cc53bc0ba8e44c59db7c7274a758363bcb4982801e524016f8be834bdd21908d00c1fb0
z4444e1e15263b3be32d07f8ba73e6dc77d8e68f1c72c1b76a7991cd4eb5eb7e5ab0b879a00a0a8
zb412fb70a95ef6304a3e576491fe83c58404169f1c9a00ea44bc4a295cc0ce8358f78a89317555
z53ce7fec1929874f74ce9502d511f32c30980194c57ed6c727841a5d58c03011a71526dedafd79
z3663b56b82f037169a86af92839223f922912a8c2818e05988542c43b0bf04acd0f11d27f60710
z7769b8784aa9b72df7ea1e10451413c4b67bdacab0a8f524c7a58d1a27b05d24d1527bb7a84ef2
z735f5e4e14b9b5a4c051cfe47426a059533e8b503140e8f25f040e8d1111d6b9fa4242b540224e
z7c05775db949fbbc7d58765d274b23498d72060c052f4be950b031987d588705edc8475f7a28e3
zb90cd62f6f1b003738c9e9b410f70ffdab5fae87e47851a068a214709fd91e652d91e27d48c0ec
z478eb396bf48e1cbc0312e2baffe6be93e363ff86342e1cc29daabe5d3e707357ab38078781fec
zc4c66caf608a0602e35df54dc936b58f67857f3d4e9ce9cb44631a30a32eee17cbf09f0b05212d
zfb37202aebe218cae6376e98a3f38aac8af458c76911cdd8f2ba9a9784b0944a0f6639c84cabdf
z9c87eff90ee499839c16e386389c58454802726fe6062f2bc4881babf7ab661606d4ff04f350c4
zb0b46c99567157d3c1448e13c296d9f98e7c8bd36f5601fdcbb703c9e1d6d6d04468a25d2078b1
z0c8949a01af502d089950675277e8056b35bfa708863ba1083c716d29544585e3af706b8041781
z2c0133866f79c091be3eb0661fce036e3e5ff2251a4acaaa25c07fca4a30e94dcade42ae8f8969
zd94de9a949b509cd57ee37a0c99cd6c40c03bdfc503a9af088055fa2466c4ac26d6b5a95a0b675
zc22288b2b2c7a06a72cabb83739f335774f7b0e0e07afbc58a8465ffaff1f55f93b94e03c8330c
zc9ff63ec853e904fbcdaae6fc41974035fb7d9c1afcadc23135dc87a52e2fdf061f2e48d0044e9
z91fde2481297b887be4af46fe1def051d112550479d7539569a730567157bc072c8ccf3d5164c9
z6b80eeef290b8e71fc5408742b3f74c23df559aaca5e20f294a95e1dc8ec5f2418ddc946780379
z55e232b960b8f4484fd7ac5d0ef4cd0fa9e5be8cea3aa206384538536318ebc99c09d9d9ecb3d9
z78903e00678e8f713881fdfd981eda1869a46212e885b222117fbb46082de6a8111cefdde8b215
zd7f3e5e91f2b993998e0db95b97b4bf258b2a0766422b98732dcd8c8cc5890b111c2ffe1b3b511
ze9fb8ea49d01f5debcbf806d6389a5e0ef7ffe76c6676c5c6b29e2175174e04072073c496d49b1
z003e461513970e41dc1ee68a17b57abf5687aaa820270bbcd986c8e8e5226146a39dab6aba46ea
zfc58d2db7add727f230a13f470c1b9fe54a6d13d33a6db8e9b2aebeb6fe0fcd2e35447bb327a6c
zfdfccffc385eae1dcedc57969580975b33261f43e42670763d8714431a729375ccd4f29dd41654
z3e0d33c002c1d15372d324ee94742f9067d4a4d844689497612f4dbfa62b6d94c2c4f46d4e0cc7
z88534ccd55a2a5dfb776f919bfe9d77be3255a5df3426f63911385bf24b07578d46fe66bcd9bdc
z8b0bc15f490860b7e753282fa24794afc8dff92a9eda8022a2dafd7ab3afa1efde1915093f60f7
zb8cb8422a12d52a8a749f874acd4d31598021b7c1aeb526cbb7e33edc3b6a611aa56ed8f5deefb
zd71c468d6acbf48e28426000349bb582e69695e70510d500725c54cb3e7de6d219a47b954b6b6f
zaaf35020bce0ab32997b35470c767c1bfabfbff07f5b6f364adb77a48fe29a6cbabd57c6693450
z5445480a225e1a688472ddfb2923df8dfcaa8e6364e3282a296563b16f3863d6ba7a0cfad9ba04
z1446fed750e46bb60107d726eeeb276d37bf8ff34ba1294e3459507751bd49a06c97f5c86c95c4
z66371b06c2f677cfe748ae27af089c7a24b2a9faa40affd1f1002127574291a0ff24590df5fb2d
z2d6601454e617c4da7289c4e7bb6f3d87603dbd7217189490e8db7998d33a612d3547aa2ad0a6c
z61d8aec15dd92f9d205b2cb04e783373f87c826bb047426f59b9167b9429e76e94ada997a1d0bc
zc242ee144c5c5c4ecc92d7fba89967a2d86407dcaf7652fc5fcbbaeefd74820edf9ecd15afd1b9
z9cfefe5d6d3cd8620e16ce5c29603258e58f7731299bd0c50fd930fca7b5ca9791cd2c1d9073d1
zfa1774f9161d2514a6142dccfc8891e7bcd18886127f2b709a7e9878f5456aa3ffa90339a1c712
z12244bcd2012c4c5b31a603dde5c6ac8b971a31cb11bb3a5c3fb9d0678c1d9c4d1f8c5840dc5c2
z7b8659578cfb76bf90bddbc1307c81e5ff1f03362fcec278a1f820699c10ce5d757312fd1c143d
z5f798b520092165bde6b83ecc37c98d57db394923a7b77a0e19c690c77117b75ee0b7c9552c928
z8d4bdc729db97765bdef1a411524e9f4ecc0e7866d25702c628cc39c9acf0c48879cbf9d82d302
z40eaf56fb0485139010502c73b75f86079bd4e4dd9328f09d8c5ae62b2e45f27cee6382180dd08
z58057128f610029ed38658f08f63d73a0dcd32eb5762ca4df836a37f977990fccf5ae2285ba794
zd0aeace4efb7f207769d98a2c6f449b020a0ef9a4d135033623898814baedebf822264de689a43
z3aca815058bc291559892fcc13dc292529ba81c7397d5ebf649cf3cb9da0cf0787fff810388e90
zd78adf715197424b5031ec55b630a7b01381dde80a079cbc2a0e43b4a21f148f07e3fe0c69397b
zfb78a9c0e2552ba99257cea4d9749d9caca25ba01f30f83ee633cf9d05884d2242933a474c00db
z0aecce29f9e211d3b4f0036632140c6b9b2930e8e7c3ddb2291c68470849c38d136e2ed8d15ebe
z6e77e29d790474155eaa423e4d1fd7a137b96bd7ffa9d03c5c8487c146b12d7594a069058d70f5
z05059cca0d67a158997e281b66a22a0819490940f5b9ee8e9c977a16429adcea10fc166cb656c7
zaeff972db17e4eba9088ccc61a6bccb99565d4062b3780cfa641f395693401aff46ba123919898
z345f356e5295a348d56e440560de7cf8b01f3a94eda9d010798afcae981168cae8167211725e21
z638b37a04b89dda1adf8265d18c8bae76433ef5bc8157a5e5f26a505688b8981d3291363cb5bd2
z1f9e70de956897865128328cf9f89d7f1e7575a6050ed899c106524387cd82f0f2cec8941f5b12
z9f9ca16d7638d41d47bef24fea4ea3326234bbdf13ae87558aec62d1276acb2f9e08e0533119ce
zda2f36bdfaf51aef851d0a3b31030a16c72f1fc9b79a6bf4003879338cadd506a2ed6a95b87cfb
z1c99e3ce1d761254b6d73053cc1c88151d0e69035f31ea8d6d2a322f9e7de1455b30899792c8a0
z6136f490b6faefcbc4eed890674f0081c33694872ce91954b9c6805730f14d29a324299cb29be9
z575206a6ec376984132e57909291e31f27e48e8613f7a1c71575dc484ef6f177e7dd812ca923df
z162398faf62e5e8caafc7b75b4d86f3420785937a0fe365c78e42b57b1cb724b42c87e7f04b21b
z01892914316bd2de796b0a6394478fa6bb46747a9fcef1e1a9c6d4170bad754989ef1f578c9125
z77fd8800168d38cb097df9d734f1ffc19681e22751f1a45ccb3ce6f1c1aab6e04463e047a18633
z7d6f1926e15ac0f3bd170c084e49c1e1a3ef5d9a3e5240104d14d27cda74577b21538b8cd26918
zc2192782a6767c8402f23bb841f1c007ea736ee7179a81a63a7053e746089ed028ef47406503a1
z11502d4b72cbe5eb8704475cdaf06cfede993754fa3cefdf8ee461cf7b18b355d450070b59a991
zb49f31ef0f267e018108227eeecff4dc379c1e278c7571ea52d6aad9c61adebad4c5639fe3f275
zad48d6d4b9f96a10f464017724e4d70b6e7599cb7646e5c77d454e9965bc4bd0a3efea8961f5be
zcac3090d195d2bab1ab8f6a3f070c78474419000ca1d9c611a1248d9d5cd1f26f527c79a0da4a5
zc91f29e7fcd0c005ccacde16465bde636af505f79feb659b52acf48255b086bc12b939b56956d6
zf4b9f0ce22452cee15beee6a76eacc97705353ab92fb352577e57d2472c6e84937f2ca43dd9205
zbab89c1bec37793219cbadfdd63441508369aae9dec968ffffb4ded43b04b0b42c8795d5243f65
z1206cec985b81ec4584216e88468648633e48e8ad28f8409ff9b5d9121c7b377523d7fef678ab0
ze5b25695e373a112f22e84d9eb155a6e90e6399e2af6f01706298e357fb0b7acc6639bf11b70bd
z40706a00ce3783cf10080b48fc13205e1432e9a9814b979b2076633626af7ef988ac2181cc2e56
z582c9d029ab6a2b78bddd075bc22c3d85f749f43a8466f934416172563c82fabdaac2ceb8e830a
z28b1d24c1d3262dd45324d28276319942fe2aefaf5c2f3a6916abd21cb692620c961804af88ce5
z11eb52338fbfad48d8755f52e8be8b26ed588738b38103a45715d1972b40b4633e5e28612756b8
z2d26bfc77970c2991117db066481e1c0d5b6da8be0d06647a9d2bc95a235728a28daf2126fa873
zcf0342641766731d56f9dc95430b140018cf0919beceae6e3b94ec607243e2cc89f3b95f30b4fa
z63c4d13fab54fe1cf15854b631c3fda734e055474dff33aad2871deeda5232fb50fba7cfd89d4e
z8869ec5d4a61e45f049e8b9740e19e3f63f6992f95a968e7b0a77ed1be3b16a24b94afd026c21f
z4fefe29049636d4a054465b349c699e8ae38acd089854ce4dfba9ee24010c3449ff32376947236
z45d30f3aff205d9731c32e73c12c4525b448fdf274bf0205fd6d0c675f295b3f72fc9ad6e5e71f
z39776279b1e7be7551ddb4c8a3b843499cade7cfbe13a0f585d6f9cb6ecfd4584f3efb7a78b0ef
z58673840860c2a18205b7de11c1e68c04b7903d3cd3424687d020571034f1a9d921576c8efe9ff
zf37b334b54c53cf83d38bb3d225c5c7a42a4fc352907cbe9d0a8fee408d2c31a1f8c372f13f3db
ze7505abd8fcb90032707e25c9be9660b5b663639b0661a44218fcc6bca663fe07b67a068b079c4
za2f38d3e69d9319dd0b8df28fe32d99910cbc253559ecfb6bd32282d6885d8bd03dae35d9f2f78
z24be292a304a1a1e6d382fcb0af6b06b31f41a25b3cd811ae8014df5c938a02a36cf6f5ceb352c
zea3998cc2d169eb65b60cc1e02322af71803202055758405c34131c8f1aec1a1820e7b10c08f55
za10fef4997b2326c86aab27053b60165c6c869124d048d2bd9759b905fcb925a51aff2d8df552a
z227f643f2b33832736713ee4d55d7cabf574532754953de4ef9c82a66492f796cdf3d281a84442
zfa2cb1916e3f819c220eb8a669deff00b4ca60dca82ab68d816b48b050a4bc4cdc76c2b8f828b9
zd91b06fcc521deccecb5250b9cfe877f4e8d9ad0baeffaa584413958919194de1f8998fdf819b0
z180ac77720c7f51587df18400a067f7e976ee8f24ca95fd8270f6227dbdffc9c9cffb737f2374c
z3a598041c9d644cf23c5e54a9b95e6e2e5449fd157658d68abedf231167105582d18122f258c09
z05b82b188197ba5412549104ca0a3da50a6a6a41b88d2fa0744b5ba36dab180ed578c074a12f41
z4af08a1b16a0a93e3b8aa6bbda764bffddbe2ebbb2dfbac76f541c7514be36be3e6bf73ef8946a
z7a65c8f1bef8f9ece5261ebfb758bdc20ea5f3407cd2beeb8d1b002216f7431bc2b00f4cd1cfd6
zb0b24a31112a959fbbaf08e974329b311b1f835a6ff1c5cc67e826e9e4a25840be145d6bd56114
z7bd6acc36ffb02cbc2473c619f3d043a85bfa0a0e5cc81b9f3c803a6325b35ecf1801662bfc51f
zc6fcbaee13484793352308d6ef083856c6d666e42aeaacc252027ae813c86ed4683c48d29a144f
zd7ba5d8ef356d0990878272d5b6dc4a4ec116542023c4e25068001a3c338e9d2a2db1a77b4155c
z8dfbab7899c440bbf8e2c7f6644e9a6bc0e27a10ae18ac79f3b4cd94f9b2eab59abbec40f7ae30
z5a47e313aa11f50c2ec60ee627201b6a2c7e0a6b3ad81fab2bfe8532020f596ed074895e3c91d9
z4f2db5b83cbfa7cb908bd6cc6f2a256b5003b24aa53511511c316852d6f4bdfbe949b64d3d799a
z27c3c1bc7c5475ccd1f12f4d92048c94a5a93f0cd314444380f487b28133d64b4e8c1f0fa872f0
zd1d386fa67a00d311dd2c3e463f8f5f2b4ee46383cfde7c4ff72f65ce96445d24d88f1e06a1633
z2596e0ab7278737007c425bbe4799ed8a8b54f5fe9bb4a0887e855616faa54988f780d63ae7b29
z96c2988548c436b60ec80ce507aa58d304485939ab1c040254cb6804aea27105b0b020573e6ff9
z91a2e7dbdd4297fb74d29f337a39bc6868ad651f31ac8bf4e8544e5a542cf7b987e7474dc72b73
z97a52c7ab797d09d0210d18fbd0b195cc295db87f929d4cc3d44077e2ae1426e55ffaed0d76d15
z4f9570d20b427e6c75c24fa7f22e87c98a084c1843eeb2db02471207545ceef555ee9376a059c0
z7a0f646e36f4d420da8abd18061653361dfa9278b10388c81229728d2490438cf82197093f1f4e
z925fe373899db0629af5754b1d4cd0714255a7c6e82b63a948a6157500cd163868a33b471445e9
z75abad9bc2b3c35fcc7d52998f0f19a1f983dfb0790716757a771621d4715d6e8c1d7ccb508422
z46fa2724615d09aea717f145a086c089c7ff6a29fda12fabcfe3f453e2fd5a31a4d8b716e02b0a
z271d090fae27f68c03bd9fa60db8c32fc5f6b517bb6d7fdde7214782b0e8fa3298e9faa9391de9
zd5a42ab5ea90c602922a268f1c1e4d2f8f6c1126f053c4a9644108b1557e2cb2fc0d27f856560b
z94bc36f34a1c8a791c7f267a89aba6528a04659bee0b28f3f0d54b7a466d8f3d7e918fa6b8c669
zbf92cf5468a79e036af2de1bb7ba85b37404b1143fb5202a31d651250e8f8b01184b9b307c3e76
z47f1be8a883ea3add50cb48dbbb3498815838f6fd64f8e057040141d40c9b0707cc6252a78c488
z326e398e9c4eb5ef7f7b289b2a62bfc812b519fc6d9a362b2a07a2b0baf4dcaf5908a19616cb27
ze1c620de569ba6547b13dfebeef35337c8503a0b12c1c615999540a46e3151f531255e0f9d08da
z700e2c8331c0088925156037d67894ffa77ebb0f0e17da0768a4f4c49b5dfab1d2dd9d48ec2dd6
zb9f5f5a8ac5556c36653bac514fd945edc20a9359d0833ce25222efbc0bc1b43e7c03ca87c70f4
z25f871664acc18bbab9d44a20b1a3d3bc2cac404e5e2d15e55d76d4af5a8ac9151b929b5a32d26
zb34f292ff158ecc1dae3e8d52c4ce1b69b6092a0a480c99454b3ac1f1f59c9035b1b026db34948
zc913a2587b172290ba2a5ddfb1b9787de0d8be95271c0fc7d34d63b119151d707673ed1daf54ea
z66b14585d5cf9cd82dd073a8e5f73683588a704c80d0a052b18d4bb3b4a8e7eaa5a8fcd7d248fb
zfa447ee4e7412bd21f6af86bec4dc42147647847067252718a804723fbae14bc5e2be367edfd8c
z538a4ef3fa56c984708a8cc30f2b23d2ad3356bfacdeee98abdd15f97df99ada86274315b018e8
z8a2d6509a2b72747b82572fc0e77f4663c5679c5f1a1f912860f208232445313d95c0ae35a4eac
z1e7b106b2f6b726c04b2cddd4cc63caf6f7e2873f14ce6f650dac641f4454d6a330ead17196901
zdbe763cf94d01f8809844260a67a3583640d676abc925432d0b467364e809c22f70ca30da0ff31
zf9de53c47863ef321547526fb6c1f71bc4b5fa94d710e85cf920c198dd9b67ec77934fe33343a8
zc41bd3bed9fcfd7282f86a12cec6489a60e2475d5d0e44590139720e4503e74e28cd626c5a8853
z491c7f724014bdffd03a903c91ac99edd8f375dc1a4001000a73ac76a919ad4fe14b37ecf95628
z862b4a54ac9aeacf94ec64852212b5c168f8c83947f460d4c32f8e27238791edee00eee1e0adce
za92e0fdfb9b60222cd302430538e47616e3350333e85f356e50dcee662b826dffb0edea92a437f
z44a77dbee7d71ec52b72260139f9cf62c0647533c3b11d3339bf2b0f16ec24aa01f598a5d70e2c
z4e4ef735f1115a5b2ed3ec15f2f91120498b23bde26ceeedce2e12e9cefb55f2ad427802b3d0b0
z2db14f2a1c590c883ec689ef6082141e390d49bd4fdb7652598c21193e5b99019cba6aea12cdd9
z7e63e1ab873e9e0ed884027664cf7ebf197263f8dea76f724de435aa71afacd68a0a475c2b1db9
z0565441ced3b7b19faf06aaa7320523e9baa3dfa007d75c7b6ee27f536f25efc486f192c0b1d82
zd64a62bbe2ccd1bca373b4b5ac0315bc76d56905011ca2e2c891cb1aba378e0ce7155612ddf473
z8d738dc40d2b9c7ea3349306edfb3e8b642d80033bca9001061d3d74ab38ba497152e2357d1af7
z2044e7cf8ddf4801a24525093e78a61867071c41edfdce676ee2a1e9296f19e4dddf1458cf174d
zea563007364a89e95bb37b2434449ba76698b448f67e0b4c9a2d9714383f6256c27f8bd5e2580e
z77ae5a009182160d24d401ab8a8e69475648eecfab1de15ef719d8224b8af87905536c284a84f5
zb1e857f1fbe29743edfc5df75f5d103abeebcf2d623b546a4e1df424326c153b92bdaeffbfcb0c
ze6a8c8a6540ea2e35919514870e08a4313d873fec65d4749d505a5ec414a00ee81180245c400bc
z74bcc855859e3dcaab0f80b786a02f094f05da705010305b79b51936809a8242fe6f25fc0cf903
z7f5e93fe0d847e157e8f97a0ab98c61db6f409338b6a248acd8ae0cebc2c402dc6ab4052bb819c
z610e11d9dc3e5e24bb183d461580453b74647ba8dad7f5d35ad71dd31eda8ceb061285670cef6b
z5718aeadcb0eaf743cca91fd3fdfca4c3bdbd23a75cf25fda0a02ed33fa518704853b7eb5c1c60
z640e9c36f5f3c5c004c265441118afdfe350efaddae9310d91325791b4915a73509b9b3a97b8b9
zeef72845ecb01feb21a121d9a014643c37f429abb41952fa4a3d040666590b8a90aedef3a7890b
z6ffc4d14672655db035c4f37b5d5a488aa71712199ed0f15696aafb93e9855abbd09a6fcda54a2
zce7298e228098ec676aa7b357bb89124f7e86380246a126c2a5e5905388725917c01eb2c08c98b
z07b016f96719528b49677f531919ba55c9880698da2a931de5b30491cc3219818167102b29bd75
z15251f61d487fe59e86191ea82f9b1a0e087a367131808e6f9c2f31534d896381218072e779b27
z0a7504c4a30657b76b8220554debf06a1bdd44e5938ed88c726b9062bf076ae35ba827bc69402d
z35e7081c9ddff05951fd4a4a0570c8744b6ab696a8ba80739a7fc0f64a57b7632e5f05d1c156c8
z27cb2e16365ebc11fa7dc84e180a0a1eaaef4436ec0c3bb10b328de5709929ab3f25531bda9d3a
z6ec0067f684fb89d991460317a71e9b9447f5ae1a38efc563f92926af5c9ca42006ea7ef69b133
zdb50aa0bcac55260efb55222fe512da2eb89a09ab5ed02dc59b355cb76d05bda234594a4503174
z60a2c6fe14d389f4dceda0628c4014f6702b12ff46ad23d48b96db0ddf05c0e5f4f90b48b5db3c
z6158dcdb6a25657695638ed059656d98d4008d76307d270e20abbe5489efe671f6e8d61dad4b3f
z6ffee81918d6e61e72b8aec41b8226bf438f212e3c6a8b1df89512cc9219aacdc1e967fc16d6f1
z335e8286d0d4551acca7b20b15a9b5b83f037eb9b0f7578cd3da607318278e629fadae49e3b2ae
z05a3d9e30323cb875188b378a1bb90ddde763788691caae2471efdf9e564ee094e464aa1123e97
z7eb4931187f62f21c19127967ff268bb58367a2059259624c34d29660fb7e014775d9adce57121
zfc087276ae22532ff9801bf9e8cdaa1c7c8162172cfe1d244dcf343719e7b38225ac88b9b3de0f
z8748c33b1963dd0032f843ab49a60b27e3d67191cc96e24deee41a835c8a310bf3b4c74a738991
z1774cbedfcbad8037f6bedbfddc2fc9cef7d4028b7b62cba64366678529d75219e8381d6effb06
zd5e1a60bf409659b6aa501364e435bb6fefd4ef1a084471ed9bc8c95993beb5a627fff0ab30f39
z4d13c47f79f2e52f9cd8857ed6d2caacb90ec2c1d3fd7eecd1416261b2e1dd3c73a302973af3e2
z82da6b71f6f38508c653f066b7a773ef932b18a9d75f088303108e163e26145618684597b89fea
z25c1130778dae940527f3651dea5cc844cf6203420ded24978bbdfe5ae7ac3b5c82f91e65b0ffc
z43e7ae5f9dfc5f8fd0ea32686919f5e6a8b1bdb90aab84bbdf6be3a7df382dabfb7728d91ac73b
z5685d536b0902bd6b79cac836b3d0f70a2eccd206650fd3c70a3887d0e657033920ebc9c9e1529
z07eb6287a6ec1170b4d31f20bb761391f9b06010dadddb4ca4e0badcafc2beea58fddc1f6f9809
zac750efd1c6adfce0857849bd8bd8ec5fc1d2481064bf68b9164c4731102993841f68a96d4f84c
z438de9ecb6639a4e5725174db8f1ee24b95814314d3a58136475d3411a80427e37bd4e9a579afe
ze2367ff0e03eb6f35c6a91b46b5a9bd63dc098cb06d6bf689d366c024458bc0a8c242f0c93d0fa
z5b06e990307ef095bf825148cc7b62957fd992dcad69eef3a54ce850adf2fa5573942a61010979
z0c95cc1989b1faf26a8a5f1f40e92712c2c56a0719aa38a38ac2479907e8bda331c94b0f2c4781
z6752dc164d8791e9edcdf1af67b40d9782d8a46651afbbd89b516b46fb892611d36d0b513708a2
zb5d8a64429451ca6df4f2483e6a4152d081edc31dc223f237b868e7fc68951b281e1dc2e8952a2
zd001be6ab6630f4fd3b391e69d524b34f60171e7e8cb4c8acfdf1306e5e8633809ea9a9c551286
z62816b5de9db7e9a631ef5623c1f63304b46372c8a841f598660d0832f3f670a99099ad7686ee9
z00082437071e81fc27e3b25835b8c8369322cc3ef2974d96c9c3befa980900da11e08d357b00be
ze7faff4c31c1bfe69d09e932d2c446460cc771adbc8c9a87ce8dba9a338ca9ce630a15d23050cd
z7d98db8efb5391226a5536f2429f153300d51f054eafaf0e10589c82c63573079068d4dc158a7a
zff7670247a4326e7542c5b0e429dead12b9d57ad5a4739fa3557e40a662f819e5b64515ed26855
z39a78cd2996d83636cab8dc4b385df65955628ba95f11896c53be655f600de13e3278e6fff6e76
z55cd028aaefe7a6288dfa303ba9e1094417c07ac5379982d950d243b6db648af680f10f2fd2465
z63d094096fc3a1fc5357e50c795b82a177f8683e6be0de60bf25dad1de94642d2d8816d3715a07
z1a7fa82ede1ee4b44e036b647cbb47d48b98e5062ead77cf4a037e28e7e9dc116f3edd2f855bff
z7785f888fa447e14d2b21c6c4dba0904ca7445636b61fe544c54323b7a5ed4b15e70adac418329
z6db3faa697c09067e9f50e0691977eeef2c79b1d2bdd6437977c87cfb90e47bc764310c81f65e7
zc223ed091b151b1e88d4935ea36a07ac687b125a93df189dd424b4f3c746baa634486f6d0a1dad
z38e3bf1a1589f18db39e5f7de68dc8ea8208cb9dbeeef38ae10857d572962240d3cb189f816a34
z2ae736f8d1cb25bfe4b47449e529feed139ac8782e6f446ac3a240f6f83f889a7a6b696be4c31f
z5c2b71c35f88c8d09b11d7e829400b9c765a9ab7d75c6c8193af3aa2485060955eafd999748768
z2da894add78ca0d9efe886129ceeae89d8d08b5960837d7977b68d995779e0040200b4605932bd
z002c79834031f402b3d086c798c1eb1873599c4eaff37caa5a1f5a1f180b096359088cd946326f
z7dcf1750cb844864b70d4977e67bd1287189be5dc3c4a51574f86e2e69803c7205df05fabf3082
z8cdee460b6aad84794a8366b39b8e421fd4326403f8a1235441d9857b9f693f5ed10e5303d2bd4
z4cde984ddec2dd219438c9e8439c4c3ee2186606b60ee32808e52a1307378e69cd274902420eae
zf4ff8c430c4ad35c8a55fd62c21100e917983ab8beabcdba0d55c485e076fd977b8357d5d5b36f
z1a02161a99ba6ce27591de1a770d8f5251ee52e23a800142ecf1131f80693ff2a39d125ff0015d
zffa2e9a5a05ce56aa336bc7de3e8d3b30c79bfa3597ebcd189b3de9bd100478670ebc2d57e9633
z2faceb3e0d7188143586cb12f551083d4bdccc1654e65a38885e3535b528ed7119daa33c1770e2
z06cb05acedbffb38319f100ef0ec3dc47d9e92a043f5f6451a63436472b33e26eac3d98e9527c9
zf61393cb598595f8dc5622500d3a4c3aff759c9b8109f716d3aa364adfb0094181c005588bc9ed
zdd81b722f33bfc0a2cf10bcbae1deddf267f7622dc2fcdb3120333202479b01fffe8f659a23e2d
z2b048929a0ebfc1d160d88c3209f6f3c9064e49391a8aaee468360e75724ef63147944af6c8adf
zb27e3a2e9cee6507dd1907f2eeff7874fb9daedd4ad7a37912dc2a8abfec3305836481db8121f2
zf673763a34b00fc42c22aca340d26901c2c3289571f435d41f26c9614c433a85a7f9185749eda5
z37611e6f26849ef92ba367be9de4e03a734ca4c01067a101080a902913c112826e3385489616d5
zc709cd0667dce17e24d06b0b6cfb377dba2fe9e11485048924f10c0daad432ff1cb869756ed025
zb20ff7a1508ee993d7f770a53cd9e51f0657e0d59ccba4878f2954d6c02ab9ee30825f2f01346d
z4a8d7a8ca7886765ee6a36205faa2d528505c50981353a53a681ec142c84ce0e3fdfe05c35f28b
z88c71d8971b845b6d4b8c9d1547c1d8c91ae905b0bf81c19b5f1da91b034670502d85a81e89aff
z6ab1b4afd8052026946020584f81f847363ba19980b2aa2c150e1e2790d1cd91f67e8aaef42fbb
z65391c5655e865b2b1ce3f7f4ceae6539b2ea005e64d68d259bec6f7485675a3fe91a3afcae5f8
z149c1e7ff9db48af94d696127873184d06195dc9dd0f8b9c5f1b6ffbba4330ee91064667a4b63b
z68f681bb7c8f084c8afad3a02b4d8f14124f9928d1d7fe3204d9576fefa79375b696357f59dace
zf71154d41d746b3bd4624c89b4dba43b9801cd00d7240b1f7347692c8f59b7f748f95ae5af4549
za1a8f331309b633788097d013233c8a37fa1688725b16693a0fd3ab3256ae3788fa6c4e1a843b0
z4e83b3c04aa5829f11958f47fb714566c578f1d48b39dddfd9cb399e18d7e13f925d25fabee436
z37eb9e8be7cbcc88e1fdf56062990d7d1f14e5c99e76e31000e8038a778b76e98474cbc709ff8e
z3c2ce099c4fa9c990e958252e3ce4a3e57804c9d13f11024b2629885adb71d95416fa1ce4d8b35
zcd7793ac255fbba49361d907a78b7c2e21b07a19108d609c729fcfba10990905f4852010ee800f
zd2a54dcc2343d15dd6be6914eccb8c68ad3af6699e74befe2de5d8bb4ac6ba86549538fe765c71
zf7e1a5b811e818c7affce94ee6cd19e2cd95326ab6fac9273d9c4bdbae40c06ea208a0672524b8
z6c830f3d2d31cd5b565a81dcaeca6a92d96c1e990ca62359f10bdf4391e19dea4e3077b8f48eaf
z40c656091d9cd3779c849c4c46fd57a4ae1d3fdfe29f59c76b25dce362ae68ec0e0b7b78ccadde
za7b270a78d15f791de538da323969d6083e7688898e71fc15365dee67896297f9bbde8e2e94772
ze0fc076cea2374fe0ef415abcfde28b2e70b5d2647bc5fbaa630b2751253b4b0faf74fdbc9da4b
zed1eb33df9bcfef7b431e5e21a03f57d0b42e76a72fae8641b73b64194c95ea9333430593bdd3a
zfddd3847d0b7f5407eaf7bba503d294ae367d1cd354d6fb491acddcaa3a3b7f8319b8266165e5a
zbae7f4f7c2e2bc1f3c1ed32c577ed99fc39f051d1350ed62a3bd5c2247b254492a75f70616b365
z6c632d39c99ecc615c318069fcc8a3b690e4d3e003760383105718b5f7faf6fd6ec7288a7aff05
z89b1e6d0aa60b6addeefc954cb0ce68fadba1ce1197ffd4a1fd14b044730cd6a9384e3461d420a
z10df38e4d3ffd234d46890b8055b43313fc1d766d99d1c083b35307518894f9e13225b087bf5a5
zccab192abdc3abf6777a4205622da096c2d1fc225a5313e802ffc8a02b9bd5bba0b1272cdb1f45
z02fe8f01ab451afdac3887089e90dd2a4b8ce6fd720cdff7c4949cd634c79d645d853a505e4566
zfc60874d5c2c8fe477b4f53166ee406d5a7ce37eeffa475bd285f0e09bb00610d867cd5534a294
z33deb6f51bfc477149624385004ccbcd75e0719652f76a4d8bea2c0cdec573488f6ad981a599a5
za847875e5441fa6180966c12b1b8fb5fe2204b00226928deb6910a90a748fc57833a674ad5f393
z725108b807dfc3fd80ad7a5c694b831e9fe6e9656f7b50dfb7a5c9c5749557bf383a0e3a76c216
z88b03e92fce227861fc551c6878524f7e41403f53ca73a6f0a2f6f135261a5bfb06e67339d16fa
z1d4a4a8a2b9326a72ddd2559b5399b177cd7c9ab186296f32c054deb4e71371fe006e00710a4b4
z1ff0fb1772680eae946c5a4d14d3d0a92c48c01280552dc38789a53af36b3ca7dd57a26042faaf
zf370a6c1f6a594bd00d1d5272735c6bed9d6155f1feb0ecf6d6fd5cef3324f36464abb99146c2a
z418abb2d4a01d95cd2052f5d0472b20aa381241bf260ea4dc5713b80d096957edbeddb24dc4043
ze9f38c37f583e3345c39c4d07728ddec0bce992c0d85b6405508921396706ac0124ba11f012368
z0a2faa14d1a11d4c4a93e57b684231875e7dc32121adc20342c17459d91dcdf5554e9c0021e72a
z05a453bdf60acb52dde8f9d308acf3a33a688cd347cd5a90b1c9109b9f6a5f678cdfdff9766c90
z8e68b04b1c232cc72692ba03f04bb09801172402c40723c544dafab3a43b3f018d95ba2b0148e0
zd00627ac43615207ef474aa978544cecbbc8690aad25517039802bb309f91f4ae6db2dd387d58a
ze723815be75cda4f06fc6fbd189c568390807ded1d5e8f69cb7a9bfb89d1cddcdf26526aba4042
zd5d24a0de101cf63ae32d02c2244d6768a925590aca4258c53341113336f528db9719b2c422f50
z4ce1e9380b114d749c60659680b75a5f6592a06b86240db34f40ca787c364e1f74c677e7b4ce69
zd8a1654fed928d38e5ea7916cb9355bc379f872a6beb6be13b6e2740aa0dcb57b66574370007ef
za69a72514e31cc5e178e41b9d08ae91e9ce80ff6eb24d039f62194fb5450714a696a858a9a274b
z0bc309b05d58201214277092ef4683eefacbad6af3c34009de11ad5a73cbfd271aa97c1346bcc4
zba752704ef2684b3fd3bb687e464b2b6eaaf9d24318e9898daffe72048d374060ca48460b0ffb3
za0df17cfe0d199f637604a9cf84c5cf33b104bd9c85526ca97d26f8f37624a36a1d7b5cba48fc8
z153da9a6166abb3c3eb45a16a50c81191b0e32c9f6e61ee673e1a1479fd0244ad6190e574fde4c
ze247e2eb5802802d17d5c534b3b34bc53d4867808f907c02b53e3c94841b91b0b4bfb89c8266b1
z04883cd6ca984710c8186ab8ae499d4e4fca7fc920237182294ed2e6af456367175ee4eecff6c5
z025d37e206948ad55f06ebb150ad84c63707cc2ddaf7750cf4cfa58da60ba3b88cb60e35550b30
z0c5407cb2192a39ed745653bd1bd2a0ffa75fe17364e8e92e3a91e14f4369e8234a87be89d61d7
z9d74ce7821a905e771dd6f2527bda51a4bba48f14bb881e348bdc3f3926b088cce0a572383e24c
ze52ab2c1cd00c982e4d5f9346a947a3375fc89160e731c0c4a9362d21a483ba1fff6e594c2b34d
z7f374f32f9fa2c275dc9c7a6a96eb4e866be2d8e9018f12520f9417b1c77256887b05fe3d23acf
z907e3d817add9116fd64efd92593da1263f19c761c658768c9f8d3107d871978577d23843ae4e8
z116d5b37e789187ba978e79fc1afc858235b41ff5e18e9f7eb0a2f3e4a2d300bccb02df226870e
z002e93166dd117454f193a2615afbe36e68dbeabac8247f290cc1251f3d12f7ff52ec60e1832c0
z6e9343c345c822c09ebc094bc1dbea4fa6309d124670d1471fe31be145632a99c72a3f859b9511
zace008b3d0cd16d7f2a1b225140e87d31dc71d8820595176ad49fed5acc73dc46d0a8f4031c73e
zf2738b33c3a73148da04754363dc58e634aa0d8db8c14deb9dab70edbc3572d5959ff3544acfec
zd28ba5cb061f40dddda1c5fc7545b48230e28eb8812c6df1b6a326b7460da710624bbdff4ab1fd
zdbb5a3490f6904abcd03251d3c40da4511fca77cc2c5588f538865f8c4342f780693678242cdba
z5798b6d2d5b00e187afd93455b6e65119d47be6d97493307df5b2f0af1693206b2a8812800c9d8
z1cb0779171e394c7dbccf03764045dc4bfd05df684c07c3d22c59d50d1bd491a15391835a3b35c
z3e8c9346a55b97fb51c9bc0572ec2ff57214f696f4328bd57efaac3169c2d3ffbad2a3d0286703
zac6e07ff50020afbe1121a68d515207dd4ee9fc57776767940958489d5fffd23e4dac67110ec92
zfb604d7b79d2f1956389d7b82a350136231749e14fea3ccba33ea1d974a38e3fbe2a127049d375
z25351cb6698c516c76020ef11f6d466195a0d2733396bd418b97bd7c9ecea14357d1757c36f84c
zd7787cbd6278bfde9967f2cc3cc7d5e9cec0ba6d960fae944707ebf3c95edc83900b125f67ed9f
zc4d8efe51d7957c4bfc3ed9f21794a65ac646e4d34b485920bf367c0d9b6caf58e6603bd5bbae8
z336a57752699ce3357bc29fb457b652c58bb34d36cb06000f225f21651f275dff3cb5265dffa9c
z741405919d77206112d4eb9a03f065454c513138b6ffbb27219acf6a678ec22a625a7af88b6982
z11086308112cdf98f99dd792b6aa9fd1614281fedec9c868e306c4ec4716da5caba2a3d27ccaab
z5027c0ffeead24e51c245748433185b56f7c52bd5b263526cb5987bdc5bbc3108959e3ff836f4f
z42f8bdaa41d3993ef17ec6962bccde3abdd0d565e6fa03345919d0eb2182f7e6264e25e550c83a
zac98ea018cb47065f3caac8510b5b0d25cf7c3ed61e8a4fd6083df5e5e1003965e075d75a64041
z2812ac2313c6ea5ab97bb3ef030f9f5af0e932708c9b06955a7ee2b4fc96dd642ad7b6327704a6
zb856ba47c1ac3a73f5a4415b2b89361c7e323b14f97f31aabae140445615a403ce45d1c5eadcec
z4bb1346e2900d4c8a37b622a62e9ea243fe301c84f7f36f591f5bc0c308aba1e6b6be6b5dcff02
z74f7f95051eed5fe55a377044aa37a5db9b0bd5394da77dd6387144512a48f9303471f93431e1b
zcafbcecc91cc526a68a8bf159293b12cfb22de0256fb9911db88b6477e6f1114145d9a96d913ab
zeeb08e9112d81efc38f3767f94b7ca17ef943a388cdb90ccb87e9161d674c875509e3f2d32c9ab
z19867a81ad2df743711a609593142ac0d192e1614b4264865aadbd11bd76762b7b3e7c452c0090
zfadecfef5ae01997c053ad8162ca08846a0db619445aad9481e9aabd636c7daa6c49135e00515e
z2c8548e8db2493bcbf88843f23c3ce943f62f426022d726fa05bda0bfa6a52447150f6436c0645
zf596e275ef6ad09c76f1074a80de377a10c92ba26cbe2c0c9958534b23b85fe5fc3357f9586b84
ze33db97e0cdf22fa0093679479c07720bfd303c0c189fb1a7b69da0586de33304309c321232127
za188d2bac7e0f0993dd76e52f2490563dc7b69b59dba283f6267e5ced14da23dbfd6a3f612fad0
z48716fe66e22939645022dbec68198ee6e052b3082d2821b204cf97be229774d6954b4551e8a3d
z4e19b2bda28abbaba8e2d5f550e5d7c591a4aa727298cdea507092e9c701206c8e59c63ac79b89
z45d4c003ff170aa9e29e2cb09704fab61af261c4e8a462e6d7a0018250bb296281921d454e172c
z28b01c0683411a1d42dd76bab2c6fa520e2f1c751e128563679332857d56ceba182a50003ad269
zc042d7c98e2fa3ce7d538024df8a67701836bc033ef756eacb09802a2e1379e596150f5ed4a078
zc90286a1e3e40bdb99afece7b89e2437a040cf6babceac542297b3afcf6defacc078f7184e61e5
z64acc55ca3c3cc4ae966c99916c9cfb41b4a017a18122c52cde738a06304c933ce2bd23299e24d
zb31b1561295c4932371597448824dff64143015c83245516f67e6e90ab346e07a581ac8264d1c2
z3d1871168340ab1b15d012d065f7b94539903e7fc1805f5bcc3c76c512971d56533cbb10fc0526
zd0d336b67b84073aa247dac032f08dd6dce70321894a8b9cb8682dea97c9b3c93183afa6d9d5bc
z9e3cb552a83cec512f0c2f400fdc852df49880fe77830b5105ae721354784f201d51244bdade5b
z369b39710fa8b93da75bb8aea1473786fa3bf2f5ee625d6dfbaa5f847a377036efdc0fbcb601f3
z43149ef909cec14ea5e15f1102ba85f90bedf50b1f5ce9d6af9ef2cb59180fd8fd62fe1812e460
zfe1876b9874e08ff324c23843fb5643f2f010a2c2f995cf62e27f29eb98f91613891fcd570f79d
z57a2d69fcbac1a7db5878d8000b088f1878fe2aa75ba3761f0164b24eaadf144f0b099fd9eafae
z0da9224e884f21187e7efb3811d4aa1fbb43101b3a0059ec0c61069211307a53b948a9689f4c1f
z8b2a0cba5f27fb06df9cdbd110fa3dcd42cd58960ef40f837c1510d883dc7ebf6197174c7667bf
zed39b6be1523b36091beaf52150a0439fa4341915ea160486809d596ca70cca5603796d84b9957
z71bd42e6a24c2ddd0ba381646f001c371f2a248816f430c4dfe24be1b37c806c315c3d59690b67
z05859819e587f3941f7fed46cdd61f254ba2158561547251c67356afd87512c616ba154622db6c
z6944e0d10212a63619e24b32aebdda7c1eb9372b3342b116f7a6efdaf80f1e48186d6ac3a1ecdc
z0e3a71d27a0460efc2d7171d98879fdec42f7d1257dd0c1e97d276a2f50553351a247a32972ad6
z43b9a0902b4bf557904ad4d87743602e28cf3ae26da9b8e24492071553173f43ca2183fae8f194
z1ee76caf4214bc7e52166a6fa2582625f71ecb967d22078483fe5252f1783db1c38c4ab93d94e9
z8003e3e23528ced0a5bdde51c2bba2c667fa69c70a1bb458ab35b886df0714afc634e2c9f48056
z93de9af0c3b959d93e82d0d8606d8856fa1016876cdfb25e669a4755ca898a10aacc370d52699e
z065da78b6023f6c6392456866a849ca7f8238bde9f00396f987bdca722cc4b0c8c82bbe402da3d
zef85930189230d321908f3d941fc1c9b0a25872ce4980ed98810ebd9c28a00abde6ccd4fcc14f7
zbd0a6f791c70ce5365f21107868b1f8f7ae7d89dcbbe22c8bef7bc9be4de0a727577fead7a3fed
z6f44f575daed8660774052c11998ba3d056c08788d4264a1eafc560abde78f1f9465bc71ca5fe5
z81fa1efc3ae74db2ad11933a604b294a482e4dd1b6accba9e0fecf3e7d7d24a6bb4ed2c0dd0abb
z5c5f77864cb5685b7dd70bc2688a007f3cba60cf78cfde5b6165674ee9347d58e1976a335a689f
z4424f4073029c37413d86149a0878ce1d8eeb7568a5f19b00491c569225838031bacff53ac92ca
zdb7d920f2f8b876789ea3cab03d3efc1689ace2b3e476809c34ad2fa607188afd398d5dd2f5289
zf706bf7a8062dd09334eb8a09567b79b16bf7dd0614206bd038fecd15ca0f74eeaea6446d02580
z5bf248a12839f4c607b9f3277e5b502f8721ed430fdbc2573f4d8a9b2a3cdc96e88c0c30e50dc0
z73f703d580a5235dbb37cf031e3014a90e22687d5a3c3987b62cb58d297669b19cbcbf3a9ba470
zaf894d66bc4c921ec72d9e7bb0f6989d828d5098c0e9f245581063c6b9bdf495fe10f2f5026326
z916ca543e7449fb15f35bad91973d762407db7bb5e9343e1cd5d7cba3e27d7c26b740b23b77795
zd939f2905876e7c3db15fb1c65bbf1dce85d54f8282016567d94cff6f79ee6a9837e8e6fc038c1
ze83a7a0a140b5308b832c4eb1232f3841a72f6f6b1f414cb13ba7976b9fe3fa7b3cf519a8fd631
zcea281231d1a4e5df3d5daf2b4aaa4ef6ca2d0c60e4c957ad83c2225e4a3dc0cc206e3ef944f48
z823e5314937ebbf7563191a9d297c6a0e28cd1cc829fd15f041851c0672f2c8615d0a5838c653a
z1d08725edc2d5c7f2b978c06dbbfc24fcd7704d7f26b8d45039d8fb80c659d40033ade1ff96670
z46d1ecfe6ed6cbe8f077c5db3323cc7c132bde09bb1a220bbcec5ec1e00bf3b71be8cc15ce164b
z286b87e39828b972307bbd009efe0ab563e613e52a9866f340f2afdd334c09c587ff28f146a262
z0293193ea7d87c1e2faa4c2617a226ab459089cb0d962c267afc53f3b95870aabfb8c288d3566a
z3c7cdc3b4265a9e6afa74e20eb38e8c6c8b2bdd627d06eab247605ae3b7ea6d8c799867c67052e
zdf9236b6142aa41c5b6e5d1176a5d599a6fae9e8dcacfd4013c7fd527c9a498f0e8141df9ddcb2
zc9ab01c2184c8b501700370bc35eb0495b424d17a0423f530f80be61c798d404fea2f97f7b83c3
z8c519e008425f9ce81aca3524a9416d010984c9c29ca369041b99b1eb1332da57b1f1c4ea5a644
z8d68cf6288ad4904d2dce6c9428ab72ff21e02d0d3890594284da0e7dd541620c882f8b8074651
z6f189da9ec34f8f48687ba4c589dfd5e7505596bee9b201f56df52516742afbae448597b4a2d23
z99b514ce9d0a0591f0c7816870deb355ac2877509e74004a1f7c08efebc90b93d5f59e2c346ef4
z0d1bea6502408fe526d2686fe7504aa8150a83159c6a6cf1cb9010227535d3f9535c6a61d7df13
z2ea5cb8208fe5bcc07d72933727f7d3fe95fd4690ec6562b727403735411247dc6dd6e963a7e40
ze59f20976d68e2e82e40ce03123f6419e8c3ef46e039434ee2e64e3911920113a4430f3d29fd32
za4968965c4d3e65594817382f1e9fff875bedbfa312e3cbbcd5b40568b9f82f83efcfec60e810a
zcafd0a56971d1788e29867d4d293f7155ed9037b0965c1d119834f7bbd44b1ba764a3e2162849a
z387d8a52dae4a0a46935d8974e8cc28f233da0c0480d6abbc50c3bc3b36fdd292f83837dffe937
z1705f6977620b66ce043fdc448b5e6e31a60c25f3b8a3d3e286dfd695680ac52554b34faf645f8
z1db3084d1176ba59011f534ec289885f6893f9f189d46091a6e24cefaf2d991f95d6a2f1daf71b
z0c0846bb18695b5524501cc4cbe01eb9651657190cd73f2c6d50016c8386a24a3ea043aa241213
z333cd7853805e8f12f7e4708496882a456ac0345d436d7719f8da0ff27d0656c346439969aebac
z48d880276840177d0260f9d9e1df8fb0417025e285cf3b54b411d2bd1b34e38527fe98a8b72f93
zb74e5d9838cd4a52d5503fc883c8c991e38ee9e02f8c8b9816b5ed716ef4a7c0f1085c7ce90b63
z7cf16d00923fceaf00466be711e30ca73b51f7e0649379bb30e5d0d36bc6b8832add29e36ad947
zcdf6d2898bf3f59361e9f99e4f147be58572cd61b8ed7be3ae43ba097602096941deef3daa69ea
z5b61a01a098eef229f061c80f3a77cdf3a1835d8aba63352f5a44f9b5c49de3ff623defc23a66a
z0a1a19b23993db9fff76971509cbc13d2ac68ea689d96d04388973507720d749fe144d39bd6e79
z012c85f6055eec91a0883017bc3427bd6e81095579b9e07ba795284bb320f60e4a1af99dcd48fa
z4e7b14f3908160c15bf121ebbf80eda41985b951fc2d92735b4febb9d64cf9d8b016b73e6d8920
z0c079808c044e131b2f22ba34248495ea667278759dbeab0d3e2f2848aff59b7c28574a1a8c720
z0b94a204cfdbd9b38399656f5b06c3538df98d9e242959012c2690c836c8bdca169196d47fecfa
z20b9cca22338b5de609701e716dc30b0b1b5aac43689bd71261ab1494b1152c1e2e19157d88a37
z0f858a495a44e1fc3e7408e9f5376892b9ad003c7f7ec9ead2148387a4b5baafd6339aba8ea090
z0101db9c242af5e2f38f7ef82d374de28acb01ff3faf71f54a3af7fcbaf2873917212acba157be
zdc491e044e4d3532a1951a60d789555f88b962c9bcea7b6fdada48f0524fda9eab6380b1f66930
z9db2079074a0ee36f05441fb33e0b26b619d2d6baa744aa6cdd9c76bf93aacf47b8fff375c65ab
z2ce9f5670e616b0aa7a3812e66af5a72e1bbc4c28c894f08c7366ae19c8600c48e74c36615b0c9
z71a6a647f5aa02dae65bd2d8d648d9060c8249654108fd6098bdee785da393a6789728793ba35a
zea01ea7572959f90a2c37d154fdbf603ec40561fb0ae8388fefe5b29c5a0462b09e95447a92aeb
zd22787079757e939ed6bd52476dfc7566ab740fcaa7ecc41962dec336e6cea8cff18e7ccf77a1c
zff6ad8e341b774bce85fc538f9dc4517a5f88f697790e85f65a77e158a71a6e4f2b559ad7a6bc8
z629504f7b3f0e6bd89580b68dec2a1c054c15e071d2f1f759598b30f716148d7f117138757ed8e
ze9ae04b2290895b2ec1dfd9a5b7169d937509bb66305764de24989f5567f507c8a0f790ee74040
z5b81f71ac9497d5605e742fc600f7638cf616afc1dd7434b4e0cf32a12f16a5f84a6f8a2067acb
z818dbcd297c76cd8340b2f763e5ce9577100b8832e54c86f7dc9b6cecbcab04414c53d3bdf33d8
z06174dc45d820adfe45e0a8d4eb5f5947dc03f05856734c6e700b02df947962d26ec3efbfc3cbb
zb8c60827fa4d2ac762c8ef03b54fb7c9803d723837814eb143dc3bad894a12ba6cda53b9add311
zd36ab63eb26fb89bb38ee567a0149df435a342580490b302db37ff2682e1b9c1820537c199f0bf
z3ff763262eb2327eb4a25840472d4700224aac3b844ccd298df119d665815f7d33640ca5d6a086
z4d0fc0027ae61ba06b456453799839549e962f2d414455d217d3c62dd18d59418bef7c0e580b65
z261576df12e7c712908e72f5c45a45edc7232ca571d8a3bc95b5f0299048fabd24c9d0211ca0aa
zacd5d19442a7507fd3889c924a1dd026843fa4ec1b76b86a46792c6294566706617ea3787f53cf
zd4ce6f40668a00573bbd1fa8963e5ad8ccf4daf252c78ce02034b3c13a6035a7d8778bac0c4865
z155455eafe6a86501a8b3becfa2d1763abdcf8263202148f5fdde8e1a5bf364ce96cd9cf0658c8
zfefc1a2d772f5714b10d019e2dfbfe8240fd782952b7542f3f0073bd01f0181118463478eb2907
zfdd5a516419b8b5e9a84ab0ad949042c86509b1a488d3864ab8ebbe05862aa47144eb5c23a2ed7
za676c6451e7c1822d0f9d2718ac708acfafe67a6e5809875b71d987e425d6d4d4a4888aed73e8e
za38d16d5b2bfd0e0e9f63d5031ad559da1c953ce60393cd104c70efd3a0b03fb126678a1740768
zde940340cfd2e2c2d12ce34351eff5d5ff9a467280e6825780b5b0256013bfdc9e0ebed4bed91f
z1dd4455b5e619bb470cddc8acb514fff6603c808dd83cc3c39df58fa148bfda01a316d04456d26
zca1c9c1fda78a0014af14e0e5e31ff0a4f32eb700a168fc574e9494521695846fc9ffa0c1afd12
zeaeaf379c300602681ec930ca00f9d08edd512806faa0902187ff36df0f0cfd4ef06ebed0ef8b9
z2b429fe44acf37f05c5bad1de2ed62be71dcfd09b75b32fde635a16a5dcff5bd59900aeeda22b6
z9557a47086ea6eedea9a8fd3afc700691e4463564d9889eb0ca93eb32a0386d74c8b77d2935419
zf772c562963fe061c7b8ec0364bfc1774cbb9281ac167ed25e1738f07a93922dabeb79e107cbfc
zbed876362f99b26c297c85b13221c85884b0458a95dcb66765a141326894ab24e9205483c9ed87
zcd1988560fe8af942764f8992fd323dd708236da29b39e6d97cd892a9ad5183b673f94ac2a87d9
z9a9f66557b252c607bd846a45a825196a4e9353ee304589b31510c231d8a8fddf2c43d64ab4549
zc55868f23858df27c12572cc63fa81875533ab43909f71defd65c4dce83a8eeb4b05bebf47aad8
z24760f847a588fbf51b435187a99564a64c2622311a37f6aa2103c1343f604e2d13b4d0b81868e
zeb881e3efd309ef4e8c3cb7f8f0c6f944d24ef11eca4c3a754a59a9889a2701fbae2048ca673b8
zdd55e7640fb975bbd2e6896f6494d465b015154a6415b5f8e4ace7f07abbfaa85176f8727ac764
z00cf9b30999d676c436fef8f61c1db38fd8071fa323a350c6da9ee31f0a4d9f5e15fd2f9542eda
z5ca009e5ba16668b6a1e090137dc2b675850a7e7ef980864364ab8b541c0718098597422358449
z3b91f384cfa05f4c441c82d922a317b80440376e44100deca7375217a29f1c76f496a708efdc51
z94a808cf32f71e63048b1120b8b50aa358a3a5f02a1beb3efa64588b02faf6bb23ed04b8cf3927
z9bc59f109eb849dfdc18eebef3de9fbf93b409caafe7e5eafb791400ea8662ae2a107301d68463
z719bf033a6f68cc9c6d7e8b2ada194e9e63d43b6791ce7360d04d094730ac69750ece56478b081
z82462936d781e3a809a73d47bc5a0e018f9562042ac2598a2fef2fa32b1e88a385cc30251351c1
ze0cb1ed18adc87b70cce5bd459824371324222b0aad72aa8d6c0ec8ab56eb8cc7c34715b2a8958
z81b0d8529d10aefedde3e4c1b6fa57abf32a3dd8c97824d559523f142250ecbe3dbae0237c75e9
z762d09dfd985e2d93cecc57604788e03b684ee2dc3afe7b4ee04e0a95f5214fc1e86ddf7d95e6f
zc9a08ddaf0d45e3fa59a8ba4adc18ab8ebaab2b45075636c15215ad89f4b769f89cebf501e1290
z8d0f9973b467adcbf653571d0ac55088782a0cf1c609c43cd350fa5882c5b395f3857b7d574103
zabcf8b867a91ae47d26dc5fb5501006b15f889151ed276eea5fc333843ff065d2231ba8a670f7f
za50057c87169e6fbc9692dee66ee360ae74ea3365ded28d260e1d5b955221bcf0a698996f31fcf
z981047ac1df471fb92f1d3c76efb277154e216a70f0102d1958514afbf1f3661443f060bbf6afc
zdbc0d98cfd4a9bb7b2eab41aef31b29674b3f8f08118d0ea0a315dbab5631012afb7991eea3550
z1628702d5ca97ff216e3aa4e18fb44b593ff5e7ae13b1987701cd8aaa0f37ed0272222b81cbe27
zbbb1fb81c63f11f913e00c4d3137634c171f074de322e3ac8bcc00d340753e0ee88d105fa97c68
z5835ba87c9d781c2706a32ece0a6bce57c0952c8f171d529b71b21623cd7a2d759f76f1cc4f3d0
z6f5314640ff18a49e3cfef41b1c6e38b41a638beb767af0d7838868fc093afa9be291178dcb6b6
z577758d37cd69122dbf217ac46b9d6f135f8968afccad07c5fdfc0db8cee3c28a0c468a0f0601b
zca655c22efcca8a0e5bfc5e7933ce3eec48913885ad6dafdb47b55499de16412f3278600b2055b
z5a10ef88c3f4dd0886f7ec86a6af61d3b7cdcbfac863fda4198d94e746fe2ba49c889b43aef8f5
z4cceba28cb461904fa715f2d938a5327cb504be647780739f067ef76dc5cbfba9819bb0fe82bf6
z4c01e5b8d05d70ac8a78ba0e50c6e8d28bc3d8d4a9fcda04565eae704133583eab6dc5e7e90590
z80d595cafc0f916fc310f252a1200c50e24a87b1bd19cf42aef381719d2f6c24cf7908a0a19f81
z1d562e61bd9da781c403d96c982e91e33da2c1e6e435318965c6ee9a10fe0323edeaff9b53185f
zf5fa6609453e36e6429c86b2521757206a9fc0c8b6ddce1c059417f4e277c243d57dbb332e0f67
z4232590f679c014d3839efb775026424a4a3b3d9c5c954bb7d51a31d4f99640e2042f64580e437
z2520bd5810264c812f327159070b6e64893ccc8b5b4133f00b6256cbffddabd4384b64e305e022
z02e1bcb7e490449bf21817c983c5d5d425577f31a0ed0b6cbb668eee242e389acbee78dcea5129
za2e92af2914322397a8f18e9bb7826cb3a1a185428ed1aa2eed91958ceb158f4455c94f222ff68
z291cf59318a4b3a97d28b795927cb1c801ad2fc1d724f5b1f90cc7e2da0ffaa9448d3442c27e76
z7aafe748bbaf5f4f434f4eaf47175e72b1a867af0bd281c0ad90bb2737e64e546d1ecdd8fe66fc
zb5b35670e49d59d283a01e7867a16682369b4160bf0961372fb31f47c7754e1087590f242c2270
zb170c92a5bb1987c4a90cb45e003be963aed5d7b1314a3c12b1e48575b96b18a933719d63ee202
z4d1a6f0ea37d67b33f838737e815a480c398dbdd4f21dbdae004c594e8eccab4a62678ab65bbd5
z0759a8e6b9d0627b7345ba58e01a13984de8c2b7e1e2920b9547b7ff6b9f94b5b1847849e03747
z1978a0e849b02a5b2df2bd4e34b3531a04ed6dcbaa5f59b73462d6aa450ca66b454404c77e036b
z0336e1882ba1579633d2df4ac265e501cbacf9c47c9c93360582ee0668f73a0ce32d5832bfd096
z1a86621c3902d8d3d7e53e2851226977ec3e5c75638490b1fc8065af8ac698168a6c53fdedf4ec
z4d90bc45328f6069c0caf3b5fcef0dfc29bd8abe58e1d7123933767837a57f6450141b4939ef64
zdfd3386608eed9d07f103ad029dda792641cc186f4c032ae137354e8d769741e8d0cb9fc8f52a3
z100b1c7b6258802f679613c1761968f5ebcf56cdefffeb92203a54c060867d35437c8885d01646
zcdf045e7e4f3286661ab9de3eed28fdc869fa74ae0fd6fec076d95694f6feaa34f4d83c9dc32b1
zac0067e6612a5f075a224cba2eabb7e1c3eed4a8210c59a801a804fbcb3ed3bcba384005de174d
z3de3e26da5cc63a8d25656ed47e2841a95f8083579cc27978ff40d206f6dbe6fc1935ebf41ee58
za59092eb901360a53db0dd15ac896b1ffd340a81c9a5cc3884a693b3ac93d96e69b4eba450e451
zdf63ab54b68fed60b747869208cc9ff72de0915fe908aee5ae634a8cad77063442ad0bee00e3ec
z1dbc2508a98b94408678a97484fd7dcf9ef1d302adc49407ee74799b7f7471cdb2c8d7d40d676d
z1ba7d31ea2c659377a3a7d1f0eded07220fdec866710017e363477daa472b0a4afb617b7a51bd7
z685c55c0824a844c70b764bfcb40689f89228f03a02be431e914153e81af926801b2e56b90db6b
z6f8707f5d8adde0d06ff844cbba585b750957417a09b764b62425be9eaffc8e44d18daf49aeaa1
zcaa069a2ca1437dd12dc62332a010b4dbdf71e27d550fb40f6662d6b7bb588c1d3a027da212dff
z8f1aa232c6283ac8199d2044e924111d755f09b263045b0e450c3029ac6d3cc92498eae47cf50d
zc442044ebcc58b9cbd711c9e3fd6233311e1620ff3d39aa8b9c047abe0251a6c7bac44195fc7b9
z0af5d068ce36b88ea218cbdc23c47e836c72e676a242387170b04346193800393ece859238c052
zb613105088431168ef0b7bcb3959a6656f35b4cdd375227990f8bc67563267413d0b9fab39f4c3
z357bed8af1e9489eab4c6dba037f61f0c924e483db3ee2133f8c5ebbde8d5a854deb5b950061da
zf201eb22fd55f8cfc2737276faaaceda4dc5662107e554fbdc9c879fe538acc336e0a188cab7e3
zf6f77f6047b065722fd586f4933034f5ca3ca2a4e4f7a7e9f7e38b214dcc5650a86ad61683070e
z6ae2454041f04e90dce0e5b61872f04c02b2baddca0668b14002f6dc1d738812f905157d1bc89d
z5928c55d63815ef81263bb0bca09fda6bf05475fc20d2af0dcfa44ceebeae38583f869dfd6b7b0
z8eb52158793d84113480750246b627adf96dc940790c844a68b6a457814b590f5f33d6e8fd349c
zffb31a66bef4cfffa861b90078f4ed5ca5481682766d99bbee133197138f6f2ef3cf23085609e2
z0d44e738e4db4753897ffa1ff91329ecb77e97ffd545e75f9e3491dd3959bcfa052bc9a6daabb0
zf750bdc2e8177f45641d1f927c81520d61f12f3eb94103ce133999d308b2f303e82f48375081ef
z3c3f3646f3a054b5b36af39fa5e1d3d95860b49dad6b8fe86d568913ac47871891cd2494dbdd36
za42b9c91deff85a8866fc84d0dad5eae22266b4f94ca6a09d176a80e96386461cfcc9959c62c11
z129eb5a28f3223e53df5d913ae8911cfd9dde080547265d0f8b0173017490e2431a14c8978f55b
zed37d6ac46592ef04266b83ffad0525f0d3ecaec4576db6d58c14b98e858f784cb713e44f289ea
z4e0d18fbf01fc197c0d9b8a9a3b168727c932c1a2042e08ab07cf97f13ddcd65ec5e20d26c7085
z217c5db1b930887c7d17d6168cf5d36a007b4b1cb4c050aa58310dc26862818d5dadd93c23d240
za9b093a1c1299b0f5efc5ed8f40a969cefc4c5552913f8ad84f5db094a0850e0b5b59572c76cca
z10f7567c6820fb2fb6e7dcf9f490ad9bcb497c205b887d8a2a87a4e50eca4beb218f022a02cc39
z5fffe1f505ed394b365a1f17f9293a299496f5eea632dedfdb79b2cd592681f70c4f6e05d076ce
zc6caf8a7a50635c79a60d16dfa1e68a56a6160378aeb0a86c1b72986e8ca9efdd32a404859a48c
z1920f5399eabcc389b1a78d48293fa83c462f70f8467fb01dfe33a1f113d202a88b645922cfc56
z0de0cc3f50aa161e5647ec63ae49ade7c07338417ffc9973b54bedf57dbf2de54ac2611f62473c
z62c403d8169c24572ed98053fbc336ee606cd895d4762ec69c3e22a0aae7c4ee0de54433cf6f27
z9cca6ec62ec574b9938807f11e95ffaf759b34a622407aecfb7574cc96a32a45fee02508bbd728
z18cef8eecfb57c50fee61b8fe886902022866902c4dee12823b67c8887e5ed96ba2e19766587e9
z6b4e0ef71e0106ad6ad467234217a4e263403e95a41464262f68fabccdff358da87ccac0ac55db
zcdb0b689d6402315125620e39e35604cf90e985b4d000dcb4e44f5e7c8be2d59a8551c42105f24
zf40baf5b44fa7e80d541fef6870726363be064eae2eca06a50808e1e46cf00be8b29e917fa151d
z3ba2d579710a8a657a14acf98543ca823e4e801a82ebcab5f94a527ad564d7387b69d76ca1028b
z7f6648a7f795f6df5812055217f15aff90fb3b84428d5b3ed01dfa52f11639fbd61720086d8d15
z41f318e5c1c9c0edc23cadf5a4db59b09360631112a591d1c0c4169d7d76ac15f4d6d00a74d037
z4d798abf5a2fd5124c76b49cd31f4aef7c32c83b71e47bcc77afeefb949dbded7f3d3ac61e5dd9
z7e7458e83d83111047b9baf735c960b5f9ee3a36ff612649ab89fefae21cece9e1c8e82924c939
z9a8a10789c7f7b73a046e04d3fb3c50b748d5bcb6946bfe7433e42c540a6d00a3e38fad26b8463
z6998ac2e57caac4bcafd083b40e8f01785a633aed6d75997040a50f71f609df5d1959d723f97e8
z5ba621e3f7cdb0f614ab546072b1942d721bcfb2b900952912231fb68d2f391f491163d03e97ee
zd6bb8566075d825f823d5d17dc5e635fa7a61c014ac5c3161292fcc4c30d7a6a7803979680eb23
ze7258776572d90abec19adc14caeeb04151427b8758cd467abef972c28698d4860e2c04e71d5ff
z1ff69840bd0a20835b1b6268026a71d8b012d667c05738895e573fb5c45e711a7ca22312b5919a
zeaf6f0820dfb8c3aaa1a01919a72ed5dc9e457726fb315260a5f799488911ee9b38deab716ef8f
z91e50f16904846addc9948104989bffda116d2de8188ef940f8e38acd2203e1a2b0f40b0711124
za2776d80c3109c9968276d808ba552ba1a42ac66744a44bcbf3dbb1b4e1944311b7cb6c17230a0
z26fc2151e8877568d99af569760fac200c5cdf396edd8c0fcd5ce0b96085baf4ef673b1b70e9ca
zdabc2bb3abf301fdd178f7b8b27f5f9c4f4f8e9cbc60ca60f3ace77fb4d4272d4e4834792a1263
zed5e95f9e181c0f8b0178a9f47a21d79ed4bc678a031ff3c84208bb04ff339e8212953e0d78f96
z8ec40b613b847665a6ef41ba0c13f9c7b49c1dcabb004343f77926b8aa81e7fa2251d0a64ccac5
z3f79c8132e3adff6fd20dccc84aee5e13c48aba4aada5daed932f6e2882c91cbb768061fab3bfe
z20ede2aef9c99945a43b0263df26525eb19132150d4f0b4dcdf7ae234d55173f331daa30baf9f0
za483705bb6f9467893da7884049189c5a9226f3456bf8b57510eee1ebfebecc8dad6127ce37d07
z1ef912643d1c4a3113c4025bb930ca62e5c787591f7248f0069dac341686a923147e6d8576de78
z0d46dfc0d1b9ef723a23c4774351f0ce52bc4153401d451b509899645fad941bc39f7c97bd3469
zbc3658da06bd27ea8b1b7f72f5b8bfdc8255dd6c907db78eacc9b0662e41f19dd6cdd564a2e5d4
zbf0e26db1bcfc3e5fa648af80c1a7292d9e847570951638da51d61daecde416b86ff0130b50e44
z31aad2603d2e3460667f5f41a402dd2c2dd22d63906ef1c66962687bbf3ce148dd097f612e60b2
z57b2ba25a07f4a8e186e88d2a8b3ee2e4b545417dd3495ff8a22eefca1b401a164eb3a27f8d0ed
z7e6f7e6d13fdfacd3264037971db258f7cdeabf082ddad5c316ffbe383cb7799df9a938af05769
zbe8126e46d84a13f4e1d16cc36077dd0c03a0f575e2a638438fc5a81e3fcac51ca4b134a656f1c
z3cc160052ec576e66552848006df0f913149db9696d1b85e7aee0a4dc7345b79107d2670c02b97
z7210b9810509dc626dd633bec1df29639c3ad304a71df0eec8ea49c6b6ea86ba6ff2f9d43d003e
z56901be4662044d6133003d60e4d56bb2dc215735150d010d396b45de3e602d6c315f5d8056295
z5e643c3712ed457ab6af2248788e0c678ce54cbd8b715ed1a0b9a7c01f1ec8db22179fe22ef7ea
zfed1c3576917946fc26e5444a2d14959813f66dbd5319d9157df551d4e6fa189c7130a2ebcc2c3
z5149e83a48046aea32829869ae5598eb862aba2aac4dfb068fb7e36d5f391e5a1646aa8fc99f6b
z0bf36cf7a262b844134108fb487594d061068286c28acfdd18e57eaaeeb530bca19f3ebef47a32
z317d6fc96ec416d4c4847350c99bab34ccc9ce52d99d8036925efe68b1ad723baa7991939235cd
z0b539816a8930c47d67c72f1de7b8a2248a9a550cb06eec2b18392c615a301c06c8e3964205e36
z9c3122d291a80bdd41545190610f83b03bb7b67f260593936c41a4c48eabaa3eec3da1061b04ae
ze242c314e298c9731e0654e5f028cfa8e9450da6fd0631cb8e42f97f747194a60cf1a9d8722377
z182f23fcc48237077438ea04b19bd6482cccfa1fa8f9c00cb173a5991ad704448e20f9f5d13592
z081ba22b2dff2cc6e36d85c39b3fcac2bdfc6a197d633cafb51d6c46107cf08442dd0191e7ca05
z866357c69d28a25c13a8b27290db90d4b812800b0d0b5c05caf83dffe3ad342e52fa325e6c3da9
z09266e28b2bf0229108d29cc03985b23eaa948e11f05f4731db6a1778bbdf224b19203f6663234
z9a498b71eabdd4d48136afcd8cae8f2be13f1c4bb9127a764f18bd5711f4f9b0abd9d443468b49
zeb620fd910734f3c49517f61af99c6d1e933bdb77ff19332e89ca12ce195807d99f5670b7fe356
z6ace2ea7be3d65e5aacf2963d4fecf885a74d0e72ba794b0d35efa3409af5da1934c047d015ed5
z437b3cbca4777ca1495540f28d4eb54c3f8bce73c00beceaaa80515845011c1240295def2c913f
zdbf50dc22b7dcdbaf1514cc0f85977a70a834ea2f5b8ed88fcf48b5a9c991573efaeb4a6c27dc3
zaf75b604d7ea6c35d35835379c2c1457c2fbd8f5373f621f027facc14eea5349a1137d6d36628d
z58afdfd68dae7194142ec763f66900d6fea7cc7439f2db4ee09d22fc95f63d50247eed961722db
z132130eadb459cec2adcb56a44ae467ea39412e64bddb0f98d103d4962d44f9b7830779d0bb730
zb47aa29cea368be7d5376e6a29c5671e3261e4c071e5c1be7960dc4ae829c3e0c6c7fac7333e46
z989f4eed7dfc26ae523e2fcd1694e20a5fe74b1bcbc983a6d024d39db8a15046c41c55aa346d41
z8c614ed9f80ee29e0119b552aace1f3c6cdb4308dd2324c01765faf6309bafcd638fbb2bd08397
zbc97bbe9aa2c9b569ef27dc85a54cf26f141387bb5beb387a8170ba89d2ba10f4491e3014c30fb
ze93bef1bead6ebe83a491a6031e165688dc1cad5517afe60ce2bb9e5b3f6faf28dc11d6d91ab27
z9209037a3f7d2fb3f91e32c68eb8f3df831447e679dec256a459b269413035c852ca1d8e7b57c3
z63a904f7e7a86dc85b506d6cbbeaf929697a399ef48431dec18786795c74c6ff5bf98174bfe98c
zda3750363632713494e0a5ce0dcee447b2b0049380a6dfd393384564a9ddc623f1c4d154b3f15a
z4727df29bdae7341cd49bea5b30d4b20d78346b4c81a1b4b29fdbe7b48563e883a92c12e773755
zd000edc21fca9ef667bd92f2e15e66e22258b911e708c7be11d941b3f698f8950eb57af3770d9c
zc4480cf26c7ddc3df3600249ea360b38c85c1856a3656255ccd986a260259ef1954e3958b0f173
z3a67dd4cc4bfe0b346b5c3d4310e9b4f759804157eca552abeb6ff613ea015fb9bf78d82f9b666
z4dd97cbd46e87e7cee956358e10504fc6a9ae10565163bd1f83975ec7749593dbe99f53840338d
z531db0109b1e8f2f3dc69d8f4950c1ee163ba3c56b400c2fd586b8716e38b948ce100f2dce6af6
zd8e9dd068c5899aec55fb67a1fec7d1e18eeece22e5c3069f55555940d27243a6dcfb1c536b8cf
zda99d3fe20efaf4b37746348ca3d661c27f00dfbf8b1b3c9aca79448908f312d6b11893089d735
z80f0e5b26cf2c730644373379039d5bf7f77ea8a30043bf24c9f4631a066b4194541d54e6d4462
za44b14ed84c6c9bd5698fdac8feec2b766bfae8c396162a34655b75f0d05804c408ac68e54d9f8
zcc1a2bfe3881a64c3bf4871ee8a8985e1c80339a571c95de08ecb7ea61ef75fa78b07d2c5ef0f0
z94d8b2c3083ff02b26ba50419d34f62808d46dfff08a54151c2cff27487f56306643fde2a19182
zcb41638aad128e677cca91bd98e80b9b6960d86790a5fe429cb70168bf746fa1340b2f018b57cf
z3921979679aae87f7aa44ec5b579ab7ba56785ad228cad103438adeba567dcc466e146a58295ff
ze78019f565f33e0803fae072537271bcaeb81e9f84816398ae1eb08577c31e6b98f5af1c06492d
zf6f1b736de979eda99d29b4bf284e0e64e8f2b4ed6a47f65f8e0b9546520461189eb8d9e29817d
zfc7b74c097453e7ecf66640ee9f3445658f3edb8413715a7e09f24ce964e995408df8579fd0a15
z66676649ba3cf10b08817a0803ef032a922616264cb7b0ca6d4eaacc216873b581f204dfec93a6
z21041ce911212e0612f4aab004d8f1bb815fb2330e2c646b5910c0ce33ae1d63636d132bdfa557
z1a6f33026bba8af61afda954235e9b17f5a39d069a86155301acb54477340fcdf116e6bc13ff97
z6c07f944258f6b08b85705f5d7a88983e05500f2b6bf0712f54bfc0f14b0bc00e6a0a9349cdf58
z9297ae2826980b5ca61fc9ded2c64893efbbdbd56b28610588f6c86e9b2839e658578553732532
z61131e43b7b77c2459240dcc6770023c8e24b918d3c1566a274272d81a8f5174b2a80e7ed5c024
ze2da32ec463ef5567f06cedea28e2b0013ff2bd5c803eead1d84af8d1400d45b0e578ef8dccfe8
zaa961aa2bdb134d142621f5ed9bffc3a90106d06d5efef08b1caf636fb717942f0e8b0113c32e6
zdfd9c36c67154c118eec8af5491e3d02973d3035eb821e3a535e2945f00c593b9458c796d1deef
zf65b0ea10293c949456388ea287bb85b824ad819a1c45cf3da671e26de2d5eca60bd6df3f68597
ze2d3a9523f73f8058dc87d06823ace8cd5e871ca4034bd9b443dedc5715dec5b44cf615cf80883
z8b74198dcfad278c7ce97dc4660c5d9b2850ffde0f421503122b3409389252833f2be560477125
z7d46e27139717af2b60dd1e9b2538f8777b48d5a1c2c51232c4eae71b70ed4e9204e0e0bb77f5d
zbc03cd2c2f1321518df0a2233816bb59cef8dcef221c7dd16ffead82a9d48f801144d6be581a0a
z68455fa1a0edbe89adbb5327ea35280d041d10579174036aeffa8f7275a18f73201fa826617821
z9b7d125597a8eaa4a3c67f71f5bccdf6f4e4354bf995b581e5aed8fc8f1d21e86ee6e9f7fb24e8
z283cc8c6eed0330c983ace019275dfce748754bb1f4a324962dbe0f06cf5b720e262c49aa784a8
z95666e88fb0bf507a64504596a564d9c3e5dff033538a30781b7ecfdffd0c20df24abf8075678a
z1e325eeee29756d197d2b2df47b0a1b0a1d57fd1ba238f2be8a1d090959b534d5ab6e80a29498a
z130147d6bdd85cfb2a2473012c603517bd796bca958d8e8e38dab1b0cb73f754ec327a8cc69a16
z81d1454d7ac66d5696a16f9dd09b832ddb1620d427fc71342254fe17071a98a0203c78ce9ef95c
zfb61f4800894c77365fa6067ce08cd0dd59b19c707a54cdd62ca0cafca22ff2e58f8132237399e
z98da7793f0b542742d2601487d96826b7000ad9b6ffdb5a0f721cc0f3c3b2dbdaae0785ea0c702
z765447dc1cc15052293c9207d2ec4c38eb2a769ba45e1bb897a931d410e0771e8cdb20cd2f939d
zed9361f20f203806d7db5b4405d12a3b793c675dd489f3031881dd01b97ed77e55f843ebafd032
zbedc85f3d9625834333cea75db25f2d4711092c6980a5e0366bb0e7ce62c00c2ac398470a662f9
za83fe8d0d4a95438e41cd2d79cde17358248f2b707bb190db9ccdbd353c825537928fdc586e03f
z7a04aac9f7a6b82c92772bf586f6cd5a04b21c50a5797b54e252bf9fe3562c244a724ab55365f2
z69fc1ef9e943233885318bd0e77128f19d1fcccf3978e55d2df9ef7486cace6d332054e2240be8
z973495ee7fdb2302fd1e3090b393dfb5d6630d29f86905941d0dbd069ec728cc6ee979b2d0961f
z5e23ab6ef4ed2d7c8d4e6ec847f9dad4e0a6a91112cde9c7dea3bdaaa22b92ced308944c40418e
zc61334f0c3599f6f1fcf2c7e5241966eb6b65901225c0f104cbfcd80e2a581810db849a9f92c2f
z4f562021bb552cd218ab061d313d6268714d422fe77fa5239d8ee200e49879d19ce5e47859e7cb
zbd5c109ab3d462b997176e30ebf29b413a3c2cdd1a3686342cf7336e97a5ac6e0caa0996d0457c
z37fd6edbe9d3d16b6476c2e113e5b22d71b064667e4c373886ac5620d5672123cb5b47d1a6fee0
zccf28fedfde6a057cbcade8cf26907d6b975dfacc2d3f96143e5bc59c1b435501b86941a33fa64
z71a53058287dbe3f762520604b3c93b4191ad1292f9abcf3781e16b1ccd7005039b115d5eeb72c
z6f7669844cef5245db7bd3ae62bb9ebe16095dcf73500b77d10bff87f6a8633e60dd616f7b11b9
zb9f4c4f967a9e142b5d3783e4057e738a7ed24d3a924e06a71758dbb73a647f01b439e8e251546
z347c1cca22981ed659ae52e59c184961bce9068ff80e22586bf8b991543dc4c9c27b8a1cb9b7b1
zd5e9de88a7b5630c4df1e316c188af350e77321d6fae82d224c53ba018eadcbf203c9dbe3f6a4c
z13d786156f1c799b4c302424685ae07b146248efbc29478180ee73bed627a6282be8922f88261a
z67b45e8325bfea98852565dc5c7e164ac168ed709999fbb68e4f6b57e834634f7516481f7f7295
z839088d25814b09b23bd78de7d164b31244ba8511b9bfc793e02ffa79bf6f16168975033d5f426
zb2735fd6de3e32173f5dadb3d4288b653cfa0d9ce69e888ed6ac4bb1ff5c9ac389e114856ed864
zdd0fd5e5ff9e2155d54e85861d744a5e875bb673b8d1a3a2768c5ed1be16c8cfebb9d3212f332a
z4f446fbbe115d71a767860fb07ecd04ba68136dacd175e0da81f2c8e3329894605936fa01555cf
zd1228e3ce5fdf876f0144bfb03d1c08600baa1c455ffc9ee2f88a16a7c0bfcb1bfcbaea8b0daf4
z252e18e8c6670faffc7c08165ad0c6e687028de065381b6204202a4e8f18402eb6c4cfcc529adf
z562979faa9efc8d29cbc1101b24db1c230059fd6a9a438af4918cbe36dfec0c1e33534ce873d97
z58884787e22f89fce4dcd03c233538afb78f73bf66c915699965c7db7820993ba6911e096d3683
z828b4c3523bf96215905ec79897c64622b97168ddb1deec18347d715280be63f3b5234d637700f
zb3d46e5dad6305f7c9e8b20c55277a4dabd06253ae0b87bbc2c0687f8bf37b9e1913406aebbf23
z0ac02593d765efff1fde585c8452af01ed26a473dda35f62ffa57995f98b0cd69910ff5c43489d
za1e3a6ebe55ea75f9a70dff6ee16398c2e6fd55d18f14b810050270e0e14389ca68c3c2c2e65b3
z6b04ff6e06d2bb3dbf18ee50c888e0cb2e9d216600884a3f13f3ec398d624c372b17a94829a862
z0e6fd395ae81b128f8cdd4867b867205576a07a1b422675b95617ae4f561182055ec2fc2ef32d2
z1b35f00ce326c42f77c6fe42f212c92aee2a7514dae6fa36ba23ed55848d0eae8a935bc6a911cf
z0b0ca97c30d58903fcca55360a573150e28bf7ea29a68aae39f519c49638b095adb88a4fec5ae8
z2349cb4f8f3260ae974eb39681dc69377bb5ed15e89e5c385e290d4737135e96cbd85dda344b99
za5b9e4aeee6fefbad6680252424e436df8a994ff28eab278acfedc3eff7061437491ec084fe3cb
z2036a3aa71811f486764a2e60d2a8d48dd83e870429e3be852391b5b7b698dc42139434b6607b3
z08f69cb030aad51af55a6813cd1d2568b1016b2c858909cfaa559c20d97c0e0a53d4c89fc92f7e
zaae5df9c9615a60f3140dbbc1173a5ffbc4fbeb977140e393fbc074a25f255875921be7b972df0
z0a1e8272d4dd78f7574d9b4e667fb028fc11ea6239b4361a14bd54b78ae7158091c67c6cacf4d5
z8b9f0323a270cf7393c0dfb9f6fb6fbca90a9cb7a40880e3f27687c28202b7f12e25f6e0bf3da5
z5d55cfc306f8006160e167e23a903519ce873d54e9be1f9be9c4f361ab7be850c796c903612211
z62d4d511bd52579b5a00e5acb12c5fdd4fea0562a2f6938d764d1265a0ce466a29116285e3f551
z192e96c862587529b35af087a9b7a695c81125f6bebaa8e0c888920b74354c508316df2c56cc37
z2ffdfc517d5730428b1b0b8bb267c3348815c48b8d6cf89d2765b0a7ccdf5088517c5dc38794d9
z0b84003b7557ceb295a714f695c182278906566c9ee4c4d8fe647c992fcfcf67d7c95fa807f68b
z3b6223bad1fd3c0676572bf4ade39e83669a1a8b163448f436a4a4f22ada5dfbda412b76189849
zdbde17bedd1a5003bddb681ef687a6f45d397e1f1e0f1fd91768e1c02988b8f394ba4cdc1e2d23
z83b53e378bd2d0c9a0e3277d29bebd16f4e450c890704636d074cb122ed142fb52af24f05d2ffd
z06153814d8b39c34075694bd8ac4b682da53f13dc8cd1b18d9eb9be542ed9ef46e16f1a9986a08
zd9dc15fa718a00c1721a932ba86c4d8b7732bd8d40ff09f474e6fe7be56a5c200a53ea5eb25200
zee51012170d79b9cf7121fdfeb0db09b3993995655997554da79710a1b7e6f4cc05db60f23c5f2
z7f0f61fffc581af854c9a4393ca1587bb91890d8893b0ecfc86f1bb52c16d8c676afdb6335224b
z9f287828ffec193afb29c70b8b573b108451ff49a67b8950dfa05db3eac80ab065018638c4d438
z2704cf3415ebfedbae9481975956a27f3a2925eb85d2f11852e23733693883fe0814994be40775
zccd8ede4c308358a198809e5ec962a2d608b28048376174c8cbfffd5231258ebad81635015b7cb
z38590f4050b9aa46a027b1b4ec2ac4f323cc03181ae83a9bc14d0a78a138eace6be2be87c8bcd1
zbf569b4bf4f743719f8666f11eec51811f3abb88b7c10114b21f9f855f7e2f0a263ace9819a94b
z2c559a1770c21b4b104d2d0441a5895d0b66e2a0dcc6cfecf42d48ead384eb280e74d89487b597
z042a50709f8317a2120b9ef5cee7ddd270c5bbe8c7fba5d4b4af1de63dfdfddc0e802527d58542
z635a360cdc6b48113cb47383398ac2a712384bd2c2ae7e2df4247e674c82c6afb16615bb32d72f
zdc905ba37f334be9c742d9f515d6c015e36f889983b2ab3642ff16e509a6999c261c53db621f74
zc22dfd6afcda143825f94e69284efc36a57b5a2aa1ef526f1b0faf596ca793a3ee05bb30fc8476
zd61e13bc6df6ed63d208d133a6446789afc25b59e6f2df82427190d0b14552185e831c69fd4858
z6ce25ada2933067f3fbb6d6026f1b9e662fb304b96138e482f057e22fb08104aa891b19e34c1c4
zd3fb53fbfa690994933a9c6c4ede85c5eb8306bf9575e46f46cc6ae79d44eb44ebf64c2096c2e0
z050e018e882ed2d7b8505a3b8069e9a3e08037e55879ed3f1f6ff305998ded4d6eed86c3f036da
z845af117322d4ba14970e5abb70c4bb02db34adaae7f75161949a0a28bbf02f5b619c17ac02e53
z3172a5e69113265da304fb395fdaa84ee809e0acf16bfaef4f9e5155681e3a8ac35c5673e588d7
zeaf03adb48a118e4ca02bd52e1d6065b52819bc134cbc4e9188c9374c80ef852dae9e10250f8f1
z69957b5da24ce0cef51c7021d9ddd7953b7d5a7ba6a0fa0d08760f1399043fdf6ef4b52a1415c5
z6c405fb1dc8a4a55cc6344ad47ae5db0fbcdd42e4f6cd1425afb9e6868b2230064649d6d528c58
z39d5580da4271a2679494a4edcc4149cbbf78d6e3c30216b5a5ae0095a597e84dd6975754c7969
z6d0ea57bc6bc206533fe6f8b7d9c110765ab583edcc9af70881de3298a16731455c3eee605024a
z8c994072ad49f22cfacc65c81e240ad4d4c03dfbef0a8af5f70495947fa2a217db020f703118f6
zda55b7001b6c98f524adf334f317d7a8d603ed51d35735117f90884ae845a06670c8803a72f72b
z28f17fce6825ca6702d823c77505f0861d28d985af9f1c9f8a327d3102644cff11a5a71f0ff073
zcd3c333ad08681abad2a3b8a26da9bb93a41f3dbd7403366cd72f0d74cda3c1aef87e1c096031a
z3f4b269f1f1ccb87fe5264b19cc3bc06f114e6e4e497a7d91a3308dd151f539f17a005a0319a53
zb9cdc12c5664a51d9c8d1046c9e6cc171a26d65044b263af4b26b8f0a117117009cc046998ffa0
z72f1305b81d6fad9bb9487bb31c7558b3398c85f4c61bf6354f9ef5e297f4e33ac04197b432379
z1d37daf38d2bebcb672c31f31f142789233dcc1734e3ff5d29331ea48f1ac6cea30f0cef09618d
z7eec9a85ec74fe8021976080b864aec78fd6a0072d288eb66ab0d2707dd637a02763787da06401
zd554c6045ef5768d819883b967854d534e4c1158c984c14284ccdb0eab8514370a71921c817c8d
zfbcfc2c01520db9bd7cd4dfe667d451bf1b261ded98d77fd35c880f5df2876498292108ff4af32
z88a6de3b4b01d9875fb6bac35b698c266ec1ef85dc73fb84eae9d0820c01a781bc1b8690911251
zba4d4dc572eea5b2637c34fdb0ed095d368a12a03d8f9c749fc1f09d0eb4ae81d068875b01bf17
z4436a5e86fb7583d6adafe74f5bd3764d7b3eda71e46bbdf385787ba61d00a2a8f4fa5c9e574bf
zb163a5f6ceef45624397e9acb65b4be477e1819988d815a117b8042aaf38f600624295dd7ef269
zc24188d80fb642b7d8e4ba60d8572f7c7cda68f35d8b3a6c01d8a0d2bf59a4a5d8b04fc046b5d2
z963805e1b1444b7f15f118d5b6ec9d67bf34f31a44837c01e773d574e81d6fe0eb857863cac555
z51803b047009e91bf90a1e3cd9f8fd2e59117673d4d87d66b5295606be2cb9558832e34c534b31
zb6755f3972fe27a7228b380b90007703422691f44b6cd189631bb4b668bd6381eec1cc02502e77
z6a6f2b6e12c012e53321394417606393e2f8d10058ba76b88c1143d08536c0b25b0fab41364f6a
zf41216f53d400753f89b20b28edc00c0ebeaf57ef2ee45c1dd1e8487f3bf878f6dbeeece614b1d
z3f7cda707ec02f2f3e72856a87cb06c202e50359cb51322e5fa9bf2751ed74139844455f39cf84
zf593fc1b9d905e17aab60678fcb5ef96e47bc10d8445255331ae42fe2a5596956d9a4e6f950ff2
z800571b5d800d02ea6cdd1ae60e71c8be40416a0c1902ac796084e3e9d446b7b5e9c731620f1d2
z24427f0950c50fbdef79edee1ad7b99c11cd0513b0c1340fba53940d55adf19b1c3d63c563a885
z382093bf49a1b18765045c7286e6e20ccc4335c2742df35c23772627f72685ab8b72af44269d17
ze24731291d8b484ea0938a0179533f6651e76de12dc711e3c66430127954ba5d765b9ee6a9a52e
za2b8b958d88d2045d65803ac15bb445e18b995de1c3d48d74be215b5d0d8e4971becce6780ae8f
zbf385bd2458800eb0bd4c9a5f1c64ca6f5075a415f99ebe70ecf671d78b652fae19a6ec3d3a135
z62a1bc0e07b107da76a14a862dd80595002569d47db0abed40818ab638db73534819e3d3df9b85
z404a246253402eb321b6d154996c207e4ee207469acb9bac2d43a08493ea887a27b5188232aa8c
z6efe0d0ed9da83dc1cc3b4d10d8d1fe4f55695a991ee05f3542761f7d2d8b180f72e4ca5fb2207
z5c6f5e4c27d9c1c65ddd9cd2c43ce4a47c4072cdf67d61a2ca5a9ba9ad88ee0407b412bbb6ae99
z07600f93144361d790c806eb0e356248fbea2b5448179c84b8238a5d62b4799ab8dcbdcd1f6f99
zb1dc16e8817fa0233f680f95b84941631ec147f07df535a727dfe68183e93054cd02a1ba3c2d65
z95901e602d099b6a83b8556823f3c642fd565fde94b9d30970ff6b896d8d19f39f50e43d7bed63
z70373b728847c4b8ef712dd03ba5a8b7cf8ae6bb16fe3af737d606b619d40383726c2230fba44f
zc28c209c08cc54b51f1804d6e0d9a95a4bb0f27d6e047bd2191f3c283f5dd9b31e450cbff44818
z1dd007b27f2cdc0d5d40cc848517484abfcdaaddda7451b741a807ead6a19309defd434206c64e
zf3f53b9fb7e01b66eb83988e32b2c431adcfa1fed46a83f6c7e66c81fb9e85dd428ac67a2517dc
z57f2711a61c4e3bfe54360dc692680665722c32aafc35e51ed2e4785895736c023c399a8e6c9fb
z70896235db38ef0d40c806d6988516a0d4c3d218ccd4039f6d990fae94dd6e02138d81f3f4d785
z950c3c1cf1952f0979a5a87db1ee07058fc83261f56f787866a3bfd89c8c988ddcf66fcdd34391
zfb371196e9adea596b251c8f9b9ba403f3c7dc161c9b2492a72a36249ad9c4046e2d7ee100f41d
zdc3f44fd23153c58e74dd63caeb5757c019bdf2d15083081eb92800576d6a0026bb4d0ffcfee78
zb321a1a4caeb07321499abe343f54fe06e14e82ec47a6919e791ce000314a9a875dd3057944393
z06d2b10c6ec49baf325253c9e09059a8a89ecc4450d9de38c67dab9fd012a54829268a68d142a0
z5594fd745cca247aa187b94b061d9130098b15a9020d5e4aae78d23f2e27e1d65b5f75c1213d70
z33edd6e583ccccedafcecdf8f0a55be6f871c74c9b354ce1f6faad98c761b1698e9635236f830e
z07afa3cc2745519f71cfba0ce7c574b3ebb071b3ec690219a6c33ae0f24af34d7aa19e93580939
z0623628a35cc7b736a742584288a533d7deaa6bee5e09c75176f79b9b7d271497b47ac19391493
z8e590cb55a9f89606e4805ef574e16d7b6792bd116d6a730faedc9297942e3dc00ad134b5bd2d6
z0f1b5d38014f17b90ed1411b113da0054e809af33a7b5b4b8b157069d581a2ce4d32f5079da571
z8cea38ad02414002c78a5b663627debaafe4542cad080b5336ad1fdac6b32553f1b0c9fd5be5b1
z0238a7c67ac4649c15ed83f8733f3d78f405e21c2206e914b74088d4f754a4dbf97ad94bfec17d
z02e7978e07f1f52bea7b574a5dff8d75f95d31493f666adc685cd33c16798e600ab8311c806593
z863a99c6abd62612e2a2922427b0da53562ed1040b099d77d9c4fb46b39e7f57c263a4f1f6c428
zb7f389317d67814ede25a340323691b5a16591ad519778ceb422736f41b000f4995eb146c6addb
ze455ed47676f5947a2d1f3f615958267aa854cac1d875d05c02c006ef1e19fe471e421c83538a3
zb030f789181c3618f1608025aaa80c70ac57a9e0a8592683df179dc289257fd854825c81f2ffa0
zb87f45642ea19dfbca09abe8d58fdd68375e88e9a2ec40e7eb939f3f78d98483369d1cc463c57a
z0027d1daf3da4eb2656f49474665fda5bd835b68065ffa1c409fac340a4bde196418975bbe7583
z571cbc68ed43d3fba2845c70329179e689c99f149d345750685641e6cbf367c6ff19509ac7e92c
za64c8def3680ddbc974dbf101b2c695a7606561fda68a03e7e7f433f530604eef9f39e1707cf40
za5584728b4f5cb35374fef77ed5b6c64116965458b61f65eb6ecba1c0e276bb8d17f5236ed9cb0
z923fb0fa44982c3ccb71257263ce8c289cb6e6a6f73f5d6f5ef534f149856202c01fd613a621d7
z746583e31b4aec4b72018ed87361cb9f9740461b2bbd062142c92db7aaca8c1d9c5ab71081ee74
zaf7c144249abe6a696d3d00f4b46a7fe789c847d32c0d00bb410a27ca788d66fa4b5451d7d9e37
zb62f609c95a5cdbe70e824d26c67a5f591692d9838c4557b726c9be75aa87d15934ba3728c2920
z1961a615fd9f52d0c15ad20533c6093b950066eb984c64a94471f0f4e71de93bc73315add311cd
zd3818feed8c1c902926cd9456125998c3b872b3e475d1091c6ac81d2e6f15d697b0e8d1f548b47
z2ba96b428822baf1ccdadabd4a2601888e27e07f6ed68bba9c974a9c3a2fcb99e7f9ce48d06311
zc24cca035d717a4408b737f7f7a6b11aa5ecfe7999f63c0ddafe4642687d7ca3d74cdb4b59f2c5
zd6d8fa13db4729965f298327b5650e5a80291f42ce3fcd2cd77e57a38ee36e7da781570d08cdf2
z66134f5eeb76d6dc54dd672a335f92e4357c2c64fb15a38f34c7cd4f8012c2990ff621a9b7d1f1
z9e0391739f5103d8dc640be93d0abfa618efaa457de0508abbc3e95f7e36745203df70aa8cd2e3
z8d65448a4f553e6a759ae9c0773a0bd65b8702e72a7fb8b01238b61f65f8a21b07b91b93a904f3
z95944407d858ffd92fc6d9eaa216b109af6828220069c04b4644f5ae790c31da21035561d5d244
ze8a92f56e1202c8301f2b3e98aaf43cc32621e1d197132861be5bf25155226255fdf1e49a8221b
zc22311b64ef2a7948aa9a61d5fa3f6c1578309bd78dc3dfbd5e7115faea91d2619c187919cddbc
z43c29c34a5c33f2ccdb7892d4d424e64cb55f028df5e945b2f93826f65ac1646a35c819b3db4a0
zd1c077cb8305570b2aad6e40e306d89703fd1ecbec2944a109321641d7f716d8554d86ea000276
z70709eff2c73a823f9ab5ebde93d4edc4ead563e69aa5509b331417c2e5d89523561943f110ca6
zcc5f206659e6e3dc39b7c2c9fb2a4f378c7410277fa56f93fb0b4a26b95e0c5ed9d581e552ac86
z77499932f5880a24165b1ecd8083c48ad6d066cf3e623712948a4b90e9cab1c1972bda4d49c605
z19466641fa0ad485986f4c3b4287dceb1e3195fac5401860afa93d5240fcedffad623b7cb0f8d3
z4e2c85448b55bdb9b967d0071e25d0688fe4ff17870ad5dde1cdcf623f41f99916a56b01b1bb23
z878999055ebdea508e1a425b4b467e1fb94314a88c6290e35dfea5e1796d8ff6cdbd2e44b31ebd
zfe358c9903f8ade0a73d06a9d41c290a65109dd4be96a8da6dad5d93e6bf7daf91d12ea42f640a
z41887955b29572757316352ee5f94f2a07c42a5d48d4e9424805d1dd07c77c600e474cd060afb3
z4d62a426a0a1e53811e0993c9bc876af79d1a32d83e52c0acfbe9b54f798d429686ce8398613bc
ze022210a6a6a6ce23adf605620af43f0f9fd2f243b2876db44d06951a22cf3e16711bb70884af8
z431c571efbaa862dcd08d03867ec6fd75f95012a1dbe56a7c25fdcd8a71858ae525ac2bd357cf1
z567ded1dc643b9d270cb9081a57e8ca6aede7653b2a2cd275a134be2672ad38e946159a6b58cd1
z9c12b5e154c64eaf50bffaeab32fa82931516e754082c49b1bedd0c167700efe2ca9a18a103ab5
zb1b280340ef1668e23d6db9e4e15d0a418960051f608ea6a42a313de17162805a48d3579f886e8
z2626cc08e9fab35792cbfd36c4fae050675c66ecf8f561414a764a0d5c1759bcce3b2688794107
zb019d4271d939703322bc0df7b3b05338a687cda004deb8f125044d4b29a2eca33188547b4a335
zb2c84f6c1c1cc31142e58ac37cb274c9fc46336786e3552c9ce16046bd5f04f36e33484612ec26
z75890f4abb8756d83f9ef90e25664618676684b05f6dbc9421eb50fe261e6f89687cb47b68d24b
z5ed6213d6891248bf88711a557c1bb82ef28b0c83b23ddd323e2a4ab2a5e565261d404c3630ae7
zc3cae00e2f40c1991d59ed3ebb675b69afb84a2bb4793d18b262068e1fa7297ae5d60bb927b4c1
z28caf170c9ff747e1590e9d905e2bf92f14d70e5c68373142d4bd1dd262ee8b47fe310ed7da958
z739918dcabf0c15c9cf11117a3303a912cd999bc98df6f0cd6142880499252b8ae30c0a1482d21
z6bde9d52d1518e1a730577d3b51bd204c48ae15fc44dcd6d2aa33d3df3e5d5010e62c77819b815
z62af51607ad35b5730d83eacf020d6dd807c8a4c459024e3e7b33a61896db5a80100e75eeb34b1
z29b879c509b6b3ef53a0bbc7466743dc46af8ba08e86548705dcce1e3cfd0375c8d2b798ab83d0
zb422f73c4e917ed2f88715847f6af0007df06db3c11232f4211125394e943d67c4b5510148e32a
zecaf17d38803177c34564779919f41f9724c841f2202c1014a6c2191edf3e8f2ffbd37c6133ec2
zb99823cdba92da7010be9f60c5bfed90f70444efb5fac70b84b3a6daa98125b3d97fd7ada71ee4
z08d9bc62974dcabf1cb860f398bf2f1a5f9e97409008adebd0d24a23a61992de27c4190e3f55fe
zd299a4599684d7a629f3fa12130af7ccd358191eda866b290e1f91c579ace8a8eb698a32eb8fb7
zb762f28220452ec457590a4c5f234c8aceb3749304c2b46872780a466c1d36c369e978e5e3d4eb
z9ff5afb2a27e280e7b4c5d9a490491afc269661658bee59d8d170ad65f43b006c7c6e51544dc59
zeaae8840c610488fed412b33cea04b93c7aa503cbeeb775cd4be77b65711489bc0a249ee0e03ac
ze5e01331bdb85d39c5cf0e37f83dafd016b653c8f95ec95bcddb6b31674bb5fb5a6bd6e9a97efd
zff74da509f1363f4cffc9a6a759526b5dfa14a6813acd8ad7ccdd219a2a18ec24bd21173ee6e15
zdda6e072e0339cfe44acfd94aac92f76f5e7d2fe5c13ce4a6474e1735fcc415e67cfd8132d994d
zcf712b90c19d9b6f6dff9b94016406d5bc47a3736e5a7ca986769d774068de6fce0d651069f240
ze7220f531a0ca8d0186cef63059ec5c21303e62ade304618c3a57a7a97f1d811f87926aabe6891
z32bf82ef5888fc7cbb01a9a0712b24f446035dd98ad131814227b4bd0ced5823b3274d78b88bbe
z18d7998bcd18d573c7ecdf9a1a5e9afef78dea227fef3b4180dc60c515408df42b01456850c37d
z656397508a92a285ec8d41cc8d41669a4c413eddad054af181cdf6b29843da229500862c006434
zd8f056a764dcf6f531e4109a4baaa285508a45b30cc4bc702f8f475c3a9a1a9cf7e0f825445d83
zc52f49e0e2596c6f602322095fef530a3bfb25ea2de51a8c4b42361c88a955a8b8481cdd082142
za6d40ba70a84772113a14dd89c9a66203c04cdb5686aa2f9ed849aa78b65251e4b84cf01b07958
zd5045bdc71cce90e4770d60876206b4ba9e9b369aede24e81ee58bc339624bed765bd2bf3e31b7
ze012e826049704a2507b9514a519520ca6e13f5bd548a3ffb21afa32d97d649d24bf833811d616
z6f5e415cbbfb35ca11938195a86b3ba493a209ff60012361b1e8ee69cc3dba30ffc5c88c574389
zf3ee6f18f8ccffae83018cab56441ff0e6ffe74d884c159ce8473adf2f32b5d8186cfb5289b2a7
z7cf881209862422d512c7e2226de37e10bcc8a823fbbfbe4fc45bac3b14f100c2090c5aeaeb94b
z28ea64cb7f9ff202a258d76bb81dcd7e7b44ff1271f7b7efa79407c1bb1cd8642a0b97b8ed6f08
zd1b6736e62b58b70b6b8e2a7518f13ba7fccee08bc908fd885f0390861326529fbbd524525f78d
zb4b07575527967acd00ffbf9e29e51b7c033013b2444774345308ec6ce91384305f4a529f2b6f2
zeb791b644114ee3e0be8b82730e4f8bd15e6c4291848de94c0e374410bbdf7bdcd6647f909cbf1
zcf2ab43cd36a0f9f313b0029cc333ac39fb4b24bb070b8329ebefe069e824fd729821bed4c2e69
zd5d89a7b1d9dbc6f288aed9495ce9f129c0f5d71e86b9263454f69476862ccfd438804e010ff42
z02ed25d815fd6142929d36d333e8e8915c9032395d253a471c840dcd73d41d5fc162b536bfa30d
z63cb4f0b9880653847f42ff219edfd86301752c3749fd0897b27008a23546adb21402e6e9d5c4b
z8ccb29a468bd47de2a7631d86ca2b1e1996ac98625625ccb057417003d3c3ed2cf47c7f6fe38e7
zd93f9d746fcc79fe3ee63497544f0be2beda8776e253a75d53b60b8cb4ab573c592e2f321a2d87
zf9ba3e4246bef11b73593c8a16dd84fce8515901339a3299bd9f71976677b3643e327458712709
ze6dfe6188be770154343c3cf50688d398b2d6da63d1e824da2234bc1c46b93d0eaac94729b0db9
z68a19407a7d55b15457e88dc88bd48aa37bb7a21e563a80f976961897f7d763457881ef4f2fcab
ze44b93a95e0d322c4e27c7787b40ce40311aa7197ebf8340a196744493d548218f0354ff0234cd
z19812c215567997acc384f998800812cb455e741847eb53cb35d25111461f0c0602194ef06a4bb
zca87716133ea096bf5744c291784dd12372ecf83b1d5331dc4d8fdb8bc3530d305d0228165a709
zd3f2c1c3ab7776f233c40f779c1fa6abde7ce1e26443468c07f264d0938e13e792463c83288066
zf1cfc07bff4e2e569b15ca0af9d98a80673edd4c0f302c8a68e964689ec34052fbd5c2c4ec4d8d
z8598928018bfaf7ba458571533dedcc462e86e2ba9abc96b25343a30336a9d722be1808bd5488f
zfcc13c9620bf0e06c4db3c98d1276b533bcc9571b9fbe33ce2a00290d0686c8335f61f64272a61
z127941df1b542ea32d06d04c2af16d0967c7a0175126db00601d7cc97040920354edb5912b669f
z675081da9766ff2969cab7376e4ed3598ff30b8a5dcc904f479ac9912f5d4e34d5a09353a9a82f
zd208499fe02d5255fff5b25d1f3a6bec40669edae8462a6adfdb4cc15217e3b6a7e9adf0d903c4
z86aa8f5b5e486b98d56e10978308d7261daf9a294c393de3d6daa54365e6f1f23eacf8c18fe8db
zc95b6389d198e3505637b1b95d35abb6728f78c6015d1242640c6453ac2a81325558f734406cae
z5a66ca0638175d577f0bcb77fe17c3d3d653c15942884e5a4573d46cb1536748167e6333617436
z08adb15efeb5b134d2ac0a3fd3caed52b529e11b723a7ad827a5d83aaa54a8df75bf277cfc0513
za434f1cc48a2840a9e0e9296617e8aa6d510d558db7911be26d9cc3c8396843a8d145d938eaf05
z823dba67ac8749187d89d19ef9897cf79c3b5b32495952a7c8debdd8c0c104d030e1d314ab36fe
z24ba580c8e0415ade2719bf43686e71049a37197f8f92fc28c9e8d6670dc9ce9d43181c2dde3aa
z43452fb2b07461ca4790d4df507345f9b483d001a35a31a89f1d8085a5c553f7521239729d3b6c
zf220d66f301c9f43a4aa30ef7f818809c9821789849209961f6c4e11fc39bfd5dbb32120805683
zee6d29b2c8090b3708f3582e659a61f42c7f10fd0c31746cb4d34cd7c69bfa264e77c7c4b6eb40
z6f36bc87ae212c9586acd5e2569a4fe0f291e7f7f96f981357d5dd60d2444adbd832e586c671fd
z14e63e436f22ef727a23b79743e267229c6192aa78d4df0225dfa7d5ca37138ad6d7d68bda3165
z5c48c59c4a3a93b9c910df7de93430235244fcbc3dd4416f7c0eb53970b4072d9daacdcfa29f2c
z8b22347e4c71533fd3f68cd181ca5edd86abb0844547b4d2e298127f51d35a31ffc7e6c6b8848d
zc95d7d2897b822521803ab57a89ca65275127b77c04868581b34ad0067b33ce8c031d4383c802e
z428a4f9ff7a28ec769ac205d53681e610ac71cd9e827453d65ac0e9c1595e11b5492c22f237cd4
z73bd808dff14ba73b5050c7d90b05cdc22e21d4478b6e78c908caad5216fb73594518bcbc9da4d
z79b3de26c107a17ee48c5bbe26f9f7c9539fa6f0093162bcab5a0787efd20484c2b5c2766f9110
z88039d2317de50f410e886e58b8646968e189d8d5313d4c3ae8dc755b55174e65f44769d0acdf0
z7dc6895f9f1cd512094df83d34852f0ac54cb33b8cd3f9e23733b4e2fa70072a95c1a939a11201
z9d58745bfccca17d29d7fba58214dd17d8696902772a1d37db47ecff8fa406b2132728020835ac
zd29f04efeebb9c4e46cf88882acca127eebc1fab13aee3d0603e87fdd80fcacbe1686c55368906
z36ae36ff3d9e3ece7df7239f04e6d1b2217ffc141eb57a6509882790aabe4f66ca6da610ea1ff7
z68753e43099235324bcfad00a01ed3b285196b7a053507285f30f476964ce5d9f1f9a3c739c2b9
zb8483490fe60dcd170bbd87256e80cf8a7c4e52776d5ec567f4f14224b18b3005d30e9dc2c8b37
zd2d333c359f95b1637679c976802ff0dc06546b9c5de477990733c21ff31acc9f9684624c18284
za229a06b241d3aae37aac15bd655f623578d223561b543703300caa99ae69007f77b171267e922
z35a2bc5f2d69e6707e365863775c4130db399945be52e654f52a3f766ecba210f9ad3595c630a4
zc82a34ab418a8e507493baa5f25e6fe23fe1d82ac41827670878dc1734e496950ff4f3c52cf37a
zb2e4b58a1cce81a4258e125385029883bfa6b5c55b347fec025f752711d24e820e8c695614688a
zbde6c3f84b61be636642d7232fc68ca546fbd326e42d6d872088824206cca741c9696aa890197b
za545598d3eea042d09ebf0edfa3058c71223386e9eeeff2f447ea86c3f5cb675c61bf0684c53ee
z916bbe294444dc45fc8136166b93ab6dca33c2a6c3513b40788ae808833ca33525c635bd7bf241
z4407a64bfbdbaaa658afab90f35b3e5a68208e12fc4925ce122f77c3e8badedac0c5d721483933
zca1daeb28bce766533add1c657eda9d4383c91ff86e171dd3c5ee5c5a4f86bbee276c8763e4684
z97b7acd815b22bf9ff20fe7a9b55533db64f23bfe984d8637a8e79c1eb162b7be4b7f7a1b6823c
z2ac0e0cf622770d5dc83819fff098b88c914f8b31b5d080c1edc0b7ed27846454bd19c127ca431
z5928a2c6d109c46a09aea26a3da9dbab970f1c698bc1b0201e949bda389bebd5d77b28671d29ed
z0f9010b5bfea0674b7406d1164101268208544b2064e54c58e2efdec2724419f43528ac9349208
z9741b74dafd38287ec10809313030d845c9818c8481585f51328de071a72d7f08f9efd6f0667ab
z1c92b71d956a7ed3f75e69519599530ce0a94607ac1b13542913ebaa0aa8b4d49fe94c9a0b5951
z87f5c6eaf35ae8755cab742b9fd3b005bca37086eaf9fb84d98462dc658bbddbb5e819b78bf62c
z9fafd119cd5221a65393d18fc0e0d917e7a2e3c1a3076104d8d5e35de76b7422cde9631d47d20a
z8e29a067de09e36108f067e84c1d65a40e90903b11b67b5f7469a330ca3989be08b3ddd9d4b146
z0a0b41dbfb5d072548e527d7a555745e704ea7ae6553ebef2062e6bcc499811ae5f8fe0b1e16b0
z1e966c59f4b535e2413e55a6b14a1a186e6bc8aeaa2ff9ae41c4599e926e766d97ba86bceda640
zb5ebf458e72b669bdd73dfd02216f30400c4ccf667bc25a28716c7fa62893ebf5a02cf8edf58b9
z313f292013e21f64bb3cfe3cd8a6da4e87bf461054b0d5fed16095021f4200a6835505b35c0d38
zafd9bdd4e265728fb5a30b8b92ff1efc56932dab7af1633ba00036f9579cff86064b85984c1d8a
zfb822d371a53a6390980375f6f762aa02697bdf9429a7df27fa6cb4ebd7b1859d1fd461ac3806f
z33219924796985a38fc8e9c7f2d27f47786ab90e4dce90b6d0f100072fd50fb18d5162f92618ba
zb0e73b0dbf26640dccbbff28e564c75bb9b2011dc3620807410122170bc27a4b33f422b9cf9310
z675372a4b43c4c42a75e681d594aff72d2d757d06a45782e287e23dfbc629a56b8a76337c1ebd8
z1ba00b93fd110cc1a0f2ceabe4bca471e4af8bd5fbec8f766187373279fef463cdf304a0de9e8b
z4aa6a70dd5bd23a4f36d58aaae4f87331f2cb7a20a36d01de160436fd3b5b86bab0507252fd004
zf243a39cfb2f2d9673f7e4eaee15f6162f4bd1130c0f61af38958a42463d58a72f0b79c28f01cc
za5f929587bf3a9f5acdecb2f96ae222388e2d76c90e28ebdd0e57397d08eb7c3ec800458180e73
z609bdcf273e3906c195a505a4f04fefe82572e95c1277d42daf45e82dd292883145ac627e99085
zeade6f6f5b56347db95468d60192795cd07e30d317b4aaaccf90ad227a7a22b75624560bbb6685
zb61ac68c09aa8cdf265ed8c803f50840ef5bba5dfa93e192a95bdc19c49887c8362b447c93f403
zc9f4429107690eb3f75c2d6741b0b739adcc4f654881988193230719123c457cb1cc57f2b365c1
zfa9ddb50119d47922634e359862d264d92361e4ac8cdc3f5f5a304f9fb765296984a66ed4db7a1
z0c731c0ca345cadda4d81d72fc04fc8b39e58c94085761d0bffb5f6d4208a55d33fa094926e2c6
zbe99b87be5525e6cc4c48d3f3849b354a6637c9e4f42a52c286c4549ad74737390ccd0e533aee3
z9b5531d91485b572572ceccaab8bf18b5db1568fcb2f8416d8c8a4dc3c1ab39a5d9b9e5f9faefd
z70bbc5f12e871d7bdef9e8d7f980ec74c5bced0eea0eb4865d175714a362f3f21c21d7244508a9
zdd88bd3595d25816236b61cf5ed27829552b7b69add9fdc071854f20a981a8f0a57953cb856c77
zc44de3f26d5ea9674c0c6919b7484ed6879b455bcd14cd71d4cad419c0c471a86c54d53e08e12c
z3d3162d4d1037bbf576db76beeb928267f89a80ffa9dc8d8393e47d5828a726e19c207f75b7ed0
zd0bab86cd0ea5dd1e074d3c811e88c2283748635c08b241c1ead19720dcdb22768c55dd68d0040
zb761bd988ab11c3a3e511e40deb730684a11142e70d2dcb333488978cab75f322e29021174f203
z0d861851cba6f68bf75f3464009c46e2a084502dddedeb094948c9dd64cadf87e4bf7ee48a800e
z24df505a47d8a1a93747c1f10ffa6baee468dbdb1d22650730b6429372e0a88f01e39dae1663b5
z0ae1f8e82fe0ea969c3c40343a4a369746256006872ea38ef710c06688ef272faf7274133d91f3
zf48ba1cfddcc5cde2ccf007c3785d65ed9181ed319ca8b9a6d4af32575bcc63cee783efc020304
z3f1c5ef75accc8ca9bd1c410d696d095d8c471f5fd79dde65a7398bed769e64eb6e9b929a8d12e
z9928893483a088310e64098c7a025211aeb277c711c34f20589484d260458599acadb2fe94e4fe
ze9f13ebc0a9ba4c1ebc7fc8fca179d8b9e6491a0b71b9b0c3e2d30f44f230c1ab409e21f83a310
z2ababa2efcb5d5c63b4c5d810d348f33f888afa6bcab165cd7d6d783c0af940bbc0f6adb96cc06
za0b7a25a12175105539005cf240f593f8e0b1f1fc09ee4a49ac2487e75186db07efe77c89c0302
zec7c6f0224021b2ee32f6be16b342c19960c040f99e2c0d2e89abae3947065a34258f7a29fdb5b
z80830fcd13745aa83a43bddf4f7b468f5e5c5ed6b4cc4c7c05ea78d64fa094899990744f2628cf
z51e5358dacbde230a9c219c7686b56963977bb187124bca588facee9e760b8fa22ce9600e1f895
z092f2f94759e03183785eb3dc578af0baf22e08ca59598711c231248626908853e18ed09393b7a
z2a6005128ca529160d07b44020a61a4627cb9c0a01dfd6d4279fd1f350c64fabaa429f7fdccdc4
z7fa0a805490cd65373a2ba154810cf79b7544480d4fa1d83893d1f419cc9bb59f999f17193f87a
z4b07066394e4a2bc0d38f67ebc865c6e66b40aabb39f869c36365b30be8b32046f12c056104cae
z6dbf7b2275311ad41ecd37d46acd7fc3c85a5abc52fcfb74d8ac19a08d3dc96ab4dfa6094fbf66
ze7f4029845c173a8717415e267e133f006973f32ab8181fa2caa2d5a7248b8b4dfb937300c6e85
z6bda3b188b3055e4451842b2945b151f46fb2ae918edee780e5b1b10a882392dbf0708b14c2ec0
zb372c783e03f866aa6fe61b8aec574409d6482a83184389c131edbb8394686200b2a6a3a872138
z3675612f478eecf1481c0ac2da299f927835acd7d411c9e51255ad33ec948f81dee44133fb505f
zdb2764d68371b87a59a1a7d276e76d26e9f32b6dcc3bfe6beb3ed2b2cf4623725d63f3b8531408
z68cd440ec4de9fb021b5de7a606fc4675ebff8066431ebcfc4a2c9402d13912b4701ec5f250aaf
zaa49ed36c119fb36cda4516b60a345f23d7936c1c231f919d1920a181bd62971ced498279232c6
z28c14ffc0f562f87967b7e6e37aa9f8118ffbaef93900457994272b22556a87fa8ac5856fe897a
z61be19a9f9fa85dcafd526311e455dd9e3c87d088791cf2d288d5aee70dd5572935d0a8b49b1cd
zef1af6cd6be1815135c466153aff928addeac1eb8d56851fe2a34f5857bbf2fb10c30e7453281a
zaffebb68e5fc2e93a90f5fe43218280c298778caa4e9a754c19cb1dc2aaa563536c6e8b3c47380
z0a5f77f181d1f3a2d432d4d279e83ab0b31a6b06de99559b2fdd362486126793d099aa3513c010
z0b48651e845e3670ec6481d3b01d417b58871a1d9635db0761696386d19a4777a353cefdbee6ee
z3a5c303b1f4dbf5c37604739a98344ff3cac37ccaec3b6a473fcbce30c7ce81cdf485f67f42903
z96fd87769f660aa7365c0498183cdbc770ce2d505121cc4ba94ea858509f27013ca14f75050486
zf7cce85be4cf8c3822e349b2f3216fdaf25914d9489f1e5dcd86492b100351bbac58c5a855ee66
zf7129fe195e63c1563240062ea7960fb73cd5a7319420df973f206fcba661f1d9d01f658499ea7
z67682361aad77f35f78150c8e89e1a5d089fb8a4626605df147e25b77b0f573b5ec7651e810acc
z9776c8151b2cf9ee33ff60829c8079b371cfab3dec238c14b02d9626cd8dcfba730fff1f7fcec9
z614e78bed3f5f27910ee88c9cb0ba6f755632af633b92464e6bc8440c9349ce8d3059b8ee645ec
z2d1a0e145a254cc2307e8c932ac7b1573c69b4220e7d21915c521628e099aaac31d33eb88f1881
z43935bf7214705962a91515a99934cd3ac424f5064791c5ee827bf46d4a9dc027c6a8ea0734d46
z110dac41ed14efdd3e3e555f179f0ba25924e59756da9781fa4934c938995796927440b0af183c
z4c6dab0f1d2575348bb10f20f45a6ba07cd06d248cb64c588673377612ebee64bfb04a56d8decf
z5980ae37a5f6b7b840177f666eb529594792768eefe4df3639ef868d8c035a474de05943e7b329
z7a6d7638d3919edc4d33b85a2ca1fd0a3b1c6ee69c9371952c02da74445816e541f5fba94b2ef2
zca619a176045b31252501e6b8cbc55f5f64a64544661b39011ec9ea8a4180aa4e294d6fbe8494e
zb8ab72c68d64fb771612aeb8aeae373cdf165f220d11edee767ea78174d7346799dbd7245f4273
zdd06dc69fda4ef2dffa97d58253698752732b075249546c3bf601534ff038af8544a3b022f8d36
z62be5a6f1542ddad5ff7d0f8868051569d251607500fe86e9cecc85bca255b9ab61a2d32b6f779
z439d42d2b6c89cbb805296366ed62776abde36edebaef7a63a9d033d264fbd386cc3076ccc9ac2
zcaca648a7176bc3347e2f0091b315c2ac26c3d2a20819306c8c13aff026533cca7303980dc00d1
za5b586bb43d9f19cb614259bff886d7b35376eca87105693a45531e1455dde29a71f7118af2ca1
za05d81133645ac8d7d12a528faeb3ccefe625566ba4444a265818a2c2f64ccb6edfb7caca1c370
z403705501d5862efa32ac819802c911ec192ed781134f0a0b3783fa84c55aa94f37733f670ae1a
z9af8a56aa2a8e16e6f0f2d0c3034b93d0fb5053f11647c82dabc7aa68325fd33d0cc8130a0ded8
z6d6919fc61e1c47a6a9d6bc3fc9d18539035f7224d86726d316330d746c2ca4c41702fb1eeb184
z023ab33a2c2c844294cfc63e60b642379a3b7cf21501150a3aa5744f9b8157043aa561581a0fd5
z15f940bc1e437d3a57f7f0479f87801a9f41a42f49118e7a4d8845462e61244e08ff0c38d98e14
z3b40b845d4bc7675702a9b0b07838ee5d4dba1d3d6335dc5684f0ca19f52c5b4c2b0b7ae3a2b58
z3c6c985dc54bb1dea16d3343fe88dc80beb5699154d4b6826167a9fdce4d3c854043b652a51127
z174e184f59c59d375c036f4234cc61e0f0233228df77308558b11fddabc6c10924042ae653d0d8
z3ff0e08605a8a9841e5ec738c851f4591c21115bc15c8facf77d01e5a33d2e5788ef95ae1ec322
zc71570e262fd19f14ce68ecb9885b642fed86327e624d139ff976b84489d4fc276fedb45e03dfe
z33c51eef54145abbd6480fcce508f5d9fc4b63b3a7a64a2d08c64ab806369cc814d9a3bf7f0fd4
z96df7e38cd1213a2e56311216b08135c6fb080bc42445e68ce978c264390ae39a85cb3c0195526
z131aae4252e27acc440afbb6f9934e06c8da5c8807d0ff00008cd55941ed72e126122bc411e2c1
zbc6c192c41cce24cfb53197c973e529b45e2d48dbf9478e97f4f88956fa1d58bc23ff03098e615
zc8db05e342fffff541d1796e339c65751e379cca2f7157c04d187d49759f7b0fe69bc467423d49
z61d2bf05cf010ead29f1f627ba86e3026a13d52042f6a01e6c048ff44a43900bfcd5acf1c0380d
z04f31a32b5d4fc5455307679eb252525840ba34e2ea4b79befaae386241303facf5f4e54b95228
zd8aef9bf3bedd9a6db3fa8b60de69215c8b4fce4abe7e9c3a0525613f914c24050ed0f7c931670
z67ebbc38ad1c5f23167eeef4dc35761763025c8c4e3510ff98a265c014d52ee5a7b9ceb58aea7d
zb8ce84fc89335d63a9bb32da9edb0e77bc18a37a9920aabb4ca47e3fb56f44449793af8e4bd920
z81a77c3b722788ac9bfe4df23e618e9fbbba5582ac84f3ae45e5af7082a6e425bfcf00d80bda1f
z1a0559618dc928d013c0548b7885155ba9770776867c07393059eaf95e60ea44d88d40f6141d69
z94b5212be46360ffc19690a1dc717c44fdcaeff5d8882286c32751ce39d492bf4e98ed40fad6af
zcb8cc949f0e2d3baa27d484d53b0c7bbe04709e0b8427e3b1235f8d28d2ccd7e1b5da04bad1720
zae1d3f08a6586305522a80af347d6c6c59fd4c203b4ca880bb8c18e0b8cc1cb1e74184d586bea8
z86fb58ab0222a54d29ea1a7b0b3d89c8a8471fbb8a71b8813d5276007ff292e1f1d8c0689fd2a2
z78348bb274e5d68bf739c974d62a9379106dc73672575776b5e20ec0d2f0cbe5687bbfe46682f7
z4b72d7cb741152ff1ba4e2a0b3a58d69604645d1329e095abaeca1d094064d14fb98de576d5e32
z0cd8737b7d67146c88b8d80930eff4c6796f66a8c0adf5dabb6de7a8235e48b0b5270766a88dda
z51001ab3ac68e7d719aa2aa29689fd78cbb50cbdca1467539624d5107f0709052e311865c78efb
zc36e06935ab968c1b22039501516867f251aeb9263d63c694073f5c73f9833a5c66b30304b707f
zd7c7f3cbd7183ead899d75c88cb088c9c6fca48e4f8a48131d3ed0c7adc56d0ad567f75ee063fb
zf6e689c2901f5448b1d728809417558e5e4bfdd3be32f3413909485784ee23de84d15439511c01
zd9d1a33763f92437a4af48e9350facc9e5aeef328b0d4717facf873c533de10500c4d91f1ada31
zbe13854ef57e89ff8990920ca2c4775f904c575a722064fdfedbde245634acf329d000d61fb55a
zeab5a9da463583641f648c08be0843e22c939fc72d88a3974b46f0f911aca3ed95bd7f28286933
z7ec558d40dafabe1fc6db7314917f543c4892df7c2ba9b65ea2ee12bd2f2a2e151329ee281b397
z0606fe07a505f88f1e52eecee9ff41cd205559c959cfc71567976f0226702fef429c70696cf979
z021f7666065071cc25841702a618310206b7ae8f1490032822f382620f4aee9b4a94d800e518c5
z05171d63d54ebdc201ce96a16c9dc242fad30e9cde6e322da4a924e976516b3016df98e21966b6
z774cc0f11811dbb6af9676c2ce0344e02ebc15ed305ea39e6a7208c890deb8640b72dbf62fc6f8
zb56087effdd3638d6b568a17af044e622d1ce9396c7109eaf0423d1783eae747127bddc8944ecb
z5f4da4210e86b6751133013a354732db540e870d77fd9748b59a4a85433e342c041cea50811a2b
za07aa207e3cfcb804cdfdeadaacbd644a0234b9540908490f7edec6c3f6db1ab14961b07f1e2d9
z296d979b6140975667dc528852a50b63469b50165b4a1c56b38c80746df2fa13b2eface10ef588
z1950f92801bcec40b7f5b8986e77ac6ee3cc9f7a064248c2e57c9cebc2440a2d0e2d3ade395f2d
z75f0c97b5ebef41f972e7f3d05b4451419d40177f7de3899b66c285015c1a10a9896212c8c2075
zc6f4cf3a7dfc4f11afd2dd331c04dc99ded363f0a2327264853df7eed0c0f29f0a55edb715dbeb
z4d9925d267149508bbd187cd154c5170f0b5e6ea41372e2c20d1fd4c50db01439b504519cf0731
zf0405f4dd3554ed76f54dbfdc160af79e2c1d43cd3de01d1aefc5900a1987e434d302e3fcc233c
z62ba8c29d3614aa71c4914b8591fe946740b95f097cd085f036b10a20bd96360564abdf8f2487d
z748a7a0825654c01b02db10eb0eb5c07eb0393f483b7308b135f76fe8247804b91d524bc3e749a
z0cedd7e5ebb4e53e77bd60a224fcfa05e29c79546cd3d173784fbe36fea333bdc8f72534d7ea22
zb3415077efc93900895d28d0e67f8ebcf654920063585bd376233cd998baf4d6e5dc3e6e488ed8
z8dd9895f8a6f7d6b56b9c84e8bd389aa1f57a3103099a463e2d4f8b62a1454fc08f3c27446f2ae
z7e803a4f238f235d0953e931683de6900cbbed8ef66b641d9a220b7f24552f596bea41188b949f
zbef953f8b3b83439f485ee9327e6e5a5069b9583d3ed714e887ad19247e406d66b0f711b5e4978
z8e0732e577c38e4676cf57392636a1092799ba311708695bbf76b13a2f518058047845a14c4a6d
z34bb0dcb82b9faa85f32a4acf68e40330a0029609faaa09359dca0b5a92de05da20a0921e6447f
zbe138e9d2db67284bb0e678271c1dfc295b7fc98b09b2a95a725cc40eb05aa0a3a0eb619fb640a
z7eb755ae8cca3e8fbed4dc2ac48f5050b162edb7d3b4e14ff7f2bfe6b8799b52846cb98d7a0f8e
z3c33e0d654abdd2952c7311250a0c3c972100277a600e3c9af68a0d6895d74eafeb94f9e71f940
z5680ad4eede4565b8217f7a4859612d4374dac06383422722dedb677c43c4939bb0719e47dbac2
zeddd80de62298afceebcb98f47802c75f73205f63c039e83c515e84f2ccfbbe0270fabdfe90bda
z44afbd91b537a617aaa5508476af7b3cd8408862906f4cfaf02565f36773fd1c50a153794ed215
z446e2504a459ae99c79e7242fd909f949e0fd44ce8c10f69f37322a2e520174eefb009607aeb00
z9dc9e4c3cced46127fe905136dfa199fb6556e0970eefdadf8a48419f80751d8fae64c8ae163be
zce2c4fc33d69dfd9fed0a266973509dcb5fe578b62079b2189a5801ebe010fa2b493ce4b330e48
zdc6dddbcc4c62870a7e8edafac8511a0924ff93ebe1f30442386d0a4457f1b39ac97efdd838090
z62e99b6d9b10e67b02dc8b164752c5e3bdd16e511d4b2ad565a323d1cd451f6457748d94a7a968
z7e723d81b95c7b1970f44663efe83f57a28c516d0f8029c5553ab8156efb6ee6de9d266e11e2eb
z54f7f5d8694efe3ef1b891fce648188f5b7a6600a4db5cbade84c65c34ebf9c636e35062660e70
z3abd11c6d9cd3cf6b10435f4692e4030e33b31be3cbe7d38e2adecf1abac8680e6545c670db66e
z381651588654adb53fb55a4a29c8122cbece69a85fa4494f15dad23505919e9bfbfeca215dd8c6
zac2c079ee616ba4b7d5329f06e73c595f93229a475eb661dfba32ed72c28c048cd65591cf257e1
zde30f70a59480348450925ab9613da8ea77cd5786cbf67bce6a37364d5a57955a0dc531ce363a8
zd47890fc9eb9f24cab2dacd1dc2c138c014fd1a25b5e4c49396735b83d6d448e3f7635553426b1
zc6d2a4862ac88604a4357160a232afc1bb996c7a5be3e9b888c90df07777d37eed3ae6be6e74af
z417707b568d5c43fdb4876a25a27a639ae5f1ee126fa8e6a3c2ab2f10d9c4f0be0a1bf26652ced
z2b0e6d4524dc69a027b6d1f9efc2c707c10d60ff684ffcc753f6650e2bd2f15e24ad9512508e69
zd80bebaf09aa6cf92af410d9076da6a4dea355498775244538405c81b735f6bea2bc4067133a3d
zd664da1621a27b00c0b39c989773a21d7315306272c5cd95ed01407e7fe93e3b2de849f9fd45b5
z409aaf7e6642adefe76b5e61150a9d134c72ff26c8fc616710579eefd70c8b8ae592d7791ab187
z0d3af1ec88dd9537430765b76905596ee709617503526f59c456331c13c384f50e2c80e69487f8
z9b51aac8a9984850e347b669254f5e0703b9ee821264be7a56a41a05e692470dffdf21f9eec164
zc4adb187b4b568c3ba61db96107b77371a0c3769e0fd3e433e5b632fd9c894c0e761ed2d6a42b1
zdb70f9f20e48290aacf659106843252376ef5a12bffa2be26cc21e001687b07da2afd6ba1b9fb0
zb7c1c0fe1dc4e497dd2921858fab66c8348cd8eac35f3ce001c47ae3b1dc7d1784fd1d75a07ef5
zabe55a6fd59b05c34bd6b44a428aa5b0c3b8c8ba14f23794554307ac6169f7f8b37e19917b806f
z4cc5fa871b0376e8e52d0f37c5ef2b6054ecc3247cc1ae88793841aa272f0c864e84ae1a616629
z2f941679ea988ab8f95e98173e16412b66f3f485b7aac3587c834521837987d91a5222c455ee93
z3d43912212ad053f75f64fd62715b5ba4a6c66fd1cd589e1861f969dad91b0b594a2b7867a01b5
zcf7fccdc569101f3e23cc5fe4d5b151d794030f2da406bba19b690c1114cc930c10f6067a687b3
zf8cd3eaaf3b68229870fcbdc645278999fddfca1fc3a366c0ddbb38da2b00393dd706eb934abd0
z2e5ba2ca2f8d59c83c6c580475a994041a60f8d3253228530c5029bfbfb507353c2e306b05f49d
z6854af231164021ff9cf2bea751fe0c458979a9e33a53d34c063d9f61a420c47db969fa84c9a9b
zdf0e438172398970cf0fab450e2bef20f8cc66702c500a410824f7316ddc16426f1af06dc0d921
zefd17ac775eccfc54b3ffe8ac9daf76d67940886a52335089db0358f7fe49098dea5e377dc6816
z101852dfd3e52bd1781c7b8e05c20024415aabb5e9edb03a2e9e9790eefd7cbdfe9bdab57107fe
z9540ac11fd4b9304037e4973473fe7be6e524b94468231500da37cd99814a71ec5a8750f1784ab
z794447bd5e0d3cb405c5ea8131178b73b73ec45d7bb1100d516dc168a666434a273609cb7807fc
z1031553a1893c461543744b0a3bad9a3a8484e1cab8783a40bc59d2c713da4ce4e6f1e9d7d5d6f
z49dcb55bc691737254072939c170cb8a236cf2e62ed4603c128c142bd93942e039def24193bdc4
z778a87fe1c60ce36a65b634dd85f0fa3488b4a710c4f5ac4de9a7e1898d50949c86a702f67e296
zdbda21afda673e53c3b8bee3dc9b0f8627197a8ed235961d458d0c23ce31fd8f72d8656767a485
z59367227d3af91f6367d8ab40c5a8838e5c8b8988d19e9d7458a4c8e98880956f96bd8e2896ce1
z74b711456d73562064ccf8486111e8481f2d8b9baec293eb2d8505244f795d2a631b7cab81f11e
za8c5c15e9c4719614193456ce18a130f6cf531d64a225487adcdd625d52cd026380dd0a258ef84
zfa3db40199e50b76edf12e37c7bcde88f2ae59e16700944a035c532f28e53ef16f5416a51b54d2
z5ecb0f6ae85712c56fba028a749b0120c6f432dcf5d4660adc9f6838aea59d41deb455d29ba9ea
z4e21e2b3ca0fa0511fa36b55d5cdcb72427f7a83447ecb06340c05eb81083eeaa25188867a3334
z7e9ed7fb1f12098017021d964ce101dd57c1c164befe444cd725129dde65df8e20ef4a76853d4a
z2ebd590817f64ed9666360335f2ce47ba2635ab91275161e24cb0610315270190b53dd2df0e645
z67e041178b4d598dbf4738bad52cd167b03df8a4707cfdd1a3f63c285a7ab05f7fce1457e67143
z251c269af34f3570bb51f2f8f63dc43cb596ffa6dbb5b89fa145641343bb41a76d20f5902ecce9
zb4f2bb52d2fccc4e8d7387ec30340d8785d7b4cc521daa2f4967a8937601247d024b8dc33d3201
z25c48303052918c1587587fa178c8e72022643c05ae2018ab95f83f3a560ba2c8d054b2d98bde7
z09377cbb2c568bfd2d4cca449bb4702d8142b734b853586027623cc9e1f00461308dba54142c75
z972267149fcf81788d9bcf5ad7203e8116f91758d9c01d8c211b5fceffeae0fc143720d2d22a7c
z4db7083e73849c14acaa45e2f8826f36968e90c198a18d9809d884456dd8f5eeb2932cba003384
zf06ced9ade156b8deef231565f1f8cc6a85b24b180554456f84b48eff8087e8d7d066ff209e904
z906bfa735b122bf5d64a3c8b09f40d310d9b89c03ef218c9bc6b4fc9a7382e5806aaf6c0bc4be2
z174819f08822c29ad9bc1daca380c6ab9f86a1f038c2b53cdbd37160bad977fcfea0682b5eb1d1
z16c27182738228b70dc6f9c70c3aa2d462d529a2c42293313b39e993c221a443da17f09dae12db
zce11e56e2223ab36ac8240813d0f59e32a96aaf6396c24dfe36e5b9a0784a73ab4d099a0f4703a
z854a7bed7fc6af1d6a5cb74ef0a954ad2fc0cb2874602cf30330f832eaf5fd04f093693e0f497e
zf24a0e31b44a5d5dce844399bd52110a80a7d9f9554415cf176d4a3b774ed8a20220499d76f832
za8ecf896af757aa7c9421e70cec672e97a533b1279192d2cb02924348bc93b86fe7f45b084c3dc
zafc179a43e613efc1921ea906b40977dc1f3756cb82cae09d0e99cc4ebe2dc2a1e08997f017e58
z46633e0d792e989ba8d21309ef5a2d43510253eea6f61e2e69c21633b990e2471e23ec1ed991c4
zd689437d2cd73d622e166b12b88429b95cb307cf64cbed2b714d45d2b48fe542a032340ca64c30
zb12135553eb778ee2b202d4df0d27f94c6b7dd5e5c3bdbe4d954fc0bbe278c11d91544e53303f0
z2f07a46abd77de7ff842418ac0f5b30969266698f314f384ae9e25c62bc57dee38d40b87cf42c5
z2a8b7acb9187d2c0268ef88c146ddb4f68db29df778535a059c8e864b0613b29df110781ab3b1a
zd48a8c7e6f20ac9892a9612b834a7ab3a5d9528b3ae5d7f063f6c6c5f4a14acea59b25c3e2d7f1
zdbe3d845803706c2562267bba55be367051357bb5a89dddf58c7de334a33f2cec2d6ce512960b6
z626b890d76b9edd0cbf46c63b8714b49533aff651f0c45f360f7225dc52208edbcb22215784599
zafa6623dceeb7266257351f72807bc8efbea332b64c35292e09253dec2e703a72cf4b415c8a831
z883b563c02ccc15b15c84968040f1bba391c8904b8180991889b85a73877239e9a075f2f320121
zc7b037b08fd50f4404b7a3f2b18aa8f4199b2d78adea2aee23340ae4ddecc59c138f079c6e6852
z772309be81ee7d4f32109f2e27188e99fe427f759f8b52d52979e805ad17c3996d8320a9c7266a
z3c06443a0d84b1b7d6bf31d21a109a74059ba61459cea985ba040617d496c88694bca36b61ee19
z22a199c7f9c39e05e26bd831455acaae50960ff86302478047fbdacf57db4bdcf740aa352fcc8b
zb7eb3701b69eece6230a0b79aab131312b417cd23a9ea56839f471878247704fa038ba34c178da
za58977c33780505ba05286fe260e595918a6696014b1bdf4d10b3de6a59d0981430e5765fd6d14
zf5b2e05f1308a9ed4a24e7c0e35b118ca65b1648821f1e31ddc0713c573eb564a452e6c8bfc87d
z3119e38c39e3271a3bea2734aa56ca24422073f3ee95e50b79eea899318386182ada4c8c64e955
z8e55b13d08d32f6dc5f202c6f182b5880ba66736fa442d70ce468c9d27e1093da7c4a3fcb43d38
z2b9d6f135af464466c42f695c8a6d8fe4e5c2c69b63fc9b2dfe79b962eb07486e7e75b6b68e411
z166956debf3ab470b35dd7f7c7d80efdb648a1de2da887854ad5efc59f848deab16eac07973e0a
z16616f0574c5b91c9fec9375cff2ad9ede0049ec34f0062617aa86a237dbf27636a746d1a4936f
z582823300f9b707a50ee81766dc7d311ec23f409891e8896c94ae22befa766b43dae125e0a959c
z12c4d6b278db012283864edac7a6c8f29a7f128faee45a31c179203ea74fb7a75e9d9ba55b41e8
ze8bb6d633dbad9df854e751ed7b924da2b4c8dd8d814ebf641c9ca16d73b7dfe4911dadb022145
ze7ff7f453667389fa547d3cab2a9414e181b63478e79f6813069904ccc403e61151db7509ae832
z8d2255cc0e2028b9d63f2d0d8744b663bec1b343085ca98761606efe873db01d591566afa777f4
z1f97034b32d10c438c93a8aaeeed9427a9eb4b50b8985164655dffeeb23df1fa98c5396e31fe90
zad10b9030ae98872eb57e9847698f13be9689316e1bcf83b12aa3ead2be02868bdc5842ce91d1d
z723c25d55ddae067e8cee80bebc488a68b2b1a61455a2fdff3849e1782e571917c71d9e0498241
z7c522582be405c9a3a6f7fac75f5be622f9abebb41a17b986ce5b954d056449cc4b2853b8bea19
zb26a86aab3ca9686f1ae9d652384d18326ace0f60c4efe85e8691169d2aaa767701acd44861fcf
z8a01d87119e6c9de05845b58e322d3e0e9885880b5a36fba432e3114666480f9e03ddbb1b2ba7a
z6095925b648b735343151dda659ef2119820c06050bb4f16a368e4eb25f0e219305305b7be21dc
zfe80e036ecbca264d8bd7736dfd9ee5252089a5f0152a6dc60abf60836b65e483cd94485d7a24b
z8de98a30d79ff74c0527c913206b0584f9d2425959a171ff02cb8448e9d71984006050acfdb288
z9c917ab2812580552768c8d67b3cbc481a6217824d9efe263b5e32de6e23aac3e6dc61904a6463
z5415adcc4fcc93b5d9a2b8d56362773417b13439478690e3deb60b71391576e8dbbfb85b927e4d
zca6ecd8b26bc4fbd97b04f8821611dc79d957d7437ecb6f6cd6dec831f4912560352271b8e3ee2
zf4975c34a10ede3be0588d16f22c02aa4ac8b7a192d4c17e760c0aca6a7d5ab939bb5d3751394c
zb37564c9e9fdf16b64851d65fd0686dcba1c3ae043ed964df2d6ecd167c61ffee852b414281c2e
ze99490d6fa8a955ea0274ce50b02034491946e4260d46accad36c78661567fb54030b2d7386c49
z5bead732f2ec9c1284c1c4e0b26f292360ce688629e58b6a690228e6f5c7c2d6a156c4aa5733aa
zc6fdc3df3c85d738df4378934dfd6a38a9cf1941f493484648ca7972fd0e6c5c959b1b241f0ffd
zc90d7ac34179633cfff1f29e0dc22f8a030d52d6dc5d984273743c25d1b400cd2b8bbfb176b6f7
zf0586c7964867c437cd4548f06e649c8bde2a8b0429cd9cf173d094befd82842078ebc4b407672
z3165ad1ff380eb43e522321c97682721fe4a55634d1e41eb23e0d1846e548ccb3537930c2143e4
z7ae63ab28f5cee74bd02f7f95dba78dbc69efee2b04673034089830fbfb90459c875b0cc22c45f
zad2b2aacf1e7b5dc817cb393a1609c0c99d87f1430872649ec0429bf37b75a3e94db9b51391bb1
z162fa322a3d08bc822b60e86ff80aba39e636c9c776dcc4a6090c411ee52bdab1998458d88da6d
zccdc6a28e4c1ec01f8a5187d4c28755031b2c57532e8f67739d5884b41c8a547d50e14d4992229
zc2bfc62e7ce010cc87a44db8eb145b7bca69112501da645a1957ac6997f0572a6615964c9cf92a
zfbb899a6adf9afa77a723282e8a1cf7d7179382f2bfcb75a2bff2588a48ed54249bbf0d3816838
zb297233a8743092a3a90759f1cc01ed92301ef7ad27a6af8410930dafb5693855f8ac73a2a01df
zd72530b1a3110d86e20393cbade7731bcc9aceb48ab8f79aa25fb5d1038494d5d34dbf8bf80145
za287aed46b63e62f337d5db838409d2fd5ef6466487cc0614f16954735dd3257ab15a352e52c95
zcf06565fea22dcc54f22c4161b3e5781deaa1cd6de73784b1828b8098f9864f5ced771f208a2d7
zdd5583393d124c2dc718e42dd11873113467ca5e621a9a55cade583cfe654f5b42b54417fafe8d
z1fa711144508c449bf42fc514e765b1612d63cbfb8b7754c02d7f1497efead9c5d2e38ddfdafea
zde1ec67de0403152c3e455385db51b1942cce55b54826fba22e7641cc713c088de4faebf7431ec
za09436aefe5b36e84b5d8851f8545665eead03a557546b7c5b863dc925762dc2516138f9db7eb6
zede86e8e05dc96b8253fcaff64a654c64e700b2863aa15d9a9683a600453c4dd43fbd12e7e47c6
z7169af2e083a10aa058ffd733c8b382914a407687cdd5075efc94bb029a9ae1e9c80f2860a0341
ze0f4d66825f1ed703ab9357b175f83f8b54d47ec5223ed37094d21f4c784743859f91afaecb501
zdec453f3bee4feafaba4a467df7defdf2456b5ca5fec03d6a8b80a6dd72872160e54e9aa54f897
zdea3f38fca781cf40c2ca9c760b6d047950c653f76ec43a90b4ddbc140fa0793280b7846fc4ee0
z5c74c0097b99713546afdf9ded2773adc30d7f00a9340aea96761174be9db35f665255b3a6b3bf
z47a3fee464b5134a57756457846cb2cce43a8ba2489d304ea3aab0b93a2ad4218aff0442888820
zce114458ca17ee4e5df0649eb7e040b42de40c0bc2a4abd2ac484d9233533664185e0491b292ce
ze054b5e0845669acdc37e66249a6d25e6aeae99f329b336967910d7b5f548a849db0aa168ea12c
z691bcdcdd494ab10d2d046324545d3b0292309a20692b5b756f2fae52d874f6a728543e856c353
zeb15f674d771970df32f61a2e56e1a05868302c3468ab51287fe9ab6a922fec03dffaf11c29fd9
zd31cfd6abeaadcb2a216dbcdd9d179a4db958953c2f9e05eef160b1c6602b3a26f688da6fe01ac
zf8f6652f04dfc14b7da25cb7aeb26401b900d0867895dd06dc34b0658191f908cd3c69a14ba955
zd5729f4b0e9fc7cefe6cf4c76646409d2e8293b7110b0bce49bd47d8d177c9c6ed584b7e8e166b
z13ee108da058d17f0a392e1ea004a243ca7affd43f569d64a1113605bc67bdc89f7c2a2a5a587c
z389544a55ed38d927407171211d50822a03e726be54570b4e5c930ae08048048ee9a09fd52684b
zf2d90af9add149d5383d197a79aa9b880ad513d8dd49cde462a30eb9d8a1feed4dbada268115e6
z2c91f2ebc3d79a656d6dbc252b6ed990b95eee949f08aed0d570fd1f8709d9bd2ea8636eaab93a
zf3568651fcc311b0a7c40d8481e1949f50e85133a2e98e99314e18d72f873738de914d42367c6e
z359622f31936dee0a548b0ae537a679afc29cd5abe9e3af20916bf672179482392a23fd0e966d9
z5ea40701bd0a4d64212a91ec6cd76eff5c075488a082022232c5d1c2bab90bd9be2801f84584a1
za25b3a4aede56e283f069fa7e35c31f34ab5c005da6e3a0a5e17da83ca39b61542b8637818c7e4
zec03b248e820f5d0cce9e3c4f9086906a625448a313c88e2181deae665a4d9d0bb8af5c5fc9d2a
zca236c1ac8e0e756712c153ffeea503412ae908763cfac2d94f2159ab1b4cb7bc8de0d4c29e65d
zc42c566587f0558a86becd8c8f4da69e8e0e4e5ff73f81d12159eba77a06c60a497f5a97e5b7cc
z6e79531130b1c9eb5d81c72ff63ddd690c00de5cf931688fda44bab47eca2b4856efb80e095bde
z75907f7a5ff63d86e985fc1bfd63012e5954a88d581a273deeb9a864b496571a9f4daa0ebbe81e
ze505f7bd2cb84237bfb21afce44252c0880c342b701a46523f27faf969bc30fc8b3b9fd2013fe0
z31053c8c36eece09debf95599bccb2260d81e6a041ff70eda9a831223bf27bba8fe1df34351768
zdb8187fc5da8e8b8f02b81e6b8ea49917396dcc57667bd8436ada7fb308ae355b07454633af97e
z276b97edd83de25b6b25375989977212a350ec0b218674ad5f46f167a8f9b6b8e46bd57e30cd69
zfaafc6a3a8a855dda146db492bec1122ad52b45ba67a1772977d0d84c1065dd3bed4c7ec383d66
z1f7cc8d25278ba573a7b5feaeabb05d4108c350279bdbebae3a9cff9694ee44e0bd7219fabae03
z44386a0b9377538c9a1c2fafe05bd01f9edd4d050f17b50befa89d4b67244c6b44445fb806faa7
z60c2de0262db0d758500eb8b9350d3d2030750921ed7da2313335bdf66a625746d75854f0493b8
zd4aa258affddcab71bfca079633e8b5144bfb0422f729cd17055317edee8084c21491b8ec9304d
z16f117a8c2a2ea86ccb711f87b5e100f530317c83b7c32e902aefc5c270312e636de280e28890e
z4329e6d9453681a7a0c2ea4f001e598dc789f4f0b07153276ef3bd72a40fb99ecdcc9891ded671
zc271d57f690402d3171a2fb4c36e88d84d68d994e4db7266d15aadcea3a74434da46f5a4a4e734
z070a9ac499508c8d6891d7da20a7fa53d74a3f1d1295d817c095224aae15e3908917cdf1aabdf0
z8292ca085abc12700cece2cd01af5ab986c5479db6c0544a4105443f99a865d1449b3a198be596
z8b72122dba388e2063727cab653bf5f5351feca6ca033fd14df009937b69a6479addf81c4daf54
z46d69b387dd4c249c053c038d7c3db2cdd48fcbc0122dd052361848836801a83ff942368ecbcec
ze71b1cac61cc5a31c293cd8630ff7ed9f6c78aec9368d04e476ecde091b2fa3da8ea587dbbddec
z7191fb3422294da7a81adf5d2c4e1cef8f7de4121fe95e7714467643c5923e680fcabc57060ec1
zf8c56425310191732ad12be3cd2ed8f291494497fe476e5087952e541bdd3899c5fe0a9fedcaaa
zcaf4061b3bd5a97f0adbd93c4274ac14055d88bf7ddf3c8e6718998c5fcf88115975c0eaab42d6
zb77718500f2dfefe1b2c309b9de557f94029ab37a7cf7ad8c6fdb86d65e2f75d49307401d5a3bd
z66481b8f135101ed533e0668cf36a316a0745f912342e16a33abbdba9bfd9fec0c53112bac3d78
z0a78ce9c5e31efbce245fe417b0c68a2720f916dd5b6ff3f20040e77205f1a00206ddfa7bad481
zd4bd4943b12a3a66e7872c113d9d2435452a80d26b88970101147836585172e3f37c055370937e
z24629ec1465b739a3e9e99164f74a689cdc434a6705a1b2df57a43abcd63b2a0caa3e9056890bb
z82dee37af3a11cc73d1be7e3d6bd05363a3024a0b2efc91228d268aab034e37abcb6103c586d28
z4a0066ff6b13cab0b054b455a102351fba2883f5c8344600a263df757f05f8588b6d843425e198
z3c65f714f079da191d74eede81b7fa760bffdf9297accff01b768d7ed288637b3b39331b78c36b
z89f591dfd957a662e4af11009e12fa46958575e6d7d6f2405eaa2e9b14677c1d482965a271a844
z81b360a10713d5134f0b4869ad6d83c085fd17c493ffe031a33089872a1bc9c714b475f0cfb5bb
zd9d522dcb3b17a4ff2307cdd4b357dbfc8c98893dd95587bd66ce2a76f0548192db843b94b2c15
zbac21dfd0193f1dc9a2e73265da2fa87cb9c487e6fbe368fd7930d96d7b679a868586d981a6738
z813ce3978e37285be67baac5868d49ff31b84338338a99ed4b5dd9531e8a2af5775de1e2802cd8
z4ab7e3f3e2f8ea91d2788a5815b5c2951a574237918a4e984aa7658366af60768ca69d478a2288
z2e985a3babef8f7dcb19ad186f023ba5a0f0926523364a4589824f4355b4f97b00ddcd9ceb14e3
zc06bc812c0e13467d06d068738a2f2eb06bdcb5a127947eed808beac960dcd7a5c9ebde08d4b07
z319147486662d33374b90d38362116f9dd2842d642e6e7d1f0e59975934690cc5a80e5171f80e4
z00d8a93cdd5bfe107fed58ffb7b0e9ea630447235da9a37ba1d693b702180bee88867de3079b1d
z0d72e37e7988a6ff4592a6ce3e638b6a82c436d29e4216dd1c4cb70bafca705718a36b667758ad
z5062e2f2c24552d8da25b5df4de0de9d661e8687e8a815ba7024680d858febaf9155ded3d47357
z0bd3a0d53405db973c8dba49ec997f5326bda2a603ab88db4cad530ef16baf3ab077ba521355eb
z048a814374cb010105e188407c3e5fa847820eb082971e6bb85915ff46b9ad80c2df88affe0050
zffcaa5ef066c79cd492d1b193eeaf356fd8431e6975f012aa4ee4025ac808598afbfcce6b3d7f2
z5abad95edfb8306a33a5f38c4ce68bc3e33deb0718cb690fce81fc69f8d06af7e2559d48d25e3b
z0abd2041886c9ed547f11cca2b7984cab712cda3c4fc839393ee4eec8091a5f78943d4f30b1edd
z53d508bc26397be922082cbe7a94275a07208b217e846441d9766e09cc0f60f1a43abba02e1a85
z48676cb4b11321332d682344ecb09b0245ba8d09fa5233b2befb017aa9597a2a381bc678f1fded
z95dac469123a5fb24970e63d39200a0353dbc825891826cae54372a2162b1558acf989386d3695
z9f4ab80fd36a6a1c5f773271d4cc753f2eb9993687cbdb445a916ca7809ae3ed01bcba99fd2ab5
zb3b9ad4f10f4b4012977854a0237345a69873db1b5f39a652cd6df2322d36eede4edc1020bc9e1
zd99ed40bf156bba57124de39baad44998ab570ea8bb57aa97130eaaa4d5fcb43b6aca41fc056ac
zd688a4ad90c6f423dfa086a425397e6b779db68b8b14964fa5d02de5cdacba390a0556c4505c14
z560c00de0f8a4eedbdcde9bdd94fd90fb241a058d5ab26569fea899c7552090bbc58fdc1f7725b
z04edb1610841020d3ec50ac0d8a93c3cba3b2098ac7b972076c2e45d9ff4b84f5d26e55c742cb4
zbb9f476fab0e5490df4a68b3ebbd4192cf5f75eb78927516896b0c65301e5959bda5179afc73d9
z2d0378abb5c02ac40d24e5d67610b40c2a392dca5b29be057a9207e743625bcf632705abcc1c8d
z54ddf2a91a5ab59dddccffdb31a75e89c0fe8b06c08344a513e82c2e397f42b0ecb283836af04e
z37ba2af3801d27619e3fba34abae9fa8042aaa62eff539b3cecd48fda7680c228ba88732e82fbc
z73adc78aa76200067bff8bbc04a778d91c6ce41bdb6f01cb1b01752d36a6ef44a9801637a900da
z0d34a29a2b35c8a44bae4fef7a14a1fda0a43138601d16b95519e45cd48e2a484281b72f02849c
zd262304bf2cc83d24f247c9497ad227271174d078f61416c2539be066608d945d71122f9906178
z7c40d9e4d76dbd784ec9f9810f3e8cdbb4f769867ffbd29f6593ad4374801a06d6bfa06f57bc58
zcdfc83dc4c6076f9a41be4900ba5e3ac367579cb76931a94666797e8add3bd97dde0ff2b460ebd
z2d6272cbdbfb53a70a521cfec9db126ebcdd4b30ebb15d2de526928c60e8c5b9f9efd48a32c44f
za9ae58dbb820df23b4309f63b3d93afca253253ca7627adb6e52c0eba3bbe9717cfd505b5f1401
z3c0cbee1554248cb5d285de862e0c397e23f55cdc12ae655cf5e08667ee4d8a90109419bc15cf8
z1e6d4353c0f2a3a30944e5ab5dc8c057afb10871493025d708fc9b50fe653f1951994c8673a868
zd6e36de832a183db621543f29a9abc712d67d8de179d6e16753c315eb07254151e2b54c59ad509
z8ed9a25dde780e16f12990ecd33ac690a12937d78348a76ecbf7fe42fb4dd30106d7fb3dd20fcd
z923080724b0d89777c5fd7ca799d88cec5a7c371725996882022aa12ac247a3ce66638f0621d35
z0445faba7f3b0414137a88dea668f73ca5a8d2ca891f1730193a05634245a28cc3ac014ef662cd
zd5609dcb086cb0558d8902060edc7269bb76e4917c63f5576e43d3854c2374b37026b4475d25d2
z3d65f9f5b4d4b0913da36e2bac534858045973a22b4c665b8aeb030ce08418ec549a4aa79d459e
zbd114ff9da6deed9b8d5c4da8d49b5d442e8b351a96ab5e79fa682c22088ee35f1c02c0c3a9361
ze1e1c837e3103dab8d5e5c8be5daf16d62eab71a99d6a3ca96d7f2c1c25e65dff732501ffc31af
zfd6bd3fc6ead8c51829723bcec1eef956e472daab39d72efb97999e11ad039e0d67048957104aa
z32116e4bbe4e6605e8ff52f8f1c8db1d4d682dd11a02d25cc1e60694e1c964b1aee3f5b45b2202
z890cddfa59d13cfaede19667b5c98f4646e5390dec11d4b3da16d1fdb9f5eb4cdbd88d0acfcace
zd5d181ebe8552e08bd71166f2ec1befb1c37cc733207a71a840c9475d53a08c561a28b7278cebd
zb78fd2c7ebfc2847a924a7ddc9b2b98f846c309046fb67d91b69bb8104c306ebe2e7ea3794ed7d
z071961da0185b53bb78390f898fe265db7ca0268e6443402d6e3836c8bc15ab549105f1813e4cd
z9a8f4faec647e3c34a400e6e893205929edf805141f5d5086e6a07b2a20600fb6ab10edf3b1569
z9bffb2f9709533f296f33b25887d3ff41cff68807f4dc890b9f9cdba463172a76009e57acbad64
z20b092060ae66dced8fc6c5fdc05d9dd44855fecacde057b921e14b0cbb59a1cbd462066fe9f0a
zeb8ec58082f7cf8519355e6e0e6a659217a014b9f87f3ee3d183281915ebc03cd4f648f0534de3
z3592f18f76adca62e0c127cfe845ea1babbc95c191632240c1ba98e7dc40be42107b226117a095
zbc21ebe08335548e8b6995451afd26729423d60c51dcbf351e6f34c61e48a72a2681e3fb08454d
zf965ee080d6b221a49e8cd49762148ab47320fe82c8142b2d76db330e6efdafc7d0b6cd6d3438a
zdb23b6ba5b6bfdc979c621ba0d69e3071e7256c7e0d348be918211f511e5ecd1d3e3cb5d02ea50
zf87eae5c7abb5ce0b76056ec231b493eef3b6cbaec6b4894d3a00164083e8adefd201ba8bcfcc7
z2bbfb86e3447a0132de57696049c512afdd7981d07adb762a57de91e08f4c21de84cb282e72917
zaf1282d621b291d097ee006eb9ade1b9bcf6ee1b6b979dfc9e3d8add3c617e249530f617165cc3
z4d0341e3ab2ef20c78327a79621e50055c402db59a145421b5e0ac29778c9fcd2b4251945a1e28
zc8d2ba97d397943197675cff2009e5df9a17f4b538ea91181598b410354152cbf280190eb3ee25
z4d1802710a3efaf732a91081823ece8ebeea2cc8c3cb3f71e9fd6c5d41694e15cce63aa091d9e7
z4a8653a3c43ef8a8c5f331dda01a591494d96950ef838a881080edca99aabb8e9a9e669f589014
z7c4f9b0c70a1831a10d3f579966ec13fade9741808902d34862d4ef336ec027cce17793957edc8
z9626acb36674afbe11d20dbdddda171b83c685f8dcde5a242f6b858334db140e7c651579040a06
zbf4a854fc51971d99528f7b45275a89648279e4e29a0f56519827f0382a364a77fa68ecac08595
zb1f7d32dd2f1d36dcee33d89bb09be76790d42ebe21f4a0f0c9d62a999af34b881bf972a73a0d4
z4b9524019d7251e0f481dde9e0aa6b23e52b784dbc36f8400003f2f730ab1a732745332c1f2336
ze99d14e6d6fa3189ba02c6d738b830d6b7b5015847f77a03514aae6c4a366408fbcdc1bf734cfb
ze3261f00a1b48b88825175b848e98968dcd49fdb5e35f78eabb840bd89a7393ce8e5d56c592fb4
z8c4df0eea69498596a54085e72a4a3c3c6b4e22b995358a568619fdaff436f7eee26599c6e200a
zcb6b3d9f026ac4874c11aa6ec39dee51ee127f9935048468d360538294087263c441cf687f3703
zbd6bb08e131cb1fa16a4ad2e86a2da5ed02b85e1b5cd4e998922390a0ec8e486e48e9193f01e68
z4b7e44e732b770beb9bd72e5c002651ae8eb58d1fdb740f25f602c1d554554b52fa537dcd20a02
z46b0708193e9a6015f54a41a8536b70b96b45c14851f4d0fb0e70ee00436060411a803f151ca2b
z3fdca519fa293e39c8222fbf4f1acda53fee98791ad8c757b36c0fa1d02c55b46d065bce0a21d1
zb680f31d725e1a68e19c58b7d95036f7db8cf94197c969ba80105f2b7b256bfa5dc03c53de7121
z6ed8c024501a091335da5a543206be1105d488385a23209191b061e5543c1006b9776a30749dd3
z022fcb85a67607ab50ccad60dbbefc8cf2dc7add0b65bab50f13b95325f6aba63e4a5581ea4977
z912c62f63a8e580fff2c519cf8bc0486aa1726812b1abc16af06b4246fecdaa45d1e7f9edbca0b
z46f9dba2555b326f3e78064f4edc48d6629d2bd712018bc5ba5bb42bfe37e94154f79b5c5ec4d0
z46ddde8ef0db1876b7ad8839013223e8f2fa4f1203ed4ea5cb054fcadb930a3c7b4be48ad743c0
zcc71b1f299bae56437d12900db20534b25b10a2826de0d9a61e48a9e8fb01ec033dcba9c43321b
zb66e2f206438655bd4cd12476ef14dd80c8010c7ec27711292d31c3dc01a134f1a9db2ded117f2
z5c873da3d6504dc815c9bdf5f80c59dade47dec4e349b46b9ade365a40e59422d71a03ad6e5daa
zf0f9a82f8754682b8886da0459a1f870565525301a555e868fd274b46aa9555f3ad6ee504c97a4
z123bdccb03bb2d3cd7329a98a57276e258616288bbc4c043b93b3a44b065e1973bade3282df535
z2bc1bebcf4ccd8a03cd26e2808f6425ec6342d221f9e5e87221b6f11bd9b283ba4e9540c7b3d94
zd898815264808912b77fa580268daae813b22cca43c35064a09bfed96eefdd9e9f868f41730310
z3e4a90591b534c89de8ea0f0ccf6f68dfc141039ec4a7305665e12204bd47b2295ee2e471ed7a8
z2819952dc5230951d8f5991435901375f2dc7a702352f6b56fe5856b50330a665f79f89a28a507
z0153a25984c2ca725e6cc2ec1b932c19205222a67b09bb5bb917211fb61cb8c0c73c8a2075cb71
z028f39d136f22dba528377bc0a1a6532d61c9aaecbd58e4f5fa1dcf765214540bf950fa3ddf4f0
z68b3582a44f04899796cd52c57a396cd97000e261a633191e5f99a8e899c0b7d318950d5a71465
z719ac44973d2e2576b2e074dee35a357dc2a42c36b841dcdee89da674e3e59372abaf23e3665ea
z64b8ee8b2a02d87bdc8de9b7249688e3fc41c565abc80dc774c34a2518ad2da43cb2ca47d22ea1
zd58317e0d5e1666e4b8dbaad99045665f53cb37d2551eeff9b7303627537b91697edc1e3ac6dda
z99fb47188a240a81709e0d8fb38de7dccfa9dd84511fc0012a0f54c8780af520b6dc9e8c7cb844
ze67e60867f69389f271c30e9263eaa98f3efc42b0466f0677519d6f9b6dfc0cd4ef7cf6a5703bf
z9b124a4cb18c2a9346d33924d8b38830bdc9fa1d13ae7fb9bdc87c629bd8d675d5d163ab57aa56
z2f701666d4195c0321ae03246ed9f6cbd1495f35991b6b052d605662e4128c28dc52148c8f38a4
z8cdb7b7223d9ec7869b8a992a364f87f88aa74f451ed39c58ffe182c731402876de67de8e1a31c
zfb5e32696ca7bce54b0d3c4fb7274ce2b84fee31d0e6087ee2071fd0a71b172b9713d3da8efcc7
z72500df1cc3cd6b055f3a625fc8906ad1ff0a9f203d19efa4b80d1a66b792c5a6d68c91c7cad3f
ze52c55f390a61af95cc869d694f9594ce95dd1d6e579789c59ed11a580cf611539c502faa8a36e
z6bce110bff6f149db53a9837dd4792d26c5e7142c08e42488883d8f7537befdb89cb87fe9d305b
zc56855e48b697531f56bd398ab00d148575a36ffebb99b614afa120350d4d55f95d2e3ecb8b7a9
zc21d393bb8e644870d43a603d8d8341ff7cc98bea4d0c4402ca3e527c62d65b80f47b673d77e90
z191f80312baca0196cd258fed9434aa259699736fa679741b534c48a1d80a19f14c7f8b2b74577
za62f38ae587f268fb76ba489fbd7c8587f3daa3e0625a7640c4fc43c5ae56b0da396ca6a7b4900
zcb0a7248507cdc75b0d98c57ab3aca068d336954526f93017a476f147373331671e70b5c943753
z93f7a0cfa82f0b827bbeba2f01197566256d441e0985e317c03a3a9ea347d4529f6a954f740dda
z71722ef7aa47301fdb6811f66c69850e2d320a0b485f3860cb76ea576b7749d9b268106b188d90
zf658702c030ac349ecb89233485c8269d488aadf2ff2b344fc997d85f8ce9137341d643a35607e
z345604ff887e94481e5ac7e2feb6d0ce53e439b1f8d01aa556003321af603e921b2226ed776274
za65afb36312ff98c81b1eb48c938faf7f0bf8663b4aa9da7898f3b58a9db668c6418ee15836cc4
z4dfd7f5e57a6b1e58d02314b2595b867889a43e068c39b1777c8679bcf5d649cae88f93f6e20fd
zb690db95b3f807c2bb603e52d8e3096156d22345a147158cbe8da67f675a3ca6bee54d479ad0b4
z92ebf130804738f550302531054a85e6a03cd1ff85820084483c15e8b3b4c2526ab5f8271b97ab
z27fb9ae7f3a55b21d4eeeb97fd1108b5dc057046c5013932ec6248da3b9a635e192703a15c6ff8
zb9bf827241e3b292771e05c3530a168076a10a82a230be8b22426860674add274ae2f0e08f9b8b
z8522599c316908d1bd73abcbc958467cf7b1bf8b52366deaa9f0068bdb2cb43c2d105a5521b763
z13df27b9e8ef9d55efa77bb609a7a09f4000beeb82bed8ec000cbea112fc3c4ebbdccdae23f039
z41c6432466794ee98d2d2a0b7aeee99188d5253b06a3654f850b4579a309313c231ac415c59149
z62dab53a0edd5316341bd2805a7914dd147c20ac3f70378047e817130a463bb97100599f4b3a34
z1e4e8d85733511d9e60774358669c5923d3d0bed3a29fbc49f18bb748c1c71c268b6f9a1da9970
z8bf2ae4e4e24c8fc1619ab6d08e8151130aad4a1ba06ad886fa8aea3345edf6daf1af135aec3d0
z901f536b9d1bee256320812a4eafb000ba7c05d82b50d55f8225ad353ff71c6be7c94344322761
z314673c02ac8a9a2958263c65feb91f9e52e14cb923ec4fea7bc3750ff17251fbb69e68217111d
z6828bd558f777de1cccf6f99eb804a7178c2b2d049b5a1aa6d869ce15908d9f808ac6772e22438
z4d060e44bcebf98f46d383b665ea8c6ca159fc74d3e3ddd5aa4a125a276088103911032142f424
z73d5ac43866eada4de44ee59f2f5dde1200453387acbc767b03bb919a3397a1fe7409fe7f5b164
z63e9c9b9c3b16987be9a7de4d05017a4b5f07bab88a74b120ff7ce282bbde9c8bdb679cb54d5c2
za30b3e191dad410dc0fafec33f60204667c5594aed608f115c7b8cdfc796855f2a10a0d5ea71cb
ze6d6eb08eee5dadd326714557515e292dd12e4ead7bd1090227b4b09ea9097b0949a8beb3f142a
za48104d811ecc09ca464ae7b8c5f88e306806e734c8460d88e9993116a7a210a3c8023b2e82348
z19026fd49d36d0fd4257276d4551747d3e28f3066fcf1e08589166b972eb059ae55a80d3de2c9f
z1e70de178212eda5c8c7da9668a247f43c6534eca33f54da1420453016b1744f5b26ff8a17113d
z55fae9199aeb8581933ef8936203db46cc78773e05c689a3a0fcda8d30b0fc20bef9af7f127aa5
zcd460978b35f31228aaf2aa6ef7c36ee5deabb0d4e1407fc5934247e2326642977317169798696
zf7b08013646d70476be9880c54dd5ace82fbc4c48ff7d3188cb99dd7d2f1ed42a310215c20f857
zc83077d5262a04b98b83a54a0461a84d5bcbaac62efc9b1c0880cbd1308d43e47e7a1111441156
zdd04e499fddf1be87b653746d7d510f2f891932dfe92566708485a0293094214f7ff71735d5933
z2a971d544ad5577d21f9052070298d889caede6a78fe3511f17b8d71b2d3ffa5662025edc6ddf1
zb155ca68e611a5404dea42d581d38e3849488b3e701ff901fb59d34a981e9dde708565264e54e7
z0f7863b6f8c44b6cde7b53d21e149bd883d9fc2b19e77305027ad937e86d02dedca3baa8c08ee3
z38fa2743d9b7724c2d822f7832125458c237e8eb6b69eecceeead92f6bf37b9144180d73580e5b
zce66fe940d6ceebb46235de86704c7cc0a60bd0857e2191430e8d31ad27f0cd464f7c966048a33
zddcf4dfd6dfbddcb0d033182ec7af7b068f850e4a8504cdd6ae72f9645ffa0e98bcfeefa3534c5
z3a099eded41cb1c4e72d849fa7f49ef9bfdcd0ba5bc84fa75e10ffad0a22d1e8e5f75d5063a25a
zd3e21113edfc0aaf7cbebcacc3223ee0d3d73808c1539156f65780a1afb9aa308895c0a178a9bc
zd9f26fdd06921b625e1d2f54e9bd51a03f0bd34ef89d61f1037276ff24350474f88c76108911fd
zba5a71191b24450317dd5c70567db8d4b51e11b3fb47d9cab7f160adee1e140fca4b71d80c5f28
z894cb6be147920265df1d0278355833cf5dcb1cbe8993b2b8a6a6402da06f0b2178d9c12a23564
za5c548d49f5f383a8a2e3cd84f4bb9f2dab46ae51a4f16c591054598b8bf90b287818563ae7d04
z51f5f44d51417931a4dde7786537f2ae88b92f3d2d22fc17aa20127bd3e825501d1af0d9f159dc
zb2e55ff9cb86def35b6659e760a497427e9b26d850e45d9f2550dd2f581985c71e1c25935df774
z3baa796b1319e49bbafbd7f75bbeb6168e91b20b8c4314f59bc39d967558fec85f33a4bf7e0edc
z6dd09a44b7d724ef756589ff197165989251abc1b1970cf13b6b274ca642027d0236ec332e255c
zbe038f349d32151e9d4afb866bd08ef11b17bc42e44b984752fc2e67f1a63004e8e987d68ddd64
z437d1bef3e261c5ad826aee5d9881414e23d39ee41b184740210e2571e42a392fabd70ef596559
z29a2824cbf0630457e67d6d8ee92ff3082e85747d322ebf4d1fbb531daee23ae2102e06be79031
z66199dc326cd55d6d124888029f6327d9c711c761e5a71f866d0562d2fdb9368e36edba2dc9920
zbefda10eb8be2c4cd77bacffa648e330c07d071c337a20dbfa46a773a4f8eeaab1529e523ad36a
z20c6b7d2c8246399cb80ab60f7e5d9c862c1bec24e044964e8b179e1c0cc059ac4106cf3256242
zbece8ee0ff0a3f2a63c4a0554b16e50a627c9b70975f03a8b285f9427c3d7f0d290f61f0f44b8e
zb80d1316d20f47d210b4b137bc0f6451a3e382944a5722d4ed19bd1566f4bf3559bb5bbb73ca23
zc4e6ea5399cd30900996c4ce8c6b6c3b912d9b51261ae23eb68dbd3f67e42d907f2572cd809fd6
z166d0dc0864853fd637d20ecbb5a0122d830493b28a733e7c0c88b463883ee3f5e0eeb1bb3b3a1
z47a8a155cc3a0a2f1991d280579f292e6d00e7538b85232add786b624d4f3c18c82935f1b2ff30
z94ec00bc9b67f1ad7b5cb42bc5009ce38c8f00ffda2ea45524368757da397750c6709dc33b6d42
zd8001d17897203b2a4da86785db19af436566df34c9d6806577ede472aa99ce9c1f7b276c5c9c3
z4ae7e6f073a827acae0d9e58278f8483204c1eef892e45e09dcfb2581b5ed7991b25d23fcd4de2
z16978c02e6f7cd74d9e8d8cebfe8958269131ea1ad2d9246cfcbecacad1f57bd46db32ff98196d
za34c7297644e6f952ffe6a5e5bdcc86986ec054df8753072b51d2f0c0c889ecd0aa901731408ea
z76ce44b0b10f8d4282e1689386f8bba46329fd3bc5a969a0cb1714f304fc633b8f5589d1d8fc89
z2fa1a31220a1ed1a69b27f3bb1ba1eb816f37d8082c76f7591de2111afefbb273bbbd9d3cfc149
z18e87266ea5f28aa8d766e4601b796356f606da1b46af1c3b9ab3eeac97de773890c79a9e6a275
zb180680e58f0274d70ccca2f338826dfaca236800ec20bbcaa5070bfdb828db88abec3e745da33
z476993e2da791be5fdf92b8455b883608db5a709039c39c8519b3b25c1f25411910ee44b24902b
zd252857f930fcf28cee7bdb13320522879e4d5d96fe26042e999e46e975d15a048771e9523067c
z851d7f65a39c75a1b319ff76aecc0b9308aa5ce66229529fc2589936acfa40db1cea1e7d11360c
zbb466a2a1b5fb0ec827b1e108407d8d552081da212ce11a2d7ddcf23411ed3b8fd4e3bfc3dcb49
zd7e147fb8524d2f9769d16a1974f89487297d04527551eb78e24331d96ff5ac994b39902045bc7
z213fa4d666227ea351be38a08aa71e9c662f34fd084295186ff5076ec8961ad3dfe06ffa199fd2
ze4ad64e2987e5d3229f2105e2f2c455932e0c40d4bd4c4a78a3066d16a54ed5904718ddd7468c9
zd762e70d0bbbdd5cc9725342d8f32d137d9b5ea049a15fc01a843ce958a46127ee5f3186008e3e
zaaec91b40218cc79f615f8160f321ae14408f842557fbfc23d39031699f7ad664bfc3330b3f71b
z71f90584d16bd6206b10d8a2b67b961b03384e4d44cd89b317ecd1568620c8d84de812504fda1d
zb494f64bdc5f6fed1f989c642e643d7670bada7ef9cec723b7f7249e081cf6bfe58a6c4f603222
zc121acefb18160f6fa26b98fe49ec07e2dd9ed74ec215791620d1986b84ad1f07dff3b036550e9
z4cb7e4a14dc83faf63f2b7b6887f439518d1c01309b044ddbc253b289836209d41bc86f4179583
zfe10d97497012e32b98ef53d1b495bd8e37a28fadd409032e6bd663a43d57c93135e236a843a3f
z49b727cbab2581e1a9006a656023cfd703228e85fa3d27d944f49063b84bac7be908d5dbfb7834
za8e4519128d3541363789287a3afab9b2fc8fd1743915d316af25d622d9c86c4e98b6984d23787
z56de9cfd21dd9f45a90dfc977f670463cd8ff47d3c426f74f91b54036e563597085b4892edf74e
zffbdaaf31cfdb4d168a5a9f467c3a1a0eec64be8676b67124671aef1e9affbc7d9261dc6561a39
ze187dcb01c942bee5b9ebda02b65067b6204c95ed90e85b621d6520612a47220664d29b6bcf979
z10f722a0d9466618dd12cdfdd6cf665d88d6f81997651343c4fda80af2e0a6b33c5339ee2a3cb1
zdb9d0cf494493631e3e08e2f75ee34459b970fde43f849dcf960d3569406a9538cab9a322adefe
zb15ee698d8f404196f12e2cbab104da398609c134bf2080ce027af893b0a5922881a64a750c2df
z3375364a214b75db9521c6c2d1cd0038099e012d214223920be384bb1a5bb364afdd438ede839c
z92e76b2f74789524d41661c385d4fe752e77087050f9acabbb04a0463d5965c11c85ef1a3dd91e
z5093ad03948df97d82db1d1a723dd2c5602a6345aba416c97db02783f5d4f08e2551b4f043a649
z3f90b4e41a0db35924b09bb5824de60cafdb600e2c95a350986301618aa74189215200000de9be
z5e093e191c05557ab81d3b1a1b91db854b422286a69e5bb441925c8cbc44f2ef0942d02ec26749
zd37ae70c58302112a1ba575c5901adba279a308b3d42d734c6664357574cdce8c4eaba2259adaf
zfaf773891080fe35aa517345b16006e7772cd0f36c8acb3187ec8f1561c85932ce5fbf3c31bd18
z49a89bf4d0a17786ab1dbfedc75d175d369a3f011c60580d9631f16550aecdc0b288e79c651296
z40450ac29e94048cc78b13f999b0bc5d8fc04ca1c210a54499b4aa5e3c07dbd433a6e2024f1138
z6174a59b2e91f18f3fffaf876f30476302f93c3e72646d9042eb93fb78997773ba52c26ba6b20a
z45f316a157286041297f7baafdda6900e5900f35536da40568319b3eeb19cab207066e50b703df
z4efade5a0735b760e00f7360ee164e1aabd2ed47033041f62d1a2a49417a047f82b6c8ced37b78
zcb0a0374e77b8005074b67e88c05fba7a7e59f65a3add785ee7b761eb8f368d734a2ee6b3fdca5
z017dcd02da7166bc8c701b81db7261e8cafa25684436b7157e7f770d6536f1ec85879b3412bf5d
z1c6a233bd1567e73f80c21c99d657ce77ca7819b465dcd814471ec4ec7feebfcfcb761a9094a7d
z42ce1db50e16afdca4aea656f12194de6bbaf85dc8756876ccf5b80d8d847147916a3cbdea0994
z02c5ba140acc11e82ea396eaa127d447d28737bcdb5848c382ab6db53844487dcccecc316aba26
zc4ace50709e4a201259eaaa7096d03b7d072f8ed3ecd4f47d17b7cc564d8813d34bef27a6f4670
z39d84004e413d0712e712223f1b86ff608a4374e696ebeb7053200ec80feb9ffdc849489f2f4f1
z222fd9cd98db03e248fa2a239000439c85d71843c3bc5a8a1aedff8aa02aed0da66f1affdaec0b
z3cea216b023abf73e2d6660802e2df162b081ae5cc90e50c8e36a63d34fcbeea8cced0c4f7ab88
z3d2d1c5a9ccbd2cbfa1939cb7e5d8a1871c950fbe77d4a09cd28933da6f7477a1bb19408b94d23
z23dd9bbbe3114b4c568e1d30fbe2ccf392f9e8761252b7ca8f3011c043debf038be804097d9c73
z85e64d6df4fad070b95ae5952e9f979750ce116acef4f414efe3b0a531439ec28065d3348f50c9
z75a4e2df07530e3add425e07ba02e9a75af095fe81640678e018f7938b2c0da930b6d594d714d5
z34d4fb7cc34faa7bd61d24cdb88de23bea9d5ec63d7539c273bee40ddcc8f2cd2b2c0f22221c1e
z0ecc593a4661092ee67cb10a1616dffc2cb6d9f5daca8c74791a78ae29e58fd5c982e7ed1e32f4
z19b3bded45a64f1deca6558fe096b2045e9975fb399586c51785b236f28a12706db2f9f9925087
z928a7e9d24b6c6996801658d72047317713d5ec5aa1fc3ee8c3e1c80b68d1e5f668786b29405fe
zee4873d68f7d19aa451c4104cb4c31ecf67620a088d83d6f15e2b1a43763dda3fdaec9fdf0c054
z4abe8ab18cd973460642f2c5b07516a3ce6205d16641e5645c1a1590c20377dc518c36f2ab7712
z9d3bf1f14786868de58e2e234f6da844a88a31ac2c673111a0ea7cb52b5703f025adc501a9df83
z6b1aa5c44c5b485d92e93cb18257f3c6e33b337998b2b2ae61125a8eae137eb4d178604d200e8c
zf7255d302f94428dedac4fe7fad5a634dc6e4dbbfc67d25c1837df17f5f5e433cb0a1ff957271e
z7480bd0d18941a813c4644dbab5ffebb2b395566e44be141c0bb413416488e0af4685c67bcdb81
z0c55124176b26d5f233fd3ed8babc0fc44aec113de4a1460c7599a7855d2ebfd7ec21e7c5cf167
z6d3823f5c6b3e1b052a8e500a2486c38e46a45044de5d3c72af164c277ec3cd38a5bfb8e2d8ea1
z45954936f7772202107f5e9d6d2f94fecfcc0de960acae844a0f26da096141d8449f4eb51a97d7
z5f8e83c51b7d846e0420f1569f2da4f71bde14ecb4e1f338ba79d902e312e7fdb993b80b3e699d
ze5ba9088270098a7d621708aaf6d28bbf9bb5eab211156c22690c0ed3be9fa68ca6c1f4652f7fe
z52839637eb12b1e9316a5a3d7483a1989be061c5f484a827da3b0c4d656fc46bfd341ca3dc3f2b
zea480dbcaba39d99a5c0e8e7b9818c99da63337151bd0d9c74d1f18388f3f96d0a7c8b7be6eda9
zb08c8462aaae1e7ffb93188bdfd4ab49505acf43a5460930df4b8c6a2daf6a4c47819b6e0071e0
zfb6a741b60f831453c71020c64a896620110d6bf1668145bcc977c8c511523aa74003146513029
zfb86ffc15e6c3431e3c78d1bce3e9bf717288747fb571fdb479f5a8b4328d1f765f1e7ea9ab88b
z6a8b836e8b0b167817f3ebcd119d56cb0ea864fca298e25be6fd0a0cfa158a30f806222103987b
zdba21519a02b5caa7fdd878c744d7455aa176c9d0c9c8eb3237828066ba3b758b00fb320bc29e1
z7025b43529d2e72f828211c4d8b23cf7503e88777f781884e5a62369989c4add5f112db54de0b4
z3c0010fe7e1dc57ae5d8b099bdb97dc07e9d8168ae642e8db5700cf2f91835a4d1e4a8378b9451
z845f3248f4345d6f1e71a8e5eda1967f347af545207787c189af3f86e4b16a46d8ef3365268c92
zd434158ba6c011ab437f5112e87ef4b2b5942df5eb87cbdec662f5643620fca68a2d206dc8c23a
zf5685a8de8038bce76067f5cede28d31109bdd38e0498756e0e3454570da36c1035c7f3fa37aa3
z0a946459c5db2ed19607efd3c52a94ba554223e746be6490750653b6ae965c57d22568e1763dbd
z16be2e1560e806722568c277d1012605c6524841038988b195d168daa9483ceed5507856ee5c07
z73f3b25fda9f27c5981c5cfedfc16dd31bee4e47b48646a8638f212cab59f001017826952fc78c
z12f1b53281758b3f8794fb6043327102e63b89cb71d3019b866e3fe6279aeff61f6b6962e86616
z1e09da8105d48271e518fff943a2311d1ed3f6b167b192db86a68a42630795f875797437d64b01
z79623d553db3d5734f71c72eeafd192ab816d5fb7edf7dc01577ae607f000be9b8197cf5c9da46
z9d2f13408a7a7e05c77182c6e6c5f9781cd5ea2ad0de257ac3d3a89bee5f2c2c70ada75e17ec4e
z3893c2da2fdbbf6dd0aa70d8b9b54eb1868e7de28056918f42ad044ed6551050af91ee3da5512e
z36724d976dccf2c1d87ba5fd2e482a20c4f1588a345da049fe9c840c25c341a30ad09e473fef3a
zfd7451e72fc5eebc929b0254b0bdf9ec1ea6234612fb52249ad22b1c60dea8416ffbc221ff887f
z8e9de5119651e2ce57b74fd4bc7e1b824a85c2b2d708596495e429f563e1fd63a6005257f22fac
z5c3723269c535c1dfa6070087bb0fe8e68284f2ecfe3e85a89facc80414f28757cad85d75ddf7b
z063dc649997e773274e2ce17e729cb1ff2ac81a23a35e3dd706e4fe63445a2d42d5fa01dcac3b2
z1f922b27f2f41ab9ff97cb57528557ec4305b97c90869aa304fbcc7a7a8cb368d8f33996860870
zce37b0b57a0a847139285f06a2dcb127524a3748d8ee4175a586377afe28d47750907065b6e756
z665b7804ce3dc095570578c976b2f545c63fb4f00537b0231038be9deafb0c8a8fa5d4de757a2a
zaafda858e2773a31b49fd9d526ff40c9915bc37994aec2e5165d64dddce0ba3ff8d5277975c40a
za24d3676e3c1599398dedefd6a5779cd967d79dc784b5cc146dc33c3dcddd002e23a61986537b0
zaf1eb0a59c34baa280f5d3971a7dd5faa0000d2df3133fe09d7ab0273f780fc0e6265f55a31460
z47402ec1ea556f3e50cff75e0b508be93dd90431871a4a1cdd52e1d4a2a09029eb1f1225cf31a8
z69c841a7cc281b92603510716ca80183ece0bf8ce8ef80d9c41b2a1b1686b0645e08492c19b502
za26ffdd2465d111b36e0b145a28ef70603ec3effbbe6fc994c94f046efbf46bd8cb448db2ca758
z77917cbb7115aa17cd89fc14fe4e2a3c640a75aee68395879ddd784351d97737974ee84a27d979
ze999c67957b14c9aea4befb549001be7a575b0c8fdce27848bd2f09db4985a502b7c58fac88f56
zdd29230cd2c8f2e1ae23fa028dcf4ab2c99eb1995ac959f898f9b549f4b10fbfe3411a972d9fa3
z87b4b332233df654446565ba25b52f6be1204ec16083261fe03731c365b908d49a40eb36c0127b
zfa57213a6bf30ec3d64207bd1bcf15139021f596bf3f6cb7c5d39ee7866cd0002a64a5227489c3
z584d6e86a3f3d3f947a0674249458021ade432fb9a86c185c2c3ceada02f00fc2f91cbe69aba5c
z16dac4fa5d581d42c30ca210cca8bf1dd7c3a0490bc8466c7ff8be9bc239e3c08a20b5c97dad4f
z7b2ea0b900182933fa9b1203e245904f13c5874d15acadfaffa89fe142f178def72049a149ad0b
z91d0ba4a234c5b2b7faedaaca90572c49244d8c8a86819eb1e3c12c0c30da2b395f00ecb82ba80
zcb8a4787f71a1f2dfb39d04081552a3ec51dd60385e1f392d9a12bc039c548491ca734fe09ea2e
zaaddd9a571fa8d1f394dcd26f87892362bde405afffe95dff0e15043c3870cd390a4f43ceab17a
z84287d661de0726609b961e8dfa2d6fe3e79c64f4ce5b9aa6ff20152cbf27cb7cfe050a8a7b2c1
z44cff22f62ee64511a93c618d46886c3415b0b5a9f793aab01d43cd9d39b078172de0dc487cc83
zded102e0361374bf513d662d46d8f04b0e6f020956d73fd943e1f53ce19790cfb1410da15343c3
z4496782fdc97292e1d79b5f8e9bc18ad6569e48a67d4b4eb93d47b519024130f1a1d6168d74470
zd66624e8cdc3228cfeec52843b0b83d0f27f8e7629a451d384ae5fd703ecd69ceadb0b2e4d496f
z349067ca8f0befae63a59b69c559bfd007be59fbfc781bbda2d3d89dbb082dbb9e285f97c7d049
zdb63a99685240429ae48bab8d38a8bb7305eb89ee48bf318228ff9173646be1375522550dedeba
z667304096593144b2f8aaf9ec5a0b5f513f067db7b5869806cb49a5f6e622b5f922374b518b662
z339955c5530bc1578a2067517c2b164e731f68b9c905d22c240001a9e10e423a1cd0df2e1c7358
zefab37e6cd049f9939fb6bb295adc85fbbe3aadc487bafa5fdf3ac267bf3c6ab5dde3b4044ccb3
z60aae13af23d5518e4145dabab8ec263773f412edbb7845f685fd0d8e457ce6522fc1f75adee1a
zca6fbd8dc93509e279034df0095f27ed8cecaaf1d923d85641021052ed2eb120c6f5711189e448
z21e9f7a2a18f776c050c37992c862bec2e76045e3ba68a05ebc5aac91ee0528b7ab98693874183
ze8f5ba3bfecc03b32f4d2d5cee4301c009c7fcdf848f265c8546efd4f922ae32fa8435db53a09d
ze2a93ef0bd53e7d31aaa09efeb01d6e0956137b904ce0572a306eeed7017ed474d7387b97eace7
z5dfc44cf9bd44c10ae3acaeacf33c76cd8401e62035a4935c8a3c3e6b3b797612e32dcd0c6a031
z4482dc9d22ffa8aab059bac49210f239d8832ef9f6e6fe4ae0273311f8552234893dbf7633e85a
zd5bf1d886c7834f5e28f72f7f718f976c7a770b3647cbbb669d72a87906fca08792cc674304216
zc9842942b8515ff1b2380b13821be0747c54fda8d2d09760e718b4648ed600d187360f5a39dc09
z2b249557637201612932bf176bd38f0c025c404ae7711ded057cd70b3589ba5d414798a94ec1f0
z18ee0d24b2baee41d44699e13bdf273c030ddee6bc927252fb656d7f6eca74cd1d01098ecf978b
z51b0d02ccc5eeebc68e4c9024ad73f754bf98d636ad277571af72f57d7c252ab553473bb405eca
z2bef99927c0ee0c1c07e3ae59f208e7e347f5f0084b9dac661169260a9a87b10f1a242e83e6b5e
z3b871d66123a51d8f6d86ac19a8916167720b31167d765a9487aa6cafbde5f8ec29aae69172d83
z3a8c0fa2106a23b7f048768163b6a78ee01189fb78265b054d29f724814c7cdfba74a08268c934
zd606628a20f3f5b2e103f56ff134d4eefba8a720e03a5813d99e049933ccb752346dc340ff9a9e
zc83f909dee511408a2ec332895cef1d49de720c0b3902a1c6f98ff1ff56cc56742c83b4d13dbf1
z05f960febef40013fbf2c3163ef37fa9e805eb7d383a69ea420decefec94b762b07d9af496dedf
z85a02c35a63a24274d383f09e7e4fc0e99e8cedb83492c45401fa166ac6825ef8dd25f793c2a86
z7d56a951122dd3058a8ae50da5cc43d98d021fd990884473f5c83b5a17ffa776ceee9c0460ba10
zb5bfcba1d12f16ede1733fff08ccf7ad64e9bc236446dcd26ac2a4f8522b224e8da6090995d977
z6542f25ddbdfd1823dfc82e483e2b17a1ac36c0659c7260cd0ee4e9f678e3452f33be9d4b28bfd
z12c1b53b895d7dd8d80ea7b00831e6694431232fea8ea37339081914d335f39296ab795476d82e
ze3fd578c1a68574c7fdc37d56c3687b9896c8b9c2d8e160330cbadb82686ce6134f337fb3f5981
zd3eff8630080237352a4fa9325adb691c4a7f23370d3cdd003d5c70368b386b09faf9ffc96dc44
z6aacb84618ef6c2192d62acf2286433b1468d4f6a0d4c8ded3aa191d432f41ff84b14f0658aac2
z78d6de9a63b73e33541d677748c2821ca55ebdc81a64a9e81ad5f9d4c62220b1f9c4dfcd5fd7db
z2bf0f33c47137973871e978d77e7c218bb0d05c01d1f8c7f144085ddebbb888887f69aed401059
zfae436ae047384588958cfdd96ec46e0d5aeee8520f3809e6dbd35ad5439dbd84d3d923490788c
zbf83e64ef1890d4e0a31b8d8ddc2660aee321f8dbe6b0cd042416f55d9a8354be819dbb1334af2
zca7feb4360e98c3cc538d3f8015c2aa440e275e9c1427b03e70f93fce1d72552a461274ab93ced
z3b982750595001571535ae38e582bbbd4a002b096adb05dd3679c79c5098ce7856381a228aabd4
zc96295bba3904a7fa6e2b92395369b868186667cd8caa32471817ea3dd338e3c35647230170e64
z1301550f713bf9a76d587f5f0f35e81292fd7b80fd949d00ff7da47b1cdc06e5ad8be19f1bd506
zbfdcc582190cba98f92bdc5130a74b3d05b0abdc305ae78835a1e3b8e7c506ac634a3bf1def3ab
z5bbf0374b7f8401e071f65d995193cc866b953fe351804016285ada3eeb022c10dbd259ee3e7d7
z30bee432e3c222085e9af405597aab977c2467aacb59e67dd48d79d0093a2eb2c6e9413779a3a6
z81056d1fb3af12a5fe33f47e682a0fa8332cab6258b0de8f311405e6e08189b7f4fb546a7fad08
z2cef4a317da826331d9f1074c0b6f5681789ec1b9781c43b7a61b55e3d8d1c8a16c884e1e2b555
z106127288a379f212dc5036031be66cd1672f974acf687565b68861eda50c837cfcd256b96d3c4
z87749593aa0876b27f6d28b44f13940f017b2e42609aed1618f62a6a7ba03594f51c0fb3307a03
z245338d40e4be59aee12c849c5845c72fc6fff941a402ed28738961a1a0fb1fc377368dd2008fe
z963931b3dd0aafb7bde3bb1ff09b4815335e6bbc38c20caa2598d3734a25abb35666c1cc65291c
zc44739d2b37ca69f43d11f46a66de882920221409a9dc6ee3594afa897510394ee7c45e8ff3e97
z136dff5b59a31cad470c0ede34b640dc0a6b39c882fefba1bce25330ffc2d8fbadb33224c1f289
zd5f819bf735c8fd19a0b946682a9125642aedcfe5493ce3adb21e89fab3bb51ffcbd4353e9ccca
z18d2f0fc7962ea16a9609041fd94845b1077912657f0cf4e246b1349a61e1f029c127f2506cf9d
zd55c8affd37d05b5da99415b9ce9d5ef19e8f28b0cba6b2ac02efb7348d7459b4b1d8f66c83d7d
z365ce1a480690dc6db3ee55244fcf6aaa9c118944bbe242a7703eeb36a3fd058130f3ae1822600
zb9c81ce515b98a1e844f0a6bc35624b8817e02f4b374446fe574ba2db2226339cae157c213064e
zecd4d93d18596534a3c74bb1574b37741f24a4e214a18a3aa3053ddea29e21b5a2bc7820f91b6a
zfd718fdce89a98d5c61af7d842443acb7946c538abaff9767aa53b0767cb728d6346884b98c08e
z1e632be36490ba643a77b7ddaf2e0a0eff855aeb4b4337caf015b957d4ef732d8fdc811d21dbea
zdc09c8ddc18de9ef2b6c9cb4e343640837cf02afd580a9ab0c1b37896611b8d9c41ccc02adf730
z29264e7e88ca2cb459694d2ea111e60b727c5f198ccf7f3cb633eb4ebe021a51406d02f65c440a
zd7b4ecf2e2018207a90ba95a19c0afb629969dbb9805c3e7e3b84fddbfa019108f4d7c424e2a1d
z929db39176282a0dae9475b31d8bb67dfdacd1a8b5fca2d74d41569176901308bce0c8d86f3e64
z01f4a0905a1a3ae701f1138f1651605431b69e87e87beee2d5383899313729d33ef599a936fd9f
z7b2003e31ef08bd15f36b8f477196758bdf7be9046bc371dfe51d436882268eab77142a129c297
z4450a4d05879d862c8491c1f5d8e08ace3b11ad598b645988838aa90f90ea7b3cf346ccff7c609
z24be72cdae8e9518a4c501d9ba99603bc84079bce29ee7e7e7cd54fdb2772ce1952a6c0dbfe5b0
z3a868873e12b0b6a6f9a467ddb33593842c330799cc6386eb47be05d96a223febb41739e8e4ee7
za6e64c8160f9d9f092339ac66cafde009a14fa29f5e46e1e4aca023d1af17437f28e7db3212361
z5042089daf686432706ab6be075031d3e319fe41d89eda7fe264c16e1e761ab553cd1d25d0cc6c
z25961d1c42fa51e7d75ee347d37c99b58d47d48c892951118c03ef94fee3c1683d68eddf3e004b
z08c58b08c01ac1a852153c7f05649a2c78863b2610c6aa3744134ac7f22760320c6d3dd70f8525
z97f012fa07d3f60700a38fa7678e336f4bcf4440494b517307181e8939cc52b904e0116020b8e3
ze8fe2087250556ec08c6fc3800b456af3d5e89858fd1044a61beb77f8bb25929fc97b87924bfbc
zb43988e1d2c2a3a732a2305366a0d293d9694900abff0cd9ba559c10991f9632f831982e0838a2
z28cf744d6c7e59df2be3019420ff656bd2cfe3d8b2fafea6592f53ac26f87bd5336f73a7c91998
zf51a434455117cab00744b9bce7118e3376945c84d86c5bd49a2bd598004ee8fbe8003ecb575ea
z06a69defd1b1584edbbfa60ce0e9735382dbc308833b43b63d1df0134a0760294abe626cb832c3
z5b2c2bd690521a9fa072b3df1857dcb7ba8f584e66bb02c4ebbc73b0efe255d1bfda2c922181b7
zd3de09fbae92eab44b746fe7a25b428d35f5b10e1214c27c30e21957169dd8821631faee14af15
z8d84a064675d639dd612500b6402b2e76468d2e2c85949ff4a68bdd4f09a003e472989f7ecc4ae
z038220a343ec636c14e15aba4f027c240434ce16d5e995b40c249ea590f2b4df1c93e0a8d03d86
z6f5db33b8e8a49e48717a2af30a3869a34d1f29aec75d49eac2759d7ba1e0fc95b1bba1b0f6121
zf661bc50aaa200efa3b7bdaa8aae9a37abaa5edc73d5aeb92b16756802f7ed9df6ea4e46ebc00b
z71617679eda398f86694ba12f98fb63cf52e961efdb05d9bc9442a522be2194ed92c7edfc4e328
zb84131e73f897e38a558bc02e413e7d64f0347b9f5f8ca9b16c31cd9baa7fbe20b0db5f48fa46a
zaa666260c3c8af11f3c7d2657e0fb6d29b89bf120f8a204db97dd8eb33b17c0938515b10062af2
zd9ba3ba5aa8fd1e6cbfd37ad53dc72527c56e7da38fd569a4a28ed752c2c3d5310ca432a5356ce
za37380b3f14366366c55b6212988d89a62433b5233e185e4cc1c5d958ad0748e1f7001eefcbefa
zcf13b80e59418713775639358aa8a49867061bbd8d5b5fcefbece5fd7b3b1e3df3b1ced4bbbe7a
zda927502ff80b62aca76776a221e6089fabf837b0f5765012fb088d93ed4a744173fabab0595a1
z94a0a9b41b80d586969fe844211ad6b3e5217cfe8858716d3ed4efc72f2df93f1f159cf4ce0eb1
z95d8d76bbff07a0ca7e50bf3c81fbee164465ed3bb4b914300b2597b1b64acde3d8b82ae7c0bd0
za8a2ededecbc84a5f9bb0b886df59527584917badb548750c910be2baf602b020740c50bc6dffd
zdbd9dccc2f138c087073f21b0b88e729b9cdf530dcfffe84ae7009f3553e8c67f880aaec04d0e3
z3295bc09cac265ce01239bc63377d76829af44f9a5f9aba4c5cd9b0659694e2fde70781348084b
z777187561a90c8eba9a63a9246c650d7f06a6df21d8dcdb973d9e806533db9ca104e3c7f838646
ze253250a5db988ae610e526cb028debad0963afbf5a0b27a00ea6f592abf1e1bac38a3acd4131c
z698396e1ce44531c37c0f4f29dffa14c5f4a29da163aa75b20e9758191f48fbfd1fe5a69bff868
z73b79d313db5fa0f6349e440c8a867c17a3799eb7a08f56002206f6e5ad0f96a0c1b952eaa025b
za6531c2c93bedbe743ec802791da8832fb241ed80984d2a63def9143b14f86d88065e785dab57f
z4ce010cf32b80b22190c2b27e159d9d30a299663c5ab12cc94ca473dac0b37f1b1e6c3ffb52f2a
ze8f9cbe881d6e6f5fac500c95ff321a3f21c6299a2eb9df5b66b05e0a97e24c7c5d5a1ec255fa1
z9258b49879e9ed81a6c4c27124ce4fd74d1af316ffe591081313570a7547b3fc50de784564262d
zc0a6823d59c4c36ac71da5cf1ce7c1c990ff7b987d1523d5e7f33cb9bb3210fbb244b0e7adca6d
z0e4d1fa0179bf4ec25b320dbee12f571b85bec8c6dd39e9fb4075fe6202abe4a27628b86387598
zd3222cf7e7cc93140079dbae6fd59e32544b640f2995b192780c33098df078f54b674a3a1b47d2
z1739f8229ab6216be22deebd78f7e530aaef941392551876b92342d7ec6820c037f0b874d6b848
z2f867790a247cedb11a1ae174687276626ad776da38b54ca9fdd3aa86622ebf5edc641d8b31ecf
zb5e2426cbaa96931c6eec96229c68b2c6f2f20922f90a654bb9597ae2fafacd3dc4b53f8db5504
za1355611e19d4c71f2c45579332351fa7f5c5b881c8672ceaf70ec83846dacfe5843b7e0e8b7e9
zf94748171623f5f7f1c677ae95a3446cf44abaef0d30f4220f23b901e16629c63c7e24c6fcd632
z667c63173289c83e40f570586f2f7858d97e9b8aab3f21ff37985066deb5181034de84384ad730
z33abf726baf51868968b0cecc44410d2b6500bbc64828ab93849d35ea2654591e06350eee76c53
ze5edbb2456812caf9069940794075c18d8e7bd8e974eb2567b5c23f6fbbc0d8f63fedbd0f8b317
z135c681b015682a3ac7572752c5bf8074987e0ca54bbcb09f7ac521fefcc94da7e0d66a22e72c5
z51e3b95be506af92b9b8799b9ea820f124e219fabb12aeb23b6a8653e335ab119f2555a03e9f74
z1336c44f3d5be185d57fba61ca945ae33c668d535f799a344de757733219de464118463d787221
zfec5682dd4e8d9a1766d914ee5a9de09c02ce008a3a7c77156cb3c76d78c90119c0b912ee0b691
zb5d2e625d24cbbb154ac5d2a97a37385e25a84f87f12b651a774dc0de879f8c5547590746a60ee
zc9b696307f6c4098487b462afdef685c59df13ec203fc4d136513224784c413091a30101c65b48
zed93b8a974c1874d6309019fb1c9875c2db2941d88e3e5544249baa2e122420db809ad098d02c5
z309f763bc15eec44f146ff39ec6569933129c5a7d52643d90432cac82e9ce2ff85a65d00ad326e
z61b7f4752913d803e4b55f56174e034563f3c12cb1f70992ad731eb4d452e11a811fbc24cce1ed
za13e59850f7564ba8f0f73d8df40befc7e71dc1053804646aa90efaf9aa540b5b4bba0d2819a4c
z378d1753383ad1815b57f07be05aa71ceeb750810e2c9575fbed2ae43df442b6a230b8d189fa4c
zb2f684b49f275fe0b5b6b205e092790bc134fb333b920e4217ae35fcc3f0fe7f1771df666ca641
z08a2269b8c66216e1742402cd3533cd23fa7d4ec3e7e7074fc7cf1b2ce81fdb9579f08c3d9eaf1
zb0d5111aad1f891eb624c8fecba37466c65250d6328a29982519b0af3e1ab3ba44da71293b2d8f
ze16bd44647dd055d9aaddb9252117b80bc089706cc6851485342715c7b78b8991f76e144accfb8
z394a537a8fe0aee199a2bea98b48ad5e2a9f8e02242368c59a7e9c77b525201aae233c5c80d1e4
zc619b64111c82b62a779c7f30c68139fd82ed48ad6e287418a213d7c02380a4c4b8593734aec8d
ze658d95481a15ff68508ddb870ce05bec04602c99c6fc93cd20b1aaaae8a69d65faee6bc7468e4
z9e7f2e9250571ad937fc93a163027e7f7c7b13ad3991cab56261561804801c7bb1dd5e46b1407d
zd9997b4c9d9e6c9447dd2f9eb9ed334f0e0f5eaa45a83a3cf5c15b97f78edbdd8a9b24a2161a4e
zc0abcc729f9cf3ccb6c0a8085edbd17058ce30bb588c1abb8fc6a314ba6e55a3fdc59183b6dcd1
za0ee0a9b95b72031104a96173d86a162965fb58721b25924702a54aa7bb12d90ec938d371e5e65
z46811e7c01a80a354243b0adaaf5f63f7bb93cbd966abed7cf4badce7fb7bb4a84b3467a965e87
z027a145b8e941b6256f22790cec92e3944e7a31ecce7ccca517ea63650bb93ac9bfce8e3385a79
z01439e46b08a2f21ad5008168737d64d821728df23a2752238fddeb64da49872bf6133ae00db2d
za96a014f6a3ab5325263223687ecc2c3f23b29540e0f36bfdcd95e16191651013d2eec47b1038c
zdc6be57a5149024cb150d260874dca91b18dd44dfc3ac770541c1213be96277224f2b37b99727a
zb7343c045ef7b378ed765f724187b216db55cacd86acb63f3c8ca8ffdd6c5959c5f9c26e145147
zd731589a89619f9f6da1a303b990fcbca6d85b9c1b25cb345a86cfc5d56c2184430e60038d35c9
zab781e5c94078d154f2ef6929f370f1821a282b1680d36f66921303821a2a5df85dd09bcdc998c
z155f6eb9ae814fcb7b5834e5af802f2b35173d41b065ee6d111bacb304982a4c275a91329abbb9
z9055eefe74b7def219e7087d5d53f39f3a844d57248780b5217bdff4b8387d60ed049cedbf143d
z4df47602782b8072363692f2b97ef79c89613ae380f1b2a66d969d7cb4f0c01f0c5a2e2508079e
z9684177d0de14a5589bc1e7dba3f4dffd2ce6f47da055c37cd575a7cb15a8d361e7ff753eff065
z12e85101ab667bd64aad228bf57a135788594fb32075938991e99087460017edae4466790dff9e
z79d2b597c9556be6f4f235514e132f84100a187043e49d3540800092e187c1e1b4fd2f37bfa65d
zc64065edacb0dca0a774c2a92b1cccfdeb8c248192c94890938ea086a2826a4a09bf6cbf854457
zf1ec05ac133de0f1ad6d4e92bbb325240e4d0088629a6da295fcda9d76e25f055b937ed49c5fd9
z229cb4cdcf2d5341cede178586afdd0104cd53bf384101418c1b9188da670e4eb9877d8de4e943
z99071fd9f7714d60ed225e082a192dd69b12c6e43f10c12a57431f30c120902ce659ed3c5a6b87
z9888a2887757d1c48f57e3049e3b15af4d58f120d7170c2d6614c798ed22154837f6f1e3fd85a6
z46c617b317f307915b106b7e820a85246b32bfafa69e6da10a31ae188737645143d31a7933012b
z159b46c03663acaf6f4d1cc5915f521e3f901c3098441536e84646d1984560f712003f76a6cd72
z56bf85fc91e8e325b7949ac8a7e422f8367662f81cbdad5669c028dde499cc6bdfa974e9c40d3c
z9580812652b65978b00e0757f10e8ddf969548c740b7047f2781ab572346f1fa066cd57a54e98f
z5f07ddde6ba4dcb9b951adfc7de0aa3502bbe5c854c0ad17beb20b9abbec4c730e31af75215a5a
z936f4022891395facfc1de32e0e96a0c4a317bb51caae97d484e4a7df2edd88a0faf0947f1e411
z6556e928b35a0553c3e81d4ba00225b3980f273450dce01ec0008eff91c11d86707db4ff710882
zc06d090775e72920537223c3bbc2c28363a1d0da9707e5a9f3b37e2a55a3b40d23e47105577210
zfe7f1978c97e57588c948a56a2069525c5037efe8db8cb268a014d2cb59280a38144f95107e220
z04c5f3d8591c7b9fb99aaf9f051747909be6e5caa201fc4ffbcc2f311a5beb0b2f4362ef826cd2
z37d127cab2eb8fc9e1dbc45dcd688b815108015b8ed12bb419a54e03fe091d50316fbd17c1d7c6
z56fb6bb12a49ce61f80513b5a9099958d140562d4109787c2f6a6a4a94e6596a0ef55df0f92575
zeed5adab2e87bbaf385b4d26f8f531af22478def63ca3fa85ad74b2f13e0c5798783372e038a77
zcc793088cace1d4897b82ebea491d512c58241f89fab9642613acf19b6e5e9656a9ac48d5e82d2
z7b83da2ae55f3bad533ad9669e0e5cd4f2c1e56e6790a545dcbef852d752c9ba18e2af22b6029c
z465ac313d811d9f56a57a8535bbb75577fffd03b915348cca01b6011789bbf9085d267aa660b2d
z0b13cafd1d7c405bad86b2804db009ca823cdb63fdbfe0c0995e981eeca41904360bfdf2aaad7a
z19d9bf29dcb0db8c5a810e120b1a9f1f7fbbce3773fcafb442abe5625fddafa88c3d57b0a3ba31
z3a797700691173c4aa037cbe3a9bf018435d2f0116675bcc2adcce9d782a20b9e064292d09c4b3
zaedcec38d2c5fba93d35af362c537b90107784aafca0ed786f8de849fee73b998980ddf9c19280
ze8569aa6d4049df0356d0e9c0a893b37461f3915b683e42892217dbb944dc38b6e258a23166a90
z334253c2e7af48e1dfbc9bafbb087d49e652bff8f62a01cfc5f728c7a39003bae86610413d4130
zff89a22818750c0fb95c25fe71c6da181e7929ecf1c78c91e45c7b48f76f962bddaa5eb7994689
zcab27e88add72607edba2ed634c9318658c8561c1aa64b86881819fdae2734155de3e5ad46f36d
z573d351a990e85c8978452f5ed59f9ba3b3efaac8bf90d8bf42b85a3ce42e4888012c1465c1412
z7c7445d50e7de70f192988e3aa012b3f8973b46d776c65748e4ba28da66a4fdcc0ba44a9a274a2
z215670203cf5a224a230daae3eb7f2ab6e7b5126ddf03cec68f56486870114354a98aef83e5ac0
z6c754650db89959a9219602251f24f24dc369d3d21dbc9134267e918ec632c7274ca68ddfe0558
zfd1526fc04cd4b275d550f471f866709f078378e136a519a3b4231803bc0a80d2375e86c1c7489
z05ec6f7bdc7d66a12a8c5f5f25637c3d49f41a7b5d4551046a3f1c55cbe053b1c404dd4478ed65
zb46e23510e8fa77d20860fab32be9774bff691d20800aa8a20853f4fc828292edc57897f13a0f2
zc54a31d075fcbf5e3b7dad84f785844101a2e823a3a0877f4235dead03821823480725179faf8f
ze8c5fd7823c9cbd2455904999455ebcdf7a08f20a4f8042bebd571e3d88038b647d4487d6cb196
z9537cdf40cc015050375e3995681e0f1170b4a991f95e11c29ea582314c4a6293a818f5f4e3a61
z5cca13a79f10138ed9d0d5d182e880eedd25b19dbdf27199e91556b190120145583dc043baf9e6
zd25702ab1b07139c4c8796df0361124b3ccefbc715cfbf051f02ebb28922228ef8edb36906716c
zb6d3997b4704a1858a11ec0f8ac6fe27bed2484e10ccc765e6ed0795f7a50dff57217b469a8729
z09c289606f0011d3e6535909da1ecab314c649515ab63beb5938fe12238bfbee1e21ce4cf7920c
zb5ebaf39d1c1c52db7f9edc9e53332188cecbd32c29fcc9fc912c0f11e6e0bae9f74f28e0e3c12
z54067e457a33e89ae2644dfa4b5508e347fc0b37ce96bf49a925a22f9ff4329c4030ea854e97c9
z859ba27ca4c125efcff7c05ca7df28bd9984995080b4b72003be125d277fb979ac7a26d13592b9
z0878c00001d02206f66f4cc8839dbac2273f5b8d8bc295382cc44acadc7c602af96f9bffdd61ab
z5782c545d295d13e02f0cee257b76507592551aad896b57d07ee33a65daa6cc44e17b1de21aa38
z8de1c5897e66a0da6687e62bc28bd63d2b0555f7016281c7f624615b6fff5f311cbe0799416363
zcdd0f159959d8be48e2153ffa6ce38679194e6f06baefdd7a849573858300fbce60642671ae64b
ze1851d7758aee0b271fec024052e0c7a68450b8cc85ad6c5900f6d60e61bc22f546ef9895aea9e
zf98fd0838d31fab3b39439a80a7218fa12db948226e69aeddc87f1e21e3f7fee1fe7d075143f49
z9d5ceb83b17afd1b46b383d60f558afdd1a78fee0e4d646e494a7707d9dbf21504f7dc02bf988b
ze05a3999cead5da0f5fac536de04bdd153477e41ac85dde830314ab68f6be8438d052b3b6ae2f5
zf71eaa7d694de88d4c487a31a639b5bbe40e0992120a5e90d5d8d3969680a7466c13cc88151b90
z609e89b892497ac8879fe5cbff69714851d6677c3ee41b563bdf4664cf50f03af7d461f7d80cc2
z3a78d845af69a37e56a728fe4844d2eef77fce3c40b7038a2d347bba56911d23b4484e38aef3fb
ze1b6441d276a9068a3fecad98ad4b4b31bc9da68140aae853fd203bcf4e0484981d95d1070723d
zf0e53df783bb86abb42ab2fb119525bf7b8321125a3ed271e7255b916df346b674a6d99fc26856
zcdc2d64e24766c41f211e24bb3aa863445ab1812d05a4d8e80a55cf169eb90460a582676047f7e
zf151bf3f651cc4d4d823327fcce42304206d2e645f0da8a5c15612407417f609280ebe1a830032
z9cbbbf760a32cc58ceb10ccadc2cecad1de04d05343d32d02a415c21bd7e38c82cb66cca9cef94
ze13218c0e93d330b5fe508908324312e94aee027ddd2b852dc56feeb95951c86fa06cfb4c7ff50
z8c969e91347ec1bb96dea89f67af76d87b9e45fd00e867128f564bb18173da063fe219ed05c748
zcf3bf0b06ee2164451e1aa2f98974542353c613e63437f0653a58f0dc8f3bfe437e02729939219
z3216a49aece8204870c40955d34f1da9e2d5f5520d1b6f5b758609a444c3a08ccbe6160dff1b26
z3cf451a15147b974d24d59821537740ea3eb4e271102dc92ba434a6d5773df85dd4b49825e13aa
z705566a3a68bca2ec7e2edb76395640641770f4e12702181e83e39734933600f97d6db0317ad74
zace2396ee46868fa9e189170436a90eb240e9ebef1757a6d524f7113caa46bf11a747df283f068
z6ba747cf2dee71ed86dd12840f7231a06f6bc8b7b5316118e6985ffd36f039ec46f37437b3294c
z808ca7de10ea52115602e2d6d35b4f7d2f1f09446f04d3a98fbf608a65da12b8d0aaf763f9de2d
zb6787692d4639c27fe6dbd714a77c988eb968b8db2ecf3c2ec8fb42d5b241d21f2b5f8d54245e1
z90c4bb8829c120714ebf9e5a1259a835db5852e0e8560f306008730122f8380799be3b6ed619e7
zf007cac4b2878c07b3395805a733af9da22e32018e56eb726250ab42f9d1f8e5299528968faba1
z21eebeab31e42584192a3026311732a517a86767ebb5edec2977d121f74a442bab6b10f76e99d6
z9902165852d0b54d6699788f56fb5af9cdad34f92b7dabee1d319b92314c2a7d2d49573e0aa711
ze9863d266288d9f59d339b46a19cbfafc6b3d9e1c868ba4d24b89c1924acddfca4c84a1f2316ca
za7dd6bac947154c2ddc7e83d83b434a3ef96d8576072ffb0e0099689e8f40949a17999b1fa38cf
za7c29cbd8869fadd2fde79d939601579c9eda1ce700babe8fe468c21cf65a6211288140dd4fbfd
zfa19c0429579ff358067584c0009f1429f69421de1e1fa9bc4ca6bbb26fe3291ddda774123bfd9
z53cc0742b17ebd41db38fcc7f9d91b280ec9bc62bca291883081dd618c132bb1478ff9823bbecd
z8ff7d7100cd0e3e6a514edb0437406effad25600d2c6cb0cb3b1fc2bd68d0e848c5651732e439a
z6091b97430e6f4f6c07e12e856e55e1887b5b899a3dc729175fffd171d99148c97d1e726ada123
z0a4cca01f02dc799d3ae92ea03055303a8a2f06cfb9529136ebcc1e93bc9feae9152e33af15270
z0902c64e35e1bd0fc5eb92fa4dec6377b85c8189ec307a76e412f7498d9a75c8f2945c5b087a56
z5a5569541ead560c581f86cbbd3aa8e4bcfedfdb2be00848b8ea41f577abe7922c1971b0e02e78
z0874a0715f26f958a0b17168ca10f925ca6c3f1e141e6cfa07b27cc2e112ac5c91c218a253dde9
zef53b575463eaa499d1966c9a7aaad65c3ed64e5d451a1e106001297840a0f25c755ec96b54163
z6d492b80301c02f1cce6c2206029ec1207a5b1c6dd0cc4331852fb0cadbb6a059597f77d2062e0
z862c7efd0727c1c95a40d3ac946cbcb3d406d53e86d77c6db57cf1dc3223d9c700faac0ee0fa12
zbd4680ce3920d1564fd3c6a7587f4d5ff4cd604a895ff37cb0b76db5ae201376daddb1312c3380
zcdc4782cf618154834eb9351455c9e65b863723db4b9828d39af2ca135b743d9d0af7688e51ac5
z45b516fadd27682c8021a5778872c7c530465d679ca835578af9261ec7ece718a69fc7ebd20585
z5469ab367949523e15b66c211807ae1c5151fd61b0f619249849fa4881138e78b1299d4038af20
z03628ee44d694fd1dc5841aea4146131ea20316da14acce3d9e58ff862204788496c923c60a5cb
z12efd76f1a9d5413477bd2f58a8423d7d5bcb481adfccf662088ff9d8cd400eeff4db1ed7f4be1
zd23b9c33d15cc4511d27b5f8436d9664c0f27a7cce27c1415f412185610fd556f07f83015abc6d
z2d2906fe80d81ac35ccbee9659407b485d4d543e81407a1d4e72d4801ae5f4e9f2c325648dcccc
z457da2fa3e73e1e510aebae0a3bce34fb3b44093bc0d778893f79bd31082685fc0f68120b10a15
z6ce4e84db76e6ab588f75a25ee7665ff7b33271df8b2a34198efd010888e859a19aad28d1a3e34
z743a74f0bd85e7140569a2b64bdf783c93384a608610defcc257590200250a5b9149df66a5a2a9
z44b443174880230f3df7aad1fea532159a4dd8e3a9aa3e3cca9ee3bd206ee8611144b8e121f11f
zdfef498fbbb248a505ae1b55eebaa4e58375826f83bbcaba0db8eabdd1762ef16c78c5ece52203
z4ebfd16d66a6d1ca9a4a51a018e10a549de7240a4bdebfeb55431ea64d0bd505b67d8e5853d3a7
z5d1adcaaf8bd47c45739cb09bb39c6bf6f0b19214110979f24635331b01c17c30999a949c48887
zd1c319970e9ff2a9164827c0ee467af3aa3250ade2de7874f147784a3ab5dc6cdb2265ce2511a3
zc7898589923e2e33699bcbacbadb25a8ec115764e30a56107b5d4187562cafaed22b59325988bb
zb771b2b1d6cdc6176606dd58b12b9a62bb8ddbcc95a084796dc3f42441e7f01d4e7844163e56ba
z135a5f3847fa093bff7cfaf4b1e8efb657251558e2296a0d3ccbe6afdd6ec9b6ac3aad950ec37a
z68979cb906ed11963f8804d47e07708d4ccd894942843787d78d75228e6b3c8c426d28cd6783a0
z6771e9cd8c5e1e8c78b2cbe6d1787bcdc5faaf99ff65977272773da8e13c05a178ba2ac83321c8
z5467264a9aafaaea51905d43d4821968e5943af7813061b373dccfcee064fd504d5c06d586b773
zf273ab32a998a0b338e86e012af7bfa1caee520de36ced7ab01a6457cd303bb9e6151f9bb14f70
z8f88dfcca1050be702c79eeb7acfb6cbc201988f1c0f18c2b72689cb4047217bd9d1ca7becb0c9
z9c07bd2f3db328ba7c2a345a6fa3b9a5ec1fe11d4315586b48c49c6274eac3bb720c134c1c992d
zeea99dd1ed9f15e8b67c3374a3d5d9fa78340e1b5b9cc2717b7c9f3e549bce01e6bdd764cd6980
z8df4ac6a8504d162843675aae34354429f6f889a3ea8d4bae0f1b7601f8823fa4cffec6312bec0
z4a5421334ddea754001f1de28cbe1974b0c42772e37e3daf2739d2bce4525d87dc4ca60a04f613
z68f2e0d8d4b21f10b009e3c5331f0eb9444c154b1d2460d8efd6b4775a16c3a48d4ab536eded08
z00a023ae8e0d81c0e9355ad513c86777703b35531ec9da77b89c6e0497305676b0349b413dad2f
z31f91780ac8e7986d0fe0d258f4c2252f6e1a8f696e30993e99ced1caadc2994334fe88c5a5b89
z2d309d6ebfb7306690b0ca24a229e95e54159034876b5d0a427ccfb62b076996b824dc3363aaad
zf8832379836f4d71fe4b15bb07ef93a6f79022aaadf0c55ae4c10c1623b47b505bba163fa33173
z7b2541b1dc07e0a191862e4aa96c8faa67934f2960b124f0ad3dd5d8f1d5918cd165ea5825da28
z97035f1fa85efe8fa8c6b7629eb3a3b0cb95bf63ff2f4ac21e0ef3d238b90c8d3a91e203612a25
z5205e6a3e10ce29a73f91b09d545b82f66c8356d63713769c043b48b457215abd88a2d6f6b0b6d
z605917055bc2460e17597687733c9fab2b7ab0cce669e99b204b8edcfcd4918e4961f027592a22
ze3e216bd60c2aa592ef597078e02f0a811801d79dfb8bccde3039be7b9fd24c21fbf0a8ebd2592
zab988dcec3abe307b6abff210786bb7a0d7a27aaac90571c34a407ce32fe4316a460535901d5db
z37af5918104b94ffb2d48af84f5be4b8797fd06994972a20fa43898c36e3e00f5e9ae27c52ddf2
z8ed64d4260da40607c33baef5ce896c82913822af6669b43257b786465950d66d5bd954727e362
z69c72c373a37b5201ed0775d95ccaf30c539eb7cc0000b572aa181c18ea35dc7037ea7feeb21a5
zc67c26a8a9ccb44ef9c576584a651c69bfd99c2dbd9c0c08e8aa087406779136c17c71f450610f
z14cd2b2ac8da667d5bc82f092de5e29158d0085f77e4420206f9d76ce75183bf40760bc6ff62cf
z5f65c10583278b0fba56bea1ffc92bedf3984003df8464732a801f62d3ed9114195294518e19f4
z4c5ea82473f25f923a6f7338f8573de7dbdc7bbaafa52fd2df84bdcfc48bcf1d5cd5b42314eff5
zb092645ef6cd21b96af1caa14903609d440cce2d98ff41356c976155eb85ecae64d505ee26d68e
za0d47ff4ffc3228e11077a055b6b975693acdb2090fdfc17ac1db5bbaa31010798fdeb54c98a36
z7e6c51e760f371584fdd416a20d2f0a6ab6ca46f34f596c06b2d38e953e614bcff2f731f9085e5
zef891b14d103995d80932c77b5bff191584cf338d178ab0534225e53913eed1d49eaee1a1ac0d1
z10cc18ebc04929b66cded0fd709298396e37e4319dcb424c44df86a47f0a9f9948ac7703983f6e
z70c6d88bc3fd163400ea7808adfa0bf6790f59d9591c6a835255f9bcabdde8142d5530af70573b
z3bf594d2adc1beee497059099b8502ec1a123e0fb6500268aeff762da2ae3c872885287bb8cc9b
z517441abfaeb12164e90354569cd4af195129b9266b111bc8bae984bfd035aae5e37c9741aa4e3
ze4ce54dc95b30d52a184009cbe2f9d2f22d20e3d1c2fe769775f8a9341b4b0326577d5d7f2ac46
z69900656109ffcb6962cd17164783a372d21f97ff17e7b80bd09a9b00493fb0bb3aaaac70bc01f
zcade918436b31a711a50840ebd43c2a538d5c1074588a3fcbba3412b97e2346febc59afbc4c502
zb263391e6f5bbeb68158bdf9d33e31fd09278b456f0c3f6366e26bfcec70de817e0e33e56eba1b
z38725c6273e352588e8e2ca5f37d9894282507a6ab1e0f852aa87554018fa817654985ae12d809
z7290459eb162c147c4125ec0d895d36fdfc1aeff05f0454dbedc1c831508110949ad0de77102a5
z5c1eee96f6963ba194a0dcc4a1317feeebdd9b79b8036041a3f00fbb7c957bf9750a96132f9c84
z66dc9c61ae3d537f5fe71db220862a35635c7c3ffa90c9f915e41a46aa74239648c81272077eb2
z415ad2e37e8bfca738f961b6cb4bf55506ec8c61a65bde5bf89278c2ffb12f1d306522ffd73636
z1581b2747b4cc64bcf03ff4cd454dcad520f137dc538a70ce99f9205ba7f6c3f52621b87d62ebe
zae25f34d0ba5c172d3df163e9da94e7a94c1515f258b4855644a1e605f47b66ccf00624acd8bed
z330fd3f96f5fa03365f309a78d4965db382b47fb911053b6c41b23aedaf0ec8dbc5c5c4093eebb
z6f0647838d3752abecbcb3f5e70e851a119bcc055d77eac0cced39f00792e7faddeb64d846f99e
z46f5291a46d4fad4d13918497a6cc71f18daea52de6f8715e018707df0837cf4a64ab4c1194885
z6dfe5b2c2537ff64b291b427e3729b6bd93390536a67106bba99ab1a75fd1898adf6092c1b0b03
za6712e8e2111a532072d3507d5474001391fa066f1190b2c508dbfff6da60190ba19014891eca2
zc2726f8bfd3d1e41979306bd3e8ce5f150247602194afb2f9f79a3f68cba2f971a833d3c01ce31
z2e0f17907b6c1ab79fc1ee9cb40330b8a97a98ac9d1c0c6c316b2b91bc9c0bd9e4b6c710f8e0f9
zc1a3562c64bf74bd73d17f0fb67ab4c83483139cff379ca51639e0b07c06f4f3c3cfaade344a0b
z65a4a8b4161d66ecd4a7d12d5900d7e1313b2e2d1ad033d135b4dd465642eeb9652f9c99221441
z048f7f7f3d662f6496e843a444d48960c040686ad1f0a7eb1d1204b361cfff26a8988c19967912
z851b0e553d2b140ea15c11b06e75fdb67d7e7f54e93c34ee2e86d22ce0f3275a71fb268e78a4da
zea7af4fc3fd55f6ab8d98d2d5c830f73013585230cc7a448e803b4e0c46b28075d9e66c17cbca2
zce81e2e54b4239fb7e7d59bdabc3d438fffaad4d98942dae2a0489322f6f0ad80f716ac77df75f
z769866aae52321d4f01a26cbbc6b214bfb6892264309235eb871a352ba9f7be08ed4af50ef641a
za1a483cd1a1dd265339bf90d241a1810ac73539ec3edf63a01a443be403cbd78924cbb1c214c6d
z6964205543eca6f964ae99cc1bf6b6edfe992079d944f8e3a4056d417ecde4ff65ddeed3845575
z8617c105edf9a828058759b8ccfeecdce8805b9d58c643fe1f6afdd22d8d99ca1d6a159cf3f57e
z276d83b55001396abe7852599328a3932ef060a58fbefa5bffd0b28de97e2e220a1bef71391fe6
zb5d5cdd498a5aae3deb386d61a6ea4a1dd24601d061cbbcbe88a987f444bf627af32d07300fac4
za6a084512f1991237f559865250d181634413673011d1a53f8ab917c03011ed9dd39101e5752e0
z8ab8b6ead344b720cda08e32799cf61de9c7657ef0f9788a62e2e2b85cb029e872cfbe0490e68f
z2a4c9f0b87f78debd4e19ea5944410ab021d8a45196f95885d8eb158a0a4a3e0599b9cb3a483bd
z9a9c0ca0a60346e4663355984ef0746dc6f84a5891c28c50c6ced10961a60da49746d2f5937570
z8233c7c7e9772e37e8298dc261f38670867b0499669bc686837ec7f44f360b7422570db9619113
z43aa83cee9fedc99d138dcdd7a794224108e9da8da96593b9d7fb962bd2c37a002470af2531b9f
z221791309226cf438f076fc973d51ccede9ba4f2f405ae7d775bf04ad8d62c9ce44e105b010ca0
z088ac8864385bd8a0ebd8c60b5afe4ba82e56a655253d2f11a77f255915ffafef78fca849a076f
z4a9b614559657cd0a971d4a1dfeb76d0054c64285ee14ba78a2d9c353c7234a70fdae8c6c5ea64
z842c585d9c23f3b5185cb80ff82374c2483130fa9138afaa29dcd3275c2a23336c62513ea6397a
z574258fead5e5a56c4c48c934977b534ef1c83a50b3893ee1b3cf956ba6c70b69629eb3ee7b896
za288992820a1788f1863c5c75921ea0a1feeff26c1474c29b43bdb1f587326ff8fed05a04896b1
z58660f984ef459834d925d90e0ecc3c59f89e7198c75f0761b06ea79bde255cf9caf7ef70fc08c
z0b2e3f57e945c12d67f3ced22b6355dd0bf282318e3907a9588d13065623929db588d326270b0a
z3e448f33ed2a2dcb88984bd982fbbfb3508267d1d73643a10f6bff3f44a1f23101af3abdf3b9a0
z97e2beaaa2fa38a5bd8e4cffd9e6767ba1c76a889b85ed7f48fe780786b179b43730ef85b704af
z4f2a769128565b028ecd2c3dbd6575567b3cdfec626c76b33d7c9a067073b320c33cb4c61f90d5
z6dae1f2cc0c4c200891f92eb78f46325b6f47006128907d2806303dad8641c9939b4caffdfdc8d
z95a7c2e0320421f5c26594351dd8205603f71f11015bd85a800d6b8f9470e416137d1e50a6cf90
z64e97618c6762f2c2b97722e38134350e1b60ea90e513ee7a93c44ca6ba9d7acd32f71faff61ec
zf2a8e68e867c56b335d8ba21c741cd5869e2368cd39c41070b75315496a3c683bfec9ad3362652
za49d5b05f7653adb5fe8192c25a0caeb34cb197df06053f84f7a474d8717f41ac44fd0d1c875dd
z536a3dd067d3418116503b3a2d49650d2a98f219339c8464b24679a1250550685a6ca980ac2dd2
z0d73d137fd58aad37bc25edf88e1a4bd50bc40759281de1ff064578c0ad616a3b637201572464d
zffdf50794596ab2a584b5fb8dd492b1489c62a7aadf0e11d9430f1a93ee461e0cc9631c92ec2ed
z0447d1936fa78bae3cb2c6dd1553a4cbb2951a1ce2b5dbb7aa58b5330f4fda8650a138521260d3
z048c9aa8faaeaf978f6cc03703eb735aa796a3839478730f445bce13a6ed7a3a9613d9be83e54c
z4b10dfba49e570e56a66de9054e54acadcf2050eeccd5fda8a4a4fef0620d967b78c1e7fee68c4
zd3039859ea4b7180d4f22541794e07ae9fa7b6cb682922859ab66fef501713198efafa728ed32d
z27119c6926ed76308966dcfff012dcf0944afed407b4115fa8a3d7001277a26f6083c78d87389f
z576a48663bca2904ce8852a719fbb2966a99c7d00f95a6832de3192ffc27af6678c2a0c03bf17b
zd023955a4701643169a8d921bda5c53dca8c63ec98462beac6947b07c0178d285a76627a0f1792
ze9be684febdc991fcfa4d871f70bda5a60d9c6268c22e2a144ef8239a193375dbd2c0ceba45736
ze13993a268c4e2de4d6041e2d72a0d571e221ddb5e9941c0c9e739997a4f28fcf95bb759d6390c
z39edcf6be46231ce70d6873aa9263c60cc9878a22f9393bd045d874562633b11949e13b0fdc703
z2463ea92895f75f2f539a72a1c88c3197ebc070424607c98807fc789812290375f17757645c2cf
zfe73ae741689674f5b2e5765d1890f9dda1dd6d33dd34d22f51b971176648fed700b725fd88ad7
z13ad68bf5908a17d35a3b633f9dce81f61a68ecee64bf6c9af1c74eefac5987259b6809b5d3c96
z8a613357791ae15b379c565d69babdce2513a9594d87a97b8d4fddfc3478b056ab17b5a30c191d
ze5ce530806fc54e94b2cdc2fc0dc1d292eb75c027bed7137f00d2420c3066801a11a8923c5f9ca
za510a779c5eae4bdb2dcc4a1ca055a4696f495158e972fbbcd3fdbdb4eb5a2d19de14e16f65e41
z297f6914989c09033141fd3951e12fc7edfe100486d31634d547247c59b0821d50366b33e5a31f
z02060fc81c5dabccc63311d00156ef565dfade6559322bb393651465e703fbfc875c07912458f1
zfe134febf6ab5aa51075776ab7134be88fd6744bf0273d378ae6ac79206ddcbff185ffbc1ccafe
zb8cbbbe700a8a98e31a621ef0e2a10a8fbf2a9866ac60f3e5ec8fffa83a7ad5e0cc77f1723c3c4
z81b9164b4fee0860eea85f7fee11e622c773d061e92a10d8903a1c7998455dbd10e4e26e2e27c2
z51a1d7a0f39b11c16e5f566dab99e8d964aa5b9459b6636491b06376416026c7187b1beb2fae32
z3fe72ef44eda500cb9eae39496e99345182e8ce33ae8c1a04bdea50e169d5d12e9ab0f6ceca5cb
z75d22b02ac0c0cf612fe8e3a7a69504578fa18e815978afb53275265ff86be57be86456a63c90e
zc45cfe64f6e1da22f468afa6cf77293a166cc9ae24824c83257d2dbb24e90372913db9bac7491d
zbd85df4e6952e369a6bf8cf6939d540f1825a3a8034cfc0e9672c8c03c5e952e1f36c955ca8c3d
z222c223b3a39e42f193f6011b925934a7ab407ba9da0059dd3691c8a4304a5f1208118340f493f
z7535c85b0282b6ad4d2eeab204ba0dd5f6903c5532be9a97c02805e8850f0d6ece0eea22e1b546
z1d7890a07fc5ffc74004600dc27df5ac0a849cb3de01d58a85bb69ee9f7b3769b6eed695d6202d
z1c923859a4a5a901d70a1edddf8a3c7adb50523d1d29a243ea5011867e5a23d8b782a322bdb5f5
zdf2ab0ff18b84c5dea88dd083217fc56d8b6ac47455c1c0845b118716d0698f21d26ffa15e9638
z4883f4490a6ecb001bf88177fe9db3d00e951d477c8556a8e005dd841c4a1c6dab8b99f01702d1
z9ae14b19d1b2494c4c1e1505d9e21eca18f368ee4ac48368dc4592ff85503975f9ef85db727c0c
z063d9d75930770eccfca8ee9f82d77b3965a756cead8fdea7180fdce2aa056298c58d289868683
zc5ca06c07367183dea768c7798e10657bed78ff5b5e14aec08508edafb08c928db7a74b70f3467
zaeccbf855ced6dc3a1c447514da012a655abd81faad6074483d4dc6c78acb9d42e84584b3d5621
z3611d1e02102128c396477fb8a35b7eb60880f570d9b150afa87ea081f3205f2756574e971adbc
zcd52f9e702c865c0dec2694e096268a9d22b28b60419037c585ff1d9ba4847c3f431ea6e468673
z1768fdc434811341df4cb136b6bea1b9f956b4d61e07f2dd9db1099bdb716c43318058bf57c8e2
z7efa0a244edb3e65a2f08f5eab3418de51638a49fbea141a608c3a3f06ad4c513b89963ac7f63f
zbc868f887a65308621767da767de7ad0ea927c30dba576f66f5dad2a634ac4bf739c8c4137d4fb
z1d8646840c51ab4cc03b2447caa903f46a2e4aad1445500e76058d399eabedcf0a949c1fe641fd
zb59e1b55dcf92aa93be450200c0ed9f1ffd4ca246b765917a4372e2949d409d9bed37411b16ad5
zf8c7e010fab53ff5bdea788bc72b25e82344b8ac34dabcb9314735eb68670b0b843c85ee696402
zc813bdc4fbd98bce0b4531c250d4753379863eb49ff53fb30f9bf5b1cd5fc1b0c0aec1201aa1ec
z56b9589915ac5f2572b7187eb0412ed6c3a8d0b1410c77dc87f2fdbc65b10d40dfc8c1feecec9b
z7e76b530d8ce82befa463523c3e70324fe23eea9179088a959e9b006218035511a83948a511e93
z2adf2c1e2c533cb424fcf52dcd3f5ea5f338d57a85f020bed915c3b5a955e6581328b44bea9b8b
z480f73a9f517aa928efb65ce2576ab2b2ead19a16a9641eeaf7441160d0bd0c84ed372ec255aeb
zc8add0b1c681c005c2576383476f24f0e798a9f215d4ce95af050d54eacd5e46f6111c137db28f
z0b6024317cbb287ecb6227b5d161dd7b6fe8bc2d4921689100c6cec3472fe8117aa388cd78a1c3
zdba6a9602e07ba0a88a8f7d460ce64213e29d670a90dec61f64734416d666a3ef33ce772d5aef1
z08a0bad36f13a14ae8436f9cf15e16eac2ecfa59dbc1fbdb258c138c83f3c75c7a1ea277278825
z1c734996dda74391ebe4bac9265304045a23de7213651fd169986634a61710890e42984dc452c4
z4856aaa4a44382317376202ec73adbd35630c8358f8648af3ab85720925dda5a161e08cccefd07
z363469c392e8e7930b40516a76b0faf61ecf78ebce33f0c55bd00ddc593f9af29370a7f913b334
z6311e398e0fa7497af306440219c1e1b117ceab823d788f80cacfafd2537c90859f57b0422f6b9
zb3778d3fde7c1be2b3ed83a05fce0aec06d5c406d3b66f907a43e50b52f2619421517a767b8b8a
zac828fd2c9be3c7758cee2cbc759e1072c99654d2f731b5a86dc054b0bd85ce329cdf38fcadbcd
z9dcc0d874b4cc710fe73a33828f90050a9ccf2d9b27e8e94d54beaba4b40ad573d15a9fe80725e
z48eaa9455301724a381a7dd5f618a0ac123fab229bb97472d07111473034f4c7476b68d9c58eb8
ze355ea857fa3d933a1f7fb68eefab6ce5b2b56be002d93dd7c2f4c1c14055ac1342efd2e770701
z9ad730ba0202c19a3fbd8a0a942318b42b48abb896d1f040cfa57aedffcf9a433d210dbce303bb
z623490cbcc182e80c44fa28a79d21a806ca0e2e13430f36ef7c0ae5d5fb8952e9271ebefb61b61
zf231aea7d14a15b1ec9db22581b25b811d9640a0d90ceeec2f46eee2263f7671724ef8b04dfbb5
z56fb19a57ef76ad90e80600a77825a2d65f7564f7e65031561b249a8dff23b3fb2be0f75348b03
z5f06595fbecf17727a10cc3eb9600857fc843dbabbe68e63633cdb5098f25f15487ebb9964da73
z903e4433026f0b5194e92229ae6aaae7ddb9d52257ebee88bbd3ec481cb789b129202e296d4b8e
z73c1be9c7e17ae76d567a4c2e794b263de5e0a8510e615c443150c9aa258642e1eef592207ba05
zfc75117467ce4c771dc4bc01775aed66ac435d2dca532be1e690aac96017aba6938dd4ca8127d2
z601d81e10cadc1b1fb76e5cd0dca2e33da633240134ad2ec5d4ee2cd2e3cfef2221e50d08174c8
za8bd0849ce48582485b527bffebd8966db760b249c84a04bdcae2f1d38f8cb96d03a5734a07d47
z680f5f666f377c67c2705d595aec1054df1f5ab1dc1cad88cd06c08e4b47d0815fc4d3a757b520
z512d7548a5b5040cc777b5b1544742bc8151dbc628539d014b33f519a47f2f3391f24124e9fc0e
z688cacd10bb009d49e109f5ced93ee469444d228fb5c4c20662490aac9f5505ed29ff891cfb385
zca1577ea4dc1bef81f589bcc76c5584d188b1c58646733d32d962f8918d9a5baa902de6347822c
z232546079d49fad1638a4e2d65ce44e98b6040487fb5d0d8a12dcfcfb6a2bee0c446aa50c9f4b8
z7480b4a5eca787cb47135c328396ce201b77fca9c6834c82afe9e57a5afa1667a754c917c2e3c7
z15419f11641b24a5ac4c87b3b572ea8a152690787118011795ad84385b8e987a1e01a911856d1a
z763a8850fa19f0732e9081aff3dab0d8fa2a5bd7e6e6cb35a0dc530e8b444ffb5a0c4d1fc7180e
z0914961b53457b2185f7f41af5445b00fe4b2ec5fa90367af660de9796ead3c80986a17dfb50e3
z0dac43c4ca71c1027299b264fe3361c75821f0832fae56509f78df4a73cb888bb15916d11c833d
z18583e8a916bd9baf39b04d9f66e337c74a7b84e0f7371d4a6470bda45a261e820ceb19422a451
z190c1dc4300ea12500b16de791ab8ec8abbcf18d223a0297c058dbd00bb1d7f32c9fdf859cb213
zf76f26e521ee23d34346a0569d8ef91ea1fc55c204dc08f5246ed9493162db63b0ecc9c8814046
z9b26d824fa03ceb58000f593d28dcf7a39bf2c04e8caf94363ffe65f807b513bc3f33d934a8202
z1e3f7620675afc5b4b3012dd391c2a89f2ba0c75ce3d8c2cde5d15d0606b8f8e4b0d5ea280ed42
z749914bca6cf7b4d3ed7f08141504c3c76067650392575c0f9201757287f004fc7f04fcc93dab2
z995bbf4d61263d60beb81e29321b150d9ee09004d6202063bf0bdc90b3166b5e3e3044d1a36bb3
zc679225927b7dfcd11e2c22aa78aca4857e267064461a8539271e180e124e53fd6416dc1931b77
za2ededdfc3fd95042b050e1910a5ba2303bfa4af2e7bdd8814a7fb9a57289e1ac8358bd1d4927f
z186c68393deb84f7dff98810e2236acfe7cab7df7bf3e6fd82ea598399574ab23e2e410fbe0ebb
z5bbef09745b7d617e519c36d245fff3413889c39651a33ed066d1c28fe800582f4e610a616e0e2
z338d4e8452ca2f5ca78168aaa90d668f12a1ce670de7824f1573121792434017fd41a081a4ce88
z8a6423bbb4d181e21d5e79534fafd461c65c956fac06cbb943eb9732f4737f58717c46a62518e6
zb1825b17bb688085c2178b298af218edf7699fd44876cefc0226d53d56c5743698aeb37315fca9
zae0bc132784db17af3d94b6f9c82b90ed580d99c6afe70a9a233e2e001d82e95e6c376bb84ea32
z009374ee348300705cb9187f252125ff0761ba295209c0662b07976939602068d6f53e93d4ac33
zd2b280b7fdde488254006ec459f64bfe151c51d35103de2bc336f4e2448077351c76c779ba3019
zc7e339e685688b0dc65d5c6cee280f8d66a2e06d5a83638c6f953b3e121f4615bab082e0a751f8
za981c8b669f2af79c896f088207608feb68aa1095cca2039ac2be2b4851a91db04d0643549127c
z2aaaf58ae5a75946d105cdac4f2e625060cbd3d6d222cfc54ed5ef1673c6744b77158cb2890028
z19675c6aca8de96395964b3e0a15dea4024cb02cf9aad682e806ef48a98253969965055277fd20
zb21492cf10940a72703ad335608dd911173db345c545d8a04b009078f9ee0fceb0e001cbdcb5b6
zf7f0fb8687f8985ba86e04ea2183ddf7f5d40e402eaa7becf238c6abe5bf429a3efa408febe7ec
za2493c7de9125bebf59451a79a625ad386862e9e9e056027c94f9d0a80b6bfb39c3e7a1fc0340a
z94cce022ae89957ef080163ae7d85bd2648f081bcb39a544a86d4e6c8d7f9d98c70bbe0a26d719
z0b286c36cbd64003271876e2dfe5c668dc7654a472267b619a463abe05f8204b423b6f0df7a3cf
zbf50795fe6e47e864fd23b9198ff96fb5911a5005ccaf5539800d75e2fd7d4d1fad0ae277c2865
z01c0d89cf942d4856a8b59c4ff7f474f220b4f754f46e89c56f179c103aceb4a14ab6ca17108ce
ze38e40a46b4421cce1a7de6c3d57d0dc5c6ed0988c784e70ccced2161181ddb04aa19f2c6b7f69
zb13eb98c8af2efd05c3f0985f20a73c99809568188ad908a0efbd20b0fde2bf42d1a969b147e7e
z448fde1eae59ed410ce5887bed1ec38c3c5bc868568e160dc6aa5d2c3ffccc37c91ae9bbbc6c04
zdacf312addab56a79f2c26984fd38955eb5fb3e5e54301f2cbdfdb326a6d49e522aca861350895
zdff8201264175e9237d3136b0ee0d004903ccb7ab1d718244117346338cc3f90a0cd791905806a
zb01a6472062ef2cddeaffd40749c57992743934f677465b153d79c41a5d15ec3558dded7c5ae9e
z781b1fd986973c778a05df3b975c16eb7b4b907eae6fddf9bfd71b314a5dc380531f20b4d299cf
zc0fd679c91416589c0ee51061c2c9e18c13c56305678e4141ceb89084187e266e484fa460b52bf
zdbc81c2d5c277406b7098fcaba604623d4242d06c2bdf029795910c0a9b644546dd800648eb103
z71fbbff4acd3a4b2b2336c0991c42652d3c251d024ba05a5be0d78b29d581eefda8400980b51d7
z023c9d475011fef97452e10a6faa53214ed9921850556187c550ca47ec02f443e5fee4a5b1fc3d
z0d5e636be4d54cb1061d6524d55942d5d08186d5245917c229cf0b1a890ba1d000cb50d943770a
z8c163d32882b0fe7bc2ef007d25b1074c65d4b3c11fef99f5304d45399cbb096a9b1edbc5fd16c
z3994b50ed56df5c80013a2b8efebaace2f396c1a81241405d8ba81d593b7345c7320f8321d7989
z527d9ef0b8db09af265c93f76ebf57d2bcb8ceffb0292dde13b5b26bbe80239491908002624d9c
z1b5a1720706c503b9c520e2c03116b6b2061a2b8a1a2d25d720401b3b9dea2edf7c19d293dea15
z23b5a8572bdb27fa424b86661c6cb615f159b35cbcaeba5a78a45dd1d260697f5a3070b3d2ac27
z89bca433cc6415aff6e03bdb5586d281dbf9f0d3ef4e5a57762840aae21b8771a63fe3f147c82a
za960ee611f3f6214a79973bd0d715a083f8a9110ce313bf82a36f546b28b6027a009140f2a4913
z617c4d64db4249037ac41cad5a347ed29b62dd0f2b9f2ced234898e2e9395064a68e1b23ab16dc
zf8a3b0acd316402a5e2b6ac211682232eecef06380df0c0600753f75657eda957b1eab580250fc
ze18b99535c0d571cf93fc17c35cb56766718399be12e24e27867a2fd2379a675f42d0d05d9b849
z21045b3795c35913dad6f5319d96741085c4be3963c049664c2a72d789e097035ea864f324e432
z8abffc974a3509d2f3b358630adec390308ec1ef0554bd1e6becc1609dc82899659f9af450be3f
z2655bf7e7a31b7fc1e66ff50aa4710851ac30c0a58dcce243e21744ac1c8beb62cac9fa5a52128
zb5ad8c448b5428758e8f12879f6b00f7c42674f3af334b7e682c0307f937d0acbb282dda69efc9
zdd2e492a2a78e7c54fa81806e960debd71ba5770b7693c0fdd803c53b8cd301ae882c6b9c5bd64
z442de5e5250217ad62d79f3320028bd09fd1fc6b530e13b0c4a4af3bca1e341ba2d92fa3185197
z3a0ca137d5f7d7107726d19e9394eb3cb5446323918f16a2fdc9046b9d5149146da615a8f3ad5e
zce15db70713f414a06a130c0bcdbe05ee01666e958862c43b304632aa4ef4135cf8fdbd7cc8406
ze298b4ab61eaa9c875a25c46466689755fbfed0c06d1a79add9108f18f35e88e8c312154d2fe7b
zfccb7aefc4bffb06aa562f7371a1631be4fcf1e204c4bbf7f598c75fa22385b89ddc8471c06e3d
zc1fdc77a8a3312cd19ba926efe792d071c0f34cfc08b212c6d9452dc7a358615a911baf008c413
z53a57b571af1bb33072c390fffc8a19f0a4dd709b02e7c7399b7507a3c68bce4167891d5c89b5a
z024c3714a78ca7d6299b4da9a95fc2539dfd590160980379ef46457b1425ecf4632a833c5e6c2e
z10f84fb26748ae0c46a830848a7fce3a882b887b472b5a26d923b25a396f367c16bc74ee83c873
z3a3a95fcb4bf4d6d4394e647c5cc6e0f1c52a3171b7cbdc39aac1ade525ad4fe290435214c1b14
zf516a944885059d0df62085717e5aa735a9a35aeaa67175d6bf52bc49448bb6cf33f9fcc546b39
z950c97c15ba1e380f233fa5ffd58ba700b61893fa8db1144e7d3e87b5be97c7654753cc0511f49
z7a82bb0798b9fbee03d3aa76bd9ff651a266605b77f73936f7e053702b43144dfea4f7a8aa2a64
z3b1e8e0b05a892ec07eb37f2766ff06467b6a29d463fe2b99503e757a533c72c785287b40be9e6
z71caeb2a5d1138430fded76db529bcc0bcf43346b1800da7ceef0030b8e1ea3c1b550d92695b75
zfea9f26ad7745e16a1c413c7f52459da71dba52caf5d933f2b56624b5fb6a72f2e61418853421f
zee36799767dbdc722758a424fbf69d79400ee9738acf55249a7812a29f5eaefccc534f52bdfeec
z148fae6a1b598a1a14c5bba6387aa1a9c25f3f9a46072fcb004597b519f2df2c64304d1bbedac9
z86eacb23b0a709384e4a8c040d1a564c238a729ce36036dcdb2930a0a77df2e4824022604a3884
z587f64b046117d809f81b9e2a7c8b27a72d2fa96c3e3199bea46d0cfc888b1dbb6ba157b4405b8
z4a3e7ab167da45da2df96fa003c679468fbb8ce8f437b8af8137d2a89b2a012bcfcf0443677d73
z5eb44f3b55708a9a188188c292bde33709a431875443981abc17a0a9049d12f0b9e0cd731ccfe0
z277133e23c7696711381fe8add338faa83fc6562d007109d53319874feb65b277fcd08f6b60b64
z0315429fda5861ed5dbe66c93bcf2fa77c9b746b37cdf5b862f6f164c32c41fe966d2192fb0376
z95a2c28dff15e08090efeead05fc80159645b9dacc93d7d0185394f202440b1b541d663b06fd19
z37a1b72e120a8fac65d032ef249b74c41ef000039557f61f9e08bab8ad45fb5ef0d67b2bd05595
zfb669bcb99cba01bde00e9621c56cb33f3c78bcf194b940c045363a47fa16514ffdf81a02006a9
zd7007263169cd81adc53505ffc9185c01603fecdfba779a4100a6485ad30fbc647b50c4fd0709e
z9e3a3f7a77caaee2f8f38d02e75b68040f723f0c23ed6af3da4342764e86447a0525a9ca974889
zc81ae8bce15cfb3f820d75be68d8fce8fcf8e4f20c604bf7e47b59c89337d4c88a47b99bf3ced8
z8e0371e323b6294ee549eae7693b9496ff88a1f106f49a476530f72908da757bde8ce985c54124
z3b0d330a5225e21ad94ec790aa0863508e7b97b412052adaed5ca62a8be2367211631da47413b4
z45eb382aef33490172ea3d65b7dac70ac56a22ed66076a4dddb981d3549c87c859a0df19305ff6
z1eeeacef8ae58055964e92d9b59bc6654572745b96b1f0053d7300150416ef254820c1165df151
z324c10385efde1bfcb5ace72c26296d0d14ee12daa5ab639e74789c7f2a1b2b0aaa0d3b1a87552
z79190e779e8ba507d5b70986a025b51f67cb34b122fe66384692387ddd61af2f08c168d508a9c0
z244ca2d617448ef4269cad48c958bd88d1fdf9a8b9dc295099e2588f0317013b481b407f63fb52
z1690e79077c20fd27a46a3d0a314b38dfe57c36939a652638bf8f5e3b8016a577b41a1e2a9d770
z3ca4ed9533dce8bd1083b9b320bb7110924f6a85fb43eb2a93ae7bba5139a7e7e563b3a08e13d3
zdce233deab4b0b54ceb668460a9af8ab487a32fd23baa54c978ecb00343f9c51c601a91db9ed80
za80f1404d10b943ceb8de69fe394e6f7ffc6fbc1164a3b983e47d55a60cd93d7eadcf34cbabaa1
zaad322642d6dd97e8c7ef698842dcaf5daa3ad79b0f1817aff848ca33a20fd20c779cb646ae4e2
zcc9907a1b752005e3d06eda022bf8316899262213c5ac461166d45c1b8c0ad0af879d14d785333
zd4447e4ff4b4dfa695bfbac4e82a590ea05cdbd2beb6a424e6da2ab3fe2fc74b0cf18ad1f1a7c1
z5b09ad91bdb6380640356ceb18d8b25cdf8808b5ce2dc79d37bea1cbeea5c48fff466bc949040f
zaaddc1559890d1e06db0ed4afe165b2d699ea2ac08705c4e8d0db0bd805aad0f0ca76dd0a237f9
z4c941ef2e0b59a0fb8c9ad5ab788c9ef49d6e562e7abfc84a80b19d799fc82a87bf5a889e8420f
zfc3700c1f530c1426b0b275d1d30f8b48162684b86c3daa99f517fabb157f9b9360a21953777d7
z1a2df6f0613374be923e567f08c1535abe6891e5e09b1457a5c8415040058de631b932a5a6f44c
zf326c32d1a8b517aaec9be158d203c5b7b5645dae4e6cad250dd699670649d7d945da9ea5f8aa1
zc38a17ccb36e4f6528197c1025d3560e01a6adad5e102b460ca385f3208fda80ee923949744780
zeb4ae8278d24a7d2d75cc0010e24f08478ed21d1f38f72c4136fbe706370fddf5a7bb24c60db0a
zb49a9845971e30faa3f077bcd40e487973a01f1316327d43b51dee300eef1b937a45bc1e946d3d
z297172696b77d01781a43a99552462d04b988f38348694931f7441424ede7b288647c73db13849
zfca4cd71eb6172ca09a25d7a36701e2c198df89dd4ac58864659747c71d8392ad19c087aac1b13
zd51e290dcfe970d9f4322aefd9f8c1a7d5a652c5aead1c4395f64d0247168577e4b26535665633
zcdc7ecb6301eb0dff8392a892cd7e7374d11131cc24c9f0e5d1630c9b1cfc9784f1be55e7d90e8
z025d796e3636c85b6fea8bf7dbd360d3a5dd625b3a1defe44e81a0cca18dc311e54917296e01ed
zb9059ae9507ccda0b8773d985c13beccd28e36f92f0e564e09332f520b5388980a8755c5f22213
z55d1973df85bc3efff38080db88902318cfc01a54e9f1bc38215d8ba5b1655af29257fa4b626b3
z0c34179eacf762365ff7a22641b68650f7e9d4f5db859eb73458cfe664743b10b2fdd7f7b66291
z5da67185d95edbd6b9453cf424867be3ee19c4c9dd758aa861f6a56b6e7de55d1fbbab9d8a9146
z955db6f86986680f34a56538280cc56bc6eaaa5ae21c732dedeea2464c3bbd4dcde85da2357d77
zb80486a78eb993709194871eb71efad8609b624591c969f08ea0c1ede35692d1ad3e9feb90e995
z10287668efa4323d957f8a8bf20f1795a545d39f43f0e0f8900a70146ea440646bd66a399e2f0a
z98801544ec02d607448d21ca89f42b907c2ebdebdd3c317e73acf62ebef7fd6c6e95052d35baba
z60a0ef612e3c280c55a97c3cece76ee649ed987a8f94d7095dfc384c7c1c805732fcf1c9f75d3e
z2eaf391a0f0091256e8bb68d22575e969fedfa0cae2a51125d6556c1c6c2d49a318f1d1f9a8fbd
z51270795fd79e533476809368cbaba77a75c37eac39c09a755eab844549878129f16d9c4153641
z1f0f011b65fd44a9f2aac49f3654b581d0aafff3bd8c60f35583e0416727d96af903625363c226
z5fc3faae6820df4c6791fb44297e622cabad05316aa3aa247737bef8284fb81be83ef700246235
ze3eb807e383c23d69f22b3fc9323cb8ee8f6e1e4f0aa8895964680e6176d5bc7248d55bf6de752
zbb1c562283d774c7ca03bc6d83e9419d77a4cf81a1a671a7a5643bda066f9c5a2e622b055bbd00
zee5633be196c885631f7c26f4b2c694093df65c6153b92b51e5320aa33cc850edbf709d4317868
z9948dc300fb4b531062d259cfdbe3d9122a7696a2a66342c69ca0f23e0faf59c96bb5438ba3396
z08086e5f18dc7d0d46147d1b554371c92e8f9abbbac1ea9721b1b671182450e86be733b26f170d
z8793928d0612bdb9c74d194a5440ddbc84ae51f6a25a37adc3e9a65fa7aaaae7db1b267227d39f
z6b83865f9eec8131d71e5bf7a0c8bd28a992ca13276c7ea9233df94b2a8e0e0a9e9f32b2d546d3
ze8891d3de42e8282573989891117c548ad4d6996a7670ad1db11156c333d32021abb1600ab8f5d
z86ef50808630f96fc81f0a5c87733c5e41c5da00d1e80dc2b20c65debc0e342612ad6b630fac42
z64a64cd54c05db6dc3006ad7d13a2d00ad6b096d6a65a2d8590397491c08aed5276b8f31e20ca9
z89908bf513efd90a5aee33a6149f41af4708f26a854635cfa6803ea5591eef9449cf002402fe6a
z5fdd946b86553bed329a3f97613c06ee08e54dc7b5ac145a67ff4e7bda9c41df7c1684d01d3666
z258415dd6ac623dd400b8556faf1569a68b3c59d3dee5781a33d82440d928c3cfea010b6a77fc4
z96ad2ae12a0b1b6c785e05ac2f9b094511c88345a99640e8f7c45da698ae509ce1f8caf9d0d7c2
zd78790c381061e61369cd8729c8cbb363da565a911e19e3f014a6670db484752ef181640e38113
z2ec2b17df49a6c0204eb5002e49ca493b205b0b966ccf8e02f49c4b77f9712e75869acba8fe5f6
z6c6788f0d71bddd92d92799e20d37beb9b1c36636cdfdd0c69a8c07acaf4b5b7171e1c1552b3ed
z73f90bf7b85b24f2c3ddbaf3867c78904cef22a0d6939354f11cd594022f03690a6dac58259b5d
z73a5640f6194befa491533165431d84fc748907ea7c38ea8e4eeac310abbef041d1ac5ff59ae2a
z641efaea10347bc64c655ad966ea9beb074f8123bf5e8201d55c2749502ad8cc45963c16714065
z13423186d532b14bf1b65866bc262378fd9afb4dbce47e5a961231072c68f46e1e4d62d3ded07f
zab1a2b02b62e0d78198fad84203647c4f9b30c6b26e70fc68f9c36e29c8ffdc80f96d120dc3e97
zb87dd45b02c3e68ab6b66df60ba88e2debf8eeb0fb64153a274611631e01c9667504758cbda6a7
z016fcff4cb389b81f936ed5c6505920371274dd0d9bf1d8ff299ed43e092599c0cf849cd83cabc
z5fab310c2fb78635ebfd701628bd94339c64063bcf4aad0b0e97f980fb1f68108e8a91e8833f69
zf334f85a79c2f1ab18912c49e2c249b52bf0edbac8c97e734833b45a2c5f3b801e00fa9d3fe178
zb9a8852881c32cafc374260997dd11f1caa4ee541009b23d8e138e9812b9bf136f58b7ba53b893
zcab35f5f6b4c5781f36e8dfe830e0de9720167229f480435b14cfe1184ef1c6590a0365a78f978
z4b08cc30d0b08694018689bb5af2f6e1bfce19ae522ea6a7a3a7985af6cac60bc8826f91053986
z9760c7e90d7956d743a19243774198c0625ca6b33de94f48e4f18b30e783386aa9910ff98c7dbd
zc875f9f332a3bd2630af77d4af8c16df8889961a7cd65f3d1c09c2a269810da74005d21cbf1f84
z6e4ef6d085ced7244b8498f4477d0a7f30734be2584d215b596c069de1817d15bf6bfcae4871cc
zd6096f56505bbca8ca89ce9126d0d9b674bc9615b05ef3b675dadeadf743c544219db0e66df98d
zc7fe0754e06fe54f76cb91f9e1dd2cfb0fe054998b77b2fce5af623ea68414dfabe04e910bce03
z95b107350739a804c6a4439056d9f4e4fcdccbe75e91ff2be34ac9d5aa9683e309b972be5ad678
zef66b2598faba713e20b9f8c056052bcd4bffc1ee658bb3c8aee75a46739d53e196173c3c549d5
zc4b6ee434a3213474fb1a27df2f5e95068b4305b578ba5991edcdebd7179bc30fffc58e923f209
zcb905c8db45165cca95fc5a0caaeb8d4961b747dfae7dfb67b0e9d4c9932b7a06f6476cf674a55
z448ae85f9aac9d753dd45772d54ae0c254b2cb6b5189572b80dd595e6d34f53ff4a4ba393a9f2d
z9ae2da8fc783ddf9a597f8bc7ded3a6ab8277432b84532f42d902edce5bef9b9336514029c0f87
z9a26e7f8aaad306653cdeee3c3b2560bd48c867ddb12d34d9355f63a7bba0ac813a164ba6460ba
z44c641626a66f8363d3735d325c58507274b412533f115fb2a4c19d5f7a73a931e7d191ee9f0f3
z4e33c15a828548cd254474808d70f2f1f7e55f168325d06d06277ef0833f6d5ef8a2159cc1dfd7
za45c4141d65dc6f469e89c7dba3b5ec5585a6195d377b68a0304bdecb6fd232f5ccea7d4962ec5
zda62bdba56d12f401bb0eeb9a54fd7495f991e626eb5540e2bed59ee2de4de6ac26d7d71797b54
z8cbd024a8ecd7feb210cde10305f1d9c48755cdb8ec62e3377dbc8b0b8e1cd6ced49cd99c92bb5
z0523e9b03fb4178998e88a0493da0f84b1d495cd01289f7ab5e16e2d3957edade39efe372aa119
z7083ef9fa88bd28d0d245116b571fe5a83055b73b8495f362d189476eae1eb11d5722b329b5054
z68465263353ecfa4ad137c6756f88c65d0402d92f9b40dddd664a1185ced220ae2e815d4eea955
zeb10f80efe1e9e56ddf25537a70411ec3e63ce1564bf4e3d974d5f3268919d21796f2d25c066be
zd9feec4786bf9fbcddd3092aef46fa1df54c8c5647181789fefdc3b249af00448559170857b5a7
z726557d82723f9ac722fb5c90a80bd08140154a0e9d8c025fc098bed1aee5f2ebd0883616b90c5
zedf98aabfcd0a901fc7f46be8159f1a20f173510147907691e423b6f64286f86eecf0fc8f413e0
zd69b4831e528787fee83b476cfa116549165abced0a60d1b2313aa005d1e3e35bfdbb246ddc02c
z38ea40b7de9de7017bd0bc8c3c6c591807f9839a177ac6282662e7096b3d5da50b2ecbff80f011
z806b854598ded834b42f75caa765a8f3666c90a6737b7ea54bdd6884c7a8a155a49a04b2d17236
ze38491adbf7a7b5a69c7bd3cd20e159d6ec96745fae4393e5581f10cdda8d0a046b31f47a77152
zd64c6ba3c949b75d30d9dffe46c2846a4f6a6147625c5dccb154fc095d9d8a94963c310522de2e
z5632218a10cb9dd4682964bc52885699b11f8eb7a1e3e02026e3d54f16090fe77af8db4aeb7e6b
zf86d69490fcb3640415bd9a986392a7cef63e1822a1616639080ccdbfcd1c2e3a74b840643b841
z726259a6b9fc0e13afbbb5ef8ac76276255c7afacf37b5b7607b22cb2f4cc6cec6d7654402aa6a
z2879228b4949e748ce1dccd17d3515fde051fe07b17abb7895369394ae8f6d68d7212676d638ee
z5053259bebabbd43bb0c41cc9616ba9b200a9027e1f568b0da3069f98d5e0dc050d1f6f964e4df
zc90f021e53b2e9e411e75bdee4c61ced9d8a63ced487036581acd311d9d99ede846bc6d42894c4
zfad1c26d5cae165732c053ccfe469419a9dea0e1864724f69a59d3c0f5d6177fd7e049c2906bd2
z3fa0840144da103be8754cac08dbff823b54189a3b3eb6ed05d43e6ba5266fd7e856585142b73f
z70f59c2189455f8bb9af09b2ea8a3516a42f2efb9a5217ac58e79e870bd80eda2cc42c0c8115d7
z1468685037b4d97ac59b0af8f1ddb507432770cd5184bd08659840344233eb7cfbecfcf8807355
z078699d2809af96c20ab29b867f440990e953afb0ffc068eb4f22e909b56b0ebfae055afec53a0
z71ca9625c2ff592b232547ad3839aa7872c1914e5ad3c6dcc0854a3e4febf6954be8eb97f8753b
z8e9973942a63eb81a18216fdb167f59339a9b8596d43818f59b24a5e1b470722ef5646e3692254
z3eb16aea8e1bd97cadfc8d0a7e22e37befb21ac3e5978d957a99826aaafd53788b9251909a1a3c
zcd0c5aed08a7c6e8d03c1cd2e24fb0e860f566be9085b6b409ac73d34384ab7308d2af04552917
zc21aa5322cc06402db371e86ac107fa56317492e30e1afcd7cdb409c08257ba44adf965f2dbd06
zf00a020d9f95ecfb8a1c061b9dda5d60e688713ae3bf57bfa24296cbe221dad87e48cce3403b13
z885cbe1c25fa07e62d643d36dd65ee577835cdfd6d601ac05e65ffd626ec9c88ebe5e1fe927e23
zfebf16da50b3b9284c8b689aaf753cc335c04d8070f10df097632009fdaff2ec4ac72f7a6b0350
z38e3d049bb0f9bb167771c586122058873d013f8836d6251f4fa3b1dea0c3849261b000e0d9fb9
zd3fbd9aa25bbbba5424767d4c887b41b75a1a055e6c0fa0942edc797058097c3026ce0b3e67522
z0f04714ffddc9d0e977fbf06b6d87816cc36397dc1ff99e938cc08fea2c00e3617351db415e352
z533f2b76947560598b26b15822ded0f4fab3e063a11534cd74822c53b45638982b7e108a8a987c
z06ed9c5292b90ef1f22113a91aaf2b310170c7d025d15a7f230a02673dad53b7273097846e4a95
zc25a2c97f0b4a64693044fc9eea63d3749cdf2345b5732945dccad56c9c55c86109c4be060354d
z7f111426e83eb110cf95b2fc68aabaf10f4d8623a3dcefb6e4978a9f40c4d2a404da0f09373644
z28859ea92a1cf72d014e534cd5a4efe7fd30357dd97efd15f71e43a22505c248fddd53f888b4fa
z309fc7299fcefdab88814b51acf8fab360dcb6689f04a0e4e7e8ae3204d8780bd4f6c54537140d
z6c49a27eaff85644a54bb4fcee05ccee5d58e07e3e2bf3103e8d35c042e4b7a9ce728524ccca1e
z260c926f6e7657b2cf281f813d2a3a071e144f9008d40d6c49729620d876b6a04cd421943959e8
zc6dab316abc0dc66e3ede068a541b59ad2738d928eaeae8969dd278a0b7f82e99102bcb057e4a3
z00d87d4469c005e99314f2dfc16d451048d54b3825b9a301a434698048b79b078d817f18acb674
z4d6866b386a9fbc1ec1239bbfcdecaa68ae8ebbf75582d42da5fbd86bb4e95d244c003c15d5b24
z50ff1a4a7b0c9c32932bcee6426a167b8ee5fe8ab320c844df93903cf547b234dbea13c08840f5
za9ccf6b69652d0e663598a38f0d9eee625afd0738e666028aa1eb3d59db91ea35ea8ce62aaa99f
zfeb38eda710546b899eb6347e8735224595fc64117fd965702d84db03e8173dcbac54246561295
z8cda26eb72fc8d6573c3be9f073df9f280f88c2d519778457f850db21692b270b211fa8fd0ec26
z339fe5a066a33b1dc9205788b81d690b7cc5d215614ed1b1de8a3088a6b671e1985c6533eafef0
z6bb6be6a40a399980dd55a37633d07b54f6d4b99a293d3036f3a600d0ac7e5c38edd2d8e29d194
z2a535c13a2a21968b81c8180bd5414b53e2912ece81d06dacf0b2e21f642171fa4f1a3a93ecb8d
z9f4de92695ae89ee25b3230f3913100046fcfb4651233d849608e1d5d5111c9d5292f48c0f2193
z459c4b41bb04d0e1c19cc1ae3b23e4363795f46e3e8152fe37619f03be9fcc030d0ef8443ce190
z1eb17fe9df51cca807f2be6a056e2fa205eed04d4184977e0e08a23b823be83293ae65896a7ac2
z3083d4748b9112a0eccbff5dde59b119f6d3989244afca3a0c6c3ce7056a56b1ba6b77ac969e5e
z2b0806ed5c49417f2d6ea40581ec52426bc0ac37ce9e6a5cfa595fdf1e4d07fac0f8bc754a552a
z66a6abd3def2a06728051b16564e4655afd9bb0daad38aa290574efd830f62f86e991a3a29e9e5
zd6518743a493e36bba3e5227165529e91398808c13a4d62134a065b7ae7f50cad9104e9d8d4e3d
z8ed6f89e4bab91aa11dc90bd01c1feba7d85434bd2d00e0594f11214acc2d79bbaf63f9036a316
zb9f5056834c23b5eeedc91c0bacb0f2b6c2bc46ec9e7a0d266738c01be251b320018c9375a6cb0
z58f41ae12f3ebd8ff615b7876b3cb283198b26a9635b9266e28d36ba6f54e3709e96191e3fae05
zc0a1e7e43d9aca19e98cc18ce6b56f8e4153b187c2db5dcf04ed7839daa900ae044dd47ada31d9
z490c99ff17c11f2560464ec4024bcd8fed3286477baaa9534de1a0e0a8d3e703dadc4476da7d7a
zbc3d042f8364703adfd785c9d208003472eed19abc0211d7f67ae268d669dba0428fdfd0269374
z619b30316e4082c7a6d09cd55b213289fee8d9ef74b1f0405f175abe34baf7aa5fa25336f7cd50
z8e4ef1c3191f4b9e83604cd596f0f5457a52ed10312e7a220f2318e43d575aa71bc18a9b616a24
zeaf3914937fcc63a83cf9b35524c31c501924dab541dbb9008feb596cc14fe66d3498301180481
ze0c30f6e94e2598347a1b9b616671ce7aa9d148e8331684fc25e7dfa0a9d3c7b69ace6875b43f1
z90591e1efcf784840911838fc5e2394160a0b7f36d1dd7fb12576d7a067d166759cca72f3f0056
z8dcf1cc1ea3d39c72c7e22acbcc6e361403413f405193b4106e4a9572ad2b18d36efc8891b2901
zded68d43bbfe932316ed1a13e1b84711827f5c1884670d09de5852d3f01bcd07a8b975939201b7
z7784496753d80be1fb545c661130be506f528456ab5df2cfbdaac6a64ef3226f5147b17de0404a
z4baf7e7f4debf1111583298ebc591bf446afffb456b4a1be3509ed7b3b1a6990d9f748693f92f0
z72bbad92eff91d52f9b4fe09604836a20e10bce64bdc516c5398aaa08d7d6b097cfdc41557231a
zdfb2ca6085daf61d84626c1210e265982d4ee1e7cae2270b0de06aa5b7c65554a6c7d75d7ee3d6
ze868869145c1b6b9088da200b3c18a663ce8626fb0001ba45da9cf43a25ce1a45219fd0a34cc66
zd744db6c4f2caa912b62960bfd29f813d08e421ad9c062a3231bfc9807c8a4596006b5a4d19e6d
zcf10b2283a9b76fd12324f7a8943322dad743fe0dcfbb780f83cae461871a1e9d31af654489a3d
zf266f5bf0f5993bc2e2c53745488b97976874af022fce546b81e33ccdcf6a96c862f310da796b4
z9cd946ddf3e2b3cb989b6157a18624c7c0b646d3f8cb44189bce63912bf1fc849d11cb118a7c4b
z881dae8288d8835b873bdf6dc7c9c03c9692ccc516a8ffc6e1aacb5a9ea86fb27808a205f8e22f
zcfadacb9ce3c02ec01f94e494f4c1fca23ca2dacde3986487acd46e06fcbad582a6d74ca7847ac
zaa0124256f7e0428e0fe78f29b35a579a9ebdbcddf549be799e6805c7d1cc42391b1035e0ba0dd
z8fafb7d65c9e79a78fc6ab1398a6aa1326dab7559a173d64e7f6ec34fd8c52a402aa5399121f49
zc531eb4f95b7b57f47f7ebd5ac7963bd725c0409ca5d5d40f3e19da9f4f1fda6269c20d77ac2c6
z94cbf90859de4b01f33cbb7887cf97310755bf20acb4aa174adcd5f4b623e14c7926b0227763a1
z082abf84c0ba5c11844b85bd557dff7e5bd15375fc021ea6d92a917a26db2b33e6269374c34763
zaafff08f25fb2fd7d72956ed2746ab0e996c901726ecd061e2700ba9baf6a3cc4848801f507d5e
z88564271a049afa18b78d74bfab333edb214894d86937304a3b770b6a24661bc1367b16b6247a2
zdffe75320e9fc48378fe21379c957d0b6afdae5d582440b5b4dfe48491c5441c6d0b13918d15a9
z43bd1a3c8ef5ff9897e350297b70aa65ac531264f5bad4431e0aae36d3fa8d81fa37df276f7b9f
zbe81baf39df550e369f2f568f7719cee9027c4ec4f8a928c330ac32c168a8176da9a2dd82ed244
zd58cb9b631b30bac10aa3142e691b3c09c6523108249b3e1c59db63a813b0f75d2a4d4aa10711c
z9ef9261e8a05adf24647c6c56aab6c3081117582f52f993bd3b496107f5cdb4202c507bd4bccf6
z2106f8941354825e3307f98bb558819ea43f0810c626b935ab27a16295d10a92481ffb6246e07e
z18fb5ce65cfc25b9ca6ae42d8164f267ce8966cc85eaa584ef062cd95c479181d495a36db07e18
zc783c18eb0cb974618ac2b9e37113c2e76b34ba3705b7a69b7eeb8ea9c2b638f18a36ad2dda229
zd2e149cbcec9619999322ee3136d5e20579c02785eb6f44ed3dbe95da3680e58ac867c0736a413
zceda5ab127e522a54fc5ddbcf0b756def72cfa3d6c22310575444cfb72a5f9a0f9f36175ca3612
z8d966cc8f49323bcc3617d4d145e0ae3d80e81f386a76b46f18ba241d7bc7f7f80394327fbd9d2
zfe40f3001fbceec87badd20668e7846b97ff4d1c4fca6afc1d11cd508f5f2af871bec46a7dc952
zcd0c0934d724ca3d0737cc4fd08c79ef69ea01b69c5411eb6ac98c1266a8a1324a0d9908aae551
z02b3da4f6ac4afb508425235d9bd67e2e3f586511743e42591e3e352bc6cf90720dc44d7d48cc9
z7941929e2ff4ca6c3ed94f20d958db937d924f88ee60858b85b3523a07ca4c81ae5ba62dcdc93c
zcdc6f4e02bbba780124cfcf7c483d7601a8a4fb858971fb564007b2126c0abc8dbfd720cbce3dc
z2d5d72eadda4f8bb6d30e711a99f5870973f2ff592c53cc2bf3768d7e3ab3e898a231cdd09b554
zfe2e512bd6fcea9f8e95455c4d0d525ff4818fd79e8ef0b32466b2cbd75889e0a8c9d4c37d32b4
zf2d7cf518b9ff75461f39b06f4e3f86b17a6d03a5662d319f815314f2f7f7545bee000342b2720
zf98ec537b72a0597efbf23b6ae444153da1fa0cf018d967e20e1b286a08e10aaf963a2083e3aef
z020f0f4c7aabb69dc2bb9dfd15e9dc616735c6effeaa8e65dbc248b151e19a456900cc68bf8103
z75c386ed11b661b8c84c8656b80ff50a49fb1648b560abc27b59376e33fbc82ca75ea246bc52ec
zf43200111bdd39bbfa0ea51590bf64cc54d387b6388154811b38834f42862381a1e798e467e8a2
z39e581f4e7d1f1b99af24777472bdf3506e178a8fda18ed30666d96aeed76dabbe6cc3d68b7736
zb92bfdd36de8ec118338944c9352144e09fa4144474155dee4e3d1e4509eb4fc251362562011f8
zd94087feee73d16014341d11f087ec72cbeab786fad12522b1f46f07e544c8cc9ae5fba4888057
z754160b94276aa9261420ecde3efb6e8e77982d41458d8b1694140204bf664f04dc55084b59ea7
z33d12fe82ec6a5e8ddfe698eb4c32d8cd0c32cb2b6f63175fcbc6c032e0323ee4c21f0ca0ee3db
z259d4c3edc8c8bbbbabf7c579285b8ec7a9cc12632af73cc9949ecf5ef00d476964261c42670be
z50758625256353ff46ec184f70f8d9999640162bdce6832cff4882166ddb2e36ae643d3403744a
z70507de3409f75f478365177b3ab615045336c8768cd57424470c6b7411847e42637f170d770f1
zb94ff09e7d07d4ac5dcf89daa595c5698dfcfa8dea1123e9ce1a9a9c30deae20457ad66d893f83
zac8005ad3ba152a48091963752968f829bc521e0cc079bea47040c8ee2a8d45f81cc3a0ea93d37
zb53b56bcce73b55f798e0b50081f2fed94d41d271d2ec22a25ab5161baa240db30baf99fcc662f
z5fd3721265471711c1d177e26463ccabfcd545cf5a501efac77e855253b9ca84523fbca2a593d3
zc3bde2ac375549c7878348b7b5bd5e4b3f224083e3e87e96fef6553d033aa70094127c738a8d19
z935ba31b0c22af71c38b80e293f5512a27b30b182d64a1813aa3d8936036effb009ad09727c410
zd7142c6a6b88e2312f62a0f70fe812d2c028a7e24b788ec40ce5f047f614542bdbd47e8349178e
z90a13ef8561c9bc9561f10932f7a3dcb9fcde3a084b866d0b4839c984487ee0ca2fca757d1e67e
zeb84a3aab4b39110377286f1a4343868b8e0e2e9fffd246cfe9514c47e3134c477c910fb12595a
z461535e2233d584bf34136ec7a8809bdc68dc3678f6a6da7b6b0d48827d5a5ca8f136695689dae
zc330bc0dbe9572f165738137379749789e2c787d1f68d7b3e86346dfab702cef22b394d7d51701
za4aeac140186087765f99831fe879aaf6802b86544f3db854a87e7c64d4418c4e904e2410bf326
zb41c7cbbedccff245eea8b4c0b25b449360b5544d7723c56683d5ce572bcbbbd8369c1ecde407f
zc4cf3a347ad01f50a7f897a3561fb8401887cb3f7de1da0e0bc22fa3c2f0729632477194985c05
zb8a7a03d2df788b8f17634d841a0b5e337929a4547d3ebeec200d3fa8e0cf5992d9a3980afb895
z85c15ea3858233451c1cbffd41aa1d401beccfedc88f1acc0f6687683e109669c3bacc5a757429
z8d075fdcb9fdaa746d3bab8b984f5309562ab4c1419efe5461b79303705a814bc9cf57e9068d68
z349e7e79e95fea0ec1091e3ab7cdf27f2412c0b317643e50b5f89b9d074f56073224398534b762
z7542af240ae96e1d73785661ac1713285d501fe34985fd5e2c9a594833ac8c24dd94ac7d1a8915
z07ffbea59f13196f859bc9a7a4c8fd7963fc62bc0c3bb44aef672646dc9dab7d815e574e2dbfbb
zd870c989209b17a6d5aa707a4508c3e73754a1e47a4223567140259cf65dc77158cc3f5cb3b8a0
z61c977e7819e2db0d87876f8b7943cb6f794b68ee38db323fb45f180fe16fedb420664a7494e52
zee4427cc43722466fbaf2f9a31249efb1012b4d11874717e7f707d0dab5367bdd5fa7c272259e9
zf3c86978a241d6020a38b3c6f935e2fc5b2968f88bd945c809c0c797ed649756d0bc561512148f
z4a59b9a7e83c155cb1c61672c3492fbcd3d126560339e4ea14c8b8f0bb0e2ad3a021548174330a
z7d3b0a8ce2c7461e6d17d6d18bc9cf57a4c2f023a51068e8ba46371769503a5a24996c36d0aebb
z9791143567a2d612e63d723ed0ee7583823472f369ca31c3a931ff98e887c30e0e699c8550b863
z61b6fcd49db780e9413b2eabc0428bee06ed6559cd3b5fdc552c6274791d1efd1789102d723ac3
zb5637a3d80d14795070c7c2fc6eee6dee9031abdc538d12c22a83d4206bf77e33edfd5851b5f4b
zed22d6981fbe33a8d96b4f6a4e896d9066ec35c10d83ce376297ee1aff86b7efd51e0e947c5a64
z8cb09f8464914c9f98b2f44c71d46e218318be76a57d0bcc0caf6d9d509567f8b196254c53a6cf
z37e2016abd46b138bdfd6faf201ab029ecd3dcda2a886389f0e1b2a5a0c55b0ef9f48a51d886e5
z82bc5ff8f31bd4fc39da5a4b04cb9965f4d374c28f63916e610f341218cf38db57e947fd612056
z5af57f678269113502dd88e8140a5b688974d465d088a800c30354a46c30cf88ba9e0a507077e8
ze4dc19efacdbecca332765fc90f60d13586280d9c96d7c280627af04fbac549b682205f3f7c44d
z57a5247bec6f7fd0e671cdf43bdcf85365697f7ce70806d36132e2341b24be690acb6056c23e23
zced786fc6efd722665ed538f35bc9c3960408dc57f797bda27267626dfdc08f55dbdefc3d26b8d
z7ed456c74df852a12b471de7e6652203dd63f0ad4de0edbf12d1da8bcd4fa19d8e1c023c08728c
zf02e002f3a89ae274134fdc1cb35185f356872a3cd66a2411c0e6ce68d3a80b6da847cfc2e5bfa
z6ac199e5abdddcf84f3b18e92c9cef29ba756836b99f4c61c353450959b7f56966255ab8842acb
z00eb5a53e540a72798ab1b86a07fc96a9eb9d7c45d0490c7a64c9d0fd1de1687ce60b4e243911b
z45abef499aafb9b8d47756e93666786dc485d3e5378c59690004f3180ebe3b8eebdd779a2d81eb
zcad0ee427e4da5c42171c29ede85962d5f6b637cb1fdfe8f9ba0253b4c4394ac08a164d71e8808
z179313ca98656a9ed293ca173fa42a11a42d11a6f55ed2733f00a087b2351145037127b3b5fd3f
z931f9e897d81ce747821c09d3ddd3c48e6cb14f2037a6e6f481b77b871c0d8ac8cd818d81fc3aa
zb739942382e5c430d6458fc6de4ac1602011286e740c9685a480480b47c13c23af7083d3eb5b8d
z5ec5daea4ac10a10cb96ee4c60a5da0612a64ff305634f168f3e1ae9de1750e6cbd99327afa4c5
z0bdddc7199874bdc041e0eace309bb5104e5915dd8fee1da5e1204191b964e4d43f71e25e8f27f
z94e2394e371f2db53d69a89a67e4115bd78eb82682a33b32b87b5cd653d8ef52211267d9737386
zd0294935e1e9db79d8a975332c8ca4aa5824c78fb75fb49c009d6628a0dcd06a917a5d71358ba8
z93f88f29f7476bb21910106f66937eca9563e38a22fb97082ed3c773bb4987940591ab38708377
z09dd0e79d585eb779a21b2336e7f7b2e4ce06c23ee22aba5e248e1a2ce70c2fe64b64215ea0bf2
z44eb89f3a32087b78004c65708c202b6fde9bdeb194c61885ec62a706fac7f4f24f0e941791c67
zcebeb197acf2389380d90e340ab8ea8297264d81cb94ed3a3a9e97a49735b659b5127d5dc6a095
zadb27e3f461b9dd8156a281f26712863f610d6d39739f8aebb1f502da2e7270ea5eafb3b763bd3
z947e529110154eb539489684c9b9dbb25a8c295fb1860d11bb80d03f3ad242f15b91d9e46504fa
z2a9e3deb437e5fa2d91f503fb97d082500cad0ea1d67ac0731776fef5c7fa45168cc4accce0861
z076707045d0c0a4b40849cff93521293c5c89f339987b126a43e45f455e76ea0e6c68eba9b1aa5
zce762ca080573e23a7c8150d80663c1cebf2b3d1e1cf41e9e6933d39d588d01bfcd42382bdc197
zb3a1b5dbf7178edcc3a66e4063e6d7c44c7e2faefa761463717f8b025a2ef1c563d1309c5aa1ad
z257bf5db9a4569a4b95c0f48a26636a7ac4a3661c1c268fbc3042c35f0097e7c9d0bd78371592d
z1694b6b96a517a15f69f1cf852b3cd4984a74e2f959d3c82e9f08252c9169fd21c75609a8298c3
z0ef09ddc2747288ea3a51a53a18d171470f9766ab4f76cf855d2c07a3653a1518022a5a897bc1a
z9eaf68508be7ca85b4c92b4b647b40ccc29d4d53e3ad7c70aac64bcb2cbb7de6ea4672dde4edf3
z1b3ca01627c1bbe82a41fbddbdcbf68bc151d55e1e02ede1de2d4d0d87ce8482287a3c04f606c7
zfd23986d3f54a5f291933211506fffaaadda6c8a82099ec36bb7968f3bb4aee8e0340f1a31c09b
z270f8115c7c65f55f404ac48a40e4c89cd59e82fbdacea62f45778b1edf0395a45301ddfa431b8
z7aeb3abe58192b9fe562c29998f93d5e767d5af08682d886d8f2e78d23f5d1164e76883d1395f0
z8b4f4f5090168de6779c63e8247e3db7f67a906774657bb4e5e9adb6de31834f18da0381dd68a5
zc565ea4796464acdc6f3d4c147ad4f9acd097f937e875fab7eb4d283f1951a91d37fa12bb38321
z7f6ad4be6b80097c119c34f3bfdc6fee4ce8d1fce5db45d2aa4a4e5fc87bcfee83df9b66703825
z4e5a2c14fe2b1032bab0c18e1c4ccd83a406c59a607b4142c4c9d29dc396d25ec16da9152fcb10
ze5bf690fdc639e1e46977110df2adde122f1959120b189d763abf452bcd2c2f98803ee24d4c964
z5ee419190d30aca89b47bf5ed50252f1a6580d4c008b4a88d6965b9454ae952f82dc20331302b4
z734bf647645f4d384559f3ef191f896077e5d00531b0154b73c3dca29591d8b17a6766980ef166
z3f3e1a3c614cd9a291ec6d1b1bd9a6cdb7b477e9cc92c09b1a1e079db6119df5c451afdbf57952
zd4cd1088b1b10030e917247d34876e37622a15a00608d033f5fd57404aa81b816537fed544cc99
za91125f7b5bdf5aa6e7c55358b2d2d71bf35642108979d34fa57078eeaac55a9a6830dac93ebc2
z6c681fba13f90e0940308f1df9295e7225062c105c3fcbf1271da3caebba54b013de23265f0a76
z33fe06a35fc2124c6b7002238f42674bbb341f38f1883ad894575679490f44e59a1cae0103def0
zd0a5c900dd33d9f7abe4018bb2ad0a5c1d7deff72b136ca265805713d33f100a33b036d173899b
z9af8cca4ac1ce3715e0422012d4d6df1c5abd0cb65c78aa2ab36b1c0a9b785d251cb9fb92c5c53
z2e102df0c627cf97f99930f283f1336ee4c3d5468b821f8bd811ce5e6ba9f65a9c2ed143172409
z7d34484f1870db0ac7e6853eef234d17e4ecd37eb538978b3f1be5add0c5274e92370860325eeb
z8ded928b9dcd9f7289d2472dbe42d14a3e0b89ee5546dd96481d19a5fbc14542e2377de9e712ea
za4cf85a6df77fec3d8269dcd799cf201d87e7eb7b9aefab29a418829a192de8a240c42abc65ec7
z3f54f44b3a67143250e83685b498a8dac0c21681976701865816e88e11b3e15b46c01ab194f494
zea9d729f2ef7f4b2ea1347e9bab3ea58bad2ee89a8c66843268b76258965a30be58ad702811b51
z75083a9b789ce4f30c26d7deb8844f5c0b896c5213097d53a5c1df46841f78786fde10b469442b
z9a94d750d3b1d674d2d6aa2bc1fdfc97d31463c91e114bf5ed34c712e535be270f4190fc06b640
zbd6e7c322deea5cd4390fc011716c105fe51b9a98b5fc0767a4689b2e2d17d035fb294ef5f87b6
ze4372b60b480f6f2e937551e66653c8522d7e4375c39efd4168d7fc744e5f76cd090f176746d26
za47d393189ec31d7f46ec8e6f6940a8baae9ae8feb6958d2976d2aefbf1c4557ee871d5473eb24
zf17ade11a366c2d4a11f0a6d9ff6ec6f371ab93f1f3481c7b213e0a1f7f6520c0c1d827d0f4821
zce05dbbd8475d622220033c73d7857d9d1cda46912e7da157795008c5512dd21cdc05a4192aad4
z3a3c0cb37736451eb7fe55ec93cdd258d582de49237b59c1151c905cfa8ab5ae9d514b7288adf8
z4baf297270a6a7b35cb426a9b77513de8010d48da5993ca819c215c68775323cac80c9e007f11b
z45ef042da5d5545f12d6e4fc94a02f29dd02156f85da3ad3fe20341b12c280449236c3feff47cf
z155989e652547497e32cc8f598f3e7987c846026b2ce44f815ca3a68c5a45bf3508956769cea89
z7261d1df8feb1b64671f1d240e57220ea07f955085c988aeba670deaeacbdbb47040e01e26bd3d
zaeeec9de94d402027674496e01ff7369a6e9574669689aabe2459aed8821ac41835a2df90db11b
zae9b705b4f250e9a027433c594fda3bd81067e6ca19918363e23b07827cfd6ef43cb1331336d99
zfe48b03d760f5298a53fc649f11ee94f1c19f7c008199e25680ba1cedc1c77034d33bdfabb1a46
z2c38f12a9cabb0843d3e40e6ab8647528f62558400083ece11ed49645df56db1e0db183b2f0e97
zae398debc899cb66a0dab4d972bc65ae840b834f078aa31329898a96a7b1d83f3e7b862e1127bf
z6d679db7023d50df994e526ca5f68ffc8f5105a2168ee387d6529c5be5e8dcc7049d1e55d00a45
z061d04596ebbd27cba498acd0903872a87befcc92323ff038415da6b07c120a937084507f10aae
z402e739ed1e4b8fdc25ce6b8bfc318e0d1fb3bc0a75ff4efc35a2afc042507edaec64c2c0d40b6
za4cd84b7f6a02b924ee6ba284ec08a2b09f7c6d7007e43fdac53460b3bd9d376d23b49a84eb658
zae3aa254cf7293b25b82b51e2d68abf5cd2299b0a0ec0ead741d8494d56c62446c8e3445f4e578
z0f0e056db7d75e086986b1ef9dbdccf78c706afbc18f1f57c49d8de44b47cc11633e01e8898cf0
z2f9e5c50c9247b797049d5aad9173569f87a9c4fe37cd5afe385a9bf7bff7aae590c62252bab87
zc77bff28519c24dac3ffa95aba55578f92a6e99ff47b83326cb6e8a53fbcca9be2e7d981ffd1f0
z8eb85d678e30bc1621fc4b4fdfdaa9db998388a28e660762cbf7036ac0ca164630a6f76281e8ab
zaac689629b88d4c512afdd5ce4d5e4a18624d9ad00e05cc1ecf90518a3c859d9a30fdc3e1b60b1
zbcf4778fee43310029c55ca4914990386c635987eb6ec662d323055329910e267bbd3ef19f0076
z3326b94b1a922313bcf5c95adb6ae4f4e831dbeb9dafe8e338c91e640f4f05c04abe9b5d1b8063
z32d9aaa92ee63355a818c6ff9d25027c7d4ae6c39a06a9d89161af16419ff965e139bd33b47cea
z0afa50ecc13aee6ae8bd93f488c4f9a11358ace5659681bff67198e8f2a7db1c3115d199927126
zb1c56c4f776dae15834b3f09b17cae7898c16776793b4a09c32ba45e9357d0dfbba38026d852e0
zf366ecff0ebffe416c56d7d5b0f0a40184e8f9009a439517fd64aa008612d73920f50f3c8e68a0
zc637feeb6c1d5a6fc86c818f6c0706f4bde5688eb1d9abebccfee67209803839872d19c4ed4dcc
z62e1a9bbd009c75495762b87be83cc397703ea2322a1c1241568ecf669d851a33d50f1eb4361be
z39ee5c30360a116044d44ee9a494b7ba78b99601cc8097773ebb623ed34e018fc01ac857e578a3
z26b3545894364280366d451615ca2f5262bcb54bf6a25fa00e3b00a1c2d0d7411968308a9543a3
z678d9291e62492d53cae483f5cba4838895b31d01bd6414d11579113484510d6280e78216c36cb
z84862a36629467f5bf44a0ce3ddc2b28ca0ace2fef5a9bd178d2cc1d6bb3dc7f3791e7f9ec38b9
z659a3fa5c661ff4b916af11ce15f136856cae30f92a3a8ed8ad5a73b08d0950f5bfebd3d8a87a1
z526cd21e260b1e19e2422022cf3af88456b24a84eb92e9116dd5013620e158ab470e04e9aedf6a
z3fab2f1fc0ba0a3518b8a5710f9fca77f709c32c95884d9dcda0315cb4cbaf4c942f64f3df259f
zb17a01e9184f5e27e9a5255f746b31e13ca70c32b386f40e79a31277d455f8dfcf4a3e2fc9bf28
z26a82d0237dc74cc306b8c33b4b60f6688640870e27a9070475f009f687d04076bea9704dfaf30
z7f1d7447f0734599570011efc3ed739549bc8b63093605f304a6453bbce40b0ff6dbbeada7a133
z15a55d26c4b04fc5a3912d5b260adaeba58faa1f6d0781b38769474ae16036383e9483e77d2479
zb529b7a90b71220cd75507793792dfe4e395f83e528e27b5647d96204ee791a1e5ed578c8ddfe9
z79dfa1d6e38f8038f23b28b5477dbdcfd58ce98ac31fa541582a6d4a8529ba8cfe12e5792f825b
z34f3b182f670a4fc2e6e3c849f78eb97c4c5840dcd339418a31ab2979225067f08220cf11ca51b
z9b0160575d2b8d102b101cec0e767193c24706f24099b7a28f776256f84448ef2b4bf72b8b3631
zeaa87e1ad50aa21c1067191b13782ab8d1e1d7d094ed8939cd8ea9202d557c09d1bd82693ab87e
z7491aecc6b2151f5d576a0621964c490a8b31cc1293de46220f273b05da5ef3fba785c1063accd
z69997139fa99d6d66475cb97531aac27b6a8aa2d013f8bd8cd7485ce625bc0ae1bac5b6e7875b1
z4ab9fe16dab19ff7b4cf023fd2f00a9051e98ba0f8632b6767f538933661ad4beb02bb9f86fa0c
z8c532fb473c09bd3db7a68f7a44b7f98c878320e19142ea8c986f3c62a8107da752ab7a4529e60
zdcd226f4701a313862487cbf0e89cd89355804b82b9483ed8d316ca59681a11d82f46efbb1dcaa
z093f30061efba2ba3eef57aace74f932a2d43a053e2c6d70284d33f0ec2ca4046c1ff1820cc1ff
z1ca74b313287408356fd5bef6c61ed6db9f9b01569f13698bc526d4c1ffd23694fb16c1d9ff213
z54f54ea727fa40b3478d9421e5cf22dc8fde0363034efc28cd2b9d3bb502670b62f77ce56b0d9f
z2a6a7fc2da93e1a23cbd3686ec2a478893d88294173fae7beb4db49995c28559d9c99c0f3da634
z33a5f806bdb5a599a41fa58601229e4d54b58661a1fa8a105f57a1c98ee811772d10f1a9f58791
z4c1e84779c20ccff6a575e28d5f6d0ca61d57fc87f00b3f5332a5cae7601e4272b8f7aea32b0c3
ze73093105e91837c00ec62dc403017fb5e27ae5e12af29de1ce820367c558a33aef6d17726bbd4
z6077bb852e4294742dc5973080585fab95bcd270f2eb7889f21ec4a83eeb1638e005ee254e9fbc
z6fff689200260525fb63b117817a4f10e9385be9bf13a2d1042e8d443afa7da378397ce06ae4f3
z93b980dd74bf0e44cf27480d21dcb4d0caaaad7390df850725957de3adf6d236bdc094e308279f
z0b6fb33cac70be709fa01abd844573d2f9f91b7e209293c8a87adec0436df5c676709fd1bccc2b
z4fd30b5b586adb358598e3efa9ef842047b2e4f8d7da7aa1a370d0e4bc4f7abfbd59a947eea117
zf783a002d6db099f02d1d4348ecaaf6f86e26601a09b6d4ba1120663ac41c72f4e436b59023cda
z164bfa9d703dfe7c71a474d3d025242f2d9c26f0eae3da9fb88c96969a09db13a82a5d87247e44
z78836bf7ad3937d11865f977bfe8d15470d9dbaf4aaa7e9984a990c9fe1336a887521cd721ea76
z10da52a00fd69528202cf81379d4ba2f7f52cf5a9e9b1fdf1c801862d96d445aa9941761a3e9f2
z443ef17e8cf73c56ce74a8f4a3b230048cccfcf7b9eb30e655bdf1512995d177c8c427c8dc3042
zdbcba6e60a8c53a95b5b19c4099be471bd43afa8ad108794b3165f456584bdc053f32ba8a26fbf
z64259db7a8c893ab1c0d213f6451a9d701f9d02a7c01fcb33a0d3404924aac8d461696fe07ee91
z82108189a9a175900aa11c2949be55b3fff88b31e873b45817f44eb154e37fbeaf8266585713bf
z64939cacbbdfa6352486b1b758b562d884c7f91154157ba130497c3d2ade0771307307191edfc4
zc04e2cda7716525517070f0b84aea34c47b4665108395a79a2e5adeee4543ab9c92fd654eb53aa
zcc173cd6744db1f3ed1c95c7af17cbb2f3a52a387e8d7e54ff6c92df2a8513294be5361a615efa
z018d119c7b20b2e564745abb7a7bd5f05b7ec5fe9cb2e90a1775ee74b8d94975f09a42f1b54ed7
zebcd00da05b16612f2b6bd93baf39573ff03b9589754fa9a1a912b0f5166de5c901f06927931c7
z4256a02bf342a2656b28e5d5c5c9a60caed1f3f73b7db289a612cb28398d1583060f0e0d4c38ad
z7a7d466857fb015af3f0a831125a9796ff47723d963e27c0395fc4f4fec414a4a51909dc7e93ae
ze4d2b04ccc05721d4307437357deb81f201da80211156157f4b5364ac8a7a8cf113562dfd0e290
z420912aaa684ce3b63aee333bd346a79a685cd1d0059d2dd36bbc003c818efab00e5e9c8475a24
z6a1d7e0b2494515087c65194de370c75184378f6d61ba8e2d3f4070410f2df724ae4826b434d39
z2ed556b2e5dbfc8d58ea3f33fa1a26080e6aab4dd8608bab6d983e5f8d8a7407cba1b477b552e9
z63a962e7c5614015631020cc89deecfbbc6d7cc4d34bf7a16803e8d85373bedeb84da3e158bb6e
zbe11f5d8425ab906d76fa783d45d821f3a571680438d22de2bc22dfe5ada737ab35300f4dced69
zb0c3f9cd880c1698e90b1858fa2c1ff29badbf920bbad5d2ec8002e76ff095a2c3a7bbe7de9da5
z6bac3211994c894cab81028290a1e48129fb767d7a4d73ba312ff46fd4bedc0770e2f89c5d5695
z57459d5e480642f2e1c32afd1f56cd936144807c884a0dacec7ffe30c6591fa81d05af59bc03f2
z57c3f56ab1ec002bd33add9f99a5719330e3145aa53a832b86247fbd554139c9f5b1f324725d97
za09ecdfce7a0fdaa682a2f34f40c6bd256b2ba3f4f39927ff25d647be3d7e41873415c34d9d787
z177092ade6c96fa14d4616f0e22a6a5a9e0c5c9019172d1341c4ab3cb11e117c9460efaae5f7e4
z156cfd437f6901e7a93d8e34c0b4f4031e5af8a8de468f8bb0764ad11bff14df91c080f52b5941
za1e6a73b3f20623b92501ef39f23deec98332017a5f5940e9fe14f98ba423c444014cc19524a95
z5e4c1ba423c657c4c01b44b3790734cdda44b96fdbc3414e6feefe741fd68ad21d7f107889ccd3
z2d621f50df01009f0f81af3888edadcc57c5c157ae7c25fe14fff06ff2678369b5a40ecba29af2
z101302399fe6491cb76a2a46f3ba442b8c0e7760e43ea155f26c9c965612c9e9e3d8cd00dfcde1
z40de0b57a7320bb302c490c8c69bb782d57437842ea09e2f42e06aca0b729567df2150d755e717
zb9c7d9bdc8300b5729c9dc8e9c648f7302d2f33649617839883cdd91797a3526e883692329841d
zcc97510d978ac8324218de5fe88235573086cb257febbe02f4dba3eaf48578f05143973a36a454
z20d140453347987fa720eb72add40fd5e2d40cb0070e4f290f0ccf0f6c6224279184e2fbde782c
z6192eb0423c3de94ac78d9a3cab7c3a6fbb66833447a22282f8667bfad3379b1ded4f9eaf8e88d
z1909a2f675a4b9d7c64f87334b036cc66400e8e6846215c90210cb5a75ea7bb9b7918276f3d92b
z4c765e294d2f7cf81d11812b4e442f54b504a27aa912694a4e6d379782c001f5bf355c37b410cf
ze7bbb0a9656676ed364c713aa35a0e6de5cfc7e08a8053149de2c381261b3d535f28bbcbf9d80e
zc5bf38ca476cc2ee056a06ef51e4c0302a4daf6255d4da1ee5a54747a74444311af212d4f9f60d
z7d689c48e4c6a1d80c1d1996a398a3b37844c9570ce38ad8354c0c42bae7d5ddc06df105a7ee1a
z41c09ee2cb07635acb7091f23e2dea5ef3c3929e3a94f710c56d543fbd64d1eca88e5be81458ee
z2ff58c40549bc7561c890c829d641b9f3a9303ff5d6734ed28204ed6635467c5b17325d20a12bc
zc10ebab5f84aebb34e741ba22e9ccd7aaed2a37111bb93779e530d52d3346fe5c1ad09586c97cd
zaac35a1279a06624d64544c87b1410783a34b8a449a0aebe0e652f661bb8b32160bee75436f661
z8859f84c218f2d5576fbb33ba4b0f1071dc1a3d7d46f2c4cba2d2e2380befa539c645c7c984eab
z6388f1523227f320460ca6b870d3ca26ccae500c46de9cd4744868598a09e5f382b3ab0111ca1c
z5a01e5b19b8a4b4118fc3cb0de94af1225649292feca38e9441289dc739e12c6b22111ab76a931
zea63e5d5900a27e7ea7aa0cf78bffa14dd0ee76a796878ebe5119fd71a6f94bcb8e32a4763ebe7
z63d8fad5b2e86de1d9ce11d4cf20d303bf4739dbf1000774675d1ec2fc17aadba282f59834f13d
zd3d4832b67a63c1ab70f74a6a7e203af2285b6142de5bcb5b36ee2d1c4344a3d0fe5eae5bf7c91
z3ede9bad1fcc94815c34373b40f3b2f12651355b800edaf3d7c5bb8cd9a81c01ffc0926639f0ad
z3674593d781944659d6ac67d35ac8dff4bf57a45184837c2975d1ec9896411bf1d533eb30ac1d2
ze82fc2349b469fbc181379eb87bf54ab159b084d22037c7cc4d68198379f7d629107d1927d5ab6
z258ae1e393e5d60e6d6d592855b89aed00539d6b7ee3870bb3ebb8e8cb4ceb9a6eef71f7fbe462
zddcf256e0eee6a235511255c320d0ee231779468612b362c468fcf3a6b6476bcec2a699668cd50
z5f508e244b82e8edb14d2dad2e0e679d59f19c899198d6993a0da254e9b3267e0363445eab130f
zb05265693b68a52a0a88ad4513cd20e9fbf774c36e8bb25231a6713e7a3af0027203f58341f3d0
zf561251a5269c7624be97e80cf0ae9843ec68b97d595241d882e89c349cc30a1228343cc11c659
z52612938a6f630867004d3b3d020f02ad34768311d47f160c664c3617a58b855de75ed01597a45
z3da89a49d6e5dfc240e81947878f5fbbcafa98c187a8ddede6a4e64394b043795e364e7e89f23a
zf38564b47d1ace27200380ff995a6a1d1c32104cc419b966c63a068eb142e4b61917726ec3009d
zeb79d204b7f615d0545ca150d09524d58796377eeea5bb5a06808103366e1fd3ac584e14c39c05
zccf679b1b8b445d2ee7f3c2f11acf941b3599d7ae9c806f287c6c4aace462f9cc5f3ecdff97e98
zea7a103ac7286e004e2f5efb4c1677227520f2b0ba9ac826f61ace30199d3114a816256943f562
z96decf8694c727d99a36c32926551f481425a946546e8381b4174b8e01b64af8e1fb118c0ef8e2
zec9890f829ddab8d253dce05a60f3a49511ed24251e5186fd1d466b2dc104fcd8b68a47725fd14
z91a8ee00dbda70aa1ac56d26d4b06d771e73dc17bccf267c657ab39b3d5ea1f420a53a202a8892
z065f35226e7e8dca1956c2eec656ed474cef8429ca8dbe343aa401e266386d447ba94257e6336f
za001871653d4f3c4005360c6431321c47553d9ba369f8d7d5246ef524b4c609df76898d6d0cbc7
zcda9977c79601e822b64ff8b860e4620c0278712a117afad4130b9122962303e24bb00f34b3623
zed6a26ce864006f8f9caef378cdc57e56a68aacfaff6018a06b595fed6ece157d877b828089183
ze1a809126fbd5715e12422db301363b03810d223e79b1b1e1a36197c4276a3a67d829c60490303
z368d31c72d8dbe0af5341c0eed954362e8cad0fcc619078bb6600444a18c7cad0f41c348e75a61
z0b63663137fb43c286aa729a2cf082af7afc23f366a32a8211f654506d3894c49564275ac770dd
z01519bc138317b79c2cc5ce5ecde8a1e0427ed3daf645984ddc323ffef52b77108cb2ad080741a
z2e4d7cfccad2e2031e89a93958827e97d019544a5da30546d3584f770083058efe36beb5d27731
z65107da7d069b369526960ca868b895729726e30fc402d995d34136d4431e0be5af0d7004a0229
zd0b46e7cca0fd4a3c5710a9488ca8db3c4ef21858ceb08cc3a4e03eba550635c04c37883b2d0d9
z1103b7aae04155f8bcf88109aba18a0c15a47dc9d21a517ea794701cdc46e2a6e0a308ba1215ca
z83b48053a9c993e8241d5b357b7a03568a30721af42d6a2467d6f80d9804870768b138518a3c4c
za912a27882ac24ff68212651ff64393eb969bc61f2faa294c072a9505552128eed2bc1f19f6104
z11fb2432d951bb6ef9b337783b63e76c142e2ff5789a83665e8cba0ff64c96e4f82849dc61dd95
z875f0f1e752428710e3e4511558381d84a05c3db6c91a06b5cea39abe643c7befb550a0e5bf039
z8ac7aeb651c66b8efe03e3f6d4cebc8eb8bdfe66f8dd39100d3410fb37a67aa9b40b0e94fe285a
zaf2aaf34975e256fa8b6f3ccad209f06a7c9871cdd0066478c542c26f6880a2b681d1d81218db3
z3b31ae374bdf40ebc0d99ea523268cb36590ba24f3d4381af920f89678bdb4227182e2e8c5b224
zcd79b6ddf90cbc719655877d466ace87713cef382a73261e6d7ff04531b04432e67e9ba549c490
z975a24efec417fd6acc1360d8243488a41a97e6bab39b7542d89c60000bc53c8dd38e76cd2387d
z2bfa4e73bde5744feb848de01810142e06aa3853a4c2b214afa51afc119fba2f909420142643b4
zb44d8bd239e8ebcfd5c29cbb85182e1f96a459f6a42c381c10f78aa6ec5837eed0130eec9a710c
zc57dd99878992d890577ab77a0dd98cd4960e129d50cf66347210e24a0ca2ad7f63db114cf76f9
zd279a99f03b4d21adba2dc62414ad62f0c5c7bcfc6a125327be610bdad6687e6fdb96e700b6fe7
z7c0cbe87c12629738e553aba8e12afba64eb7c4e3e49a20c293307301a55c6c27b506a6ef2687b
z768b4f70d06f1b890be379d054e2283c2dd9352f70d72da36bd9d7f79e5430082da9171f48703e
z254a918317d2ca45963debae808cd90b8560b7d8d5cfe911c794b17c2063d84cc5b11bd41c174b
zb8f79608277762d8b7eb3b668a5d31e17ac523718edac354881e8e7e7b353e9c12a60d379814ba
zcd80c1e246fc5a2b0ed5e2a5aa228e1565c75f3b343941c3a8552de739baab037168fa3633f726
z4148dc79005f13bc08db80d2cda58d17bfd1a43a0f8542cffcc58314f5e1c90c3c68151abb7320
zc7c7be833dd16fe038afc54e4267f581c5906bb755062339a33c5343b5ab095a5bb71cc73866a4
z0de142cf930f2665997e72e70caa4bd987fcf6c552302a3703ab1da2fbcfc0f5db374dfa05a55f
zc5c8efdc4a91588b8f8edd11d2dafcdb43485b5d8cd352e1a6ae60682b1a4cb8bed95bd537555c
z17379eb600706c24e13e8d98458dc7a5e583bc850197c4207b96a6ec0073fd4a5276085c626243
z7bf4d0bb20cfab517b5e454a6ef314bd0565b0b09ba553c06f71a4652ca5b0dbdc2503bf7193d6
z07401bb4cd9b0584f2d76d7c0ebda2b289540d25bae335e9326c0a89529fc8791ae2ca9048e312
z0ecd146bdc21f01198f24fe0faacfb790c3158fc063e1da9ef399f2176428b31f3bad55e32bd68
z014bb20c1f37be9aa2f75a5f167aff193a894af591e1d26961d6ca7143dace1bbc7940682fac63
z4d1718090dca7b3cb8a8e32f34fe436e10f8e19e02a40e46a4c91b0eba73c719a9bc8fdeec4e6f
zfba6490268aa91d12cf3c122e1979f0b13f2d707ad6cd4a478b9a2a1687c1c0aa8c3c9b7091d46
zfe48680e8b776707ef0dab1b46ab878b81494ba91f81064b9f93883cb3340e6d5a6b8b03711fd6
zcdb2dff1235e3ca9fcc99dbba051e39e9d5c5166dc164fc86ce74d7a8fe27bb18fc4914dce27b3
zf9ce4f056924a766144e675df59e0b2a52f1745bf6f43ef806410f785269dc582c58d9848470a0
z1ae832ec0a08108fd71509e861afd2fb2f615edcd138ef5e94302a4b9ac04afc45e409b1725390
z4b8ae7b371b45aadb09f6e7e204ff61010abb53c9de3226c475b567cec07211c279b7997695f97
z2518eb21243a5b1bd26b4cb4d3c0e6ec69f50e8a4e6ebb3eecc94ebd31516f5ecc517152319ddb
zf224c1bed1f78ed22bdd89af8de23c7d4a2fe4f6e8680eebacdb3b96370b4b8de84716e8c74825
z9e15937958e295d81b05483f52b44a84047388ad2829be32f1c501abe72549b428824ed5f1e0e3
zef8dc316e527a889ee3c68c56c35df3fdc477be6fd423f8fcb212f6f7f91a592b7895c2919a9e9
z4703793ca026fdec631c0c7af5bb69f53509a7dee438e9b8d17eb944de1aa9ce18f8c8a01c3b5c
zd6fcb6b5b092ab7234f6515c4dbf2b4359d1c0d735c8036b515766a9d7750e4389225c95d0cc98
z63047a1e9eaf26b96cef0db36d9fc161003c14f9658e08340f1ec4f515f6fa1e5f021e3781bbbb
z52c649ecfe2292287cf28043e592fc111c2e860a7b10578180a177276bb71f462176f369551377
z57fddd84f4368e0695c232e7a6d1fcd808643314323d05012cbd6e934eba16e3ebdf92432e721b
zc66117175048d846b0be5d8ce15267d172e51d6b6d27eb5ba38c5ace0c527ad70510dcf929896e
zaeedde6d91a70669a8b3de8007b7ed7a20d32c820a47116b44decbc4f64c63c511d412a81acbe5
zeb65ad18c804f12d65ffd3d7bb04e2c91a83bc851ee8d93da998eee81a96d7a19f239babbcb388
za27bc3a5f1e763e23ac61b606a4c9eb0f010eac8e418565c2878fcfa1638ee13b14e8c0da76d9f
z752b4fd310f00ccd02362889ede2c10e7c3a9a059a596513f6e9b79de16787239f2b9f4d150083
zd3576ba6a696370af0b871e530c597ec09e10a7377feeb78b6536bc89301018bef4b56bb19207c
zf095fdbbbd11aec1fe3a4f09b5b2f8a0cdb2fc2f61b64aefcf0ca23596d8dcc2a50998c25b2cf9
z49b1b0c9d3dc5fd1d0e71fcee3a730567dcd71529ed92b0c75d9bf3bc9561c2ef1f74553a99f8c
z95b306d8d9c82f17801a7638f800c8047cf9350689e1a2ecbd517bae178339eefc5499beb30089
ze132b1dde3cedc2f5955902abb3ee4789979a531a54b72967d6160adc76d9105878be49fc810dd
z32c55a9b8a57f07610376b1045c3cd508a8b0f21eb5b452051102f7069c61d8b1f0eede7f2045b
z461289f901964017401d2ba3920c7e531c768aa1f5de422a125852ca85002a995a021c8d06d0a1
z25f0492ba65b4739a40a93dcc770f9e533587ff8fc5e8600833709a6afcd232788a1306640437e
zd9063087346e722c7249f02837ed3e249583a42694c51442a04a0fae89af96c0faeeea012d3321
z73bd5852ca73248863df83fa97066f1f01a35dda80a124c261d42e1937577229ff7aaac198a5b3
z957d0bfaba6ecf22d4f7fb86cbd10817245d829d75e79f0f96f610a1cb5fbee3b25677c546bc91
z0c6d45e6f41571987e82cb79b645d4d18cdf7618d4890cbf50ef70c894fba0d76d8648e66398d3
z0812558a0f9bd3967bdfee2096c62f3ec9b653aeaa6c4ec4fc787e0d07589008f0be2487b38314
zc33c6c3f64bb47773616657ebb9f2fea1e5487673d10ff990707d1e14e7db36076e84a33c0d3f8
z9b07a3d8344d852a57920377fb7e62e8d9645268755097e38a15cc24f2d3bb84b535ccbc065aa4
z63d6d0c1fc8c3ec7e4b8c2758cb32b7862ac9dd342e1560ca2a9e0094cc18b98db779b4acf2d4a
zeffd49ebc04d15b950592abb178e46a18a2710389d0ccd2375ee6591f074de57f641fe6610b948
zeed3c4d2ba7cbc8698d7919d45bdc9de62987cc35307505df6e54ca4e73349db924c556e0b07e6
ze126d7be3dc6180f179a83c3ac8e2fdbde102cd25955c70e51347c2125ab736a7f78c9e9b8fc5a
z1786b876fadd5464586b4d2a021ac9570296c5573a8f5adaa2b573c9c0250706b8d761aef7ffce
z9425caced5e1f800b8bd344964a4475e7733b899eaf63fa72f7166d81ce42e3338e6230a891b5e
z44bbb8e10de895128168a82861425f63f02c59ad3938f06ae4acb5f010381e5ea1f63f5b1e0c19
z4b8e344e86d489436301eb6151f8c9e60a866b58ebe980942ef24570f5b4699f69fd0c77a15ad1
zb5ad72eb789769ebbca8b406541e82625a1701a740f73a7054e62fd7af0ab8cc1b9aee91179f3b
zf40616a4ecf61ca0ccca768330b48f2e7ca28de88b216c31d2c3dfaee3482a39d4731987c3992b
z55c7d36b8e45dc124c0f5e40cf3a51067434a7abb3fe2f8d1668432dd25c49177f8590c821c910
z730720d8c9273702844a5ffd22b02d93d02b41ad9b8f3901aa0461ec79fd5908444dedfc6c437b
z8749188783db02c9c5a7ffd7dbdcf81c2ffa7ba3dcefd8cbfcebe3ab1c8f959d10e52cffe7df66
za22a5c77bc1372beeb560d4dc8b4109c5167b9f5bb251672d9d54562780146f921486fd4095516
z3017a7c8e1922156ccd1a0abfeedab3e05d3aa43ef00713eda7690600289aafe6eb54546d4135a
z6b61cf2459e340153e46cb2f2813628e27d5274044988b9982ae19fdef6b6bc9637e0102468a83
zd07b54dc7e1a9e23276d23af45cbb8ebd28996a413ff1f8122bcc8a3ec868cfc4eeb940b15f065
z00caee24c7a45cfe6f71ed634a3a81453f3094c84fde5291b0c4a0f4777587e0c0354839da0efc
z0cdb7e642e407458a6e20569dcaea28c39666c80fe8043882365594716e87f62f5da8fd2b02e8e
za8bce2986afa9c6554b2bf669efdb29c2e7915c9a23221efa8a89903fae011092d0e727d9ce529
z5e12f2d64481d664f5752d801ffa345866c27f73f47337c7933211c8ba27084dac58fad92b2bf2
z801eaa4e43e2f8d2033150eaa3217d87f12f65cba51a4d5fc8979a550001d9f00dac0d565e03e5
z622a45106f51c23e06753a08fee4626c40abd4481b6b4022ea1e05012f9d020f2ea30dbc04ec57
z44ec430a4f5eb65af2b9a4026c14499a76818a6b5d14d57e4782eb8806d05e3995b47ef4b3a573
zd27adf8f354e1430f88c3f9249d1c52819623bcada59b352e44d8e18dd443378fc2e057d03543b
z467e4e1da38ffd4503a9256e093b1443b662978af61dff4f46d4823d1c3e115abb20afc88415c9
z2c85898f220ea5fa6e203f1f494dbff78686c2a948508b117e84fbac3f35704a6cf6122e366795
z93ef2820cb60bfa417be5ef840f8ba005a239f6d0fe117b7c564f5cf56f4216e7cb86aee07e649
z4cf0f6694c25e054a4ecfd61e6917a09dce2f04c88208d2bc6b7ce2a8ce4425a97cebaf1e35aa4
z24c75e36a79355ff4629ee08c1a0e5782c6e8b8e047e48bd2eb67e6bbd3008c9932e87d2decf48
zce59baa377ffb96c944099568cd32bd2e98911488f7298c277d06d3857d8b0adf815ae232b811d
zfc6ba76b369b0b684696bd855e2f1bbb3ea25c3546c4ac2852e1ff9903a8694a7f2fd3f20021ae
z927bd035040efb3956bfd47cfe4882ededf29294be32c479f691cb4b8ff12c65f7297cef50f666
z00418568ab5e4126393d6c287bc771d49aaee6a77ec8baef351f02aa1759a457f08d00cd54010f
zb9e8e3f2400f466167c2ceec558a1c49184a5892d3d79a9254e50bf0770fa9cf38baf9a29bca50
z27497318c796f097cfb2fb00ef4aa8480aa1358c92b18b033c7868c14b25147c63b0cc1dc7dd51
z728d589840d66644967b31b7b01d67e80eca1711b478012629d6dbef202eb718774c10a77b8b95
z2be56ad9640a0d4f8e2d8c10f2ff748d7b596db4d54b0bf70fe3c7dfa70d71847b8f58992395a4
z7d7c07478ada5d006f32b935d7e9e552a8f334ba33ce6f46c2867deccb732a8dc4909ebd0751c0
zb2d11163c90d03c2b034c4a753a9b027dcef1df986f040ade8dde6c0d65a50f613a8212c74b9a7
zbbc5692dba7daf186c11354f22d4586bcda2070930c0ae8c5f843d35ae35e36fdecd465a228a21
z71a8692256ca8d100701d157b46008c809548a716b5e232d083b9602973ee6c006975391a703da
zd385ec1103acad38edb383b38d3f925474ac46e8c12223a4083ba41ac1f7e09c8645205a9b0463
z099750841275f7cfe012d20407fd42f9a0f9f7eb4ab0ad86c354306ba3d619c19df1215ebcbfb7
z033af8bd36b5c532a531e8f8b4c1122a5da349251e9914a80045a2efe6075f31bf849c3b06715c
zbf610fe709a466c2d43ca942e21ca9705954ed8fe069ec9bb4bb7cecaefd310c870c607c200b29
z80643c53ccacb4f42370e4c41855144c0bfd9a71cb309289292bd2e4e81272bf1272e1082af5c6
z01644fb5600ed50a326ef6eb675bbfbe162ab23b365669c039d18ff5a4af754c34a2fff29f3a41
zb33719391644d303dc46a2ffb008e659b7929cdc8b9d5eb910b990c73465946e131b90ae98a02f
zcca25ad7af21537626bd9e759c563f3b3e060b6f10326ecba39de352d0f348d97b5e0d81a6b6bd
zebcc04c49c5ec273fedf883c04fb7964f2ce9fc6e972af71b1bc4a3b4f68f3bd2b34f431ab45aa
z12bae59917be0bf9ee3b7a27d8acfb688470061e416641ecf0d1b1b85f551020ed5c4e1123c6b8
z873c8ee19c9c51ac6de1f4d2a493a817c97ad0ce40b4f6e5998048c45d626fdb9df42666c065ba
z050204bfd1ed439694fe05ffd52d3e1978556141a9d4a6b82f1a2964b47851c9cfe564f3aec6dc
z74a757bf26345ce67dba923e5d908da10c278febc25b5a1ba1d2846b34990f95cf01c6889b6315
z03fbc572353620b72ce6870bf9c6aec94d5232aa800e5c39ba92edd8b3de29776fc6a7355a795c
z4e5e40e67bff2caddb1c4c98ded378add01fbb76bf7bce718873941b7c1efa287f3775806caa1c
z7156823609ec97a6858bf4a9a35ae6df743c578e42fb9341febfb447663613c14f441af736aee3
z64f724d5b6a6fb8769d6aaedd9fbd104762c6572e692050f665d4ada5695a63d5cc524885acb96
z41d0a0ce15df515c1b800b6b8f2589a4724dc562b5ac7d7cf887683a6091473a06aceb3d2400e4
z0f99867e1c6a19b7bcb74233dd9fdb3f531ec6853d9b758bde741e63fac02532b1504e91ef422c
zd208c366ee5b4320980a7b3059ced9085a0cc2c49ecd7cf28130e645b0fec5383fa6ef36569748
z01458cb5bab3fa2e57c70aa9b3b391fd030d826546601d6207929afd7149929911e46ef897da31
z3599a09b1db07fd17344faa00f44a9e0d5616bba5431d8a4562fb136b53c22a77e0d71d025b417
z102cbb0b0bdd78f02d814d7e0eaf2a6517f19122b8696c66865f2bb37f8699b8a7a158b868562f
z5652a82d9a088ddb99b395f01baac57c8bbe5d7206baa43147b22758edb1d18978ab14c457f474
zc1688846bebe146d29f8a9301569e5853205693735656bf607cf02e65461cee6c8313e6578bee1
z4f0f6b1b9836c7aa14b8ea2b71a3b7589aa7b943819ac5e1e9981c472dd9bb987e865010b1fb00
z5f7f590ef1cc3245c140d5aab5a878232e4e9e7f636c5884dcecc00ae4116af6480ffddc2dbdbb
z6f8439fcd913cff73b57c2ca4f90d9df0608b57f766eb09f925d7747534e8977d703dda3902a74
z984055403f4ef67e440f28b5b6c2537a5b5eaef20dc6fcda830f2f5351fbdf720e4c60199d9de3
z85e34a28f5c8e994f61ce8d4d72f010404757f94fe5446a21897c8e5258da9b27302238b887356
z313f120095357ad33f7a06744597a88164393190a6f3b0ebdeb211641e7394634a2e8c26c5ca3d
z630ef1022177a41ef92b445f871d1b881c65b6d83404826c28b77ed174cefb49a865039046df7e
z85b16c434f7412827554be9f75551120ea312f5ce34eeda3418e464012faf4d390790c4c4dc952
ze0aafdf0a9499dcd219bea6a514c394f4944e9a6c255d2fd7db170edcad55f0b827af603365f0a
z94cd0bfefed713543a845d3ffac861b43aaab2f75f5ce5f89af83a13745942c0af803aad67d28e
z74b8ab665ad5c34b4333c562e71f27aca4387e3f12980dfb6472d38587bd1e3e820daf2774af25
zc414eec1d74eb5e39c4fe17aa6c047fee435590c6ba8c2fa41cb1f4afc6ae2c2f68236400f9c5c
z5c93cc80836a07943a5393c6921e08e30b2e1d71a3df19d75dbc26f6b093f24eb54ca35c2d88ef
z32f073cc1a83474db73379bf78ae2423ae87b028a2e03238389b75ffa5b92640146fe5104aed6e
zd5317dd9f3d5c0f13d016401b1d29ac07046dbd5d62033ca8c2fb071747f9440ba008e96a81513
zec2cbad86c767da34be9d4c071bb487cc820d387c3556b9f29bc5950d4a7d851131e8dcbfe8a06
z816581c08cfe10fc6b3ba29ca9dfa1baaaf53a52e70c82b4bd1230011e521f3d9531a8829ae21c
z468e8699bfbfaa7b53b76dbacb63285b5aae0a772b0200c1ff2590d83d6d1ac9c183890fd129a1
z36d2666f45598ddd737197b768712455ef338e93d10b0e36741989081e24693de46c1f649dd3e7
z69d225516486f5673d124186a011cde0ac968a73892d8be7d7fe3ebb2040b7853bacdc7b95e162
zaca4044df5088724628f9ae1651f2db43260aed3d441a0383f5ed5abd3b16ffc159eec233f9be8
z958a6921ffa1d8f61a647a008044d2ebf8a4c2ffeeaa0040e165941cc4e2fd2c3c75ce5a959fc6
z2e64ebf546395ffdf0cd7ffcb80aa1b643d97efd540e67fb49b3e5136297734a1515888a4d4f4b
z5213190e822ebbcf9f246ba376aaf16bf75c7995a4b8e5bcc6b39c5a8e559363ca04ab21abdc3d
z636b0b913ed02dd22fe8462d7a2f32a123013239c7bc8013435b8004a5c40a2b5fe3aac5352b16
z59ed1e496e399025fa548c4e29bcfc299c2ff3fc126796db8398ae1768312359c53b9ce454ab76
z81d8754bfeace6d4bc2b4d3fc8bbfda9c60d1b458afadbe71452fd14e34ca6b48fe590198b6b78
z2595f8602ea7780ecc9abea149c995aae2db37eafb7e89010cae6b8bc4ae2250343d20da0899a4
z5fdb1740803d5832b1eeddbccc6955d695b8fbd72061a2c65f6e51e8886da724afcb09fe5d9125
ze1e9ac47be9a7c1acfb4fb16c111c08064c880a72449ece16bc953430606889e28c4335640576d
zf3cf5f7b618109a21c1f22818f1d3fcceaaf3b1b8a76152cb4fc971eef3885396c6b8190a79c28
z2b0c61f5925e8a67a446ae9f95d192793f3ac2e72700275b32969a19b49a0ff6a8d3a13190dd1f
z4ed8b0b58309ee06e0f88aa9a5ca0697d4537713eca3e68436e3c195e7048746bb1aa0bb92f21d
z3a8f9d047dbc23360f48107c409a8d2b22109908e8a9846ff1391185347225556580983cdb7b27
zcc09c3455f500f5d518dd0946cc7fc9c8ce1e1f3d9811c344deaf49a6819d07ab5942301763639
z32b228a072365a152e3a7510f02b2d58e664d9412531c303bf0d9da5c490779fa19e1ab7b74568
zc8a31d5078d36ecdb0d504c54100726a81e9c0965b48e685ae463e2f74402950c888e647b844b6
zf164242c3bfff50b05e97d0125bb14f2076cb3746c58f9c5f2bcecc6e93fa8bdca2b222e9a0dfa
zca821ad7b11e797b6e51e1c8a4df803521f85c6ad01f81a1c5601fe53e14d07c2121d4e267577e
z0a812dc5de19b9d893c7ea148c37f4311b96038bd7ae5624a8797076b211fc23a95788d91278a5
z97a49c6e54c64a6c4c6b457207e222e0f199eedf85257e9cb4ca75266ef3b3aaae8fef26de621b
z2c1a4f06c2fe329502d3e096fc0e02495714457f2d6542c26b81cdf96474b9b743f458669e564a
za47a17b7cdcf5b2b04955e4a8df4b5c95457c93ec8ecc09e9aed355dda73e5e55bd88bb63e2eee
z64ef468c6d8be1c2c7ce95624a917a08d97b2f38607549980c7f3180f38cf27a4c134e7fe08a02
zcbe89dcfda96636dcee1b25f4a990fb510e4ca0e7817aadb1c022969270c4ff3c15aa72c77551f
z72163639fd196e9b5f6414060e49dc87def826b666fcd25c506ab9a1afb03de410e1c8258dd3c3
ze80c50c6e5f9a0ebc4ad973b82fbefedb88a033281ccd637916e83f3392ef4f800753aaa11a2f4
z8de5d828f09b2ceefcf16f91aa1054c16b38e67f993ada4568520be6968e3c8e4c8f0e21ce7fc3
z53e0e8066d7bb92a43553716bb61f1d93780ffac5d1a442444955d7606bfac5ec7b465382ca6ec
zfd26781da0818332143eac2184e93562a843baba22a7e052c8bb9bb7762ba4af7d7f8fafaf2a10
z95b2369ffa033843fbfef9194db8336e6382c287311a4e851c96b960d39dac4652d0bdb661af99
zdf79852d54a933845bcac62a9e6a7a4e4d2e983d289cda54f74fb72a991607c73d140876b18587
z431b524cabb200d3da70c07c74ee06a6d0a524bd5e722f897ee486de2809cb27478bedafe910a0
z9e3d77e295b1583cd3d3d79f887d3f4c00c2146ddf71bc952cf48fc11a2e1889b42e212723c569
z7b818cf7fc4550b4c9c618bc5974387296570087d643d0499093ba8b03933b78520ce1d1e23176
z39862f2c5352e7f30a9a61e8252de4e6bbb9dfb36e3d831cb355c5282e28460916a5e341c6b2fe
z1b766c6a49514776f2d8ddd93a8d3ad4e86d2f16535d4a1b2a84ada285e4b4e8d0e870e754e3eb
z20ba64af36be6449b80a0c7e6ead1f876398b359da850ca6a309992260912fb24bbaa694195e96
z1b8e01a5386d277c390d7ab402d36fb13b2588fe4819614c6863fa13b885b8522b2cae2c248c36
z5f55bcc010a188dbdcfda93e410a142442c4bd1cd057935d29efd3c22e74fb85ce1d02b2a6944c
zda21f292fbb53af3420b5f3c266b9973dba5cdf76afa65abc03927eb6bbe7cabf87b79ce3686b1
z2cc4dec5282d1f2e27447daa7387b5957322b52f06077eabbc509d47aaab3e01b02850ab44359c
z5efb34e32892648c22b51b18e08d09f46322e9214dcda9365f4c2490a759400a6d72586aaef5ad
z7ea9853d4d1787fd0f7708d5e6ec469831b68c40c98852ed5da8a7dc3c7c091b040dfae6beb1e7
zab4f9c07c592c6b5f0b690dcbf576295754b5af3e8357248c785d3c1324de899a40d256c56a073
z07d420248c64896ffb190278c57924252d7dda18377540b3742dba56aa8b467768243e1c7db3d2
z8bb4b62fe60f5974dc1076556147f1497c25d733d2400da31f0eeaf341ba48cb7b07e1e9703c60
z2ed75c7791371278fa7a085b230119055fece05cf5d6482670df6e72debe25873de8f81cf8013d
zf9b6c121aca449008f5cfcb3d334d66b300de4ed69505399bbc54e024042296c6ac724997cfaa9
zfdc5615cede98bed47540f57a8610a58b827bebba7693361639f4bd48d2474d69e2bf75bfa0905
zf1c37ce748c73a218c28a8816de8436e552b9559318ac6495c0c26a7983046a4b59873ddd091e4
zac881c0d11de140840c1a87feccebd6e2ca3a10370e737e47e269078d88232d539db2566ec82ba
zdef75b9d75550e0564b91c1fa111b0cc50e3347f5336fced0d186b2096a2fcbec1b29d69577587
z858b4fa5664f00d8f2471a8de0b3556b6c8e8ec123fee565d4b29a21c0fc27a63ea4454ff0eb4f
z4cccb2fabd1d41a6dc62fb9f1f5472d22705d93188430b31b7bd8b45a5be12bab199382feb6ea2
zd8d1769d8427e84f72e61c3685796215a2552b2576f4c3643dac531898bbe4c97441ae96ef3bd5
z344b7195ae76a48b5f5c8780ca3691b27c3e3190e88757ad9206dc5e47d7b7031cb24baba4cab4
z4f3c9f32c02f72963ef2e24722defe712893d41b3726a57994a9127f750035f0512cedacc57cf4
z69882f1bf5e15af5764b576ac10b1ff12126635e0400f6859693d17407a687312d322834aec56a
z1da709f89ddb234142fdeb0d001a81a787bb0a6b037f41e3d53862526f3b0a0e6e871fa6b04a01
zf73c7ea0962a449d4dee08d13b43c1b08bbc255ef4bc25693cb4cea2ae0ee755ffe24fb047e317
zf24f43e6d971a420b885ba27e1257482788e11e6e3c42696a5ad003729f6a55089a990a6dca352
z325073d47b51746212bc775d2b523daa5eabab6be51359046ea7eee2f6622263d0d6d278d25b1d
z0e5dc632c64856928b85339838aa636f65051ad5463cb6a8194d005f75b5696b8823048ba781e2
z03502fe119de889a9fba6b3bc620687144a6829a63e1493765e5065a10c77ed503134fee4de2b0
z19109f21a940a5472fad6267d909b9e63685624099dd81bf522f617419e1339ddf69f3873e6eac
z21db62324b13d62d741ad81742b9052945aae0fe075f14defa0b50e5dc938c62ddc69e17edc57e
z9328896a04a13cb947b6b1846356bd9ebac9405bfa3c4d7f1c94928cd428c99b7982c5ca5ffa11
z61c7e82b2ca22447a0d380e1790c790be6c9e0066a7df156162094089b8c4c5f77db5efb2eba12
z1aa670d2ff71a5b243ddbabab75c0eac2ad994f246968a2962d77b9c5def896acd2b9227f06986
zb13024f963926bf3025ff5dbe814ef63c2ea8f40e03e31d4480aa30f7c36859916b6cca01e8702
z44f259e24eee1769b4ffa1c2ed2a2d188b25f7cdc3780e3c9dd5df64b5ec6ab55fec83485cf32d
zcf77a4e063969414060877d05bf7ae3deebbafd9ee86c578dcf642dfbfc78e2d523fe1d3073def
za56089fa76e78a119956cce4ba9c16081801b008ff2a5df5b3ca01d9f42b3d5f6e626527fdc865
z809cfb014b2d6eb5a832de0637cf1421c6c632e194deecff0024b2a5aff822511de68b11ce2559
z5a9e5ff842323ef6c8924c729f9d8877c82f5f36f4a5718cf15627c44d0c0456c9e943c89853c5
z979179972c9c2ba186a43a409165ccf6a303712533dc11ca84d5e1c0bd49a87585dce50e905b94
zf14a9c005bbbbb22cfefcceaf860d98434b7cc1641fcdc4ce9e2479623e5aef404277cc2fb53e5
z1eeb9346856cc316a7332734c1dce31ef16291e22e0f6b97765cd7d60cc6dfc1bf0f3de6f1d230
z91896a4b817063847e718d12b04861b6613d6b171e03ff9e21147c49ff460ee95050076d0cedfd
zec3f1501de91847f6a8663c4dca46dd11eeea06a412d4f955b24a28f61884b873011fb068e457c
ze0547c44e1ceeed2ad5fb3c1eade5542f3e4fc6691ee7e90dbb0951e45ac55e851a5b277576217
zd858e3efb1f251ee838d574e0dc4aca5bc42710c9b34caa05c0a19fa1234a5fdb66f15dfb8558e
z6f3371edb2c2151ea244ec52fe1bc09b29b6272ee40d918be4677a0ea1c99d62a8eae201fa4a69
z42f2ef1cb23c9398c85e2af94398120172f0a69f45299406e8f41197be4df6d319ffbac0da8aec
z81eda7ba60a79d88bcec796703747609363705e14b942af1d007af826201df2bb682902afbd5ed
z68d2619bc4034dc1a3021d59b7e17332c4bdc9394e15838cfb76638ac87d8f23e9625a948b7146
z476ba621a0d83df590d0e51c6ad32231105537cd0a80f10b032151cecd889b4ce27a0b7292abb0
z199c17610b21fa3d5bb7e67086c8b4f1378e519771a0f57ae64e02e1791f67236928ce4405ac39
zf3d10c38a38704670c062eea9f1be65650093d5d918abd754876d8238e7af2d0ad0441b12c716d
zbaf16373ee994092279b8489a66f854f6a6afecf9378916dbcc0736d255d0d2b0b0c665b069815
z3f7d0e6439de99d0f465d64c33024406af73d2b2c4aca90974d7daba6b928c117a3db3f899640a
zfc48d0a6058798782f4dad1563bb3badabc3a0d701c57c2eb46f50a4637c0eba90836896902622
zc0f9403fdf8cae3fec924096e1bbad7787bed5536892e3ba0e290f0e2c0010c03b7605616a5a51
z4ad8465f777893bfcda9d13e8e3a90e2f05b1c03b57a1538281f785ff248d1ef6113f6695036b3
zd5dc3052a5eb7dbf059fbaad36444b6c6ef25cfd0f11b833bfe6e13729e9a13a9301c108358816
zcb1763e62cacb37bb6e0270f0e4c5a16a4384ad5495d3885c6aae0528ef35035b9b60f29c26848
zd6c8d6b3abd527f1603c108dafe4d874c49fad056e439b6212e55ce25bca7e9ff09feddf4ebdc8
z90ae0ebe447a83cc1349050aaa9e46061247e6d90947cd0ea0a1043423da2b7d7a5bd54f39c578
z2ea346aaeb3bdfb34971716c6c85f6b0668803e06a237aec5778f7706a98d2bd6aa6cd92f425aa
z0e99c9118726484afa5840d75d16749ef1728314a2519cdced74238ec45794694a1fa8c642312a
z5fc583d4a9d933981397db6bb1f5a0c0bcfbcd86378f80f75738c7b0ec691d6226cfd7f255ec87
za2efa2e0dc782964668a340b572f8357b658fd7920129a6684b7ef2b0a87fe34bd3cf7e563036c
z2b74efc66d3c818a899a1999b12c716755d592d0946306869ca97c4103d90ed17017b4066b52a9
z126837d9dbba25873c75d88da45e62d5a653f20699a5b03301e8a24cd471683ae948482fccc38e
z98b4dcd6d3b841dcc7fb24958e604d702e2508e60b3f6ef88b8ae548ce18b06e8cd76d121a286d
z9cc839f3918060440de67b2499817ad7ccd71757102bb1a5dafd7fc0083a6fa740b1867c02abc5
zaf7d1cb6748ad3d05839ec9cb4045ce9e1c7369c6f3c7532273ab0090737bceb0da54702f128f4
z9046bc9faee132c79e5a177ce046e2e56b464e6bf89c22dc468ef6ee7d4c28d3060767fae0f0dc
z28695101a54eebe9e1394e7e5a7065be70dfaab0e6f30fb23c48a7f8cc53ce3b9cab049fe2b53f
z930bbe32f6f10108300ef310800ee78ae5650df7b21c33ac32643f3c41e36003e3f4fba48249eb
z78bf8482002a9d110e7b54d9a80f83a6081040e946fb0cea180e4cbbe64aa65265db37e3a9b624
z6758418ea4f60b469c25201a2e1cd4e816f6f05ca783342cbb015c9c567953db1568524428dc27
zb14c81465a08ae9aef87d4b35c664c5136e62a7b90a425966db9f34c87f595f5e3793e20f62de2
zb3128e91c97154aafdb0474ab3ab548ff85906dd481aa02f0ed7b134b7639268a1d15f6252a1e8
z1556a1beab932caa8b40a9aa4b6d021b85d1e3e7f283352890198ee18c28664062fa98d3cb1d87
z844d2d7ce2e61c076e71de3fdeb544fc429035eb5f11a621fff855b17b9eb458fcf67655ddff97
z307b933bf9f7c9729247b73ae66761248a4b46aaef3e0f1622385dcde044853acf3d1c46a87bf8
zb561af07cb5e136ed22c7bc16a2f7623c4b202a66de585358d8ec4cf5edcaabf31be89534cf8d0
zb9a548fc7973858108ff45ac813ec0a9bf3e2cdb67ac87ef6eb6cbcc1bcdb8521257e7b39d94a6
za3b2737f40d143513f164566b996ba29be1cac226b5ae6575d555d7894d727d6b3f7f3a8b20be0
z51d920121692baf7f74314371cee81f1f585319982b8014a1cd5123027c8222e4e4aa292a497a7
z450d1e9296d006efea469179eaa53611b705853d96fd351616e7d84ba5402cc35e2c90f8a0f2bf
z7754c052f29f968c9bfa5e48db485f739453cc53ec7403b0ca3b96535c541b092938c2e81f731b
zb974bee90643ca1eb2d78c9954cff9452b29a67a2fefb7ed2d163f54498fd209988418fb280834
zd1a9613380eece26697e7d6df34cf7cf25c202e804f4ab823cdfcdaa44d01d7af01dde234c5d65
z981bead295e68c79b68ea9a67a24a465bb7ca0be51d578904bb387d56fcec0d5349540a8e26606
z0c0b81b374977c2ffaa01e02716975d6d145179adda32359e0389d9f3eeeee4bfd13384b5298bd
zed7a6a302a40868afd466c172b263e6a84c7b1ffd5ff341a3ec2c59c7ae3e3a71a0cf0189881fd
za854f609869e7afd31728469cad02d5f62d99529d2665f9681c3765a13a3d077ded2da07e1d082
z490d883b617b5cbd54427eb87d097f017cec45ec10f80d1a70cb82acc66ce9c317d485d71a2835
z660a6c7ce07239ddc08cddd660f5f260c4ebd90af2101c991c00830edec8c757751dd4b5d43522
zc94231e13b9ff15b7fc42e588a288be514127139a3a557b335f9a550ae6acb21ab2ef7b4e8f1b9
z919095a94e0aeb1abe7ef0374cb68a928c25bda02d54ccfb1ebccf15772d59dacdbbad53da7625
z5cc1825a3d1f5509d43d67f54c353f02f646cf8c079d572c29d79c183cd0c9eed6822deff43651
z05d55e676a3fca6de2212c52b15035793afbf9d5dfef69b6ef96ba821c97b73e7953c4698a0742
ze71d94b775168145af1a5b3a12ed6e47781a48e9686b744434733bee77a4cb2525d909a8fd9d44
za13f0e56eab412aeba8bf9fcb10811f4409a7643d50b1ef4828251644edca51b8ee06f47fa54d3
zc54487b90c6b7b2e20bbf30d23d808e2c262d9b171a49e033757afc9128dad50c3d1e853400a25
z32cf0d2d369c171d27582c5a9cb5a5c6cb2814a97f80690e5522fd693fd13ae79bd325a51d42bc
z15023d6940a545df6a779de19c4b5c97098dc33fc62df4c67a3f605576bc057061a57a31fbaa1a
z3f8bc12babfbb37126f4a6e325b4511ba784d23b3430c848d11a393227c5610b1ce146f968458a
zda56049d554887f8e51d159406b589bb8b91747b4b45e383c6bd693bfa677b1494da3f54ed2f18
za3e4ae24c0de226fb967207432a5a734cb33e5fb90408e23ea500d8a762ec929de49184deacf3c
zc32c796d848ec1135c253d7fc94e146ecc535965e5717d6267f6d4f4798ed165948737e3119ade
z4ef8b069ef315d10acd3460395d2952b8ba2d7d60697d1c6fd61078c90824c1853ac9ce73150a1
zea4ef39b21dd4225751aa82da323108e8384975199ca4c44ec0fbe2f77292dd43a65e3519d019f
z381e796f1d39798f7407203f5b88bb7b3a14ea63ac9e573ca08361777b8f4bd480940cd247cbbc
z7b2fd68c377cba73b9abd86aca685c10b6a812173fde56c84406bb06633012da272d3372a33651
z4a5d9fbdb8ca561dbcf04f93182bc3aea149cf13e80dcc36d7e03e77be54f301cb22235f3305e7
zb9f3f781f878388e609e94fd733c8d247298a17bbe677b6ca3e6f3853598a84fe698fae5037b73
z259e47a476fcc7b2af95bed71845c9df8e90791b117f125e1f49509d51e618d05a9b5585bec2a2
z87fc4212768ecf5ae8bcc6eca1ca21b4d49572f29195730ee12a0cb96592cc125784376b2aec29
zfcab3d694f261db989baeff18774794ee69ad0c376db727f5680f1c201becaa90a819efa4c72a4
zc7222e3fda44883925aaabf5f8abf4790840a1214b9613051c18fc74ea4d1ab1c671dadf031a11
z4339d210e687c321cd4a20bccf0eb399029fda2b0a91411c7a6f7d0c989ccda21a22a935a040c3
z404c1fe09306f003e5f725af68a27b41fdb50e02b9935b0f342d7bf2fd8560d1b7f557c1bd130d
za391dbb71654831e2c14d28b44168332edc99ad798e612055c1da8d6b22a5dcf790d8209b9623e
z214daca164119b7b27c57892498a2a4aefd1993b5106fd5cff244b4d29e2302163360af1bf49e7
z2da5271002183f316d15b5e121bc9a9b8943eccb8b6e208fb25e0273158e297eeb8a325d212baf
z4b42c1db7717174620bf2013957d0c20f0dfbac87dec61549a293c556c38ed0cb0ed19fc9177dc
z6b70f7fe722f2bdc9aad730cc4aec5a3ce230ae4b9efcb2b10dc7bbaa4fa6e4b23d835480a7ee3
z763449afeb8e6737fa02d27307f176b7e833501af70dd2fd7b2f3df40c8aef84dc68b24b192b6e
z0157d22824e344d0e8fe3e13665b12165aeb385aac496a2c65ac9cc97c5541a449cdfbc1f678c9
z50c3de6c8a85875e5d9362b36b454cbed831d62ab476dac913167d8f40c75b8db13d0a19559804
zee92725b6a206f5448782b3b74c61e83f6bccfca90fc32b545115e8f1e8e236396b721d44dc026
zcd2d464e868967e38b9c1d4f9b15145b97a58039663d864a9ce00033d76f8bdcfde3a9838fc8f9
z3dda2e4b0b03635dcc14cf5a9d4324e82f37dd6c3ff8df6db346de53ce81b0233cd556c907d5f6
z4b831630220030368819f3d92cf6c56d47c2c8a67811b0f7b77df61c1d267bace5f6d272458b6f
zcf4521a298bdf90eda643314b71b29f505ddb42b07c0f54c220f92c28244b29b9ec53352e50de6
z71caa09f03820fedcb8062efc7a4649e9993b4f0f4f23ae8ef5d71a85832519e7250918dfd4b8a
zad8fe85db9ade739469a97f38b15826d50781c04dd20e4f107a375a55f8ad8ca6f9c0b4a511e93
zd2243d03e7812bdbb2332d3e69743d81c47e323840f1dba7bceeac68ce31666caa70cf13edac2c
z04c372f25659d3f02427ba241792318c2751cf8dd38840688d1c2ad56ce61fea60bd4f54be4cf2
zb8074be14a90ee4137759f07bb488e2f3c18d5fea22f833a496327469fb3d03491b2d83711236c
z09c5ebb1bd63799199ecc22adcb9fc541c1274bec294e35515185f4f0ef4026fa8ee5b27f50f84
z5a8d74939cb1d6fa36b0746c42c27fa2f05556f8946c4318a068ea92a4e5f84f6e9b372247dd38
ze87ab4edf7850f795dc745b9f4de45b548216441958819f503045a90006e8ac1bafeaae9a34de6
z00ddceea62221cb77463c404443d7f81588d2b5aca29cb8b2e9ef2eafa293ec6091b7e6831fae8
z1cf2f9d2548744e1f621f758319fc396d079e20cfde071831360837ffc2122410a9421bfed15fe
zc74559fbcca1542cd7f9e0bffd6414ff6f2508cebb16964696ce4333eab9f94cb0c6143333b240
z5b6075c60f02cafc537e29db9d35a86da2ed7b3988334bcc431481c6fb04bb0d118f98bd748009
ze4e724e0236708fb9fe6900242138795ce5a7c029faef7d60241cfc8bb4c335048543cbbdc8f39
zc3a34a66904c08c9de4bdbe0f447b8ce95b33ca569146ead479c254cfe9399b5b4f87c176b86ca
z93f048f66ea49636a90b9a6f39cf2f69dbd6422400f668e3323e1ecfbc6c5dc5326228564e9ec3
z346191b50373183136503dff0c4d1cdab4679a7ed5a6dafd51537a7a023f56af1778d7158dcbb2
z9cf113da154d36b11012dee66740cd7298e3aaeeecb4946263df8a1835e97d7e83c2ac24d71bad
zc237610ac18531fb5a5c33f4830103e7c0eebacf024217a7561ae47df6bff682b03d111e8ddec0
z1aeea7d24134fc23ed8469662581b44afa45eb8a27129c18b9fb309e86e125ab4034441da66831
za443988602b7c8344852c4c45992c4b110c47cae9c894ea9a0f5c037ba9318a67cc8496771154e
z2b8e856ef0cfb108c3fd2bc172e112d2e77946f4b066617e98977d207ab4134fda345695be8c2b
z04ccc4ebf04041c0d59c24144b490f5d9cb674b73cdfd8f560ccfecc37ae21cf7045553946c68d
z65c0155c03f2f4eaf3741ec2a32f6e04a6e76d6796a5f8d934386791f69649b3d504770fac43be
z61a153802175af6e5d8d0e848b4ffb9a0c4423b2eed8cf35e09e464eb3db4eff6d5e6ec5161ae5
z808a9fbe5abe34184ecc267e0dc4d17df46dbcbe50471d2dc3ad0f5898dc2a9f9277e96e8e1186
z9821b90fc4840a74dc6c5a8e64632287390b9e549f86d67eed1a1551c83d407221b6fe1439c717
z4f60c1c761db559b6b59de1c7ae06cfa2df645fe42e8f19dd0c3b0faadcd8cc0ec69ac1cea8c1f
z12282b6afc057eb36c8e447b03638bdd6f2a5986e63849310f5382b7b86834eb837ad9faffa43e
zbc8fc7ef86b125fbe9859907b13f65c83d66f9bd50ddb05700e89d49f0a41917005378b9bfbd80
z2bc61f08793820246559a8099706c75ab678dd589f39c61e714b92faf158d7ef640b07b35d1322
zb654749b1a144fd96787972a8d6ae4ca55fada059c83344dd3be66b9bbe71de8a13eadd79c032b
zc924f1d7bb8808a1b97731bccd5847c7d3f3141dedbb35a7bd1b2214c9d2b5bf71e7ff3cbb61b6
z1b9e5d6ca606b4ef09caf1e111887000c66083fec8bef829afb265f0cb6ed1b40e236087fa0190
zeb054051b468604c292a0fe412d1947938ff588224f19d530f1266a3f58e9deff3918019ca7cfe
za19094a72c06d632b7c6d433869e6e3467ab3ba7ad87860ecfe5b226740d837578f02a27b3a012
z1a1f62d359fcf086aeea851109c085b60262ef4d3c1c8efe37658d458a5784c9a14acb57e6faf6
z7e47c244634b4c56a3cf2797f0d6e3f76c33b5a87f5d16c42145a4936b836305a2995745d47371
z617a228362f34904619b5d6bd77fb04cf8aef09511a005ae6fc0dd54182095a0bb30d11cb06a07
zcfbc0dd291ebb06bf5ac21e3696d85ddd6602db233fc754fbc7e702848c394ed85b5806e64a295
z5fd3f2e1eb4a1ad01a6497f7f8d5d7812301c8be2931c14216d8fa477ed9a969ac57de9a7ba8ea
zb6d4bbaf16656dc4b7b92faa476d3005c7e154fc68e0dcf8d0bc3d7b23d38269554d50fef7f003
z6307e025a79b0aa577b52bca560fb46c1b272c81f676927f6e0bbf6e84ef43c9772f4e3e3c66d7
zd36cf86bb7d1e508bf7b6972130e4b590b10740d3e923f1fac76a65119a4c38d7d99c20eb29e24
zd52c592f7f6c1de6fcd40b32cbf2d5f2e78731f01795ed4d6f263f214f3966094760aab338dd58
z838f14b853ba12f9828fd158824da0f7611eba05fbf450c0c9d4b0906a16625aaefd6614f1e48c
z7c4cdd88f8a91dd0f84980806cec879d4ba9de98b745ca7056c87aecc1513e9570052654704ab6
zf08c964591d55df296029ddc7a01f8d2cae5162ee808e7a9b2dbd64515b88a1e6fa457f197172f
z9ec7d090612ab231a33651140c56d799ec671285b25bc4ae347709fc498db7c2a75067d422a724
zb7d9dd4becc6630b0ee693b3b86164e881af262f0c8361a86944cf81b0f0c4b4a05afaf58fc2c4
zb79381a9457ea43042abc6c720201da63db7bcf2bfbbc417ac2dc8a8a01b48fb707271a7900184
z76658d194ca8f903c1c0cc354efa96c64204f57dfdac4ff5307a524137b04bf32dfaf3419955c0
z3b745d2cae4013a6ba5745535699f05c0ad04272cf875ba0a06c490d80f9a685c5c27aefac4204
zf17a0fcf59a9720feac3301b11cb2dd98833ace99535fc25c4901f20a22fbe348821b7c4414f24
zf1fd14f0353caf57d6b117cb74e23bc0dcac4b20ba1e266fee6e0709a8adee2584e1c93b2dd5fc
zd8977b89d3ee1bf8135e48dfc13f56f6cbe9e86dd6be1145443ed066128fc9d4a3714ffdbb24f9
z42c4fcf44502c3512d07a9fae397e735493d67a85d6d417222559f4212228077df0973b58ca8f9
zcab2cbe17c678c959e6f71849d5fa011e69464e75d703b856773e76b5380243ad4f881416088b6
z69217569500e40b0bebca0c94c2d4da53f0b825c05e154fa4cfb9725aef5554959b64a812f84e3
z28304218ec7e815271b00467a47b9a7db7a0c81b6d90481bb814db4efc88bf0c2b7e6419c4a47f
z2de6648ddc744ae36364bd071657ba0434327c3d7d8eaffd6ac78eee96c98958b1a5408fb7e28b
z9078dd0089ba9b9cb314c7c06cd5a8eb5099aac1629caf213fb967dca8bd3778b9643557a9206a
z19ef38aad93214d7502d938473b8f2bca05e6af9885f30980b9dc50fd21daca265c9f79c5e3edd
z1eaa405b45773f789a405955d0c1625de2cd0d1e9a4e853d43aab253b0491ee88ba5787a32d188
zb61a56f2226ef13d07ad925f61477938917b18f32e17be5085b721aaa9bf01df356562367ff5c8
z5a19e8a984d8615f1a6b1f7252f14adc74deac8ed819cb621aa8d2a566d6b640cf455bad2ecb53
z8bb9956982a1c8d559039d9e838ba63aa200a6fb27217fa4a88c2a530ad2c0457bae93132a8eb8
z57d8f63780e721bd3705ff10d757bab4cedd15068d84c5280af7bd1a424918a68163b0cc849c8b
z7b32737c4dc50f92103ed15eb23f0bf553a355933b845834ff9c877753344aae05118b12902963
zba75859cbc1bc13eb9a55a623c18829cff772e349f0dc0d4d0c344f5ccfa40af0ade5ca407a018
z8cdb4144220024e37255ec65997e59c1bbbf339f252c8e7b4e920fbf08ab48be86f34247ef8c07
zf2f3a876f8a45a30194597e172124f13db0aec8b6f995bf3fda809f0d2fd04540e2c295b7b1863
z8d546f61e10254b7b7fc8c50b6218a1a1657e1686e099276ddce35aa3922b998516c9e859d428e
z455de32070605ad2cc82dda6c38f8754cd77209d1edf20e6760e45f23b059a244ee1dc87c2b6ce
z72d30a719d4f8a12e38fafff2714cd1a2ef5101665c5bb6ef49fe7ff0e9ec2668037ff9653fedd
zc93a2b957b38028dd9033e4cedecc7fb394f1ee2824e0e807b85b2fe55a59dc68d0e320ec41ed5
z446ced12b71e6b6996c9d9c4c4b94ada60852d902dc88127d8ede43a4ba2045ef48bafb58cce3c
z28d7fafae5570991bb865afb966d21e8bb2e2b3dececdbd459bbd1b84ea99a5ce61d98eefb35a8
z9b6fd4494cec854922b0d87ab6ce1e51e16fd2f0235612c0d51b4fedde0d9577080039657a3f8e
z74aefa0391e3e8b5f0adf1434ee4c45ccdc7c80c370df107f513ffa55558a6ce4fc39a1ef16344
zcbd038ec4c4503e4ee1beab94c02645ab711d75d4174645590eec4ed4205c055f5b03b8fe34ef1
zf63733b21558fa0f381eab978f43f76a0751ea20fe65cd90695ff594ea607d4d8a2598f3258418
za4214720e9c7d648251871dca4e86d062d46e01df416667e5712eb252b680fded52d40b4f3051f
zae686607e78d980b275f7c9ffbf9e18d11b95044c26ae34be556b46e06ada9ce677888e990c5cf
z87fce3e90747a43198359eb5887bec59381e895abc2d3f4cf31b510e4de0401ca1a98a7412c5e3
zeae6133873bc55f57ab26a4358f92dcd3a679d28351903ff83332e4fcac3ee659ea6426b6567d1
zc9c38b8a6c89e895a0b83b01af2df02f74f2941f1510214fa594d1e356d1c1e45f3a797240d00e
zc1a9cc7473575036fbdab16435ab6e2c7d3177c8bde9ef54015d0e28b4d98aebbb96556e18dddd
z8052d25b016c63ff311f81005c3db572e27c30f68ab475b2c4b0c0bebdb522df6b5039d2df3c70
zaf21d7e14272922eb01604a8b0f397a838e2183a584b40d10a9646dc507cde8f544f2cd78b2b5a
zb3c29e85e42e9975ea1d23a70abb8358dc197ab6b55b28069d51299d7f8c822da14f9ba23fccf4
z7341525144d2a88348e8e2c746b5db2ffb9a4f8ec3c05713f462d7b2a42eb9bb792de3d11ecb4e
z3f5ffd7b31858a5cba4865d19ba0ceff13c57fe32c0c5e6bf434216cf99df6dda2c24d1ad7c64a
z1696f914380bd7c92e26825bc2e7a3fab45064dab8b427fb55646b9f881299a9bd0803b4a586a4
z0bc9e7b0e2c973a3090e273dcd85416f8d43555e724d55dea2aa980f945d5148a40a936b798e26
ze6c68113b6f90962655331fe3c437da46c96d22fb2f2e2628e0ac25a5db6ef7019d49a466bbf00
z1917e061f76381b3e82ddea274315a381f8f3f3bb43f0fdee07b4c8d0cd85509c65927319a522a
z2a89de523725ae2a55bb2ed806c7155f0a37d6adbc53705de6491413056b93d690df1c25bdae26
zd91dcab442f224b11d2abdfb238687489ab4e5734c863ab77ddaedf86146171923bb0093240ca1
z2d2d4e4886a270df6c231ab8f5561c7ceca41c93480dd09f522a80fb76c0e772e494e49c64a17e
z70c36a4c0050578db5958e2c18d7964f621bffbcf6266cd81271a70b4ecc95b91b3dac6f34a261
zdb5185455470281363e7043a29184fe1a76791f6f680812471a67140933016ba41e2d7cb2ce744
z70cc45281c460c07e359d60c98972c7bc475f56a1adc93a597eaa7bf2f1bd19884ab4af9912982
z6528ec98abdf8e878adef8845a615917cdf7d6d3f96a63f9d14788c2663df678a5dc0bea6c6b59
zd67bc60bea860b66737ec1eb02c5725777be9bd354cfbeeb74d98a9b348d90217c30afe9e4f78c
za276b5f13cd274505c54aa090f87b91c47f7643ebc97435b16de6393dd9d915b2e0d05d59d6136
zb76c8d84de3fe5ab2b18bd1f42864931687a73ff3ccefcd252166212a5088ba64cf3553028b8c3
za59b0091acc1ed98dbe1f7c4cbf54cdde7775f5e59c8ef885eb5f88649237fdb683696576122bb
z9b21c8e0e4b2b9d8e95a2a01f95eb38a84ced5f9f54321f52d5c27f136b8471317fca845f40e68
ze5f624eb776887993922eb1edd88e9ce849a80c8b7da151c6d5ad7ef3404691be437d1e96f70a7
zad72ddc258b362edf48f86a3fa42470a0197f5692b7695a00d137422122c4cd78666a12b084e61
z72df8e52015ad43091f7187811a8ae817b67ab37b47a1c4c33d241bf1ae76dbc7e2da27186bfda
za96265402b89062df2852098111fcf12c55e0ef05cf5dfe2818ffe5a0ae31b6e9ed58654cda5b6
z0be689791d1dd839ec80a399f579bfd32ce849b8ebb78b108262f6fb73244268feb373b195abb9
zc57fd082734423378eab40cb84d1aea0cd498c568cd957c546a13efa4f580d5ca9efb350e0b676
z4a2c9259609da51b7cdc2eb1669db265db3be0232df9bfb020a17c13cf4586aae04155745a20ca
z7113dabdbc2d61fcd5a3a862980dae3a572ac21df32f73f12032a2f2bdf01267219ed116cf56c1
z628dfc2d014101562cc931bd407bb3fd70373eb17692c05cf4ed5b6ea5555522399e026d3f445a
z81697d64da75a397e9bd7a6db3bcbe8943f63ed86bbdd11a561d64ed7c55eb91c1ea9b2271f6ff
z2f69b35f8e75d9efbc9dade978fdb7de5576ea99ad66903c7217c418198fed811bbf20b1e27dd9
z0a2c4b03d392f143d136cf526299f999b35faf8bc85224321ee9b07832f1eb8198c5e7a6faa3f3
zc5cb86e14972a9d67cf0dd47549cd9805da5cd96726b2b199d513b2e3863361a2c2a4cf8e46efd
z452132999482786a9b73e7ccfca734eef5623d783dc27470ab07cdfb93c15083579f8ee9777c5d
z154368794963dcd50d9f1f4fe49bc6a7be28bb8ef474543bcb5c88860962e1943d80911c90bcd5
z23c0186084c59ab9b47813e6bbda47003890416a69576edfce79f0eced4308c01f6266ef510341
z4368dbf78f8da638f94b6e3010538d0e22868d03cf56c12bee29fee90f855c71e2944a11b4bf0f
z5e74e4eff7788fee36d5a73969180e9fe7ee56b1dff4c41bfdbb6d301f88f726238f01ecb5c175
zaec8ee0a69201a02bf6be2ca6268b57d2249971fe19f3cd05cbc000cfb9d0dc632c1ae309e38b9
z8481749e0659b7bfc6accc3b4272790f45b39eadb7442c9768b935697098b8d644277f5da84bf7
zc796655e8fc8a98181683b27dce1244f36cc98e3a62824e9807a36623fdc9a5bca524a8243544e
ze3d84f3b356ae9e6b4a06d63e18f4145f9ab086323e769efcc0ece5dcf2e493cdbbdbb6c2c88d8
z6f9ea27c2f59cf09ec88284d6954b8f8659708a7f57dc1e88532bcd1715cd5376fd0dec723b5ec
z61c6fb811dec37b4abaa70294e6eee0ea04ff2d56ae992a11ea2a8e755d4300c87b5c499575941
z639435e526ffde83b819c00b1f20185bdc4618f60f0640dc17948bce5aefd2be31b830fb3d6242
z570af211edff28f76b563dfc81d5242e44c70c4d9a0b5ef56272475f3c18f966a2aebb3bcfdb91
z10b4f07ca581ed7212e807b793dd57d2dceeaf0ec92ae4cf9aef18ba22d99e005b1bff2b0e7e89
z11b0b3e2034d47ab78c3ae6d89bb21ffcd01cddb3544e496601f55b202a84ca3385cee95ddcb80
z960b8f22b8c15882cfafe122edc77324c8737ef4cb6924c48e37ed3935a5ff59b34e2c736ade9a
z0b9221519c13f9e86a0476fe805b69869cef3b5f04dc7bec4a004b64aa7373ebe1f10fa7242959
z527bb72e312da7dd3742cbe3b172088eec844d4bc69704c9a7c9f4a0d4cec4ab1ce44eef104780
zf3a281ab70295c43b9370e544b228920e4662c08ce766830d7b55066febb7619c8c82253c01467
zee2a00d40b1b2569d58ba066fc0955c7a46e634b0f71979292d31d4f1383f26416499c2c050f22
z48334146bc74a39612970131981acad608fdbfc45acd027b2093aef7c13310a31e2ecac32d8c09
z4688391766c27dfe4d3558f33e2397f9c8171b3a94ec395a3ee5b99e1b1978335b7095aa04af3c
zca67fe208b0a04f08ef3b1fc075aaf32ee3522057e0f39e4d86ad3da8d1c2e97b39deb5e742f8f
z910268cc33f1ef1be0edb08b6f8be4efed52a1a5e11aa5de0dc01a98d45cc71fd469dbeef6637c
za44eacf8c167a1b5ddca0d4e045d41b70861702c8a2a1b7d44aa1bd325b5f5305adc610403028d
z2618b9e61b4df4feb49d4c0395cd3639e8467006b673f7341ca682556f5ccfc342eee78306fe90
z424177876a998868299524d612b5465269504268a31da79e16229aa2350524d216669468680b5a
zd1f6b63b5530dc8a363b2754fee76bdf5783c41c12ad10ca91180085a7d0d6edadccae33fa6ee2
z8d4ffd61a60161b3544a88b0882ca13292d58d0709f0f41ff7ddc277b15b55a94d7bfcced81b25
z3f0f09dbe6adfb40459278d0e43786a54b8d5db5c0f8cce47a5275ca4ad073fdf172677f155162
zebe2edd7ce029ec6ee010636a87937893edfa2be91637cc0982a1720e43d5f3c096373e6669e00
zb4f00b2febb175be0d6d950ed74ac8a39be487d914ebcd1dfc3f2f20dce49ab750ba204a378cfa
z1699be35dfbe5b9b0ab189ce9643d3cab33521dadb01080040f28289bf70b6950cd2d995a8b1b8
z0454ddf7b5b3bdfcdebf33c85ecf64f23c35316ee8457d498dd3957ca7ffbcd59eda0f9a05ff9a
za5d5d356967abf83922e4699014ff92aef726c6b3ac3fdf4b9ac0240073d928b72369cad6bec7d
z48619c6527bfcbb9081b063bcdbd4bc4b2f2eff8043fb5ae61375b4546aaedd1fbcdcf55b5c2f6
z9ca6aef9d1f7c2da31642300c0debde2fa9a3f97f18121b038e00b0c6dc0f1894b81081672d6dc
z525a779cb51dc49f11c801c69777043e6d659323290da420221951eaf50fbe4e91bc4ec818ca51
ze07c3daffcb0c524fd06fc8a41204d1b8e634200686b1d9f6b31961ed1a6602e6bf143a08441c7
zcc17fdb57b7976c6acff4d79264def0584b21ee680f3c8e039b1792aa241a63d71250f6fa7d3c0
zd786ec3ecf46e8951f177d8fc6674e8cc17cada55fa5e451326464ffedc45c963df1d1065ab2fc
zeb19c05e4200cde5495afe447ddcf38b472b91b899264734095e301caa898d897299c89e4dfd8f
z803c2efc44080e754a2f9187d94eb386cc5fbc8f7f0360dcd75f890fa896ab29b594e2ec53c36e
z8a955b15914458398b88cb3e7cb2bac25927c5ea080dd4b9f6f3a1c3099dc99c62421a36d510b5
z1f21adf742bf3156dda20bd4408c7b5cf19e52fc94929d510d8c272a4ea7a9c9ae24bf1b40a96c
z5065312a481d9ad24029f9fd28498a9d28f896a21a2403659f61ba33b454b108e16042ac1d5697
zfc32d1dba70aa9a7e68906ec159f9918c8beecb217047e9799015bf490f60a145bdefb2adfaa10
z787e20664b60c2461ebcec0ebbc90b274670bc170db1f14c452839e2124e8485cdf4e7c589042f
z27adb8b9f53abc233be0cff544862648c6b18accb17121362fa2e7a07d2c18e51bc9ba0c43bb23
z4a08df0350664f7dcd0e1092882d3a97c88cef9346c2b3ee13cdfa86a73895fbbcf27e3bcae479
zcbbbdd7c3647d06e246490f171ecb874b4774a6585463e00c48af8905bb7ac987884ba9e8ea9a5
zcf897f6f49297ef8d3c5ce8dcf69e0a9d5454cd52ae0b5844438b06c7a7532060a978e5a39f3f5
zb0b59485b10100e21949e36f6647164e0d46e723f09570cfdb53fc87c561cda6927522c56c3c2f
zd5156912abcef9ea7a98fa2093948b61ab4b7dba08df3f12afd0fea31631f5972476db35cefb09
zf64b94504eeb2073f5e0d913aa75beacb90f6e3c10b478dfb5c25d0feee7a36db3be9fdb3ae1d2
z9318838e73f8ca3c71fbce5143ec4829dabc195a4342a95afca29fbbda73bfadf21da16543b5c8
z35deb961d3ecd028f5f7ff5dc107751f0548ddfb6bdba57a1bfcf3999f4eca32604edee5bd57e3
ze2b83408efca9e0dd27a2bb5ec01e875759163791ec6f836e5f300a189b76c41010a481458e471
z4dd0cd88f1fb6cd6ff34b41706e2947d7f16d6ee05c1714c70cb5e429df2ac0ce9c0c0e7ecd42b
zb2b5639934af2d80bde26bb74818a79f2ebe2bb7ba155723f1c3ee021f010a54b9cb8535542270
z35ff92fcefa940663db600f0708fdf57c1be4903013f291371b71d8ae86f75732a2a878a1546ba
zf15f98e6bd6ab16503eba0549eba0464087c746ac90c488fb7392e64fc66750eefb825ff45d5bc
z733945755e751671c25287b05abd6b259137e7a81ed10e5dc492062f78fbf43e15c9ce4520eadb
z8fe623b3a023bd542a3782549756d7c10eec3330e4e97c2de86222267d1333a7fc17b17c1a4d9f
zf74bbef08b4dd2e1a75b3dcacf6ab0a5110d23152d3cf123d7c7527277423ec65109b95ac1b906
zd3513c1efb8a8dec993471a8c7a91836aec3421ba1efe7516046cc9260a8efd39955822c8d1131
zbccc15f940ad76ec9984f0827a2537608655455d7d5d6cc0706de281c818aeec6188626f5a1f40
zc4a0d8a223d83bc7ee64aa8467e81776e1a1095bedf8a729e4b607af11df73d0e1de009da0b5f8
z50abb42aa0876113bbb53e1e5e1039ddfca943fc232ffeb634ee254eb023d540db79292f48e8eb
zd77cbb4e92702f5bdf1a369bc6ac7fef66d358d86ec1edca4954be3ea55a921cb35ed92b6fb4c7
zc94ec5073d2073c16b2636a39336d2b77898130341dc5a7649a15a2cbb7f34bb2faf1054df64dc
zd7841374a45da59c8d4691667a4809e65276de7bbf178e389f1d3e73cebcdfd3cacc52887cb11b
z38f321542d5847b926b8964dd892de6cc9eeb5c4f62df407e07adc1df2478a0972fca234df4aa1
zbbdf88cbf7c6f0af53fa33a422b2e1b595fea2bd6383b4da9372ff32ee494ae1c4f5cd90ec2368
z3cf5465e2b8406b519d11150ad31a16ce5a23e881a6b66fab4b1524cf45d4034ec03e46714be69
zd8c705be5ae80ea94365b5ba259d42beb3ca06e90a19d3f84524d0c4ade473ec1bedfd1091f663
z7937311409ef83ee2cebff07f975c9222be3385dacd38bf9165df41a8aa6016de3b468d74319f6
zc81c152f2f7ba668a35d2340533ced6bb59c6d66daf8b8fdb39171abc88ae5d627a310663275d6
z42418a24e9d26b48e01b249a5053f2db2a16dba08a59b0493824c915c68cff1d1c25d03bd35d60
z3459a4f22e2a71102ba8bf572522033511102eb2a2d224665f90357a19f3adb163788488d955d9
z3537aaa247da700ba27d45c3d2757436f15fa030e7e307ec2074472f69a833adac96d45c4d3aa6
zf7643df2feb9cc7a0d8d574d3df9bbfdac9d9a9dbd3b44d3d859158b5f981f45298cc99e56de6d
z4f0f8f4f0b8c0915b87634ea2912a3991ac55671f376417c9d734606ccb9bde27a0037e0faf3dd
zc51481efdbf8f6e4b23a8dd44c2a8a80606846bd6a02f1b29cc8d353a0fa3aee24099996c2e8f0
z870ff74a93c42d74d286ba19e277b612f8cc872cc9cf3e69366260cf4d05e065ef2177d26f0d15
z54e0524f6cb05f556da06d4253981eb2f333ac8e9caa268bc38c0e21a83d27616476b0654b12db
zfb43c5f78e91774a36765c7737c5aec6a8e9c3e57afd3f751a5e61477f05e7e61f5fce664eaf0e
z8e46c518dde9865b12a770dfee08b1d687d1531dfae0ffeb9c680855db11c308a6e36ab2dd02aa
z2c353be1b1f397d4432657a5a53cb86b7ee64af4dc237d3f57e7c86bd6b627674d787add7650e0
z88b5f8008408ed7069677984448762e71f79290b76f14a94b80566f01a4e5d62f5668511e92036
z796f4cff84aecafcef2eb0099bb775e0c1ec2a692f3db649248b99b3220a195242095966a99d96
z6ee94ea0c15a87f4acc02fe7090f379bad09d5770ab09c5cd54d8302817fa267735fcd046fe52d
zb91ba9c8a8e12836352c954664afeabd716d189d897b703aacb48ad4defce04ce4d4d374316fbf
zcad679219dfcfacc410467883d683b4452ef82ea5c3891cb43327de60fe6c7e56126830960dcb0
z9b000ae2dd14e4c7086996e021840c3d37301f191457e420b1f5adfdadfbaa2c610175cccacf9d
z71ecd330f3e48c49a2e31229c4337c2b95611f4f2be43d8d53dffda4e5613a8bb2bb84ebda2d1c
z45204ec18e280f5a7bd53d2ea06b572ca0a28e0edecc18a7a17cf2563ada5950be2f1eefdcae9e
z413ef8756996badb773e8bc40a2ea77ff8e8cd2de804c49ddef2d6155c3af57a5e35efa4e238e2
zcd409f7d25b4be2632bee03ebd9ff713ba0a2fa3764b0a945792a59cfc22392ada1efa1e7efa50
z00bdc471de97b86539cb8e00a5759c76dafa2fd3e7566a2f31956fb53c906ce0271a0f5d034c73
z73f0109f6026c003a5e67f00d5dfaadfd4a12dd25696406a4f29043c5cce9f434f7b6392f79a48
z29917ba13053d042a74c6b0c205e61199df4d2cd5c2207dfd92dfb61714cd9ea263787fd6520de
z9b8514dda23c149153a077e3f079e0b5857530940952af9f6fcdc952d11621e4c22e931afc6e3d
zdbaffea5ba70a8dc9e6ae386760d3c7abdfbf4fb414d2513f883ccdb7776c64c23e2159d24f773
z0e98881d0b84bdade12688461393f12fb040586a2527b52797d72fd85cdb254e8df5be6eb82396
z1579378932a85748e7c595e01d7b084eae424910118d18d823682b867b15da208258d2246edf7f
zaef7c21e57e86f1e121b56f14d685cbe949dd0c98f5e1fd4d6eb56c71ea23156130db7557cc141
z3af52e408df1cd13dfdc1571c86ec8167ede1e9d746e01ba8f376c1bbf7dc466e4d0147eb0492f
za2048056eda13f2b429e801f6772fbb55282e50aeb5db6d4b48fb892135d04509a260640e7afb4
ze0ec4ab52a96bbb48631eb1b980738e8a3b60eba7d4b71e5de55c85594f4e0bab9fb0476f68f6b
z70e26fc49e905a44ad0423fd1b8adefab61f26bd83113d41ca7311799d7bdb70a3968e0a1855c9
z87e218a5fc7763ae3643532ca059abb6b05e714c5fc8817595b34120a145415dcc825a00aff5aa
zca79b418b917271e00a44ce25d22270150973b4f890de47c8acfd5fe4efb0ad641f47b415eaafb
z0084dcda16616bae6c45206f508abc6745d0a70a8ff21b8f42b7002c1a23a0b9e3d8d3009f160e
z31b0e28e6a93465a184674c79ceeeafc58d969b434aa802f777f5bf2c789984cc47de6cc3db104
z41476921bb04136a7b22f6acea2b7528db818c3aed2a404236b2fe8ba14067f2ee34b36af00b39
z00f30bc943d7c77bacd6a212ea087e66ceb2dfaca64e7e34dc47edb47aa2e46b3b387103c5bea6
z01f3881f09fc4f6275eebe245b4cd6c7a2209daabd051f56077e8e971798dd3f179a24d9edfc41
za1415697551110a988c65271fded2edf7799ea073ebaa10b4c5aa527a41aa40f6b7b3e7dd88b56
za86893d2fed9e8d233bc071b1a7eb470274e2b03ab96884e544e99f9610315ea9cb053151d24c6
zad9bba8d646b9f85762f8e7f9e5af05ed00c08151d006656d272651aa6027f3c61faf29b3fbe44
zeebbfab5c7104ad3e4d3a6eda64f0dc4bb68707997e3a7fdd7ec0c197acb10caf41c592f279ef3
z373ef3fcfed3baa87cd498be1cb8eeb540898ca2c480e7b2d18fbb4644368e3fdf3f7766544706
z2b82cdee7bb2d352fcb91a10cf3276b38e95bfd740706c0f279a1d0e4b214d95f8f3eb7dd4b9d5
zabb23ad7794c632d127dd501740d92a6d21353bf746497e39e53980e53a8193bcc74a8141d088e
za6e0abad105af35d46782d7286fb5574b63cdb4fc9dd0baa09af1d111543194876668fb372189c
z6f12ad24e5ff6576d011572b79f61b11077df7224041efa486f23a5cc7c322d3bb1de0c3c27737
z75e06e08f0fc5ebb0c120aa70cee989fa6b8758321bbf6f7b4c931b234499e358e8812ff2d0b26
z899a746b2aa9c66dc4d402fe391cfc085dc3054ae19aed04168d7d223ffc84d0e653cf7eb53f6b
zf2d7397312489fac55dfd9b9dde1204e89d3b18987d8a118865cc0b936f47d469ceac99d1bce0f
zd6345a4c199e54a511e7dd8b37e2ab2c73b9b6591276b98860e9a1d151bdfbd36c43c7c0b337f2
z4cf9e91e878d2658588e3bd70e21ea6ca423ae8a42b714a361de4060ab099f7b3215f0c406ff4c
ze48d633c9088f1b5e69ea48fa5dbae1de0921a7b1e01745c58bc6500142419e971b03840a6cc1d
z8d4f388bf6f127dcae98dc7a220c705db636fd6777ae191283f526603e1c454199dcd484ff7bad
z31be2b40e59c0def6c8157eaadfaef80999f3805934399facad60f5fb410d5f1e5db54414d8fbc
za3065b60f14ac91d7ba392640fef1fe406eee075fefaf0f6685c1e02698985655cca7f5789dfe8
ze0a100d177bbd549933829d25bebb655ffb6c214ebc662bc62748f58c8ce05eb5fca0ce3c2d546
ze9d9e76f40be0cb3e2c8777dc3bb34f1daef56b6f984468428b15accae60b703af266be7695b06
zbcbff2558141e91c3814820dd5e06d2a6f3c42c767a66b107f797cf1921626f34f6d9d9c5b59ea
z376ad13ccaf693d7728cfe5cd213b24ee1ea9b7da4e0dbffa4be8f66541887d9f1bcf228e93e44
z19c12dec6fea39e203e0533e657d9a54380a80b462ae375a8f82fa3b2cefd178e9832b61a789bd
z691c553f8f917000aef70587f7cca50bea188dce2d3c8776ab58a8c2361f38d9794bc5ab91c018
zf33e15ecab0546ddfed7851d852a22628fa1e6b913747ccbbb7dff4e1434277db88355a64770e2
z6a28442c174c74a8679509ef610338483a977b40ee8feeb71bb89d2222456955cf2fd69859bb1c
zaa842541ff2258742cf540741afa630183389bffa5458d8d1d30bfb5a3e56329480c141899fc75
zd9a59870745915682dac714bce9da36dfc2ee4dee414dc43f6125c99b8c06829bec46f65487c8f
zd9a779033887004be2073d8919947615f8b0b51ba3777ff947fb2b746e9c5a37e9d493254883bf
z5e983add0426aee69fcecca5580b36aee44d2a4459d3239d5951972587b5867a5cc2f261799978
z34789d2741371637b612687f83784e062ff6dc442dd2c27c60a5250e96cbe089370905d5a948f5
zbe253fd5b266a595b529cddd7b86ccd4030ede3c94416a90c064bd31926e51a45330aa49e86b94
z7291a8403cda66299fd2a90473917ffe097126f94242a871204981713ad97b58a2dc7076e8b502
z723a20cdd39d2364839de99f6a1d6a7b0a0f2ed44592c25c896f1549c44d551dc160d35a4b03a6
z31e7e43d125ec80a507289c163e5602bff3781ff606c78fbb759b8fe7593041c563bea12919395
ze7c9072c8af9ee3118edc0bfa71deae1f2eeaa846c33d5a6d2cce4931d00caaa744633d11692a6
z4ead091a4f9ea755ab2b0f3062a5ec6fcb28ffd0372faf834901e010bfe21ddf09498ce97efeb9
z86b89fff05b0d99e7b79cd34cbe806d97f2abc7fdcdf7b84c46c1dd08cc17e939a52ef70084187
zac5aa1f59cff1effb11ccb403523b0f6e93e4db6674e04e47ce9dd1aff632726deec4f3f450cbb
z108f9e36ed211f8eef12310b26405ad552efe9488c42dc4453ba3dc90e46d65334158be8cc137f
z94bd043fb0117001aedecc5cb849e4475761c2e0042d45f9bd6184a1a9c56f7add8c16c07edd98
zcbb75a96d1a4a709a946afa7f59dc3880b581d739eb253e0b3a1495111e13a4d691bbdec1ad32c
z724421e7b186a15f383ab341dd31548deb526e66d4faf527b813522dd3c344d53f4456c5a53a9d
z70bbf6ebf6e9dc59554f2f43b05719b0de6226a49dbf229c84996a8710c691ef513be321197789
z5be74e9f759cc040ec818e49b548b81481f7064655e5380014a15997d97be8957a4f376d648e76
z438df811776439f9e19dde8e375ff8b652cb3d79c23954e46846b6965610f2eb52b5edb966ac80
z0121ccca88a5b85c30c7a983052ab190905a90bf8e186c891d727609decb6bd9c8d85c4cf020e4
zd8599af223521480c1387d8c41d5c3cf8395c5925ae8fc206d2d3dc4dde5829b4c7399493a2417
z04f217a3a2c991b67204134f33bfb6f62170ec5700187027488408d342313f393d2923b2d119da
za343b45615044152bc25a8fb77b91495b437d0f9d17f2b284bb51d302de7a24b876595a43d2de9
zbcb1be169d04974d147ee3a35022b49f33eaec3358af179be363613ef0deba743ee67cd04837fc
z3b715bb7f05be1f79dab7e1e02bd4c1373fc14f2064af3378298e0a10d5796bc9f588c6cc94658
z2507a97fb02a4ab74d7f6ecbf818207aa471138ecf64979b8efe8ff6dac0fd66ef7522540edaa0
zc75bfe99f2fb52ae70dc604a0ad1de522a9a9a5bef628db1d2167a368f1fd2e3fe5f8b6d00297a
z2e8a4e7d446985ccb98426169539d815d9a2a6a2a621ddc8464531baae50955653cb595b3104fe
ze9b023f060d74ee58a8ed251ab4f6c6451de2bd1ff538eca4ace6f76aacdee2ce32f5167e49db2
z99d85759dbc41d72b3bb2f176c21f2b2b3804c6cb64028fb810571e5222906f59ae3d1681661e9
zcc21edee7677267c3a872f57c707adba9fae743e5bb32da500301938e04d28233fbcd36ae10668
zfafe31d7bff4722cf3a8cb2d2e9af9584f5d67005125ab5dfdafe8651e580546d8346d7b06ba3a
z2a5d6a0478e629fb95003d2143295059b14487c445add8e69f8b9f9e830a1c6851604f206b87e7
z173d0a2d181be7b464be8c4ee40b3fd0726a23b72c9f26bf9ec09e5a85d411c346ebb81b64a5c3
z2be76a6e86b8a08daba729fde2b220b1b9bc403a0a0689c4a3d2d916f487199b9f54c984b5ea21
z6b868d5ca426059f75c3b0be0c2e93c47fc0b809fc123786720dc8697cc1cc14c3e6e926dcb3d2
z698398cf0695ee74ebea0ce0f4a2262dd1e1dfdab47aa788aac78f52689d6528e0fcf60ca8be33
zc9b3cf43dc270ec53de2adeda324d2866aa19ba06c430454f034662684d894da97f8e69562243a
z74adcee0a15949e43cc12e9d03f3710bb22d038f6f26a6f52e99f68bc4feb18b84526d22b0867c
zaffade9bb35f27a9967e7ab31e6733219265c8a0f1600bdbdc9648f411cb88c5c733374a29217f
zeebc7279536a9a345cb50f814ba0a9554fa4054420f789998f5092473ac2a4298b9aabc1a28e43
zce51d011360a0324cad8be6fb81fe2c73764436cf9b31f5dd852ef413c999b0577d28f4c62b03c
z1e2e3e39148a05f2b0c071fcf18f40a0f5846aa88b95a5485a4ebc26597d2ccd62520194d2ffff
z0acee10a968cdcb5694e52f6873b6d697a937fd9211666f41b12bfab7ec3b24807be86ee979fe5
z7966e155d1297476f0758ae942ad8fc9ac1c94214b56dff347c7b005bed0f969fce1fe8440271a
z0c8ae7879b0639dfd4d5c3137117204db7dce402050c30e2daa6b695ae7e2abe8f6da0b9283aa1
za669ae59bdff01098822a7584b549ce805b41a8641b19b0161e4c8fff8cadd5a3ffb8688e007db
z4bf5e424ca0059a5c804efbdd3a382cc4071ae3e04149426edd535d825d8b1fce0a08982860bbe
zea1c6a7b7612119d6864975e7fa54a494b7b692ffaf4de75a4bb63271d6f44275391ac76f0ed23
z50f36e1b02fc432349602f8539e6f49143c7eb5c825f93fb850724fa0f8d6d6848142a222d6db4
zafdf102c0c68a975cc4621a050680eba597e26b1ddd2d395b3d5d2dad2128f0500a28eacf216d0
z42c6c1489eb8ba93238114841eaafd6960303e4f4a114aa1e670508f3cfce77d3219eb794abf61
zacd20d5e82e4d66b707af3cad46c634b56685a0b3c371a8eeeafb6f9ba764ca9d2eae43af13309
z3a0fe0d69b3d58b5656fbd7ecf49b7b0a722c6ac3d12a764d4c31443b76f46aff2ce24b1e03f76
ze4a2372636727a0db550a54b41b663c56a9d92a60a8c1f43c6ece24731781d9952eba719edf7d7
z716474f69cf673255172430b4d178b1be0c0269d1b4647e45a72a6b9e84e39c9da32a3350f4cc6
z323d046b4cfa1c555c940a536bcb9359aae8b7b67e91d9f39e8d22fb7bafb91d0e972adfc85f86
z4b9f5407450a9f696888d9020e8371b1b283fc2d39b12e2738cb9f9ae7856ecff2367c31695c03
zca0c904ea2cd522c5953b2b5b4ca81ba8e6ea2b6e96c62bed782f6d9e005542bed3dabb562c4b4
z71b140d2285fb17ed80ec768091a7bca52130c48ae82c837c3e2216923622d23797fab71a7c246
z6b38f390526123dc0bcb2b77cb659fd942fa3076a9df9850b4b7ac26c6751a3b63bc9708930346
zf07ebcf9eb965707a226d02976deba1558068d4984332f2e1bc80d7a469507b0bae37df840902c
z3cdd4904643aa80c3e69ef24512d54314dbc88a43b82e167b6e222c878415c7b5b7196c1810c76
zbc564557eaf736da18c051ec7b6e47d7a612c5bfa29e39f406dd189b0fdf620f4750b223bb3faf
z700dcb8b8f94602a22ac502355ad3e619e5aed13a465b1c7a84bd74cb05921cfc6e90e36578327
zdb2c5eac8678f0840772affd3653dd6412a9ab454f098a5ed79084e9da34d994ff12c068029983
z5f8cbf93b311ef52dfe9ddd6f876314cd229e3d19643b8a97a6c69d0151f626f202693ce3474a0
z94b1fad360e8d69b220532e345dd8da1ec1c2fbfb31d334f04a753fee8bb9c94848c6ea4880708
z72b9c616bb59804cd89eafe4ed22665acfa2507a3265c279f2c48940d2ba137210d97e01be757e
z0616077fc17890f49b5625fa30e11f6c0827ee3ed0afd024d4e4ee18ca7229ce65984df999fb9e
zbcb5c301e66e486c7c5919a1cfb3238753b6b42db68b08a8af5b3be4a90de2ae003ef64cf7c4d2
z54b358c0bd95af4999ec98571fb0f59ff1b1f97e6da737ac93fbbda665176d1beb580bb9c54a5d
za7459f7d2a1e2b1262523d7b949761a09812a20e4fa9ba29209c90ce986da7dbd3f55fba5c5f5d
z1bd2b1c50afc6e16668f55f0856786ef09dc936f1f5aa79523d51648c62329c245f773abe7f86a
z5e13a8bfc96ce9c691fdf385c8191e7911dfec51d6c34f6635f7410401cd4724d2c4c525003642
zb1cd4434262885531ad1a18f8d9e21deb7e6129bb1fc8474306694ad95ce47ca8366f6caeb2b18
z308bee0cdd627c6e019295f62f4f6c89922b88adf2e6d546b47b9ebec79ed2a6058464efd5c486
z009efb7db6533c934b5cfd7c3c78daaf9fe045f3d2c4c6ccac10bb2e58b931da159a3f48f7b388
z3a4f862e8e3e6fb758190e2dbe89cc3296b4c1317bc24c5f2760c5915f361d183334861b3c2306
z165f2541ee87be568c5b9fc824232aa47c42e41d40244d9eff16bd7a5845d6a9199f86ac64cd4d
z4e36dab551f1d6912d4a56702ddbed01e049a4ad4ca7b2aad91481e1e2160f69f4b12b2818748c
z37e797cbc73160a5ce72b3f42d80294d1af8b1d072a7b36943223b09ec517516bceeb650093f37
z625a360f398cd9d5dbd85fc9b072a72f2045c4a634e85f811beec9e44c133ad7e1e27b9af9fff3
z525bb12f6691bf109e3c8a50bd50d15cef80332093b03eee916d51d7229d171a92c472e0a95e6e
z521b0a2f6c8ba3fdbd5aeceb6d62332fefda2598bd842de4043f65665be62d9f9e3866a2e6d10c
zd5fc072d3a12f7667aab1d236e76351ed7235cb37dbbd23781e5461c84d0d371c44a7ca8fafcb7
z55c3ff403b90f5428975b9c301dbeff964125d816bf4154aae12c361e46a39919e21dd4c501d82
ze4636a29a2462b7398c1a4f3a22c0a3b7502714890306eb6cffd7b290955d1604d89ab70fd571b
z8cd81bb5090707ae811e267bf0db7850bc6404895ebd7305e15d463121ca0924c190a74dcda88d
za23c4256d9ab5bc5578ddc90a4cc9bf9671fac69cdb3ace9f79be7b6ff18533b438c71c023ec2a
z9d5d8ee1a5d6bdd90e1b46500a95c0c246b2424227250643d54be72ad7c7571998b7db20eed4f0
z5a80a69bbdaad03a89037c305d67df0b05da539e76a3ed54d1623bf1290d6949ad32237a9f88ef
zce7e828414f0fffac7ae669e450c7207e276127875ede0d78e74ffcbc2aab6b50e8c455bb78463
zef3efa0389f96776f0da7fa5a51075cea287be519450f02264b476da4f9554fcf9f2bf91199c5b
z5877ce8178ed668185c0f844cc8cf50fe0e42f32ccb1089469babc210d252d9c1e37dc44dfc104
z5cf06f7b3e9a27c5e0adaf267f1ef00c76d8961be2ca713b45d6b1232cddee8d70bb36184714e4
z1921735e20b23cae90d1973dd31b30d3285e986290ad0f2bc76334602a465921dba2813c84b876
za2fc928d4344b597df41ee9cd2efd29509e1a8051e9b35cb0c6d3cf392fd8d0d1294b4354eead1
zf9f27b11738d8527ac1aa5ab9aa6c912a1e5f8acad3aaaaa8a3bd5b7026f6d67a7fa708bd918a8
z89c282c2fbbe230e4998fef72fe895ae9e156d248e49418f449446feac6d517d295fb4665bc3bb
z723fe2cae5d9d3085c0d3c00943820c697e7405c4115c35d58cd0cd514d80c7f68f9713ff2d979
zea10a61d47ac2e4f902de47d20b8b9240b89ac398d9c83c66a252b7a248531f1704537bc6a10cd
zb1d3ba492c2cd8d5542df99e1e252d1bfbee2da7ccc80226fba1c81a12c881d0bdc3805561d9d2
z11ef67635b7e5152e40f5107661f2ed72de9690a546dead84f6d3e1e6997caac269f499c43da59
zd970bfc5582a6dfd889b34876440a11681b9a6cfb47e836154d644336dd122d5bc6241bec486ac
z660c69ab6f90acb3dc32f202477d6cdadcdf90d31e458389c5c4e7a8c5cbacfa236f249d015e53
z1088370c392564b7362c3ecdd661f6db03460f577577e05e6daa2ca7b51cc1ba8d67a562c2c6a8
zc53cf50cc34d19445dbbf9cfb9e55cb7a96582e16d674b5a63295cba8b35acfaf3dda13132f2b6
zfa9509b3e4bc92b03900e74d6db1bdeb079dcabc2b44bba7e0ae206a596e4d0ccc090400566df9
zb20a53a5f952958157779cba9ab5f254bb5408c1b1bb466f03ea249e685b801c6a9b583916c787
z98d8d87716ccf5d17cb81289dfbbe67e87e24c70b263ce523d56bbf91d95722bd109fee2da2938
zf4f02b52b379a5ff8a7bf936cdef2c33c83986f37ccae3ccfb4c72a84523ed400f6a4fac87d52e
zca7d986636cbd1777bcc4564b0ca9e80cce14810a87f3c5cb0b21424cd970242fcbd208fb159e3
zd3b326e3b9d57104053d687c95ec33733a96c2f5f772b6241027318def7316e081e62aa58f2bbe
z3cadb297c42da48e89e02bdc971dd0319f667ff0cfbed99a159b98f8c7d05a4ef14e1af67ba2c4
zdefa073bf7f8280c04f2ac74ae9ad994914c7d74f8c1e984825d6df3500414c8da0be7fc82d369
z4544b35ba481bedd5f8ec68ecf2348a4e22dd608d6247e25a3abb19f0b6e95c596025ad311a92a
z56016d84f6f9a070562dd2409d65c71a047bf0bbc557ba5226edc4bfe1d86959395334166d73e1
zf6adbaf15cbe1a0dacc5f1f4138eff2a846ae419ffeca4a53020012bbcb02213a0cddbadec0fe1
z7a76ce0a6c0dfd2d14e18f563480bc62ff5a5f149cfa4575078be3dd86969d2f3b4a3a2a72cebc
z05831e036afbe3e8d72aa65e17d870395b7d3866b990adf3db2bef999a2c63ac33af9446e2abaf
z9fc7f03d32cd4cb13e5daed6729f4048336fbacaec46c33a27a40420783f85aa15ee2ae792eecc
z680ea0066e868da184697cf7c2768843c9b6603ea13531e5f03e0d97ce7ff8ef31e29dedc58d4c
z923a02669281c1a27f643e49e3e006d205ddfdb0812a0e9283d5b70c05f899c7ddb51c9a98013f
z880e69a361da66f550b041c9a12f605431aab11bf2577c5fa010e834dd96d372787ec942af478d
z3f83dca6f56145d2320cc0ca9707646425a2560de698756d75508724b0a5bb9fad7093b3b8a4a5
z28cfb7e2b3c494ebf6243104140e8aa3e02221770f722d94e61f97e39c8b4d5358415fd1aa9ce8
z9191fb0ce4119984794923ff2f9862dd34127a224707813bd7b077f0caae0347399d8ee7a96e09
zbb5b1cd6ee664ba1b8b3c8f6e413c5df1f5214aee7365ee8783a30458be0867aed3f9f8576153a
zf8ef6d72dd00ad7f50ed1cdcb597e707b6cdc84c1a67d9d7a60172ceb67be14d9d290e421ec778
zbf0b2ae42a4f8c8ebbcc181144ac7994d011e73f763788eb4fc75f1328ec8a2718e624802964aa
zeaaca7691dc1f0158abcdaec7d3616292fd56f444169bfdc2b62df1b2979be3ef858968daff496
z576f61fd7cc58d673976b2551794a41418e98aacf70fef9f4b8ded1fd8139616c8f4f8b552d4e1
zf7ebad48b54b6143d642d52c6767a7987e9c31a7c9081649faa6148625c74cec63ad4fa564ce45
zfd3918b7005c8e1fbbe369346914dd28b7a19de7818c9193ca44d055a578826aa7fd8bb5b30e85
z016c04926b22032a46b27e34482ae0fffd9862ae7500fd42c9cf0f29c466ea878257eaa208dcb5
z6a3254af95459190d8f03c7eb5576270889f9b4c04ad4cd3ec30ca9aa243b91184e3726955dc7f
z34335d6b5515c650758ad1e4ea1915898a9dcdd6e8fe6bf8fcc57f1b7caf14d4bf9338d2be8f4b
z465e993739d477ba9b89260299c6bf46e73b3bd1eed66507257b7996ae568c89087d83dc6fe963
z2a1ef63c81e1f4363d6a90527925721de60a0197fd7b6e9a4125dc6274da5a7fb63228c048b586
zb2583e1c67941777dc2cead6c36d674aad6771f20afd0fc4bd8e5f1370898408cf285f634c9186
ze8affd6d5a971ac32c6460e18cd162f1e4690063547f424f7fad461917cd18312f4c8d7e3b28bc
za0f0f66a17bfeecac368dfc8f2e99e50903daef189ec6b74d4b9bc63f030a15b918931b9fc7632
z7e3da125bac3130bc0b45e3d20bdba8a498a21e4dd5b00dd09432a4b30a6144bc326b54d8a5883
z2d7ccd201c5280118ab8b0f99aa487645c641378776dc7bc97ca9c52c9ef394884237d64756621
z6216fce2bab2cb93f9ded92a0d3e86636280fff87018cd7c81c8648f9e1910866baf2212a56862
z514612d2c2bfa104a4cb8098685de30edf125c7ca4f7fe439f33139caeeb1344e2f30d7d64001b
z39427cbe80798ff3fbafd83bfe745f3109e73fc82284cc51bd0922f271c010648be38e1c6c10e2
z05f67f5afb0dd356c34318e8a39289539b36dcfebca11c05c5a9241bca45f509936edc214eabfb
z4f6118be9b8347848274ab3c37cbb9f567994c0c6d3c7f5e8e3b48691504dc9d858873195d9ace
za6738bb6ccbcbf359a8cab4140a6982885cf984f13b8fcba409a2252269425bb52ac6dee1d89cb
z782cbbfbda21f9c59b569b585e8aedf702c79c79c10c1f19397d2ef9002d88777c36bc763b11c8
z609bcfbf2bea9c310eecff3efb31e8c41a093b0feca7e08d27be75ff21b443c5d96a4474f07462
zb6d5a58dd5995bf5667cfa1a2f698d7f7bf859f08b3b5bc628ca4f5301167327e075f07ca0eb1d
z5714f89c528f88a743ee879d81162a130a1598337e503420874dc16e85bb182cb1361da0da51e4
zd1a8246cd46269fba57eedfc03310e27ec3699a0b6d8d620b2c6c25b9e454d35cd6eb7f3b9c447
za3e735dcc4d7c7898dbd01f9984ac1533cdee86caa6c3143434171e6e54473141d0d3285b511fb
zfd8f2207acdfbc801ab47195394b86b2739568ed95288056d5e5cb0948235c1581f64a15fb7171
z5d53370d3950dfd75959d39bb072f5031eac1ad43eb2154c90891ebf4d2f48df30e5605694d388
z571e43829ed693318746d692c4d9b9db444b203453b03a285025dca490bea1777e4df35fc75dd6
zdae0de4ba6edfde70e383c69365ee764bb9c2b6a75344870fad442d673bb9de8e6bac89bff9dea
zea4276ebad5ead6117e999872f5452563d46bb9d324650de4ec689b618c7b4af4332f3142f926e
z4296c8ceed68c0208d87c899e93ea2cdd1b519ec86765af00309037a9c2345eb1ebfc5a24c0332
z679b011987e7a41baab5602bc39e85be2ff254398a117782c93c0e4bd85277b5fe5fa4c3e80467
z9ad849978ac5d48a169e538f9ff9d824da0e00f9e4ef1e3387691fd2760a30cde77b4b6129e33b
zdd40e16e9ba2bca9dca4986ba9c9fad38462c33014b28df38be232781564e9b8b7ac8c68ea988e
zb370e22323d9716d14e1a058b3e217eb419764140324d2bed31bc5500bfb31883b1d44e128e3b9
zb3cfd8a8eaff5299789a61d87cd4aa05266229415f95678cc366a741d0fa77098e63d820290ed2
z03b09d0e14dcab46012c2424e25cac2d5ad18466e3d91f97733c9498167c559dde52cd7b383184
za5f4b587cd30a75c0a276a022b543e35386fe50c47db8985023e3b55892b6f84791e1e41bbc79c
zdaaab0cfb42e8fc516910f753b0f3b81c0edc418861580ae7f846bc87d1808ada117f6a4d3a600
zc119742623b2a4a17b204fd466d671432ff617a0e363c698e5014e0ef8bab5e76bce8571404b75
z3f329b12f5e762ecec4496a4bebd0b626b1ff33c8ea41c8771167ad1778d7d0a88ce5b3bf91d15
z88172290821637161d7ada9f830f934b0c6ab1c01e072f04761056d2c0a81676be63b467fa09d7
z282bc76f0216bd56eba9c66eaee5a1449d9c4e828827a5422f8a7fefe2c4e1f75173f118484930
ze8a89330b0ca39d15f18935f17d10f31cbdc9f06a8e1dd693f48743b6552a7848d6acd2c3df562
z205aef9939971beb95c09a1bfcf5b8c49081b290093644c276938acfb0d46488da30e044ee3864
zb645c49cf9f84efaf99620a6f6783f2143091e4689dc27c295b69c81f72d9f04c9df32d6aa3899
z4f1d399028f38de4cca86d609e5df6606ece492d3f86bca8263f692819eea5af0c3e346c08cb84
z5a018c435e529f3dce7530bb129d3170a1e22be3aa7a6b568db17ea79212cc8c7fb265b9188440
zdceca513c48e58b6b5657fce1c53cc9872c9ef430a1a23a524d1f1d7990fca0e9528804ed40fa7
z42639074927dc192dd2c825d45d69af940b1c1ba413b2dbc6d6605e529277684e81b2771958743
zda3bc9480545f57e92aea220eb971e7f31654cabab75fce32d7b051aa25474e9d75a62cd02f2ed
zfafd43c16ebf5ed3a7c8f43127f0dacaef6c211bf596596a98350cd30f3dd2be58020c05cf2772
z1770082f00f42d84716f5b6a950dfc2bcaebfb19728986783d63fb1c08adb4c636cf982260d3e4
zbdc90f4805b50e78422fd0554daf7ff3f68ae75080a6b371eb72686cc3f4cb5829e22a755eaa0c
z9456d5d73d45553fed3a1482cacc78916e9a16727ac476fde87366815dacab78125a68f8147711
z8946e5226241035002a32be07738e414579a11b1ff9a35ef37658aa1ab32637329986e271d2f9e
z89e3a01856ad3931da4bd0ca083e774d5de0e568bbaba5a1b48d775479d5b813394034e82059b1
z39528c25d3f443c6ff5a9cd8675c16ca6869f70802f35603ebde9cd978bd9efbeea799ded52362
zc7600b429b9de7352cf754098b38ba7e780760cf316cf197bfe4ea5e4416c16f06569b2fc79adf
z8fc1de86efd769c94c673f6ea82f434594db7d4c9de34ce07962bb860af71fcb8ed23fcf7838d4
z44bb3e9b9fc6eb57f071ca1d04b3e27f5de79625e136065b9f1d352b19ec52a563ca066c2fc281
zba90308baa14dc6e761c6ba973799d967e200d35e0dc6d32382669010071284862bf17b199edac
z807478cda181625decf8544c71d83e5d3d41bdc397559a2239e1c3a377233d9903aa046ace2a23
zb5d6c06a35a43c8593ad8acfc388d4604f6b5d78f2e5e2ef0b64cedf7cec7ef9f892cbb96533ea
z3c806d71f7f194e7160ec1d4b0e979305ece99d5fae2fcb9a3c72785e6fc89dbfc77fe84046018
z9730d51f6b37db182b3ea54174b6db735421e301fb478e659260aa615eeda2908c819c5c86732a
z6622caaae9970e877774fd19633bbdd0dec4d87db1635ef0b7ca83cad4118ebe7756ce7cd4b354
z665a1564ad2e1d940607a54b67873e09b54ebe59af2acae51a92f5c649824d8e1fe6381421a379
z5fa7807e0429f41479030bfb134301b587d3f76d69f228de07a5d19c5d646183ec8c5116032948
z3d7ddfd21164a255e6a85a5f50ea4d8449971fadc224c3db1c46283f85c2b55d9085984c4276f1
z3b130b358de258d38fad656ddb23a4ee518d7e87e63e2c470ef635f60dcd086438d4f34252407f
z0f296382076d872ab17b508295fdfcf0b578d0e8161d25b5ceab369059d05a01ac7b58f31efc19
zbdeca42a159919becf5b78bad1b2c080806422530fe2ba78be6ea9e1c4286c809987f29a00005d
zfae565eeaa669736769a76127d07322e75864b8b29af61b54817827e4aa8c9bfb18b3f8ddf607c
z5dd4939b6e886e7bfea9f54e51bfda6ef0771db1b6db97b859809d8a82405f4d5e71502bd8ea9c
z015777794295bc7bdb6c9be96b4211ce9f713aa81248454b6fef4d9a64c07e03d071bc02f2c831
z08ce07932884da284d41a35caf9bd183c9a8b02d3cca55c34d14d5923c38bf5716494032817884
z0f4b683c1fda2af5050c6bfc86efe33552a60bd1829fe70476345cc0f7e2113a5453d3f2cec205
z21fadc55c3a49499f4def30f888dd85d7eed74e9176bb08d9ccf48ca862531d648c425bf2781f1
z58dc12decf5b0bddd5692ec79949ef72d0f7f31acba89b69b479338c19564ece476aaa80469d06
z9e5ec54174d748ec6164197606f5a0df1388d27549cf9624aa4f80aba355670f197cab5dfa3925
zff8cf92fd89d3c11b775c978b66cd70d744402b97006077d46cacbe6b69a434e1bd18d92b25f8c
z7ff55b9a3e7b510e8f1b1f89aa071b705e87d60e821736e9679ffffa39cdad68e84c7ba4ca3668
z34010a56a2fee5126b5c0156da506fa88b123ca65c7dac95697d98d4db336ca7302cba1cfe69d0
zbe2dfcd36a3e949a6c6b63dc873f11f9927ad34146c0596fda44547adfaa84da3ef2983e1e62c3
z6dcae7f99f6a07e8c81ee307e14a27bed813f1ddda187996c24788aaa655af03fcb8393cedd162
zc6693d98dedeb0b662761873ba0a6e67b63de6daefbc497ea8b0ec5045ee65ce64ed23ef8aa3d2
zdc2469e8211bc266c65e4cb00db6dbaa9f53a8f60abc759a2249d435b50ad8bb22048120a957e7
z88a52cd330e5f12f75a1063e27bfb6354aa2b0e1aff05822bf0139c4353ed3467bb5b30beac1db
z45b7254848f5fd6ca01caad8327b66e0855ca5220603d267067ed10d219e4cdc25e786437fd7c5
z5004cbd8ac0f7b6692a72538934bd86ddac4a570ae60b38e78038755382c0de07afcd82802857c
z7fdeaa7ee49aa504d87ea0b6f039fb69f976f217a7772f36f91d91a3d139a8c26ecae714132b1b
zf733628812ed201398433e2f589d1ddb14989e9ceb0ca5ec003f9a386e8c9de4cb329045ca1f78
z5413c5e889bab5458bad907e42c2ddbd7a420b4bf45971624b04aa0c46c17eb4b0df18dbebf55f
z0e03135e2dd9c4319094fdacb16d12bc9938418f773088f6bdd6a9dd4fb9d849a5c709d239c1e1
zc044865118a3d1d31e99a9dd63d5ae1e159ae203fe0233592aa4beb42b5ce4307d766eeec02eec
ze41f11b479dcd0effae3a4dc4a3a852b5d560c0a1c572c5f57a3eafc2aec35f6f4b56a3461c3cf
z2c5372f8689a18786148281ba5680a89f4cae547532e578e99f91ab1441e22030210f2df0b3766
z4a1d1956c27432d6660279a3815d8eeec668e55b6109b8c3bd750491a74c19e8e989df72d7a63f
zcd822ea7a3b86c30423c96ea2d6963144dcde9fb2a41ea024d67dd4c70edba5617466ccb3ba0f5
z10a5d98844a67e9c6f6186ded4569a54f098778a24f3f822f00ccf4acf074d03abcefb23a02f18
z31b016ef6b5be695e96c2393e08f49ddfc9e79a9045b1999b82d2312111c97aebfc9850febcfea
z1fec802f28f52c2059fbff7338b727ed668a5153cd8fc29a92d5dae0a6c0438c77afbf88e2e82e
z0fb1df9bc4d7afc80474d0060a2ccd273fce6bbc5bbb3658a3eed409279db26ac0afc02f9cf52d
z94c17af0d483c08798227e8e79a2dbb0b5d91cfe00320a7357b2fd48b751b20648687b9194b086
za68abb8a706a6f9ec7ff64ed9e9670a1e930656ef26c52e55d663f48e70da84b5af135b30fb575
z5c9d754b0f0f7515eab6ff695b68eb40565a5d047097f0d4701542263e8192e073d0347118a71c
zacaf362bafeb1e4a0f29e742c31542255d6f38f12798fc602c497bf2c0257875898091beac4af7
z2d469e5caccec71cba2fb65fdb80afa38c113fe5a748354739f47cf94fbb748c7593e420225a1a
z677824a82c1806ca946ae06789c5662c04bf59558372a3f48355174e2ed0babf23e62096defd3d
z927c1b9dd73b3f766ae94a2dc7c2346681e76558ddfa4c9e938543b8693fd17f6afe25eb65c710
zc6388394b0b43bcd82e9d6a727b82238ca2e65350578fb50ed0b484fde855642a2cbbaf0ef7c25
z021c09413b99926c9e831d3b4f791e936885d4d59cc6b20ba8c70c0f6a4f073427497e07b81e36
z18134d7bf786534c88a1c4aace13c693961865b160f444f30266bde363fb84e5d7c26816a8b61e
z9aa01d509c1be15fa0680208fde96fb64e5a7cf01547fa4e793273eb16dbaa037f03d888a56c11
z55b663df10dc959fa832206229ece2285d654fe48d8231ad18f40eb946b1fb274d9c6ac77f14e4
zc472efb1756d68c4a8d4c81ff4fb61d9b688d80d021e82ff0e90152b1f7d83d3812d575f945d71
z5994aee701d0a972abeb0d3c57440509688101c3df034ce68537b19be04402cd12981ec9a356c4
z64de0d6060def40d08c1ecacbdc5856e11eb71abde55e55b43011c471998d102e75e34b0404cf9
z15b54fa6b8cbe8b250db40ce21ba99174a61b0726318f8258b8c01998a11284933edb758bbc950
z6ff00c456837a8e049045f2c60f73be6a1ba6fe5cca2582bb8cebae21c76252df8811c431b3a2c
z07f5baa244ed1ebeba7e19cd374c9104af4ee46fbaa511654c22167187a0f099b9c46a11b8ad76
zcbf0546b8348e96a0744991168df3a629e4ca63fe2bf4940d8069894a7a4c827dad3a4c2481da0
zf974b2cc462428c4aaf288c21a40a45d2cbb0c22d7b4b838a466a817747be688f834659d7ca456
z88b0e87c23699432b1e3f7f9c331d49ba6727716f997e376d51306cfc82c5906b2059c89e25341
z633e368ce77f9810a9083124baa7be382d4af0d501295607f298e46b4f1239132aa9fbdd20cea1
z6c681068c14e3ed9b402bb7a65335bef5a7740a80be65775f2a9c20d2626960829e12423beea6c
z327e7acfeb560122b80d72626f7de7e62f51a673d1eb4c60c61c97d44d82beebddf10ab2b415b3
zc4f6926d0919d8a08b06e5ce9267eb5bf1d2d37d869e65700826cc113ad6d806116c764cdbd6bd
zf68b099f3ff162f5084d556f2a1ffb57a404d75e069e2fa79f1f0dd069eead00877c213ac5b370
z3162c509dcdb9b90b131eab5e34c8b21019af8080476dac1d2efe445aba225f7c37372337aaef0
z55f1cfef7a1fbabb9eadb3f2a0387b97c17e6792bfc01135caafca880d3544a9b1ca399ec1dd62
z3a012cc580146ab8dcaf44494887a474dcc398ed47e0c1d639a9b551ed962c0b7b4995f3ad34c4
zaeda6600a9083c7cca01e9e9e2334aca7f5b3fea0f2c11f7be0b1757d334435d1b375f71d573aa
z6f3563231014dcc16a03b3ec25c1f95dafa4f23c210dd8a14c077fdd58d142157312d469c1d514
z0b1c65c9fc23dc27ddfdc74ba4bc130bbc01e5c222dfb59224527163cb979c533e19aa747ec64e
zce508adeef6e68f43066b1a5f273de7b3fe9c7888ab517d22c05d77cb575f3c397017fa62073af
zf4b04bdce453fdbed3d95f1ac49d66bd7073e3991b146e89ffca24224be1a8f5414ee428fd9f2d
z9bb6db7987c36d0d291a03e01b84433130424eb6ae9da6a639c619e55143bac93b3ad20593ae65
z326dfbbf75808d85d65f634c85aa4fc6a557928b7022fb9d8f72e5dcb66d2bd775d1cf29df928b
z251c0b634ddd9c9be3be6af4aad78dd3ca2b41cf63e3165c2bd67e1700d53b066b95f5bab8b158
z530e29c078ae1f47b54fb001d0ca9f5fb3f4b6645835d9f2ac7a32ec91d5c363800dd5729e23b7
z6e7fd1640ae3316fe346e289fc30f8fdb4f84813d9f82e6f349a25d530a65bced341b970aebf19
zb2c2d16e0cdf0c0367ff5b756de8751415bd8f9c10e85f93cba479af6f6097c2d0fb6c586adfd7
z9ad011a2b66ee8201cf05dc5102793730b464709aedb59fc247653c0fd023fabf44dce70b6c8ef
z4c289dfbfe870c5f518f4f539cc5b416ed90a09ba929b8ea2bfc417e2032b41bdea9d271dafc43
z334bf720ff396516aeb2785d55227630810756b40548719a999ebf83b6d8c07228c28f0d5e9648
z9bc3abed411c5ce278d4b3532e5df7353d4df5fd8ca912b0d1f4dd94015820b82b4fe54f81e757
z816b0c62e9d6fbf3bc45c61b04c44971f16db45e82349f46a468bf4c2a8c7ff396741c44027bf8
z549c881668e13d5f066f4c8ed8b7654d1b751566050a50e2c12def1691e35e51c19d8dc6f17db7
zeaceb31e9f4bc8a86049665afa08b04bdc721a2c34a07fcaba8d6e07a7d6cc027264ccdb66db8a
z20b13d8a94c708fb52fa6ccba37537ed0660b311bdc1312464b20baac167df4a09dd825899c077
zab4b94323743a9916fcee835f1225ab6f0ff0cf9d7e403d4c227a34d69d1628c5597221c2fa451
z2f7e0d72084d2a5aab01bc446e3cf1d58d9e3d3be7492e14f846ed11a2c5cdf115a1d237f8eb62
zb0ea97a76170990f72aeb2544b07e2a29cf6ab4fedf697d8cf4fd5f6d00b6885a452bcacdc0ce2
z7e4923a1bce8ecb403fe08b1eee31f637628d7dc012f69fdbc48192d1517c9eeae4f3544257eeb
z3f3407217ee0e536c9ceb017fe28117f83411d30b3b678bf60ef836af9e8e22e121efbad3460ee
z55a0ed40e4ac9c22c2c5cfb23c67ff35e280a17b8eb109e0f2979a32eec10fa39365fb4553c7ce
z3c99f64d4e171b736da500281f4a6535bb6a388f85a4869216453685be5126777b94bc282d8bf0
z164d3d6843694b43de04e116a790f1c10cc0cc64d2f1ed95003d9b69f437363dde58a62ea46bca
z52c3fe3f474417f2bbdcdb0b48edd17f1901e4a698e6e4d861d1717f1e287c0115f4f1a1086acf
z0f82effe17ee80d5e12a57ada3601b1a17f0dd53c0a45f04f309abeed4164576fe5a3d0fabab22
z5c194ca279991156fea8b33a0c80c820f07ae6d87359f2569ef6de2fb6b5ea5b5fc52430b3a4ec
za41483619021c67df4d2e676bf244ec99fdf1debe77c66d251144eba070dd2c6a76abcb9a1c0eb
z7b34f757323618fb186bdc919f193fa514bfa40f5117b71c26a726eac6a3778b4f833ff4d9e631
zd960d002ed8e18e0e5aaaaa41e56d005662cba2f18dd092baf613fc1d66376a9a01c62b11d89d3
z4bef7b549acf72cbcc2175c5db3e2f107d3784d27f01f5bcf855b592edbd9e6a077e419d7fc0c0
z6ea39c11875f945737c9c853a933666d3d1e6ff885e724e51cf621e87ed9b7c25bcb754713be09
z63d28ebb531e96161f93e0650c95ce92075d563c3c5e70f51f6d0f6c8a02a3c6f87f00d0bafddf
zb03e3a2cf5a4f5561f76c4c0ed0b17f59745d166040d766fd445fb420efa76534aaec2c02d2962
z17bbf222a2cc67571880c8ad4e0302e3403a686a1ac894acf2c9f80f5b2243240cfb0a97371cee
ze640ce6cca20f434c200106df2982e5365bb1165a298bfe705bc9187dff40471366e9b1216d9fa
za38dba27548ce75274dd31af8a207780ffa823e4a68d371d42f57933a466eb693c26394c50cbd4
zb954910b742e7423aac5b923bd1438ee2546add2751b1d63406e65ddbfb87f7beb54f533293e58
zc6b75b025dbdf658be2ea9e2557107f22d9dc1afd5c5b2d32c7e3bc8a0e4a71b6a981ede2929bf
z5ccf4f25c181f48cda300a0aa33fd5525f24fcfc05447ad00c71e99663b7bd5bf6f30a0215e530
z24db2635b8b34fb330383123283d79d0e8d8cd1e216716c79d1be0f528746699b20c62b16188cb
z3b88e6452a1e0babc64eb68c8e8721843108d636793525eaf4fc7a393eb44112b48b8811e8f8d3
z52303d1ec8519d26274da8c92b114050bde8e8f86e22618a3622ef52feae77ca15437f76cb08ae
z28d36c2943f784383d8a3c57a87d308d3b96242f6e14545a271a6f72619b62cf4dbefc42d8fc1d
zb546af1d7a8ad947061b15a0b7136fede9b77b2dc8eff8fb2431e8653696be7e52e02eaa8a37a9
z4e739bf5275f03914f2dca6594e5d52ab9c258365fe3319c31763b893f4dc6282b281ca20f412b
zacda7178aa631048fef78b85d53cda1114ad612c5e44383ecd649f499e35498a058521c17a9e5e
z562ce5a029f422a4f2aaaa549a7a56eee42ef3f86862b4dc035ef174c759cc111801689d6c61f3
z09103872bbc42c790243d94c37054d4e8a2759741b4154670109a51e6356e1578db0f20d90b024
z5f5c3bcd4d8758b582592968274da8de28b87c1c59c1753bb14e697dd59c335cfb527871092def
z573dbc02135deabc46db05fe912ad0701ba3645934e00b61c833a3455d6a496f65274b149ea24d
z54a9eeba22e9ef4d9d04288ee4c229c260f3dbc9704522ae5fcd6d2fd72aa0f933bb012385a16b
z5779d24454e27585246a4897818cb7fa016b903531c1d2c3ea99d3b6adf5fbb6cb6887319a314e
zd31b2a6ac6da830bb0dd1a4c54a852ed4c8446a2a2f2de02c8160241a1a71e0a959ec2ba00125d
z3bd49a788222d01ece47c34732edee2dc3d595b742b781ab5e85d5de5e05254654ecc246975cfa
zbbe6a00634e63d6a840f401d2fb9907d87568030d562ed912d7e9179d1872873292fceae4cda5a
z5919550ebddb0f96328c10666f894ce035f81daf5e2a4f2f416a61c275587c359d04307a3e077d
z7735aed8654e1ceb1714a763d8b19318fb6fab3f177f8fa5b63498e59fc7b95e2f7a071710165c
zf4ee6ec9a991bd9e35bdae56ecc5bff2443545fb2352e472a6d2ecd9f79d5e644dc7cf205f39dc
z2e1aedffe00d073f1ae4dcb50a8e0cd89eb64dedf0281daad026d6531a1cd1dde2589f5590808a
z0cae7b3d1e0f6b5af8071f95b6e020b1c572dda8879648438e1fc9bf3a5a5ecb0848d71e919505
z724a30687e385357727b325348645b3c5ded672fd590a206d71007df7bcba6877db6973033af8e
z726afd61b8129b538660c2a1ac4b4625f89718baf54afcb6f5c8c7102b161726bd96fdcc5dc844
z00917eff4b30414a8be3afdd7a5a20820b07e7640f4261e17ace0c20afba9392c2c6135711887b
z3d582ea8f0fde0ce37d75a1547f868454622318dc67ee837318965b945351653c493883421e078
zd205f9577d0c11013052d57021191f58a89015354f4bbe7cbca0ffd884333d472c937756070052
z86ff9813b17ed290cfcc82130197dfb99d367dfd95d143ba2511a2b138a366d763f9cc6ee329cd
z0d941e26d70374a3e9aacb5d209b8e19a1228c039779acf2398989534096b152e7bfba4162a223
za0af907c8824c55a6dc436fbb3ee60fc03d940f4a4a5bfad0ee9594d67b9be2d477bdd3780e225
z255d6df95c5fbd31ca2d3166c7039c367fe729b21917375c137a814f1415a5ad0ac424b7d827fa
z3a0d99724f404a1982e9bef62fe36a7c620709e52c3d773fe9b38f229125e119b98a7b2bd2aeea
z73e162fca5516cb10fcd5305e0858b1a6c1d312ffa6894f8d6a7e49a3a9e61b7441e5fbc35c5c3
z20472c965d940ef29df8189ce864ab38b4c956f3fbd50912daf313a0c284ebbc292d710f5fddf5
zf572683a0aaecaaa367de1e671dfbc75e5ce2243a032aea6d92f8084e29894ed57e0a1898e6446
z28532620581879f5dc928cf92b978acda19f529d9e52d0a03855eb6d8ed0109d9fbad0ca1c52c8
z352212468e783eb4fb8a6c3d8c0bc233da8f528b6b4e94fb7fdd30ba17358da6d67bbdc0f26b87
zc9a04a332a83f01788c34d805d3d5c8e89ac5ead0a8e31e41f3fe6c1d292ef01b8f44a6abec17c
z66e12ae12f28f09b6016b7b76560162e26b6a1e3e3aa03f2aeaf99b48c0bd25da995c763d0de40
z788f01fa8a5a919bd450ee0cc3bc34b7253aae70a71cedbaed07825bb989de2e0672d15f0d751a
z888305b9c69c21430fb27e4f76e4d55ddbc3300b603b0c6132e1a86a555b48accdaffabb3987ae
z51d1e5b48947ce572b39a5f154424d2604e80a604feefc1df962f4f5572ee01d43b1440192f69d
zfbb5665e8038633fb8da2363a18c4b1b325986b7425e27ed7b4b84e203cedf8e027b6d982f50a8
z1461019e60ace39750f31391612b12172742db488ceff147f9b69c851935315845267aa5285966
z25e727a8a3b076dc3ed8aa77411b901400470c679b4a2093f4bf75bcb5dc849e99d2a6eaa0b225
z527bf0bcf0cd75f746d88d05ec6efb738f27a482db59ecac578eaa6f7b7ab586a2a74398fd48e1
zaa20ae25eea282fbe169cbd03f555e55e62ef8f079ac6a0456c5b181c047d7afdce9972cf9a698
zaa7b2d10e8bf2f7bc2f73ce1e3c9e4c04866d36dcefb60136595bae4f2020840c4cb8ea0df4142
z9593cc67ec4e85ce813d95040d10f56111b8a0396f1dbc03d1d34cd0dc513d16a2dd6d885dd687
zf1818c27b6e04b75e7ce508e7568e2a75b6f8965b04ededef8c80b35654539ee89e26937e1dcfc
zcbb6bb59cd1b9c9f8f961af9f15ac37a7401252163058720a42ec1d26e53df7785b0d0e13b0509
z5c61a30d0db37d26dcf0c4a182c8a99eb391200ba4a8e84d54e4a33a34194432dee41605665502
zdf2adcf37fea8b5735d1b4e6d42055ce5cb7d61665c966904534ca05562119ac451bcd00c844bd
z92b7ea8cdb65c2c8d9b49529535a9fcd724ade7b58b926686086e54e7d14367c7767f1a3c43e46
zd9fa8ff7a81faf17484618a553579335792177b8cb990c8fd09031d199cb3847f0f2697898cfd9
z94a00d84cdfcb711e360ca5ef05a00a49125778d7cee1da815e7a980b089ee858cada29b7418ea
z1b7ade4d561c99aad462919d168c369061b4c444539e0d7e75d9c85d1270bbccff44147f68c749
zf5d555b3794681ac13e52e41b9380d33920be8b1c7fd4923ee566db679233e99354933a7e34062
z66346be727609d3ada4e8ed928885ed901efeecdfc10e02b0f65cd66068cda8db43ed93c73e3c7
ze1d5d5c59f5925a1745bb76030fd50007a6e71d697e2ffff0e311be3e1e456ff67263dc61146cb
z0aec922a7691ba63f32891acc9fa58410df1bdcd4121ee8c749f210ee9b683637108925e3a67d3
z5205351cad066e68600621e8d7dbd2ca32efef521d9554363f07ebe8c140d398635b21c77349c0
zc892138545c3542f1df69e12435e636d69451a30c2210e691128bd39106cdef828a90bf80cf31e
z7b651d413959f7beffdbc730341e6787d83c3fc0c3c2696c269ecaa1bdcb04185833c9a2c34e4c
zdafa24e98725a113421121634f2dec5340dbd27d04c38ff4b345d5465c218587df714723eb9bfb
z7820e841348285e71b801f3f42f735d4e7787d78ea021eb79685787931345493a5958c31ce550b
z719b5d697c22dbcddf37390bb464efe36b3ac46c108db1dab219ed7fc7a0b43032fe94fdb33071
zad6d8ee6695d6bfc9fb501fda0480795330aeb754e4558860252f367658e5a6fe7c3d0f9c99001
z5687c6e0c0498bd3d63539069ef4b19b49bfea849b59dc8d0fb26b1943abe3147aa87243e06c75
z2373e0fa977ca7382cb17739892a217ab9f7657b0a42fb7b9e7fe63e2dfe586175de013547b10d
z8941673f1d049438760f349d323e68f6626dfb7322ccec10a05b6b635baef8a324434e590b576c
za5026bee16a7297699455b99d0eac39d13f28a83313846ed1deb781cd49151e41b5029ab5ff15a
z545bbffdef62f6073363c288a4097a7e376f7e1911f52d16625c059df24be7570efc4b29c43cb2
zc8df30eb42d43b7b484f97fdb768491eda67c0b8c948da1eb335c35396a21ebcfd9055197a2c02
z67c07743a8ef9d20ec9f548f44471ba40cd8abebd596703d5443ecda692ccad601e7749950ee1c
zf2bb9f81358faa9d370caa4fc4ee1a09f3f0355685597a35cf77a9c02885f5ce4507f0d14d1536
zd4f0daa4c847e9ca625f984e99655a5a3f19b5393aa2cc5818778d15dbe9e5aef68d6ded9784b7
zde2c38591a0803ddf2dca4c9f26a218fad859873b2e32e1f3c94804932a5a9f67aad19ab8ec283
za58dfe73dabd9565c28f26aba26e71fa4c166640f9535af0edc7d3145f3cf28d013fcfe5d051a3
z373f97884eb2df2eb6c9094ab6c7427431c73cd1abbc9ae0f7af21fe9e61e89a58a5ca7d3e3d26
zae44898c9e6a9484e9bde6fede870de6328cb3acee24320aeb3b74eb5d8c2825603a51c9608fa0
zcca65eeb112d5d34573c69f5a898c2b5ad53e25029d5be9f379a8bb24be80a744ed4be8e3c635e
zbc5f990512a6a8a2ef00e74b7f4168c7fe58439b2c8a666245f358934950c2807ecef0d4c2bdca
z6a0e4e59d4e76d4a60e3a62abb8b979564b4621fad355dd0ccfe47e7eac40c32bfcca505290ff0
zd7bbece022ded3ccfbeae7d6a4f9acad4e682baae7ae253c04d4a754672fa3f09a3f9672fb0055
z60fb422ccd022462fbecbad4d790d2587a211731cc92bc7354f10c880f6ed66f92e4f5d54389e9
z25bd50df2b88181abc2785b85973cf334e15933c42382530d8ce7fc4ec3e7a0219e9712d574767
z575b7dc1bbfd1a11a92ed2c550d89bf50cfffec32a4466e77b729f73e94c9aea9647c873bd2a37
z062736d1e455af3230220310536fd2b78d59479f51e594a8f32c04ff12326f87d2416faf1b7249
ze351d9f22dd88730ca9094bd32ac9606b265a48bb0e2542e2b23ee884d7215163073728373f1a4
z59ddae020ce3ded2db4f5ff9b0fff258d68da4cb5d089bfc9f9d1f9cc8da0f332cc805aeb0bc38
zb511f8b64defd4a8cd06945ed5b566145cb9fdc8bbe7fffca1ee2d3f85158dcbd87a7518367fcc
z808542d848936e7b92559bcf3d6e1a92a8fb0ceee135b0a91bce829d7464dc00bc0722c9c4308e
z5b0bcdebc717365e7f5b578eb5c8ebab6ae9c763a92f32648a178674ab84bdec73b480bb9fe7df
z14f73bb82a78ab1cdbd1fe7a4db95636c53bf3ca715fbd8b345ab616cc2cd211f5c7ac4985f673
z8f0fccfdb76c1b5e754181eae1bdd36f4ac9b5fdace8ec893f501b67672cbad6b764b18596083a
z262b8560ae4b34fee3469c98efa6c8019fa87ef891e71e6cc444757a729757c3806c0b2fa7d310
ze57f117ce1015f4abaa71c3ba1ce0edb208be489ea0e060c5e0f7740dd7c8b04fc6e64d550c1f6
z77a79cc375627f1ada14f7713f649767e3fc33e757c9abbac535e308a2a0d5c4f793d4fb463014
z045381edfafa0ddfec16617ee498e61b7e5bf112e8fc90482e2f6ed2f85f26e4ca548888b14117
z82cb68f279b8389a88c291f4a9f2905666050f012774fb0738c5aa3f4f39a7795880661e5ada33
z6958764f581eab705a72bfe658ce39bdc26c031eaf4f1f61fec2c6534a6fce8159b6aa17a33c04
z61e1657ce6e73bd8f25a72e84df145b433115c728e0892a4a3efb905b993e3f460f78aca411283
zaec093d7468150bcf34a680e670c80a1c843b6c51e26a8c58dfe663bfdb4d0b2385032f878bcc1
zabb6d7cbc718bdd45b51e770e054043b7570f66a96134e2a950d00cce90cdc7c91ce2ef948d483
z22856cb64c29e2779527e4198e05e6022a307081877bec04909b066bb596ca4a9a364ddf81b4a4
z94d5d748175525908ce847cc692414db773e707d14856af92ccbb62abf4a65ea51f19c9892b486
zf1091b811f45063523bddb0e962f2297b7f5c24e6ee394d2ff77c24d2430f603e5e3373f84eb9f
z75821142019d4bf37ce640073a6f0da4daf114a057088c293e4d849d516c73d90fadb3d8cf97e2
z0df292a0ab37797269643c7cb7e0165ba6f3ecd4a500067691ecdea1889c4a727fc318f4fa8df7
za819ba8993786f0bfad575c79f31bcf8eb976e6a2917131fa0c3b359a53873982d7f9edf395e9c
zcd8cdb6629b81b122c54e420b5d78f2a6506978f67c1b0742035b6e4cce0f9262a92d97eca262d
zace0d76c9ca3e255e4c92d92ca4ec768681a5886dbcba3dce102fea6ff9cdd4a8f43866d86d5ab
za71bb8f50cbad99af36870518cf19366679fa3b90d990cf98fd68ded287c80e8c288b3f1d6f9d4
z22cbe3932c435b9e96ce22e9ca45e29e64c689ab28f603aeb5615a384d0aac563059b1e6972b30
z71be2c14fc3942dae31aa96edf202ce0970b311d52ea88a47b8e682bdaeeead5bb488eb99a1dfe
z64f5cb87366b90e5dfed0388974e30dcc53d17956332b858446bca2236f1e6059a506c4eac27ee
z93032d4b1b8195f305a362636ef6488fafaf19ae532dfd446e0f344ec16219820a5fd7b72a3b92
zb19416ae1ae19579dac49f6d774fd2b4292fff0d6658c2991572be88f2760ba2ccc70a185ee021
zb30bd7c3c1e562003adc239ee8a609aca8e7d69087f7977b9b27063777823fdd80ecac4d8f7b5d
zc59e1a60e6bef710e02108e481c6fa1beb24c210db699749e320e130e023482ccdfe5ea0a0d7c0
zcf05396926b9a1494882d09432836ac70352d8561815a5eb8363d4ec11222fa12406f2ab58ab64
zcb2636b025e33078d3adcff8258fae79d06c72abf91e1ab95418656e2fa9ef0ce7e62ec536758a
z14f521cc244a3c3c2bb95b03819e028a9931738bcf06e74ee1632f4efa6c0138dd9c9e35fe8e7a
z621c1336b1530be18abd10fed3f4d40dbd8dfa3e0709bbfa14878ab0eafebf5dd8ff172fd1aa5b
z79dcba08814cb8261f951480b70d2b7776bbad793d4c7cfed60ed1d23f172ff6b26a3594b46d4b
zca82c9ce9205e92649dd5158acc2c3703d7446dde4847520c99c26e1fe733caf1b3a1dd731516a
zca2b7e2380982f19b489ae2e8c9ee8067229d3fa06feebd5b99378762a4a5cbed1e65b26494091
z61859bd4713db775e79b51ab450db46f937cb92511006e11927ebe596a33255f6f685fecf03499
zc985aca19674bb7442483c3aa76442a83c51c1b007b7f13a9fb1ef2dbe1dd66dc362d38a54dad1
z6aab7df9b5c355855c0cde99aeef782e823bd2f367337e11e15bfad86d75eac28240b380cf4962
z9ffaf294ef8e7cdc4f0446f4846b80dc6a239095c19591295ed29e6b399e7f291a9abddb64ad0c
za5398b609b07fdae9b76eef99904b83d7f92e7353a80aa813ef2c48b5468776ecf22f4179d2c1a
z926e5f70904e0dbc5f12372fec667b5bf10c31df948bd45bd1c30678c29507c7f737beae971ef4
zc9d65e46d571b04de0be1b9f9f3710cf922ad852b2aa821c3a0a28d6a19207500d1e6d1ac07378
z2fe4f001f3c1036e638378ced1febf751769cd326685569fec7ca99116c5037dd55986ec25fad5
za8a225fb5c3851327e0bae08af6f1db2a1f07e4a369236108b8a76007b249784cfda789aa4af3d
z854485aa3fdc9aff58019e7d54daa2411b9a7c5c535d887a351515f4f6eae00121212056171297
z55eaba10b1d8d8fb5478a97850f17f80271ac5e93a4890dc75ccc91d3a1899d0a821e9f104d51d
zf6cf3bc1465e4ccd0c2a7b3874f16c10b277589935cca12840d1e4ae42dba82fe5900eb450fef0
z92a13006f955840177b2c029bc898375383a472af80824f24e8e1e31c49653d4bd112fe6d945bd
z7d4a5dcb51d2cd295e803204f824a20aa07b6ac0e91ccd2b461baa7dd5b40a82521f37d98c3391
z4c0440f588132efaee761c555ad5b57ee9206ea51fc6fa69794cfd5cee076f3161f11254ee532b
z907d1504dbb8aa13ea2c411228f7db98d02c09c18fea9312848c6862e4e37376cb37e4d0bd806d
z830907b68da74a06417ae30b713313de60b7f7d2cf0ddbdc63256646a2729cf3369dd9036a9b35
za9b5944b735bab68995dab0718b8044db6c3cdf23b9a9c891c26ee3d5f2c7463ebdc497826c53d
z43390a7a9ad59bd2e9dd8e453d8677e918a907e30b47322b539fa6dce9ff8412f8d39f2847ced4
z32486635052fcfa9706383848d79ba6a03b532d6ad2559eed1fda9f1cd0f7ad992453d72af8ef8
zaeade42cf21bdb9e831928366c049f5cfaf6ac9be89d661231bff41680e2f0f8dfeae1eb733785
z2d4581f33ff48b0bbb8c3ff221f2ec17681962d923646b1ac63ca709e2c00c55ca5fbe8ad7b3e4
zdcbf848288f0eaa8763cd41f6bdecea46a4c8681a4dd5bf951700af9d0f6e3ea88ee1d6bb58aff
z612a3df9c554b1945c752598b10978af5128106dabb9923f35a2f1ec02e29c7edf76666cca2158
zd52ff7deba06092093d8488cb4e422564c00dd52e051a7c4e2e70373a632141e6ed9a54e37dc83
zc1d9cc14f3c586df54ec223eb9e956d933460f182213c339a17f9435aac6a2553a7b52ef98d18f
z3666e415a0d36b75d56965072b8a81e3ffe8629e3e3b6e7c232fc72d0a87c9add16ff1dd7c364f
ze72c2a55116d663520237fbaa4f18ed8c50bfa27422f32f01431ec069e4eb6fbf4f34e42f6b9c7
z6bcd33d0f2adadfb0143e15394bae1ba761836d427a2100507dcf3fc48677dc23f21eb9c362c20
z46cd7c4926fccec66b6b3e95add37f9ea43d3aa1c20aa3cd08cfbcd702e334ac45b0d9dc9f6b71
zf660beb64da331e556cfbdf57164412745d16fa0189e280ae546e1c409942222f872a583e5fb63
z17580c8e7242bc7e9333f9fa5102f784c9524cd91ac4226639389c21efbca4d8f69785195e3059
zd5d026db5260a0101a39f29a0eaea9278a54e301089cdb3f101761a0e9d08a9930434b6f6f5b94
zad5a36f849cdcb3c5e8a6576c8be6c0d0af294de5b7d32148aadcb2237843434c9579bbe0e1a16
za9f2578c08f6dfbb47742f297e8e1c00500b42d382ac08947345dd995130f7978bc0c22c7332f1
ze497a6049ca4170bacd9a2e022533ca94600618f2911147e49141083204eea2358dd801c691e15
z47c8b541f9f2fad15351a36dff3febb39272a81c9eb8c9bb1a27eb26b2ec62f913b92c7d8f2d95
z218a45425c966a4440a4f0208f6afa49e091ea327aad9aa750bc3c512cf6b87eb31ea4deae12c1
z4c0ac37d3791d44a42a079f44fd8c01c236e12fa35a59fbf33a1f4acdb46068665d69d50fec189
zb6b14dd33ecde7c653e56fd8e7b0bbe8776bd36dd564c4091a04191adce0167c83e17ad93909df
z2998cb292fe03e2eb64dc880af0bb3743e7e461a29268b7f9bbb671a2dfb4f7e7150013ddd80e3
z66084a7d8cd4c98222187a64a1a0ad2fd99816d3e7b8260a6ddb21e233582e2dc226a203d1f584
z6133ed202c1c52a84b32f1726038ce7b2b4dde276ee4189180396e34ff87d7bbeaf1cc7e1472be
zceeacad8c186ec09feeedf80fa99faa3e9ce15f39379794d575daaf646118562d3734c99dcf445
zddbdd6070fdb8e7977631b8119bd80466d007acac5b46084026ef9d31f429a762856d99480f907
z04f025670df4627abdfd57f27d8684db45f9f28d781fdb1835df8674796ce663a2d942a61aa6ef
z65a95a0a1af8a7f1dc69c2e23914d398e0a2693c527cc5122a69f91ac5372b1e3657a4164fa68a
zff4134abe357cb579c8db2c250f3dad9ec05a886db899ed6e1ceab87fb860cd30dffd816cd8301
zde103c103b3315b8f8ebe9876b1fd3133f459a3235ceb3d8827c0e1d4110f4c4de8a3c8340223d
zc128674b4e037f15edd65ac52cca31d588197d4022c6ed2b3248e5cfca90f34e2ffa2b89250d11
za3ed6c095b6fa5fb1d0c8097780a8f9b596b777d0adb4a1b3bb9ea5e8bb2a54297b3bdd9e16df4
zf8a5daea9ed9151d9dbda4418de99a4fc22bc652ec525c16f2e52b7743901424e1f207463f9679
zbddcc847db2ecfa275c7492aa24dd4ebee44943e096064f35ed9929cab7c1496b6015b711b44f4
za6113de75822cb79ed7d3ac2c8eb488bd2dde6d2776d9e906005de547b9c587d168f590afec6e5
zde94acc97e8011bb2ff9004fe30d290fabcad5aa9401491ae3a8783d02d8e9ada87c3a6a346edd
zbb304a50e9964ba819a10aae9040ec18a2845fad335471dd40c14c1fa4d2b3f70d39e27da1810d
z8a3cbcc332982cefc9209ace85aa2d8f8bccc46cf3c870ac9db96781af993e25240d16cc9238e0
zb21ba7b8cf26c7c90ac0509a2d1950446df079c44ed4256319ec17900ee3a6e4dd58a6849a51e4
z2a227d21d5fb24f19e7c44e1eecc41498a2e97371cde21b8b8d4d9e1795f1ce1c4de2d5d52d106
za817999105cbb1128368adca44c0a6141b062dda89fe5777761dc1c1960da871ab31d7a0251c25
z60bbc4978c730d71a2f742f380b4b73b05773710dd3644819237a3d3ac88e0bdb17de0cf0572ff
z9e973dd781efb6478fc6a910fdfbfccd09dc68421b1d816780e5d9489a4ee2bbf760478c9b7e7b
zd8d124a06f3577baddef44fd2924ec36d2591da81133dea374e085a05aac199dc02aeb3e79bb25
zda4ca3d14cf4ebd1e6e94705124033534d5119b2ab775c63882aab4ad1f86b4f56affa0faecfe8
z23afdae8230b9ddd00e914712481de50fd500ad89ce306945b70f63ad454666392ff616eac679e
zac7f6ca91525cfddfa57caf56f9835e093b3f51ffed2d0d40e0dc1acf7b64fcaaa6c1aa8b0a713
zd44447d44982a3036478e172fb90865e50c86c5b471fa12d6a861ba1cc8e0594b13b3714a4aed5
z86f3a5b05daef8b056de8a753eb924af67d1353e72098b87e85c9b7ea810f750c394e211116768
z8eab1b26b842dbe7f8d4ad429c25729fd470a71bf8f2f84bff9343ee197540476dbb438df3d141
zb1649fc1bdc2b11f02ce4c6e1ec531f032d7840e88b75d2e35124176dc5cd5e0ea8e6d0c902159
zf18951d75145cef3014626bbd35f676755f383f472d6662b849290ca52bd3be48f7ab0ff1d22d5
z7408acbd10fe316806fc46e2779fd1ef79ef47110304ab5e7aa66fd314bce02b467b33e87ab1fc
zadd81e451f508e0a4ad80f2b9517f912f282e79879017708dd757936dfdb8476efa6d3e2ef97e7
z2f5307be159b934788114ffcdc7d3e3bec83b9d8861d76af0dd2326f962c8dd380d44a6513f779
zd439cd74f2d2d9296455a648a38d6651ac6847dde3fe841e79451c68a31098934ea65903e67fff
zbba3c9d40d89fa57c56a90fda3f16ba1cb9ab45146d2713fbb056e2c7f6a242a47bfcfef7c823d
zc5792ac0589dc5a22ac8856e75f3bcb1ec2b21579e91ce621562c68c7a0b2a0b97183d379e8714
z683e1a988ca2774dba599362e54e4eb2aae9d37f9aeffa5fa78cc4df3b1ca2261bff63a031cdf6
z1fd8f23ef56e8acd3b69e7e603f96ae281aa73137412046ac6b31f81a0b8fbb897b754ea35fd69
z48a4c6102d8b528ac46212363cf5138cd787df06b5dde7d9b17b3190a264573a517be2e6d7ad81
z669c8e750368af00a19848df47da189b93b940bff35cbace318afdcf13afda88a9a4fedaad59d3
z5383b07c79bea68fc1fa5e70fc4b2825858381cac42981ebb58e436712f22f03bedfdf7a22260a
zf8d4dd802b10e589e7e3b79fb63593e6f052d221aff4cb2cb466c8c107ddcdf8fd3733893362e3
zc8a249ae37841e193e81d371c0840d52194437d2c417da08bcd6ef2ad99ebd63525e2f2e616374
z4860da50af86e11e638b3c294f79edf7015ad406a40ee3595c655f6faffe14b34050427bfd8aee
ze7c4238a69dbffcb8bc41767f8e92fdf73e72b1ed3a205b3350204e40791e1053908328c585121
z9c6950490f1f21a45995917f9cb823b2f58aac67842e4222008cc337dad87668dd65b6ef051f15
zb95a9ad3b48ba89f8f863cb5b4f69b4b68426bd06ec5dc67b0336a93e2e56b7aa88f9132d47b05
z4b7fd57a1ea8ec083d0599996dccba2e99f91b958aceb74b4ebb158848cb4cf31496047299531b
zc828674578347f44ee6bbe71e61cdee82c0d89b00e63cef70cb15f3cc030e54ec1e51165c7f145
z7f5eed8bd8651d6c0ddcdc44b48b45b76d430e8a53dcdbc828a95a701fb524eb1b3d3908075e4c
z0a8f55a038f7b3890fc3c85b1aac3c352028897870614a0b7a407f7aecf210aac4a0edceb9127c
z0f278194a420b2722373ab3af34999c113615648428a509dce1f51ddc4aa6f8d786255edb28d3e
zd10090543f9ce2f85cc6081028b337dbfbc1cf55b9016c46fdadde391d53f23386375bdf63cc57
z398bcdb506065fda841edc1055014bf13c03cd980314202e6aee994648266654b522df9b3beeda
zccec4dc6cd886109de22f2d264722b22524103f66c15950e099d00c457bb8f5657ff265b435a7e
zc51222e0fd540e368215f68ae5ef2cc9a160c80ce5398b01eb5b85f41b0507f5f732cbfd47552f
zcb6f592491cb15e232ec8ba8379749738f5a5450794ef0f501c3e2d245478312b36f5871c4dab9
zacab971d0f008cee3e2076a84f514862f18f362dcd7ea3d07d4175382823b9f9a0ab9b9d264b6e
z6761f089d8dc5fc687d748c78f59420002900554d306f661a090dfed12021bb24772d3e83f1e58
zcab0cb2b171732da16465288a6347a577cdc14f56aa8d61242e726e93a4690f653c44bdd6d76f9
z72bfb3977c766be7f2f9c5eb7d6123beb599c7c7a87dc96f7516bc09fc58c900d2e54430286340
z43f61506ce32c8f6051850fa649bb345312b7a836c2d435f5747f83dde88a50dbbe4f732228e2c
zb3be946041deb134c9cec1f2ebac66ca50a41a978c699d4776c50d297ce9573e5d84f292a43e74
zcbe99fb70ce65b68f6c97d4a9ad54c3349f9bd107b0b24b93bd62a583bf2244b2ac1d82cd3d980
z5dbc39022e04fef100ff63204ad24050c992fa43f14e823e2779e6b128545fc000bd20e824f8da
zd084db1a7911d9cd3009d4d81019a3a072a06e29ebe395827a8bfd3d25eccfcb768d3cd12802c4
z9161062a37800de3f3936d38087ad8cf3b1d18061f1cf288fed226143b071e145d28647358a7ce
z7baeb151a7131859a760494c663053abab51a98814f0db159c9b1d28d0a73944e443dfac56ff14
z7e2bfe1829869bc57cecc3561831821458878b04c5ce6bf7c68a19e0cbd913388913b6ef6f2858
z70d052ba7842bcaca53b9adf74b3dcb204c8c29f4f1e2f95a94fa1e3e7f4311392a8956f999266
z45a5ac0a79693c934ab5673ad6b94f2e66f16aa9083a9042e801fe6fc6c6194f81a82fdd29f460
za1c425a9b8cf65b77790e37132b48e2282bddb015f6c1664a9cd201c439810df915698b5a8d827
z7eea6632eb8c5c904386a76c33fdb9502fe11ccf5bb00cef067c43384bebd03f096665efac598b
zdf5df1d47e625455a9535eb7d31a6e4cd026f18324ca24708e6f9e079fc89c1a5c552140387d91
z86c9fc982c176cb36ee434fc7ad54002554dd224cf9398f4d02d781b8a6ff63511408038cf4b23
z65cd494473117aebc19188e85f1d282858eab6ef997c83cb226474d8810443583f22e511e65f1b
z9cf853d7feec9d85508c3971cefc65a4bf96a400ba6f2c40bb15d94b791060bf3e0efa706a1f1d
z6be2beb3bf511a9d4df04074196de9f82aa5f1f16b48d249468fdf78b27c4b2228a538f8a728e0
z34596d44619322b66dfd33f8651d97995bf614332e61b988d9848f919b36e5578cce5c207b03fa
z9b0a2e256d706e1a36e0f0ecee9aa5f569fcf920a10bfdb5ab96a66e2c7443c68d9ad6341d6669
z7a89ef810e0d4b0bdf9faf1b6cfa2ab509e0949df05786f76f15ecd86c2abc158e65c24f9787ab
ze5a7cd4e9a70459debbf8451426d2e91fb446055da6496b61cd1a01373d8d6deea3d5d812d0553
z575cc539f10285383f9a70a871d6f3b449f37337b0363627aac76ed96ba5370f3a5dac633e633b
z7379d120ad07f72b8c2d2e567835086a9e144d5ee155f01f1e7a872743bf96d0f4c88631b77e5c
z3514ae17659aa539791f62a2468e88c9b0f0701f8fa31e7b9c3defa346adc375da8e2c099923cd
z32124028e6e17c8808f6a3a5a6645f1ff58bf9db24c6f9e2732ef61a80b366e2a1d229dae11a06
zdfb41bee2e3b30bb2a615f79dd618436af0171b0f33aa703c45dd6c8cdd56f836a60ccfc0b566c
z40cef40d747ce59a55e54fbcb76bfb71f47c525db720304dc47bca812e35aacaa2d6200e928e57
z3772e8e9b77fee68479af71546d5b93fc0b79e947343fce7a6cd9e3106639c67aff2ae028e6c05
z92c464c3aca27d9cf3f569739b3863fa00531bb2e26a0767088cb03b6c744c526ecf20920586af
zaab65e6424fb41a1c5a249198b471fb96a368b514ff8617942c1a9616adbd3b42fa658de95b3f8
z7a5d9b5b8dadf2fd12f4210605d20dde6ae398bfffff2e5181fde5cfd9358df7c8d8fcad7eea9b
zcb916cf3eadf69e2f6587ea985672e2bc3ae25f1bee882e26a9aec7da59a361aa56bed21657ce6
zec31ab4ed204d1c7a8f6ad30e48cc30315a36e34c7371578f1ae848a0f5b8e80a8f9120770b105
z0531441a2fc940026a81c4261c88a94aaf15c0aaf3faba94f890a19bad117725f659d92c8894ed
zace161c510e5d840ed9a3fea8f413343904f1093b9e8b7f5634624c1b04382c30faa8f2dcaace8
z238765b4280290950299035a6aa86fe2dc5c5f23b26fb68ef84485feba1d157809cc41399c2d28
z6ec6abe33b16f643dee956a2fada64e915ea230171ddfe14dc15a28b0379089f4e740e868ef316
z0b357399dfc32b13c95ce0d7c89e324b581975610e820071e643d9a394e4b512c0fb22a956c8c7
z829d6a117012bee3c2180b267e6be863ecf9899d6a839685dbf4c4afbd256576593144542b366b
zfd67316b6c742f7d85b6d8bd1fb02496481bcc2ab57898c112d499342173ddd1a0813da6c5fb8c
z1371960f5aad40679654526e4f1327e5eb744c0df1046ed9518a24b77ec1aaba22902b7c28751c
zf019fb2d7d4e2df89e1a01925a9f50df5c63f9488aa186f3f23fefa4601bb8bc65cd64746eede6
z32172b51e7099b410fd684701ecae5ca2d650d0bc835704ffa234ea82b0337f07752b9fae07e14
za85bca0f232067159ec7f4f2ebcd3563cc38fb74fef4e0f96956a431bfd8ea7d9328cb4e4be5ff
ze8d408eb8aa8f3fd2874f518d25bdde2ee6a72a45b40835b5d1cf5768d2bdfdbe9df01cf4cccf9
zfa7a739a7dde70ca17a7e67f850679d0f09c01527c4b8974d3842eaef029e7b1ae39e612a17b1f
z333b4fc58cd8326c6852387652238aaa725b0fadcc8d29e874b552000fc288a7eec6179d01bf7d
z651223945c20f4ebd6973f51efb8e49d4181531bf2dadabbc3ed2e5b77a9f1dfdafc71eacf8985
zcda872cb622d6fb8ab6ed58ab38b0f766ac0c79c774548187fade25e4fa452d4409738c263313c
zf2e7fd79e8b1b7dacfd4aed56bab03791f00a5f1a914f2c998744c4a81f1144a2b50f1e3205b10
z60acbb72f01ae74f0c5eff25f655699bfd67d10e48630fd17e2a682e4953d43ae71e542bb1e552
z6c66e5f2ec30882d961cfb636380000789ed2e3dc6fec5af0ef339df840959c6f6e75cf1a8d66d
zda7a306946909c05ee6db841279f21bd8f4d44331cc3c64982138b99827e3cd04bc4ddf3bd7ad9
zad7a578a4a2728fff5b97cdb70307562b559ecb7f869afb4005f12fe5d55148b475e9bafc17313
ze100858b69e39852c8a25ef9ad765168ec73d5a10f0c6964c51bfa270a8dc673a4f62494f925ca
z176c602fb0f69ecbdb9c10df5bc188edbb1abea1402b7626c1907ccffea6837d7502bed89ea060
zd07851bec3e6ffae62e56f591d059c6e87e3baec2041949e5caec606e6945912d90e5870a3a754
z4d67bd910393a1bbce43d39505e7c23ba8b3296c0826d833214cf691aeee686dc48bf224bff415
zbf7d1f4785ff1a6d6482e21bd90c7e240b5a1f5706b31b82bf821598347a755ec769b925b9b038
zcc99a2b5c765485f60166c4490a8b21ad239a79be18e7408dc0110aa0a5145ed894eb4aad920b3
z21a1d7a5fb65561318760d0b5634dc9d2522e74267682a3437abcfcac211896f69f097bdbc2dba
z32d84b2606cd24e51119156aa853a17a86a0f0c77bd4c3961048b27f2c9524ea6d3bdcd6b02f13
z1afe7375886b57d63afb0bfeff8263c4f7d31b75de3ac6dc034c31c58203ffba81c26201d3c63e
z31d201dd0abdac0360605734d341178ddf438cd7323fa2faf5a78efb22db2cb05de5b68d270198
zea8e44b576885e434b9b280fdd2de83f53f0e35d4dace9322dcd5a1de042dcb8023e2dd2603ef6
z2bdbdeda902f7d2d0e138a9b3009887361f523c59953d5b25df79acfb11391241248aed62b31c5
za40a5f1680e36966fea0c2cdb4dcf8843e37670c9e1ff9ed42266f7899382209d1f68258f5f7b3
zffdb3e3741a67ba2c45580c6e6bd274c4fb61e0ee77884d61ca1aa54f5c4e91fbda505215811bc
zb49700259ccb15904683967954a25f9bb0d135b3f941bdeca5b28a71ae7f6700b30513446c6c06
z01e16e250a8d4fdb050cdaeff7cc200891cf14532e185504144da1e83d903bd9fefdfd71f098c2
zae0c666e3ad82316fe80e8064619a454356e363ad1655d488df6f8fbd02ae846400a1ab0dbcbde
z7f5c1105db22b6ce7ca1ac217f58299466b6c0f43458b3df3e1dcd269ad4ef58b2e05fe09b3c33
z10cdde3f5ad290cfdaf3920673a41875b744cf50ce27b4d3c28ae79d2f2bac0c50a71c12545982
z4861f4515c1d69062c9906eb7604f04b9e580d7f8032c79024fcf2717b4e32d91a4919f96212bf
z6643d9c00f0c0b94f31128ec3e17d6b3ba2a22328e67403858b453e784f80ef845356e5d8ea0bf
z36e915f7cd375dc0ebee8a0c959a57274256b6f45f62af07ed854848e14676dba6e3007bb08ada
zafcf5890c16d26a838825f4cee8ef78bc372473a9a9b01ebaa1fe4e889b48df5ff73fe6de5ed2a
z1479f26617c092683469b94885e577604dfc488a605c39f6b4d58f6d101ca38a657b82d55a2ced
z78207e00de4b106fe501c67d56390e42674cbf8d41114533cac23f3775742bd98a43d0076e92f7
ze7504525b4ab866724be95d5d8e5f78b32e16b95b7a51c1a198a9a67fc03deea8934cf085304cd
zaad4eca0822148e3c518562a96001a28d817e5e0b04cbd64e7ebf3a2d35c898147366afeb7cc55
z60cac79a8d6e2915cd94cf1b65d5dbf4947e08139063f828fcfbe70fd8de506aba15eefaaeb5a8
z051806209e795f49d8087621785c73a59b7af5f4582cf9e1198dc1b3a151943746c44c273b1348
zf378e4cfa31f2765786d4be5297efe317406b7e1df6c064f52d8d72f1f9b891976a0b4a2496a32
z4b12b67e0c488f5fd6736cca13f55e05220ad2de58b814f397b1dd536db08bb4af3f17c8cd0933
z13a570039c991bf6c69097fee4947a4f5992398996f47655a9223129750a7cb6d968245807a427
z9635f402522bfbebcfa6ee6438fe8188fda9c28e1614101e9d7b40261fcbceb2a15bd2726ff40c
z27d4783d7ffa667d30eee0e35864ad99e0df6b8121422aabe8928cf5c098dee0fc998d872bd7a0
z1a747bd54a08adb7089f9ab38fc9e17efe1b75c6916f75f0afe0a6ad8c165d5730f71fa10129a0
zf20419bacd49a0ce97522851b3720e220af3cb4fae6cf7edf27b143c4d016a843ea1ca011d3df7
z03ddcb5a62bf0a9558356c766aa2fe4988022ef378b7081b864316f63264a8c9c626b4677d2125
z3936412e838c9ae3a388de140859bc6ecb8c9e556a0c27132e93cebdd34d49d6774b12b7e495ed
zc93805758e2e4f4ecda898e6380701cd3a93af7cd3476b0167468bbb66ddfa62eebb99ad9219b9
z0934cf0a57a488ad1cb5aaa026dcf55fdf967ec841c3f17d6d489d241a1e22567c8c445aa2ff4c
z4b3751b244ac1b3e6c00c246c86d84d0073aa231b8c8f7895d94d55297d10ae3a795f0277a307a
zf45e3044d98159f98a48608d97ad71ac4585bcffa711aa20200d1d2f18bfa12abc120128c7e74a
z18dade0970033295be8320c127535543cd13607f389ac2c6ffcea67d1dcbee5d9cd062a5285147
z982357963bb14597af19b76165a884aa66750f47b373aa8062447a97756ce8534364f51a9e226f
z35ddead4a32408523c32d08d52581e60cef5e8de9ab5a2e060dd9a684309e70bbff58cc54d5084
zcb1bcc32ce7b8e167e7241f1c28a3700c7f668c7f2d52015cc5ae53b2a3d5a0dc35dc21bd10dc7
zcf04b7ac4c7b73ea2132b5f2fd446bcb16afc3c8bbd58d0b8a38deac63d879167114799d855ba9
z554368b7803d61d4f8e5e752544ec8b8e7b4767b7003feff916bfc098d1562cc75cd0ff97bb7d8
zdce9f4a97864e792daa679a2f2654a4264028c4670b99c2be62bb4818422be31119da03a8e97e1
zc7174d0c93724d9c2442499baa61c5f8a0cfdc35dc210bc06180a599f8f4c9e87631df67780d8c
zb8bf122d875b702422afc22bc522a79a8bac3ccdd737b24e3f5a38a0f8b2fbfd9a27708dbe5dd6
z9c65a9a37bbacfdf271eacb4fba03bd8eae89932a34a310b9698c9dde198617109f94389241407
ze82e8a6ac42e67e7b13f34151cf88781958ef7cd4565835e576e2c972a9db605ff8d6ee1708872
z5d17bbd0311fd27744e24ba22957e5b4097c4a0fbc44307d9fb70eda7f91edbec6e487c71408c7
z4efe5e39921d8fc04d871337c472ac22cfabc9b5087295f15c479acfcb6734b0100a4d433a63c6
zec09e5dd49e1ffcfdd7e360f28c044ded213bfda94796bed39d30bb20ee173aa70bfcda70738a8
zbaa776d1f24f0a7ad562e4fd76bda78526d7e773ac25862b2be3b27931621ccd28983cc5479b98
zc94705d64be09c2e883e7b70a0b0462fb0ca24a1bbf6e4f937d24608df350b49657fc314bbab26
za9764436744affca85c30d81217fdc5f28a172cdef4963b72dd9799699e54103ac926bfeb03ca2
zc05ca4100c5bc03e286774cde0d4b5296c32ff9f0520e2330b08399a9d89cce558e0765f7581a7
z7ed41d76e4c79eae1f097e49b26660d50e3192ee9881a18aaf37547c3f121c32febff81272920f
z96a754672761f2a82934aaf9427b9ff4ead273212ce17457ef546f04fcfd764e44edc1d57ccbe2
z800ffd63d00a7156291107d72ae8a0666e81936521ef1b8fc9a15287da845a2635909503586404
z6ba047edcef1299fca1aafb748b316b38c2f5cb792ac035238d101139809f474b14fa5cefe97a8
z23d31463d221f65483572f9b0e13137927fed6df9729a8c3f9a119d3f8e67382412977e57df553
z1569a7d6f3b9605ecf5e9801a7e6e20f7a2e68607a404cb585039ca66aa0031c200fa656d65ae6
zc61dcefe403f2c5f4b2300b0100482155330edf27d9c0572a2a38442adc1aeeca14224710d740a
za9a597fdb9ea1095abc687637432284f858c5ecde274198bbdee4ab61415367a828b2ecc4bdf51
zc0a7ada45eb3bdee78647de2ebf38b11428f1f2cda155ccee67287b1c161fcdbda83bfd6fbe18b
zcb029bf6c8c7978daabf34fca0f9f7637a72ae693d0fda80945242275157baf7b7f2d16a6b1da9
z489cccbf0829eb70014a8e7dd5c845b1f29c2ccaae352812f0f819f04bf758b4bb4b0339abc47a
zaa07f01cee0bdc9d7454e410d4d5e46ea7f3b7fa87998d13e994afe36f259755dc058a3bba0fd1
z6a6ac2afb6215bd7a8616f6026106cc89f9fe7d3f41403d85cf87055efc9e046592ee9c1257719
z2f7fbd4e7f4268bb94a5f952b5798715a0775e1109c59e19c0384884c2aec4959f2434aa36eb95
z5b483f19c910f5b1d2eeec3f0518eed77d90b30229428636dc338e597451ff402e8cbd49610422
zc59572c6371fae86c0c76b89f9339e96ece5b54ebce2a33cac01551b3a08f5c364606d55568c42
za511f13cd0bbb099ac61c39d4c6013d52b2843b5f3b2b5d277d9d8817767e1654144f9746fa7d3
z7cb004f88f89f1877083d2a21745df5679ada2a5d7893140a0591cf97ae71b851a9541d3497206
z01d3c8761b71eda3feb046edf3771f0c60e1acae0fbac9336d1d5d3e1a7be0d839171a6a10721c
z3f8f546b713f2d176b50c7a19afaa241efe856f643ec169bae99389d5530d08e326abfbf466ebd
z1985e0eb4b3a44e798ea4629728b2fd4edde768798bf27a324eb36e8baf60abccb0c8d78d60666
ze45a510640e0ee8ec239a3f2007bc2cbfbb32f56a7887504647808db0ddf810b9228752bde7536
z4b8300517966491d536a955e171fca4c44349aec9c4644f59a6e2c34dfad9480f4843d9e02db77
zc1353509786457e9275ca95642df92deed8337e75a74af17f85dc613236cc9caa80795373b64ec
z4a3ebe0658ddbfacd0b57c145268656a7175c55625d8258a6d870feba7b8d699d5b76d64e2513c
z6250092c9faf19fa1ab9849ba578018664adf2028ad7fa7d22d0bc7650e046529176d60d28ff58
zdcead20d8407d580d2af2233f7ed7f4538150c958f4303130f106dd073ab7fde0d7255e2188c80
z523d0905399bfa66d4bb65c2b6bc9b8c3ddc04a4466e5888fa16f8ea09da387e83ea72474fc071
zd2cc6ac8d3739d86686b1c96196a4883fdd3bd7bce1972ffea47c0f3a7523040ef621052c5acaa
zb3eb90dbb34b9b098ce8a5e5b674b0be3fd93e25e7c62d941513a08aa3f31f0fc131cf2ba0225c
zbd1f66b8d9b3a9fe3dcca1431d13f87869fd0cf77b68db9ef54a577d8df55aa4a2be0e42757e2a
za90c9eb1c392fcc0d9a559b2c09bbdb5467179e28e8268ce99077d503fd92a3ca61bcc5d4a3d68
z05fdf78b657ac3f280cbcf3477c6e0a09b5c05468c987b2aa1da38981b3ce605b6bbe9fb7943a5
z856e52163fbf8b987eccb025dd24216e3d551c715c2a93d1631cb5e7f37e2c356d6d92628b2fe2
z080e54e394e6676bbf145b3c03cfdc796aa26d9d55c240993eb9917c82ad58ecae10ec50c6eede
z66d22d36b3450e06d5517ca21c70b75e5cf1c50965878260b0a15dbe6965245722a95129b9333c
z1007dd38e8577fe35abf4fac83740453fce902c799042a4e6c9dd834b7ef482a3a7c18627c2d15
z8399b762a169b034930555f098374d54f79e0979217f12c0f54d9d21bf587fc57027eeb31cd8d3
z012e56e4d59f2ce5c1cf08b267ec7ab3c691dd0ad46bd266ef6faa159a3402fbcdb1c380bf5723
zd8f2a92657db8426d61610181d4b6ec104a2ea036d9851a10917da627f172781fa1ddff0b6df02
z6af7aa15b2d67b0d0a4f5a3e2fabec828175e0fd28a5b4080b18bf9e789dbf98d6878d82ed9576
z99932cade7f67d0f64853288122a9752cd9ea375545852a6051c3bb05be927f8e78197323a702e
zd69428e9dc11a666bb387b82784b3d8a992d9f30da68c7ed05b5e6a06fb8be5e7c1e5c6e4b067f
z4a1e3b53b2ef72477282b20ac87bea3981486ceeb1b74990843de3bc73cbb78fbc66098554fcf6
z817831bbb6a2737a46c6df6ab5142f4de76bfc30a7566f70519218511295ea1e7e3f0e9eb4503b
z90bf9c2641337a40cbaef3f636bf27f95314ab67bc6335366b3874045b741788c84117b98fc8cb
z62af2ea018946b3be30ad45aa9ef53390976acec037803429065d06bf46384e968004e2e9a99a5
zb1d7f2308f9699a66e1dfe319b2936aac3150833ba76549fbfe86c3e584dbab9c4bd058f77ae3b
zaeb8fb70cee5e51a494053785a7ce6f80dea27047fb06678fa8b6c8b141767cca99912add9f248
zc2ed0dd23fde6a70876491dea3ac18b7389fa936cc5432d74ae210e9a961431792bcb1464c4a5d
z0b296adf9d497459204f220c7af8f0214a7a7b74679dfbc2eb169a393a26ce8b7ef4fa33d67c7c
zce57fb8f0e54373fd08be52fff3a0dad61055d6141371dfb76a662b5a30d870e5713f4323b6612
z24aac092bea048e439a5c3b7de499ab32e2bff9d83be41a4f04235165c48e973f55c55d48562ed
z94ebbe045c3157981f7081b82908dc0eb381c670ea4a8f7afe75d16a98a54d06f8b370ca3b78ac
z27287d47de5e6546fffd30e9ca77a4697c2c08b9703d70aead27418770e4fd1308259489a8d51b
z3aaa623e9e48eb56cdb5ebc7af93017a18533bd74ac4a94fbccbd34eabb8fd65fc20e7b2eaa968
za076feca85b68f775d399da9451a411c7b1a51528976a0590c47c72e60e1adb4b6b294136cc82a
zf43db1722d4bfdcf5d9cf736057620c404424d931d83be424dddb022846752479d84a2ef7938c1
zcc345fad9e74f9e1a0c077bfb65d78e65a37a86064b0bb94d590f63468d2196b7d0782065ab968
zf4a4f4b19c0ebb8c37eb454ce630aa9e8cec1eb5d6e599e631067fdc761b9b18c57cf255106364
z876196e04445899dc139c1af6463f3efccaf4e820988a7bbff1d4aaf084efbf09ead589d62705f
z19909e7dd8a3be848e01e07e6614f8364a87716069a359d685012b679280879a6204ad424bfe90
z1b36ca30902cece5d76c9287a18643e1e740de48dc1cce415445b1ad38371a8ac1402573fb9e04
zbe13e566027298f38229097239fe7b73ed998b6f351a7674aafedc740b68d543bcdb3e34c89b26
zbecbc0eded0bd332cfdd71619d17d8fd635af9844af7a571f52f68aea83f40eca1a5cbce79ca25
z28ab5f860d4db832a922d699f57c83285eb539a639f27e225a282c3369ce44251a430d452fc829
ze095ad5a2fbf74eedf8e5377c5b6414f061eda4bb9c2b36fade5569ab0143edc99e601623f5441
zca9aee2597ebcfa630a485b31516baa886860a10bc8a3d9f5dda9e5fd70305a81d9274b0499ede
zc1db45e9246cae615e478c615ce66261767cae534fe36198c826e8871455ef9e729ee3d0e5f056
z669eb8a595b6f92e240a9875fe257c680c8ca00ba97219141a1612e4f5a33585d06dfac438d33b
z822e86d48f89e7308c6715a33f5316b0eb0cc2ca6d1986dbf759bc792caf841802c869958165f0
z8fe02105c7d15fc47d3922c13ca9ed273cbe1e7da24c75f0004a82d64dbfc8f920e1f35bde28a0
z5ebdc39727042427e24c4364f25c14887463aa2893a36b9817b6a7b922525276104037940a08e0
zaf89fa669cf72fcd28799fc40eb8afbda01b92c8f294d09e227a3b9416016b82a64fdf71217cb5
z4d1f370d380103f458b3470f32c3bf68fcad93fedf6095853f4328096e92acac8c6e5bea736001
zd32b7e49426506306d5e78f7051377555fd8a5c3690d8500b8992f8398071d5db9064fd4674832
z651ff1cbb1377d4bca3e7ebfd131ea1821f82bf981a80515e9b1364b608e749461fe67e68aa68b
zf6ccc1628ad7c3399294ac64bc0ee7f421d82299ecc79e1893f6a795b472667b245dcf39302639
zb2b2205c447c8f9dbd92d0773986dfc22df3d0445e4d693e2a57e69565ad1ba3eeb41645c5f509
z426a1da6bf85f47495c293bbe7021c3abd2764ba315ca589f03cd80210b1cd80f8bbc3b8d537ef
zc51d189317cf3d34b3511bc96a791a675dc23e69370f67878074e1f1bf1192734eff88a5d36a5e
z28c6cd8396a9f6dbaefad3a0e14d56974be36ef9d4bf5b1c9011b75e2e48d68bad9e5742efef17
z45ce77d28a6147c15839c860dbb2792ba68944cbfa7e8989856264eeccf799e4a2c67153b2faf4
z366463cb6c1e3ff93325b25d3358c1f7df03a27ffc52646a8e9ffaf87e624129786264a47d07e9
zb1bf668fdefe9f4dd282e5db61ccaa71d7e8a8d0f6a94c09f29ab351d9bfab3c18506b26af801f
zaefb9eb4057b379d82808750d828422268f9dec3e118cfeaf15dea9594bd31c43a57dee2ab3493
zeca255a9a2cde58e594e5fc1712abdc6a68e99d06acb80736a6ada4b688890d0e5d3c15f665bf3
z370f65f6a95f8a6ad636bbe99d5edad6e7d3dda9cc3017052ffddcf698204340aa2effcabe8ed8
zbe08897f4a9fb0041e8c37b0b403092a423f0e6519e43001c5225850e6ad31db6c8a70c49c579e
z13fba31549da565b4a15577787aacd5ee70f84234ce637898157512f44f610922e405d35a9c33f
z137103de67bd46f4024763f69ab5eabdce9b6606d4ce96478204045ac1b70cd90db4bae8a8c2dd
zfc6a95eedb4762c2604b9bf8634e03f006a2b618e1bcf7cc849128ba4ba27b7e0eb915bb9e8448
z1423095aa401529d842c7f55c62650665f3b4fde6c233c31f4ab892f48216e97a80da565d6e122
z5f465ee34adda5c17c312268d8e8a99b380f720dabd8e01fa44480fa999a924e9099356a893110
zb15502cd1675577ec631dd0cfe78a5e9b3053c022c51758339ae947ab5206ad4d70799f9255b55
zad650f5e78ba8d470a08642ea8aebab34b36783e7f6f157280b9816f8acd91efe668f743464a16
zcfb8e389e377dd6c3d7f6b227e3f9c7ecd70ead878b514785c07e84d8cf54517810b3ef06a6fca
zf8ea375139600ebb29940aef6451221eaf9791eb269ab67b25312e0963a33a8f21892bb18ede6d
zc014074fd0e3ac5aacb79c8e285446c214aa0a621547f440dbe05a1f20ed88e7e8c2273790e69b
ze7d5abb700383abab5a0acbd9427c8c56e8648ac47a273a1bf2984bd6595f9c108065c798eb180
z5af26fed29547147f5d1fe65c98641b89ccf40fc8535956690189fb48fb7d73ad0235c00c592ee
zbc1f4f905289b3625b5311e50452403b3b9f6fa8d23cc33dff842fe6cd8c86995e0d06bd895c5f
z9ee09ab638fcc93330b451604ed6cdfaa56a08262a34b004e0117304e0a462daccafee3626954b
ze9dada9944197c426bcf362ddcbefcd1bf932674988d98d548b126ef696036715fb9a495f3bcf1
z094dd99ef509f3e67edb15ac230349f0c6815c7dddca9494db21ee2a24f08e33e02cc66f5a8628
z6687343ce4169a09036a811d0195fa38e4f7ca2866f008316867fac6d5ec04426563a4eaa5bbc2
zb700f0d012cc3a2649f880b807d44053855cac4104add137527198c031892f9031b45dcd679b4f
z8b78f33cfa866f33567c0cfcd009ca1ea0af212821c8191b99545aaa6f19b7e3647ef463ad1790
z460efe6f5c346dee2e88c6e60256007b09b5c42fc1b8b2b6443f186ac0f47a834afafbf2304519
zdf7a943186369303920bed09c551364c7b66f3da631d0a5db0cffdfecdb9a7d6be2c486d4e0394
z74931a5dd825e3d7eb8405019b372a053f477673777ce9da2c2260a0af712720af1452c94418c7
z801dbe89165f94c872ecb1d74419b7e41f866923709f0a779543e2849c1e791958908a8b57a42f
z8ed2f82841baf35c18bee2b6880df4fcadd16fae98b3838883fab77d92a801d1e3dde9d3bba662
zec4b0c1370f9e0a3c6489f2da5eaec74f2fe36d4756c12fc3ed9c6a9a7c162ddae33eb3e015be1
zcd9bb4161926278893e11f039e97b59da3442d47c3264a1fee8e9c4649dc11205568f359dbd422
za339ce55053b058b25b8077e6fd451c6a9971f7f9f067dd59539795f7d0851a22c02913d98e842
z0cfa973d856b4d17b9720ad96f6d1e8c0c2f2c0c68cdc8f2a52a5f0fe6953c44920bff40b04c7a
zaeb5e727654fca77f387b1c680285725303c4536a279c2fc9afeeefd33a37e7e1aac0802a841c3
z41fe9474c201638716fdf11878c7cd06bc2f3abd189b14c96ae92a1e910e57974aceadd6e68ff0
z89d1987438260f5c85ddc3e51f3cac2ac5fa4c9808310c2e6bf21fb9d29fc9f6106a9418a55d15
zf558e32b7c462334a4f64dba7676aed7bd8f1b52f5b9cdcc2281ea9fb28a8cf80930e54746cd0d
zf1b6272eb9d8c9753291c5490baa8c09144fd4283f39978428b5b7f71b28414c96e7ce96324d56
z44786111e006c3ee518675bb808496b8d792f24f65091027f2aabd54765345e85ff042c7f0bcc6
z277a35cb059b4075eeec6b0baafc797a2ccaa169690ac064e4c8d7bc02e37ffbc03d4c0ad75b18
z5303ac4e660567b0b2dc986a70039dfb09667366b6fdf38dc784498870eaf4c8b81951525bee1e
z8c252ee5e9a656c0f31c470e09002b576081ef2eb6cf0f206c4a994bac533dfc0a2190143357a9
z589a9f36eae559273a52b62efe5269f8f2d94477c952e47888ab69f7439e23b0be57d55701f6eb
z6db0aa61331d4901b7cf85967f2ac5c3d79fefbac7e6d5f63e21b91e8fb1b439cb76d0d4556f1a
zc4231e75577177546c0f7953307774c4ca1991b008f7d878401b9f2e03f1a1bf55d14f187ef6c7
z64b8f947c9f0079641ad7f4f1a8cda229442304970210c95e91fcbf2b09fc553dfeb3692d2a552
z3718128bced6997895fd0e1e7db18c0379d45cb5ca6ae697e81b9d3dc49c9055cdcbe1128d89e1
z42d637638ae44877b0889093249d62a32a68be4d38b948d74c842415ea3b6f47fbc54652b805f9
zbdd2f4aca95434905bc433b08f4bc2e90042c2abcc3ba39270425c4486caf94a0cc5f6254253b9
z41dacdd8da9f54ff54c735f320b34bdfcf650a857a22720fe4483e3b6812331578595ce28eba73
z0dc9bd9c35ea95e925f7448f1ea1eb3a8eb8f27d7b7ba03e076580837229a2e377c7b91869c80b
z75aeaec1b8a67bb69799d545a4855bf2703ff47c47269407e57e811499038e8c91399123066533
z75e536d65e203444fb2b2131c0f40c4b21625f7a5681a612860bfbb8d19496215b437a11e79aa8
z2edc0e4f77561a9c6c7a75381e8684b24d6bcca92efa73cef17e771b05c4c8565324caff875d54
z09c0c458e6d8df06c0e29c07e52905140a9f0416b3c9e9a84992e9bc7fa8de0006176f4ad4003b
zaab77936c1146412cc6671f244b23324f4c797adf64d03816340274b0c2d233fe068f61dbc9f17
z7f282bf7d234898016ffecff0ab865ac98ab73d7518b8d8031a45ef8985c88e6112cea569c3ef9
zc23ce95c4a2b0ebfa4f79c4675be78a20dfe136a638c3a4b4e311f0e066705403a855259c1deb8
z842ec04bd900fee83b23314d946489a7e7f127d9933e44a41215c66a49e9408937c720327a4e7b
zc04649db57255b977f63294977c3640f4fac080b6b7598aba6c61b0eafe828cbf3e33cdf2e232a
z3d743bc1826da9fb4c1e4e08930c091c6e9c00fa33498881776715bf777d7be525b9259323dc20
z5bce411579d14c9a64a5167330a3ef04913bbd6654c51d08f027657a0751aebc6410c17c179c07
z849503432c9ed9ab2d71a38be313f6d07bb719e2526bf867fc1e62ec031dd88bad3946edaa0882
ze6172c5b776721634b1c1a53cb1ec6c2c6dc06c713d9a706fc4718ac9099581b170a5a6f68c32a
z39e3c73dd6a86dcb74adb484da9fba639ca4f4a5d05cbac0fad9754d23d2f63d0da8c61d19f88f
z6844b1f298dc710a3673bbfcea0273f7e968aaa16b9c8469bbf3633a04ad1ddb524427242e3f2d
zd39ffe0a5935a019c4c1b2c5fd4d68b1f95a9608aa7126c96bdeba2ac9d245ea8710eb9ead351f
z309e484a00152f153c03767628727cd5452abd186bbb40e795679d9ac97a71e59ccb2ad08ba7d3
zca02ca489a65b66dafbf6cc3b00b453d50ab2ded08897ee24f6389576afea9de305697037ae448
zf89387b148cc8ffec076965fd19101469f034d176f3278870bd3b7f50ccfe6e3ead97270655d76
z82a423c71ea90aa8c3e09c8bea56e76436272966c34a5afea9583f05b8ae3870483cc234081c96
z498cd075424f05dc01d6376899623681fe682daa6701017582a45543880aa619445eabfa95f4e6
z5a7c8f17bad9fbff287842ed837243e2f6b4015d7e24016192f78a7d60958f992f7feb865dc1ae
zcf3fdd9f9a36e8dee82e1c875a515d7f1e0b07aa6e15da948a97bc21157c19c841aebab3429e5f
zd5e4e3f3124e51a2edd110b9fb695ee83d29adbb763643dfc6ba7f7b5e5147d8b0a728896a3405
z18f2d9d2409a66ec3034fe4b2b65da3e9819841433662167d366072f4825b22ee5740b69778569
z2d9a5a2dd56e2cad68389efe1da20a0567c439a0bcbef38256d68f80bc16e7b34422d3826281f3
ze1237282fc06f66b003fa2b64563982357e8154ba98e8f062d6a4a4840257a683546769216bde7
z897b14ccd2b20baa82f1d15f91a156020f13f53c9a5638d375f8da56f63d34eebc645a9b242e27
z86b15b906edca0003ff2b3b5beaebef578cc03d23a90ec3acfb7655fb68b1c21fbb41ae42fd4d2
zcaa17227e96c294e1c69d82bc6054d9d8d48df4737b2c3cc5a53d48a1aea8017f3cfef6ef63207
z730e370a15334b2f3a042c56c0c7d8455bee547dc7c7d8701a2da2f796cdfe9f5ca2cf8feba79d
z47156e73ba4eaf27a1ee7a6aaa89f01cb13c9cd1d2d667eec09ff42ec491df4dbc8f61c9bac691
z42003ff0cc7efa141417f8f9fc0c64913447db4b7cd9f8238ead5071c6efbce016f3b1cf087704
zbef2f95e8393017e1eeff2651f678e776434d623515fbf46039948e242839a6a96541966abd50a
z21e0ad1019e667a207a867d2dfd6a78532583c7bf118d722a005d5a1691cfee3a694051827970c
z7f4442754008f893125719ee82bfe98498c8f796f925fcad23c0c94505e0c97f14ade89db1f853
z59108d8b154c1b8619f5396374282e7c76f7b1bdd04cc51690fb51ae6a927e4ebff2d60e366f6a
zd8c44c0f9b6f964b4e0b3a0cf8a05c30e5406368e7553450a69b3f4b4d9599817b898241111624
z591ae24aeb2ffc5554c96ec2a7c2c5ef23cd1cafdd643fc3a07e623d99e9b0a1879c5bdd0a675f
z86d27a9a75afa9f0da5ba99827659d2e45627ab71ea82ee869226cb74c2f8914b8f358807597b7
zbef13eda7236d5d4e602daedca447589fbf83fa9f947e627529efb114a699bf0aaf1cd76e54fef
z82283b64210d2e03bc276dfe2a6b0a2e3042bf2f78aafa91ddae220492f8c47591ce51b81fc7af
zeba863c594639966c4443b237313f4e4777e347a47a82a700ac6069c5a918e155ce21954cf639e
zae2aa977376ed6d4ab048e10de92fb6cc5cae4958502ca5df112dce95b1d7d25199eb1a6a3cdb3
z79ce5e8d0b3d07988fad03ffd3fc073423b868e229a81d6152c37ed3f7208a83096d14fdc65c70
z70e25c05d61f04cf3e725142c04f1f7a561564d2391c48c256d927fb2ae1779382e4641141ba7f
z90caaa7c58c479403f9ee17322efc58b5c349873d9d9ccdbf5c8e9a65fadfe50528e4214b24337
z67cd3a2464b4c512aa47a961d83ff7c02da34eafe4cd1a710b1ef5665142e6ddab38edaffd8633
z02bf8ebd20ff136be35f2ef18868b24191cf05aab1d5dbb9e2f1ae69220403c96dfd8046c4e390
z365b66fdcef1ff3b5c50bb3870161909fdfeddd8769076bf9666164751b95a6ae46576af15ccb7
z119ed34c8dccd1751098f3e95be026e44050b6534f8eeeb4cd85cb709d41e057993af9d3c9e1df
z5548f692913b3af97192e34b0e384a1cb320068f8912575cfacfc9753c795c891a062a19fac567
z5ee20f05e9a07babe199d329399ed54297afa07a5f099ca333e89840967d25c819a8af95de6520
z1dfb4767b75b0b30562e85276ddfdb71caf9031f9cfb9e3c975104b7bc463d592eb355776fca7d
zadb41dc063aaebe7ec97d119ee4f776b796b8b64cf20bc7d105de2ed7d3ac803a9a63355fa7918
z2787f60e52d451b472968b07c5a0f0b4dd4024808977aad77ddca7f8d440ac6022a844dd0f7454
zdd7e2cfdfb7f32b86342d3f89eb48856222f68e38f79007680b6f785a973fa67c417cb476c047c
zda1337f4dab2dc20f53f732077b6e9c71364c43680721fbbb33b56ac162e9d0e900f73c7d902c5
z70a62ba3bbfcdc893e66d2cb97baefd447c0e8d444cf1580e54abf31c04caa4adc6f39a48af678
z4b0f49bbdda485cbead091c98769a79b32538c9103ddea17b9c2c0adb1d973de6c22fcb39e92de
z0197fdcfd2620449f9480b23a34df91f9450f2416d49e743331e6b30207bd29b023f9edf1abf99
zb5338b0c216bd074c8f572d25ecca2919cf1028c10fa9ea7375dc7028d5ae19dd2011f7ea8deda
zdd577108f25cde7c918c2bbbd7a0e8454abab4cd57edbca0d5295a421d530626d312bf64ba9c60
z1d91e0f41c78d34dcb53ce892d7a7256a3e04b94b04493cfa8a1c4ec52d886ab025bdf3cb31234
zc28e92cbb92a7fba9fd003a9bc076dda54928d1bd3b24d34cbfa1dfff74a6bcbe437acd5054e84
zee22e22f5b9566af3c83e2a189a956d80e308e02fb29c61bccc60e22aac91eb745d37ac8b500ee
z882b61f013a27a500e300c47a95b3d325c432322bc5640186e68015f6db882f366cb41c279b721
z14791d6d4fa270ec626f41c2c0f506ad178b2c4ada410cf34b265fc66d7018823cf641006c1b52
z841096aae8e359a2e76806d3c5d20f30899d64dc2dd8de774349e9af4015717c48f9fa3df5d466
za8c3c7048092bc64194240da5dfbf01e1082023e370dcd9cd36b8ad3a202ac3c771f841857b94b
z5112c982bb0d98bd847d3280f0821cd3f7895a6c7aaef1bb1e6f809c6048dfd9e3c8a4164e5544
zd4ad1aa00fc0d4576b247e5493c2e836eb05d7d543a3cdb352ce7af96783e569d56769d0b18b26
z8d66a69509be0797b22d57cf71894a7518c55176649603725d714f4f9fc4ee4d83eabb94890115
zeb7fc3e1a1aca88586c9e1ca07a3d2043310724087f72ed52e5c4ee1b3cdf3c3803cab6bac9b98
z0d06fe7cc187a490a65a8520b94a4fe25eaca946d7a8d57b973849effd425df13eb095a7da9afd
z5cd1b990b8e218a5990bf7a97e6c55dc845ca821523969f7f675d6c9715a6e1fadf270ef7a7bed
z21c564df5f27a96cc9675f76221fc3ece35ffccfde3cad36641cb658c9d1d9ed2e59396c81b717
z0c8ed883af56d16ea4c91fb76512503d3c2c1fc67ddfb9c3a98862d2d14e5f0a347009d68b8297
z3bc36c761f91b2d7acb5cb5e4cc8a08c1f26366fbe6f7dbd1ab5653de68da3e7c1c0f83c09360d
z5fc1133e4b5ba305ad4bec0ef3c3078d30e052c9da67d932985a1a4209a52252c54d3419ac733d
za80cfb2679c755b5848e81a35fc1833b2829e64a4eb8813ab9f0bd63ef467178f3168f5665fe15
z8652ea97368e3483eca4abad8f22ad97ef3abc0b2df195f892ce42272471bfadc2f88f2c834476
zaf7a93b2c8f3e868789248db4446e5194e75e39d4cc496c5bcc2f97101b10ee7885248b71c2c0e
zac2565d24b494fb4157effce3c233e32ec2a91960095935808f3453818a1f3ceb852323984d658
z95cfa947b0cca1873d21f8e95d9fa22fa27949723e96e1bc77b2479477db3bc1679062bc539b2d
z2f2ac261ced97950a0ddc255a47049c6832820b243384fb5bd1c58335ec28f04b93aa3272bebb0
z8bf172dbf08279d2c127a83c57c24a09e91f0a3c5f1b4090e56c3a34d7f214869c708683d8495c
z7e6dec2816314230a5e1474684dbb5cf144e745fcc36ea66cabbc2a680a28de401a515ecd96406
z8629aee182dc5b5c95e1f11d13af8e79c64933a803b31767667fd6b936669ba3fdbdd2e7635116
zfbc2d6ecb6698bfce6a867431db71c7f192991ea3e5ddf81a9a390e932565b8d0e6329593984a9
z9ce589ea61c4af871e25d0936a56a2bc54305515a46d461dd9cb368fa00c3c8f5f5298d0241e80
z1e45c2baeef9ba02a3d02e40dfe0fead03bd612788ff75dd0b88bbdf7985aadf271b20a0f1c71a
ze250643c15e7ca706e7ce5419a0009a4ca37f5bc959c39c3aeabfd72db1d407ecb5b24276a4365
z57abd8db25b584ed413e39220fab9c7474c6029b18538df6db7febad35e2f96f0dd88fbec8fed4
z334ddcb21006e888fbf096e6418a8545658cd639c1e9fdeea5554c69dc36186e7137876d61f79e
z00f709eb098cb0eb3e46dbcffb9962c28baeb104127120ae08a98f1d2847e5da1f35c9ee82be4d
z27e30187f28ce8bb24f2b95997ce29c2dd2ae6c14cfd8debd67fb0777cdb99616da9d0597696fd
z57e6f61f1fc0b1b3e2349216dc5e59c3b4f662ed49fda89747c3484fedcd9cca46786634ea202c
zc7f6656de896863ce30c660351ad5312e64a7a5a1e7822dc8bcef62b7e422dfce3e4090ecd3acb
za97dbe68b474237fd035d2bff0e51174d61e9609ec061b9788b0b5bb17effecb7aca8397d184af
zb1f7f30cf5088f08e61f94728bb047f98158c51aa3078ddeee66454bee70451a7087cfc099e66e
z770f10719b48c5d500d061dbbba3d7c079d306f2e2f9fe61df99dd1419be4ab4f6859d773daea8
zd1fecf57740b2a1b5104ddcc7ff2216ce46f78ff2fd98e73c71b3edd5f2d9f0cf3bd3137a29012
z02d4c09637b8fedc2c32413937fe82f1ce995ed5cdcc665770ef0093bfe26ecc9514967704853e
z67f6377cb1f0cd55edca7fac83b7935dcfc9545e2773b20b9fe2a91e335ffd6fb41d3d85622974
z7fcd5763340a7873ce5c1767d0d213a8b5a5cd9da833753f56aadeb10a0d2aad7d1371e97ff2a5
zed6ae3bd0ded86faa8a880532e41998ccfcb256afafe15e398b383d42ba1a1078b4deea9c3564a
z94fa535e3714e7900034afdfe8d1c39ea09d3175444ad039b84f658a3f88aa4bc524aed4fd029f
zac393250c1545ce77c7275ba67dea7029f15e3f3998005ba64faeb3ff515c0973ec062cc004c79
z8fcfad260e55790a1699e6c0d1b66452d4eeca40eb012e92d80d82eddfefcfa78979a611e72f36
za613c27e7f8f85037fe3bacd23a79ec52ef0ab3d03950b2f9dd10669e28affd7e28b891d479a58
z2f08eac5f439a1759ef4dec150b2e61fb45cf633a9ac0b96d023421c6a43602522562c91415d9b
z8a80b9bdd37a12b416950099b6b27b3a10f2aff81748dcec622a990e19d69acdd3dab9597c2d64
zfa8b119b5c3e983d0643884a52a42a62fb66c85adbec744c2a00581915fb5de82ea0dfb9cfa427
zd25208fc1ff9a31c9692ebcfcdce864faa472f9332c2c6c2d1904022d9cc25fc2e5c2fceb49132
ze3fd7d3b8b3ced5ecda25bc251525797acbba92aef820f57bf9cc683048e3e141d892ea52d51df
z931d6b31685d89850fa9dac4e77b53cc5c5d4dfdfaacca74a18f6256ee9e9e740eb1545b0f8518
z11945de14a68a961a5868826803dcc71bbf630927d6bbfeed9d9120181896d5fe682023db7498f
zaafbe124c0342691ee41985b70bf3a0d9b659586da6239a220876e34113915d189f47c5fdb7f8f
zabdce8a86f8372198965089b24e0893d2efd37e323b754e7662069a46f6d93e415f567636f18bd
ze21cefd5648567ffb749421bbefdec06bfc2231bc63bbabad5480a5a454afbd08d876a37706f99
z4d964f1535a30014cee79b6198f41ba1378d6fdf2b9a23e6a2be2fb0543988adc0e9ce7dec45f2
z57a90a3416d5d50e64755ed92980184b6519ebb84e126fac0735b231604d213c1b79d8ec15e897
z8621c5de50f78780413729708bf096ccd67ccf14f8ae2388850067b8312148b3ae3e14314bb725
z0c8718f005d90a69814665526d3b81168c65370d3df59dd2d5fbf7e0757a4bab0eba5a6a33b720
z647b4061685055b64fdb019ea976fb14ff07c49ebae74b2b147a3f5504366350ca0580ead291f7
z7382109be2185771d441cb90765d4e7fb78ecfadfe5cc943a9eb48baa299c5244592b6d8fdc18c
z92a1c54c6ad3d243ec26fe8270d286bfcbc9cdc3e6c0b39cc9af477a2ced496883c174914c7e40
z4be2faa0347a1616912944e86e0eebfef3e12efad98746d1d3a13f4d64bbbda7d33062443578f4
z2db591a7650ee2d1f6b8b9699d632c0b83f6a01509b8e9ed09ddf319d4fe49ef311e13dcbf0644
za1a130e898a95e55c07e20487657351496e2bbf62bc9ba88bd117acb091f7aaddc44aef52b886a
zc82947fa088a7cdb3b5977d9bab53c50ac8f0123fb0af7d51b1958cd38256264d588de6ae02736
zd9a4615c564e7802ae1e82f9fd232d26f99e805c491e8fe09042818ebc974548a59eb496a5bee1
zd7dc81e5c58528752675f3f308c563e5dc15a2f67822a86a30c8419f6d0b3e97cc531d32ca0101
zc8a29ff275ff44ff4d52f729cd2f1e0acb27a75ccb13d1fc07c22b83b34f5c4aac5fa235603b0f
zf81992569481686f3760f2f98151a86b4a1978ecd4db1743ea53c5776b556b04350fa676ce119b
zb83c6e64a2013f63dcf3bc74cc14cd08ab763cb3e741a24feec1f28483c4ad285c8f1e825d01c9
zea8228a0595ae01635d77936b464a3e268241f8129303ad8993dad06c2de2426180dcb149204d0
z0a30dd4d6c86a4c209c20cbf740f02112aad61259c23574265ea1f284840ef5d21fc8d7e3da860
z3e4d0eb2b9e86c9a5c0e47f0ca921e567d8bfa637b45216f43ebeea73be8aca6808326269c1adb
z9c21edca03cc9de6404eacf0e7fe7a60045e9c383329465dc0e8ce436e225ff14c0ba86d8fbb72
ze3ce665bc1ed2a0107fe8972813a7974926d7ed3859315be2c443ad0e4eec74ccc080c9d3861dd
zb976b93e19ead7b74bde6ad44b8cf85b86aafa0dfb172ee257a08c7c1927fa132f9458c6ff547a
z9256e75fde5c13a7dcc74077e984502a85b99fbbc44bbd9bb53284d7eaf9e16602f9b8fb0066bd
zc6c7a02b34c62f80ce60e467fc4e34d3dca1f15e61925a4ce664f89989a64987a0d43e2aaf79a9
z04a40bb987325631f72de9aa3d72c1deafe69ec7e828e4844ba19d33d23bc6bf27fe41d698bcf3
z80e7f0e2650fa6c1ca68b791ca69ec7ed6b5527445a9d52ac5e15c89bfe39bb8cdfbdc3e736ca1
zf945b37060b9ac8707c33db89e68e7580b635abf3ad96eea8b3fc7b5b8f77954761cfb8675977c
ze682ae2e9f5445a5d731a30255c8fc22d1b48d1670ac6e01add5082e29a07164d1918d9b4804f8
z3b43d40c0f2f4253cda5b013030862b96d30dee9c7a9cdef04189feb6bc4ef4cb1ce0405a333c6
zc615f2151da2147167ca59572a09c696dd93fbc8c7120adeb5982587047c35ca221cd6f85011fd
z23cff69b675af1882d5804af25ce879bfafb2efeba5c301867722e66f4d0cf462bcd3e62a4de1f
z35ad5ced78977d60229c8d6cc74b7d8db5f069df7e296085f75d732e9721397f18c64dab808cf8
zb2a05689ceb830517582516cad271c011f94a391913c2e8b33f1b3189c6358eebc93a4b8092b40
z696d490e4afc115c77b51dc2f13c5a182c84a0975f8e5cf9ac3baaed000a11a8d5b62fe7d92ee1
zd6c605e4713b663c0f285b7471e33cf62037c41bfe2dd5a5aa697c2e9b04e25881b8855f643f5f
z76e2f27bcadf19a97fd34023c41c3a859812a1f3dab1530953bb51f6c488d0b2793276398c8337
zd2960934d7ce36fd6524c44cbbd1921c3eda26d8754f7d3d0afc6a360afd7779d1986669096cb2
z348ed4d680e02f3dee07b12c29c395c1f147c7c2117681a7b2e125c0cce056bd6d38fa4fdd50e3
z0bc5dcf9d605908a6bbcf6aa39bf520c2859fc7ef5a5af4ce57ed99e34e86680fd83ebb2de3c1a
z657b7af953f7afa792b3924d6b7515bf3d02e50d4e2d4e7e9a515cbc79b7f202140cda6b9018ba
z170a755d82c93de51a786f8a9bc1c1330ba7a48c7378746f035c61036e7eff40bcbaa161d159f7
z40a5f086b94619841855139c7233289016bc41424dfcd5e6c8a4d1e1f8f1cb69cbe029c19fc36f
z9e4b74e7c0dcaeb9a5a75b33712514553d95abfc04e11615ec72a56cb5bf8bf5f4571c0176ad15
z3aa83f109a4342165abd4a256a38ec3d2bf97e9bbfe9d77922f59fc0dc81638bc364d814ba52c7
zf88dce33dc052f18c7dd3e2e7c0d83285f3ff2d077894bf6ce970b5a83100c5c4be5f738ade922
zd3ff12d467d4ee41b73aa5b7fb8940472ec8d1944d4ba486243b23b51a11dff74b17b12337a1fa
zf7be5390d12822cfc2816a73f79d135ba94ae73efc2dbed3a418a7981a08ebdff9cf528af7f460
z268b28389c2e67254cbe1878d639aab372a3b2e30370c44b89672c2a961bfc21ccff05626ad6d8
z2aa114b05ccc8ec44fde4767b6bb59585ea88abd897bf41e6e97451a47708d3b0958af93ce8823
ze842ab5ef95fd2e0cd1070898a93448663a16c2ce2f9ee3cffbc79a25ea2a823ad27c60cef0f1c
z9469888d57b1b484774074117be81768a4a71a4a73286895745b375bf2e1ddb661c280fc1d0013
z0ca14fce45ffb84861027d71bcd9ea0453383266c9fe3298db3a9cb2a5f6bf2244ad120e9d24b5
z925fa6587a3b5651ceabbb404815e84fa7725ee615e1e4b3c3a0662dbba3c0a14c4291fb6e8b4c
zbedb1489d69ff1a3d92f3ef2e3d01d4a4ea8fa14e868a0638212939c73e8ea13ebe6133c700c86
z0e033e47574d35e48f9452d49ac157ac1d85d32168cb431c4a91c40920ad4912b723e312b04d0b
z57f05b118bba92ea460f529b7c5c4716637c3005b279974d61e85c46c5caad398ca715bab8612e
z678c58f7d99182b4799e2f92a3592d9f42d877f2edf802ed4a7ef9cfe27023f505039549a10104
zc311cb772e0ef3f4c98159360c0462d80e75cad2f63d38f4392572c19dd36976493c34297ade18
z786afbe7865e13135357d14ad62ec6143dee8b10f2b7770ca93c2bf1ed4b6c3623f9b912ae6714
zdd212943c129101e911957370b84cf653dab70798095a93167a1806ea9a08393a41859a82d057b
zddd847b3f2ff985fdc41a1df3b59f3139bfc66d336ae2eb2e91a5b3ea1cfb6e1a97b93a27267d9
z44894459e23e717ef557a066cc1a9e3830f624631b7e0c37e03e366ba92e2f1bf8bbadaef6c7d6
z21c7ba3cb661daddcd963bd79185efeaa1c7b9c46ff7418a3a1970c6457f4b0198d3f5e1ab6bb3
z92f50c56005b4bef412f933060e0e5e32b8a5f29fe603f9da71053ead941785b45f269b5fad13b
z46ac17fa33416bb4bd9901bf7fbc9e9d903f141bbf81612fcd46f8edd4d95631247f08c41117fb
z0aef426a4e7e5e5886e94d1c0df6301c5d218f82762b89a0829d9b688ac7bcc60f3302569ed3ab
zcc0b8b5536f5957e07b78fd6ed83642a29e0939ff2a00e98cdfecb17cbce1138691307783b76c7
z812fbb04883780f72c14d094927d2755771457d4edea7f707d3835f067f2d5dda86af2ba8e3a5b
z8380017415b7be020e49c161158ba6c934f2bcdb85f6afe1519a8d009fd3051627379bca87e141
z5a8871dedc38e3388fa0346d1761b8e8e829b10b96aaa4b8248ded21e42e190b191205bb26da4b
z1aeadf60b94051a1be9dabe104538c82d272bf99d2d829edbd30988ac8870616f9c047d143919f
zf2c9804a7a9743892cd580665ae936978ad6131c67063814cc7bbca73bed25f48ae7235bb4b481
z5dc636f443941e8a55b41d0fb07173b93a7c08b34b2f685bdba3db7f70f4167885f2aa53d38c16
zfa6be81be9fb805b7b9aeffb13c5ee6cb63e2763cf8e6fe72205afc86fd0431edaa3579fcd4481
zd98c53fbf762f2cb7641319b11b366fa868259c2e99c9f80a44b4a7c3d8b416df53a3a696bdd48
z482755ce3877ebe775aa0456f2a8a1e02a4cc945c2f1825fbf50c2313378d84a9ec48473306018
zd7b33ec785bfd737f0df20ee389a003410510fe64480e068a88d2a572b884df06572f33069132e
zc487b45e90325f5a3b0613ce782c29cc7e0840ec3000bcd887e01311c481602ebe74d5e106452c
z5975e9ebefca323735b1808af3728870ae9fa0d1dd418c58eef1c755515edaf97f863d3b7bb1f9
zc5715ed76de250200652c8f53c82a195d6f5a5aba15995307fe4641878576d9cb3249829eb1c80
zee52936a3f2e50226bb05056617cedcf851c7bf969ec116275014f882a9112de6dadec20eef9fe
z86d0f60b8ce51766d664b0c1091528075f8191e12e0e1d3a2f88fc9902655184990b401cbe3473
z2aedc04037c3e21b9435b5d6f3df31be3aa309fbc9955df8d73d279e319b2740f4bcfa72cddd3c
z68c6848077105abe71350f907e3d4dde283fa4c5474124384fbcc403679343cc75110dd667ff95
zf16cc2017870b33075065962d5814a6619275acfc8d5648bcbac1dd2e821b276b00e7364cc57ae
z3296d56610685adc1cc60edd57d4acadaf3977c6f0fc86643f9df87fdf1d5ad7938ac01cde7ee2
z9c35f17b3fb82635c0ee7a76110cd9afb50e5c3755d2e1d90037403219b129227287da9ab48a49
zb9c99f3ff1bbfb72b94e57c44075dbee9724ddc736897b3617b141652569c61a6fbf4ce16d8d70
z6ea0d9ebd0fb59cf85a79d4c9d32978aafed31e00511a3eee48665cbdadaebb4989068d30e10fe
z04e3f9ad72df37986258767d49805c967908e6948ac7c6af5150be033b5f1d6e4375f4ad17b99d
zcc9ffdce35257ecca46582388a458e841473e22b21b07f060ab47a2d4fd13884d183ba0f8286e1
z2dbce44f96c2fb52030ddf3e77ac82d937bc1272f0ad8465bc30c79a6f7ede91bc8be6624d768f
z2c0133a3b767d703bd60774ce537b25bc31de91c35efff5eeb76bc59b9ffd28c9cc27de9a542cb
z5e810d123bb8c1966c44885dbda95a58c273b111c870644e3d98a7ec2ada6b2942f48f5fd85e02
z2945ff548b07d06fa1fa46e5359936a7bbbe6990c33c90e6580df51b8beb36932be7ece3fde868
z82aec71c6a500da1a309a5c802cf31e56dbeb3ecf92d5daba6ca35746e4f895f2fdb4fad2becc8
z7f640a6ae2edda481a315ae43826f496920474eb5fdcbfc04552fe6cdd17f7d505869c5d61a76d
zece061304ef81da12983f1c0b9eddbbde2d05d0edcd5ced35efbe6ea006a341bc7c6c5ca505715
za8fb66e4fee6feec3d0d0d8adb67c679a5e162eaa209964a84b0afcdc998ac61bdef3a44e66276
zff9b30fab72460f7bddf2c5e03a111acd0a9a6145b0138101cc9cad5092bff5c719ebcf159c0d7
ze344bf476fdcdda358abf1b80e41f3a5af146082fdf59c19064f6aeb0c817ccf0bb88868ab7a3d
z4cf4de3adf05c3398932e1d715ace85a3ea086e94853c9ab2438be057a02ecc2b23d9e21717374
ze5ee7b9d09ba706c140072c962ca0a7c47e9a05535c7f1576efd2bfa33e5439e08ae2506e765aa
zdfb10435226b492f453e16a47c6f45edfd48894eef36e004ee839e8abee782773d1c6b835c0928
zbe53713dc4734397919a8f06069572feb067eb0849f974aa4fd80ac41c38f17bd596244c575146
za7987b0ab4d8d98e23c36605287bdf62f13e68044035528fb2b85f0d3edaef2f3eb1405739acd6
zbce0a81eec19a34a67937f5c48e0eb503a51abac8333d6d44bf653f7572e620666b3fc40ca505c
z998eac9180a159610c03fa753f7e0497b125384cd394b4fdefe402d01b331d4fcc83b63e9ae651
z0c73d02410782ff7e8f17104a65ca85f95c40512ceccb9fd638f22d6ec8b3f142cf7a2e6e84504
z628a0bbb9506fae42f121b1b8c584a582f438610ffdbda24fcd2782a3a56ad3aaf01d9df784a33
z9d61a0677a6a3293e8afb9b46c46392610e46ce3675cabbc538863910bcc5fa0a3b93f8ebb5756
z64329794f973efc431c9d00610d6af948e4081d26e38e051fae7f19938c26fe6011b81ae4bdec5
z3d2f8a3f094dc723f726b1a22e2c676b2a73193190e4418a337afef11998a20e61bf6879427e53
z7af7e7ed1e424c71cd92df59338ecca311837673bdf615b872c84cd7e27eabf56244addd20ff99
zdd3c9d008633a3cc7b7c85c3cad40ef4dcadb156463bf405f0a233992bbc1721719e8f62a9c7ef
z92494a093374bf844ad5cdea95f31bea4c0328e850a1d98800261b251ef4f16181462749af0e93
z4c2b6afb289b1c47e77c328fbb7de9851c82620b90b35c66b79ff6e7c645be1bd8865e26d8667e
zd0106a27694655b07de0100e9ddcbaca4decae1ed05fd9fdb4390dd638f79ae0b109cbbfff80e2
z24926dca5a6564551db70d359670a3a008fde1d22fa5987a623a7dbfda0c1d8babc5922fa98018
z2a16cec14abb92aa8d00842876b6e9d2c32c9e7eb64016cc715a960b3d08ca33c0c81314ac6217
z5bbd6b84dfabe876e5c2d6b507e0e938528ae003d0396ef7a7c9b9bce667db8c37d572a99a8a5b
zacecf8b28e6b7b656954eba5e00a92a1afd22daa008327757db7bdb1494b7d8f4c023f7c3b9039
z8a29c2673fd28af49760eb7ade161573fc059b407d2116cdac0a92b579c74a2b4083da3eb96f3d
zf29f83220b8b66c8f353734a1a19dcb6f796bd4c90200f7fdf64f8c0230c4f2d6699bff25ddb47
z59ee5cc36146ce1eeae6308a6e8a3a9a7e41135b672a05ef16c13ab4f902b743c85d3760aa9ca0
zee05c434bbc33026a25d2fc4497b06f6778b69063b06041a977efeab628ba2483396930089c378
zf80f0a7276be422b46c13f351ee631f1befd5fc7bcf6dbac0ec7aa0fa94498684e7d079ac07e5c
z7117f0449d90b2512e617a8350166fe84b21145d05e9f9b940091d7b7be0a0c90cd156c8ff00c6
z81eff42220971e792ca3e681c73b8b36a888cf5c1a1f745ac7fd0c02e81e39271d49fa154a5e88
z36f83c42e1ab5367d2570a1c948c3935cf24fe5207c71ff9a6b680bc4887b70dc980580abae2e9
zf5eb1c8a1c676f8268b2e0c63f82f19d43b8c231920cfc44be47745539bacc4875d837c778dde7
ze9fb99cd7d9488a4f74c32fa84ef8e1d6607d604d6a6b7c46fa8d24743067dcca1d8fbdc8481db
zc29480fbca3049a50acd901fc22a86c56bd7744f1b127bb8685c4106b449e870e1036cf011ac09
zf86af941a0a29054708a79e6ba9de48f0b283ee1bc51f566bcbdad114c126f925f65580b46eedc
z0ca7d9107ffb1a642295d40c2740ae4e7056daa1ca8a8552ff9c2129240e50b8c8295b2f100e7f
z6da8e0a12653029667aad08e0c316154b8d37c751e72b73d8d569c6fbdbcf4de574114ba766e1c
z4bfc496538f18765bb4541daff80b105d071d598e37b653196c45cafa9e417ccadd46c27b7cc06
zda5b0255dd7016d43b7e3602c7040c63bafa88850edbf9aa3083196fb63fc8efd0f87b8acc9363
z4f1bb3d04c62b769ad338e12f1945a8a6e35d9b8b0379d8c84b07081f0356bb84ac0476030852c
zd045d04c10440d49731e51790e49620ca9c9c1b8877c86823c23aa2f7f49ae5d9a584590e2129b
zde9f9b1f84bc0900c430fcbe9e066ef867fed40c3a8bf2ff1d46313f89188afa45494372410322
z87423c3601e15ff14e26d3e905b3b7d3ebc61af831f861dfb062f54270534969d9b54bc0c7229b
z6779a9cdf20fa629bb57a66dace6cc5d96a6cda05f27bb9c48b80e7911c4deae3c03e1324bac45
z793922c9341c6ba99ea8efbfc7a7fb0f35f6b9097f5d8a2070c46c1b4854fa5c2045bf8fe633b3
z2575f9a656534663faff2964de458cdaffe3e1dd9df8775942609ac4306e64b5d429b1bfb91cb5
zb370b2a4df58452d40f835d0e0f07e5fdbfff0a1aa4313928532ab056eccde52ee8e40a0ebbff8
z5aa478576f214981f188c0e8931a744c38f249d38527c89a7950a69f6f0d4d9a8af30ab371af4f
zbe83b7bfeb80a17a8dea0a30aea32cff77a3413138b7330bc3f42d2f0e135617c1c10a68fa7875
z98ffb7de950db60b0d7bb0e1958cf6e1533af792eb0e707182adad53ff39fadcf8b0171e5eec33
z9937f9c47fecf83099e944eca9926e78aa14c44333e526297e59e840d0fa6a7d83c177e495a648
z71a7593e77f4b93016afae542b6c413d734f37ac3da059c85e45614738812d29cb48920e5b51ae
z6c853289939281a1049e1d2dc9549e75aa93fb0efaeeb4d4307b41337e19d7e2781eac37f13e16
z58cd5b38e143042249dfc32467da09a680fb7a9dfb0e7b0dbf8d935a582fafae3f0a6121b82245
z46d611ea8efe4f398b43d443cfd72571ee36a0b327925936d487973de7bdff55945d25d0635e87
z8282386844de52aeeef0eed9516db01b1e619778dcb7e3fa58addfaeb27e323295e9d8e4d97245
z7869988dd76480966b76c8bb13811938f2714ecb265a48e5fa0400bcfcb52b0aa77e731f30a5ad
zf130d2d8ae3f9552efab4b330a4f14bcca7c5f2401ed9c6237cd2f0b74a78ad34567eed368002b
z73619ff2342e0977b78fcacb728d3e519b735ed566fe19cb5e3d58f2935f6a9e6cc086d5e350c6
zede4b0d3b03ee203dcd87dcb3b0df0ea8664321eaa7d2963a525dba6c6e5d794291d506da1f68e
z3346a0f5925f619902d622ce3e881ebac6616f051779309f12d621767329591e5b02a28aa75935
zd928131222b0c0a597fa726e736cd50c45b821ec8cc8258adf7b334af29eb9b1855f062b2b6303
ze7608d0860c96c1de2ef1fc573ebc9ec24c0b65ad7fe463817ec00409bba5ebb3016735f33a70f
zbcc2c1bb812a862e5b7cf6400e567e451253b1be973ef223a73281cac2740f5365d757671b84ee
z9cba4dc8284fc0c489bef866888b0599fe3c29e40748bb4805d5ccc949915d52363ffe31adcf44
z070567bbc06b5cf791d002041b08a5dba180b5427581dd15877ee55e482e30446cf4ee1548aeaa
z14a41796f9af17acdeec458bb09536e1724b555cddf2a82edfc2c6298fa95bde93b786ebc1a534
zf3e6e20b36f8b2816338b8d7c4111b6e681fa4f0d69f37ae4b78fead5226f50e5ca5fae8c14a83
zac962a1a452c200aee6b1de4132932c415080a9538bb2caa2c44759f685b401347161eb9cd4d2b
zd6ea0ca65f860623623f1d1b5f0f7f8e7dc461f906b717795712f2b76c6e37f30fe1736eb02a9a
zf8e628e078e028714af379df8b923f032c2b4ca7bbbc29441def8abfb58cddb02d7cdeaef6a609
z56b898d2fcc0c08bbd06bc48a67f8e74bb72382cccbe30ef188c8824290f3a6a5211e7890a9551
z4c6ccac2e78a0b38c69f591b0f7b57a343f86e3ce6d66970326e798886670af205ae69192d9d6a
zb691594b9501fae6cd857a3559960d2848fec6a6dc06c0323beea82c5e0666d627a0ce02a7cbb0
zf87cabfc127afd62073a60696d6360811cf5dc2a9263ec372113168efec9cf5c9a79ba2d8b2702
zf7a00f85671e56e0e2c64bafbe1a93c7a55e76d28013a341e4f7b7c7b3ef1fe57ec56f9e611287
zf2519e1901cdd8de91c91d96b48fbeb8237f068a4e5c42a8faa77b3774ad4aa12a77c7ff3b9374
z5b17530ed942e5bcf99ce985747d6e8c6b4d18b8796db9dfcda6b901f5f7b2a01ec579ef99b0aa
z3309642e7eee29ea4f41d4e883809462d6bb99db2781aec475b9e88e72b2002f8972e9c0bcc3d6
zc58ef72935addd1cab54af8306b0cfd50d737baf7570efa3425d7f4262d1be06bf7fb875c423e1
zfed9cc883ad76fc432794cfba5e0041c57b239abddeae7cd36d190325047b9fa222fe2e7ee4c26
z44651d12cd72713840eb9b89e8a7f59c99ba5edc581c4800dab6263883847da6ef989017e53e65
z39e295ec53f746809b87447f019ca7989834cbd9ca7a65eb77c103321797c4955d9f6397ec61e3
zd60fe297d44cb05bfa55bbe97791b2a1326cd0084c86fb36b5d72969bacf4131ee1b296272b6ec
zfad60b17fa9ee474238a92ba4f13df9c13a0a0a7407234a57327066f189403f1d2bc4b0647e3b9
z013d2c0639558a4174de33620ed354fea61b061e0806373ebd6936fb860c989f79045ce197d8a9
z9ce7378c572018d41497d35ff8d0c1bc89619d1510405ff136d1d913d2160f1ae14830227d670e
z663fb0bb525824de38d4a78d5b7f47a2f4c864182207fe2e40f0e3bfab1f99485c65b54f4415c1
z6ce9efe7353429bb5e753d2e1d68490ad74076e15ac4d6c870b49696debfb5991b619e652890b5
z34f6111ea51bca72f1756a97c4ab79bf5c26559114b65d7bbfef4b93e9a68992aa539aea3cb5bd
zf452d0ac85660c02a8b96eaca5b37fa5d9f179ae898952ef6771e70f87f39a90c4a160a07a0ce4
z76f0f803c4a8307e9afdd01da83a33a54e1d276d01d1523396509b4c74d0425640727551929612
zbe5252ca55577fa9ef25193c3b3504f29677c44c638e60edef36c250c400f7da9e9d0a60c56031
z4e9aec1b0a34156a5128293224a77533ab0a73d4b32f794d7bea4013d3b19e26cc74bc072a8b95
z2b9c0c46bae7c6f7f5a2e84bf1f454c7b85515443d2584bd212b8e66c18a9122c16fb710b63807
zefe076a82edd23bb95e3834b9a0f73275d0cfa64285e96aa248de9ce45341166298459701235b7
z95c29746693380b8ed9636d9e86dbb65b13a004a532d14e858643d56bd8ef7a0e40f8871532a1c
z586997e49fda240b889a483da9c39f202d0b418e1c805e2a2f8ff9c1cfe75b55498d468a3fa1de
z3b3218da3baf0585b9c7911c95c9ed2f235b3ae9d50e9431f042fe19183c37a4e96cf900f399f3
z43e5bfa7df1425ee5a6a084348d3791364a5c166e3d8b6db8f1480832c956398fd3c0bd84e94ba
z10a15e4ac9a0e7020e28b9ad608c72c019ed60be3cd512b7a109d32fc9ae081833e3d3de833094
z04115374d5003319bec72df3b8c8cbdeaa103798abadeb32142ccf814e7bc89cc9a8e770dcc3b4
z1d46ec6f139223fb3b3fb4238a9074ad1ba8cb2f9f53fe6691478b570f21a05957639e90b7f548
z8249c029e0dd01c17bc354799a310d990d8271f4a4e45fcc3ba36bae1af7b62e4edfbda5f0ec33
z6de7fec862f78e0fe9758853977c4b908c67bfe17b5823be74905e34bb3b783326f24c7a67174f
z2763b8cef50749aab9965ab215049445534f6fbf0fd4463be15d6e1f5343a34b346fe45603f290
z366f38d5a375451eba1503d108868e44adadb9d5e6e302ad8906ba2c64ce386f7e2bece26a2dcd
z1665edb37eb965ce15be49216f0d9019fe770fb94cd5fc185af28376e427f50d952ba48d48fe45
z71f3745fb8f636f8e5f8a2587998eb580d02983755fd36ff17044c70a1745e5438ee3b23edff5b
z9d878f4053d2e0ba436f47db91523c8173ae4cda4ccc0af832dab5a97ce5ff6bbfaddff3fbb9b0
z1010da7e78172634b29c74063a317836d0c6b2df58562d63a5ffacef0c75c60d2355ce8fd0192b
z84291937e213fd273fdb0fd8b134aff65946767d81dce559ee5952f9d2ba741cab77a24f234b6c
z319aefb6ff291c20abf6a59cbc8eeff6340926942453b62b214bae6ae8474fd8effc4c1a8b5f85
z39be575013dbec3c72b2346c9cc48e74d6a926520f38128d8fae5fbf4359c107895565a6d4f00e
z7f096f01200aef8732948bc20263ee917b0224e75a77e2db6b1eaf6b4cddca582445b39176d12e
z90be7ea68cf91620344779bb005e6b244b6f8cd8a91973945f60ed93cbccb9bed740fcb842928d
z12a5b2e5baeed02a77726e209e9085167d62421e02113048cdc36d136cce9be78e644b3ee73e3c
z33dcc31d3e8377083cd03597f0307aa93f96e3a9865be0c0284d5f26232efbb159dd8d257bdfe0
zf3ec7978731ae28d4cacb9f49c7b86b9f0de985b8d9c976401e14e5726f28100c49b6089015f35
z2c38ba04fe9a1920687bcebd29ee33a9d3d74579ca21ecbb36f343a387b4e8cc5fb63ce8cbdc0b
z1eb2006df3de1283828b8db518e7aeddbc7781f44c71a4eb8ca6c47e521574135c94a8a7af6d11
zac7b8a0fcf574b8da0768111ae1a97629029d378061fdb954b612e27dd747fd98867765956f2a0
z0b300232b6ca9f8166ffd13aa6833d23a4f4de812e09afc8d5fee66beec0345ec5455fc0c6d87f
z12c34709d2f06ad911589c8cf9bba56ea36cdc084d3d1993be0f7d472fef4364078f11050e2b50
z3f85f096b5c01b3a361e664acd008bdc3725f656d9aca1db189debf694b0c011554eb51df1fb08
zc014bd75cb662425107f285c9e9a6af62ebd9e5c8f23353685ce833e569e34d695d607fc29dc89
z4db27c6aa91e93a8f859531b6e9e6b376fc898671d4ca4eff2a902824d99624c7720442426c6ef
z3129a9a0ad7f9cbad8c3d0130758d0d72775e2420bf913b760d09ae32148962e9daead665d5d06
z74869cf838808aa6393fdf13b7bddea7e051da63c2bcf145f91541444cee023f9bb020ae47cb90
z60b3ace3f3f38e637410a6b6325b2ad12c95868281277c62080d59ddcc5331097f795d2b989690
z79a9b3fb76388496782a9b6392a0c1dbe43077ca7b842eb88566e653908800a0fe5daa6ff1ac0b
z244333afbed1bbdbc6bb9058d923f29fa727b17d363bb24383c02b43f7f5c53f14b739119240ff
z920427aba3ac789b4f8af47d35a9e82c32412409c600ddc4a7a4f195a479dae1af4196d551b4f7
ze66ce3011e3d3a4d91b245a77f1759953629d06d48b738e15838669bb832ba63db4a991eecc0f4
z09315f45e1daf0d6ddbffca8db34578c6466625bbaa9d8ff23e1ca100820c0d36a920bc42c4fd4
z8a0b7e426bb95de6fce673ca5929882ae35f533495f9d9c2a0ff1dfa3eae96d979fce0d7652513
zced3b67db97abeeb78afa920e32030925c17efbe63027535e53614eecaca5e8317975babdb6b3f
z6fe2a2951b7381ef91be07d7340ebc582d3fa1c5492d89e8622cf7e04d2f99e94d9ca1d86ed1f1
z10676052667f747f4ea22fac83d7bf3a5df77dd4b1aec6954e8ec6b4235495f894e207f03b3a95
z9383946d58ccfe1e8cde26d5e466bc98ee5240374010b555632ad9eeb610762d3318a9476a85e8
z421ebbbdcf2deec7f27a5d50b11040ffafe4106a4c51c3129adfe2e4d6afdd22b0d3a8af24e4ed
z3e36c85e0ee17957f89cfb956aab25607f17f6b02c485b40dab2d4270045b65a9c5b1fa2e4b05b
z7f7e42856669b88353da6e6c03dd2ec6b9cb19cb4dbb8628995da6f8a09c90f78be2986d2ae081
zb9e069446a5001b83c9d9cd3858dd7ac0920d3f23311e8bb6bcb5023ca9ea4f95600e3fa220074
z510cd14eab4a1d671c782f725dd89c15740f517a4deec9beb670960b6089b47f84b99863bea709
z38d7c0e02ecef0b17d33d11486a2d5369231121aa6555c60e681b27b1b4e35a929b1236c4c2fa1
z8322964a43f94b4394e4a2032c90b7d36e11ab77ae26b269012bb7b05f60f693cd062d048a22b4
z0035d17eed4583fc9b503a53c9a87fd0f1c72b3a153e5df31e7509383ad88f4daac9f64ed0a684
zce615a82ddec5e33c94367ca2285875ad466524d41308d96def1180c8b457e5f1873daac95ed45
z67b06c67ac80aa33d209edc479f6c0a963b779c6c705b1da6369cd8459dcaf9eecd7665538133c
z7ba43f2c5c4f0b01262e7992700332120649bb686a9056a8f1e5da00c80619662d2d875efcd710
z96de03f84728812942ec0045356d516f53478d5e01543c17320716ca7322aa7288f166f90813c1
zb5a4eac5d102f137a2cda237e2a996e1f59641b857a0b4f0bce386cf84ebcd98d00ac274a3ca5d
zad8f8eeba0c0057d6b06b467df64f87e1b7ea49fbc25f38046ab18666b4f8ada5d6b279fbeecf3
z4b98d12a7cd5782cc822beebd95066c213d5b45914ffd5a5dd684c26b93c722f157c54a78a2f84
z28aec75ab0437010da1fdfbf9385237aae5d1ff3661aa1d94518450d9ce00521d6d3af910899ed
z845aaa45956f7d8c0593d1f5fa749a3cf6a7d75afa2972b2b6b02075affd4194bc35d7c1830d24
z07f8053ef0bd8a1f9c2a202664287bcc7268fa9f2c2d6007114310b6f8afc63bc7216b7b99dd66
z128f33deef8d9c766e6c044aa4fefd14394d03438dde760c55d605d571f71c280f63b42d89406b
z10708828eae660481479c953831ffca45a1cb2f16a5bf42a946ecdb43f83c19aa8c50192215a04
z5ddcfe5a593886bd13b7b35949525d2a7eda0926a02053a93e7b01e021fa5ae5f8216c7f6447f4
z893dba52dac265f8983285caf84de88b4d570ccd1d302d1f0317e64c96a26161c2e42779f8fa3f
zd678554c26489ea7b72408efff50f4a4bc8f197582d7cbd84d496eb93d9d96362dae6599eabf19
z0b02efe18119f1535cd88f26f7769d02cdfc5c8a20066aeb4d4880cd63b8ab5e0551bad9da59ea
z7cf118c218f9b2f03b28eb7dd3ff405b457fcc7a668ed8327c73a0754d826dfb6c408b564075cf
z7e210a8c2444778b0bb0b49622b657bb5063200323111b8ee55dc7f97645cb35eef805192f393d
z0f19a7bb0af85dcd6861bd0c91f556bb9c6b265aba65954f4dca30010eb344741972890de1f2fb
z1d26b222d0000ac749095a4217d17adbb41b8067e1b9657c665c6da13771113a1fb932bd0181e7
z410ec86e32de076eae5760c8618ef47034fe1d29fbf32d27aabd51626c831b8962adf0cb84bf54
zbabd6fee361a99c639f19029d327a0dbc9208d0f69f85dc5756f46ed2ee06d47a9173bc175cba2
zb03dadcde587d27206cb7f40903ddd3497915006cafddf4a95991d9c55157f095ce620b7a34f23
z015d65ce0fbe6eae85bdffc4455e9b3be00b9995a3ef1ef775a217a05ff9df591e7776ec1c85cb
z7712c2177c89dccdc330025e3b8eb7974dafc2c6a096a8d5884ec2a0d4db0f9bc052d98385539f
z2f360032df1fdcf45d1979e7a57f71760da5b71f89fcfa36dd0cc0f11fedc39cfa501e16a2e21d
z200fa899a427666c3e5827a1e6584f3eaae953a2c7a972d86c5ebbccc5f6b6aa412a66746cd918
z87bb8e2254dbefd206823be674667d2de1675b562a88bbfde52104eea20ef3229b434de4bd5839
z746bcac6cacca3e5097942e7e3a05e32f20fcf50de4b1dc39399a607804de590cfa93f4c19b374
zeafc1843833a6f42f2905c96ed6fd9ac6037621bd82c21874b40b7794ed326f00b7ede11b69bd2
z656010844e766b2e76829c33500d4af6fda01fa0eb5007860abbf3dc10ef441e9ca2b6b72544e9
z3999054ee5c4f1df6a5ec0e18d196506629b54bf7a1d5120c43d9b416faf03bda2388c4175f025
zce5162641a745a0125a41707af78cf39feaa42f95e4558a72b5922207af8220ae79c03b7e58190
z9e9c81c57696fa89a6055a3d461cb9ef3b99eb35f3f693b071c30f38a272fbe39e1798074ae51e
z6525768eaf146fd75605c975f35cf067b02ea0911d9e13423ec4656cff02a33e016a3f6787ef92
z01538b47e8369970d47fd9c125481b321bec0ea0c7c2e6a9939de489fd761ee68c13586288ce42
z37c6ccf968ceb8ea11b55447998fc380a909e67dfade80616569e762170380799c9f0a4146d933
z3b113657ed46bb5db821b0ed7bcc9ac28c13dbcd26ca8fdd6aa6466a5f647ef36f611e4c1036f3
z55c8a6d5e9f461fca0719ce0a5510be3a66ae9ba3be6a4b91957e66e2c4a17d3fdf6e3a6e4e9ba
zabc3af3a4eabf34d03416f4c98acb270a619fb5e1740c103fd1065c74e2b293494488a9264c5e0
za537705c970c5f6b172256188babd5f13d366aaea5b2759d260130755c04b407421961cdbc0dbf
z25c727e77ff5dc065ec73e72c45d0024d3564d870579eed720b788682aab875ad35b9df43b98c5
zacf406e13c7b65c828631732d7f9b358e1c622b40e980a6cb17024b6895e8a214f3d0364efae64
z98396cadb31706826dd4c2ec70963c0a81ad96f8689f2c5c2c8cbd9f452c76f928ed8fe7a8fadf
zed30ed7a916ac0b6cebf407f3363cd2233996e01d5e5bf16f9b184edd78478ad445ad4c5274fc9
zd919ee693f1c98cc3c16d0c500620cb0ecc5d0aabe769e16db15e54fad4d82f4acb8176a31f280
zde4366d8906d31a6855ba1d4a4bd81b5e4725639788c7153ed7efaa5b010153c8d0d3bb19215c2
z2e1a736f21cbaed844bdee5b0759ce1952b625d80d37b411ff6ab427d5b82e53e1d03bd738a922
z18aad29b4df6bb0b2e70d077e5fc9001e768f5a465d836553117d136d2971855a4d1f037db45bf
z900477e063f2e035ad30e6c458b86e48a3149119d4c9515cb3c01695eb59f3050d6f035fe3fffb
zcd62dba4fbe35227acc931319d8f1928a75db7e5efddac5b9fabd294129fd3a012775d8cc0a33b
z7f0ea85874b1c53cb8ded6efb24d894c8ae98a8d7c677b7e0dab4a1c185aacbe0c1b7146ab9add
z627c297aabdb9891ea7cbd9736aa90ca2b6cc68ebc93e732d752a6e78197b9936db1937faabddf
z23b16aec1445d01800efe2812c257759c1f67953354343955aeab8812b5c443a9c3787613c0f5b
z6ba23912c2f1a30809726d5b147fe608d704020d1c0ca361f6ebb4a80250cdae72903fbb01702a
z746fe42b58500a67b2ee8956c44424a72d0f44323d7725007a8939d12f01d17e7d7c5413a522ea
ze6f1885747f8c46c80952c2d4d0e7854c88214072eae26c4780d7fea48cb0f2353cc1974cde786
zc0488907c92e1574a0ade75118a15cad7451a1a467f24c5436867430801bc9f74ef82e0e9300f5
z42883cd2ec8b08b4d79f40fc30707dfc2980cfdacb6095333e034c5732b5309ecb71f3a99dd1da
z7da69170ca33deb04d66fa9011f5902a3cf4651d97da15b5a204160a8335a95ac33b40586acbf6
zdb711d06dccaba7f797d2ac64f9300558271dcbeae7569399954a9faa04f0b7ebe254c9e78f2e0
z1bef5619b77394b8db803326baf84bc390fd0a7f9ec78bc5dd2c2af9fff027df6b0d2dfe3117e0
z036be8b7a6cf046eefd6c2af1eee829c00a494dab5c1a55e38ccee16757db96bbf2038acb5c177
z8af6ba4253e7b28bac3fdd7f39aa943311b2792bd1879ec248fcfe395e92084b5b431349d46da5
z4adf5d1d57b9087a0aebecaa7b559d846243ec9836f5489fa4e4d304fd392d1b6afe3805c4728e
z4b0eca49c119a30f4017e35de740bdc289a3dcc74a4f982754773bb167ea84930ed763f6556318
zd83d0b477faf73bd888263a807ddb62df4144b25acb821721ec015ef162affa2fdbd9614482708
z4a37a586f9b0d89a7a5297babe67bea31c29087af2197436438617ed2a63f56b2ac6ebb14c5937
zb682899d62673f23071ed92aae4be959b27744e14fbbecb9fa80bf9d32ad22f04125737366617b
zb6b7b693c0439568db055c392854197605ce2ef66cb63e46f0254da1acea10fa976a819bcef3c9
z71219405fbb20d372b6d3f3751bc0a4ceb78143a189f937a6200402e4ac947ba009cb21a7fabeb
zad893ba41c337efcdaeaa51d1a4473d751bf3374087dbaeff4370eea9214709e8f5c0a19df5cc0
zd549b5557e85ca936263eeb1e70a8b52c8d88a4464601798885872804e6b15bab5876ea23cb16b
z6e7ddd131cbd4b3d9b3c3c6005a2a67aeaed7b386be99ca21f425bcb96c3af8df644ff3309367f
z39de99e1d298b2e9456b55ababa87842ac78eb1daeb153554d7464e3e5c3e816e11b0f5577d181
zfba85a2fc232de2dfc7bf9e22324677602bf3a1c2bd72065ab5f90b95463357bda97c726c83a9b
zcb9b6a5304aa9725b3ac88411501a897511f8080443613b5a5172d8b8cab502226291105f247c8
z26a48402e16ce8527d25c85579dbd71f3f6bbc98b32a764de2d30195a4b239012e49324f804282
z8f15414c21b975c1ca89393b84032bac9571a1e704b9d2281ac6076c862d252980d749e133c748
zdcd850a8b9f4e9eb2ad0eb66061c72b62492fc8485ac95ab4ebc7cd60333c33373c3184340a70b
z4ad6953cf00d032ed3533370e7b6a40fd964d47ec93f04f82420dd09f89bd59ebc3221a734ae75
z5fe098ddca9ecf839bdbddc2b1e776b855a1b5675e79069800959abbf92d8dcb319f542d0567d3
z00ee1b4479aa30886a0208cc5a493af936e7ca82c937a4621e8a9633eaf52be4f9af1fb42b91c2
z562f0ec9d0201a11e639c1963e28eb80fb827b5631b090f5b9130a20c391f3a1c2e374a1854e0e
z2a2bc8b5bed72d2332b5e0fee57df715ddb8944f5297e29dc95077ad04445dd3fb2cc9eb2ed092
zb8ba4da692333a1a8a37e1f735a4a556eb4b4e18b14bc8a5493e3c1f5cf0475c7cd9eac58611d8
z6fa22e49b0e3c727d3588ff958810377c640fffce3826c9901100c42080420e5a3e72ab1e70266
z5c89f1041f83f1ae39c0a7dfdba086e498de158d6e141ae4b4a1f64eb0ce7198a26683001ce699
z09dd480823e117c1816a319bc78560ec47861d7176623753e59d05995b99395d2e45d78a3b7bce
z4d3a9d52e5b32799c9908212b3c80aa2b519970c2c0d5b87a25b507288db7b343120a07f9a26c0
z954d6d907abc6429f41e03426d057265cfba560e1f0264128c8df25d9793721c27b16c09fcec67
zffaf767653fa56967586c9893d3dbbb80e4644726011d045b5a322dcde1ad834f1ff1a100283bf
z3af36e40a05d870bcd94ce64e30cf5dbb0ec5e0e21ba2492f1777e40642b47dfa358db49aa6111
z5208cdb37f72d353fd18725277c4ce3a119e94063a9af3b9c159d4a781ffb97451c580c729c4d6
z36ffb2e6644c5d97fb0bb35d161c2942bae3e0e7c4c01a7ae61ea787c5a88f5b959abcf6076293
zaca603bc538c7aeb268ad789b1a483b1aa1e66bcc11cc86cc1c9267e5df8bc98c4044030b417cc
zda2d6781b24f34f31e0571592c227f1a9696c2255c9a3602c730458242e2887083ab8ca31a2c8e
z7f20d7a2e1e8f6efee076e2e5beb4224745c5c7cd3ead574cd70301864de946af4a4918181193f
ze142dc2f6fb8e789184c51aee9dbfac94f80da02bbcf0f0034af21f254112dd2f9c5e3b99b81a0
z516f75686a29b844f4259c6314a99de126f9675d67b9d576a40e67424f87e1a86cb382459cd783
z92b8c04335fd5c6f8d57384245486e0c4175fddd49b97e3a560d0dcde546a0a74dfa322c1b7ca0
zf4a4a26ad0958860a7b38822b8e6e96d3fc2ef7011d5bbf4442b4a5682c75a11e3252e84b36eea
z04278b946d84afbf1f3de023f22b16fd3195c43aa6befb9bae5cd08b44c3a7c14c224a8ae6f469
za387e0ce264055788dd54b0358eba5e0b4340fc353baf5ef0b1884a893fadf56671009a5bee8f3
z883ce0e2bc7496b887729e26c8f1d7dff0a61de6d82747a7970b7c63075c04579d6c1339c6b957
zd12f8063e59302c0a86b26cdd9459bea0d3f18fdac9ae9010f3f2b27590fae25a1f83bbfcbc925
z9849e742ec770d2abb9ab0c2a6b1a5123522f74b3a4397da480e443f3ce603e882bacb6cfbd641
zc598ee11d17b84744c326bcd964a9358efa037e2cea0de071b6e6ac7ea3109cff86fe689a7f114
z46d6d95b493a7c49a77a2ff248da20baf1db5b60502e84c6f07d50abbc7e2a4d20a8d1d4a1a55d
z1109c1f07b32f18a2b34138173c1547db9e88c144f46a0977290f607a72d910fe3b87ddbcc29cf
zfe34ddc1720d09d236378d02423ce3366affbd94497cd5982715125dd32bbf207a5d868eb59cd1
z399ff9225b5b9961583dd69b6fe97de4dfe10cfc490bf88c958fe2a905cdecbff07a248ee19e06
z10ed047069594bc28cb9d8fb24eaed5126e27effe5431c7c0347ec1dd30e7804f854c92da12d36
zd000ad142e791d76574ec2c2091506c49bb2d51751964ce8fe0df2439b01dd8f92203e75a61d53
z7cd5167cf07626a7f8e5c922070619c69dffe407a3235bfec9d76c3c6f47bf2190db36b5b6a426
z326034f4390c1e95c74ec82914cf100adb61a3ef38d76b0dde37942a1ba53a66d129cc38ebd1ca
z5a1ffb3882f1b18f02d22db8e96ebe778dacd2f69b5f2f5f1eb59e23656e56def93caf20ce8291
zb9a9a049fc74ea9d3e7f9a0e9750129373670aae0b3194bbc31205d977fc40f646d48c4e2efa89
z5997b9d051acbc4e163808ceb3db72559a846479277a5d4a419933349e105c2ca1d3f93b7c2f5d
z25662b1d2f3a8ec01edb0971f31f006ed0538986ebdf7f4a6cdcbef4e3700d85fa2c932febad16
z0158dca01cfd1b386924bcbf3f39cb6950893a25b9d533be3816b637fe6d0a673123723ca93fe5
z9848016d06beaef7120209a54721a0deadcd15e9f15f68d17d3d95ed7e9f0bb8284c40cd60a586
z838fca88f8e4145d8fa2c07a8aec0e3ebbec1074c9532b5fdd989f3ed4e477160edadeaacd342e
zfca018dcd5de5447c0e5768571af9bbabc5f38eebff2cbe2c90a4f4d17a01deaf5c0f707862cf9
z255d92e31a79715d987c2de6eb12b0a105bde72dfd3a0844ba8b387e2ff69f6a4bd52e48192a87
z9ff985b81948683ba0aca940ef5c3dd121e2d287e9c9ba79559737ff78a9f45b162f49af253386
z1d3609d17541c7343384d46e4d6277706a43173dd6afef1943e827f4554cf407a0eff9b78d5b6a
z528b16d00cabe1235506745d2b678f9bbd1aaa10f6cbef034d21fb3a2a91b149c7f394bdbbbe88
zee29b8b4368e3d1eb3b42960047cb16ed5da3b6618c34ba21da06ac2f48fe2892a1f735f71204d
z017e8637ba5a3be69d2b41d962fbe135fe8fb142eb4e99cdcd4dfb32a16c8be8e6dcc91e4fee99
zcf8f153af4e60d122c48c2b232ed3e7cc5d5ecfe4c78250f1bddddefbe9dceff473394f398ff30
zc43899ee229535b6672308d47b51d9e1cc1162db9624ad8cfa4fe8d106a40475da49cabedae599
zaff5c66ceec915b3392fef4f2d4632bca601d8c7212d580ef76a8d5c839f503c5c7cc347076df5
z591c1b5560e1deb3b2961310ffb809f8a4f37dc46bcb9ab233544a9b114df9c005463c59ae889e
z7b113b31293850a632f877a0fbf42fba789de83dc7d89a2ab3b87b0c0c95f78f57925e1c8beaab
zf4ea4985423a2b2adae4fa0b1629fc59247402a590bea2edf1e5f6039bf8aa84afc970fa1ef784
z5ea4b09b3db84252c3c7c4e2f36fa6a5c5f6d679d1b6980436bb5c925c284f9f4e9b129f365a8c
zdb1c6239276c00d91b2b00b6d2ca72cb95549fc0159b3737216fe4cb025cbc79676d9e0726a94e
ze9fc1aeacc395c0d608a5f0dc17e804cab209e0d2e866d5ba0e16060fd3cc26746f377bdde0d69
z41997703c72a432c6350da4ca87855bc9929d1d02c97a471046c23ed9c741db1e052c4839e7a1a
ze2e208b12b04adda220f5cb3976ee8d251a4910b7a9b5a8e6c055202f3ba26b3da9182a4639719
z7702d72dc29c54917631cbf85299fee319066c321419161068693f115adba9888263c43dd585c7
zf9753ca57cc4219b9f2aa5982dc502d580063dfac6a7b61f678b0ea3e26f0a58e0441d52abe061
z0a36ad7d33c7b5665b8f5e24a961cff4524c41ca1a65b254010ed5b01117692d3c80472dac59a1
zf8562190c9617690ca9fb5b026c64d079b838513838a3eac30cabcac37fd52537273446c8f9022
zf3e3ad387b73fb0a04992430d60b5996fc1eacbb67af6c144438025fe7379e66bc0fdac9c22005
z8e35a7586c54b1f8ac8394410171b3fc82d24650346b1c3dcdc4b13c2ab5df0879da211b9345be
z9bf2762ac2abd56295f3e98c4db1e2a270a6c732e9d4112542a31397fb2ff4f479e928c5129e01
zfea07a28db1297ff307095d08152316b1d83e82db6fbce663b6bdf327746abc561b081ac01c07a
zbe52d56366d17c6be3f8625c330c94e5d5021d97906dde60184bac2f748fab19a519f6e1d3ad64
z4d70f45c1a5a8744ab63047b4bf1251a8ff2b626c45905a1b154f01adf074f87cb8eff2e9befe6
zbaf02d1e399411ed91a8f7475d6b911fe649b8224860efa64c1b8fe7dc3757ae0c1fda9786c109
z6ecdc8146619c330af489e421de7f173c8a6c13a2e51076569585e26263450b6bb9c97baaf9d31
z46e8d00e884fe0e71e39991806ed9415d0de7ca9ed7f8401a573518696c84f49c05680b9864651
zf210586029c831fbb517e662e097be12e86c2533d1b1fac8e9a4d54e0862e7663f1da35cd2d7dc
z17795b2150d91324545bd4feeff81a8960aa1ac416ee0d36629c64bd4a4216c8cd6448320cf11e
za27848174e0d7be9390b5fdc3577d8380f6073a0f19f284f50a54dc1cbb8b3c3688f7e5d444726
zab1fe827dc771cc741933f5243f85c34ccc4dec66eb5f141c357547f8c6e6fac3952a185d34d61
za20a665925fd24b93e6536a06bf44f7674efff5b8402eb9a4c38a90be2f9cf6ee5a7ebf77dcd40
z57a8ce72eb3bcec2f30d8dba75900c7e811616a836ce322a135f52c148c1fa04c79b16427e364e
z9b83a6b3c9f985df8e64ab85cc1497b86eba4fa04f5b1b9b42fed823e4f825c37e9a11a9101ae7
ze578574bb3c9fffe3d70b000f60b2209104d65a9b0ed37b29c774e78cb992a9496d173a68214ff
z7cc2b44a19f7e531c854737cff72bb02401aec33aebc99ad1ea7d32b43477df0348e302b28773e
z03130c6dfd6d1736fad75411f8e77f7726204d91d374d41db569c38971ee32d50a5826939d5b2f
z0a1cddf9ed1dc081913b54699899bb1f9593dbb3f164df5fba06acdabc9e999c029bbd3771a8ed
z17c69872057f58faa6c7c3012456426ee24e5068b5bd59d046823017530da55fc171de3e0fcb0e
z6d1f596b410c1f04845e243ef234a6a77f354e61c198ac15d6718768fd7926a62e19f24575f79c
zfba541c40b0e303eb2f99a8a1de2e930312e132abc257d21a7fff13dacf8e423f865324a10d04d
z187c985040c20b1bc25db818c6d751626e08ec03987e29b0ba1980b34d68abb375759107122dff
z56de03bec781bd71536d1fdc425b777063dd46a923b837314b5db42fd0e2cbdf3ea6ab17606b7d
z701f79db2cef2de6792865191be1ca648b92522cbb5bd94b55ded28021087e2911b56e628bb7e2
z9302dafbd96dab79689feac0b51f5d6a392be8982bd5e2ed1d62f4dc13a40aa28ae772feee6517
z2701f093bcf3887bebf66d5c3b536edfa39dbac9e96689d1143ba347dcbc69f087173a4e1aff54
z66b2f691896179975d4319407d57c2658a7896d76b30d7f08a64eb0b38f374c1995f422fa3942f
z793533788b051766e10d90726356e6a0bb440170468212b086987e6881620ec7c04a737e9b6075
z44195b4b9ef193afe5b7479de59a038c8299375c12b90736b5849ad717864fffe677dff8ab99c7
z3e37fc37902ecd8ede2710d0215ddc95b5105f64fd50ed876935a488f2c015b8e80d90348478e4
z093e9c53f4a3d7e87340fc883cc0db4a84b238ea687c7da8d2e85ae876a1ea9e76bf30df78d5e5
z25e75cd65ac6afdc9188238e02a84f77c3d93c77ac1ed0e0366028d06961fb0c59d95354c1f9d7
z467524ae90421696a2eaf9cecda3ef5ac10b87f6d2358fe02baa0c93262978141f12cbe02222f9
z16dc96ec4edcd9053e02c5133cbee2bbdb607dd6a03c274f406926a0e182ab5cee773ce648d393
ze64f3796077bc5261fead0324641af77cc3d2b8bbf4095a0eeaabaefee2234d9882a4c10ba2370
z109c0d1a372dc944e97671362d882b37d2568f1aca53621da11c7581ee831a1a85b6eb54077e58
z804e5967d58240060cf4ae76d8dd2bb40858b7353a974b362462b354c148836fef75b22d54a44d
z6229aa17e588d36f0dcad002426ddd4dca1eaeb502186aca100bd072c6cc813219b61f7ff24365
z21d0fe0f603c7f988af0a6ec2897bded46730d2429b9756c483918ae7302bf6afb23e144518dfb
za348b153a3f0b02273e1545be86cf8ec552411321457fbebcb018a68f6246d5f2e61690592c6d1
zc1eb253177aba2542c0c385325708777e6837d7d46f1875daa6026240a4fe495cfe11d7b3acf59
zb91d183b1f1a6b116f79c1a60afa3d7c218f7b6fa4c77e6ea30626604cbaadf93ac4737d01fc42
za24ff1a36f58d2230fbab54e08f7ac30306b2ffb296130c93f8012c442a62660835cc1ada5510c
z5d313e1104d43cdf37e49a4d7041f115c10fe61f6965274c754d85c99740cca8a59348e5c41731
ze27afc45491f900758a560189d87015bc8d01b3c58e018f4e495743b514293f53a20a0f5071d34
zfe8fabf3824bb894afda17ee898d88893f75f2445bda6b45dd0ec92e3b3ca39545a4cafab350cc
z7933cd963413bc24ab82e608f02b84016053740256a6d5a88a6aff22b7bb457ab6036cf3be744a
z07e223f18f4cc291224b1e9bfdaab12c07a76631122d2af3e354370d24cbe002c0d64c3f6e6629
zb210c00f04387d9bb405c3113b32484789c5582be85875ac147ef6de41cca44bdf7228a6adadec
za7db821463e391946c3a6d05a5ebc25377b47f204285a2b29619f1129ae9740902321eca11f9ff
zc18c17e3b26183ff169fadab2ec5bccc0fd9229c4616d951a401eb5847662a4e35e0ff539bde9c
z696400a2cb7ef151f6d30c5ffe43175f7f6cd0ef32606b63461fab24492e3131af9f67630fa8d4
z114aabe6d29bdb74c8a01eb6db7980700779259426e9f71895f77a57e85b9784d58615c3f80727
z10ad67a1bd40afe406b6fbc4f991c87d285dc5937f9ad7a661f1b6fda7d0151afcd1dc2d014192
zf2128d80502e8132d7567415aa1abd456d25d7e58a6791385c06828cac74182d2e6261a85e9011
z9b3f8482e7048dd223b81e4e01d73732c2fa4e392762a9dd610422763fb252b35585cdfd8dfc23
z5011e3e91573ad7542874317e67ae3ed08376893f41f8732c42ee0087b259019314a8a7307a7c9
zd6112132b31c809932b046d6b7b17b8856b5c75037aa87433ae8da98ba16ded7b5a58da2aad232
zbe3109648f78f3b89f910753724f77ffbe102e0b5b97e854b9b230323690e3de77546ea170a77d
z61e5672b13a1ba07619682f97f787f41b44266e183ed2d8c2b72199808cfdf551a6f6ec5bf30f4
z0ad9d54fd39285376fa0229b951e8c8cb4855b0a6cd116978f4a138851426514d5cdbfcad41990
zfe2f6e11a19c4820b6d72830401a2ca3893b9188fbee7b0d0b8189662f90be9d6c385c131d7012
zefc75ea1816829f2ffbf2645c64c5b13d0e53a95d6abe4478e4ead377046ea9686ac18e259b462
z1321d4d841c902de2bd02b0547273caa4cb34ff103985584d4ca0eaf4307f27fd7316257b3b7d8
z258198b6e7621f3dba1e7d4882ebb1a9add706c322d05ce014bb2e5a058e416e46a7491cec902a
z255d9e645763c81fe69d8e308f03820027289f396be635b8ff1eab92317e973a6adee3bbb7d4b9
zf542802b3ba279eb7428a5f7cc484884a86409fbe52362a3241e6f98d7f5c591c459631aaff50e
z7d71f4689c8c9f936733b8400417a9065b5e0515355df9f8c216156bc1e90fd50df86e00667b52
zae5f86158e5685474f760917daad0311010d00911ba4a9d9ab5fc791887c45aa920be8104c12e3
zb157410e9ce3fbdddb58899c92345db813cb7e2f217f12beca0dd65b6f25ba5e5057355a36fd22
z82156c4fd1f7cf6fc10d374e2d9dd500199d06c69a1bcccf292f5587c8b664e83e9cb7c18ac1e5
z38a5f9289806324cc16f93d4ceef8cf449a84df9539484cee5f678687a852d63d9a79330aa7afa
zb8e90157b0bb188929de806769462a1ff1d5c19855a7a132a0590980b12852002406b7668524c1
z045cb804a788e069059e54a4e661362bea25223495903d6c7172594bc82740a4572e7c5bf79041
z7eff2df75ef9d5a1dd2d2e3f0808f9e4f1593ee8024d053778104ed80a29b476ff3bdc4591bb94
z6af6498e1a01531f5661eba4a84c66aa4875b57f0b0d2cf364d8499954396441021d4207a6fde4
z0284ede118f0af1f42039c14fbbf1df4e3c8fa046fac5b983d894d2cd63e0b04686de37aecaa1e
z5bce9c6eeca54fd8f1e7a5daa9f443ce7803936f3e794e159498e324902acd0cd9a796b7dcb582
zad1dcdd529b1410b5b59e4c87daee9527a41958db2d25806c32ff959cf129e8ad504412f13b436
z62c707e661a44854a39566b639561d05421a92657950535b40a2e173a6a0442383561ddb302c4e
z07498da3844118ad44e9385905ffccb93cccbd057c2cc9198b2093ac058d1d899842e6cfb5a929
zbe719f77a5c6fda2ef615160bf3ef08ec864f4688ea791b4b0c87d23a8e3180304d732fadba8bb
z0b058f550b0fac1bc7d95cbb1481a7998bb7c5ce77cdbbc2bf7ce5616e1a29effcac36a2e2e656
z812d10819c4f5bfd768e014fd20f1e9213e1b251fea8086d210ea8a71fe95ca7de491026cc7cc7
ze89e260b9dc3742fbccb03e0a56ceb97e37346be2a426361211c39d7f2dc9b0dc0cfd26934caa8
z6c8561c0c787ed1f2961915c869134b122b30efb4656d40ad9ba3b446e3b720eeb33f6bb1eafe7
z76f2bcc2fbac8380663b50f32eef4cf2ff90d422880786163eb96d50b3d02d986955bf8fdbe9d5
z99ec388ab3da38873c6941b36d17a03ce241a896959e0b27054ecab710ec817e3c6a8a3266030d
z0d97db608b35d9b397996fa85165f71e108206fca5ec6c0ce13ee5be4c228a09d1781ceaa273be
z21e600650ed98b5d84d5a7f2d659ef96bfddfc9abf0299345103ddd1d4a248191b13a36517f61c
zcac179d9339fbf883193c139f97288c741c9b40b44db8c6cd4f9b10b24faf5a5b250831a8ad695
zefee5b9a9caf3441d760afba263a68cf149f939635a4c110f98e7218ed0b7d8e2c9bd264110e1d
z6cf24bf0e36912e6e9e558ec28dd2bcff52ee95e4e2672e3e7e367eb5c34453cfc2337848150a7
z416a7a6e8d59509ddc949e61743505108ef327d5cddfec207aa918e12bead57d3bb577c4f9ed94
z68e321e77ed801f81c1d71255446cc1a19b30d5b4660501f272974d0a2b315b765b358c13f7554
ze109369e4122af5c829be536821f3ba8fa5e09e179a2e5ea723219caa756f62fd5986468a0d1a5
zff1f00deda1b14934fcf944e625124757829794cd79af5bc4390cc95cf14ec0269b90bd4b011ea
zbe0c4e3b6001c22253ef5680c8a63a24a009cc6333f3bb28e02366247ec81d4a9cff9b917fca97
z683f4b057b3210b780b110f0bf84624a3aeb482c709b87471a8f1fc8886462f67c85ebe2ae4f9c
zb13787b54514a482ad6641707fede12f79f3dc3216f648c619ef317c6af21b1284b770c37fec86
zeb8007c397cffd6b0028653a7276ff09d460abcf44524d39305466dba16854c491d2977bc8ab1d
z0ee72cdba356b0c2a07160e86b0b9f611d6d019fde298938de4f37408be380c86022beebdfb0e4
z1a9de00db0b7c059d8131d1ceaa1ac3f57fdc335c84d923666f54a65885f3b9f0dfcd92c391bc2
z5d77b49cfa8567252b6cd5e5e2bf3435782dbe44b51a4cc6e3bbe40c15d380714a2889efb8f8c7
zd26fd80b304ac525dd7855b6ac5f44b44d9f04f72faab45e5491cc5873b7d4022f7529ab65cd84
z8e0f2fd3af2177279cd1c4255edb3f553e4f3e1b23a166df3021e3a6f868407103a982337c1cad
z9110d79ee59ee7916111d969b5161600d850d0b321678162c5442194e5cb7c3492e647e7962fdf
z2f34a9dce4ec2443dfcea50372732b44a79ba69afd81a9992c9af80347aa6a733c02391aa6cdbb
z61c3ea584f25a75a95f3255a6156ae1a7df9da0871619e983754d55430d8fd02ad258e7408eafa
z09b3658d5b97c12f94f8daf2cc52c72c14512a5b889159f0f4428145492523858d7b1b62c7a328
zcb86dc94516bc737b31105a03c03d1ab182febe6df818171695fb601b77f62814f1f101edc05d4
z99d1ff33cd27a951ed8f0767f06e1350565c5e1139b96554086c780018de6641a2bae906020080
z4b3ecf31dade0300d70489d4b18ed948d23c3bd51b241c223520217de4150a51bda2d6d9175f95
z87c45b684790d41a63e9051d8a49b26e9d45d5cadee459e77d6da8e94622d3f8c22a4c1bdc5795
zd416da849cadf415b0cc6f9d0620934e577c89f90d9de44eabefefbd789c5bb4c7e771d7a19fe0
z17a47d0c60c3c7605b0b6f332ef612a399373f0822c93c6172d92ba60a30d958471c2e0c840b44
z230f95e001301e32bc816a04700ebe350cd51fb47d9723ff68a2a6f06d76648337199033392afe
z30b9b0fd5fbc4981653874ef2bc858b10ec52902dab7808c92a922a86875b75c244a5069578340
z68126b6a763f5c726059ffdae73b8f107d869824e285039003ddd4517512d1ff43947d2393a5ec
zc63ac4ea4c3c716006bde21a6ecfff0156fe01f0b92c622fd9d3d7e432ad83580548fc5d3623fd
za12836e269ad08a35cfeb009a65e233ea66a4a3e8c0d2a5bfa81d9c10b57750e9eec02ad36d71c
z46c2f577c4eab115d46f70adf104a74f706944f1da41a74c109e07bdfb6226da78f80675e7a968
zd9b885a9b86f2c08b52614b431475f1994e22d936dc856e6899c6f4d7fa8f254292113f205c6ff
z302b26ce03521f36e6b2ffb010527186e9c998e49c63eb74f2fa5073759abc5935676386b5baca
zff17a777264db3f6e44be8239c28865dec52bc5efd6c8c875adc6308f921ca5e51274312977747
zdd011dec970c761fbba034b390673a7003ba40ce9eb0ca1bf6a09514771c451bcabca1fac35ede
z6917e824e0ad9b36d597f791d404857dfaa1a3bdddd9f20e9249bd829d7ca8ffb3806502e928d5
zde46f4c9185ba17088c9fa9f5942c6d58aa61f0342cb4199ac2c63d89a0df7be62f772f55f3f54
zd22c04cf6379d98f25e41289e84afdb8ca1399048418b20562ffef2ac7972d3bc7da5d4d08fd83
zc04a428641bb4a2f578d5ccbf53862e9e7e82bcf1eeb54ccc863f4f9cbc17dbfabf4f01dd69cb7
z118adf509a01f55b2512e34e58d8f80665e35655e20d0c95f67932e9d1d46132c1b60234ff6cda
z8dc3ffa5eee4b1059ddc4dfc1510cec04b36e74446560856a077c35329047878672970bcf9bfab
zd1dd4ef93f277a869b3b5db9e2b0e6a48528bc6beb273260ee6b48877bba84a14170376a131400
zd2d5d3f496131a337a8ba58bddfaf6ac98e3efa3a74a3055eef7eb855cedb88b8e73faf9baaffc
z0057e2ca5366f3161b9b9ac365e795b6b098cab9d39d0c11c85690c076d92c238668dc6b1c50e9
z2310ebfca6ca057535c6bcc50548f237e0b0ea018492a1cd4e8cb9c4d6a3ab7cd481efa35bcc9d
z5d96277f05c0d834db9b453046c02cb3b5bc9604208f311c0e8dfd60919f9b63f02851f1e16f43
z24b8a5c90d12a062f1c5587b2be72cf7d498375b41e9639df6183dd7995e406811e7b0cbdef689
z0093d2ac4c3148a354c01b244cccb59fd28b6122d3ce57bd78c60315fb64a608b87fc8f7a43bdf
z3f3a4ded355b7b53e7f52c1ff806b0b7fa8e7d3ad392becc01fc6eaf635b12b56d2d943818e68c
zdf135585ec4ba46f1589fd1f1daaf546e3fa330761816e24a52f93d48fe7e814d1aa7263a72730
z8c55fdc7b929888ecde52fe59607702affb077050de4e7805f79c3b3f08681e7c76d5c1c6ecc09
ze0ca68c87ea8fb9fbd965b2f7b04bd248466e45066436ef49e67123d63c3ed1d60bb5ca38fb609
z1bf586c7728e4b2df2f641601713129e65b6b42396f5d9770b5ad2703baaef1c512c78449ff463
zf175228951b09cacabb365c087314e3977d32fc676790440d0f587ab0b51f904d54e6812eacf69
zb636ffe8cea1da69b1068f66b5dfcbb41d088cc1091ece11aec365cadc2925c5e2556d0a62c359
z92de36ff67f71740ebb83000e4bb7318cae4164651761b27070ee7eef28ce9fbbe02a66bed1aae
z6eea8f2b87b4376de22ea22070035bb0eed18751088d19a286720249430f4f1faab900155ee2da
z35876d435194432f48c6598ac59eb5761e232edaef5b90c61497dde14e1e010cf396dfff6841b0
zd1dc3e80060da0cf32c1dd9c16f5c562c83bdba9de72dfc05d60ed0f475fdc5392f965ebe7387b
z2fd29bf6adaa6a6b801cf854ec8b575700d31be71c08772a258546045b041a2aa74d127ea14fac
z290be4b2fc98897c57736969af8efae2e01c1325e8fb813eddd5fb071e32cb5f147f8ebace4589
z87d0bd18ef67b4273f8c5a2c5eaab2867c515a2a145df1f15893bb87327c430789945561b40258
zfd57d7cad61c1910948f9feb2b9e9f91a3d2b5520aad93807de1cd1c1ff4db5d25499d6b882866
z8c0cf1b31ef9596f0f021ed85704af4da300466cbd1a42a956e28a56201e60342f40ec656aaa2a
zec42bc0cc4b5e5ed79850deddffca5c15302766feb47d6fd5e577121d0308a2e4cd26fa114b15f
zc2dc0372c602b135971415fda3be584e1b9f106d8329a7c4e385820542753f0fd74e46eb74665b
z87a12836ce62febb2334a02574391ed28b1e700e8cb34509a4f5bff3c112817487c9bcfe5b1b67
z6e1d88cddfae9f8382d7c633030eec4728c6e66da2b8e3995f67109e04b20efc0b54c308360d81
z2ebd8e5aa64b3ce18a36adf8ee701e9f48297cb805d5ec798145cd660f6f568c569b4c3a344779
z861e5f932430e8d8fec852fcdd8a879c854ca1d0e98025bddb61ced78f67647cfc1befc867d535
z42e0de1484f10f59136dd91f606440c8a72237f5a467549a6e7e5cd2e77a4fdf47fa276c3e151b
z2828b0efa69ed3320d0cf95f3abcd59de215b1d8dea514a55833fa964b0fe59b640e118b77bba1
z51ac68caaa58a752bab887e486c2beeb6537734059d11f80c5b05ea1e43f702b3846ebb5d1aec1
zece5a44c91299050d07306c6f4ee9e1b3ee126fddf3ba3982979b38077a7fe4f5291fd76f1b0e3
zd61491977883f5cc2b01c519892b0900cb9c21e27b867a89595b97e44fffb0bc355603217fe87d
z8be6873a75125bea631ba205f85af35e5e5b9cc825683634a0c521067398a6eec96682904e73c5
z295697390f9417841971b3965a99bf31096f1f4607db942124ed11e1849b1132c0b93a6ffb2a15
z2419751bc7e517f668ad5d64c93df3aa960867c69ca18958eb902c3d8e74defccf50ce67f33e45
z35ee8d72f4c1bff38255c9f1392e823b17361d9c6f6fcba97253d59780bf9134213ac604e81b25
zbbed56e9cda56cfe73ea882e6bb9ba94ef0ce5a9e5b8793087c28eb9611e7e7c2ab32e3b77d52e
z41386c1494110016f56f9e5750413214bd154764d6ab77ff3e06edcb9f331d21cf29a39588a46a
zdbe5d4d15ddd585e015ab63496964605f25cc9b7e596e5394a907bd8233cddd57c167f71d9b586
z8d6b28bd92005c3f990d49fcea77cc4cb0c2bf4e35ebe46fe9d9f60fec753b7f7215fc133ff27d
z56c487e236f7894b08a4f12aada9ba2a67d3b8e5e43496ffb6af3da4befcfd5f987245affa8ea8
zfd8075a8e68c0ba0a179e7240d3d5dce5000cd19b3fd2b3259e94235d7b2a770773c46e74bb785
z42810c6fcb5003af8d6883921a6498db1eade42b450299a4342153ccee56c426e26dc462e8d3b4
z60d7047380d4f6e7d86d8e2530fa771b41c22ef84f9006199f3ce9b6e55e661982044678a8d3c8
z9931d04c2a0111ea6406d7d543d71aa045636f0500b4689259fe706eca7adfa4b4110927fd7abc
z208dabae44cddc4c6499b7920f21cb96c95013ffd6e6ab1b1f0d01b32306c871bb1ccbfde7d6c4
zd0fbc5b534b8a98677d2c9f35bf4d627fd79b60417761ebb0030afe0366faa33c25180250647e1
z3a42afd870af4caf3a21ef12b2e5988f719bfecb358b0fbf24a15fb7f9e6ecc6af9767dfdc1dec
z424c29508d1004729b9b74f0ab5e0b1ef1ffecded2e9ede20e1db92ac7e29521bf0dece3604733
zaf650e4d72803c7dcaf65c722b852cd5d672cbeb8d61b6ecd28b151c81716b16e46acc35d338c6
z6f83a1c5a0badea0395a712727f6eea8f1e823c9a5ab11150719b342f28421fecb22c44e503563
zff08a43646f2bc6274f1e2671bba84a235c9de3651114c937e3b0a2ec6456f1d63c9fc294e9de6
z536e37b35d5db706f8f51613d1898a1c5e60639e80e4ab14c5003f4813c90b3dcb4b88b5c13458
za2f51a675c42f1227686cee01971b9ad256754def2056105ce0362fe42d5b4afc4eba3359c3fd1
za3c8c6557fc3fbdba8c237d54048052109835fc6b782ae8e98b41a54f30121817e8c64af1b466b
ze6b5ee1538a0018a50f6f26afb502dc22811da6ff66d58535983276393efb82888f60c0a83530a
zb41b3c336d5c98cc426acdfef7310e8f2b4932f6ea170a017b90dc3aa62d556dfd924399ca7af7
z42c8e56ccbea0a3e147893f297dbb6e34e7809e207367573d984766a37acefeda44394257d6b41
zdc30a2811ef7f68cfe12d203d4dd10375444cae14e5a8f256d44f34e7f13466247338206fdc423
zd93b60511f91eacff9739b95b836b96e26b4b4c82ba4af2dc560323b73ea2284f301ef2732f07e
z0447ffe24d93e25b93bf34ea74b0f37ff7f27348081884dcd0ed513ff3a080836015907d37fd5e
z6f0336daa400e879f636278392aec54f7b1ffb334327a3267723ec054e8e92a5fc133ac7397d9c
zafa5ff42cb71dbf4f22b2fdadac9129fa3895ae9a74801349dbd8e018c4622b2bbf84c6b5fb2ae
z3b1334733ce2f45a6c3662a3a3c1eeb6d1e3e026407330effb7e09d850bca5a54bd61bc231506c
ze4ceac84d9b4c11e87db8f50fbe6f8080777098f8bd1a53b4bb02ea489fec152b3911eb7fcbc70
z8481a309975218ea0ce5b8c42b469c9b39afb65b4533319f60e0cbb00b46f69f072106428789f8
z443ae440df16fe9c282c093963ea832c789e8e7961b791246b8c3d0457a22cd77f1769f2395887
z6c0c1c4bbae61bd2d89c408acc76a63a8163d4ac2a813074922ef07ed80f94b089c64d241a9fb6
z3ea0fd093cf99725e7704e9154c5043ca89cd78c798a760ada70d4a066e56f0b18044e6f6e7f42
z74e44a4a09cf6a5a6d440d2cd06f097cbf743a6688d1b2ba2e06c90ab9619f20dbf6c5f6161c00
z4c404189853eca3b6638d635fb9da825359b9b24b991b17209d41059616bd6f5fddec163be6edd
z57c719acbced2c70848db5fa687e9094905e881942711d4dd2586d1bcbce391aa931c78648f461
zed7498fa0ae899e9bea1c14741b85f72848ce1aee042321e3e61618abfd2fccf38d8074d691e0a
zd7a6b994587fe70a330b3de92b08adc68b1bdd664627b5283ffc5fe7031f1597bacacb8c38d6fd
z78f2124672c9d0fd365ce12151514eb16e1561a38fedad8ffc23d8c57d68b08bf2d078d48c4d92
z59c1ee8e9f5c9390078319b944d78f0aa41aa7f9d8a7bddefd969f68a9e7c35d7f7e71014f3599
z75a9b11de42aca9956db77845e54c490f4c6fc1bd8b0e0babc8aeac103fbda109c097f1c359d89
z66811ecd2c81584690f31ccac416e7af903b4c31183cf0e8bff051be8a6394c038382b390eca38
z9adaac4f034f0bd2dee772797797f276f89bfc664147cc3546ab851fd0d106b4155c3f0f362c6f
z191a122f1c91f1c275dcae5a4997fb963147d6033474ea2f06de564f515c9ace7b6c71c6ed967d
ze84e1958dc3066fd3b077a81ace9c12bfb96959f05dcc948353f92898aaad92aec172d79533012
z8f53afdade71e96b228d1b46e6f18b55da41e172fc04a0b8f82566095f0af45502d70c8a70bb56
zb37298eae0308f37f6c2e1f42643551be23b9681ecb4f4a8b4d974cbfe8074bea19b9793ac730b
z04c65390618f5e20618d997fbe718390d530a6577ae1e6a3160c821850dcb5dec13299abf7552f
za551f1c6d6e3d708e0769ffa116a93ccc78801fb83faded8625bd12d72242c386fc9417fa7c010
ze3d79254a0890b597136bffe45684015653377e40a1beb1dd86a35dbc82b8ec8de7e967e6a6c0d
z4937e420b660620b10aa742a7c3b94a6a0c774080244b2bc550b3df1257f31d23cb2d7706550dc
z709271b5fa6e48d990479d6d74ba4c2eb71fcd8c04c1dcf8677419aeea90bf000e5931933f11fc
z3059d40917f314f67a4ec0b42df2d75114f0f0a5309c33ee46bf93e50fef5b8ec731fef496e970
z8e66e439d6f4e799ad248390914e8d2f00336b932c07a7641cdacd827adb2adaa5f9bdbe73cc0e
z0ade8bd76d9dc1671411da9c52ab2f67054a937aadaf1c1956ac5575b4a2e63e9b4d93e9a5807c
z3a9fa6b4f98fe47fe334460c6514025bbcec4a13b9f8181c5785dab6d70857b2f8b696a06c7fe2
z8a4a99bdf59ce6e67e39034ae3f04e2bdd1c49be7280368883dba5373075d67177653ccd0d378e
zf4a4a213597e40426a95ca6e91e31cd1f0e390ed04d78e9cb2cca5ada85a08890688e6f7ce50b9
z7bfd17d056ccf02903a2b09595b452fe1acba6797e5728138d1909531901aa61168a7a81a50e61
z03b7dd1d12d15d352a977aa9ee7d5cb3c2f16a607161bfc65e5f33a946ba64707256b96ec6afe9
z2c0365910ed9675882d79c8e4be655431806143159c61ffb24b3194ae83f1205355c72b9381a86
zc36fd6061c08210cc3b2cbcb73aaabad0ae4963fddf2afe7c6b65a2f3774344eb8a12704d43c4f
z6f1a228d2001e58ed5bd8eea5d7a0131f8c1e4c65adefb77985ed146f4695435202f5da67301b8
zc049fdf78cdde0d93a49ff2cb950eeb21a0189e6d8bdc89ebd825eae52c227769cf37105854774
z9919c7082639ebfe1e49ce01aa7654ccff13f919b2e3943fd1c80c809ec65c8bc952649dc0573b
z105739ba89fc69e4cfed6e41370c2b991bbe1043e173b4e5b1ef10fd4a41adb52fd2074862cca5
zf16a48c8f5a41e33eb3b828c6c8baec30e631c23fb365f18aefa13819ac7631f069508a9dc3d92
z1892aa494b1147cc23f822da10cc1f34a34e0b99543120f02ef4e76fcc588997e166a475fb8caf
zad38367f94ccf7b7fa5e2572636d13cd035c41476f78e016c5bb8433080a955fa765424423bf95
za53ce568cd2f549f2c68cbb3b33f1594c25ce898566b3951baaf8aacb1f2e6b31b781e8272b2c8
z59cdd2494933d499deb078904debc8fc6e26354a3bc554207ef53a35957315c40ac4af3337742b
z8777c63d2c32f6d460d44bee6ab2184cd0d4c0ab181c460f7e5ffb700e2737cbede1bf326d748b
z3793a4e70f53940b582e111019b0371bfbae0f8186f73418669014b6997aad5a727cd4ad0626c9
zcd673c765200bc27859d11161ceb201a0eb7c4ebe3e8bebf6cee38b5083950a4d40b6fc48dbc51
z14e8d90c80c55895c0846d4e55c01dd8b2e27161b3efcf2915fce12ea7dbce1d6d3b3984d995ae
z172172dc48cf4cbe966daf552ba846a709d998d002392e1b20d5139fc60cf96f18f648abca651c
zc8a90aa44d51359673000ee2f6771a3b12f36c3606b9b609bca07483649b2c10231eda76d255e8
ze33350ca0982d4bac67f9a3f59d749d21c001bc80aa14c869a300eeaccfe6a2468fd3cb68125c8
zfbd29fd5576cb0484bb92bea500ba2b5c6d7bcc5bfcfacdccfe463478bffadaff9ed5efb6bf39b
z11ab38dda04faf56919521c5888a01b7fa5db903e46a249a75395a43202f4ffab19efc034d96df
z34d7fcef8458c5d4f4110c3047496024d227807e38154bda85c180c6b22da17413887706d85471
zca781bba398a85b5d85297bd114d9fbfa33b4bb526e55bdf0019cec0d58a2302479d0c34005998
z673f74c82486d60477282044c5cae7f6e0e3986fca2204d6ca5a8e92fec7fd6eb6760bd44fea2a
zff498ffd1b53365ca934d9e1ff4af04194026c92a8a83f1d84acc68d2755de41422c1068540e2e
zda86b18579ab9cf9e35204321ae456e57dc1616ad30e82e188295704e88d1a0c8545c05c47e0a6
z9fcccbede1ac4af8f12581a9312d3e6194828b01d64ff319b8620b687d6488a8d212c711d23a6e
z054bd9313a8c831416b0f905c264ffa9c5159ee10ce7d9e4382924367145ae5d750f99e549506b
zb9d199f15006b6cd1ba104c146bbd31bd7f596ee16b86fbaec3fd1cc80334a70b87c63747ef207
z0cdfe478144620f148e0b773899d4b59d3f3e6a201740f5349c21f8fa79288d3f48e59056d619f
zd10f6e3dfe488c18ec4f30cf31012cebb2b7bba3ddeef3551d58b23317b44b0f5ab2d3c3b3a432
z99310208c63cff43d4879d910f4d772dd7bd6e08c8d21592e84b9dda1bd365cf3d1451870bc589
z5a2fa4201f7e09e35440928ef3240ebb4875d9898f9f71d0b811feed55e41b8c3d4227396e7269
z8130d1b5ca0ac707affe4c8c81567795cee7e9e6caf0ef619b7deebcd163ee85127a86895ab423
z7cbb0dbb3815b23bf27af1f7d4187fe1ec7506750069917f616e27125574da23d6a2b976408564
z8c31a939b66571ffaa6e7ce921812c5231dce64afd4730332a2cae00598bface9c86454499347c
zeb0e75f92ef002b8d998a124880d8be67f6525c33bc525ad1ebd7028147e1478a9c5597b2ea1d0
z67935bc044bd71841cffffe4b7ed1e2bec18e201c45a7ffb02fcafff016839443711688b6070d3
z238a8c46a679d380fbc095623d5aa110e57a919f1600b095b9e816322267423794be75591c7431
zf2b50e5f63059af76f1c9427714cadbe862e6af8119f98312e50a3564d72b37d65227e378a8675
z4274aac8e28d886da6a8d35f2733dc306177921711680cc07ba6eb23e69e74e5bcd649354123b7
za6ecab54262759e5fb78b88a51137a801b5b51e4244dd48f3dfb2bbf5e8054d53eed7add534721
zcb53c737cfd3fd49135fb518151f2ea0803833e31952286d283bfebe65bc92d894db6aebd08a35
z7e35a866edaf81a0573cb231a776f15226f4020a4f29c94b64849262e13c6498d6230266eed764
z48a0c29f777a8bb23b4526391fc4e980c516befb602ecf74e0bf9398746af628b3bec4525a2ca6
z8210d415060787cc0396c48acc743d213b9b2779ce0d20abfedcae7cd725944322a54157a180a0
zb72439a1b8fc05d229c9320703c3ea7b4ed4e5ad947e77a0e77fcdccb40e1be9865cc75d7e44bb
zf710367208aefdebbb2af161e16dbd01fa7d455d02d0260fdfececaf552394f03f0a1344be89e2
zb436b7c0a1426710523f4ce9ce75815dade4558f3bee406ec26c008313bf0f056c75ec2eefb4be
z39a45b8b7238f9edc0984c03958cd18a881171304b11dd2bf5f1341c123bd11cd538f5cf34f1e5
ze2e8a73835c8b3a14a12e21c69fc67876bc4c25dd3a657996cf37151dfcce127fea0bed5688a0e
z0ef6b2667e5964250f09295efebcdeebd6c2d2b9a73aedc5040a9a91b710c110ac05d8e2969441
za3b3dc7374a27e6f99d0ba8aaeaff27bf32db4285c5b7166dcbbe4fb0545b180b0a48977c91e99
z812b1faf9d3e65e5db8a5ae1b9d2770ad7c6f69461a9f06e8f6f542e43ed53a3a96a5599043711
zddbd711b6e79320e203b8bc82b3908dd3119fda03cb190a66ea47bf52feef3c5ed8d61b82baff9
z74ff533f04143033b9abdb6360bb92289c1f79413927e0c43d455b44151c2e472dffa94b52a0b8
z075533628bedc79b0d0a4cd471fcefc929c61fe20b94cd894b8b1f0ab5fdd3a9c4466207725391
za65a0ac1b25be82f912568a208afbdb34e83c8058f8a0b8c17648305fa9f20abef5325fd5a948a
z6490c6f11f4640f32bbc6ceb27e1595cc4b7515b2ddbc302c75363bd9f2d82ef2c1b23cd09a564
zf6f1775fe12ee9dafbb6b4b887135f0cfa78b3ccad74603588d060a04e4183b4e9139ed7c56b44
zadc42396e2d51d3c316f7d4b00591ce27ee88a5a4bf62cdea8063653c82c84ca7834ad6bfbbcf4
z9679246ddf96349cea8f136483ae565990c657e1ef7d4ca5da28f95ff80c3270bf9bd7a5403a13
z82da18043cbbab15f8cccb5848a54013ef69f261904cbd5ae216c4fdbd4d269da2542eeb2bd5dd
z289f5bfda28e6910aa76a3f1242b6035998b0f1af2a4e07fb11f4f31d07ab8c2b06bf6f0530f42
z59d966b7959424a5c61c5d666d213770a3791144adbcae5fd2241b385eed55a784ebed92b0468f
zccbbd5e1e66bd43899a36bbb27f02b92e7f68c95ad615bf06bacff258f73853267709b39a56b7d
z18cee22f55d4f736a8ba2765821c5b8a31019cf7d6d3eaa466a80d325006812701ff484436cd64
zf3c4ec218346a24c7d36425bcb20c96b6988b829c290a9d543913700bf10506cc72a920517d68a
za36b8f310afc162856101b08c53e0aa3af9ac127493dd3670bd9abe487d2ba28c0959089319ba9
z7151acf579e49c4a8ba2bedd1d2d9e6a92673dda406f066a548604d184758e502b02352bf26331
z69bf8599b67828527561cefffab03cd6b96a5b2615342ebd8ed5d7966d5a85fe760c628de6ba98
z563e7cd93f6d38dcdc0f3062389010364211a96234c21de730d7df9ae47e3901a6368c22b8a2d9
z61ec60a3e978006f3803e4eae288368e36e7a77862f3b83512a74f67a6853716fbcac9216920af
zbf89c0490f8705314635c7c12d00bbcf7a7fe60c2d9e650e96a84a6ec6b0c3ba8d66e0490d55a2
z752c33bbabe52863a5bc26f43710b686d9f2b7de48ee5ec4feeadfcf65fa9297b56e3077507f1d
zb9c6d5b2e631e9b4131488f27a2f2ed116acf8eae70ccb8096eb098b457772755bec3c78ad5eb1
zeb7c7f486330c05676f098ce0fb77989ce4ffe41cd1a7ee7a4046f93ec92abeedd520ab9e2edee
z8fba46c5ef99082c0bb49f5d3def98913005c238be1482db75547194ab5b9f887f4c1f015cd1f2
z584ca7473826f436568fe2f4a1d09cb48f0ef66e5783966d8cc637822a1fcccde42e8ff72658a8
z22b4ef1033db476372a762a14d8aa62886a45897c5884aeba10243ebf747876e49584ad4b2dbd3
z477e2c20215ca72256ce20019d37b928b69b0a2616148b73e1f975138a7c1736250494174844f6
z5f982f57b1bd3938d9d6557897e4c3a5d76459ee8cfa50127fb399d6be8d35f0a13a28aaa8b555
z63815ef24d19c924047b29899bcac18a96ae721bc89337317818c9ed20f5bdcce183bb5b499c2e
zcefa306d400b1dc56808c6bc3edfe0df6d52d11199beb4aded03ba5686340a674be2537e296478
z27b8cbb5865ee2355bef1e5bd6a74990df81793257e5afc4a1713d98f8a3613a737b037259751f
zcd43a6a3809e283c313c80bd6dd4de51189195547561c929fea38c59c3e87ab85072228d1cda10
ze3df9a5b4fc1955ba0ed6c7982c7208415b2331df710c80b0068e64b35fb3b55f58b601a6238e6
zb5214c2c7d3e56a989a081482b3dfad7575720d2031e450adf95314de9096dd19efb9a4564b978
zdc8b9ec4d2faa9b5904119944ef6d71b3339522f5f34c669525faa164543deba0545288be0cf06
z63034ed01943893b540b0986fbf4793860b7f15b8306a8862a4ce5bc5daeae4bb3501d26cf59e0
zd34284586b8633bbc0524f400803ae8e78a68e235de9268e79a9dec15a0516cf421cb11577bd96
z404a3a8ff3cf5f4e21f5972d80417fa63df1a31b1d4f8055c0f87930bf5094e6302d1292d0cc2b
z0a31386cdc3919a33f8811e9bf6828d2d2ff73da1f91001e8ced433f96a5cfcf62d6aa5e473347
z1a2a022ac4e4b23f36e15828e405a856547ba4dd3952e7bb1b25f4394f59995bde00d1c729352a
z2b7ed58abff0a33c294eea4cafaa2f648b9862b3bd597d2b436c99dc77c3a4176d2702326932ca
zac74373e770e4c775d80127764b56b0db6d9a8d01face13b2a6f5109fef7de5772e16a5be0005a
z07fccb83765f3d0d8a6a2eeba1c925b489da6c8a7029a750425758a73b4d5fafcd3864bd9e997a
z4e55d2de23d9e4fa306588318d8e9ccb29bae75dfea216ac2879afd6f78e662cac33bcfd06a214
z5e15863dbba5094544176b4f806f76f9a6b7cbffac951f8af3fa3554b9e4a750c2ab1255074c9b
z85744cbf21a78147c6a3c055e2484324dcdd447ecfbbc8e4ff9f67bb0e8029f869a31fca8aaa14
z12332508adc1f8eb4744acd71b40cc81273f35995d86ff7599cf62abf4576eff278d9cee160506
zf16c05637e4793333f41ff427bee4e8bed1ad348ff265e57c5f782691d3234edb2160f82b18d96
zf9833a47ff1f29dbd607929a22a0e17cc2eb29bcd6bb48e893633d1d76f2c0aaa29920ef6f518c
zd6159e6c0b868a25e38a4ef3d156b9490166b423488e1accdefc08f381e9457154b79b8b78a39d
z4a8402add807a9e7a7f39d02fcc96a0283b4c359065c9b6d6ddf50a266ad6e8e8903f6b18552a5
z4f46674155cd47874390eb8722387fa5636b5d9faf3cb9cbaaad4ba4e5e2ae610c53bd3175b485
z7317127b91671fbe49f63a826cd726f4fb1264458e6f8635aa15f544c714171a4c4d1e6c91d9ad
z2b0142b3b2e6d7b459dc28da0ec385248f5ac7b3ae1510ba742d1269a66923cb125f244e1effdd
z956e0ad6ada1a55542993373d9080260a89bfbfb78e53131004bb47153684029f130f9fd81d5c8
za1b4401994402ad6b56e77f9d73162221ce39b2fa0bba91c7ada2d1d3eac56b2f927e464aec498
z46ebc7841b9386315b1b125544d6bf3eeaf76e588975879c75d808c788a1830b5181bc6b1b9bb9
zc7563317d8602c448e1188e0487ff9b207fdf98b5ff64ccc739d054a3c95111f6a7435e4eaca4b
zb6678cd0c0ff1f245d205273bf6dc42908b9761c0f876c9e81aecf7bc89db2869485bec383e3e4
zb57f7c64998754438362b92ec95683d3890809542e3faa3ab8bb79ffd8a4f3986e60e0643c8ce4
z5fbcb7e992de1588ec9c0ad49664729153a1184c08c479323924567522b83b681664177d44e195
z1466743e94d0ad4bd95caba1b7b2d6463f746f41c39a5b2291c1599e90ffb0edec6fba55565400
z5e9f3c0f683125ef2746f71a6a64962c210b2ecaeb0d5ae7bf6ae264c9e306cfa78429d95a5842
z29a624f26dfebfb4107fef9efa70af007177619bdc2c90a7199fc31fd245a6ee0d1ea092cf7bc0
ze11f75064b30624c5ef86e51a7c75389121d2c516f74a6d3e61a782e553395de8955b16fd9d97f
z816f0b5d11747ac2d4d95f53366666d00f7e47095e8a7f533a07557d58a8cafa48048eeaf183a7
z2a9c7e0c73201818fa811dc43a1ae2ec22b2ca4373f96adea2fa697032c604d86e2334cca93b93
ze12af8e284450d70f0ceae43b67a60aed07f7dd82c872004ce9762ae0c615ac4878e2ce1df7773
zfbef6b25d00b577f46f4ca0707cf9eac0ea110a7685d33236bc09fe2d66f6a2344da199b8a8414
zfb9e0d6e39ebd53a4d78af58e728efacf2fcf6a972cd071e67f5c1b6fb8758aff3324214121376
z29c5331314564dc1b58eb7db8c1055d27fc236531cfc6b9b1e31c02c8757b413c4d2e5db6a9a06
ze65290d741ae94a998ba753dfb064de345fd478f94b446dbc62d5090248db1668035bd433705d7
zb63efaeed2e014fee747c4334e8cd6e3e46c68aa6212055fa8ad0b70ea3037f26b2b8bdaf0490a
z200a38031a2584cfff13b540c9f4688d4ab02bf782a2ee43d566d4fcaef7cb247bfc74906b58a3
zb646f12d0beaa0505747f4816b77abc95eed59c6003b334e4052c7ae00d542658999443178dc7a
z41b5a07f76bd09409d5410dbd7a4fa26cfe1410828e1e7154204aae427a16b391041c221f63126
z00939ed1070e61e407ca2b7b9635d738db2d1fc54d7bd18e11562cc166416d82b69fbb1d83dc96
z4ded863cffafe24c18c65a07435f2cba8eafe27ab59488f390823f4fb3780fe3bd69c44b5558fe
z9721526a2874103996a9496892ec70250bfe18965102d27613012b43abb613cd568dcde292a530
zdc7377e9f99ea9724785e1bbf3718cd288b71bdf2d1b3742fef4ce6332daddcabf1c263744f1ea
z7a91178a822029c215fb70e9624e247525e798ba3b5ecdce9678a8036c39223afd4e91e336a8f2
z285caca3ee020f19e02cc4af134d964623184ec078e3c12fb46fedb94ab75db382e6a661a95948
za4e467a02dccf117b82f1c160ecf60c5b0a01a325b435744c6209e0cb366f7483719a5b8edeb85
z15d90986b72ba28a99666a980c1887d5c56f84764f97a24e38a0f448d26815e4581af8ef6b2dfc
zf803ae8b5c25ab80ad22f40f6c017d5bbbb251e9fb01973f6f575583d2e9a063e81ceb36a66e40
z5b1eb89ee2c2aa09cb18db6087a04ee53c6ab5061734660434237c5b31875fae326c2f93ddd9f0
z8f1555f507ed7d711738d54418ea7da4521caa253b7314dd20d0ba8aab75fda757c17b8df5410e
z2c06bacef28b624715d26bcde1c270d6838bccd7090671c65bbf2e67f5bccbf744b95064ab4b3e
z13113b73fb9e07e2d64b3442bd08c0170514e7e2d2d92540c24fd7193ab6cde520ce4e912c7edd
z280f92edaefd1cf92538c7f6c67ba33432bb568975917ca81b4a00db91419bb6a107473a787c96
ze1099c71f77ed3c688075a641d6b5ad45e9ea343e99c54008c63fc4e5616c5f9660f4eda7b1e7d
z8c522042aa8c46510397666f10b08459f3e62cfed38dcd4c5ad238b23d5f9bddde2dd05d255476
z7887f4e4cf84812efc1d257ddd06893fa7d64596ceb7cc81215477b69ae051f975d302468a8d26
z30f55f64aba7abc546fcf206216cb5a1d37433a90036725c7e6451dff5b549b309bf28ec727bf0
zdcc732f5d80a49e761e32604b668630b5d770bbaa2e9112da2d002275feb37fb73d047b965007f
z84965e2edad1a62f2b0d9a66fc3a41bf1d1a681d09dbeb3c624b9a6a88632be7798ae3d4c019f2
z51f088bfaa514da254c81a5ff7b7c24a3575a90c994222b3f9a52c849536b33c9a9b5c5f6d5320
zb1be518d97f6cb3bf12ff7cd3ae4f4cb863e3e84aa5acdf48c981094e000831336ecd8bc6a3bb4
z04723e76fbc201d264b34a1e707e1272d6eabc996194e752ff680ec4b9944b9c6dc1f89c643a1a
z7ec661f6bd6915340daba19c8154964a44d273363f41cf053f3d746a0f27c954876aa88586c9f9
z85a0b3f40dc8ad7780b6abfda381091a62a3620d65a43254b09d9b232f0e1511570774c3765cda
zd8ef82fc9869bb4d249bba5095527d12db0f1cc96e995b8efd6ca126d529c834972e9e218eeac5
zac8467f847f624ff9a8f8b36acc3cec8c51af09a3e7c2490679ad305be91d017934265336a2622
zb7fa80dedef56f2c00498236f5e9e3c9118e12937c14484b7afe7a53761145075f04e8bf3b2aea
z9157d260cb8fd9ef55aa5ad97c8cbf726427ebe79c5a44cdd2241a8518a8538f3d70da79fd25ec
z42976fc005c8f9ca803967ed7f33fcb06231344cacdd6b67606f1b1d6f2fd336ea5d0271d9cb94
zbe7d1b87718779d83c7caabad785abc556c4ba92bb92f3dbe45563ebb6fc038c5ae17949ad360b
zaaff8748f039f353fbd1d33345ce43aa788c79cdfe16962ace21b848835253b6c812c0436a8122
z3fa7d09931fbc94ec4bc98904ef15764de025d4dedfe3d09a3acbab42c42ff85447296a95db3b1
z5e1ed1b9f6cf489f0a42ac79c683a80dc5f77ce108a423dfb5fc44007de4407a6ac2a9b5e50de9
z92d44385691b4300874236b63a593b305b9bcb85c55b274a4c682188099939e4eeb7eacee5ed94
z7c2ee69a5a79d69980a27dcc2a09b1308c71f4ed6c055628af433b8456487cd40c4b3149d8f58a
zd05012164ecd2a82cd366e45e256703d8357eb725d179fc817b9ce6e6e72f325b643b7bdee684d
zd48d4ef976eac20867af07b17ec42a2513d043944b00b97c64a4bb0cd05536fbb41edf25fe7851
z6485c0b25025b89a4a53d0725d7885db742d8f75b4db8f1ecc0247f6208f0629e7d0718be9db62
z7f4366f3cb07a7fc40661e39fbf51a480b4aa0ecc09876ced8e5acac66ffd6fa9f60b2b1a3cbf1
zb8a3344ded9ceec6a16c6b720e45a10e763d97bae9f9eefd95bcae63b91d081dd298f3d408ef1f
ze82d3d7034ee4c7fc638b0ad848394e3827577cfc08332936a172f562ee3de95a2c83ed5c670d2
z6131aff8ca981b4363bbb428674a92a03f39aeee8a58003c1fbd05a422c0265fa905e0ac374048
z71e2ce8de62629151aab3f84326f6fe340631784031125ab80a624967fd73604f47dff5dba7dfa
z746adbe340cd63cafcf4b93f52a90ebc58e036352325bac9d290ee7c0dd1114dbbb48b8f2a72a0
z1dfb480eab3a705b059489ef612cc2ebc1d853fb14f0331040da95bf32894c168a205ce8e1b229
zc0db4207b50d6dacda8f2a261dc6901367a9738dcaf310e79500a6e34793912ca351d2bfe6b2d3
z5364698e4d781a465cfd86f988e2e8f9b66cdbd214fcb51622da7602f8d1a375d48014e4b66447
z620f92e6e2d928beed2bae7e9dab2593930b58127c0d58bba0bf1b73f2c0aeaa52c9185a13e623
za9e178ca05302270616754a9b95b3d8c0116b0d9fe9b1bddbea041c3c18b89d5a10bd2b59177b4
zbaa8ce4e682d5dc05c9f4047aaae20f7691b95036a87cf57575b519dc6a90f612cf21f3363d501
z5582e9b8c0324e453427818d6c79c69ec6601ef34957b012f41b7e2b9fc4f0f7d00cbbe0679f0c
zbb628c9bd427be457e3d599067223e0e77fd2b64e1920d097fd74d35e207d4517154af82ee5ab9
z514e94df177ca21a558cbdda6a0dc5866e9c8b396bc99b01d1f0b222eee1eada51f4938a1e1985
zb4ca1635b6f8b2eff8b35bb20a2fde643c1c8ac2bde998f080e41e5292b68de3c50e7b2538e027
z95e941d2fc1ea1ba9a6f2344dbeb63da0392e6d0d8be09fa775d6fdf688db50aa760ffbcf55f5f
z7f793bc6f6786f463d1b82fe0b8b03b62ed09c98858b6ad3bfa3b17bd18f0e204db33a238110db
zb1eb35763d61f89d143ff51305b8052799ed9b9aaac5770fa0681ef1f4ac3464b0257a12240cd6
zf5f992c250d1b4a861931176e69c67e977eb34e198f5405bb0b5d2422a49ce18013d4f75dcce5c
zd5e499fff4c757a1d198b7e1a013f78e452dd2f54728ba3c2a38aeb819c99b3eda416cfb4c33c3
z9fa65dbc3c0db8ced2535fd16929e22883bee3d9e256d64abb6e1a8a6c2064aa48f64133952190
zf841fbb5ae6825861a6936893a30de9692401ac5cdbdbfa7f4f9bd0d1d10ad7d91e02c1c0102b5
z2a05baf09b40e5b61d6afa7ecfd280bc0b4ef9b7de52cd96af361f2ef0169bbd27a0ac24ee8b65
z14970481b8588554e3e5ab7e31de56581786709657d06e901785f2c040a10e7be43688860710bc
z4f271b40c8d79df076e5a0f721fb0c114be6f314e5f8605452f9e503618139e60faac8578b65d8
z3d8d3ff830c0fba4e57afed667e7bdbe5836d5c1f9dc9a2e88f935348630aee43ac9485b81e457
z00157ebaee13bf6c6fba6431f88501c01458d44497629e50a54e518eb268d412cfe99fd6ae35d9
zf869b689af2469fdb8416dd3064ac6b913555040ab5b82a445d06474157e15ddb1074e1b6a8cd9
zac585cabc0a469f5384c71ea1a7a556d958e39972e159c3e4db6edc9289a90a6c2e931f9bca9a3
z21deb2fef48689dad04487808ac084bf3f211cc9d7621243de613ed71f4cb8f26d192922bacc2e
z50f6a6beb9a936c073a2e47bcfe4b809a8edbf14f7babeb860991697a94e45055623d8c6c79c3d
zfc7fe5fc94e3bde9d6c22e80a927d1df037d8935d1ef94fc76495fde781d19aa78abf91a123174
zca3e9fb75bbcfad774f7e882ee508d92e20035d24c309473266f911791bdc15f558c595413d659
z04dc5f199c4323275073e4f9b6154be67155153357dad98ca2ab07890007f729bdc0b14c174943
z4e7d70fd21d2348e19c7140bd3f31eff3a79cdee2c65b93e9fb21bb21757e31abae76be94313c9
z744adf3dcba4a03957045e2d4e35fed0d7bbe8d3bee17c3e5a9302292e78fd82535bc8d670b109
zab5cb774e55537239d011f4e0e2458e6c367726f01034497317713ff0f66bd13e6ecf8fd474320
z9bf10de0b21b0fcd4f8ded1a97b509d541e3178a0d787767dcb13877435eca48d8e35b85c62a32
z6ad880407c631c606ab3a8a42e6f8ad7f792ca5724d97447bdfd9eaac5d518cc8b8352395c29ab
z25b72504b3743feb360f456e52a2a1c9216a7787655c043f67c579099bff58d9603267fbf94a7d
z700846c01b610f20267649945ce67df4132a33a8538b2002418837c4789e6f5e49c21fcc215946
zdd6443c80950054be8438923ec4a39e7fd8af491cf5b93e0712ff591f34e7fab276841d8fd7449
z3b41316ca08e686c4263557787146a041bf617b9b7e868b08a9a5bfb0bd8e8168b52d71fd4edeb
z4a1aad878f6222b157eea355a80486229aff8eeccab21b353b2d8832ef73cd76425a6ea30f7463
z7706a7bfac6ca13e08473842e77d98e637fc11c50663b55ce13521694a65ed042efbab5a51df18
z2327d75f8bafe1e151178fca8874625530850ff900ecc308b09711d054171a6b09ae77e6a650a3
z116c89c4d8ddb84fa454eb6ed517d44d102b31232bb1964ca9c286823ea1527740448ee99746d2
z4a7332eb88bf80aba937850312243f613ffae2d2f15f4f409e495b683c32d7fd58c6d2cffeccba
z80b646bc9b83c70d568f947b9e282d03c2f790cfd92c48328230bc114b2d0b53a3ebb5030d0b2a
z365399cbb51f922d2b4f467b0b9eb6a3523ed59cdc843e489b43c861390dbc0cc2137fbbee1f3e
z4e6d5be7e3189fccb484fb55d72931bb06f9e1ab6454e1ab7a288a764bb774e62552c247556c32
z0aae26075da9fec88c949f3d38111a7b22ade0259ad1c41f951607bc2692639a6ce899c4ae82af
zfff2228c56afbc8ac0b682a01a0ceddd37788caec7f94524c001537faf3b99e11a7da498d3fd62
z24b8631c3866f2182ca1fdca5ef111fe236f0a6d04cd858275d8de11c04041face4d5053da158e
z68fa29fc14ac5139b61de9534c4c886053faa7eb4ecfa6d849943fd4fe9d49246159954b4ccbb3
ze50ad976a1e1b326af374b0503a1ea3291cef3f85080e9031a1a59fdbb5c54d31b3e2db7f7273a
z679cc885dbbd8439e156b389738c2f013e5d9633c48d50563bf16b5696af1351111a25cab9fd7b
zd2f830ccb28910d1aad486118c9886af8dce536d33b9bd399c8e88faa796b008ed818d56404bf7
z8fdb6ef1e71fdc51f64e84f7e57b9c653e958037f4b04802d99c534de74749760afc2905d753b2
z439d3eb769e81321b0245312b8c127e05b87ec94d997cf0b2071dd2bed24bc872d8f428c807dc8
zf4ac458541ffedd7f518adf146e8f86d708bf3c7bd1365002223045696fab9f24f72ba6ea57313
za0b24182660fabaa9c3c25fb8fda5a7d1efeda619088f966889aa2d70c826cd3a85c080d0f146a
zacfaf184f9dc6ae9243645db19f416552a68f767be2cc0c39ab5cf1ec9ae664fb3986e9f94a3ef
zceddba6a76853c17cc64c00727a9e07e5a68e33f693535a3ec29ebd6bc52c9c0dbeddef70f9917
zcf87072caa2a24b2dcf50ef79ea0edb9255052482cf4299d486e0527ab5d4deb9a0da87b9e69a5
z10d933a4ded0db4eb229ad22a2f54cc3087fa7a265d773edeeb1cf1c2cbcb8d92d21266f609498
za61160e0ca31804087624de15961258ed5fa99798994c372f6414ffebceb220003f71cc8a4d01c
z855fd182686dd646dbe1d418ccb91528eebffcf76e5911dba53500226ee90f81086047da336827
zaa7638a8959fb611254d6b5968a78653091078fb5da34d5e9bcd196c3e97cc514dca55efb863ba
za00a264cd639e6a4e2170caf72534e5c04ca3a69d536dbe4417acd57abd0b5c154b756bcfcdfd7
zcdaa53a3586d41de8571c720a3cb84c99982687d53a03afa1a271f0ba0f68d466a5ba63b500bbd
z2713c004b1cfeef969fb794cd1a56545fa1ab60b0acf9604a485e876a70980d372c9b69fb86510
z1f9b5cbe3eea90d661bc69ab3f2e2edfdca0b44bbbd73673dc3313677834655209a2347e128a1d
z8e65f6d559a9821578b1756b17f9f77c2b43ae5eca7a62f40fa4ec66a05a0f3c4a81c5b079933b
z0162ad8e85347aac8e475c3d9a3c5e3efd899c6d85ede6c19bd393f2df84a996c3dd573030929d
zab6f93554a4e738085b36c4c03b2114007c7647211e6568986a8f82c2240e0c78f9a7526425801
z43d7fde2455621822de1c64f4d3834faef22ea708858a4e4677d8aa08e8b4bfbf0b098e5881137
z04cfa9e11675cd4c642b9ccea7c8b6a33599af5c3cd270c93f8c20a63f96711a6d2d5e258b9a4f
zbc432e679e08ed803272058b327a9752d3cb2cd9b8b187eb7414449072daf46eaf18d33172cd87
zae53ed6bf1964dc7f71a22c045c1b467c098224de8efe69ac34148be966352d6f343c76960f95e
z5806722f65936c72a0ade39fe9f810728bb02d7ab76e3e3297b1fdcdc6fae8837daa0c4d337756
z7077e319308d5f8549d924b96854dc29ff222b7195bdf12ee4db3d3299bba5f8d13207835a3367
zca93f9b3d9b644c4b9733666dae996a45e62577786027d3595b06d6c285ccf73a515eeb776c7fa
zdb2c3f51757f96b443bd9963824f2998db13953a2c039a134be65ea75e0b6359fff0a811a97c11
z0609df6949d0c185a53d5b881260ab4382ce5b35f371144e63f168889e6e684d3d60baff5ab48f
z554288b3a8e2372cc512558516ba22562fae299b1aff476632444f1aef99a0dfc61d0a55cd96fe
z8cd2f864f248ad9a8a7420371e2482f174e788e74894d10a16f6a53f472f156eafa351c8ff0bd1
zf25f078f40db36b95383b6543ea1548959ac8e2b4078fbcf86c02fbd82532281215740593335c6
z5c0fb25a29e69da5e84e8bf1d82eac6e748d95d73eb7f730c5bd89e83a609faa8412d390bc4890
zf9cec0f338a5268c4896366c031ce3883e0ffb620544fb17c947c0b2a2920d8ba34b917878ec62
zf77bb1b974a2963680220aac6d28de40c5abfa02799e91e569a3755f63edb0d3a2770d8096bdfa
z8baebac2bdaa7b8ac6f2a021fead91ee7a6d2f2c792c9e92a28455559eeea58cd479cf9053ef7a
zc381e9f612b590aff5347324d4ddfbadb9baf8162200cd67cd02af7990df036a0d7dc19e8a6c13
z2f136ddbecb48afd0fbec088e1cccf0c9005bc13180cf63f397f0fd7a3fdc9ebff4f95ca8534cd
zcf671ff7a08510529de7f050c959e400211b05fe7588de5ca82955f81aa39c68aa27e56b3a7b4c
z551b5d1ac58bb781318355ca5068409560f169a80bd20fe319d856e71d218f144831f412e89186
zda391da3fc5c8f02204a7509337b0876ba8ff87eb63687c269ec6cd6e434828e98a8ca3b96b593
z33a317d7eaea04a5ef016e65aed4a87f2d99a5e519b1c5a19577091a15d649a4539f40dace8df1
z15d42f43b5419918544f9df46a56c85157370bffa13ea1c2b45876357fc9b8690b4e0943b64ac8
z8c1835cd630a2c244f48279a80765096a12016196efc2f39e1275cd019be497322eff7f9c6f9ba
z765a3eeae178bade71e05bffe1b5e8cb2959277466d1ebc1381a63f1102a060f101387e8c18e63
zcbd145b575cc8ce551ebbe058f0bfd757cdf8b9afd9d975a71692fc8858a661fb407b7d56cea7a
z1d670a25937e70932d9ec4cc0cc39fd2906606fdd6ee41cbb32b2374d6eaf67b5876319206a191
z5893bfecedc0ae4d23bfe1a9325ccb7d6a993d90aa6c9c50fa20826bcaabd99b70bf0c1e55da0e
zf0062eb24e607fab5064d87970efdf306a3cf7af7857f99f76b1cee4cadc59822e8d0abd48fb5a
zeef76b17360324e55cca7d9235ccd6193f9ebe752cee5e3d4b8aa347d4910fa4e90d08ea16071b
z442159a9e7a0cb5d1ac3057a4d696df0d9019d7967480bace483ec055116551bf5eb45a57f8e68
z3b3ab1dd4f825cec75cb805ab3bee76148c0d80c64faa3f3a5939fc05379d4c033ca5eb0f2c4c4
zc4d459855f44143b8b10ed090c327490e47fd05144d60ae72f609aeb4490af474e24d0982c88dd
zb7473d40b25ee22a6b43de37134675aed43be7adbc0c9a517665e5899c66d813d044950aee8058
z510770432f17ad39e24fb94abfa1574a8efacebf85ae2d3eb1afad18baa9ba2dd0c92173c277dd
z8454a8225fac5224e5766daa86f50eb22a585857b96b1458f9f06de011008ee3f832cf56084d17
zb8c3da994a8270c0c1883180a3447ebc643660d0407d3a605af8339d167e3cddd6ae0e6e328563
zb536fdfbd78068bd09ed1113887a3c0a80260ef2bb76cfad04e8e26b23334c94f7ebccd828da33
z5ed0c1158a73d0a8bc6d6772e3d2e7b33fb721beb3fcd9c8427d811a872fa1bf6cc4ff335a0b27
z654b50cbfa394269f0e5b98516e167217196e05318b2af1e4e1a075efbad12f4a3c096f875d981
z828e0a29d410d7912e108273e8784a0c998b2d81494bc54ea0ddccd8fe114811418caa81a51b1f
zf025c4e3762e5f1621cffd9e2234e1b62abc7ec461bec577d27c0425012c3ae62fabcccb3bede0
ze7a80fd18325f13aa93e9fa45787be06d01083c1d678e6bb1b61e898ef655bfdf7ca222ba91010
z77715667ae77fcc22124ea4b2e0c4532e2393c245f0ea0eca85c2786e15e5fee9c95023c588669
zfcc3b1ef88973f27bbc1808f3c6dd6eb86bcf891c640f60d94c93a155809e287928102afd4b57c
zf349540af03a4884962a8ae4e5361a92fe97eb74e2e1d472a8bc8441f003f6c5f423202ea64f45
zec0a2f4723c325772069c33642fce2ad0a3400a765c674ce8337e6b40121be51a0c9a238a920c3
z9456be224369512c4c0a54a7327f48d5dcd5858da0840a2c66f6d9d1cc57dd090cbcd6161a241a
z147291429eeaf392ec5afb8327e73b50bd7888479c1d502f1d709960a0f73ddcc20acd27e17075
z8a81ac529e4a501380b638062ef2db2bd6378e25ba6dcc27fd2e956954f6ae8fac32b83c51c1e4
z199b46df5c2ca7dc48a4a4be5cb828546c59a79a939c1d1097b55ec24a17aea95184f353c335fa
z5fdf85b2f67330dbdcfdf286152fded2e2886fbf9b9696898247501115ee47a68df9bef6a63307
zb980fd5ae0bdce12172d2c4831dc5708f9323071f94b49a5b94eaa0921863990c6d0617553e5fb
z2ba942d8787d884d475a746b8df1c1722074151cf370b6a1b79acd81024f800854358f685d279a
z4c6f95103ffd1597505dd80cc8df11ff750ce12ba5ea479bfb0ffb5f9aabb6bca4596327259240
z1f1762c47d1d035e235d99c40fe0448e8ceb2abac2a72aa0ffe0d5290ca18ecd0e014e504adcba
z95238bb008958582c7cff25ff6fd95971fc3279ea569f9294a50b6b9f79bdab81c3b8d5281ceb7
zf229f3c903edf2c1d5561d59f221f583bce7f6e76d0f6cd3035fd8b17c396cf229ec31355d3996
zee0cdc500543d519b115a1c86383653bd0d7bccc06aa332fb40e377d6f2af7e29aa65cce38e6dc
zb3295c0e14f5444d80316916f437e4185ee8c19c459ea05ca5e9c233c198358f3b13ee352a38a3
z76b8975432c5fbce947536d80593ac654a540605d0d1f228277d6dee52958f27f963d7e04c35cf
z21b10085338a5e7c3abae43e3ea3b55e54b6e014cf74a52d07966f7fc28aae6d2efcfc921b74b3
zb08961bdfd383191cc138f5821f98d031022395f85149bb3e87fad05f8d91ee5f78dfe7029c322
z53b1bf3241edf97ef3b6692a14e8dc6d6975d8005199acbed723ae3893ca23c1ef8d566bd54c81
z721ddce5884a11c6350b19f4bc0cdd3f4a41e3facf73e15ff335b703663d47687ae352323d27cc
zc271700c52dee60126b77d18810881f4d31a87adf40c3920accae6470634bf3d950a54f92b0907
z414fa0e81a7dc0948585ba168af2b7a0efdef91e1dc47d362287b0e33f982cc12a4085bbe133c2
zbd51ef15785b1d19cbee3fcc26bb30d5136c77a7789ac069051f8f7e3c990222f841052b95c960
z491c7d42a3091e701671996facd4a7d3cc1f29319131665312babd460a82cb401a586e6e3a99cf
z83208636942dad64ad4b37b8a06259c81c305366c44ded25957818d18b847d6b409373e2f49da4
zd330fe3e109841b86dbc45dd7d49082c2c0d983ec6184d5427ef60f3e2c12e764ab0f3ffd3c43e
zd0d00c892f11ea7ab92bc6b9b5a30937050250dc86e24465f191af400d4fd61b40b1544d2751bc
z2980f6b8407366387704b5c69d85a61d52f365e6f796d4de2ad863b56dfb50aa3238d41163abe5
zfbffaab96ca5c011c7ac7bd6c9e2ad06f4982184d345c9745878999f7c8606e0967124bec796ff
z3d9b68bca9f881bedceb4f305c0fe7e1885a43cfae542db87fa41a6d02c69d9764792f2ef04fe9
zeecc5388e2e07b583eea07b2017afacf69cc3e1a3097bedeba337ccc93201c03cab63c454fd5f3
zd6cdb3f321572139ce5a408b7ee987d18eb04df39dab6b91c5ce0e3a76f84808cfb6fc744f50cb
z5fb54da2a26456b8efdc12b83d54892c19989457027a907f13d3d7317b07591703a3b98ac8ea19
z14dd1fa6798d1ba0048b59c8573a407a81310fb4d662aedc61810f33c7cde169af51e0e35b4cc5
z4d55689f38de835316e594f6f19e1aa4917f538fd7cbcc39c759d457a781b1aa07fb0564c0d6ab
zf8d0efef6b24907f18bafd65f1866d29a256c617946dac06f4451a9efa5113e8367d64600cf6cf
zc1ee85e6a857d1dc6ae5fd6582e786fe158ba43dceabfedb6c840407491ca0d0e87d2baf03110f
ze6ff33b3b2851ed65cf07693ab8925ae0c1d6b697e9fa32ba9c2af1a337d2c6c1a4bf96527441a
zf2ba6625a75677fc6548a0b42403f1cd31ad5c2f744d5cdbf03ad48695a704625d62b60b2d0cad
z94f9161e8001992a3d272232035b327807c83ebd3fda256cf13a89c22ae5e1d73c29863f423dbe
z3afe63527ec120681994b8926891ff212c6a50910edffc1effb612233b4cc7e55ccfddf85b8a27
z5b595607634b6c650ecc2f02ff3cef4710c141db80f13ce064094eece41dbb2be231878396e2ac
zc81159c827726872c0ebe33208982e5277b5a2eb23525f923a13ffd9d83f7350e03ef79153c292
zf30841a6667a53075aba256fc65a9fba4979bfc375357e98f839da112dbd4bf4c0f52ea32c47e3
z1b74bc33d6f146d9de740c39136bcaa3f6be7d02cc4fe4dc8b82424418cb20e5a249f0b85fabfa
zd2d7fcee19d12f82d5a2f02e8330c6e6f9c13218705ea31d5be70954dc9a2046a8176a629f6d4e
z5ccffa98f0924c54f341fe7fa3e4c3be942ece56f5d01c3b3d9c9bb1f78119da2b96044394e540
z2b31735c7148859545b4a8e3a101f07110ccf0f1ddee719453cded62dcd76beed17b372b635d11
ze940eed4cae14c275603fb979b5f8d3e4a9f682375334fbd79ab0f60f6766bde10803242e47a8d
zd813d22e753274a223f2dc858d97cee2e3a0089be7086af923cddd480c9cf21830855b40a257d1
z27bba58afe0949199fee86aca821520bea25c5c7638f49c7b55bbf8cca54f24dd89040565b2477
zba706840828ac1fece24c6a6906bcbe1eecd0acbda5ff40f8be217ea3e7954479c11a21003aef8
z0f77c9b81c45f0cefdd9dd20ae0baa18dd26dfa24d6184977832318d0eddb5a1ec84010d10e473
ze53ac04f0fd44befe9d769cd1add47a2c0a43104dd971002b31021d74fbf6e700a3209c182d9a9
zaf4a9585196a2541d54d2c8a4948dd590bc86ceed68df43231d08ff74e3e5047cf6c9958499e9d
z4e4a697741d60d0a726632f695a33b0ceebf839360a8401e91642f64f07e76ef4411d9336f5cb2
z00fbf9c508c613ecad4443fd35dcb8fd07f4bad8373edf02a6020899f73509fde05f1ed503c4ab
zc5be2181ab43e7128e224294fb4f483be8bb71ec3cd639a4cb9a00e44105de1538d3c0d0943f0e
z7a45a62100f74c4f63531e20d05a922b143771b25939a7b4d75fb37a11ee2f15e43dbd4abd812f
z45d430878e296fdbca613b8883de35ce7be2fbbb09f61ffce7c55f9dbc546bf455da0ce6c82784
z7b7bbb60a2d142fdbe0d109392c9b39287790d24cfc79207180c7e3605737ffc392841aaab3ebd
z29b27d8113026e33efdfa253992f293818f031374ee8f35e5c6fddf3fea80e7038c03b44aebaea
zc0b120ae82414f73cbdc63fa352e38bb7c9f54e27564780be49058cff819c8885caf280333bf5f
ze81a0176397fce6e7c6e15d297eab64c8d3ac626f2fbf295175f7b84d0662fb9fb86e2c4423bc1
z5af52d9e860b4eb969a3fe50ae7b1817e30d2df01cf82d8b26d66733a259d0e61ced52eba965a9
za1c4209b1aa475f2671dd24f849dda362e58dd6a84eee1c4bd4368e1a2703cf48a467c3405dcb9
zd8daf0540a6caedcdc2f67ab40d1c4313e49333e53b62ded5369068f78887c7a8a55f712be61f3
z259896e4ee8765d3f813f187d7f5bd195cf702b2c5d888fde36acc07df387bd2f1b3e54147597e
z5dc9c295345f6359f249fb1d9553353f6bada0641d633bae2d4588ef39e768e7c6cb9eeafc52ba
z19b8562b3d9511f8eecb4daf5e40622f8fc221b5a14f5ec20121fc0a63036071fcbba098bc6e7a
zf5886054bf7b7bda64060e9febd7509b38eae42d4f344a2627b229e4494295bf06ca3b5c66d788
zcd0809a639277b4507a71d8e00a816c82372dedbd7a0bca3c7bc8b5971d529156aa86a1fb2633f
z2f36dcc80e2d7098142139d8327fdc31b7d06efa8f73ad730fa5662a84ac6d67db5afaac25e066
z0fe84d039296d1fdb0a9897caa9246755730492fccd275277544807905ae5cc4fbdfd1cabe0c4d
z84715adf82ba534de3684cb462ae5d9146da2b816ad7d81eeef610815fe3ca4a49e84f0b6c020d
zaec8ec830c273bbbe8022d2ff9e9e772031f9debf577a6a5091a4c24d4adcdc8d97efaaa07b388
z497b4366abd26d4c41eb754f838463d7182ee9ed161c1f9e0408cc3db82087d9204621f036a56e
z053682103bf1b6985157c19fb916e879dffcdab4a93abae2715ef0f748cdaf243495078f5fa66e
z5cee19818d723bd655b695829459e8385b675a01615c385ee1969b2ab2456a367043427304a64b
z3e8832b66b71a132a18097015ab3fbced0eb8bbce66c7909d3085e30adabeb66de8996de540dad
z648e248c9a8a2e112e1d67098521e0c359d2886a533817cc41dca0e25ae041441002a6bfecbaac
z1ec7a49f51f475cba7db698e53c0221583755b9bb4955d803ece92335f7edf02150a4b001f919a
z22ba2a82a9c59297c8911a65b19c54fc2b2fd8de51da4e8599fd8190e6cbf9964627d268c9584f
z046734dafe84b39e4081959d409ae4d649f38c8150f28d236d137b072eb5cdbae65816a1120f70
zf4b116fdd2c16e1f446f33cd649dfd6206b1d7302125c473fa0792514e8349886e005fa0c1c3f1
zf828089d178c2644345136c01ae1e1e5cea23377e26f4a997c08cda499724097b5e896c0ac2de4
zf19ecf100d9114fce4ec2ec41bcb153edf47640ea9c1ecfd33f44336759adde4cb6b68627e5f7a
zf1e681a778d2f45928c70a697f2e0a4d0164538bdad50ec289802cd6cc5e73be836ec4a5ba2cad
zfc87ffc1c194d17dbfa41e56f66e8d83a10938d5a965ab6c649073af1c471a30ddc4c7929dabfa
zcbeff05833547b84e6e7011a8a9bdd699214f03eff0cc02f41b896844373de3c5ae46aad45179e
z823b8ce768838388b32ae1ae90f53fa7e194abe99ed985ae635628ac00e761fe4fcaf8195e6130
zf1c464c8bf7e17c4e168fabc5e536f0b9e17c71f21ba177903dd9ce391b079cd7a1c98030ee9b4
z1beefaf6c48f4346dd4223afcf31cd413d4dc2b9f722664fe40e50e36dadd8921114369781d5ec
z46f62877676818ed3594d2a9a54dee5e76e3b55bbe22b25707a04eedd001a9f2359e43aaa9e2e5
z1222377b66e88fb8c8fb400b384357982dc3f17c516182ee460ce5d91a8bc47426758a17d7d2bd
zeae1a28c958cb10e72ff918754cd165fc18e1091576b7947df342b1d76427ee1c1d287fb7fa920
zcff26a6132dfc2a084057e306975daaff1d8d6ea58153218c4ae4f87853bef168f19c3dea337f2
zcffaeac0cf3637ac73b0795f127cb49a2c3459ddbe9bc34e68530a7a85ea4fb53d66ceed644367
zde9e3a3bd082beb56d013259add8bfe19aea44b81bd37a254d446489b3116cbe40497eb0c19334
z8623a7929102b696127956707d9a94b0b8c68ffb4d7b4b42fec44b697541ad5364b73de7338436
zb306eee04a5a29ce1f0118b34376f57b66a9a0b1a0cbbdab40901b2face55933add80e14ad9cb4
z775293079d1b264d95abb57b581fa61cd74915b8081dc02bfb880567159ab5117b1b332d54be6b
zb9e0563fbd23b2f049496d823a2c23e8a9c968f27f98252d955d17b888ae1fd5266efa0f5112a9
z50b200c2b82708aeb38141532ea3cd5d65be4c7182ac356119e6ae061c3a95c19a121a2014e2c4
z174b0ea25c2e93bd8f5eb5e6ff128a53bcafad108136993f71a69d68a970beb54729980788daab
zf4eac1dcbf73532e90f1bd0c8ed962348646067605bf8df36f32ad8648ee45d8c5c5c62c088a4b
z0473eaf558d154518bafd85e21a019a17b95b3796e4106b54ea2934a5ab03bc6e9acf7c5e26efe
z90521e1b999da6f52301c9b367f6e302ab2f63f28ad2aa18bc454b795b30ae4ad1c85159e52198
z072e5817ab173a42e3d8c9af02300725ec5670df9cc76daab64f59dc64084625964f7c486e405e
ze9137d795c8e5981c420e4bb6ea1cea3543591e88de583060917737c650f0126b15fb9731a602c
zde38a9a09f761e1465ee2f6e9b9a1bf5e4b37fd1f8ac60047237526fb5a265c7ca434d11c5e6c5
z7c60ea4c0fa93f9afae95270e853cff83111e1c3c0fcc01cb85c43a6ed8cda3d284762ef7843a2
zb3fae0427c90a0e749b847475d9d4c00459ba4b9d3c6bb3830f395e4b85542492515c40c73aeae
z7f6f212531deb46a943e97cfdb5c066f720b20160ce44a4a8f1d83af77ed8e95b425535d685990
z3aea85444e3f4968fcab46a3c24c03eb8520ef052be3afb6a4029d8de1c6b6bdf35977cb9972cb
z58b2d6162e8928eaa4b6344db8b3d10802abb47565054f9983dfa9e70c9b24db0bcd34cbde05f9
z78fe9d0a81bffc21078918805daa5cc76ed2d4cec674708546bb68da25eb98ca67cc5c2668f371
z9a9faf7e42df0dfd5e7448741b944d7183289f7e7e78f0b8659caf4a8cf0b46130e3afa0751220
z48034fbcf82d991b723aba7f76510c28cf7def09e3ab3f4fb9b8e0ffc89de2514d114383222d9c
zcf15990ef8b4d2b86101020147ffdae8614c56fab496413cf1090bab3db38cd62296a5c0b5608f
zb8b3a6883ebbd5d5f9a9569e341ec4f2dc78a1976dcc1c9edfde119e8aeed799391ff4d8e81d9f
z947a60c1c87aa85089e75ca385fd46ddac9c99acd306654d5ea4643720aefb8aabd40eba8286a5
zdcb3adfbe9eb2c3cae1af218858a30bacce2c407359cad2a75564fc1facef8ebef98c047c53e6f
ze6bf09d13cfd0c24c5390ca0a67bc1783b94e4bebed738fc4c65637562c247323ba1c92f07dcf6
zfef6c5368a26151773c94cbc98b6991b3c56f16a4fe600fa036f973164d518ce313a1b7dd8711c
z75dba116c414fc9e81b05810cc129f5e83a560080793555de0ab5e199e22d7473391b5e7a5d063
ze4978d15f4b415612dabee698c24aaae7f1bc21dd2ff33255f38cafbcc7bbee6a69c91e732da96
z7123678e6e3aba05cc0be08d4fda607c167ddbbb299dfea5e319bc7b04c47c4d6348e060c84647
zb2f6f1ef6c5dca70da9003936345689a1c108c56bfdf8af21de21c2b50f92fa9113cd1e52dda88
zc2b9b3030e4ee955ff2fc71367cedaf3533a2b6a35bc64c1a51181d0dcb4dde80fc87a4bc57331
z6c151a0c364b1939fae25436de4ecd3189ffe20e7cb8a5edbda2db408097448763dee187752702
zb34551520633be8a298a4d124e7787d4eb7af33fd38ddcb25118a28b968b4eba16882e0e793c7f
z4b4457af5b644339e0f23cb9c03f6e5cd9afa33d27205c2da5746a183998cb19eb13a0fc57483d
z55e3591ac636db994eef867c499860cf97889de7d0029ead78f8de3f7ce491070b684e782d1df8
z18e11c18731690fa4c2d6e46f8e1ed8b9f35745e2b017bc9ab75e785859902357c9ef23a356731
z777dcb9c1f0bd408dc31932d8ebed05c1f186a55d042409a9072c0178012526cb4f07d5feb5cfc
zf097702ba541e0c47ba6cfea31cc25891ac4ef61e48ea9ddec6cee027d65dc725ac67a908e93cd
z4520370c459f8dd417597c388ebeda0807d1a4ded0ddfa0b56a433c229441ad8b79a6f97d86381
z8e5dffdc14755d9cd7aa6c1036929c7e9ef045aa3c93a6f4a2a36ba8406ffae05e80e331b11312
zd0d6993701fecfe31c9dca19ba3a5de3617c715a1ed0600eb12cd8fc657c3eca601baa8972c262
zec27be30119a6dc406ff77e9f56fa90a8efa30485cafae35ef5407f2e835f3ca76d17a0fa10d36
z5edcacb7b3f6a54822fe1e12379d64ad8017f0bbe3b801ce9b39dc707e9fa7fd5e603a3ad6dfd8
z86aaeb13864dc430a3c443e061f9b3adf399a2337345b704dedcf3077deeed52b57723b26640ae
z4248c31b51fb74189c0026666032c6d8d8da69faf5f38ac9640d0708e403026a00de8e0eec540a
z8b7531b087eaffb0587c80b4ecb7820f00075a5b08eaa06e0f2d028584da6e22d68452b5f0278d
z80d9f755f349dc01256560d1346c85bbd898cfc7dea188e4416734f6a628c54b62bfe10cac65bd
zc8858c22515af0b276fe2fe520b25bcbe78a1d0092e4f48d47d591ec29ecf05d4a023e0d7e6891
z61ded6d984a6f0da193ef057ddc443d93616431d8d54c513422ef890b48254bdd747e312e99015
z538ba75cae2ea859a5f3c1b8e85393a53546e8026850d7d51ad161900c4dfa69464a6bfa686a1c
z57b0a17b1abb164fb79417cfa7571c6d4d5b4cbd9abcdfbba662d4d5be1144bdb7e6553db8cfae
z212393ce5848a04d6e267daacff7c976ddfcd465b5aee8ebf43693480d3cc3347e02249683a9f5
za303ee3af178dc9d31173e136dc9ac2d1994d2fa1784737a19ba212dcee5c8fafbb4894a39e23a
z24e2ddbcb8af3f0b8347648580350bb2237f26ea956b9f5a5dded75e6bd4f9409a4d8e7d506e7b
z93ab26d37adb647ff038c4347250dcdc323c6c664c4c3823220a27bcf3f236514bea9aaee3c1f2
z0ead3f2c84a8cc6b101ecd027e3fecffb2d405110fc90f45031c9bc0c4faa8781d2537c6339aaa
zc2b1a3e95b5ca1de8579fe29ca69f7df717d98de41215b43e12dbc3c34d32b60ba9f261c9686d3
z5b7b8f58919127200d61d48b6905c2306d06e0718c27c43991ad023df608d321def5e8a0f4f518
z0198e582aab3bea0092d8844dcc8deb0f93c4b95f50aeded523b36bdc1cabbad54e448411092fc
za3cf8bf39dc41fc629632c37f143e629e385dfdecf320d9bef4d6b448614f223aaa8a43a68f293
zcfcd76dedbd5fd3e887ad44b63e06ee86286676806581eaaeda2b5d1f617121983984d4a49a2f7
zf453bed0980a71fd00c7a45aadffc2d4f4ea74b16be768d0a04a7d51e4faa92c92bccf009bd7b5
zfadb3eeb0ca65ef953841bf20d7518b5151d6940e6017b176b7b17f75901d870d5844a64e4054f
z9e38632a7020e5bd5a05da99c2d5b80b68078c039e9052d2d6db7d6e3ad495c9f2b149b43af41d
ze650e46937ef8f68d4e43e204af70a7063baa57d29ca91ce988178c3c80c481eb8d223666db0d8
z13f9a60550132afa1b2adc2c80d876448facd1a4428ad7f30f40d58bde597d40b54b7ce02dbd0b
z4aac3e69c84ebb0a1cdd34f5538d367c83c20df14ed19738b28588f47b3d68e2e5fbf32c804a3a
zbf10ff3cc4a005e4ee71f3a5e6e2c834363d3db065d8557c24ff5acafdbe2793f9f0a19f178fc1
z6b55c16f93597d15a49681dee4f51c04917848f85065c915399453d8dc36cf2c196346fb1e8d5b
z972464437f9b05ac964aa1909cbf186eb8eb64c23be5f4fad7896191b0b7ab1344f53aa7ce4a6b
z220965d2b2f5b3ceb6f02babc102490d240075e5fcdd8be8ab25de3226624c8cccbb484af3f8a2
ze1d153b86811eded144cbdeedcaafef160ed286f0c1b3e879336a32dc956fe9ef3df5f87841d39
z4a40dffc388036a32bacb9adf41353946083a6c7e68caf35bd19644e777eafc7293d0d3cf244bc
zfb0d25144a9ba32692ea0796b7ec6b2d5e1bc32ea0e971c65f03eac4c76abfd67ff70398be789a
z9bda83619b62bcb64027e2a3d3f4b9e29391836a674454909b0033f0c12594077eb922385bf562
z500e2288778d5c381abdf7f82dfb3f28c8ab08bb33eebb0ea0e3a889a5f7f7b0c6f553d03dc0c3
zf655a1a289d72f459cd0d50e8993dfc8838c31293f6ecc7d488d01da0c8372e8df13857db014ae
z1745d2b991f86c9d6a807fa4e4a90450b9d812a57ae630106b07f385c640492f46e5b3b88c4948
z6963c78abed617b03d35e91e6cc7728f12895ceed034cc8eacef75a83bdde26125c6baca19f310
z5b88ea4c439e89f66faad3215ae205c7fba3edeacb088b547a87cc13790dfb6c4c53a7c52c58da
z8dd21f477912112617fe4d0b9b5ff39d2979d95afa080a4c802bf51e479b23dbc54eec35cfe8be
z348bedde0d80aa956e388355fe556864e0cf55f4ffc6625a3bfb1d174b5d4a156ef6649a45df8c
z7e6104d714e4b3e1a7cc338ae12e88ab3d508fa3be31e2e329cf50705fa34bd5a979cd8846799b
z483f87bfb8478f93327cbae92ea76b6940bba3cecf770bae77d31a16a4e84f9ee1bb542e982d1e
z874537c04aa7939de01521da37f3352f9c462c8507d6891d857470e2b43d250b1f99b7a635c3a5
z9f2c1660f5db2d7b0405faddb607914f0240050596c72949aebc1da4389c4c03b26cd984aae7f4
ze510c680e7b2cc5e76c69e274d69808fd48e9961c3cb8f53454b4e90a2ddbcc5856dff1cf3fed3
z0a1a1e60dd39b1fc6b67d3d99ae467368aff92f48cb3ed0189e1fcd90b09e089bd3141818a2911
zdaebbf7e2827e7a9c18a958899323db6d196309cd3b65530cb960508369b66828acb440b316813
ze6b5cb47df2d8904e062f33804f3c3ac94aef08e8298b0989c3ad28cfec21b3d386a3937f3e25a
ze4b9fcf96843bff8cdd208a4640b8979ce7c94e1d8d27f89a5746e0a172fef7d3ea5dae9930edf
z5804f653db8fcdc9c6b56b111c83ff413eb30a1dd2b71fd3cfc8ec3a80f0162a98dd1f21892e71
z4dd67368ef99452aaa1341684ad98469352a17ff0d0ec22281691922772377dbd27dc16ba5ff41
z5572716fffa35ea4a047d5fdd4b8661dc5590395dc3e3c64f190620be3ace789be7a4a526dc39a
z1bf871ddb88581a7ade66937355a0584d10342ae9e59fbfcdd0da90958040d4dfa0da7c4621066
zda4dcb657475c3cd3591af1e1ce0b3fce753a34ea7d7f6755472c661ce5d21769f8498cfe28e59
zd3152497dfda8fb29532259de5dbb8b5ca0e88e166c4b95b9e62c15e8b81dbca0ec38cb831c7e1
z433aaea1df2e60254fecc5db243dad85509271d28481f0a7713b6abd075567c79f37ca69b000a5
z181d64aa74c0f3a3a98e590b07559b13ee04996dd6fc1e6cef44685169513655ef72deba717092
z75d5ffad5f38f18e1225e74b979f463decb8ed86697d8a997618820ecb3d9c19a5539feccb3a1c
za33aacf614bd35069100bf67b0e138a00a7b58ba522981f87a603a7e760b15b40592addd7dda18
z496cd22953c17d6ba69dffcd1719098f53dd89f75623cd4629bc4ec6a0c3c0180f33bacc5a8c70
z45d6f8a80c9da9e82dc384e4ce1b11902994041bdeedb209ed72b353d74c224b80eb93a2223b1d
z79e0f1490716d0b5560204c826f00719aea0325e454a811be56f3802efa3492808a80ae8c917af
z21bd509f1ab4d0849e5785d43ec9aabe21b1002f0f933ee2a51be9d6fd6153d1fec10d25a190ef
z81689d18d09257bd72040aae2ba8b9981a674cddebedfc4596e68415909662ec4dc2632adb1314
zdb7dd549574438f7a1228f43755be27a84e3d9b9e1dbbc62662522d84874aa82243ebfb5d8103a
z3382b63815e6f3e9736b92972855a562664f8e233a753b8ae485855dabb94fc4e14093e92158ce
zbfc53495c3a9a1527f7834fc6c80ba93a516b680072dd892e26a44cc59b633ab65eb1d36c5284c
z36515cb253b73e653acda7d20f9575eeced31bd2045fd180132a2d0906c3b7f1afc6a13e2c0559
z5ef9af0412ba22081a76ce3084b7bf3fcc6be1a9297d8b80c08e218c78bce5375228b3e6997d4f
z5f3843e172485642baa4b17fb11e482f0eb6f4719ed7d0870533939cf80803b82b193ab49a0a44
z9b4cbefa01f650dccc316b1a97b1051786532d883941b3049b1b649b019d7fc56c6730782e110a
z009e29eecaeba772b2827f36351a7e13de6111f39d02936789374c89403923ffaad52523d17d73
zb8ba9925888b24c2e67a75a2e4abb07a8b9b7f31e8b378eba6c7292d1df26c7375fabda15aad17
z0c7ab46d6d32c30051b74256df3004b171db57a391692cfda0a895f165cbc7faedc43ef4e17e65
z3e045d06f1fbeeca6c1cbe20a781a3912c25f4cd49b58d6137ebb92b56512221e79ec1069bd543
z99dd69e21b45f9621aa1fd277c1d4c336287ecfe5a714230fd5da600a8d44126517d93fff6e239
z089cf1401f5466a0805680dcad7f897a9cb2ac867b40ba36679e2f749a0e9509e3688a1e744f2b
z84463df21d3162ae545d26169456ff17bcc9b1c0e0772b5df785f878b522b5ce217ddfb8311f8d
z1b66154c1aa8f03d8265d012bb70bab83f827c291558404d3f10d1cc2a46c2599c17742f8b18cd
z6202d5141dfcf9cce2aa1af8e1a7cbe6eeb1a38415656214a542190656aeba909f0aaa02925eac
z742737fa12e1acc5e9c0bb8e82373b28c3d459f03f387fe4889283880a1e56e2e335aa9121dc44
z80b06ebb7bbf9b622cff8287bd2e8a30a858a60e7e804d8aec25556881a47901e244dd1d12da93
zfbf89e1ad22bc0814c9f7692b611c201a9ad74a0e0cdfd34aa13df91438ffe04df416bd02e91db
z02a20eccb47fc7db6d19ec1bbf11ab5e7e9d5e7555c343a2d8e8ad3f8075bcb4f719122249e4de
z7769893d9b697974e6f1a4d264f02e104efe6715ebe24c87510f2ba100859981c64397167c6a33
z6e791392e9d55ab7257c7f2d18b2ca1dd8a1d4c1055ee7239c201279d0fffb0a6b2fb0f1f14616
z6ccb5a62729930d1a41a60b47398fa51c5ab7c3549745930f43ca26e8ca4e170680bac7b6a7c0a
z17047ced5ff896797a12333fd4efbbc3d5b4ba19269dbed7488ffe51d469c6bad5042fb841d4f0
z6880026b33791b09547d38970f5da66289da6ebe2d3e4b46a75081def9baff5de11513de91dd6f
zc4bc4f77b775b3b38f8a3015444688dd1fb5057521c331538e6870880b286f834bf82b325b58d6
zb3233f9142670cdcd05068d186b4af7b4f957680075e297add1321907f8c8afd344a14371e4028
z8f77352e1ece5fc9b03de7ef1ede374f0054eedb1a5696b84315e37d6ca3526240d4bb74da99e4
z4ea7544e9fe46bef671bbe6c908adf07b1136efc9f1b2a6e4347a371f674da0398c59e4aff6065
zff15db3a458cdbdf4ae98e845988fa62cdc3cacd8d4414c37ed24baf307074a71fc771ec4b6cca
z09f5cc6969d39729edd2bd86c6026eb10b9aa3b652ee0a037d6e58fde0fd3e24539c27ad714525
z0d18dc574180f7ffe6219c3bedb8d8590140b37375fb5e122357f8adafcb1137397e318a9c0b65
z099218ce3f015dcdbb1006060728672c6d396734b6b8408f8eb2a6d4c6ff74c9f096ee31aa00a7
z8c6fd8e7d88463dfd2d6ca902008c7ee0982beb964ed321a169ad6fd24b969476946def2a3f514
z551610ed3cf7ea10fba57751e5b6fc9c1591fbfd42d0af6279743f2aeb00a89d302b94a3a3d3a4
zff8c5cb616880c86e1dee2316b35311e20907844b0e591c54c10e6d2099f52488f7a00bfb56320
zb89cf9febae3129f2969bb3c07f7054f402ff143290fc169108fb87ae608d511d25c4ce366f0be
zfaa03428c923e96957db4cbc7e567e09ba15a20021f6c394236f5ca0bd1385fc2f83185eda8146
z059d51cde9114314f9424a3ecca384eb4737061380a5de4156a426263874a6ce598ed763526566
zf2459395607c43469378cdfd3b34454715f4dc666960dda25d224ddc2f07b21f2aa1b800333817
z84b886fee9ee4d18db0f2daa8e0aba997bc58c0621b0f04c528786e840a8b7865db79481838fe8
za0ff290a0d95ddb9f331872ba0ff7df5828e797f1caf3a047628d4bc9429fb223fa48151181479
z05640bc13e2c57e85d28a1b7f75f45115ccfbfda2b84656b21be7010393053def4857b1f1574bd
zdc259196c6c89f9ce5a786bf3831b2efee2ee378b91bcdef249c05dd102f29dcf890c88d56f679
z842f493f0b486ff0acf631f845b6f76bb6439ab5e3a3cc541dfd575e67afa46e4352c66556d6b2
zeef3b46afca316d07bc0f6a89c9f6a9f81d501bb999620de8cf459db62532a0508b632c43f917f
zdf425a2544d228f357b147ce899722ec8287be20a990c813b7145c9236c418bcbc942444e8ff1b
z639ccbd5b90c1f44d40a91f58c4904cfb29fe64b3dbe55a95f53725433163338b92ca7abd9410c
zc0de82d7358b50edd8579666bcef17cf193f8725601107e21c0c38933e502878d7bae0eb5fb1dc
zf19d7ccddab4b186be08f39dd1ba80397864dd9f0c78eae2c01afc1c276e02ea1d5c88bbc31f9f
ze8897df5ecc1e0ace1b8462536fea8bdf44b7cc1f59cebf8c31e02c2d0265a9f60c356d7393206
z1b046efafcf4bca8b37cbbc51c8fdcdcfecd379a3f95ebb9bec04b2c73d8e6270f96c7215b2309
z4db7464ec1daf0c619294a8b5ccd5eca294dba09a0005c5a4ddee15d4147da3bc935fcb3db5819
z1813158b73bd5310a8715f654eaaf042710818c55c691b577926e3fd55daa1c3ab6ec38df3ce4c
z09c47558124e23e62c49786147d073755ba7181899b1a28ad60867cf7bd0a7e806c37a742e9d1d
zdad4083c86029a31709243981df0637f71524d30cb31506a2ce948414ab3329d4329212607d402
z659476163e256030fbe2111c64058d667c003390986c546cebedfec5f681cd7c054cac67846359
z40af7574e8782ed949e6deda1225b99449c0324d6cfccd72d25d9a1d03ff7f95a37cef8745e567
za602f3ad2b2263c55fc8fb98af9cfbd97e91cf6cfad028a0abb6953918aa209de8b2433e6a271d
za92e84fbbd364c81e01f5cff3c2468a0cf7a7ae666956f44f0153613c9b94b820a87e95066c861
z5e9c1c6a141a28d6fd6df40803efd188936bb933bc0c32eb3b329e07753dfae29d43b57a8e36c0
zfb1fa1c3b2016217fa5fcdb76f41ca8b18f51b017d19cc9fa4544952dbf3d089ec7a2e4c2ad765
z6f4c8eec53e912bfcdcd64f10a569238d68252aced39a125d0bdd322723862dd2906bd8be2ae68
z39d4ae10f93514e5d4e38a7ccb55462bd41e63d3e77c646c228437843ce6f4de371150c26c6015
z4db4f3d0a72b30901d0c465e518af0cd66b81a3194b7e30ccd53ded5daff715731b2844fd6db7c
z984d2b5a3d8def4e461b9dbc0263cfe4f6461c211503df2238329d1251c6131459691872f57a07
za1ff0232f21dc063192a11d585083630bf28e1932eb98c2270fd7260c79978504007b3e5411f2f
zf05e95e8949af5886e40bd757e1b548f348556d0ccd11864554083b6b7b1001a89f7c916f418df
z8e159e41a2718239309ac3aab93a551fd562a140738237ec67336215cff89ac0224d79b09e57e2
z841657df7f0e55e3da5a2aaa2e269f81bbe67273b43376711b5c02332184783d89a1167af19d79
z4e137d8412fe08c143459b9a54e80047a934061d84803a272d8e6d38492a07bceb3a7121626eba
z65b65d7dc8b2acd1c147f91379d455a2d830a540237dbcd857542106c66e216427b762d6e1be70
zdaccc4754ef5aa5fa3fcfb943fa5e8d5bbe7e9f88c12fd62da8a0c903e5bd62328a05356a596ba
za450d0b9b715e3de166b0a2eb11846a4b160ccab35f873bd4cf75da9e7f2eac901a36a6e0115b3
zc81a0b2baff3ef31ce1e6a42edf0814ab765aa50e9e81f6185659c5b5225e1a34e47ca63412ec3
zd3828aea76aa618d7ce98e9e9b8a930cac2dba2a931f6aeb9cf13826c0466d990761e8bfded4d6
z12952c451db865f0e8389823ae0216caaa7bc16f4645b58f75f965a8720a475b94cb5d7156cb86
zeb5553b178b35f8b8940feeb38a95d83a3fa0a28c8229c6954314a93c39ff217f39d9a7b1d5a6d
zde36dbedf0c28003a36ccfa4897b08f12e718b01299c06c833e3dac68551b3464d2df776073a7f
zb623d8b0c72c7c9c3a396d29229818c44f17ea94c15677d9cb4ecb8ccc95194bdb8e353937cd90
z4bc067214bd7473f4955028322fff731c427722092560c3b172a6ca32a55738a756cadd0c28c4c
z776897b12aca0084f1ee6f70322088d1d7eabf69fd13d15a48393ada63a7733d97acd62b14bec9
zdbad199268831640f3a62ab6945c0405997528d3437a9499c736d6910965e3c3db95f32a55c028
z52460d2f1de6531eb0311036de53c66906e938f7b091977aeccd8050ee4f73d6ad34ae4c093a23
z5a947790823cb2a2332e772b7e845964118f593dbcfb60dc609ab05e781b63db4dc47890c22e80
zdefaef488def22a36500f745529d4fa551d8a9d689930c7b21fb9fdcb849df0ea2bcab8dfabd60
z46fc7a0449d00ee397c7fa1da1c57ca96343d2c9551eb789f076d1cb98d78de1ee8d108d7eb520
zc3b1c4737e366e5f2bb60db436cd52c0401c92b27c77235e97ac85a7eb28bc3569a609135fb49c
z4f3863c1b58267d180a8f2a6635018ecb7a7aac2b7c1d12d762bc775e26095220333a6aab75663
z53a23fe6d6d293920d847a3c418c21043f4260db10ef82930cd22337eaec5e8e9a833712e5dc3f
zfcd59616ef131852c4f985be262d6234841e009c46f9f19fcc2be36c5be6ea39ec28b7f1208d6e
zfb4ef5a57a470249d04723d7844c17e59f68fa2925e34f74f0a1810f02175912019747e56e0392
z97c1adb9fa8199836af05fb48394914a1af26bdad824fd205ba4a1ff335b9f7f89fd6da5e70c64
zabc363933400231b0e495263cc88035c3c92af1138b61bd3952956c30d1ee6a53264396fbb6da0
z1d2c9241a8a74b0fb78c86f056cf039714ceb2a3988c51a31965939708385bf73c4fd4e5890aae
z49b4fc406823ccfcf5f03e7a78d256573919855df0dfbb0c517f51971f125c92ec00bd6fdb182f
zbec6ab66e20902718fc3da8024732baa3cc28f5434841a688f8f632cb15038783b3a513e02f5c0
zc10e2d2c477b0cda86f7e6fdefd36e1a276e9b449db50f893468594f365bf44b1f3b08ca69496c
z26f7505cffbcc14443d9acc1c4c9daa7df63e0309205b567664e06654fc6a2908f90ffb8f78e13
z73535c649702cfbc862d6d91654740267a61e3905544f16ba9b6549a3f3a8d33da9615918e5b70
zf4245fa3111db141af9aa89174fea3767b92dae73dd55dd4c1538d5cf20e6a432bef1e57273f75
ze9185a37fdcfe75c67bc52a7e1121822043315d99d0d54b91f07c45e00eeda63e95556f0015f44
zbbf0bea780db54d761c26f0be2942aa93c4d43ad895e6c45bef15aeab37cc0f69832719c8a6430
z7ad246241560839dfbcdf2e684e58593d521abf55116b7a415d8532e5b097677fd9bda382fe112
z62ada6dece8b1702029e9823b2072024e0ef5e23b264eae4185bb3e70cc9f36536ffe35eccde64
z629100255fd14d69ea4f7d7dc2bc5fe2a1a5d944c92ac39bfa5aa7bad825ec3a1403a4b9c6f57b
za4dd209d23a5d5e6e1ae03f1a7afc562d74020d3b5f846927393882f6d889a8d12d6e6b4c03796
zaf8efddcda5cd1046b51ce2a4dd2739fea8b4242cde195f51c0af685cceae15dfdf508ef196c6a
z978d7266f955dc58c49745166c6361ae7540a18033f064d761f0b4228d1ee2e7ed7f26bbc1ab13
z90ab07332ca92a7afe1820a18110efebf5fd5972efe531fc8ce8c28218d34f4fe0892c68006fca
z3d9022c5a0381bf338e5abc1479aa8db351afdfe89396688d7ccf9b2be9dcc31d1be8f603b68d6
z927aa4db06d41d95a71ffbbbfdddceca72525c833d2358edae3153fd2f69349aa0f1b89a6aaa67
z1b8603e409c6012ccb6d32ca7026d00eeab2a0bcc916c229c0b821185931e3a44a26c46fef748a
z0d7d6c147a4a750ac688849e5d6c7b06b842420c484c678dd8c28fae60edf6b1799012447b00ed
z6819547090ad22d29ebf6ec197b850b4aaac9538ad77da42fae094dfcfd0900ee40862f9ddc490
z77228f591da81b723653b402af58d3989585be10e25925945a6d917d70df47e4fa4f994ee635c6
z52308e5af9fe5de0c53feef08466de1517bd4e48e5e9adbe48cee27c48cb7f9e9405fc2ef11f4b
zfd090a2bcfe28f9189d9dc07a7ad43352ddbd4905f7fb8ef70e3a4dcadef478104526cbb261963
z8ba801409e902bce47014b86ebe52773e59a2e78b8074709e106cf40ee2fc4736835c3b0d1830f
z6dcc8bca7e82d75ebee5320a290346424c95a27ae2c86f30e63f5532b7d64d80b172483784fde9
zb24081f63abf71d71560ee8092be7c04f30782cb14c054076364e5bc3e59e63f0387846f9c69d3
z0d8d21f23ee7b531df79ce0f6c6c96f622da0328d004eb177a7a0095ed56a56a089684090325f4
z57df4da525e6dc89e9c3d5e30b6582b4a0131b2feb008f7f2222590ad1cff5577b46b20cddae64
z8da60790122ed811a8e6c8d3be419b00c71fccb6c64c63899b7385ec491ce8a96d3be4b952097c
zd43ae5a27124b8fce016a6517bc298d7ceae4284f3b28c66c53ebf78f03d7d0b39cee42e6e77da
zea8be028a08248842e750284d21d3d436fb6081a6ab19b4fcafd04c6ccfdb2e7e55ae1b224d4b9
z5b99750496e3f0e292379beeee36ca300d14916922dd839e8a2c7d107b6687ce4604baec237e37
z34d5f6b22f252f45dd4279ddaed7aad6583da53edf5796682a1515030d4b8b14b077b542eadb9d
z4e4e67ddf760d3061e95d4af2c5f234542864728807861ea47bc8292ebab7857e5ad844d2ea029
zb9f46004e65efd75315953b6975efe96d7afbc73608a7f1ddc6151b75d081e2bfd012f80ceb5c2
zc566b722d49ec2bcc25692e89475f9f62dc8da82062dd9c5524153c84edb999d5641d15f44913e
z69db6466e61c80df7760219b49ac018edb07f9a4cc57801170d84e1294eed7185250700e8af5fa
z4cfdb9ba31ea4a6b6be6dbb0006df3363e6428e47d326eb3cbdcfc204141d415ea5a9cb3cc6ad6
z7e310e7268df92843d44501a1ffde02c8fbaa02400c2ef0d562995f424027aa72eec3b57b5e322
z14d062b38a10f990d59f22ce27e6a7e0d9692f1a9eb7430f52ad0c170ef00c830edc9d0f47860e
zfb282b1c366fea22223326129bcd99cd3365004717a0cd8f6e51431be210081cc3520ac71589e4
z9e9547b718a8c6cc940bb0d626d471ef955c7f2957b849954d0c00f8b93b2e12f235d5c9d0efa3
z4e3a6d5fbb8a53c71bb4ac18ec17856f449a76c1010e1e883a3bec8bf8865f338b7e3670ee0e43
z4829c8325f5207ff99d49d11a6da891f934d83e06a627e6e1db996f742b14e1730c1585dc3b0c9
z13d92f544faba0038cc1bfa9dfeca97a0b5eb9833b436785671fd00031d71f7539ae2a631c3187
z5aa8c7dd658324380959c61c24d3944831e44fe47aed653962dea270b7e0b36f654b183c4fa493
zb00e1aef0d16b219827108f7a03d2d27c5ad896c3ee3ab10ee6cc728141947b25d9f90d531d587
z5885fe716659c8d8025e88b095ee4f80a2dd8752006198c46bf8b3677f94705dd0ba51e3a91e6b
zc4c43b891ccb41874fbedbf61d4b6ea02b1a7861d8ef65adfa4514a0f64c24f65b117648d97747
z4bd54026a0f6c849ce17a99c961ca85c9d667163064afbe1f1745835d225ba136ea023d53b8cd3
ze47a13b865eb0c9a6642095188f185a7db15a5576c9ccbaa91050ea567b8323f1f553ddf6a7dca
za2534fd67fe388f82b9d1faeb6fd5c589f8559bcca0d3a6b4c86e9ecc23a5778562d15faf0bbc6
z6eb41dbe8aac19c36202607002ca4303d9566b0808df73c8ef7866f9d240a2d62e014b64c87ac8
zd6d1826248d27ab11c2eaa4d7fdcf22b9b2079db54a32c34c6991b830fd4eb39f63c9396d81848
zde2df51eea8246c1a643258da556ae578891e9c3b066d3f3080772d22cc036e9c4bd2a4e2b12bf
z61b48d39c1fef6407f06abc4f99dc70dc4f022c9873662b98c3ba1dff7c217859800dd733f9286
zc9a3fd8d0b7b499792006ad7eaf99bc8302d8a26bb5a494d094a601a0ad02f7e4f8099fa0c9fb0
z14a043a355a07de3f2d7af5536707e9db9e6e07cfd511c25f8f88a629a95b354db57cc9c4f0cd8
za05a51851d1d4959a912c47b2e2ac08b62ff75d5cc11a8acc16375b0607a58a41950e7ccb5879b
zb871149ee415b8b17bb27ccb7796f0a6b2f4cc41d74b4807469e1eda4a6487595b2dfa1d7d9200
z7d145feb476965cadd41db2b1f1032a7f159a4e44864b2f0d10827446cdb2faa9de674021ac9cf
za6a4aefc2f8b8c48871e29b634bd8d79769fc28955e994947c0bde7a7bee5a9dda1a72be3e1005
z298ed425d017d4fdbc9d5fce1bf2b72333623728b2effd29850ae45f6c1b2673eed966c61ec1c6
zbbb5449832237dfc19c9401a9396872fe979ce8f33956b82c9c2b3d0f563b313b579313e2729ec
z374e4d3cb1db86be28a2b989a45c7079682178df4695d9d46a4b20bd183cd5de28fd9e479a9cbe
z828ecac7a57fec4360832cc54b6b864e589278629ee7ebf1f67c40d4574ad0a557c427a77ac0eb
zd34fde3cedccfae9dd34edc0bac77b60595c1c2f70efbe690e4386d97309d392b1035df97a431a
z9c0399d2481b5893ad7c22e60538ebda9a9e362f5e044dfe99828819c6c4d8a049ff105c8b568b
z26743afc6f925f7fc5cde865c5ec41cc47878603d2842af5def6a5cd455197d9fd375f8c04fc03
z2b4aa07172bbdecf5cf840af7bbff13c09d92c76d2c85f6c836455f6df66aac0a74bf5c568be58
z3baf0ca684799b2ae2bcdbad507d299854034d5a73a375873972737c897a497ce9e2d53b7f5140
zada1ea74538f4c842a8116389973f4ec201975ad310f33045e84c798191994f3a0c87bbf957077
z39b1b2dca626d39bb3784a37c983c70b9bdee2a22ddd6e77a9b690ede171a06fb281612183f3ff
zf188e395a51d6aa598646fbb7a8db881bb98a0f7f6a8fb8005ac94fb3dde9c270d94e4c8b009b7
zf7cfca758a199a70dbad8cb7fc277856f436b9571fb31989bd642024e7e533653ea89c1b117e61
z279393c651579410f43cb41fc569b58131808f90edc509c3b7351707d489966dd0c34c49a73bff
z16d4b4f5e8cc4d4cea583353b3b1067936d45a4d804f969ac9d3f9517bbe7d348399c34ac9d3cc
zee73d52704abe95688d7e78992e3d3867adb7a5cd6b7f2d6336b4f851d08595bd7c99f66f47762
z44f4004045ee393fae5563f6847870a1cc459cb8f38c803d9bc191e34a3674b45bd44d95458294
z1508c47be193463c33bbc7126c1dbd4725e1d3f045deabdfad4d125f1b397d8957305af0a0666d
z3c60127905ddd4f7965a0cb889db6be02a7b8b73c3b4d567013a37afbfe285ab2ab17d5e57ac69
z004ffaf886541c6feb920f073a99b7751eab846169283557999c3b7b5892126a23160cf5b9b918
z1c6c3c909ba47454593d7ace93561ff9b7a0c1a5f973b48e7a50f1f1bb5730593fe48967aa2f31
z069d50d3770dde96a3b7d6c9d359fb010f1ea568703628a3d87b65d5f0f35fa37b4dca598041dc
z6bed73d0f40660bcaa7b5ce6fd5eb7df8446c8ed7712ff194038d6a15f5c3db276157f4a493ca5
z30fd15aad4cf9b19319ea5dfab51516c8f600fbc00b658d74b4aa7b31c5239a267401c7c8a92ec
z7947e05e200198d7afe245918e727988ae402dc5d9ade50c8fb66bf9f036f7d5dc3cda665a207d
z4d43c8b56a345d86584ad4a776ef6201ccdc8111c524e92877f4948da6b80a050e95cad5155e25
zb5d40835543ea434544a106f088fa2fd54445c95e78ce4f96b25183cddcaa6b7423413c5820a43
z841b8443ebfa2587155a6e925aa5e75e7ec6e71b2af285c1d35f0c7da084ea016aec0bf17cffd0
z51e7797c372971ed2f17859d7194934fb3c9f6e7df16e81b367f5b317a26dad6741d0d7f515c6e
ze3ab5c3aa584639ad9ec74159094d60cf75eb3b4b3df1a2df10d8163ebf2c1e1aa786a583b1daa
z3b8e47b9ed82abe76403acbd154a73b9257babaf699879819f8eea9a7b78a1003487f53e638a64
z287b28c7643e7a995bb7a381141e8d675350aad6e069a0e5ccb65fa5b1b34ad73ee2def729040f
zce5c920b4fda1879b738f626f63704e45530559213b0adca371aed59c625cfa2558a412284edda
z50873634c51617e40ca5519716e26b16cb253c907d9590df3a30bf7572391401c07ae76402cd1d
zee1dd52d4aef8541e493d12895829e19ff97a38be42cd971e388a53fde1bd1965e59fac5022a4a
z4d12afbbfa5724a3ffdc6ef17d2008b3fd476b9f126a632847d3ce1215105a083f6f1d18e1e191
z98eadc066e8e773aba3677c2b75f28015bdc64f2cf8f8746327fa105b30b569315b80b273cb270
z1b93c03decd347fafe2aa304233fc695503a9cab454d5532e90879209a4224fb0f57e85eb70332
zf493be9bdb2af8296b7a932c0310faab250c099aff499adb18f5315be1a60299a5f35abab94ecb
z712f0780c5f2aad0b590a7851e1432dc804f68cbde04879252867b0841b577165f76388cfcfc0f
z4e1813d08fed8442775d4362f1436aa6409ef5120476b29b8c98b863821a89da07c5a6a74562c7
zafc1713f860e198edd991b585d60a1294d7d911cc9627612d9d42bb444344d53c89ab20db64833
z6a738d3ff5b3ea397ab2fc1e94c503e4e138a908be2aff0b09e63021054711461ab441873eef5a
zd4003497619a9f41c2f964fb33dbdec5cc6d817e6528321ffba9b4583b126859bb5d17b43d7835
zb35fbff8cb1af6a90f152b5ae01563e535e6937cc989b07e07de98140a05c1ea2d35de6a5ed1cf
z69161eb8e75fc9fd233e12bb4a44938970a9998848baaf695f2e7bb6bd1866191723329e639109
z945e3d54d07b737e368d467acb57459af081e61461c8def6a879191f5958e955b4cd91333b4d7e
z0f67db56c80440f994fc34c252806e410fc5f6d1be1e1cd070513a55b47d06716d70fd4d7c878a
z227716b467d08d04c2ef075e56541777d56859ae45f3a1e10b4b587a327608ca855551b5ac3d34
z0a7b606bb8563b6ff61e383d9297c39960e54c6a8e52f34ee1f2f08d68846194a452700f5701b1
z6f8cb19ebb3ccfe9bc683ed15e0202daddfff0e9b139c6ea51319fd41caad4ae2baf4ce7a4ebf9
zcea52e15f3cea83366daf0d2f8d7f93365f868fc7673c1e3f129f13ba262a41a9e41bac8e5a540
zeb5c8d3f06bbc4c755c9f74c1613ef65728fc69efeecdd1cdc5bfd0accb724beeaacb94f1fbe3b
z2c6c9cbf4f2a86402a3576d4f91b2ed240f8dce08b9ff7652056f0d742460c9e6f05592b5060d0
z4b4caa643c34a1f494b706b58f52c5db5e373858de870a6ce39db0df43f64d0091ccda6159f9fe
z379598ef5e4634cc21a33acd3fec176fb4104b07b6523a74b6fdfdeaf68b0100a981ef5bfdb15a
zaee4d4f5b58f46e7ad7b1963a206d8686e65dfb48ce557d1c0b82a052d1aa6d43a013c39e4672a
zd61b849926c1298c0336171765fdee0a1281ebb9c7b261aad0ae943f4a5e78a670a99ea2c301e5
zbadf4ecae12ed393c5cefd22a6116e62e4d34bffd90cc455bf6d7fb120ec6836bf158a03dde626
z87eb49730bb44e878823f2ed1332ebc4e8f115b0e6e4d5858fe74a90ab8f81b3a6c636853ab68d
z3ead559d16d458e476b50625aa773d4e8b08416d87d55ea156376dfb4dc84b4140287bf509bb0f
za56f4f3b1662b7d119cf0882098b346416226dc82b97a33a7d10ff2bb4cf4b62887f329ddfeff4
zf629f33509ccc184c760b35da91fb697eb82cba9f169f50a6884d5d90c6592bab0278692095549
z1dd93c85fb39ebe64759e35ae2b4ad017171e63c445e3cf95800ef3b567e857769e8b195b0471c
z85dac4b94841331b79fb5f058060d70d9dbb63ce350bf1fd38403e5f501004e5f19a69c73d85ae
z94d0d73cfd4c15340e84190fa452ede782a21716a73396c66e8534d3d75a8be4e71f098704a2cb
z5f2c2b607d59b8801ced565c053772b6580a53fdb95ffa5eb308325ee86b76e6bd892aa5a861c9
z84b3c71dbd29ccb7967a5415988ef93f3e85b4e3f13cd9ba317d40854263c17bc7f1d5f43e6e9e
zdd5aee74aafed561c6f8f2ab60607342568628a0efe113e49ee7b2b0e1899b2a44ea49f1904fac
z6abb40db38851b568b700a5ebc6f5187640236c709c91c48731f379ca826285feb697325b22049
ze84cf9ef6be1b8ead34d4e5e6134a86acc853def8c554ac86b6dba6824935d1c3dd19e033cad50
zd5753545e8af7efa5f90cb5c5c0fd84d63c9a8858cf1efef98d2167997931ca189ab8ea76465f6
z6ced2f91a3284af8c78ede8544e22199c92c676b5cdd0ef93f69bc12a4da093472ec57a5b29849
zb7863ded380c852d401f19e3f3b38de74d3e76368a065b021cabe003460a3bd97b0251df063563
z4b11e8a1631b5cbc333f664b5c2c7609657b03896f55e0f9e659a74514806a1732330e250fcd1d
z6647e6eca2bcc8c179c41e3b20ba6c25abeef0f0d05522005b970b7752a05cbd91b53023e00a43
za23e2b87e2eaf782669212057ce34e11effabe591f500e5811e692c136d5f245662f88996aadd4
z5734edbe41cdd4e5bd8bf03c86a83179ddc738c84feca6a440dc0d6101d11ff21acc307084b62d
z7d20d8d8eb65e1fda36efeab72e630d7e64dd5e5de56c1ff6deef851b57356e6ad2c9cd9224007
zc94e6fa225130013e52aca968bf08890b9c6b35e00f074fd5b67e41d3db3ce0104b20c56d043d6
zab8b17c1e124cf4ee7f3a2ac82af2aadbeadedcf69097d063c81baef61b8d9c576e224ea2a274a
zfd3783a26b0b47daa0f31a06e20160c4d6e4110d1a24c9936b435a7b114fef5de5fe36c7e43b4f
z87cd4e207dfd376b147c86131c519d86ecd7c0fbedc296e65624f87cc356f8b0d82154b0e4e802
z40a6ae3fe0c0faa37bd76afb266722761c9d260084e0ac6fd28b397ec9768afd40b423dcac3aec
z275ec0675618f81e91452eb4db3cc2fec94976b170b6c999ad5303969c14b792b217ff5131ab11
z5f58b0dd09fb14d24b8cbd37e123001472f379a09219c6298358aafb842a93dbae48bcc87d04d0
z3eb8f8945832e5b4f555aec840ad27c30be42623982d9c68fe27f21adc8d74d569b55d4913fd6e
z3aaa9288bd571d8a83273f9fa8d3b65927499017061862b6cc249560394291c3893bd36d38f0bc
z3162f54e7bebc47e2e3bb622bc976c450bf40a244eea2902795220133d02c41bba8f64ee60d34b
z30542d09dd82c45d72e544b3bc538cdb6189c1a0c48eba9ef28b00ebe9d53e12da49e6ff450679
z9322412ecb67a348bf142576024a14ca1b4a96a6c0865b2b5e1e1204f663df3da3f2122055cefa
z8b2350b6d5eb40485cee14a66e1f1047924f2cef087d8938cf64c97cc255488945947bff31bb33
z705b98025a03650ff75ea9493ad62807343c0762fa152375a526022a3a5e2413cc2e180fac49b1
z0951e2a2b7fb6bfd4e90de5dfed5ead277a308b6b5588a313b8c080667f9541e318a46c7ac7220
z59227b59bb91817d6faa9c10bb2d741f7175d90c99b6d5b3579af84855dfafefc026d454530a56
z530c0e5a9034f30cec0004898eded8009e010137e9fc98a81808ee5dfb64a7398dfd5cf491ba66
zbf242dd9e052879470c3599696b8f9bb62b892154ea0a7e87f0950d1b265a8e1f2f9c807123f7b
z1d691d5c6d519fda7f15a4d04d0b36e284eecfb47a207086a89e653d297e7d10e659e29188b17c
z20bc361bdde4f2e035cdf004315da9c16853606a7e886943a3cc779d46cb55ed301ea4d1d262e0
zec9407df6b58d6e976d6d190f2a50bee022d3a0b1fdcfb97440247c136b5d565198cd45c58291b
z012230c9acb6b95b6c7f3cc0d1e630f5cde56c3cb5cd19333a51b0e4a456695a9d1942895d854b
z9a3c733ba1c63efc19fc941b0dbc865e0ee369588dabe26089f8a8d33f11fa7beac3e53808eb11
z39de4d88f3e72895aa9650c492c196379c37affcaad54e1eba40e305dec1e23a8d2e5c7203b8b3
zf1cf24ca65332d8a63f59c48ea4d08aef8f7a5c27df519222a9d0e849f74f99bfe9a3d8eaad985
z96c4f89454f18f5212efcca2c4ab68898004c3abf34f4f89cefc7b6f4eed97224b8fe648497ef2
zd4d03debaf14f03c5b4c843abac6f1559a3fce5702e6538eeae01bd6e74a8740089d1c26282706
z39a6a4263d56f55e153de4fff0580488144e958f216c09b09bcabd4ac772ec7caeaab81a133ad7
z11ac0d7753df1ae269cade158f2769efa56110d28cef424f680bcc6603763e81dfa81458fa6c27
zed3fa7549f3c86371472aa6e0380998063200c5ca68211f39b02ac8bd9337c0250bbbc6f4732c3
za88ac1e12a3ea3886f927f441a3a851bc65fba9cb38ee825c7ed0f00f66cf2f0f636bb50b02a12
z2f5d768510abf7d4271b799e57908296a5f26c01423b78a78284d1e48235ce252b10845d40369d
za0e2ff6b3b443b9d73458cbd53f7bcb18d21cb4dfa91c9ad5e130ba50e6f6e0af698768490b5ad
z05e00318051db364f72b688539c39289193382419073dd2860c37be93f3badd45750411da9715e
zf0b28ace91ec680f9d47b55de071f3ff0da2b3d4c903e5e20baf83369e978b00c6fe400497785d
z3354cba2d3d167f0965d15ca34cc0b8ef5faa53df4cb98ad229ce7a845929a736600e17e70cf6a
za27b70cb874351b902aa869aa8c4e9498b67349870aec6d4e3f65840fd0ccb8af078a4a3bdf602
z0a58c42935b68d3c718cc23fe37a99f6bf9f2f63b02a2bd42022e63d7a97acc35d2955f799d1c9
z3356c0e7bfa4fe794e4019e71671b914ba13d1c56714f251a26126fa86e766da310dde07880aa0
z226be2ed332704967664b6fa8b47d960b60421d5c677e055488589366979a38fe7ea58d9e544b2
zaef99278741233f7dd2181103c7b716bd93b462831ae700439b7387578578fb665657cbc849a9b
zb4b0bf444f0a65d49cb98278bbbc844b7a5303fbcab439c0944b6d67b939dee0a3e51f03f62e64
z8e377f0bc8ae418de3140f22ae07142101c83a8f5ef2f426be097854c3123faed283c1936862a7
zf1091ce2d9d24d512756959b9142737c702838218b1321d61195dc75eb97c3342113a21e7a3ece
z274dd1dc36e133d9d1f2d4704c3799d2b732525b01212e259d6e65334173be763e361868fac240
zfabc9769008c3381cde4faffc93ab1008452218059901774957236f6663ccf4cb207cd794638d5
zd40bdf18e7cb82803de70ff84e758728144df0420cd46ee4bb5cee0c21c13921b90a7cc2c4a3b4
z97638eb0ec459d9248888a211a363774f025b3c8ce3fa8a8c60c4ca9cb20a90dc29d864a8d52a6
za48dfe70a7d4afd09f4f7eccafb965b13517ca15d812b4a581189ab543da849da342af9882b8f0
z502f325ca89d1c466b8667ded1d5c4412553718d3070d516bcaf4e6e7c0b29669e0f8d8fa91a44
z40b2578e16c48b15c2ebcc8811ba526ad78e85208d618380951596e3fa481cad70a9c9b08f6754
z5e2affa9faa3d814ed0ba1b24f37257c3fbcc82776dd7a405e2290337a9c66e2c6b81096265acc
zc87a576227342b4e98dc72724892bad9ac9892b6d87778996b2ddd4f0aefec4e6318b11108903f
zf9614ab8149bd23656c6691fda9462904516b1cbd0018b35ca687a8896739d68b97b3c0cf4f3a6
z45ae64bc7c4211c41b33a7ceb2d2cf3ae7f4864c318b77c71904da83228e6de961e6c5df4f209a
z9ee0d4c2eec3445a18061dea4a5942c62386879d3c97cf4c1bd6bbe390b37079b1d8d98ad59ea2
z99f5a7bc10cf21f3d73bc53f27c9f065269429f0245d1b7fd848ac31ab71095003947ba8204e38
z58408bd5641c3f72ba4305192671b10336720c1d62e4bef846fa399169c534b81eb76c7b5d67ba
z989b80ef1fe72fef5d381182b2e5a25d3a02c57605e7cc19b92ff2ed7733c850ebf1f0702f793c
z2a0fbe090a626a08ee358d96a81c27aff1ae8dfa0fc8508e9173d2351ce85f8d1a9522b7d5fc7a
zbafaaf686a99428c6a842bb7b25227d6f610cd559cfea9e51a8315421bc24803e8519e005a06cc
z6b75ed836697688ebe11becdd6352cb9505be23dd5ae9a647f9491d0528ca26f6bfb1945b7c418
z21c1baa7d52d4be7e1745accb3b3cb7c7b485980b5bbf503b2109f38718a2814898d4761027422
z97c73460da228c2eb215465cc1e32fa0892b0c39e9ff30e37fa269255f1f0da5249486cb4d3dd7
z780894846c6564d9ab60d5164c4a653b31ceb1801b9b4b09349d1d1a2a722a7a46986d1f906066
z33e3895de98b9452f9b2e8e200d9b712b7fe507e80a03f93e761aca1d7965f847b7e46da22aaef
zc1799569fc61406a8a47049ddd1bf3fd0af06b6560f9ed581941534a2f8bd66fd659b15a435046
z52f9c61587b4c9e49577c16e911773beb473ea02d7a6e2abdadebee25f24e39b01cc84789355a4
zc6e57e4794dc757c45d7aeabfafc4785c25de64ef7da7fa76cce512d1efbd348aa417695586c3e
z584a5cc087b314bb43f4d7f8ae9c8270a7ebd6f8cd341f3dfa99078412509eb3c65db0d2553d37
z1a645979910e763009a54747823d04386b040f83121176c53819eda704e1d89a339212f09c9a95
zc6dcc39c91ac739c0da522954e77ebf2d3e6abdc55798a7dd16a512f138fdae996b8e3db5c15dd
z965de8383fd57f2a9dc721c16127c35fe1642d3974ecd3772a1f96240154e56f41b13c983a8cd0
zbe335f7b1edd7130ca953e0fb88557debb4d8ae1708af448e135cf554f4b7a2ed30dbd7e4dfbc6
z8b64d3c93b60e819a142b64039e0d27c0572d8e519e75042905eafe237fde585de2adf2434d9ce
z1355599292360f8f79ce321e9346f3d4581b71a13a33c469102c433cb23347e4f09c2004cc30ba
z4cf9dbec0d8653b1545146c964db3e0ae5610db767a4d299e08b27a51d0bf05de5a597469d04a4
z7463ba3b6a6a15f730bab67fe9030e5baadb0c3d26ec92ad8579ebe13a5a0945cc3476df26a697
zb039155077dc5fdc67db0a53cb055bf0384a0dea896f82c6a36f568e2922ebe18ddfae5c264df0
z8eb23ac087ab88ee3da4c5f040f62c1f96b42e34d8b4a23aae610b3b5e3c35b9b558051829779c
zd28be13f8b1893e4104d48fcc0abebf48e6f0557ee30c6a1884a2fb3dbbfec18af88886164b6f7
zf8466ced539e6c4617fe5f8b174d4a229198f5d47d847960dc680ceeeea0c4800f9c866f1c7fec
z253bac254b710bb99b55a88a23ecef7dc287dbc1994a5d4f2e6d5cb32ab90d21f2e3cc51387f96
z6be66b4c31729159c482b1a0410008d96963b659f7271c3f89a5533d19a60137c5daf27a06f256
z9ae482a211f56ed086fad2f6f5b7a5e89fbef69d41c500f65d21bc04c82b56e8ac6764f9ff1a5b
ze6d8a85bafc3cf2c34433eacdcb9372121e0bb12e36c2736ce32a9ee7c4a10ab18d7960d3c4a0c
z32d8cfa7de06ba2f3f4b80e4eb3cb723de7ddd4b2612ae398fd9b076e5c5864d8c0c80083b9cec
zc91852f6bfcf076a9345f23627e237e95af3e56c7b45fef1383f593a83b28d9d07d12eb908bc47
z7a62f7a41b410dd61c4ce2a7c08036c40991570f047ca0c48167ac2d0755f6873ad5e3ed64881e
zd3eabd1c39f735fe6e24e9d552efd8585a7ab0af9391b6026e3a89f061b342d8549cdc6f458464
zf24a36d0709aba0279511d99b860c311c0166a04eb387554c50d095c9a44998496c6bea1ba15e3
z3124172adf8ef74ddbb4714ce3533c74cc7c9c0189d03a03247beac1bc308c901f5de0afbe43a3
z74c87541032636dadfe496328c03132f82bc8e083c64318ead99e23899c093e6abd9e733ff5d0e
z4111b0639387fb94bc4d14a654f96b5deb9a0099bfe99d86da4b0a610987f3479f385515ea0a0f
z362a43a7621fb92ed2d985adb47884041db1d42d1656f719e72ac4d1ffb514ba704153e638212b
zddf4b0d22b942a3ec0ca233ba9fb203c495cd908adc050de2c0da80782540a7bb72ecc37e77b3e
zcd2d295839773f09cc170f2f2081f323ce6f4dc48e6942e4488e8f7d9f5e04a02deaaa04a7b475
zbd60caa088471ea7d5076689dbb86b189f4c05e69ebc6a392bc461d7758f100995a57a530cc9ad
z4c4c971349c2b5bb8fcbdffd473cad0832f193cbee3d921aff128abdc17b35fe796b9dead05972
z8a90a88e3865c8aec2e4cb7d940b5ea22b8144da85dc76c5e8e102e74c6092aa53dfc2f869b59f
zbcb187facd8f603678e3e97ee64c0df26eef962edfad38807593da6a2b3c9826a58759746b792b
z95c342fd737c79a2a5eb172cac61d246a3517317a62a5f87f617351a687291cbfec5abf54b5075
z094f15c5a150a14164f06c4cae2170a657d560f0e85b18768a46051b0858260f129d0ff64f60ca
zde1cdeb8887f074a1512ecdc5e44f93e61e23ab95034bf057274849af8f9e64bbd7c3bb09969eb
z13d263cfdb51c48cc8a41dcb8e283d4674fffe2386be8cc4cda5b927f04a105869ed278e81997c
z25f3eee62effd16ec304cb3e8f8f4ad219044dd2597a5d93797c3d17d241a38fda3a462af1c3cd
ze4e2f69601071554638a015ccfbe98a77c4afae6e581c1b9b7068ab16145a9d821f80411376533
z7f81c005f223d96f5c6d75a3484cceceab06d7964977369424ef1779ec13d379f73269fc90d8b9
z88b70df37f2023808d76e28a48fe9c2836f7a9a5e961630e9edee34ddd11a877a5ab1509aa276a
z2455dd85d42299c1456878d3ad611c0eb2a7d59cf0ea2a5aa3170f8f09a80bca4237245a645987
zacc6599db7d1e560f009a8cddfdff9c22d08b6e9f175164255815615e2911693bff0a4027bd0f0
zc70ca9945edf9613135a2357ddff1c06b7d03dd64712daf3b066b977eda835633ad45955bbd959
zfdf9d87073ad3f96549910301ffd53b33b97d75cdbf19f5a95d17b29ce324512e15efa5e46b2ed
z6045d61ebd40dc92e3a78588f856807eaec318b8c3556cd15f1fe9e2d75cfabefab0ed4e61acf2
z464df32ad789832d1c94a7bb239344173b5a874941752b74e116457403cdd946a0219524f76cae
z738913bd668a0d678748f63758b0b7106c6c41eeff25ddb3f21be2c6038a79bdf87079831aefec
zea4fa0d1e269b23b875156b2e41986ef060d6f8a9ed8633e541c26b3a87aa16d4ee7ae312019a8
zeeba958d9f7d747079da10e7ed96c9d50f67ffe1a9a17b6e3d6acd2e31b16a8171e4f621daae45
z1d9571e2ddefb35784eece61609fcffcc95a192f046d725cf4ded560451e4c3e7a2b6a74524004
z029981230d3f9040ebf31b38fb576c4772cb6923ded1eb7dae7e23773f81125d5d2555a86e8a1a
z02a1fccd0155ab4d52310e379085ec0f26d4755908a47d47b69dfeceb169b45cc8fd7c22ea29e8
z3f4ec0baba1170aaad5a129b00e10728e63a16baea9bdbc74dd43ea58f76bd98815611d44eefbc
z8ac19dc88fdf646c1941002a2475fc6b923f54b801b70e2fd6886e3959125ec663a4bfd40439b1
zf2b2af53c6d28906eab79d80d4b7296324458cb61e35ec47d9efdf4b6ef863be25be6bdd544454
zdad2042046e783324e9933937701f79264321e1d7ab587cd860204df38134110d9766d333cd13a
za1df0c0cec5503f29853a1705f615ce1c98cbd72e4c78bf207488c62e8705733be4af296aa35dc
z82565643c439e1a63d7eb68abc447d67d3ec7151d5238be1d9c59aa38ffafb69cc107f7591b143
ze0b4f8c4ebfd9e84ac0fbd386dfcf068f7b11560b2e4620b7cd844b811be68aee0dec561960757
z12aa3cab60e219758e10a28d075966c1595b6699bacf5e71cd0387a1e0a1ee6667cb0d8433b735
zb9d0bc9735cea6162d5b8bc5fb1c05de285d0c9c76668d023f332b693a37d54bb073e00e4b239d
z4d489026386ff2bb477460e0fed1ed311ba46bf1172629741aeae9f365bbf0ef3a9dfb725c9462
zc34883a9ac17d62456f17cd80c49bb70ebb2cdf964aa898145f565cdfae39d71c2403dcdb1fc12
ze9b813050fdc2912916ff763d7b70137121a249950c604894e0b9c932269d9f5e663a6e0d45453
z79789d5e2f3f9675266653e765b0036a413afd999fcff1c183e806343a79911ed880fa742512b1
z2a7abe66a6369bb8e14b1f3abd2e20f87500019678a7994c0f89d3a8766bfe0aa0679445ca848a
z7cc73205d21e8419d704c42d41e0531b32402b91aae00cb42d0e8fac634dc955a73a89cecf7cfd
z80f7486ff546fc70a351cfeaad1642188fea174925392e1c052ff952c1b2341fc9c43cd71995e1
z31af3f14f80015eb0855e351fb18e3f06bca17c5a256e2120b6eaa222f2c8389f8a909a23664ba
z54f84820ff5d373382faea1d3d5b0319312920e487677c63f60b3be27bbae4796e263311c6539f
z1bd44c5ef286b5e69970ca39615b653d86c14c7af90e6b07b9eca8fc58485f5cd9e70441c6c175
z822f2cd4d7e0b13df6a742dfe010e1785d0ce1801d8a6d1516ee60a495ee94b78c7cf9b2f0f407
z82aeb0b19cb24d2383f956f68cea06d2ffc33c1f08dccb7f60380d2aa97d0587714d748fad0d34
ze44a5a5add613c5c1791445791549923b8db035a1cba4f5892ce570e0ec2d27ca8401af6b454af
z83ec15335e7e08d8596d10572eb79c827410034c78fbe6ad6942a111e3a20c8ab819b2f93ed556
z9a9c40d61570813ff4e6543dbe92d60c6ca592733fe99a0ee439fea6cd4b26ea498b642cc80fb1
z041af5759ec6d8b5a2c58691377ff50ea5bc148377c984a4537a35bf3361733af2928ed98a12c5
zf3562b9fd388150aaf748f8fd2e6f6260eee68a58d6bbe2cbb61792a5b3ac8ead61e491c834435
zf5d93eca8cbf589db8faef508b35da7cfb43078ffd5ea2e0681c64c7a5a03f731cc2d7fd0f0a32
z81ab1bded8575d905cbfb9cbcde77a2ac809f0ccf97486fbdc1f2ad722f12496b8c7b35fb18617
zd4e1ea26178fa5fe35c3266140fcddac8012f39113a182ba16ddbf76dea71aeb9071d6a5cb7a5d
z05b6e4fc9716fcb9fb97852e530013243793235fcdcb9054e1fc2cdac2b2a1aaaaa878bb611757
z67df4003c617fbf16a0833e2e9453eda74e2f9cbc757f232b02204eabbd0b0e47ac5583d32a21a
z70b1262f8e722e2645d50a243404e6b01a42b43d4e0e9b4419dcce2e07ebe8825117eb382ce1cd
z27f5ee56dd454bbd636877bfb9f41eec92e8aabef50fcd475ee3414d19e6e2edcf451cafa017fb
zbd27c758f70bf0af91d8190b0b75d95eedf712ee6717f4bed07e79fa85ba7deadb0f360f4b67c5
z2a6643507fe23e08bceaf997cd76ab546ee53c9377f185ae335868bf12718c3b10544a1961629a
z888bf25ee69b20968ea1d965424bee5fa589c06250a99f8c3f76e2bd47472506668bb3980ddf81
z0581b94e1431495555fc8b52c80bee1de54f4deafe4d12c1a77e5fc059862a1e760af2a1f38f7a
z58135ac81d86db118ef23f1d49777b1befd34a3ab4f3335139e3fc9b5f7d59257154091a57092e
zdf312decba7ea09fc6fa28c93e68a146ea23d10ef3180d32ba96afd988bc39c0b8523694a254d7
z48c6b1dbf5a52dc740b1c33e6552a703230215b31b361c1874336bf745631523fd9792eda5d918
z3f2edfaf9cd5b2250b373aa00a905dadf2be4fb5c53cdc3a013563428faa976c54634f5ddb8e48
z30704629821584974d85a002beeb9f01c49df2602b6e68f12430b503498564c7b22cc68be1e5ac
z82b934462dfee3e4ff05190ced5c9b2fbb4d12b15264af5ea0b495c15ad875d565b10e2b201472
z24463b5c3cb704e3a0642726c4d4b6587c9a0bd33dd5530693ed23820d6141a00ce8282a5322fd
z2de60ad037eee3167139fb9a2e1a21f6d38586938f63ab5bb61315d04898a2454c848b16bac14e
z9ab656eb14c1ff204c5faa35bf6fe720f7a51c62446fc73c9625a25d3b898573def2529d1644a3
zc76f18624e7463d495f157cdb80820cfb2522b138a5922f27aca62e62926d25dd05b1da7d8de2f
z4f8cc2922045a1bce01f42f3251bea0213f22a244c975e99fcb1e45c36a7fdf51be3193c2cfc24
z45fa71a407bfd67daa6c7770c4e05aecc29ce5c2750af11f06e55ff88185dbe384921c70b2cafa
z54f6c3d9c542c84638c97050bc8786b35cf60bf6407cc90864e39790d1625b21936cb994a2c165
z26c6d7a713086be0b497dc3bfe112e0a9c09aa471909a937da4c08a949d729f9d6234f2f9cf391
z8d5a94fd3a302341e462f773d7f9cddd421accb0e85aff2d572a7a793a3ab4ff3170abaf230917
z78d4b1fe12f24babdb1994ac33fe5bde74e2988b0dc0061178f15fa3ca39c9cab75434191dc889
zbd4cedd5cdeaf0d1a4561ffc904ce3566e01e522f6a87d0e1501ba19da8cc5e8e99492d90cef5a
z8589fd0c1131dd726797eb741d0a6cf53d23d85262eda2fb083ae8d3bc63a4e3cd9e3b9dacd0b9
zda5e082677f0458168db51d947d3bdf7d13a1af97fcf5f80870aa94837729f5b1dad2ca0807df2
z7a14a1228a983d2c7dc33c5f9ab8773787e2f1f02b7f6e47f4b6168fe07c07d91ce96797da5cb2
z93a060f884a5b44875521cbd7359269859e5dad021b0b7f843dc184b7bddb5ae61fd475a5fb548
z52f16d5dcbfb9cd34f066569b252ea57061dd2e3272d2f75c1cd370b8a671753fb56bbd8e60c6f
z022d7dbed0e9df12ad10fa03329ae8826f19c90e2c8c2382d106aa857a00c68137ce5f9be37afe
z80e096e5cf9a40d8c61c4053b03b40d0ade96b69af19d19480b80fa987dc1a01c5d763d1f78944
za84994469ef4eea65b26ad4d6c506822e98d193068117588ef0f8cd85d76c7ec1ae982b656e575
z88046c21ba2a576d0181f4e29d6364a0d5307af9c9f49128f7c94439aeed13c8a3cb56ad678c3f
z95e1be9edc2ad7dd0aee392a74709dddc020e9bf017621d47ed38444421fe674d5dc49bc44ffec
zf5d64a8f6bd21188462602260e690fb2e70f0f0e5a6d0496d5a1f67eadb0055469c887481cd935
zdb3d04f9890e2613a0816548bdc2cd44c3ebbb9bce148d002fde592a66af61e3ca6e1461254d57
z9b2748fc44e18e06494e639953e242f9af87c81a2bcc8e0130f37b9a974a2ecc7ca113f48922b1
zcaebdd24b9dcfd7e210146bd5b9e358c5c6f669fb9ec8a492c6c0a458b1fdc28a2fcf23296b19b
z66b16a47f94e644711b6ee4b4f4b83b3309bd43db95d1b2efa94944bd939be739b4b25c4453b54
z7476a3c70bc0a07ee4dcf4f3984577fd967d397a4674a50c68ea6a6033fc120bcb57fb3af5cc74
ze8cc30cd96c1e981872f9cd087b485508347b1da4e73659c37bcf5167ac472c1b9860db9693170
z2c5221efe06d08559561a7b54b005ccb81b015a074aa537834e051e174bf8c88a0d4d14770a76b
z2d0609c20e15219685764abba88d9c803539351635ac0985d6c6360e2fba3b7fb51feab872cb01
z3a1daa7cf18a34af428c5b7f7717f9bd7d6f8cc88e3bce1a3547b971075c28e0883f1dbb84da14
z880d12b6e99241f6f1d1ef2a2f534c6ba6e236029de178b5af3c645226aa0d6e2a5d0066e9d3c6
zda457af0dd1a6b371db8489af1ef8fd8168cb45d563673e60945ffe8cfdc1acb11c17ecb5d526c
zd2dea3762b370c3d86a7626d893a6e572bb19531070c6f9204604653d0e733706ee7cd2b0fc2de
z96503dc628fbc18a47e6abf5645b21379525c9e7085ade59569dc428f9a6815f667ba38ba11d4d
zde2b6d920675a45a55ef1e8e9ca4c54db94c3d799a8d6281bebab7547b54a58c40b1c28de0dedc
z523b090dcee7bce1372d1cce0beba5ddbde039dbcd7398642341b8d5416cfe3f084856404ab016
zb2ab05a8f59ad467bc466e3e98a2aa90459745175209b30bc97dbc6cb41bdd238078f79bf051f3
z4dcf4ed7fdc5b617d20863ad8f897ea4545e1d2738dc3e49ea909f84d4d1f3d1b397f2a2a85982
zae7b6aeb113b7af0c2ccb76d72398240f305a6f075ff37f057b061f43b0e814e21f477535430c6
ze5478174f97f5546117c6b1f7da4cf484e81558f7023687729f77af2288c183993d46c7a1a9d5f
z4e4724f7d1f54208c8eeadc837675c6f1dd8933b3b717327de55901cf1babd252c72f63d585639
z327f717f5c21e9997c0de361e7640d70f0ca83674f0fc4a8826a4fb57f5f1ed720b26532c05b45
zbae25f986d3652fa6a2eea4aa794d0d0e6a1f2c708c7fa4e6eb3bec9a108230e6e01a92e38c6d6
z88c7dd85245963a9223fbe080b2898937a2820a66afca3912a892a6039390531d61dde0eb5f6ad
z9bd6f4fe0b1188353add82ed964c995083ba72b7dcdf028b052d9884761c022062cedded58aa6e
zf2aff704acbc3efb985f716d854c18b9c02486d5c27dd0b4f3257ee19dfad2ef40208fed59ece5
z65baa599c80c3f93472d41eb27b6f8a6bf16c42ca02377a0431fe2bf1e429a66e71f902c6fb3ac
z4810180388d3b320196051cfd69800845a81746b183e744482ad4a287e884bd983e7bf2caa160d
z882c2683470d4beee477bd7c937329f5a6ffa382b71981295d15fa3245720f579db85469ee74ee
z325b783b278b2bea72197a8af44ce78e8b3157e4b6ab8cacf75428e5d25ad40a91bb35031dce77
z255cf494adfe45d70ca4eb4ebe89fe87465d4b42dbdd565ac301d2d1cd371e37433abe7d41e662
z7b4b1c19e3bc26138cc4a700f5e47bb792cd885ddd17d0a5f80d0569f9a66277c5b42e9db055d6
z49aca1f268959897bcfc801f2ec15bfe7c46fad28f52c0d00c6a732e99e811c44d82d4280bbaf3
z537571413c2f85795de457076c6084d31752def6243a21477fc4cf570ba13375bc557a4712179e
zfa0b26362593e656d6a975874df2c25151d6f33409731f28b76df671b5f3056d376a5eed8f9efa
z90f4e576bd9b776c9d3423812dd66a7b18eea8a39a6bff9a7d6f18c0d0cad74c843e20200a030e
z5c0fc4f552becad992786bf77f45dd795b8e42e42fed3441b4bfa7d70acc64093cb01cf04af617
zec515fdc6f08bd044761b66d457d136e78f9aeef8c5cf4583f9cdd32ce0a8572769091cb898d63
z170205d6e9714ceeae6492fe2b409e028d60a3b7e6d88f5777563a518bc577179dae35237023f8
z0f0c0d4c29f317169ee8bd8ca8464446bbb17ba696c52277f8dc2451ecb03fbb187cd8c49f02de
z706735c8f5972f1789c1ab32f994726a5e4478686b4d75e3d79620538334f93a550dacd7b5bb93
z9844539c851e52c49572ef7965e8fe0e4b09f4f6ba79eeaa6b0137034a65b06083bf8fed7fdb8e
zcfb197ca00e35ae7a40d51d4314f66b9524875cefc56439a9fb5e74c154b32e34c39a408faf4e2
zb1b5a560870e3aa6000d144f8c7a4e2150f7c99dcf2b4c298c43728a3dc1da780bf006ef53d386
zf080ad42e705ce61e0c8a90a5d402a8b303efa17ddd9c27dc35b5bb8750bf5f0ed59386f4fa794
z41a241a4f19c43402ce61eb466d6ec8512cb6c3fa95b8e56d4ec66c0e149d48020221992b9a134
zbe93aefcd6874ff927648d78ca5d02ba8ce7e57d204d461a8968f34f56fb17fdb418d83fcc6340
z231733e5372973548c455d189395f4269db65e2512a0fb888fa4e352f1ed3426b700e9c46d7a39
z566ff4dca96426835dc732a17c40f520efcf93e9995fb440f32bc105db3ffef69c6eb0acde54fc
z9ddee5c13382543b4c51f13fa2d33fd0e7087505320e77235361d7f7938b5b5bd2e8e76f928107
z65616579ee14f0ef2c49969e9e8acbb02afc9937870e9744ba22ee038d8a2a09f10ee55683455f
z18c1a32af025b30a4c831859b7fc1703bd87801307342bea5d78a8e48ade59eb6caa6ec82af31b
zbf877a978b09fcf274d1bad1fae9b209a8ffd6bae9d2b9c727b79de83fd806dc6946426038fab7
z93ebf125faf84ebf97dbb5ff7c0d0a74e2ff87f3556b6608b176f5d40d1730ef024082b08e74b1
zf55f75d2061f2df6ffb179c30e19ecef31a9e47bb4b98bcf20d128b16d6dc9a138737faad6deee
z1e017911e8cd34b0965b7c84382a5a94b8e671417090b351671f5f6438f0446f8b94c69dcba072
z0287c07e4b6bc1e6ea1fd61109701eaf7734839cecbb675acfba78f36324e3fdfe2feb66c4f478
z03cc2be6076e88fdd2b313a08af27900af86ab2b2cec52cff290a1427f2998808dedbf52812cd5
z2fca8e59fa4467a809f42b02fd4afac5da3d510de3fe20292b4770fef8a9cb5ee3a4a52165c535
zaf0e5d80ab30ddba8f17f9bbb8fd5ce39e0dc24631e8044201e97a6f6336251e3199d4696f194c
ze25b47191890c8db26d2956bed3f8055f5c961b10596824314ac1975e441ab0b5431fe532ed62b
za5d7ffb3888b051be65330f1f684000ef2eb317ee96507c1175ec4b2c19597c62a928eef523d9a
zd0776fda5fbe7c96bbdec2e03348f7211e6c5239b619ea274d7a20ca08b10b5522c35d0ff921cb
z0298300943c099ec0fafa7f6c441d669a2f78d53df4c70e3cb7373bfa48c704e33cf27eec2ed55
z4256d007acc927cee93aa27e6ca4ada35fdad35dc9fae782fbedbbed25ac0196c5455b569059e7
z3d0cb89df3a6c68de9ef87936e64e6eba953c97e16b35f6316f45f1e9999386bd31220d5a78465
z98cd14aaf18dd2c5f484c6981ebce50b88d398ac921b7ebeb42df255233fd648d2e816f313c08e
z09a902901ebcd725f30591108fcb9921aea50620537380b74ae9712c19dacbbe58b7d1c9cee351
z26def25c8bd51f2bebb136cfa0f8ffc8a6943b92baec6eff3c214728558b2d3c6c53f159d32622
ze4f8624ae342a615488dee32688bfe9acd78570c2d4d273a53a206c9009a5f43ad647521920cc7
z7abd5ed4085eb32b7e97c0b0bddd6e633ef8a6e86fda664613edc9082ade61eaccbf217cb208eb
z33550aeab88e8e7c3248e9834c2ed1faa420b5e2176cd01eb55c0894d859ca481b80af9bec34b4
zcbee3b7845c620871efd03607d479500f166ce239de424b4d7db31eef9a5aeebe1b5bae6cd3f2b
zf463c40b9372c41b09d812597d4ae5c7897e1310028dab7ce8b46436a547f7319cd764b6ee8364
z0d8bbbe030d74839a561802a3df288e95c90fb4a97eee07fc0085e33b36e42e697f300234459d8
z38f79ea872e2a26a06e4234a8180e89cc5fb554fe9985168c1e5957c5a4c6f82437f59f9896193
z9435e9d6ea6d9423d627a892d1630cc9c1b6ab876f485736f326e6d30dfb251cfb64b9ae24cfee
z087403888a4c5f2e15c4798bd3347996ac314a437c4757fbbf4fec0ded756a23b5405d2a5e4a74
z6147b30b49278fabc662f85c1f37274fc60588a94db9f5966f7361689325b31af2bdcf0c85a163
zca6aa4df02b59059dcfffef9bea617a480c7eeace469114ee1e5b7beb3e0038ab8053e9fa2073d
zdb7b16f43e68464083467e45cd873444860411145c27424a36a5af0f4a6dd982867adc8638bb7f
z5deb1877e4910617c7f5de2c09403a967ac1fb0da434cb6a289fa769009708466a5e36296c69e8
z9773c424bdd9e4d1758267158769ae73579653693c7f99d15e51c2d4a1fb9ec51d82002af42908
z0f2a1e1ad5d474fd4d3854cb907e5b65087fba072c736c82b0ec9dd9e22a37c3a0ea405042d1c4
zd7e6917327ea9a3c3443e0b14c0850f216b16cb4d48c1d2348717be260957efb7aa87355f2917c
za414e736305e93f97d935fceb0ef4517b75224b76cad5640577704977610ac279a986777d53e39
zf5a17a0fa715dbc57436f89cf5e21fa0a0b342fac11381877642632643c4511a971632d6ec5525
z97823ad7d365f82ddab5636a8e23ab981560eab69d79d4917d228f97fb49c9e7915d6a0859cae2
zcb77c47643f433caa3f677edf57114480a98e71cd0a41c4e2d7da4f8b32643879d1236d52255d8
zc8e35cae80409689603de28451f712b4698d800e1a16ea4a45d15fd5cf06ac53c5adef06fc0f1e
z1a7867e0fb9646ec951b80e5466df4766a4a7afe63dc80e7ffba9d37c273514a8f7fc0086c9961
zc5f71d267feba8e6448f7f58740023d77eeae9232235c7b2c924b90dffeed378a56c2858b7f2d5
z27e899b98fdb3020ddc8931da276e0b3143c0b570f14a7a62ad83d24851807da3b63369c361b27
z00f164a1d8c1fcc74a85a780e3488e099ba4130562e430d40e503b48c832aa03c95f6480edde0f
zfacb8b55c289ccfd5be02aa78497d517e6a52fe6e5adc2c7da006fa649a21fedf4cd5e1091166d
z3f69e8808524c95b29dfb1efe0bf879c3fabe7da1c1cb73aae7d57b1f49a88dcca52f089b6bc0a
z14d7ac26ba853e2f01a2171f8981706f28b619869313395147adce4c68d34eadd34e7559c3291c
z0fbac2c77819bcb6edded71bb4043bfbf4dca894171999f281ae2389514fe827afb6dbfc31d5f7
z1a02978f2a9d2a424dcd631e97a349f8657c4d7f1f3a6aefb70ceeee75be196463bfdc2fae074f
zad05fcd415ebadcc183ef6a73ff880a7de8ff863df8c9781d5676d3e7876f9d65b31e9107b5c6b
zf9b4c63094847d916c4e85b74eb4a46ee3867de2b899f4afdb40d1a676687dbcfe76f0fc4358d0
z8e2176cf20d006e391ccdf4b9bee11adbff74e3d17ca2975e819add019c866a14c48320baaae12
z599b72ae2119e9b29c988a5b73bfa29bd7ddc66c00313ba348bed359da020a5c7b84ba7a8182e5
za23ff0f5d4e68072f9adf012d068a78cc02a78effb07346809b1ba7139c26cbc2da6b740500e57
z03e994e52137659c030dbff90372b11348b8c26953b7e2a18c5c50948baaf879430d6addcd991d
z5a1200987ae2fc2d2070ee02569649e91d260bb00aff8f5d0cefdd17626fa104228996c47c76a3
z5d8804402de29ceb97f38b944eb68ad3c292b4b47b909951fbb39f96d30f0b4fa55ac98e219e75
z472b3bf40cf50917ed30858cfb70887eae5d3ddf73eceb82128dcf8e19d1d0bf3917af61171d69
z39423b280e9cc2ef8b0a6315c768f3435cc84d217213d17da33c4659b057a1cfb29341c1833632
z3f64ce3dd9feb6d1e5390e790caaacce52531a6851efa5e7bc1e45ff624b45d458f625d02c5589
zeb99b93efcaf6fd72608f2afddcfb2866c1d2a8dbf822be1d5f694ebfb871864b2e85aa6842cac
zca9502d48e7b110024dbcee6d1f34a9b393ef08aaea5822bbf7a2d27210d688ffa1d559ebdae4c
zc0c5897832f91a932efb70c3d3691e29d2a5353680babe33e4172e217962bd982de821dd63cc77
zac7a6bc3e515767c62364e0ba43f1271f9b4cf93e70a5f3fbf7b435fc83cb305327e851e146a68
z9b8d75d53ed33948fe7e5705cfce5e0dec6fda07f771ae0d72e64a28aafb8b5484cb63c9248942
zfbbeafe9e2972d3c21eee8c7a79f28d1277eb1077c370836dfb3756606ee1e029d256aa4dae31f
z936448d2646f29079c14c0d620e88e960c8b1b21a46e57c018c965de9c5620bbe36c8b7e372cd4
z77c469ad67a30ad117c6ae45bd11d39d586d65a9fb9b17e608f1683e4a397ed5ad83eb283c50fa
zfec656847c75692cfe6fc2cb8597a68c01edd04741066c39e0fa046f55351d07d608e8bac31edf
z4b1b113e22fc1968546799e29c64b3bf5aa7841e9cab26e3003afaaa9c7859aea616b416b43d56
za1ad8f84d207a277bc7908b489c83073d74b87cdfb67ef510b7b0fadcb1a46fbc281cf1e6c13c9
zb0a217f3deac218bdd5687f4270471da03a0e488a2978adc7f1a05bd8735eea06281289d73b162
z6616624115f3abfddafc3639ab76f4740c0d82b0823f7d9809e28015a7966ec2d960177c9b1d2c
z88a9b1b378bfcd08b3a4bc1367515cae733ab9991cc7f9a46abb0edaaaba6fc9d9354b9a5c67b4
z989ae09a2abced885d1a193e343059d8a5d43eb22692e8fc38f1a4b70b24fa5f68b52f7a6d6ddc
zb2a1fc4fa7f6e55703979742998d7dfb301f277ee7634089663f76bb2bd04888b2305512895486
z65a317f2bbf2edc0ba4cf69b9c2c86f8e9c905aa1dfc9519cdea987bf0a047cabff65dc3bea427
z7b66319b0aa19191b51442419f051940c2907d8b50e4848745e2aaa390eb235f1fef584e9cd4f7
z0415b926494864357f8b182b7041c9a556c3e5c2d276c21a25c08eedfd7c94b68d52ea4127a41d
za4e1dcdc269ef413fc277c5f514ecb8548d2005729cfb42321d79c2320d5d8dce81b4ca05ddb6d
z902c2ee740acf8fc5d9afc33922970b6f5c4a149d3d8da6d9f67dbd4e69914092327783c04becf
z720c5044462ff58b040230dca5f8c97a02c59d0f14291dc505db9058926781fab1ec239a19c20e
z150687406fc6c6b0890301aa75f01bbb3641765cc0e98d3d756e935383ce3ddb7e491249f4369e
z40e3017d70af23dced505a0ead67bff81db82186bd6d3f445dad3fe52df0fc283d7b7007a9cb58
z843b6b542aa09b5138faaa541ec049ac4225519dbec7e54d856d5d9109c5212db8bdfbca8a3c8d
z55dab6e1e6302bd4eef5d22b19d914ebf139f068a7aa35b178eb0ec34a01d703d9b68ea340ce49
z87043ed7c9a8178d676faee7a6169596ad066f1b1e0ccb3a90a60de8edc56d5bb2d83fbbb9dd61
zf0cb6d281598da9cfb25f4969a538806a5076275404d5b29bb350cf7cd8b36a4c3c6dcb0a8d734
z8b89640c77ab5c37ee69e43be888791a7ab9831dbde3e30238b16abdb574c3f90bfdea7cda0ee1
z292c9b0955106804c9d187099010db7e7b686b4f384178c9dee0b4ad78de2b9888e4a9b31b64a1
zfc45eef6b7d2cfbc873dac292361d60be6bb7f2b8f914b30789c2ef4377d05d06853c256d418ee
z5e1ad951de72b9289948bbadbb5721d3868427b13b5faea55e0202f64a465e9d74a37b4757ac40
z2d77de5bf6bba85583b52076e26ea5e091ec145d6335d1c25e51adfc7b5574af1c4e75dbd5f87c
z4a5c799493bedee97e9c2715487cef6c92dfed1d93abccbfd1049762f8c50026e51d2074eea212
zab68106a08fce0d4ab2e43badb8c9f0e17a3c40b64e82821be0869a75c2e89dd6af05302cad774
z7720a8e966dfc8309f1fc7cb0a71105eed91ff453d9152ec370c82f75c3f57007eec65cd541ad6
zf9ca594506ea9c66a9cc987d7bdfc053bcfb6a1397c28aeb79cf6cb306492e5da6d9ce06c42ea6
zf8b9f566f14de068acb3f1d7c774ffc09e3f2ecdfccb69b2038c302438658c6635b25cf1ee4380
ze264069e1496518488ccf47c1710ed831371c9669f581a09ac9fb1715d12fb14f74d8b233dde45
z398a3a3571500761dde1da28f3357c4ea80cc14129577fb3d121b1ae96643648ea7325707ddff8
z988f30e72c417888e32cb8d7dbbe7cd88f8400d718159b0f9cb2a3a8af4cb501d1cf5d221becad
z8df8cc4af7cf4da36c9f9b1cc885d52f3580899718a3e088fda704d9fb01f4c36855b3b89abd36
z854087180d08d178666cf141db5858b95a04f2de1732d7b03e7fd43d46429a3baca3a953b79378
z9798bbdc4d447103e914212419d2e94b295ab18a265bfb55d116dd6fc965595156c839f5a41879
z45e27425972e014207e7bcbf8874487bee76a081f0dce83bc8e4280eaf2e83554d5297b21210e4
zf4722cce226964b16af72ba8c4ddf1ec25cec74cc009dc20c3a5c21e70d31e4ad362d0340f75ae
z66d67e21d583b28de22519bc824221c41b9085c93247d5658539608fe3f36eb935bfc6b40d548f
zb08f1fe79c25d1daf42ca5fb52316eecd8945993e77d7e1dfa640edd779b1e4f8f68cd9126167d
z2f3646ad05330d6ea5235ef56c14f7e20d2a6cf751034af88ea748b8f67494608b1c06a71ca795
zc9678b29c5948438ed76145a70cc86f5cf2197771d7e96c56e84eb03c52ba3e9f558c1cbf168fc
z35df27e59493b6daa882a0383c9b6ae10aedc614f6f89844486bddb8b6a514452fb27ea1d65d91
z9f32b63e65fc6204fd7b0b2088573cb7184d47e5e587fbd13edadb5892071ba3676c04c758c601
z4150a2cdca03b075a9a0eaa4667a5c42de18313113044c5232db8d61bd58d1ac569ae4353fb9b4
za3703ce263bbe0c581051679071d529eeff3357500969dec03db1754af5a182b5e614e9f0c449c
z6f1a6c8b5d21fbdafc0ac97f93e8efd69bb4bf93aecf77b0562bee564c2473fef878b2f2980c44
z53d9a0e1a564c137acf634670e693438687f0bf248da0b8ac19bf62b985cfd016ad9959295e447
z5b6c3f23a2cffac31a803215255620de7d1353ae62630fa534dbe6790c44dae62f7f0f2796213f
zd4a16d50a50921c8c8a769b8179e5cc8a4255a2b594b5f7892b860f3c2e778e56c83777b64805e
z7639fd0bfbcc4784d0b282a2ce8cbdae3d0f2b7b1f0df5d9b97009276219da38f46432b1312deb
z2207a14f6815704909a8247332a83147751176af9c58bc8b04b5cdb78e9e9beaa9ded89116a723
zb92e54c84e3b6b66fcca68c65da6cf874ae6454bfd82efb86abb537ce0fb4898ddc1115f3bf769
zbaee339e24526d6d4cb0e229d3b57b773af4b8ca8988bf2dbec46d6c5dbb7b7ef7052235f91707
zb1c64836782e2d6513492056fcd2a6d4b9298eba10ce52efafd8595f44f26af1b7716fb609f70e
zea607550fca9ffd989019acab909cdf615d76689bf11ebaf7e771d71b72a812c7d90ac93aa893d
ze89a7f94cad6de23d934d3ee98a347ec699f97d0602ac56f9105083d90e684f8878efd2de41e25
z8e0c0f8883e68cdabe5888873612b916e3a5fdd2d0fc7faaf147164129fd7c79f2704f963c1a29
zbb553f9375a0cae9b51cecabec8500c11f4da91f28a478ef2f656614a6bea4231e645365216e60
z4e50cc24fa474eb19ee552e2d96b32b96e248263a1b108c8138ea3eed11ff4c08ef3a977afcef3
zf34b66a6626d1cc3a90f01594e15267ed968482af95d573c719f869ece2c8785f93b148977751e
z610b9e783f4b6e4211d91d7242acb9157108a205e8b5aa4e7d63d63c1d8fd10189a6e9aac945cc
z907aa968f3dfa49540b5a0567b9ed6a0a806a57a64f5f7f3e00ccf8e7af1459f09c1944e3cd4b4
zbf3d216d653f9e409d0c1bedb2669880e55a01b4c22247ab0501e499305a11824eeac86481aec6
z8d18db55e33ed6dc48395a7c2b58dc7ad6671315b94c64d8e79aa720b668dda1028509e6036833
z5fc752e6270b8f1d3742220ba242f8e1d6ffb5a1e6be963fe8d8af18ea950e790a500f476233e8
z5dbb9624809580770418d1a901472529f2dbb3d353b8e331f507b06c39ce674f2e913866306fb7
z44f00eee9fb162739d22b81460f09a1d5bbca8af519078d30278b8d94a5e0bf8e9445f61702853
zf0bc72b6ba9148a6423ece446f79f154c2dda71270d4920091c1e0939527f69e5f95c4e1e0732d
z04916e75ae9e00c51de35037eca9c54fb22df849a2039f1bee2282a6ca3383b5f84a7eecb1dd13
za490fc9114cb43b0af6dab9d7874b08a15684cf1b28481bba86975eb61402066945d5dfeb495a8
z995f015cb15c85874c42e4b1e7db66f12b3a380b5293af384918512fbe1bf86b088acf516b0bd5
zd9316392295fa7970335891c9c4d925cc4a9275d1551dc21726a2dc6a269d00f350567852c4a8e
z5b6fce9a7b551d3c0694b7f5a3446088903cdb4fb798cd13652c311d8d6436336764f5710c1a9b
z47d96308fc7f3905dc544e9837eee823bcc54c9ecd225badcd78934a868722916dbc5f35a2fae2
zce06d16a6704ee0fd6035284d0fdda977d070203275ddc29b3d009f3f36134d5870d2e702044c9
ze8d2e6ca10013f84776e5d6c45ce7b7fc79f0c89d10481af4a9f9b033df5ae1699991be93fec72
zcb6eaca283ba7d6a118b89fed742a567b75b4fa660a52b840902ab9a2e3f3dba73a5137e9a2966
zb58ac27c83edb19fc97e582c13e46cb76e44ad6e2bb0c312a04f70c9b0f933298f5deff86f599d
z9db5fb64fdc7cdc6c72a278d1fa7b6c6bff7bc8bc89b57fa93cfdcaee5e04253d2c0d0c63f382e
z72795b3005ce579956d31561a39321f01380b492f6f9032624461b3c432efda3597296d527b617
z20c3f35165e5aded0cbfe654851e860db9451fc31b14ce5323d3af5a456318dc26af0db49434cd
zdcedd6c99db2cc7913a136014760cfe62a97ca218211e4c7ef9273b38b08b7e636ce010f5e231e
z767876a1e29035e59737f0b18f19ca4048d1543f5bd75588b111cb5f9379014331c000311e05cd
ze58fd587b28e5a45b21cc817c76ce149ced8d1894f6a721e51282013a34e63da92c2f7baf8e2c6
z3e499ba082d0b2eea495939ebe3e54c91d16e88a8751325b8c61e5b796b01d52875f5709792032
zc70aed7093fadf15674a4f5e0ee0e7f463e26eda4b02d600036e2469c4fb00089e74827b2391f0
z6a6cbcc82cd8175d490fceb9710eea45cf2dbc38031ef158739cec95f9c1f124d243d6af4f486b
z26525fae92886585d5a59cd0174c0f56620ed38fe354bfb63f08174e9d133b28cb08c081f6cf86
zc3556767faced794afdbf3efc8e7c22801ec83a34b0c7c7a25b0412d2876e9fee04904a88cf673
zc8127b91035b19599a71e9e518b4d28890f9a67ef637aafb1739e190173af7fd21f4deb0ae5ab0
z93e7c923b520d3ef4aa0c193fa1bfe05a9bd372cabc2e8f1672c5c7dd285693e2e3da458f60965
z51abcd767a7102079cf92eeba0512e216f89ebb9a3e4bf7f0f5955be85e2ea06b15bdc17c91288
z8584c5f17b136e188d34822a09a83cf60c60d149b0dc1bed08405efbd9fd0dbefc452dcec1fbb6
za453f3d114bba83164a189175f09e68f7303e31f7cfaa41417555686d2a26c88c708983b35bc1c
ze3cdd5d75822370b5f3787f7e4f833dd63b08b07dc89b4094309f7d510ea5af1296099f24bc332
z0dc2ce64c9155a0f534a607cdbf44cc3df646ca2e52ecf242c3396226ff4a93c9eefed842c214e
zac1c24594a43442407b6c3928e80cb6f1b6f1dc6ba5a46b7eb736e15f1a6cf51b9fc2aa21bd258
z71a7672fd04eb6586989cb443604ed24fa437b67c0f320898961d7667c259998bf0a93b5a0858e
z27f204de0c4297f6294ba8c6f7eb18c674d6d3d306cf964dd53f3c804bcd1be69b7e52bfb8e9e0
zaaa8e1414122425d362373b583dee7d757a10d651bcfc238a987120debf40ddc0bd48a13307e7f
ze8092323f7a15d3a8038596aa9bb256555c10dbc133e609ff55fe53992713fad9846d1c75bd452
z63e5145aac2f93e330c485f13bcd2589cf2db53c37333bc679b7169604566b00d4b14dc9599114
z94c568ed371f3b9d414adad106c828a37c8cc0a566dcd2acea63120ba5ff1864f46c13dcd34a49
z7ff736932d598881881772b8758cb8e4185171d2279d152c658a009416a62337bcfd5bb67d5f89
z47ed9b78a3854c05d0fc2f30e3120ea1cecc37b28c73553eaeb50101cdf6f0a6505feb7234323e
z15ed9bbc5b56fe192406be35b3e2b58702a0fde72b892bc9ef41479c263a183db84cd204f0e789
zb0b282a898f46d06f00ce9d4d8b24ae521f13437afa717ad163251a912cdc1c857c87f1594c0e2
zf0cb9733517162bf6d51e512365effb49f5bf58d49318b133fef2fadcf966b3b54b1e105f56b3b
z300ca4df10d2f0b3c3aab9c272860f64c83dc08263ead218f0c9bdbda4ae332c5fe7d3706bd66a
z232f26030c967a5edcaa59bf6d6ed324998ec722e0121889da317eff281584aff3f45a176047ca
z6fd4af37c6ab5bb593ff61f78846396bc1024261a18d71b780b16441c6f31d354c09325c51a5fd
ze501ad0cc3fe3f809cf8b6fa31e6e1677a74ec4805f078b1e20014e7dcf8066339d1f7e969e9de
ze9a404da1fc41b2946248b7ec07df7aa13a4bf959c8f969a976b1627f9f1ed1f17e4d9ef49d211
zda3bf688e830a18be46f118f651b22834eafcb30d7ebf31b8d3a0101b7b690156516811d57dae9
z358f5e08a9e84662c9a3ad332d5b008e223f808011a9c5b4409b1a3ada3302cc9a008c97298936
zb0a0edf6d854b8b40fa6f06de0ecd9c9f61b1989cd4a18d13201f30794dcdd6b87a83c08a6fd37
z24751db9f23968ca59b4589ca174dfde64bc284d22c0e30faf41b68db0fa7bdfaf4c5f1f7fa776
z7d9e1267ae52604a85626e25562e6b9e75b0c6548eb2855ba3459c9b2908818e9b4afaae3eca56
z0931f86cfe905d84452c78b9ceb61318d41332e82c2dc263d69e6d70c9c2780d7cb1112eda90b4
zfe2dbd3e5b7b902e81e5e58b8f85ae5ea3f592d56afb27a9a1866891770d60fb1e3b89c43e5177
z112979da09846de2211f29b75f0850dcce56c6bc39146391fb089d3fbc1add024e38c1afb4b231
z80cc6eaa1eac332ded5ec3a2fe22377e59a5e526307a78599b5a233d449e0e8b97b3f96590ed52
za1f412d99c47a17cbb6737470354b755587e379d6f57ff0aa840bbf58d9ab7e6c072e2bfa16636
ze675ca95f7434b433b4660c7f05e516d31233d464915c631f96d7abcd3f45c4f1e2876641ad73d
z2ec2103f3926d89bfa0dd5cc9e63591fc11d37c0aae291051aa7741d00a82f4519ee5725fdd8a3
z8dacd6892692de5557dda713e7c308873ce4848ecc4a024e1443d3b04984b1c8c11a56ddc73372
z5f831bb17f484c9c1afaf856844174aee2623b6370ac9a4a3e171c95214294e2d128d346834385
z9547610d679749f03f77c7dc2f27acf748d110f0dd75660f8b54d2bf8733c327855c943b2f869e
zad057b5ffb5fdc528822140b85d0cb064bd1565be90b1c1b2a1c864fcba870c5322d1a76a48fda
z4295ddbce52c8de9bcdcf3d77b475245f851b0ff1e106aefaa26470ef4a8590e0bffcf60907b00
z4a3eca74bf5e24e9f2a6e4999a8ce49ef565f1f4ca4b020a5e189802dcb2178a24809df232b7e4
z2c10550eb8a288d73a66064945335e5bb7f04b83478b1d18f4b11407c61fb9f1f2832f2cbfa441
z963a4e741fb09a174ea6c322de784603e944f3709b24e409a2e03aea006bab39e3c2678bdcd9fe
z61d7c8d33d5da48171175a364369120cbda7cdafbcb7ff2409e9b0ff4018c811266e938b57c235
z973c9d9ca3ff213dae55f4476045b60ed4b1642c505503218f3a7ca1d8df288a6b26e8f51b54a4
z14806239b81f115ba9f8b2ea5e4727e4cf43faf9d5156a6f8bc402a29bba804fd44b7c9142387c
z89d4d87bac8a4c76b06e332b24acdab30844a4f125446bca8cc068feb9e2b95c71937db99b24dd
z74743b411e4fcaf2f2646ce5b489e65e758db42fe777af9832d786afb3072ad826907f0b3b79b0
za4d1e0bd4103a4ed3336a95d5f95b52e34e19050f5da185c6baaf9c31f629ac51a8b63baca3b1d
z8dae6e4242edc274ebfcc27f873402c73d34ca085329d69b5a5d43231eaa26f5fccadfcdf7c445
z9af86fdb9303335eedd46c1df094ec9766433bc8d793cb2524479e0261d801bf4d131491f1d55f
z3076196278c4e3b8ce200767a8965d3c43aa5cc9b12e104462fa404407acc07719d0635028b28c
z841060741dd1be5009c34b97893f75429257c15fee814a1273e81f1fb0584edd3e915db2d97edb
z04ea849eae43a47376c7213002c32037d30b96c5d8fe53e46b73175b9e7cbfc1e34a7778ae65cf
ze325a9015ee1c2e99e8f7f3671b6669860d425dd6df26dcee1617a68fbda8ec21b2689f794a819
z596c284cc5f80355fd67ca551780bcce46606831ca50a68cab426844cd8f8ae6f7a531e00f113d
z3134ac51403844e05b0bad6fb8124f76de926a9f5abf5b3b666eabaf7c8cdb07a6a2417c20cf5d
z6be05ee642a3bcac80034ed6c0cf45b1340df67cae043db4c5a0ad9301a0fcab12e4eb220a75cb
z8f171dd8ea32698caabb9d4908d8f88530bb5a963c2c97e5062f7e3d8ccf7d9b57b0a9f14857b3
z74cabc4b1f5a2bd8f4568884f2fd387971b8520610de786c3cf9e592979e13459df2da770ed5a1
za755dc384dfa2fb6ecf29652051c6cbee882ac545bb064b8acb7aa9fdb883642946f02f835cf3d
zac5fa15e040710633f08b4b418feeaddeaf9a48ce0048229d9275c09383840cdc325aae083627f
z690aa4f67270cb9931218a2ff84ed1d0c786d8c7b9b4dcfc2691e536ea78456a40b2bdfe0e78b3
z85926a38cf23011305d5d347662de4dc0927444d507deaec7faf4349b78952d9f3f20bc009d478
zf175ae4869ef79319173af03d6f111ea93729ad357e2781e0b9e88d7d55c47b02a4afd3a29c985
z99538393463ff9a3350893e6ea34e19510a52217a69163d3969d3838ac7b8ba65fd87aca129271
zd84f2b0a6a5142ee6923923f4e7480cbeb634ad42c28d907c8f189b9f5bdf73fa051457a6058d4
z8b9b6833d1ad2d5be636629d1afdfd8582d575ea5827903c3c0a9a7255e052f1a758ccd0221803
z1f5e9ea904e0922755ad068c4c67afbabdb12d50546cc60f8941196fbe67f3c4385514d59b0d42
z4044e8643ed2f3b15b4fcf59798ead472eb2cb6cfd4f72c757a00b374c2504d9531ee1c9444ac4
z1e279bdc55da521e05593461196da3b471d03f40a5cfd0a9de419b4aa260d0658ded3420734e58
z0306c00ca8f325f7078d1d2bc59b967efe50d12c278eb0bfd3270a2f6873007064d9592192b9a7
z8e2dd6ca5c741bfc3fffe99e7cf808399dff5e250daa77d560c6fe093c4966acc9f594f2138aca
z02e8259867cf2cd7387795c24f8e51afccada5ddd9b60c2acccd6341dc905f8fe1dfb393e3b5ef
zf4de8948b839d08a0ded7b3891bb386a0a15af98019baf67b4f496f8078bc6d1ea4ce7312d603f
z19645e39580fb5cb51638f457e1b519c386b4f3788b847161300264b61dd334504161f7bc86e6f
z042dea1a9f5950ee001a5e1f4d2040c511229223adc5950dae77e3ee5962529cb2f6ac16b0df30
zd304f08208fb37c55789333509eada5572367ff9511ac33bd8ef04284e864736f0b77a2d8abc60
z8886e62779baef36f7e30e10bb36f0b60789c6ed3f3ed8faccc93d0786c72bc8dd5d2a5bc3fc8e
z738c1018daf5f32a4f6010057b4d3f013be06f7bc3e0168c62798e93735747659769aabfa1f831
zee8154fbbda0af2db9f802d5f24e9bf7b9bf1a9a407dbbcf1eed2ce7ad3f2f72f9ac8ae61af90d
za23060239d4d135a9d7ff77a16fb2e2b902cfd92b2329ab9ada70dc27b1d81426b82d0514510c9
z32070e41da1dfa6601f324a5a6a6403d43f7457ee3cbdca4cf0a2faf9110bde74e8e0d494ca6c8
z355c3c0742c800b34a2081bf7009eea98e2bca3738a1418d15c984f7ceade1fb323447dc6eadd8
z1b8ae43a4b5f1d2ef014b1eb1be59b62392e3e583b2fb36f3649677d61229a4251f50217b12207
z77686af8da340bc85cb5d4cf732d0a957af07d101d8bd4ab12738a92cdc947c28d5f44e5293c54
ze51f9d510cb66256a7284e5c7ccf46f3ac21823cd3aa9784f9e10864d739f06857b589d0ab22f9
z02f6ab545ca3f670ba0b9d28f831edc14d13c2fd5deb35377a683fd6d947e85fa8a6a4efbefdb4
z31c4b90a6ee78ffcf00966c3cc93a6490cc66e2a8e8da907c6071cc68ca4f6b8f4d8ecbaeed8e5
z8b89ddc0bd7007bee85ee49c3e6deee5484260d4b9ece4103cb55a4bbd9f8e123a7585f188ef73
zf79e5e0ae2ef4d090da20f99cab248819d3a1ca1795808c4dc98c9e7582416bd1102cff0d99821
z6f281e48bcae5aa3f71165feb1680dde17cb3cc8eaab856374db2544b677be54f54686ce9c2ead
z2f46dc74e92ce7385bea0dbbf60202768eb878aa28657bcb76a62bc8483ce83551ba706c4040e9
z94c29fc9fcd003b5e2d4863fe92da06c4594b30827685c030284f3de6298c14ad93e44180d00d8
zd90647f5c87066c798822a83a9ecce839a48d733f682891f81b250ddf3197b565e4daa01b33b9f
z5aae0e778a2bffc342b70461f732bacfd6f15e7d18f6d4cad3f0a8ad8d73c7b92a28d545688312
zc7aa34866162bb6be1ee3bc7cc9cf26cd8300b7d402fb6073bcee2c77f295ed1b5fc4a8bc115fb
zba7b1ef8fba09fcbc117fb088b315d6fb27154e346346ea4d118c75f713f9206557ec0b599f68e
zb3acdc87c76025f5485761cfe274e8858ab1622c6359e17c54b885eb4f53b5d3c5f0c83e7cb404
z045fc3cc539e7d45ebf9220d272e4a65f890b8f665f11b7e727486b6d8c36f7bc591f95a508efd
zd18c249c000b7337aefed0be776643a5594570db81e868bbb4867a1d6b7a10ad0806fbeee13dd3
z7594a1533ad282a301a43e9f12bf68bf6c7c9a23b9e40ebfb8a0590a8f76d49c3cb4ac8aeef970
z99078d0aca103c3f82f2f0574d1232b4625bb251eafaa5453dcde932fa0adc557671444d225b21
zbddd1dc4992ad3a8fb7aee95e93d368ff4b4da811358443579ae88f03e816f4cb714a7103f47fa
z22c96d4d22aa8c12ed8cb2c9be8210d8c0ca2c5386d53d736c87b53739b488177da6ce8f2a41aa
z0d750e05ee267043823bafc0b31fdb72b990b42e4afd9bc01e3e2e468cadf98cd3282c392d021d
z78ecfecbd2815210abe79b8829ed8e43e4f7ffe3dfb29948f69ccb728542860ac89914ceb5ccd8
z2e55b93286d42c3b64579270f42232ae183431108aa96435762d10af3fc156ed443e7472ab92db
z10a9a7c759049d9e03832e83fe6aebec3859e9eb9e62be0b3aafde2c0af6b9212b3d70be7c8f25
zd46bcb0e7e48db21544583e11bf58305daba909ca7e454c8b5662e0892a97d060c8c61cd7d18ef
zc315f5afa08901f477bd2b5ce4e144e638e379caf2b6e51c835915630d9d4c323dc4ff88672a42
z35e2567fec2c143e7149aac24b8115665cc539ef61d546972d306a3a3979803f65a8f42da52f58
za669e8d50dd2008c0c20254d2cebb085c4f2fc4efa1b7dea0c0c5ba5547d584de17427e6b1b4c1
z1f74254999ca3831863c98bcf7aa159d3b76f5635bf1be9a8ceaf1aae40bbd7a283c0cc14a4cc8
z85df98fcaff745c314738b1561f481d4d0853884fee0b3e3c24f2417a6afd05fc3775c4ffbbb77
zf586c0162ae8a14c47062aaf78050e215a467d30a96f38680de1f240657234c2accb8079c4d76d
z174fda7174c69aafe7a64eec64d0155fa23cb92984a9ee4b0bff584ab63578c74238ee1f4ae74d
z544219c8044314a93249a0d9f5bd2faae383f692dfd86f22e4be66767cd49bd4bd1ff5f47a6db4
z2a99ab4c80d4e39bdee70a9320bf2f5ec365670d1ad596ee0a167a343ae60b7a4baae4bf4564f1
z1b6c24d04f4602a33b35bde1668b217cc60c41880ae6e280a0a18277922ea3514fffaa452f114a
zf6ab3258cbcf62e4a7a5dc0a5e84ecbddb40a3de7ccd3e49f1ad6afab50dd18881f499b2635128
z40d90a019ed9169c3742cb46dbe1302c62419497246d7d565d457284147a4b7fe49b42c69e1fee
z3ad527c8fb7fdddec74e7ca96e6d357cc714ea2724944bcbae9db073864f49a93cc3563d7f684b
z457a982eb704a7fc802c1f47208cfbce498c4e26fb774af7535a8ed444a64f97f634ed47b9195d
ze8bb702a77d067edb17b7a3ddb47d8fc73f5f851efaa3377a3451e291bf909dc5515f770d265aa
za889c2c3ace55386dae8afe4c62287eef45a02f49e42d3aa940c6ad8a8634d53cdf747301f18a1
zfa5b6c974ec6551788e9c8a61eae95017f1b5d4d99167645e406d9451b30935cd332b1b741be72
zc3b106b521f37d427a4c7fc27e929fefb9139cd342ad194d080f82c09c8ec6bb3ef53f746e8871
z9d3c369af01d76836a02389deeab6c1b97c512a4bf0b210a42eb63bbf03da9e0cf1d8c48cdca9c
zb6d3e8a06e8133b870ab54c466aad95cf316d921b44812fc088cf60aad403a0e054ce9e46f9bf3
z6cce5ecfd8cdaa7e037054218df3800096b48cecac21aa309a82f8b82e89d7a22c827f54d2578c
zb90da53f4292822dc3496ad2c9ba01af248dc8bf0ef7d86049fbbb8e01f5f27328bf280bfc4e3f
z2ef57638c9fbe2bbf77517b7f8f7a644b0a63054018297571b44e90247f15f29c49db49bf1ac3f
z1621ab60fcf49e705395cf7e90ed67de8ac56c5be72ed53f355548399636546c37babf46f72ff6
z00bc910c46d9dd4290b02f9641f8cbd447cd84bbc1ac3188b767002eb269c7da8b43425722e181
z80a0268bb45de74fd96826f8547c6db1905c4341329279659d958609bc5a9b2534b2b2c9c405a0
z9f26d94f18e0d8b05cb93a15d3487a758e109fe626fde557f4d2577faf1b6c06e2907420d0bde0
z73fd711cc73dc8cd6c4c529b2893993ac744bcc028fc1b71f8e61fe86227e6640cddc68c282b09
zbaccc4bcc00143ce9e9e756c9d0f71f9679c50ba6453be3239af7163085cec7158276a13dbfd86
z7d9493121de8ae11f17620fbdb2449b770c087546166993b2c17838a50e96b5571608dadcbc036
z875ec33096bfc6e33800c290021c7814c6d4fd449785ceb71ffdbeb22be8dcd14a48e008df3cc6
z3596d4489768c76c75e41c2419c7de53532f99fd1c333b897a983de39dad1df7156da5a15c2592
z277426a4189b3504ce37bf12c9c2acf487105549b0e7ac0e8317be11df73d77132276fdcbab5b1
z2d535c66b6cf949709fff7a4c73ab749a126f81d718890eb3c1741469b695cd652306a5e9b0153
za44f1b1d02cc52df2808950e9cc0b1796e2fc1b73713f939c57aacd66bbae8492517a10e53b471
z493a383cb1697c5b29463d5f8485ef34bbad77d135b006dc1a92b03880654438ab272d6579d0ef
z36cf883f2fb7aab8f2576ed24ef502143c8868020369bbbdbd5a111edb1a6cf64fd304880bbcc1
z0b0dc84506e26107e85c23df54561d08a3993eae5a7c3961eb447757c5cccd8af896ac08c7715d
zd0af2755dd5d5d3d9b40c5568b57225fe8e5c7ca9f3f632aeb8385b160d3a9ce3c1f7b3b5ef34b
zb0a55750ad894468fea0501e039cfc718d62a201c6e84aef2754175d8a703a4f32a249771c96d3
ze637acd23242054b53624c20a205fcb74f8b53da8395cd132f07dfc5bb849d31931b2aa8082d34
z8d9d42e410b20ccbd481995739b566fdf2689eb33e994acc99d8c97e970b7a96ab5a0cc25b0be9
zb65b815989aeba96906e4f3b46d40f385da93f9906e4268be5de69b6b1326a2dd21b5fecda00bd
z09730252c7233d3adc57e0767ec04b5560b88a46b8ccd1ab1db31269cccc470fc7f71581603c25
ze4cf9361d5a6d74cbee12e14af1493e2f58addaf404c6c1689506e3e48555ae266270ea451a577
zf37ce7534f2cbde102e1e400050af51640e1c2661521707321797e0bd524a3243ec0348cb678e6
ze2680ea50ec7f977a39694fce46bca4e646ad00199753bfff1f90f331435977e66fb2c2b5c15a4
z2123d56448dc53842c40bf08a07a5e04ab3f7405e8f7f9ccdc7697a461e0d21d30f814ac78116e
z822d00fec484e9355a07b664292f9d5312e7769814ddd4d741346b4fa7959a78f573e3ca0bf0f4
z0ea9e58b1218aca52d402dfd7deda5b80aef1cb8fc5f1f2b95b51c9b619f9940a99f938f2f1974
zdc52568cfd7ef4819f37024a3dd55a59a76baafc1fa8ced0e3c39ee9be72844ef3d8d4db3bce33
zd195ac3e70d39af553b72e545de17622f8a2005b3485d8d78c68178219732e4ddb2796e3e0bedc
z832d94549475f2264399df4a07ed9b46287180518e56c7b9a670d1e7dd5a9c62de46282b63d604
z52816848558155b3292e76c76016a1cca3152b53e0ee12f1daaa661fdcce024c7e59a209c28ea4
za2a487a32fd3335bea2074249bf868aa4d10eb86693cfa528cd3d4ce749c43a8b1852577376ca7
zb5ace5ef69f738329bfd7059b38740a6290445e492ffa8129fbc1bffd4102926f8826079afef62
zda625686ab129ae5006e1b532bcb3563f0d4b6dc8e1a744f1497a4c06e8a599d5947f85e03a0ab
zbd168a35264da5fa7b58a7029024d4a93d37ea71ae7dab5d7df8715f955a174c81c7a3472a9705
z61c5dee91c98bca13f92ae9e29fcc2bb8366a0694bf9f22d8039c9459a5da5362260d2aa363299
z07e6aec3ed11558d6cf4558ec98852956a84f6825755cd1638183b3f8fe03ae1797b836f684575
zec7345bae2a38d4570fa135d629b24202cdf50f77eba7048bde7324ca1b180a52d77ca1e3883de
z28b41c7ed934615152e982b5c79a048006733a97c44f18967247635ecd599737e2714e840b7513
z49e8dc862af36076d55bb55a14d4d9056ddb04ef5121dbad5459574591720c5d3be98703b56be8
z66d3adef2bcff0422f75f745c18e672f3bd263721af5b650038d6d8d611e7704c1c994ddf056ac
zfbde9f752da7f11b18990546f04392164721bde9988455c572f5a9be88d78d392fd43217236e38
z4464eda97f00603b128aac447731a8349dfd987e92a3371c3e268c01221fa3bbc0566c824c2922
z4a717a89dab0abe6b0a50e03cad1f61396a0f4d70671a5898efe93851f777e319740856c4d8a34
z2ed77003c1525cec0128666c92d7ecae023f43cd91e03f394417098400007e5c63ff031179fcc5
z34f7ced2578ca55428927fd64884a9e1c09085438c88209784091c6fe8798237b8db7861011f65
z1c49e30905821c0812abda0d5455cc503fcd1f1b581e949fa29ff6b433c85a83334b279e519e5a
z8f4dcfcc272e782133d3215dc9b29c8e30ab0233c821641f9cd17ee272a800aa8b2ee2a164bd58
zf2328b7521124debd711f69aa2fe4c8439430b5191194ff8592e923805876831e5229c8d3b1267
z4ffa3b79bbe4f272db1f493896bb7587f236996cfc0ccad081928ec1d7a8671deaabac6cf04874
z4bd4ad2793c8b9b1cb585749ee788654d74857cf1736121696b729024152bc61cdfee2731ad132
z4f9d5b30b4e292bf73c978bdfbc70464f07e5ec7ea6ed84f9bec8204b0b62f50d239e8e6a2df7c
z0c137676684130be6914de233ba3db5ce5a171819cd407a8ea4f045bd7018d3e617b5526aeb020
z9f6cd8eb698f9e5725314835eea7620937783eeb6c2401f7aa6cc277a2b9259f00efca37a92d44
zb45066619eee4f62ae1b2353ff48832c7dc833731617c5e1e3454641f06d8d88ff532eebbdd490
z1105ebda9be3f668a9062e30e6a7582f8764f9ff9af7291cf53851460ebc2798bc63da424f11ca
z319c94a2379359bcbf381fb97daa0b9cf117e9f8ead5cb46620dbaf9a56c726d8f697c65f5e3ee
z3f5cfd144f9e0599a813b6474274392b068d54d98a8ebcd9d5f2b3f988eca37ca0ef35ab868d53
z8f409a2c2c79c9239875a6b4b496c138b029be4307c882915c65d0394bba5e89455f9729a22c4a
zc01958512d93415e34c195dd24eb3068c24f6cbee887727fb2060fb2377c6fe026fcfe6d321ae0
z68f1627b036d1108735b64df630d3a0bcbec42c63507baf0d1b993bec65a25666aef88bfa337f9
z2a60d3426219cfd3edf0ec4fb599f55f1edac83144f0c9490605700e762cc089b728e0a3a5a540
z1d64be51db79ae8d4ecefcc0a95fb420d8a2a0fca3a5092d917007262dc17540bacca2a316f00f
zead568a6cb3588b7a2bffb802bb1bcdb31958f2532131c630bc57922ce218b3f4bb1b1603cc1ee
zb8d60202188aba2eaa6c9baa82197dba0f61e329fd1d0388cff267c46abcc35721d2157b15b395
z4b95e907b55c75d8465e1914b97f7fd6f09a4e322e42555ca21a0849d232155c8e9a1bc01f5fec
z7e6c93d5b4a6aae951dda1d85d2242cc4a28d841400eb9a7337bc384b4518229620cb0da2c4c38
z8adf9729b948f3dcfb810f0105c71be0b96f179fe40ab918523c5758e749820e3bf666e338a875
z7a0a2faf9487b969a7c54334f9099d080f7766785afe5d60224863fef1283bd7db32f5d06798d8
z8fccc9a3a64b2584ea702b05f0303acd1a24fde583332af6d6e4e9adca44d3fb79af076de9e5d4
zc6265067a958078c9f24eca79d5f8073fb1eefdb70b046ecee91809b4976cdc141546e7039757e
zd908261ddcfed945ff79e4cfd914a93514769997d2e747206e9403c0e739874f83451ccda64540
z63e6f18bf7fea8ace9d3ce52f11a6d65165cfac7b097fcdb18d7120f6fcecfdd6cb967a382f8d1
zc39e225b88ba34853b981ff5a8926e079a364887ddca36d9fb1d5e7ef6d245eca627682c3d3d75
z6a89defcdfe1a1c6d2d58c1292d615fcdd4d9acee3ea93b692659708e9719e7a9d65f81dcd06d7
ze25b6001de8ae737acab2743170e453d5665f15a58be6bcd5a59341a02751d722ef477ddc7906d
z229b4a6505feb4243cc77db2335e79969564ba7e706219284cd9373873992c775c98d2ff283c07
z31cde2344935a7da3a75268d6ad568b766f04e67e3c0970e4da11d1176e1a6684f7b717b8c9dc0
zee8e5981d814924e7f77d9743acac627d4da09bd061a9f283175068412005c04bf1cc2864bf56f
z25dc457afe28bce64a8c3a9b27aeaa39fc3bb52b8a472c7f1c6b1609584da460176ed58a5dc594
z3ae2ec23574abc1840e6c585c25153507b25a514b8bf050641bf7d14dc90dce897b048157950bf
zd50cd5512403e5d6ae7b3e7742f246162b0f44b87b6baf9a1a4cbeb0f4d8e3df78bb65601f0070
zea6a36bb93313bb5181f55a3bcfb5ca318e39f9ada5b0c53b4a5e6727ddc4eb328e231088b5db2
z9f9f1228a3c6adebbef911ac5f3dafcff355b75bf1664d57899ab8e420d76c20df186aa00a5903
z83ba89795f381b332731092e5e3e58a8447488f8eb5736e62dba1f9760ad8dbfbcfe94525e17cb
z8d29f22b1b39b88ba887e21a37b35544e44e9ea6db3c2fc51f3f8161f57e9fda3b469851d17028
z7909859c49673771b19729b918ce84fafb67777995d55c0e1540206a317f16476e51ff3f4c8ba1
z1a200e2d037719b2d329d0e5715df32d038e666310057691f4fade38baf4ae8ca779ee8a386444
zea413e29c57de05f4612f438e14a0a4b11cf5075e4313e9d0d9a627e9ef3fd6a317f29e7012097
zba25566f2d2a3dd6d7b85f442caa76f6e40009d4ac26714014b00e45a420917bd1b4c53759f41e
z50fbefe6bd189bfd86cac19948adecdbc572280e4435ee9a0410413fbb02629a5c403b75face93
zd4eec0e39abe9de197fc79ec22244bba5ec56cc656b6f0b0dacc6f487ad3678aa8a51664a47abe
z7f995bdcba691bb3767b3787a668e4426dcc5ccd2dd1a02d0d3d5cdf886c9aa4f745fa12baa1af
z9818c3915b4ecf32678f09d5f373b6c5eff659d81d0924915ec834782eaa74be67b67a1c36dee0
zea23d2f7dc1f5a16998fb239f85b69c2067d8cebc01e6271d18d5eb8f9f46f2bf81c7798486fa3
z025fd1b9e80a0081afce86aac23f1906d1070c60c9763d00fae3ac5624f3e0437760fb24d02500
zf9d7fcb35073d8adf7e3c040348f1e9752ded8026b79235ae6508d1e9dd3178f7cbdfa9f3561eb
z145423154805f0417998e1c512a41a24e0032e391978ba6077cc9d0972ca370e4e8119dca91cca
zb0ff0dc98e32b3263470bf15b620a2ec14028d21c73cb81e754fd9ab4cdd602e7091f7768c14d0
z8770be0848233182210320c04c3441c8528e538a78d215a96d3b626a0f885ddb3cbd45ecbae5cf
zdbb4fb2fee712b52371c89434e7034f4b74d7440a395b7810fb0b40a596fc28714a3a080bf430d
z9343265c70c0fb111403e9b3b341a5bae03e5445c781ca964653e9b415ed347eee6765b6260fb7
zbaafadc5d6a14a68dd70ce7084a21094f593a8f7c372f172fef32ad4253ebaae6ac01c2b5a9bf0
z7185260f5753cf78d76632ac5f1a012fa5435e748fb565d3a9be6681b492be00b2cc0bb348a383
z89d7f4cba8591a5985980d94a389c3f0a7a60d5dbb7902e18dcff2d48318fce62061bff7994a30
zc23ffbf374390977f3053129f2d3b643b893162e4bdb860dad9da314ef48ab4f9cbdd6d54c556c
z419b76ce4b38ca5754cbafeac62e764cef7da0bf28e959f1bbad2e1221d087e8ece3c02b4a8dfc
z355b3ffd8d84c3d18db93c87dfbd0e4a8a43bb9538e7d2384ce8b54e29f243a68f225487966058
z96c6097b0263af2efb27791de5d05ff64cd03da7a29e456efec4839ece5d54179de42cb5529070
z34ed5ac00356e4be50549d11e9dc0264e8c6c92f191aff9a6b0361f2d342a5a460ec93a33b5154
zdd1decf923d3d4d4fa048f6fe7fdcf5d38afda1f59ca6a7373e15bde07bc636170a7d3e219792f
z9bc8e2dce83ad3d1ed80c95b8bf708002e795cbae0150e099b9686dcdbb6b8be7cfa19a43f902e
z71bddbbbd7ae63fadc066c5ff54c77f053a0fc8e0396f695e7af8f828e327198064402117188a0
z69b4370dab452a6e53ee94556cacf83aa13cea3804d8a44b776b785beccfc24c84ef6e13bd572e
z47fb732ebff8a3168d673104ed53a0dc8c9b46b1cf38dcd7a2e35e9af94d04a601607fef0da499
z301a82cb323303a101067c79e97aed06b3acb374539a270c456e8cb725c3851b82ee97d0da835d
z13bd0828ab692f9b7743c22370fad80033cc31a53a2a9c7be43ffed81bc596a632ff8a9b81cc1b
zfc0b0b8240d7f5debdf85b8f78df6122f839cebe7f91338ed5048595957016a78b3023ec0d1a8d
z0ba8eb7416ea5c6a5c7e1b17ed84f64627c3a7e5b776ad07a2489d4f8b33a05b1aa7b268c32cdb
z8891dced33cd5f08e51c8388499044667e28ce9493f8360053a7c6e3232272610b9cfce2a9f9fb
z732502f13404f49c1c19c4b73a2178a8355f85d1caa72bdda1e38903e57c4655632ca52f6936dc
z145239af5793b2de99b4cb8309e5dfc299303154411db2fbeebd527077519ec8d531d7d0967c77
z0073af482420c7acd8a35124c57fa178112306c1f2530dae10d7b95d68c8f4396702f01f6c8b0a
z2433f2bec3be9f6ef0be5681d9790e2e7dc472e5eab9d4835a8cd61e0d5824c3b33492527569af
z9a407113fa4588319ed05fd6edb4e4d28e6d36a54671455d6c606c0df966b4ca1fe6c86e22b9fb
zdd1f5f5ffbec8754cc70e95be23457cc5b700c9344b89b498dabb9821096b170a564f26caaabf1
z703ae8781bf1a9903071e4012ac3125a6ff635c341ef090b540f5b1f7c2a0a56bab722270b0b45
z04bf5f5c4c7c7c20c08676c10f4bbb7c4faf6b5780c27d4c801c765e53fbf29a3c41adb739d17f
zfcefe96e62e86ff3191c8be065aea1178b9f1af22660d266a88db09754f859e52415021b62346a
zb2ed24a45407a7f9bf43f5aa5ea22077ba884a5a89a9bb78a94c59fc0c240855cb9a342b6a6120
z34ec9600636f3263115e8203e902a9c87b99ac0f1e4da8c5e251fc746045a19e789ed49ff60f83
z43c4508b16940d9ea43b17e2cdb08dad78488838fd9d41a707d5a57130cb0a9c24d9024ae0daa5
z5b1eb4f4df13b691dbb012893508d023a62a44d30cb5ae06b1e04b03caea313b4de8a14d44e4c8
z65ab1008f7cd325191cf2ff7495d19b8c120f19c405f4b05eeab79152d5c4bdfc60bbcbbd5a4fc
z481ea5c391f64773a35b6e2f5e6e4f3e360083b7b4731bf2f0f32a9b51d7aa9c8a1d0a200508ae
z7ee75acc779eac519ebc1b80f282b76399a1340c189265aa50f8abfeffc597df7503449f87bc33
za8d899ffe6145940dc6fd5112cc61881a2b22a19c5eae1621a7e3c2ba4685bfe549c598ea85b11
zeabff4215a0887f25684e7983ccb211c3caf76bf3788f41f5986a41833f992e411c44d8a5322c7
z2ccee2173c01ac35776fdb231e22aecfa264e0e18b8060953f6a1f1a2f12521b08380ee386789d
z6668788b2051b85bc45b7f5988e3715b796b887ffea986618a5864882f67a88f9944e739f5c2d8
ze03f74f8cf460949717a276c1424f9ad8687f67e6070dc24d01a3db2fda645dd8f129d881980d0
z2abc90b57dd5eb4a3dc9e86e4fef98b2a10b956fa2b039d98a62bed783ba8fe1b4f8a1df96dbc7
z42423300279a9996f69580481e22b6d4ec8fb5523195877efae1e5e36c8a31b1e065e083cad42b
z1591238702a0b1757b4ef1348018423fd833ecfa45c897c5b0fbd779d769dd24290dd92cf9e93e
z2df8d0985e8271aa0ade259b58afaac74384e705ae239bfcd34aae05424c90113f12e292e30e0a
z03ca54b5b33dddd6809dd203f1c9949f24ba1f568d5f720f222e22dc82b4a9247f20bbf4c656d2
zfd5fed6158934a96996d6c5a05903932ad79da4575e66511c606a625b404be56496b386359c2e8
z11c81916e3bff18c2efbace8f36a8e96cdf595760a9b20565542daf6ac9193462e427aee3379af
z533ade38e0aed922958f4c1b1bc46356e0f151b19baea6fb92985010d4ee0a6161541f979b60be
z24dca86d79a47f84673c9de22dceb6733563672153c8ff3907325ad54c035f9216f9b2f8ad34b4
z5bd74ee8005edd2c0d516d340d1ebee98bf9c3d12793e2b802127cbe269b9b40ad0173a3663597
zffbe7353bbd4d7c55adf83d80307b6225b68a23c0d6eafdea2f99c64a358ddc7cf87510040fed1
zcc6e7b3a5c1ca9c50725052bde440b8369d5936f6279d7f42aa5a96dd3b6712b98c19c6349b20c
z5782269777cdd9b5335de9f3f94527892361f857dff07b602590133aeb29f1865c916760ff62c9
z86d8c9471c637e396c9afcf92bd6609a01c87cb26104b3746695868c261914b1983f80e3e70421
z5db12af7f7ab9b834c71797b14364dfaab6321b9889d5808e052bb00293269a0fc6c153ed9f92b
z3748a2c2bd40965e086036fff7118f0149ccd267d01bc909925a8c76ff6cdcb5c1ed8462914682
z641eedc782df97cac547276289e487b7b75d33a347ad33a66f089503dbd422cfdc4515afdf9405
zad7dc2421b84632136a44f3630b0e682f97c7a8f71a83ecd873903908bb7bf262afc32613e96eb
z516c5e23ded0328775048a03ad7e3c392a228c18be176c813de39cdc04e5c5115d3dae319edcc7
z1ce79496e71e18be349fa0b1e68ea21d2cc630f16ae48b4152b2f5328b05d86545da99544d3555
z2acb8ef475d8bb70d3fec6eabcb7eecb4965c19ca176a1bfa885262af9619055a9e90613d6bd78
z87c5468702df2c83b13788fe1bd26fe25a6a4822b872a5b336d5dd1eeedd5c22f207db7d9f52f4
z35e39ff469e097682dce54189dc30cbd647fb0f3b95f45b7eab0c28e85077c0087461c50796e85
zb6a7653ad09861f2219d356916aed976ef82c0f7696127247ea9d8a172afd2c4e6beb36f158c35
z0c94f6301aa9ff5309bc1f9121a1e741a655b7d5bce01bcc71064dfe7968237316b2f0c79e2da2
z0c14e0c8222f6f4f99fe9abc5fe08174a43083af017a5d1aa8de9043a17d6f106adfd96260c2ae
ze8e0a645e303ef640f043b21e791bba06eaea1a57ead055da2d0d26c65d84df1bb7d379ab68c3c
zf1597be3a0a4a57f99d28da2f0d5c5f2c53dd13e351251d02eb361f5f8ea9ef696205c931f3eba
z71d359a97f9d716e928d3e0008ab76363de79d5127068aeb1f31d4dda866a2cf180c332eda827d
z30adaab37f23bed04b8724ea4031106f0c32483a689ef25d34868e69143db49ab4e99f0ad50b60
zff28f490589202210c690fc702530ad74aad5d8c249618a5caeca2bd2de8162f645a2c20c9cfc6
z5d179cc148d3e8646c2a641f6b69c8cfed3f58f8c3e6b5c8afb64e19b22099b5e924a8a0b8c4d2
z98a6e70dc84ad1928812407bbcd2a53815ffed4e8b615c588c915f10084546ba0fc7a66961db4d
z6ab19ea528b148abc87fcd7123a24d27f4b1d66de37e85b930f5b68c7c3e52f657815d5e24e1da
z200f088a3e282833438c13cfaac47a22fadea014008a0b8e1f3c364130b4c5951b83d5a2351286
z46460a7af5943a83a5a8085e0563433188b33d12bec976bf0891eb9a52d35e7e586e78fa0782d2
z7c77a1bd7a0ddf0f1ed3e534ff5d1d6a3fa27aa480f6137ba3311034b64472f0eed3dae353171f
ze11641039eb52c02c1a0232fe8355a2c83d96a820910e802a93e88985b8e01ff06a9411f2e4efc
z5a99194a3eafa88a3547d3733520741ded98e9212d9cb1a7a6a94fc5e54e6d0ccc3439dc76985d
z701e753d1be7070252e09fda6e284b8b5ddcb2ebdd8dcd4f8a5eaad51c36386c441f90b5b28db3
zdd35ba66219aec5554f795a5a985d0124047099dede728eb85f7bc69165dc61dc4270c1a3045cf
zd7d9435498b829d5e38abb435b142c59f9743ad576665635295fd05dd2f4d7c85e78c1bed0376a
z871a7482de41cc681851a5f6c00c1e5cd871fd93bca1e7822d5f5f454b4fbed983dc366c070682
zb6e40ce20804bd997e803ca8bc30e5a0f8184dd747e4f6d5a242e4d1eb7656369b21f89267b3cb
z6fb091f846c7ccaf1c010dbcfd5fb417321787a80c2e14553f12613fc72e4576d9a2d46fb5218f
z815a5d39555b08cd211c2f93aafbde91599bb9dfc44327d997a491c4fd175095d192036fdda85a
zbbc6d923392631f390b3e370e31d2ee4c3de01ca4b8af159046c9139f7700fbcce7ba4dc427c6e
z1463e20068b5ca2c32473ff00ed76690558f020c921b26506da36b1b37434dad50b806150ead71
z43a1c2717fc30878b00d1853ddeb8ab52bcf7b4f4931f2d9c0621af112c9dad3365df312f9a2cc
z718df72cf130f1fc54f85122c3261143f57c56c2c37b04f3b62f1af8b089d4e889522f903a371a
z99ed71f44599446f78ff0492b7eb08943edba9c74cffd516fbcc4571144dd1027cfc6fb9e899cb
z94445421e02bd98e27833c0b974fd3dde05a965cee77a56c3e064e9f61569ceeef28127c158bfc
zaf9203787baa3a7ff29d6e258ee506763dfb720aed9ff88bb37f948d381e7f760a5cf2087fb059
z9436559bffd5a2337824a9585e08c3c6fbaa79daf23d4ed47cc9eb38c84a530bca070a1b623055
ze9098dd23f41d18e5d749c78e6b85ae48340e2730f3e82244cecb81f9ceb0f4b30d2d3f35c271e
z87c186e4fae3056d0aac957164e1173eb1375ecbefba500b37733e052930c0b2c9c6483a5f539c
z8f1518d90a9d0674b15e4a3064cad4fe009c2572e1ff5c18736eec55d2bb338c3b20d92187eded
zd878de21a70128e1c4b85dfde3dc3800a48b2245defcf64fb4c090d501e1a8ea7fd9954fe29c4d
zc146295a7a47dd330c202da967e0e16c63fcb5ed6de4b50233698c7856785fd4ed5f99d936a62b
zcb4fb74d8eb413055b214757eeae0f79d86c34313cdbad6aa66cede47f4914c5e023892650d263
z47e730b14c8b42d986df210e017cc551d8f3018f6cb82dec2511813f3692d4737ecedc8bd80432
zf5c5b28db2e3a92109193b13ee462ac5612a155014d28549bc3babf7264c1f01f44a4618167c70
z048a4230ad4e4b06e8a576b51ebbae14d11936cc906bd2a496fb4f82fbed9dc41066c3224ea93c
z2027dac60d8285d8cdd7b8cb0265e55a35d64c56783767c437b1183c1236ce41ae2d64efde3652
z4cd8cb5932a35d4b46230e3687bdc2b4131c670c1d559f1e753d944be1e7eed1e151c66917a483
z9274d1514afe838a13d85854d59de8d8a62f36147a218b62b7acde99d7d0e6bf37b7b563ef1ad5
za2f4a80a5045dff7e011c953054acb75ff0a32719b97fecb8473d083b0933430d099e2219274e9
z666464d4a34788b8ce7c324434ae9ab84fb8783ab63170ab173e1386d9baaa64175f489aca6738
z958e76cd79c599972d7274e95775d9203e0a3d627de7ccc03573c6519c0f82ba6b459e5d3ee571
z73caa42ea3b5ff0cd52e701250f8b43feae1dffbe1a4b64f51f3db2c38a75d5986d7e5738694bd
zc97e769156c394b5eefec0fc33fc5f1de970a6ecc4ccba0cb77bac99d391bba179528d6e699a55
z9fb3b51eb44bc6cbdf004838beb22a4f765b5cb81cc87b16a2a4cec9419af84f29ef74c3e18434
za7bd8cc921b6ee2a7e014a84f8dc9981b79bc27edcf0ea7098262fec47573d4c0c35af63a801a7
z188a2bd95411c5e2568214962c7acb14774d68bba2c54094249aeb9310a1a34fbb5827b8fce854
z627fdd0bbdd3d96328897fa6cc7228753dd96c1bd980da4693670dfd3f197c856b78a8ff33000e
z7b6fc71fa2ac9b85f08445d729d4398c2662c21a3f2fd17558594c1e7c8f215f08689bdffc4859
zdb6493d65c13ffd8ee433109b7e54c0ac316ce0ad0706f04e15707d0e73ddd555f736bfb2648cd
zf4fd1426edccdcd3902f30208ca37fe3fa2e9715e6f59674e63c34d0595fbc21670ee2f5716166
za045e58ec1113c87543597134b3c405c9638f97b6a191b8b9ad591b622142e7a58bb61370b10d1
z9e3e3a5e1f48dc1c1cc181fa2a393ee5ab99a1d946065783facabe99001c956bc3b31be8d05970
z914feb885fe48bc59ee6334927e374fde57535ce802441f6db145644496f1abed6b5a788e47e84
zf2507eddc13c673be094d190a3d982f912e2a6e19d189fc3500252947653c62b6d99bf3bbf2ffa
z658e48deec7a8374156675d1733b41cc06ece6218d73058941492e7d6bf1272acd656c492b3fa7
z7f04a2a75e360f74581dca450a9c805bc0136c1c2ed5a6c4edf4eb1b653dc1158cab5091c74223
z49253014a79cd02b9bad545a14ec1fa1ec143392765b9b4a518698f67a6dc8115d11a662eb1656
zd5d75d5c81718fe7754e930f4489f34925df7815d8cc0d6a97a21d0a8878bdec873e3e6ab347de
z84c5ba3be458d109e06cc86aaaff746f2de1cf54c81befcdd69ed9a5f47a7a80d9fbd490d2b95c
zaf1b92c6f748df78c008ef09d50b338aae4d0430c75e43fd64fccfb3ef3b7105def1b9f2d11468
zf2d04a1c4212533715e41b80712de982410cc78e64eb785dd37f9c0ee7763a89881a66e7b56656
zda74c6df33ecab7c38b5e102b2a31d70de4eb0dd54aae293134c87fab9fb61f59a452a682fcbbf
z14ba08332cc71cdf318bf948599daa85cb31518c74df8879d1c1e202828047ebbe79270de7c5c4
z0457befca168e21570ee3dffe924760c0c088e98b170b0247f112ce0bc6fb0c4b210312539a200
z399c317619b27b412a518d6b4be6343373cc71a97c5db7d684371e17d853459c1d3acc1dc0616a
zb4bbfb02a2ba7e14d55f0cb2682111e6d398115e17eb40c76652d9bdf04c2778ecea685b980d36
z29673276d0129dea03b313b15929068884fb505d12a985eed37d4bb09aae6902e7e38d1f3c5640
z51520ddc87a8d569f104e426924916fde6129d622e0dfe2d655475ac5491380fdfacefa85bef1d
z7918b6e76d29d92dbb59c037480bfa96ff9c7e4b5f13d1c842b911d7f18d6293bb4289073b5268
z8cbd1ba914b8cd1e947df0932d2d02d9c9ae9402328b95597b0433b71a312150ecbea1a2694596
zdee0ca6ac7407e21045a0ba58abac73c77dd1e612aa2d6e0a21efa7785e8eba5964bc139956f45
zf2ca4888b663a95e2bcd2801b5f57cf406c703ad55ac8c017ef429340383f0fd54bda549284d35
z8f41170c1f605eb3acc8316aac8532db2c8dbf3a0f7ce1ef65af5a08f179d8b923b72b6616a21a
z3fff7f2cf1f26006735d2518c5dac0d40f2716e7e2bbe8bcce9326de33b132872239a4fe413b15
zcf5cffd29dcb9d0de23047b96812aa1aef177a4df32b5ed20db0c6540e7bf37779b79edf816a4b
z38190e6172aca469ccf06b2864863aeed8a353cd54dba0cc852518d8653e69ccc347e13eb3b558
z5c568d094928c5d5288b5da6df586429ec223c34ecf1a116faa2911c9fdd64829e3351c6738326
z298ab28d86ced2e11297388aa2bef9038d3a915d9da55e072e5147b832af03f7d765901a70a0a7
z2175d980d960fd781b583d3a9574ba4506cc7a134c66f48ea4baf7046dd9be2bba4aecf6106580
za23f9c87b90a9bc475f671aad5bb50b93dd1f52820e2bff8e35b6bbbd40c2ad4583f35de35141a
z44536a6b89fa9d1ffce39946926ed3eb5da67b2ca8c2176d6fb22bfb78542e68cb7db1cec998a8
ze2dc3e30278a73adb53cb2c70f6ff607542d44ccdac9b7b72b9ae601aed788d987167beeb5ed3c
zd98718080d46401f694b4bf81aa05b08a43e4a36a878756b0ddbdcea1bcca68ef987906898f58b
z989005e1cad7c029ec008d9e833becba4a4df3130251bfe0dd1256bab4af7873ffa27caceda14c
z19902ce111dfb81cbad3d1ce312d413ebfe3a959d53c67f583dc3d3872544d837cb129b959b6e5
z42e6c18d47fd1e24fbcd908f6d4388922a26d71df517f62e25efdc9fccc1c2a6e2583bdbae98c0
za6f5c0ffd6ca49548b03a9c01be62915549a54e06115023c9c8762a56d664b12c4cdffa7aaccac
zbf37c1a580d8adb7f44a38b883256b0aec0565b644da90f8c7f0052fa3f6036940bca33431bc01
zc15ad6950f64297c32667ec4b61cad4b372d0da07c2f46ba2f23d51b0a03d7fe87c5e34d1f323a
zd48e6411385154e802417274162a429f045c31986846559667abbfab65e70257f7e11540d609c4
z958471c7583845baafb6d2aca0e2619c77ad2f0cd9330bd9eea4ba5c32ece0957a2e2a92ed8d5b
zc93a9b50ab9e0c78b76225e277c23d96a1160392786c485017e69a3eabf68e60e0c18b8ac410c3
z2c51db4a93e0ecddab5c7e121a4a5cadb9521be5eaa7a2fb9cc55222f1a8379ff152c6279a7dfa
za6c0023cf3b0ecc168728969e4e982f03882b279c11e15320a70ff3192b8e17db1f75a78772de9
z43790d7bdc7c98508dabf6ea749c786541ed02ba21945eae41043086d63e8b72f888f8b39f67e2
z8db93d019c0eee88aa5efff495a566cc429f7f3583e91b2f7d0386197587a7342f72bb2e9a30cf
z2c709836b55c37b5006fd6362a211a013e816c26923c98f606b4ccd7df9c444d4fec412964e477
z75756e92116a44b08ed7df7d7014876f1402f90a064b52a65b80ca63adf92c631435086956cecc
z5b9ddb6e67e2cca21c15d9c371a7e4f69f526dd832aeb3be8248736e080952ad77352c2f87dd91
zfd427f822047021f14caa69431950100b7349721066d07ba1dfae51090244d6e08998aba7a2f3e
zcf9c8e59a7e9939e721c7f1cbd8f8b9a0cf870a8bc9037c9dfecab541e295b7bf56ab3606027b3
z9c834f89bebadd6860e06485c6642f44bcff1a02d083b11ef6ef8122b55cad38e150d9640469cb
zb73212359b29567bbfd8af584840ef4f7d682a11391889473ff015d2d9adba13a74c2b817b3104
z704f0d87f8be56560f8297f939cbc5fe81a8df9574fe699d29e4cf4bff5053a302de80531e85ab
zaba20cad7772b0966d2531dfa9a17943dcf469bbede0f354fa1a179dab4a4dc79183dc3e406ac2
zeb9c959b4a60d8954b0b545e2391a4f019480dff9d798031164fb90be6bd0eaff891aea9e5a3d7
zc4805c738f811e0eaba4662acf38ae48628b727b4b90f6e3431bb3c78f91242b8035e2f2385c76
z339983e3cea5fc028edc5d4a733d01ac892ba00ea18e3b9bde2d6d9325c1d3ae6a3d069237a0e5
z06d0b43940f365da2ee776a7eabea59f1c50c1d7a4b0a7f48cfc3e59df6f933d44f3d3d3cc4a21
z81824e658bb66210d1023e1ca4f583c1de764e27c54ebae6a16f9c830cc999df4a25a0334c3f4a
z0ff74d4d9793c593f6dec3ce836e4ebf9b55b54cc1085d7850df8739e228bc5313ad2ae5f1b816
zf44fda0dcfc4c4eba7ee82000545c243f0c342c416e3b87a9fefcbd6a1ca360d9498661e82cc13
zb5df46828f80a7a27c9bdbe16594c5cea7c81c2064d90af2c1d84b8f7b3702b708117aad7308d4
z07e5266549618254b5fb375e6367db8eac5070bd1366a7487b862ed5bb2af9bab6cadefc7562db
z5dc3263828208311c974436945c20da84e7b26e957fc31b93a5b6a720ce3ae25c850e5a33ff34d
z83e7df38a292be7111785ecc9a8a06da3fd7d867c2b019641f73ea52c1f2c3a51d2c67781a5d29
z024d731f19f3eb5748a8569556f1424a01f60ae4a36cc21c840221ddb48b179fd675e6069608c3
z81bad96505c33686e0742ae44a640383666c82c21a4fec01c17b7432469c5df9164c25e3822e94
z5110c9286da581a4c93346cc953211d3fd17be611397d6e7c56cbd21b164fdd8c12894fc38e8dc
z51f39d7099b012e5ef5ab3b58f7067c1366489aaf0d10740f5b99641b6ca9f9606500d7f4813a9
z22039dedf3224c3cb6f1e6999db9e847bb8a1480281c7249dde816d1c76e923cf1c16f07e64cb6
z9a90fa75338efca61d4e0497d7a9789bfb1701939361823a37de270605800200f22e4e0f7c2b34
z8485ef4afcb5a62dd252728bd38b41fe5770738525a69633cca6befb33eb0d546044ac343a05e0
ze9dd357544f21e99314683ecb8922cbdd69c03ed6a5dbc6eadfc0414780d98376e265c430d8752
z746a8732a6186a1bac25584acce3f7ca4accdf19f864a3cd96322a2584595e968546d4fe53373e
z620ce7afa78d5118a5dac12083d49e4a60efa81dcd98169714a68e2aadb2922c8bb784148ced64
z5a749e010ba781211dc051e85aad1264be20bb4bf370bd2d1cd038cdb7d5f4c92fd4dfc3517235
zfb90d1c23dd2ee92a2ab6e1afa591584821420dc98b85f725176b8c8f88a105e1f318b39514c45
zb9fbd29565127181923a5c831b1997a00868fa570fccf11bcce8ec3aa737b168dbad35a6008003
z874b35180b44f4f80fa597e0464c35fd8f7bbcab52312dcb9073ba525954a40a6a3568af094895
z07f423cfb32e1d40f2e2fdfedcb3684c2a15c92b59f08336f74c3aca1927112490998360e90891
zaaee8b6528a3bbf8ee7878ba22215876532ebd7030b4c17ce1ca2f5e39945b0c71d13f071b1da9
zcf652f3653fdb1bcf2a25db7e38a88e0f9bf69c0aa7ba8162a4c354303d1a8eade8a5246e59830
z987cec1f3dca0abf7afc1d8d0ff1d35fd12b43a613d4fe0ca156510a53c19dcf43792b99130134
zad4e0d4d0c6d39dccac5174f63c0a251277970fdd7922fc078ef68f20e63ab0563a6921561c511
zec70870b9b4ca800fb1d5c90479a47a462fc1f5249dbe97d6bb72c4a354f8e063349e876fe31f6
z46bc840d4f6b553b150a2f942fa7e40cd998749b3bd2aa19312c98b8d905bd2fd05d46ab1d3a3a
ze10194bf038fabe203923e9774ee00fecbb2d4032522b7339283f25bc434d9a170396e273d44b5
zd65e8274396a197645661ee08b30495184057344959d32550406c4e549feaa702a4fbb7dd91ecc
z07db8cc4438f94974e106e81c09d6edb7c48129d30c7b3f09f1289cd748f7a70033a22bb4dd6e6
z4315fa53e49d3490e7569ddd1b53ac892940dcdc225c678f9570c4c1571fc610092aa1addb3e03
z7080fe2dc6ba1bcbd1b7b14cf0469bb63a76e0fa7472ae5b0bddb7d7fc5571b590bbddc166cdfb
z87742dfb012451b8dc5d13934dc7ed28656aefad09aad13a2b06df9bb6edcc03b6646638aa1a5c
z1b4c14c2f1cdc2049dd73e140f7254a7d3b1a51dceccd69e33fa8a6a38a00b99f4ee58e1a3254b
z87e66c4f812ea92b6af9ad7d09d7f4d1972acc15d01861ed169f31c4f0b2659123c1cc6718b307
z8faaebf00f02d4859b45142b6f103ba5ab5604b60459af6cd06f1d35320c1314597e7a9ee87a8e
zc9e3d7e464d2b7ee13c6ec62b21a2e8a3b72ce29b08b83a41504cd32f5c27e70bd57ee35b79534
z120c97a15e7d7ba74da5de930ba550d6491d58adddee0aa17b9bc1f4621249acf14d1eae6dba94
z57e5e59571d09acfa5a5bf9f0ad2fae5a4531caeb082164d74eeb8cdbb1fece0d2a70cd7397e72
z8f6a9553a45bfede5c910a3e56d7bc7fc415fdd79db5ea4f4040ed0943ab7f4a22285f2f6284f5
z33997d82cb5056fe7b663e66b9cd3523bb37b0c092db65cb2b62f0d25c7676edbc2be0115645ce
z536b7aa6bfd33a29f7691f1a4b28efaa52924ac299530079856bfb709ab2a6d1a66760bb99916b
z21719ec054e14bc8218ff446fa75bda308f05cc029a533dac514601a2cdd51c93a98277446447d
z2e88c0cdb2140ec7ab04e8f5ba8363396feb4136faea6decd58b94177d904f171297760d4c10f8
z2380989a7fa0cfc6d41e6db72d9a44c6e936898461f2244f4e09a475f1d76ad405bcc7eb216a20
zd64c90241de8724b909c08998f3600e05d84ab7f98753328ad23cd220bfeb7350e29406849aad2
z283cc52ee60fb712edf280e163dd9f10f3f30224c51ca9227b8c084785ba188b1dfc55c2cd6976
z58435e8c706468da8c626627a3eb43b69b3edcd2d3734734f7fb767235b98977dfd83160d238ee
z2e8d3b60479743aaf2b992c685df617733895fb981140c896af193df78b5c8598087e07204c580
za9441d20ba65c424fb6dc16a9a9509097f55d43788a2b75aad68eb3f4cd31243f588e4f3f41cfe
ze9f65179d2ef2c989c3c2a32890f5d581430ab8d3525a7925550d22883b29d4e7e4e0099fb5eff
z5cd3bcfa538683a4bb0de8f536026b5999a4a6bd90f17b9758615e735453f3f2e87b8f6729ebd1
z1fbb83b2099e9674b90107902303cca332218f48bee4e80ed264323a0528a6fed596a75d71b591
z686482bd464e4887dca31e854377acc88ae80d755b7c8fb7bab90ee33a04c207ed93c5827425fe
z9275e5321edba19471ad822d98de8c856e441fb95c62a6fa642a3ca33245991416198bc8963e1d
zca38276ec84422d99370763618b9a8922088cece96c99ed3ce6fe13da7d6b56c6ef7ec6001edd5
z6f1a0fc84f54becada5444c7113917f28edc53652475e3dade67108e931f95b1bf2c8d0fcfba01
zb9ed998c253756dce52f7c467ea5211af52ac51be5d1b6808ade01ce3686b8a640a922017365bd
z58680732ca52501a16f5786d3f1f71f4bef6cdea7434793132d524ab619e385639fd96df6656a4
z1ae5c60d345f08095cc319b23bd57e2393c703279622304523a30b815f0ad49a7f1e4704407ee4
z43e132c53f253ecf3e24e646f4c0e459ab9e1306a45471f06336cacb3de39138382bae6115b119
z4a388388481260e60f22cb1147f222a01328295e7de333a8fae8f1c3b70dc73b10073be891b354
zcacf184533306803d742f3a5b3101568ea796b8967cc674b3bd529360586c9062825222180ac13
z29ceca3fa6924eb16d57745c68b1c0e079976317d13823cfb99faabc2a95b6ec0c39f8d5570237
zf0e50ca273a7fa254c0016ffaa395367524e8c554120f0ab449a48c0839e4159ed4f6ee2c5f0d2
z16b4c9c64b805164f945b011cf9bb9c7172bee468f2d0327c769194696eaf515e3d30e0b0d8dfa
z1bd55fa4cfa9a83241e592a9d80ca5ef1eded2f9cd867f18726a63c2acd71acf9d479a4cbb3ed9
zb1080b54fe9be112979a2ff4ef78d1ec35d1f7e628c42c1eca5f41ca8b307d3e6817567e5c2a15
zb28adee5492388ee5c57dbc2c15721bf1f72115cdbcbbdf01273120ab2f008fc52b2706d432c5b
z7d260372d862893e795755eb71ceefd49266d0e69e0b242c25291e5a182383f6dd579546dbc19b
z72f503367fb9854e099a3793a47909d0cf311d7f4e811ce62331f6613ae445c897cdfbb59f5030
zf764df79e44bc0973a43151be1c86c73672aa394c81ae7167c2428c33be5df5896b0f9116600ad
zfde1102fae897c46fa8228f996da7a07ca699e76a0df88b67d84cf95417f1189bd85316f995a49
zb7c654f7a5c7b3782512656c4d722127fcf096be07b9f07fdabf52b58f7cc7fdfcdcf2ebaa4c10
ze08124c2e1dcfe000c4af621f01e1dcbc14a02db36b8565b1a293ba81c84f17bc745d45992b315
zba392d84d54c6ff9fa99903baef8aada753066c84548a413930df1f53d902dde54f29f35b1e4f8
z74e7a12f3383f0f4bbaf1f286fdd93269b741fb26fbac58413514401fe0f3ff9c176e96a76b187
zb29b64fdaea99ab611d34c180f8646a62c6b1663b6964670c79965d158f5b381b6d79158dac8d8
zcbab3f81c6d99cbe86111dbc4cce6cfbd844645ae55d22857389bd623ab1cc7dbcad4396d12298
zf76bbaeffdc1739f937326bbea2c941cf7ce79ffa4132046d6cbf57212104c7f791cee86efb06e
z57847881b7b703d04a2c5b42e755c42f25562f40eada9138ac8c6087b927fe025a2a6370e8f454
z77a59894ed1c5f19d9320e044b6a901aa92749db40d1d43db74adc0fde2185faf9630c507662ad
z2910f3ef535a0657a4cf4bcd46a8de43f557b2167cdf7176c49c40d53b6e06100221a9e17d4437
zfeaae15c4e3e5e0f566f4484be5d6d5bec3cfe9f1135c1491a6cd632d57ad3026bdf5eeac9fdfa
z53092ea7da6de3445e2f21adf548b9c41d307d9e48a292702a5f9ee6501077245000343d047c45
zfe14e703526451bcdc2e2492606676fabeabce782ab707412b89bbdad8bf5252b8e7aaef2ff41f
zea14b87f9837b78364ebcd3b4d5edbf91d137fa5987369cd659ccdf8120271b0b63f8e483e862c
zd9b3abeaac2273fa113d2d61edd0103d055c3df0dae8be0826b4e66d837c82b2faa96acb720b8b
z72484656c3cac92066e74e42dae54cc972cd2ce1c8c5886adcc6dbc39591f162071ee4396216a1
zd89035b828dea267e463cbe27f394e90e30ba84d98ff899a101a9b2e3285523c6b9b1cf3a7db80
z887daa92cd4b8b7364dfdefb4e2c18faa7930592df15b1f32c6227c95f5b60abf297830ecf05a1
z714918612b82decfcbc65de1c0c4edf624a4cd892fa6293fe7288a855ea927c700b375a0b80501
zc7ea28e6ce0b41759093b9942ba3644e7033236b0244d9f2a718dc1b8cea709165bda80383695e
z727b6a7bdc423295b0a91ca5e35405eae4a691947d2ef3144e92a15c672bb8a54a7947fce6f77c
zb405dbf6cc648ca7679d8dd51fe454e6fe71b32613b67eaf26dcee7252199e3527a450cb8d82fc
z90640acf6e11cd37a8e1285499c413d357640dc1e8dfd5e482a88d235d6d8cbeac5f087743a74c
z0a4203b025509cfb5f91a4feedce8e1bd2a01c5b0ac7c169f0cc8c8378767fbcb89e053be1bc1c
z2e5e99fe2d2dfb620d2b325bdea9a04ecb816b7a5b3284334cd9f0e36d9af5cce672d16918ac02
ze01e64321fd935dab9a0e981f7d834cbdfc474e0f4e7335efa080017ca0e8d4af27c0b709afcbb
z3662fdd469421d490727b0e5807bc6edfbf543e8e42ae5d38c50bc6d32b3995de487638ce5e074
z53524146b2c26de9b0f692ad5c3e6b8d68af3b125fc3fea9d0c870197d34be82f8a31ab0ed5c50
z7d9046ff91cde51585c737b41ad922d239fe42d2c6fef4ffcb24fa040ade942f30806060c33d31
z3e053f318ba48d667e5da33b1023437bd01be48ca0b0ffdb262ad8df37e23f69f52394d70ce378
zf9191dad09db9d03b15bff5ba35b40c9354c0c9c879ab735162ed2e3c145866dd12cddc0d97f9a
z9708b5e5efa782c8b767199f7d1968f6bc6daf46950537b172778fa3a725ffd403de8b00347909
z4532644f5a764a38155be241ac1ee53c7df05fe2802fbda7cc175a6afa771c1820501a7533deb8
z96ce1bedfd1c179d9f07896cce894c7453eb13600f53b0a441d4779f1b38e994d682883d3fed52
z84f7a4bd827b9d946265928ab17db48a45aa08a93c53ad9e726e4f15db11693e853eee34bcaf43
za1fb706523ab8b3477f0bff7cb78bdc95a26e79ba36f2e9819fc89d214ac299b73d49a582bd43b
ze24137b2ca8c2062c62ec581cbc26ff26e0aadff9e7fd8d8177d17c1bf2dd032ab009e1dde2cc2
z4101d3a1cc9160253e9f5bf001a63edf636881db2941861ed65637d281a209363e293759a43e8e
z264488e50830ed754c105c2a05a447f5726d0ea77ce94d6f0cc2a2b646b016cd2eb30ed01be817
z6d54c392a9499cdb1d0107058872f0df7bdf956f6adf37c16a9732b19ad8045971941f32637948
z4e33d0d2a2f1a36ab8e753a09ee7a2264dce6bf28edea261a7dfcd22a3b6d968d2db1eb112878b
z023bc4ed47e0bc6f094d7433c37da42c08ef9affde97a4e690f672cf0801d4058dcf984f499b6c
z532b2d2182e5f37c5373656aa62f251032af7c68e02949db7a12b8c9586d463e94d32f3489da08
z500b74a0cacd9e17ae5e3e61e6ef2c90d0be7c08bc36afcc9ed030ab17e0dc10c3dee337c3a175
zd26050948f5b649695f1a833515bb70e31d4321fcf468fec6cd683fcd4fd09e046c066aa2dd605
z7b5cb2c0ea4823b6281afbe47db9050307e0244eb727d25df500846066404729dbc6a8e59a8b3b
z8359bfb6d597254770e51a484ad39a8f544d36e4bf2cfce0728a86dce2256233a2ba5274482319
zb426ffa9d9dd2d292981792cecdaf99083beca21d5477249158da086ca912ea7cb0e506b6cb620
zfd658a251d3f7224d890ee5b5ce2a63cf38ea6caf1d9beee1db84d6f6db8a7231474bfdc59124c
zeaf80b23942b5799c2d2312bb8ea87c81727e836e3d0e50e85a9cb4374d60ccc0ee4a3c32dd4b1
z1a417200692f5faa4da8fca31a86f01d1ba2b48c06cb7003992da633cd3ae25e01cbe559735671
z37871e28a0f65b1265430b7236cba1c29e6b096c5c2665c95fd3d8ca52a1902f654f20566fe9b9
z20a9e04502438155949753999249ab0593d443e17853024b87554d50033d561b20266f23f814f7
zcfbaf57642a0c1c51ec83efdd8668a85f3330b06754c6f07d4e66acab5976a4134efaef1884129
z6f95543e357ddd6f455f6885ce7c14f38ac3ef4ca0d7b55e5096c2c0422a44a669b76541ea3788
z7920b1db99deb1e1307d5fd46d48fae9c2a6e8be980918ced894eb6df56bea969238e4503c4a93
za03bc325c67207c9696ef56202225819b8e406f834b88d3d477245e45da547797ee9b4a5c104c2
z685500937b620c5e78f99e83e7cf053f69b5c0585b4aa4070aa50f831098dc92ff2d1a9f11e053
z706298c985ac05b9a5123ed093676cd2f18235aeac22acc1706ed1753b9a8be03c0689f7af64b5
z6e043c708b55cb06934c8aaa8f45c328d586f7daffc2e185aebf3ef2d264fa22c12872b90883ab
z59c35b8c62010db630a53eb48d788c2af384ad69cf990de78eb3762aaceb3f1dbf0f0986bbb28c
z1f50cd45b44060b5833ea9bee55012d72f1abfbad20bf38a60abe901887761d31d603051d41835
zb43582ed6e209227001212c14db219dbc8d9c1c7e8754da3e1ab31af1ae242a1ed63bda6e8cb29
z211b9e19e1ab68300d00bf82ea6b744aabd28358b65e4eecda8b75ec235ea096d07231914902e6
zc1ac894c936f9e89dee2ff1006012113a9a9d2923d031f73d7869e63911f3bb3668ce1e9b7661b
z17b5add7827f337350c708e13cfe3952686a6fedb3b8f97a0a1ebd9796eec76e9181d994edb042
zfb895cff3849fedcaa597d9a8ce90e7367903a5e601fc1cd06429b27f927f7773101746d0b30b2
zf2df6883b3bae252ff8cb3a727095b73a9f55a298614396df28b2193d73efe8544f30e2965587a
z097dc421a1473ca68c7239a1710e86c0ad913676791597319abad8ed886309347ea12246196e77
z7adbf0027274c6a2579240b360be215c9d2caea6638d5c3ab6dcf45ad00737577a12b2c2e45002
zb6b5706a6c105380e8568b28096d38c9b7572bbcac69de34173af8cbd84013066e858df0876cb2
z59dd882065be2b660a465002c8c2e6c02e7797b4a94f0a0bf5943bd711c44d4f597c98e5de3887
zf1c554a6935c9122fdc507ce59a5c9787c64f29633c60718c782c413072768b83194d18b0b2507
zb1b48b0b9bb4e02d28ac5430f750658a7a1932d3a7716b60b43a228a7d89e3c37d438df5bdfbf3
zae49568ddac55e5593467e75dbbe549593641356d74628eaad0a68866734beb2ae1f5008a205de
zc9000dd89ed2e3b9b4587f2196ae56b3aeb0c961205c99bbb72ffa27e8c39ab766958b361cef55
z4a8066215596b34c66a09bd8ed91d60e3d10b45043cb9db82852c4284620047fc79847aa5d5fa3
z27c3bdfe3d4162ecc9adb170d01cfd6cc2e7a97b7e8ccf3676dc89df9fdb46e0dd55035d64d321
zbaab4cf15d5198ec2bfe9a81b99ef7836513bb6a4f562fafc724132ea4e3e181b39cb368dd06c2
z9a64fa84d47e66352bc67dd7bbc10434447c4c7f8b38e882066f76b76f77805d829654e30dd095
zae633679b29591a281e05e605d8accd4d0add5eeb0ef399efbfe1668dbb1607a024f095fda36cd
z6751b9eb7ef1142767cb819baff93685e1dae1aef998b9bb253a3bceb0a89e528224ee98cbb85f
z0c44c7dfa616a4e0ed2869c7f6ec73d87da480ba15ecfd9b8b887977ed31366f19c477a08c14d7
zd70ea1c6e082ed7bf29dfdd18509bc11d683f63eb53ace411576014b421c3da32531234d33d87f
z4d2dfd25398b0b3256b8af8fc1f27fe45cc1b8d441ae7b4cb4a1e5f70ed807e68a4e545089afaa
ze8ff608e5e972d4900815e4ae730fc304dacad7fe5541071453445e73e8553b3a83abcf451ca2b
zd82b2287755aa045ef60363989886dc5855f3c8e24784d8edf9cb5a63f8862a4f3d4e60deb61e9
zfbe6c9eaadae9d9eba2ab3134cdaa09e00383f7632f6a1ae2d88ef8d6f83ae1ae2427e53faf12b
z4445754b0db6714b471e978bd013af567853967a001da98e926c1d8d36deef4cc4116080019988
z4aa8409b2484fe0ff74edc409abad02b1e334ee1f2884f54074f07ea9d2b5b48b650c15c623dae
zae1983482b6bb0b417ba51a093f005dbaa1e755a8ede75c1c108623de581431c991ca91a2b5c2e
z1f64ec9392b1e8447d348f627f749b260ad6f38b52f2b86c83ffb885b1190d9c048b2d2b753902
z8def430874f1076600a89ac20a75a10743c09378bd95b7c4e1b17c0a1dc8db8f648f7eb15791f8
z911d0c1c4bc11099685db920262ec718562417c5aec17e0f75bcb7c1d15b9ef95ebf0c0c94ec45
zbaf46cba0cc498d791b136ee945c2a268b4acbabd222848c24a816aaabaa9c45d3a39a716f4892
z35961a2af7b41e10991dfc62d1c553e08d9166c1f661910ab6d4ff76984497709c3c9ffc4f94ff
ze4837b484ef2dbf0dbebe4c85774627770aa30e3ae2215a5cb37e1052783993e9f36bac01a7c19
z03e56f875238cab264b4611cbcae7418092eda7bece9087eced8d35f5a1672dc27005173d848e1
zb151bbbcb31016217dbb4b9ad7ab57e93794f5e7f872e4c620ecdea85f26082bfa0a49277441f3
z482e00750e7d45492212f3f9c9cffd38fd823012a800ef929b4e2e87db1061539d0eeba2c340d9
z73ed90a28b1ca02ed88430419d0648da5d9f18a2bfa0110c38ec123df9119c703127c43f7bacd9
z9fc583b6acf3812b8d4378d8fdf731af5d0a735c4483f2551146004c2dd3d1973a05d21688036e
z606a0e1ed53290c884476000860c32eedda1ed3b54e5553869aaa6eeb7c23be8ec985d86b47218
z2239cf635ea65bf8c45852e77804c10d36242e6249e4ae330e38a0c31dcb4f68a8f6eee1f32974
z0456429436fc35b098eab15c117d65ee8f56bd861cb6e5bb9713bf087aa3d22647b1ff907f9154
zc3c1a30fb7e582a07ce096cfc90558950ce7bc1f6b134a6ac57129cde70322d4ab2ba01511308f
z475150ecebf92844930764ee6750cb0d43af972fb33c63f15dc884c94c561294e337470aa547f1
z76bb68c8126027869f89c85c635a13744787cd478775751e213ca9663c23933af3c811788c473b
za593fee5583921b9a0b6de25807caf6bf25d5657ff72a1650496c84cd0702a112864da77f2f592
zafe866a4ad61ac1782e06efaeb85035f366760258a735dc1d5ae20379a954ff831c89aea5b76a2
zf22a84dd7da8e533aaecbc1b8e43d78ea60c34ef712f93aed19a68f263b195c47e1187646b70f3
z6fc673868c7cf5955ddacd7533287ecd0b2b6c44dfa4a6630b80d336bb8f0065da619f016cb733
z785ad77f603a2881d5aa839d1a33556490a499b131f91f94c9fdab04330e51a161743429caa9ff
zd6467b77ebefe4c9f763101938ba26593197081c4a899e6bde172314b5f55c65f7de6853cb2c0b
zda19fbd5ec2044854bf8eb9af403f02a94d9f813249bc0aad7d4480f02a162c8b847b5f6357495
z46df0cc569710afbf671fe59fb06123194c19bd7261f028067ff3b5f189f08ced760bf87151342
ze10c239b7f4cbb3fb50b41dfbce2e9b1e80df93a5fb70a7c97728e604bb9e2618ad317138b31eb
ze9bb1a135c28b5a7ce5163ce068c21936edbcdaca34796d428d3217822874226b0ba0b8fe3f8f3
z541b595d061d01fdbd6c561a382d237cce8df5bb6fdca1c7c8f7667332c815cfb39405880c413b
zae81b7dccd41bca2a08a4b600f0280cbe04c1c3c8eb3e4757a6be78f68553e7c6ba7f483f93f33
z0efcc00440aaed1875c0c3e42725bbab8a0b13fbab0b14e67ab21d7548c1a9437f945d1488d677
z1e84af73402d45c1b5fe29fada19f91194e2e3f49bd5519a5b58ad9358e67c06e8b4bb52c61326
z0e21394bafcc66802ebe2c8b2f128d7e5059f77876888d1d63dff91d2513f951388772ec5f46e9
z53ac1cdbce936227f0e0fbfd236e87968c69d362908a4337ba32d8402b6bc7beda0ed281f4904b
z61f4e5185a65779bbec1eec155e4609d67b2a93b92a7dbed2c053acdb311da493041a34cbc9d25
z69aa02bd5e26b5f03e0af7e9843c4662ceaa5797a59d3184300f2b9c9c0736f9487ec4cfd483e1
zf036ced41709a520562de9250fb6cca466d4ee8934612129ed6cdd5c7d5ced4f1a57fcabb8887a
z532f5f1c82440ab17200b26325d6228d2c4596ff85b97b9cb545d165d9e97a0fa1e3a0cb59be93
z161467e2f2d45b7dc0f65722885b97f3e4852c02fef37ea15982fcef35693bfdf8f81e4e89cda5
zd2ed6b751c1d92e2056ce2def4e78c26bcca9d678e7abc2ed120b06b4b65b33b4ca09e1f1ad2fc
zf5b0f914f282623b1ed7cf85562f161aaf7d9a6bf408ceea173cec53dc62512b0005cc669e4e8b
z93fe57dfb74600dcd48c8e265346ce6ccfc07465579bd855d18fdb0ed1d0c1b130f10b800be094
z36aa97bfa3b377fbde866cfde99108553a7e232e1f8a37f3d354262ada51bbae2eed5b1b19443a
z28e3744fb320acc7c4ee383180b7825e61e3ce0ab427d5942e8cf9df2028581eedbb745b4c9343
zb4c0258e84986bb004f7447a456ddf84bae1554ffbe59848330e0787d3b9a5c72e9a91164d0987
zd254edd0b44c1fb85c17d152c8d99e956e88174260ae2236d7781e69742d246d6db57f41a0acf3
zfc67fe71c8cf06e624559230653582ca8206353fd054cac0a2673186a85c999811b04285151e69
z6a58e8403b599b6a0ae40ffb64bf91160c1a0cd3d93bf65236f160e5f7a3c0ec7d34f964c0b63a
z8048b111f3721359ac2348bef57bf7ce1e182d174bfa8fa794ae9797101888e1a56e40413deca0
z57c4c1ae74efeeadad1c0b00c0475c0f9561aeaa3184579f7e51afa4637a4f9beaef5cd1c0d629
z652700626e3c5d7a55fac6ee06902e6346303a8dbca1dee5ebe01901a297aa4e48d2ea7af995ae
zfdb20f4cecf019c28fbbcddeed90e6e686fe9957ff8206561d3cb4c7a14060fb94991fcb263298
z7c6a7fc076f7ad3607a034a84e9b711dedf5eea871f9d14bf2da84e0cd4796dfaabc8e3746427e
zcee963695d12cb263550055a3810a46ab991f290e731f9fdfead6f792c332eb85e3f89c46669b5
z1f0d64eacb85aa34ae2c19dd6ad884d8e8eeb574dc82acf3bb051277a1bf2c50670e4e550d73eb
z4c425b9398c5989e20e1703180e31f5ef60f6e14d40bcd7bec96e797defd242ff2570db6ed4aae
z4397ce7cb40bdfe38da0ed460fc451afd7127a4f54a59937b31c43cb5c2836a75879f5070531d3
z0cedb3ef21d84a7bea29e48be603429fea2773a665596919f30d9312e65f04209f8b77882bb964
za97722e1be39e1ae88aa9d8eefc5cd382f3485ef2ac4f6cb6d04a1883b181519ae79d136bf9b96
z5b1d6fa29a5361da35c4bbba8e0080e506233dab9c6cd44494003427f2097dbe091dbd0ef39336
zf34a50033155f3a9f63f910344453ca40ae1778b2266d5b0238716459f255803bd2604e8c5acfc
z33ce65369754d9dae8cc2ed920f6a2bd298a1247186fc345088efc8b1f07aab68179e8f4e13557
za74f3e78db50e65bfdbdb7fc9c4f1e3da30190c0d274500344d3557fc5b20bbe5a8cf75e277740
z0724985fdafd1dd876f1bde2e302381ce27466fce48b92670d34124e78450480c1aea4f3af535c
z3240ab10b65ac2db7b732ffd40e1afd4f3587e3bf53eafd3f062a652f886f10b121c54c4c2ce58
zb2b8d616712ca30e915c405fc42a2d179e65845c07d3321cbac2499c762fee51e69051a34d9cee
zb4ab96a60cc71e84a8225b149627da697f3e90ad28ed8e41edce0e5ce210d0ec00fca84815b4fc
z9ec757ed33ff4e03a3366d4c58d3493a30e12bb898849434455b05b262ccb0948300f17dd92b65
zf5583eafbcde07cdb4f74f51bebe45de87950690e7f6fb978b83db08b206162fcb0293042b1df3
z9e3953df4e908fd520c7796bf75ec1c7a98a40fd6cdf8e29593e750f19222aa738220ea2d57c8c
z30c16e19c2606fb9ea6a32eba4bc9f06d32cc3160185dc53e9131a5cc26f95411f643730982df0
z0a9048450132485ead24cf4ae26a0a3ce91871d832f81239da4bf594a5bd8bb889147d2cffe37e
z4991a5905be54b2d5be128dff1c6b06a44ca78ade5f5ffa5c60264aeaf79b2a11749d96d6c18f3
z2956dcabc6e07adfc6ce937a06f99b7b4a770fc293cff69780c9cfacfef101bbaedc8dbef78796
z4d4dfb1bf133653628c0f814a3a80f0cc594f4bcbc743a9200b7e4f5b55fcb5ef9842b989a1688
z744f1d05bb2f8d5bb6d152f0f08a6581c27111eaa4a1f3b1b560189c58304ec52ac2680e1ad935
z56a6a7ec9a2fe2c3ba2d653eb56593bd3c0a42faa6f436ea7ac6d417a57a59e2716fcec0209f20
z40a649bc0b27a7aab844ace49af71a5b6b8e25d71944184b469f7eaf51118e2b3c5a0b91f10051
z7019ab937d1a59a6257fa3a8eb73d7483824bbcb643235e138a5213ac8a6c71c2f6e4fa80f9f83
z8a87d4800dd6c238247e9ce9bb528244d7ab0f521969fccc639ce31ecb0e30484d7abbc3c3cbc8
z45ca10b20b2020dc47f47b90ad17f0e9f86d173d2d08d5f21fa6d69e58c96e04801c5dd3d7268d
zcd73422185b00ea79c83a7278f37e4a0ada2ccab3e34e0e982ab6f1e3443859d466f60e16f0af2
zef1d84a891cbe95e4080235a13585e64041680347f72322774c246926dd8d85fb5c1daa000ae14
ze6e8ca1b72fbf5b5917aa2ba13892e3948c7fe980d928d137ca580a381471284c4b07b6c0927b3
z61bdc52b9ee0ceb4e34b2fff18704ad388e2205c8bc6c8264301b58caf9190db22b0e31687aaa7
za06c0225ee93f60c3297e152baac742d1340c21d7db35516441ea53a7b78460e6c19e0e7cf7ece
z6bfa164aa6b67469e31312d77d0cb801bcb829e355415bcd1c93630dc2746211c0b94ec2f3b506
z4dfd4e474dabb46fd31d90dd6e1f90af2fd55eb2f06b5decf2de4721ab207a9678d86d54b767aa
zeb4378615a65a47e6e58231604f9bc0fe6f7b276409020ca6a8e4f2bf711b5acfb7b2f7b844559
z0bb298679480215051229416291e8a18d8a726f8048b150d862507b0bec0363f5897e95d2501c4
z8e22f4e127d8316f73d4531f62343214beeb7089abd03f1a58a30f1eef27919416ad57cec36c80
z0033e91a5c9bf5b0a6ea790e16dcf54b85fe957b257b15e833ad129f9e7355242ffa8ff450f320
z463a8c420811dc504e8630420b72891291ebfac6b737441a1167a75089997d4b3788f24c6a83ed
za7ff63c4e5f815606eb0128ef735bfaf4bbd47b569ea24ff2662014232b5427baa143eafc6e75c
za58cd569363a5e427d1f8bedbc31a80908744777d4106285e117bc3a5dcb494f4557db8f3e9800
z5f44b219cdc7f318d00c10f6b7c8ab1a430a88b029e35ff967b57abd62ae06922ba76cf0d4c88a
ze00f0796b7159ce1279832fb9dc5965e3db13d6d2c0a286367258ec5ccb2f3dfb33518b8527f98
z3cd7c1d9ab66adfd2827283860c5371ce58ebfd6015b7a125c442032baba4c01c73b6e3ad24e2d
z2e4b725a371fd55ebf92370eb4637c094b1dfbe589c4bb663009680bc9666d56e3c24a7b00de59
z95596b9bf10c3b360acbc0e0208b9051d82ea9076deea848e3c35027c0526531c5c0456b9d5b6a
z2189cc0ebdd1da67f01a449d63284b0938b881badabf7c0153f3b853fef126c3065061f808eaff
zd1613434a41dc56337ac963926face0e33b23c7de3c7967d11b2e5f06688e09429843d6dca7be8
z51d4e6455205e8c6244c7d10b91d7b4e1570b3860dd9ae23349b73e6e142c02a95e36e7c8298bf
ze65ade6903e36468a5c8d5fa1d8a2f0604708583bab2393c04f743fc8a188f56af5fce8a757095
zb98b799a48f077aaf4a5f8719cce0a59eeb6c864a4f553a2f24629273112f4e14061350f3dac88
zb9a5eca5d1b0eec22233f988fb0a48b17f7b416f88eec2dab7818d521d7d8e448b2782129b96b6
z81ab3d11d06655de8ecae28c582a5a3e4adf4618932b044b61981f40d78455a528c2ece37a9558
z930d6d41faec9a6b4001c8723fe4ba95f78913869b338f0d6a21c8886cc27b540d5829c7f1346e
z2a73fd9c6cdf2256332ae58f0aa4a14907e74f9da1031fee0fda4fdd7168cfa8c3078ddd5dd25a
z8ca430caefbfec1777cfb3b34ba3836e4a6af8461c0cc21b86062bd060a7e1a4fe77159dd3810e
za879d2a2596a12aef6bd77558d6e416cdcadf55552d3c87cddabfee5f06493d821e32e7e1533e0
z556a672ad8a8724664f2028ab78df1fc19a316a354eabdd45c5d84ce369e8660cd370be44e9a20
zb4edb7f8450363d5b76640f427cdb29e7b9c28cb803ae4cb6924424a6083ef0763e12a47f148c6
z77ef5053c188e30f56f07e3f9f8ff8e3d5ca3cb1900b301c9156ebdddf338c38737d2ffd52c58a
z53d7ebfb783a4536e0f29dea7a26329f92eee75aae51ada6e07dd7b75eb32457b53477c48c9daf
z7b3a434044b33b67ea80037be1d4eaf0afd0eb6088039eb3e6675648908254be44b07a3f18e8bf
z196bf61010096555b75e8cb73b67c3d74b289f3cfef35c95d996208660be2365f6258947ba0d3b
zecef9f73689e29f259646f9e3825979d8c768279e2e98c6ccb3feef636be0cc7182e8d465de057
z662fd286d3d42e1c82cce99a09d558b7247326046c94360a12bdf09850db49322135dd616b1f89
zb73002e923fab8df4db28d62204db20de77047555b49e8f11f1bd4ea309d81c8eaf75c59c116a8
z5257d2ec65157b427c77a3530da2fee80ea104c82b2440e0b011356d37053a9d84041af967741b
z9046c7c1fb434269c4dbf5b8d93c9ffb9aaecc064dc2ad1a8a41193a8376e5e03459c5c0378241
z696ca22aa3d5e825959e677a8321ac28c96c7be2ae77065556d62b3545f91a683de62447471a21
zb3a165c7af79ae20f912c335052f09420ee2d16d4d93d23c6d2890b56c22e564cd5055cec5d011
zdf49ad61b92a69ede47cc289dc07d4dbf79ed01bf8ebf7a433299b3ba4831431176b7cd4271dba
zff9b78ed392191011cea1478768a79d2f3972560223a9741c4dcf4fef30bbea6e6b088bf69857b
zf8a9e9976eddbe4a98afe13cf94f10da84a983853f80d584e8439400f7999fe42c575965b91010
z92e1b9678174b3ef67234891f3af7358751c18dbb765f5e3f50583a9194f5c72a611bbf71ffbd3
z0abe3f84ba532657c0400ce47944d8847c5df4bb27c57b961229e4eadfcf20027fb30563de3aea
z1fcb1cbc5de168e2308a7ced78871658d6eb99d5bd033c92e7a2fb68eb0ba0cef3c80ffa32001a
z5dad6539c0250b5fa603cbdaa628131211b2a47c9d89ecd7b9611d659e4d0c9eb910fc6c8901a9
z4032cc25b3f86408778e8ae91f7d06039577e967408efa71034cafb6d8acbe7559de4c19b5135f
z928dcef3cb78cfb6163a712baa02a9baf2a66544ae6d64af6c1a54cc1786b54d88561b8480521c
ze7a9f8381176af38b5be22a2f1df2cfbb4eb1b1fe68b6d74cb0aae3263867371ca5d220a17e76d
z0d1f58d79e2f29d14243f77505a2348f5e66713b3452f45d4fa4096bfb3de347068f57b366831f
z70b65163da72e0253b00fe2df6cc1a318fb80852a3a2a5fd3ab11a0c1556f6360d0ae59f841a34
z79da1ad9ab0c5e2416d555eb79b30037465b83f32ff60abd9088c60264ee9efa3280c60aabe9e6
z5f4afced30827a1df396a978c7d10858143bbd210d07f72b9d22b94c1aca876a8c0790eff2f5be
z4ff79aeae9eb7d52c38c84d69ff55a73bd4aa545437de93308e624c6dc2dfbc5f883d58d4466a2
z67cba3a613cb1aea24e8d41d3fe227cbe4ea027d5ba03a4773684ad6d09c319d94b91b4efeb772
z1be4fca3ea6d0c7082726d78b474d33f253c0010849864c8dcd0f8adeb836fa78f8ee2d0c287a9
zca9dfd22915e6ed854095136e3a4b1dd8b9e73fbe39883c3c1c7985185581bbfdd0134d06f6821
z8b8e5244451ec76a6f530536386b1b1d916c2532189dbe4f829a38785dc87d38acd1209fe3bc8d
z774ed3e7af0ac747dff18dbad7f117b206ca7c71d6f134a46fd51d5b1ab6e30b325e57296e4729
z6bbb0d4202eab9e023610b6a044117130b123b140c098e502c741c4b8c53411142ebf3657e949a
zabcaeed86084ed01ae3fc9f93c7f0e90cc411c8f2ba926de934524af886eeaef9854e72ed1bce3
zce40e09337c15d99fa349c3327915956a149fd0e80c79df93b03eaf2c6772ad3ee2e3a8a39e1a6
z22823eb969832731dac0ee62875e7cc4bedaa55b082136e79ef4ab06fc0a2a2b91d7416fbfef87
z24964dceadaa3506845f35b2e0498540ed99ee6b2de5d39380161e1e86d6f2a98aa4da34332b92
ze72221f93616f011e0b3fed5ce34dca50c61bbe7f07914a2950d7e753c36a4db6339c87d09f482
z9bc35b89fcdd225d87aacefe3a4c77920938009fcb660dddfa2cce2eff5677fd6428d9f2fb46d6
zf8d36a1c6a1142fe728c43ae63ff8238e39e95dc0725a500b39b51bf6856e8d4bba152530fa6a0
z730b8c5d72450b5ed53a6a787eb991988856336ce188beead656b5b8a3de95f1d8a86e61abda43
z82081a84940f4346ba916ea2e203ab9b811586228dbb00ccfb8bebecf5b73f808aaf230860c1b8
z23d24c62c92d5470dd5deaa9632baec21c8a3aed8eac69262e8e2817e8cb428e20c08c57452341
z9faf7f528c34f2f5a7c4d26ec568a3b289413afa452ff3110ac4ae11b319233e9ef775332db6f3
z4ed70e9369d2fb5a2745096170f6407818d954ef365c32bfee946733855932654fdc30562006d3
zb85bd438cf808d982f92e86006d2599bc3c8d21bb941226f4b3964d0ac9abf0d38f787215bee13
zf2ff5b243dd03f28aff8c6109ea415145be28e907db4b4c233bc211b8efa85ffffce73d951164e
zc0e1569eec6f46da669e6df90ea860f2cb839e31c06746d1ae4b07a4990f5b5dca4c725d9ae5af
z5bbc1436635ef579140ff88e707f6f289e8694b6380fa0668df0b9767422eab9fc11407e1cdef4
z1ab9ca6d4879b16ca9d4069ed862c0ac92b95bdc71dcd5504e87eb753662c175b7064620fb9ea6
z166d4cea5260b428cd87cc7ace68206cff042c982f546120697dd577e7f2ce7ddabec23a539d5b
z5b10234381fcc818610770d9be33fc6a20c205fdba9afb3d77aeb8a63587f7e77febc5ad52b58f
zf540f1a24c46848a5687229ec40c85c1dd9f84fed5466d62bb4377d8d69e5436581f004ca1ed6a
z01cd5cf6d48d43b80a50728c8b0975a37f8a839e4f4d637f5d9117b7de31311ca04ed89be41a07
zbb989d1ded4e0bd5a9d6dab9e4f830f9438b3b7c331a8b174a86cb77b7b53d90b689b684d45069
z1d0ff66d3760e566632ab03a32c9330459fd7fa5907199a6ad5b0fc1f90fb3c72462a479ea5ee4
z7ec65b34936c7ab09975c604abd50c536454fa7344c61fda0960bb0712067bcc97bf3089606968
z8863a75905aae201aca11bcdb39a7439489b9c92047ac1165a8092283f34772a97d34b4a6e1980
z8c1cf77c6d139204166418b4f3a9fb3e5a26dbe03819cc6ca297b9e354c8166572495ab5a7cf89
z9af37830db469271b0240fa9a3b55c7512584c1a0332c396c7a3ae812cbd7c0b5c67fbafde214c
z3fb1cc0969075eed0bd883afb4a6a8eba179f774fc94008cdd71c2a76f6bfad698a7b1775629c5
zb5910d197b861ce968d752e78c88a22c1307dd819f4a355bb3bac1dd14e9ef799849b5e7633bc5
zde8d7cea7e70fa8d731ff0129b81d5a7079c391f89ca4ddfa47b42a25ad852afd44a1d044cb099
zf5368852115cf715a189b35315e0aea060cf20cdd499b804b4ed5696decedd38eb1dbe466730a3
za95c1e9ea049c2a9feba9ab0530a3df5ccd5d4747bf279dd22d2fc5ce506fff225da093f632a12
z3e996254938437daaafacfa8381e294f286ce85835eeb94ab0b5bf634d91338672497371c0dd99
z3c0ab81cb634452ee059ee96a003f5b4c348876f0d9a2a347908903e34ab502ae22ef2d33e5e82
zab36177408428cedf106949c7b9ff5ffb0b676520bdb86f97499b571ea9e1e7de418001bfaa00b
z77513909f4130103ab908e1e37d97fdc32a82a151d0207dbf899026014b026efcf4e870511e2d5
z7a43467cb54bc50ead5169ee1d1045e6d48e40c66df559f212025fac72c0eb04b0dd32540be8ac
z2c155b3c1adb1dc5f8ad3711c23da5bfccbfc7c65e7281eb35c69ed841ad7480669d49dc13e724
z2119d88835052cd5caa2fca58d6ab82033aa53e3625f846c514507cac6f7dd4f84bbe60399466e
z009ec0965a3b0f4db44e7a84339f7183a1313018d768dcb8e48a799b1f524198cec217fc4f0755
z7ea72a4e249c34301a7bf90ad5c8486dbe6ade6d14f3b0ea15a74be15dcd2e1319881cce5ff23d
z549e558f2806f3fbff6cce809930efcdf68ad5d15e1b44c25b4b9a042789f4834dab74dcc41c80
z0daef10fae88fdb5183ba3cb20f224d7fd3605786150d8fa1b306ccf6792f340203209f8772660
z817553e123e6212ef8314bab83172b988268f8e9d984fa54df12120afed77ed0f33003e6073d3c
z894fab14c462ad07282699030964cfb6f2d9b33d4e616b14ff2119b1db1a78bd9c9dbddc52e15c
z4b6974f60d2a81274c5e449bb2c33e0e6926faae12845db4887decc3131801bb5fded5103d2c2f
z833f5c102b6e99f7c4a69958b71a3e0830b15e41665a918ebaafe4e01967c9066994bb586b6c32
z2e5a8383866c9bc3c3b9dec5aec4da107c9d1ded31de3f2dfd90fd5810a3f7b6df5a23920dc2d3
z0c1d312d86eeb26fbf5ee01aa8bcb866793962cbe31b7102add7747274e2fcc1cffc342ab08fbb
zefb97b32156bae6cde3bc0311a80f55a01ea48c53900a779f3ffbe6b5e04274fd2a3b07fbfba70
z874de7d6ee98d0e37f16e9a56ef1349abc9de995c6e1d04b986beec8afe7bc529c1826a736341e
z9207ab534b4003dc91e1ee8db023de4b0d456570ef1a78410d1a46e75ba0b5a9b2e723475989b0
z75a18eba95f3c76a8b77afae68129fc74fbf2a9516757a842a176c1ea6e81e4da952a99d6fb3bc
z76b2f5fbcc636dbef8f36fdf7e7c6422bf719cfbe6796765a47d950299d75d112c098670dd0d23
zc01405fb05e32b144e85a5e13b8027fc83d136706c70d0485a9ee5dafd6cccd299c779d4b0e537
z0400ebb8f74ce649e18826ac8edfdd58fdab18d5b77de335643ed244f7bc0f150d2cbfeb229b2f
z783b1154d62188aed5cf52868b281735330c4fe3dd94ae4571f060d1c1300a29c4df4957c2476c
z697c6a37c32d84855b9fc3083118a105df71931c98d3c449bae64df3c22d4214129eea77890d64
z2305531124b36a757462f711841d328226d3d1c0f654b031322ed410cb0873694a33308a210a06
z51aa46e756eb9f28c0b492c74ca4ea0a8d6226cc0872dabbb7116b96baf696526473b0133614bc
zc505d2f77a0f9d875be89b4e39216400ec76f2d409df5f7daf33d055d83d3269ce7ecb6cf2d296
z5302ac90348e2241d8294e334c17e789898ac4cb629a267729175c3a06dd7f382abac2903a81f9
z7273a5c63e724c1dff1e38657d3fca3250bcb43eec73a3942877d0bc07c27c7743ffaf73a7a23b
z26f0e6b211bff6208399f867c5cac9ed3cc3da4652dd5b579a16675735ea0e2e371b590a091f41
z410fb0b72b1426f11131e685be4126e4533e25bdfd06634d7f3112cd3bc93de0ad5e8b6a863aa8
zbda25fee5d4d36e173cc29787c620eebf7767443dd35ac9a7b5802e00000732d24ae4c34132881
z20d1e728acc522aa2531f94ea15fe56f2f4e3e4979d2e76a1c3b5a80bff6127285548c8fda929e
z8228b59aae7f8c60e03eeded7020c7a77134d43e31e4c58e2c16f1364b5006ab3d6066e57d8c67
zf2fd5ca0550ded1d2bc5af9dec12c0f2d3bf25ab7dae39f9e016020fb7c1b88ad8008c06b15d35
z80476d7f4fb2e86ae674a62e95f3a3ca1d5dab9923998978be00bc039da7358581865acc3aa6a1
z7bd71f25bcd52ac9374dd246bd5379be7989fc60a5dc25ef8a603389ebea6e3ebff450f806e174
z6a9865053dc1fc8f954623bfbfb2444e2ef61bdd15d6ccb5994286e27fa2479ee25051055a9f39
z3c8e7f8be5a1b233935ba1f09007153cbb11ffbfb0d3397f37cadb96124c53a6e5223290ee062d
zf892d0e0279aaac09c2d1ecac2640bc5d508c5477672b645663db5e74185ca10e02554f670a6d5
ze5e2d9da9966a645a995796dc2d5ca100cb9a03ac39cbdb1ef8b0c7fa39c33158d299612e0781e
z96717c7273484ecb23a6369387d27366d8f87e37b22f7bb858cc5cb94a4a6c6605edda99373493
z5b9b5cbed96dd342e460159e0666ea85ce1812effec1f30a4fb467b095d6eb3e7c086b8206f0bb
zc90bf60fd2a6dee2074054bd0469e315a83e969fced246184686cc8db25035fc7bd3561d969c1e
zd4a470d2587f37367a44360e03c0df8ddf971ec580359c7d37614d8c90180213aed8fc9265aaa8
z75722a6c6bb1ec83a807dbe1fdcb274174dc8a70dec5d889d44d49201bfffa0bb56e10d5ecdfc9
za8242fbc34e21d11ff7452b17fbf3ac15130008ad1affac304763d4bc0f28f8742cfa39bd34633
z1942eeada4dd1beec48c35b338f9113ff5f333ca93ab0c0c122ca7cb769e9f1b21eeda2dabd43a
zd9a7a611f3cd9c0408b86e6772b9eb1346355134ceb6655f19444341e2d299d4d93e424d8c24e3
z6081e2dbc530d485e28bb1b1eb5c435be18a16b7c201088cc07ea5e257b2e2df64d1efe65384f0
z500a47b0b06002b32afe562bb1161e01ee25a17c91b1566a69d32fa541cc8a064261537d977fe4
zf2e821c08d7ef26a0a95bd34e212e5e298b6a6da9e213afcf0d9ce478257055dcf9bb7ea7dc28a
zec14a9798fb4d66ad0d0a1ad0c2a5e5021b2675108de4d5127d3bfaa8fac44b8682a7e43ecadc6
zbfc7ff7fcbb1c655feca9e87e1fba2a562c63484c5e9091f21fbdfa88eb654413169050de1fd36
z4f0ab58439567786abfb8dbd8e96b298dc4a4a2ce9c9f77b29d769ac62360f65fd8aeef11696db
z6e20870f49267074d294b06bbd31b34e4f8665246249f5ef82a7ffc05a84d8555eb1398fb65a38
zd3f4faeaf53c14488421219bc30ff324ee243371b847a37aeb8f81b8f00de51c97d60411dd9d71
zd63cf366fee8a5c7c8396c9ef281da36762695d9033d8102dc0c8a1fb422129fa9766656e0b9d7
zcfc6587a575ef406420e91d4f27e1ce6cd3bd55fdecb26af8d4fcadf3271dd338b95bc436acce5
z46f51212502d6b9dc8eb1715021fcbb2006b382764bee6ca6ed5954f171d134da80bb1c3f67dd6
z01eecbcfc150c6ce9553c4276efdc7258cd6ce2304561b2a4d31c482687130144687a72f4284b7
zda799d6a4f1e36fcf75100eaf1f7c9e8c0f33f37734dd8463a033e526de965dbb5bfc8a3aa5567
zf1d03e85fb204c247dc4e14f380f98320ed8ee881b05a19df69938336cec14e194da6b495efabb
zf89dc6c96f3f42038e5b8b2d3f883c1e7246ec9a48257907798f0b71d586ed7711dabb79774cb1
zd54c66a5076c3f5eba05680c168caa1fbba60454b1e80c739b1d70ef740a86cf0275404b761eaa
z0ec383c2b4e2fbe0c8cb8cca0dcad95b357f7a215b2eeb0fa04bad13f3d7bf524c71333ff81d79
z626d6841fe6f37fc11683c8a6407b16b04f950a06ed32f000186dc7f7cc339b449c44d5030a8cc
z7b64ef9c893961bc558f5643ec18c6c2995035ac56c82abc5a471e55b101e4b5444ce3bc719be9
zd285d4ffd0edea8b809ae9685eaea22cd42392186d8247c308410b3e55fcaf9a4f263581464404
zd80070a0c461029ada0e60cfa51dd598631856abf0842f7357d5c73b607e81f53ef8888ec833f7
za7e6531d95bd10d81447d2ce6a2a845bef49182ced85677b1d6279ce6750010799f906269c68a2
z24e777432b29f5c2cb0a0e9d3c06b0f540d90d477b24c5922198e7a1f04ae7dd8c0526756332d8
z12f9de5f56c3d1de35f7303ef4e5a8264c294e22949fe9ecb44fcba4ef7619f799e24a4b70f846
zf3bd3a0075606b9c51d35f0a73791aa27d463b07a94b5a24f6c1917ec4e1ed0d50723df8440aa4
z511491e366304c6cac26f5db07855b9afc70712df38a7493b02389fdfc7b994908f40e1865080a
z63ba497f3e483954a24bd83fb8b3f7f768b836e56a7c789fa28e6e38317765e24ccb13d1e2749c
z523f1473d4e59e7eb7ed969670d704b6c9f28ccd5549c91dc6cf6bd6c7dfe3de2a42327070ed32
zef76c232b1968c80dc54d7f4b455f2a11f90855ea1e0bdf4fd5485606a44cca25c1ea4d6c045ba
z30a91569d0ba4544b009256d1210a51fcfc77dee91b46ded2ee7c0a1d91cdbcf54bad02504a793
z2da088530d8966764b3df4ca332fa1b6eb85a7a248747385754dd7f22a81a51f68b715a2e471db
zc82ea28253c22b4603fe6eeab22771719a04b486b90443da2fc83fb66432437d88b567e5b0e916
zcc7a45a43c50083f50448134c842b40a6064f23aa794befc9ca59e915d30eed5c9f552669738dd
z5243dbd0d336db943b23c6b8dbfbd051cf09585f62b0a42a0d6dab8939233555e4ec55ef71facd
zaafb553afcae7e46fcb110c1a64e90772e055a8b425564055f6c52fc580ccef6088ff4b9bfd90e
z2a531352cc1b0470cf8b8d8d59812e84e9f3cf085a6db3ba175f15a85aa8b4b8966d4aa5900798
z7542a63318a78eabfc9c34516eb459d52f64f3cb40c58482d6be2a6bf686c21b19b3558d3747c7
z34f9ee31a4c6277ee2c995a47da9e4c571a39ae6364e35a79f470a5003e3128ce865fdd073cbde
zfe7d23beba5b6435cc71c32caf0b92dd40104ff351b2abffb62d204e9a3cff614cf48b4c6f8399
zb958698552cca5d3b9b0c465e0cadfb26f1fb0703e2e1344bfedf843d23f56176884753f5124bf
z8852a0321f3e213aa153b47424e8c1ccbffd47a7567c17744301d012877cc6c2f9c012048c79fb
zc476c9ef5155fd50999603cc6932e118c9bdc357743be770d057530de9608ac4cac7c35167c979
zd674c76c7f798508cc27a9dcb0cd2bdfec2e31abea8f9e3d0e6831fa6c5438f5b0c827b5400c0e
zf75398a68e9998e04f88a0a071acd080950b64621c8f77b1c16b440b027a2f48b223c5fc84bfcb
z5e036c4c44b58f895e5ed2c40edbaf47efa9c63c779a3df95b179b13528d8753d831f0fa4d6db4
z1ca7911aae7c12af31f7bbd334ae59c49a6b39b4e98ebe9039585028fc2abc9925f8c42a359831
z1f555ea735feeb5f88d019ee737629c16211ca339c3d24453e494233b1a41e105a07bff7764209
z91160369c6071f88ff7d241c08fd3a80c356168064c6ad672c118fc41f295aa8f6c4711f5e9252
zda4fbf8517f5ddf585c718324bbb386759606d29241bbd0d4f427399e1aee0826bcf5f9afbc4e2
zfd099d35c063654b8733ccad5f455ba883382a56f7e8a150707839aebc744189dac3def86230a5
zc3f2a49cf3efcb7c1b28cf0880c3807ba1eb8ca6e90b8301fe064d7570dcf26ce8f42fc3a47260
zee0f88fe734fab89f75b7bce4c809ade10a2118d1e133a48d3ff9b906bad012b1ffbbb1da357a0
z40d467b33ddd1df599367ff2530d2f520ffc5a5899e457010b1f5d0d21b5c295491e488c636b7a
z8685e7f1d8197760a884068a3f8eb052fbc79d6a929c3a929969a99667245a31c57ea5685e6b70
zfbda038a769b4cf71f2b1f139a4c8d368ca103d01b2794285c55d4be147dde2024a5ce45455893
zd6906c4935f8783d26e0dec786eb078d6eeab5d925c300fd56ac76563850a297813034e8776eb9
z9fdc4da4b66721099e644f7a82d756162bd52e9c3e4cc7b67ad7b26c9ccf34c40a53b19e1d21b1
z8b7e6aa312c48d81dc4f25ceff85fddd5d6ed5388dbcfd71f0842fd3f7477da4a24bf62f40b7ca
z4698d9a52b31efa094d209beeb591578b2b94b56d8197b1498acd1514637e0eb9c6a5a94de2288
z1b172b95467d843a37515e4507634234bce37b21e1ef81713e649c0c5af461aed3c3b46ad0d080
zc4c3d8d250c3dc1055f09740c3fc108929487852ed46ee385131a87457e16a577a3ae703e5fb90
zfaf1b8267eecca4fcd12b6abe7c4f4f23370199148646a054e0ba6d54c75a97a0640812e74e077
zbd5887aad104f2bda9f5eda686d8acb140d27abe35f41f636e816059ac68ec60705dafca39e75e
z6b20518c53749e4fbaedc0a4c7f98d2a4afe50a4494ade1f7cfd8c7de5a342cebca06f93176482
z2d685002b1e4c346e2bcc08eb3508b788f51d2224913e571c3341f9119f598e9929d4af6e4e341
z46d5d7420ca1c047c4967231b8e79647c27f43a546d6268d11485e27c590eb6f93be44804cb108
z95086ace76e6d63806752af78ee0e3898aacdbdc88c026a7ac8054953245c2c0d8c533be5818f6
z484832fbbd3572fd934f5a9eb20424c214354f1863f2987898899ba39179674dd44b3f3df2dc0e
z16a9d9080a418394e96ab8dec1da364c8615ecc7fccfb9fd5a9c195f199994e4bff326721aaf8b
zf7a31a328fa2e34d77ca8bcc5c85f0e030474becafe607ce53fa28a0364de42eaffc60017944ea
z610dcac82c1531c58ed7bff49020459c596007f06323a178a466aadc879e115031ae3571c03020
z01ffaeef439ca6f15e09fb68029bacebc393955742f96271768608117a82bc852682b2737a5519
ze961ccf6e05faae53f4307c4c314f0d73f5f3884d64d00cebfe47acaef547f3529b0326116514c
z5b4f71f57dab08870a3ec34077ee094886605972139d5b2ad72c75f511e17615530d3abcb81557
zea7f3f4fa47e431b621439eace7cdb4a1b532561aee4dedb40cedda68d13aed2d45c6f5a2b4316
z26148a0f9238558fb6e76bf0d8a6d3c40bc79bf06193bc00a9fcd4d2b73e8efacd14535b5de8cc
z5dc0e625b3393945c6f6f281ba6af77d556da93cf325d8ea342b0e4594b573595917e00ac5953e
z8c7695e326ae3b4897c3c33c3c9452b3584ee590f14282275a3f1df5329cd99438f0e11fa516e3
z3ded83e9466adfeb4e82aed1cbbf086e1dda10137fc9e79da9490d66b8ac5bbe7c84f2a3ebac70
zc69d02d0ef406abc0dff187cdf64d48624088223368a48a7d21ed93831ac3a01fd87efcc323ce9
z12f90a0c7856d875ca366b064e2fe6f435bad941366684102865eb22219b3babfaf052cea3bf9c
z9716ae517f62e3b57228f9a4f65a4a0abf8f7a5bb6496c0802fa928671781cdb007b5eba144779
z77587f5d972d428d810952be30b4b99fd150bb422002a350286010455be73f8949f0b37fbd9d63
z71e4892f2891c7e8876f55779a2373e1248e716e9c0182bb81d54afda50e84d4bfae7207ff6637
z3c3a38b3fdac30ceb1c5fd56e5e7eb2fd2aeb3aae35f25657190179eef4ca8f15be06d72027eac
z55f7d203d834cc7f43a18e7a8b50b9cf5485b009ecbefe08b17838d2f2719466ed50941ce478d0
z87f334008adbc1937513b72bd1fca9d7e5285c87596d90073c2bb2221481edf633a727d4d1e3c5
z947b49857475d1ceecce29d0af2ce0899cedfe65a7a340cff1f6c5439135d418386b357f803a76
z0d92c7f89452ec315c31b64adf9dea491e3071770547cde54a347d27511f2de15eda08ab224531
z049ff5abc22260f794f2d0164e68579eeeb766a227d8b2c55af984f41c927f2b4e4f0c211a2c31
z62e471516f0f61f98c8b4db51e53767fd31315ea4c21c2bf183f54e92a2c1b369ec8167c802d60
z71a1668c2bf66561a102cf73f30c8bb31db09fca4580501caf9d329e1cd540211b5f4b7b946197
z3995db6648b96ce84b1d1308931fdd91626a5cca4f3ade4af4667a76eef630344369abc25f728a
ze7b8720d5e73aced880efa90b90972a88ee134d8304e0bd9c1eb3659e11a7a49b98199e669feeb
z86e512f0b8dea536d131a5ee699326f33ddd1f113e9b2dc4abefa7d5c879b77ec85fe2ad444412
z5f4ed1c0001846e07620ba1c5253186f1e25e7b8a9a9838730a95b37c711d1bff62e8befbccd4a
z737b2e086bd0cd593dc462d8a1d75a596108c24a3bef345bf78120863f5ab3e4768c99f68b3f48
z486f826214d02edbcfb7b653a937a6627341a37a109ced563344ac87b7b4d8319e93d740d54ff3
z0b79483c8ffa3e4cef71c747923225a417e04fa908899b5b0f504ded4357e3eab009b9a74381db
zd079d518bfb4de84b975cb74ac326b34e79f631ed6108788eb13c2b4d696c0aacddb6ec0354a00
z2bc489b877e42ee79ec8a3ca85786bbb90b932a6012ae5e6c0da3ab59a95d38f70b467ba849244
zbd689f71428037404ac72db9c2980aa3f0a3582a10bfeba613d4486c7fe1afe2722418f5727326
ze74fd5931108805170affc14a20f6e7455a65d733ce9bfe4eb97f39ec27335d151abdc8a1db46f
z6f54db31f5db5a243ebce4f90ec8d7c07d4a378be27a294b0080f9c9e4edab374616239360c64c
z6a501557c49c2b36c8f16dfb126f6a9dfcb20365edd33001f48478b93a726795673dc493914d29
zb9cc12eacefb7076a407db8246bcbd2cd84298766117480bc60262d327c0c83f214daefaa7ec48
zff26a773bd1a6c2a41dc7baf43696708bf1cc0cb25af0096a17e3196e61fb6e4d7d7cb80b9bc9b
z5bd2e09653b71553cf9d19c8ca23101e7ce5ef13f26d748971ae2aabbe209ce130d0909a35a42f
z931913b2d9d2f1f260b4c08f14e202a9fa35e0899c6f26cdac8c5171ad8313454441dd5038029b
zc364e30bc2dec7e38f3007cf9f60dbc76c2b50932d1b450357587ba9a558c9b8a252b5b1d5a632
z76d3916b4714b42d0bd21e3824b68d43e71fe3f3e7f091db706d17469c386fc2109f127bfe4b69
z81102a7bc1dd608b6549ee48cb3789baa2ac01ac9a8c0697df70e36a5eb1de8bb5923e0e37c3e7
z7a75afb84a0b98f434123ae5e3d512302e9219570b6843539e4af722223c1789e93a8a3675aebc
z650f7675f414c1ccfb59dcb106aa481eb866afbd713a8747462fd12a26da52d3cab3ff1465cd32
z9a018057310cd3a73c665dc4478126ba65faeb9d4eae9270e00cbeeaa470798a362e5d35ce75b4
z5d8ec8781fd326523f14e906f09e463e596c69117ff7c902830f2c73b045b0a1a9e78b5f11a071
z52b1f6c6b76f4a5f9177f231ef2ad1934fe7e7f134595ab1548a44fc48179a7e469e3470f9ec9d
zec2c6b68d5c2fe8b2f4608e081a282cd4781a213f3ff8ddf5915691315918de909828ed9ec104d
zab68958d3c855ebb606bdecbfd41a85d068c70f8e25e5ead8626e98703dde176513e9cbe4fe3ff
z50d0c6f895c7ef5a5a4f18c79576cdf857ebde6edff68885d6376c6a0697601b9f6e28cef025dd
z3a27ed314b0b4c8fb460fecc029d4db66b3c6ebd890f4c1b652a47a86fdb15e9fa63c9940e7e05
z9b58f9954c0df8587d00f796ac78807372fc7d5f05bd4909226be2a0e8f5653cc6ae499e4f1535
z192a2ed22b4cf92b5e4c0e49a3bdd84b75c565d994ce4902cbf26382c9166986be5352d8fdb633
zd2744f285c098ffe59df7f891900295149cdeb2b373e71db901c0dd15fffa26105962ee98d26be
z3b37982db64aceb52ef997157ca59143f6aca828f50f0721edba2112ca89468dfa93558822ea32
zd22bdd38c2f949f51fca027d417bb315cceb2dd08aae97100b7e549b0c973153bc13617cddc478
z5cebec4aef7ac2cb54f263c95a8512afb0f54626afdc7df3cdbe9dcf1146b7d8d0e96543a363a8
z115a24fde56ea4228d43b08bfae8e44e975018508789f4ff53e558aac63d6e660cb5cd42f8fbcf
z43c506e31ba30f86819f124897a6bcbc5430342b60e7a04ba72193d4485cd4781e01553958d80f
zc0507d759d225b69ede1ac9ea05f0b9ed4bf79a067523d025a41ac0d17233a41f69ed29367b72a
ze4bf9f9b34297f31eed9272c917a4b03a7f34038ac3541f7cd8efab45bfd3d8b11649c2c07b425
z645a31758adeec5658f5c22170529c247f4a4c79ba0f00bca8ddb7c96885f2f04d6eee110a2baa
z6f54c3b46cc49a96e137e16c535778ae4e45e4592605ec0e0280004cec883e7a418cdae4635581
z2ed57f8c06cba4ffb129230af015052f44c267e96277005e269a1e1e7b9f03e986cf655c2a8f15
z9da139ea3beae2ace38994b2493f711b8f278346d6bd491b9c17342830000c17f83a0476e19c96
zcced70d8be78028a86813953a70dd5465f9c7de699d842120c219deeab7999e2a832ebb3f76422
z971a035c7e99549aab1f80522a3159d2f9297f8064450e9f610af714c2cca0b98fec08a6020503
zd53cbb1bd77df76f6acc6bf4c16a8a55102f3bbeedeae448fb63f395476eadfc49db3861aa7d52
z24393a1525b56e8d1ccd120baf74f9c67b040654b78147f7e4adde9f55db230913f122310740c0
za5e5c06ca9dfb44ab80dce28c8d6d8df5ba7696d5529661cdee194c7d0c8b3aecbbc1c7cb492de
za4a0e44c6e598ae02d3f9e1fd84fe391622a4fd6eb01588875e7dc2c7b00cda497e2624f6478b8
zddfe4221be108b79d93db02a9df4f4d6e975b5d7473245a0871b3408d80dc1cc1efefd589fa144
zbd1f0e4d40032f8ed148fd9937882688af3c958626a31d472fbe4e6cc2505460448363e80563a4
z59b5234571c17c9826ec0462d4007394df934ca713bc81c15fd8e953f608e7e2c23391c3ef91e4
z461bbf24fa1482000e472896d5f0b3ec7e261c5d6bea036056864ff8ace53b9578b6862066c2ef
zd4172de3e3ec7b3a30f74d8b1b02f418bf3efe46651c5bb1c3add8047455ce4b880008ab7ebabf
z02961d71b8d554500e527315bad63d2c2441aacec1cbbbd01972ec7eb681d3966332df8042effa
z12382b817f3ff861b8861e62dfc4488813675f4595c6a58d563cdffcd0ba4929475a895733d6db
z7527df039d8eb2733d7878a469781e13c7f428d313348adb6ad8412535a76de03a4738367d250f
zb697390de994ed09e3f0472f1952a803acb18302615fa4fbbf704dbe67185f37361c1cdb4871b5
z7e842add65acbc18693583387f918492777a86f07358fca1f50e5157046d084bf4f783788df9b8
z78840efae2f0499c474f2150e29971fb6975ff1684f3b06098355953f837b7a95a894c0a5cbb31
z22b6f0d6fef6bcfa833d624f1fae0c62850433f1c92d7891484a91f4d5f85611bbb54bf19c5997
z15e4c9d047d2ed2f172279ade9949496047d99bfd47a33a0df4f7f6a6395315dfcfd17131ac8a8
z2e407493b6d3df68a593d3088589814f0a081cd914266939bce20f815a299f6abf6d4c0db1e36a
z0f145dd223d8eb529172f177ef787523db119ae4a1f12dc8c0948c6db13c8cce20b57fc009d640
zf696c2f58e470ef4469ef610cbb52242065e7fb0f75c9dc6a350c92cbf7d1b16ecbdd3f4f49e60
zf53a3e79276691394e3086c27ec9c05cec8d0f83419a7655c384476252bdff9551c263e0c9eaba
zcf1732689fa8c65b416d46bffd78f4467080015f87737397fcd4fefefa2a59206522c663db11b4
zabc7c14dacaf2f6c1be8a8afe144e84defb5a449cafd18aa83f779bad4fa4e13fedf38dce5c2fd
z5edcdc477dedb11cc52cfd3ef854af16590f8cb222c8da7c2b6b6c6cca3d52aa03937a85761fec
zff3b1f3602c37bb2b15ecc77a12bedbc77290f23eff45e0e670db507958bfac8bfe36c6994a04f
z68687389fd32580510a02aebb76b0a9a059f4109101848f64ed976d1091ac25a2852eef0a80b40
z93b53cb76065ed9e0fa117131a85ca7061e8c4d7c54f642e53583a68bef59e47b811d20a47897d
z9c81c36f2b06c1c1ce331ad035c3a44b06a807de75e96babcaaf0df07a749472836e557cd1b8bf
z1fdbcacb4628a7ad4c7a0a92793b6be5daa653cd8d567ab90271970a832216e6975a79694d43bc
z1a49b805efcca306c206ba4567a07361fe999874f18ba4aae466689dc70f4d5bfe6f1f535b66e2
z7368dc56ab5e541e2ac29cf244b0bbad0052abed726b08c8b0c24f985067f3fe29806507dc8703
z61fa48d825efb6ae4f0661adcbf6a3181a788dc414a67ccb650a86c20f8eebbc56a24d2becd739
z95006933de3687d9c79bfabdca77846e7f9e88c9daf0648d1d842db16649e33224c552204bb5e3
ze9d013485c8f305701306a6a0f5135461a519b27ab76f19586d6c193cff870e9280f885a902c6a
ze8fcff535a00f1f32c624fb5878e5349399930a0b9e11234edcf968a068f37c08a505d94a84218
zf420174a2bd06c0476560cc6c4a4f22b02b7171333ff11e03fe6f975c3d105996b9dba25f14190
zc252e11a8f1f04684870befe866e5cdbf16541d7e107e1bc38722baa96076b04a8e43ceb65b6e4
zfcfb568a01e09a9eab129f7af57d48334f7a0dfb3beec0b16df8122329f0f4d7f93923a13928d4
ze6216de9531efbe2acf09e7aa86c7fb2174760ff3ac9f191d4812dd5600f59e62abd4026ef0cdd
zc2cc5ab47b4755b255b0e10b14481644ab8d5cf805e0a691d74c9e87bff005a9ecd74e8acc028b
z7fbece8eb1fd0e37da277de6039e0b3b218f23433772df3cde19fafbaa8ede6a962b6a2767397a
z982f5a637d033ecebb7a05f19d0151163aa68b2b1db2eed39cf15c6b727f32e246e38de38dc60a
z995d0132d11c9336090a1c296d531965537b19c9746e402f68d19da015caaef1921669bbf51ad3
z3d536ffb153bae00bf3bbf2ab847f6dd42b090feeb36bc465787c62ff1e96ad6866b8772bb87ed
zafe95c7c321bcef03e7dd4d0b99a9733d51791623910694b6faeada425a2faa732fb006f1a5aa0
z2d7f155adf88149cef288a7accf774ec7be9eeb1a686cadfe4f83a2f6b7ec7c9941051557e0671
z655d8ccdb874e6b8550707ae9f0fbba6ae06174206cc826199d21421118da66d4bb5ec848ed308
z4796ef93d33151b1300309052f0eece50bb15cfc0bb90b299ff65fa4600c68ba9e2f11ecf1fba1
zbdf475d13d604a5f6a97e761aa0577566d4d81dcead5fbd1d0a00e2472474d16b62da893777830
z33b7dff0b1b4d05e342f6e47eef298daacc8c0c019e2f0c265cbf79f896712c69838969ceb4b96
z57add2221c26bfe605fe7d6981ed295e6fb61947f7ef7b397cc8e8eeffd7d5da527188e6c2309a
z531ef0c32ce080246e257b85a18dc6369da118dfd9edb3b037e4407ea52f9412972152e64d5454
z7dbcc859c1964be3d46a056b4e34179cb7b1491added12fa9ca8d0ba450d1a4090c4e5129288dd
zc737807058762debc27b83003c14932d199c1b7fc24e0b76f765f1ca8d2c18482c14400441b878
z7a571b0f77bbfa5e35d4dd0a52229e46d8063dd808cebe6e4c10f13b6ce6bceb35d528d556354c
z6eabeafd264342d346bf2ebe3dae8d0723e8296b5e264ef85ff108456c0a9ead3c231a2ef8c26d
zaf576fa608554cfac6b52bbefc872422fb6959fec52119f3f8dc5cc2d1738565fe74881639f166
zd32f0e499c08211b563e075d2abd6e617708092a3d6d6d81f65f1a4d29a71df9f2ae54a9aa339b
z1cee3cd10123493a32cc69ac36de1042d05f3402e3d8fa3879ca38a9d8c693d48d8dcb2d506079
zeba449dc9a3c381fbf05ae7c3aec393b43afa77bffed0a500dc108abf9c869e72d8d2b34065fbc
z24bb0e82f8e320ed780a3e8722a5d5368becd666eae378a645d2f6ab3376a23d287689cd52d74b
z39d056b10711315bd5d1bc05fad2437caf1e47ae66739a1e8bf8d1646f15d33b6071962787831d
zed07cb3dce13b8922cb58b914b0559fd64f2637016f34d9fc8b2de6cdef26bdf98e35a616cdf39
za631acf6a1ba72c7e8c9b1b757bacec746ff83aea8f9830181d79a338ca7a504e6b432c1c0fd0b
zb9128cca841376b85bf842b3ca918fedd38d7a7aa65bb2b6dbf64e85e4d32fd32c11e1991a3c25
z9b3a60bad6613d229df8086293ffd97f888c72e0abdcfd28ae8c55f2be7c7b836041bd934c9ce2
zea8a72752631b5e17a424a3ae27d181c13a3d776c8e18ffdf10b48307ec04d19e47cd566e7d7e2
zb3f5511deee4bde35e06f1d9e773a547a7291a26d0664818200c304e856d25c68ff8990d04201b
z001992873b4d14b28d006f91386495512fb4ca9394968fa49231e71ed5eb8d521585a070454d21
z8ce980847d0ba97aca6f997aedcb88109c6bab031342ce6f5f9d183f2daf3dbbf0feb479d37d13
zf659b0297430a18042a743a38976ee26c317b133858da751269f6d03db022b4f5830568379b70c
z0617be8a8cd208d0e8f8ed58b14a92685888f2d930d22e29b26f9d826e13b1fa48bcc08215143b
z998957862de6b380c68d1e61c930e8df0c2b2a8287e8558df57ba8522bf763f3c7116c4c7e3ff1
z9d5f2f774acdc1525f72b3899b414d48786331e58305e5b970544442f8bef40dce83f8fddf960b
zc82ac3be8434b0878192c48a7325633b950f6ca814edcfa2c7eb4eb0ef910289128c713f91d090
z70e472d38f84006e5a0599827d3798681c9edb38968508a514fc44d2b431f5872aef49d4ffe85c
zc0c7d1335077540cd1448518d3a57bb95c8b5dd6eb06fefcc55b568df0dcbc38b4e6b735ecba2e
z4b82422ac559ce6562e142d5870f6262d7db5ce08b578f35178f86061effdce3aa94daa2bbc255
zdf6d4d5788dfd1684d40d9524fdfe90b0ee612e77a3b01e6376f16815f01872798dc8ed922800d
zae1da3beea3638a2ed5d700082237c5ad87692076d885aaaa47a567af6c8b50ea0f7d3a44cdbfa
zcc8e3f22ca34cda7564c66f2975a6502b1524763db0d9839fe748d81cf5eb3379f56d4e86cea09
z5eea8e77a30c752aee22365498c0efa288fdc1d39495517e308ce283cb32a36986b57d599f054e
z4fd64d03e04886b4e7006708cee96b42536ff60e86dcdc6cf213b15b0c648d43c61b72c614bc8f
z0192a90a1784864a7bd2ff5397cb15219eb2c3d999902b987fc5c5810d66561892f67032b90096
z9451d31ec48c170444198ef1d6d340eecd7046586d05922ee04ebfffadbca94a721ef86ca580a5
z5976ed5a4ac0ce5fd33690a424f7d1f576b35a3cc296d35eab83299161d3ce31d032fd75d6ce7c
z75d47b83d8c13f50cae32caacb1ccc3df0c6b9f5f8738e8bc3eb3d5dda4ea914e3b370674a9ad1
z0f728750dad91bce0ed54e8033a70162680414876fbf10ee9850127f2d59f9189093d6b4009492
z2cfc4cd03f3a77f3faa99bdc486904fb2a1d41516a564a73bc43825bde5d9daa21389671e7240e
z355c96a4859602cfe99cd71902e313905df84d7cd3bb9126fadc6bf272f07486c6a0e075237b47
ze63b9c675172362764f517791aceea7d39d1cfdb55d0bb57a77391557be0ddc36382d54eb72879
z7807ea2b549323cf7b2a8a4e51b3ebfaf24445dda27d039135c607a258a5b22524accfce856489
za73c33cbff7cb4090bd84189c3fad80f097742f8b30061d415be59d696e674d51b2306741ea6cd
z29d300dc4dcf0c66c0a814ecc9602c4b63e03a92e7cfd7f99b810a7039d38809ff827ebf933c75
z436325a6b0512809c6fe71a2bc48d4e3217bfd33aa75d4fffe53ad6479f7471a7cd27412c0d262
zf3fb7e6af3ce95aed0407f38aeebcdeeea2278f448a27d10595275d726f99a23fc10cd606c6625
zd730180b0088f6c38320b14fde12ab35e23898f94aada59c47b9af94fc35340ca7b7c0e63d249b
z81e7936496d59c3b3f6a36262570b54343a68712feaf9a1ddbf857ba1500c19c0d7c85286fa6ab
z451b0ec232ab4a5afbf47c51a9efe2f6b1d17fd177f0905dced9e273a22794c5c0fb3972c20d63
z001c60d9467dd539c311527d5b9ce5e0e1d03a550f4c725777b0db1eb62f61f4bb103819f92f91
ze6ef6fdcba44f0d61b660d57320fae10b8ebaeb29bcc8faf3982867b665fc51dd5ae90d10c83bd
zcd4f43321da5e0dd060469440c00c5b889751d520194f61eff3fbc45abb95c6dd5859dab817291
zbde98f27343b47fa256b93b08dd347904493f653badc1104ac801acd24142a825eb47395da02c8
zbc3cb0bb962a2ca7c88c8cdaacf5287e41f3eba97e7738add4f0488a13eedf62f78f168892d227
z3e4ca897152b4580e5e4303d30f74148f37a6644213875a4755758e22bc0c706cca2c68b140391
zb010973ad7a65a084b041d28b82d34e67e665b0b3c56903549be6f5f5f8fcda58634edab9f5829
z90a1368c1d8cfdf22f410794bd6ebed30e63a92f6025e1878d6cc0527edc6b464bae2eed08c076
z27ec717e8bd6522de1fa8529fde9ce0d26acebae009df28d51a87481121ebd31ce87ccba5e3950
zdc5961a3cab1aa024d4b6c5cd53c518ceafc28fc9c02adb9dc3e9e7f45a096cc625e20ece76f23
z210dcf89d49d7a843dfa19440ae23f664bf8cadeba463ce74e8425b7fdf7bfd21f5738f41c2199
z0c73abdc713e0a1899a09a4bb97d596c3efdaea491b4edfb60dcef96445616a3b60d9296b9fd4b
z0fedd99bc1bfc8f4d640f3f7b3c92e3685bce30eda618d88a6e4ba08d4fcca9dbc8dbf1ef8ef80
z0c0c4b1c8797a9c61153f2ffc9645f002613c7187def159088b004152f6d22fb12c610dbd77f51
z002f8457c75e8170681bc755878b20c070079a38dc7033ff3a5c01dba43be05cba9cec3438b938
z9cbc4fce3ab132a63a14c12d75fa6c682e64fffd9c754896e83c124d485a905104224f9b615dbe
z1fff05a8632eb049131711a24ee26bd8e300872ea87e061e4d3b09e721109cea7a83aa833395f5
z19dddf129d1a2fafaf816207158e7eb849b7a73e4dcdc5af5fe9411e788ca8f53f66ce89c07a9a
z78ce672b025fcb785595891b8487609394c101d7c13cc1a5164c459e9630c7af13e509f7c77d77
za882392c8ded3aa18eaf0869513abddbb63860602fa05726f31059574610946666837a335a4018
zf24c9e42e422da81777ccf6c4dc440a85c5f48570aaccc656e02b50ce50baaa5e6b0e63e94d2b8
za06ca563d1b5f991efae1a2b040eefad54b3ac9dadd9f383acba9d629ac7641f80ae8657e01a4f
z7f7dadcc77cd2cb332395a4020957308ae407c8c78f6b40d1887e97b51d2cf512a414fe07ba6bc
z55808332d77ab296eff64c40c1b5a1ccb417898aa3087ab9315229c3dea24cc7209bc55dbb142f
z89942896e3064e54f0ff6f869f7b85165128f1cd8ea7fdbb105f221466153161ccf59c3db7c48c
z9e78e41c6c2cc3a0a2cf30ca76dfb08e54ee2fac9b0631bc0544f4f4ee2284364f1fa8d269017f
z87c95c01cb0b11465b9a4e21d9dedd20cc7b55ff2aa50ca0775f5da2364b0aed8ff60b669a70e3
zc1c9638a57b336290729a65d06928738d9b8bb86733a105d4729b82c0e48bf62877eae3e450ca2
ze2bbac2680e1ce6a00683827de8ebd0af31ccab5c6b270b7a5f5138db0aea40eb6c28172c9afbc
z64ce3c030124b351e35a89ee2156adf2aa39109587fb5ebb54e428dd2f59f437aa2e3c03fd3b0d
zc49549b5fd4ee3884316fed006a5fa45bd31b9989802a62fb574cd408643aa947270e5284adc94
zab497fcc2065eaca82a7b11a81cdfaceab6bb9f44507b37e446d9ba9043d5c0de666340ee8ba98
zf4f8ddb87c313493d38d2ae055ae1ced33f2544f09efa63c3a1d0535c788f1d4e594dd21e0fd05
zf47852a3f5f4c66befb27bcba5dc1acd9204351ecded3014f84d84b6df7de8f7cbc2dff9924399
z37230aaaf62af962c65618bc06b463b237b55c6a9330b14d29bc391d35e6d238e528baffb06a89
z627aafe14bfea09690b412e58da91b67b3c5ba417268c455207279669cf8778c99d7a10ca380ac
z90e93bb176e68ca259f2c7c48d2d2f69292761e886ab9f76902674a583e71752f3fd82151dbeff
zedbc3b12df51cd1d88ce196b5105f7f3ed9f042a47d7fc77e578f0499ae22cef952b5be1ae3f89
z29a13dcaa71570a71bbf163d3c52e14c2021fb7239034b3823f0b3f274b347249a832d505b4d61
zdafa7439b458218aed1e7c3cadfd0e8f5cbeb386aa7195843cbe4f89913b0d116fba310f319334
z9a7cc5c2dd03d4d441acf212c557a26dbf5d61b4249e228ca8f27c119c2985d0fcb06abe091e0b
z6ccdf8a03daa6a96573503e323ea11931b134f9ccaf91be7e97fac3ad3dc24317f71a49cd6e080
zfc0b1785ce3277ceb20e92689236c2dad1aca5f4941affd33bf738f06ec1dc9bcd0bb3ef4ba938
z5202a50a5974e7295afd2f5d34b71f5322a35a5dbc936fc0fed45e83688a81b8bb33186e63ddd4
za360cb1829aeabcc7efcb247dd3f07a761727c3b70f434a569cedd6a6d681a66405fb69ab77d1a
z06d28caf3fb089a3d44b055a2720c0a9a86c0551b96a94baf07e56a41daf8cfe2f0e66d9195776
z36424fc3b09ef432046c32dcf80137627cbbddadc707317045a9fab9c369b43aece4d7b8b7e5b8
z88eb3f9009727b5d3aef2c7835ab2fb7ad58d931b3886e02a70ca0f111698f2324880ac842ee2e
zb2c114cf5be0151ca5c849c330806b1c3df8be64dd069f27e11338cc75f79d52cea919c2500610
z6c98309ee13ce7f4cad5c5e1256751c422612d394a1a961250db121ad19687a435f8e4d8ab5a38
za5ff30932e774be12eaaa4a10c110299f7eb3568bae7e5dfc49d0f9378c57f39d9a6ed9bee839f
zc2bc4b3da50c663812ab74d1594d73dd17703eaccd9a8a312e028413ccf079949e4f8e677551db
z36408b4db166a73b7349ea22a7cb8c9fe7832ed164884038fc357aee29736b8b92a14318f400f0
z92c582244bc49b322944d0583b89fbe474c2268373149e3dcecd5fbd8a5da9c2326cd91d831583
z51ca280d045db3c55d447ea593be49800f9931674b919e86336aa6d78f44fee248ac07d8b28f90
z3e3945699fc7d51a519aef551b5c009f5ed9b3caafa3aee001c6d038f06fd84e1403031a3aa564
z618d23fc2edc4d3869958d73e1df708536fcbc876f00e2c7de4c26b410db09124b665f8aeb2d74
z37f9d32460df1a7ceae5f76469c4919dc95f2085fc3e2aa131f0d9514dd7942bc59bed1f3e67f7
zcdd93aa3e524c8e318a2640b10179f6ab6b50fea02ea25a0697b9a1865f143d51e54d1af551e98
z07c21da13bba5284e106fb8be530068b878eb9be7f5acbb876d1575c9cb4409e7d9dca33996d93
z140fbea8f52021ed2b1b1fa4e535e86274bd0a28c6ce39322baa89d5e143ccddd87768c6c04218
zaa38500e6b8475cfb2d5e47f9b4f785ac6ac8b7d6ed275a9fee48d40fed7e1db64e1a5e6c84360
z01be57074e1f7a2bcfc4acd32482d6e8b0bc0700750e3e04614c76dc14dd0de2dd2899cdbef117
z2c8dd65f9fb6728bff22d9c1b9c348db6635095aa59f9c2ba4c472d0ed73ceff93b8a0327b4a25
z0ecb0f04cd994ed39f4305decd3c37e8164200748da5cb8111e1065d3364df44a1c8e3084f4778
z86eb25d80bdd78601c20184c5027898520635a1e2463f48c79a495596f32b703aa115936f37c6a
zcbc90430acf7f2e1b28cb5bfa9cbff4e502b2757a78b87ab18d782a0ee431e922b9a423ac1dfa8
zbeb5fa9847a11ba3577b6f0e2ca89ac0b01c9d5d3419aa37a69b1ef32a094b8caa9baa1822faf6
z9cb6fd75becb3bcac5f32e9de590ebef6fda175948fa121771fd887b3bf3a766def691778c554e
zf85e65748bb9ea7f9f63d1184d1793ec15656d93a8dc5fa35b5ac2f1b40286cce9561281371c1b
z02f53d95a237d02c5ddb1a9439e78b4ce3b9b453f110c51222ad2723363182d13407c4024395c3
z8fa8578af84374bbd4c4884a423cd2faa4fa77201ada8059d0d5eb8173bef3ac5f849c87da625d
z8ee62bd7b902332e645681061fcee600e5695e43c24f24d2496d298b7ba9c46a96639ba2ffcc19
zd1a0b2bf09e96681fcafd5b72574f6433a8aa706582b19e6d69736153ef0b935e0cf9740e330b6
zf7a6dd85a467ec66e1a2a07341f8ebf5b4b67ea0e524119e0180b8cd9b088a8fe3b24c450ea55b
zb5899284d924c72762e32a3890a89bbf9b96f889430ee92dda1fb3615dc011661833fd9c1053d4
z98872948b1730d014010c119847d8f9764c25c2be13b824eec99a719cb72063f5ecf874d0febde
z8a2fa1957fcee87f82b1350af5d333592a135641e2ab8b9b97b80d1bdfaecc52d470399eae7ed8
zcb3f310784a2cc5ba0a4334304efbec89873ccef16024e0131cafc7aac24824d781544f6207f13
z533ff35f61c2c1904e6077c87764496d125af3bedd55902e5e7adc7c2b35a638f68be3bffff585
zdf07b6e812432349a4f83de4b889a6d7d3657b71499f7da252282e3d762eb57ed28e7e16c57f71
zf7ccefde117e5fe61591206d4ca64aa9722c7f29d65736eb967ece6c302bd9312bfe82df4897f2
z4ef8412e5aea2aeacaba4d8cf5740240d57e738d747e7408822ea8524bd8cdfb3c935891965f3e
z2eeb5b7961186229658aec478837e660186218d9182eb4c2d4e9b415ef8a06652393afc8f79756
z07cce5f853e497c96a63a5987f770ba0f3fcb5fe68f7c26d4315c2d69404f4a56ce708ec408d23
z9ea4d21dada0b8af1576301fcc43fe6e1381547bee9cfb7525f2ef204d158843d5c01c558ffbc8
zc5bbf3a0380de2281e0d9dd5caa215d1e5ee1c17e784e2dc73344fc2fa6d63fecb316fdf0eb01a
z7e139a9a630c2d918d8d2e8d176fd38c7d7302b2cc68357c8625ad464fe64162f4edf86e66365a
zb32a2668d945a650d6054721fdecea58b86e8204a3e78809e27fcd872d49eb07a5addce85323dc
zfbaff4c78ae1fb23ce1be5f5b54acfa72f3bfecf527892bf565b920d2bf5a62a5718039a59ce08
zbd64e007bd086b590a48876bf87f1cd1274af6d05ed0f28c472125d71d19eac5a1cb1d4dde8e47
z28c9873aaa99346627ee1582d2007591171dfbbd7a93a41d1f5704e89a7a0f9983cfe76d8323ef
z059de0bc857464fe1dc16d54f91b313b1f42b72ea559baee71caf93efd0a22693833c2606cb254
za2f23a15c24fa87d5e1b37f55b9cfd91b70ee12a1146b5885d409bedebce04341034b69ff4cf90
z6089161bf9bd098a6248dbc30704b772aef74c3cdca8c0d5bb251f4ec9dc1519d857192aace43a
z5cace51c8e4c9e0cd45a587a46d2248c3eda0ca4e606aa58ce40b33bcc8d85eba58524dafa89de
zb21db497eaf1b96ce0b936afd06093f8a7d4899e88b2d2af790c892bb373cc26e2a108e168b25a
zef5711da3dc39117c665f5b296bf5a96694b7449e530232378401c5a2b9199cff54666dc68b255
z28b52c6ad8e2d76bbf246de31cc4f5428a1e31a76f86afca4779e81c3be2fe3bf7b94d6cdb352c
z6ad567e12a4d9d6cb691c2317a6bbc99d511c4da92691dde2dfa81ec6a94081368c14d757fa3d3
zea8984de63006346176ce23eb466c827e7974daf8778f2d380df465c9e7539d62bfdfeb606c5f0
z41bec91c6e7fdefe7e63f8763d0a8611b0188de9eb9fac0700772d79b4a10574dbab708332cabb
z6720cc600f54b15706783e52d62822603c4a0545b04d5128dba0c7434abc8c2dd6f5a64b1eee0e
zdc0e0d4a0ea0ebc202f504f2e18ffd5b23a04273310a59db592269348541b4b540b245410f4bb8
zc32deeaa2d553ac2f433369044304c51778a17fd0c7367adfe402043b5886ae4e8d89dba6b8227
zd880a5772a416dbfefdd8e96f140e23bc5a4367ccaf6d076628c201b805aa2e98026b746e0748b
zc652189c957411047fedf3831f19ef2f6577a88a94f1e84cbf1c5d7b10258b754193d2f90c5812
zc54287c4dabba0586286a7af86568fa6859e75b82892c956644458771f0956e3cb361f6c1889d6
z9734a3d30a14cac59d3fa47846494d630ce51fa8ce629cf3667ae2d9c2e77646136dc60ce896a1
zd9cb2db02fc3e6271f7e83945b9fdcd0f3659c2f755cc4cd7dd9a543c8995693a07d84a8901b1e
zc5057975883aeab27ba37cc325fc6fe66850da9b6878d2e5569d414b54a6afa950df8b2ad8cc74
z8170facc5b3f93bbd0d4e0e2c2ded32d05a727d28a65a02d1b032800dbb1895b6e184bc01ed2ae
z3583ab760312510ea24b9bf55240b5af6421cd8cd4c4af037d1618a826cfe9d1bafe5c3b6df98e
zeb686d017dfc83bba84ebc66cfedf882fb77655b65fb2a9b0d513dc4e385bec7fa87193c799bfe
z245939937c4464e820762b90d79553c58fedc3c31029821b5a38183f4be9fbf3a3b40538ae9009
z9b451f033acf09e463eb136e98a9733abfea406b34c855f2217f35633872728ab227082f173a59
z32f481d9e0215a081a1393d41837c789d771c6e4c5b08192291fc3d9ae00038490ea3c34d93564
z6717d16bf13c9efbaceb952c540858d4e65c7c3e721c9347785aebe03483eb345937b0e8a95dc7
zfd5a0401856ea3a2a2889c1638037e497e78c8d8d8dc69723f47c41e681a064a74b8b765a2d36f
z1e49726efaf4dbb6920665a5316d148111e27295f77d0439c90f72ead817f0ed8dc7602ef4c5e3
zebc0b15d94905822b782ddfa7d6d816608bf6c0f15f19529773d2db639eaeb373e5a682216cb9e
ze49b408739a29accc582a713b0bb4b1697467fc0abd56562a91bdddb1973f409bfe7def3c6ebd0
zf19720e4b63faeb49d645ea24ceb5ff6dd0564d27bd1df48be8e6a46a4c01d3c617a3f4f4ee9fc
zce0dea5d897a473af7567d22ea6f7132e77d2fb5a9c448817b57764a1552b2f68995515b225934
z2573f7a2a021b5f8749c033632110363dc588d1e230cb41d8bafed78a81a5e73bae8e7b7e04878
ze78520f9c651664a61cce45661108d54a52e6ddb89b2ed68c3bb1457e7a20041b2087a914f9dc6
z7c4b6700b748be95aaa2f86261ab5efb357bb8c2ee9bd9053320f5ddaf41327834178f1973394e
z200f94db5aa3d7553e68d89c001a2daff30202f15300a330b9e16cb2f873782044bb06c22b97be
z1390bb3ebf6617c101c6d9815e900850149aed9c5117f57eaf1f44a27d57142f18697aed4e9ba6
z00c2a0f41a5985bab8c787f107727ecaa852cb1623516e66e30960ced1fab345fd11d79ac9367f
z9315714e7a22bc3da40a07ef754f9365de1468e161bb828a004288f1a9c7bd97abbd1b1066cd9c
z0bde75fd4b76d5c134403c030b2a467b3f37d2a98e62c79ca6ebdc12c435837e808d6a3d1ad5f8
z4fe6faae81bf4994297050d03596e5a5667b5076e05c9900efd137593d1f15b26b2593e2b9e604
z8aa797cfe0d671753979a043ceae58bcb780292c820dd8138d4ad67dfda78a2ff927f3c265acfd
zd995476d14b285c65a48d352ee1f6cdf77e9fd85a24537523f3364c4eaac10619350c945afc6f9
z33eb7d49a93a5d0de28f42309f1aa3e1df3931345e568f441ebff354a8e3069044f5583a35a791
zbfc75c569881c8b1835cace2d09d5c07461ff4f322de03ecc2f2e3166ee17a84356a1a785568aa
zdc3db418080b2231a427d579cb9382760fad3f880ef8410dffd1bdec1fe8ac782469cd26a363f0
z392c80593f003bfa633dc5253261fb8f5b68e3c2723637916616e10a78a79710b38a15e391e2f9
z030114025a8e297e7113609df1496ce5841be7463ff813c378c21a732bfe18ddc950f5879d6ff2
zfc6efb7cbe0a8c5f13eec89a5fc8178efcac409c493f7a50893731821a2bc80d599061ba110548
z0625e1ef9cc4f64cbaf90dfe407913f515c8443b97fffa6770ca048dae2c2713bf1eb14b0487d0
za7968cdf318bdf7a26c4209595f880d3b855ec5a41c75f177500701cb5f0afc759bbfba94d6746
z219c278df8cccc32dd74f54ee26fb5c01ddeca662e582b06a86891e1587f1ca67fee4c622816d5
z2ea5f0a08d08aa5a11caecd3b4155d2aca291af796111af01a491e36db71548d01efd57a9881c0
z98dcff04521ed836f6148d1c632551713286c44a195f77d3394b4f0b87c51a118f818163cb33eb
za9f5a6a00bd34523a312bd7f4345a4ab3227b436ee4f1ed5ff6f1bc9cf59fe07e8fcb63bba540a
z2cd87dcfb3507ed4c7cf02113d6ce7d92776795f2d0064c7438207c8be7403f0d33ab42ef0b204
z4f3a57269905359bdda6206f5eb68301ebb4d89ae3d30de623498277e583bdeba52a3630e00164
z6c34e80c629b9612063ca2a3a125993ec9b55b32bc3158a6f96b316dda2e89f855ccb313395d67
zb63dcbda4401c006e66cac960f26eb217f2bc1271ac2a70f233f1f5b5bbf84f520144e2e6f9757
z63b9c52065b2e358d31184a81d3a105d5314dfaf56520458efabb565292d74ef0f683e2baae360
z6d89c5792a0c964c0d68b5707399e7598aa99c82b4d3bb38de86f7335d2d8d0d45d6b03fbadc00
zaa20c2fd0aa2891d3131a3e60b99ad493e98f2084f13164dc45d8de041ffed4f3d9e6e44b4915f
z7fafc66f5e199463695255285e4b319e32bdfb6888f20c21d39feea3ebd185da0ee6ff5c805a26
zb4bf263cc0e8b59cf64dccf42d54b07c9850da0e5626ab9daaa947cf2a59ac0b5c2350c19fc6ea
zdb06ee3fc2f34f9f4b32eeae1d02e5cb8e1e154375ec6811f88ec3828a05f7062ecb4652f50598
ze5d9d2315c42d665cee8aee73de432123c9080320ca8061ca2f70b46d77e7e16ded938f7ecffcd
zf112605337a85185279e42943b262a0061cfee515758fe423940dcef212b016905d2f09e097abe
za9b0557fc65105dfdabdf85a5674295074de846c6cf2633bfa7e9099991d147654e5cc55639921
z87095d8a061728d65472e101ac168361e1531d7589adab5b8a06c2a862509b2da10b9c5b95ccdb
zfe7cf185266d2d9a4e1958a5e0cd617ad9d5266256b1d8c3a6991b7b5ec06cd41d34c7279d1a8c
zea3356863f2fe17153b00214f5d26d043c8abb46e9bb2a7ca4cfe8d5573ddc12cf2bf0a6862802
zf2a00fbc15ee361ff9a283605265e111fac1b3c67e3eec57e5af48edda03ba4740506e4e69683c
z79117e9c8f875e5e4f7f8e22b675e5b54caf10a519d9c5470febca44e2ee9dd6254bd8c7475aef
zed36bf1e4310833a4901402e0c2fb95c77a85fb5d3e116f6480a8fcb0b43319a9fb4d73f2b954d
ze6479417fa09202cc5792c78b82f9d035c9a1ba97714404f4bcf424fa267ca16276675d6c64611
z623b05ed2964f7c9e2fa169a82c11e80e9324f2330d840da96e97a85c9dea6432e8b47b34a7101
z6c1021db5694d35d3412e9dc5a77a1e94d5fd2d09e69ca7cc10997882a2e04e9fa380955c8a4fc
z9c9c2f539ac3cec616b9fd5524838532ed3a7c1ddb7dd009162b1cc29ab4db7c928b82501b54d7
z1ab5e0e9b0d68d1df8c29fc014e91ab0ee0a00652ba944e23c765a5592e5e58267beb0c8883e7e
ze77fa4dad911d466b667b87e6a4291c044d18928e0ed493c09796cbc98ed1677c6c0662284588e
zb9fd5268c24669c07ac5a53dbc7a13969039cad56d9e27d053a91306de8a0da45c72f70e6e843f
za76b105e1248a25501b31e4ae05022c341ae850ba395fe6e45c967d98f57a708aa5b9f2c6b6a9f
z3fc7fc475c5b9e767da6e7d012f68e7716310329fddd2aa207c1ebbbcb8c49393da6c4a3de9ea3
z0647950e8c1e6a990879267969cb88ca531f48377d54721207ff9dca449e9410556a3a91364b6d
zbbc862db48c41a7c7c89b10fbc574f56ba687c507f3fbaacd934d9f248ccd34c0ddbf8dd059d0d
z7f138c02cc489525c0c9d9707daa854546d14bd925149b1d8ea048646c899043fbc7a517d0fddb
z6e16121c29a7756a8abe05c462e9a986938ae668c8d774e173dbe933c2a96ef6948ce065d26566
zdef9f6d3289a8d9a88b3e5491e8b16fa2c62af49eed6104148826ffa3d9d4a806e81aa4aa99114
z285e56e5e9b3d5378dc6d44221d6e20d382996bd5b87331f6d144b64e692339f0e4f5e26b83452
zc2f167894808427505c408b195ec2463deb995b7ebed933737b670d60ecceff89a4a670ac1eafe
z855a36c63f5b718deebe5ff3546d0e03637f0d7ed877f0382712a3e315e5b5b9a63d007c387683
za810eb9a7124ab505c8b2dda063e16a17b7a841a073d19016e3ae97438a6cbbc131e1b21e2d923
z06eb3dcf5bdf75e1bb211664da6c260bd1505caf0943ab2bf2b23553ea9e534c497cfaf2e4b3cb
z56d7ffb9586408fb9797c2624d508d24950903198f6641040d7790ca32487590b0353bc1b790a1
z849952b4505b85de270037dac5f5b6cdec59cdc7b41c861ae2a4f878138b566144581cc579a207
z8b6d7029ea661a0df85e4eb2ba7b71484e0ae999b2d5d87733246adecc7eea229da7d104c7f26d
zaee613f3abf7337e5f3dc8f192693c8834995656a72d824ce04a795493912bcf77b3ccdca68183
z3eeed108f795b03f69f8840f071b2a76b687628bff998148154149a3c068be53a6861aa091277b
z04ff16aa7befb9d6bac731925c90607486fc9e086456974e5936863fcbdc4b6b220891e4f7dd0b
z60f2f31ed7e26fcd7c23d0102608b42c0282f8027e4a10a9dfb997ca17d573b769290814960513
z03c8a09d75a2f18bd648d09f49efe42225356968c5e1b459dd58356077dd6890458b811a19f0fc
z820ef45e67ee1118236747f6aff9803a7561266f4c63c7f532224ba69e40aa28fa7df0c11f2738
z03de11a5480d020968782096bebcd484f129678bdd668d098816c39849a3a838b362b806200ac3
z5fcc34f16e3b7275f7a0ad74a4eeccd60c833ba899e6af8d786c6040bd8ede296060796b00482f
zeb3d566c50e6f2b0f190161687ba4887a9d3945bb07795ce11cd2c46973e00cbf7e7ab440515ed
z9898865c470ea7f949d70d9225e1538b221872021592cde30b602b67bfa8558a8c2baa3a41ee71
z51ffe866c2c053f38d1cacd4e76102ccacd71580aef3436b53c31518541fd22201257c459e5a49
z205720f5e57cd561bcd727894d00e62dfef1a92f7ba4ec8c91add18c6fd80372fb8f046cb49be6
zd6f0b0dd8307b63daff928836f11f7faa3bf57fd8a0a7ed6cbea40d7b4d97d54f8fab780defe61
z35f9b7dd288eea9ae45cd4b1b248c301cbe49e7dca2a2e746402510550bbeb668ea1d33d6560eb
zdb59320f402b5bb6b03c95dea7feae2ea1d2463d6ae774d4efd0b04721db452c274db45ce1e2c3
z1de9f643fb6acbdb5ab062961cde3926ef0d98d93effa806ac702659001216e90775fe03901ad8
zd155c15c0c1862ed665f219a1a672b62ab8c0ad82a3670ff29b8ba6289827c51ccc9a42ae8d494
zf32e19a9268756dd7e6051aeb1b8e255c414224918857afb7c1a88aef64a34d07558be17d3e318
z974bbceaaad3cf8db32520ff61bb368ad06f3dbd650919db655c917fb4760cfc96d13eaa5ae566
z874195578ffe22065a79b21a836a7132f4ca8457f4b487a893a5976d838b02194c71ec4505b8ec
z3efa2a9d72c5d19b90fcf39653c5e219a6933fa5d5a8ccfd2f6f2e90f23b1c3328e6071c3c262e
zf5c67bd8cae2b0e811329fc58b901bc62cbe85823dd88c5f9da9a8ab2822a06761aa01633bcc00
z445de52854ad88df415200e70df96f4d5fb16d416cc41cd978c6bfa20723918218c6ad92a9fedc
z1d0e5e273b67448d09657432403bf16c484c4de82c4364ed772c7fb33678c3782405adbb89b499
z8ee4653b0333688902f7b30030919bd8adb1b0c7b57123cc9dd9108e615aeb20919f958874ad81
z572f9614b9bd66950ac205782ca10b68a0babf9d0f3dd55c96cb3717ab6a778e33a2e69b0c889d
ze440bbbbe738078f8055324565dee90967fb86e016d0971946162f398513a2696de995eeb85e34
z7b28376989dfd3319096f8ba44598e8a93c8e09c52d369eebbec1723535b9bddb90f9e945ebc2d
z868fb51db4c4cfdaa7d3e2b9351a18632eb16d10a7c5e19649d214f1120793ecd7ec56913020a5
z1acf7463f28a673a43d746edc7c9486acf5e3d4348d0a2e99597b956e413b88ecb5c54cb1a53f3
zf90f5be21caa76c7c408e902f9259831da109b6e80db6bd93f47d29b994f86a1b96465a376cb6b
z4d282104b8c7b1c347f6fc1d528e92931bc1be6d635e40df4e4019bb343dcae1fb1acec79d3415
zf085f9b0e1253b33dbc872ac224674626804e3998063b08c21a7267eb13bbfb8aed9603c0b88f8
z8be47a301a53be1517fcc0dfbaec88312975a6c9499588c6e7ac1d5747c7b93763ea59bbdd610d
z2bbdd6c9069590a15b09fc570778f4c5ef3bf3927f476d788a76912d211c911e11ca1e8f279afa
z0d921cd5aada16e5a821563a31460c4a710824877cf628fb197556081efd4b7b8877ac03ee2fc7
zbc9b7a5e280f420b347a4c8a9fd68fd7fb9f6124d451220d463e61f13b13fefd98672dca4f1db0
zde0f29a85e899372b425aeb58be4b35d0bd244b18a4e979607663f24d2b46e49e9fb7b54e3f444
z27f32eda56fd7c340fb4b6bce5d88fd199554266ba90fca50564456bc98721895c5d9882ae725d
zd591b9e19a9686f7e6a56d06f08f67ce0e15d0fe56f0820b786f0c810ab9152076e252f9c6d3f3
zee6bbda9985e29f726fe8501ff80d79867181b3ab8f9523dcf68a3e3c7253015feba7da9542275
zd0b6fb7814ad33ee088f0d8ede6be5fef1171b685c251163934ab4c19a26d0d2732b0f9b1cb02e
z5a40c9e1418338b44fc4c222ddd530aa8579c1d80ada58ed521a4bef87c78cba7d293a8764cfa0
z319997699f11d031fefd2d1bbdac61f246d56816ab1a33462d767d194d8241f412bf37967a0d25
zbaa9799f7efd287e50292dd7c8e7c6ac9e1b4a65dd10e8ee5d091c40544e83ac8a92315acc1c5c
ze53f7f2bdaea6a19497727ffeeb06cd8512da930415ceb4ca618c09c01d56e551b2b72116cb3b7
z1826032dfd3c27723ad6c2a590520a331929d6ea903282126cc604a3313339c93552d9cb712dd8
z904fe312c73a8a71952add4debf88a8bf25d71803dace97c052308e6b627a3501ed1398c92f523
z5949fca1966c9ae9d003cecaf23006e592dc723e47421d58c552f7fbe0b21640bfb8ae7470bf1b
zc5048db6535ae5d1b6fc2a60654a437afe847aa465be82a32093bd0a3ec1fd67c39f5ffa1237eb
z3c078268f894b10cbc439c58048ab1541ab96f2eadcd7cd2006e2aac490220719b13d9b54749f2
z4c40d7262a4287b979bb7b840b90881e3a1fd85d192a21db75c3d8fd80499e190b1675f4ceb69e
z28fe0f0be786c571e0cfc022c7a49f11774599833755ac8df12baba14f1abdb0ad4f41054a56a5
z9a8e325e3534b80f58d116738103e794bba2daf8cca7bc77a381c0c27830a7dfe80a6777dd216f
zdda306e42adca8fe930c11a82b5ef4aca5a1df8561bc344029f463da1e1b76306ee9584213c376
z9d767bf42bdc4ac133f2e4f1dd060bd024e0213860432843cfb509880da72c1f3cee808cf42d2a
z33e003a91aa5f7efcadab260bc0f6ccc4004e82648e7f6b735f6b56a375cccc1cc0ef3e2a32f67
z6035a7a9645bba1bb045fe8bb756fa2d2d2451c102140af0eb4a1f5051957a78f066593435d862
z33288bc1f510c338d93e4b66aa19b6c668baf3fde654e1c3621d11bf08f4291bd5bbb2db2eac1e
zb2a8f04976b3b6f7bfe302a3c9db644723de9e37f4e324f648268eb6abee1f2ba5612e76fc17df
zdad8a651e6174481910fe499378ce3adba00a8bd8db2597153d92f0fdba6d0c63b97ebb21011e0
za830588eced27247c3acf17fd3b0f3f51f281cc957f905c999818891a3c9c521a0b34cbc85bad1
zb4d13f20c1008e3f7c45df206e0611313a37d05b05007dc6ba78408f88051ffb06bcc0d5b572f4
zdee69385a4b926b2867c52aa32658bbadef5e0978950e8d6e96cce479f0f82e796dbabd7bfd2e1
z07d3ee9b3f028166aa60246545835c087955535af6f4499a82b976b2b1f460b2e3809a7fd2f04f
zffd80b4d75e49d214365072bf0eb71d7765c9e1aa451d9f56be1cb3172283c333082c1dbf5092b
ze17a2b749c4630380379324843636a9b62fe8dd3ada8621995308d46ffd0b4dd6231b416e69026
zc1030b54f484bd0a22ed18314082119613d7be11f5fa97e8cf089df9ef875a7222f89848d34455
z8a39b83b2dcd403f6b31a10c55a05f66adb94e60ede8a59010f3e37fe16c9b8d6a0aafec25ef3a
z57359b2eaf3a9f8e60d7c57f1dbc7d974eaff0f212a24fe2a0e6a9b91b166f65533c379801a558
z7b3f82cbdba60f608352971d40fadfcee5d960e134bf994119e4f0f1850f146aac8952494f70ec
z2b9cc210e714e23b4385d64c9fa776ca08a48d1e41e0ea45f991073f2732577fb25983be26f1e2
z45d5a77d0247c81d9b054282b7e859677664ce3445426f9b0ad11c0916cfa5c04f15e522de9b63
z22f25020db1295f914649edf53291d09ed05209278ac63e895b70338690994a1f41db30faec3ac
zff23c4de08b533e129fc609e81c198512ef4dd4bac66ff3f7113916705b5525327e31a33a0f1d8
z80449173f19d93f9d6c1517caae0981a4e39fbbb6949bf6fecc9e48b281403fa75e847c1519117
z7e3f16efd2e95142f2c8e32c074514e6e6c75c61f32ed3e0c6d2fad2a958e12fea9116792024e0
zc0a9aa5f6df168f1722f729d26ef769e8d7003afb0f90573841f5fe53b56e454666c56353c0f69
z22aa07537c7492a6613ac5ca968c29cfeb61cb91be99922bd4a23c61fa1c44be233cab944a53f2
zfda722bddc5b262f69974325d71ba10d7e4d1dd3e73ec3aa2009ae9fbfcf65c71714f92510e9d4
ze8765708221dd61eb4f356110f1da3e2f47191d615d99c0d93a49990d162846a81c80261a0d16d
zc709262f9dd146fe70cd9cefcc0d5e21fdcecedcb8e080f1dcf07cc14bde8c5ccf1ee75caec038
z56cccd2cdd0317412c8caafe78802dc135bea6469d8b46245c5cc1e2028822cd063e7f7540a000
z656a56df231220cae79b8816a65e182fa6aea3ad54cfa52dc0eea05264898b30ceeb067b872b35
z803d0a2e25decbf6e2efd301aafc65e75eed5f1c0a43b1718c94436d5491971bf9f20ae18227ec
zf7ab5966b0de954e7474ac47c5283ca09bd7f3a0a1c9888b0fe0d93612b25b89690a78f9cd5f39
zdba19fd3be4a900de2d340bc651b215bf6bf059195587bbd6325fe261adf021d1ed441f852dd9c
zc83bbf2fe8983c03a8fdb450a10f742ee4726f70f52b393adba8b7baa537668b565f0edf318d5a
z917e251bcbd844ce8b57e29935e77612214bc023ac7def98f4aa444c6e03bd1abd11ff2b9a3bff
zd4c6e2bc61d576f4a99412554bfc6837140323d6f9553b8275126f3d6b85d3c0905497a6275592
z6ec7233af7da1f4eaa0248dc99b050116afa36738ac0768c12c6ac1f38a5ca74b869aaf6aa496b
z18463be8f8bde05c1ce05de3fb07256f9fe24842613ecf3c7df2c23877f47094187d5f8fc1fd2b
z052399016d5c4fffb0ce5184fb4875684b4bd1e0690b92b2d87d3ba6588bd36c114a77826d0485
z14515f0a0798a860c5cf441b5723fed408eb96569ff3264b76ab7d11e4f811ddd79d6d73bde10a
zf4cc82fe333b9057d523ff6df50595c743613d57da78690ce1eb13a9ca237634c14aea889c1554
z128e3bd9c2547fea5b5c521d7b5ec46cc10bde28d1fc0d0950c3c183e60b50c4831bb397a007df
z06763638b652dcac00c4e623527fe9a862ecf817eec70239926059c5a6ed8c7f1b5e1484b33cc1
zc4fcd1f8d4bd5ac207db4454661bb1aa24143d3bfde9e35ed089ffd1f04580a98c03d4011ab383
z2d50660cd4506057c446dd73bb853c0869373203b9df6cbe57168c56757f1a05cfbb441bc690d5
zfebe9cdcc9eb8d3c7beba53ddf598cd0aa9a0548f4f1fb4e73990b4b9e8b67429caaf1d7808330
zc693801cd5c8dd738e7db02ae09e5d80a25be50db49046b63d273af7b916f7552b9164e44e6eb8
z1ec1751c29e635c74c1ed466788c4f6dacf70e263488b375174e420ffbe917eb3d8f520d9218ed
z115cec2e7ce421e4fea4b99dab4cc39697990670b5be93190027e00c9d55bdaed1c0b89b89ecf8
z549ca945d13a8c0dad00bcf83ca4e84dfc5e36c246bd8674a29a06cb318853b985edfc718dddee
z941973d2f0c02f8dfdc2943a553e26431f9a1185f1b26de27d3ca7bbeed4b20a4df9c59bfb0aa8
zac40a6ca497977f12ba5abd4ef012848ce628127d736228872677c2b96cd4a219004224666cd43
z0b5b82c7b6b0ec6a44b2c31302e38d198961f51f655156892742a52e19378ba16a416d88a4c1af
zc2d966ad69a62d23da48b6abcaf1b066e0883750b495daefa14beb85a311bb1a5cfebf0a737f3e
zd918a578cb454964d71c2ab329c965f998c83f430d6b6aa98fc03a4bf9725c684643548a34dbc8
ze5cfed2fdc3786a19b206b5858428c274a8dcacfa8d160b638bfb7e4a6fb5be1d225cf5cd8ca79
z256c6ea5e7e162a9a34a78316434e6ac4a085a5c70bb788775ee47a55c437dc7fdfcaf2cc32618
zeb44ab5064628e42bcd4acc8c1f3045c964702cf69a0bf372bc563b6a90fa328f4731d1795d0f3
zaf37d68ef16f87b30dcc165c47491d9fc66f26d442095ef77cce6b9304c385f13dce9db56ab2c1
z538cfa1148652f2d8b9dd10dfb82b19adb2d59adae5335ebb5c878608ff56824fd27927126e7c7
za0896e0ccef09e74bff91f06ddddc0434ce25c9ddfed788d57c0041e56cb916482a117d650e350
zc82c04da2adb187c68d301e87a3b3ae12cb7863a8892773de18d7c28bebf9f029efb39898939f2
z3960dda160e0f6d04b2237ad090b53e50ad4b218be41ca116da8d6a7d4cadb98da23d280a59ad2
z17f4b17a3e3c6acf4284366e2657c920814b12a90fefcb52f660da3644a0910b5ffc880c78dc59
z9836d5a86443cfd49d15221356829d89d5085b688627b8cdd419ea201357cebcaeb182387d28c2
z5bb44011972d5820a1fcca517e243c806768b693068e1c4b62d9f38c0c17120d7cb93a24d277d2
zed06b7b0f837244f57ed7ee8e0d9aa4f4ce5f9bbfb13e81e1f1d6571f25e52868a73d2e4e7ac9b
z945ac6040979c0f6d2a7946769b177c6bc853d044dbef7e66d337060c0d5e5b8a0f7e316a333ee
zc18df529c88ebd54979d06323199a8652e8cc44dab3251abb684361237043179919d35be4adc79
z5b500332fcca9b7dba2edb5445e9cdd5b8f6e4292f4384cff664e720155875247c27d7b0debea2
z5b46ce47ab2721336e19a5b6ea317b7227e28beb5d26607ed35d2374a8cc014e4fa475cf7eb04b
zeaf2b777bdb48cef947a56a63ee404abdd784a8f6ffb20b3b28ab439a02c3f18ecb58a9c59c873
z67d6548befd178a41c760ade70d4cc58d5c6eae55ae5d5d47e6e13195f098051640b0a9e350b5b
zf3981f6c13ebde5f5dbdcbea5897fc982fa5a52c549f5c2c03bf4ef70bd3cdbce0b5f0f992937e
zd570f0c28ea9b0b42b31129e426c5a2675824301ac7b28b77b31ebd4adb83baabfc25961a5504a
zca20306a865863e5e62c14fecb4e1d8b26d4b1e0e1f92eaf43f6f49353d3e254094451a51d6c45
z6f2ddcdb1aac9613179ebf5aac87a49a9c237844958116adba85742309bc0618e9cb398e753c1b
zf409cfeedde666ac1fa844d71ed0208fe4bb0835d64a7de200b20015c6c840d49ce11bb4aa6cc9
z694421d88695b5c27c1f2358d6e667da40a0ca5309749f08e92feafe92f85e1d34d019107bd1c5
z7969020e48f6eddaa5b7f29257583dbafdd9275581865e3bfe356951bfb712760f8c73f7a0db08
z9e1b340a7e40288e7506bda5b46978a4932c1730caa2eff8ccd0af9f0cc572fe7d78247c232af7
z7affac34003e4acfb0fe46500428d9e4a7cd86590225e115b63ac8fd2af2b7044da2240d636a42
z3ebe433135d94350a03e69a7e350618ee59985b27c660b16310ee804bec287eaf4b3ef9f5b2c39
z9fd23ff52424cc9fe76c6a7bb29e6f919015fc63bd6f837b1ff6f67adf008e90221772ac601f35
z40a9eb0282330c3b2144a05b3260e45f68e4882feea2bed787c61f08cff758265bcf3c6ffe00b3
z55acb9f9906a8ad45a8c507809a08abeed6a30b393dd0facc059669a3b4739539f7554ab5c5689
z468c42406cc8d1b2e9c4bed3accad81304de9bfbbf85c616ee0e1bd5fb2a90bd457ab8f5689805
z45ba3e6c84b33825d91d0fd8db6b4654c36b630f23d7e3a82e63c3ed1828e2a2e2da2f4df0f007
z5b00731439d8c69b3a8814262aa406a5d761f94fb8cbe9f75b05187b93daea930f339643e371d5
z59fce5b0123416335689c1a2fbb217a95c1609d4b5438b646cadbccaf781b44a9a94b31aa40e21
z2859d4a50b774f7f9c3ef7fea07271d57ce0b90a7b61e048271430ae2f51833f8ef709d336ab8d
za92ea3df92684d0c995bda286bdc4fc5bea5394d6de14993566bae1c65556fb80bde045312b189
z1aada89d7915e4d044988428631164fe57d7c3c42030e999447b6abf827b54ddff6f7c0facd8e8
z09ff0a260883219e2e9f14873396278bb0d30451da0c00089733f3283bc68f6d671710af6facca
zad8cd97b82062ffdf5d3d361f2a7e0249b6eb9e193b378c3270936e6760e75e6567389dd499481
z4bf04ca15449bfe35eaa6f41c85a7bf117a3e53cece34577775d970fe101405738065bbe8312b5
zf620e7a420c70a28794e4979c487e4d2da1f730ebf0f41d02cb562a3f7c8974e920daf739fc7e2
z21175525ee722b18f077456a0df58f15b3aa3f554820bf9b1fe33edf122f71f27720a9a1d616c3
z3aa687f034a1bb31903407d36bcee287e6af7efc0728b2d8b877c71edfa190564cb498ac7b5de0
z642e5ad2e3d91c145873c1fea7b2fc6bc6c873d6d4b42a780d02642cfcff8e2633f86a59e33526
zd8897ee8a63342704306722f3c846c0da6bdbc10d2765515fbeba4e1270196b8a28a718e1f7bfa
z79e78fe50398527f4b24b936fa5537988c8bd91120ed636c43a5b8445f89f45606dc59dda914fa
za1d41b32346fbd68ae16728a32c6f8456b0bfa8944d5f8c39ec4601d30090b4abd744ece590322
z4a185da77d7e2891e4b2d88eae6faada16e1e65b7e36f0fcd9d31152c9c93a8816c9a5e5e5fb1f
z44238587aa0c0dfed5f0315620e0f37bb986f63f2de878f62749432ecb22998fcddc7cb4290cc3
z7b93fd897950010d5f25693d9866dc808ad5b3f03f0a5d1f02ac95b2fc4369cbe1642de0a45274
za23e17675fa50126bbf2f1767d74f59b4f6046118294c2db109f0b00ebbf0346dbff66a486c3e3
z6b729b8cba19d309768a0161b56f94b2fab442b1a447ad3377b209c7de6208557b3989eebfdc04
z5d3a2f98617f758ed84da415bbe296da49bc84e3dcd7f8cf08684ae3e2bb626ce7e013977664c1
z673aa91c525a983d580e0079b259d63ca02fceacd8bd03c30285ce273064984f13fd08e0da0bf5
z16ed002aef598130d0ea450b18c9cf4b3708824d8210b5cfa5d35e7cd64469ca69326fb9276d3e
zf062223097b3ae305bb5ba72d852cec20e7f0269fa80903cc4c9b8c6743fbac11c809816a386ce
z70f547b8ad1332617ef882b7f286276cfa84dfcb8e50445f9dd5fa22a9ad7c8937f09af50d4515
zbc6e2756e0eb2ffde5f8569c86304282a2ff3f95db6e49f3519ee2aaed03d35662b557871e7364
z84b3a215cfb1260f42cd8b6163949066a06d6cb292a1aeda8f161496714ecb37cf5487cc2c9b88
zd5618074f234ba7de181828953d72ddd127f31128f9f56591e6bc0109cdc55ac9627b12fee228e
z98b4a922fe8446ea552a7d06f4efd4db14374308075c27e74edf3c2c6f643d1919e2a605835ec4
zc1a85fdcfa3cc4224e12b1e666eeae776547be250d471d6cfe92899dd81685450875416a6676fd
z6a0d9c0ee10c107940b67898a9e18f2545bfa6f9e7038eaef20365934d6e293fd17232f21efbce
zf76cf7dad85e94d5d0dff1edbd9245ddb32fdbf8475651029c72507b3ca3b0a08cf7ba8cb94076
z8566b3fc55e30632c103797dfd18cfc5d99dfdc7b5492d162b2617218716df90053eed5de8ed53
z04c10cbaf8e564b0a640200db3420a920f9a505283093df8434ec4727ad41943cf133ea2efd43d
z4ed61d580ab57bfd298fd1374f713f8920c4ff3b113a5dda343326b276578654a09d31ce219f6f
zf4d4081f23925ab272c042856b1acafbf945bf290118552c9a07530009a2c76e1425b701825866
z7ec096c087a19ce373211a9f450e317633d67e7aa2db8c0f19a39e2e14c7c3aa79be89dfc87614
z565ca15c4dce872a0fda6a318b0ca51e3de2e63dd200614711fc01647468a8235a053cc9d4fbb3
z21e08222a9f9daefb3eb13f6362c0624a6a6069386c780c4fd5905381ec5c6ac85c4519682c3c1
z9421cd815448d75bc283539ad046af060a4aba635542cdf52d23649a4cf066de91afcd401f8934
zdd9fd0c87bf694bb05b680b158dbe38b193af9733065496205a825bf047dc351d5a851e0b3d3e9
z368c6a259eb97a6c206db6a7cf14927e5ee2b6f81de755597e75111f33bddb83f01c4d8a36cbc2
zc399508c65e8e8833acdc1d4d97fc4248728eb24feb5b6cbfc114c749834ced5408a163ff273ee
z64706c36e49ece817094e841edf8d227bb8a4ac67aa226930913ec85adac8ecc5c92430fb728ff
z24ba7e7dca8df58d4098ca5cccbe2c63e17b216fe73335a567dc8aed890b2ed48a2db001c7d866
z7d9aedc5a9fea037a67a4b3de394f9871e6eb8542bb3b272922296838ed0878a80f28e615f1542
z79bc4fdc4dda1f5335725365b95e9f01f0c9c6eb25e01bb0769cb245fe371cb6d760e5f868c7dc
za8f492cca345824b1dba5a23a21e39316181e444239f9aff3f6d86c644431cfe93f2c1db418d34
zb5de8a073becbd6aa3e5a8ca26aaa36c3fae24b0e6e2e44a40817c1660c7da6b9bf7f8f5e3db65
z09be5a8bf5d7a26c2a5ce7f87d8c46a6bee86e3269564d4778b89dc117bc4ad744f68b1f512c39
z745a46b2aa3f9c4c939f766c701bcf3c5291f982868a4080edefbb26bc05f64c564d678edb2b1c
zb158ba0071a290744193ef585a105999b1fa86e683bc73db3535c2bd630fc71b12fe7a907e47fc
zc4474e056ce43e565a6329de63978c1472ba72f47aacf0b002aef4d6543c6d33a27c7b244ad87f
z08570a6aa0963684f9a8d26609dd237f194be0ceba99130c6d61e406251f6b7ae92d5bc25682de
zf416d4e35dfc762a6b1dad00420c0d44c5f34d4e9a12a40968420c9bb6489628c27c351b8ffff2
z116e631f5f24ffc3079c3e8d773492e0e425e9beed885cc108bfb433627401577eef91dd35bf64
zeed7b2f6c257489cc68ee5e1370bda00e499ae0d2a4612a39ac7ec51b9526331a9e60d222397db
z88c32257976aed51a9e470aca4fee78b9de853567e6265e4a849c310f342c5c5a8b0684e161064
z9baa09ca9e80f8ef2a6657f0b86d11499fd067dada3f4d4f5947441252625465ba885414d8dcc4
zfc8faa32bc212f6f15dad4c94f72876c2b06367b80c16d2d1ab9702485d960904d483093116f1a
z670760f127caf3c321bd638b99b65ef1cd5a7339fc61bfa0f49093227502e704c899245bbd45c1
zb93866a80f7908e9a081f82298952e5ef6c95144e25cfd3429d9da61dd679eee798645370be31c
z959e703f18d9404e82dc89e76cc790f2477f94a3139545871f817844c1403dbdf4b83f525d8be4
zc86e3d0acd01a8c8eb0dc64e047189efc7ef66c8ab9c57616a1161b2f1c39cc8ba639076db08eb
z9867075c874e0974709bbe65b98798ec0fc02e36b325189a3b5baabebeb244dd04b06f863c4662
z76d9a199825620c4909a051055c9b7fc751fdeff541a83896d03cf2f2e8577f8698e654de0da20
z09db9bdc4de20d39d86e19ae2436c2b1c23b7cb47135cd78ba82f76e5054a7e509e1cb938907c6
zd316a0030dec7eb91f3c9d686c7d4841caa5647f884326327193a5ed2d40fc64a3d04aa6dd7541
z1af99fd45c011a6a5adaaf8b747896daaa496d36d47bf1222705af72137f595f0b1e3a6a53d53e
z0668648896318349e7863a03240a9f1a62c2376974bf19ca11df387263d74fa0e614b2a2f08e12
z665069c802466f556ce17406888d1d78b73eef69c5d2afe7e507606fe79c9adf87cedefc661992
z43bee64b794faeafa2c1256a6e1ed5053bf1aeb210535c623b8283767d694174874383bba817af
z2d62bd67a27357d5afb915bc2b3b0e002c956ebafc901cb60087ebd8b57f76ebda9f459e86fc4d
zfa788f3dc461ff47a61779686529a0aed09edd2d0c0e7795394711118d3afdbd6396fbbb5cb7ce
z891628d096752825a71935378b6281f76acebcb147009a1e71f38c338fefd96b50fcbd324ad55d
zca9c8fc1170f41049dba487bb0308f234a1d0cea8843f200094c7a012c2986ebf00824c1dbe6af
z3903dd21b122437a764d7cb0573c4b4538fe47ed1bdea0f788950ab0ece82c9aadfe9a25e5af9d
z0d61fc0c16b5f1920f162ff526a519257025cd74b77e2be5de7b270f6a7b1f9d12254275cc52b6
ze2cfaa0ea2afb01d66f34c041d31954bd180ff26b04ffb1b2af2fa7ed8b0d2f053e542a618e032
zaccf502b36d32a5a0477ee76b1909f5a2b17645f5897865401feb810819dc72b522c22cbbe24d2
zfaa477f6f1a0471eb833189a39d3aebe0190353fb60d696eb709ac558b675ed0ee245ff1805fd4
zb42b7e40e069abf9aa94038ce9246df6832d59e29bdb4f4600af9ed491259394e99c68678f7fb5
z3a634f18d67744ac077556c9521e2d1d4b84784763ca96491bbe59a78e0d459962869e1c8df051
ze145cb7e1ad693cf1f329d3ba1863e7b39817cb7c48871fc5d15cfd1c72a97a5e443c2bdf1c3fe
z64431140377080d486eb6ac23add2dc014bca3182e6fb281000dec0a0b29ae043995aa2c5124cd
zcfe6935547931d9fcda6794aeab519cd565a553ef3e8f4ec673059e91e60cbbaf5fb7fe0fd1f7c
z7a050062248dd4c9d2613abc71cc927530d58169f47db34579cedef2899463c1a023f8f5d37ebb
z047440775c84ffaa7d5a1bbbeb49582ffafc0a9474132397ac616a6e9910100c7b720913c18571
z00c659787bf12af20b7ec7a7ff5df133dfbbc7c490af776da7b2c8ca9e2b7c052f9a58d1ed8e94
z092ab549d5f2027bce96158a0390c53683e2aaaac666cef7347b0ccd557f88cf80399520809baf
z7b2c31a40f4a335fc997bd65371fedb41def298c4593de1cfb5112d528a5476b865e4da17af9c2
zd2a68a04a541cf14114ba577562278489df9b627fcca623e3542d9df2fe4b65ae867c423e59b50
zc0ac9b78e7a3259e5a3fcbfa9b1b3a5665e7b933f3140dfc8da27881476d490b11fd48d7e51814
zf4dd8fb9a595f85faab9319d9806cd29cbd0e083e0df2ee64ec6175a44d599fc3de1f248981b4f
z6ca91bc479c7f658bcb179369e0102c1b5c35f95449d57300537b3dc39b652efa41891222d31f3
z5b83cb95da8d55d324659593a432135595f9965758a2141ea701a9b5127746aeb3c5b5fdae6bf9
zed0af60eba15587fe4da04a80f4c16723e690d537ba548c2b966eed82bad4ebe348ea259bdc58d
z37b11917372f4d1849b13069c41451a6af581be54d40ee858f8bf2bdce8c692acca3de3a961cda
z216e36d78aa29bd10f6cbf3275ed28c39c609d99c172850b7e6bd066b6c63556c6490fb49ad438
z5c5019ebc5f3771aacadede3312b2341ce2383fc6101ffba1e19bf8fff86acf1b47b097c13fa6a
z48faa7765c2ee8d95e5d09d288ffa37783f3c140b47d5d17c31c4fd0e773d42d88248e6f270f93
z034d2f985ff553c0659bf1166b5e3a898e8fee766f9ff171a151ddc78ac4d1f3b3603b13702b46
zed9c0e107e2907b92a3aae1dd7ef762ed283f812d9587a0a69e2300d9e39d20f37caa273a8e09d
z8623ec827fcd6cc87b8fddd25d58be017df1d26c4460187c0ac12459af8485057e5eb991cfc661
za5e1e415d8371a3b34fbc1d0d2b112c5f9ef871a88bb987d0e5e29602b2b5347a64b121d424511
zcefdc2f7b385fc2adfe5eaa7666bb1d1d00ed335e07167c9153c878bcd39fe8e7280134d7c7084
z0fd3d5e627f04eb635871eb6c7c086af115645b87a81630b34d565d63f4ba78e145e237aeb94d0
zf5b3acfcfcf522cfced13108c69e203a7316387195d222aa176eaa28829c2b3f7489733413295c
ze9fbf7471ea9dfaf64b01ca3451f19d18b4e5504e14ba85e39a42ca36719124fe76ae419fe7a96
z89d6696d3ae32dab00490c401c77948318dc861e36167669bd9a021abc86fcfd1f3ca2c90b946e
z07d12d6b6b410c02fe798f5c2ac5f920b07dc45d0f11c60f2a0984eec8b8bdc9cc733bb912dcd9
zcd0ef7911aaf723225b9fd18604b57b07e51c44d4679a38aa84d8c91dabcda4b83eabec9b6d006
z4e2eacd734dd01c653e1789ed53171ed3d9297b4bdb77e9cdb20f90431a943bc78a1d770578016
z41c121eb47bc2126a71a0d51d455ae177535181c1bb3a309a33e91a6a4b9aba93ab3ba19f3ee24
za3a859afcaf287db69915d3169bf573f9d30d66a90be6dc840bcd85143b7320d92cc0d788ac912
z36910ebdbbe60c5840c7e1b4347f717421528f0236ba052a3b124472f03d0861675d0e8ec43749
z9176abb0808a735fbd3cecdc22889afa34c5a1b833c88452f6a444f4b73b45ccf3a0e19032b98b
zef6202f6964158e731cb9b6f26bd07a49a0bcdd72f7e3a51834cde00be5d635529fb0a9e4e5d86
z9615f92f6eed2aab82bcbf38b99cb408ee13578d5778d0997d7dd0997c2edc8fc42a20cee930a2
zc53fdf59bcde201b14cbbd145ecbb89c66b91b02ab418a372bc6e7a088d3a264679efd9f68172f
zab32ae482bf493e54dff60cc6137317d19cff13738bd8b4c359af86293eeb86e9dea52d7c29003
zc5bd4dd684f54bc4ce4778fac1c6262cad2e24bd53cb465a21b2ac06622e406dfbbecb57eb6c62
z90149322841fe88ccb6291aef420ad1d1ce038a490a4a8218b3c13f1d8e75440037ee627badad6
za2c5096398eeefae61aa4955bf74e05f43aa98ab3ccf3ca8aee3763726f3c70a42698e0073fb79
z2c8820946181484716de83e3e60adaf2862761e5155066b9c36a7f9a3dd9b4cd0d6d582832650c
zfe7805acbea5dfab642a33d8aba5ec112ee0a54e9b4d0536c98703c3a496aed1443d0de378185d
z2b6b55c0738330aeb438e91394cbae8c174f19ec4df48c2eb550cae009814edeef05dca0084c95
z2a589554cee517296715d767ff47529c5864d9599fc578d776d9c166acda89a177af04ac6561bd
zdab41a775a4c316e7fb3c242a594d90d357f1150096ac930544fe98949bd73921f7e5510d91863
zc96cdf89d2e8e333140cb340b98cce8fdde369b1e055992700760382fd769229093021429c20c9
zc8d34abff19a213e7ac44341bffa0e18998c319b3c9f6afcbd6f76b624fc365097fcd05efca2f5
zcf6a917e1eb9c6a4dd4326a250c38ea9e5ec23ef3e238d680eb63f470dba238d0104200d9acd90
z699107804e1e6032e78720110017cf4f2bf0820a4292575c0f9bb18f076842aa662c4d082bf020
z44ce9b4fdca07ccd5a20e93444b383055f7a683381952b725560ed9c1495df81bc609ae59377c4
zc0f65fb592a12d6dad4aae7d32407269815f313e3f56d79a971a913e79c7cf450d6cbf08529ecc
za51f78c36c1d45757ededb928fc6507500b955414dca32fc848be4ef3a4e194fca5455d61ae00d
zc7ec665b913af3fe4a68d41c944801339dc15ee1c86a863187ff8bd4337f31c58a1e347f2bc010
ze98349247586730939642241575e9ca2eb4f3352188cb7627a29545b36ac3f6da1f8dea599ac7d
zbe18595f4caeb00946bdbf09e167faf2fe3a84e02e9cb8e51c9a9cd94f597d916cc078284bc681
z25e139b2b0901f0c4e04300e9b466ec9c8a4005f4560d794c2ddba99c1805e04258b2084a5e9ae
z9f01d4dba7dc2c69ececc76fb79179782021b60ac1fa410931d05b8b0d16f4a38b2deb602c5987
za85e16a6125cd58b2536fa3a5350a14d3e17918fd0079d7725bc8b68619eee388bb951cf68372c
ze8c9e0a209f4ae6733c58dd7fb704178a06284acc3802806118cd8f563928c3dfa035ef7e332a3
zeecf0945dad583dbb6860f78df22aa517a86e36d48658f123b1ced7db7f8ed85f64f53a28adeb4
z05bc4ef5e0143a96c740abdfbae90bf768f6a8764704db3aae6e26f70fad209170bb812c793c60
za77867de27f769186c573d1b29c594ce41f94440ed32a82a8daaf091534116041b70e4bca46bcb
zca920204adcfc1fa51a073dd48c5245069b36d61afc46aa44afdf8b4929cd246fff1905d9125f4
z5e2c861e9f780bd2f26422ab6fc37f8f8c4e97f387a4f17ce6da6e6302789067d135aeb61ef6f9
z1c6e526b4d8e66e96132d543a671acdb8f7757213b67a1cdd8c49a30abc7053665e2f0572af186
ze0508d5cf9b5efdeb3eab6e0255f44300085ad0c4f3c16253b0c41ba5991abce2dee72822cd6ca
zf8cd96a4c43f05f6507cc643a3b1444b424bc86b3b22133c9cff90f290d4686f230cdbf14bae12
zafcf304676ba9d1dbc4e99cc45cc4e72ece6e42300934a652a88ca9c1081011f74157d99f87b50
z1f1f680a06f4dc99f0c6977bb74999eb850b6269061a3a5840c9221fa5fc0e833efb8548a7d294
zdf8d1ab8e41d3166cf2a4a80dd2cf31d96bfff50f0c4a33e6534914827a8cd8a65af64dd7ca308
z663d7febb82e4b1c6d2f19cd121fce6b1dcf3e2733dc243d1a7bf916119ffe6aac92750d4b8b04
z9389c3f6528c1847fe499b517e1cbb12ca06639e9ce125ea3b9602fe41fdf48ed5561edc38c58d
z1b9852c49ac95b604d13482e5a9b9d77c9b98458de722c855b295353bbacf068c506d5eebd883a
zef55caf1c0cf56b02dcd1444a585f4c54c4988779c54b8ff058fb5272a7471eaab8fd1c6ee1396
z90d772749d3ff1eb34fab35f8d34986c1733111779908b9bff619a9015c45563a822fe30484d02
zc86bd98fb2016d579e48d5ec9cde675a370b1554c0ce2e2312b9a8e0cfa71b3b9eb215fade701c
z5a91454f93461c0e04c8c9884701502788626efa0c61af4e497c04f70b9807a6614760b24ab6a1
zc8a5e818067734ada07eaea2acdd00bd03eb20408e23c711dad49fbdd3039705589adb5bea87cd
z7e78c17a7a62d49167fb9cb9144a9749656db722a72bbe206a9e5a208d8f1da5d41203431b8c3a
z7c1d350ab88b3383640762200493123bf9cd79561872d65849e81fc4e1dd4e0f103de44fa8901e
z9c43f386a522277ec07b3ca97d83f7f68757a0beacb9eebbee44452c15b02fbdbae0e6d1f9cebb
z9d8a9ec06d4fc30706423ef084e82ad0ad5abf7363b0008ea873cf7b0988c311a40e316f251fbb
z5d935229ad35eb83cbf398091016ef6a5c62a9098659323e218d776dc98ec5caca5701226ab065
zd4ecd958554cf90387301f783c300a64d4160ed44885787736f9e2a9b5d48b0726a2961ff375e6
z577b09ea6451952692b02ecca6adb80efcdbff9654517faab6c29d2978ed862705a7aa2bd66c3a
zb460b5d5b6811d0c53f06499ecd2904307c7716de34aa8b3e82a1576659418de675621720fd7b7
z3dc001279caaedd13119dd6f16d6f2cffb5cadadf8d5a6ea432bbcbce2312a867ac5c49d0b6331
zd7e29e64e37dd404630e24badb887230851dbed75befb196021eb674c91292d1f3cf37160d88e7
z06f09c8b2ac631635acb9e76ce526096de5f116f3f778fc38a3ffd280783e794c419139be95fe8
z7c89351326da6ed11f98e2383b6580f961f7049850a6648a047005ea1e868237c89492f9703f78
za102969dba4339e38b5310996149ab7fcc62bf44f8af9d169115b531cff9ad7d87d05bd3eafbc0
z938b5558aa6e74c32aae86f17c8ad15fff847760d79f086a7975b2ca8dc6f7a1fc7afbbbe84841
z00e674bc9bc6ed9f4f27d119ee773e4552fdc377bbd15ee616791afd7e3e013192bae413bbf8f3
z6d7f2617978277feab49410ac9d9fd0261eef18c176be8a55da25eae68228c568aed755cefc828
zbbc2a50c56a7c8167cb3828d1da56575623faf228dce5b483ad13ff64873d63363ffc54dca7d54
z783533fdfddbe8ccac50fa10df049ace27bca17e72141cb7c185bceedc1891f8d22c30748c35af
z5c46aee873018f06e4b5fa629550ecd2af46faf12008f4e38f9326a44637000b9c57f32530d0cc
z9376d7c4798f6366c7edc505a45ebe1cf48f0f7d3d4e8a0210273d0497a38a658fc397c38046bb
zc47e8b006aa1736918e0a8bbbf37e62deddd69a63a06004348e99588ab7ab7e0c15961df1a3717
z7d6987e042262ca7e9d6c9d851cf6ad92e27b369f01b9a7eac394ab9e6a745f817e4de41f9305b
z25d9e4cbb5bdf3c23bfc68fa1303f29ae01a9d3b2360900579e292bda0b989aa2f35265b16de12
z6a4f80a3dc710e59013b22c6a2e3021aa83a8c791c870172d6c5d9a0d75894053b1edf652c3a66
z0d97c458b72934d345e3f6e60f3f16b72db3bd3d834f43f38d8fe0187b7c37e55f52453cc93059
ze89dc1c522be0d05b49e894d0250fef6ab7947e03ec4de7004b8f7226072d0e82d531bb403def4
z77f740676d541a493da697c6e827e8117f518f11988d12712fbe6d272b59686b2a560de0deb545
z6bb56947815521f1bce9f04b5eacc7c33016a0c6bd6269b9b806ac25e897d4f34fa20357a30787
z16a4a62fbe5f6eed425a308b409cb68236c0342cbf96b08734beba6923354639e28844736b7fdd
z53f2f1dc664efc2e3860523db9de6e426772c9f623ee824957b21ce3f47539131a7af2c707773a
z304e1d4d20e4ed4c4ed75a3df31f5acf3eded40d2b5654789612348b09fad3178dc452a06a7023
z04bdbc69737415db17c26613590c62bfa441529c3a5f8834215529a2be593c1e3a696f82cdedc4
z54774badeb10f9246e7c35e8c6432e4fc3dfbd5e7425b3687a82665a5c66832bddba7f91130edb
zdb478552cfabdadbb16b7e2af0e086a5090430ea2a277934a0083413490d04d078ed30f3a3a4d3
z7874e160b64552c70c086901d90ee369f25762d166838744dd175f8af7bea5814a02c0bae963ca
zf1f84f7ae1e690c642fc300740e3067177caadbef33c158626a31fc12a83a6a41b33b262f19bc8
z938aa84e2cf626442e93c80870521f5194522f497d06b62d3acfd293e614ac4355ec069a09fcbd
z2c863781eeb3cdae6f44d3e946d52d91c89f9cbd32149bd86951fb900757676d5084ca36429721
z0dc1d7b6be87957473a90a454cf890fd6bfdb6457890182cc40846a3f2c7c13b120d1bb2facfa1
zc95e380c064b523b89b4345ddd5443731edcaaf20203ff339396ac57afe714515d0f86d54fa8b5
z757b691a711a49897983daefddef8fe8b149a0bffdb8fe97629efb94ba773eedb612daa191d630
z685f2db8189c93f75d63824ce7ce7d8e65cf854b4fd2f4d4d16564cc5cef7132666fe2589c6000
z3acc79b52ba4df60939a5d2b7f33c8b6af03c09dc694f61ff2f4964404b04a9fe51b71765e9096
z512b149f5202139284e72ba7bdcc2a19187c320b05871fc81c6a43aa2f3b7040cf34331526034d
zf535ed3ac5bf6ffa352ed3cccdfeb8ac466a9d4300d76cc871f95b8ad123e1e9c7770159029417
z74f6efa6cc01b4fea1d2e091aeca43c456f89b27d8ba31b071ea258b5e8aad20e4bd42da5afdb0
z14629cc52988c5a4e684fd09e89e732974afd5d4ddc6b27318727e66e1c8d98b4dc4b2c9e79414
z384a1bc2e059cf238053a55fa2eb05ecb41ae04487aecf463e7fbd2e76c3cf2562b0873bc0d10e
zf703910bc3d87252bd2af82b2b868825a9bb1387c921de0ebeb87dfe69669cd8832c65f1559f9f
z818fbd70f1ea78d29db1498fbc75ebe362ecd4a8a2ed9f301dbe944f154eba529560168274ee7d
z317619abfb6306e66c81b5d2b40c97aff68e15f7a7b55e6863c27181868f9663e1d94b040c0bcf
zbcba8dfe8155ce782a389348b9eea0e43a61a06649ef448d1afbe48778714c14c482c9403eee3a
z813ed4767b07dbe66dd465f6c43e2d27993d5d131f77f1af0947b2b2d18df4fcb74f0f8dcea9ff
zcac096896a181ea7489ad91cdf6c36e86a390d7d357c0a67febae9e8bdcb9c8cf46989d8d5c597
z10ca9c022bdcebfdbb77074b5b46e014aa33ab67d3dd8e348ee9f0976edb5970bdada1ff5e2827
zde78b0521a36d7959280a8876d3cc941846bbc50e15a9e37f002b840249fbba11d339b05b2c5d9
z3365d79298738bb1c5a56c241dc82952844c9a2825f555f6030f22a47f7ecd41fbdb8d4990d20e
zdff5bd756c58c2f7e527f51a17c843e26948dbbbade379f395b7a5afde976d2ff27e2c53a8a890
z1e621cdad936bb09bc1465c3cf6535fbcef7955e6d2b04d24fc077d0cfb10bd39f1901b00dfc8e
zf40ce8f187929b448df424616b33442d44f62fa9d2bae399807b7dad74232059b87d88113541f0
z9a48b497a392aa3155ddf7239c4bf9f65e9d60748e00757a422298071e4b0a8e8af2eaa85af5dd
z791e6e993d09d25bf08e8170238591aa36783b6bbb9c2da5da531f0c5b44f67678aad337ffc399
za8f4b882e0f65c05b52e6f7bad59cf35cdd2a8de70699c3c9f10a0af026da41a70c29d37e8581c
z5affcc2d25e7157340c38a5b0f070955b42b7dc06e2a7b1c1bf8c393e6683583f6b6707f879150
zfe0a3f664dbd6ebf6106b7514ee7646026892fc5ce2be78f2137d00051a46fed0409f8c6953a0e
zc65dfe06711c6fb3124d36b7d630066e25b8c91b0a44620ee338705d2ffd4c9b160dd7d9fb935e
zc79f88a6fe26aa0bea353b4ee21e8b0ed2d3d52bd781b3faceda1da1215f637ea8bdf1b7a1bc02
z6feefca0ddb60fe5e328e9a50e7648df30301b0ce5dcbf632f228a73a39ce21e1a5d9a11903a32
z0619621c453bf371dca4f2ab095f9f267e524a2d9bdad2d38d2a1ec8fc766ae9a27cff702d6147
ze67bc3adfa5a4db4a4db248494b5ff3c13f0fef950eb7cc87d123651132258f3faf799c878be9d
z1974bfaab5fb16042211f11db31215f159bfa7c2ec0bcf9f5cd1b8bd70858a7bcf19189b089890
z593545a1c8d77b8992cc3689c50c882b0a89e07735ba0c2fe171b9a57590c84114db91b74cf492
z3685fae0c0b357da709be7261e6114c0ae2e9e4189ae172039bc078a07304d75d209de68d4a839
z0ca4d33decce4c22474c9f3a9edc46874cf2adb403f3ba03765f97fafb0b3e06f18f72c1fb7a28
zaf95e4b5e32230fb93888a945c5fb914e7245184022fd05d8c81fa71ecc731e53965cca01e8c5c
z70ce6fd34499cbf3e77cf350b1ba84954a28867f715cfa2a3d75e8206df47dbbb67d1183dc18ba
zb227b2e135a03edf44f2c25da4a664404e91a9e975e53f99cf2a60a87f1c78b4fa18bcc4f924e7
z5856f4da428db5881bca4e2b82b9d95494cd8be5c3f650c631a4514b10094c450af6c7521234b1
ze7a3f0ee4605123f931f72c0641b1b37b7a3afbab768fc2ae9578c59bdfcc341fb90b5b96225ec
z018cae514aaed8fa46d2504d8bb837ed78b34c0cb72fdbdc3f0c03afbed7b53cfe3e5be8a96cb7
zcb2c8907299d7dc8be3a86f5c7bdd18d488b1d96259e0b025b10e395a23bb3a7ec8eb50e641b1d
zf04acce5a36b199d8f54a30ce24a0a4d248c473cb693aced613d9932d0fcdd163d70ad0f8d7644
z239fbb50e6349a27b4720535b12f4a6559eb82dcddf01cd6d11f8163a1d044621d8ec77df696a6
zd618447fd959b8f49aca9fb5c1201f5620a53f758d85cb48d889ba68fdfeff476c63deefd75747
z18960d5d12be7a205f9670e2e6c8b6d66e2c09b098c4a54e0f0944ddcface3e9a322c6312a9fb0
z9435c3f7d18c0ef09c19d16cfc9c394f940d3b33692eaf0f7ebcc56ebc639b2c95f44ecb4f5e3a
z38592546b398e9b4fe156eb7fed9a13415cca14aeaf7ca4794ace3bfb26fa412d4a180350f0f81
z601d94068f3fdcf48205ca7b054847fdce36db4945f6cc2095c7debab46851dfb625e7513d96cb
z6c4432a7969aeae5169f0ff65f17e49088c0b506992697e6eb72cd6d42fd4821cbe5805a0464ac
zdcea7c2654b68abfaae6333f70e0a10185d1d002e56c36d2a42a944e3ed8838cd9a9f7dc57149d
z527bbe7b00254f5fa0d41b149fadff74b255548887689fe0faee427ec17ce1567312b22125ac8e
z32967d8b9c76be2cc1bb874039ca7dd4a79a2939ebcdd9fd1c3927a2d593e75f30f3adbbe8d54e
zdd7a73500de83973673cb155db3410800150f02813a8370b0fbd38549a051e2a0c721b1f50cc41
z66b201154f0f703fe94c6c42d14e91770c4e237ced6a69b112b395688f4c9f50e36ea63377974d
z981633a9fcd10ded35c71c49ec0620c53a37c9aead37994e9b026c06b377af4b49e1234be7c379
z67dee8dc004621ab79ea869fa0fb57e9bf947f3bb4e5a2c5779dd5e31427e2196506933967ce0a
zaa50127b95e60953287026480d9b5469c5553f2007a46ddc99e147c3b5d392003f1ac31a672d0d
z68e4559c72dffe02de648720ad7d47f958ed3f26904129d6f55a33f241e0de37c22eaa8c82ea06
z2e91e8af8b31e98222fa5061ec4c7f9a2a2f907c94c6a3189c16e8037ebc5c961edf3f30d3dd4c
z0faafe1d516804a88b378d9d2aa6f923c29e847886a71f9c4fd67c19d85369b076452058c5496b
z0ee380b163eb0a864add6decf1f8284ee8d1f263f120657e73ee32a3e6e434a89119de3c7b52be
z08afbf0ca8d932811ec74312f2ef373dea23307db0160f4b4175d5853877ed775dae09cbb9bde8
za9a98c06410a35da7b9cfdbada4ef875b62426723dbcbe04ef55d173a43fa72d016332949b82a1
z48eba9241d5904d9739c00813af54f45edb9c922e7ae0cbdf1caeb93c02e69a9b5442536e1db92
z7ddb5a5248633f9a23f58b67c67c0c67064a5ce7431ccbb3d6580f61139114d7cdbcd00c76b2d3
z186e2456aeec9b333d55c59f5ce84de5b96c3d17eeea02f635d412edd703258f2eb98ea39af873
z582988f9abd285c97b1638660bfc51c63357ea8426e001aee4dc979ae2bf373706c2fe6a550ccd
z44a9537df5b074ef180d81918f68a425486e09124f14b407d70c21e29edc30118931e78fe9276e
z98682cd8c0fb7cd86c38353c0394f7167fbea7e294bb5b84b92f9035a7a021434c3236c89e9e5d
z8bdfc9b423d561152371cba28233e91d20b1c04daeaa28666ca67505d1a4d8c58600c8759a5a42
z67b72da103752dec5926286d4261413d4de905cab633ca285c6fc788bc197e8d63cdef1c879707
zc42dc242b979268670dc8809cac96d3a51c9450a50a1baa4591a7e9bde8f5741294d8647cce6a6
zd357d4dcebeb3833ca52b3905cf4db53c9065ff4066d34880f4cb13c1c9c25803d945c00c895ca
za69f9e961b66e2bcb15fb7190a83c5df1f613ecf429a537c33743640af8ab8cc8a22a7b966f360
zfef9b9fdfef32b36f134713c9a0d2819fa622a2eb89f39a1e539209645e4905e1fcdef82c94ce4
zf99b1a893558e3b67b6e9e20a202d1541d0bad68e9f360e5e1cc1294c0564de980dcacce299a73
z64cd3d091285c2ca2d9d739fc93f19b4bdcb571e1df3b1f19b0e59e31e1ab3cf258a762ecb48d4
z23352d306e9a6c2ff5a34dba03888e5da6416560499cb8381ccef7c0ca78d300bdb8f44895c1ba
z9f0a53677662594553d8a56638add172eb82b83a91bc453e7aae425855f2209b2c2790b0837552
zb68b3cf4dc0750c3791d0ad56eecc3faf8642d15ff57ac64b9453a3601d9cd3af655b519cc7728
z454d889343c921d543e019148532edaa69c3433e669bdb04f33d571b5a2a8149ed4897cfa51097
z87ccadd3155d88ffaebd9b38c1115957c9e7727bea62bf4991a15281f2ec93a1a8a940a2351fe1
z38e88d97a4a45fa3eaa05ddb8b57abe8fd1c351151559c190bfb1be92979bdaf63a3440e798bf1
z42dfb029f1693ea2b8c3a8a6d7f5e649979a78c4c0b8f1f7ececaac64e9aafbdaf5d25a48a5ec6
zb0ba0922d8d591196718b6d7708edf52956af41725c098b83d2a9c41b76911679bd7db30586df8
zd812dd25001ff75f9b757e27368ff95a24aa54e33f6f4f49c51f82cafe193bdddc8c26fd3d7c5d
zfcd02a1ad5331427a76f0e83719b524b695bbadfd00ad01fd70cc7248023ef9683ce1295452e51
z9c53dc9e2fc02ffdde8a820f0891d7f8d47174dbe9ade4822625c0b8e3529c51f6fa3fed0a2826
z64e5c4431846c0a0581f1f3b81bfea50e2374b8df3a14c6859088cd97864ccb0c2ae5e4c75fcf1
z258595d8a4e05269eb35725137c26acafa892e187f55a38858ea7f0f27ea82e67b0a8ddcf1e8b7
z81f96b5443299fe36c482a18969642e7302b2a3ea06e310e9d03e99075b2c524023a36150c0540
zb826d601932619f22d0b7708ef40706b6bd5e21d2385315db2577797acf91bfb6c721bdaa059c8
z3b870803d0fffac35e75636ffad27e79b78027ef915103bb8ff92b80a6d45a8374b1ff60dc1c21
z2b516408a912621b224ed8fb4de43a7628a6961ad26b18743ebf615807cb8bcac7d95972c9830e
z8f6a18d3bbe5a2ee2c88c937844eb1f408fb31f3f4cb860ee594d6021397f7743301dc342e47cb
z343be02d2b0860b4cbbcc6d7d80dd1751cedf7a929053e3cc1fd33124469caca7a6c78aafccbb8
z501e2120a9b0195aa926bddeae03911798597cba853475f7f402fdcafeec921152e833b497e2ed
z8abcf113769f35ab124d3c8fc32400dbfefcff12d188712458a693ec214abf09da7517b9c7998c
z8c7e780fbae6f4689cc2c026653679d7125c83ab24c668872c7d0d47652337a8c224e5d78c8fe1
z014b6f92eaa4b99303c1458741ecc74e2c6ff54f80f7efa140c869c6a933797fd88d874db53e29
zc6b05d0231e3adae054f09b3f99425cbe40ff18c5444ef020307413dad0ec5386b99a544131fd8
z8be9293ffc9c233b04c61d8d091a30e73f63659bbc1d0621b13f5dfd63a9fb615b1fcbcddbb76f
z3afe25095b50d900fb301e4e51b1dffadc2cf779bd960ef705bbf21cfdfdcfd145f6a78764153a
z6ae7ad0cf90eaab3e974e16a50338150fbf7a50e1688bb2baaa3963f1a843aefa21f9f08d6e0e7
z4d931df03908c457c6e8b1d27bfb8534a82ab62446b75a52e6dd2c394aa4873a2d9b161e9a42c0
zf834535e171e97afe5d60afa44c25c715ba60399b8ab90e0ea5277edea1cbdd79d89d5bca2cfdd
z3d5b18e1b10372cc4158a9259a2ed8b94f88830b94b393e76606d0bf7a58d70c25763b57b3ee20
zd67d9d08f68bc5a13cbe93b3dbfc3b427e538feb7f809be606f5568da26b9af8a696432086e6e7
z98a0cdf664caaee7c846881dffd72559cf2ed0936910675c86c0dbe6674553ede9ad2c53c82277
zcb20275ca1a5da706fe0e8cdc7acb7e07ef5054165b022b6c5efe626571a698e75affebd48434e
z6966b6e67374a1e3a9014e619a65336a103b1e184380ae4c23f8492bad9fdaa9d3d27db93e8bed
z42ca4644fac5243373e2100186fcb09d06aebf0ee3b6a191c833c90d146fb46cb54133153cec28
zd8837d5503ac01ecd2e1ce7db2d2b31398b08e8646b269231aeb968e304ddb9076e2178d8c198d
z68951705635eded45a1bec1150a835d2c44332471cddf0ad93ebcd7cd75b33b81ed66cc80e6394
z8c3aa3c8d6947a4ebedf37d5839568bd8e45f9680b4f5b80d7c30391fbe4dd45ce26703cf464d4
z29b3b541a2e879af6b18079662f9e793989be043e4024884cf9d9344d42f00651c9de02c163b56
zf0f8764254a3e8412a331b4b4a3d2de118317a11d64f7a7e0b09e590e71c4df3bfd2c18bce7c22
ze47b344b36b713e3cce8f7da12edb3640e2f8a051d7e4a4b9616e55acb2c9c6bd20ed88fc1aa30
z941cf9ba22be70d605b02f62156ff27a234c8c7c4ed75da04835ad92712177affcbbf566a2b362
z2f3f2c2c237d837562bec1f7ce344c95477968a792e3907c39c2250ed9d4927da35b3694b58712
z4bf1ae1fba06d0dda9899149dedb1b48db4c84490fbdf9fe45ba0d3e86e31653dcd35a87dc8fc1
z11280f5a2af8c11b4fddb24b430a0ff8b73020025a2d5859ee0fa58faf0a48545382bdb96484ae
z22c4b552e69e95a52950d54a3302977f2e5d170ec897c02a0d3143e6b2b8a394da806a8ad90834
z19273b4612d9da1a9aa013fbd4417a97eeada78cbdca076fc1b810f0c759a07da7770762ffe48d
z01db175d6aacbd43212ae3f4d2d855bc631ce6b2f2264c8e4e8b8ebfdf6a9d57eff2f5b52d4d05
zffb6e5e46b073e79b87821abc0a397f17287006b818c601797007e42fa12a013caac1bc38130d6
ze063a97f2cccf455ddf218d0cb51c0da232d61801c5565a7afe87e57638c79aa9223e70a8da151
ze5cbceec77b88be929158e41ecdd90df1d4d2eb0d3b95605e9f09ddec38967029f60afea6131b8
zfcde34bb3de5dd908e1632face050d52d6aeeec980349a65c998cb3ac7ddbd9b71297fe521f6f2
z86b20457ffe3ca3a98b02b66d87cb101a813f574a89dc75697014f1b699a6c59f0e97426cc8d54
z05146af1954811efede82ffc486adb02f911bceaf580301c9ea9d2841e151b5532dafe9cdb4eae
z1c9b71a5c33858ef4af142f7cafcd306bfb3ba831cab3649bf41c15668aaef4af0122a0b7b8f8b
z3487b24cde4a241d5092ea1728b71e5f199b7df5d34a6303e321ed200a682d01f1778cbe97e28d
z38602c1541fed0774d2ca8393123dea8a10a56f0f5817f9d8685fa6bbc4320c7abb62563a775b0
zd156f3954dd3bff441f6d4ec4f274e4da8166321c8b1fcba1aae2e7a6bef7615713a1a8a805fd2
z30b7a0fb35a2871ddd
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_sas_link_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
