`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026201628cee5aae21fb892db766c4
zb5b1406e11aebfd6dfacc9da5ec03b70c276807a3eb15e28ec7ab1dddec42388b9424ea285623a
z248195c9f894b36317ca6e59c86f11031163f5f5bfdba36b10b435d36514783bc1c6e60eaff7f9
za2b8eba90f8fd9a9cd7c932ce34efca1757e6b2718aa68644ba032b1bdd74efc688b935cf38d81
zb1f311df3e5b8e4d46dbf459c824f309500192485674c175e61de609f1c94488da73614dd500c3
z680b7fbf510ef6c68927870992ed3376661d943d2a929d90faac51228c485cc4f90c0eee6be4a2
zce41f6565994f8c457ad3f059f0f75d13b595288a756e41a6033f636eea17dcdf0844c8e225d45
z55436586fc78f7c2c04155001676fa3f49b24d3beb3584c63daa43ed80ce015162ba22d33c9763
zba142d3955797e70f433f00a9ae14f9d776b76291d31153dd23eef201b698c8aa3a640b228a83f
z18eedf1d37da4b3680484605b10d0117d140a2fec482eb066a6b3e23701cd7a6c894de53e39ac7
z965f6450c8b1c2aeef13e4dbbd2cfb983fae62219cce167861d4291eb96a217f8c834ac6d8cd97
z3fb107301461c673b573fe10ba27feffb84003be8504678bdeb8fde88ef5ce321f88cb3311d3e4
z3967093b4d555c4434ca75af2749c48959e85d0c3a9fbfbebcebb6494d83e27e01ac4c667ed322
za3b077f2f69273f140dcda394caf8c2a8ce384c08761d34cb8c43346b815742115c69db52129ff
z5844ab9bb4552a6ecfec0617ae18cde60d8143585820e4d584bc0146010ee65c6367bd4ebb9116
zdef9f83ca5f2510db14e3c4c3159d928e5362e7283c09d5d7d951a4de11d8f04b9ed9b2a912a25
z32a274bfce4f54e4cfed937ef40e4a69e595ab44bf66b1acb8a0fa0b91302457e1f4d000e946ac
zda0de85e09fbab1b7f7dccdd45b53c2533a3082f08cc0bafad1d4db319048fcf4c05dc77412102
zda864d6fadb88ed0b50175b782181bfaf3c6501b089c03267dbff78d772e9ad5ec71919ffa3a8b
z0297eea20a6dc97d43737912ddb87addd89af196d58df0ea2eb6596b2d61512b550bdc2d0e25e4
zbd1ed43e87cc5488c07143e89262f655b5ba02a907500c83a8562355b77333d42f2cdaf419cc0f
z052fcdcf2d96ec830cce129dc934b3a9b255ad6245271f167622b385745cb23209dfab390ed023
z6548878399244a4dde01d35bc70f128b2e6766f4a97e2be95d7027c3f59e6df0b6b8e470db447e
z604ed1987145739b28a323859e0ec35945a04ece5dd0836832d2c7173114d1ce61ae7a1b2d4d4e
z135402d9779c00aeace2c84599d517892fd7501d4a53afa9d9f36b658cc40c7d157a0ea4659f77
z93d7870ed99ad90b393d28bca30d85b3e5a2e4638e5b734435c93ae24e41273794207a9bd83d3d
zbb627bc67cfc8c92afe8088c645dc3c729ccac0b64150b5a2ea8ec45be020ea1f60fd92f0c12df
z92a84c7b5889bce16bbdea4f080314a5fae63273d84efc861e3db1e7833b74c9006d3b5fc72c86
z946076df62f85265a2b0b6e89de592293f6539c64bd27b1883742693773dfb4e6ba73ce3f80ede
z00b7696fbe9445902438eec0ec8128bf47230d4b4409d1966fc94454df46a90e7b60681196897e
z61fe55bccaf7672bf403b6911f99e982d14b941421549c47de632e95e5904ebcd1917d2c5a1a78
z4278c6ae7a7a171a0292d393e7abfa1f75b0a63dfaed6c429aadb52e099cceec4bbccf79194aec
zd23cbbd782c50d701ae18fab0767c9ee872fdebbb14ee9282d43215fd1af80b2f3c60f723c6dfc
z971197b408ac21d98cc44c567c6a3724d0a3db9a0f58e1da1d6c87290b19fc4019a2858fd3fa81
zcffcedb323b855fd9937a6dd586cf28f63ddec94e70c1aeb08dd33a6e323976edfa4644211c89e
ze424979b14ab038e2e5295ebc27f7c9eb12f9cf849a35012da657ea66eb23c81c7404db1bb0b88
z98ee0810c88099e0554d7d077fc78cce2411522cc90cfd232a9c67a464f8ada168965909819f9c
za19a72b66c01121640e391717e351c149138ac2dc805bc523eeb65673a051734b218aeeed51ec4
z8f94ad1354636335f16875e7e6a9040a23c9ab8b0a1bbe0234fc936678454984d1efd5e7550731
z7c569b721a77f2a0cc870331fa3a52876335a204c19d6f24044e2698c6303142b1ddb817e9e2a4
z100ba0e26591bc870e95807d27cb736c1c34f421038323a21f2654506feb7fb23d41ca60e1c317
z468c2fc6d0f2df6b5b9df43a89e6802a70da55da9f31bcde5ca28a20f0ca51a1e4999fc966129d
z60d7897e24a541bb37034f8156c40f8cce82a26cbaffc93163ca2db266406f94aa865733e16030
ze149459f92be7690a2e5aafe1b439f6e494889f46838f04b851ea01b4243a9256fdf3ef803399d
z3437adb1b95ae7a698710d15cbbdb6e8a44ed88cd4d7e8e25184193b5cf2a867b68efd17449409
z15487b4c6751e3d452870d5cbea8395fa892d18677059d8de4fad71a8fb09f5c8b2aa0f8c3d7ab
zbfbb5b2090d69110e86b7180a69b3846c879558fe05b139f7392f52a19fd127ff5d499855e4d38
z12fb6374b7b71d78823c56b97e2906e1810b96146a98940e8f60fd75498ffb787dcd45afbb74b3
z3412479ff6f17151d89d1c172f2bce989e15a61315d851edbb53d9a1b8e31c622aba1006d7837c
z9b80756dff81c7794cb14032e8e44fa1c5a9d042742ec7ffedd0418d6b8eea85ed436ed332ff29
ze67c1be075b48c937ec151835b08ceab0b58ffc03fc30e92eb75f78f14228bf071d6dd41ff196b
zbe7d6185517fb1d6a9e93ee0ad15dab1fb31e9148c8531a04f1cc6e1ba7724a3a51c76b13cc9d4
z91993901599cb08b7ebacefff3c8d0589222eb70559ac3d3d15e6f8446bf4deb87e5dc7d09470a
z0f2a403361baf45807c4fdea251d1786a916c63e7707154e5afa726d12150611e3b55ee4b57305
zbaa4f89ab8f976f77c703256dca711d8e03fee6dd1d7c001bd8bee1ca456e0168a3f7f33c44cca
zea56babc9d3046cfff80f4b11677d9f4346593425b2b0e3c08ef60f83fd2574d53b4358cfbeb01
z04b191f73aa1c97cd73d8bdc22e867b09c3796673ffacc9c6a948e6c68fa8f0c9d3a736e22a691
zdb9fa8002f3151f536000991748f331cefe7c2be2176b0a970917c825c0295c731ae309dbb1e26
z4289b117c5857fa18bc213f0738f721fe9b03a7c52a9fa01392e348e13e7957fb78c5aeef630bb
zaa14ec6a9c1c3e30fdcc90bcf760b037625ced920aea5334fb905051034b5f46526ebf9005c1a2
z2cab37ac9a550592c2a8c35470b192a28160b2cc42d6d2def60beb558e5d01d5149d52ac53d663
z185ec4ccdc13ba2ab27cc10453f0d3df47a45dbb57a1815002311c9f5af0344b8dcf42af61b48b
zb0e75929269e8ddb06e23aa9634dd485e0ee02cbc8a5e91f4a250ebe68e20acf826748c2a25f3d
z6cafb85569c89263b7add34217bed12658bfc4c35cb9155b1bc39ddc59be6191d846b7bede9d31
z59117adee5e9a0dfb894cae3861f862d9d65e40b0e56e4b903e07e7ee30888ece8d9ddfbafce2e
z3fb5315e06fae7ffa90d9be58db52ee2232ba4ab70466cb87b5fe7e31e7cb2657a08f584a46a20
z870fb3007fa7bf96057e1ca128acbcbdaf5007b0aa3bbd7e32063190f7f309da55861d792843c1
z2f17b60ba44c9dfdfcc4bd99dcd2cdff966caf7721e891991b30c410282eb51f0b5befa44ae0fe
z44dfa8791fd8416e82aa691d8ad76a510e9a7831c3223d871c1ec3fd0537f529f3eca73b7dd1f1
zd41507f3d9fa9f5f891df1021997b56d4439d965f7539aded61cae241741ae6bf73d3724e845c5
z6810a81ddad475e87246bee39a9e0e4fd7f8e8c1be5e72fa282faec0f1ee21c397307170ee7b36
z276b9691ad80a5d77f12ddfb4e0bc54c2bd8258e8c7f29beca106329e79164e8064a0b068f5ad6
z3aea4423a91acee3041a11436c7710eafa450ca99d155f28413eb774be4d647d95265260fc3476
z8bfda78cbb3631f719e7ae4cb143103691fc1857fe1b9ab7b94bd72ee01684cf57df2a157793ae
z5782afef76eeafbd6a27e2771c67367d64bc7d0b655349aa8a68d98f0bcbce5d31bb008eb776d3
zba532dc6fb1192936985c042053e59bc056a38c9910480a97f201a6834a55011cf2d22942c6089
z94d189e81a95585e1c41b9c1595f6d0dfacddb08399850ae86e91120bf53390bcdc987a417f938
z1f9b34365d73123a76e0b7583465d55e3287e1fe679e34c6687c6f57441d745afecd584536cf74
z1fd7a725920c24d3f618732bf6afaaeb2169b6b93776ffcfadd53675d4ce0fe897311d5f1bf621
z31322c4111a97a02e6bd1f7046c702ff0db612f26f94d0e57cde0cb2eb14c6a42bfc07d9360cf2
zffe0c3037d807a3d4303b7c4c6aa72b7420ead6a5529ddfb44cb57413b5c4e45028042dbb29f6b
z605436daab53ac561a3cbf399401b1046b79180c72961196dd706e52b4660c23226e1f381cd9b0
z6c5ac1889ee3f05c9054d301ffb62348904f4657e2c43f16da9770f781c58cdb2f9ab81faf9694
z1747f6829a2d3160a99e8a3cef4eb30ee14c36a188f2eee6676761bf276dac2bc6108119845adc
z77497ac0c5cb55f50cb103ebcae3f50810906441ef1162bf1160b72d5bff887570865f35ab6fdf
z7282a8be44d962e81559034227672b9530fa197ccbac8cda2586ffa850f3014d2489050e9dd726
z080dc2ed64cd016794d7835d5d187e3c0a4db40a3bd66f1c78b35db8e738c808367a4b16218849
z3b38cb89c5d454870008c97143eb2ffbd751a16b4e4d0fdcf12930813a0b9378408f7209307f2f
zceaa83b6f4f9cca21bc535f4819b91e5b129c29ca57aef6287002563bd8c98b5e6e144a249e87d
z79f1b3bbd56bd46c31c4148b021ffef16438c53cb5475abbd58564b661a9a2d5c22be12a3fce8b
zfee1a47085cbd754715654de2380549bf85e361a319f1a687f73e0eae22899c93feea3c522e42f
zcfc6f447ade89b28ed25367bdb2062850e1319e3deba92f1772dcd2b7522b7a65d97201ca9631f
z5b544bbcd94e365597164cc90dd09ec00c1da4332cd53ba361614c28c6a72090169b3074727047
z1b0593c0375dbcfff56123708519330690de192fefa2af3d9edb38634fc581622807312277df95
z33b40b67e617a9dbc793eeb79124bd266ad89a31d20da62a2a3fcef9208cd5e1ec832bd4b684e4
z59e5d67be7842eacb774c26c986c2c94356e6e2d428261073392e67b6a3d09ef27dbcf8c70ac50
z7fdc630a10fab3b7fc3b51a1bf1dc0193ee7adf47d2cbd1abad30fe04a97db45f4aa34693cb98d
za187341dba65829ee4ccbe8281ba84bd3195d294cdf5a9a731c9f46f8d7fd749000ee02181e03d
z617ce0dd64629e1e70e91536467aca515c53c64c44866cda5e744bd82fab9ca30624916a81dfa8
z2a063d2f70551adbaf91f290f53f9313b774674a969d4d0083e587ae38fa4d559c04115c8fe11f
z39f5cd28532b6622af915327eff41877b215cade64c45e5efdb5f29c11a9309d406f7ab0e3ffee
z4528e5c7e85a14df26eaacdc49732a4c346632d6d5c993bf9c6c81f8479555a3fba42bd37bf5e0
zcac5e8dbc639d22181c04a8de7f52d63e4c98bacd127abadc870bd0fe2cb9b2a3207d85f5504e2
zf2e0dbb2d41db8086623fe083306136d9d7ae742154c5cda8a1fca200172c6d0ec073fd7bab246
z8eb9cb830e02aa6eb92b51a94bc5bec59a8e8c34597075a70fde50c3702371649bf5096431b00b
zb3864e9483feb8e30cd337e10c4e318f88c8ef49c7f712355ca3289a0a34e781254892297100fd
z5fbbe2373415680991d24c6a8ea9b654d1c2c9c862986be4d4b13a8acd0e7e4341d71367493db7
z4bc4bf1f53ea249d286436e9ccc8c6040e8c3a4b63ac51a020041321ca6b49a0ab6d6c97898939
z0f23b246114b53ec5b9bbdefe2ef0eb8fa83b8448a9934a2b018150c57d1c8e8834b5a6a80e4ef
ze01345a037906724587d450ec505ea910a8fd289b39a832c1f9dcb9ba8164181630893e73fa4fb
z681c37bb9e63d4d6ef4f3efa27d1077a19a11faca326932ae656069ebf7d4fcb7445872dec3a1f
z63b308706fc0c199e7250479ccf44d5ecb1616d7f5f7963a7e848560af15abb0cbba37f6c3abb0
z022f12a9a0341cc9cf1a1c599a8f7a980930a916e9ade15411e15a65798da7c2ddacae4684e10e
zffe51d8e92c0fdb451bcb710b2ccbdc0acf1c61a9ec901700ae66e492af9c943e2fc5f60011324
zda611aa64787c16c6bb2885d3581690ed7c33cd2437cedf2b5cdb2db8af0bb68a68f4b50b86e34
zf174fd46bdf4a541fe485678425639b84f7f5766e870da970812ab36680ab022835f223eccd5f5
z13ab5910cd202b8f6b1ded7223615cd716d5ad3009e21fca6d5caed104cba7cc6da5cd0a4be3d0
zc430334b4ad8c283dcb8183e46d69eac9b8eeac9fe6bd19591ddfdd48dd291c58ad9baaf139164
z2a9a77c1c018abda29ec3f685960d8dac2268c2e9cc58987faf14bf40c44f2da90255d294eba89
zba2df3cb73eadf85171f7613bb41b598f6a97c38ee32dd944ecd9df0d05cc048ebadb58b2bf9e5
z5c08b3cc58664ca0db5dcf5bd642088f2ed0fe2ef7d51d9c290ea13fb53530c6f98dc016d5462b
z06cc702d71c9db404916a89bb0c8a2267e8194ef6d6a21f7c8c11bbaf304de920c9abb185690cf
zbfc0750fddf78cc40eb5260107405f9c48c7a8ed15acc4754ec2d87cab2e7e11e6bab9e0715f4e
z6353bc91da1516e41489fc162590703d370a8b1326121fc29566ecd1fc48488a8c50a5f7737675
zd29df57ae000b6a34d46d302a52d67134d3bf76da62f7c9f260f91aef2670794c3887010397bcb
zfe6864e6606c0ac0e5ef24b5c26ee27564317557e6ef86831aa60fd063962801c50e7baa589a1c
zcc9961b84c5318ef000064fa59a2e11cfce1395eaf81f28e543b04a18051936381ff772ceeeb7a
zb6b5fbc5750eb65331a262c42e688b26df88d8da067625f1040f198a74653edf290dcfcb52349b
z47ba9a91e029c8d5bd740bb014fbba5b0de858971231005ee4c69c582c69cdc71e00118e6a4340
zafdd82be698023479d1058bd36b27f97f50b1d60bfffffc58b483018194b98da52a2da19803b9b
zd2c12fc419f341d9a965f4ce585fc4d3054734ab058fca4b63f1399ed31f88ea0bb96a1af3d7c7
zffae657dae6a55acd74103592d9111610cb4cb9999fe83bf840eed0d3500295a5e8872cec339b0
z5b10ed9e1c84cf31dd5a5d24a9a6c522830480df6598ea7491ebd6ff5083390712862f5adf6644
zed9a1bcfdf74eba82ec2fec1305c9b2bbac752f83ae590a4d081ca9daf7c28cf7e26e26680f298
z883b9788c82669a1dedfd9f895a49e3bd7492a2c9b5425dbec4f4f1632cf7f6df93c8dea41e3de
z2fc98e106f0e797cce21cd0dbd5e76d8f6c88857a311da36b412d47c955d9399a55c2068523871
zfeb5a87b9a6534d4084a89877a6f4a3d59e123d5a1d4b71e3f9d0c5e900a45a35d28b7931581fb
z26ed097ef70adce88ea3bda4a3a2934d7cbbf60d40d93d0f9b23081fe20819fc6204a1be9d28b5
z7bbef77b0b1af52afee1b98698a30db2a2a2bb752871e36c4fbca48444adc4b66a97ec6c4b1204
z5bd1e1f09bf82a5989b9beb58efab5060bf74089bc992efc41b3e5cce30ec374e0442b77eb33f7
z1947117854b7406b8c879cd1844a915351c1f2b13e389016299aee85e72b429268cf5f97978653
z05b2d10577bd077781f7f84a39fcd4a228b7a486bcc0c106ab4d424311ac65c01530ada30ce91a
zd13133478a96efff866fab73aab7e330e576170c13bd6e8ed90853b449da53397574e3a56bbd66
z011ac26c8cd818edf7e68734ebb67a4bc4e81e43728c9291baaf60103f4467e86da25bc4dfbea0
zcd7cc6379b9105fbbbbfb189ebf06ad5b29e23298c9236451688783c93653359b3372e525a8cb7
z39a592b2a4b52ab45e848faeada461350bac92534b0aaf954718be12277eaf1212636c31f1bc5c
zfe8349d1ec926916a003716a498e817194a7268879d30d12299551f39e63b76e6c6fadff38cd18
z9a62fc61f09ad1edb2d0d58488dd54218fcc4471acd37752a560029078260aab3e5e8e3313ca26
z132ce1d8919a2b0636a2da4d96b0126428044d525c19eddb30f5fb9f5546063e2718aa11d16102
ze43a04700329e0427f50bb83b45dcc7a1f7d92ee69ed1e581c8cda6ebcb79c0e4b2220453d9664
z714c1533a4bd562c21df091610fa9239ca10855172ef5d07163d55392f5987fa01f000aa66b112
zd4cf4e40b59cdb7ffefba6d6804dd2c6e675fd9a6705d539f6022a567c04937a0dfa562c04ff1d
z947d7fb2f153ac3ac5043d8284de3801e4742ca024ef70eb62ee9250605552456a49a8784eea97
z82c5225ddd49df5de829a0f7939af1f6d917724e85a8a47ece0954c07f9d6d1461d6d97b73b0db
z9e14e65876a19bf52a4de9a96347c885186b112dcf84ae067e38cf1f8f3b394663aed5793f3b7c
z757ec32a879998a548169b785ae751d7973dd12728cdbcc8c87d669ecab2a2bbf9b841ce09e93f
z3177ab51eb992c2e9e0b3904a0e46bc24486d161fb61914440c8c03077ad5107a9b6027d57fed7
z0082019d1eec6de5d8c4ef8e78f40b83f8e2df280a8f28f162886732fd4d1f735b1bb0fa6b9591
z358280a3cf2f82a3790676c07e8bdbe00d7dbb4869e2e8361ede383b5b06e8cd89bb776abb536e
zcd2b417f2ae98e1ce75af6a78fa85cb18a992d9d9d787a96b6a109fc32796765a84c7a8c6eda97
z7b0f3ce8578c1bec929e5e73720e7ef33de01f28ccdb6096ca4776517b786e01d4fba010c2e426
zf5795599cbef6a76145184f5c173d7c88700c60a16df3024b7fb81112108fdddf6388b92ed0e5b
z29e6475ff170be9a13499b9fc9d6305296b091349cc712d85cb3c7ed423919f729e4933114e016
ze830db5ce9b4735a67fe19739121855a2941d04b1d81f18356483a4ee5256196884260a081816f
z8315c0e6363aaf6588b7e2cfa67359f674a2894c27a7d32b8e9ed92ddd99730df2af5e2af880be
z1c9021aef36c3ec66dbb74775a2f95937e5995fb598310e137eb8e290e7b4998962e23e066d26a
za3bc8d95733b168f8535b7b0f456123d67ff1b4b43aa244df6e1504f7d7f04104e7a2cc1468ab5
z644a45eda3dbff95a026b00ec648d9845f0e79de50b68342337529ad473d7af7cfa15928906d67
zcf4c15f56522176fc95ed1d6a120b0adb7b2b417122e233560154f87cf2369bf5b6c2a3a95cd1a
z76fc6acd6adbd181c3758c41d50cacd8f0603e5526f8eb85574a307846f9517e68bbc5763fc100
z5260ce169d0f5de1f15853bc01f289678ff8066ce50197ceee8b700522d4b77a06a0a7683a9657
zbbb7632a7fe0e048e0b257828c794a4f880418007919174b5c02b86f7c2678786fdae805caf647
z86660106797bff87c7a08f6c546f23a4563687cee79a744778f69da5091edee8fe8595bbfc74d2
z466b374994381d456b8a04ea0c0e3a27840ffcdfa86c08351ca2257f6f7998dd281df83704c90e
zec2c47c82664a5d9f7329ffb2d06c057907e0faffd47db16bac08a8e4c8cf1d5c8798e5248ed1d
z615b7e090332a7280d44d8ed8bdf42af4a56d6dadb871bda615f5a662858ac236d9b0217454f49
z5388efc1e7919965f9be0bff4c0f30c127b8959735cae05950c79d071c3bc89b280004c54b8714
z3836edf4309fbc2f0816ff8f64098f99346c5450224b11f369df9ac90aa60bf471dbc8b8e62c96
z6ab9e2798d87dc49e15bc9244824fc88cd0cc10f5c9ae4ea697e638e9fe6196e2ecedc28cebe36
z008b3865d71a4f5e9f1e5800d329a391c6bb4b09442f3597011d36e53c1a974f4d5e48ed8c8928
z0a55ca3df0678fd6404304993c852ae3f8971a2aefdb2df9e1669f05ac2749b046e6fda1097ad6
z2331122068b811e53e23c4c040a3682d9bc3c49a212f79ecc5f56bedaba61501d549da679030ae
z82a4b529a3d351203369118e53d0fb4599a429561876a4fa82fb07b14fbba14a09301fdac38483
ze4c5fe8ead797003213ee02d777b2e981cb2e35980ad4d1f5d6a38114d8e7f12c607d7a37659d7
z243b7bb4a0b707ada36a0ef6ff7ca0627056e0064ad253bce060a9eb5440e3f3f6cab3a15adf93
zb78805087d61b4d42b61391a51cefd57edce2ee9cbbe7f3bc9e2b5eb810ca6401cfaab38dba478
z1bda98f3d9a072882b2f946786261dcc29b29e517c28c9f46700a3b0fcf78b0012d92c1b954452
z82358a41117e65191af162de0a759c17fcac73669091f4ee673a65e8080e27bbbe1403d7a3dcdc
zb822da5b25d97a4b0f48b08e9eec0d5eeae29a8f55ec6ad4edb9320444a337993e144d6cd45509
zeefcbbcbacb40300c94db2bd1e31acf879a03579309bd3aa868a01e6eba7509282d445c21c89b0
zcf556df2dee94b1e2348b9fe8714914b2c89bf09e184dd9a158860605fdceaaa7f6733195f871e
zb7904fbca1c0e128d35ba91c05576df7d66a839749b0ae887b2fa30df8c7541f4a6115e6ffe2ca
z4c666f8e1419c276b2763a5794897e442480487fc896bbf4044e02d2c08c986621d512609a4e36
z75f608e0f524f4e189dc08905d49c29e0377a7a7dee65ca27dac779317dfae7675d4ca050b11d9
z98f7ffdaef738ee3ad97fb0cbbe0ba0d4bc157a5f2b3c499e2aa52e122e8527d71642b5866aaba
zcfaf9602c89685b2d31fc62d031938408e2655702c52347d1b4ea9ee69ba9dc975ce3ed5e02185
z7d30639f1143a8138e8f29b3f8488054fa7c677eeef5bf7384140715d6ce4688557e5b9a077fdb
z4935a52400ba72fe7aec9a3de677a9a6399fb280875667accea14b845c2847a561619b02fd97e5
zca193dbcd37320dc8a1eabfa18580111144e922e177fe3496216f02985da43e0b24de5cd4d1409
zcb3096b12b73c576253f197985b7549e9573e6a9e94862f77a2ce7b649c8608c3d6b383bd82fb6
z8eaa70a9f26da5ff38239fe743ab7801766d313269a632d3a9db0751b867f7180c2a60ecd01728
z8453c839e6b5bc6212a536b4f72c576a51f26a1ea21544c33e25d511a4ab651b8c23dd37803db5
ze795bfa64cfa0504c8309f354f24fa57293c5b2c78fdd7b6c91356e40699c2bd9624113174cc7f
z69dfab837dd5d5706b6ce143a57a82e37cf2fb5175ae0df2f475c21a0fcdfde04eaa7bc2f26d6c
zec4b7cf990d2221d3f4b1ce26819d702522733cfc459133eccaa3588042d25f0b2647e4a7dc2ad
z0e4dc7abb0b53c39d51f2cca6452f9a5af7dd75504cda4b25d41f890fa5f8b86d86728d4bde458
z666b3daeb8b4795680dda225ecbc86eaf160de796e6f4952b49870f37e0d25bbce523ea155454c
ze3c4c981abb958170d32a2839e4e8e7dc4d3e7ed034a158b2f7e4168395c33fe73323f8de9e453
z39ec2f29bdab4470bd37f9f8beb18e9f983374828624e8feeeb396d0dca525a26296705f712cbe
zd4328ff8e4481a9c6214b18acea7800beaf2bceb1903c92d36397c5021100010ff4d25007ccbfc
zd42ac0ed94761e84b318b7591253e830050b9030c6c90e1a267dae2df9be42520bed4fd225df85
z797a3b17af9233bcce84962c5563db31f4fd81c5543620d1c681cda4408a0b8da88daeb9ac13e7
z8678139a8f196716f6e3cd8bd7a60a8b00eb713967499b2288db1241372f200a971ad2615cb1d7
z38924dc1856ddae5f74566762767b9fad8684a7b07748ed1ba7cc831694b44b32aa964c8dfe485
zfc243fe65ddd8513384fae536b43159dc64aee1e004e53b38da0351d6d7e1a9ea9b400dd8fd6d0
z1f928322805b78aa9a4e9f004cc48ba5ab5b295723c87737163874ff4fff6402fe6e9991364108
z5b39c479556a2b78d5a24511f14cf44bee3fc5052759b20098b5c2e9cf2431f09e30e554458c12
z9d12f6954a9983680508dadfe704b2eeeb31544c5f9d92a9003b40ed8b47606ee961167f7c81cb
za11f0e70bec2b26f70869ebe23f21faf093fd1f5fd69ca946f84f4a3e0041bbb26d8ce3cd5d5b7
zb0a7231e8789889fd46efd9e08c96c97ba1fe3ac7218f81fb72b45dff4e88b19f3e8b8473bf802
z91cd9718425151f348c8196a2144bd46d42dfe60dc6b9d4d854a4c8c75c234c429448b64023b6d
ze9619485354a873dc20256eccd3b06fa08d37decc39da1da9a667426161880cb83fc51f9f07e47
zdb840b7d8b02d53cb8f5e2d821110810508074228024ea39a0c1eeea484f03719e876592d0700f
zfd53f4bce1c28d59254c56017a6d35856c0e36f976303c7424be54d7d88ecb2cd6a3b668f9d3f5
zdeca11208ed4a41c27d945b6cb126bef51f25d4368ab66891c89754d6d5496e9db1354172e5d81
z0323720f48c74d712638f77c4e1dafbcd4336fa419ba2bef1460b41a0705ca6b315ba320c39ca2
zc2985e0dd6bec5af38a993e812e3f036709f7e592cbb0ecce641b5dbed02b640f52283bac9e029
zbf200b1c9d9681e78ff96dee1a1e1f3c755d0dc37a8e7aa9263b2844c7061f07d4f24dddc2712e
z9c0067fa6ca4473e7240a9ba10fac9ded8ef7d0264d4e13d7f9353e7913085dd990fc0a1fd916d
z47f3cdf9a411dc22282415534165ffe507430cb8a17763c8a14ef7ee53b9e371950d0f3f746a75
zcd5182c8d7df59c06aadfe7f25c1f4baac1886f7b7bd1907e440c17b901dc25a67e590ee682a63
zf1ae707cbe87bbbc4b0c0d8f18cfe80d2c3b19852d36cd7c918553970d1387e4894491a82b5107
z5d14d9d08cf339243ff82fdb8c79e46eb62db2d760cf977fe7c86f1cbe7fc395f14b008ad3e8da
z89efcb95d076ffc47f38ec79725609348200dd8bc3b50f18ed2098da2cf4695dcbc275c238a154
zf1ba39848e0f3eb680f03896c7398304acf2f75c5167e4e046824e95ac658f2d9e6054dac8bcbc
z2d449e77f058a6355af3baa2ee6e8dd61992baa60ae60331faf4e6e3ec4f4074453bfde9082758
z11c8b7ef78b78fc2299b0ae3558342a4d179a489944d3038d4a4ab0646573ebd4612262b4352f2
z0ecf81dba2abf3320a03d1851e194d3a281c06afc7ae764e0a3c1cc9af8929dee0d05455e4fc05
zf6c4e3fe3e946ab1af61c6e977b3d949ac57831487e41bb6763ed38fe95cf6c6fb08a9fcf3eadc
z2b9171757d281ab5d2c16900566b7b58c467981c3834b8ee31e2070933b63d90732bda5b7c245a
z0120bdb239ab4cdb8134950526b215b95e913ce2e3ccd7d031f944fcf198fa0445307363d79419
z24d6161fd3d04325c16167b8978931e9a5d44569c0da5e47a0d4ad8e344901b7bef2a1540d13a1
z78ca85b38158206b10f2d4c0149ecba832bdbed5652c4901ec3689f11e281fef21b80543b7b7f4
za626737ceb9ec16efa0d2eabef10179aac0ce74177bf5dfcce79767e898339a667fbe886a483d2
z60cb61e5e7212042e3a41a7b12c92081eafd5e87ffe0da73d6eab94d132443942feab15ada0edf
z08195df652a154f408bd12fc9400c3bba6d33ba5f6da57ef7cffa00c156ffa4a3d476bac8ddd11
z3b41108403b147c54ce50037b7abb70928f0ba46ec70f8ecb10cf6f6d2952ce0f893fc11fedd21
z4add9c37043857e2279d5744bd4f07a37ff58dd6ab2147fa8b4fce371ae375744c41e5a0561324
zff0424bdf64072c42a80928e8562086acb7869c51016845b58ed94d319d08ccfb99f6dd7296dec
z5b43950009f92fda90f6887e1bcfea8bb52d16f8df94caa399055c7ba2a71aea23c6c29110ab82
ze62c5ffb66592246f9e905d767abc57075181a58c608cfe06dc39387e6ebe09b42cc8df672fa9b
ze9220ca87e6f2a0cdc03fa0834f16b5d542d79e7eaad1682e2163c4fda3f2e2e25862929b52d4f
z07442ca24e16843003a57386067a610781f2e86854e00d19fd599cda0b1baaf309a82155522a93
z98f31bf97baee572895c198ea9b288861d21144b80042224ea41b3088cf92e8a8d2441f9c5ae4d
zb0d44c39e86b431404d2a9c6773bec49c0775b15e54cee2bba4a5d1ca5e2099d69f0cd52559015
z62722dd0d5a2cdb77c5ddf97e2864cac8c2aecf352a5e2119329fba2d8cab7c32631528b42a379
z3436a3dce1e7e566076f1f78f4e43ee3e2593e1b649ed9fe146defbdcbf72b5496ed49e7923540
z54ad3f369c4397ca26cd0fcdbb1a55823cc0a455d7990324e7574747ed8476fc6a86bf7fb987d1
z93ff0c35855a0529dd52232cb65dc28eb9400321fd2cd18cbe0389da437fa4022c0cd3b36ff2fa
z52fd6ee2c007b7a16b23c96cd1b6e3fa572d18799ecce72713f1136ed7d542056c040871536119
z7cb74924361d5181a41b5a3a6e09388356427b8fbb6bd835ce67b5d24dc585dfae4bf351252572
z74984177902dc21fd7c4df1f496b219fbd04b489ceeb18f5c9ede0eea2755a0940c53821638f28
z0405391c76902bb7e0dd80c3f81c2a33a4a127879744b92e620069a100ae56530842874af9ae24
z9ef523071fca077852bb4d1fb3f811f97c5ee8601cef0af272d9575be3842332954190bcb859aa
zfcc604e60bf51f1584e207e6a3c2f81ba27b25bd491437343701d249cbb1bc13323efff9562d64
z7141cab2501ae0584e16f7cd1c12e93593934ae012fd442abec08b8ccc340ebbb45647abbf703d
z4be1a514bf7b14cca621ce04ac27ba188326f9b85a760c87372d3bfad067f333f496dd322c34d5
z1dc64489af1e1b7bbe982987b6d28ac680819aabc621144849a4c17638a4ec1e3d27ad9826c8fe
zb48d232e79cf3866fd4d404e3adfae12e87639ee7549d29e3f61c09baf1f8097fbc817995f4b73
zc13c735010fac62cba5b105c88d821598762220886045797ef0c0e02ea988a2f0857e392f0b31a
z4d7c2a3526cf38bf1b04e64a1e2ae9d103e608216ec5c8dc6642c83f847471ccd43a1b614f3e25
za208c4b255ef94aa7ba5d1b6f211edb9333220c32613686ba3ea2157cd12f8e40de505a7d88dcb
z2ea45c4680f935049a603e95af37f75138d0c8add98e96a222b95a0965da74284d55cd2656e069
z5518b2b0f4e4ae7883d761923b3762c4bd5314287ad871d0955cef776f443067622c2031267336
ze980dd95c08472f634d66048a448150c9ea66000e7a672a30268e4ca06934cc9fc38ac7fb095fa
z6af9ba5d5c5ed2718363e42406cd473f6f7ac60198b46b655689e845629e01461de36acff99614
z22f81ac58f3b5116e0fc0c2eb27a33addb710cf0f3fabcf4ab9ff507ca9f44b0498824f8d958fc
z47bcd4b44947a509f4891c19b5abc4ebdc6d74b6d33cf33ce3ecbf3175c740b451a1fe1cf185c6
z94045ac12ba4e8551c6c1c4e1a3ff58d0b3cc4e35486e21bf654ae8d00cba168931d7fc96bac90
zba789214509fc42815ac24b68db429f379896ae3195150a74415a97ff5ea1e277eaf06e8c41b5b
z0fac55e20da1d468f7e4a8911c08d895c073a524224e04a4632f40c30f0c0fa7d92aa5bd59054d
zb06a8366b486b866c31654a93418526ff3953696d214aadf7ef15f6a7677d29d35de43ff26e21e
z7f4851732149cf3c7c2b4f484289064a0c10b36527c70e757afb23cc259d9e231c66a270a538d7
zae61e99241756c870203ffd6b22a63d42501b8654ea615933be63926b3564f6c5c643a10611439
z0024d6bd7febe31130d3ab4f96537e51d70da2206f7801958fddca61c06def4a5d3b745522b8f0
zf2946182b589ef3a32028c327506459ebeb18bef726ac334430bb05fe7cb4105847f4bbcab6185
zacc33cc46d4c8b0d4dcd4798ad320bcb44ed9aed95405339dbd8c6a71eaf4ef6d8eec8367c9b31
z8824948a679562c4e3d5c047f6eda1eecce3d3b8458db15a57d63906058b7fa5302e17b2ecfc30
z7b7084fc82e66f73f9409816d151cad655476202eb848a7658cfb65b79c2829afb5ae93e8ecfad
zada70d919c164c2573f6530576b0a2f5ad1755ef7d7c6bafe4b71163371887ee2ffe7d90bf4beb
zee9700e0dfab09ae908ef428aa77ba3a68c8ed3ef4d0234ac3b3d6048cda4788d2393aa64266a0
z96f66a4f5cf670b526bffbdb8aead8e68066a91d081c259087c4bff9232a56cac236fea3e7dde4
zae9e3769b1253fdf473ca46f2cd1e54372640a5d4e378e54de2e6a7c31efbbbefe29b3ee490aea
z671546baa01b931db36e948ef041336e796e697f2228c66a410975d524bc5f0ac8062b45f16f6c
z2b97c5b495a1e20d8063dfd4b35b0c1a252e0b31f3cbfeff20f0bad705c80aeb2584ac8400d56f
z43e62fe0ec7ff70d7188568e4415f0284b68cf3fd259e196fae56cefd018ce9de621b899a045d9
z0fb46f801697fec4b8a2b5801fa24d39c7189de470594adebd5f6c424232e6d68200aa98be9553
zd081400b5185778612d54e645f1f830a9fd8c1191d700c24a7b29185d0b1584fd79eed92e2e6ea
z3cb37b1cd7ea6652a64fd0c2a3a92b1bbbcf089df78b73bb584284d6e2554eab33d8a3c653d564
ze5f73982103df788da2775c4bb29fb618ba097a63c08b23b6fbfb74712788cf0aac6fc58b3462f
z85fdb15e5cbcd7e75c56a7c39a7ecb2b1e4a106a9c8bf01360316d1a4d51da7db716d880d77aaf
z332e0b442adc460d83a2906f118c756d908755d062e31180d6d5809e653ebdefbee992df6cdd4d
ze58ff29e6c49e5b9b5bc11335b7544e9fe537c88d755293b3e1087d28afc98c0f569bf6a4448a6
z64173472d5700c0196a23ab3be3dd6fd2c973bf4414e562db24ae1808a7a9662a079b55321687b
z51953a58bbcc81d72e27718a9d4a8c1cfc628b046d79cfe0b0798f5522ab0d7832b731704744c4
zf7c061b0a999805aa3ec90d22fa960c7ea8b87785e3ca3a2c95829469ccff705a0433d76d66b3d
z66f9a46bfa89f0477267c6fcb02390b466f6d0551a549b566673eb1cf510f06c2bebb66fe070b4
z7fd083fece22dbdd18aafcdf9a025fe5db19d5e9626f308cf90ffac92c50356727df8dd89f4147
z261eebc5c3ce9d33d2a93552a249bb5440b0575d6180c0f3f427cad881ba3f308f5b805d6bc632
zc689010944c951eaeb93092bfe5e408b39e36fa8027d4242342c49de2b835d4d503e8e2217aa4f
zdbb97695ecfc5e8ff20b3fee2b2673978ee0c1fed45295aebf41de08491bdfe69d3ca0c96a9d39
zc6af2fc72e5c584c02b1288074b04b01910b427b00b08e2c273cbc60d41d93c835d378196ee59e
z49a0be34ccb273791bca5e8083dca2133f2cb248e235d3bdf00ef267cf9adf90bf2ad806ce810f
zf96e2aef6eed70037b5e867cb6139c24b7d75a4022f80ffb1e08f278537680ac0dda12bd9f8848
zff5c168aa17c5fc2b9c3c2c5f2e8c4fd62cf5d5f32615acd72a97cb26f6157f8bc5b0d7ae0b9b4
z10a03c8511b9c41fd7a5c55a431fc36f42bbf152213ac86c289dc2573b7695ea452c687f88d525
z8c78adee4b9120b073818b7822d4e1857ea12c2d85d217ed7e9d8a75fa6006068b06e8569997f7
z6ca6700b7a4a3f7463964a72c752c7e915a3b3f5724b2aa4bf8865d6555496172629d58a9e5260
za345f857396f7a399377955e0811d875905c1c7e26b4633dea6d4e63d2a7d77b5ebd91976f4476
z1f92b724f4f703a224fe07bcfc066c72abfd1728b7492d8322cddd9e85d23d83ed05301a6f7709
z9082870883d103c015e2dddb837487546128ba6ff206043885f881887461bf5d231017a1161b7d
z350fa976f15574e8b430bfaefec136f2522bf758e54e235807fea858480b7e17457c51f48238b6
z070eda40ab046e061371172fdf42d73e822ae7fde588dae3d59999a102b65cabb503b8a22bb3b6
z06e79a651b14c7c47944c016fbca1813fdc44d9b8c0bdda4376d6bcd981e027257fe0f66949053
z48e7100cb1c9ce08eaf28df07b2ed44ead2d22a3cb66a1d6198fb0dcf0a0260121e48bdcc76cf1
z7ace20c99075b5c2b90181f0b4035bbff3a2a72ec6038287429ce4b0f9eddf748d83863e6cce86
z1071d9fa72aa81646cafd0547bdbe069a1060c2feb580bb590f5d11dacb78c22a390977d7eab4f
zad4a7776998dd04e8e77b8d63019c4bc5d24789754d97132ff654b1886de7e78aa01ca67616944
z6d4eb3fdf04c98aa08913134501a9d057263aec2bcb0ec9c1f5017e60edadbdb1cfa164a3775b7
z3ea02afad251f3d26b045b113f02bf8884631e4a5711d318c9d6fa307df266c6ff0f8e64c2503c
z1f35ba4ddb7de99fcdefd1602f8cc4ced7655e3299bdea45fec934f4432bdb22958f1cf9244bd7
za2f1b5c06446ef14beb9b4b93e4588f61139b83ac6f3071472c752db0b6c8d879046057846ce32
z90858bc490c79bb9a934f7086905f721061c870bf52cac91eafbc1c022b30006f43687ee255cb2
z16935201a3e994b3906c35a22736c0fc754e70b1f0d1895937205f2a31b03ac2b4e302ff5b455d
za3acce113f4c7f24ab851d871bfbad4cb56f9f82ba0dc0262755fcd6045042159c98869a91e1c8
zbbdb560aedbef6bac0e673aa8de60cdf1e978cc96c10e6ca74a9cf0a41ab7ebc2b5aa556badd71
zeba7be5a94754ddde6a79e5f1e7084a3b942fdb7e976c06eab8a9eccf22ce7bf1ebf0361a604b6
zb52075c6bdada49cdb3a2129b05f350d0c9b6642aee42a031ad0d54cc83c67390132f78b8f1eaf
zb42bfe93a6eb65aa10df6206a4cfdc05abd1b45f65da00fb5c53651362b15f92925680f4cd4f16
z70fffc1b70ea11f36b3aa457c221515ea3a42b8948737e1f6497e5e4de171b73e20f995eedbd42
z5338a110922ed24127329f4521083c7c889da5bec0cd34322dff9030d32203d0d1bda077331680
z03caa683bd9bd0a80bc1ecfc41be243e096a98ff8289f5cf0caa8485b21176bda28143fd33a831
zbbfe780e8fefca173d05c73640e33f84ce03a071fd130642aab99d04271b4e37e74e53c84cd2c2
z7143c0c32745e20c2a3869ae1985414e4702fd59ca26ca6dbe8a68f573d0a521b6aaca7ca9f16b
z50f8f88e74814516e6ac84b490d648908e35ca34f0d76afb6e2244905341b49bba3ad0552d76b4
z9576689dedfc06623ffb2a1a477c74438e34c815af10ddf18c7506a2451368dc17beac61d6f82e
z8cf7e52245865531e1f9b18d60181789c8ee1a0465c480fe7413e99355e425c7d8d3bcbc1e3b6d
z5d0f901c9661b8f253fadb88940f94b4abc5991f205134c154f6eff05512233eee69b353e353e0
zc3b97db7974a94ed2f5e54ad53f63a312b2c4360423db0b511e8a5ddb6e0932967af7ed9a7d844
z1cb73b4e207c7bba9a95fde8cae93af065f896b7ab752876d80f8f137b32a30b0165f13d069fdd
z21a6fade58713f5b2de65238cf20ae15aeb85f64b772dece9f11a8d43d34b7b3dd524867779485
z621c1e1848448475cedf991cb77ac14bee9fb2a1ce5ef060725ef81c50727c1d6e460acdafb4da
z8bb66edbe98fe691c81c58fbe3c7bd7244435141f2c22170255b53d533254f4256fb151c6af22b
zb1971952ae408e9f5a75c75441e735aaebbb63f70ee3a500a6c97d9b1a356c07e21b81a324bd6c
z29d4c63744590d438c32c3b59a0712ff1d1b07f2653773ba7f29f2d1a48feeb841bd571b7f5d58
z0ed8faf4fd6d873044a21c6c8687b9cf4ca85e83a3dab445b64fb328542b321d186acb0a565300
zbc0302142ebbc385d30f8a788ded0e23c11a2b9b3f050fdf8abeb817fe7ca455e01d36946ca039
zae53e74d00e2e14466c69b149e59555c1f7bb0e04014529e753d731aa621a6c1ab6dfc0713ae03
zb6cc3168e693924db2e76066c562b1da0e47807feefb807c3b67be51410dc6a1b332052f0cef19
z92d7e05881bcb5c894b96439ec51bdef8aab66b7aeae4b980025c9cd445c1bbb8c86b7cc7b9599
zbd226deb935ce3aca8ef751ef9810e83f2ab58e8348bf14e1b35d123cbe73a0f7cb60896affe50
z7a12a025088afeb171c191191d841ecb87e027d6b729652fcb945434e36d186850ace541b53793
z8b41bef52ca41d6ba185b2ae50e1c25765b17ba2163278f5dae9d1d722bb8250a5a530c35234d5
z81196c489f05bbd3937432e3be398b21dd027463b8393a08650be8d7905d0648a407b7d5b6d121
zbb60bd960d9c4a312a84a9cfde96e4c5652a26521548d702a97e1899c57d53070a0da91c77ce71
z5f054545a4b7f7b20e236699272a527efe9d7f6918829c716a74af920c482278113d73d2580dbd
z0646ace7142392db7ea77cbe753975cc76a2edbebf336822d2b6f6fc2c61db5ba13748d50b52fc
zc2f959798c5db57c550ada07b1fb8c7af11a17752ca24b093a46c95a3e483ef4670ef54942e972
z8071d2d6e2cbc02510d207d86b08d4e07619dc12e4d63196c6bec3fbe12d6a27d6ac23e011f101
z9f8a4ae94097a742288c2c372bdb06d13103d73d1b3d58094474d2793ffb96a682666261df5370
zb4722da610ac98fcdbbc35ebe17a737cb2cb457e61b9dc23c7e584ab7c0187f5eeec9a26040357
zd42161148766b870905a0131668e545e574d54c201bb6588de078ea657fa6f5f656fe148b2d9c9
zd8033b29518665c6016b6166fe8e48688a5793a4c15e5e1c5a16292a0f0d018af1c5dc7e866f35
zd716e75ad321fe7e9337d59619605d4534bd4f35f8062b72521a22a418e1cadae7b597030added
zad5f4f1fc7aa82ffbf4e594bfc828e90b1fae565ef832a55f3faf0f8f4cabca0d7782b7b11da5c
z82d9228c829c6bbb4419d3ab6df817c767d31e82b681e7de4e7b9ff95f75de1b02f7dc6d0e0515
zd0d97bce434c75fd56e5fe2875fe718d3d09e79582282e97a155ce366e85690d1b13ebe424cd12
zee038850e0849deae2223d3d3398fe3da27760ba350a4a5a5a05850619c587b9a209f368dfe114
zb2b0c4ec0ab192e95efdbb2c0834047561c1aa1b1f200bab2eace6c43695606f9784551fe8d095
z2b3ae584d5f5620ad9f22b47f55b47ac792c76d0ffa6517e4a7381d872e75155a87d9f09ebbbec
zb3bd5245f0a13ffeff47711151bb88ea01c0b55361cbde5efb64261a215637efd65656e256a2a5
z9e986b04f7dbb4e178e42302fe67e0de2d323a22e52b0320f0569b622bb6b86fb9f77ac24a8920
z416253e44232493122682eb2e03eb4196f4f5d5fb6838db7e6a21b460784660f667f0ee5b891e1
zbf654530fa0c35ce3089022d9b10123b7386006d45842da6f7521ad459adcc63a17d9ea7e45463
ze7d0439418d46e9277305091d25401ab666b55785adfb7b2de1bda27ba0747b2b23a69434bb654
z60a8903e8ef73f1e74eef816f7c567fd4df84647f9f1f1f57dd2ed157a68c2adafcf365da2bfb6
z65e7df9b85b36b1b491ddf79cab61146040cff9a8762f87e7c190b4dce6dad29453e7f70f8f730
z89b646420569b24f24ea12ba1057653afaae4a469f501e4e578ab93331bf64f7b943cbf0179c35
z162dabf43c3f4447d29cbff3c752052fe58b28754337bfe506d817c22d6808f01cc16f714547e7
zed6be870eebc3a951b2a4940218917e3c817c0c6ad5547e5e9dcb15c29d7770a26e1132963bac0
z2036545c78415002e4d43c3c0de9ce1ec021b875c9a602785420081ba813d63cb3441e9bd3db88
zd88350d183a82698fcf91ee5bbf004e048ebd2a1e494e10433cf7b8d08229f6fb1fe55376ad67f
z12d034ea999b1daaa09719519b40ce36c45532e327e9faa325b233a1106b68ec76280475941704
z6d36682b6faaababa59f2b718c1381c7ba9b17d78657b63a65605ca9ea4199700372c20909fecd
z7ca4a27fb74142a18a9608b27df81fe1e2058e9b06adb1c84f166b51de0ec79d305f4e7c92b701
z6ea9762cba9c74b876bcf683e9cc64f33100156bcea7ad162663a1e322d209b39d71ebc70ce880
zc08d90b75cb57d8318b52e4615941e702f503c021091f8abc5a6db76978ed68f2a2cd2aec3f654
z0289654c336aa4b9a511965c4926af89b0a1f182d621d1e3ca794b7a2c745a82c3a93856ff5f51
z017f2361a4a55ccd9150fc7d52a420038da28a1adbb5648c2e5a494b6247850199bf936840125d
zeaa766a94172bcc98e8ff92c7c3425eb11297c62939f63222bd3efdcff0a8df33f18bdd8da0185
zfc2fa93ff93eeeb66a757cbad5e9b4f88e3d62cddbf710778a646e987869e4d04395c50a6b0bde
z36c22f6f3ad4373037922f9b5cf30b6ed5a6e1f22f1a6eeaa96a6ef29f92fffe466403041c8825
zb92f762e91677032557a81d8d9d8a2471cc7ccca253d81ef8dda8f57428433c62da349915c2697
z2cfbf01a0714e5f58ae5c62f5066015156af94f16e466639ff77661e4390c360a8a6e0a441e492
z05d30eba8e52387a57d8724e866287147563e854134639b340829c0ae679f71b5729d2bbb9317e
z17265b78150ced003161ec715987f8c7a5b273cf88355f42a63c3e2956deb7e868af154a14b6b4
ze510dc74d6a1970c9255e6c51edb3d498021aa7b6c89d0054287b987609310b16add1da80b6de9
z33b58b2ddeaa5e0506b5f771ad7596a1d763cb258c5985c81a1685f13c18b0716518f649586dbb
zbbaee98eedecfbe615ac93958e9c9a96985858e51c37206137dffe2b210af3cdfdf32ba5f91ce5
z781dfb8621a496a72fc08cfdad9b408782787987ef8c4698b2045ef4ee825839dfe72ed92265cf
z3289a55b3b29aaae28c0cdfcad47145f719940ab8ea56eed5de8019a0391fdf5fa8be85103921d
z5f6b05583564702a82fbf7481d2a9881707adca353113673d95faeb3d96cb86a96279191bd68d3
z7b5391333a0bf8a7afd9a2979a88526260995fd0afdf2853d2bca434124eb8bb409c3bc13a853a
zadc66210df5d7bcfbbaf572e777348c20f1b43b8e2b04283e2ca8ae89ca369b909b39c46a267b3
z3cf751eaf1e336901c115d4f9da7c6ff304a216a6fbc9ca507a8b193502700e08b1f882dad699f
z26ef498a7feaab1bb03a551e1a89fc505331f9ee9e54bce28eadcdfc940b85a75d26e9d35bf552
zab86471906aff9699d41b78466b3c0aa2cec9e25ce14ce43157e2e2629b241a05d3ccfbd43e6c6
z010ff38207f3d446a4b867c590f5ef777ca82b637846a58597b72f9c3827cd35273f7540e4f59a
zea0c53c21fbb6f8d7dd55a97c4f1bf008f18e95e47d4c3e060c68405239aaa5db727e094acf789
zf2cd2509fb9591a755a5231da3f727ca096ac3acb0d51f3ee5a21dffb0457d4d49a5a80f96de81
z848b7a7e393d6224e4c818bd422162379813aecb86c11ef1dcf6929a7b1efc3bc50f674486ce90
z09c7a7da13cf291e1e170fb6c9f63d28ac8574d5c48dac463e043b394df0f408407eb3dbdc8bc4
z6361c09ebfe19325009f2878e59e6422c6deacdee28daab76e9d0fd26c9c50ec4e82cd1138f68a
zcd9001b59882c2827b4f881e30ec5c741123f97c713640a13db48e31187b87b5eea97536e7fb01
z08aeb878db621b8abd1857789c80fa4f7071fbca0711fd8eb7c3a9559cc07de40973a0ffddd03b
z15ce8e26d092851bef4f25040ad417c9722a84f4b452af7bd6a13ab8baadfb73e93695a3939f14
zfc8291f8fd03a789fbfca9589a61ca12133ce367120aad52a37b548c782e9d412091bfe7503a74
z094579db6904aba84ca405cb245d08bd0cafec515bf1605e378b7ef977aefea6851c0b81188c14
z4b85224d886f70538fffd7763069311864896ba649d63107799ebae2478ab475d4bb14504c0c23
zb8fa308670308a95ef134f79458915ac1118384faf57801d1e0556658553499348512d7e738339
z79ba440b17c0076e1774ef61c6540f192338eb7858b6467715c268fd32becf1c96d41c898cd718
z9c85ced9ac2a4cd672a68672353b54057cee804dbeb61c9c336396e72add8c546b665ce9b87ea7
z461e3b03941842033006742adb17a13f155156dc01c39216c5b5de9bdca51587ea33ab5354f03b
z26bc0b0330749642c6e370dc41fd9f13d83a94df3393f366a03b224ac6ccc61308a4e3e7441dd3
z2f4323c16c45b2e25eafe3e4cd2d2e747af20ffadd382daa6d8f4afe632050b4608b878a2a8365
z11a607e5b224bc8d5490103ab9d0d3f2971e10f8cb991600a08c952ab5a7a5aa7a7086cd09d29c
z20f523d38571fd9f02f169c8b9568226002804dff9e7900742a1ef2c6eb49f2a160aa629d793fe
z09473a69528b8841d920c309ad2ea9f281695c5c04c366a0e46a3666b81cae6f12835913521021
z435637a7678f86f19217b910189cdf2524b3ed7a2816ed18b138e81ce1b7a0fd762b9f20d2965b
zbee26ca0cc77f722847b067aaf573b891b134846f8ffb462aa8ae126e261d0c7d763ea068c88f8
z59e2172b6a5a79c91c0da868b04c4faf7b756a8fbda310b20d2f2b7a7f3b97f6ccb5135d39b40b
z830a0e0579c7b0a1fa8e5b0b08906721a7bb82b7be4402024b61b755cc41b96864c142d0431a91
zaf6e1f728666014f9320c764d569edb29daf0941894a63e6384bd91bf75fbb77387ea0c516955c
z6ad3aab79caba403192e84a4d98322e2467626a1feb5400e8ff93945158d0f7ec51da58f98029f
z014fca7b9160f4a0117c6aa312efba6fa79813d8f1bfc56fe2a7c0582a54eb1e04f9cc54ff65c9
zea9a74e97a4169dd8a0ed9bdb54052187c18d16a542c2c4f0837515de84ca5c20026031a3d3eb0
z64e8edd0bbdff27e1195d05a03364319345eb462f3bedde3a8c9ab53c0c78d7b792440e8b63130
z71b275c90bed9ed905884082be4deb23e5b55696c492d7d6c172d43afe9343384a1f60b230f231
zf4aed514df9df36ebc28fab509d8e6e62ca7c88beab653ccb63067cea6591cfc4010ba8e771047
z83a176c7f5273025bc71928393be9b9e3fcf639db71d7bc7a78f477c1142d3c498a3e55ffdbcea
z22a9d68201b993cd4494e1ddaf87d67775f99fe545d80f9afbab353ff40c1ee14524e58b773656
zee73d3e6c9bab9db6cbae6df84e9a8d21c9a622221cd88b730b8e04661f4fd55e0fe7236203550
z5fde347531bb98e7523811dae2515e18d94733fd5cca38b0c7b6e95d31fb5105dff37f7f014b01
zd8b5929bc844d238b8e0e6eb53b7df5a65f8d4c9090a1ca38882fc0d4ce4278c55de1677f58c32
zcdcea3b32b17491cab8c3c5a25200fb124753465a82cbce58bf8d2bb87bb8e5407ad3a533b9779
z0c9aff2961cb25f19d7227f5568f04c7ef9d504321b5d31c97e1eb4996126573e532c565db7845
zd6de0d6f530a4b42d3c124c2bf769d627e154ffdbc77a5e907ce3e01a02fb3c2f5ba4dc2e37655
z99863484b5f052772a2c5a4153b8741bcb642f073eb598a1530ddef2062293f0fae6611f9967f8
z6776862ffd8063e0dd0b3dcff3ec789a053621ba1e6e22199fac3cad1ecf6cafce6f67115d38a5
z4dba2d8808d744e9ca605257901a906cc0d58696d26ef42101013c456568dc20e6c13323faf97e
zd37b6a8d5efa22037314cc097b1766557c205be3e688f3d3825a095f7a1fa5b7cccdade9fcd498
ze48556d5e2ea4d1760e9dd6715994a508a0c52a06b37c38c76716eef32abe8fc973e486fbf714e
z8122db6e7cd2991598118467a55092e1d6698f9f206ec09716ab161c8a5a907f13ee7f0391d2b2
z4f7339aefa2962ab3dfd616dc9590fc599f679c21942a8fb2b6374a29eacc1cd9f573aa85399e0
z17fab78cba82b3fc1a73c1f089ea5284a202d0ec41b67da88112da8d25f38a702469e543db58db
z1a6b39d532e42a658ff5fefd24fcc92aa9a872dd7327166a7edc1443a281b36821d44230ccdc08
z3325972df3c7f47c9cf39941968d6cb3fe3abfc37c506f49df81812be8c3a309a2923f9dc6d287
z359853ab8704372230610b39ba100f87b97e1c161e32a889884dab2d3b3747a6793112c1dbb4a6
z827ce140faac003173ea64ee9dd55c13602378865bb57ab05bdd46dd2688b8ce43dee11b840088
z2873ff84e8f6036ff38709c445d1970db33abe2dc0c40febf513de780338a922672ea8d4d290bd
zdf48be60efff8eb7a2ac250612ac955357a5e95bf013af2ed90e8d3690c72842238a512b54ff5b
z06a1cc0eef4b662c3b072dd3feb1a659d139178dda88bc00301903d7f7d8cc9412670c50f74024
ze98e84c2b2b90f6100a749c0001b12b40d4c1a15e284341bfedbc0c001a389d25815d0d8f9c1d8
ze2c93f6f52ae5dd23a0b0524346013f1defbfacc78bd6f3d0585f2087ea839cdf181c9055e675f
z395fa6832731b778d13ab30ac6001b9d8dba25a03b7a45c87a383b58400b63a5a6ee2dfdadf9bb
z674ac960821a1515fb1fed08be740feaa7dce7e8bb74adc0dddc45b041ac759b5fc0e9600113b2
zc13b5a42f870819a8322660f923be5e9e56004cae355d44d12221d06b0eaf83c723c0ae40f1c89
za93d4ea4499a9d4f3df8288e16deac2ef1f41d9b7dd65375b2553d7e49e09f08b03f7f92f735a1
z8cd9195aa2e49c937e7de765325fbb505a6bf42ce04de2da87f46cd6c8f81e0120739e0bf1d457
zaafa6c51caca9270c37712f8f4b5e497a0ccd8f8de510671446fcaf51825a7f989bd2949181e33
z3a7a7e137d0462a4386794b103b217ad8673d984314359511128e497d06868a0709aa2200c3439
z159127b9200cd8c914ac5fefe3b62629798f443f56edb3f1abfec53a91f8618c86fba1235564d4
zdbd4e59060f328e42fac3ea5543e3ef21427f25df0f511c0ef603b4c1a0da1d58945ab3c5f9f37
z0b5885cc0db8d24938dee9c85928575320b1d7d2da69ea27d7715db15063cc0dde5bc67da654d7
zbde3804af2ad6a1476f572409b27f57e0960456af8df890ffe00638d2ba2f042d17f94656c09d8
zd8254b96f82c6a47332ef11459463786829b1e446b85b5f19a894d3fe3ccac46909d1bed32ce0a
z1cd2bd08432603ffc4ab70a21ca2e34912739bd07b3f1d69596274e6930b00db88cfd3e602196f
z95f1f4ee538c3b8679061a248346844761fee47102c94cafa970d7bd6b96eedb83dd5566841360
z870fdf346e68320ab42a84f4f87a8aeb1d5a6d7de8e3b81a9d6237a4ca9df8a591aa67f5b1a9be
z9dfba8ed7759dd61e0329f29ce85badce5f4590c6f4d20f769e2742b20be42e2fb10667104f02e
z17b87d5e25586f2ccbf284d58061b7504c7728874d0148b14fb832249716cb03e0df7a6d068e00
z455086ab2fc47998c79c062647febb22697e156dd07a60d9c1f27b5b08728b97458687d2ee0216
z5b7196222e0008242f2316ea10e12166cfa94def7df3661de582f21f53b9bb531ade746dd59897
z33ed732c6e04d1c3efebd681acb107b4a1409ed55635dbc01bc4b6fed555d3e4b2f2ed377959a5
zc3f0e04cfa02fbe4209557ef80b0c873d955b8b47613c03b3891db4b66fb5cf99e1067db9d388b
z7c5300724717605a31e152ec63d648d991d865446bcfaa1034487422ef668b3e3ef37fce6bbe2b
z52b89558e7a383af10f385a9b988beea6257eb24556f2fba7a2425ad0043cadfbc0b25fa8aba8b
z2c717d908e489a73d3822892a1c464a94fb48ed1460dcf83b58902163b19bd5543caa377487e46
ze70de495dc59821fc6ad4dee35612a74db41358f9e1ad960e83ceed05d1f64fc6acd6e3c98abc4
z7a3ee8fed17c0686483e15dfbc89f5cd3200a6d495e75c5dfadafb8032bbaf2e7eb8a363097982
z0daec4d33da187963b4c52cbf2bbcd4dfc81abdf4e788945e42513bd15522048a848b1a8b3ef76
z3abb219e73653a8ef37ae4c10420df43699b0f660ea938be42f003772c16f28d529c887d83c52e
z12c295f950f1878e23becac8d466f696dd68a3c803e1e9268712e321ef66502fe9c8c6229c253d
z857e8af8ce4a1571ef40086b021c00be2b76a824de3e78f8997ed51dc26de7070018a949c88933
z6bc1c0e10f2c158a52cbb76c8028aff634c3947134d87aba892cf5b6bb6065b5c3cab8afd803fb
zb42777eb9ab0428c4991b084127b686d55a76bfc9e44c5005d89f19ebaaff4d7ed76b86e10613f
zd789b4f9e27531649e5d969ac9f4d83fd123ad0eb308a112273e113be6814f1ef41988ee5783ea
z44d514989f43dceddb63043a239253f71cfee90ffb4c247de3fd78b8adc727628720e0353ec065
z6db24243cd50fcd08443cadc4e75212522974c03b679e4190439c39e0fd9f7aeba972ad79f67e0
z49ed0b0a8ea460523daf10889d961575be3c8ce69ac410264ae486a17afa979c1168a890557942
z0b3982ed187418e2dfd78fec23069ef8b1ff979b070f59961eae9baca28dd9c40691f066471bcb
z7b1953eeb9ada2612fb6cd724b167acbe8de1453b444d2934a8d79e3e8c1619e17c9410c072e13
z8833a5a7e9f3060e6e0d21a21555895e5c15d2d7a5f392d98553fbbf2aa2301664087f0b8e4783
z21f28e3a2a7a50f29e3472c4a15e2d7df6fbdadf719995a55f6ed7d162b18fe54d56df784c3f93
zbe37bd85fa3ed505f1da3c5a1d2264646c015afe91fb1de83338f8d4cee26dbede90a0e583c64d
za56b50c2ff3dfa1524d6add4fb510f29d6e8513533c281c5209ee0d36b2f2304aa2862192555af
z23ce24b96d50071944e4350bb819e9f6364251117c6f6995ceb8ea3197a5c9f280493df983f54e
z6d9197d1baf3f1ddaf4c1d92cf414053c3a09530933ae0be116da9b8c86deeaeb9f266055d976b
zccd9e12597dd6c4dc23d146358b8a7740437d676a1e14fe413374cd39d52eaafe606d47d9e2a00
z24368eb8a799a7878c63c5873d136f193c8a924b99eb00da8dba63ffbd824489d10c92bcb6ef57
z7ddb3aa2ae720cc2f81f36dc4411beef58610ffcc964b403df7f3b8ee1f68dc9d6b5e22a5f164f
zc4f455b42fbf4b94c8f14cfadf64611135f7a3e53630544360a9071aaaf75342dc660efda4438c
zda15d7a25150a3874ea73b0a92f8cf5ac88c50847fec7839a59eceb94ce5ca8e3560d62c3c1a8a
za27037a6add74456880f6eeb32942f8ddbbe5ada80f22ba802d60114f680127b102e1552a942cd
zf1b501e54fa8b01688b2e271bb00ccb5145894d1d6e533c4df4dde497556d2d3569d40510de592
z2ca5c16056def7f369c3d3df9405e4f7353255e092baa33af342c653f981ca8b902de4283149bc
zc0de1bdcdf04d11bf3d817d368d36022c88a2ac63649e99b7b31c5a276c2e3eaa24f015c6d3cb4
z0d05c7c97af70f5ae155a3d7d40a028c9ad7335f987a4ff1e2f6d32a253da4eb282193615e5d05
z4c0f7de43387dcbd776988d468f85e00e03172afc0abbd9cbb0878a1828f20dd56911832e20ed6
z231ea84b25bb326f46e5af25aaa35afef07a7b13f4f54e9f07396855f1235d51bbcf1f14caff21
z8459f5303b51d6f97e9754edbb2a3b2adb5502bd7366889a1a73a74a1a734a9aa8c02983dbc942
zb99978b3b53311bd479bfe8bebd3d5154df887ffac2326b8aa2029db194927bf9f1c86ce88e480
z6102ccdb95d731e91701a181bac89f9b7c76d7a8e3243adca449a59ae123dbbd21fb10697abe23
z396d336eb7f8bd9b6d82d0c54059cdb3620271191ef59ffde629ca4ebc713e20af24d5d6ed891a
z1351906dcb77fbc1775b22442e046d3ac24ccd482937514b27120567b0bdc30569e274183df8ad
z76b1f28f4c7ef738e88d8ac22e5c336e9e085aaf1569bab5c6976ae23bf7cd4616966ac2dc0f0d
z7547ba563843a1ec6de5c83bea2ea1e7d633843a584c2d78b3304db063e77a5055aab990d6627e
z35914e3ae3449d291174bd7f9c1137d80d4075b55f0d4e8e31fde9c7b24eb65ad6e37571461347
z3e32832edea94ab3bfa755ef334010c7f5c71d686015898b04655d3955ac4f7b6146207a769dc8
z6df8c197496651288459b76212e521429c3277dd3e83403d54941666205ea1181b336338160f50
zdd9324e1e2d04ab7eb775aace47cfc66a441582083886e69dfb70a6ea143a9efe2c8d2a118b78b
z668e2b835a404537fbb11a9a147c9d77e285ba433ca9832bf33a5f57d4f090b479dfff98be08f0
z1d7e1765a9ac81edbdf74accf7f5f11f19fae48cf15d3f89de1c46f5725c76457c492589b6c697
z959ac3bbf3a8b3ba2cb8b6c82a6fabd03690b9df743fb9f011deea544684891a5ac98f4d4fe0dd
zcc703b884624cfd134efe820d69ea47ce1ddaace377db5a50d84b64d22e1a3b51d5dd494d44365
zea2cedd3f53eebc7b92054d9ac491a602c85e0ec7e3ba7edeba8ce7add1621e4b07d753ed047be
z53a001fa675289bfb495e316491206b32ffae7e5dbc607772c69c90dee26d735c303808fc5f46c
z04ec514472972a60787c3392770e03f284a94589ed73571010e64fddcdb9497e473ec2153742fe
zb46ee4f538abd7e1c26f7d32ea1204784ee993d48d1601b423ec3eeb851273f0b775b2ab3bddba
z1e88c94315ce59ff5d27a14f43a96d402093d75a82a3afe95a7becc89af747f455181778844158
zd1a666ab217d880c89440ef4b5550eb0c2b41c35aac8ef242d144caec93c2fa3d84717b39d175e
z5ddb437c0bc15591287d1e7ab56d4969eecb6debfa33709618af28a4fb57264931d9b754122b65
z05b92568b8546c452799f682764241e947dfd0ced3878d5048712229bb78d006bcd0aed1ab894c
z4b6664075d888df7e64e4c705c12c50b6754fe59fe13ba25d69bc21acc81622060bf74a41c9a08
z6ea38db7453b225b9175039537b495e7b77ac2649b6d80fcbb7e4de5ebfc9e1926220da37dedc0
z0bcfdbcbff9e0bd9c309dad27d4586b01fbaaff874390005a0fd2629d92595b9776ad77d7baaf3
z10eace62ce1bdef0f618d54aa3466990c377a71b5cd71ed7f3d57b3e075c2e7975595f49d31f10
zc22d1f3c2e218c40e5cdf9bb1284712cd8643768e583d3403202211ca839905a05d12d4bf3d249
zcd9e0a2e9b80ddfd015e4be0efdbf7685c6c28160bca18ce95cc970289dadc7b75615ede0b9979
zfa522506cd7c198acfbc1c9aff034e8dbaa7bff392aebc2d486d6c2bd36452190cfbd7ebf6b684
z648d0d880c486a96af76670494e36894a3da700459cc6eee9e7d1e55a8f5e8629d7f02003f5d8b
z60864174d181bfaafcd3a316527f490ffbd1303f20d0eb3a5ac5f47bb60dbb7a4001c28accb1b0
z033fa4a19fd271b822ccb601521b32962d27db7c086df6481604f2a6d2305e7b4b5a5dfb8bfad5
zf2587b8ab628ade2afa5869be363c79d5c9a6795160eacdab32bd156f33fdda9a330180faf2f04
zabdc55351f98e70c85ecdc4d7e6ab81c3b69053d3f4b319bade51e3cda8653e234ed5e77ee4633
z7f8aa43bbf04a10c62aa7e4978e68a399b8f96e4df47e11a384511d1bb2b5ead3d92004dfd472f
zfc45a28be69fa00e65a93e5e94fd07483dc68ebf08ae508593f766d24fa9bb03c1e232e3b6fb4e
ze68085de3755807304e70eb9b5a09a053750daa9baa1fe85c98bbb3b38c9f746d894f6816befda
z3d3c21f999570e53ec64326e28bfe89794e558692918578817bb11902535563a20bb1b1b2593bd
za86ee4ee2c5c4720f0f38fef3d140d2ac8b37f0e4d4c2e344ee6eb4e253476d8e1a42aa56c3658
zb2dd6d7413461538b99f59e421630d2b01154197974727c465e92a1163212a280fe4611f060f6d
z7c38f708de80c0d4df09c664722b3621865d974d673e779250c132dbc7d9301d12f74c0490159d
zaf9a9e03bc804af76381ac2535c0b2d6685a34a5ebc2a812ac9cfe1d00e69b4f9f5965bcb4c574
z8c7a67c873172ce5da3d95dc9c403742fdd73747da6266e8914f35ea414f0ed592e36613ed4a86
zf2e6d2bfacd661b0365c5c323966b3999f641b3ee446fc9d3ca97ff8a9eff1509a2873c1e5114c
z6ad4f485478800f1d85c60fd536941d1f2c861012510ddbd9cb5cab64bc139c07ec599269528a3
z31d2d1106cbd23507092096bb148cec651765d1811f7eea72bda400aff25ec019a5983d93b8ab0
z14934bc65046c0a9f8d0f5c8c0fb2af44d7eb93a4f1f4eb8b34e9ec5ab249de2129b74fe4601fb
zfbeebc267a7d880ac8705727700373da11c914303da72ca34558eaaf6913b29fbbcb3afaeb4edb
zf2e2944be07106cdb817a0f15ed0c0d3ada0183b3239688cd9e09ef8d33c7e785fd2ac37a730dd
z96b42659a2293b651824555ad742256594c1dbbe5367ebb4c8171cd3bf95a369fc6fd9d6b3632b
z30c56e8da63c33f67a3853abaf409629a81fd046955a569c4cf5a57f27e843690c5c4d1f5ddf10
z043feb614dda7d35238e4d4c88c35795d7dac73b1b45402bdaf0248dec4fb38cecc199d2f3df6d
z05c61308b91b6b4c50436c568406979d4569c0162c547ad0341f175bf8a297ab5934e5f8577bc8
z731c01c591ff2a09b9481ba7005aab6913bac0e88e142f14134d43ec64483fe0283df91d75a718
z45dc3abe9b2f94846ae6be98983f5b9bdaef68c99abfbb08a98d2dd7ac9dcf16a2bdfb04c62195
z3c4f189291913a994a004327b304a4b1dde8714ec9bfe5786cb9639bd3de7214971c3d516e48e5
z0a47f87e0e6aae5be64ab8f07a0b5430f66f61a7595b252e7072cd675d87577f75659523a250ad
zb4b4023f1474a4de84a04b091a64d88c81eba678fcdb6409c6d759121b08c7c319882f4c136234
zacf3b4efb63c77
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_sas_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
