`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab30857016fc53a
za25afc8341302f0c829d94450c399b8ff9b0386c187cb854ee330605b7b59da379b1f26f488e1d
z36e675f0b1336408b3a1ad87d0723054f952fbefc8d5a33eaca6ef5be8f42bc59870a29a5cc9dd
z4fec09ce6e44cac279651402e7e1f590df88ce49ec26ab39f12b4a02855703c6f03b1e85c797d7
za357087d98e5b1f45502e45892e5823d6fa4b762932009620038c05d74efcea7c3fdb38901d620
z36515d0824367e48d1bc182335f158c262d396cada6b0ad58add4f945eee634c2dceadbfb5118e
z14969c29a743830a07124bfa78707f3952b96b0db7af7c9ff36f77137d8c490c4f79328328069e
zd7d5280e4f95742c9841340368b9764f0f80413adb175ecfbdf3c40716abca7b8cef6f7fe92ab9
z6bd2453f1aef7f7899c5365c5c83793cacc7795c269413f6cf0dabad14d40e9285afde8c01a47e
zb61893788ec5060288cabde8fb553f21b02eac61ab0b48ad3d54f4d1d76508b22f0c600861b5ce
zcb30ba708be817b1f50f59c0f6fce449203e7355c1be55b662fef3f92ba58243d81537761af8d6
ze27d7864d2dae99372b2b75bacdc0437a4f7e011d68c3487a89759e3625548fcc920ad06471ee7
z2d701aabf726859343208b0a543c73eeff8406febf277e3babff437ec820fb49d6b78e73bc2353
z884917487d35a6cd06d7d73ccff5f05355122888b886d1b7ae29679db6c9d2d7f218ac9728369e
z0ba3297b105b1781345d5dadc1077db50a0833d4730649f7637b2138ee147e44110be94d8a1fcd
z556e6119eef917699f779ed0e94abd74240fc4193974bfa70d60cffbc620c55278c9e1e14e5101
z31e4184911f1dd9ba3e96b7e8c03693e4ca780a30a1980561a5e6ff97b136902ca7e3f829ee4bb
z59e124fe00f67dcb066f614537b5610816b86d91593518c97555301f13cdbde2409249a9dce892
z43c9001a08d078bd75e7a6b677dcbb261cb1980a517f5000a478fd3dd8b61e5519432dbb53cd07
zc003c318e8669039e65c4240fb4025182b71043f55233245f67482d8a6ec31210efad20b11cac2
z07ccac77b3c573c8546151ba7b181277e90eebb747ab0458760014cf6031a3cfb40fcfe82a54fd
z803dd7485fb0febc6460bc5a210feb71f13e99dca62bd922d9ea809a69d119a1c4fafe35bab7d3
z9c91742229ff8f6c0ccbc71ff838632d297ecc5cdb220b1e13a74d861b247cba264018bfe501b9
zc05d911bb16c248ac7eda4a6adbe926c807c17395092a68e0749f0868be60912956cae8f915e2a
z9017c06a829acc9c29e5df3123380dc2e952e3bb90a0a1079b777dbda523b08d3fc6a371414895
z591d22f472ada1e263db1e5ac76cd003a8fcd32f58bb915b77fc1e99d47a49a2faa767de22b047
z887b4597262d6d21bd9e23354a9cb6ba826bc06d8b3cd9f610ac01a1f3733935ce4ed03a2866c9
z38821d19608be5f8dc8243b0b05ac678e46b3f8f55d324629e6da80179952fea4998639d37ab8a
z3862ce6e79029d7669a6a02797e72d597eb97d500c28916a3878cdd2b960010d53767fd7736008
z984ffac4eeedae5bf73d1cd53b9e33f46cfe12868846962a1cc1e5cae49b923c816969cde60002
z95dfe88ae58fdfaa1472cc1dd0ae99b50e8419bc80e859ee7c1ed6329add5bb13e953fb810f370
z12bb81fd2fb50f22ae70d80aaa687fa51068c9a9de687014959a99c5036aedaf311272b49c3711
z05a18d8d811a3a18622b323a643f723fc828e68a7eda1669def04b021a7927f8822f11272d3cda
z1314104a2cc83b00cd22cc49bca897515cfe10b208d333f69f4dfb569360c00a8b2eebb524cb64
zfb31499dfc80081b2f063e6100052c2475469d917b671993a5a54d67a447092a1aed6e6781ddfb
z9b4d232fe8afc3b838f70d370165539971497d865d82e071974910bbba0ad5ea1755ba3cff26a7
z4b9a3917908750ba31227e106b080e3f3f3a4ff2ad2159d3fa80ccb6f622ef16d28e1a8ced3a62
z796e89a333875f964f18452ad95175ef52833e76ee5b0612dfa40286fae7fc243b8c0457f8026a
z7f8b4cc17a704ae041030d1787ef7a5ca8557f8cfdcb34941df8269225522bab74eb357861a43b
z7b934bde62731667e90c1df7247f4e987e495cb96e06ba17d84ef445473e72b8f58ac4b55fce13
z544142eb7e0918a41e5f097979422b2d12850e20810afa2efe890711f814498447219aa467a66a
z9005458e2237d089c32ef42089aa1a946eb256668304245296376769ff5d7202e206f7e7a871a5
z0a77dde62fcf249eb91847ba170cb351f11f97b81085940d9b3152a62611b9176569acce21ee92
z98febcd18a06d08237d20e7299d61bbfa6cd48c1f0164bd3b23d6719e67cd77674099520bad7df
z52f17fc4a0f77c2cc633066cf709c5dd0fb5cb94cf46d7f30c12190750dfc0235cdc602424bad3
ze925f006cb93a17a0a9506183f5c87cdf21409d741b159691a7569e800a17b884f298603c9d527
ze6bb66729c644c5cb8d351118e7649669c9c49283487ef8b5781b901efc5dde89420e245cdd100
zc879e73706d74358cff1fe092880c04f583012b8395c6c1d741bbcb305f2559a550e289dbb166d
z210fe3986a65f2156ba720c93910625fbf34fe4028fea511a44494ce0f39e81c0d31ea29daff13
zf37d025f250f9e1d437748a36d03c3026c757ce220d23cc18dcdefc98d5041133d847dbd7deb25
z9b86784a8936f1cfe43393aeaa3e924936e2393e019e595c73071e87fb4a46feea33c0f18fce45
zc155cb6e2445597776b523707555a7493ddbc115ab8478ca19b1ea1402a893dd180bbc0853a955
z291fc48bd344257033c9b9b6be86288204ac3da89d0d07380e5dab1d312224b71d2329ba74388b
zb614ee530e5b8f2ab07192747f9eee35fa25a046b659d606d585a24ff4fffa0b3208c745a8774a
z8a9a376e673bae0621a40be26d5eef2feed9e2c22879f83666b49d8b09c60de7fa4acfe5fe21a3
z9f4b2618d90cc2356b6c5214aa7e4acab90583681d9fce7685f51f5fe987007ef7ca820598c759
z3b462188b82136d053b08d5de284dbc7bf00d1446d06fcfc2e946402081886c08cc062c07029c7
zf55607ecd0a6a83f7cb1c03139cc6d4b064bfbfd88b5d03a5bd3db1ace4a6be5050f22b29425ce
z02361beea1330183cd89d87e87c336f9960e6c9c360d3c2e17c6561d999170e9093c6cac08491c
z21dd1dccf0cebe24226d97a3672513d25c07e46e7e58cadacff3289d5bd534631e2bf6f0b1a002
z4e1d04e6bccfaf2fd70dd95f24795067d0b9e24d64888412577aa32edde199ab5d64deb87d7d41
z89d93f747fb83fb159daf0d3a5d0699f8619d6a3836e0e1f9233bd9b7af4fe094cc21afa7fc117
zd677f132c44096c4698aa91bd1372977d27a85ae1fb9c0ad35487e116a598ed6cf0900b555bb87
zb1c1fa88feb8b9f053b89689a63b91992a2e9350e3ddefa998dcc7cfece0f6c1bb6da66fd854ce
zdbdfdcd68ad81fa0bc25483938e7782cc548ed38043ce630269c5287729e8107d354aad9864e1d
zb6e2745c94e4f2778c27c9365542a2d7f012d25328f7536d53ca9fed1b9450a185100b49e9cedd
z27618fe2a32296a6d4fab0830c36567f8b8d7c536e8fad98f7384e3ff90662f6889ebcf8688993
zf0bc0f16b3d08c6ac8282d64a2870d62e796e43299af2a8d2ecd0d24fe6e87f92975c13b6ff379
z3c2539c84a4e8b1e1f2a45a99c11a44cc26ecb632feb6a0b6c3326f9af92f40d849347fcc26952
z73698ef263975695a547342efcf23076e3650a26eb128c01f91a8abda4f73db5dcf80df4ec530d
zdadd47c7273f18cf3915730af5b37dfb157fc5d6d51aa0d185cb0df01afafb66bba6e48609ff78
z313a80c163a92523bcf169f6992b2b30759df3d3c1cb3b1da8a89f9b141f897272e02a957f667c
z6f53e23859464a1ba1a86d593d11c6e689bdf9b3b004507152e15eb34a85e47eb36b13a2e882ed
za7d9c16bebded4fc2c0ba93852cb7d49dd1451fbf20577dece6e2e9be872515f6bd35dbf3c427c
zbd69fe068f99325628a5b0ac30e76064b8401b4c92f5f0a1f8e073728f3b9219ba05e99a59e1d4
zf1f6334f585f897bfad60337f16309190f912374f9b63ef577e0af6fed2500f67ef10eb4b32ff3
ze7adf085f3f9b18cfcf818f1c62b8512e38a5f481aa236f8a42238df5cfc5383cca140ce201466
ze74e4c086d3d50bb338e4a2997e8d52cca9f72fd3b474c7558cf24b2a91cf78ca740b211289e24
z08376382e03417770a73e11b9630e6a0f2e9e160ef854ec35ed1be54551d420784ecc76c632d0e
ze7923d03c555a51b4949355f46ca754a2c77121cd33da6ae726ecce809fd247ab7c8479cfc5494
z8a75e246579632f6842852b259b96bc68071a92e869d12fcde21f445fcd15ec7c6b6203c989a3a
z3e5972db878f14e207553ea565aa7dd0bef669a164b57be6f532187bfeef617f3af3d78c48c4bf
zf5b4c49fa2af2de4e91b45471fae38c34d34fbc9759add6ba340fec210866cf46eef9a300c1952
z1e216c5eafb74c3c205e57a3c06dc77eb5cad3498ca85366be45d6c744ef0bcb159111ec31f7f3
z3db2c4bc85749ffd62cb091fc0eef4bb9ae0144b2284ea7738fce4e286890a3357abca04486ed5
z302640eed6b3b26e4cea43b07e9ff5c7134d5dfd927d2afa75886fb8d18e5141f46c14bc74fdae
z2b9121d1ec5056ee4df416430da4c030107f59d6a0277ffab1cf131bcb562a82d714c2c078a9bb
z3c472cbd8f453ff86497e15af650e2735264cf9041c23a4a7966073aa287b764f47a06f293324e
z0a30d34ff4bf7123a859018b1fd7cc2c88ca98c6385e7e47439aafcf674acea5da5cbd476b5c64
zf4ef8bb0cfab4dd8ef7eb3ae8959f867bc7cb91dbb95e10ccb7000ff342e6d8487f434e6d92167
z2c797dd416ac2b1fc03a60aec304dd63ce98118a04a9afcef2c2b77db1f95e329446e47ea3184d
z0f2c677e0ae6388195674c6a1ea9e1794f14a8cfab1d730306ef24be3e03effab0d86923f88a4c
z43b4ce08ebc022869a9f1857f4e45a5704f6dbe563d90ae298aa59dcb6849c8bae1e29051acb99
z1539d8b5792b393a5ae9c6635aaac9c29372bec36271452a9837de2e05302841c5fb8441e91bfa
z3976a258c1b261490ea29e083e77eecabff6a30553b9fd47a960dbf6b2338b2e63fbd085e39412
z38d3cac750593e46ff76c9f39d2f73dff3579b6f2f3174cd359e3249370fd13cc57a30960e5ec5
z59802a2e3fd69386ba2c2a45c4622a9f83df3331e8209517198d72b831ca4b17339152f0a7b78f
z6656a4b516e66672f95245a6d22e270a427dd515de9e93424e6581014a147e3f4b2d1c61367c97
z1e3d69f7b08efc7b9b37d18bade7f0c5ed50f4c4f084b735ed83186221fa03e179f134f8e21aac
zb39ddcc474d53cf4d2f147529e958522cf3e503038bfc29a5b490487a5a097f140fdb6fa16d782
zdf1f641f11b6585e5ddd8857d5c90edfc0ccf8f176c254324dc4ca96f555292aa915274c147dcf
z428a59b0813d3eec565e547ec26cdf713fc8b38fc6de73eff53eb4922074b6d5a379800e666f8d
z14cf86b893618dca182961042e8d12255a1c9a08acf5e3a8e8985e1bb9833d35a80868b1784555
z8c80d508246bd23ac0d39ec0dd2a2efa3f1a3ac6e348c8c09cb955453a72cbb407bb16968962c0
zadf60f5a41aa018fb5c4fff48fab3fb5796b40905f5717e1e637b295926085865b6a4aacecb2dc
z4bf22be51748c53f1ff0527d1171e9203207c3751eb86014f8e72d12110883b89fe4a6f7632a3e
zc08018292e280e3521992fa7f4fd107c1ff8ea124196879027ec8fd70a4d5cab8b4513139e8bde
z4b9da47bc359f84bd594996cffb780d3537d68dd5d5e783567b89cca7bae967a6fb2a7ef0cfe31
z1de9f6b25818107bd64478f5376ed219d9912556a8dcc92dead821ca0e4ef81f47a72f88ed3eea
zf1f9772499bce92c1936bbb275d16e0823f1c17d06a1b0a947475968b39594f5dc8800b55e65bf
z4220dc68fa48e49fefaed790c44ca6f67479fe11d4f6a32e2e2f90bc30dfe2319322f0280a9b8d
z19d25eaa2eedbafaaeb92fce058aa3941ad5d89a4e195444719b6769969c53662dfb17883b2683
z2833c53b216dcf1869dd0443ee349f120867e48608e1a0ea0dcd7a464b465078df072cfe72471e
z588d614869188450a6971d73c695a6ea4c903e92eb260cac4cacd81d4d4ff69e3a36d96db4e027
zb99de39fdb0eb7fa0d0ea656900f83ddae97ace8d5454779a20d1bb2bf612a9471c9828109be65
z900e50661b0dbc5f66c9ed8436a66056e9530f369cfd89dc74e1d8ea699b92fef54a5eca812d14
z8b79d74d675cc4299d5573837b54342d1d8e80a515fed29494d2b483f7b703bb31459fe9c361f3
z630dcf8c0bb201801be1a535cc2f1c6952319199acda764d9638f991aa8e0c6acc5adb54506929
zc4972feb34c48cc624feb4a58d2a00d1af051da416bb1ee061fd0f94665778d4de9f37dda3d682
z278ab20613c9b28b498096c34b443a009216509ee12751ba8c84d833cff07e9abed9dc953beade
z4cd245996d58d17b166c1dfc0c92dcabbed965368e8aacbd0cf1f45d911e8d382968db4957877f
zef49370db3566d6bfbd36c3a95a5a0fe4c1b45b5af668d53a01f1d3fbadfac656cc6dbb68bbc90
z8a538be4b6984cdc1d9ceff39c8c448a06715f2cb134bbf6c67362a7703e878e6a55f2645d3660
z9f0f657e2ff3f77b688e0a5606af2d9f65b33f44c17ba8c9b8170bf8bdb13b19e0f2cc079f45a0
z9f229bbc8f4ae420bfe5cd5da6c952231481f986cb2022e70221eb73586a65eef0ec3e5bc87f47
z045442e5d77077790b196139719de61e48d4f485c743101568052ea2c9427ed801e90d2830c052
z11236193cee1b8134a607253f3bdc2bd11ea2f52eeadc0d617bb3c696d61beb074651d9156b5e9
z279ec9d3487058fc7622c5b6521d60148015845678d16389dc4243a2a8d374053b93ac4850dedf
ze666d3aa43691bcea23e3f5d5edf1c77f43d681b0cb30c53ecaeff0ef6cc17433d0461043efa2d
zdecac0ac2d96bfc21c5f9a686d5acff3ffe0eb9592225ea799022a24326f68dc149dfaf87a37be
z97241ccc0f00cf9aebd4837680e4fab6603fedb4f6be66217f9a53aa4b9a9b0d4b55d349a55a2e
zf095c6bf82283b3d6b154640d1723fc4ce4ed104d66d922fcbb1c0503b58798b4ae10d219d4b1d
z5c91b5c3805dc851e99b0a7fd8ccd863a92ffe56c353825fa26135295d195c071937ef64449b0c
z110c702c7c27a65c4d766a340dc2639a94879db2afda8e38c8f4a679cefb88ec914498fdd28a20
za4726f17b5a39ec365887fdedda648c2114adde020ad5b6d5781a57ed8c0c3999cb075f4b4ce4c
za3eca02f05ad85041f82312f61841e4b537ebc727cd8e66901b838dfc32458ed384eb722fd81a5
zea739b9e11db5740f950d46885334183eb26f8118f54176a24438c742231763513baf5380b7749
z59752253f2121c05df51e950e140bf2a9ee8327d869e4d731239aa719135a935a48c6e82ede8c5
z0382f9d2c23df2668b265492bb85fd58cee29e30fc69d6c4c2c3ce75337fdb94765c5d443d39eb
z40074dcded531fb5064d8922d1e0460c742c9aac76506bd36f3b8b5ee12e26902bcfe6f3195e7f
zc9ae5b0ea71bdd6222ebd21e2617e3873a8b75f0512796a080e2217e2b104ac84732dab945bc49
zf8c1f43aa255dc58029f11add8f4219cb33017337027620e3388c406cdecba1691775dfe7cfcd2
zc3c1ce06095cb5dcf0786385f4ddbd68742dd9ee1077a28ecf8fd110b740026a829a1cd6335ad6
z305dd7d6da4c0b92fba3d692def3959dcda823eba88ccac6c05627a27e195f0ddf121c5ac1c903
zca3b2bfe0f59390a745855d7d31bf2e6b89af91905f49520f3abac18121cca1e5576552f229258
z5fe051212e179c682dd6500ea519671f2e21ef6db678579d7005fd9f0ca57c8d4bcda0579009f3
z6881a0fe2a68e63fa894af1c80c8c672773098a36f11636c822a34c161b47a0f45e04748a1851f
zebafcf4c809a693a2da0a5cc7a3d5b39a61646216344ca078c753a3e7089a7d8bebc600580d419
z0c804e08d9b092c63f77198e4f7eb7737937c9546e13d12db6ad5aac39b7c15b170e357728a247
zf55d890e92ce25e7e0f158ce0380e80dd153422e1a2202fe051bcaf7ccf94b096f840c0c6a50a4
z7ed499f0e0c8338595c2240bd04467d14a15859cce7c170aa3cb96ac73a9d39ddc25fcfbec110a
z136005b8fb671642543b174f7be253ea2d243c915de8db56073b9bb74b66c37d33b624811feebf
zc69f56ed90e7ebe8d847097f63ff74946843d34a44b6d0e53a88e07691e1de680af99c63c94b25
z393a590b24aa1ea21b84938b7d806896a7070be5d69376cee949013a0c6cf34e08e1adbe59b11e
z4159cc3f8518b232857de267c951f96a58e9d837439f6232763f1ee942fa53fbe62298e32b5038
zb94aeed7caed38cee307b8d6aba58be0c329236b66088dfc67c46c0d70577e3858c3700db38f9c
zc12e9003d217567ec219e8794ad38d407731c42e50246890c5d1f1bd9ff4157fce1b70a3fe822f
z11b2134681ef4ad86fd3ec1a96703031ec244c342dd21a3619fc536e2f5346735e10f2c15c7d2b
z56664558a85ec63cc22373a611032d42762dcb67418d9071e2bf080cc81b08a8bdf1e175ceca53
z4db60dacb12d96d680b2158cf65cc5e065dd0d97a198ddbd3c427abca5de8b1251c62f4fd31b71
z5c2485bce899b376ab376a7bb9d6a0998a501943174f9799c416c22fa5acaba8401a318ab61ddc
z28cdfd9b8db34edf1a6bbf3a25c325686242e3b0669677422e0cdb841232f8255292dadb31953f
zf559f5b9ccea82c81af951dd3d420a68faf4e35d3c820bf38f029bd8d58bcfe899c71ef5ec818d
zabe8bf5f490daf522a2a05818b5783ceeb181f2d9eae9e834e0ac3dbd837ba89c0756afa0425df
z8f2b0a4a015982bb0b32883fdf05dd03ba40f0276ea5348c17dc9b68128638e5fcb36f9dc5da7d
zbe9fff752f1b366aad8af001d5df8df66cbbfb965fa8d41dc8dc12d9df81103120498a728a9572
z35f07f10c1d8bf3ab7d642690274e71d5075494b80979aa755f298c9a9e2816d9a031fe3858846
z6954d14e17a1846c78266a650b2a62af13fb39fc335471958c75ab035c2b9a333036118e7e0b5b
zb1295cebdaf1a1f6c6914368383a7a39bdf9befa2d91ca28b041dc7b1cb982172ee832179dd22d
zb47df1b1148b63ce94435b0c4d02ddbd47aeb85c5415d7184b7ef730e55838e981aad147bda6e1
z0c79a6f3021ed8cdc206a5feb36218028c223b501e344f2dea44600cceb220bbfe13685cf81364
z30dfdc5bbdeb23c3417fcd9fec479f63d1cf825191c0671bf5a777e95efcb3da5b01fb8050a870
z3766d8e9e0f7a2815c4e2fe6c8ed2e4f21f8ca7788c247ce0403dc29be58ae782662bccd70b168
z4d2193ecd33c674d9e24e6792e9f792c4cf47e045b7024c202296266c4374fd461fb705d8c0b29
z083bd2e83149f396224cf012aa1ed64e7c0342dbee9a3f2ef3a449db8e143a9d7130f2328a9d5e
z82696b2457788d6da287498a01557f33874120981887b9ece6be5bff544c496a2e347afd789321
z40896761be75e2824cae33121f06af5c5b2417dbceeea83addb30754dcfe3a3338b19f9ab1e74a
zfd512bf168e0a36e3a8b7b4a69aa37c8d6454d9b08d2a86804ae4d4e6eebdf108c635f42b65ec6
z0202c1a58edcb89a58fda8291fc4e8f9a53d1260f5b01fc57b2fdc9368bd6c0b454134e898ce83
zd6901dd7a5f94b256ebee718161d191b66f8d6a3ee140898d70b788c6997aa3e20df1b22ebcdae
z896fbf17d561ac783e479151b7611c8cfbaf5fb1af28427ee2d043ffb600c5767bc76c214e5ee8
z5521fa19d613f70b06ff17722948ba6b2c93c7d017c72acd1cb88863825c51077ab5552ef090b0
zc4dba892c8894fb75b37bfa661c78ad60f9a0539cc925208985f255d85ec186d86ee49998c1abd
zd6cc73362549e3dc1cd06d11a07d759157a4ef516319310519dfd5b669f06837d93622aecae756
zf2dcdb2e90099fbf32df0f9222e968e83ce14fc8efc916fb1a889e311ac8ed57b046576e7772ff
zbd87b58b0fdbe70f9ba7955bf8780a1493708de86a0dacbec7d660a2be43b67771f7856a30024c
za0451b3ff71fb85efa52bff1294fdac057b2baf652eb2aee993a085636a74be47353affe9162c6
zae5a769fd328d7e56a03a8d487b2336dbdaa99af552d77f376701f45cef4390908323531ee144d
ze0fb113dc10c7d03108826c6f73adb7573529fa63d96ca598894e3b02bee35f975d83323428403
z16537320a8cb0818045338b980588d1cd97ac0c17cbfcae1188972e33d7829efb79bb9d42f285c
z0b835e95beca2baeab82895f27aa02faaeda4c085c2bcf92a9f7206faa4e150ff07e28790d5d38
z91839c79d089172ccb8ba5ba30d93045518aa1bbc27c8ea24176a02ba899adbffb817056835565
zcbd0d222c2ec26b83f5b718820f8f012c222d5e052129f8ff2cdb7061984b96c0db79ca495eb71
zb84fdb507a9be1678235aa72c1b55fb3791e5dd4352ae5b5d683fb64c1462091d0dafeb22241f6
z497a4b1c15188acabe382c6b6ef6569d1fd820bf6730b98f2582a47e0c5f75567f81f02be280ed
z0184c30edb4ce1a30fe32fb60b7dea0a88c3dc164bca3416f3ec91aab8f44c5375b23a551f027c
z2301ff00e9dfb09db978a4c33b709f86893ee7f540047121137f482f814949a921d308fee63e4f
zeb702c6cdc8fdb02fef9b7a29e44b43415b9a0ff04743ea760ec0d9a227e29ff32d6ed57cf73d2
z7da9a58587299602469c72471b8c5997993cf3303c7938dfd29e13d7d4c43e32c754565cc21d6d
z7c87e55cdf4acaa43aa53387b9f83ad67dc13c50df4c919555983180cc0ee24ead3192e81dc43c
ze21c55a33adc599fd4a61b590e20aaf84ab272884a805567ef2fb6a96dbfaa138e72eb504133c7
zfe19370547dc1955516f9a22b760ee1447ce4cd8f5fbe1b7ca5dddbd91ff31d1bff760301d508d
zd50ef3497e577ab9dd35730d0e87b6501075c8a1facbee6e1a2e4de75382aa914eb073865e42fc
z6ff1f20398d630ea89bcbcc3e28aa21264ff820a6787bf8adead7276bfec17d2c6d47696a9d9f4
z6e2992ca4f2d9f09002c0c10122b265e596f0d07adf684fd057902c9043645274f6fd6640e2e6c
zb05ec0e82be501f6681249773ed866c27110547fa63c83f4747127144862d26daa05643aff9fd8
z84ba3ca760af3dda5752fd468bcb328a177ce19733fe0f581359e797ef296c4e1ce732a979ee15
z162545a6fe6bfd40c788b1c3a4f87b3155bf5ccb115ef87935948f970df8d31956993c699e8946
z0f31ae232eba1b1be556a4eda732d7ba95946c79d0d34b9a5b590a87ddb9691d61084db2e215f0
z1c2f30f962e2434c68d8c1a53f94a0de2c60c23e0048e9df14533b863ed3b0cfeae39a8cc27cba
z336271f662510e06267ca9f562e9936e9da043de1347101058633b73b74268b3bbcc7c9e0eed0f
z16ace5a0969c854fc90cb2899365fb07defa648705a73dbdc0432b57ee65f406d07430283fd51d
z78473ad982912b56cac0bb362dda788e9d21771251dd835907f98b83a918d614fbbe942a724b41
z9816444cca0621a25285d9a82aac1c402fa779d01c0dcbed001b73332751aa7ba9559167ed61ab
zeb15c969d7a3b1a561ff9c181ac4dd4e6da84ecf86e16a3276d5baf4a7ff0d886b684fcbe92dc1
z71d74a8f54a5f6be4da2ca804e594440c1595e1d90ee1201c39a20139e1f00cae8eb5d2db4e889
z317db5fb639e91ba864e36806b8d36eed9c75fc76b4a2f6211a4f83295196b2ed6dcae3842f6b9
zf9b4ddf645e9586d7d3998d017abdb4963f1eea1635b754ed3b82684c75a81caa918676af7f22f
ze9b0ba771946145496673d8697392d2e69c9ca533c25abee35051647b16d9dff5ca3fab49bd8f4
zbce72ba0ec06b929a3a42685b3eec9926f23d37bede5da0f8a596153fbfc491ddc459e9013010c
zd33a3c7b58bec4d1c33be69bacbcde57dd9c6a331f65755b854393c350d33ba5d5a794e6b6b3c0
zcc4663d5cf492b6ccae791d2c99cbf743e4bed76ab897b153644aa3f9b8b30c2dd34b2d1bf57a6
zcf295729a907220031ef489ebd4c250e577dbf11db7349dbbdee6dd8710f5bd404f36cd0b70f14
z5091a0352c542c740ea9a44de5c0bf73a4e4be7ec3163836b6ac452805c4d566b86f9c3068368f
ze132fb7ff4b3bca71c20597f1c4d1d0bc2de4e7df7cafa5c23ee80576a40faf0fa3ae3b6d355cd
z201a7c3696da63d389031b699581735ecf91a87bfe2325528d05d03a5e30654f69ccc46f35d8cb
z2a5118c78813af60cbe3e8f2c90bfac59dc355f8096e0e9ce54635c46cf1446c6ef27b98c3b16b
z825a248c21e02e17abff01cab74a8527b96cde96de1cdfdf7e4d4d385569eb568a79e9a0197ed2
z450db76e92908b9b137ab7d0fe1b6fcacab90ffa5853274d064d82dd65f056f012052ec4537e9a
z6e52a016a6e7e0a936e8fb71b17d6d12ac2b28da77f3b11b298fcde01837334d31ebc97bd50b34
zd165db1da1bc82708e58211e23a18139af623466dd238fb457925cf421651e356a78d324283820
zc9426999aeac87bf4f165b1df6d54872d3eb994e4d6b6ca37d78871347bb1ea7762453f0b41574
zc7439152630e772faf164a799b0cf1349526b39024017f6f3b5b5e36083b9b4d6c59282175c55d
z7fe98d84803df8b97a8bca7ce1a2cc7db874b9dd844013fab83eb686edf6ab47a826c925d1d12e
zd3deddf463f5df36ccad7107e5a1ed8fea6f81b2d04d004f8973f1821cafb88669107e9934c336
z9b1872ecae14b66b608f3e8bbe60a3badee5ffa10c53ef0e9aa08b4852cb787fb7de4e8757c78e
zd03f2630d0d95ead23148aa8702aba60928630f267ed569ba7b3d3990d9f79ef4078eea415a0a4
z79e1d168d1677f21baed1c224963ff51450ad9321a6fc90e634568d5128261bc1e8491087a06bc
z6cacfe92a1f58674fe5d576a01dd85fb8d3fa13c9146e4157f9e4c7a253b92692057d061415bdd
z1e83c90e116f4a2d1f5be7aa78a70246dde687d1b101ed3876d39231b126651f7ada532b7c1749
zb6f4fa7d65ccef998f3fae132257cde638df4bcabb25ff123916800dd35f72e60aa1d2eecef2ec
z61a790c509adbeeaa08dd7ff47454c1f655bc9b6be9ae7f908934677b5565a028936a40aa5f719
z74ef7926c40d3540869be03a70646cf0011f8f7ed4ee6046be1808492c6f789b5b2cf8d9033720
zd599cf74af0cfed286d304908ed94f946c2356394185b43b5bf1499d68ebea830c3d6be0f6d62d
z54aa54def8b63a5b07f5ecf3b486ac076619d0b9ae349017363b643cab5252717ae7612be0cc9f
za120cbd5cf97839f8fc3adba00fdfa5f03d15bbb99bb6d98d2ec2c0cc68d5250a8bc5fbdd033b6
z919936a9c17f0bc308177fb2064fdd3d9066c07bab41a2733a926894aa84a829be74c5f41974a5
zd60dd7e2b57ff20980b5a2c67ac584318ac8be75638eaca1d6f0f8c672de7f3572f4f15d517436
z88f8c9770ee683929bcb22f4ec1226f0a8ec6ac43fd1dda3d6eab60918f1e76d9aeb9d693c896a
z085e53d9b6a7731479064f4541ccfc5a1d0dc2ac9e78f5059a75f447e009ee3fcf87bdeebd93d5
zff849be53e93e42a07229aca0efbbae261178c1d92884bc4325c052d7a10aa2f67dc38b3580e35
zacd13cabb259ee156eda427339a9ee4f25999411a1e56a68c3bb70ab040f14904c466423699fdb
z039f1824439c4b2b99e8760487957666cc2067cf0943ece024e87fb507df587a73d21e392d9a3a
z2b5ac3426e73f0a3cf413c6096da480e19de2d4b0212acee4848f50eb241f7306f86f1f1b889e7
z5754bbce4be985ffec22e74bd0bc18282759af59bcb58559aa0e2142985b7e4be3d9b8ffc652d5
zc07965987fee8eb198b23f123aa21e74773cec7b1a27145beb44682621c466761754cd94727611
z896b9f26b43c38bf0beb09aeb823049de25721cee190cc76883097aeed58bbee29ea5035143e5e
z2b058db66e25e8e7cd29d0ac9f8e91d5a844698963b60b5ef59c1f03595be7cffa0e5b96847f96
z3d515b7252b5cdc1dc3015dbd63db4f3f29e974961d355f84874f3d7018ba09f47f44c46145b8e
zb786a28b22bb47eae66d796e6ede7b53131dd589e13bfb86e9626797ad6d59ad535a2ee1b628ff
z3ae8d8d73d7fa34b43c3322a367d32f3168611d4801138669ae7bef652d51bacfc2f0c0817e217
z4d38dbd103f6511cf71c3d6275901d11a00255ee36c413d93c34cedee54761abf1be7f76a0c579
zd6c86cf839506a9712f947bcc31bf890a664e843f0bc1aa14ac52785dcf4457902314a98dc1a33
z04a23ef1a021b4e6b46c615f9012d4fc17cec152a8cc61d89932c02dd3a84943b052425ee14ca0
zffc1471b1e1dba214942171305064a873efde34b8846531c48360d92232f962aedfa6fd779850a
zdb3077ae22168b2819147d7ffdf8a92d2814474124675b9e3371b1194b7449e8a950eb5ae5bb54
zc6b4745ecb869ec378dcd1f92f23a197b16c59fbb03b1c300cef44d41df10409fd802a5d882399
z8078bd728818dada6f13e13962c2c82e5272f4303d53422524e3be620a6dea4c2e1d5529730e7e
z65d1022c3af4e62ef29e5996394d9c714ad8867f14795430a6d1ff75834586e199a9e51be80776
z8b67287ac7df5f8f86d86e2c77a53a57912213fa8ca2b364c90cc0e2070f6373e9ebb3c2b75905
z25764d1211eef086da99beb119a4b40163335dc211ebf55f6684290d2b222d797edbff560f781a
z4ba8178cba06e73967f76fd7e4b00480b7a2e0cdc937bd5e56736f2c4639e8341b2108173f0d8a
zef8476edf61c1a5a48ec8081951dff59a243f69f8736770868e3d10cad82a8f948ec1a080fd595
ze0cdc2349a1eb55fee98f13f6d3e39b3e81ff4b2d41051a2e2969ab41e217d8ff2db6812cf90ac
z6487fbaf92a6f4df7e1a8cdbd88230f07b5ee1487486ae50a6a68ebe74152b1484a7596b0873e8
zf3f90e4e627951c0a92ce3a997e670bb5066b974a510784e8d5f1f2e8d5edbb2af69237cf3f865
ze9cc457a82aa4c496be2b6720ad61ce929259ebf741dfafbe17b9aa31a3c669876452bf08db4e0
zc5bc0baa9ff470158ac62ab9dac2e78b72c9179d2f8d0628cf45ef64d05f035a930a850d4eef1d
z3c544dda0f75d6c26bcfe14b33a21d759e5ed37d8692b6dd0c71c116699bd20b7ce45fde90df7d
z81a5bac28f594e084fc169a14a6dbc18603c14f28f6dd83c708abb2d5a06a7352735d2de627d4d
ze7df3f501000b92ae46726478eed9f0f74b3449e364409d737882f763b5decd1006bcf7115d718
z8fcfcc64e7d433ad2a16a1fe97083a010ead34e1fb77d7ed6e1189e82efe933e30b0d0b209d407
z64eb376fe456b91bc21c493cc78a885ad3451eccd46f2f767b43587e5ccb5ac9c25562e5308fa6
z04b54e3eefd26a4722c810a5ebb85169ed469a8305150088dbcfe06027075405c775324524b4ce
z7b033254502a31c46816a2cb95dc5871fff3ad178dd4cf1a7cb9f26e64f33816d1eb57230636b3
z115b116d2465eb98dbf12c138c0ac57e795d5d6ed6931155e091dca13c35813fb690574cf56101
z539e398d848edacea50dfbcee00f26b0ace978448720187e2c5d016d81b34254443d7841ece26c
z017d8f18635b67ab831a91e5a12c7efca62b083424093ee0d3c8b95f5ffb5951ca1dd32f7fed5e
z3e7e41bd26638a88163dc3c90362d3224b3597515dcb623c94be66fc904a278ccc062f92269f8c
z052438e95fe25fe4eafb836170fcb48ea1efd6d8845bd0fec8a6cec07092dcef9ac7e96b173006
z22caccfd609b38f6bc8711ae2799ff8efc490839529497f91d0df655635cda6db722b9af4dbfed
zd1ecb8cd24ec93e757da7ad1a77c7b5eedae235f4c8fdd902a17c9c87ba5925406ee218a6e44f4
zc6c9e10df4c62852c44ca48b5d0f57d0d6973db30d67a53bad4e5d3b3f55cfc79cd441ad54ae5b
zdadbf0da9b5890d66c4ab1e35d8b63fa9707de8fa1a4ec7265bc851d1c3d2acecde5c33779c55a
z42933632b0b781e927aad058d09163ea80a57db80ec62256818e90c7c0b3190baad0580fe14824
zd4eb1e56c06d96a82bf84a7fe5754215558f2dad61635e8841625ae0a43cd69086f51bd7c930fe
z3cff5be4ad6e767a9fa0d78cba4a191ca8cb64ccc7597d0425fd0c38a69634ea7b23732dfa190b
zb32bcf682d5d4965249ee0b7fd4499d8b0866921fa3294e7dc9d8b3a60a12dc00f7f74217a0ee8
z839bdd857aa146e3336e4f016faf6c1b7080bdcae333ebfee89d5f11dac1a27116b2b593177910
zc6a75ec60bf68ae041624da470ca8ce189a484e2bfec37321d5c554aafbca72fc72f9f0267c532
z288fea11d2e237b0cdbc1eba8747e4c395ad601650c3fb77ab2514068bcd6f4457ed198b85c805
z2d6d7ed91f09df524c7af8732e2784d531558a758efef08b73a3806ee450c058eceea93ef1f736
zff9cf1fae2a1f40220abbfc341440ae2844fe906495ac0a887c17e6defa726a6458c91e508aa35
za1ff662b8916e6192a2578754b081f8b8f9eddd3d0603512a5f534d43f54e6168e209a91c70e09
zea8056cc3f85bec5f5a618489d66db5d1c4b9cffb24fe0cc0b153b627f7f84c4a71c63f2b95703
zcbfee099b91e104dfdcdfe73e322a52bb8acc0e324054532b12cecb2af77c075aa37d9c818e5a3
z8d7c9da1e6549164ec62001e1022b63cf27fe746836b66ee771907bc2ff540dc8cef4d9c0064d8
z837139162ec754e9afa02c62feecf82846bcad39a09db7546153ce8b533719dc7cc98ee7d2f6a9
z6143abffcd996245c9a2d8253f625452df2e600d8b210063e44ec6a2fd5b800e147db5589250e7
z2ff7ecf89c124e7db25061d3c9714a172d100bb9cb0e755c7d42cd4b666a08cc42577c952338ba
z4087270bbca65c78c82609e2b3ebccc65b228c39ed7bf17d4ac0b78b90fab465f33fb5f8643f0c
z887aff7f1773917acbff18c1de5ea7df12deab821e6533e4ea2e733e16992a9519a7c41cded605
zc9a360cc21f31d906a53c168a996fd90b91466082526a9f152f7e2910fce58b49d036fd34e3d90
zd8fa8a97b029698beaad16dec464f92a98c8bccaf74a7edd3c5cc0ef63ec458aac755c0c67dff8
zd71250f1a44bc8278e4b0d64b765f1bd6db2def5c750311c0e57d45b9213afa859bb3c5e0d53cf
z994df23404716811df1287afd6c5a900d2a90ef6f2705447261a2791f08fd19cbf0c907420fa7b
z90a74ca1e14fdba04f6f2d99e7e81a91bba5a43d02193c8f82d2c8165c9d24bd04b414e6752fb2
zfbedbeda9f8d76c347c71caec2c0db73a0d754225c5e116a9a5cc69c50878f472337a9e7e0bf7a
z2c375c0292f4bf40ef6908b40785a04428df16fbb3816ef9ef3c355493f4985f649a9ca127b2e1
z42f8428823f4a894c4b17738774acd14a9a5ba763207228c64fdaba381af2a1989fd307de54989
z58b9353bfcf8d6f8fffacefbb1beba83a312bfec30f559a035eff563a3ccdaea92a1864b8c49fe
z343587ac7f049389db3011f3fdb7f4be0b8bcede221ab05efec1006d248d28ba689a8a40052c1e
z2ff8256d929b1a01a2a8d0f1cf7eeabb5658e18ffecb64a82ccabb1fe6549da1b93814471fa30a
z06190b1ba329aaa27de0b50cc7e1dcce6e686d9a1145a4b1fa83a80ef09ef48523844c8007814a
zc272fbea283363a796a30d94753e6ba540c859c71654b8a72ef56527e9fdc59a65f868916a1e08
z4f595e53313eb88a3d1703d6f6d08d1226b783168661615ad3de71ca213b24d1bd2c9e21cb6b15
z5e2fbdb9c21f66822aa2154c1cecba76cf9d6e5fe05cdaaf0602899366d178f18350f859c367c1
z987dd143cd0db908bb168c1a243c97bb6278b8d182d2ceb22a80e918d78518b12bf29077bfbd9e
z66649e6cb6af1a3395b7b223c583f453e6810c7e30d4d6178aea29d83f05f43dfc68efff9c3189
z68f912e3229dbd42381bb79d3d185746d7cc2c054577acbdf4ca49a246def139da21fa8718e7b8
z71d16e94fa726909e448abaa7fe4b77e565c8cc3338f9a432be52f54ff8bba5668d27c43d29802
zd3ec101320dd0f1128615de5b55c3fd1b4005da112c4c63d4b3f9365e5c5ff073f766c0f3760d8
z18f90d135d8a170ce5e856f9ea60a3ee29061e05e922fc6a02695457ef7f30fe8571a70a2ea552
zef0c165d37d94a027b28536c8fdeb5dad87f621188959fd20f5a10d087d256680cbf7607fb361d
z0f91619428a9ae9a43a32e3d8d56b4c49965c9bdf0eb2017621c7d9696233e1dd42c213e8254a8
za5909d94ca85dea9a9fc05b57e8ab8c226677bccf4f325d2de4387cc458457de22cf56b87b98f7
z61f4d57d908741ee0a3970c81eb03d7466d512345545cc8ca48a6ce5b9c30ac0da76aa334defc1
z430b3cf9cb040e78eb7c147ae39b673210d2a14ea68074ae657f65be256b9a4c0e7a96ac7c2a79
zf0275400afa28cef4af7be6a7497b194b157e1dedfe4b36bbf9a09db20a8c348036fbc22f0c2cb
z507d54ec97e219029fb87d6a5fed05bf8f7073fa29ca7c7b5559d7a39ed9d6702e425530fd8858
zb08f159c8015e57b253162a81576a3a40956e0f55a1c39229dfa0e51a9fb45a23ca4b3c86e8960
z9c453017a26e9f049b3aecb16e636c192e1dec8d9f6d5ff1098d4b674714856f3c783088f41209
z43d46db2b103363ace788c1a9f4afa78777e5e4babed53c6022983aa57329064cf1b0e359af6d0
z3743a40107da06d9709834bfe47d464eafb4813acbc636aa86a4cc8231cf40ecd2879656ebd76b
ze5580f6ed37256bf156f4a637c04fb2c183e382720b36a4eb13d5c264fa26acb2f6452b93819b2
zf1d68cc5e42808f45c62a44f72b5aad144d21eb8c1fdcb2000df4f8cfec1caf6720023e1fc3639
z5886bc1acc4561de73bed051e6ed59e2b7bb766d99dcf256f5195e99bc9ffc90ac2813ee3e0691
z48d1af6bc7ac5632f8210850c7145670a5c0f8cb35bb523ee8567182a74b0465165dfe5af8316f
zcd0de27b3ec5d93056710cca809ca961d8132009c948513b2e60b73206f33f26c1ca2f1211b1de
zb686b79e694f8386c61310efcecb76d54f9286faa45c388592f85671359c39f78514ed6e2d12a1
z795affdb1bc2332904721cd5cfc741005a0a4e8bba15921fa7ef135cf7979d6ba3ba79b88bd0bf
z1580be9055f9a9e361bbbe26aa6295547effade59112dd6e849cc474e155eb2d6743c015e54834
z4c346cd680a7559efdbf486dce4e7f87dc2da511e8c1eb54d550bf8f6bc37464f755c2d598e9bc
zb90361996ebece7b39814286569f920f534a6884746ed1eabbc61c0f795f01027f08ce5c844d55
zc78aade6bc85e75275dee9b3fbd8a9614eb22b989b89c1016ee48201093b0582536db52d57dfbd
ze1cb6bfc1cf1760ac9a694578dd110e7d3be502dff0fb2251a6a997b756279957d2fa958a989c5
z4dddf156a04ae6fa9dbd55567adb813e8d99dd30359c659f54e9443eb0bde0de3ec25d58a08b97
z3ecc162814ba96ad720a8361496f27b641f2f234c369f0ccea5714cb03af07ab58a4dc2b458baa
z17f518fbee60f20ce52992652e50ea153eead1427d967289a338bc58312056b5b78ac1ea246b0b
z6e6e6f5eeec723b3ce2e79b7be16b1b908ed4e0cadce4c9c13428d9031cee38c250bd5141a3ac1
z8edee6a95626c4090fe151639bedd5926a6b1a80d9adc7f31cba48f344827b6a8ba95f5ea084d2
zbbb23f1ef05a53855504616407fc2d6f147a80f3208d5c230034ed08373e9bc14c972775972e42
z545937695f025f55d73f45830ecdc704e98180cbcf9f8646455ee2e8f9072cb78c424d73
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_timeout_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
