`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699166942afea5fb71013544a379d857e14685a03b77f81ac
z296de8f163f6909d2cea8160366dcd1069a4ec7b3eafe2a3ca97cb83086a74bd9bd0fdac0291af
ze44ecbc1f91d60b48acdd3afca719670e39357f5448e977180eb5cfab3de63dff72cea566f1646
z0120c08938d14dd8a38e1ee382ccf375cdfe4d19c75b0ed7c629c009781b4c8941f40c232e5f43
z17b5146380d9fd3edeb219b83674d2b7a1edb607f41678cde95cb4b47d46df23a7fd46ae218b37
z0989f0ea404f34e59583bc532b4a5e4407bd70c0de32180526897537c1b3224a441fc88708169a
z00155d21c0df2df5f465101c77bc93ab00803a4ee64bc17033a6405a312763e105117b518d5594
zb11b72507d9a6b005514b8b6a15fddee1b21a04a517c72efad33b87a1f2b9456ba6eca4fd6a23f
z539122fe8615670ce4e20bc6a14eb2879d240e20a895946048d9091cfd13c6911629d8f4c21684
zad62f70f250bd7deb0d6f359daf6e4a6d84087684f3c28a718783b43f040717f11f23555680682
zca7a224b3608699ad680981b35fbd4a767892ddfc4508fc7ab58af7ca1dd43542edce52216d2c8
z9168a4e192babad85b34d9739353ac4dee29ccbc8a204441bd447f1cc60a09a939e4fe53d66be8
z44b73bc0d951f02124da0d2a6a44eac4c1cce5bc3780ab2a8a4564711dd46acb375da42a8f73cb
z7be9c655909357183550acbfde5e3847260331afc908d95aff58de325ca9d3258a2a0a32c1e7b1
zb41ca01c1b0664ba10eb1ac386dd269cc930227d2c6b211157a028660679535a53671c88dda26a
zbc971d50243fde0f73d8692216e4ecf74b896f19a68f9b2ca3aca5b55ba05bd5457183d6ed7ff8
zf560e42a5cb123c0f5ebccad242f1c7c4c4cd3b147d0cb212042457f25ea567466af2a63edc1fa
zb2e7425b666e6945d6a3efea85ac48b9b8dfce3f01827efe3409fb9e53b9040a382f20c662a800
z23f49381cb580176461ab83bf783ac594b5a239ce1c57d27db1146cf6e74475b84e4574a032401
z9b23aabfb517a7803e6c8c07adb9e9d63a561bfb1599cafa9c0eaff79067f4fd15c5fc1948fa94
z8b0c53457b1aca651ef7911af5d5a91d950c2623d27969fa31408147434ac29759adaecb86f67c
z61c18a5fb08904ffebf86971fb4ee6edc3af721755f1ee9bb2b86cf7d81944eb594e6d89e63c46
z8acdc824d3a8b646da46d86a7f457a932efa1ad108363125c8adc994828b687d5682865ec5e2f9
zdcb37ebeb8d520211cb2274d36d667bbdc6deb6fd04dd1f222bf000705f4556ad7adc5e338cf14
ze222bbe0525d2876834aa0d91fbf0c328bb676fb05ac97c8019f84888213d91bf7d5b1cba15bb4
zb72305cde5396256e0b40965b557a04b8ba8acc2384ca7f096e6223082fa0b324803a218348fa5
zeb0679311369b34382b1048cdbbe596945a4ce07f8e8ac3685b8ef1a5255cfe22bfe68f59ce325
ze5090775c24ff7ae32311d59845be858fef2f9b6c5c8dbab3a2f6c99e2c8f953793d15eb34e5d9
z9362815c451624512330154230f73f5660110e1c2bad050641ad884bb8cfc6ebb2b971012c41a2
z0cb0781393fcb2141fd6c4a361708b3ece7999dc5de45bbd47c80b85b45883155c8d313ba86d89
za231e0c7120ea0c6e12f4dc4393330e441f613bc5aa53299875d32a8de6e1850b61c8f02c38821
z0a887c7bdd6b2e42217a473ceb83582432e8a5b5adb3ecec6324fa6a88a183cd374759170b82c7
z7348dffa799b718bdba22e735271655351e67cd2e45b8bf2fc99315be44defe2bbf1f5adb54b3e
ze5fc80953406519402b7036e4123cedb9f981525a9c1d9be86849cb2239f00a7f70b6e97da32b8
z31bdad077e6321d970b0933b27a38e75fcc56fcbc0ace6e87fa0a85acddf1c4b6bc2c664f4f4fc
z53864cac42556b6cd56dc3f84b7f34350b158f163edad73eef36ca880f7ce955b0d5c28dca832f
z3e51b8e52ba480e2762d623148071e1f24fc7751f89b49b26398e1845156c89ea2cda7556bf079
za2df19ce839f4937d4ad710a41e424a320290c5951ab6515ad71f2ccea3f4ce04b5dde69ac232d
z52fd7409117a6ab01ccd653f7be2f15441775eee5725142b1426a550acf393d825df6d8bba0b30
zc0d853340e17411ca1a83f5661ceb46d301bdeab0c0bb9cef5e519068613ee7ab8faf36a981686
z2c59f6c639ab950c18be7763086ba66d84c5edc5bef85ec155a732064ba8457d02a92a819117f8
zb36a85f40af5c583b95bd7c42b870e7c3c9369484aed495fb58e63e75c732aa2aeffcf82d30670
z6271b0579fe2fb32c75c5a49f10cfe2adbd67f02678ff614b7d3e12ca3c059dc0aa883ba13f187
z334786ff74680ed248eea8e3297b29856de6b13dbd0c0c80a40c1410597c9fe35be63dc97de4d5
z160817ecb83b2e6c23d4c117296de4bcc1af9e520d43fce07ca0ae6bf73f9fe74fb8eb0bcb962a
z61d90045b47bce15a65df6334ad393cf2c6be48a32850509bdd57d7e690b7fc8128a5d106eae12
z09865f42d05a2f30733e3f165ee9b615fd3ac240a4296b0ac7afe32252e3c43722011867802f42
z5afa33c457d919c0416aa6da1775e8c8d25310fa0cde1c06d86a9f667fd77a84fceeec70315eb3
z564dc7832a18bb5468514364a66b4c75390a26e23659cd01208caf6123b2b35abf936a81ccbc41
zd7d5dde35e45255af33e99909c909ba481faefa85e9201b9c2a08a28c7b1de8d03955463bbb682
z69201139ae262a2a2feff4451ae757560d875800ee5108949a264e42674f3f56a4d1bb25952061
z7d340a578d47f02860d985016e31c48ebdaa6f724a5bb53aba358fb12a6dd221b7a151055f72e2
z5d58a9d9f49e58b780137237f78406392817530191123ab5b274836be9ff04e16cd664cf265993
zd441723d0f8043f4bb3b34759b4858b8c3404a602ac43570138665f93965a7147695837b997216
z37d8f35f42c40443c8175b4239e203f60c8738bef4a9979df8d96023ec0510e59343dafbbd2bb4
z107d13bc2284221bbd2eaa4a25663efbed58423dbda5c3e5d7597a154ab55eba2e975995ce0d51
zf64efa9d504fb690df795016bec479f779e6fd62635336adffcb532621495782edfc9e20d24b23
z2f924053f8efb7d14e004bf1c070f573fee4c937b15982e2cf71a70e893486a8a0342cf2a3814b
z9315dc654ec555da26e3f11a434434f8ec7fd842e17e7be44daeb11eaa9fb9e81d4195477b3c90
z59663b6fd46d10bd7e636e4743ae9ef8d2b9651a7506a9ee4192210c9f0270661585aeca3dc1f2
z8c7bcfb891a3194c2e24c6caf579c8682fc82f0eb548b5befd2c169152d1ceeb9c9264ac252546
z63f479dc037c78582a81b4991b6a1d8f57f0ef4f16ec0600a61a2718de23801bdb9d2889a839a3
ze072fbe3d2548fcfa8004d8ff310aebb6b32ea2945cd87a367377527853a63a352c73e5e22a5fa
zd057f6c9b949fdd5881c10ce4990795e69bbfbdb939cdd440a4272fd821584b6c67d2be3c02154
z557422c4f56d55696673360000c9d7d44535624271af716486c522399866576d041d0f93864002
zad49b3c8cebb6728f5837ecbe20da39a428ee81b13b108912d9cd7ee2967001032f8f02417818f
za9ffb040efbc5c49fe1749a1bd26e758bc46b2f3479a650118ba4b88feb7e46faf4bdc6e26550f
zd49822ea1787e9403336fe022216fcf7bb3d0fb44d0237e19439b6055c1d820cb1760c1270725c
z19ff168d9ceab4897c67fece4ed25884926a697bb53b5fb54256e0888d0d40b6302a84123aa858
z666cb5eacc64aac6fe886db135d4f7b55b9807817ae07d35850dd4de98ba9b351749ceab8499d2
z2f8383ca304a0b44d9ca7fb5f2c663ec43d5beba941430b8e1466fe2843b1ee9b932cd3ca08335
z29239d7f9ec1316d52943412adcbc447ee52aa631a9b755cc577f33ca33bb4abc0ce553468e9b0
zb54a97d13a7c8486ce602e15eccff56d9f868a9dfdb0d6c18ebe9ef5c2e53ddad9b332be675c7a
zb06cd48d8becaff71bcd6577bcef8a853e6326ba9fd3a11055bbaa2ad9243b48f359ce9d34c00c
z4b64a06d160631aa9c0e9b1fa2e0d4b639ef61caaad85d5d1ffb156a8b6879501cc83bc4579d22
z2e6a4037b30859838dfcde0fa0768fe30fba8fb29cd22b13020f96c48c6c8f0e5b6f4f989cd197
zd1614d97352185112188cd5c1464c41e682df11d2f900b0f53c8bc638b2936fe88bbef5fbaa89b
z08c76deec3f44de3c5d10fa551df951932fb964abb1d3acf28e74c60a158624ec6ce7314ad087e
zefbb505c7b6052dab6eebb68a86a5eda220a0619a45a35787c97f013982041bbf253d503f11c76
z3e539030857ffe7cca1f1ec194953c528cbb92ec6f759c0698a6d4af4febf145873f8bfa78b532
z024694ba2fd6f28f0a43763de47fe269505c72518f0916bf5e640548f29b4aca93c0bc4b0d218b
zfffa769e231757d987fdb8831d23b6c6f22e0ccab81ec5ae171460af701b5bedf0beb99e0043f0
zfd04d724c3ec4abdadc52bb0f417e259fb2a192b898edab4db81e5ad1810f994e1d9990564aac4
z42281a6b8dde55c48a3e25fd75fb639fc632549ce02428a98f7a316dd4496a7e80e08fe597a931
z19de31e08a6200efa89873d5bfb2c697fb85ce8f34bede2634f35a86b56abb7deb39cdb7e3adda
zc77db85822fb2d7d60a4bf4ee9e17b663b6df6ba6fc21fbc1286f1e3c8424de3f643998fc598f1
z17217482bdde221c5c4b19a2ea01abbb1c423150ee4540846f5bff8e0f2a696384936ea6b03da0
z524995f4e7b1f8c67f7b47a56630172c2b265fa633eba725e811165ab5bf7d474ed13b5341206c
z085875abaae3f0b24dc89125b838ba3ea28377e3db399ce648394ca998ee174683e92c1676f08e
zd5ea8718337fe2eab44c7165bb5f2d41728edcbb20ceffd4d4a5a345f4bc5e753f2fb5e91030c4
z25503712cdc3e1b5cc1407b4ed69ce4f0910486017e5c6043d52858501608a28aef1350a096da3
zb94eff65303c6f90f6139c072c21a9f68f279a802ae621ec0ff53ecd460f4097bc9056dfd034d7
z45910289a2ac66710cfb35494e1b3dd6664f63b7093f7e4c5c1ab74e7c2aa41338c894d44ebc5c
z1cb409f44d45a6da3808318a81247eddee30116a0d400c241738f77baeeeab4750c351255116f0
z5e70f3e4df889bdb18b70fd94552115352c113485c82e50b6458a46c44b3653f276d8dcc316281
z195364345c1a6da40b490771774bc34a8495a64e9616929cc6829aa80d64178e2612836d3e1ed7
z6816352027efc6af0719f1147de1be651fc0e9937d3f0c22f8d3d930ba7f930570f6649dc59e3e
z7fcba956bc39381d74f7c3404f36b9da6e682f1f1b606e6540dd9ea66b0f203bb1345a140ce591
zbc02fd8295b15dbae3e0cced28eecb8daf772ec68c25bad4600902a29f54084c3b0146fc996126
zd3fbfbd470333a077444ed960d5b36d3afcbef3e9c22f177cc2b7e12e691dcb9921a8083afad5b
zdf173493aa120005739fdca6669a1874a65c15339675ea6d21ab0b9ee47642ea1d6d7a9553290a
z6eaf572ecd6407eb58ba83dd7e222702a0b8f4f1fc2c893c30baa0c95c378d813632718e71b664
z48e06c684eee16367570a3aac2f982d9f43d4e14f0f821f8e83d79973bf11c522d496d8cf04b41
z212d079a0dd4a39d1b8f48856a6e913748a347e8bbccf30e56c7e1dfc3eda9d56c0e7afdcd24dc
z82b148ca004be33f94dfd254bfdbafccef6d9b384d59abae8e01ba26200fb36b5e7e17f2f047f2
ze7bdddcee16d2cde574a1c9b5ac0daf42f423d674bb5c0aace6578c33e5322df16ff9da0ac421d
zcd761945597b43b5ee55f03bf70244f0469e5c98198a9a55fa2b3bcedd728c9353f6e03b59f2a7
za99327ddf4ceb30150a3253c22e4ab573ad05c8e49b231893a891b062ddd80db984a1a136cbf9d
zd85e93e75773541eba6ca497d0fa4e756807919e78e2279aba11c527a4219ff36ab925cced956c
zd68f6665943a279ee5f5dc845c77d882bd5f28ea3d601eb56fab5274544d9dc7a71b94e932cc21
zf28d6c5c64850feba294e6e57d0cb06af4d0a79007d0894a4edb4a6248465b77f3ed973b56ccdb
z8f2c3de5a30fac429c402aa6a7b4387dda2f1f5f58ab36260d8e453601846bf52bd52581c6edaa
zd95a303a6d8d677a4c97177476fe73df08cc6d340ad4e633dd636e21c8cbba85e1786fb6aa3d16
z0cb28858aa9ae7381e322c7b769a6c16b36c3cb9bb7400cc8292a607c2e3534c1f0c87f47e8ad6
z018ddcd5dba045dacbe861919978c2b870e03c04ad9662f6ee47390fc139ea790f9cd05b9bcd3e
z1580477e51e93d6590b7081b08d3e469c8d19eec96a658f5b1ee9b62f308b1368f06f70829e25b
z2bd0abbef4045448f013bf0d778130d1d90af040d29c5c58183dadc6e12d80912f066bcb90a408
zd2dbcfecaccfbaeb6aa3758ca3cce845c491636872c81734717bf2986cd3fb393066b42fd3c123
z21f6f8663201d0cf37432cb1d18f96f2f7364b5744b6d2a8a63f67f2854236fbf2c713cce91dff
z575d48bfe25a554abdd0cd836ca50a3fae086d58b829c45a601b4e9a237b65b0094d76b32be210
zc10c2f31f6d312587873030c4df29e1b60884b4df9d574d1fc6808a93ad199f1f028dd4e06513b
z2650ffdcbb7110ad554c04827b3e7d174a76eafdd24e7a0eddaf3b410a84ec6ab322d8d341b7c0
z1bbcf185c12b6cb9cb1101b09ca3e9a91d3a5cb51bbde9e4195c0aa9f2e80da5e02beb950118ae
zd8acf3d476685670ce230443e6d3a99f7ffbb62c554924d81fd430ad663fc747de0842b33299b7
z3a141a5c2c5228573ecf5a4ee2930d82dae0087f52be6e8d755432e1e8babc4660127908588afa
z7b2137a179fd22829e6f88423d0c5c8bfdb2b691d00a8de882dbb4a4d397dba58d63aece03719f
za7353859dda552c7c219100cc04f54eb8fbe897cb3f3efe9bca3974f078ea54a20eb995d87dae6
za831ef239e3ca5c19196144a00f59b73d870bfb2f0df6a8d02d785e92d91e2895b6135863d3e27
z58a93a9688071eec870592f5d3ba6578e1c87c1f8d1ac87d8787e38ff1fe4a998853c102798c9a
z5edf3f29645a74cd42bf5b684d5b1d5b682d14c08712a85b06d595c5e6a9db6bbbbdcd580644b4
z03e75f8d5016c89c50c42cd7244df7c6ecca504a317a20e889f8216a0ce5612b7bc2783cd5c2de
z285c6351ea845ab17f054933714b45c0616e84a3d5a367cecc3a5ecd3318ff20580de92b16949d
z288d3ed34f26f8eae616651eb26d0e4ef6994fec561a224516323692b69d20025db5a0075dffd4
z869fed363abc8f2e43532cf7d5402c6f6b72c98bae375a611ae9672012415e5477d8555b7cc6fd
z1e7e5025b7b6ae66ee425b518647865c34bbb43958ade8ca3b774681f1b568552bfaad929dfcd5
z773a8aa9e450f774a8f5186838977c3e72138a21b09763c7920b23db534901e1256d07c8273d18
zbef2be8bd1ae997ebf8f4bd911dcc606336cdf31c2d8ebd3bebbf30c295e07fed7c4f1a666ecbf
zdfd1354a0de9cbcb4afdefb62ce3e99ed2c2aa6bd1738467047661acd1212e66bb2f07f6109245
zb3f5468f97d761497280a9a43ca1f0d80d86a65534fb0eb15d9a66166485443d52122ff87a9a15
z91135e181b25f4968e202050d4b80c0be407ff48d1953b4ff17f8a72cd69d4e2b59b5d05b4f614
z458f48fb4ab28bfbce30e96665f5f9f7ac263ed813d1126fbb020916f39850e99c9bf30f8f2b4f
z4e1ff2b714ae7faf9f1a311a1b24d5cb8d03a39f6e49b8fa2d56a6a0b61c0cca2f3d2fc6e0ffc1
z3d1a110602325e8319b071a6ceb222225285e31e96437075354dfcd65dab02b94f69ee34ddc3a1
ze311ca0be68e8098bd191fb9b63d9fb2ca06b7eb2b9fbebf251ae203e60911c8d98e8715087439
z5a99b3be06868de760673979e8bce5fd1c082aa8924d891240a30c58d0d438f5726300338195e7
z77f98e3749a4540a37325b4ec040b11370137d2b15b454d499273280a01c5e9e31f01e057d41f2
zd4b3be0c5fbfd80022441ff6f0721b124a9cd7788cc057829af817f6e615b7ec5c30a358bb5f5b
za63c4083ed0c2831da83d04fcd0ba35c45cb4d8a1710428390b857bd461147f20f4fd7e6f5a08e
z8c6b5b5138fc136fd388618ec0acac45f68b8420e99d7d151e31aafd1224d075f7edd4d3537060
zadacbc5161f236a42a14022b94ee409f3a31fdee7fdf083ae30adfbfdc62d76a881e2f36a5455d
z80970ddb3772778aa1b85365f42d93db32dc8d65a841410608f5eb0e982b12b027129a45bbb289
z1b1dc987d86853fd5eccea8bbc81f6d31460d5b538f00991215eac4b35dc727003be0e0fa139cd
z7e417a016da7338d784f3449e1c000181277814c9b75d8739a3000f48d85e1f16036d65519f336
z16f293a1115cb84ed39342e09e24f16b99c7c18b9e937fe5cc41c9c5b7dee19772b30f0568770a
zdce3e24a861ad351768604e6fad6d53e672c23866f148c7900629df3e1d8017bec032b4139c6d2
z7d02faa119fb6fc3d01ff973950cdc31ee10b53704892640858022f2bf9ceb976d1beca1c28129
z75d29927db5f6fd0298c68eaf4d8d83890cfcdeec53bef54a8e1c9b33caba160c0bccbda987d17
ze72874844f45ae152efd0babade9f901e71c5c461b4b7b162a20ceb672d086938cf0688da2c164
za00ff72e325325f604b71dbf22e11cf780c221806b1b9deb7468e39d3ea80a3d48b372fc528f5f
zbf6fb2f15a04793237a9c4792fca682a3cf258ab2a5dfa87c474bb38ae8a4c6daeb83ce1a04bb0
z386ee7be298efe460e93b3b1aeb849ef2721b00c96b7084a20963ccc9711050fcaeeca252294e0
ze5979e0dfef48c1004cccecb4577b69aaef1d07b511f4f5bbdf0296e472e16b834700bf88492d1
z7ce95aed5bd9eb52d5076ece3fbcdf421f36d4e6c95977f233de33e88e39c6824c094eac4ea480
za171555e4f40d1fda91a3226d44d5221f697f754e18a107d9181a0c7db510a7c2b19022603c279
za970d20c1cd375bb8146e07130b1f7b4f778e95838dba5945985edc44277c83ced2febc2f43c8b
z5832e9a7ce389cf1960760c41cac14852e2f5bdb716397a32f117235e1353ecdde397949d206df
z2852fac5ba6c69a8a066b7d0085a8b151fcdb1816bc2a757bea9c0ecec68209ca29736d001c82c
z7c6e756703cccfa657ccc0d79ffe3de2e7b3250731273052e8824f8cd9ee5b30973cf1c1aefd43
zd4a3ae710d9ba883df6ff0e4f005e7ba33bc7397723e5fab4b614fd1b46bcbba0f482b165bc610
z7ca30a01ab0f2763b8cadc4d9292563aa8266d22fcf492d896efb58a4b9e98f9343042ab953c85
zfb3a829a66d25c7494ac856865cb2cc254e31347f0283c15e94a0af2f85b4c2740ee271213f185
zb2c0dbf7c69f14f687ae91f9a6746c1d03f0c9e627db7e9bfcb3fde2b020fda6b45143cbecada1
z09f67289c8725b2c55ee093f8c01a2d00b2c836b47f5f55e25240ddb6c0b4e4b4e6598700313a3
z9353d980316bfab9da0051a451a878ebba343c0759fab7b85b3fca1564106ee417c18d576d0362
z499bd6e90d10bd4e2b56185ad041a58dbe4c1b591db5440bfd931dba80a3d4e8bcc89b0d2b9772
zcd413a1a66f0bfdbe0a97c36a99779e580118ae5a032bd0ed43c45031d6ddd1fa05ec5a5e22fe5
z55767e86e5428ad9c1c58afb2eaada8fe1eede88933f563f64c3203c39146e0660616a3009d02c
z4f47f53a5020b3685affbae2e02d270b919719b7f8370dc60cc419089cb3a16e3fc01de9fb209e
z07d97b57446f45632bde87000fd333b393a236728613301b06577c6f349b306ddac94bf686efdc
z66babc4c4f45daec65687b2a88660ff85d25298441313747e101b46f4739c4261e7763a87e1d4b
zfd970294222576b239045abb0a314398411fc0b616e70284b76a69beec58c4c4d06d91e6483f80
z92febb54be8d99e35b2703907238c647801224e00f28a078468180a160a1ca0a4c637792742c14
z30ab992eeaac032522034db675138bc608f02bbec612ab65afe15f533790062c6d0d11ed7e8fe3
zb8dc95379bc0043398b81bf93ac65876dec03bbdf9141a281087fd97121d77b784bb18523011d0
z2798c3790b9dee2a27df41aca3b558d137b11a880147fba5fe54256bb9c69a86324f2a0d0ec268
zbb39c868467b1eb610bc841a28c0436a9c39d79390541a4527a8cc992af7034c8fb127041dd91e
z799849f018a2a465b1868ffa0610336b1d974777180c03bfdd7f8975fde0e8ca163a40abe48b16
zaad809ff22236907c8991cfde486f90035dfe754a136f86c7e0b89d4c07d7c841acab6eb6ae4c4
z737046b66603a4cb85271c4e17e42dc1be26e4704510ad33424282bf451483464c204da2618ffa
z647d5f66c21fd5c663e704f0ccc8f844d49b5d8dd0e26bf71b9f1739b80482737d3379d36496a7
z015a55286752245e5e5c6ef988cd9913de1fc50708bfe4fa1333cc41e2cf4a45d671fa9e4d1ea9
zfce2817a78a8452a0ef4fc9bef791f82444af02d80cbcc1c3272e7a498a7b05a6856e912b3faac
z20033d887d6f461c1d4573460f17708d28c470685dfed780b58f91340e7fd8ff144979f5c8f80d
z4efc5749ad9970b758eb74bec2f8cd8823317b099d6c34158d1e4d79b3b04f21ff4eccff61b28a
z2378bd7398338492726cfb3139b08e9a567c4ef96c9cd652d931d1f8edf8ba796673a6511e79a0
zb13ec5e523ded1daf8ae32983eb2ee57bfd33fa8669aad94e55e648bbf0f2ce0fe6bd3ce817c69
z06dda66d04be0e8f619f3206c129b58ebfb51fc5f4160318bc7567056f53f710311b15f6fc53ff
z71b94c3b940bf01a340dcfb924b2e649cc16365adc1dc0f386ce4f00f1f24278181e97547c8ff9
z3d6e96ea10a8aec6e94d2663e2ce2325f147f369488eb7a8c3d54cda4267e3ddea903e9f082527
zc3aa7460718f10c1a2dac109065b6c0e07e5e70f3e55ff68c943ea5c262ed85eb3137958ce0c32
zaeacc6de83c2e5f6bd5ff726dab8a5af96d2a9dd84663db68e636eb2c52622a56e74ad8bb165d3
z2d23046a9c4c5c50fd3836b7a8e376ecf230def78ad8fe8fd787ead7c1a579f9490e2d7351f3da
z235159ae2faceba68145725c36be6c08bcd855e576697f8032068b69bffc0ae9e372d207c007a3
zc24cf5df5da698fabe6cdbc025aba6ca5a93627978b01e43d4063ac3c0f95deee22272bd10e51d
zf8137d3d81ab2d9d20a0b36673f12ae020075407bc680ef00a37d7f4626163914c7e9fcb3e9a13
z72a09190b82c0f3d661301fb6e657a525abee5b3278ca4fc428b2a904e6ccfdb0873c1a400207b
ze5d83a333550b77f5f1b86e194c65fe96851c1f51a799ff03a9e35fb1fd4519a27c963c2511472
zaeab54f12cd06c83c86977ec558b4376bb0d79833790e54a5693a671a59c38916790e4c7297c13
zbc0a5275346032ee4f9080c6286d2c8ee68e0f1596ad314ceefd1a7a85fb607336f776c6a1c790
z337db1157df4f3cea1c34b6c26c44b61af46dcb1e99876fa024fd65b235bbfbbcf51fb1956fcea
ze7208229f21086724021be3b483a8ad1f1e4da963fb8cbeb4e734f141f0c8fc17c385b5112eed1
z686503c668b881bd3a297b73934eadc6eebd9592f360a555ec2ee18a5309ff7d4bd73695880c09
z18f74009b8dd19561e842fcb02baf96930576830de8d31bdf1f6f6d5d170e391b9377af4edac67
zfd2e947e254feab0433f5bd852bb1ad579775bb06a489158738773c371d4383eae4799429ddaf3
z6594a312c56765a3f3a6c8d4435d150fd54e2c93594730722e8b14939d1f470346db0c9dc4f414
z3ebf4d4bf64e460d107209cf5e9c500d49f401999ce0bd1c5ae11df9f6ed744bb9e4b479a5cf3e
z67d7aca36ccedb3f3d6353244861c39705ba1c5e730e027f697a0058c414805f419687d7032406
z8466812b4c5121f65c7bfafc95edd155efd5bbbf5da9a0639a1beb49852a4512a85275b1f73d52
z05f32be708e94da186d1e8e5987dbd2f830284fd205b8fdf9b54057b5efa394a3c635e1b404217
z831e2b72ee85fc36c9258a72349e98bc76bd62e0700289e0d41cdf059416cee58299f080f1251e
z2b77376ef31ad9aafdd9e61c3723ec9394f86ee65916aefaba22012fbb0c80fbf51142bf4aa9e7
z9bdce87e21976166b56d3a76e3ea75e1149efa2185a4c747b5fea0663ed73aa8cfd7934cbe0f3b
zdf7712ab2f44ce5883eac7edcab03f3ca324497e33b3d2729d532c9f7ba6df784b58b08093d7ae
z0369ece1213f4cda1726261283bd26d5fe64badea78b92f5064715d7eedb9187b0cf0a753998e3
zc8fdf444d9d7a8a209c13ae0eaf58314f31d9202874e8caeb65850f112f478f6545832c7877ed2
za02b0201450ee792cc84d9a2b8c464eeb77fa0ca3db844d26120415cbba9669790fff17126bcc7
z4403b99ac0b6dfbe57acc994d6763e6098b91ad53818721affe5e92f7fb2b043622037961c2e49
zada4c17cb61908571896914fd63bac0246fb77462ce614d5a56af89859462537f42382d26a5be9
z3e8448164d8e8e1040890271cc836b3c899ea919ad9d4e1c1b0eb6861b7ab9c6d1a62a50165e6c
z607fbb12f32a026939a645bac1df073fa07e7cefe05dfc1def1b318d937e7b2bee79ff83d85c09
z8d9d54098c4007e851920ac09ded36c181081ad73cb52737d6a73c79148a01a3cdf19665d704de
z8b407362a94a7837dcf8df6a4acda2ce6624d162f1dac72dd8389585a0649904bf2bceb73174cd
z7d595fd60399bb3619f0c0ad32ef27fa4b9a3c7a4964a0be6139bf0078bd96423d8b7f22e2cfd0
z24bdfc01838f7a237c0c66f3778c2a1944eeed800cdd73e6198b714b30f2dd4ba91c84a308dda4
z6e571bf86a54e8c95774a53033caba34e704559dbbead369caaf66980f6bcaca2b97fa2655b832
z92e09ba1a578909b997f9634bae9230f203205c947a72c5fb70b3affa62e4f579aa0ba3eaf981d
z50078dd6bda496a470f6d3df434bdc5391ccb54cf0c417998ad472cf8f3d1aa413b45092557477
z99865628fc4807ebf2562adeaa6911fa7edd6678086ee2c0f42e556abe648c1092cedbf7ceadfb
zda93302cac1606acc4d3d041dfec851423219e18c06199a92b6bb5df3058527b6ddf2518a815f0
z518fc8673cfab8cee9aa8b37c76a9e3f85a1f88fe59de3484f827ec42d9de5ae9ebd4651b3fbce
z14b13a52f953693f1f424fe0c96e72da43892326d15658f80323f4edc33704bb61642ae14b6ade
zcc2ac8d2f39c11ade03d22db76f12cfe408f7c3df9a19f1d6ba64d23ef8eaf753ca7d41199e754
za3a6620c8a73654755bda09c37c8c08b9ae5919fdf588c10e79d474ac3a066a2c8037b58acc6dd
z778ba582b37b6f0ef3dab2ed06f160025a5251c0b78905fcc29c01575e62412e802642a823bf2f
z3a03a78b97151ee8ac52923d3c5ded3a68493308b9c4aba8a4cb7c282a27706269056cbb80ef2c
z8c57d4261aa2ec3519cb45c19875bd420d7ba2c7f6a766a23f9c92dd93b441e3b63c16e89dcc9e
zcb554d5ed04e35222cfb78de290162e9886ed83368fdf4929fedba7b3d59e9859fffb0bbc47321
zbaca7f5a3afbcace52ce55a218ea8b7838be3608a69d865d0db2ddccb31a4dc220a578e3fd2dc3
z93521b4110487f52b9da3bdc75a019abd402a8f1e79fbc83576bb7ce68b8b2f74aacfcac154e7c
zd3b6f21768b6e2f16965ff2c050e73315d7a83d641126861bf8e4ba7b5a0d6714c592f996b4f22
zab957113f86a5b633b8d23891cde73d7afcf511ab1d3ce6cbf7ffb98a16b90e3ba9ae179492e52
ze49a501fd7befcf642e7d0b365614ff3eff27afe01328c107c0f223db89ae8e35542755f7dbc46
z4b6f783d4c87f08df3d69758ef96eb2fdbef2b7a22e8e2358c9f3424f3b88ceaaf54dd80733a5a
z8d53fbdebab22cb72b096d6577172dad96b35712eeb6f43046a60810fb911be7c47b3b0473bd58
z027fc52ee8b3a32bb304644c83cfae65dccf70f77079523e2797f78b9db060c9cf65b22143a863
z07d4ed81f6b5a769db1fa0c89a6bc040c203026b030517ff1616094b8afa7d95a4b0245ea6efc1
z10135b9b8ef787925c2c5f9197a639c272fb1ed0fefc4b5a6d81e9840a6d5bf5f90d96eb4307dc
zdb174c6fe07621824685d81f5b8def02bb98723c71282acb60f9136aa81f721ae0fe809e5a8701
z49402bcbf6c592195d67a5a48eef11563e0976a5a3d4f629dd12957692bcca256ff1a11a0d9da1
zc11900df0876696f7dfc00170a32022c328c77578f703de05e83bb4296d48c00a344bf929a9a24
z541f7098275bb3267d955ac7e98d1b019f9b016633a147e58e8202a402a299fe763505f02bd419
z13aa48880b9e4df335bbaa3845d3acf438308e630059567a5e79848d827f03601c166db1cae054
ze4bcd3ee597350b4d6f353fedfcb5447b78865ac0e924cdec3a2ab9f1e375a6c1662d4c1c05b3c
z57c01b961ba533474ee733c2b3146b61d818ab04a622f70ed749a6f6f9ef490687b8883c8f9c2c
z42b380054194271eb6bd232ed0a647da66d66e88ef2cfdf1ee3d1ef4ff2c7bbeb2fedbf619b924
z6fa84dd4f4dc0747c5df33f09e41c7e01aab94d12f0e74637cb48435bacd6db67a417574dccd1c
z3ca58f5d7ee67ec19fe17671ffd2e32fbfa47d1ef4d6454e74d3641f17bae6b55d1a6f35f08110
z6d2f416583760a8c98e923fd1d70f3c52a395396020afa1249320d00c0be949af768f7220c08c7
zf3a08ba1348b2bad7fc8b0d059d8d03b63fb99a3d4fd5872effbdc0f8fbc9e4f8bf0aa6917d7fe
z9e7d06bc099639a1da25dad5ff92725a235b2cd4425cc50265eae218f91c43867d8211e3de9d02
zb69a6ffc5871bcd831a8e8f224c0e6878ace36401567049e9b6c872b2212aa101e27d571d8d195
z1564755962ca7d8598a070349c82718627e8220a2c753c63d9f994679065a7eaa6a24e38acd767
z4da59365d300eed06515d80e7cb7d02a07f1221a23a4ac84ddf52412b8fb53817aec46f48713e0
z516c82595921f14f8979fb50d2448c509309f1f88537b774eb2fdb7841b7da5a19835984192944
z267152f573a508882817de6e82210982e5c45047229bce69117893a0e7f7e88919ae9fd4d3189c
z865620a190851c3cba14853247d094309b0d5d04aad6d471d24f6459dd46866cb88fa449373584
z41f5a8aba0c7ce498f731399a15688c3a01ba023d0c0315ed91adc034a61ebe21db361fe1e5490
z7a11c0fbf86122fc5aba59ea228a7f178f0855d34dc22cd7cc474b307c399f3e00534818b677a7
zc1fa96984c2c3118d7877917d117853b7d841884af5f380ce183b98f72500b6a4aa9cad1bcae76
z50f2410ba0d1b73d75a8d04c910751eaa1b0b0b675f831c0b6a3b1dacc835d116a5eea55033e05
zd059ff2871bbd25a964d6cc8bae812db3b1e6cbd2718777dea508f5d6aae8cafaf4fb2f6e17c43
z6556b4a6cc55d35376776ecb6987da6b3e3ecbb8b7f03546ff8325f63df7a165f0297eb15c2462
zf82d8e841afc7c97e48c2d8971773cde2ee6261867fa2dac9a6395229fed7c73e798b3007193cb
za4d6a52f61359c6a3dbf34ce7f1887df6be29b37a6a2cec8656fb4d13cc7adbd4b6fab207e660f
za56ba51812bc891e569dc75fecc401dacedcc57369ffb64973d4a0e4bc5f0fa75b3a1c80ac0921
z9ef0e247735e7055ed6751a7c5def1bc45b28b7b637d3de511db3ae557894fdc0f8374b9063d78
z6f7a961eb317a0f13d51b7ac46d40e52fa3710e534131719b0a8f5099c1f9fb404711003401115
z4d7e34e60ddd4013ef38eaec44b1457b3bf5f4da60a3086bd0ce3ef64b332f1de54dd8fd585581
z269727504d3f9aef1ef2884d4ec1aa3cfe2d0b4c6ff11db48a03767a340ef2ce241642444f3200
z0e5beb1e23ad39c9b13fd644719a583c1551c4e43750fd9e7ac1f31db44ccfde9ff656d6d74d43
zad52254628362c7942b49f746b66c8a719b1a01974e444683e74b649dc15356782056c50e383c3
z7f1d9a2eca681eefd9d27d77e65e007a12ba90709023673aef6534d6afe152739f4209f25bb0bf
z581c0255950c9c02ecf05ad4620142948a7e35584e40d8ae7c34d0170c80a9f4ac65b1155c82c5
zf3abeb1dd31646b6a9b49c2e39995cb813c5ec7aacda2b7fa2aeb9a20d02d04259e8ff25e5778b
zd27844e64e08599a5d8f4dfec3bfe5841739a1e934887d841ecdf4987e4954dc7c067bb733385d
z8dcc79054a655a062043e4fa3d5fd27c0315d4efee3fa1fc88b30df3826988ca6d0e51d8b1b559
zf08c313065f22222ed2a70873434e12669b540e554bd58e868f34b2e0064082203a67916475f20
zb0e6ef0811942500cef36c8e4c9abee036557dad98ffe15e07af2ae92957924821ec7c88d66724
z0bf9f4196cbe5a9f42ac696b83ef3696fe746ea7bb8c9391f36c7f48bdfaee5ff58edca5f9f2e0
z35c2892c8bf57990f9f8944d139f7bb2b7b2e6c9e9f49cc575a80046f8d45fc4c27357e0166c53
z9d6424fc8800650ae0187a92c1be5cf389a3eb8de795a6285007acc2bb4e48dfebf49e3fa1dae6
z3604ec3de540f5c14e8f4631c4cbe3978c93f84ffacd5bbaedf1864710a022161da27b40aea0af
ze2f81097325ed5378f8b63a63f8220a2c8edbd6b0f2f9772f136835955ea0998ac8e26463b02aa
z1a427888bd326af7e2b467f1eb3a67bd32b2cb94eb529a13f0ab562d0008ab9557af311f1b7779
z5269db3fbb694441016f6dc6cda2e0c9406889e9e847dcdc9d8fb963ca51e3988eb4c92a364cd3
zdc776f9bfc3ff783100423116613a4cfa55ed0545779ed2471f8f3299740e90cbd941a01366b08
z947ee2152890a3a83ed03b6b235bdaa115612021ffadc23925fe12d075f2e6da186302df743681
zace612504c60b27a49c7e6b0b96b14b634f9decfc65b7ef9286ce8d1f10728c64eea31f8373b6a
zb63b0adb92cd7914a217012555ecfcc9d7f5015a128fdadfab9f0bf6f28eb820416ab5aeb38f95
zee4f7f9dea062697393d182a0d5cbb1d978d1bea2cb6a4a536d192fe1ae808825661d22bcf8073
z4812d082801097cec611822c27c3a3ea8cb94e4048f62f8fdc9d3561ae0db2e1d23b723dbff2da
z2a0610a9a804e179ef71514969428552224e8dc4968e888ae48299a29bae7be28775b4b88b156e
zaa4585120ad21935fa1d80f58663c63205458d2a8b15c565858a536a4d8bf05f397576982abcb9
zab23aaa5700491739484d34d7b211a5ae8617453562f5534644d42dfd71fd441f7cb6a15bd9ec2
zc700b25523ef470a3140e3f4ceaa350c4a2b615150d9fd5b87510011d8b2834862e0f843e4db3e
z8ab3c5b826c78bfd5a69f007f7dfda872b679c8530b5778df1f637051e455d42b88f3eb33d1744
z16ea96de4273bd3eced67e135dc85a10926a8f35554a4edd2c59a5a0432b7eccf760c07f330428
z604d154322cbfaf4a96be58933730097c1c4442e9c0de937023c37a7d2e5785fcf90ed62bcbfe1
z837853b9120cc8329579a193bacd3bdadb327dd89d7caff7e0e59027d9042ef85bf0a782ef3f58
z553d8045a25e73877f9dd5edb52e07a9a05e53d75b2db80fe7d5bc99070b65756230c6ccab4321
zbbd294588d6cfad8196c29f01f45dd8ba797776f909891a4444d4226b7bc3c110a2f1746e8bd06
z430c43ff54045ab24110d252ac64e85e027d545349a0b9e5a97220e2ce6dcba8c7a27890125604
zacaffd437696d33d8d881b0aa10d8568bc6e82d026505a4b0d3b2e4a8e5f5ea8e4eeddfca05ec5
zbbc90478f8b2d6856027822ab16aebe89b9a4a758bdef7312364b406bf99fe1b0b5d583f2a95b0
z4259276c13f1954f16bc56e08cc798116c3546a9bacaf183fbd81a5cc8a64b4bc67e915a3e387f
z1e2a8c8e0b134be0d2fd41fd1f32fea70f483ee7482173d8c2eb6f07dc34adf2d3dc5afb789012
z5b5130514f20b30d5fdfb8da5af66b5032f2ea0e15314a2d6c763eedcc438073a626eea36f07aa
z606a9c523cdc93b359717d4458e6c4a2c348502751143259c4d52e02e5fd38abe8849443dbf979
z5d8b2955eb6a0ba3dc285318bb3521f0e16cda92b452547c4f75c8f9fd94e9892007390e4a21a5
zc93a78e2a9a34e076af063fa2d1b0661a007693c3e0e01e0147f37cdfd677b271908fe8d668a08
z42e60e2bff8f8f16df96396ed39de5acb1f3a509d8431ae308e19eaffd8e021789e589d4fc660d
zd99af085c5f1f9f31f83bed3aef95f2ea052bf8dc53f77f89ccb5005fb762f2c031e2a71bd6161
z9acc987d4205642b2089e6d73934306332528df0ef3beeef1564eb73734956f0df5db1bf447079
zcbf705cb704273fe4cde1117bfe987357347ec057bf283c5ae940d536a9814c548cb81ce844ddb
zd2423d24eefa5f6454958d33ede0850251cadc90447157d29a53469e2d8d1ba8472dbfc54c7ae4
z73873b13d15d4b922a606eadfd8d03a192e5d8861154f9c6086b10e10369c5cc233c2b87ba0932
z78f35840f419ed59ea4e56254556f80aa37bacb8412cfa5f6fcf72e66137f89310e3a7a4ffaaed
zb1580b83521813465d457a058e1834acad8ffcfdeb2338500bea339c2ecda02c49f3f9126b2b43
z9573e58c31132214d307dfbb9cb53603151ed9ee867e8e933640cc6be8ce5c7fd882aafba0b087
zbc9030f48aeb949a4bdc2d629050e67757d1f936c2ad3d467ef620d5169f931d22531f3e1c9cab
za3e64d0da1854acac3c95b396a68b738d751191deb1dd56132ffc73860b657d5c4bbb8fb6d12f2
z571517b33db59230c7f2d5aeb0e25cbc5b51eca6cfbd4f3e55af7e1acd962fdfb31f52dcdf9dc8
za311958972fdebd928865a405898d852611f4a874abb7bfdb9ed096b60435faf1c0159e8a118fc
z0795421a5b588687dd781dd3e1fd78e090acf05cc43c485f5d107001cc68340a0bfbe8e1f92aee
z7276aea5a265da8cf27dba9c4c8a32c7066b95674e6afc3ae0101224a54d04eca7c37886a4fc1b
z46c290d0f24e7667523973e19c0e02039d228d39dced47aeea61d593565a35745619ca6343a68b
z690997bb6b37fd730d174a4e15ad47a05f832564efdb00f013f89f1261eefa00da106ff2f9e631
z6b5bc6450d16d846d69cd8a4f85a159cd9a145a23926ed5b25738bb402c7fe28de8c08d1a1f2e4
zb5cc6d49fcfb049f05a93b5a0192aa3f5343b2ecd06c8a90f2ed983e4bcab1116967906d0c9e70
zd790bdfb1ca952c192293d6f40a048ce99d656829407136011c9a588edf94a9b921b15a7193410
z4322d04367dfb5f4d43d2596b25dbf5e35cd5df1fc7f30456e970bbf48d932f648b625dd081529
z1489c5c6d684a3217262c0dd8f3c20c618a671a20c72a5a17f12c3f6d217e97da5ecfbfa7e618e
z58e0c009a568a3b19e0673afeae6ebe16866e32ad7031a23e1083ac5a13ede9242861730a8d380
za55d67d16c23f126f5df52e5967a31074504aa298eba057a32bc4eb8cb7d3e3486471b37d499ab
z6488c67de3d0f78a426a05e35bdfee9c321859ea5319d7da47ceafb06055ee99b9ad4d18783fbe
za1e2c8dbc6d607d7bc477241c5822828e76cd0243a098f1f83df2dd4edc0921fb675a3fc921444
z0fe31694213dabe0e05437702e4c19e48f54c88f7073c6d3882181694d3ab0912a090978af5a09
z83d60e7ef2179b95ce4b34da223b3ae344911876377d4d6039dec16431d81088959fc9641fa3de
z1abf7a846603fd15ea15eb1ac7305559c197ed778835c760dd0a6eba47de6a0f772fdbb6716886
z979890ea24885be57a87d93b4f69324f3f206e5a694bff512394f9ca6ca6578c050f49e8827d5f
zcc0bc038166eab351686a63613df64459d9cab552f1c584b62a666868607db002c7986d7ea8f3f
zcd0b46b2564ecb9f9cde757426d96898c638f8eae052826ae9ef0bc314e122d4fc0213728acbeb
ze0c3c5eba7328dfd3eca7d0d82daf22c96acb4da25c4c5bf297fc58c74ee8d7061b17d0d14adb0
zec085194262b642debb6a6ca7bb812977c10ee50c8acb7b3eba581d43d77dc3903990836eafc76
z00c739a2c26320d59e0768c26d1cef91336f1aad3efc31277eb45fbfe506c3eeb5bfb512b7b04f
zb18c9e60f0fd85725f88edd6dc6f8cd8d4a5b0632734862546d0f38dbbab49270fd6f03e74acae
zec22e5ea498a885e4d0b6a5ebc97e51de0ddc4076b2fbe85ba5a2f5fc1688eb0c4542305a49e0e
z3d79088ec0e6b0f53e7894d4537eaf097812f5aa4e404edacb9cef78a567896533160fbd8dae73
z06cdc2c0196034438c1db8157fa63f838691f756b38a02a88ec65be9b4c3dfec2bd5080721e778
z893fcc04425ec7198741bae91f7b84979e6e03260acecfccc6c8f68c692d99972574c9be39b70f
zfdfecad1795f91726a2643cdfd189aae6de4b93d90cb91ed9955f665b34f47ce5768616b4a9721
zb31de450f7f0a890fb873a2e3099d790e79dea69f83dd9d69a95f1ca078e89b18b6b1bff283767
za4a14875937f19cd9c7ca5b3a27ffdfbf7bccff95f61c6eb8a509e2d94f42c9851fff52d4a1248
z906a1e8da8fe0e48da7810b2b24272097887e1806727635347dfda3fe39d29a9e1e65086807104
z4daaaea933ea8d0aa164a6bca9ca18bd266bebb05e9396ddfcba43c82dada0390dbe6100fcff8c
z95ddbab368fda68eff5f4af0a311c54addc3e77fda416ac42a8f0472ef86fa5d392dc0a78f6126
za6e169c409b44af802ee9ba5cfb55fe8091edd20c1318637710296207b5d3e8ce8a2de971a8424
z603355fd8241969574c3d15ba7d523f027513ccb6d56cabb9b23a77b0cf886be5604c4d26bfa8e
z3b5b16fbd2e52ba36b656454efbfd72393bfdc87a903a9abc6389e6adbe27fe6b34a1096eb71c1
zef104adfbd3207d056756ebc95f38b24139b4d0b382fac645c8fbdbc84829b35d6e4aab6d8b0e7
zaa7f3f61c880ff195e3d9c785f0239c3532e5a06c4bf3778a58493cb3d75bbc7d32700d8c5e52d
zb017b17f0f8287be9fa41382933c0751550b6d42d91d29aa6488ec8d8cb8e892dea12f498e9ef4
z3538512a72e49efd5191648b7d6f6f020f8be78c0096fc45d1eb09f1a7eb9f7278e7d6a6d7e525
zee53e2323a13cd3a529c48e8a9a706b75d8bae4cfab6c598e00014e5a3e2c4ff50474ac5945b95
z182f91573f08f004c18bae73760bfbd66f8b7af3c0b18ddea16da1caceaea00fb8299e94a98ad4
z3d6e68f2f9906dd6c1d3b4b5d256f5742f33135af737a99f2ae3c08c9801aa3e8a7ae06c1703f2
z84ffe94e76b53565109e00734c695a72e9b3d6db80d10cf6ae33e4189c0fbb0de60e7e06fcf71a
z2e4ca2f9a6e60e1c6785dc7b7e158f6836a00961677328c868c7aae1e618fcabe2b1c3a91e89dc
z238ac7ba974ee7fca0f3fb863b63339a78523397eadd40dd36b14d9279c239c5e096b4098eef72
z46caf8d441cf19a6b82f8d6a3a5213a570ed24190d6dba7f8d4a6c0f1fb8a30f3b5856514c2af1
z812b9b77ef06806a0d15341c03f5edb0b95293b2ad3464da219517af1ec102d191c4dd349af47a
z4044a394e1807b800b35e968bf36991549dc79360b860da275fbd9a98bc2eadaa01285ceeeee31
z2ff547c8b08d13383d42b46a5b6525c77c2862a8ee2c53c6aeb298ac9f3332ec2668e8ab6c3a67
z567c0b82794d2b25ef2a128f94803ffd068c794be5741c5edd2fb63764f448183e2d6c6e4d064e
z8cf1cab359bddd697d1ee343575c5a73485e09e4e00cbd2ce053fdec0ec0c77be02ad319db3ae4
z03b7c45e51a90cfb01e1c822f95f7afad1ec227ccdab043844759eccaa9439fbe8824b2ed7de99
za0145a49f180d4ca4d12c1c5b17c971be10852402a12bee8cf2aac2eb203f9f9c46de7b24b1d60
z460f7068b407bf206a577dad88dffbf30b15276f83d38e0e0df97ac0d74e9f69576dc619ca8f4d
z0ff9ee0cae2b32dc67210f641b70f8a1b7f663bf543245362965c415c1bede4fae3fae9dc7233b
z95e0e9d7a1bd59797d7f33eb9a5212592b87587b765cb4df560e9de42c024970f1480e837cc091
z787144283a8eff2636be3c098e7927a7e96eff04a79b7aa821388a44e8f46530a810663ecd3ce6
zaa6bbc7357c5d781b79d66cf607103c8924571287723268dd1801aeb66bc3dd611d94f5344c932
z669c8f5338012b1c6da6312f6219d52597778995c0e9dc3cc79b88e2cd7c898d222b9d685d120e
z6f914ee1ddcf9fc442eeeca2e67cd312b06e55923923496b3752fddd51a2fb83a0d7de9552f276
ze8c2b4b52549e656741a7432d0379ce6008c2c0b45476ac9bcaf8e984f1d3134820c2ca5861cdf
zfbdbc31abecbef7c73f5361de6a735b962aa340bd07959f3cd8c750816ec373796dd5931e5b633
z80d8b270b98931875b776a9ec700eb56e200c7c80afbbc5b317f1d77b0bb7ee3219e0692953bbf
z1a4b103b4e071d8763c7ea4bd0ea6222b5805de491f9429f80f2481c684b6f7e1295a056c432ef
z0af1ed57da3466d706d11527488fd1df977cab0e48d204441729b5fb0a633c18bf9fc3f53dc990
zc44a1c2340a778b2ce047d7c94af5580272e1a33e7e0f1ccfafda71c7eb2be17e70e1471e10c7d
z36e94c635ed5269f9725bb4db4706d2be2ae6d319cae7ab8a7676452782a46544de4aa7adf0fb3
zcfbfd1e8305ef38936aaee6bf946972cf9498e04fbd4baccf2005fe5ddf3ec884285d68a893be2
z1de2ed71af4983f8731222c8277b3f64ec1d63bf7ca527607e785c2413008cf21de72a38c4dc24
z50f1e500519e650edf1f21fa133fe5c6842d419d23c58c174bf504f245cfed57812f3c8897e82c
z9dad15b2b53331eaa056f870e8b65d9133e8031424706aa7bd06e0b405631f7eee1d566fca35b6
za74897947469a894b0e5ac132402f86438914255889be30ebc69d94bce9121fa9800a092e6af3a
zbd79d358f1d17635cc5e45606b13dba3aad2696ae8c1a14e0d1530f00a44545c92ddf07cd22a64
ze530bdd82b36630034c495bbbf8071d6cde38fa7b171bccc2815905172a44322c05102e72bbe4f
zd260c873574f1674218e80ca985e46c51c55285380abcdf91ca8daf0afeb40727102013dee0f36
z9d76afdd151ddd03ace1dca63c2887699b50f8f466d81f81848ed195468e58032c1fc0f2e4f80f
za08f18abc208e469340ceb8460cbf58ddb3367770ba861acb13f2a94964525ff4779265807f869
z63554971b86ffbd1545ccd82690a1b24cf100dd6bc450d5a14adc05944efac4e7ca80529401c09
zacffbb8b53d13cf81e509085eeab132d0e3077ca9214a55b0a724ee07a9616ac0f6f504fb62e64
z0769086108f2a1e0c6de95fa9e123fdd00ca53a74eea302b540f0132f0f4221c55feef7124ee56
z88539f00fc884683ee3f8f6cb218144e6f1228162f5d63fc5a5faf01fad8cf7b178c99853fa39b
zb757157d3f9046fe0920a18107b6074f42146ad98166c8da83488f0baf87d39c9c7abef36a3deb
z1fbc64660116bbaa2857c87d21845551b4d628aeab89ec5209d6281a18fbdb752c701d2d3fd906
z2e2ad8298c43b68ac2a9f984eafa68c2beeb8e175f0b8d6579c60552f536db5dd9c1d10253e83f
z56f9b09436c00d5c6e31e92c6fcdabd3f6a98d7378b013f43c80219a64e8851fb40c34a6a08124
zdf71de0e17218efa5154b06317b9d85621c739154717966bbf1a7e4d74d7f994f6294f7b94a1e2
z0035cab14e7d8e7663dac466b661e216963f5e361f722f4df91ccd982ca1ce1b0d221478323551
zdd79221e833a0c7f8bceeb0b9b7716fbe0437c5da79c03934e4c1033e017d76a2e9b1a84014eb3
zf506fab29183696a53a26812f1235c9e68c71798c5f3d3452bd18b1edfd9aa17a25c3d5e212c39
z8e2ef21c0405d632a2c517affcff973bea1ef5cd0803c6ab55663e9aa3c0d2e2b2694898f03130
z0a89601a1d0ebee0fbdf1e0a24a0fdef398ce56c54c0a844104417c7d8a371f4e25c8dd1422e07
zaf0ddd78b90dc1fa994f04c9b9eb9536e58fcab0c224e0ae0f06dc129bb78300e9d29e0d9493b2
zf36a1e49b07f01e8a393ddc7dcd9598c93fd846cf4422beb81482847ac994b22bd3337d1e2f837
zcf490b28e09236be263a59ed382d25295f610c1bd9149ef5cca1c5fe19b69c3118d96912a65331
z705b8cc7061859897dd7e03a6f59ea1d6ec9b400878400416e8c9450cf99f6e7315bb3340f4d6c
zd14403a33d2c30e3ab9f630fdc79b66ab24a64e866d77502869a9c3592580a1f83f74b8d56fbb9
z97f2603a469d8dd260d3b84f270209423f058698376e9589e15d6adafaf54b41bd4140328c1b5c
zdff97ab04779addc645fcde1611d2ac0299c03933aa843fa5f76300e84fd73cac6758eed40f40f
z46c66f9f90e4ec57b36473d1c0b5d4c8a0d9fd0c386c738a1cb865bbfd70f88971d122241a2b64
z5e7e867bc0faad2ff68c0f1147a2520c7a2dec0929c71242445e6d44f1eedb5d92053c129ee570
z8967c88823763ed48b3442648cbfdc68acfa42ab1ba131e5c96d4e13ba5fcce1c9ddf7fdebe6bc
zc2a87c8f5c54a2278c707d3344d2ac4958380c6bb6fe6ac2e1fc43c012190c5b12b7c6ee3d55b4
z36a8786e62057a81aa492dd074a88e0bca889ec13feeea0926d016504de9587230c0ae49c086f9
za9eeb355eeb2f56e80bdde66549038cadee76e8d6735e74b9cf941faa6550e9f654f05ed0d9b5c
z149b3d1c9259955e2f03e76ba866753581b36b848f56cc7888d921777b798b97c5c0a37cc614c5
z5d31426dc1cc5abfbb1815c444125ecd7d112b52afdda30d6f0d30681f697cbab7ab959ff38576
z5451ba5a3e90c60aa4988dbe327d0e1440628b015d87b5e148fc1171646d1eae3e6d48b1e44739
z4be917c2903a00db865adea0edb0c96c85a3aff642879187f08c7729298ebf3f5a14a2220bfe52
z1ae460529a876e376c5117939b5275d7772e0528e8da2ec586e793e7ea87d1b58458af00b63b13
z48db6d57061fe1febe5160f55becf9516bf4483fb899ffbacfabeb74bd15117309cd8d40c42355
ze5e89590cf72d1a77773805b4c76e42e0712021887784d27342076b397afe2bcbede692447bc8d
z197fdf60b6ae7c1d6b9515db038540e803988fdee70a2a89eec872906cbefa310f68805fcde72c
z72ca8a6fc5bf384a766d83136ad84a05507112c45a313ed80e4b459e4588f405a99f12862ec0f1
ze8cfc2fdf841b250552c97911f421376ca7840f197bb0dadbc08aea6dac1834d054bcfb2842c1f
zcbe51ef749162938f313f5de1042c14be9f78eb84bc35f3ed2e9e579b226214243993de8038069
zb0f44b430b9eaa589ae0e3f98dc8e683dde4e99ea73cc56cb04d1b3f4eef82c37df61c8f8e2925
zf0bd17a458c946364f36bbaddedba78020dfedcd5c155a9276457b573de33207e096fd6f5d4843
z28152aab9b1ead07ce27ecdc3e7bb5dd5a9532c624246e3413d687cd57f5063894ff1a065a6a11
z4ecd42d4b6670e70801f3e1c15e6add2b8a97184d41f5a735c4d5a9dc6ab3a6069ee94927be119
zf6bca7d081d13124c4d153fed32d5ad39c1d38602c02f842df5c9c63f84d08c44d6ee1f9793193
z2dae68a24feec13baa13c1718c2bdd24182f647212cb15bfee5afb653fa638b7878369cb30ca62
ze4d7149aae0f9ab53a083c1187d934990c1f1dcfc5529714ddd2aa4ba5b60deebd2cffb7d7162e
z0aa2a89c2ca87b731768ad2c39010f8f21046bd85b107f6fdc84964b56b2ba386ef5fb9ea07e5f
zd43e151e5115065d2cbf3860c3d7930b2d9cec33d3cba2465935dec5477ce3a419b284b116ab51
zee22f05ee4acc176e8387e6e13bb59d57047d06df9b76947ebd78b0be5bd09996021f03c3c128b
zc9205196a431c15ce85f21d526f0609e46b1ea1c2a994111f48537a0c362a9298d450003a788de
z32c2fac8087004a05b765791b77501e46aded8a3231a7e5a70f7059598222d2534cbfff72881a2
z40e84ba2207fc5a025fceac0289ad5e47cfaf61e2c8952f67eb128bfb73ccf11815d9b838f025c
zd84f464837334065290a720623af2578e6e3cecebe1ddafd88bb1837020f66c1a709c6d9608d70
z0af569286ab73c9485271d80082ff1dbca309e13e93ffa110cce32d3d6ba0f2c5bdf948a588895
z40f70db0fabc7d9b454d0fd053f77017467ccf034003ee601f32e321f0f69a03517ac6f05951f0
z57d4360be1a7656dfdc88a7e41a1429c84b575ca8ce3f056c42d8c2ec76007b3edb62ff2710e30
z64288dc377aae6a6506ab62cd68576a39f5adaddc1c79fb55e99b1e7f122b8b670757301a835db
z388ddabd7ca7e384137f5622e24fddfb44a18e5ccc8a5a04b7b9e6959c96257301cad78ae66017
zf62c052b7f2b192cd802ea13f38a2c0864df3bf5aefd3cc0939a98e2f13b0735b83b923428d103
z7a28d9750d523c34b576c7275dac2d10f28b3e3168f51e173864fcc12279c6fd2ae5b112872499
z2c8df0cbff77434535eb65cab6b00f186b6896ec9a6c3ec11dd963df8de7b953e67f4061fe9824
ze034106baec6d828fc130d7d141792658c2028d20f59b098e3439e5be451c1e981e4d22d2d33f7
zc9c959b5893c56d005ae3ac24cca9975a210da8d6399bfcaaa903f6e7793f1f57b748f4ace9626
z87c4dac3a37a5b366220d4912829f2b295e2fff484cec33876889f2022a29eb1a71f5a267910e4
z0cc667545232c6650462dc8458e5ea167d21801b3af8082cf68414ab078757cb84634c1a1be9b9
z04bd2670c21f5cfb3f82464f42868ffe9255e8b563e620ab23e26094d0fc2461ee813f79f3019e
z33b92174d1e2e0cf97de6c02e316fdc8a7f2a11c4c00e6f00036a167ea8960ba570df4b7d0bce9
zf5b739016eb7d556406ff5ae482aa0f907d24b42799f582c2fca162f47dc8fef8b0e6ea3d7f27e
z82507cc1fb93098b5ca372fe4c714c43c79751f21e7e4c00c4f91d451bf3701fe7af7971b62ede
z09ff943e8eabc81d837e94f25f15f2d124ab6eb7dc097619293e1f4442b8eb9f6e511e181df0cd
z914dd60fcd2725837e2f8766327edbf486dc6b893fbeb20fb46e26a3c8c6cd07c4433ae3a290fd
z96dfe980ca3f0f5c5c8321757319949a57ae9a967837087459607ad43b2b431a22083d7fc49c45
zed6b8ce923103ea2c8cb34d2294cf0554907aef5e579a50d278a890ae0bc65cd52466bcc669357
zb6b38d1044494de80c448f0afe3272a7b4470935dfb0ef59311021eafdb9a335a3ad39a5fbc3e4
zc37061da342cc3a85227d6d1fba9ec6fdb0414badff2a4c589143435d59a7ed6796b7140409ad6
zf996fc0d5a897c1137104b26b9823fee09f50c92abe5b2801cd592bd88c736cb806673f2f54875
zf3fb83fe962eaa432e3e2fab91e57e3e5d493ec6249123c8e5fe68f3f7e3dfc68cbad101564a89
zaf4561095b20ac30cbd58a9e28f22dd72a617f228b30f047f010e8f42f307ffd39ef6f6f6a3738
z55c9a2e53cc5ff9cc5f953660ea98c872b8b3bc41180a2351a556d166acdb67d55b2c6f35d10bf
z22f6bbfc5d26d426954ff949d55c9475a38f780e1bf2458b8f953876f1ebcae284c94d3c9ba587
zaf22da2a59b8ebd017784fbbc5ef6caa7ce1737695523b187a69292052e7362253ca89d1e0217f
ze3788649eb8645929e3353eb156e6f3b68907b3284657d414fc3582def428f70e67e2d7199ddb5
zb3cb029830dcdeff85818d9bb61f6f5b0cd76dd907352d7481bc4fba35e6bf7dc9a0ddc8315f54
z86117cf1da3286e728a2876313e5fc2270548d8e6604ac33c204d34b152c3e02f1361ade567478
ze73f4c45b97996542551fbb34c02ce8c2713b27d6f00d17842110148596a035ee984b455fdcb32
z07941623fd0c6ec9bb5eed50b128ae13230b095c91f74807419d66617019a292fb10d483f6bc1a
z9a3f46bf0d5ba9f64cc228a16ea6c99feffcc9a2be4362ed73b78d45a366b4aabf3a2e555e2d12
z7a1b9ccaa94f814a85439bcdba7b5d31dd7650e62e1cdc33f6c5af39d00d59ed80e02b07e7edc0
z97cb66fac0cc31db7f83773fb6916d3b8bbf6c92fe7e29f89da8e43b74ba2205a2b233186b87e3
z1b1453f94d9c7aeb5f73e04f652af4617581a4b83a28d24df54d6b8b2d459d1657ff33f83cff61
z7d6ccb50d004d0ee3d741b6221f11698fea3e3dd04b3fadc7a7af058448e825fba3cd91705a2d2
ze9ee14cdeaddc4adf908a3366e9ab9a8d83d55c3f1c52b5eb9a49787264790dd7682bead8b37c6
z5345a61b936149e346ff0dc9d0565168fae3ffae944a155a54837724abfa2b364df8148b1eac8d
z5bd9e0bee34edb30d1be8ee96e41bfaf4a53b5731357f427923fff8977ea9c2ad0b2de4e0003b5
zbb4125a69aa4bc7d3063d8f1771ca4c2d801ae064365ea0ae00fceda4cba6e15f671b2e165bc9a
zcb0fa683ca963e64ca315788fd6d19ac47fbd4e566b3dbf5c1c0e295dff6eb20bc32e8b688fdd4
z70c54abad9d74199e03bd62075b2fb44f22c301718aaba9b0f0141d8c0a939913113e18a620818
zdc8a999951f192ac1db6f241fc633c57c20cbcd223c54fc1612e475da2d81e94c5f8786212bc5a
zf1912b727327bdc104e24af5681d0e8aaecdb2845d9f655f3da0313fc65ec79ad15754d80dbe9f
zdd2dfd125602e848e67b60cf1652746e9978636ac364f2a55c2fb40ef5a3179e323aa7c2ea6acf
z2561cc844626e8f08c7caee2ce7da63be6b596ede13c6f1b0c096e903c19525f5a536c4e6db3fd
zaffad5bd6c2625bc7cf41e4476127b29ed3f45dc9d52e5347fa711cf943bee13acc3a200c89a30
z649412f1c73846ae4d854706d249a622d070f95f6715971d544cdd89414b791c65f32decd9f4c0
z1b9e561a5cc42f9fbd4142e9b3429d051c36ffc0897652df835a79c1385fa6fd7cfd334b11fb7c
z3d3367f5d4d42e8cc71faf4138cb0dbffb4882ac4865f1f3822a585c3436611e89374a1f279477
z4c569ddce8d0f96521394b00b7d072c8ebc63af61888bf18c57cb9ab1211f1a659d47c6075624d
z09ccc5ed9723d1fb23320fe338995a75562f3a48e3adb71f44d45c2f37c277f94827d746436295
z83021e8462a50bb97099c524b9b91bf1188c598ece1f03f6cf762c811067cf8c74156958ce9059
zaf4e85c175aa13d6309f161be6ffc439c2e1615b030413852e2c662fe2166d39d9098c29c70ccd
zce21d17277a5c9bfdcd00a34f76599c4fc94112715af19f94707a3a7c2bdb42b38777fc994707b
zfa6c03b29f1f67047bab393f2521fe84bdfe63df521b103be61ede289727a1c6c3b9cf60c80efb
z6e4db498ee9c5ccde6a76c733743e96b244fcb22f841e1786905c806d36370c24f384d251b25bf
z3bd3d5e7dd195edf91c125bbb989424023e6e1738ec47f70363dbbb45401deeda98fa4698e79a7
zeb6fb93e9170e511d924f3a35d7813c8a5a5463687ef9a6fca41d09df9d2588e8c544bf6a8732a
z6b33a2d56d4f9dad503421206a484b6131cab6f03b1c5b8abf3fa09dc2409670efc74cf2f49db2
z929656ca790e1ac0840251bf7809ab7443fecd21fdbacaae69e4a76426abd11c6b1e7695b2b56f
z977c0b8f707056f39ba1e8056927b33a7779205ce6e0da4df84385aebd0917830149a3cbad9f21
z95f3e9c5b4c6e8720aea02354c68151120dbe292b37c66a824d2a8596d0d3d483bde12f7be0438
z02139f7c2496ab9ad8b95ae82b51fd7e28962d8d0d9fece945915cab3f2662bb0c5e97cafa67b9
zc958f5bb8bc421e6b9a692d86046ce202ca590919fd3e8b860afa16673fd5d2af59ba322b661da
z931f08cec9f360ec729646cc81d3f4a6baf172ad71efdff8546d09595f2cfbed8ff28e30f1ea11
z249ebf57b1910382d6802537420cda6e16b5a955413d76645dfbfdf98265d9d70bf9432284a6b9
z7fa08072cf7014b7173e758fa12f3dbf0d1e3084ad4182e7de373d46d5cbddac9ebbf98f15d2f9
zc09706dd254d7b451c9882dab0ef64080aafea3101387a08c5cfd1b670c2097dfbdc824bee16de
z1baf2124afa1d98f88c6640f0af6e821bd0b419dfab139ba2592c0b0ab0074b0419f2fbac95a01
zb42484113a27145f52935dcee29af186e2435c4598fc569d68f760c857923d704f7a6dc54896a5
z8fc2e492ab31206211ccb0ca59afcdcddd9b21d4e210f1832db8a5501ac01f02e93354c87c4378
zd905b4ca68aaf0afeebb970920c5644b3aa5017c8b9d6bcdf61866bfeb88888437e74dbb08fcdc
zb2bc10e024bb7abff6f56d5b3da2e3abefb1253cfb94b4ba7984da4978022d6f1a5065bebefcb6
zf5cfd462493c6e00c8adcb62707b6a3f509247fb012b4ade48f108a8f3e174fde2d85de3c6fe30
z529a0863e1e2ccf2dfe436b0704e53c39476d0e513bee9da2ef8ba3ed171c05f335b2b1062fd38
z753e18f1c040f373a4a31d661166b74d72b06a9fe46cf7ed8bc8de7823dae136b29658f50bf483
zd3c751b89f5c4ba15a2ff801de05519a8862a068e11cce6cdf37d9774e4d933b5cfcb31492a240
z14a620243c698018833007a19bfe3d861ebab2b6290660771f6345bb58936bb671051ed0d2521d
za8b5195a28be115023c48e2e44b2399cf2578d6d1d04049c25ee2c0d8b28747895a938f732b62e
z2e5423e0e36e4888763027276c413cc020fe4f7c4f60c3900a2c01d68ae43d73ec74fc3b3ec210
zca4790e28a3ebdf5c78225e2e5afd69b695d161f99a033dc2a9f9bdb9cbe070a6f7150f8407ddd
z81681ca42044e20f98c1db8282e287a60f448e53380623b52b0c7d3870bcaf1759c4f7d5186e43
z99e3a75f70f28256c81e878dd13b0aa5c2ab1097c2216c1dc3bbcdcc6dc2afc2d6fda9acc67777
z0d777ffcc2bf69acee9f5007e3b357857d3cd5096285b8a92d1c4fb68f3b0de08a290fc5f80c8e
z77ccc14790257b1de797174a7946c4b3b03f496f0c9a043a4a27d040236eb23eb5743cb575df52
z00658d527ee3ef3fcab6e0b97e8da59292ea9862c0aa7b1fdb657042f2b3fc8d606a82c5e6b66c
zad8536547a8f7d876540fbef42c67792b17fe2267b7062525af3be49028b84ed309cb014a7945f
zbd58edaaf3ae7f342dec1e425596bc83d900c0d45db9e6f82d107bfe0ffdbe3beed14a067bc0f9
z6462911c570e33c8654cbab0640fcaf599b69494cc9198474835d9d2e9d80c35847caac92a381e
zecda4970c0772b01b2913b0a1c330931d25e5ac0e33f138447c51bcf91732feda054a99a6cf4fe
zb18e726db8459eeb79cea537280a730127cd8f51430b72b9a24c95d1bbd8c13722795f61b3c96b
z99e85d471568c4aec16495aa0a48ca19fc4b8416929936e296ea85e70e8e58a8661ffd38d45eb0
ze8933cd20ffd561c642946bf5d72dc521c5f9cdfa3c30f89d55de07a47be1847c9096e306b8905
z0af5977a01a1ce3bc52d997438cc926293f090b302f0ad54924dc1741ff265dc3c76fa56749647
z9edb32e9b71bba48e736400906415c30af68642300fc6683837c99ca4af7644264002fd6099e47
zb35e2dbc55b7dc774086a9032f5a2c75d119a897c31ca90d3612b9d4f126aa90a2ca59c76bcd69
z243bcf580a6106b61111242369f70b349424a58ab25ae1a3a73b2da43486088cd753e80b3e24d6
z2f06e81c93f0fa878db55cc3e2309a9eff09090680c4dd2405aa65b84f228fea06ae277929dba0
zc8f656755a4bec337bae7012a0686d6ba7e6ba8624afbea00c5e4c440914055113098f5b395399
zad1ab336496540d6b0897fc9678510dc07f5b0a2c55d5935935da548f01b7552d2fd783e8d17d5
z06495f2c7c9441e48cbd43ef6a6ef3d30469bf7b77392c7dd452401932a15f33a1f94e42c2f3c4
z02fbb09b064389d1a9964dddb78b88a2c324ed5e03093c0afc796c792ea9f33752b2a4cdd5f083
z76196a4753ed35ca00481b85f83dca7f721b5c8baec6c5bb08edaf4b2ab2ff602b1149d3b0c6b1
zf26fea15ce71335bf273d19e0a34bb85a56ffbd4316367a3c20021de8109d335e6a6daef7a89e2
zf4638edc071d66a66316805d4a0d2e9bde548d265045f5008d661ed544524954ba30380fdbdfd6
z882443b7a43165e09d9800f2ebe49e68630652eb7123df653900734f1c9bb28ee7674e8c5c51f4
za743f00e1596cba14917be73cb1aae479a7224c18a9e170a303b1bdbb4332b5ecad466603d8742
z1b5c1bce979cc3fc4d3c6205534b2e4db2765cab077d981e88b84bed81f0179c3d2f14a10bdba8
zb6a21c35f5839715cd4d1109264f794240d391f5eab140d0ee1998da34123afaf263948c8be48f
z36ed668b568c1ef305568421ab341ce9c2f30219470343259ab8ae0a040a7b3859b36822f1815b
zb6779bcee343098598ad81f92072c9f5444e19f5240c8a01543a2203ae890dd8ca0d0702f35f6f
zcc756406e0fded1a539a688ccb27d771987aba5d8391bd64e6c8a2723a957d29fcfe5841482541
ze6342d90e3bc026baf158a2d17a86c13a9c7dbf6d5c9f7e4bf078276a1dd8b6bd9e703ea18eec7
z8dd1fbc2ef5d78476d56b3115dc9af04ba9aaa72a93b262765751f910b178d84515b50a6298fab
z78fba6f184fc4687adebbd591bed0b3d3364d9bed1c44fd5ed72efb59374c5a3c8c6e3102942ce
zf062c3d8c41c80b0a77c98ce6295720b280722d2e26a6fbb427a075abda04c0c0abc49ae1a1de6
zc4142bff82328bb8bc789069ec8ac7ac248d70e4ec664f36acabc06cc2bed680d9e61624355faa
z17e5b5695b0e5eb647c6afce586346ad8bc806cfe505f27d22b82fe9c2cd34f5af73ae4dec34b8
zf8104eef92dfe98aed3a1d8719881457b849b8e7fa744a91035e9db3d38e1fb6cc914cbccd3ecc
z16922e638e67ffe77e696c8fbd85b4d354d1d2da28818ec79f1a3393af53aa6f845f2b538149a0
za4374ae33df4dd294166f3744209946c56b90a54e2c2b35237e16a4566c115aad396c630709cf4
zd8c51c22653ff4d907b8455a292198f837271f5075983d4775ae089687d828ee267eb90f065acc
z628d68f34458fd51839b78827a588d97263b3374bc0447b9a703d372f1d4382c2f7a8c60d97278
z4056fe30faab4202336df5f6f23b3465da4b10ee11dd1ba285b9e9515d1cac13493a36640eee09
ze88f2d83d39b7d06a9872975ba54fdea9a9f75b1abcb722c268c95342e6840e44328f6aee503e5
z3954f744546c575ade0a9f35c034c558e23450928b33c306c30761a685379509433dcd93e9e2de
z817c26ad2a6877feeb9940fc112bf4b7c7697d00558112314df253d2af1c267d2266960f29591a
zcfb20ddfb286938f50027b1bf3ab40c53c015b33424c3aa05e9cae29effafc12de6905a9c653ae
z1f04b11dc690c2c7339970a41522270fd48b5229350df21f6c89d8d4ed59115f0272db9cee1e85
z5cd6605556b529cbc8204b56439eb5095b4db99fa871daf697171ebecc01979ec46603c586e035
za663b64ab9dc69d37179672315b999e9a1577cc558e4231e499a5a53abc929baac95aeababe928
z19076e66d6a08f905fdb1e1cc6ed78d95659e235a9da3522504f12c298cabf9040f6bd258db507
z864f84f67e3606e3b28f1cdfda8ffccff396569055dedf4bcd15a19865f951d237ccf90f16cf38
zd0df8393ec62b6725936c409f86618550ec92812874b3a31aae873cfe712555aa894
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gigabit_ethernet_rmii_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
