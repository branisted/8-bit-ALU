`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc3904db24
zc5b0040322f5de9957e599cc94de9db74bd4c19709cb5f8f887bf3183c78c7b1fecb712ae25fe9
zbf36c1aec3f46a9970eeb408b685c353aebd3a89407438d6b759bfe8b464c36335c2c76627192c
z7e21a060402679c6ff07b0b7a557799de6d1284daf4449467462ecccb08901828ecb0d1bd81b99
z36f041416d5a1e41723bf473bffef4db8a80676fff2c16a0e9f4e6850ea24a4148e9706e1f443f
z0afdf7f0b1786d24e5d05a79d9b90256093d957266c7ae3af652b7a2930e103e50024052d9ef7b
zd3993af204a54fa525702fa2059a599e41f91acc7cb1221b69e2ccf23335962914195b9d362b05
z4d8b8449ef941dee2e243da961305ecbf4340ebfb053a385c3e3d148439c7c05e2a82dbca0d337
z4fbcb69f16c2bb83f3f8c907f96d48bb03e55ee3673f94c569a3170f68dbd223b63a5e1bdf4549
z959236d4cc9fb76ebdc0410f3b22054ba0ee19b0ca9ce164b25f37c1b3f85208f5749301e3ed50
z6c64058044c78d7bbfd4288a35b8de9b97aba018ab1bc54567bc147697142a3f93d667e2f6653b
zb56cbdee022660987d8c2312d1ecdb486f2ee3acb5774f48f73124725c92ecde6f013b62a3322d
z1048db368c70613dc223b732745ddf28ace42d8508d473d05379a4997b08ef0350bac9aa9a9af1
z69218c14fcf702730e041a67f466ed89876e4fe96aaccd8d3b88c3f41395ddda611886e83baaba
z88810dfd5d25fd15b204b1f29960e07be7cdee32e5500ed6398d2e7bfedf799faa2b60dcde5095
z2f7063adc0295871b598536cbd418b62c89bc45f2d63444e8a41808a91299e0f405681bfed6a62
z2738a485e607030157660936170511ab25dfa6adab73837d554fd3d7a013b5fbbffc31bab5d791
z203cbec8e5b618887f964ba56fd19b549d255dc0917257fd3cb8be05cda66bcc4f65aeedf4f574
zf4904bf360ee0c3550917668755d8023a9a6fe094a6c574d3001549ec817b00edc4b648fe052ab
zfb7cf0fcc78861a8edfbe78cc4e19afe800c203f595cfa6e3418868971366842deb3872b072e32
z26688c0b574bd7591d73d059e34a2dafb97fb24ac0ca999c11571a0e736df2af5a2440fc390a61
z10f393619cbbcba35b4646664f1ce5d0c6c24a8eb45c3b85b79aaf3443eef2e3f4bcf39116d406
z2fbcdd527db05ad1ac5d2f76aa375a2b76f493bf19cc44890a668b34e9618606dcfd04b6b8410f
z0d4cbd62562436626d77a3cb0b2e549e08d391ac702486a0f3fa2591b6b40d9553ed3fbfc2fa7e
z5617e29cd6a75973d52f74b339cedbb3f49018aea03efed5830b498e8081072738b5e2adfbb33b
z12612b025931f2ac17f17333d3f2db90b7de7e4c048c3aee8476407c48c40d7aceb8324939ddb8
z460860a53a2e316a28362f358e91e13bbccb116a9859aa086d082cd6e1644e6e4cebd0ac454c0d
zb68b512450db528180d2dc60b7675a09e7675bf245a8fd07ee8d74c568bd7f2bce4313e12e2881
zfe7a07649564bb0a9e92fb03ddeae123171e7e2e81be0215e77a0387ec62e4cfb83e43bd91ea1c
z4204c0990323c79bc1fdde170874c93da1284b3786b08ebec86abf3b0176e7956f9c1145fac1a1
z353f8c879b7a02abe89eb236b61386830319fb6344a4c1794ec61414ffc1cc7f88bb1a3972a229
zdd67732ab3eb4793bbf97084bebaf2622d3f13ca38c706ae5c552defd1eb9a2ad2aef27766e639
ze4166f3929f99a9dac03029a2181718bf975521a4198ef9774f978823e0f328d608f8e01407f71
z4a6725cd97d2f1b9cfb09be9b8acc574083b1c0b80cbff298ba5c4e71be400a098579d54eec463
z17c6f296ad96003d1efdf02993bc7fae5f21f4aa25b73f3df7bac2ff5013f669c049032974a5e4
z21ded60dc8b2e4320580c82197ea6564e8a6ebc65d44fdc7fd91de7f14596bb6ed2705879fa8ec
zc8983005ea3cc6d00d8beab4516ac1884034c476fd16209bb2e15d171711fe6bce74b7aaa9683c
zea75848c84ec9974c37fe600fba6ea574d9883e4ef871cb3b6687468e94b33a5203fcfc9ead779
z7df29830b0ca199c77569bf6150b0983c8408621457e147de84c3d3fe8310672e1795ab610106d
z057a1c4cebbf8dba02f5f039bc021a6ca9a852346034c690047a70b69013f3aeb02777d3186756
z9a69945f641a589d3241117ed23fe4d7daebf98c4b0c472b894d72d52719f0f5fb031a7cbd0611
z01e7877b7916d772bae41d4189d4ea5cfc60ef6052d401586269dd8fd6e1ae46ca679a994e1e5f
zf00323a9a3eb6d7c0699387383c227d38b97f3664257bb37a0a13b7280d066b9a304c31cf5370a
z72c2c3c62bf119dc1098693382bbd1e0e2131dc11b7931317af0f0fb26e809b0062e327b515c33
zbb28a4f160ebde3699929c12eccf2d1210397862db7f679a4a18f508f5befa5c14e5bffe0f0aa3
z6655bd43e28914fea8ac70fe17aa0d0203ae8bd9b08e15a3b6f31c2c3923987871033980bc0155
z906f8ca669e08c546abcf1ad8e1078bd5e014648425c22feb5a48aca5763b5088dc8ad1917f55c
ze2abb801b759292a4cad7bb4e04e8c0b694f4d6a603f7a03df347252878c76ef42d3f957e0e5b5
za621d894fbc8c8b613d993e341458c010b79e9955cd475b945bf025cc714c42e014d091d2ec703
zd47188a3946d5c87a964ccd60fe1f6e4f08f2d64c04c0fc1a439b9a15523b084b0a1e1dcb0c547
zd9947520b4a24e49c3a09aa38395e17209e92ee0f63e483dffbb7c56f757c2845777203e2e37ae
z69c2225ee2ff6b9089e576bc4e9590ba8980f0c53fb6142523802b8dc3572d4f29346f9348db8c
z28ba25d4b98cbac8366ea5bb81cff70a1f9a16adaf84983db9020775f071b711c38f7cd1123a5b
zd48fae656bc534db0986be2a0a09fc1cbb7b087d89b843894ea905aad2cdb458a54fa802e43539
z52e8f097b6782329e2ad59cf8543a1bccda8f9c725ee1f1b71ce2c9063388fe3450ce905cd24c2
z6a3a00aa02ad693e2f23e49298cf4bbf9537f43de793de0007f487042383cdaa3e6be740fbe5d8
z8d740345e6f0a72a07d8e3c36ba1460d1be09ec0575497490d9915a2f5bcd2de5891caf7d41cc8
zfa0fa252657f8a88ce9ae6e482caab2f984dc792a02a505e11328b57bd8ab70d16d906a38b4022
z1bba8a83f1b9a3151238899c0981f488e680a4582309ed32f996c1581e9a3f8d7a1a5f8cffd1f8
za6225f86a530e496473b6399928a61409c851827719c11eff5432634c2a06c8e5259832eeb8b04
zdbcfd4a3719cb2d7ef92e8d167d7fbdd8eee9d5c21f7bdfbbc55477528c8c7ba437e8aa637e7b7
zd7c67c2f6797bff43a35fe76ccfa292ffe41ce5f109cf42f7827fc8ca2d4f46e3e4c69477a39fa
z9d5051cd7579377681cfa50bc8cb310e7ef838f34da272e12654365c57f949c1426d379263cd1f
z9c353d4167b280f5d8251ef7cac8f472d2e3add15b1dc2db94a9d127e686e73ee02d74b0b79864
z5248869bf16f473985765f25eec50f2faee7eb3f27e0df0048df040a557d2adcb598e6507d5c74
z2db4fd802fbe63b63eac831f0952755f729fa75e0389849b15fde8abe529889f78fca2dbb47e98
zb4718669925eacb7d8a8437fb2b94718c99c0bddac01795acc9ee3e4f2a4ec1071d643b419133b
z5411134624dda1fcb5219a9d61001c47e90e87ff57df5dfeb6afbecfe9be91369b01bcbd445e5c
ze3c66b6dd6d10de4655274712e0af88f5722d299fe390b79571e760bd07e5b1b860fe9b82e9179
z13b85b302cee140505aa32fa831cb14674dff056d9cae372ff829d33caa1a73240e808d2c8d27a
zd5a48010fb802ab27bc336bf0269219d3ba71fc23e1c2d204f12cfc7a3c2f58594260649a5329d
za2a028098c8cb07ac38e8b4fd98d2af43099b2fa84116116fe7df6ff0ac7229eecd8fc77389644
z86fed630e0b4dd6741a861b2627d77d5a9655d50117ef39a734b637974bf19067d877f9befabbf
z1bdb5db35d5b0297b1dea5213b840f30758400ed8ec3c7cd9955a1a1c8b55dc4af1ffc538bf843
zfd2fe1f37172eff1bc6ad0aae1a9cc55ea9a76b659bd0bcc72d90ebe9ffa10798b1fdce6c3c445
zb5e47f18f0975f8b2744bb53def33778a414b9d8b30de07eab4f014ebe48d7f6980b1cce3fd26a
z79160846cad8781b0914c6857a9ea863df90c7595aa1eb97022a526812b682b2cf4b40d45ff830
zdbf2960dc4819190164bf081253facf7ac5d6a5bbd9fcce326681741a3e64cc72c8ff33f9aafc4
z6c37b572637f8697eab9d6c7f009dd7eadc327615079b0275243eb4e19336ca155c15845e25d0c
z1c504fa5034629c3ca3b3e043dc048d32a1b9d5e41f52481ed8920b2f850af3b5b32bd11216d7d
z86e52a5c28e82c22d8aab5d159e7d18c0baca389bd6fe6b521f316d0db6c28473cf028f7f67ff9
zadce61b5b5ab30b28fced6e73365d9dfeb02ba91970941970b2b70b3c59ecb012aad1a5ce2fa88
zda81dca4d10ceb0555446b766357b0d854bc4d22e2496e080f4daa3d889ea82e3192635a83e89e
zca879bd902ac3435c85fa54f8b5e20e2b9d46ca5fc4b82280410f2d2a85078662501f322586354
zd7c22720543f0598bd8dd1f94ccebff1d9d97cb42325943d6493c1a7b8779fb9b0dee121377d0b
z58e2b52d9239eb498acafdf723427feebde1bdbf5c8bf51f322270f153820fee3fe3140395ae51
zcb13d4848c2d8179ff39d6a804830a65102c42c0bea16f71986b8d53fb043ada2c80d64f8d6351
z1e1ebf453f588d52c81924f460623c8b0950a2df1f6dabb6caf983b90e9bbb2db4fc8d0b5778c7
z9552e9efbc536d23ac851eaa3cb38dfd0b187b45fa5bd1841c0a7c109cf893cef241d9431cb459
zd40b4d08a2b03b844ec056da67eded8803a0352110a8a3e1d7970f143787bd0b9aa97f4c35268a
z2cbfd2ac488cae443a523747c664bc3f0bee7041891d1e9320ee07bfbe58fd04bdf07b68cb512f
z952cb559c752ac524b60d968e886cb0189136be5f79a983eaed6fc7b7e1b8cfba6c38d21710e8c
zd97b385d7332982bab580f80e21518989218f76a1a8515badce4e44c674c828de8c39b7668dd44
zd9e9cc72781d5e72e55065eb5b75e25ce7b8add1c6a80e32dbb6fa6d2ad4dc8a1922dff1ce58da
z3b78b702444bf6c828d2ad304e97fd3e432bf48b0ff9cf1ec04dc537f51c5aae1ef607b3944e82
z7f1cd9063dae5748a13619d56a6735152fd7857f6a4379fc0ec11e42af63e822e9599badd7e834
zd2a78b7f8a8b30242708f798353a100324dba5121025a7602e648069813aed20012f82b32ed30c
z54fc7b460a8a661760d3e8d755d15a2737536b6e98cd2bfaf4e52b5843ad41bc6023acc3f3151c
z6fd94c1e141699009693c23e16fad6e6a87ec83553aea5edf2add567ce71ec1ebef27781a900eb
zcd788b387a64c0da387cb91e00e55e933d01201c46dc8667eaa86fc9d342180ab4621818d00eae
z615536435b32d1c9758bed2d9018522b5e73734ace44c7b43da7dc1c4c6cabaf29975729959c07
zc4481d00183986b0ebd1814f5628043973b54707a69ebcd32b3f38bdc355ea38adab9dd74d1f2c
zf4fbea922861b68202fc9c0d836befcd4d0029f6ac7934219e74ddf81d09f20e1b86ccb5b0886b
ze3ab3676ca68ce2eb6b2285bd669b6e80e1d7a9b29b74221decf71045967810674c1415414bcb7
z00b941628b042a4e138e749676c315634fab3c74db6e336964d9fa8d6b8610064ef13cb3efc996
z373be6d2992d1b92a9baa25a47c88cbd05e248651e91682ebd141b8148540c64eb34a1c543784f
z3622916405e6f0e44d3e9e1bb952ea0276bbd894d1a999fe1398b223fc99ff5ec70e34bffa1797
z28f4d615be1d59e9850a42401ab1f652d0eb3a9307cf49116471087a1714dc64417b41b63a58b5
z7915a204d8cae06d84bc7a99166983d5e8588dfd568f2828058563a5cd1c54e3d05bcddde8c9ee
za526eb444f840f8f73189c19b651ef68710d5ad28cbd24c06e8b720e6bdbcad03f86f059229472
z254e680591abbd1a14d715419dc829876405260dbcb7fed885be0f708af80b984b4a09e6a5f0f6
zd96b9b605df11176af6c5e78417299c18d5c6140b1ee4805635ee87bea46b9fc45525789bc69fe
zb6ca5bb83d29b77fed835479d40d9570ed917b020edab256f343e337190ee49cd5d0990cf9736d
z5b293a86206124b811bfc0cc995a2845e5811d58f1a63f018df57cbe63017b7c28506355ec0921
z53ea4ba4591b0ea380b97ee2b0b47c2a871a86ec479375c28b94b02cede08025a8a3ca9101f55f
z0dbb411846548e3bb9060cbb9f03d9519a1540cbad813bb9897a372a10d73da50e60bec3c61576
zf6747a00609ec259f5eea0611b2d714739a46d77bd4df6e19db3f7a31d36b26118101c728a6363
z38dac19b28ddf76cb6c456200da51ab7461b0979876882a4821511ca671f80456c8d9be848e037
z660453b26c2e211f5a7fad44f00f1a7384fda0ebce26ee3083708c4f55ca8b44385de79f973e9a
ze69021e3a0b62b53e345fdc1f011545b1ad70d8bc8502afacaf2921e026b281c083f071996657f
z7f7c3c346bceaeff574a7ca34f32ae339d19a9fa9b42ab6ebf94341b572ef92cc3da9913531c07
z7b32351f9d9d971f0bdf993ec28ef5c7873d76df7eed3b6acae36415c7fd3c4b0e9d58016c9187
z00b08b9f125544d9c18a6dc291e9d7a43694b17abf695f88d64cfe28ea40c2149fd72d4bbef59c
z0b792c9a35f9dd3c4fafb4273502e93c338ca25659f3c0808660cd63c71665256b4e4f3011ccdf
zc74f41b75a2619785778bb0dcfddea3104d0f235978202321906b247efdde4196a9cfdd1ecc671
z9dbb026ee10649472bf7ec6255a99e533b5da80b45fcf23f1cb093338c4a4dbff2e0831516b334
ze51b3f356fd66058635b9996df9be7aa36de9368268b260f50fdf3d9d6d117a992a1a6356ed537
z62ac5d4db9dcd5e1bd6599bf82b52700b8b280fc0fba8ea8dc51b4951b0b34316d83502bacf3fc
z6a23bea3b745048875aaff8f4458a992d18fbc3f26a6e01da99ea76896c59e0eb8e7d656f386b9
z30d9cfe47e395fcbaedca170d432fc5933b95fca81c651a96cb74b56610b3f6ebddd2268b60c28
z31e396cb258bb8c6c841ccef7475b8d9e65dfa9c0445cf986c4da331f5a1168843a20ce1e8cb16
z162067c1e1a86ce623b84c664c806c6d1e84eb0d59a00c5e44387d33ade0056b81ea54b97cdaf7
zb2aed63db7031f685e1966daec81915a36fc1a9514c571d79d60e82e2889c4e2fd476744e259f8
ze596cedcf88bd45ba66dea15cb9728103a589e1a731018a6913be56f63f68dde105a411df4b9e5
z0db0a20a0632c89e2eb1253a67a1fec0ed8133f28ba96b1e4f0530d6d0beeebbffbb742480e6a8
zcc19bb3db51afe3fb7b8455b9b6e1726a56525d507ad44f28193a02f06768a40593e20fa515d5f
z709e12d833781950e60c6760dc380b286ef177268332f282c564aa7c3faf4f5919287ca301a227
z2256aac726043c2f5ee6927ec4e6cda18a45f7772d57770ed8d6f3c812aa71b0790331ce626372
zb63bed678ea58e493e30c527dfb6b23cc49a50933dbb3cd9eac009ff8386978df5c185bf711d54
z3374b006a222d7ec3911fc59dcc3941f4cf464e9613309e72aee1608386079513b3c50a6902594
z728a93df07bf73b91ed142b9614b32ddce0c0d7032984e830d18357994ce42fa34c45d6e547f5e
z2778343268d58ffee7e41659052aa0f863eae485f043fe650aad45c294a53a931d481c0a56c4e9
zb28f0b056c36bdbf89e96d57cf9257ad41b07f4e47803ef7be20e02664c29de64761a73958561b
z8752988a39a5601b7a54cf3500d81a65c188248ddfb2d6714dfcf3ed881a6dfb2ee101e555c0f0
z77c22d402000362e70144bdfc3c6ce5ad273574da64e95d041a5df0a4505f21d2d5e37e5f3bacb
z03c98dd624bf5905ffc3fee7d4c43b4a5b14c1448d85149f5f665f3622689ab50b663e6dac6d3a
z4d5faa37335957785d9e4e6e0088f70be7824406bdf50e3dc5bb1e7acdd51d6c9be38a00c9cea8
z95b4fd0b1a4c11a64a794599f16db0bd7ebc3dc7cc09557022a0a50f01cd109a59340afb1c0484
z1d9d903dd8b64fe198e90a210c65eef2f552fd4637f6255da36628edd6c20037342a0519b6f75f
z8d1de0f1d82f4f4065066fa2c899dfeecfc317f33e01e5f57007c93ba7ea7a26bc6f01bb6a5a4a
z824e3f18cfef27aa486d9d07185790608c8ec7b7eaa88be0422190fea3a6a40e2b6b171f276425
z7c1751e83862a15b0344ac277c3c6e77e45d7bad10edaa763c59fdcb114ebfe92578325f14cb58
zcdc42d0476cebda85099bd6e164aa2587521cff133f352b4d7a14c8f15e9fb26611e1a4b4249be
z3874f37971e7703b167d5ca9761b8d4a469c8de6f41af848e1087fb61769ac33bbbc626f8c8769
z18b4f5d96d453a7ac39648ede20ed42d2e95b11f45531a6b283c2c16f5d2a0ecfeeab2e05ae291
z779405090a1caeba82a8b770f920c4ad3c7a572602fea5ad3caa72258c45292b57bbb06c33e979
z6461e266b0baf8f43976f0b2859051e5c464fe46754f57e009b1df763226cd4cbc72dbed03eb03
zf484f1cac606eab0bc46ea07f55837346177974a12f57bfa17219053c0216c845111afe328642d
z1bf818552c62a0b533324e9a898a79f3507ef89199b21a825a1120665b93ad8c1a407278a9e9b4
zbb88ac0d21e511f70b5f12617c30d520cfe709d50682a69f9f2a31d6ad23782dcfa60864314c8d
zd4240cbab9d32e142aa5b6782448a301b3b3b105a990d7e2a77190076e135d737fdd38662dab3c
z87c3aeada7b2bc2511cd3c562dc37432b1957dcebc39c257c5c4ad9a10c3d8a37bc17eeba967f5
z77c58bb7de67dda0b9343d9b9548ab6c99e03abef0d0d0adc8e64d260be8a618ac291caad88c3c
z48f43472fe7f8838006e9f27381160e077458df24acecc11fb9312ef30cc37b1a044fdc2efbc0e
z9b4df02c0c54886882ba806082b5b7e67a66fd836292b1384abfe629cd1bb97c989ff56f531ebf
z161279f58d9c81901c39f061cc07338dbf10659bf66a6f90cbe28a5ca0da5c12e66b4bdbf31d28
zcbf8ca5512bc9a0585d5e59f9379e4de77a686809b8e9de0891ede72ef70f09853100579822bd4
z81754b2224470ab4216b058aa5cba5c45d9d5aaf4dca5f5e8f090e143342f311a809ac77404690
z35b1df1e1d71995b0a1dcbbbfa4a7237290304898629873f30866c564287acb48697990b63c9ac
zc4c96e8d82b5df2b8ac9d589c241a731434462c094092e19d3c1245d116ea7b9f7beba212f6612
zf9b301d8cc4916929e0728ae91e7d806685100a4f8028edb3c9d221784a59a891e969654728ba3
z50425a13cea48275dd84e8d3f1e9c165d8ca21d946651bf5aa0b780b31e225da5784bb8e0445f1
z67fc51b489d1329492e5ce4991604a9a1f09c27e290c913a8525a3d3cbcea71e0d1f3e28470067
z170181dfaf7b097b1465189679700ee150ed9273c08b5c243629bfa5317a9b06564f4e2e8d3b3b
z76f5cf8331219fd8834349713fc9f533869f821767ec7a3bf1f4985053aea6a29b269d37652294
z5cda0930f82d1201eb3de5b924a0c2dfb35cae73249e5f9162accd1db3baaf90b647198ddd60cc
za1ad75c23bee57fb713a7e7af76338d5b5ced4aa5ebb758329211dd8973855d53287219c88f1f8
z843f1b8d5368d38a659097846c6174777037cdc087e3ece8864aa844943f79fd67c78251af8e63
z5ac3aeab113d75c4d047712b666c2396335f5cfeaf1b209d8e362ffd46f0b79f6436b6beb29837
z91cb5db04389c987ec6a1423e636b90fae16a6a0385d00e5a374ef3be2efeb5d820f14627e4241
za2d0dbc61b448f993bda15734498e82b1416f1b00fd710f1c643ad2a65fda07514f32e387b0e8a
zcdb46669bfb9fa2018d00635c57ab4062b70cd918a281450bb4a6a50a5de32c77949c8aca12f3a
z95e5e35e36b07d227f8bb69c4659720e10289314c5aa6d642526f0a96f2dff32d2808dfdeed661
zaa736c24eb6bbd836b32f09816e9f164262c8e73fefc969abf5a7fbf51614c6794fc6533ed5206
zdde9fcaa4b51bc86e798b7bd8aecf9a798cf5bf143ac2dfb9477de407ab171053cf5b52805656b
ze73f9f838a4e4e671e4871eaabab3230464a31544ffc9bd97c4de50d0cc71235308ecf97f7d0e2
z8e69db607a2b2b45e7009d43424d6eae952ce10f33516959fec490ad317eec29dab7010fb1ff34
z28b081d2c5119f1fd567cc1a85aea03789517a75174e73a1481c80513be08a41600f95a7fad3fd
zd60bab03eaa7e77246da69d24d7d5a4d14837873a28a9f992433df0ab72ee43ce356b182b4f7b2
zc2cf6615b4a91ed287021fb87e74da17032231b068b28a2a6878a650a15356978686664dcdabca
z7c0728b8a8beec89812ea7401546ac0f3ed976459b676225bbc16c00391ff101ecb665d33bda51
zf1d1631b2fe0c522d86ce0078f2c6d649c1f09b1eb36e7f4622031a071efe1760f833288c915ea
z4b4bc1ad22ce4fb3851ba4d86adf672f247bf085f4a3b6b82b12ddfdb331d06f3df3420913d11a
z0a3d9e8c2deac93911c8662c63b5e90abc0d84f18c941e28780f9b29e8e45242047d3583a289eb
zce834de80af0bf9be2a8260c893dd6a4418764a31a1956dd5640facfa1d4bb6205f63767b0e260
z4c253257ed8cf4239f6031259d8505d78c4e8eadfceb486e7a57c1a42498514db68edfb8e7c3fa
zafe2784e20a730600674c322c25436d5ced86dfd938bbb88aa5dde2272c0e987a16d9b65f18c79
zccbcdae2949849384261d22b7d4a3a33f186dedfb53a148ddd16b1616d04072d8d1e911e26d568
z5b3e1cf8929aa28fc7f098f3f9a4833c729ecc76bcc9f395aec081b33c68eab098d790dcee1b88
za58416e195db7ca3d2a89a0b4186fd6479aa0b1b03af36b2951aab919d22fe62d7f6c7c5cefabf
z8aad96cd6ad87ed35cf6d01861a2254df009f266a1760a40f8f0717b16052ae5d5976310f4de75
zf7dc99a89c98a9488336a9bd2e65e1f7181c8173b23fc70cabae337ef60a34bf54df89bbfec3ed
z116b9210f6a10c4ef98adac43d166022799d8e8c89e36adbf293d361c4b67852b37d90be49e455
z3c3846c219d04701c45515f3bfabfae0649eba27f7a04f12b28cfca4d9464e9619c14faba0e747
zcadece518ea1fc329ce75940305c6f4793ae0b0066d1af10773ea4bb3333d8b892a751c53e319e
zcb8b613bdd15fe0602cd09c4804721196645bdef1ae843e991875093a0878061ab68c9a764dbbe
z130d7de60f28ea2cabaddd00361cfe487d74759426c10c69c629cc433b0777fc074cd4b5ffc383
zb23629fb7afd3d29b2afe0a9f58c91e54a12eb816014805466e5baa0f197c523e5fa500e397b53
za9b7142ea66ec489e2f563e85e3eba44162d2c2abd1956b1db7a2a0fc400baae19b4d18db7546b
zbe73d8bfe4ecb9cdfa3c9b0b5c383c56e15d2d0b126eb7bfc7f7b846bb4466239eda8a82101668
z31aa8cb747336683528436e75d2900ec8f059fe95791f389b29e25ab221dde4757a638928f73ef
z457a7c0183fc9d39438800204e1aa5816c4becceb0d10639c53b5490e445342154d732b7d9a58e
zb9a972ca24322089a5b9983dbf1df440eb599097741090294ec21b21dac096400dda5feca27a13
z75fd489b6bad5919b59b0ebb7d7b93cc877683b85fc245e348c64b9655f2b40ac7319961e52beb
zc3f490c3cab7a69e2a45a0adc8d00c917c40bf19549b299f79165b4d55c8ae2614e99affd4a0c4
zc456f5d4bb7f3482ea61486ca0c7baf76b14efffe07e4ef2cf0565fd6619b7a05d627e626f412c
zc2c925c48fbc750664181aec43becbeadb4516935cf9c17cbb55114622d28e09a89c10f1876a74
zdb7edbff8cb8c331319164dad1b5c710b9b27b6b3f9e98d2ab6e60aa4c380dd7a6e04229354438
z8db84ed56028e185d1a9932de0e7b80e22355048106a9bd7cab63bff71aae9d0e451fdc0f3e5bf
zb68150aea01d6b4373aeb87c4c95d7f693dd82b94dda4d35e1a2d7cbebb99ae65ce450c3005fef
ze55d53c712c4cab55609f6a29e47cb3cc5db0bbc1789201b3c2027c3adc02acb6f040586d23a9a
zfceb47d87e51a8c4aaf83b5db97536d78c27c51cd773b84ca66409141fa1d079fca4cea61b192d
z38e54073eb2d3a2eecb316dfcba46878362210f99163220fbca4616e5f663cfe6a77f9f95a801a
zc2f81a1484692b9760d8666555954738785a8401af4380350c96ff4720181eb5b3473e85b36051
z0050aaaa171579383054b96e14399a7f758e890159c5bc6712be95dd394d1ce2871a7c225d873a
z31261c50371fa64c0a7e0dcbeb968e9f86db819e8f11147137ae1efe6da210fe1fadfa31dc5c40
z5c1c2b165c1a6d623b5622c7e95090579a8bdffd40c303fa58471d4c099bee9797158b098b636c
zf4a197e55ffdfb9370daf05d4f342c324b81f55c43b825998aad0419335f5eda382f7fef8065d9
z8c5cc91dddcbe1bbc60cd1a5e644ceb878e8393aa4bb71c87351d7da83dd881f97dd5b9086892a
z8be0ae869e0f92c691bbf0805ba1a510e7e3b6038564e813ebe743b0e3c9917c1748d7936ba308
z05824af422800ba97c3887eaf85ee770bb70b6f466a57c9b784ec9de7037e131d734cd84f858ee
zf911c9450c4c000939f307cbcaf1cb4de264531ea7b583159f926aae3b81c43f5542964d83b32e
z4d35d0eca0265ec87b988f449b12c4bfca6141d3998b57f86ea94ee92e771842659f1bdb7be6c8
z9535be535be51a26b0cd1a01f4723b700ac2b96268a6724737e6b9988a17defd5debad501a4bb3
z12f051fe08b5d291833cbb4ab0cdf60821b15e4dcd04971e7626e722f4b935d96b5d6122804cd3
z53dca9fc2a4e1a9d46e5a8231b4abb1b3ea93a5db2613759b7b1cd73014801342a22fe4654bcf6
z1417037af2f33ce06b8ea189d5ac68b3191a47d25ebb6bed99d6bc9e4b5d75e4f8132c5757b9e2
zc05784df9cb08d4137952c9b99563276cda4e893ca5c3782d3ea39303712b8c2a77ac8e23c21d1
z94f03c9e3ea96c2b246a542fb5135fabfb5ffebc045c27586a800f60c697fd6c2e56de37974370
z72b393ef900324d33622143fa78986e03057434547e16d4ac708e2e3d26a3c7aa1f75807fc3627
z843e446c971d38c731ab929539c27d16d9913fea61046e3d905c3fdb51051d94529798279f256f
z4fc701ad8f1c8f9a29d30ff499d000a603d6f2975110bbaa32959b4bb4e57c0dbad98848660de1
zb712e54c5114f129a71c95529146f77246855f03c7d60fa93600053e274c04f59ff34e52933fd4
zd155c1a4f0043561035a5a3a3d324fc838db7b4f45216a0aa17ef7d8e9eac9e1847917b4996ca8
z348e654a2326d8770cafaa35229da575bec533b8dde650fff129c85d82aaed9a4d0b0f8cc29a4d
z61aa3693469f324799171c7eadd1a6c19e5794a534a5b3f3041f886f5094a2e4ae4bfe5e7857a2
z979400188d997196f0ff120a0a8e19a5285de46011892fd29e34ebe0489a5822a7395c578cd232
z2ae9bc74439f9cc6f50bb107316f12bc4de09cb3c0431f7cb43865cb80d5134ad877a6964e1a4f
zac4c7d489a7260984204babf7bfda4ebf86a1132731b468518374b84a153d5deaeaf88e76dffde
z6777e40857a9dda1a98856c7d39acd0066c1dab722817c6f902b8410e765db1d058f9fb08fe23a
z930eb2266cd91998a9d8a5d95ad7f69aaa904c777db921c5e7902ecb557fc4d0437f699e07121e
z9d2f721a7905d86f0da23fcb02379f9486d2ec7e069c7874b588f506d66073cf7c099cb48caea2
za88519bf256706b0c95a8b57785819ad3ef31f72ba95f479fea0090f1f1df1af08fe94139b8eae
z61c13832bc434c8c52e420d36a6b96a80ae6d30c145bfb9fa19db98099d29f45a0e137504f22c7
z09a23c776e12707dff6c4b607de4c4010ec58d40cc936f9820d3468241d2b361d81f506ea7810e
z33cbe8a4fedfc2d1a52f43a6c04265d20018325ebf19e51cc332c9b3f25a74e1a6e10add18cb35
z1154d413912d87f8e937549f1dac4c554ec20087f78f5745b814517f36ddd4c1a0f1b21e250b1a
z0acdfbfe7c20a871230d508ab8aae3a0201774f30a8fb5b4fe98376d68b0927a2d670ba715f7ec
z57d7d7b6230580c5b0b1547117925e85037be2ad8e0229b128ccd91bbedd4a183e10e809790eb7
zfe5ec1640b25500054290b76b98422552090acca56d423f06051c405bf85f1ce06a4942a7cd4d0
zf4c6cd808c509849f0fdca74753a9f0ad448fd6dcaf0be8881430ee11a28937055e0f0337bb916
ze8e71404597593b8215c5e96665c3f5f153d75564acbac4256aa2c6d24412d2773b82245837b58
z2b04857d4e4773eb16d56890d1fc089372244e869fc18ff623528bd73bb8f74e90c4f1de766d38
za44f5f5eb1099981fe4b86bc0cbb0919914f1fada1b888f0619cffb7154f433af74cb0b7aa1ec4
zbe1e996a372b7a294598fe9aea48d9544594c003a917cef5bcc918f33a19ac63414d936f56a5d4
z213862c2f58dc81d28ffb42d695edb2322eed0605de41d97b37a451fbe76cbe45b997950279944
zaed70ed167fef56b2523927824309f247fe6f98c5942c649ffe620b88b929ca227bb6a544774ea
z0f59cc2062a6ff8b081c9d2e1a9137549724e024e476507aeadaf90bc9045cae46c5c11dc414f4
za7ad0ffb56d3340ae4b8f8cbc999db780511cc5b6bcabbdfab9e51e713be2c6fffa3b39904c298
zd002a9e0fd942b0d7650f88856fa3bdc628eea62d06c54abb7ab2a085974c972b478cac7b53100
zf95f6135be87cd0328f528eadcc0cdabf198fc3cf0ea96c0f809bc18570e32ea841f3f85c49bc8
z611f1c4f512df8ba2eed129487610c252c03aec67bdce21d4a4082ce683575707a301cee342d85
zfc1dac7823c49d76c2682e61fd6f517915660fa71ab0c140ddf5b78d676a948cd15e5095094082
z32f512afb07e2fc6fac60db3a9b2973d4fea81712677d8e27cfbcedd1d5c2eb43b3fc654a34e1e
zf86c8f85f13a8606bdbde53505e760cf30215a46aab6998d75587e10732dc4aa9b24e1328c85cd
z1dc550b170fd8e68ecb1ad0c7deb43d755cb844d44dc7d68c604afbec03e7092a323a04ed297e6
z1fd8297816407187a3663d81d0e3ad658cdf6ef9d1d40be69c4af6fe1b45b6e17629599cc87c52
zcebaa7c020d1b8fc8f83a81a1c7c7f5fe2876c3223ca6ef0e05338453b8d63f111cf03ea2ad27e
z4708f533b9004eb244849004c56771cb5ec99449e5bc94a726838e798a9a47916b22976fb02909
z9af0338b194ead5773bbb22dca4afd2fbc9283fef7795be66e69d57c53592f4e5b0e9d7015f4eb
z1efab5f7057111e5f4ecf0da2e02c40c2f32b11150a863ccb74b1ed71634be45e30bc7dfa00933
zf78e1ac534cef6c8d368005aa174cfe9ca9210aab48115354f1b2be9799545ca1a8c1b3f9b889e
z3c6e44de8791e8dfc44974c14594c36be7999776f0bf457e860f04b087d13d264331b3fbb179d7
z37bddfaaac9b21748d196691f74f2a27af002e0be13e48cc2b374eabb6ea518fa8c874a4a87d06
z326b06b97db8f6f47d46fc934482e478094393b6ea353eafb8ab59db168cbd69394ccd1c2b2aee
z2810c1f15dd019f11c5ceafc0025e4817296d1795cb256426b2be10325a61266cd04d3bd024953
zc5cf147a24ad2f7414d5df077bbaed128fd599559f940b1cc886d3880600f7df350808e6527ba1
zd3355ce5180c1d602044cca0273aed37d0a55b44389a84f73d7a2512a4c2e5ff628bca50135173
zd5b696a1cae155134a9d58b9b0801bc7c154a1c5f3c3e8f4fc6eea0f6f7803a2b6d0cead059ff4
zc2432a5464e634f9af92347ebcb238dde5940c8a4611b263890a375d06438e51375e7a186f2788
zc9abc4d284077a4d597d4e4ecf6a553806d4c37591c0f3fbe0ae5bdeaee4bc4b8ef8691e4c0674
z61936ba2fb28c11c9e32005aaf1484711ddffa1acb6ca345e33d18d20d0b5c879aedf6e130814b
z9750a65f705cfbab389119c8217328bc207a9d7dc9bdcecdf073518953ed93939e453e6205043f
z165977193a20ef6143fdb17e6a2d46c7c2f3d5c884d224f584082e8d779e998064f3d5d842c930
z24607eba0ac38ac007212d837004d7776a7e742340c1465d0bc2b63cefd0c1e92aa1cf9061fc33
zab58da78dbcceae8165c0e713b184705a5ddf961014d9da9c94e4f3d602a24980661cea795db0b
z1939fa543ba235b51ffa8f39f4057853946bbf91cb833e60997af76c1ed543eb0fc79ccf3f35fe
z83e5f7fd65e559d3e65b7c69c0fe80b6d33f7389c3d3d27968c5d4594deaee8941ce5173fbcc29
zb23eb52a7ef746ac4a317a4002689fe2c43fe9dbb206164a426670c29680d0e3b7db045abf5168
z5b079a2860e0c75c04b58a4646e21eb1bedf2c1b41a28d4b9c9eba4886fce982f8ff0ed9cc0648
z943c0ac0dac5f12d5c52d7ced2ecd585a3eff3aa3e579b8fd1f14d70466ba8d6f5448db8c09d24
z3527d660e0b28ff1fc8ffababc2b33c735b7c6e0c46f2c78a2e8e96ac91e5a778d49c8cfeefc5c
zb35c604937b3a841adc37510f70ea1b0e6fb69344a454ed253c6b88cdd7f2b66fbc43f7bcb2e46
zb8cfbfc9d56d3e47915ca1496c0493d778422ca1606bf5ff2e0728b99eb0e1f5b145dae2c733ba
zf0ea4c43e67dc93c32d4a915185f1064bf73384d0a76cff674602f7d4f102f879337916d00a9a3
z0bdc622659da8253ca54d07c8844c95bd7b2828e58fa78b23a0c5d6ca86a9dc119152cd529cbfd
z8cc71959b1a0657f39b8ca516453762163a897382926c601ee215c7539cdf3a2054e84df5a5aae
z064a8c7a3da2196f0608cdc25394cbd26c74342ca70525caea181d302182e8e487b9829617efae
z99c544a07c0c3aacb9d4e7082605b745a904bc2c9486159416bcfa54e1808a03abcecc34c90d1e
za5df7687c30d3a86a64c175bf74230f5dd1491fc1a023fa65955d0af3755d5424e00f25b7585b9
zb5fb25d1af2964b4e4d85827178ed28e77ea7bac9c0bf83e7ae670fb179679f214da2d433ad465
z59b33fcad1a0545e0d206e7b16387e98246bba6dacdafc281779eaecdb09262c0630b20a139b1f
ze2484c47d4f9bfdb6c172e8bfe77ba26fd04ccee3a03dc299b8b32f4732ca861bef66da10276e8
zaaeb68dd45304519cc197c59fa1ff1aaa6a1847f23a98df33c98ad0bc45c344ed037dde96728b3
zb2e01a8921dce0e78a193e2087dffdcc4fed6938b24311f0f406cc71aa35294a5e87e16b81a854
z1e47ec429e88d0136baf99322268d52cdef1cf7ba00876d0bd48c4808591bfe98f70cb0aa39c6f
z5fd1a8a6bf729a0a691dd2200e22b662203e0a839ad98d86598d85c688a063e0937733a36cbb31
z4b7cf3afd728174e8b423845778be53be5caf7e8559d4e4949a81da48c5c732c59f53bde4fe9fd
z7e70fdfc675b0172b3bd059ee175b9190d65411f22f75818b84fdc612ef9ae2a56e2551d688837
z3db94296bd8bb35c4455aeb6e18fe0e8fd6516f2c76e9a935efaf6cd7566ac7225c0a0f6a5c183
z9081339cae15609727b09574873863fd475ceb5fa463aed67c6031897db01cc9b5429da8dabe70
zd30161dfbd6bd7d909c0280081175a5e6ad3bba6dfa32c74ce24d3a188b496a879fb340649e7e8
zf48b39d433b8e382da55cc1ff4243ca00ee2b1c50b2d540858668e8820b2018f08f54fd17c1721
z5acaa6a263c066ca560e0fdcff831591841e8cc883743927cf17b39ee2f5254446e254a63d7a36
z73600d19b22362d1004fb7e9f5742dc0139714b1187895adea972f15aeb9bffcaa7eb38be6f48a
z16b9625558fd3a49cdc1dc7b81f88fcb00106b5cf09e280b967f73b141949cc6e7064a76c1d948
z41b4cd35cf9b5e754e6efa9f8adc48afc4a6405cf071442d349930f2147382d2f4ec2671dcf701
zfa659d9d228a9cb68cd2cff8630933b1d314e15f428539f9e914e15ca63b6fae8f287d8f49cfe2
z49d8ada870f03fb7d23f01470efcf983a23713a416402d664b745b4d362ca540f8228009a280ba
z0b8c5c8c0cfd2d1d7067bf0aa0bf63e2b5c59869a9bfdaf329a92b29d37930ab23f6bc375d95ea
zc6997f26eca9a56caf2a5edba445d4733417dd8510aa126fde73525704ca681efd052064902fe1
z8680f521f87f2cf7a1f6651845516f4da1c233ce39b225da8943f0b65fc2373dae53ae5c715bf1
z6a7afca4c28b377f4270886d2f14788fea60c3d4bad860e10b66ede6459e2c06ec1cf1573c8607
zaf68c1607a8a9ce48bd73fa746a1634001c2130d61e01558658483159fc28ed198fe504e088549
zff7151666be1428e78205438d61bf59455303aa47a82eae43be379c7fe22280caf8305f4dcdfa0
zae3207723d4bc4fb6062af44877ce00a7232b166bde5f50769f0e21a4733ebdbb7b897a825273d
z156e27f9fe2ebce4dbdfd622aae4996f4e5211614bd948b639f7008f7a9d5523556e43231f3f33
z915695a5e6857e554aff42bf62c59762612cbd525e4df1610efe79927881117e7e990214433d22
zcb225096b5391bd701681c75bd247b317531e81e863bed2dffa69d66a948430f527d0686c68167
z49ab89a5f1ab6d5517063bca97031701d0b9587b3ee50f43f58133f00a238a531867eef1486234
z13d90d59debc179563fe82d5b0ab16a75c4bd6d925cd92a6b3592b19a1574d0c51e2f71589af08
z663f2e2137672bdd2a4a8deedfcb5581dd6ada4d9a2c7ab3e4ff64b04de335575fbea9821d0c31
ze4ce48a9de4fa94be7d50c7646d29f784c3e4f1781c3fbebd4444814ba37fd0d6fcc4e3357a102
za667c3542f1cf31b2990656510c5fa9fdee921daa0c65ce695fe6972d98ea3f9414e1e7125a49c
z9596ec7640cf20a0518ebba62d5ac92e4a1e3556410b1442950e946879a27ee04632180cc33917
z7fa19d0b0b10cac688bb257d0006c25b83bb82a2cbcd66ed64658cd0a1235d31f7be66f7f31fda
z56b6ebc66a00360f09f9dd0174953854acac9b1f302260e84d3dd089c347242f186db838a882f8
z1e684249178eaa9b52ced45099bd89d44637c394411582f26d76c63a5d90de8e6f6eb1356fc3e3
z3c3d03e08b6a416e9d286414983a7ffceae058682af5b98fcc1b1f738ac6bb4e49a58174f50000
ze63aee467768f4cbc441f1e9b373be2f92e4a6146234424b8c72434f3c9c7786016bd4937389bd
z26f285c344f851a1867e3be65677ebb28839cd9299ff172a6b8fad4082da67b951af3d2afacc28
z60ad80417c5dddbae50d8b01182fab2d425d89e7ee7d651d06e5d67a915cd45e361a1429d3ad9b
z555755b00d308ae913f3162b0d2877f18404ddc3a6cc99f56f1db58c7696e6ee407c562efca5b3
ze1a8d911e059a97596ec6b543e243390d17a9c1540c10ae8d3c6f11009e7762f55373b72635506
z3fa83c6e7c643230dd213c9342b36ef08278919c5f288ab033bfdb735382176ef83f4d0af8cf00
z61c0c2797a4e2fa3cbe921614a83c8cf258439a7e496d9443b6272717e468c4dcdf177ebc6ca4b
zf6e60fb104a905b960381caa58b3345229c9a31a1af89497f3668b97cb9b8dbf803c0ba75f5d57
z303a2cebd47686b37691eecb08d94af6509f7db69b1c601bf7048ca007515a7bb6167c801b64f4
z935cefa15f5c1b2a392c300beb4ac8cb48024450b8cbbc47010b9bdff865405117423026697d95
zea501807f4595cea07efc36753c3097143916d8e4c6b7cc0a1b0401e49dccdd0cbdbff0f81dbd8
zd461468adf77a341ad1ac2613ad2f3a27adfdaa327bed7eb93937a813227f1d3c63a8df7ed748b
z8efc5a2aafeea7967a663a91aa1547b6c5f4b8643cdbc3fcbc2ddf8f5d28af078b54f2c91dd6ba
zb75fb71b1cf777ffcdcedc6a44b59c940999ac73a40129d2a27e87b2df1b814765b2d46d2e9423
z9031535476bd642065999c489d09f85139fee676f7fcbd46cadd7d441a4d93068b82dfa649fafe
z52cfb08446502e224f54324d37a58bdafdd698d66178e13b866b30220004f07900e777031bfa2a
zb9ce7d4d536ccf9a3a14d8462b78b1d4e37307ed92af32f4b4bc28c2b556b44e00157e25ee2909
z649c3b296e4d180b6e8107ded0faa5f5585005c319f24b4f6f5b73976fe2aba89818676c3bca84
z3ccc044979fee410ae68f1abc8b3b1e1bccca951b918317ebeb63a5e48303967b743229db1e5e2
z276eef88cd4c032cc15ac4b2363b338afe89c833b10e3207f61570c6a4f2fac89989b89eed14af
zb6ed28d3dbb5bd40e3ecae448cdda4f6ebd927c834f167cfcf3b4abc549f7f4384a4d2269a9b66
za9ac0fee2ba966e832637b97a214b6b74b6f378d75cff85d310e40cf10c94908cfb4a98bbf0ff9
z9f2e48e0ab4f4cba28696659976436cb7e790d7079c5689251ee870ca64ccb95272d95ef246879
zd9c98a7fec3dd7ea64851d5e0668d12627dca5d2b0398dfc2c172e57c84592dc644fac575b505b
zecfde1062fabfd29c6ca494945e921c57dc74dc074443bcf42ad4aef58c48f426895aee76f7fac
z176fd7e976433fd7e66db2d4bfe251c5c35741bf0da8e275f4c2d8b38a8eca8f6d907e999a4914
z835c22b761786505d71857ed7cae4bbeb4b5e4f8d875a9bf82eb7cfc8bf8fd6860c83bb3257f7e
z08dd7f3c9583a3b0c63d3fb19d4ecde73ab98d2a022c0f8848d2f8ea2b894805a6ef6913560c80
zc806450ff6204cda360543ad33635f007cc2e69ef505e72011b49e8035d34fe272a8d1efdc2697
z0793d94e19035b4bfdebc2a69d6fd27a3a6088eb0c7bb1de1ab49eedb5fc2bd3bb4100e54d2d7f
zf93410a815abf673baa5f3b1a94d29d51ff9b53edf973a1d692d54a26a1ff6ac4931b07121058c
za6b3d6b115811a35984b485d5933c593f542d9228234f988b71c90fb2e7e091f7076ece8b00e86
z794fe86123b117c784c6eba4269d7509823a14083974d71b764739c7b8f0ee2e9132607ed642e5
z56d256e19367f85f4e3fe9819b3183a75d82bddbb32313e4ac8fb3cc86660d92713309f24c8282
zca0708630e5301bd65dcc3ba1f20b9a88aa33565e483fd53391f0eb692a1f22b89fc2805a4abda
zf7e3d4df534d2674c3435885f13617262ad8ed1a7ec466ca242bc4d08c91e836d06570636048d0
z11d23a306437c75a7fc833112fc8973cba32b6dd01e8233afc504d3e6e9742564154fc5e214254
z100d1d0bf191fed2b84d1d34c35c1ea52b8a89bfc92990d074c68e40c2d3985d7288cf9af93ef5
z7d82c6d64d4793f36d86c36fb3afc97704ec10f27d385283e6beb7e0310cc2e42320b9ea259d48
z85ac3a47af65a47ca3511bae2a5124aa72bacf0b3b148639260ccd72cdb500351b883017e623d5
zc52d985310d7a146a2a07f488f29fd0e34acc808e52563bae4e40c00cfde950ad70477b9f64bb0
zbf5cf14f1c20a6069fd26f7f5b8837fcb0d77eded7148a21defd85bfe21d8632cc3cd0f95d8420
z44039541adfbb55c6da2443a1a8622f5d3f1749d66d718a0bfe1ed48f41ca46d6b61be0d28de59
zad6a42086b2743682a3eec64e58ad0b156fd401e109c7f1808d90a9ee18568cfeb5e988b6b2697
z2a1dc93040fe8b24bfc5ededb9823eac41b655deb01b53f38203e68200f6ee8d4a529f6986ae64
za427025e9d82c9d4086966755afccdde8a2f34c546c63208955b2d69fb22797daf5ff71bb31ffb
z961d768c22a5697e56350d9939d468f01408b6712dbd1e77d534a860d501080ccba564b7e5494a
z9b632d52d1bad6d69cc7f611c924fd0ba701e9e566472853e2f1ca667d943b645fcda1ee7215f5
z6e23561ce40ff8377d7ea782121f320e03e3b9e2445c3bbec63b3390f650c1b276c96cbaab0e8a
z20c30e9f1e1679907833482ca5ad094ee7f1f1e07d3ae570b49bf31cbb45b8076bacfd5ceaf93c
z36ab11608ce4e63771f9558a6501c22d75ff031149c88948a6033bce98a5dd255097b4a191b499
z8e1e540e081a058fa1f83dab0eac82522de2bcc0a70f77fe2c793b84831234b3761f699524dd3d
zb50c39203b2bf17babdf589b8d5158261f1bfec625c3469fe99100490a66d2d42da20cc8ae22fd
z8be4ffc283dcafa217c88a779d11ca8712c68da3ec5ce3945af35b2f766d43c53e1aac63f1e12b
z2381c82937b80f05c9bb8b98778d36993cd8c13abcd611d080ba83c4555a978c1cb543f3138199
z6270d3e4d5555c11405b88a494336f2f8b0e2811f37ff6c25163f90c45e87101e25cea664fa806
z05b4d5e31846e530e7576e97b4140dfe7fbe850bc2d4c5fa6a04437fb20a5e6ea540614f5800e4
z95caa640c1f4647dc413bd1b2b86857b8a1af9f19c752e76cf3d02e51c7b49c39b71dff3a207ab
z0a431662a375f0cd7f30b6154ebb1a147225d1b14afe8cb4ab98b1709da9ad37c01b9b2ad6bcc4
zd82222ebe427ed3327f37dbd100eceb379c3b798d15aa670eec8490694f193be712486aa0e5fb2
z779214d07e1f078e625755d6431320228095a5cf5c5725bca1a66711af10b5c09ed1ec3cf2f183
z573bd69f6cc4e631051b42c28bcd1da7a0d6a35b95f59aadf662249baf3c9b7c8034faef1fdbcc
zd4b29e1aaa521d8f1227c368857a39b841ac707dab8d0073429902a432a6d3dbd6b64b0811489b
zdca5d294ab59b11b8ba627769c1cab672e2114005a15cb2c73439e19fd62cd1e248f4059f1150e
zeabd5310ce0e2db2ac7bd2c3c25bcfd987747e3e558265bfeddace41fea8b5e48cbc4d9a6d1781
zf295d1843da99f36ad7f23b61bb99c3b10e89416b1cc1ec2080c568abe9e99e097558ff26c680d
z5530230b96cff3be505d621bfd588a1fc56a2347ad6d16b807719632600f9cbcb3a9f9fc07f16d
zcd56ce05ffaba8e53c7f9870d0c8dbaed89392860624b055af5e4420e747796421e82c65df7319
z4f3987a573192dae25ee1d35e1264a88003db4382133345ad35a128804143d02d50bcb5451f6bf
z5516b661287e0cd9e6cade43e875516af7d03da3c7f7c7040429c3e659bdd93684b9541c232807
z20c7be5eda8045b483f0881784e2986dc97fe393301a94940e2f5a6799f3d08a9fdd12444a78fc
z123f5af7578373a8894afe99e263d276fb0abf1cdf37a7bb5ecada8c10e056d32ad1a2149b1614
z007f152909cca54ee7a4cf4ac7d1bccc553251861db4389377e2a49dbce79e2763693ddf91a931
z189f9b5e5a4105b89ce50607d96b89b0c08d152af92f819124bdd7bab1630b8e67e33b7d724ed1
z1cabef03ad8b29208cd40837974326bddc6844fbf787f1f4b3797df8b41dce2f98d38e83626253
ze4551e0e3746a703c115097ffc930a06a8400f3ad983937e141f15b3b82129010b0bc1bc765da4
z44220089a58c92a11d918c60a097896f95fa2016559fdbd9c0787941cf97eeebcef866bb1afff7
z2255c687d5c039f0b1643777e095855fcb7ca5691cd27900bcd18173f2dc643ab060cdbd554004
zf0814e3e7af0352a418fa4637aa0b32cbafb3058a8fbf0147c23c873191ea796e994fb5ce6e6c3
z8850a56aafd877089ad4cd68091e304215ef92e98f89935ec64664183daad8eda47df395c827c8
z309d9c1de99edf9af8f5596a442f9ec7c67878468c3835427dffda01da956b54e94cb3b5489e73
z2a6b6225ec9e80ae84d7d0fef7c552b847126e99984ec2d8e444a206a29f23afc56fc11882939a
za47220d76f62de75d5c78e02a40575626e1dee07c959a24393b52dc0bbf754b714601e240ea2cc
z81f4ab26e197e8a6c2f6fe6a6e53c17f7fef72734f463941fff25b2b4c874992e31ba464ddd3b6
z66278b25c5a8808b970c352fde05de055a024619255497b105a13b93fc0a71f87e4b2ca3f7fba2
z91a5bc5079108b14bfc1a9c87b1e448beaa8a64984fd5fbdb8b2527243a635f15b8684676e68d6
z89508357432fe1adb05b0f53aee39985bdad7abb9d6c76409303bb03dd525726ae7afc664ec07f
z1be2dcfe58f87a2708ae89eb10c5a96843d60fcb82e8118c25435671d2e76e79735fb887e58195
z20168c9e7bd000d1ed404dcd8db4d80e4683efe0d4222fffadfadaac0dbf7918f58b1deba76f88
z540afcc47c9be940bdd72cb57e887d0f9763c2d6e48479803501af1b56e120f63055fcf94ee5e5
z6e9b1a1d90c81216575efda5636ec743e9a656ae7c81c7f3c81193f777d1495a4cf3f217cebf4b
z7eeafda5ef304b24b93a86da10e5b3318dd153f8f7a4ffef4527eea317c0d7f2bbd4fc227dc6fa
zb8409da20df25be26c64e76e98544c4fbc8a74e8616cd626f709dcbd7ebbd20c3fe2e17c428adb
zdd109a59a6d9649f376b024eb6fa9bb8683d65622ea83b85e121d95a2aaf901a7f21ed2d2c2e38
z3909b2703e9145798c4849b74687f5f9f2adc2d7b42f192a1eb361f92a5297cab6c043c8a30890
z0566de9de1736628b0efe7804aba8165dae23ded13b65ade1446641dfb4dfa3d2808eb39e2bc0f
z7bcd6afd8602206eae2f344bf91ce9c91a019f9ad7f0099be3d57017e9561fd2a6ad0ae517f6a8
z4ae20cb854328bdfb040e5786644ee246126f7de95da5afe3314b7fb1965a363ffc9d1b13b7c4f
z4d84ccddf9243d2386c44833f39233bb41762156330aa6a97f87430c9163902795dbb5a9cd852a
zd674595738f04e35de4ff911d76ffb59ed253026d013340f3114195eb9aa49d32e3d0a08cf0975
za1b8b1f4cbb4ca797559c74b54e57b3bc6bed19940ec3a5d873aaedbbf971382ad0639d8966279
zf3a90a3dc3dfbc4b3f4f6fcbd3f1c985aa8b16fd6d4f322a6587c672ae33999a988f77a666cc8a
z172137a7232c1f52fb58b982afeee7fa503a65e844de013b205613649ab89112b287a61b98545a
z40c0c9a09b538c6b2bc29bf67e1fbac956fc8ff2b313e74e57b77d510cfd4d6648d363ab14ff42
z0f3e9b40e8436711fa815c78af79921d96983ee42723a1a6001734f31c046d605eba4f46ff2484
z78cdca3b25a16b3b9568af2b29de331c0aaae9192742b32d38ce8cedcd7d9a2e7db49dc76cf0dd
z07213b23fa81065722db240064e276123c6db7184c47950c9da3c9a809cd98600a989718e2e763
zdbe2a4370949b1405f5bddd77fecdba1672286367fa72bbfe5786d6dcde3c28258a06192847ed8
z56b91da2fcf891d32dc47ac60576a05c83ee7028d70c46cfa5adb494c027a394d37d204760b6f5
z86ab03faf80994e23478db4ad7bfd7749517d3533cb2657b0d1489f091556ce6c9f9f541205843
z7911ae9c6ffcd2d5e484ffe14ced646af97ce35887c8a4965c80f0a83c0cb50f8436e2371c2887
za360076eb6912574be0a9f42ede8b0afd09feaf8b05e21b525282be57afc770a3d16d6295f15ae
z99b073c22d5536ba5efc6fe3c99940c5a375199cfbf702b1a916f2e15fcb5e5bd53f6f7487626b
z470a1b4a9a8143db914affc5ba77727d84b5db73d4a09b4177bbb616b9a310cb34c31abed790e7
zf35dc9b8046b337c09e108ce47f4233060168c14056358ab443f1dedb04db9831e56df543d2c84
z5d488fe35a5f3cd71989e7fbb13023bc8f9b6e8c34d6a5cd8c32e1370dd8cbc91f3ba1a6c06f0f
za0dffd15c77e70694ed748b3d408c9c4e7785cbbe63f008110924f18f51a1ef046443f1062f2ed
z3d4baefcdc0544cf9e7eed0d60dba572e455a6f0b7c1742d29ddfe5f27c185dbea1e1afd7d2327
z3d78b55cfb5b2c8b49e6956397de702569e4aa9fd4d211a6805fa08c8f93e715a3bb057274abd1
z9f33d5bae9670a18d8e2fed38edb61db2ae2dc4f24179de8d9a10aa93a3782e0bfe90253eea5fd
z7a75ceeb9dc149a12a90ca2aa4fdf1f3f895b385fd498b95bff1c96e6e346e8027b0c1d035fc90
ze6edda4ee7548f1757ee0f94d0937d5e4ea3a2f5f97438b2ef6cb51c6be848e2f6300180288344
zb9327b5a994b62d775957ba055f824f1075e3dfd4a50983c7e3fcdd0c48ebc08d202219571dc1a
z12cade7d96aa8cd34c2447225b5b75da91ae791efa65b4fd5f462884fd34b0be3609d34f72223b
z4d89d49e20bf3bb2daa70d74c8cdb81661bcf78410157ded74ac5782f6f69695107b2b69f7da05
z4906b3075026548c5456d1b29eec956ebcacc8c8bc78bdc3e79ad396ff1b3f916be6825a0ce23b
z6e58d85fa101ba12bdf33e5afb2fdd3e767438d1e0df7ec894df411ab420e905edab8a6001cc0e
z3f69aeeeac6a9ee36bdd2b299340781ecdcdfbdfe75002219a01322e8da83f199a7b618334d958
zbfa7086748aed96b46af94c8422452730fc97cf15a9f8ef12f831bbc0d30f83c16093428942408
z8f97ccf7f13d0ba47f13c197482117578afd5f07d70a6b55059a58d701d61aeedea87fe8b34a4e
z592b69d00c3f34a7379ee147adf1d367040104e9a05eadb032666da318ae9b2645ab85af1cf507
z173f4228af07c00bb1fab95dd886e6e106d9883ce117c57125cfa0137ce5e859f7b40bc1a48db8
z0411ece32208900fdf6612ba99b4a735d0a204977ca6a8b09a6b7f1886bf0b5dd35c6e52162e2c
zb4770d2ccda89894150825c8f79747fe6a694f667b80b8b0d81a333faa28b0687bff35b31851b5
zc2bf86b61e6b4e7196119b23a1f204e93cfcb3c6f0837a4270461376a04f5cbcb06dd664cd2ebd
z86e9ada8f99587c10cafeefd48538b5a99ef31d48e6d474c3060a2f0c7dad036503ccb24357950
zf0646fd975e265ea556ba0f6360006231eb9258b062201728afad79bcd2071cf1a540b428a1f8a
zc14d81f0c536bc1db49d706c798225d7504e1e06c32c63d92726ad39ed96894d13a8a58a2f443a
z94de9a6fd5fcb2f539deee5b308fa65e3684e649381d724345105763b9ab303405739509c1f83c
z515d6c9052f696cf4d224ce4ec250430786993185edaff694ba6722751ce004e246aeb7de20ee2
z825429d1d0e212622c8281119d05537763f2401590d3a29a14a4a74122a3624186abdb55c30bae
z2776204cac2e9fd3d66cddf2d422fde4607c74ab1460dedf7a56b12e07ebeb7e9c6f79cd7072ae
z17c4eb74bd098a98744d26cb78a9b3d8084056ece7f00305fcfaad1f1efa9a54c321a8cd79ff92
z044fc88e343288b0110ad2e5f8dbfbf2d52849bd981c701a171839e17fb25b77f715414cd451ce
z7ceef36a2d2cda56e8d5efb9f80d072090f9b38118686a3d98073cd8165801aa512b1a9e08cbd2
z9c66ea13824ba70020aad9d318aa12474096982f66897b3fbd5a62474abce542057f749a30ff41
zcc6223a07b67a1ca3a16f7743b38778ba5c3fa3345dd56fa263a44705368643e4be0e03eaeaa9a
zd823de048bf224e6e56d3586f7fc1b6eab0a53bc48464c459bcca908eb75cdb1db63f8e58e9cc7
z40788859d1b424b022af202efdf7a4339d224131b9287ecc014d1eca54f219c7975d36c9431ade
zd87f891c6e5e0236a16efb705b14aac1f6c6dbb7d034b1f03d7798f13f6e9ce9d83ef6880d8498
zd755448fec64dc037ab75e085fc7f61acfdcbf8fbef37e9f93551e25ecbc7d8a567577e4c0e503
z25e262b32a60befbe5561cdd45be903f6291db4e2d13da3788ad1679270d9bd699a54df0670dcc
z52c80a55da2a1ac969b02b703ed53f7709d4052b82c4c59a97d3cbd84fb328ae9e8dd700f50541
zd28eea1f1c8131fa39da37f3d6eaf4d0b72ddeb6c915eeeb59533ad98b37d550b5f95b0a8fb4c2
z84c3bac241f422bbae757abb832f5e574dcb85d3b50b6aa785100cea61ff59bf0a238659ecfb25
z044375dffa94d4575369918785490a52d6ad0a3cc84294a5c04f9da4a04fdd2c5472dc230e9b04
za89b815876f8310dbcf507a55d135b35423a0c30cd64b46443fcbd1716cf8abd069c8561a2e2d5
z8c6d27b4324ab93fe687d3237fa235b588b277fe4f0a66854631e81daad450868e1864cd00565c
z7d6630f1428b51a61dcbeec2a77cabbe486e8babeae8b25ce47142ec6fe42a228cd808cd04ec41
z3706a9d65c076e360696a0bb545d162e05e714da1192f348109951454a1c812eecd7caa698ee1f
zbd34d0a73004c384fd84c874e52885102ea249b5052e53efa4f3acb074aaa3d631310987717588
z7091451f94ea511ddffb921aaeec0ed5b699a1698ddba2d3b5a47f12d9b8a046089c6cbbeed724
z6631d9a7bd77e6ca8cb41b662511c3df89bdffe16569864f8179b638efff764c6c801eaf95f991
z5b5414208a21862211153c7ec3f0597da2335efb22c251f13e05661d6a3aa431f683b6f8c9260c
z01e9a34b6ef9e34a5918f4dd05981ba6d98ce801b007259ad4d2e2ae25c684459be30540e565c2
z98511840650168315cb03e1a5311358139abf760d9dd5f1838db4dfa7c67adacaddf7ae767a12d
zfdcd6a24c99f310bc330ef2c489a406b4a2f2ac01b1f7d0f1436a1525c3fd4e2f8360ee0349c8f
z30669c249dd2b703a7ce4a2a505832e628475a21c30e729738a6bd51b927c923e239e403be9ab1
z57f47e48488a40ec84253c72d8291730fa24742f04cffed06a6bfcc52a36cc31749a68eed4d9de
z438db947cfd734a7b5a704aae1c8260827922abc6feff3ba36f1dd9d4472d8b75816aec6e996de
zcd78637a47744e729af254d93b5a06c26c10ec69d8e45e86fd80c4f0b42206da25c52a1ec7ebac
zac18a47003383ef0e6956b5abfb6eff494bedb6acbf4655f40f7c3cd6f9d43f243e29ce51d5063
zb8f27d03fc0019afbed24d4dea4a2d047273344af0f29ff606faff099b6d558533e3b2fb605bcd
z5cfdf9a8133f524757ce879bb2abe659d90b753445cb732dade4388d832fc91674df3e39d1374f
z5e5a4a93621809fde8cdf7202f26ecdbfe2b774c4d18b509f76a3c1efc789cf20f5e825d9b127b
z21af3ab4400a5faee454e4cfdf3e6b5f4aa74eaa592d19abe8289a668ee3b67a9d3dfde39d3ef0
z7c2fbea447d8224f7601028ddd96c66ebe4d2d2945546f1810c8c0461555303b157c27b137b783
zb016facb88269bbeb97fd40edae78908ee9f2ac6c5d53ccb7f06578a3a7680787ab03d4df1fa5c
z3f545917b7b2a07a79c22c04536792daeeb64616083517294e088644d4896115b333d6b096fe60
zcd40dc549291ce9c6f2151f7001eb6085e97ef76396340809c60d908668531cc8f49b88b0f4fe2
z21b3f8afc72b15d305b2db88a0239e77512df1ce7f3cac8a488004df652145a7310e30eab90820
zcdd738fe8b725c1b5f23c2b36eb9aaf4f0d0bb9e78e77c0b947a232f4a2cf316ac89f40604a68d
zcdc716b392a12fa3c539b13f2b08d7821b0a2805de748a2feed5a221a12e6c3036d7978838e333
ze6e25ef5ccaaefee82d8a08e5fd2d984a44a0ff349f0e7fc5aec1cc057e96dbe711723e60d385d
z71afde76f2e662b08a01b7c73504bffbe5b7feacb0e40dcdfd399b7951c29526278d2be4cf212d
z41282dd91241580c10b87b36085a1008b2d5048e56f2ee22fb4c13a00fa7e89dabbc80a9527e3a
z669a5a5b9bc4ea295ca614749a367caa2d919d58a22c872a66edd0ebfa6277e88ef2eb2f1825d4
z1e69fd762bd4b1fb73b39ece10118fed5fec30f2d29699dba72997209e99f040b2b968a0ce6c7b
zc4003a97ba562cdd60d4b667d0276513a43a52850c7a0affdc6a577f7c5576532228969791f454
z9c31e7ee8da7c1bf54a4240fbbb56b74dfc0f3ed5eab85f290e7c1e599ef1146d110dbff549b7d
zc5e34080fd8572fd6d19fa2d9e16e4576716ea17162a6d2097a3724a42340a53bc5a5b62fb19a8
zef0425c9afe77b39a4d9faa7a9400ce8c566d15e123f75809529d901954f88762c0fedcf979684
z002965bc85274d5f86918fb2fb9cfe60fdfa20c510d40a6745ac7137d8e79b4fe72f7405c1aa80
z98ae3688e85bd334fe0695018e25c502d30335eeeff5cfe52681549e21316e5fe7f94845c87c88
zf8e1045c8f85e28fe3613a50982311ee985e8f9ecfb3a19fe4c4a84dd25dc8d604cd4c37fd3a81
z48b315b9e6eeff8205f6e16d20a6eaf08d5c20eaa11d9432c6ef57dc9ac0c30167045969393ee9
z3b4ad3af4e723667edece601caeca79a1d351d2dea7afd25fc1c32d24ba9f7908ead42123ac1f8
zacf403a1172a6975b61899be99e3251b68926143d42b33bc3a2da87018b1872141618d76132ad7
zd4961e6060597613968e39201900dc2c518b9aa265eee1c3eee02ff9f2c2f87210480a0c18432f
z6ceb17be69eddf4327988672af3eb5d8e534936a7aade78cc66019edfe2d2f5203e5dcd3322144
z81759138ca03cdc96991260aefa8cdd43923b9cdcbe650fe9cfe6bb32da9859b8b3e87250fd429
zf132f5087fa0ef2415ef47e7255e89958666acaa00322f212d2777058907edd78d6a476a6296b0
z33fe869a9440d9a33211734976d878c29df7a8d9d99669c95420d1082b2547a87725290c7ba858
z6b09f8697c5eb3515b7d69ef8de8fd650778c7dcad20d645c8803a74c03c9815e6e0dca6201814
z2a81b559eff17d2913f0bd966bbe251119d784f532c048329dcb7f668eb58bd726d59e3aa0b846
z0a38a746438bbff0fcfac58f7851b60fff873bcf0c41af280adac81985b49f1f1dd2d143cecb9c
z9c754152fbee156c448d6e8e407d2d16c38357df43a19920f142714d244980e310f2d25179969a
zc1e02d684f890ddc82d42799750db58e3ef39a09b433eede8de1d5e0504a63a6ad557520875a90
z25f048155e72c41f7ae1cd48357c5bfcb66e4e702409db8e11c0976b939ea02f582c8f2eb54eee
z402161f77b71775d7d52bc51b1a12da5130faee7662751a41a0a6a4435b8564c8d0bae32e9ef25
zab0edc2c81378b4f594e613b8115a869472f5b46519ae3703b6769c28a37475a4cf35ec8175330
z74d4dc004404ee7a481d136aa8101d792213eec61a8b29eebec1c48cb6f2204c5b60bb4c2ecacf
zf7979eeecbeb7db2f8af346132b4fd9b7e829da29a371ae1163abd74f9f4b53c7ae516d27ec3fd
zd26faae85d1f443625e63cbfa8e8d1f8cc65e2b9262fb338f935a251f3df19989c26a3f5cfce83
z683128167071a49d9612219323d1d10a209ec6518d58a792343015f8b7c8c568f49b503ca669eb
z3fe21813d7555c58277530763135545531ee00cff042edaa44ec4d66b9a8eed2d8bffa360c508a
z5d22bdc242fc95afcc1eb4727da06318f0c1088d2078b7c69ea696efecae26aa032112420bd6af
z85c6e82f96acd63271d71c9630f9969241040d649f2976b1548b6d40d70d014d6b35cf711b1d59
z1408faf646fda6fa500f247542946695971b0d1eb3f8e4306ed46213589d305076b665135120f5
z9c824ab346cd57e78d2618b2ae48e089da3e6bd2df48cd2691b9973f69aa46666d38b7ca285135
z98fe5670bcee008a95cbed209a4c0dacb19137924ac8af8f18686208221db4daf3af0e20b2e278
zd9a899499f67a4faf21a1f22b382ae670b429b815680ef68f776d0016dc805610740d970546c0f
z88d998c7926b56c721cde5d9f96d03eabd31d46a9dfd92be0eb90bec45e220d2cfb2bb1c39ade4
z72289fdff184bb1db6a03d60631f1de7783fc93926a6a235ea4af8e2701760bb26e80be43ac2f3
z0e72505d394bc7a37f30e7895641b16faf58108b075dde4565baaadb3137a38384350cab82ba64
z2df03b42ee6c46955cd33c24695ec67df25d4504040bb623530d1a778367c12d5e3911efb9717f
z1220216573de2689a8913a809e5f8cf3bb124b6e69bc1bb0c22b2b3ba61e170d1d6cd5d009fe3f
z7f03538824de75a43be4c508508d74894dcbf1aaeb2e10dad43597d41bb3b4b1027878e67da73f
zc5d6645ade5c378ba32fb9b170f6c45c2a891132c2326c707666104472c6ded7ca1f2b331d61cd
z57d17639bc39c0d3319592ddbee44de706245ebd920d2278f812a7f6037673f7b71808d18cd836
zc0d50a4f94b60545af450995d79975c068b050c99772039c005abbeb6a5c4e1e92662c4b805d03
zf44278382eabca6151c54229ea33b3b95f0ec47f4de104d3c36280621936eb8a72c996ddf560ca
zbe57b5de50ce7d82500626110af8d0b2f1124e046fce79da76d174d5f4efe39754d6f8b4ca53bb
zb4f867fe978b9b64563d963c1b7f713960a02d540a4d8244e7a89ec323b8cdf807022e56d8bb6f
z5b74549b6fb3b8cdd78120e82d577fd38972d6d510219b3890b472d42ed819b997c97b45083d5e
zf9073575ea9501862c07692c4f68c6b885f7eea8216bc80eb621497e0c9bf5f7e1f2fa53a3aede
z06f43fa9dd85ecf919752875cda85a424e3a6ac8e2856b667d52eda548e28aa303e22fd76a5571
z9545e857d3a3b9801df020fe4fd44ee9245aa868f3567c98d613eeef66c71be75ad26a53d2277b
zc9c36747aed52675f253351be5a7422ea4320cfd93acdaabb63c81cbd34a0f2daf6f5a79a6b186
z87e48858a030c68cc91fa0f31deffa3198da108d49a6c7de8f1e63b068f40336231ec0e65212ce
z75f336828a71a1f75ee0608919699057811745bad45b80760fe890fb9d8212f3b3cddc5f2764ca
z22487642d708059fe47b2fbdd715cca77afebbd002532256c8163990a32f13cf519bd731a6d0bc
z49b27d0b1c0060d9f951cf821cbff30bf7528d729d55f4bc1d799352f1455c5b7c20ec648ad71a
zc29a0b5709c0ad7cd3c73aabc323798ec6d83cdcc228f0e1b1394a7cd20efc55498f92e823073e
z1af275a4dd8c13ca899f44752dfcd2e85bed896bcc42e88c94d3c8fbe4d3d706aa13c45add9c18
z72f7912741e3a28c2eab080385bd5ba1a4b89342c3915e19cc4a6e34c886f827f89c1e033391e1
zf7af3aa16c19fb7ec49a996a20b0425646d5adef48ce79fe5d1ea0d73c38cc343d22d920316437
z26b8638a6545c09c8e3ed5cfee2617b801b0f19ca428d41cf1ff2a54d534ae992063f8c80ce98d
zb0fe7bf37f357e5a119a2933432f6298c2ec90f48f4f6bc55404365a3adf220ef8f8a451d75c6e
za72c1104d04b2170a71eb6653531c8ee9aa6723456f5345d85d7be3884f28d1d7b105db730ec46
z522286132cec41439ebfde36502671a68711229dee6efda28a9f15567db3ae0044e4c8517400bc
z306752aedfcb4023242c72890f2b51ec59f25d5d001b9b567f76707b3fff34a64a8ee7fd549a73
z18245536bd8653b74cd2e89a6ce1e29990051b8b4313aff570357a1e476aabd2a0fd2fc135ed00
z7118ef73eca730fd0352e50209f1468b79c694096b1d8bf4ce9373c5936cc46a4de992eed1aef7
z1dec17b11d6c613669f06addb8ddb609e5da5f0209e41a83a26ff3d5782ad808cac5f2b2bd8d18
z08961de7dd277214697ea5cbdbba348752d1e51b12a1cb7308dd3a51976d6abe571c93420653fa
zc30a43bbce2c83d68ec8bd9ef09eb993cb032a003504646aba4080958d4934ac79e001247317f0
zf215915758d8e78263aa93d1df90a1db8eca4206c9cfabf3cd2b2805d3562c1dc1ef2a19680bd3
z4d9c45b6e5691c635d3848b291eb5867e98211603db5eb141a5c0acfdb6517286ef387615197e4
za1dbc020337c0110ca9635056ab16be944d2bbb013818960c0561fbe087f9a7641a13b2cf7b560
z111cd560df7245e279ce576ea0ea8207660fa0d4e0a4a571b29678181ced91cb7d3a4a31f7fe89
zdeb1a173ed70c6e89cbe9fbe540a9b1ae264d886fc0c6af34336bc036f6ade529f01ad256fd2c7
zb9dc9386eb4249f834677363bcf1c3c478a37cdc29e30109f91eaf4c76bb5846e42d325ab66daf
z78e3f57f809fe9f25da562b2798944adbf9473d91229588dbbb3f741952a4ba7322bb9e3206463
z3156c8f33281f684490f67d6b5e5ca77a02cd96dbf7d9d3672540ffeaef2ce7c505e219a34b031
z7a4bbbadaed053f70acb3afaaaafa50de48f31ab0ef7b20f967ca5556f78891746fff6bb7cb428
zb007ca9953e220a2e5b98b86f8c046a8ab1b462d51ca763b88b6c2d49dbbf91a47428371d0afe5
zd684a0f942ec807359ddf30903f51238e6ed3e0a374c961ef40f86933e3acaf1fa40d327b35620
z9ae7a638f2a4866fe7aa1726e913d3ab080e362b8a1a55dc014a47a04a4a287d13e5fae11a5132
zd26bcfaa00bfc85dd7aa9ed3a1e7e2cce238b63c892783d69b602cba79cbc6ea2c7d07f5b68d3b
zc194fca79008d1d063161ca4577bc356aebe1dd055cef4ae6be45c4b8b3448f15a6e88c7077ae8
z7f93c3e54bde0cf4432a0de5e9e2ae013b7e293860bddc316b720ff2d101d3121e1ed0675dc02e
ze53f66f14506e3b4b08fb1a2908a9ac8c347a15cc9fa9c50de88b5416afcbcc12de1fe87f01c38
zdb10e1bad4a20eac7b6a8e6088f9f58a1763647d7133aa9562cd17993714335497017beb1ccf3d
zdaae291b9a05897bd0e988929c26a847a95f8f713cc06144ef83933183707bb36bd28123c9f3f5
z0e9c37e4757e868935d1f4b830fe26c4f38eee6078eab83d6879d852f87e55e999d3695f9b24e7
ze1d36b3f759a921a61327f13a48771148fdf303abb33ed4061b250c8895b678fd2b942ca997d21
zabdf134e64026564545bf27e7971cce5d6e5cdab2b6451c6102b2a3e7d146ab9a21054bc6c4146
z1b1de2bd64838f835581000266837b0e3fb10360b69dd803bd70e34d1f20a6219d9b826d0fc9dc
z5d64aebec1f1bac30d08d7c4c1887bec46870fe6cd80fe22c9498468cf15c78cb2b4936f756302
z63ef4d1323a4597c1a336c6742eb82b4725b0b39694d3ee90c3f81d346c74427b9e4de4e19fc6c
z27eca4a27471cb76437d9d26fe55134d4547bd6a045c4ab0c6b7efcd5df7d83434e443afe5ed96
za4a64d78af0ca2861bbeb79ab6d12375f2d9a62e54a67d61b95780068313282cf48b1f0675d8a8
z122d5098f2264b454313b381f1e6a65602b5c57bffd383c2b2559acb7c9e5c179941b96f7bb776
z72abe051dbbc58888e9feca9846fdb1ac2033a5fad679b93a86cb2cef8c5508f737b009a2ae78c
z6d2f0cea0975832967fa3f80447f560e954a4b4205690fd5d564131cb27c4632881faf49d52e00
z18dd70fcd2dc780d27fed78f530b0c47e73afb1e25dd1143d87178c47e18bd5a8abeaf74460b46
zc2f962346a55b261982ef24882b7c8b895d843f6c8924ae73357580a6e0412d6e37072dc4aec98
z950fafd5a38f908fe94cd516b8e7567306575886b8985b4c841d538abdafde9cd754bbedd49846
zda8adf2cd07370e1dea36b92113f56342bbadcdf4ef0dd48ddc5c75772832557c0679a2b54aae4
ze5f038c12f35307bf06621d00364999e8145128ff24113aa36e5ab0d7cae26825c39fd8416fee4
z093efe37c128cb5bfdcac507706b3c6e1c6010de5a0a0b537f3b72d0079c9aa883349e053bd33c
zb7a168a24ab778c92c58fb4beaa09fd44c09bd0ee0ced4308309de4ffc0d190ff1316f89ef7a84
ze9d35e121fa5ed47f40988edbe759788b84207d854fc8ee8d04b6a27199a3c1bcdd8526ac38fb8
z75ddd0a7c57c52c8a3af9aeb4eb492a70d30e9ee5a535d405ff440b8cff279385d8e3a8f3f1217
zc23c11651418a2ba479ede1c39d6530501b33b13b9f74b9055a95cc49dd30fffd7a3a33706f60b
z1b00e80b729429fab1b0a1d5889974744aae53c2d1e6691cb6f157d4d77a9830cc9566c99f7959
z0d19f3373a4215b7cbcb60904523595c9578290d57a316e8efab96482776b90bff506d78f54efd
zda0429ce28a15891749f0a5613ed585d215ab317fb71cdf10089e697c6bb84d018b75866adc22a
z3536d0cb0c945b5b02208e00c193010fa902ecb68b5b5e92498f79ab020d0995577aea480b3846
z00c035bba460f1781036b9b4e52b984c2e330120f60aba18480b6e05e50c7670fb5f941f80e070
z514a9297826b913828bf60578e09d76067ff1768651000ad32baeb7446236e8bd9e5ccd1369b9e
z729968c672ab0545eae94fb9f5630d644adac145e531a7bc2e8c3e2ec3dd2962e5bff0e3c80559
za17acf520e1f70f40b5a90699aaa734844f9ccd8315953d8606f30937e68b0c9f97f365446f03e
z5761f554cc6d4f81673d048585260be93d3782929c86ec1c6a50d233b24c37e7ee67a79cbe0a9d
zb94c8fc792a940bf85bba50b6e88988398325ca62a0524ebdd2d902ff90f416f75c422b9bc1f96
z7b2711e8f7b19e98877e0036244f6c04e4bea848727d85346db7a866dc51875ae48c36936e21fe
zde1425d2c6acccdf61b6a8d749527aeb74e63f6452fd747fa7d18655be4c630cb89e33d730cee8
zf96e5b0fb3d919f57c2e3e95021a5fe48c6736060ea86f5b794d7f73ba85bb75e38d760aa36bd4
z677c1a456ce1d0be845b747953a69396712ae119660b184ee590fc1068dd4c987c0995b599c5e6
zb7fa89f542dc22a652973319bf6e421195689b923d1904e371c3dc6a7b1ee5f7a9d10686ab3f51
z35377c4ebcf771984521ae6671108539b0aa5ee330d4cdbd85d44fd5ea1edd62f625063c78a22c
za75b75d345ccc4bd8ba3ffee00285167add5f64710e23101479b12a41f207ff430e8e0fd957686
z2852791526f3db2772fb412e01d1960fc56037f1bbbdda81b6ce89fdf61f2f0b8400dc0c49bc72
z5f5cc71e207370f54d4312e03cebf0f6133dbee3a090a2f1399fecdf6fd9f7f25e5431e0d7178b
z0cdea637c86d74f478f524f6cdabd812458014964b5e6cb11aea3cabf9df518be2ef282172612a
z121a9fe0805d7d23df5c55b81eeb233ee9fdaf085d0e978255eac474ad0fe82a59e2b8d9f10979
z1657883f5ad785b252c48aa3838e9dfd743641c63458c893194860752a0e67b14ca6061c8803ae
zb5383ad005db12dd4b0ec23de3a9d5fc39c761c8771406ede8c70945d7e0399c14c779ad378180
z9224167a47f9018440534ebbd44492d388a94434119bec4aa21da2b024bc6a95866bcc561b93e0
zf71e382052153a1c8f84bd01294e7a3d6b968fceb2629247f76929f36bb29e079c154d65ec5047
z630386e1fd5641eb9f57c6615d4e16dfd0a8cd79d758cd5ec44d8886952009a728f29fe1c8aa93
zcbc4a1f43715de028595ad6ae23e7372957f88944f76b4d06306ed34b9967a06c490937de962e4
z0d13407a4b4c05cfc1b57803627f9da504daa893f38ea2a1c5e6ab8840eabe031a17281a4cd549
z7bc611ff4578612373341ded09fc9c023b0da622df35522ee88971d5803de51cd38548045984c8
zfd1331d81b7ebb3678a23f15a924544d8d39a17b87df1ddc6f0dc5561826b634993caeccabe92f
z78fa9c09dabaf39afdd9c3cb4a832619ae3044e8f149deb983daffceb6c7c63abddfc45005d7ca
z84aec52506f6063eabb31280d219524f3b6d69fb0b84f91e02208c4ad7ce26f46fde959267a96b
z68bd32b0bed07d5afc3d9e3ec86210a345d900e8e033c3c99ebfe864a75cc6ac6c970642984759
zea62ddf4dc5fcb4f4ec5ceaaf7a33be41a382b79efa65f30195bdfbdc30513c580d3992f51bd8c
za516567c2ce3e401ab9a79000f01b55736c02937f629f0673391f34777072fe95efc3178d2ef7b
z54c3db2b6f7325f488043c7a5ea2ace3e821b47787503acb8a04639d0cf955af5f9a3e0c3306d5
z00d0ee724bfa6f2591824d31b9a124b142ecaf47d9498c8127258f2c6935b195ba4c64620add6a
z6ee6a1e857554b33af8308ec0c5213614d98788b5219967507a17ba31ea69d52e83ffe7aa8c443
z9750c9e263bcf7400afbb6c9b3568833c2d6e0bbb5eba38c2e966b9d9b57912d7f6440498f9274
z4cf323648904c67bf4c9bf923b3d18469d144186e22ec3f9c3e3a94bd330230f6befb125abf889
z61d1574a33ca1bb2d7805316336b796588d8a80faee48f80533d54499e7ccb3dea921c2b679915
z3396aa98b0df46cd7c6c39ca01b8507fbaeeec593e333476f56263e540af0244e49ff534f7a61c
z5b44b230c1e7d839ee315b2c20a642f664785bbf3aa607a897f21de8f70b36934daab22e58ff8f
z16f83ccfd921b7116463842effe67bf46802293fdd647d4cbbd973501e6167485b791f132437d4
z91c60bd80fec65634e01b758260a6d13f57b021529530daed453e9fe5ddc7dc9d0d67e9d2f7927
z7e9a61163a875349ebe1eff5050bb5e4809fd123afca520edd396dd472e41e121b9990a53b1a66
zb88480e37ca86c988a629e82dc847376e81ae69967aba0e51214f45a4446a4838867de1e5ae676
zf36a92d252bae1bc0cbb03fb8efa7fc9a15186b2f2f5af828d1c71c7344f78843b78ebca4edee2
z7d0cbe2b7c6b3d51465e11de61a02ac10a5861eb40101056ca82f84638e7d9b567bc917a7708a8
z04a28a6fdcbfdab448deec9c8e05458de890b322b4734034d2bf4017cf7cabb424073e7d2d6972
z0fb01bdcd0bc84350f16559fd2d1fb62e360593a1f1c76d375aee996bef6340314f6a071b4af30
zea38ea8d830a981901fbd33e5a397e840af426fd0c27f3316916fd6dae80b1fbd9f55c7c72e2a8
z24cd95c7b0dedd40d1292ccfde34498e9aea3dd5870ca27f9465528b79433270c2170a4806792e
z31d0cc3521f4b69afabbd428a9551fd0dede196115f528c9e0143bbf9f8f1f051a985092df1e5e
z9040bc042e935f187038694c63d306d06d632f94b8b20fb0cf5f2aaea4269df825d71fa1619ebc
z8d4035ea75f753c0e129f6d95981598f143761eb0f115b7f4ea0b72439e585e6f4cf0083d03c77
z3c1adb6f8f4a4c41f272c8263c02bc7c7c0d30cdb987989628d3de0ee33b57214782c0e1dc8c17
zf8a6147118d787f8f1c0c835cbe1940b5a9fa97d935d88976561dd2680428b70f62b0f421982d2
z6741dcbfa8ba35a9670e3e8dfdb86fb617f21506690c119fdfdf4c56985c4b09189870971d94f8
z9f60be2b3e115f889fcf45edfb787adad3e03653a85839ce8a3d787baa14480708ee681acc0c25
z11437346fc9535e0e20efbe11c898e96ae04a24b3eb85c60b53675dec9a5f32e641aad28fffe6a
z28bd6b4b4bec810cf995eabe4a5268debe22e8748817ec4f8298ecd6e79316816ced11ceff871f
zd6cc82e69ced1fc340a9ade12c1847fbc8f8c208150cb5ba8a9e971858fd19d31e7a3623e81aef
z60612ac5e638de29fbb375d5e6f00f8ee18c1b5e0393982ede1c9368f10421a754e002c0699cf4
zbd249a537cd318cfc62359d97161fa37529139d48fe2fde5fb2bb3b48e1d2e3fce3af2e89a6b9d
zb7f28b0d1d4ef194d728eb1d91818ccd0368b335bb07ae5dfcec2a9dfdb4a9f1ff5caa61317bb8
z33a089277ba03e7e7ea5530d03ddf3cfdafb36569d5175592b28c748187eca87375608cf0508d3
ze7cdadaad121b2e3e4171ef897bd5110d18f00a19f0a3015ac308ae4a28975d6a97910b5f2bbe4
z1ca8e45f8d4d93c97c7c018efdcb83ce3b948dc1751b1710f70953f3663f535a9c3d32602edb8b
z057a24e7a8d015fe858bf0d0b7c0848063f74159b8cc25deef9e859201cf636feef66972a84d41
zd05100831173ae757d5b2f3cea6b572bae93d76db5fae1f853d2d7c7e6a52495ea63b4ec13c90c
z743d9216fbaa30ffaaa9092ce0d49bc181f7f00d022027d7303bace141afb74f2da5b76f8a0b72
z2aafb027c03eed8e477d6af9b2f28554d76cdab34246e0fe07be2af92958c57a49b4ead5682564
z6b860962b28ae9d3f90ccf56fb96e1c8ebc9709860f1aef7fa91fc7feaa323a468b2314024327b
ze8e17af9ba071196f0ac1f1dfb315b64025f53a8b66ecce2a6d3cd1d927077264d6a99808cf756
zebf10ba3443a71228b5634c6d6f02f55e8ac92f47e0e854242e2b37e7377837c32eda6664e7ac1
z94c0e7f5ce757ab97dbacff465093155bbc348b715e590e8aaba9ae07446c13d3c20cf3e006098
zb045ed00067b4588270d90675431851d2d8f489dbacb5b072db36d7591e3bf7e6423b523cd9dd6
z1dbcc49163dc5a03fd6d7060f59eb3f5b8f90f228e668455e93706f462be9c569ba4050b7a73e5
zeb9c7b4774698f608c20aba8fae2743071f8d435ff56e95a3d8a420aac238fb710bcaa88177c56
z955e45960a7ca1a64b160b30e23092d4b0a91d7c06b9afe69710e56650cd28ee4b917d13dd8c84
z781463f1cca2747b2755019591691b04471163cc441426b04579942cfa13960ac8a605b5019972
zb944bf168eb531082df6bf9cd9584e1d9ed146c609a59c65611c567b4e7d8a86aebfc23f7d5ad8
zf07fd7d61e0198c285eceda3c10e20e7e3a42cd4093951de3111ddca8c7af9d7caf41e88c52f1a
z65d4dd8700436f30f128ee1aab1906ce467f4493feb9b6a281cddcd88f9439c432de3870403a86
z05d3490887f57951976f84ba69982df441368182648b9c4f42588fd6153e4137db9f5450b3a0b6
za103354909e4a73a1ecc1e1ec95b5509b54e914c5d6eafbafbd3142efcebff63b03b4b0bf88185
ze1f3d30c8e799e824b6d704d2b17df2124db8f5e1e8c1305e677b9590abbe43209451f832599c4
zd4e04a0bdbd423c40d01001a70d2c01019417600f3f6eb41a4ee9eb3f8d9f498e6419d9d8a5df5
zda6a63983db802ed43e48183d2e9e24feeea5bbbafa29896d89793beda7a4d3dd5b340ebe24eb8
z02801e44b729563b3f927cac280a1860bcb4a59f8ff8358c94aafa173826d23b1196a8d7230a45
zc83537060fc0d175eddddc343e0f3c1902685076541a4952b520b03c6cf135110b94e078d123d5
z5fd3d0fbb1493e3f4960bd44d9bd43044312efd90648093829f5e7fa4bf67f24a343e6d339b97e
z1d354064902bd2fbe5a3231626e13a6f591ac8e93e72e71bfefd5ea3649c57eb15be22c00107a0
z5fbe33cbe7dc72675926bbbdba99758f96b6aeb3baf90beafac6009cb74269a2910d6007c2a92c
z9c7b4623a5a6b41cea7e468fbf813fd7828d62c2550c2efa6194e55dc493bc1330668ed671ca89
ze07268bdab72c89894d30a6449e5210bfe6b3cd1a6a44595b9d597c51003d24a4866ebb995b03c
zeeda7bf0449e5150560bffea5f8b3d7b6c145e13f323ac3b1af034423a3c7afe4d63a014df1235
zdb778b57de675d824967918ffa111898f5bc6036ce05422afd12b05fb0e4710798e27f7a8a6769
zfd2f3865763f30799d70de1d9db875f7e3dbbc164f840d72d789842189a737997e21bd29ce6f06
z5d56de145984dc4d670fc1632565675e3c21ae921f6a9acd1b35baf1ea37f87e607dccb7fec4a5
zaa9af41645fec5d10ef7be3f1d204a9d73d60010b84287e8f3edf1beab98174a1371507533a1e9
z31d10714cebc91eb101611e228187e00fbdf8be27e7c7488653f7540407fe54b9c0b4faba3fb04
z368db30481266348ccbf78d3d7e048a8b9f1cad38b7737490904990315626ad88a6431bf21309f
zb168cffa5ca70d8ad99f86daa0b0c05ad5c5e2852049cd37b856712722ceddf6ee063c416115fd
ze8d37514c4af3307a03e53d82e5197302488413fddc09d8d50af500abdc7878577a0454f20e7a9
ze20526a1249db43e78316e7c88c7b96e0e6f426f141030b0b062304a3cb6bf25c64611029360cf
zf9a0485b00e3ca820a2338275e6b85049cfa395e0b2f7b0525324356319fb3a5360e82eec080a1
zc817a83d772e0a8f82ca65b5c4db14dc69581c5da506505cbd56a9c3fd73deb262181fc3422dd7
zb7e8f0ec2d7e3ffd7578d8fa14da81331308646223e09ff2af376a85fc8959a8ff554c02918576
z77e3f7fad493c3de912c4f58b4c20e886712d27bf047693a1e3fd10a6475ecbacc3da2084510da
z5164a92d2047cbe268504e56ca20df2dff2c7f668ce3c441854240dc3f200991682cea9745f916
z87ec623561f3791fa67f52c6128d98c4a74bccf236a291873d076064af71c66993d2ee8059cb93
ze2a05d05d3f3a0643e6a725358553e28598847c7200133603f35835536760db141a7bc8fe87a3f
z0d3a6a79473715496563bba34197d4ff39e92f389351a304fbce5a8534d8cc2f96816ed9082896
za2936176c323216d40170bd165060ba9b824c270bf8c5d03615a2109be8829344c775e26e750e8
z14599e3d381334fda17461da3b69675245d086db50ad6cdde43cf91000a1cf882b754498d58e30
z7ecdaaa34315c7e12c0e977ed2e554b1c10f20041af1487dfbd4073fabc4c406e7cc3d0a505e0f
z619aae55a3c709ceeee1d18731fba9cdb628c2e8eda5c802e9decf8dc60cb3dbfd823fbd5246bb
z1d52070e060f14bc6ba1765aa235a0e48dc664f5ca39ca86b7e920fa0a4029e68300df0b96274f
z1aef1a75c1d066c5a9083c5c6e017a66bd9e2f7ae14f8340994b5e0ed9072e60d1abf7767660fe
zda5298b4012f4f09c6ce1c4e785f1fc9459499724371c7cdc9625d85507bbadeacc8033385a794
z053b734d86e48d28c55f7d3eed04daa3fbc70276f9af2eae31f9e0fbe8d57a804de6c833281245
z6bdb7bb792d0fff769d20a055e6a045acc948494b7d53996305332885ad630f703a015793fe90d
ze00872c0ab96781df08c6c85c09db53535cbb471a590aa0d176a9b144dbd08c64c0bdd7e457164
zf6abcf95369af94ecfc971d1025e18f8e11962e8b9a21c6f8b72d55dc0d626ae73b266c3e2d878
z2679919176c46a222e515405bb213427c0271341597fa3f0edea2834f05e8037d82e9a7c624152
z91a0186e8965113ba8585892e24cd4b3eb68b7bd58232298560ba1d2bd70f1b7ae398e4e0de9ac
zf63423b4dad87bedb7ea83f36b3214ed2c51849088ceea35c2d857bccf21586e0b51c6fdf88009
z140d16758ede32495f2bd3c8f59741059b562e47e59ac12b8e92933ef37eeed02bff8dec4b0af1
za7be94d20559a102e61c8f05e610bc3914b869208be003fc6ad247441cbc7d38468005915bc3a3
z6edf0831967e312559890b48efaf3f4e170decd8805fa911749723a54596cdd482b97b3aebebc2
z7f50444acc82bcf40a6af42f059ec32fe75342f6cdbd9dfe900ca5de947f0d75b41509aa06ade0
zf6df72f6bfb216c95097b393766170a522802e0280e91f02764c3317749067d37f243936c5d5c4
z9e809790a0142ee82106b52f332602e6f0d3532b30fc6f6c2a51c616dcfd434ef0273576a8678a
zb909aabc2b7d006637373ccf7d100989852ab200961883b287856400659dedbfe55373de97809f
z694fe0bb29529e20a3ac85ff4bb9f30d4d5671da881ed59b7fc69c3964467c4c10d0443561bb6f
z8b1de20a9c2c20b4e187ab30ae4dcd4e4eadce2bd61680c4f46fed56fb7d168984e85bc102c885
z57443947ef2ae33bf28962674f48af2664dc48028d6699bbf95356ae04b60050eb6836892bd952
z3a3007173a36c452d1a5daa2047cecb9bdc235a91e5a6b76c26e53bfcd0699cf6370cd90c8e848
zab62cebebac57345f91298b486c88c19f032c2adc565c038070cda079989a1b688d1ed68dd3f98
zd8ab256296a24654a080deac9248262b94bf4afebd20f5a7693082d7279cdb783b887025198815
z67af8aa555197c3f89d4efe583c8dcddd0126a0ebc07c2eb33a89f97b76fc1dce491f90184c01b
z3e3bf9513275fa162f6ace69850334118668cca702e037704491876e520c96ec8567e5aaeaf930
z46274f9ca624901c2f906e622e200caf8cc4f01dbcff4520575d6eb0c4881fb6a10c2a5ae3add0
z482df610120a2b8f324c7cfcaafee3fc5831ead1dad1236a103d1fcd31ced7acba99954088e48a
z500232fc0221dad9f96828a35d328c5a65a2fc66b959197552089f57448fd096dd31a1e001b73e
z644b92490743f9b58fe75f7d3bc1c1c006b07b17b0fe1a7544d15727fa5c231e17b350769ce785
ze3b234691e2d60f6cf25eb5cf320f0a2aa066ff54d1806d6dbfcebd98604646df519585404c94c
z8ca5f56ad623d8295f7e6012948cda4200a1a46ff353e5deddfba2775a823e145f2cab5181f819
zd8b7deb7ef87a71d5f400d355364bf42d6905831fe4f7caadb75e9e8eb5e4b686e3fbcc1e38b03
z2851e214660d7e572eccc70c5959d83bef20b1f778440cd610a1d413468e110c542be714dc79c7
zc79036a99264f3ee62f275ecb66420beb445ba84ed2d08c59f47302a7b5803387560cb92db5c02
z7e5806a2982bc631eb2b187357a29752ad39076afdc2bb372e4c36952d891d391a72477ae694d1
z483957c80a677b6c89ed84fd3bf66b474fe9b6be8f02195d47137336e0eadba0ccbd39c9fe4d69
z63bd7bd141297023bfa139acb67b9266ee5d0cd0646ea02fb230553aa88494d869a438ac4f8a3c
z4a766da472f05f36472cf9e4dd29fe2a0471b861e6527bf468d7370af3a96d05caa4598073ca24
z0b3d581b4bf9d06e9e1195379ed56ccf9e55de87311a61b9604a35df564147439585a9d893fb6a
z06d8b5d641b6f75a4277d492858798b4ae6f9324ab5fff0a209ceffcd8fb111654fe66940d2228
z9b8bca77b0864bd598d931bfba3ee801ee40b51e34120fe411f0c68e8db56a13bef20311144b78
z2f49d660860cae6e3ba31d5f2c746d2bdd6e761e5f8b94beee4bc00bd969122e69b28a14763b08
z155aad35d737f4360f1b266d0a46329c4b1100a41875086252bca00ffd161f1bf4e1aaaeae2ad3
z7b1339b4d7ea943755cff7a9bf376955f8d1d2ce9a7417fe983777c1ccb6aee211c83857caa2de
z6480f8282fbd9b128d9f9ea2e71b3e481b29585965364bb226c55e74aacadf523ad73d5a91c8f8
zb761a8913ad34a2ae18d1ec45ecaa6936c38cf51620746c747cf591743912b6c3877861ec0d368
z349c8a7d3dd77953c70797151038e9663c3131a758f3d8a30e54f81cda47e44bfce15653f11fb9
z72e332bd8488564d8e2699d58bd6e4e97f20700da56149cb69d786a6b5561ea0a7b07190e8f29e
zfeaaff4afa665d143a1ef266496c7cddbbe932f35dcf1235271b1d5bcc4634ca7ed9be7e69afa8
zb73185af588ca325f7769fee33efc72c2d7353738520795b60d4eddbf6aadd859c81173dece43d
z8f275ef7e0fb35553684af191ed71a35625472860902d1f7c5977eecc62ef4ad7344ede617d0c6
z882043e8b94c1eff3506f6184c1a595e8aa7f48ecd89241525f87da0539da0caa34713fa036e96
z2554f4aafdf1e17438d985e666d0a0ce980824ad36023a1871aafbfc71b8f3de97ed468cbe6814
zdf8c010c99cb00ed123f32d09b8654367e40482df14e6714b4ad54b1521da8426cc8f24b32678b
zb9907dbfc03d4b14acdc4231462731351c4d03f22e0788569ecc86ad4c869a10e2ae843493b7d3
zde7bfaf90a53c4246a8cf8eb7fc84fd0f820abf99fa07b353e107c361a9f55d605c1bbbcdebf37
zfd11a0d3dd53268f31b32e8d34ab198b565fb94645e99f450afdc65e4854a6f271b01c2e31025f
z9d231404400378997f686c6a4de7394f30ab8e8e950a73d6c5d8dadd78aa35c955632908e173e3
z3048533214b6a006cb5b53caaddaffc18f51fd2f7976dc57e9227e816e36ff71ce14a31ea5aed0
zd8c3fd42a72208fa246002cbd105f39b46df71fb03a401c697156cd3108710e438d176ef6908ed
zdd7ab44aaa25e6d92509a0c5bb8c79fd0c433f191953f7471a78ed31c939f8c2b2ac269d652c13
z944a85a408b9a957094e97648034779b4a4246f254250719f8f30791c5d5a51fdfba4866f9e932
z5466b43d1029371a912aca0dd92baf99a28becc8dd3060baf6344ec6ee06674c1fe92ad2816336
z0ea2df2e91c2f87024a135eda68b1d721cc16db25a716acc0faf9dc8d0712bd8121a4f274c6b61
zf5c67ff828df825c05fd863e069da655e93addf62b14905dd09d59652aedca6d26a71c6aa114eb
z345d951ca11187fc6332bfe0983f8fd7394f081dd710dac80e80fcffb6d675f320995c4998a5a1
z8c739e00ed9109f26a9d1165cec4cee5ab23ca0365f9c661e69929fa7f737c9fa438985cdc09b1
zb2d80138d1a96365fe0d3ae389509882e222d4387a6b5360c5edeac1e73e67448e736b26067756
z5cf2d4f7ba44ef58ff16c6fe2e6586edcc5670f35b21e0f18926fdc452824360db22563cc1fe3a
zbab9d44e643ab9f06ac138ab6c3c75b37579b3c54b3a52e0f485c7657c2afb2259caefa6728cbe
zca6e7faecf2c6a3a76ee2ba503f9fac90de7ab1d03db1c10adc61bd629e97afb307935334cc1de
zfa11debfe4a45740fc52ad0d8e72aa70ec0e9df550062eb1bb9f7e18e16252bf9eedf954feeefd
zccc065d85696d2a0b99b5d054b5b0189f7efafc19a06c35bee78bfd502b0cfaccb3e99d3df0371
z3630b7ec358ca025138776f95788355932733c8e824598540d8499428133cef52e9e6f5bccaf5f
z47f9874ba04b0c552fe02f7272a4f5217cd54ca4856ca01164a864211625956c2200740ee4a0c9
z336445b5db8d99df0fa5235509c9dc5e32f4e2048459b59f53ae647c59af1eaef7f529911e9fb7
zaaaf8d3dd42d28a589d1da61b3ec816fa17a1dc4bcdd455aa4cc058f7eaa0a5d20ca2461c476a9
z0e1c2fc7479af3baad0e2f4efddf31360ee4efb9b6ea32399cb9ea543d7cc0867f4e8995c4bae3
z469cbf9b319444ba9ed49847d4b09be5f850f2d3c9b60f5eaab5fc815d9095a354da65ac9158dc
z6256442fd711601e1d18e44b78d642c42a358f7adfd2ff6e951fce893e2202d4c8506b60a1c9dd
z86ffd72b0057444d95b5a5d49f5beee4b6b2e65f2d6fb9d3bd1d4c4efbabbef0df93469e68e5f5
z473f06940e58690e70ebd2f4ada64524662178560eb3a6dc90092f9921b15974047e835cad04ec
z22f750a0547563650a829038ad000eb78259b0fc7f6877a76c1aa534a2f80c8fb10c0ab7bd1516
zc0c25c787dc95c2bdd7f172a5a2e823ab5bd94adcb08f7c3a6e0910d2a9fd34998cac86ac4e36f
zbc6e7fabbe48a7c8cc54f7a195605ef274e045356ddf36bfebd1360f29b476f837cf87fa087c02
z1a1650b4cde502068034c6c594d4c8c531fc93db6d8de1634feaf1b1891b7b5ac7bf8014003d74
z49b5e510a2b9c6243e600b05b6e31d8b2988e1e82d213a931efcf7d8ea0b53630db50d17650357
zea13131ba5f2a65d0d135929f9be34a997b2d3b367c06d97a6d38d368d80a495b93430da442fca
z296f8ffa195c0340e17d31b79c3180a23b5cf7db84b9363a3eeae63e2d07ef926de635e7ffecd9
zb0a6229304bf90f800b66bfe3dc11cebab581caade76dd769d9ee0aa1cfbffaa4a3df41217b37f
zb990ff7a4951daaeea1649cdf56b4b96c98edaf0c40d88dfc48f5f6732d8f8439023f72c969699
z04cc6cb312d452ea7e070b814336854a2c81a941fbc76d9a9eec1040a1251f9a37bef36dac33be
z99485f79c30594053675aad856fd26fc0cf1518476058fed68c162f7ab2a4135e1732006e67e61
zea2c07f947e7e7e868d59037ae63c9edf75c84ea9c6c9a645e2e6c636bc1f67d1375126f2e3402
z9c5901fe08184ba5dd1415d349caf74a6b54258c29cd3d0e678516e81bbbe7a8aefb93de674478
z0917040a39672c3fa743606749cc72806d15d069341b0462169ba6f3dd8b63e7c2dd4d431676fd
z6559524515afa18e1cb90ff12ecfc26c7dd62125683d703e4a39b2c0c3198a889863035eb5329c
zf116dea835b0e25f0319bfba84b1020271648d0e711f90565246ea7e4a600a533153da56168224
zea78e9d6858ef48b49f9ff34884348375c76365f4c065c70763c624e9254c1a0ca5f58dcea3a08
zf264becbd9afd5d80da4324836198a0ca20e9f63e65f313586358fa6d0ab6b24dead34c38e2cd3
z6696d01fe41418cc275870179a6a12ccb141658e82a9396cf22e9ff714b01752dea03e7ec706fa
z88c1c86ef4b62586ad7787a5318f6f4f9d1426d5c74371be25ab17fc48a7fe999755aeb338eea6
z477a09339b57caf6df5e74601f9de6720dbaf020b3415d8bb782678e653ee800b51eba46ea7017
z114cd9d4a89b98794e79bc8d7689044853d3ecb0780d413286ff9e368a4f82f6b5bf23be2d2cb3
zdc43b5fa89b61c4d3af3e0baddad96a9dfdec68f1730cf41404f1de4f2dc01ba729bcb10aaa64c
z49f5b4365eb20c871d210fb0263a73768159e6dd2d810048c39fcb209ad3bdbbcfbf25528207a0
zfb2ec3f284536e7298181c0ca356349f620a5fb1ab0c80706cd70b1fa67453d7484d4449fe844b
z71f04e08877fa8a55d93d9856a6b4122a62215e36a4644c3bf5e6872a7986218d1dba0343bd8d4
zae0fa28e43f44ac535f0079c72b6f436631768441ca709b34a5d4ebc3384243b19ab07e8ae8841
z49a957a0e4c65d54f86492050d570b91de3c1db71313387fb16506bc2a61fca056d989507a147b
z2ddf507d7745347c75ca16cb3c0a8812570d7ae431faa87c7699fe8ebc19f091da941d7b11637d
z50e11a44b42d67fc257ffa8aeb175c8460e8ea6bfcc6b70ffb1facb973d958e6d33ca5468c786a
z62d8a002caf55c849e54afc92149162d18da26624e906d56b137e38676c2781011ac82ccbd2068
zb8c66f22d194a8a9b18c6a95bdf804b6ef35ba792746bcf99c44f88a8d440b9b75f9be79564328
z84bcd9270bae385ae0a34ac160f73b7329f7be62a5bc994275ebb705ba0f50d7211ad38b559d7c
z85b1741ab92b643daa41c875157ce97c8a92cbfdd54b6bae47d5ddbaa099eeb687fb563cca7472
z5314e8ab355df0000b95e239abb91b7a79f2ec00c6f6c536d2657f5d635205572d9fd31427dbf3
zb4a96ecb754b05a55685f2fdb800aee5df597575aed7659ec24a4e4c01010e35f7ceb70513bee6
z227a6bb69bfffe198428494578087bd2e2ce014de2e0d068a0f643ec94502f36f2ccd0ed128854
ze9be6da2ccc28d849ed30bbf7fa509622c31dbef8b0e58a2a396a0fd9cc8811d657110427b52be
z0011364e54c3be00e09e2a8b9766e69ee97481c9a90362b0f99e367f3081385003bc93d05037c6
z8d7cd7dd56df1e97db15977c4c253f940fa7e4bf93066fb8abe485af6f17df1364c9904b04e7b5
z3d4056f916687852159ff410600248d585f8d33441b0ca25c7a5b7da89eec080317ff76cc9ccc8
zf99c0baa628d68afed0ea98b11489a348a9ef3207865515809712ca6fd3617782e9ed5b85deb58
z591b0c5f94e2c8264f7bd98f18f6dcdf2f1102b0057aab3ce1c1cb28da0019c84ea3ab198bb5ba
z0c82e0dc7457fa989551ac3589c56f9827dfa9282ccd108c55ff5b442c2ec1fba39ffdd8262e28
zb36e679d3253358c78cfc87281d0e2b5ba4c17c7f023db8ba3b10cc6e762debb7a76218291241f
zb249982df8e9eb9ac2cd501875548ffeec4fe133f87a173bfa59e4f60a334f09961f8adc9c2308
zacd086623bf6be7b00c6de90bf944315390374286676cafe955cd2807ab92d58475e142a2c6ab9
zb71fd994add95b04ab258a5d00689e18ec675c51b718e1783734ba26a92166557ea4eb6adf3453
z4e7cb276518308a1e9525ae41841f219ac8db03129f864a2b125a1e554265e60cd9a53ba6856fd
z74420481e164f34d115ab2c075c524ad325a0e95dc9472af289073bd3fd9686d2297c16aacd631
z19f0d1b2ebd2c77bd4729855a83862d02e6344d165e8e64578aceb85e64f348b13a9b4af15c603
z8ef0e4f5b04e3b34b86720bf317738a28c2c7be6a676c8c161aed2f77a523adbf209efa836d993
z8c4f84c1854da125eaf396798fc253c57b2cc40413579d957a5d790957a0577d88913f32fed7fd
zbc60336b41bcd98fc39996c132c93364500267daf7f6cf8062d0dd0e6c79cbb45b294a58cb077c
z2f71e3657bccddd77e6b43554cba98aea77a20e33fe2b1d8793fba08dd9b0174a4bf1075a3b71e
z22553864af90af32b355710002dc4ddbe3a3e39050652c77f86a9f1f8e021609a798caf9dc6ae6
za7a729de6cff7f511e5a3a76b06ad2e146c1f45bf8372d2c2dbf3ef502ffc16a0db23cabecc8b4
zc3ebcf5339306a39b1a806994ee52c7f56cb47657f577d763f82f08691ee1b098de6130f14d681
zc5370d5e49823b519664840f1f82a54590c84a599f2e85a9d37779e1bb6fd9c2bac34e91c593a9
zaea2f07e45a709d7ffab9884b16b95015e0492c047014eadf6a9fdad753502d2d13fbd6a163e42
zc329b386df55882c29c412fd58fc83da53a944538ce06ab95cd6c994716cf904e454afb336181a
zf3b1e297612e58a67cdf571605faa28a856ac246430ac423cb23e4d4a0849fd003d60b16b5fc2f
zdd8d38bac8ba2cd15e5259594b5026227336f2a3651e728bfe51a9476464460affd46619d4ab5e
z191cfd909540c9d37d3502e66f12c9ee7a466f884930c73b402a88cb8094f86dc03a82411c99a6
z5e0a9c90e902501560a23d5e921c5e2296b8b6bc4ba4e445ab3755f9de3d10a565494cf80bf2a7
zce3c97f6e7ea58b525b2fc1fbe9c0a219c3d4c1117f7298c010355317569f1f5ed045528a4c52a
z32f832a41104b477340451176736f1b5fe3b5be55cb2972ab02a9751fd58ea73640cc09ce120db
z9ea0496cb3b8690e16a8bfac1ef38d4e7e519347f44b5f226a185f373842d7a8bbc9bd00dd2c2f
zb0e645758adb50b8b5995a964eb2caf78cb5a7744489459f61c0c0aef1950aa821d9fe97cf1b94
z36bd0f5705911947e2d6aa028ca595dee8a3abfe4501e4730c6d6d9a36919bde2eb82f25f49ba0
z2a0bcd0189e8f27c03b5ba2cd2761e7bad4f4b7478a8fc16a883ea98e7b51382278d16cd22ac36
z536b6bcf313bdc6efe9935a71d92192455ccb3bf69b28095f1507370b8ce758897b39265316b8b
z39ab4ea3b5938fd23b51ba49d7ee308fd327f85f0cfddcb28288347746aac2d342cc3febd4e1df
z27a74595277df23d200dc60fc113cb5185c39e6bee18aab9c69eaa033fd53ee3d9465442923aae
zc5819c685de3c9503e56784060efeeadc06b4a06caa06c6bf8b621c66c17cbbcbb162cf0bec53b
z21b63b1fc4d4577647e364e8b922c992e796df917159a29984e81a4121045874ed4d10c9380e8a
zdeac1ddb0ac998c7a4a2e03c49dec1bfec54be3322e6eac1e339898a3516166163c3b72dd60558
za6701ca53b2b4a8317a8d7429e304c6d375cd58e9fc554564d98741e3e72fb0e0a00fa80d663a9
z7bb36d6c145aa3aee1abccb9165a557642d293c743e005c1974e72f7048de598cbbf8baa6d8e5a
z171177e988c5d8a3df9176d3906d81d58543597b7a86f040916cba4c97d7d524bf0c841107c931
z135d4686f9358cded0ce9b05335a9ca1c292e8b387d9733ef051861dddadd886e443bdc9f56be7
z1a5e071eac0be92e8e9a6c4fd9659d28e19430b76595ac404685402323217be228305098d6c450
zebb7bd401645403b9728a6b24c3fd27d8e674b6ff87f8d98c13f53a2e88ee63e7645feb9d88878
z6dbb23d3a40908dbba4563428cd1da78995b3b95b45b9f56258bb7e743caa404799227c7b6f9c1
ze14fc033e40141a5223adadf6b130d3d387ca1d498aa981ffad0d53434058a6a66e2d088495472
z4b3c336e9698cc5deb3b052fc55afb35ac0da15c6a77949639e148332c6600ff8748570e07ed99
zb6ea99793d15f3c011f462889addbbba06f22916d008b7813134eba1e51179097d880eb4363d9e
z6a375ff6adaee3e92a561c6a64922afcd11ed333c20185cd61748bf0f4b5b8060973fad6af60a1
z99e86167328c007e95f26e223ab8f6f84d18fa9a30456bfb225cb5f02e77226e660ed704ba3891
ze25280bd1c13ef3b86a68ac6ce8632a905ac6738193d82ad3884591c11d4fa4e2e8be9e5e5ac8e
z8cf11dff9cc8c7dc709d55d22df960ebfc9a8cc167847733ae2045193e4a081bf97564e1cdbda5
zf24e0b51079fe2b0f3f200a8413b75246fb1bfd68dc88c17e0314a661d83db003465004747db4c
z6989e7165cb3729d1ca27e07ad8cdcd908b900f37cc9316b6c9c93388e478fc7ed1c98a30dbc04
z34239f8fd13ac4649cb4f73cf638eeb4d89c7d558df9f43e09716088ef533a6556b4fdb9a6479a
zc48aa82f8cd9e20c9dcdfc6b5a2c009aee1b213dc2d8ab750881b595a859b4f511d3fa557240f4
zad1566a0865a699259b9161d5204d39d1caeed093ad8caffcd7533f20390ab9444e4636d4b9636
zcc862ead2f6ab5d63e037d44a2317a51e96073189187ccd028427775f91e37395837566795284d
zbe41bd3d72459e11a79f8b0c2234bdcd40ad950eaa2cc834721f8a27c1c653a8145c589ac2fd2e
zf99b562dd6b9c056f62232bc02a30ef64ed83d9efdefb381c64813242bc701ace2b92c0f3f2d00
z719d4fafb7d58783e2c98da4525a84cb3d903a1ebab00ec8debd17c6d6329a3a65853c570f1552
z65364cbc7dc8d9164a3f0ec37dc5544698d13f9f209993e303841c30e4e419e37520380232c52b
z6cda07644b37a487d063db7d3a529fb5fcfc483673cd22140ee095f89d1c39248a09c9e591062d
zb169c581f7b72b28fb92febad13bcbeee2bbba84a90e98fa64e093c4800b1b8ba1993985df9f85
z305145ff50e60feab559d524da18fca011f0d501b4ec3906341a7c1b7f34776ddfa890758c0bfa
zf95ba6394d2aa8f6a9ceeca9f5000fa6e5be31fb6c4de9f6c2b49c3f81ece01bcc6cf99b7fda16
zd943bac761ad5e39b61f8070501dd553b07f48e88d1ea499c279c9c4c5c04919b2cf08f66e62f0
z15cd8ea69dfa6f46103f7993aae980533ae6e372556e02d646a155094fce9d30fe64737e99c8a4
z656fb497b82bd10e5d2fde9311bd8678b86baad7e8ce00f883193a141212e16fae8ffc3c47a3b0
zf01b9e841bd5df46f25a27ddb32ab463e2c8a4b2480a15dfe9ddb21853e0f0b0198ca47acf21a3
ze6aee01a7bc3e2d1773041c69c4d6fc4b3d59125e8bb74db913919b70e2732b77ff816dc3b3d41
zfdc1719739e1b8841b8e6161634b9f42349c9a3597185b432fc91075366709ec2fe2f26680c2f5
ze5fd466e542947d17c58c16f98b564df47fedd05daf194111a5e359c5e6578abb4ce9bb392b7bc
z64d80415721af14b2df203a64f6b55baab1198db3bb0ca731c9a28ee9bcc9f68d7f7aa1d6d0657
z267a41b418c6c61e0906d576ebf3e8d17eb098cb004eb969029da6edcf5085771f56e9b5babc39
z84f83e0fd94d2d24f5403423f6d583ddaea92b6bfa66d33496883fde6b729c008001b0d043ebec
z53a270c648b3f68998e57d0795052763949b6f1de88cc7bc6d9ce1721f44791c01fd6a363be1da
z1725c183116a6895d8cc5a2ba4cb0363414c9b528f06c739910fbe4eed55a27d980f9e453cd629
z39c4f2ebed193f2b7be61e984b791a154ba8dcc96a3fb7d80cdb398cdd0801943ae5dfb93a96b4
z2f372104b8383e6150e5b215743e37100fd1f30f59df213ab57c21af61ed369e4cb601f551cb87
zbb271306fb9d22e3a66e12dd931238f8787585d48f7e0fe59300ea317477ce450eeb5bb93928fc
zf80e327b73b6beb13c69c521ef44e9232a39df1fa8ec73ea2feadeb321c61ce25f5e4797cb75dd
zefb37d80d22d4e7de0a98b8108ebc8b36203bc50443acb3f5780dc87ea95bf98d7cf86b7bddd0c
z3e0c8c422b0292129195ead2ed24dc88446f58f81bbbeceea811f4fb886bb08147aff5f76b8a82
z8752de1eb03803b17ca307d477ccb1319dc23e8d2a74d8a968da98e4bb04f451775cbb98f7df1e
z989c933f23ba2be8f2dcb9c79e1f39186a52bd8523fb1391d6ec7948ac5e0ee4ebbc46919bb81c
z289af820cd0453c7a402293994cc9999a2edd8a350a80461ef248f3150031d936276ef6a2abb05
zb7de15d60fbce4286a68c46f8fc3fa6cefe4a7be36e00e63145f785fb649b6c3b03ee73834e7dc
z1014696cfc607b3c9934f0514c536b1062928123b86e2cd40e9fe2091733e5da347b7635ea8faa
ze76814e1a373435c25b602f13b0cbe1487f6ab34da1fa7da8533492c9aeb4dd862fc63bab47009
z5ce4c9b8e10fd60d7c4663c8d004d2f672e406b0f142e2b19e6fd0b1c7bb0f0ddc08239675ea6f
zb244095eec7b41703529f1dd2c297989a6c339af4bda3aba41d4fcf83a5957ebd2f616a2ed717d
z653a39f89a5282b6fd60469502cca4d9bae11b33972d659b5080deff64663d87eb58497c8ee408
z8aa9924b113e04d46e9e816050f3e2dc08143db52649403b468f7c509232501712bb658ed49f02
z5df23fbb312370ee9afb06bbe6f6ece0ae8ad92d627f6d2e002f860dbec02a34b3d2fa27951879
zda0cc17df65b0a9b35f6add37c92633aebd1b82ab4b7430e0dfcd476792c051de1b2a8d0a9f763
z4c7a55cb6d6f3bf5d23081d1f896f6a6b45cce2841b9ec5f305a0dda4786dcbef2931867d1cabc
zedf976e8c59f29f2b291b7312f603c384568eef41af04cbb3d896f2cd6ac8006579d6110f57145
zdfa48044f6a63e763003eb7fdb2738fcf71fa055f919cc6a8a1f59c4a24c763c1a75463233221f
z2d41350459fec847aecec06edea669411f2a62a2e7156aa5bde0b768d9d80e9b55748271079ccc
ze2c30a85f4f92c11885e241c3a8e4a4caf664443e01501cbefa15d400108eccc874bf46b9652f5
z319152733be306385767b9e770e6c82063e2496763cc91a02ca43dafe8d27738ff64ae175691ee
z3bd71d14299e2899f78bb94e8de32b42b60c61a454b8bc476f60b0186f69d7ba47087734d5ea7e
za6f23a1179ba8cc5603e8ce71c0a072211eac8435491b0e7662a2d2322e8e7a83ce55a24a959d1
z7d35c44c62fc1e9c4ed20f3e8e2cd55c2cb221835043e930f1c7f7b9ce41fa9a3cc83329e6cdc7
z6163085c5cb9f1b1a8d77bd51a0a2ebbc4e25284d75c57d68a0b30d7c8706cf08feee2995978a7
zf73f5ffad77d8d4cffcdbf24f834803ccb427b1ab19f14e7f9b04681ee868619b8c00b432ef657
ze566d2bbc9c00ef466eecc57b00f5958d8ddd26fabb477006e960b911574c577d3e860d3a41215
z1b205f93fa57ae5476601bf92af244f4ae6bb02a027fdc8ccd6efe98aeabaeef4678a962823b33
z78f0e2e7d28088117b8d3f85b591eec429c507d9751cfbcef038e5e7abe9a3ad10b2f90c79f7c4
zebece5a49311ab566a2995dd84cfaafdd903a7939cfab63c19a55f6c153afaac993036c5c4ca0f
z901625ab35c130352c326de3da0925ae1e27c06c0adb4f1e60f3f6872ce4c70567682a905666b9
z4688e8e013e64df040dfff8888aed44a776426b53f702ea6e6b5869925693cd508b87a192b81e2
z2d02eb95eed07992017734d4002c5e38b7ca2f0cc34ce064ae07beb4d964ab9193d916db5fc2fb
z787558214736e63c1e29a615d25d7fa9020ddc7cb65d2b00ff642164773a262d2e138d78cf6a4e
z989a46583082d9a9b444e74b73f564caaaaee5dedc63aecb4247450549599242ab37ecfb08ae46
z239d214264f01bff34325aa6c28fcc59ba70f0207632dd81daa97c07e0ca322db1362c21680987
z2426649a0528fdaf96dddf3c1d4bc6f093512f118d45bf278ede9f56d8b529c644f43342dc5c4e
z2f41978cb35ef780b60f76d054b8d303c5b34536c72ba4e8ad1d05a226ed34dcbd0097876f7293
ze8ce49295613931de6ec5ed7169199ecaabfc1ace731215eff007aeb616db5c40f534bba6fad11
z93be5ebc966386fbbe8c83d9286344392fd3c871c609b17b3a49355930b06dd37257b7e0145c27
z908fbbef8786c0eb5bd0eddf5ca6b405cba6163d1a876ea4fd53ac42b227a66a3f0bc0075ae15c
z681e0d128379013f00d9796beee03300619e98f0c47cbbf250c4981b142a914f8a303f3b622f52
z13172052f05dcec2c28ac09a9624191bb684871d640272bb8d80936575fa62761eeca130ecb4f0
z67fa4b39840d6a982ae3d31a094cfbdda8e7d187c1d7c15208f917607f6c827b987e036c1733fd
zc7b3d5180b9f6e9f493c8328ac0035a91c703d02feb53c202af7bd0eb577f7a5fad37cc3fdd84a
z02ec301ea3a53a584f49bdccab0e7aaeb73cf87893d618396b1a60dd14b8f2ac10ad06c813fa9d
zbc5c052c2c3292c593a2cd76ea406f3c53e339cb22f7766aaa820bd45c6da56f6565bf36c4079e
zde9fbe6885803194d452c3b5b0cf9466a99462ee36d77586685e2b8cd85c906ef04e47255cd667
z7289cedf15866c0fceb85515db7978b7212f11601a1805a53f8640afaced6bcd2761e316c87043
zf10e8f693e0e99b582056f28d31689f2b0c728220d4b58884eaaee1df8dd7b6b09a5046b82c77a
zd30743ed516ee1a3ddf8a9aac22e09397e1096fe6263992e90d6a2b8b5bbe8795224cacd7e921e
zdb2db20c7919bcb5d8990d33c15229d39a9650465d9f66a509f7e379e3f381643c12cf7ecb2d21
z682900de5404bf364ea05f09f2ec7438fa79f05224799e3bdd7bf0d34b3af3afac2f923087aa44
z2dc9081b04cfd0c4bd9ba8c84e9457f6d5b8d89c3c82bfc649ede02b53cca8fab99552ce306f64
zce50bc4782caa67e40338665dd2ece3d1d6d6b966faa8ec7164bf319706c91e0b6f54941af7cf2
zf4f6bbd0547824c1d8faa328a29875ca4335e604ded69f9d6932236a207af3dc41cc0965e1bc92
zbcd05e2d642bcbe7f8c1d6aa54b20d56ef5d49851ae961645af3f1dc07f1818349149efd96d590
z9af7ff5f5e1709999337fd555de41d059aca09921527b33445c6775b53bae8fe1027aebe42b1fa
z42906b0571806c0fca33ccf88edec31b7faab81bd5cadf5e6070afa5098c7cf50fa4cb415437f7
zcf3c9a0bcf72966e47198fd8f3b635841d6996786042de553535190138d2dbeba9753852d0e58d
z7ee5384801e72a0e22934f967cf74854838c94dcb7307c9b7e8432909fe17fde77ca2b4bf759c7
z31f36f6fe3b5c4a704d06f3f3ed11f8eec6ff52eba7b9868e2e9891333d84186a18ba99805f7cd
zb0b49a4391e071ee0a5e89c79a79253e88d3879ae3b557429e69b96d48e8b9bdc37923f1dbad0b
z2cb655419a04af92a63ebe1cd58243c8bba888b86e5b3574afda2a44fecd8e09d9431d816e9141
z66584238f6cc31bc80393a28ff0e90e34f27d068c14bf017176e197003e1cbb0621ffc20c4a8d2
z1e8ab55e65bc9d250e8b229704d748f1fb9cb6f4b902ba21368dc30f92112a2f4eadf4740da8ce
z97d06dc1a0ed30e4ef88dc2f1f5c543769b15c018c0b6ce9be353538860453411330ed9f1d930a
z087f2bb5c573d3b6ba1a8121105d20e949cdf6225c478d691a532be914e481c3c602a051a07814
z1960dcd5a4d5edcde72ca547b78cda7a574504f29710b705d932fd22763d0ee3d19102bedbc29d
zc58e0d3a82120a51d018d3c68277c488e9bdca6777954b54715f8067ed9799f97a7dcdd5900eee
z4bf7b4faafec10ad93cf4822be7ff183297c894fc7fa8efceefdaf793e4949c39645c05fd30b38
zc93409e4026e3548f25aea12c17a6952b004dd9bfafa016a82943f13ed202854d50f6b3ae3d656
z237370f9588b3edd06b013ee7fb96ad80dab5a790556f01be66f1acac920a26fdad3e49a993f9b
z2c5d4a4189a6c3232772094682f4a712195247d084cee279d3bd80511ca9c967babb236ecff5b3
z2b7b38a3394e786d56c967099ceee825df828758cc72d2e9347554c9b5e4fb630129c06ae5e31b
z42639445cfa0d72461e9df85510ac35995787f3e2ae2712b2cebeb6f5e215724e8b3103189cf06
z5983f5091ec19dea95bcb713b3440dffcd4edaf1e59f4ae4ecb44b8595130801599d16808d753c
zcea9ea9099e16f06dc62f4747b0b1edb52c23c0b89a0a574489c2115f18ed4462e7f7d22939088
z8a96398f3ef2eab7b5fd1c490018712b39bf585db2829c4e160a16e701ad834674d38f7ce2139e
zeaa914d3b9e14fd658445cb5640f51afa227a249d9cf53a15826bfdc94cf2bc1b29e3a2ebba937
zb17f2b9c57d5ba04441e43d4f6bfe2e3498e91394f20dae3a95c0bad9dce41eb3b764b3e1b1b73
z7f88a0ebfbb23306fa66a4703bdfcd312010d4bc3ec6a37b1e02196783988a3c0f7954fe1370e7
z255ea1e98a6109d962b6d19c151ae8d70b04f9398fbadfc595f8ac37de769942cef5fe4249659f
z44e5280d4d03480c27d00f1c7fded58b574c1bc5fa97e4982077da058e3883232433f32f1888b5
zb8b314eae33ae2c0d73ebc8614f2646ba39fb1e0139ef17f0ed6c210ed881de64d9a81c97fa3d0
z82517b54fa87a93628725c7d2f5f752ffce51f7a0e9281520d19f50f9441d1aa6e6d04fd832270
z98eef6a7bb36edeb90097a96ab245445177bfb14ce9c223936269612100ca30c6041014a982568
zd85795eb707526280b3d5c30e3c16b532c39cdb0e2861cd9089f4f2c7e5dfc192899da92902cfd
ze6b1028cb9b4b930d959217d02614e1579cfbaf8d04046aad1bc4fec75f76901c8d3f83ce55df8
z8736d0ec21744d4b1c2e640c358c337bccf34a2fa717f939e0a54b714ebd63aa754e69e8235f88
z8411be5c7ef6b721ee7c2e5f48891388b81787053faa2db1620eda56ee070cb82b20d2ee63844e
z06bb036efe59b86ce0a8d72a0e63bacbbb6e77267e4f72d3068927ad7e1acb97be2e57782d3d97
z597b54a79c5ca3812c983ee38afccabdc959ac8935ff1f99903c4e51cb0d3c719b51615eb36759
zb277561bb3f00490b982fc473ecfa56f4c8230c0895e373356341070eb5cf127ea793bf7f3f2b3
z14c7660021002d6cd0f0a71ee53a7ceef0bb6ef66bed8b4adef31613f2371b8f50520f90008baa
zca09f36fd17a666b311dbbd4649ce255852f0844646263bff57a382e63c7ab21fc5491ad996551
z750f993a0bf342255013efec9d83e6836fb33d775974fe570d6ca48c30d616518e63c1c505d5bf
z0776fd4410ae5eda6aae352987b00757c4475da272b471277938998b33ec33058c8ddcb49c95d2
za82f86a6230c0c5694fac82b969bce7cbd7fa69a4a8ea50772e4c7e59b98a6bba312de9669b942
z9ef5726d191eed7881be9eecd7358742cafec163d70920b82d9644fe11d03e3e981ba0c505ffdd
z6d13368a86990860b2f199b588ce81adb363882d9784112f4f3dedc6499d44918e308ea889b96f
ze4c592b9e699a02bd244616b58a1d0327c00d854709beb4e28e7f570a8473eb0a752b3c2b94a50
zf1a59147a902ea07e06ca517a1ef981f15a67c4884e764e3ca80131a7cb6817dd4f923b825b0f5
zbe2b615b37361e6039b427046e12fb441cb91bfb3973ac273cbbea974463d13a4930939d833f03
zaa386b9756a585a8adf228c78f9fa3f4cd51ebc1da077a728a15c63f78a923d3f2ffedcd04513c
z4daaaab9706f541a835c7468de4c070449a08c05cb79e9c9641c4cabe0e4cce80022e754eddb8f
z8367353664b9f43379c59a569511d73c47ba146540be84fffc88b35d0ff26b0a0cddebad57a574
z4d7abee09756f8cf4c3bbe5bae19551e9ced95c39d452bb8f350d68fc3ad0beb6cabdd35517cc1
z3cf2ef7c853207dd40c788a9b88d99a9a72209e0923de4e1ef5aa869213d54a1dda2f37c1f0007
ze35e2fd174066f4706798914a347cdfd8f72ef909052122ff472995a40adc000ea8e4c9b84c9a7
zadd1c45f2330dfc952d67420ed2bb153075b34ac7d7e0cba270c07b1170ea583b512a644eed62b
z1b1555051611d5b09634b7bdb465213178244f1ca6852c50f95213471ece9d29c18dbb22c88b7d
zed8c3d32d709702a34d0091107caf37d126bcf41e9d00d05ddee528d67c8014fe46112303a9d93
zde7870e78f846fd3901dc1c0ea59115ee043be98735d9ceaaccf4e54b418d4697cc835cc740a0c
zdeaef48999b127c6820296eea120b73ec2f3801cb4a27f8b0323de27c9e4bbcf9b2aace5e6e73d
z218e08685cd518dc9e9b4898336fa0edd7fc71e024a503679043a35cd3765990803ea4282360e2
z9a36221ff8d6cf730849bd3e3c1597e2c937949d4ffa0321098ce9413cf42adbe372017420b2ba
zca9e47466d01cabd869b270bce417c3c8796b3020427abb3a49fb77c0c3597b62a383529696f54
z554a627037ea2bc11509034268647ced9ff778b4e9f698b51c347a3a867c97e735223f1a5dbe92
z9e80774f04eac692cb4abda6cfc37c6f232d9b5b8e6f0c47a1a3bfd5942a3e6479efa86f9331e0
zea9d625ac25efbd624a887bd38e2a91e43a44931fb0c9c81df00798e9eb74e701a8d4a86da686e
za0a124a621f0bf220627cfddd41c671c1302c7698a60366d401fdafcdfb961ca8766677c0914e8
zcd9173ce6a8e9335de4121d2655ad5c14041cf83901938af01a3670977eca2c6edc242cf9a2272
z30262537da8273e44a43ff7557ff43a223159dabc2e79160e40d43e86f3116aa2fa2db82428212
z73e5538177993f5ca2839c67a155d832adb1161469043ea737f809669ef71038369d3c186bbf4a
z7cf38994854128c0f0b08f73bcac40165a30ae6febdb8f0e3c5363330b81de11e4c87780632040
z608a86d424945252a35838633e87dbf277ad5118d90b687342c6065a0b6e0dbafd90b15343f5d6
z3e1e5b9a85e9fb68b008d8a6bc0c8b5d11b052b1b79e40fd49957befce33dda1384f69edb9f724
z4b47fb32f93a624a9fc5ca1154f323daaa1642397e5c2a737514ac40945348f6467e190a20fecc
zc576b94a5b36f4272c2056c11b4b0b770fa0b0f2642e6a97da609d508f82ea76f1a2962abf0fe9
z61ecc643b389f28c5f13cfe8db6aa63357dc80c9a8979499f688e8f498916453d218569c4d8c47
zacb624e25701195f42ce22abc82f1a131e84f61c44cee98749294c86fb7bdf4c87ff22dd7cb177
z18394692e50b97c5c736b32fded9c9daadbf854f2f7dc67199a131411be1108b377f600215e7c2
zb9afa98a37b5b3546e6e95bb66f9b7816ef0fb6f95b692844f8695dc86596eba72209eabe40c5d
z2f0ce00e427e8d46b6e446dd529d0fe0a3328a5d5365ddca3d0f5d6ca16724ae2ba2fcf5ca52ea
z22b0445e6130e575a4d7603064a46f77183a0d4679c2e6f627b278e9d50b774880eb57bb3cc0da
zb0853637ff981f6281b177ac6cce074aa430233ca39411842017bd869694c911e2aef803cfca5f
z8903e96e641e788bbcf8b3e27540ba46d81aa3567c2db1d7fbfa057dded9e0e240e8490c4acfe9
z0712c35bbb2012e2739fc875da0978201c00269abd2777b3f56b2f628a727e43d2bc4d4da549f0
z3c1851198c377602f858ff5ccd15c21d4be3280f22470f52882455faf3626892527776a625877f
z069c18a502c234376ed6b7af5eb93a9b644ef6cc92c3fff269478e28ca70a8a521ecb94a242ff9
z2e8bffc7bc172e5de726afe7e5e4cfe5665feccb2df5e5d9d0182afad292b7e4382c969c55866b
z8f650f4f5aaf8c32d7204c86d66dbc6078bc19de5e4ce9007e99c8148b5cf2a79384d5e963d95c
z0a42a72f89f3c73b58cdbbcabde0ae32e5fcb29070e9f940200ddd183ca346187d05f48e1101ea
z1126eee893a91a10bb5cb217858b28d6b27a07dd1bd1c9d8200eafbb65a31c392fbb62523b2ef8
z405ecb69e249fa545963c2d49545dc8b10220b87d49d1bc9399ffea6142e2bfe70838783f08ed2
zedabd4c1a362e1676661bab138e8960cf3793185908b892dd8be9ddf332c56e4e69f3c098f32ba
zdab03156d467661552994fd00d1c52d2faf89560fbc0da794d453288ce1668990d7b22b093cc15
zc60c5838593273c6235aedd48ebbf0f3a52d03fc814ff361e418575fbdd87e7f4b2f96d0df98dd
zec033a8c01a80b6e24706463ac4a0f622b9fc6348cf791eca88ef2d21b85549ed14aa55c619ea3
zbb0e942f7a84a2a66cb946d5a309bbfc784afa8cf4db49a252bf9b71d9e6793ae3f7000c95d9e9
z9f01b6e599812fc911bd42e36dcf14df44e864833daaed762986998c514614379e1d6ae3a49292
z40dc1a3bb3ef30161a34ec9f7e1459e09bad5107bd6fa9a7d79f6a3f2b42e43133ad217be27269
z8b2475face54dcc3a515563082fb71b2fd04fcba8ef47170cae5f469e5345e7c481f63042f61b5
z07646657856db7f2dd8a5e9460828335ea240af444b3cf4f7568c2448bedc81b6b0cf8602eb330
zf66946ca674742744d3c34465138609127457ab1dc885479a50a231dc53026a8383b3ed218351f
z7967a11808b061c29941179922fbdf442e6efe62e17d024f03935eee21e7b60a5ed1666bb28878
zec11b75082d04b6e32cb8f6d41630212761c775623b42cf20bb681b46ced7cdb823caf3caab41e
zeb3b2c0e430a89fbb3883d3b1fcfee0940fbd8c27a02b2bbead13c5646cc0a79b73718604e1b81
z6d58211ab66a125c992bd298fd52feed39227d63d1298ff1205d19d414a9ad10e2184d02b5f18b
z99e64d4b8aa2cc9cf60c296ed8aba2be82e0c6ffd4be3e42ebac0836f379aa52bd95c59aec745d
z632cd8d0c6133d8541ea4b8337db6b1540b0e08815830beaf84ff0abfb07c3ef38b95c80f888a6
zb5e97ddfdba228a64064924f48dc972b66946f64474f71cd4f3ca71ec1919379fbb762db24fcb7
zefd1c62c8db686cdf779e34511d4f928e6b7c25ab7b4f6d308e1c7006e6fbd10c8bb2f7bc71ab5
z6ffa47972e5ac51ef099e48209e475b0da5ad1fd7d76809071e2663596eca4dadd5f35cbbf5ebd
z52cb433d73c63350c16169b02561012913c1f3a250982283072bb568f4bfd7a4cdc93119775b60
z12a8ba5fa8be524b86fdb2c7c2ebb3a2b1cb8f2a491ce140c5e87e23860f5ae8b807112325b059
zd16c022de27601958ccc656dc1124773649b069b0f2b55c40fab8d78167e632e9537e458145087
z52696d856350181edea30ce9940f421d4a4842c872c256cb103b7f3ddb8f207d381a3dde7f644f
zb7a8d825bb91e8802786739389bbe4e9e674c4b5c67581582028466cabc6a549a6a850bbb7b16d
zc8518be542d7e28677727172e1ee6cae34f6594bb05299b188701660a6b6dd62f961e5c21cd33f
z6a3a59c7783e02ba11807558b485e44152e61ad57e2eeea40e757c87c76c2b69b717c5c79a2d0d
zf640f9025b1d2cb22b437d436e3e2fa5feb5eee9128a83462962551ebc7657b6e13d7832cb4280
zd961c744700ef512cd3a8a8fc35e037bb45709771531731802d41cfd4898b012234cd44b083c05
zd79889c4613a7f5376d3ab570bb2dd977ef3471f95396d61dbc61cfd6d3df20c1d0c8a922b05a3
zec7691cbc9ede511a5af5c9bbc92a51232d122bbc06ec01b599e240f9ef6cf7fd0baabedd9e823
zf3941fef23c8441ed976211329b29ea6bb62c22bebf09a02e00bd37f2752275bc8ee6efb680d28
zc4474bca0fcd222281a8da1851b74fc9a0913cd4f5c1768dc17d84ba697bef9a427c6a48ea4767
ze057ff482d2178f84417bf1108090dfa37e007de2896b66b62484f23fc9b444e1073c93217e112
zc28fe4fd6e467fc48eaae932103ee6a3560e51066cdc14503d89b38adfb9abcf9cc732390eaadf
z57948516971f9affafaf39792f1856e85ea6fd02ffa2169b757f773e9fe8faada30fd559269ee8
z17f20cce38104cf500fe4339957b564fd42bc9601739ae8cd58c6661c4160cb0a33c7299dbbdc3
zd19ad8d841904f40cde542f535227a285ad329fc8e793d70738375968e6a58fff4766480712ec0
z164778e972b7011a8f199a3c699b920a581984d41cfd3c4365eb387c6fb5c3954476ac610c829b
z9a2393f44f1358212846b78c698527901e3a622dcc028a8bf59a468bedb65871f283a7f4e1e85d
zb09f364ad8b77be5fe3a6fc2f898a63adc06d7a6876deca97ae7c43a172d4c8eb1e3e7480defc2
zd72b9d568bf73bfd4f51ba823a08d3bdf73bde9cc19a39617f172f5b909e8151cd9b2718aeae64
z5a22dc20fc20797fbd9ece3a4583b94ea7c2d9eed33b00daca81c172afdec1b6dd55918c086958
z01ea1a545244661031ab5288f3a8603106998c7017d337a2e2bb56185692896f7fcc70e851b190
z1c93a94124a474415d503c72acafe1a820cd1ea3fb63d3d215b076bf6a3f97cebf25c6331006e4
z7a87a213f84ad0320593296d9c68eb8b47e10ebfe18e098e20408a414549ea8ca10025f5fe50eb
zc1786cc0d801798d88bdc3206cf07e4f83811ed1ca277f43dbd0131198d3722b6b2e9550510b0e
zab38f142db1ead811130a707b83a0187a570fd096cc24c970591938410e939be04350a23edd4bb
zb7f09962c34883276c10101f6dd072511d9bf0695e8af9484614225141abbbb605027ea2d6dfeb
za58764cf5731acac7f24757bf3f7ea728a9ae87f7aad038986ce2d68e80e7d783352cc8e85f769
zba7a2fc1019f0fbcab9d6ab1dc4ae2614cc66ad4b2a752ed0cb77ed4ef95b5b6a492fc0fde7859
z008198ef317f9285fc44ce880da2ade1225fddb71f0136223542606192e3b5b3d1b4a42aa7eda2
z5a882607a9cf9f5d2132368bc59de8adb36b73663ebbd4778ce36c27d882fc91741bf6e44a4ff0
z2438680113256af8abb5a916a122060b82015819ee1a965a9737c72ba23f89902d1160938f398c
zda38f9b5ee10b74981c960b770c6becdb8645d5be48108e8952edb45e9f5e3b07f208685504c33
z5dab3d4ca68ae8ea660c20b417edb513e3aa5be9494a45865b436930275934f3d3599a3844bf8d
zd288db2d71d287b8516bb90959790e7fa6a320d8413cf64c4e42562151a6d40ab163379b501ca2
z18ee3861c8fd4b56d340e02ec56b1f2182ca87c80fb488c91f54194c0b684ae00fe05cdec19887
ze8cb3a4d71b63e9301492f003536503ff47fdec9a0c27a3cb3121c0b32d2fa8574df08bc583587
z555e3ab55773d13c89d39b123dca9d17ff70949f16e6be508cdeda861134629b1393d42761757e
z21b38feba9aa6668e1388652484401ecf699b103161368c2f943c1faa9642990879e3126d0871e
z9f07f1c2458ff52fbe7b4ef8cf44fc115a5e09472fa687e1fc9d935a87173d8335650d5e48fda3
z9e9999081cac86705d2267bbe3c0ad12c3cbb5cc24c086ee2fd1649f4eaba1dc031e74a68675dc
z4593507b972321930cd828a29eb9a681ba25b39f1d58403a402b3dafbe6fb077587e37b71ab841
zbe7037c241aa3a37bcb2c38f101f705cc121defb12ca7a426d174fe6cc0641e0aa32fe596ea48c
zbfa245abd0a385c0d9798d30dc206a21bbcc780e667042d400c0b6347ac09bc2dcdc92dc545fad
z80dc195c5083db835a3e50dcd0e1a7945d746daa6b256914ce1eec525dce08a61e98fedd2ff939
z70442aa9ae6ac9d8d9d34bc4171a8c5cd0febc7218b1d8905b5bcd226d5ea1fe39c92580aab39f
z1dfa966b6f0e6b0a7cf50ac0c407d62b10894378e8e61450536138199cd38f215d56abd43c8afa
z11aeb2fcfa75a5b69bcffe109274f6cecc31e030530a9085cab0366153bdfedc13f26d85c9e21b
z36829508939b5935ece4650888b8db600223da79051f1fd1f694441ae2cc92bd3c406946ffb901
zc7c47b6eb32f906f82cf32f6a6426fefa857e7b9c8bedef558dcf3425f33b9317742e2e69781a8
z7a5d6b479512f460457f590276c89dc0303c0b4e43de665ca72f6452ec8dac386606de82155487
zbca73ea33d66f3326750da24ec85109bd9448bfce89f8a0b6cb570845acdf532fb01649ecd72d4
z48152a9bb0a71ed2a23e68f88d36050dcdba3af08fbe86e3620659ca18170fb98ec05bf83e6b99
z25e2d1d6c4a5ac93e412e7e2a69e8f47048fb8250eb7ff083a486922979154ff796256a9e5d038
zf3e4443906a097f36173443ea55432769116dd29d9925c584d2a7c7b07ab671591e60dbd16035c
ze3c76c70e01cb0a995663abff19fa97735482fa42ef8fec8594cc390c765868b42de203f8ef70f
za2787f377d4ae237062cdad9d6ddede92359148878fc4d3a1fde93049ef7486b8be14e98bc9d93
z90e50bdfa2e00d18aa2cc50fa8273e70952435e3dbd3fcf2b0917bd382eb42ad6204dc828a91be
z70d5f44bce61e75ad863957c7256f31211d06f84b89e76c59f7c1f8141c205d731d690c73a4eee
z0ee4b0d821eaca742fcd2d94af0cbcd23334c98a4b180da47e75fa724af6b6937b8ff158adf017
z366767674e1bcfe82082a22ea68cba5b3c0e67bdacfda4fb3f15fff22b2f33e717357d16602c13
zd49b6bc12d8d733d09589ecea23f6d4e6f713cbb66589dcc09440dfe8a77d8e9776fcc70362b10
z20f96d01f30b2293730ad776fc9d92f9d08975ff1f53a99cc85fda24e982a997f33ade5bc48a23
za03ea0d1d2e8cec1d7005c38655066841dc262e2873f90c381534879713335b0aec99fc585b418
za3d47acf3625c897069a8e4779c2df79b31e38b3aabb1da1d6dd41a63a9ecc8addf05ebe9de927
z850cc02a4c1d26f0d43fbc4fcdd6019869788e06b01a6afb7b9b0386daadf35398e2874870b1b6
z24c604e6e1f8fcd0635f8208f4e71346a2d76ce345a7012f0111aca49de6fd88e086b0c9d40bc0
zb4168df1ad71032026ec789731f7fafc3c3347324ad598ca69457cf5b7208c8f5a2a4ed2894caf
za02894055b401b7abb492b55fddb856ac5ed07334171f59aad7d1c27d2f05972e3b56e7cc926c2
z1a0c3d673f54005936f8463d460aca2aa05612d61de6cffadacc4263bce3eb3eb8a079638f29e8
zb26fa5608b69794930aee8b1b20e2150223161d234d48332ecade1e13b07b7bf9c077af7ba7b47
z164ac6d96d82a851b2bb5226c2366d4edf6f3349949f006c91da35e8d8476445d7a48501e4ccac
zbe9eb63a0d858af2ff90cd1bfd23832173057e5123c2d8834d0a9024228b0f8102a0a47fa13445
z3878f318cb655e4a74835ebe3a80354449b7faadc32725831d492dfe42558a9fb4e69c24756c06
z3a97a89601a9555d25d365ffa31cec494691ab63507624ff035c764fa1bb9bac3876a2b969510a
zb6709a332941963dee8b4eae345c96ed0480c0fb1567d52b44dafebacaba5be3b6f63a405fe0da
zd50c9ad704abf1cd330dc789de2ccaa2cb10c7f9ddfb2ac434ddc5051603b0129b49673513b1a1
zbe525457d39ca8386ef4a78b45338f94c7ac937a4a819f966bcc6198a30cca06847eb9402cc1d8
z3e8447927ee5ba60037621631ce0359d09064c4ee58e30ac2580d710b0d6323c53c2cfe9b6a9c5
z95d67e1df9fb608f9ad36a29d1c40d82ff5903155b0fbef5152c992b018271916fe9e6f085c1b4
z137c5afebddb778f05101affc3029ebe8d3c92091fea7aaf2ca2e74e2c67a1d3c9a4e40f81103b
zba70036165d8901101735b4e82d8b2b2b4b3745c9b2817a2256201aa41128ea43c78516b2225da
ze609161215978c91cb8f70d63df8a5691412647b5fc34b557e915daf40d62161010450d21c82c1
z32689becc66f8ab8a1794756e0ea0c5a0f6651598091cb99a6e32deed22c8d8214891e32b9215f
z62ead2f7e4b278a1c79d42298767ab05ba0410aee12ac300edfc37cd668e4dc5d044187f3a7f92
z96acad6932c523d92eada4681b3a354a9f67513378705878bfce9219aa28b7d649f2eb0c5283ef
z37ec82be245c5b9f871c24deea866a7dede40da3b51f36b0335e7da3ed20a6d084c10879c2a560
zd0af5b65254cbc4bb071574ab1bccee111f62d0a7071963f36336882a205f2b9fe642f52e3414a
zd9e7346a41da60d73b73482f4b619d6402a58efc00e225b324ff51fd2d97d894d730f61dc4a4c6
z0bb9fb8716327f43cf7e35ba53a8b3bba09cfcc8ab0d5aafe826e4b995b1f71039d54331a31ee8
zaa560c4a17e5e7205e981226255e4e7e74e838aa2415aeb409045b2a0d5a29f64e88c75f75798e
zddee9a503149755e35975b8d260b3fbd2a581e4316dcc8db7bec8be5a066ff089066be1846a664
z302ab510a845e7c1d6a260c32f18b1ccc634ca69fe16953f488018d20f60dd6f9d78969decadea
z99aa2a5b2b85c07f7bebf03b744906f2540c1e6779c0609fffb7c3069f8949101b6e421f803a76
zb989d4709304e1956acce0ab3509f99231375fd936b0ede0ac7c9290cffbb87d4bc996a9999e7a
zf58489e8898ff3a18e3a35b869024d0d5b864f1273e07b87b4d64b7205a1727e8bd353c3aff6df
z6a4026fb6a3575d7ccf1c2e3a8050d3d14156cee1f341bd55b4c18d8d53b2c75babf57ca747753
zced534ab975b2719eaf628dfd7a947d751a8e3c417153cc3476c3aec6c5c8df3e1baf61a545a89
z2eaca83f0f589f230fbf5898b6d713d2d61ca185be3ef6a2f85e9fd491a7f13d43e1446def74f3
z24771625f4f039d2751f03445750069fa01707fc445cc81904701f08754d224679c607d7aab350
z89acce8cc7ed33d2071ebd0c13a46d95ad98f443b27f25f878a230a63ba952aa23710487e42acf
zcc50b4c55538843a71120c000f80f2545b32064840bfb050f95c782ffe429757cce650958b2eb5
zaa16b5629a8a8e2c5ac06df47c17ab3f4995223bc8cc0ecd06614e433597a9d4d1fe69ed9cb302
zf20039cbe143a57feeb5fe3c76749266c5660cf87e926c62c600a46ccd66b66028f44a7e438a50
z09f98e8b38c5f66aeff5824620fb39a184952d8f1504043c753a95f859ce0e1e8c758c5f1a23ef
ze1ae1548bf30e465c5d4fb53897f5ee177662a5e41edc5e1fd1fa9bd34b85e2717ba65825a2a2f
ze3388a2c1024557505255c5517200c99ba18faa48067669b7f08c7b359625b2a05130c493f8c6d
z8b202ce6be080e8e9ff821c4869bbb339093b90764ff79e3a46258e0417c75104089f4934cc497
z44cb7e5a83988b27d0a2b04f136279bfbbfec13bf84f71a36a3e0659c182c5bfe9207b0c9090db
za3f51dd232ec43f65464f5ebf1652383e1866b277cb96875107cd85da698f426857429df2cc9e2
z7550f86b06f9dafe9ff6d4f943035db00101b047ae3d62eb0195949309634d0f5bec299aaeb24d
z9a55d0986662ba38fcfef882262caeb74af129a9ffbcd1df916f46a7d74aeab597d9e28c57ae9a
z5d506cdad96c8951f0167d0aab4296d2b2951494b79d169aed1aa1f2b740debb30531e84c4f688
z28997dc87b0848b8d4cce33c7b31ee19a36058c683cabed7368c18eb690286f9cd10223f224036
z83d5b3eaddfee4ae633bde387c628ff8c8fbd1d7af49f19b862cd7ecb64b1bb29b6e4af2e08927
z9555d7de3f641181a5b3e6f46b2dedc41f8fbd7638006894b6c405c6bc39afb263fdf747200bd6
z61ca965f3b175cfbb9d7c9f662dc729cf105ad48712ac7c53eac347bf867ce914220b04bab5d01
ze8851b451f51ce758dd3ac1d31e26acba19bd19e9f63d265f634fe57d1be0c96e31be872e06c83
zad5735c9bdf52e0121b368b2f0df76635e4e171ace8605f3a5b818abea15ac5a54410a6135eb8e
z039be7198386298d54f2755b88d7f07696a30351b87f4a65e52bcc88e1af1d6ad8d4f87d5bc6a7
z60ea70de454fcfaea8b34b2da447a65badaf663517fa84d90778b97d9b7d0e83506e17aa4bccfb
z91a919fef295964b649e04455147d3d1a542209340dd835bc5834b85d1038e752fd9b597b13717
za89c3f5df4610ff3393859d5ac732ce4ce43612d1e041bfde3414431e9326fb05497b6313c8c4c
zbb16089d5e5926ffd8a78b960cbc2017c2da35d5306bbcfa1ab131b30e037f5131321379ae2b5e
ze17bae969c89d87297c3a6e33978b6078246ee6acf9f85a7154c67fbab27a433388cb54dca931c
z69619265978a2df1564e45d607d49d0fcd7d414c680fc88e4ac3b246512286034f2713af20bbe2
zd85892dd3c1651216f25e958020fa5891654248f308f42ed61603043d185e3d0e6dffde62268e3
z111edb99184f43571ff1e17bb118a766600a2b06ca6de98eb8536cc46f40593be7c6028a6c8289
z42bc370c6c86bbbb5377fb4ffd6139ac29a60306d51b583497251a248255238068cc38577b86bf
z57512b90d4db27973e9166c4af7fe242a7b58bbcbf223c2bbcefcac25f95289649434085ca06c2
zc39e84eb182e8c5ea82d113d7c5eb27eb6f4638f5f03a90312bc246d3895258503c2efa5b8aea6
z118ea553076d2498999c6938fe06fe83156cc71f3a82f66bf4f99b343771953879faf70886d6fe
zdbe3b1be3ec6084f0b8b0cc0f1d6d1d44cce9178f8bdeecee18c24ac7a319476788f0a6a48117c
z6caff5a0cb2d0fa2ddd2ed1b1ef7527e61398c2d2778a85b7ba34b5ae16d081e4294fde57bda97
z2a66f11d66b40da3ca21996d548510dc75031982d2f417846393be9bd9c5c8b198bf50712b9f80
z29e96d0c56da122f485abc7c38cbb605d0d71e0cc4d6cc7a0b1ebf179867ff851038251bf2c39a
z2f709a727a524e9d35056ceec0e5de80c8eaa155db83d77df723681a7083612d18335216b2ab25
z2478c17e23d569100eb2f8d900168ead333d19d6dfa8159915d8103e4e2b244bc46c6d32eb3010
z37f13e65f405d2f122761cceaf34afea4addc4fee5c0d0879b3d7ba1bbff9c0f90e75339d6b3aa
z79f0810b45330c4c3840f8203d7f56c0b667e6cb3a7ee6598c0370f0d7a11f6d650580e17fe8eb
z654bb4d9dd8f9620fe555913efb2245bc4c7f6a871911b583fe6a6a81a047cbd09bd9632e688b6
za5d24257607f05539b8b307e93a841909b8175e36c2b6d8b05ee091c55cbd2eb2e4098f0341b53
z8d2e7cf42ca0e896c523aed6640a6a44176deecdcc765ccb2fe87e5b543958908138cf51056185
z83e7a00e25e1289831e40610ddc936e0522a5d01d7e4095434b5769d75d40d19729c87ce63d010
zc44b15531f01b1fa075ff0965b3535a2d79b0e4a7e5a72284fc02b51cc77ab62e6f3d67eda2b26
zfc49ca70899ac899c503a6cafa559e34d9d0a1f645beaf637cbf75eea59e0607ee95c7a4f58822
z6dba5e64ddd85a868a1f5b491a59f308240dcc9590c85c7fd8741b76de7e9b2ceea25b0de6bd72
zed605ca494d50c3d43755b6df37b39ec7d0ce4bb0f725c5f872c61bad34b08ca37fb2b80a2cded
z4f28a2589065d0f3f5d3be8d629c7b37a0e7bd73010b767e9ba163c88ab45160b709d593b2b077
z7ebe0b5c311e67c73386521c2f862dfffd1d740cca37ce5c3b45573097f992fdd2917be0a47aeb
zfcbed9359199845bdece8e119697916d4c35b9c621b13add9886e7de5c6f060ff46f60f6c385d4
z57143f10153ca769f573c388a2c564f53ce8ed9a5fe143f521bcb38755db10073cd27313a9728c
zbc05d4a06efdca307661a1a7803dc62dc2610b0f0c94320eb6051305fdd3b5a801469ce443d2ea
z9ba8252d257ce443a41cfd070e2fca4413a99d57ea7320af334513cfae777073a2d0e6745e74c3
z4bb8cc8c71a3799020bbb5d9e267668d8d5a27a3f2460e8cbd7ae09c81e047a8d3aeee38255c83
zc14cf7547ec5528048f27c3ee2384c62d4d35e5af8feb945f3fabfde264a78f45f8b1d12b7e860
z12127811c7d05f73f004a80527ddb62a931f51e62a2ff9838b0b9ab17cc46b92a2eadec3691fb8
z93cc10ecdec1fd5dc350bb8f7af49aed1eaf054ca89084fe89316774b3cadb9d97a6a91d8d7402
zb16e0a210f1f7bb04c07387512481ff7c80b49ac404558f030a2e8e08c14bd69ec052ba37fc37d
z966b155993db073c684ac5558737d0a8efadb7f0e6ed87b63e93d048ec67167f691275736ffb75
z4f820017806cb509e7ded78634aecf2d89e30bb0c72db7e3526a02b7a55e3c1e556d64b83bfe17
zcf5cbc2a4afd4c73f7c62b7604bcb5924fe6e18726c8350791a223593246397ec4fdb04679e7cf
z04d198e382f740461be46cf04bbbee81a0cc4398f3cec41612f5a75f992b8fd73db94236e4773c
z8e4c821a8970308e322f39b849f8e1e09fbe60784f707af9965aa72fbfd02a9986fcb6f1ac8456
z25653a9c8fb4d3c301032293308062b31f3dcc1052f87911737a3953d60068c6fcb9b36b793f03
z3ba0177c1e3942914fde0a3e6b11bd939966a0dfae3c9878efae032f5a38be26b5a9e3cedd774e
z5c216ce5345cbef4a4196fb5c088ad7346dcb7f28805d34fca8af8290e8704d2bee0076ee34519
z5f1627f3232ac56b8a640c171d0f72464732d0df940277626e2c45c19d49398cdef2efb92fa75a
zf24cefb671dfebda41156018885f2c1e6a7db7342cc80841c3101a4306aab87adb78dc4126a562
z13d1bcd2a610ba33fe76fa4ccb67d976bf4f82916f6900bf319e130ebb563ccc31b207e37287d7
z57604a2cd584a9995e07f5bf82419e143fa4088c0a86fc33556067be8e24291498eb05210217c1
z99be329ea6fc52661a76d2930cac25ecd50e2f29a39e92d0182b467759daef8809f2a41e076967
ze29e12996cf343abb8d9e51b3ce8aeec0b4ffeca473c38418ddbe528679ff37a495051fad2c069
zad01e45f860a09bf10a63d221551da75c84d9f440947fc2d2ece7633c718d7fe00d16ed65f82ea
zaa58351c4f9435a44f962ee772a0b71e8aa9e6081c9f70f545d88c1ae8237f0b20fe9ba7832742
zcef987a8e8bf2d4380470e4351118d94c9dc0fba8cf3b114a2e79072de570751339eed4743a85b
z1a844d869366c661ef4c3c51208a483aa69387e10509a5b664b72652b7d3c6708e1816ecc56f56
z33c6801beca69cee51ccdd0ea6a7d912a0f64802ecd3bd1f46591fad657f29d7d72116bdd83782
z18339932634ef01d4f516acd07273bc556b2ea7806c9f29043584e951043a85d0c62ddd8322bc3
z3ddad8af3f423f8d5db4ccb9a5fff3186ebe60cd306b5a7fe5132cde94e86a3ff27b55ed87b426
zca3d0f2f774101063d41cf3302ac031a6fc2ca9c631900c835dd9838d09bcb59fc1ea42ceec413
z85281f377f7f462e961af6b8512a01fce663c4368e36b0ac6102f92dd9bf47584e2f9becb748f2
z4cdf9726ce0259bdca4c66d5c9d8b877d86c9ded6253eb97e6ff04127b2f96caf1ca50dabdc547
z900b53b410de8cbb1151e85c5a006d0ac0176e9af720d2264ccfec7399b46c3c9d6b95db864cb8
z6069d9a07db2bc1db3f9803aa82e8104b5447f94e08f26a815d5db6016c0392404529ebee84b35
z595e43c51655fad7508de7e8cb8a1a06a135edaea3446084591ce6e492dab794ef1fbd5fda30a0
z8ed9466d1db148c66b9a829ab8098ed31f6abc0eb25258d7848a5b048a9e1339bca68193a4b665
z4d24f148c228a473d4e2b61a8801ab070333f1214c275511473c78fed00fb02fd5cb7aa6943e61
zb2b38110cb85d5462c378de5990513360a02c8972a8a03fd4a1a23ab4b3837931e0cc64f99c28c
ze1520178d19211288f9b9625c1e1adb40a2a1507d358aa3d4d7da21396056c214145f714c1feae
zdbbdb354baa5ace6830e3f3ba52a5b9e9945f222de4fba4385a0db24845718b49d79545849f9dd
z1a0dbc78d1e4989ac43c50d2bb66521637a442f1ead80e31937e1949345e1806b6a43fa5dd8dfe
za31388936a502ed07beb0fd60d245927f851aec272a584dcc2c5ff8099b8d65d5bd699ee42fd5b
z6dd90b6fc0e7d6e7c1d9d697340d6ad71208ed20d884ddba0919505df8f8073c7ae2315d54d7aa
za0808900de2aae1e73ea402f659db2de852ee8af9699cf96b51ff6f45e4b9a0c1136fa144db8e8
z0fc103c9fef8768275826ca53098f537882e5a1f1bab89b26c36bbb0e589b59077efb1b6dc505b
z8dd83ef493021004e8264bf2ad1368b9489885c524df166abf87aeffe5094f0a1535ddf8e96647
zb1bb4c820cad4dbea7365d9a149f2bb4200ba7df93941385b3d9587ae7157c05c24533bb356ad0
z0878e22bb24526e4a70258233d1d2a433a9a324a727feb0a24eb312dbadd231067bb0c4f301fca
zedcdde183c9d8e8bc92ab8a5f8a80414629f09a84b04260b68368b8b86794a97646d63151f250a
z166e38e78c252fc246fa63e0bfccec453775ccbf033ddeea56619d6cde3c1e0f3ccc9768f7d26a
z9eb62f2d1e69ca7bb1be53f0b263e1ecf1719cdb2747dfba84a080cffb634583d9f62f25cb04d7
zb0d8f383b2c38214513ee9c2f966e0c0da611924cb89dfddc952cd56c551ad0eb2b5f8980f0258
ze4f73cbb7dd665a34d69038a0da9d3364a73ce602e86704f6ad5d5a1be3a89eac4b5f2490d3be4
z04e068942559b63b42dd936c410eac1d1b3482e9091b7ca21d50ccd8ccb5e143b6939613b92eb5
z06de0e9f78883dc2306432d8166dd16340c3578215f310603193ec6bbcaab2416e56f791b0e8db
z5b7a41eed024bc44b952ca19f55a119a681e533e0816efcf028e4f9799e2239ae9cd5d77aaef5b
zc84cc998efd41aae46ce1815db89904bffa98adead82970e79dc885d52406e9f8f855e78aadbf0
zf6deaa077c45d30a49a20cb4139fe769a01f1601eb8d197b509a62f294ed6db2a187c05d0189c5
zde27dabd42b94b0413e606f03bc25e5f880f4118e0b03fd82330fc0f220528601de2181dbb1378
z1aea6a3ce4e77f468ec06da22a648c71e071e48e95969fea599896c0c134ab97742026232a7dc9
z662d223e19ba44d4d1365edd3b6360f62a338c6fd6ba8defc3d3c2516535df2a813903b9530be4
zcf5bca0ac301045abcc8fdfe63b0a412b0912e78f7608a6848d9f102912bb386389b767798f446
z4049dc79928893ba7d6df4dd7d09f25c880129c95a345db2947eea482cfa33b8c12705908f8e7d
zec92e4c64f64d4e74c30d38b3be7622ad8957b7a4d8b839a11c911cc31f6c538deb4974ead8704
za68e2907b82e16aa83a593de346a5193d95e6d16ce11ea3ae63826327e92084d65c4c6b3d8f9a8
zc1bc89824b8f18bcec8c14a51dee18938105255c023b5c357553f5844fa88f20893c5d35a9422c
zd406b503f36f3b8552540cac0142c6da4d9a753bf10010c6588048b567f26730f659a96221927e
z605c7ae76eb6f09c66dc88f0f4f87d22672c36c080a2aded5e99dbdd81065e1d491b3dbe2971f5
zf38401b19fa641f426f54d29e79a8ba8ab0da9438c99053f313a9c716e4ed49f4a520c1f0d0eaf
z16d9827c9d5a0a182aa3141d31534a1d959d4d7a1b282a8dbaa9a6365d1cf81b1238ab879a9244
z52258edf151ce55e3b7b41a3d12229eb5abfb0a142cd8386c05180efaa996dda93d2b29b027e21
z98601edb7b381d39d8b19f7893fd5150d48971a0cc36741240e4ea010fa6cb458039fb8637829e
zb90e4b9cb7ac441e6ce46fb000ce4d875174fb8d2a889af4fe7c7d27d03d180e1c74e9392f9cbf
z0979e3ceabec751412f48564a7e075e951307c5478d9de5c591b11c931fe32dba5ffbfd6ace529
z79490689a5839142292a7486257102e55b8a17c4ca5a5434e46f10133bd4a7b409e7c69fb8347c
z3fcc671d84f2457116df7d7df7d71f06c908e5d55e1f997c83bb7e85e9936923751a5141670fc1
za0ed482d7e902d3ab0a22ab86ac736cdcf755aa11e3b43393daf4ecc42daa9c12cd9be4928cae0
za4ac906efe564e5168e141e5a66bd58e102569c78748094dbf7d36de9789763d6a6cfe2e3079d9
zb49e3054e69cbb2489f48bcc0c3264bff82a0b08e5334480f47fac658cd91237084e85ccfd645c
z9d3efcf398793963ba37aefe3e1c607362d1389c458eb954a9e9b85a9f7385fca191dc415cf546
zb8969bce797d53b017e09881eb67fd745c2562e056a35148f5d91360c9eb362a0ed96b4d696df9
za5fd5a9f1b088a6f21c32000181e6d46e9b3c666e90bd9c6e1d0d5b811d90d4f33ee772de39a9b
z92804d45694af97f32852e2f2a1e43280bf7ab4c41e44253e492c15e4dd3f1b19fc5252ac213bc
zc59d7fb90cc5742c48e6c9a2fe99a31c5cbb5b117f5300f292d7037fa1c9d0d4b0aff28e7b8164
za43bf25d67c657749aa2f525b75b5942122a0df9889644873b233067867f5a06f0205fb9466cbb
zbe243a2cd02ee9fff388efc86dc3efd94c3d4742d15dc6347862c59e36cb61990499e354938bb7
z2d1e419e594679ca8ed8004bb714ba95783dbe669c9a834d46557b371a0f9b672198b5f1854827
z80678aa63a86e5a9b840e3b6808e98053e6db5c78ad5d027b82951a662566621d3de16983996d0
z1cd33254ad4638a0ce439f512dafa19b90c5de7ab88c634cdbcb56baaf6da903f2fd8f5453be87
z62a58c0752b138a5691460fd1d1074d42c99cc40327be887a446dee3976d61f537a1cf57c7251b
zed1519b93745eebad3184c25a1cb9b9f41df5b085730f3587c33c8868bf6a8793d2ffcfef16d53
zba19bc446ae9742f8143acfe20970e945d1399cbec77e8bade37a8ebc383fe809c11a2a64b576e
z52f8c67b01010c06efb7676254eafa6ac39f0c8a4c58d07c304bdece1e4a94d0e1e5c684293184
z2ea2b88f04adc9174475eb84f334495295b66fcbd5810db266c401432974de54c053e8becf4126
z0cd61b07050c395664cfddfc7c2472647cda1b2ec36d0c6e7cbfde699be046c56d3f5dd8c69260
zb82dfcca997c8f849a85a73e1c0f538e24b5fa786f269b1e2a3ef53173ba2f792428263a3d59ff
z46e129deba01e959a453aa965e2940787ff7b4e813421693f70a29581e5f37da56a1872bb8422d
z1f7a8c768746b0a23df04cdf6d2a53d9476e03e109c50b77b5972a28bf09efc765f2f9a9c9f2bb
ze5a35fc4bbfa26f73b8d5923546f404b98545b8def04c67de924da1569831f62dfa91facd75f12
zabfcea3203e828aea6df99c51fc05ba84c944e7f434983ec652adc12b027306a578416e13020e8
z2a1dab428290098da5875ef69a3c46093341376a18b63c531615367541d39c0c3938fbeafa69fe
z4654963c90e59ea9f84e0b35711d25972dc7ad100eb45427e2b32d1e2bde1f83ebd79b18d615b7
zd49d186108e9f782ec8010c11391e6dad52e6186f47f168bb902cc78c0078dba14f0d8d7990246
zef45717b72238c5d518672164b0c5425e7a6dff323891f2d0c959389741d502269c645e71543f7
z7d4dcc2e95bced9b0b4854942ee791d06dad05e66b67bfca562c9c1e4f84e548b44a018ee04582
z8d69ca5ec0999c317c4ed61f86e68ae5a6340d1d376f1e9ab2847d754f18f48e3bb4bc94f9d824
z3d78b126789c40fcbad90f768dcad5f1e93dc6e4ce75879ac2f6200a03610320681721cd30c1d6
z8c8e26da3352a2ba88d66f9a825d6859039949eaa4354803d8a2e733a0a193a532c93e257fcfb1
z2986c782280ec20140e82a452969ec7e16270eb41c0a1347c48d3808b082732de5751b06c18087
ze1b15caa59dbda71f5fc7758854fedb48abe092082580ba97e50d1345ac2c145c9b368e04f88c6
zeaf26dd5d57031ca22b50a426a21b73d7b206c10fc30c8ab65f78892c1b87a2c51ae92928c70e8
z496ac165582d280003b854d7f500dea5f1c93d331dbed2e21ea7c737789be8ce7426e8389d0846
zbf289c96c1a7d9c5d52bf891c72ab0c8d5a65cd0235459e1d3df4b2926316ba963fa921753d8d5
zb3862fc2e9edd98c067db60c9f3e249db310b776f61b69bcebf1f4f16368e88f1cf5389952f56d
z7959bd848a256d2797b0fce820c2f1469dbbfcf36f136f9b738acce4907ebaea11533352751e94
zcffe6fff828967001d5c67cca1204ce8b1ce8e8371a755275575ea1979543e7b15345203735bd3
z61564e0c33e249b015a0cdeb9acc39dd93fbae66fec4e08a48572350478f3c9553ba41a3cb06aa
zf2a39277890f7759fc4c503237aec6aecb63f1988ff090ca584cff975a3440e99317eefb3ba85d
ze45d07d6bc1bae7937051f3207e7de312910074eb71f25caec20821b79c38a8519ad88205a8974
z49f28538fd7248c5fef26faea30f81e1e56963663ef2686928f3fa68cc23ad98d1092556d09af4
z4344246e3779e3f444befc96af238b5a80f0c1003315100f4bd48de17c9e22d5bdcb8efd0cffc9
z7f672d54c215d915f937f72a3ba94009ac3e572fc403c7ff91833d3df8dbcac79d67a682a9e12d
z2ee65ddd84623b03b69eaf08d04051743d3a2429120271389c06173710437eaa6938f26e0724ce
z888d6d01a6a39fce9755e0d7767dda751eff6498a972a019814c060e39b8f53dd17f14d2d5e067
z2ee713205baa71794f6afdf176526a2f9073e3e26a806e2a8df5af51129943e74ae6bc1ba00f2c
z20e01d4f47a633e00289ec9edf4232d9f752477dde026addb9b61233f605d3dc62320290480d6e
z95782abb27037fe7458ccbf5138c742a9780accd7a5665ebe0811a77674db0b832e64f8da4619b
z02a56ba6972964aa3a77abb1d3c4631c60d9889ad0be7e4fad38d48467b43f4aa6b074e62d1519
z250377e4800aaec66aed30b0997b090a40fe0303f6f129a87fd68640614be4b061e3dd8e04b619
z090969647f9dbdd3fbcb7db58ac96eba9b8088f1e02cd59b5fa104200072653d65a0fadeb70672
z423e6a789372cf19fb08b16894cf891996ed3278c09e2f65d84e70a2d717988e8feea0d3024476
zfb3cae3fa2cbd28c5c9f2a104d343ef9f254e5200d90173ad05237cb6a675b1a5ab1288f341b8f
z6888c7a33dc3563eb0c2331efb2c8af20dfca7b0ddaf8b3b501866c17b4421527241f5e7ceebcd
z5a3280a47551fd9ac4d82e74bc2f50e946f95c785ace8cdc0d56a0a50ab0a2c79e3f6ebd0bb896
z29ee7647693cf5f00e4c375f92b5e85b069e13963aeeb3d0fa745fb443547d6366dcbed1a2ed04
z70367bc803f2c3080e222384028400e8f19f3905e942773303ed5da0751cc8414db13ff42f6214
z7c79b77d1c42bdf6d4eabad08c22b1f902da58aaeae8cb1f86ecc4350e88d8f05ff29719a887d7
z8766c9c77a868cb238f8e17bd42a73c458785a677ac21034322384ec6556d9d35ef99bd6a553fb
z42e066df8599e92845199182506637d656cd589f6f31f70b2d23f4a462501de5775413e0f68b29
z66173e3a62da5e65d69bfb262e7d8be712df6d799066e7c127c8e7d2ccca8a43018826aa589987
z14c44c1eb3edc02d00c56f05e41b2977d4f62def8d18782487c93b10de6d03c15385a4bb483715
z20eba165638346e836d4e46b27e5f4ced088292ef03a2f2009399810da3e1a02fb2d16854c81b6
zbdb09315b2cad78b93732067d683aa920b99717d7ddb26c2531eb5fb2315c0d675376f04f18d71
z8d46af3f12191d8305c57fb335185919b22b19d61a590e6cea2d8eac7b5b9b797123ab9f2825ba
z9b6165e5fbe8358c891ce3ff6722c19dfb6fc1c82f389b689c94c08770d011d62eb12ebb753668
z12405b1cf13e5f1dd6609a4737e0d1464077894598f57f807ffde20f1ddd32348232c42eee8fbb
zfaa18374bcfb3e795e38c67746733d657af78a3a61d767d4402e14e380b5da636ff34c55264011
z58e0fd1bc7db258c7363cd7c7ad15648e55c92e2f6a279f57ef0d95c580d2c842d64692b3e3fe3
zebf84f98d626309bb2346f0c1a053cf600ca140d39bc9455e1c83e710d440c7232085dcb3a9e26
z4f5fff00aa6625c6b833f968f5843d91904607b025105a6aa045199df2fe6eb0e9b18e40bb1b18
z4748271664c2bc7c0e8b28eb1b83399f105c7a8c6a33bdc67963f8905a10d2f942bded95ab05a5
z79f6a97e139aefd503c44f5ffac1a77f89a8a4d2bc241698b4ae3af2e6ea29c09e3b896d8f5362
zd5b90a6072a91857d092cb28c167c52976b7340153e823cbd5e37095844f38747285118ccfbb4e
zfc2b09a1b41b83bf068480718c299fc3cd92a7def5d407b9c173782348cb6cb230950f60477f0e
z37e7ff3ab9f2dc7166651ce7733b6ad365311945e0084a17e1f03aa521f9eb5cd88dec6ed0ad03
z6efb2c19354eccd5bb1bd0ea4033e4d6d39230cd4e7c418ddd9ced0a9bfd7d093619e71b2af70a
zc63db97550baf8749225c606f50dacf8b7f5e28a21c31decb247055c5f8b9d168b0ba244767528
z9824fcdd0b08c2d4571b34112dc00914f73d0853ad84f96beb7d3d3032dfc0ff8132b3b17613b3
zee4be0d5eb24f7860abe7f35fe013705702cf37ac94125910354ee75a399ebd58696e4e5fd0631
z0135272d3084aea11b9af3dd27a5d5af96a1e08b2898e01d23c62a1a6f8194ef0899cae5ca6f88
z27aa15efbd475295d557648b443c7d148b356241436b9dd9dfba945ad92d8042f3152d9a7877ad
z2b03e65ad6e582ad8f2239eb4beb91d320a600664b815c44ff60db1b5bf827800f194181cd9a3b
z9acd70bb819efda79f353cbe5619d4f572e86042cad32aa84fe8c632ec38bec4e76f19ac466711
z5f3f37d7949f9d993f8827501d765006044fe141d5a2ca7dd07dd6d1a97b3acfbc77f594884e47
zd709edceda2f57fb2cd5674d51528a102dc2afd26106ec43d40f7b83be2bad68647068ee4a4880
z9ebbfcd3d186495cbe3d430199eca3f4c6b2c81eb744125384995498ef210e0600f1de9753f557
z91c882d1efaea28f669940fab808a979274162c71849f4fbb7b03215f5735f98bf285668dbe5d0
zd10023670cb1503cff0be529efb83d5ec3a6ee549191e88022449a41b31dfd91f7de9f4dbeab7a
z530ad32791fe4804851eba97fa2a027f1496db4cd6fcafee1278566c705c1854af7e0d27480f23
z4e5fde601ea6d7e35a3ad877499c2ba68f797b632fdce565ca7d256d607e8210c39f6095f93784
zfc9a149c9d0d531ad62269f2730045588c430a45817ac5338ea0fe62e16196857aa696587029cb
z9df376a4d7ff3154f0bd9967d4e8673e39235529a6307e2d1079abb749d835955d39cef140d68b
z068a943a32f523762040cc03818c385ed34cab02295db608c9fa5b683b819eb489f2f6eef1526a
z9c6784bdffd095ab9acc05e1b9a6996bf6411bd232ad0df4b4215d7befad8092fc3f99679590dd
zc7bdf0c634559f140e93d38337b74df12595c973d6028062677d1d25aa77974b377571e2128c47
z0528df6da464b2012201daed1f53fcb216f48ce68460f62497cec63e9b86bd52c7b3f04d4a085e
z8f5e6e76828804e530e2f4f51aebb3743278ef84c5e3b3e27d0bf006fa5a3bd5912320d7e3a9ce
z2df53c2031f176a5abf0791528dd612cf215536bf6e1b33733a98663690e71063869e7c0f9fdf7
z2679a5a243a902b4e67c0de00223f972fcb67ca8345fb866c464900e111931f3600669c703d176
z1d206c4399c4663c03295303cefbb16a7fe9ba067598a6567f9656fc5b6efa5436ba164f2fd4ee
zd8b94d6fab523aebe15441ed524250a6a95362cd0a66101d24fb465d1e1b10c518e407681f83f4
z216e13d9110fe10fc79bd7ffba6961eef7a6775f4223156d3ffb6f0abece11d5b09700e9035649
z0bca035b60193c14d6256e5343bf826eaa792cbbf36b5c00cab15476c31736fdb3d1092e561517
zc76ae09a0e816b39d1b174f4eea2f7b62b245e83f9fc45458435e952613cbd1d881df0989a5fb0
zc6110bba85849f419c17f7a7077311f5d5fd3124740172d65a8ec8249cb5420e3a8e7504ec45cd
za6c8f79384988fc45bcfb466ae9826bf87c045fda0194a081fbb0ee4549c033e9e3ec3fcbcab3f
za9de97f2bdaf121ee0a26ad3087a926182d8e2779b8a2e6f2967d9417a28464ec7d00435be01d9
z709daebde2034cdad6a5acdba2e45e7354330a8f99bc410c690e75c40bf6e764d5aaa8ab02574f
z7506609e02f0d2dc99d5752060f5340a81e6c39aa37d1df2c850b05563594171f3259d77337361
z7de27f2fafe089248706ba79403cf1925a93cb47c40a7976eb3eab99ddecd329a7740f72970442
z73b3b27e6fbca4ad89a4f1cef3848a1bf017571544c5c51c5aacedc8edddf6a5dd1c0644f1e927
z35a02b63163e6118bb098268353f6b8ab1b12a50c578a42dc1f52de736d33d910532021e7bb46f
z46b1aeebc36a0c091b1ec942274a609a6a91672693eaf3ce670195e83ece10ca802c069493f679
z72377d66560ecd9aaedf76ca0d2e9c6e980f510b4c857ab4c6ca242c7ce73b1c9811be3336514a
z951379e50b8eff00a753e3e113feb9e1d4ad90e33f98d987cb0c164a63ac76722c07dc08236b08
z5d4282f57e8dd33a0bc0cf6f9ef6512f3e89f209b2d507f1bae8fac1db4655918da04030f88d4c
zc0592458f8e8a31baca3ec99b0ffcd4dfa4354f664a28d248521c6817267faba544bfb44d1b683
z5e26d8dd33a2c50cc84a1dd18bc5b6d2169d48b734951380e02d81d436337cfd032508efdf1d4c
z2fafef5c0d3caa435a54ea43ede6b202a600b2384728c83b23cfba2d42aceac0a27d0fe87e7a7f
z914071bcca17178bec4c0d189d90ecd70d86a0246465395ed590b6baf72c53a338964c718e50c7
z15494743180c84d4fa56a8e58ee50a91565261d3d070625156e0210d7afe863c8ee51334bb9e0c
z05300a9850b6a05a4fc98d95cfba9514808d188a9fb796132358f4398b922ed6c31b709ebc5ea9
z0d06b1c2e2f6b32cc6dbbe4dd58b3a519e269e333ee4b092459320e02ef2e901eb3edd48841f07
zbc842e6fe5f79fdf4c8b442ff3ff2cdea241f6ba37442c3006664eb320b8c9cce7e4e85e15cfb9
z5e169fdf62805e2e0922064bf4bae0e4983cdd39305ad461b4a1de46fa24aa7f974fd695e7bdde
z0ef8858959177080b7a768cff0ba36e177d7df8a11277916bed18f2bcb03d7757cdc718612f09a
zd3f850356f9b952ed37160cfc0afee85bddd32faa4c58b4a06a877a75e27f0c642b353b9709878
z529a655f382e28421cfd54b88616e54b2599284c19aa6666e645ab7c2f16adb8e3281301536bdd
z001b2c63e04605d7046c9074d49b6107bd26ab0d3e66da35786cc6ba167eb82618e0d7b3993d4f
z5391a71cc78cee54688abcdc7bbaf03ccff866d5ac95ae0f65a859b73d06ea18eb26b73514606b
z732195f341c9ae6ca5eb72fea129394c3487a830303548dd193d2d7600025fc2cdcf3d62e4988a
z911f455e7ef19d09e71c74e4e857c15d6f9d1c2adc1dd7a105deb6a8316ce29ebf5d950702fc21
z5a2c21f1634c0863b76da797b7efb0954f91dd8f9cf99709a81cbe3724e9e8beef25dda47f9140
zfb72e9f370fdae8993f92210b37bf8ee424ff86390a554f722fe0d5b7f677de5e7433f721b3118
zc9191dc1d69a61a685e21059d72c1615f71d2ff8b77a786dc71e9d63a43079f7213e942ac6d89a
z75b182c5c3071b7dfd9cde38a92cbba386b962865aaa3a3cc1e71e8794adfe5f146ea75d29c17f
z5beaf33ae43e7b0c755cd5aa11e37f219645bbfde3c23e0ec89948c2effdbbbf3e627d77445c86
z0cf850bd7ecc0579b5629c4b1eb8d440677c6919954b0ebac31fc12e5d44cd570538d890a8b3eb
z83dddd113ed4bec83da9cfa3c3e4a45d28430dcd4682780848379d6060cc811b34e3e388d5f5d8
z0ef11d3f8c71e991ffbcc00df536374d879ad1807568987a6e8630e763508aeeee93efdda23d40
z6578451f229a1524ee72829d37bd74c680237cac5cfc66a2e39d88d2c994a4bdd7a59044c4da89
zb2a4a170413dedda81b613f61f4be1dd43c27a172415a9ba5012d83d8aee466f600475de131897
z55f142b1a96580ea4f8fc0d29551bb36c77d0602a273af4898942ab6837f063816a4b017c1d541
ze8d377b1a23719ab7912f7fd04bd4de402d76851b6faa6abac89b20f58665e4f2688953af48c6b
ze59ccdda06b61f21d70e052d9664e058de74a433dad08a9082b3f61f62328fbc2e758607307397
z33154d2b2c83e9972c573a027294b47b0eea5c04670966deeecc8e69b3b5c18f41e0580a1e581b
z3aef8216dc8afc4a3a96de54123bb09d6568f6f1a29506d3a9ec61d38d285defeb970a00f5dc47
z933ab8963531036f9216bb3cf4e878c8d037c314354bf4c83e28cc0f417839d97a8a0e5341e49e
z611fc77d029061f3d8dc45dc6b248538067f1544d27fb27166abfb8b20221e56b49d5f05522a10
zcf141395478d7d2734bd3fe00f90802e2ace4053fc07c7f592b67eb007f95e27210d02138cb327
zcbd2989093ec8b1a4e15a18e3681a051bbfaf9a89106844708fe0af38b1fa69ecd1e20a7b8f450
zad06df4d410fdcdd8a40f662d063cfc5bc174bec73471fae7d6a2d4250b0aab4b668e6a83cd9ba
zdb31b925437e9c83e82f5d3ce48742be19482f2c35399ffb6340a3fa3e1906d933a3b84698457d
z0855b4958f64013b10a8187df8210b82133fc368f657e65a9cdb161621f6b431a679d9217b6ce6
z186b7813d4b81b701ec3dab5121005dffacae45706cc730b5e6722d7270eb6e9f92b03f19d5146
zd08668d98cb0e19bcf116464506ecd03037f4a5b7edca021f0ff22bf9076ca6a071195b8de80eb
z9e780ec6e5ea1a41a821e7ad454dd96b1ab63f5b8a920d1dc159431b34fce6eb4e553a8f775527
zb855c0c4f5f7333c252e1f616727b8b546dafe287e2b66b3b4eaa2892da65939a0f443f9859d77
z8153acb6a6e920b04bba9ab4282b788bcc1d56da072a4e62f4683d49bd471c94660dfb6a9ba4c3
z8942f0886906a8cac8eb554dc0cdbc4e7028fbcc2d0f6d2091fc8529098c958f4c313d11680af8
zf95da7f9f33c49c6e69d72ed759f893a16a29ab38a999963cf497d90cfeb0d2c83d7eb2b7cc62d
z56c4b1a1cac60536eb6b137f2a14649da1b4be01d514e40c98fc35e8f9c6b938684b0f7e587b99
z2da68e5ddcbee1f58a31f0819c6c13e244c63076ef9e20b739d7b7afe64cc4dea8ce9de9bdb238
zdfdd3a081eaa3fcc7e2dde1d19641dba2ff0a966e9b467d7b24fa1b8ae2ba678b5e0237eb28fec
zebb1d7d69d2c14fb8e333efe0c7f1147fb616084389c2f6edf0840b0e9a6042e15ec522cee12a1
z8746b990ac3d98a6a91bc84e94be41d3eb1d1ff51ecfe63968a75287a726fd077893091f34849d
z94074d9ea6d427145fe3d336dd74a20c1d4ea0075bf853800b2acf3c1a386ff50a6982afc01f68
zeff36f3258b1c40254a4294b04a73e3a0b0f20fd9feed066181805426bd7738377bee82eb48285
z40460d72f06bc1185ac331ed9174c4b6769a113dd7e231c9e126997ccf77d73e837cdae974a5d9
z9122a1465f2e6e783951c5009221119cc392f12d9055d3a7c31f6402c77e6ba109cd3acee4423e
z47c009bc83576f44a8c60066310cc0dec0b92c715620c829c71cb77af3f9c1281d3aff61b37e6f
z96c7976e37c14522c20054a8b2e71f4c633dd461c8252ad26f798eb3eed09681196568ea334a96
z39d928dd72a40cd1fa88a3af01654d4b8561fbde64654cda9071abbc28dbfc8dbccf484a9f76bd
zd2f23d1b6e603d2f9e0714bab00ea09bfd6d61008bbe30914fb971aecaff3461480715df363b74
zf93d0536558f3c69a6caaebfc39d1c958b38632e10209a64526f813dc91cd35044d20c1c1c12f1
z56771e8c5249041ff488b07c0ebc568568d10ddca1723f31be29905a03c377d67eb2c75d49c160
zc18c86fab509a0a1be1ffa5d5fd9df101eb84d1636e604c9d27400916665bbd0af89308833fffa
z31e22e0bd5a333c6bf789b77d18fa124d6424498ab94486bac04c489c27a885814f78b68698841
z95d95e462476571864c9ef67711cf240ff7569fc207bcf74287fd5a163a033994a0c0596c75ca7
z68fabaf2bc915f68c4c997403811084128bd40e06e5282a8a91b57013820cedbc1d4aef2d3e88d
z84cd2bc2cdd03f66a49b12addbd4e117deaf8313b1b46de25685d4cbc5db12d63675e56788ba29
zef14f0d5863da341efad24970e0d90141c95f2eb8def682ce31768f4b7b29a504ec55c3d0a801d
z732d67d0863e22f35ae21f20dc2e99c3f81b0d0fab3afd5df81a35fd9fdb70362e6f3982da4ef4
z524663c578d48ad25be975611c57d5429ba83ec7348d77cfe57f6f9cd9208eac2ce17a6b473643
ze0a67bcfd67ba2fd61a8d07e9b48e9e50be47a2259f443bca1f3f041ba7931651554dc610066e5
z54ada26e5823524bf4ae1eb71f1d1d0329a56035d3eb9aa6385bb08a5c4f3288d8d90ec9e96a4c
z1b4e56995989accb445896671e2890887a0ed56b4155eb9e81e0798bab9f791d1e789b8599d22e
z665477be03c9faf8e15868468935ed822387f00dfe00f143659ad187e245759b300ad56684b613
z56130e8c16ba820bbceac3f43b5b4483228c5fd5e3de0f287cf12626e1ad65684df616eaa97505
z7f6145c2e73c4e982ffe342e31e565ae65fe2c8b2eb2432d32195ee985bfc2059bef3277341030
zdde8362938caa699207285bbc5a15808929bb51195aa081f9fe6ca74d540c9ac8c3246a92b10ab
z758da80c80475b92b04692c66d1ac68379ec04e0cc1f5a9f86d51dd2c1d798e95c55540df8cb89
z36eb5ac98f39cf2e1464369eb3a1a2b475ecb8c17ce264163ceb4d1e3a9d9e4d1b8a71040fcd68
z0e76d2cd134b3bbb750d030c2acd4f0feac043ae35bde248014499a1014fe6c7c15ebc3270b58f
z759adffc738a4dbc48227d6c62a0a1cbffd303b16b6f088886741f65d474c6ba4a6fe17764a522
zb1d042bdec1bbe8100fd64f75bd24be6d281be2782ca4d1257677bb99d1a96931a201407dfc062
zc9f339d427c4d673cd5dbd761118cefa9e07d963d4da746be0c4907a0ac2c32b73689cef7aa9ce
z860c123bd9033a5688f24e5f9b885ecb6c5f0fe369404999771b39fd5cce48717d2cf3078ec0be
z08399df3680cab74d0c1544945ac9b4bcf1879571b79b00f06cdb1da7c511ca505d5cb9519c4d1
zc5ac259cf5c3db4b5fbf9ca8eead967a8e6d6f9d113aea2eea79924278de0946d83320011da6da
z402016d2393e5687bde163e888ef064cb2b2f98c17f72a0bd5a7973e8ffea6049008786703abb4
z5aa05e514445c454f3719f086c8e00598c9690cf999332fdf3edbfba3f39e252c4dcaee002b3ba
z87701c77cab6a494c09ca79cf95f72946dcf451bb21974d5345f2739e5575f7712df7e95b1db95
zeba0c5e5fe24ed6cf64747bd27ac83ec1477858863d9b995fe735f774e7e52980af568f27fcaba
zb75e3c53cf3a79a0b3e3cda5105c1e3f47615d081ede3f5029f465cddf93bddb7c49e3ad01e6d0
ze429ed47e0290eb2fdebc60692309604c021bdfc80ae9872dd9fd7f24c050337125bec8a0e7950
z04db87d7ef5be5dd2bb1a5e32178f488370e076b320a9072d006cd615b0ad52246272aaa1ef8ae
ze0ac5b9feec00717bce76545dbf4489df5124192eece1b56d259a6c9b524f35afe1fe180545fa5
z6ed2f4964b347289e3f83d1cb974fed9c63be59b883f81881dcdf47c2f60a92d33a9b0876d6df8
z8951b5163480ff52869854a5bb1d872658a0ba0bbe45c0b1d32cc1769b49ef1d3ad1bec2724abc
z275cbec0957840252bb55fa6c56bacb3f3d37936a2261c49ff2e131b3b3e5d3d9b80d8271352ae
z44dc08ff74462606686898bc4a84ef9d9bb526058b80c4a3ca3b1dd591bb7a43353cfde15118ce
z0d672dc326b8b81ecfc2cfdfb59ea2483536f4738f6fa767b551dcef6e2944f1cdad5a5ef3b803
zed13807620effdf67984a688ff40d152994b087828e3bc66a1307bf5ab9d709964ef4d95f34625
z5dbcd135e67f4e21adba11e00739a1c74ad869fefac19f2f1ab8dbcc1d0d35d6ccb4a94b4695c5
z08161fa84829d3e6626556e5ee48221e2e23b0980abcc1258d5653cdc573c6a3dd7aa5bfd6015e
zaf77d496ff7889b48bd16a20b7ae28642a44526f0a9a0993422980f8eb873f2c0e33462b4ed4b7
z5674e0679135abdc0f2c0c77808059c440a4af00610d2bda3adaa67d42d803024ba213c1035581
za6f03350bb5933d3744b59bdb4bd78aca5793a29e260e2bef7be3808a39f685200b774d4416488
z33a8e0dfafbbdf128c01897c25080fdd5518df2fbc0937cf31babc691a7a3afc201a1f32dda6be
z953cc73a70d190bb206eba7a9fb525545a6aaf2af9b7c3f2ea36bdd4dd4f813c6c8bb8853c8d63
z12bd97ab9c26a46ca3fbe6b2655b59c6676a5d4011286c05b5864b6822b09ff3a9c67bc83ceb17
z0bbef0877ec03e88c83b7025e31ee74653f164dcaff96ebad1af347f9a00cbe402434b09fc0363
zad982483216a4b03907e842dd9ebf420738bcde73ec6777f5b756811839e2020b1d8ee3b35b56a
zdcdcf63e99456e557dcbcd2be16a26cdb219b91328d85b3a67b53682a4127b5e3faeed69378be7
z554c4d2ae879cf775f70fe9a77af4e2d8da034f67590eabf66920b07ab27d5ff92d2c1ef7f93b5
z49641d1f91b0d0fb0166b3f15a9f93c7705665916fda7466d0b5d503213872ebf4d9f8f3bfd8f0
zcc4370156786db3bd0c8fc8fd85e4811302c565cffe5ab56f6f202c3111eb6501eaa4eaf5e2dd9
z2d3fbf277c1590fcb4b87b67bb7860fa72df87335b0602a84862c7475608c7c349a88149e054b2
zc12a6949c95427cb13d81023006ee976a2054f2e5d2a04d0bf65098d401300e1a87c8991fe49a2
zb375fd9ffc73fe095bd7a481d0a3be6c8a181450f498b4a22b3a8e437e6533b9055dbb037e606b
z2461965578e0b207df25e95d71b77accc8dcf5c7d33d1b12b935eea04ded33e1a56feca2bbc310
z4e3bf1c8148a6873700364cbacc26756240e9239c9860b957e2a8a94dea230be9a439b89151dcb
z64c59c8d2e50cf22bcaad45c6a03c335153f3b93120cb7a266eca012fc0524a8c4d24cdb1c0a35
z9f81c7d561d863df8cb1631d39eeaaa88546a9be5af3dcb852e18a5ef81dae8e9595595768414d
z6d4db7d817cd7f8e2f7f5a84a5e80b2a678aea54bb2b117747eea624b598ddbd8d6c0aaea826a9
z088e59676ab4af0281cf19372d5250714829f7a3d9ed6647671961efdfb32e350ed6c80845e87d
zaca925085b66c1f1bbf510d095f148b6efe5edbe00eaeed5fa430be9c631146cb663e53827e060
z40930bf1758331a0dea9aa2c9a0c770cb5f1aeacd923a8e611b1b1f0046413637bf3efe83b4940
z175fea7bdc89048b670b3c87722fcc6d413d2d0c8c816e5323ff9953ee5ae31ee1a200230b655c
zd0bbb8e845be705b5eb7b2bf347ed2dfd09dca58b7bfc6faa7c95939b7abca51178c2a55f12393
za2cdd6f0d8bfcd6c826569a764ac44fc22cdd53fb7e570f7238f35899c32010a04570047d1e5e4
zd170d035b8108f5226f7813c2923d01f03eab854513dcf29de785e720980d6c2ee23c2b408e456
z39e534436d0cc36fc242f8b06b3e9295f5837542974f8f0edb66443198468374a40ddb0256a427
zc9a4a05022560f04cf4099bffd3808d25c557f38c2fd23810c1c8b45766110903b4db57b6e15b8
z2663c3cd24de25061b47d8ea11e94ab347aba14460e35355bbaf900d8bc61a5b954e653be97b63
z9edc515db5011a23ab89e8f160f52f5883f19f5c666697816ca5635fd81c760dc3146be0746f2e
z83ff18dceb7f751eb87096552d0c73ced75efcce16c6d67afae3446feb86ef23948dddb61320aa
ze504e513dc0ca995aec8aa29c758e06441b28e0aa0399cdb68b47dfdd13c364294b8e2696663a1
z0c04b3b027f03347a753e87a92553d83f12808e1be816fd60b5e0ba491403efe93f02bcd3834ee
z9537ea586c1c5992ff5c21846802598ef809db4a248f3af2dc4824a62cbe2343b33616107f3fa4
z0e2efbe5bdefa9b731764293c03980cc9201a1678d4ad0a3ae706c8cf48f543f02de4fc5f13c98
z43f30b6d4e25cfdc5a7117e1e73de2e6a056ed5b7ee81e98aaa7ee4257c686bd4aa743e9a3aa13
zf97fee937c7aba607cb793e37536d57c23ec9646310d6dc43c602d842237b6a460b92f439db40c
zacbee62fd7d004965fb128e194e61e75381724a0e26c9b91d87ebdadf96d1a3c466ff743cbffe6
z22e1b2fa04322cbfc7e2e27170d8873f866365c5b8a7ea9c52b4fb3f72d719a95ebcf84c8d9515
z4fa2391a047e8544f75b28852bbe8f78297594b4119d786a288eb24fd4671c2096b6114da88f43
z4b3c231a70dc3011ebb336e577e35c44592cec625d5b14f891ae9ec58a6e3c80f192e533d4442a
z713cc9335b1adbe05f1c4833f7ce6c378efeb0ed32f883cf17aeb02551f73ee0b732db75756a2c
z856729c6e5e5210aac688dcf8e914c977a75bc7ef203889db0ccff901ca7c74f521c1c5cd83e39
ze2325d941874a14689e637420d6ba15d9529bd1ac4e72dd1043a3d80394ce970fd1d3ec02cebde
za45f8813fa75bfa845acc43d84f3e759b154539e8e6552105d917fd2795942ff607e3a9d4b661e
zcc35de0310b60990bb89177b76e27c0affa13782a168f03f667940f40e42ae96c5404042b42e5b
zfe45723dc40266248ce69f10623c31e5e37494ecf8db08074d9e1c91f38ad27cf9fbc7a2037393
z81cd5923aa1ce4b4a92f2066e2e40fe0fe0104b6c8851e78421538d9d07eabf968f0f5b2e630cd
z58279b45a3b4bd079f13d22e8b974dcaf0ff3f1c419157450791a8700e12608a15b80f455c77c1
z887f3f10e8117c758d6efcff096a637811247f48dcd0fb9fbc821ec051e38a81d14afba530c400
z6ef9c5676f6becf3b75322803d05bdba3c1880b53216bb50b9eed7ec4088c1d04a658329d28feb
zb793013e307182f62ec7cfdd61c3267614894d47043d347dd52fd24851d7f448cdd8c7d7a1c365
z826cc6bb5ac736bdd7d3994fe17b7b0bdff532ccb5076f5423eba9467216c7f48febb922a7cd93
zdbc9a32a1432e129fe7d5d2139a3910eea755f143ecd71bd919b1ba888bfc067994ea8fa7cdaa5
zaf898ecf573d67a18e710b79bb97fff7f8558141b359a9f774db39a86704b6e40d0b40d88fdb76
z7f799df447d8455a081eb7974b5b0d56f902a5bd4c6d0e90d536299a3793b97f4cfff606d36919
zbda754cff64b5e1f82b7f26d74296be2ccecc929b9ac0416d38ce712ffbd24b84c96c8bd2041c0
z2f51d0e23a175093d185d8c94a893f305aecade8cd844b3c0183a07460b70b57df272c8a362fa4
z362a346dca0878826cd7ca5a0c20bf4dc1bc6b08445aebe6f22b5157772355905de33dca77518a
zb17247e6868562df9bc4649fad6527690894918d18d9f5f433cee24be5110e5f3544f5e07e03e9
z69694419a7fd6ab7416f048236dad4b0926465a6996c423414a1600894f5eb37e9da765a6a93eb
zc413aca73e923234d53c5a8965f77933c94fe7cb1fc77393dcf7ec9841852a0779d92380f17a26
z2f046b2a195f4a4d44268759f9d62270fb0d63b7a92e0309b54e1b24b3f67843f0504c0e96e69a
z2543db8b15f6c39c912b995d5707bf1302744dacf4556f3a27e25319ba158c2f071ab89664295c
z9df38eabd440188dd92640d724498a1a468007b7f266a760880d95f0d9c729b873e2227994b598
zc99549aadca47e19a106a56d74149e4f22c9cc09c4bf1107a654b5c17a68358c8d44f9cae2f292
z63d54254f67158356e972b6f0ea330e73c8469a80baee45c56cce07c0d8930afd39eb910cf0dc0
zea8757502bd60bd5b936a0b028a1a320cbc5e7386c78ab00558ec7fd8fe4ab60bb2da33003312e
z2aca3d0436de4d20b196924eb18cf4807c52669ba50c4f5431bc922b13d3cb8b034422bf92bf22
zdc13606f01b41a4d335a197a7004f69799dcc62684dec55cae9bfe69e8185a2c5e88285feadf73
z47002e06f5b99add86263d4b6f768e51509d2e0e29340b70a594e33fcdbdc330c41ee54535fc8e
z1416e4b5e6da2e70f5a2f2d49e3bd3a2013aab0b5eca80d97247c9ed3cdbed52bffbd46d69d299
z8a38928c9a3b1242fae44f20865a25c072fb55adf2c457aeae9b0382ab2587f03b9c2d63eeda4c
z6e0904c404e79de71a193c5a93004629320aca388fdb76de952c6fb013ddf4b637f46e74f54046
zdd84b44281a7d6b5afe4c477757fb7d164fbcee0a32c3e426b15d278d0dc6c66765dfe27dbe138
z44c8cd2edf650b8be0e7529f19f48fa2689928aa9f3e62c981d70d9b120172dae48b73677597aa
z7a132ed4960b046da6da5f0c59c0780a6cf9779802f5e0219a7a20f360fbaacd0cdb6e2d286511
z762318a5f6cb33bda20fdf224d2f388da024635f496a95ea2920be007af4b333b899283046e14b
z827499aec6f0b197742434918a973af7161133d6ae16fa7ba250a5cd5ca126765f5340a0b89e06
z30e1309d103e82e2d756281bca0b1cc2e203f958fea4d097a42daae1b33ee28e2e9dfbfba2ace5
z78e5bdd6129f2f3b67a2b3a98bae4179d55a949ec55af844da73d57fef79203afd07f1622df3c0
z9c5b755f47ab7245c7351c1d6493f942e1eeb46bec1ecb67035a5b259d65e87980a992fb069165
zfb67cf4223dfb586fc0016ad2bdcd27afd174d7b77080903bcc3377f902de30f8791e67ab8e809
ze6459d2d02b92f2a048ee235ca57d2f503c93f4efc258d2a8ba2f06def3028eac49f58ffcab1f8
zcc0aad9fe2aa303b3ffc537efd6ced65e6a0c40e131848aa3438ff83167b9526edc3dc18e5c545
z09ff66096d1af30e92f29b70db9950eb11f4d3fbae3d28cc296193b632694551c0757379de1f1b
z872c5663b2611cb754f182a35e79c653a99dfd8d527e9848de8f7c58c77b3330c75c33a54d9542
z7ef2821d4c6851977d05b6cf8d7c944cc902c5c492de5bf5f628308189e12d22d964579717fe35
z546f200e1a918194af6d6db7a7ac9396c1c1d760ea10d6826ab813fb002ab5f2d53a9d5098d7ee
zca3c1471fc1b9d7a51b949d5e9de618e08bf17ffed69d13f8e933891be5595f7e68865f67300a9
z97b51ba28c49ae50f147d5abd85da1f1d9167df4dfaa54a742e7a7628ac67579a1901c6c931ad7
z6f4c22de35c75bf7ae6e277b9ff43e269260d791b461636d35b2807a86d9a31e06118dd8ddd1d6
z78467381e26e384b9865a92bd8f14ba94a58d4c43bc46bb6fab862ac132daaf2634702e2552bdb
z52e5fa7ba57745a4bc482cb7e1020a55176a57d0ab97f8463fb6f4da979325b03a44ab6ebbbf22
z3fe0fc88a389abd8ca283d3d8dadf2ba9f2bbc7dc6a07d5ee84deb2f87260463b5cfef5ba3db2c
z7b0891bb838a2edc5c835ad3dd9cd36e38980ac201d72c4fc80792a5620a3ae232aa6abf16071e
z22ad7189a346f160ff5082d6dd48805776fefc657c15eadddad09b8958ddc340adf750b737d86b
z27d6d8c5c08d756663fd2c569d9ce85efe0dadc55b32ab3a787177d1daa580bfb04402d2b263da
ze1fecfcf0b23078cf1b0bb155087606dd14244760d3c0bd9b3b9aa9e47e1e6fee11912b4cdf8a5
z84feb86c5518f275ee3e498392db3997ee554822e01b8694102e56dac7041ce4ca0c667a0436cb
za5861f17e1ac8cab093064c4faebd0a316d2671b89f3d456704680e79f0de7ee7c3958f0cb4160
z7408e6a81866825a4903303100abf952ef9bc9e7eb5667071af1e86592b0c35d29bae7bcdb5d8b
z7302244c1530ba332238b34773dde573119c5dce218a410332344d859d90d7691763ae1be83bd2
zc64fed35d1ea0966d871a7bb534a7c10e4e1fbb8e2ec4f7310a042d8cf0a454997238e123a026a
zf9076a163bb74894965f6d6659b45f839658ccff06a314fefea518e300178e2ef95ac251f7d1a7
z3dfaa9b322490738678153cae03b0ede2f922daf12642bd2b28d752acf903ccf9ec354fde8c2ed
zb1246d07859dbf8209279048727fe3bb16e2a4c7be8b9b24763628fdca26926f29febcb0a5ee98
zc8dcd1ef0e05ac10663ef4f592e3552622a83d5891c3573a447f03880ec63593f689dbef3d6d8c
ze50b59ce9d0315cb3e4f583edb62d37b1a498391ed4eb6f7fd814d4b2f5f4deb1496683881eb47
z8b1a47d9f3efae6fb870832af2478e88e2663804071c4a0af4adb289b02d1b3235dd9e4ab4d185
zeb397e28bd4720ba5ac38b7b9542486312a3fa5ece874afa617a205f28a349be6fbb388237e1bd
z0a7b8a9a8c9456ade220247535a7db978482d15b56497959e047373820b6329750cd9b0cc18762
z356f4009ebc58db1a5e249fb4b3378c9799c357d568ac0ab7b363c5f5ecb62e0ee90bc0e4518d9
zf96e8b6fb1a9582c150d3136c408415dd5c9278737e6f947b378f9471de36604f2fd104bf4c4b3
zc16a9a07a7c152b985292e8609dece40d47afc917eb7a27439bf0296466a0dc683245a6c16aaba
zd32e5f9eda40405fa09370236d9ed7fa462b490d8e181044bcc111f29a399a184a93f6988b295f
z7052907daad06086cb4e79b78102da03fb375fd803eea0e30319ddc53ec1facd6044c149c47fd1
zd83a335ba4df056ebb45c8ba2dc36b1d58aebc3e47bb92c290d8439cf199fe038aef484f5af35f
zf23610e422088790f695d4500f85e995fc383fb158d7eb872aea42b7639e7ae02062c8818650b5
zd092fc66159d2da08d44972cc4551c91ccefe9f0a06ed3f45647d54ed45042d3650490b81031d6
z3641df220df7ce1b109314535897b1cddebc241fb01c8d1a625ea2120d9951cf6d7a1d0b8ff13c
z5d4a2be2cecad358a292324db67400e9caf4c71f536f63743e4c896dc50cf42e61fd5d43024f3d
z8900cfe3538caef611c04816e038875e3c5db4759e1fa9923e4363da5b7dbac2158452146b9187
z2501fb312473a7c5fd521fcc0ad035fb85440add2fc43384b3eb83dfafe16b5284f23a29781474
zc2a8d686afe23fb1b956127684ab640c0c3480c6f7b33294d49375308250f71df9dc45dbb476af
z047cc32b28f66ea2b0ed16a6b08466eeec176a8a7773890ec34355990586a5da8e686d6700cc43
za52b42a1f5bcb725b11e945ca494cff04b6c15ae28339cb8a832c3316c555d62df5d3224275f4a
z6e6dcf8f6d3797bd38d5e1cb821551786b0fef6d8a70e0a4665174313bcfcdc5b6d3771baf4b85
z09343c9d90e4cef6be4e79d9f79097ea439050bc959db58437aa87f4d181036b0029b437f0ea7b
z21da673d9238b645468567724ab1d8017bd9b2e136fed86e0b073e3b1205358eb11f2e304f7a41
zbada5f4d463e32b74624132e013d1f17d6f8293b8c7a8f8815ab8f814e83bb534ef04127afb219
zde6d5f408bf3fe0b5b2f2a3ebf03e359134a98bd2becd6df77067114249919601a74337a2a0f58
z4f33c44f28654019efe27ab91d519ebe777681ed2d0e45c008160218a6bd6c5731f324e5393440
zf4702fcee068b3a28282a62218e88d9b11e2ced6df99ea8468b639c88226ac2bd85a6c38308860
z730a00704b507684c86a8157aa2681dd5f1ecaa4d5cc8b0d4ec5dc59ae9a9b4e6d98524a228d3e
z48ac8b94e7aad8be8e9ede517ceb6d0c51190a390cbda580fa0375163e4e30adfc719dc20c883c
z25fc3630c4b9f40d6aa0ad3928a8094f5a0226833f57ca7f750a590df93b3a1deb615fe620b244
z72f74f00602d6c32f447f78b42ad9e8d8997152b0e82b2bf04cbfb5253ad68f6b8398b17bbf27f
z771e24f6ecabe36277d261d66a2f14695dc8863736cb4b475152fa730330c3d605b63b44ed86cd
z3080f2690ea4695b0c7611391b3cc73904a7ce845f26679e24028170033c86239705253379cd3a
z0719e5fa3d2199b4ba069e2902958e2abe60b89a216689f3ef7ea105e9a571eaef72cb0b7a37fc
z0ff66259e1e3187ecb4df5beb8649af545307f6519d0fbcaba28b63900c9504f31c738565d2f4a
z48e151d8238391bb1205ab066fd3374738509ee264ae8d6a0f7e33a32932a24a641661e858ca62
zc86de626e775bec166f6e504e0292ed5144c0eebd2202a0ea4b405a220299b3943e096cb7c2a91
z7d7b771c271bc51a2d6b7ca5c5f1d5d2bb4ada6e50fda07e66e8d01997850577f3f5565ad39445
z89b654c014a31f0de815e564dc696edc009096a5c2f581a8edb8e8cfd63335b77604abebc1cf61
z8b6d0dcb0ee41265645c446fca41d519dd5c618acc676bb8cf79f1e6f6af857fea73f2e77931b8
z43d3f27598022e3999e8c3660a2e69493d16d794b18e4a289b1e7dad50320863a01a34fe79876e
z2e4c39b589f4a36024bff968dfeb694369dc327fca054a12ef3cde179066895391b9001804b54f
zcfe4df3b9521702b3c4618c0ddf8c992b7e9f2fac0bb012abf5ba87be43bfade51a90949e09bbf
z5b8d81c4109a07045215803b85dbb07a3150eb8f278ed2a3d5135764a90490c5b06bb59f759ee2
z3b7149b901cba064fe4f3ec267339e9ad809bd588b992803b251a12604ac6133a0cb0d07200b26
ze44392d8e8d42ea1cf0c8c23be25d0c5590003926fc5a513de2b0c52c53b9137513460ae90db99
zaab960baa35763dcc3c526a29c2dd16fbb39ebc9dd247da0e9592f70d53a38265061beef405b3a
z26498ff69d46788412268b862e7417f5fd2228c0fcfab22b04ee45cdcd996ee9195871ccc53cef
zf160130a74ad48cb9cdc036a8279dc2133888473e9eed48de81d463c8fce0f00763e83f479bf97
z3860e9c997e3afbdd394235cbc9f826b3450fff2a28a683d1bab40ea9134b9feae11d720973b3c
zac74d18a47a8863a125572d3cee9d9d429b03f79280d77a5da093d99905cd8a7c7255ec7f2ea6b
z4e67c1ef9d8cdffa2858d0a4f4c8f91925a8b3a3984ab69d763d56d0934acad42535f0f2e84fc8
zabaf4665080b638eed32cc9cbc1a4801f3dea55a617834f9fed612013c2ee9339712a31fde53be
z7de3c251bb91392586386f7d7453762172b8597a1b8bf696490384a9474271c770c3c0019d1bcd
zdb56b456999f59b11d5972b2127b5c67ed72fc01608bcba70c5403d287412dd76e59dcc83f007a
z755db9de4986312cfbaedebde29604d3e8771cace85927ccf0dd3fe4efc6fbb36c144c527e25d3
zb7e886d58646fd5eb08c21fa3e0a872076d4578f0076af17884fd4923581a539e98860f4eb2941
zbb504da573fb2de76d3950db137a012ce738ddb2fc0afbfc6cb3b376cc6d724517c9ba552f76d5
za83046e151e5480df9b4c6d9c8f0b4ebd51983c0fcb2dd8ccc4e6eeb99b89f356a24445f028865
z2063c895df5fa5ddd2a52ee2fcdf0fbb334082bde524a9c942ae05d5de4783c19c0ab974ef9970
zb4799244104424e99890525453efcc13e7d02e1c80c300b339ee2afa6cf4a7abfa422eaec55672
z0ddb9932c4844314775dad406500ff1ffa12360a2afcb558290d0af7adac67077dbe5188960d30
z04872ad3895855a87359a43a8ad01d46738c93a48db6a559dfef1b662b610a8b6c7f6b432cbc63
z6261360c0ae550517818bda40845fb71f4cbf1f1baac2760b6c9d1a1ebb0f69d4671747fbffd91
z9429625bce2dc2c1385ba555290613100ffc935ef934bfe000061099d8a46712a1605b0c434eea
zfa0f5b36006088baecb216546f300e42ddfd721d792a47a38fd0aa40568342e60da60abdf17702
z6e3c3e073a46da7e34915dd017398618f7b1d4d327df70cfce622b186b62f83150cf649ed5c4b3
z32637be5708a2f8ead91fad7b99777f55771c04d72eb41f1a22c4cab0fc7676cb2841e36801fd9
z99c2e70c655fc145f6e00ba9fdde1c0aab5da47e06710b85f363fb8f4a9bb34f4c807956992139
zc6906b6c52868548d2286bf1cb2c8639a8a5a12d3f20945a0ac9aae3ff8b935dec763406a0842b
zd731bef991e1e3f8f2fcaa7bba6049811dd508fe00f023af1bc382fcd6e84e1d47df11d3690a11
z36aafc9f07db4c30ca97be8ed2feacda04c1e3b0b0ce3df5da50431235c5bad810d60ed8c7debc
z720f66661d1f7650d12935dd43e5436df252133bfce3117711a5e6d95e2786a0526272803b9243
zc6a6025b428a9ce54be0eb6019128f86c83b5d4061e7c7e7c572c400c6f60c1682e9ae415e0865
z4d2036a04cfcd939ba41f65687ed47550f44e42bc210d09b2685954991677b3d5f5dc6e24e3ca7
zfad3c5adb8dc5406ac05d2924e126ae111a2e128c526b3245e55000e8e8664b43217c0955eda6c
z1d1202d978f05e2a8c34190a0a51b012c199a01dc8b67cd2c7af1a74d68925ea52d64c525fe2dd
ze35704a31c49ebc42122cbe423eb3bc53e84fe5e0a6ce54a390bb83824497a1e9910fcdd9b4a5c
z432802602997b99bdbbb1a428c92b18c4b317181b24d08f7eba4b8ac5e8daf227e1dd77f660690
z2cab15c35cc6f753c26b6042d3f4943727f25c67a654ace317148927aeff40d70424b4763049ad
z31db12a16eabc9b72f7171d09901c714e7529cd826c28c51de0eb71c2bf3fea08bc71cf2a88274
z162e72ff3f40589143ece0af94eebeab2291edf2e719a317f4100c4c621554826c241d3a71f8d1
z6412b0d16ad913c6b0943c17f76ac7fe3b4d0822d2696ffa2951c0a034f3597a8a795761483a74
z7717e28a7b7246e8802cab68a5acd489db35ba34dfaa7c4228c8e8487b7db068157b1b63d9c8ef
z4ff1adbd0a70f36349f170e0a9cbc384279e0223d128406f7787f55f0fa10ed28666d02303d8c7
z5b76cc29e5eb8000985672703a10a2c6b637b5e1c2e12721faa244dbfdc4860b5adcfdf96663f3
z8e75d9ecb8e3de03381bd8076980e3b50be0ef7766a9fcbf1290f364307034142896ecabf0374a
za50b9a6bcf9e2ceb7d0c130c8c51228f79680f5410bd2b53a2411ee64752579a131c868144e0f4
z56beab7ec6b6eea404545139beef6f496d0e99669dbb5f7211e5a4a2d7dfb48b1a2fae3e815b8c
z03b7d867b3c37629bdc6f5db4b354be6b12aa3f13f841342c62fa26d47bae81f94b3dcf580e087
zcfefa7f73094f60ca69f9fd75acd860fbff052f48ccdf551a80f32ec4af0f6f912fc7ebfabe15f
zad19fd630cb3a713426201af2f54161fb9414bb93d4dccc2c1bedc278dc68c17c1a8b2abc0bc4e
z6fe4a99dca9a822b24e3df4e26b2c04cb5858a820b0dec50c412fad70a29448c36a2afaf168bd9
z18b3878b82c67df45e1a01bf768d19c4c9e2d11f7fcbd86509a85bf27c9ea669b18316c07ac4e9
zee543a7b244f93745691dd129b01e8a366d70fbffa707f139c355245345a3ce2946345b849b1c3
zf83143837e9d7fceb1fae2148a35c2da49e85dfa1f4c26ed3bcbc4dd84a341ae55bc1c6b6e4e0f
zfde3be2001afebd073780c12bcdd7b8f5d99f15a928a521ecca0d35d22f46a11012c67f1ec9ad6
z58007e122bfeeb874230807911ca65db9c69d4e815545728cb87b2517d9e87173db8aae5809986
z356aafafb33df75ec4846ba450119932555d032934f00e5abb133367c1e869f42d05a67c63c692
zfa937b2e79ca267fa13d272fe208e23584a46af71044195748f23b5f6a38714c8ef83499a61233
zf614f6587425b7a05b79e808b4d6ee8633be34ebfa83581f7ba05f275a4e7da688d856ba1f3418
z613daa8a71f1436cbafa19633f4b78b476d96c7e5cf040b05e3c0740698b846be4edc1a79a591b
za7333b96ad7d3652757097957ed1768239a2ad216f73d4e191a281dc0e0cbd598067ec70d27cd4
z1d3d5f0082f04189937683e376b52cee67c9a54072a9ef68f54c61b55687b46a9b4701a76f5377
zeff39bed4b06c3b3034057637fd48e5e81bfd63074dae70b346dd3ecebd7693c009b124edd5969
zde5597a8b49dd120a81650a377dec60d32e40ed87435c46acbd5e1f564d63a0bfcd5d95a768912
zd0f9a859047f9d0c91076de1d8d8cd755866413ededd40faffd5c5b6310e179bffa5f26f969830
zb4c49fda3213535f14261d577eb443364f7745e9e65c0c05c9845422e8dfa9ac889368e8d38888
ze881cdbba8270a8cd18b946cdf378c5f10af7d068140d33a8a5ea66d064e536716c6560f192b94
zd9f6f1da58ee0264406e3998d396b5cc315c75de7ca0145faba3745ed2e407c7ae01933001abac
z3d8e300fcc40d19d595552e852b69379939bd34eacd976e8a3bc4a73315027b6aa4c9afe53fd13
z5d75a4b76c1dd12e0eda90057c48ef80bb3fee9c913a842d88d9ef0c390f270874a0ee03374109
zce184d9076fa81b645b33a4d101f614ff2f0e9c20db2ca61723d197ee576a155929587edca14b1
z83412ad62f416b0e310afbf447690c37d8ba51f11e8d8b5e810753f2867d67214a073d4ed1e86d
za304377c3e584374485bac78e4db1dd7ea75702392eb6e729cdfaf93158225415160babee79346
z8447e83c979992f9d24127aa4bc06ca0570f8e1bbc1b09b961ff545fc56c4de498648b48176510
zd7c17244646912042de0a24892665381163751f505d87389149a2c9d825e4a14d7b7bdf060066b
z589cd0e2cb7c082b7cb05cfa2dc118e44d5c84b6b1c99c34f452ae7184bdbc60e80f4f1a088d92
z17f6e0c402c57947359e802b6cd839338c764121218ce87612e67c4c762529177674a640d1e6a2
z9c1e02efc539ba7f981be2037b65d07b15c9cca1db798000a9abba865d98073404f2d27201e72c
z74401c8037d34d4398b62246f7957b486f18f350ab708f892cf9bdaf27ebbd52fc2e4ddc56d3eb
z591b5c950bf0f858586b18f96ac1aab321aeaea3278d98bb3110e4bc58d218c3e1f230d5504b81
zc4d483667cffb5a6e307ce1ea5fa4e1c69449755dff3001270c3cb0bff770cb3cff9efcb95092f
z2b1cce6078a256f6f4c6e2b5be795c0faef7b6212098b6ec4a8432e74e67ea830bbda2f27afdd9
z8a3eb0f6664f1201d6bec94ef826630db19e621dec14b97225325ca02e2c102b418b270cfe3cee
z20e7e80ab53f1f0c15f1e6b3a16d0b809a7d2fd7a005cd05b65dddd9f93f9e353eb72a4cf640d5
z1f16167c26f0fa1608e118f61110ceba9c328f847010d4bb3f16a751661c6ffb54bb77b136faf2
z14579735395fba074b044b75fb08acf26e89dbc8486e6fa12645538aaf1cf2f8268a5cbb9ff856
zfabf85ae497e35c6e928ee4c3330f21bd6ab55b5c0f73e4fdf68cd8ab96b0373e4f5fbac902c04
z22d22b91558634dc82574982b12c0a41a6326c76a57c143ae998fcb7c09c7edddcce8e2885adc4
ze5d37a7abbd5898c0358eb7c4a56eb37a2dae6375a4c588c3bef09d7617ac6b582b5b21ee589ba
z5a9f96c2dff65dd9da459ef0119f58e4f69600c6778db3e34adcf39f9377baabb6ef24015959db
zfceadaa981ac2883b302cc3f04a7b70c43d5a9481daacd38af57c7c8f3ef112a7adeed53c527dd
z1a60dd89a04a22140a2005dbf33059ac3e99592c3bdbfd1a983ef997482715823bf5b3ef5d1a96
z66a8d55af50a81f3751483f0ddd682126c8490835199077e848d34c03642e9aeeecb0e43fcdc7a
za68024902b61d72fa806d514f63a01b33d21e33e163747de2495f87666baea82bdaead407ecab6
z75b11bc6740fb7604f57ddf032334ab92a837825ce2ddd9526b2ad29cbdaef7c34bf62b1ae45de
zc210d396209f97695e3d36cdd1d3e60c85231f866e471b5f4e46ff177fccaf92f22e72da775987
zfb965625c7e241541aad2ae99750bb630248b15ea4596d7f6fafe809f34b669f6e577c97d043d2
z054a431c430977ce4b9ee5237024490715b534af507e8991bc65e4c3ec55b79498c6f12b079ddd
zd5bc8da46f3953b801cb313020b7f36b975b5a1b34c61497a8221c27339e4ff74cb606abb8c844
zb0a4ed2f05d7ebde7ab59a56b65470e6232f6129b7ffb67acdc03a34c9c7c537818dd5427db4d4
z4c1aa30b972808fee934d126a6040ae9f7e7941785ae5795e509849f04ae2fc3378969559563d9
z0334e5098c5fe307814625e186df327a5e928d228cf63ef5df246651dbb095aa85dfffc133a270
z749218dde6294285289a458e84216ac935c9a8b0ea72ef4acf296ed8514fd37f744f97bfbc352c
zcc3b26e8d350f1f7d07307d4884a2fa50397d9f2e95af4475347d9e2612fcca825597e2a6d6809
zb6a623a58aa4c218f7bb0e65617cab9020a18ad3a7856f056c775e752932b5c23fe8719aa65906
z74c96f93a78cbdd33580eb86112f90f8af0c3d938f5b3e085705f8b5b34e4d6e73a784b0c87e27
z79420ccbc072ddefbdd45c9871698aced7dfa022c9c3d3861c0421c031b2ea32ee11f4b2cc2487
zbb028b66aeaefd602c4e3156db0146927b40a26136cf8829c59b3c59814f1588d0779201ad9c4f
z2822b7595d1549b8d4a629be4c58532d38dadf194b85ec6558c39820c01b23819d12e532f1798d
zaf303839455e00e0a566bcd2a1334c727e4a7bdbc67c54a9882c71437960d1cd9783bd4f91394c
ze76fe9616e642a92ff815636df8d2af22d9113589675824cde75ecb058bdbb0186311eea559696
z65713f1a94a26819d03e6d7bca90b14407509f260af833c46cf677af10f35b0efd5d817e7c5996
z5df508d9fddc36b9ef8433f43c8839aeba4cad2edeb4b983f23046d355527befcb3265a1fe48f5
zdf0b5bcb6f12b2c79d6f25b321bda573a5a119fbf99d239457350fb6992ffd0d64aaa3b27c6fc4
z082e23300130366d4bde9bd2e30011c89c3195de9f10c8d248d85f1661081e1430528fda58fed6
zfb5a74cb147b8b6c561d0a6c1144cc3d188e093f30b06e104e1a8769d9237f0278690fa5b29781
zfdf6cd9998b420206008081ae501e43272bfff2f2189d551401f16514a5b8c54f80bdbfbb54d51
zff18791fb6204bcee490cb03a82326f5e7511c798ea1eba164e5a4ea496c786eac90bb75d44267
z629cec0bd02a949f09b1474017073c98f9acd1dcaf835d5bdbf0c095aadadbebb3846b23dff4a8
zc7c9ef9486cdb947ec90d8f58d4df3b7bf5724a7f4724b3f09b89ea0eca938ba78b8c267caa451
z3e61034bf947e02b1c6093f569e23c8c6000bf8028e06eb85fada66c6e6305ef58d1287a4a27ef
zf323656120637d2b30330b42d8d26108a30d330e3d696e7b4f1449f3e56e2f5adaafb059207ea4
za0b42babc530058759c6eca84df950384fe2833fe4d8eb8d7b796a6e9720284e2caf453cc7d7e5
z6bc02f98d9011b0cf625782100b7faad44866a7cff285f85b40e685bf56f395a960fa5819ef4f6
z0201c6bd133c543f31f74758052ba60e8c6594a2f97379a5df58304cff6e929ceb42bed82990d3
z6b44c5e057d62d1e23e67fba9b4a6b849c39bdb394829364dcee62e92cdfb86e781a75c3589caf
z60234d008f967c0bec8b56aec5974d068dc7ae1dc0737c48aa34e30da6e5f03f9d9c770ab50e17
z56fd2cfa30a673620aa8d6eb66d3bffcbd2d6f56e6edb519bae88f28f5692d35c85bb20cd5ef15
z5664904ee0f3e5a377cb005d965e4658a9a18033fe99991913628f6d85682ae14d5120f2d30827
zf5de267b748237bb7fb1d9027915307518de0b8a58a66c7452b0e0c8867a4818edb3f32a16c5db
zd1ddd7094688f17dc0ceed0cc36ee8d9419578ea1322e07393b9a4f269ec86a7a82cf1f82bbce7
z56bd2bba6b3a4f9c8d8a65b2f13e5b97f82096fa5de74a2881ab68e85ab5379cc0ec56ec1d2538
z000176922321a799a31f414be83def15eed052eed8ed8313ccce6e9e4c9a29075e2554f033d021
z2ffc28a1972d5f1e3aaf91981f1f8fd65a17ee9f3bbe03a3ec9e9cc9f43661bbe2f7c37fcbd582
z49e2814fa0f85fea58c8e9c07eb8b233b0e8f775c7df1f1e368ad8ccedabea4304104b631ab2fd
z9e385ab1c29e527a6cbd235b4515969f5711ef2bb36c9e827b086b640405aba4267192630c5f69
zb6df7490368d04cce43e79ea4bfee3bf92e0482d4d03a0788cbfeb3cc05edaadda80ce116de7fe
z99bf4e954b45db13f2b371aabd9428f8c46a30f9b9273447862cdf043ce760d894719c28a0e754
zc80098b87c9bb81c24d9400fd1d2c46572fd64f4919be501e339a0d3cd56220d6c10b279ea4ab8
zc6f6af5b8448cbea8562c64a6c3f91c8b3a2af3ba975d2e303c61cb67a5c8d968ac0b8fd084721
z297b677d3bb820d0c75336394070e1a1535d22b7be629136f314f61270f24cc10fb48648d8705f
z47022f1b15a5477bf307e36ed738f8441c9cb8a60df87265faa1f64ca7aeb2e33c24aa0bb4fb4a
z9ceb163ca2a3fb1cbf271f49735f94f7325efc9ffe4cc11c3ff5d0f9b26472ca343fd10881d395
z24e5984a7802065af75fee5c73987586ac6757e1d3bb5c43532e4f4a4d4f5ad8490dc774b66f4f
zfec29d19d909e6551e2c605393cb99ddae4e72081ddc50cf26768ca572bc498cda04a32128b856
zd85ddec0ca6ed924300001919a06578312094be58de4633b8a855000d42a2d050962c1c272b035
z997e6503d0791718625841d766edb0885f90a5742d18f8e3dfadecb8748083067619e12b7dcb57
z3df9c2334e1967c22ffa4585fb56c1ff0ed87c3f9f68df20e3cc34688008176cfb30adeb3ca8ca
z44605ff61c17a39dfb82ca97513baaf69b20e6969624ebfc1a325e5f551e8be49784395d57b435
z37e237dc86287984a532d0f1faecf622ead573320a8804c2cc8e9c8909f6485c3bdafbfb6d5aab
zb081e7a5304f404c6af918ca19f2ce36ff34f3139fb59c125ef246ba90d35b5cbccfade0674777
zaaff1bfc9b174e198ee09e84e4fd9e158445c97bedbc111d4c510283e8429ed958963d1414d4cd
zd933841ec689328f0f3acfcc4644f9c2a7c49d7ca12774b01bf0ebb55456fe425f97e31150d5c2
zba6390b6c66927c10a455fd6a6774e4817db4f8bf5d66ea8d86fd5cd0f9d4bee22e8a476915b7b
za8ca153e31214d20715221a030f26dca9684396b8378836f95237b1312d69e9a06c360ec3b20f1
zdea8cb61dfdb73c15b5712eeebd11854cdb6e7b6532d43bf3defb7320e2a65137c573559388860
z62c997869955da739fdd8ae56d41d59007b19a2e2eb2efba6492f474528bfe59a851d89ca10bfe
z6bc133c9e862ca6e4bbcc23987ca427bf2768d99a4c0efd522a2083a111b2b3d41bf38e868d84d
z0d166c0b7dfc23b2506a163b0bd38be3a851d835788d6ea7e160fc02c7c4ca8495b619da2c1f66
z96a8ee60f042e757d15eb1dd447df07d8512c7e566b23e06a90802b66a06692c63fe2f4582e679
zbbce10dd0d384b09c2c1c72569e3dda92ec66aa430f44a875504f6a242ed794b26abe3e4b28241
z755b06f1038d4eb01049eb7e18ac8eaf9e63dbd9b8f12a126fe1913723133f4d4f4eba7504e8d0
z44a395ef13af235af16901abf55c3496c154ee78d317d8913b228645443f70b654ede5f3d61864
zb8a36de69f6c008f379410c7b00bfbf54a193ca8908c0d95617cb8120e99ed8f937245b7cda952
zd16323b86338233e59fd520bd38e531f259fcecded5125f286ae7fd11a369bdf69c323a01c7311
z9ffa31463cb7f8f3662cc1a34960baa9a24ddfd79956e133dca7048911b7069112baaeb4f9e90b
z23bb6b4e6233e2d22fb1d59b714d44ebe59fd379c97384f8e093b76777c8b1ee6291be98a488b3
zd960c52017616d5b31ed3a7a7db9013eef955ba54bfc4b903f9a4317f6c39c66271f04e5d346eb
zbec13157cad416fd404805acfc6ff2e51d13df1bd979a9edd231816a615dfcb676658556e78e11
zdaeead2b456f1df36528235be1b0486b96cb355822a85f7929b084ecc265ec3198affc32d8f663
z131fe3bd8279da369edff521a0534a514bbba818c573ed1bd00959cbba7556f9e88c37ad0fef5a
z66888f06af53519b8b082ff801ac458c64cb46b28885a42c14c9fba3cffb7e85437bef47c86fed
zbc9f1915de5434bca355cb39d72855868c0488e9b6029d2575cf3363524c1b6a08fdccb840c14f
z72bc1a8c31189b7d8ccdea96b11eb197bfbd1cb0da19d9a62bc238b6d91f5a371bdfd7c5c76007
z3327051383c0b70ea0f926ba235fb32a7c48065def1a1a68c83861bf275d14e78d3e5d12fbdad3
z5237bd73455bc1c8aefc78ef2e9b465cd398edb613d8806f7c9ac457368b8208a212e121fd1b01
z11180669748155f96659fda7dda6d57511d154aa2b30d8bb4597c3599de81ae2d57d7ac03a0c4d
z43ab51e4a838078b6cfddc3abf4d967105933fc5667f8bf24961903f73ee27198141703ad64f76
z6b246058779f6cb34e12c93b7957ebdaa928acd0a8fcc665b706a6024f485161ea7f95c342c7a8
z36bc8538691406ed902189589c5b61f12cde4c43af650c2ad9c5623545edae16f23983a258d509
z302799c421719eefd0c9ebf9d5f0971e4d47a84de56e45db1115e875a627c9573385b2b231b202
z621a40ea6bd5170a9071093f3d942ab2034dfc30072f4d9d331d17d4e1fbb2a96fecafd484f752
z429c66a611bed79e12117e575411c20845471b7be12692f043ed1d4fb2f8ea01094f509c7990d7
z25df9a69e013afb891a3eb517940a84e99b51b0e3a76d71447a9de508fcd12d0ecfa0e2db6f305
z8e649844ecbc9e1eed40e97377e6d9f7eeea764cd701eeeb5a47c1a5adde6a8e0461606d615dd3
z6bb7114916857f0fd3b0b2cff5216562403948da139698136c3fd52506ac737caf20eb7d886f85
z813b40aff513345c630c76bf0ba4eb48e336c7a80b8ad6dcc424cce8a99465e3777b85566e34c6
z5a9fad691782b73611fab22a61ea503ad1bdf8051a62a24113edd7146eda46e72e844e4a3513b2
zcc2dfe004257924999daf1ce4d8892e032cfacabb6d850a13a31315f4e1fa5c3fc11fc6402d1dc
z2cf6444256d9ec31053574ce1cbeab71a88821679ddc234bc94fd22fa8f6529806ffc4d5409326
z46e45fe27f94496b05b0ca19022de1fa64075cc6fa83c7c8d6aacbaec96d6bacfcc82f53755580
z2d1874eef586be0805548b9d9c17836de7766ef41402991edf93ea803afcf27bd0dc9aee42b438
zc816e35d653553762cec4160ddbef6c00fae3291e6a29c933af93c3065c615e6128cc44e925c1b
z382bdcc5132d6ab77b3f84586f7584874c036f19ddb5b3d61f32b336e190b7f6f3cebb45cfc36f
zcbbf781f68cd5cf33f412b278e6882cd679853d64592b7ef5070fa7bdac7c0fe0741cc3acdafab
z490ec9ee46e6e99b8309f855b483c9e9a8663b13592a55caa2a6d8b3d444b934aa396bc838ae6e
z98736339a2b0358aeb36d6236cca24740db04993278444e599dab7dd2bd7804c028475c8ff790b
z373ed21d3f33bc2336c56d6f873974621e99757678ec92cd7e0bb1e08681a9ba34bb6efc769e59
z71113aa689d820695f381a19ebc40b4ba25eab48b1d131beadc1240f5654c3526e5709215e3e00
zf280182377b6e97eea5f039a28d3cf313029baa2c30d329fc467799c5c267bef9fb23af94ca4b8
z5e612d68259d3428927c14ce1e870a482a6916abfccea4054e5f9774b77046a3ceb79cdd66657c
zff26a36b68f78174a20cf882fee7f2350fafffbe1becd8920964c7fbac82179f219c9323871ce1
zf941903671a91d8ebf3d2825d2811e6e24684d35b0bb0dbce69ce98f9242826854573d044025ba
zf402bc2a10c0c6c897696561d2e5f30e09575e5a9011ecb0f6f72dc318aacb1aa36a884c4c499a
z8a757db9e5bf65bb86f34fec59dcb10fe12e70f40321e2ad8edc38be4f24b470eb12037cba1dfb
zae38f19eebdd1bd8ab2daa4f36f229b6d09b3052b4c7284fff5f19b9ed2738459a2bccdb081cfe
zf0d8b7f6cadd488e5e1f13bc38e05d48efeef417a9467df0f777fa2979c9215dfce3b718b5b89d
z029ab42f04d615766f6fc774aee9a11bcd25a7b77357b113dae0aa206d1cea422503aa8aefead3
z19f5368ff87cc165cb7ad62ae68e3bc70489c13593b8b523e13348510a9d912e43a00767094e90
z284f8bb218560ab38ee8fae470e78ad784ef6b0cd5b985791e4d6116279c6b63cd115f7d836e3f
z5833a1dbe40e6601bd78663b73ca356bf86733037c60283f3b50992536e719bf89f08f5dcb15c7
z1aa89ed322b4026809917d2302cade7b654b9157acf0ed7b0a2be715b9a33538c91390e3ab425b
zec843edf85357cdf1567201b2bad09587d8f27f30b8712d589370d5148aa4e8866cf08f84b2eba
z5404aaca0c80bd963f24796c70a9fb24c594f9ad153c7aa540e5f4e91fac8907dbdaa9f95c7e8b
z7ccc4bf525011b9224efdd6ceb69a3085e84a3e8a0a38642d34017b531f1940c3a85707933e188
z6d454cd3c04d25f2991283c14b3a3d2148cc55243356e0e2744c0f07d74230a7c5f3a312533d50
zad593a4f1fd49553f59077fc0bfd551a6eb9fd7ff237a08da5aa2127830f6b65f35b6f41dea47d
z5cfe8ac9bcf5db4c086fdd7bd39a03c5d34f3ab4634c97617d278dfbb4c1e0a425cfdedb130f6f
ze5285f896472cea048e37be2056dfc0cf0dd5e175a1e99715e0485f24864d92bc5a075b4ad2d51
zfe05a9024444cdb54d8ae109c58440f455dca914043ceda85e22483996c9c24a3add6ddf971a1f
z40658bed4806d1b4020b0d321616402aef5da0f60e6d16f975f4d8080351a029afdbec82edcae7
z7e18f59051c97df152c2ab19d400a3c14ce3b8dd7a2ea2d597b3dcd5e6c81f68c950a6a269a5e8
zdaeb6e2ef0a3f194cfb3a5bc05bcb6e81890af946a3ee9df38dd78c991f7e47aacc14e029af1ff
z64259135ef67c460b525efec5806b46abf9443790d2595a87fd47b156f5deb64a43387fb8ebbae
zd8387ad4f45d2e67da3102bb256c0e97244dc2ffc9a7a865627a94d93b8874e2d068e20bc002d7
zad2d54a487109a1481c32e017b00d9342f920e9b41f7322d2267d433673ae0513149a68169a5ef
z09d661d7e972ea315e60e6681d1ea72273df1c097d118ab9458bf7eede0ced7d117a20bf07b6b7
z9fc85463636bbdb1ca2c68cdc0ec80da728fb8010e0c8ca1986ad3882eb52bdeb7dcfb4efdff87
z0250d4546462184b110fc8030841351f29ca3ff0774d82ae335f24481a460a6c24ab92b082c6ce
z6d3ee0014cbe966af1f896421b6864cd3c7d883cb4aff384f94ae5d975595d1ff61849f9d91a07
zdc8c1e7d628d253859e528fdca9dfc0303cb87c9af7f0ac39b38f27d67cb6be756bf1fafd1b1d4
zf294bc4299a32e82991b909ede2a1b465ec2faebf7463dd6c689ac803f8b4238509079f12443be
z3d006822627a7f9669962f61dcf66bc49ba2f3c55ba168a2b9d9383ae63006ce1439ce4902f3eb
zbff76d7425e4e57a5d5a1cad075632b4ee6d71da3dba3b7b85b73c7f5f93063902554e8a4dc483
zf2ecea34e2bb839e0c72a19a921d75dbdfdda311353cf6ff1d07709b7dde40ef49deb2cdc16def
zdc8067457a0de2df2cabba16b7634b01c0577cbf0147636733142e38983b4458c2af452b8b0583
zaf04b413c2148cd2e2b5ebc7a86432e06af75842fdc9b1bc549157692f67f2d0174be4fd2dde91
z927f6b12bad290fd309d5fdb1b4e3f93dbf7424d8cfdacca522dab07690d77c350589461975aae
z3988fd300654e8521f27006118b22dfae52f8357a132e326cf659137a948aa9a2ef5d1f030dae9
z5f9f38e662574ad39f19f25cb645f11c908d7763f59055bacc5c9b0047975ed8b8dd0b54dbae61
zca2839920eb419188370fca5b95ee99d232427c8ff6f2c19fa48930b601640063273f3cd0507e1
z7906c4cdb894033286d2db232961fb60e01c110e726adbc2b697574eec5c8b15fe4cd34c9b1535
z7283d1a78faf29ec78b49fac37a87f67af0501d0de656f01485b832d956d0162a1b8da718bcffe
z59c2dec7bf79076e19219f9d14478621b37c1f85de3da178c91e4ae57ca947f98f53cb5f40ecf9
zacf726fe83981d7740fbb53dbfd79a68e1a9c085c274b1647c86cbcc5027d18a5da3f7a05c8103
z135caa4a0ca0d73d04a36811b0dc3eaa9771f491357bae552bd1cac61c3ea5b47bbb8827c2cfd3
zc93353e1761ab125bf8fa1d7058f9d3efa0d2c32694e0a45c95b242793eba6695f05e84df1262a
z75a1b20c40bff0f59438d41b62d5fc2f8e487c494ec62f763a17687ba7b5b5cbadabb909550ef6
zad17cbae75462b4bc3cfe19138412aea07d6aca1ea17efe3993194ef48f10a6a70b8aec548d2a1
zd23e292ea1cdc5ea3d09ba0696fdf5b135c898986e11b24ad63763a0911d8358d9a04764d434e6
zf658baae25987671635e92fd766e7cdfb26c8b8480325f271ad03e7bb28fd250dc98c4a5a30af2
zebdc1793c8399aa6d3c01dc854808267bf2b85aecee9daca12dff254468252bd4905c7b5452772
z92ed3ab4dead03d79dd28f89f455e68d2aa6d692b4ea0660a55d4a063476e8a5ddfb6c67eeaf9a
zcb721561e12860a3484fa56651a3cb5ecfc9323829f5be3dfefa578a3c53ed849122beed85d9e9
z9238868cc39dfa0af70de010dd8e9d483e674635b2a47b9071425fff988baefc9feff9c9642563
z89e16596309320393f3d8e15530d4453df79bf9c2a6ecd43da9d47eb7277365fae5b2482648e75
z4797ad37e17c88bac716e29b12a8bf071e0702ab8ca1898b1e1c5677ec3260061cb0c338d9ebf3
z84f0d6bd96fbd43e917c5f5a6e987f74a10d69660d036b4eaa69d2488f683893adc5daec96a9cd
z1f40120b61026f95ab0b439e2cb4687b8eb022f20b2048f98bd20e680ec67b18be7562eccc3ec6
z1098a36088586d367cdc9825dd567f44ec34448c37d935a19cf69d36941c6f8c2b7fe83ca78e9b
z9dc692e467f1b49a1683206ff667e2e1179c4bd34a5971c48c0c5d0f269647c8fd8c0e25e75924
zb9530b37ed8e374e9b528d842eb4c0418d6dd9f712179ed0055ac12818306ae91df3a592a31e08
z5bb892ebde7d4014c2480767c51c9f07ba356d2238e9f2a73676ab4cff316c83f91acd37a4ec50
z04768d7c114b18504a91ccff7d4a04da67f2e464a6db88de1e246fcb2514a1f7ccb61a40e68e74
z97527206de7cd018d1565b9219952026ae459b3e76d55ac5c068cb0d8c6e6094be0bb2b7a461d5
zd93f707d71950f77ba4657b541881b184f080ceb0309ad2b042339cd1e2037e02d8cbdc6be4a94
z38c28179531fabb66564ddb63c4717e5b70ff5b74dd7c0937419e80cb6b16fb0cd68743917bd04
z38f6dbbd488401f19f930970d2a5679a125eeae429265b540ea507d4e28ae87ceeae94bfc6585c
z9160dbcf40ab193e22c135689ab619618d8b4ff0a29c443c1ef7fb24efdfebbc9e13ac5342d4ed
zda7c6227bf5745ced8ffe1e8a2b308938737405f7b6d204a5826f417ab129cca0e8b21ed24f89b
zce26b753e412614d5f2d3e48622f92963076b272eb1aa227b6f0a290729174b4053503b3c87199
z8ff7dbf031c9a758801ff626d7b7d0b28cef833798cf3ce1ca8660b4af6adf7b87e861468fcb2f
z01e49f2e5365ded99c736940db476b5fbe18fa2cbc350b1ae8fa32bd3fec4872c1ded717776625
z9773bbfd958c3d0633b4848d43d1916e074ab67e14c59098500394e2395257e501fd27b460842b
z17eb5e1b638238c1d8f05a97c863ad6807822703787eaa9d52c06767e966d5f587c654122e87f0
z2a1076a6c5f4bcde59b437c0959681b6f0e5973c278099480abf42777b2bf250ad3e8cf58a70db
zb270a1b92d740331afcd22389536887f50f5972e65ec88f815c1a69a489ce61ecbbf183e1045a0
z082c395b13dd0b3bd8d746d141bd67dd7c48b63ff116f5352994840b4d962553f28805c9e7521e
z4754dd9d3819cde0c399b9c7c72a444fd844426af5bdb4e5c6ee6ae1199896cacf7e03cf443b83
z3412b0dd474298dd2a42134642afce8717afc99bb82e8ec608b438964a82720e24e28d4862e7a5
z16757fed83e21013ab7a6bdffe66446da6a5bc4d5f9644897453b1d47c8334b33640d44f00a18b
zef191722d2d875118f2d7ab32fc0034d4c8a4b55e6ef0ee1ed27ecc8f7f0beba96675ffc72a508
z9f59a8fae32ab4ea5b39256ee25ba7d784b6a488a0dc94febd75ed9a35a388b735af86a99793c1
z65f6d84d808d8f0f507bcde7bf45def212c2d3a4ef90db54de81542ac754ee3ee42f5865e42d8c
z305e207852d470ec3d7d04782361a4e134a9369250c0c6169c96daed59fde0d30d430a71adb2c8
z909fd40fa922c8e14c3c8c36c2ae8130bf7894d9c8a89ad1b7057cec5f821b673f52a4d94dd747
zcba2b26aef59bc19ec1e5e27497e70eeb0b196e7352ba0d6347ec2f383066ebb887684072d6e92
zcedd6eec07160f844d0c8ce6b33f166f6f6c0fc93b32fe0b07d5069b94ec0d2b76f97879fcdf6a
za6e038fcf971d750fb786f41b38d247467d5f85522164b374aa85273d02ace1ceae6ed34b6ad17
z138b0b7fdfea4e5c859c1a02578cae4beb0d2e272b832178e5136f9925f94be54ad4344b89f929
z59b31f5926bdcf49bead7ab41a0c9b6dafca1004f0927abd56ea73965c4ae778db7c93e3bdc6c8
zc5ec515f5b5b401fcdcc8ed14665cea490d393e8187785d8a9cb8df33db59d8faeaf8038dac7ca
zed59794ed55df60f03b659303f8495cd0bed7f98b07651aae4d10d254cadb1bd8095565ed8240e
z02994701e132832b4abcd77645cebb18031f2e2af8c920d7ce2dfc6a3d73f4ba086881d0b1b43a
z509e5ab58f251728b986a9bd72fdc3d728f4cfb679ac98477427b2fbcbea050517a98c8263e23c
ze10b3942d1d21eba300545cf64abb40f148b67169698bfaf2c907a71c895d984b9bc46cee82f60
z87c15d8ece1cbb698d0e77d6607b1f2dc4547b27913da99ab65b576de6f27af6e163d86f18d7c7
z7b9a41da8ddbf36ea01d48e7d7c549080f024b6bdc5d5c3145f33e0249e64ca54767464426337a
z40d89405ef74ae18e239cf045c13de0ad37860f5038b560d3bf509b0278d84c5200f14a8dc10b5
z0acaaf2c81960808af419ae3cbe2d45f3b48c9f6c2e5e5a280dcf86976456e6a6222fb5b466db0
z455fc6e6db3c1efa900f511491c887459bf45fcf4d79e491db80734234bbab99d2928a8b55345b
zc27ccf34b3ccc0ae44e8160adc5b75262bbebc32e7f8e67810905bfc631ba50886523a2cd0db0a
zb9be075db0d434be4d363cf85bb8f749c701612a993e366e1bd362a3af6f9f40ba011d455c4514
zab940d62cd61f69ea360ff818234df67ac033a37e54cd1558831054d31868b5aa1c0d49766b9a2
z3c9fa288f8d4678f909d5f7b6a313c3a8814ccce823acd76856e99053e1aa0724b7324b911bc82
zc5c08a8b77f103c80f416b3c6bcf60db9942d91921ae3eb8afeb593e0e255c3f6773444bac84f3
z2a069b178ef1f7742d1a5d4e5e1c8d15a631424bb473404395517190c06a152c257459abcddb42
z63b7544387221331ea00f451cbcd184d3e6d9b99e781283f72f48d6e218030c632d0dbbd6d6fec
z3deb7b399348a825286afb04c9f8e0a08d767d1771658f6ed894d8cad883cc482de756f977fba5
z3685d1964709cb10b0e5cc6e5687ecd04b7e5d40f8aed6c3b6be4f83899aa8800c0c884ee6f392
z90e034f84c8d63f103c91b05ee0d13f727f7dee8e933d456542634fd82887e7a661174eef08ef8
zaee4a8cc4dd4e141e6b7ffda41cf8471fe8f691554689e2e3b9e487c35d5626f98286dc2d9f4c8
z07a28cf4c32bebc752ba3a60b5fab5dc13638d6d639c3754ddb1d479c7b5802ebb246d90af45ae
z82e51d7af5ff52ff42d60658605282a4033d0bdc687c48305e1664484c3c95d5eb938fe3086023
zce345fd71742a79e4e8fb270894107acc8399f40ef3db5b84619cbb54da46cee197b74535f035b
zf4c352d4b8e0e5a5cf520557e31b0c4c1f789397edae1f2f6845e3d75515ab06c41ce4ad84ad0c
ze3850e1269eedca539733272ecf3285bd4fe99e15285a1303c45a02519b7fb9241c6293d9503f0
zbc72867997c9a9a004d348b027206a518697d45181d1525ae96a9ba786d9b5e285642a276a9847
z1909714efff7df2922d58eea1cee8e73beb3b319b81670eb5169daa02c2afe9ed3d78456c1797a
z489f9726c665200d51c925d4b20a1db4105057165544efcba8955999d44f9e9e04105d7691e0fd
za7cac1294e58d2b6d4be6b65219ea4047b9a636aae6cfa2e3738ab599d3fa365fc226cc60a2d3d
z7adf9b56ece938c2bdd520438b6f44d8591ba95c6671996ed89cb1f61f791bc4277992223f1fc4
z7262a5f37eb2c3c5c49bd179e3cf60f709008d204baa3eadaf37cfd7cecc847e198014315636b2
z7c4fc9c9fff99fd46e682946aaa98f04c324bab3b864a7d03d83ceb53a6b5eec6f0b98fefbb3e4
z674daf35717f5a29dbb6c80914ecca9df9d9f18b8db83241612d11265537dedb37b74a8f335fa2
z2f540d193ed973170f48e692128e13edd72d2d63fdd1383d960598cc560f4a4381a48dbffd8a24
z169306765e97c7fc57e48a492d746ecfc7702e09dd2ae44186cf7e05d166e1415483f022ff35f5
zc42a4951c1b8e9d93d57b7cf975b5953386214516913daf54a3981847e9ffadff3699771d85d24
z833558aca054db7e90b5206d06cd3a3a2b91e5bf99006364a2df41ed695174d798b6df492835e7
z1a046a311e7d45511098badc1c60d7d7793f63e2793fbb261d1a9feeeca1ef66adde46ba9a2c3e
z32027c9b73b5a7c814c30f6beb5d3f38e294e0dcfbfd107739c46acbbb6da83161c69094943647
zb0c637373ed38cde65948ada95ba6c23f8fd03261e5d6cea8fead8044b391ab8a60b1c2e31c715
z1803abb60191d38942ca939d205d3760d5ea92467e4bb34082b99fab91f3b1ce791218ff5dba9f
z095e51461119318cb6268498d0f08f3ec46607caaa52730164d2620b3cf09dd74163da95ac1631
z3226f59fa693ec3b30fb298ef06e62a7e0aede9a3da8f975482c31890fea57a123828d1bf9b19e
z21609097df7b60b5814a51a3e76c1e6418bdb009014850cc566d108854e3ab49d12e4b99227143
z5b8449402778eefe5d0dbd80b47db8fec369e5d485a9f885dbca742c8b73695b54a8168135e389
zfa6c0fda82570da952fa46155059d143d76f9f7762201404b091f239c144c24682e4e4f5f60b3e
zd9ab8a12701865d0de62db446970829182988f1821d4868c7807efdeca54378f0c5987e3595b95
z516c64017ac8d64ef6b2c03694d12e50892812d17897fb39901f7192acc8c1b0f531f5197b134c
z1f61a96517c60261e2083c54a57d13e480c9e35196fb2c390d02ff8e8b8f123a928a36a33ca8c3
zfc2f49556f37b989590d57839e3772793e53fbb55973c0eb303e43f94c13307ca4f7d900f5ae64
z1d4ed3c010a072a3205a8efa63667bffb1b5def57d6930e22ebe13acfe51bc68f3bbcba37b5432
zf58c3069411be2211ec7034a00492f65a05b09a32d99e60b47751bfaa5623952c7b7d3c28e9353
z7771bb340637c6c428022de67ce6a178618f53644ce780a742a77bf4cf671a8e30040bbc2e379e
z8eb08fe88962bceaea6d3c5b56220bcb928adc12ed1ae1cfe7765aebbaf2367338e9401ecbd4d4
z2159420eb10dede73c199a8a2e2868284e17a7a85cc391f375e2babd1e33996bcb5e85e157df0c
z366cdd0e783cd07c46021ac9d99d1fdc08433609befd5fff0b54bef7c6bf10a1f85d641f6d7fea
zc4c252fc09b93408002e2d132874ed9eb0c4739832458fb84baccb98e44de9fe4142b4e7f9d402
zfece984155979399be570ec4e564413005521fd38d60cfd15bead12f0d7b4cabce0270a9c17458
z45d3522f4eb8057903d3d2fc605f894e91aa0a18d5dab68834d0b5bbdea383f0621ccf6a1813ee
z8b6ea44a5c8e29f03f8ebc290539c6e1eb4182014a2cdbd0c43cda61ced1cd9ec7c8d03795e6b3
zaa689a6bc5880617adac43b0ab845b9af88807108b920b478f66b3ed74f554220e86b171456ed8
z0a0852dc74653bc0a28ca023354626c2d46fa0bb387c5f9f6e3e5e36effdca0b6bf2979b4fcc77
z5665aa7a1cd04a8e081670f42eda4ab97536d6be932abb0b4853099d390091c8c06aaa88ba25cb
zbed612aa6337ccea20f057647d807e9fd985b686d7f6cfc295ae07893ee93b9c7a3cbf350580d7
za7b9e1b91004cc0acebd214b07943b9cf3bf711fba5870082c6743afc068e1698217367d44ccf2
z26f6452e99e95d4840cef35c9073255a683f8c01511a09940f72f219ddfdf82c70e5f3f3f3431a
zc8a627f2fbc9e067ef41aa5f6f28a035b16d0c14d170ddfc7c75267b7ad2ed70e2a863b7e2d135
z894b33ef82eceac3f6538a4f25c37ad1ad22d7b529429b05483fb26ee0efa77ed84e84460733ee
z6ef58592e5d6367dbfc8989ae1eddd2ffac847e85918fab9ac0b92f6e91807e14c0ece6421b312
z4cd8dc39d248eece14db842b00e613255db3a12f96b399690164dd8fa7068e0a736d444d0a465a
z480719290891d269230e643cb8c41aecbf9fbb92ddc2087be4e2edfce2a632491b46192d915849
z91dfeffb439a1bb5689a88455222ef830c9231ca8d6ed8b45ae4ba6339bd6cb72e7a75c0aca230
z6f8e32c8b34b01c3e4a4441c448f6ef1430c8b4822fba7e8e2f314448602874186cf71d1694184
z3f10315f687678d1b3f79f61d8cd4cb35b9b481de204b930649089f82d3ae85ff8be8b9db0e91b
zcc6ef6d9cc3fdf93a4dc0860e114f525fcd0beee96960089f38f4aabe8318deb9687a299f6d52b
zc0b3cbc5acc38ba09598db43d181397f61bf7ac5d81c2bf5784493e2e9f40d6c1e4593f5dbac43
z93802c0878b7957dd5226697e554e0cef06a4c69693929fa0c80458f02765438a2a82741069606
z234fe7d44e5b3cd825301dbcb0abf208239aea8253887c63a0dbabf88ccdec3f70f032b34b929f
zf5046c5705577f79fd1ce667c5a56e5fa333301216ebebe67fa857108cd5d4d1a5b6dfa2fb01e1
z8309a81743144c486113e0b36824ff879c7d78eb4d63be3532b15712da9a700b2a00b64d7aaeb3
z24dcbeacc4e1cea9d84184adc8d5cc94e103eb77786ebbef8c8ffd7866f4cbf331c4a768084158
ze7ba56a3203b807b3887b19dd7ff1601c1b14861a189142491307ca4cf2389fa3220859db34bd1
z796b6350149fc4bfd269662dc1352bdd2b5d908b7af3f5a4d67f69a43def9ed822144d49213cb9
zf86f84ce7f30920c2498b7d9eee6b5660630ae766ab4603077321546da54391480977cce60bee3
zdedfb3989e329321d6a92e1b59134eb0921481ba0a4784a4c5a3393d1971403a100d4b441aac5a
z0e34753591bd689c3d8586ab929e65167f48e6ef5c0c5d0023a768fcf59edac483ab50da20bb0c
z4ecf728e5581c0f2b9528e1a44f0b3ee1cbd317b7b0a97bd210ce5fe57bdf0a38df7cdf59dfb5c
zf40e1b228be5eed726f22161bab94e05cfbc46092e651d2e37a3fac061a4b0f7e99fdac79246cc
z20c815f82591a301982896655cebaa40ca28a97a74b17d46d6800d1a421440d10bf59fcf82031c
z7b65e7c3aa55a541baf4bb97133ac17c88673361a17de7c0a157d701471680da0287b7c889ef05
z9aca98f2ab05e13cbccd62bf47b62285bdabbe4013d6f649ab0ab0e1052bdaa3a1bc1efda95bf7
z72c6f2e1d8253d23b222fbdfe7cf464c342eda1cfcf3d13457dff6c16eecbf735eb906689e22cd
z7968a386cff11b08225f6961af072b0af3ec06abc903f63e156fd40f82ea87eaa139227bef5c39
z5d1c0272c3f40a974716d1873b8b0d789b124623284882e56f6ad48610a78f7ae34949e1f29b67
zce01755579e0addc5b7c100a768a8d2b73af690b19d0e5cde187bbc8c4012e4e3aee5ef1c71845
zd4151fa658a51e3f570c8723313ffab6fc9d864989490a01803ffaa30bb70f2a2e70c1e7595b99
zfc14ef93a65649621df52b2615b4ae8dd7056e765df1165962fce2846d63946c0bc5f928d8712f
z3cef0dc80a2e10432ef38c47c92feca5faf7129842ef93451cd54207238470d57d4fdc803ec900
z4cf774e937fb77b763037d88d24c77c37387624b424fc98a2d2b298e02edfcd004ce89be92598b
z3ec75ae6542a550bac641f1bf46dd061abf2941e4bc02a51f4deb834468e7b75eab2ceb039ce57
zc0fd4433c7bf9df0495a684599875c600e3c11e343eb8a743aae42e75088ed981b783c0ce9e6bf
z40d6956fc98759a0d2265f677ba00dc37e05271d18de081470f6b0185d12daa1bcd21439bb0010
zd82ed7517043a8cb84f6df56491a67304aae517d61dec2afc2e6ef28c7595bf5dd39760a04616e
z9c5dd08d86043ff219db4dd6124345b4c5b29f9719056af8a7b2798dd8ed2db17de9411374ae9b
zf203c0becba6f10e99bb4ee6ca0b8a748d98eb20deec085c64f481c665c681c06a2f4f6a4eddc1
z2a663898ef322be2600843e16ff9816da2931ddb69821eb7d48e35608afbc2f7ee5031a67f0487
z72b432a0cdf286a32ca67db13cee490a545c6205af155939690317fc507da39b855c0dc69f8344
zd2d0690873353514482f7efe33672f2266e0c310b6c1b4db94e56c9cb63048719d9ace4b767412
zf2cc412d085002d8c751573ef834dbadc61838842417e28f0d403f991074a8eac7c0872f8ce2a3
zbd9725b69a1cc0269d15580d2ac9b725f4b746b5b72c70c7e7412a6dcc09be16b73211ff27c6fb
z847ed118cac9aca0410ee368c76960f6d4910c3f63e60aa0fb936bc7ad286e2e87e810a78aec57
zc7dc239f72191a8ff3e98572faa16518de1145eb1a83b099023c72331277bd1bb6b8e54abee362
z99c43d2697b8444be5d8654da90318333e61b8208e5fe6a9f219f5fc4b43962b5015a4a718db15
z5643b035b8fe0145c6620aba2e6ad62c463dcdc11f99822ca881c771cc644308c89c2f40cef7a0
zc629f91a361933d8dc1591fdc2c546902cda9b4e94d95989170f57c0cbd92288ff20046369c478
z690bd09720c2b3568b7334ec068740f08a7536aa023ff6584e5427d3454689a1a3b2df688028e2
zd0c0e59ae9f9cf74c0075bdd3a5a0e5d167ff50d14fdcec51a56d2498cebfe028543ed307be129
z11566f8558192668baabb4a8a3cb5aed5653814e5eb7a15c41a4d393c0677aae38593c0fc4dc31
z9fb5b4182528dbd1e9bbdd0f992a211377058b9191f3c34708bcaea49c082a7e5c9e86e7a3e7ce
zfa2150ae1d89bfc3a6a34ad85b1be61c3f9b0ae1486001fb42e7d81504e5f500bed05bd9487df3
z75086fe36c32cb37f0de4840f34b00100eea80cec7887210f99a861ac04d6bce5b774560aa4a0f
z2c6665159c8ea79179f15a30510bd2af9ee12c22aa049b7aa53c03ec0c1765f41d7727543fc54f
z0035566ce90dbaa62d5bff5bd92113f89139b6b637c8cfff594d583599462bbca07995aaf76164
zbee45185ee7200f56cd88402ca39e5e08712cb9eb8846a8229b992214c9ecfc0ed49113b380929
z57a4b4513e8942691644ea784a7ec09d93d0d37abfd394ca214785057bb12701a3298295057e47
zfeabf568f3071519ac760baeea54954453d916b93a67ffa99649e1bf83b7196c4e9c3269f6f16a
z212d8b35ac7a20b3e9978750d22081a5f0e6a1f07eefeaebee3a563a8403c5c6becdf1fb54bfe7
z34a31e6d23a2fd22bf19d5184bb76fb813ceb17c89f09333ac6c462a71a746fdb66637a404277e
zcb37d5132f115ddaa54265eb976a2d96638fd22b901751e1cce64862ea38a76141a259986b5698
z8ada7fc6936204420304991c9b9fcf1dcda7c7d410623ac6479d452abd95dc2755eef357e589ed
z8dd2ebcf0809fa7e81da9431f329541d310e0a15a2a94e8a6bcadb70e9fbaa709da8138857264d
z030cb7f188c94898c416b8b28fd663fb060613ce550f7a2b749d3f2719923797e4e6c10047a7d4
z07943b407d939473739910dcd84d2b7347fcffd94b2f7407f79f045b3262a8e775044fe6397a04
ze506d627c868d306d0b541d0f86229df35da67e63ddc572442444e6afcf84c15210a559200f5b9
z73cd8fae27b07f49af3e4f37de2d54a0104561fa5d12fedc6a9dd35ba4fa96fc598b5da1590dbd
z23236b73d0bf3ccd68d0bc3a7c90460328273a613cb15af3b8194abdbac7bbcc362ceeb2a5ca9a
zcb27f7f07fe231b247a24d25f44797dab3bfe855da266d5fee07752994e096f6b8410f717f7de8
z6db3efa1ae25d311c1aeabf6653a25cab41c89c05bbb878d0fe4e72e2a17656e47686339630cff
z39622890c564b4b10e2b2195c7ee5bce6cc740218bba5bfc9b4a99acf982642506ee136ab43aff
z2dc7d155197e95ed86ddb223607f45a5b717db560ca354407a8259b202485bf130c7966f691133
z35ee0dec80652e572b6f004ca4724fd80cb150f469f768b9d90433d537d037ee641eadb7de969e
zede6707290be12e062d4965709892fa1d0eabee24d8af8cce03b08b165b4798031ae7f755bc1c1
z0ad14a5ed525b1da9dee57ccb218f929fb88631ec885f0767a560428ff35ddbf755bb88948abf3
zaa884ac2d61b5d1f7c2ffee9876863ed51bb3e2bad1f36d552f1427871ee1df12fad0127a7dd11
z598a3abce6794e43eb0195c65e2ab514b21ae54e140d6214a7d22b39b369ec20417d85a38b6f44
z06097f61f58da81a844c987e744443dd684e3d2f312dcad40c9abecf97961cd493275d1bfb4712
ze92bf3a401b2e2f130323e2789427f92fe28d46c85a4a5cc57b85564321abcbb07452d6c036361
ze33701ca54b9f14cbf1edbf1bf3e0bc6b9d3e5703123e1f0d874cc8ad450813f91936201d3e338
z3bc7eb61a1373d59eb170253ac7bc75260df63906e28ed3d8561a73249625144ba81cd6c9c9eb6
ze47165ac43d28bbefb1692213401b4e8a63d5e56630882f186ca0718df3fa7fb53f5239a771254
z6e77e6540b24b13b181b0168905e6c51c378fe02204af9a76263e42caf4c5c0830e3765cb882a2
zfbbba5ee6dcdb008eb30be1c4218664615a5a044fb68b0b42e72062c93afe92a6d3206a9ac1920
z48438d495a3bfc896a634993ec1d264cd569304b3e0f60a7928184c3f0098c8cc4b84a70cc855b
zfaea11471481a9cc6bedbc99883fc406f235b53efaeda765ad2d267ac79bb483771f2bc2665694
zb6e55c20dad57caff68a50129a15759a5975b84fc4af656d387fcf7b2441b7a73ef2b504313902
zb32df636d357272f881b59671c7de8a8fc6e5bb5a87198908d312e137b14e0e61c07261e12a218
z5e28a49767d32c1e4276d4ed99b1b85172453633c9c7bae975eed939d206e80b93f9751760ba67
z407594aa5f4abd987b939b22df41c47051ce914dd23471db0aefd67c525f9d5c3f05534e3467b2
ze008b1ba34f3e311f49f8b4ba431f28235232865461c5c064247dd0974ba881cb411a45451a8e6
zbb3ebe1a67f7244680dc4bd9e0f0ca311243c50f78440b74dfe9c239ce00a6eee021369acb086a
z54fbf3a725426fa60a6c3536167c47a22c52c775d198963aade8d4dffff068a78011d2ce61aeb9
z88c630c2b7be41316c425438c7b7a91428267bba7868bc4dd1fb503101b96d6e5b6ec75b3e5c22
zfb1774bd5b19c29019d603151db80ca4b78e90d46be99629c83511a5095a7be7743ff279397cec
z6d8c3ff7ebeb9adde62495308c3d5d1eec5f9eb1374381d34184f857fc86ae15095a096111ae8c
z7554c007967aeea183018a3c0a794c130d37135eb133f1b6e0352d738d8b1dee90e4b1dd4aa59a
z437b34d692ec76e74f057ce62e7941617f2887922bf0526b1d9b5f92408e623cbd97a53d066b59
z00f435d6f9ae608a466c7a17692a3f1a4e794d1e446c112372d2072e7b1ed006dd99033da8f93f
ze45454cdb856340f3db6ca1adef1e95255438956a95a260d64c685a90c94b5843543954d98dd9c
z0bffa2cdc8e1fac74c864ce1838bbb4189497c342d6825024c49be03c2f95830e8b5220fc383cc
z1b314f97d45edb5f965be689c9e9fc9e92438320d7b39c15ae0b9e46159585b307fe8fac0a4924
zf2d002601f762939e083998f797d0691058e5a00348998b9c09635b83b4792d6a9f5daa97a9301
zbd2e439293acf98046b6a5a90ffe4b581827cb797d943f5bd5930ecc230886e1108bbb86825058
za4b7155d0e9dbf82318a31ff0d0520da9e5409edc297e7055fe0507520fd03fc5b5d6bff2fa438
zbfeb921dbcedbb90a566456a358ffe0f31e159954685a979492412504ba9ac25b7da78dca44ab5
z92c4d0cab202fb355a05491dd2a72816a4e238eb5893a0898034792922e1279d659a32b7443de3
ze8698693cea9ad05d462129e0b8d779583633141404921a064753477fe67c193cef669df9c209d
z27d3e57f7a5d1963e87856ccc0ae21025e476d26759751854124457d3bbffac3012c6f3b5781d9
z71f907840b2271852010f8707a217bf5df5e5edb9668645205a7ca7e123fa1e0f6218fd0ce5f44
z8356a11bfa05c93df1bde32abaecb6d0803155fca19f8121e24adfc8e41f4be96f81379dc80437
z5c88f8123d99f872c0e7aaf9aa898f3b164d1a3a0fd6b5e3dd7e016647639a6d2b6797d9229b7b
z108c2c217b2a25e1beed74800b53365da47736120bd825d018b2a551638b60f7195d5603fd385b
z084a0cf02f990b399276eb87b2d3ceb0068a518052622a0b7d62352a06ba0de296130c02ca982a
zcc0621d7786ed41a580993ba2ed033389ff6447adb1cd47395caf2f7ae1019b32d5388f0c168ec
z59425e5568de3a942876979021c66e4d82220ddab60a65ac0d3f46d981c61c46b29cc29a7baddc
z87a5251239406097181f46181840679b629c8449e40756164e42e9735c2980db13fd5b35e5f02d
z89d4874a7f677cab3c516940e569ec247a41009ada940b07953893065381ab3e2ec2b9b4d51098
z556c0cae841520fc6f29e18caf902895fa6323cbf7d059d6b246f73fda8b4996ad0038e4abf347
z1529f74477335fe119d7d3ca3bf428096b9384c8ccea0afa533cc096892d474c0f4b6c5bf598be
zeb85803adca5a9f5e7afc35972aec1db864a09df9c79077abd9d779b6536301e97a766d2221e1f
zd568e11a6f232587b1d43705e56d23329fa600535338421fc0992399c0b9b52c718c55928052fe
zbd3cdfb2294c70301be6ae1d845e442037d8856cd70faf3720952905f80ed9d3fee8209ac7b901
z070df15456b7edc0dfa2d19dbaca5b9d9e9497f39c41df46636eae145088a1f38d8f9d96eba9b4
z64449594f72f6e56a48c6e1bce5fa374d5f5d638a1357e13540abeb8bdae7fa52afd61a66621fa
z819c144b3b9e594cfaf7fec16e4a8160929f6068209590c4e8365c3121eebe51c45c646690621d
z36f3f541cf2ccbd4f013d47563796ca9bc95ef49c3f8b6f44cef84cb2b442212c0b2f5995ef49d
z9ab501a2b1236b658d04389e89710c8053970d732b94a77aa3428876fd8c893628a9e20a106648
z2e6567e9a9590524114f939a5bc0d46436560421ba34547ad31adc3624e553a3e430ee91297f75
zc38b6cb5fb72150d34753dc3aac355434aa58ad9041ba7a4c14c5f9e653d225184ab29df66268a
z4b9bc0a2669ea47c1d4d2a95e1daf4147c634a5daa95240b71041336b92f24900430bab9febbbd
z4a5f8bbf0c169ba244fe697d1e90470c84a7d0912644d9d7331cd48fb7114a3dd6c29aace1547d
z1246aa11d0bed4ea570697c1289b352884f93098b835da0c7f2918e589406c9e8d887bad60dd98
zf6080cfd25f859ebbeba4a930c8f10720bfe086fffc49ab4e2984e587518d6b7dbaf704a03bce0
z0e81a60d8c69346acc3b8864ac518dd8e921ecdb8e616e464fb6fa3190851261f29369ce1cdfae
z65f0692f6d2144f7191eeecbcd2795816e45fb5aa26e8b93f00233ea6006a27b56256ab39a406b
z356529bb0bcae6f0fdb895b6e95814512960f7af804e7b7b9cb2954b4c9d341e9eb1a8843b2d66
z76360fce4be297b45f82de57462447a2a5c712c28aa91ed72d94bd0c42887aca593f476eaca77f
z69efe2c24872765285bcf90edf8c1b71adad9bb06cc2220215fb5750adf50c65527926ed0237ff
z22c4d5999392a84b57186a00ca497ad6b95cbde4698ed1cce9680d0b60064763c83fa2db4fd52a
z732b2fa03c325092bac8f1e79f930ffc1d0acb59df0d78a7cdc0a03e5ad7de549e89cc4105f045
z63cc740c82ee22a07ab9e02978177db8e4e387cbe0f21803b87b9f8cc9b4c847ee806dd02a73f0
z035c76b23f4775974a60170a95e4ca1b1fba1c09eb64a5365fb9064a09f156f8f3f4421d80cd79
z32fb58775ae3b2973046621268c4b0635edda1465865aee12150573dc8c459f09c92a3ff0adcef
z8deaae4074c22ce95f044e6da6af1b22871a381707314588485b8526cd9a64bdf868de3b04b5a5
z48addf4c1eb1553bb25c9389c53db642b4cea32f7c0b5cce74babd60c2b6a5dfcd550bc461dbda
z239032dc9f752b1ee4c313764a45294614a8beb6463c055d103c84128410665c54122388819e34
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_multi_clock_multi_port_memory_access_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
