`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d5e386fdf9e2cb5152bcb6b17c5fb032793805dc36
z41bd7a6cc88c8e240d783536ae1f0c2d072a13001b8ed35ccb84142e6e072d1c8ecdf706602740
z9db7223e7b53816e42288b2dc42ebdda5736fe3e56f6430b4a1b48da20371c9e8d72fd29914c01
z8dce83b0ef7e6e171103acd22718a16c352a360a9a5fb4d383eac0f52511d326e1c3b9b11c8af7
zaee1dff85edcb97aa30530187dcfbe19c53a703b4e460d9fad9d74084da94f8968b8b917607b8b
zfdb8967b27883525e62faaa7ee4b828d2fd6b581ab98306d834537e006a532a80923c9b2fa3e5c
z8f91bbeab251133ec5823b022cc5ef38f4fc027091e74c588ad52c353852f78676a4e2a6a5e03d
z275549ffbee8f9c9f110c540ded54955354064238b9a7e47c312de23bc70efdfa66a0728d37807
z16bece208d6c1f2aceb79e1a2493f9362a51207002ba17369abb62bbf8ed2be560691ee182e38a
z7e067e0d8cd2f232a85c2f910f6f50e76a00a3d028c2d60409946d7f4553d335c025e73acac890
za49a6575d4908070f481c95d38c6fa123c5dfa0ec0a69b6fbf4acb054871948967f0cfde620cbd
z4d470ce4b917ab376ca22ada73e0e920ccb8e1809f349a1f1f2f6857c899eae927767d1188f3b5
z8feffe43f920b3ce126a943b7959c52c9b635ea56aa9cfb0b4e41dda62262dee305dc0b7e7ae99
zaef1b114da580012d25f1d7028b38af9e8fe7d5f89646c4f8f3b8009a1045ff4ad78223a284bf8
z5d685252c66c4cc9ce2a631abdee7df3fc165ff9166ed87b00b409e73d26d2655a0efddf7fcae7
z734619b01852999002d6910b76520fe46d8ba12617e6aa73ba93fc7b9485f41346c7104c7574c8
za6f09f19ccb0071d282a1c3690e3d6a194911e2eb14b5ba715e71c31d05ccd8545a4945929b078
za9476d94aac9566f8caffff83009796100c365d5c1829fec8ebf4a3be398396f644cc61b91b0ed
z10480e1d8edb0d3ca49240d17b57cdb76634f540805d884fa55659379049c1cc63618db3a4db55
z503104e7e157a83df728a43d6b33c57818a21eb721e9def2cd6960888345bdd9d3832c752f8534
za22d32b0cd7680445f0d13ecba2f4f0a3a7a6848930bdcd78677a411d1025e4200283ccddcbdca
za2d2a5c42b708a537734a73917f3b9e64876d4522b5bcb978bb60337b0ad7ba11a294d27ac5aea
z8d13cff999432f199e237fb1bcb1a94130ff243da59515f89a75b54b8f7293ee7714995f623113
z6619f5d581f9ae27415a24ee0d2c9af2548e11fdb569ae8a41c6c55c24b36763a9bd78c18e9b69
z221b5a5bacbc86e743771a0fd9a3418d5b0e5846f522c07dff3121ef58cbe16c755dfda08ee9bd
z29f1a86bd54bddf9a9304e9d8687d257405742a0616f42c1f53ad0ec5366115cdf632c96dae36a
z50e0f82654d19098c919e0fa547973b9fac58008d0fd156bb3388b59e4066ce9fceda2ad024fe8
z6120cd3ace0d36da99286e28badaac49f6055e97bc1e6865f6e9d4e57a7df9672b82ad84235676
zae4de79eefaaa68b6cc25ee8cbe08fe620e90938ac15ed8d8a8c898cf2c4f728ddfdd9232c1567
z3e7d8b65876e049e3a6a88e0c97553a7bf0c3da697af81d876e691119ade2611b2c773514567d4
z0e5435c6aff4f20cea143fb42b9bd108a3fafe7b1fad3350823fd1a2ea4a9cb64e13e655b46e05
zb38dc716467fa3ee62a203093c49ac9067c705c3adfbd60725e6579a486588d6b2118fbef8f534
z6aa408b8c46a70e230a61bd988e905e281778f7b68eb877df048d7067166ac231e26b5694751cf
z40f3891578a55eb70a6d8fb410686a475e94f898db8c36e060b73041c567fd1f865b175f41cb09
z7676ae25b987dcdaadd9479312e06b57046f201a47cb0b002c4ad7cedecd5bde73d6188747b562
z93420185b031ef6c531af5164df5d5dd0bc132e127e1302127aa6d8e98e287f62d4b2f99d22f57
z8d2c7b19d5f6dd510821249b7d812cec4eadd1200c26e8e77ce796cbea93e98e067ca1c45f0024
z7a927f62a2a9777ecb57dbf4ff1ebfda7cd0762f7a9fe116f74c8a54ce9966899dd6984be81f6c
z771a73a77cbdeaa3515ad2ca9f698753ee783a3e2c9ca47360a4cc461b1ff1ad7826404b16adab
z2b8c51e8a509aba3e52f4790eaf090cf696daf104b7458674857202462ad9efc0c82f442a0e42b
z33a534798e96eae8599f0ec07bb1525e5cbc32a03d5227322f2fd15e7cb37ce8776fa74082aa5a
zf2e903f8f0fa1cf8de002f7d3882d11b3bef745832f58c7ddef29d7113492a70da136037938ed8
za6723358e2e0dca476690b9516004100577fb7ecd8f985e6fa22fb2526fb7fb06b9c51320e66a8
zbbaf0dbdda9dc56283c72b12f850898a9751bb0100d8bdb690c8392c16a957bcd6b0b3867635c8
z733dbc7c59ac060bca5e85f2a3d39365056ea121ed4fc910c3dc828892c1f6b0dae981171b0630
z8e50b1e4644bed0502d022f115083781ec6f91483d2cabb7d6809f596a2db2060b2b19a65b14c1
zd33531628e28ac4c8d4cb3ebb64ae6a6971c63131ab16b3268a93f937a943037b81dd0aaa0dc27
z051f7351f6e7268c707ddc29920c09c825d3920c63c74465cdb28a78e24b3ca6b63aac2d4df603
z90d07a68b116c9999113d1d48796d2bd8e1ab2ce69c7097f542b46de701c8df0ca5b49d72fdfd2
z16e9d9de46f919bbd352fcf0a51357bacabc0c1f9f98ac9c90d46870698295064180398d1a7ff7
za93730787dd38d6552899f6cf017786640a9eb1750f36141788740ae4bd5e9ee72b1f304c736ab
z0071863632c7b957ff2a2f32f74476a9d99d7ef8b12c70d0da10312f3bd193e2ff4ddd10169a95
ze419be14b7bcd694fe6c3b2a84585a4b166a63846c57f74879b8962b569944656bee4ee45e9273
z0872e0e961394c7879cefaa0a0f95ca3d33fbd151a96b6a8efa6fc511f24292364ffc9a6d004fe
zeaed286060a77305b1a041ed293a08a915205626e3d0852e2eaea4df7c7fed954012b41810df76
zcaacdf3643cff6e2f2d266c6334b200db16de7fae81f6f8afcab858de0abe4bdfbbb00c14e9aba
z4f081487c5477d2e33ab586ba7723955775ad393d788527d4ed88a4d6f36b12a4cbdb8d6913471
z10943245efc6517aeae4b25f20cea45f43adc4fb484467d94f4fc90e0c98c853fc6f4fd8c9610a
z076e2deae5e65a1a65fd7ae874da62298b9c72c3abc5ff8437cd42d9762808576d238dc4dea804
za925566811ad23d8bd87f132411e72eb2038809e588261652f4e737fef4a3f8329a53f4426246a
z10aef1bf8a5eff55062572702d22715a2dc1dedbc8372f263dc94e4341391deb7af196e6f24220
z2b9dd69a35375a600c346becd3df830c58ab8a3fd30bb839e9f150a8c89095e7e1efa3625b1e41
z29e1756e7a1bac20fe56b3ef84b7c6e9b2de2cf98d9ae832ff06f3fefca4c97994a9686ec9e020
zc2e98d64141c356a044b61fffa1d48905c0fe832b656a82018a0c19798e9daaaec0987f08a1127
zc9ca5491f08c442a03241044b9b4e6547a887992af1baecd15dd07beb5bd7a7fb6561f3ed2e4dd
z0d1b6d7f910a07d9c91a7923f3776587999fc0df665ab74c65db0aebdad6b3d163b4a6f0425248
z7f2e58902f30f4ace9c3bed33e52e2c18939b1ebf1eaccfaa260c0e2ca38546229916d0d4534be
z92fa94b1837b5bf9ed86a0cc71a134adc16b7246f241005c351fd6c140e356ac9580a9c50f8ce4
z593e8501d0e8592fca6cb4d5153764ed1bcbd484bc9d33ab888e17a5584c6073b6f8a6d86b10b0
z703adfb255db9e4a01fedcb43c0d750abc284126ed59b9b9ace0bb692f802debd618af02dae978
z0ca2352d1de37d327499dd59cb7d2be7d3bcbb183991637f351c722483f3024dec6915961dd96c
zbbb305c950e23eef0cba2f5d25d66199bbad89e0cad89613f630753815f40363e0f5e5a36a2af7
zd0965cbb4367324520eb8224c01c4ebf49e4e2bfdbb0c2831f1c6d021c772ee8050c1bec408449
z819ea2c3f8031c80010e5c41d25b53b0663575add9b8549a973a702eebd15abb4e22bd3a44abfe
z87d63259910f509ae6b95514e87aad05c02f0df9dfa868715292447d3300cc967cce2c09b33612
z721f19d81d5c2e74dc2ff03fc1d7b49a88141248706ca70d74736586aac9bd0398e18d1e90845c
zfa12f200eef4d03f9576f3a512ca901746affe3043df3e88c449036b23fcbc03f0f34daff1ad1f
z9814c1e3305664eaa8770715f37692cce3155c34540c5b967687db630e97a3f1bcb3719b9cc290
z950beb8b79d2552876a0ac1ca6a5420d88ac8c7c18f60d9285ccfa19a2fd75db8c134a9115d63f
zb4522716bf1b844c73f0e10efb29e1b54f02b6593833c1d4968d457299b7f2c00b64fe2d3d574d
zbaabb818366a27ccc787e43786c85aba4bf9518fdbe322b89f44691d5333def6750f99dea4f25b
z291a465df38d72aef2a6e99e6e7da18b383ba3b80aaac9bb50ba970ba7137438134e4f67b3992a
z46e0d13efc1bc71a73ecbccb21c280d97e60a9ef82450d59d967e29548bf019f5a4d35c256e4d4
z61f43006802fea1857b78ae3a6e4df10bafba7627ea748aa121567a08cd3d54a4ed7b0fa17f10b
z49ff78380d8bb0e41d5c6326897adc72d268b0cf3dd7881c4faa0447986003bbd0be933fb946e9
z042a0120a53ed3520864116acc0948baf0ec6235565a11e063bf525a5c240e3352bb55980df5b2
z9fa4caf94c8f18845d8ba4eb2f3e562a67a179b9eef88519c97508be98650eef82a8dab8226522
z7b5da13fcd9e45e99c08675b854ff2cd8797362970aa71b79306eb2e9719310d74d6fd1804df39
z4376d8b3fe94a1a106bdb9915e20b0926c67225061080d61b6a2140889f53b4eecc5cd51725f6d
z88b472d344812fbc59889ce71a444a289d95283c682080c8bd51911c57e6d89fcd6ffa9f5e86ce
z5d1cf2efa1d6650ad10e705ae98c91c9ff3cf089ca6fd890d5a0c97e68ca591ecae1c7d567c806
zf915ada8125a675b0d48a3adc29328f475c579879c084ca06d9254bb72023ff42a1fa0780078ca
za61dcd90b035dde4bf57114c19f90d5f21adea4ae44c3348ca73fb10e9c109aba729a716365efb
za4b07320bd82485ef2ad1296ddf066001b6feed39260d5af0ba40df4643e454df6a94f07a5f949
z213589f332a0fec1a41dc7c79755586880cbd47d6ad01e916bc867408c940bd501b1bd61f83957
z8cba0de850b65ded73110e783165faa650895d848f6a4d228e498799484d2256c70ad26ae8476f
z9589783608a9ed633e110a66d5444cf339b9fb6b265f2e003c112a39c957c203fd3bda618bb35e
z5b9d835ffe818fdfb7ea94d428a1c582b14beb85cf9a1d2d97a967487b0f13ca9d6a84869feedc
ze8c821947291bd086c2569e4b443e76737223e5b66aa31f3aa96369295f1fb0ef93a0e0a1f3669
z62e660704fe9e0f3588d921beccf216d3ddf698f13ab66550447564023e8010c4a47df6074a643
zb9f91ceb3dc00b47e401ee92e6166ef44960a59d7279ae8ee12405f2ee5ad38bcdb26025086580
z8289253aa49c64891d16fa6d060a7177cd1965597fd4eb4cfb288e1d8496b7c050a1fb1a486d41
z08049441439ce4bb9b6ef193b294a45e014ae87bbb67eaab8ed0461ba1812b9df2c1177f5bdea8
z6f7a046749215dc12b1b9d546864ab24c4f666f9a9221693fab479a0295521df3d589c3832f115
zd72846859fd7e488d952d6320d22168f657d7559df930ef2554c3fcc5882b9cf461561c1f5822e
z406857de55d75585d04afcf441c80b5b83cebd06a1f8c3d3c303fc11c57267ee7af3f42e6cb27f
z5f101c9559b49ef86ffc4a2dcbf8e24de166ef41d2a5b56beb126c4adbd22d44dfb5fa38b3f0da
za8ced3b939e3d3c02ba8e10750af3e297d2c04d5a41b89660e89b8613abcd7e596bc82692be5f4
zbcf6a07bf7a9005c6cc63d500f3446ea7a786b90687d251d12be89b7f3be76a8e9abd790b5b3fa
z592d88207125e42c003ad163244825082a0954b4950f3497e40d5e8f20cf21a57a66a06590457d
za773fc6f4478d0f6f234abb13c008e77c5762a830c03ae577e6daf84ea2f2e838efad86ef24120
z06d1bef5d2259c9dcb49a035ed3f5bcd3d83b7b1da5a1a2c4d72f11d61475ce25182193f6c7e2d
z1dae753e3b4b94ad888c04ee8b534a0f080a52ff59f34c20886d1a8d86da2b8dc1db55e3089d00
z123075c5d7a0a7595cfca602b6d488f08bb280c0b99fccc23589df488c048da044ed397c2ba45c
zc2f2096f50a37b255b7506519910178164e6bc494ce7b8bbfec96709c8f8235f042967f1458839
zd193f15fa7e1cda8bda1a5b93a3ff1adfad0ec61b29c43789a88f24fd606a478916f794db62da1
z25934b5f392b84edbc3aa7bda0676af10e11ae1164e6aa2a5eb2b54091e139a0c54269a3132987
zb0b3019ee9c2ae4a8ac8bed4c70b38be0fcb12c1f33ffbc49a8921f963ec22ded3cf9cd05594bc
z924ea35046337daab8a2a4f78d10c21f7df3c54485944de8f77911f663db972ca18c6df22d9b1f
z6990fd35c1262a13a6ab6e69ac4262c8613106c3ee7f4170b9f1ba2974ef33705ab9f88e674a63
z75cf35eaff15c421485f3d4da9190ba1f94c5420ed5c91d398461857ffa94105fd718eecfa850c
za4ae65561254bfd1d9be0f1723a454eb3145831a5239c11cb2790f87a528a02b786d068a231588
zbf6909028dd490a38e6eb4ccf9e6f2c9c4bfab18d3648c09c222a57c5cc0537bf0ab3589f34a8a
z482a6a9283d52fe749cb6e82ce18d69cdcf7c32503c04fb217f387de4246f1bcd2286e380b7c54
z7cb6257bc751bb7ef7fb3f5015e784d3193f268ebfebd597db55dc0690e1ed40fa7eb41b9d8d81
zc279aed8a63324ca4b7c86beff976a554ed022f24342881e4eba7a8787bbd11b24fd387c986f7d
z43c34d6caf39986cf58e1ab249b48043ddcfd1235a1b3dc8b2a60bb493d0100cab7c71d8181574
z6109b5843acccec290c2fa7bd2955e2a046127c458f3850098822a4d87ccd5f855b4251282ee59
z24a3994caec7222921edd0334290844242f002e9e17b1342cb8f139be9f36d7db010b473450811
zb111c4b36fec6e18b465a3a0baaa6a7f4aed963ad41b53fb4f5b4a610962062e08a4178b126ac1
zb97ba4cf27cd4ae183555a528c784a97fa56e752b7ed5d715c42f2a3c565929767b4361f436922
z8f7c26d8f517099ee49dc4674c3dbae143e7ea5da872381d53fe439c61fccd1450534c7bc6ead5
z8fa22172b9ed3e5df4f1b8ed539d06ddedf21a1285cb756cf07164a68c3518c9c29decd0da1137
zfbb433c3b7c375ad0f9d4412fc6f6691f5ff3ef1644a27b13ffedb314c8da8155e91c3c63f03c0
za00700b7e7a5ff74b39737a6f70722c7d7eab6bbdeded2dddf5b39012e37b11b90356a7af904b5
z95327736d03383be85be918dad7392b6c51e9a6f4991af4ee08c07502a6a7160779ad5fc2f12b4
z6678ab269ec66067781ad99c9d77e11ab773e1784c894f5e18ab839f3d8d39d396396f51604dee
z59660a0b424506088a32cd1dec2385c3a084aae6a2762c92a9bd439a2d8f97cd2408832113409b
ze92ca476419c973ad985a2510ae3d0d7411a585fe13fa88dc78141c15a8f05ea0bb8031e5205f2
zb3b222dd7099be7149ada1c652fe1ff8ba04d6255ef9701722c83cf738b3cdc2feb4da64f0ac46
z53552118387e72e7a6cde4501ed7bf4e1ddf6971c79d282087d1b09235f7acc3e7378d6fcd74d7
zd8cd426ffad646f2c97bb45d6f1b95d7d87988cee544eb02496c01e05e5910fa50e133ba7a0c12
zc19e54352695382282f2d8b1b18aa2b019e9f88c447b6f5ab233ea89d0f80739ebfd9bc4be9fb7
z2dc0a4477e2e5397637a49c775fa2212e248f635d125993ce86d47faccd71eb06de680809c8845
zf27a12c4c6e1e66865fabc301f546e78da1054edf9fbba06cbef0129e16af5095b2fa32e7d09dc
z192d17eac2d5106e3e531b4ec498f6bd379291744dc07354657a88c80a551f72857d28ba6c4453
z8c21a04c9723d383f83e0c3fd9e6228183fd494584f4bb816d791a0c7a831f3795f54a861e7592
zdd840519e71fbed0f702e565ee9a149de7d73253270284aeae09f17a8e054a926fd22577cf9725
z354ad325bd85e521213ab485130723562bf7f425c4f3a00a37aae47649d1701f3ffe97b92eabca
zcfad8f891b29a2905507304944a27ab0695df1e4cccf8f806934fd23ed7e205e25fd4d8c8ddfa9
z6621cbdd3a1e8b42a237ba39e77f87c354e6c789210564c1aacdd701b7cf9a744aad9412155278
za9b9d14001cc81bcf3bf7bf93e77899e40e76c75b22c78494e20c4fa673d08cef1d4ae2ca08119
zc5de035efecf9d3be5cb9c0e4df85ba84e1bc38b316c4f0f397090abe884de9d4201c866843a09
zb88b2c27a162a551dffbf8ca06457148d87d56334110449c42d2ff0320e58781854a866e0cab28
z6d4355a3eeb455533f9233b31c7f41e7982410ff38f09a918085883a29c1ba720260cbbcd8cb27
z367522557079c4934b67a95bf784935976feb0f3cadacd2762c808efef969b11605eac1a385181
ze9fd4fd5b56d22677c41675af71e394b511c8bc15d94c21aff56f54d500331135531853c311011
zec22eac2a6a415ab5247d9b71ae4bc3e0899a0a5fab3173ebbe52b092ef74dd919dd1d7bea6967
za346a32cd59f28b48b8901aa3bc4d9ded4cf63f9f4a9f5b1ea8ea0f56657772c9ca32fc29c8cef
z58d156cd286b1a730309263b4d70b58d02ff73822e5f8ba88c33a27fef6b777a82545f0fc54374
z857034545206f9cb6d85c54608630dc69a0feef37e863871a5d60ba32938c7de19ac988bc7954d
z50580b1bb247a42c197fac75d47a1b6b06bdb3b39105973b287122dfe717414f663560ae1e698c
z8422a976cbf73aa98a1250906b083d1b4b0ed5fbeb7b3b25fa867f13e59c0be24bb10bf0955279
zbe771f7ab09bfba47a3649b4bdacce9135b788e3edaf2b0b19593d38457985a463fed9765f44ff
zca2c107026b591338faafda06b566dfb368a06aa57366b460b53969c23930654f26b8b42b4dbad
z81253f7ff4526669239969c9b3ac8e563768714c67188100d5718d556b33acd39792b1f6e888f7
z67fad89ddd0cc5a8782597e82032db3988b49e941dd3c216cddfb0ce58b898a2b2a3b913a908d4
zed07ec7ff8e26b39958d10a2929fdcf70fab21a4f0b6da1aa92cbca1072e076cdda1f6dcb6d1b2
z91e9eaddd1ce47da29087b9e8d47923e542f0f487ff3052d1e0b2cf5254e166149249e7b72c9b8
za05edc114a45a4b84e9878089eca6b48bc1a6000665284feefb93952925b4107a5b306236c5043
z388f1e65768f68f0078ab97cca64cc8cc11f914bd3ac27c4a2ec9ee0001ee80588301febf8c3e4
z07681f7ec95b40e346b69a5b871a9886a1ada84061c463362448c2d18c5845aa20468c225b2fe3
za3fae3d78e51f53bf3e057ab093cfb9df90065a437a36f8fa3de63a817b92804c5530a892f9429
z840bb846263635e013ae6ec40567f6a0710fbf0b09531f92ff925c3012ee311548d70864f90e80
z1795add299ab28f5d5d4804c7bd92ac830fb00582daca646807721c293882a317c59342ffb92b6
z9c8d6e8553b263bee0027405a46d1e2c139e6c52cc2c87b15b03c8aa7a4e851fdf75c3f3ace995
z07a65db0de528ce002973ceb776368d0ce1ed91109741121ffda89484f27b7219c0b2cc94b9a5b
zc38936944aa7033dd6cf6791ac828822635a4448e8e29a9c8947812057cb0ce39429a44407c030
z99bb9074b8faa093888508419778aebd51b932dd6e727fd8b2322461b4b2c8732fdc73e598eafc
zbea50581810ef868f0e0acc487d5520868dcd2f759bddbde94587eed8b2a10f1a642fe23c52f33
z3e171e3bf9539d455f4d33073244d6daea6a77e7f4ceae07ff4f0f59cc5b681ddcf35ae8658889
z68272aaf36e270e244d04ae1d2a3badba958be1ce2c357f062b79cc9cc67dae3b3b31b3e533749
z120d86d05eed15f8ddc0bb8741c1c66ba6cd95c2754ea7695c7d3a57a7eece2f9ccbacba861711
zd353fba43d2a66e75054f7d34537e75a87c42cfd21e4181d54cab5e8529c54889ad77ef2687c75
zff7664f250ce1571a0e43f7ab73ff7096ce234827a4340311dac3dc65ffb749eb2b2d5ed705d83
z2896659e21b6b1b41a5f05cf8e05a7ca055344145cb8d5566767459cf9b21f209435e59cdc0070
z9bc5900b3e96777627dd265be15f67d6b2ea006bbd78d6bca1986b1fb4476318268a97259c6c97
zd55b0129eb2a8d2cada99fabf13a8fbbba76c31b8c898c6c3156d246cdbe2faf968003ef2e9e67
ze218d1a706ba02db9fe9987965748b62e7552740b191a737a92642b8bd3c541c8bb38f9508d9d2
z98738ce0c563c1dc4b7433c01f343f6fdd4bbb9d1866d6fbf056babe9d29c1c301d8150cc49b11
z9218be2bf55439439ef3f0c00a27ddfb3ef9c3723b7e07233e542f27c280432203ca3de38232e1
zabbd5cfc7afdb158b63d39bc5a60c63c0b44e62460514b9b0724a1bf9e004d41ce9feb69068b17
z4d56c6160f39ba6a2602b17bc693673d6d01a27c13e46b55855f8dee9a6fe7ce496c9bc813f7ba
z98c454d4ae63bb24a4b0f1029eae53d56762825269b4c5f8095ca22e7d5da38658bfebe40c8ab5
z81b8a9da40fcc0b6a7e8003c40bafa73bb2c0cbf1bdf5931593c42d4c49305673fbd7f8b9bb847
z795c42fa4e791a47f8f999e9f036dafd9e300f2329ec2d307d25e711a37c4f0a5a0ca2bc21e414
z0321ba6e056947771a798e48be6515e744357bdf2eb355566889ad093204b048bba7725d36aca8
z8643516a26c936e47ca17b18641b8e8744718bf46ca1d3f09dc1c4ee3222e380459e2674879e5c
z401d69154a38f95a417506dd24d5ec71270c6fa5a4b981924cf130514573ac5b1a01e67823302c
z177e6bcb95bca6c55835f65a3cff01eb448895b69cd418f25818d0f47b47a0af547bff0d77e496
z6c0b24b6ba93abd7fdd75d480b0786d7686dbf4e5977ff409cf63064c606bc67ff50cb3ba00907
z79a793109a71995de15d2bd93dcdf531ce90b84ba93222af0f69efab6b3f766b9e8006b5369263
z97cf8cb6d37200e1f1f483edfc3e83965a830c90f773974a87e1a34252455fe748de036409434c
ze00899a0a1342f4247e6c44e7b89dc393593982fed0befcb5649f8be4f24c7f6259d3d02eb3748
z9033b859549d4baa678b348c6d54580b02506bdde02caa41696c71eeb2048e59c61479f86aafb8
z237a455c81057da552da3e6f301f553f1ccec83546c20b4c95e5b9904052ef0a5729c5dc25fab0
z197b97fb03b9c62fc04805a766327abd0486a3aea8571d1f9fd5d8d083feb4fb4ae03a7e53fda5
z0a339d5db04f79919faa8cbd33f291dde05cb07918949a30ad2d311003f3551bae14ce80324758
zf6624dfe08e14ba744f8db4ae6bd5b07441255463b77dd8e24d70a066f09a61a314c1f8f16485a
z2b2b1985b7d1ef5c40de6fc6942956f197c66ed5cbfc9dfaa269d91da6236a1da155090a11337e
z5207c6bb66f432835e88d03f38d7f9e8f006dfaae8acde937356114a25f7245081505aa1a016b0
za5635e7857c4af655eac2338da6c80bda67b55a4cdc83cafb12d008a6f3382617fa761c98b2b10
zd8549d32466eea3bfabccb1f0b5eaae2fd8cf9418bfdfc91165d7cdd61c2957e076e459ae4a70f
z444f557edaef2646ac1c6779f7f5e11c1b903790682f269701e297150ed4c847821cb9efdfb161
z9be79ebc5e06921a526620b7334e10efb8da9616eb41b3a583b652b98dcc80135d72c55f823215
z18b0e641a42b4bf4fd4d56c2ebe786ae389a46b852a052b428b05ac306d8fe25e64e02ddf5ce15
z16f4a506065ef8c83a7985b689d3acd09825262f451a853debc97a82c05e864cf6839a6c5237d4
z9a1b8df306339506bd7615f88604515dde02f0446b7dd0bea34980f4ba90f9946d4ec7fe8bcd27
z82ecf6fe7a160eca1e3ca601bb10acdf2b3a5c0fbb5ef79de919daed8327e8d11529dd21061ac9
z1aef9a60610a6914b0f78d433f903c9b22523221c9434b7fa305228171f8c73886c2abaa6a105f
za63b8c5f94fcacb4c185c1dd67b629758e86ba083bb76795238306b244ce8a086b3cdf931161a4
z396c9647dd6534f9865ef7209164e7816cb1231b00bb4060a907292b25d3ee0d708a079243bb2f
zfbdde63b64e9e184e82c9313bf5bf6d3b233f2a980ea9a4bd5966be03d2434f4986a23585eb51c
zaecf9a04d36bd10d8f79b977910fd68dcedec6675d495c2d1fce0a2c46b759a21939096fd9bf72
z24c1c63ddb199a4c27b07c0aae4bf14f9b09f32dc2f2639909523baf1e12525b15988b44221462
z49b743592c919afe78bf5e4ad0f26bfd494841f698f4e3254c7d799f648bf86f288ba99578df02
z13cfc7670bfdbde062c0863b913f377fb7a757f9a777c1591ba8ea904bed73fb4ce5ba1c725f99
z8b646bc06777a49fc2c8a7d0937ff7ab7c231f5c839428792b39f5bc7ed33f161c9d91c6cfa9dd
z9c3fc9954af92146944427fe95f0c910c82bebfe3a7c44d77e3ea924100d220e2a0d35000dcc3a
z22a7efeb74ea1bf0761ce1c0c6a42d20553055cd6388b3000936119c0a54e6a48a430d69e9875d
zdf6aa34b71cdffe6cbed68852b75eb866929bff8d4cd93df0de575cca3b8887112faa3de8b764d
z00511623c7d6adc5d283568397394cc1140e7524fe838ec14d5e47bc5678da270d6491cae2b332
zab45b31fc8925e4b4f2da00e4df85a200f7f695bad9489262ef7dbefae9616bc817466b6111ec0
z48421ebf45315d8a8ed070eeebfffa8953e2236d0524c69810f0259e87bfa7abc47d1db497aca6
z487ace9a85a3bf30f12e8ec4a123b34e8e0747edaf9d5ee32c5e3502b2431941a9dac8de0205d2
zbf561af56b14155cb5c79f7589c42614b91042909b97db71cbd30bc97e2e262be3472a5ae229a8
z06c4d0dc4a7407cb421662ddbad143d4dad0093693c9eab41006ba0bd89cd5b8513b961dcc0314
zf4098e8f45f7a260acfd9595dcf1111ae2ee04c2b9a0d858e5f0510134ede35b911f06968c3dcd
z876411582b355769d552a4cfac0a6f049d3eb025a6473f16ed091ffaf381843a05930a64f9c8b6
z810a497ebcaeecfc0f2a92704c37097abe75031e8fc3b28cdce3c3b680b2736704538a78ff8d2e
z027def7a279d46cdfe251dcf46616150b4bef79307764234e0c3cf847cc92853bb05a49b047964
zea65e003368f695854f239591c2d6311160a14e9e9a2be6b232b918caa073d2ed0116be5ddae1d
z95d6d602fefe21371236af1f98819a9b53efbbaaf25c4da68d4e03529dd8e1da00dfc2dff03d31
ze3fa430043ab7e45978ee786476a56209c48b9304923f198081287b32a4af8f56fe73280ca3639
z0caf1cdc43708581499243bab4b731ac7bbaefe82888ade9d0711056b3ed951a7ca537323b44b8
z09cc162aa07377b910f11bd5f43c824b564c8bb5a8a3abeaab884218c43f04b90bdd14ec46f09c
z0e03dfc85bd846e002a61da995cdadbcac623bee1e221e955c478a4dd2d8529bf301c2b21078c4
zc883f3a940a1dd815bd8f98398c2641c7dd841582f1eecc6bfd20e9328f8e49b7baaf3b3a665ea
z1b8aaa959bdcc32821f52cc073e0cced7ce67a22e62eb6fa183601a3d3176d92f9164eebc8c140
z4dcd9d05762a475de11bd39d47d02e133fa33f4aec7f27c04961ece906f7421ca8a7648d0ab485
z07f53ef99f543b8904a38ba9bb03c5d91e3c287d79a8ae7ffe51aeef8eb28c17f32581c38c0a88
zb1b17af400ea91ff54dfad32304a9d50ddd979be9de8ad714a1bb9741952494c9e858527813d2f
z1f8d89f5e06d3e44bddc38fbca9cc1e0d796df9f938312e82f95643b010eb892585b47e329135d
z36b9915df98ca44b5eb3e2372cefb23e51fdbbd115a08fde514557e0d4075c78f3916588a2e33b
z0075987e946c0ab408ea5272fe720cfdac5a8e0dbfe33fbf5ed1748459ee186855109c2d7d7409
z2707ab7f1d333e67a00bc0b644e31c2270e9274d7c08b840c2c04151c15a4a1b39873acd034ed6
z2fd6e86cba59a44f6e2087179c5edb22beed50559a4e16771724512da7ad3df61561b69df78b14
z7959d725005520f3b4f0d6655470584cb1a1aa2c5a47089d6b428f0310fdfd16b6d5dce58b6572
z4a34ec0ff7ec9e3d9fc2361dfcb09824654834b1573567271bfdf08b21a000eaaec9cb73b990f8
z96b22a4c156b48d67ff1a2b5d409ebca4f189db4aebd0ab8dff7f8f2630a3ede8ea4a59b72a639
ze87fa4be2c2711db1506fa9c8956529d496b11ad2d011ae6d5ad4d15833b8ceaeebf35bd117ace
z53c5ad91d963f53aca47ac364723e8227b16f828c168a2371be619e84d92bb087a492091932ff0
z92d9cc7839dce137168435c9bcc12a0c11257932329a21407ae6d73d3bc07c217e16ba4397f362
z2fb743800c8b65adb07422d7326065beae7d6856c9ad029c37cddb49a23074da9aa8249148b63b
z4fb7f7778f5c421467d71f6b112425649bb5e2f8a0cf559b36a50df4757774e158a251b29dc39f
zdf1cbf3094d9bf45e6ea342b8fd001229f9dfa0743f482252ddbd0a11a26096622c93893f5edd6
za96131f63297f692663540123c3e92a4f88637ecb2d9226e439e4faafd91d1e6a80a6c2167ba9c
z7695fc16269d972052ce277c8bb2749f38c384f35ae5456b7a246f875f3ebf97aeaf670cbc4338
z7bd700a49a6245fe2b60548102ac99fd47e5c9f9f6e05b7e4bd07947c86ec35a0e21e2a27938bc
zb725c20f9e258c936e3163e2f5c1a60f54bcf306860d596aefd62d4c601b10a2e5f0fe21a3aa5f
z5851ad8d29225a8e215618f0d39574c61cead7c43a49c580527458d793373c39c76d4d3874e3d2
z605e277a1ab3f6d485f39164803fb9a41a28e840a59043c9b8a25898b090381a8ab3fbabf7849a
zf9549ec1b099675cc811c04f2066aeff6336a3ddc07e5daae323520195f69d67cb604f8a47ed8a
z72b4cf04d2069eabd9c292eef638c0a4945e4c2410d710fa83b49709c2d7573320a0fed855de60
z1f48c1f0a4cdd8dbd2ecf27b6e32f09cc4f73e160fc47b5773dec9c56d01500747f693daa9ee7d
z1b0e3f5aaee841a2d1568cd22cecf87b840355e55d291d0eecc01cb91af42bce0478c6ef22db15
zc7f6980ba9bb71da43fa502696f7d7669a85499b113c6adf2e6ce8a1f04f9736344ce86587bd54
z67850568805727e8e0287d337d5cd7e0224c4df66915e785189b15286293070963c656e9171cab
z9777930c7b56e4f16b0d22b706bd51ddac2fbd6549a8e0ab18a51356387c7c8a3dd7a74aa3eb14
z7f6ea53fe5901ca6bc06a69cff427d4b3b7386dcc33a53662c366c98ccf2b5ba2adf1a966c43c3
z6ca44e239287a44aab926d1bea2dc1e67db602075d5501747b1b455f08b92fda9740a8117f5520
zf4e5a0b4cbe3d75184a98ddf710af87fb61ef699ee1fa881bf32bfc53633cef5bfa9c38457d1fd
zcfcaa5b1ed6bad9f069546fb486f70d7ad4a61b4059860e555aa317b6c126b36742eff0158b35c
z2b48008b38f3d8dd5f3cc617cf97eb0b892ec42df9e9dd813040b8e9c1d66c868c1d1f6a946e57
z3d3e2b82b1b7b5634f4834e9b68db798304d5f8783a740a6af7b9d74e755b26598a93a7235bf63
zebc934e63b079bfe0817c46e7feacf93a55dd27920f24461c2e05f111a5e43519c09a26d4ff13f
z665f2fd9f4209a1bd64761648edbf3826d348ae39c3d98fd22ea68de9e4da3b4353a53fb8d5ef9
zbfbcc5971a9c4ff44a2193f171f184f12907883925b5cbf27a5d9a7aeba93405c8be7f9323f9f8
z2cec6e928240f4da6f6f94254733e76ba7a6cbf8ed5e2e859f71d6e20f7b95630053cb11375352
z20535b4b21b4e013a0140cdbbd3d617ce630c01062bea26cac9202df0c91014aa77c015c28ebbf
z6406f9baf85c849b38c62d358fe995388ab0c0e7c4abd412bdf0dd71166a2642d04d679380f15c
z524f284cbbba69632bfc946c7605e39487640658d4710d74cf9a0016072dffd5485bcd41ef6662
zad41e7aa942d5b320a690ec1ff765ef580d92a4e984ac8d49907a16ccb83ce1d12feeaffe546b6
z3134081e0de8b27bde4483f9ce16087ba400ea62eb6a24799ebd8dec4d6d385236773c4e0de707
zeb5ab4188de129d86cd82f066b17d09c3aac98589e8d99065d3e6961d105761643911d209a7797
z10ba8771655161aceb1bc26a3b9d61a34ef1f77d1b98eeac73da9faaf8c26a929f0bdc8b0ec635
z22858745f8f17be995d62ad66c86c503f035171b031ece7822c843b6090562cf6a73a15be80d95
zb13e264bdbf8cc18c08b29832831f0d17479d61aaba5fca8972f804174392a73332211e68273ae
z92fd34706ab9310e025d27aec961fd067e03b1a9ad0816009b4af3b861e054a5d87ecfb6eb84b5
z6db4329742b26622e92e475ffacee0ed3a55c219f2236035e2c2e59fcf300efd707e8f4bb0ecc2
z8beb65910642f288a0a487cfe0f3a88003ad2d75f659608183b6ad73af61144a747106a3c14db0
z5ea3cf8e04e59dcea986b97e2dd6938a7e9fb77fc22231d1cbdc9e84c5be8e29176c5d88756678
z734dfc382da0e50b772d2060ad451a91193713bd9bfc62e71129cb2e41f5510d411248001f71b6
z424475dcca2be4e891559b0db09409806f65c5b0d917a8c06c6e8868192ea8aa9cf1a379dc87d3
zdc4e7593f4bff5d178826490d1db18c287536f5af1e43ce7966077b8058b6503815863038d1a52
zf97c81f0ddb7708c190acd9448895294e8757b6398ece5ae352958e0bb04977f7da55625c7352c
zdd8ba3fcc4de7b22f3d6fd733b690da760f062209e1832ba61f67aea588967619754727fb48278
z8e8b59fbf310c61329d26a0cc529dbd86d5c740c994969ca3d2f1236469ddc97d728796defc424
z09e3a3eed5ac7c334158210b69a775bf252f563f243a1d8ba7ba97e074e4c3cdfc47770f38667d
zae73f838b0f1fb00b7c9b9599f0ddf148d39681eed6ab246c63220e7b899175a3cda95d3818cc7
z34e56d808c314ee949f2748df0aa412e649b66fbd65ff1ae8915dcba48418f7efe5744d48477cf
z3f38066d1745b389dc0e1ff0e2f166054a6868d8e8e572cb5a1fd920e77452c1c4761d2c4bcd56
z2e6d0432f5a0a9030933c6350b72da0264756e839c77db4477c125e0e13d9e260c3572737a175f
za3e4858f9c838b8a8a15fe3b947c4a3cf6f7b538d50764ac29c31c2571ce115dd3010f1287f846
zc333d8f0d1c7a60c36ea59965ab100ffd67454eafe57823f08a982a99b57ba99bf91c7a213daf4
z050c98d2aa00ed91a8870c662fbe9abbd9e3196078ffe4a0899a3816c6e2b0edb4e1ec9d8aa069
z7bb5c3666e92715ce831df57441c220da6f427c89faf85cb8f1fcda3492fe47502fc0a3aadf421
zbbcf51c885c075cf49b8ff918b9bab5e457dbdca67f2f20345b35dd4385a5ce7657c9c833dbc0b
zba88fd756750046f9bf5f3edf5aba02f2708b2f4c4632aac86763db77a4ac6182b512e95e2c2b4
z7e0976774f8625f7c51016c5f05b589ea3bb15ae208bca15938df4a7ea3ceff3a46d79e836645b
zeac608035627265758f57ef868ad5a0fdc05367b691213d44416aa82a9142f7141a70cf16a431d
zffd91bcf5e08c0f6a8b78c8caf6c5fbf3051d1d12b47e3054f7eba7421fc37b270be50b92046cf
z0b6204e5e967169b1673b3f1893cd9de2f6d9b4a684c27ba01151a053f91a3da176de96d9caa28
z65af01a9d9e0591f38c1f2b0caf4bc065e779c6dce071e2c8d6a81e70023942154d6f4402cb36b
z7bf2d0023004039712746b937249f9826f800847937608300af573bf82c30e938acda6b058bc80
zac0c77037edceb52630c17c9f6c11ab2cdaccb45fc623159fd7a0f5f46b05bbfcfc6923854b32f
z067fdf8173b706d6213e627cc368f75b4980cbe0def11ed1efa1a8a8947563205cf7523e3c579e
z0b54d65b711e45c40f9ff564c1d113408af8afbeb64e1dc224ca5e9c6826e645460a6390577bfb
z49c779ae6e9e892e4ffa5a1db91d598b057d0303ac067ccb6fe704dccca92b46541e0b78b930ee
z58347d362f94513cab1694606c5ed06aec5551892c3916268d0857866d34a02e68325884774671
z78d0371276725f2c8c70e27096769af7a123e7a1770b826f561a9a5f6c13a3e5659c053a737652
z5496e06b1f1760c6f2d19d8618d02b09871e8abd4c9b65e7d9016c80de75c14b247dfc2fd636a0
zdbbc490e8e9fdd7453021828e4ab23ef57e7a17c762cfc7a86f5f6d1507b982f3b9695c5fad15c
z476400f6696c94ba4c6a7c50fdb7e17a3b2b8b7d9a8b761d05cb3eed69a8795365be152a47b382
z91f9a84cb459e10d0b5658741952b858a751ab6974cf132d038c332155f124c404043a6614acba
z0b0def736c729885d31be0dc492bec1744eb82f91d99e78280f838b4cef8b3706dbd3c9245f394
zde80399cca4f8a6b455bb0708c4c0a21228348a8be163adcd766c9d8ca89d5e6043570cd4929a0
z9b48fc4c34451e116a96db2650529edd1a4300d4cfd84574e35a75c46dbc6404f251bc3dd4869d
z407d6c47eed47052d64f2249ab67e746da500a1d64c962ea4a5cdc34fe0b5f637ab16fdbbfd131
zbbb3106b2c7a6ef7836d964cb7d44a045b4e9a6ea07d3c1fc1577634924adfcb546a266d515285
z7f11e0f7185f37d0d89282f5d0f6bb60b1b3782091b7129efb085a77728c15ab08c20a04e40647
z31cf54f092f203cb886de74ae94f0b8b3bdbeee7a4b2881407dd7a66f7d9c6acf5d228ef116c5f
zfb05689831ab3823955e0112963d8aba7e8d8118248a1897cf2876868231960485b874b715d40a
z216e74eb9cb180d649a4243b08d272b4e28b42b1a958c74f182729daa178a615eae46d9a94ee6c
z741eb7c3f35cdb7b923032f3d486ce2d1ecbc6d31bc4e4adac27feb39db10f46a867d4c62da6d9
z2a1fbdc5d701bb540fc23823eb2b4a875a653de6df9dd112544dfdc120b13d4ae1d5dedeeab59a
zfd73fb5a248f0d5a3aadd8c7a260c1a402e5ece7bc9b25b7a07509e4f5094a34c4764d92174343
z703a467dad3255f3df7842c88f1af43fd0864e89860964242ad9bf58f9739aee84dbb22b772863
z70d267bfa11bebd78a7eb1d506195492735a40d4203d30a325f01633607aa3465ca40e209601a4
za7f403527fa2475b216345e9f894e5bbfddf7d21f33283f4e2c4becf0565c75bf9c59f720ad7b9
z07f153f77d25188d5aaa0c050bbc3c2e99d062001060ea078908f5f360bcafcad6a88589ccfae4
z60a7fbd4400cb2d45eec7587760b859177bca6130754522c901b0a810f086d5d9b5dbf572b9495
z79d861420d25ffff8e0ea1f06c588303081a786c7d09490410953709e2cbd251ffa170262b0338
z6024257ca2678ec3e3123f264bc1c1a70feec705daf8b869c53e6ddca67e45329f435069c31542
z6343f31e8f73c4dffca5d486874b22def5f7b53e4c8a739f21d9c66a171456b23174f5ba4bce73
z076c5d8ab0f88948420abfb1c77192d9616fde23d6b40046ca5a6b96e974d03ff79da7b58b222e
z6037d2ee246d04d1d1274e9f0e740d3962ac6690ae61b20e338ebcb3e4bdf740db70dfabac31fd
z36bb1618b1ae236c2ab60d5332ecc2927a24b637a3757f8076a666a75cc793bb49b0a6314a0e93
z53f7aea45864f205bca9899c8dc2c9551f7c6712f772b1f678ef2a45dc9cff8cf4ae9499a6d481
zaecbd47ce53b6438064b0134065d522a00b2b327c6527e2adbc2e3f128c0d058f3a8ec6a4b790b
zb7e3153c3406d4bc8ce244d3495fcb8c01c669927a3be747166a2a0a4c937e4b7691785550f0d4
z98872d2105e320b74a30dc03c53263bcc8d47f28af167edda2130a8850b8bd7d8437d9153081a4
zdfe6ee080a89a4b7d0719a179b9cf9206e14cc955f862f3df4659b6d8651bb2b6d3d11a7f3f2f5
z8d2f959441e6b70f2a1375331d69be96bad8a813a2cc884aeaef3a388780ff14f279736d1a6861
z0c516b60d04130b677a081c384de2f728863881b35d742f89f08293871f9369600b72d70ae026b
zeea173e423708b63e766a1a378e509d8d682c0b1a3ce79f640f324f10ce5ee67c08ffc87dc7bf3
z5b9ced3ba6b3118483f2f6f66aa87ebfb125015adc3c222da9b847a6aecf1c45cb63ff30f80ad6
z8030e71d4d85e40720a74f503b8e476eb8fe809f2c028bab484f44b369949c5bbd0e23bcb6fa28
z5204dacff40195db3741d0e8609aac2cd309cc88a909537b6e648c5321037f5803ce986a98aaf2
z2c5e31bc1e5d8c40f82fcc12f99c6ea5a9c2ef9bd1a07c3ce61a88183a7b4e48b51275ad82047e
za1fd35f954ee7bf75b5f83ba3834c13f00242435e655a6aadea381a8d9b5ed714a0627ec06a432
z9ab8f6428fc1e4280066543a8c74f86dc5d4ae3e6e190b574dad469fe1f03e8aa0bdce51e6b965
z8cbe3b91465091a9e47e5509f460463d603b2785d2dd2f2abea00ed525a5b0260458cbb503c7df
z9b6169280804c6794cc11d339975384c5280222b47315223232161073fa9a94e8b8f412858c951
ze84f71a9b4759f30daa0976d476ee8dd0807f9932e731ffe83451117429f70b95ac18b4c5ae7f0
z113923871dd7335220ec422ffa5aa0e3e7ec93f0618be9b5b285f29b2ad20edf3946510a2c6e65
za5ffcc6d4072bd3e6c002da874393e76df2cc03ababe395e02e517054941711bd889117c207345
za817eb79da26bb3cc57b7d21d84940dd2471a5b53d266f04bfab3084c3ec1ab16eea20ee4cd3de
z2a352e6a72264835d1a49760ea5132f5d88a3b334ba15472aedcbbb7a03cb951c9a574d3263fa0
z2486a88249f80dbfd412f1ee5f33f2731f7355b115b63294e1358ea8d35354085750b9ac2c0cc1
z2af7e709fd688be19f7892f97295735b07dcafe05f4237445d49a489c5d2219a6411d3d4f13830
z4a968b32916f74dda7cb7b51e8022a1b08414fe2032557d68ca2e4ed33fa518f4214375465ee65
zdc41d7f48f4a56c47b88df74c8f4b80b43e3c93383faca90c248dda035d0ca46fb9623a940608a
z7ab7b89384f1593a0aaf8bb6b3387831fb1bde69ed6cbbeecbca6f134262af53127cea86607148
z51eabbea46cb4fdccbfca101101a5e8aa381fc52c9da4f071a656cfb09ee5437523d8b4bde031b
zb7eed961e9d9745351f29e0b8b759e4d017a432d0f80db98cebcb236073370e85643942e5edd86
z913b7ed94b872d26081eb3a6fe2095990d5e48d371080a52358e307e93e74e55d8f0542ff573f1
z07ebae9dd78e9a4111e3a3d3a6581db38382fa4070dc59345e87f0525d9d89c56c30dbd8c710cf
z7157cc278d2cbda438005da714ff6088824d66a14ca620d772b54ef8414e93b62a42ae0c99441e
zf89b656caf76473242e049b138286fffc8f811af8bb2fc5a8ff8e4010555ebbbd7da8201e83ec6
z981dd435524364261ae9490f590bc51ae5f2193be8abdf84b39fc88027c3622efbb796e3e36a8f
z4f772a62ece84c6e11e54a07fa55d8721f211b7a5cbe11969a615b4c7de1b0d991196ed81badfb
z3b5b8b8cbc1f1ae61fa990c00bd905a58de1829cfb8dd752c11dc2f7ca700d9f6c0c2339635245
zbeefd474d31c2759af2bc758426f5a75c798f37e617a1560f4cf73e494ac615d71174df148c695
z53017483089c9133e869924354dd510af10366c6ba241e2614ff6e0e5ca023d8362eff85ec4cba
z12758ffa194d34990ad73d94e8af65a269064d4b144c23a6142c1259e0cc57ff79b016bcd3f555
za8dcb3e21264288df00729cd980ab4995a4c782f7ec52fc8e803e64229806d4029355f08c4dbad
z03faa571d346bf1868648a49dbac3b9d8ccec501e7a83ce01a4be46a6e079f50d9c22f4eaff9f8
z279c3db3f4eb89e3f0c479485f30c1b63d54cfd6e8c1d1eb102cc8d8c858bc57552701a9d2a418
z34bd1a4af522718fb1b16366f6fd4dcf77d7f58bde30495160b0a953b5fd302756694dd087599d
z7b3157459568c85df9c65ee8f331114739ce889a884784deda17241bed204e9544f7101376e09c
z36f23c11db337cbcd2481ca35ed99b48857bdc2a9eb2cacba2274ab75b316ba86fd1761f32047f
z77f6e0e9453feb87057b9f9f37c315843c0f6ab8d0fd08f435605477a911d6e656993fbc4a1be7
zf4f4c8a11f56865e4ae5b184330fa1af92ec8bbad88cd7e50f8ae455584e52d9b86e6db3938c56
z37e8571a1ccf6a332a64fdca27af637bf65a4b80fa14c133e220ea11ae365aad867e051033747c
zc1c7fcfb951905bd8f12fcb40dd7fda9ef1310a1ab90e60665f3aff8a03c8598d379b6c496c763
z349ab6852f2a999c08dc3f8e2478350acd22399e7a7579506a27bda965ad9b93d2c68cd5b341f2
z61c6e7290d0aabdbffe09746bd7762ae81e9d417c9668d5a19e6ffadc628499e03e804ef7502db
ze3d9a7fea903d91b315699031a79ee1a78b4a1155b02aa757030fb9a1c5434a250979fd0793de2
z194c6b4caa713b86b002f951468408437f79227c31a6bd7b84d3ffd2196a17b6f407be50ff327e
zfebced55ca6315c45a459584e6b0f07cf6b055467df770b59bc07274279e665376c049af57e341
z5ae888bbfbfb59f86c7fdcf3f352bd6ed54c65fccbce7ec712528dfb3d749b004929689ee9295b
zaffc0e999ac5ee038fcef2fe5e608bd8dc4c7d4358c5f948f2147fc9eef27f2af536afa872416d
z6ef1ea2c50a46c0d08645fec6047229391f40d2b2887e8aeec429a9d187e208f8af66f4e0a0941
z77109a6398d2dc8f6ba66b4aec6c5ba28c93d37cbed9c483c3940dca57004850c0c25eef59d0cb
ze1ffc3d666faedef1265ed0d503e46fe36f649732e7797e7fc8288e79622a229ce737ee3b97fff
z3d808345f402371007a8537f17804a0d32f4724f1b0ec1bec0c298abee44bdc2335f90478f892c
z059963708a5ad4fd57c88a238fb5391ee69622eff41c05083a6fa2931337eca78601217657fddf
zd4521eebfc3bc69aeca1e2130dee3d2bf448b7e6c1e4aa802818053526dd9a009cd32f6cc429da
z7d69cd33e75a0ea559effac1b778e71768474994210163027872a58f60943e6e13e3d120db86ed
zf49d029eb6a180025795119f91072142c08477be9fb6520cb9d46cbe9d870f6d0b75edcb4c09ef
z2866aca6d67c7d91d5d0948359a8b4d13d60b609fba8a09d0f1b4c8257279ac8a06a25e2409e03
z0ecff08d19924d04287117dda82e456b77660150b44544704fc580f6ae88b389b724d8ad802c4d
zfac2174bb49a8ac36d7b376b28092d185ec81303b547694c59a41fd6314bad7bf24fb03a6a7dd3
z05b17a6f479d8369146da61a589d8e3ae7102c58cc9b1b4b380da67ab6bd93029eb7795340fd61
zc107e05c99078403a65952189a1bbad51887336f0c844ea5ecaeeae45d3ce2c7d463b07baa4879
z5cd51752ee5104db7ebbb8495a4a2d9ad00877a6d7db45b0bad5a5de4efd1251151b5e2696dcc6
zae332839b3bbd6f9b877b792b48e3c5faf481e00cabe71c17bd7afd3e136c55baca9634f7010a8
z1fa7df707239614400636a0be4a00d7a42cd4b21a19bf5773fe3f78019029748863a50007bf550
z8f1085d98df7e4f76baef3beb92f93f7b29a8a90fb7badc0129e286134b4c15e6b243c7006c18a
z32ecdaf31135bbb59b9776fb9815639f6f55bc0eb233b8cd4bdee066b4e6ef4faad361bfeaeff5
z07cae50307bad6b7ceef592a1e1d2e8dfd31fa039cf2b8f392ca60723b989520d4dec29fff387d
zc78788cd7ced2567743dd3938731ebb90c168b3672bebe4236df625458a36f1141796d2c2b27cb
z013b36856fa9d0e8a648864a9208fa10188b97397032090bd70388e29521c12c9bbaede65fbfc2
z2679583442032c03db5d498de976a9b4e1e093e8fc584c34753767d3872937cae85dfaf2db8bbc
zbf3242c0f32697f402347f0827f06d134eaf7bca8f6c3fd003f325f48fecf79d257a143f15cfca
zbbe65dea6e10c1af9058efcf98cf117f3023a4c443808ddaa9c20f607bd56c9c51f2a0d055090c
ze749ffa4fa0cd4db9cc9358027e4356ea681a37db233c2cdf78083342e2274854ae71569423654
z30cf2d2f70971c40d00cd68fda12bdfb3a20b0d44679e135059d439d41c55f7c4a2387fe8beccc
z12f004cf42c568290943eb96b7b0f69fcccdbb9289c1fcb42e1fa464f7bbc5c47d37b8a1e22cc5
z6a5895fc501e3a1e10b0ca80250fae44cbfab72d4eba8a59ea03265b56dc1b3c1353918044bf8e
z3c1a5f5be6c4d3a467606b5fdf133a036ebd4a5d862afd039146210b3056b041a5c0d4c7c54141
zbe2e325f63b5f1eef1da31ba64e3a233ee61963b410c7d349d4672b9643971bcaa2486c80dbc75
z332ed59858986965786b2e7bbdefd5fe0143620bd7dd23b7fe6af3e9b28a983f6e9f53f5f450a1
z0599e3e9f794c9ef99be45bd786aad0a515a03a19a275687ad50f89cae481ddd7b39d118e92b9f
za4b40dcfea97decfaa5693714c8aed0425c319b0941d6c670958860621e6b1b828146b2c08b902
zff0095ad762fa22d102fde9589b9665e65784a96ce0331bdb739033efcc1fa1538757ca5b9fc38
z0d3a070995fa9df7af66d91a6eb4883fed8e4ff04b69f84bdfc821f0f2efac1632abd5b3f8d9f6
zd356f4ae753ced38dcbd6bed9ba1cde9001710b5001e6ed93ce6d9f6aca9f8199539b1fb0b4618
zbe5c7ab54527c9f8f3c865ff2dc15398a9df424aa1eae56327d5706d62d14d18845a64d83df2bf
z425b0f7a644f1e4741705710a7d7028d3fd58185ef7b42b01e1e5f419a40fb2e1aaad5cef7c496
z0744e9d19c2a13fb00e3aaed9f3eaa4deb950ba8901b01eea4ab7a5a056cc8cc5b4473307fa8be
zffff1f553fa635257476716ee531d745fa963be468024c02053bb0a0b18289b036e6e697a67908
z9cfde2447058891f55787cb406f8e45d4a86ed2ec5a42c458f82a18cc3bb9f48d94a10b6cf2e82
z45274e04880550b1cecc081aff7d78d3a2c47db7289670c60c3beefc708a65790192c65cf8fe4d
z36abd351101bd71dc208394753c8bd9cd198c6fd42ac1e7fc96b28546192bb6eb67b676a27840c
z41835208ef2754feb6984fb7bd12f888afc0f61a9cd8a16479c908c4913eb4c5f063b67099b0e0
z46dad6cef23b96dbfb8bd64efbef0222692c92c7b556496b422ae494f2dc67d991581e9cf074f7
zba478cf324766b4bafe5b933b92e3a96c937aebe651247828045aaa56d6e725ecc9224517277d6
z9f1bc85f542d3b2852eb8e365ece2d4de222694698cf79d3e3ba01d389a8ecd34b09103a8470a9
zea9a7685a7aaa011188eb0e7cbd06cefaae018f5188cecd1c7918744494563ee2c4175a843d22e
ze8a4a6d68962ed15b43bea755a8210abbd44bb8ce566bc547677e1e541ead5dcc7fefe241ddf6d
z6cb95499ffc717b13e19b3800d1c58ec0c4f9ec7a2d588989deee63dcc5f1edc6a8ecf2bb2dfe1
z92c51df12b10c421962b7b5e06ce956ccf0c9c3413783330373e33db2e33104979819c33aaea45
zbb8151294fa58bfd0d2036a5153fd74b8651ee387baa644fd5708b9a28ca43302a7ff94d8b4c94
z73e730d05a47e511c50b259415f14928aaa7ffe2ada9581ca08705f47035f32105aa49b8c54370
zf6086c2cd7c6ac9bbc727a795050f1885cb10a1d7a32a846191eb2b3d641dcff9a75912eaee5c6
z67fc6da8727b5d8752452facd7dcc456cbba9878983d09e6353908cacebd43ea0d124c7084da15
z3654268d19edd356c8fbb3984ea69f6dcdeb96db33b6ce9b10199af9c4e169420c60929554b9b4
z6a7e18a41bca0a9045daf1a8e8c48e9cccf5f409e4893b9ea8f5f8e5a6b738eeede9c95aac8e47
ze9a4c52ad8e34b53a1239b8305df27d83b3d2a0db209fd9f85bdeb7d08b844116b56d51d0b04c0
z5bc5ff9d92603cd3dd775f39d3443090faa5bbfc884556290a4b8ea4fb712f3fdc5a8cfe30f8d0
zcb059d394071a8a7b056504e0399dd89b97a4e8ea269642a4435ba2b25253f6a8f37f842bfcc07
z1f005ea3531821c1de3c1b302ce50755f9bfce55144c86deb01fc70bd432481d1217f631d7232b
z9c7d853a3f78df811e43dd66570f475b2382da7bfd4a9133e5dae875ed42788ccc3889b604895d
z4e871f47a3913787efc85493c37143426ffea4176fe5dd24f03cef0ca331e55cbb3e6ecf99bb4d
za878bf404bd7e5201618d024542c45f7a73a2acf00ce65b65aa5f05f6c7b1043f911d29a4aa948
zc9ff6c8622161fc844b7b2dc8574f669db33c5e0331d34403b5b6898fb6a74e8a61d7afa43d9ef
zbc772162308ebf2121c8c2deedc36edd885d716e12097850ec89317734b2e29792f73294532060
zfd3e9166667b03886ed6c09813453a79ee30e166e954017c5fb9457238883464f137f77d186ce5
zc6b6338c29a33c160c609301a671adec8a8280e32400155748f66484b575489a1e060e9af409b3
zc10ed03032c967ff1b168fd7635b24a448dd44c398e98ebb685237eb2c3ec4a9caaaa5c131f672
z7fe92fe734a1792495c0387b1591aacd2ae273a58306c7fccb41cc7e0183f83168231fe712c8ed
z953362abab38c14bd312e64d72b74c1fcbcdd8981b9d49c328aa519275006224f01043846f53ec
z2e735458b41844ec9db139af668dd717f3fb9730e592817f89571a46a3660d595a0e20317babd5
z0ce20c2ab0a3f32753276d2b30cb15c953068e711ad4cfabb524c5f308da2cbdb4c2aa6ab54e18
z20780e9de110ddd5d6fc0fc3b43a13f39edbce1994c089c1090d5b0579a624d3c8f38b68f93e33
z4ec7357e303443b50c7e2000851413d6741815921bef66638f076ca0b93056a845c5731f3dae77
zaeac4f728d9100ca9ecb78b2569da15b9a10bafca4159bfe93a6e0a7a9a481c36fd51f71e24182
z8a92c0f05d85e7ec0914547a275f43f7f0c2d749726b5edd4ae518540f65fded3eb140fe96b7dc
zd73a044ffcb3050c022905c2f3203d36d66e7ec60815f05f6ab69a165f722a3839e1248cf92ff2
zd52830b5197d7d9b7fdfeb259fbf75fd3304561a80bc6a45f58dafd7b6a8874bf902a202d247ed
z2ecae17c1f2caa234b65e0dc7c50e04d79d8c80d41c25a5fe6c0760f109a87bccd66f53db2565b
z83a5000ad2d5c94ac3644b6c8d36e39ea77a127d743c12f2c3a3d781fac50f17e8cec128a8fcf6
z93566cf8454b25934b15cfc09df784553ce3bbfc680603ec287758bf0a06aecee2b2d6e2c1576a
z18c82a9ea853b82e3f752deec6a0c82a2e8630a92ac860769c1fd2dcdfa7c33679bce36c6012e0
z847b53d11fd667576a07dfa778c685bd48fd5fa268c103c741fdc407071c1668574c4abaeebd3b
ze4bd1dacc515e13ac467971c408b67419a2664b21581992b5db7acc404a6aa8c5dceabb72d189e
z974f28e82f2cc79c278f840dd153f197d790d94cf35a59a3be5167168304eeb44f6f92cd9a07bc
zde6d91e3e06ec509e9882caee792a0be2cbc6b65d18e58f87e59b1faf85da39d1d52dbef231585
z761915ce78123f06b7802c78b2b9649107bab1c336e524e25312dcd51693979d964152259507d0
zf8c55a06eae0e2020fb75c5c780a510a27ba2b3dac0f5985b9f2a434b580b08f4a185a684f6b50
z6445ca7beea9573aeb55bc4dcfe40f5c403f0082694a3796820c4d8ee9364f403a8b146a79bd4b
z24ad0a2c82f44cc03d6da4b125f4b074e7164f5d93880fb1a4e698fa8f043b273a145906acd28d
z481904e4c2a52be92b5f972e41bb1ab16d520be6b0e9109479a9786fa40b7cb4e5a95d0059fb3f
z4aa47482bebdc05b58827523638707fb25c3d5054fbdfaa87f63b141a7be6bdd27ec1cb3dd6db3
z0bea27caadcca77f25e6808154c91f08c74d25a8650c1550a0c551cf5620e281e62cbcad303b03
ze0a62f05dac53f663616077983e7b52fcdb9c63d8e90ff1ac8d2d52a702b6819f324ebc5160d09
z9033b71c02430ed7b8af2eb90f87de39f0bb24754278bc74e150d0655637643118685ea47d56a9
z61d350549f1a38ea3f6f50814da3d48544c1f6621c3d64f414adf0b5d2494c7a781601d34898b1
za70ac65460e51f2a82cc0607eb02b3071c356038c11909dbad873ba71c888e313c02abaa5b379e
z631f3abb65722fc6f1e37e9a54e288dce44aae7a3e68c480d3196b28991c8bc5dd19312a027889
za481bcd4534566e49ff86de5e9e61e60cfee4565418c71085719f0d3f53050578903d6db86523f
z86714067609186e91990840aa1b5f789d02d0b7e35c7c4a8ca2ffeeded4fd6c3b5821859685c0f
zb449f146df6d5e3329cdeefd1ca64b571d0dd6f39993a467515f44870c6c8180d66243b6d75bf1
z24f49888509f76e678255191c4d980839de3f34c50e73635bbc8f5f8ddc3c57f9fc988e443bcb0
zf91766c4523e3562c90c6f0779bcf3d5bc71988ca0782b0571918e639d9f9486e6c6b8cba640a5
z72e375fcd93ac2507d0c5218612fa115c2e292a3fccf2d2db82beff0df492d48c0b261c9030614
z9c1db18546a894179d06ea80397d4b1fad47bd56a853d2325787afe6d826ee1c728a9cbf029d6f
z542be5f75b843fa85f71b0f9f3e3d11ac7e8aef43ccccbe0e497ef6be328c06794be3ab16c9354
z509d4d59d73bd4198fcb50cd880a7021415278991f3ee6ef7c55e07c56b1f1523d5d5a56d49108
z26fad27373e5a587fe894b1b78c02e134c7fec48579722b0fcf19e057ba3384928d177c5ab8a62
zae1539f08eebe5594078273ec09246fbc43c1f009a19571c0b99ab63c757562979d1b1718722e7
z3aa7a5a4d7a38fa6a109fc8436561c347bf4fbc89c6e58e361e77d8b987f68e7b54c29a0a1e2fa
zd040627580662907c78386a093c3e30b77e3e471ee27e3f6440a8a0d1d605892e7efc845dec0f6
za4407df636e478a79c1fa1ced94d6a751f6ce0a0aa04e5945b178c7e020e1c83d443c693aa77e0
z022d880c72a8b4bdf63c06cfb5c4111d818c0ce60f7212589c4a98a4577160814056359d2cb35f
zc9f35e2b22135c8296b201b2de06454d87ab9387b693bf771c4aa5c919f7dab45197d82bd7b417
zfca8fec4ea51f610c5cab8c347b2e8279d4ddf3e9d8a4cf03713460f28fa64eecf4f45ecd32b31
z4a612f4262aa896c38c60d7bbb54dfcb34de353e0b790a719c3105efa853355a832c45e3e617e1
z4994976e89cea541273fa30a7d1af7c91083ca9e5b41cffaaaa66fe218b445a82e32b0acac01b5
za1162c1059d01b42f77ed53913b1662bd15fd21e850d9eb6454baf4d42e6641e0af57d4b39da48
z3f48bf2ba675b0f44121f976642619ffe47e03367d182c56ba6a026a1415f56b1a2cf8294ebdf1
z831d30ac69ce91303b2c17612174e535ffd593d4f185fb79bce5e9dc6acc46f37fbdbf532ec094
zf3de82e0f2b4d4c30874ed90e90acca59c5688a05611b860f975807f1b6a91bb5b3439e875a22e
z6dc2540fe3acd9d62ffbada67538c806e76e4a172d63c14ea12fc56f5316b58750dba12533844d
zf6f2d6604ca59521868facfe5694fbbe6ecb098f440f6552acaf2f0d94d5523f0c532e2abd01a6
zf184765361d6728bfc899bc5d6451edaf079c74d3d4ed16173d3ba4bce839271bb13923631e2df
z60d16de599a1e8a84d3c728f1533e862305adec6bcb71e8b1943f21555f2c45ff79e05337349d8
z8498f7eb104225e9a0ac727364ca7296ea1c3cdb510abd661b89dddd639f0974506c4817c6933e
zec4cccef5adabedc4ed5ae4cbb5bf508fa8b440fa158737dcf0a66d3c9c6b9c40294ac3a6a2429
zae1b87a38a86ac9bc18f82e7b089b0496b0a29e24d1b2e39e3a05397d48a32b2c9fbbbd35a87b1
z9bca34cb22baa7bd7aa71a4017231cb7015872ef124e583b07f3d801c78602f64308fcc7154702
zf3afd08d999b2454525e9b551d4a011a020e333b1c2f288689ddb83d87eab91415721d2ccfbd7b
z3ee4e83499f9a1335b71526524559354c4bab1b64978628cb8701d75070b7a5488b91eca588eb1
zd40994ddc1396949ca55865c29b3bfd6f188fd7627a9bf53d8820ce8081d1a10ff0e6ddd1cb073
z1add4fbb9642556f8aa4475e3dc6aa4c1d02fc494f83655615c562df39dd4328fe93980cbfc485
zf31df1cde50eb3efb0031c2505639562641a07fdaab25cfd6a4d0a1b1dceed5bfeb41bfe73ec70
z22f17f452020f8e9bbd33ac3999c43418a7cbed316bc6860abe614cd21d487e8df153e5aa2cea6
z5e0c49e2f492bf72946cc006808cb3b46576aba618b54e9bac8d1627ff4ffdc97691ad53067d7c
z03c691be38e484f187c7ecb0a6f7282902411946aca3b1d49ba9befc71c9810318c22a8037e18d
z76a82c253cacdda307fbe51d90547770b3014d824c6321b8bd18fda23c14e52ae0e5748dfb2f44
z6c5521f0611d1f8ba8558f1b92ab2064ef142da218a322d6c24612a9e2b7d51c3de6ab70c094a6
z0c870ed1daf20311aa6274dce178071e13d26e91eabbf5180077927320c366a5aeacfcb3016618
za06de32b4e9468a69fd744dbb7ac00fd18d2d334b38ac6f8566142ff938ca3f34e4991f04f6ee6
z46cd490f20fe373e607ac6c7b8b3
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_back_pressure_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
