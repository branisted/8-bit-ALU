`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc54b3c9b8
z81acf2d45222519b03045f223680651f0ad1117bc11c20f6367bf7e55795f5a0f4a9df96ac1966
z6065b08f032279942349cc97f8daa0ce07a74f3bde6cf66a7f7048b99b482a48bc9df1d50668de
z50b477f14dbf58431e426d8cbee91b76f6eed260b6f757546f0e2d5d635f1177ccfa702757920a
z51f9146570876fdc03fed5b0183b8742732d3c2a300b3377d42b439520304ce8d6e50aad71f52e
zf106d419d7f30d701593c37c5ff55096dbecf6663fd9a64ab33f0867f4cbeabafa199dbd392dde
z4a3b07dc39bf5e090eb330956243a9dcf02ee6a5d02444ed855f00efedd94ae21c9830c41ef24f
z338f34bc4ea636751b5ae42d80727be25aa791bc83289e08a6341e57e52284457fb6b97bc723f3
z4f3d30906a6ee334e90596b6ec74ecccbf5f4deb8b4bf0c94faad32254f75d011641a3959beba0
ze70d38efabfe724fdae3ccfba980a27180bccdf96fd78f5df7dac37bdbec5cb781f594006152a3
z0627862c288a0a2e5751449ca24425cc9ed66747430c6df01f4e9d42dfea57d9eb44b40f2b15f3
zf23caecc2cff56f4cb36d47c8b2bd548fb8027f4929a32f617b89a75dbea399e4f8fd82768d9d3
zee9c964d385fad7785d7e4a612800f9ee6a06e636bb324925d903d89fd62f5874a8c147c1e9518
zcd37f55b2d17035bca1dba06c3c0fbfe0d9126373876c2edf64fa808a37804ba506a253683b3a7
z81445199999031639b697ff6738e1bdf405eed483fc5c96e402c262e325977cd704872a871fc29
zbd28a92f3c09fbbf080fca5e02d172d18ae5a5660711e35e0d60b5cf35a6066d975a30c3b6d2a1
z60ff82020a762ee0bb21e0b7745114c86e950bc2c433bf62fdcd01830f0936c7b211c77f468511
z8f3544692c84b2ecedf09344a437471f5d0a2e7e00b2f6c9f050b586289591b83a271620ee07dc
z1ecca334abc6c399e2832257c8e2518aac3d8f78507be087a427c329602d44143df522af7975f3
z1d737ca4ea081f0c52b04aa0db940272241a175b3c1e40170d0d2a4aa82af08e613cd9858156f9
z02813671ec3a1103a4e550013a92fea88ba53ac0a54b6e25ce27af9581264bde58f2b1f8c26472
z6e111b38e528a4fee50b8bfa997c54afc56ea9a915556e61366ed4e0fd2703a5df1f855acd0446
z3d5ca416b6d42d20ffbafac1068da022d78c6c51fdba33265a1c32c067dcd70036e15fc52322e9
z3c4926609a9e587fd0df3a361a3c493c3c285eb4e077dee8f3a922c64f4170a61de6272e21a9ad
z3976180e79be51e28064d1dd600fd80f3191ab1c8d61a6391509767139645ba162a41c0bfdd7e6
z63a7fd866e97bf58ddb278680ecda4ba393a01ca601fbcafa02422784816445c9d63722a04f51a
zeda185e7476997c15edbc2b956d6f9aada40f158c2811e77e547b08d8159d235c456aa9ba1fa31
z74e92ac323f8e647459f3699ea3cc74c546664b85f6e1b2af25d087f6977f487c559ef283549fd
z97671f03d5d2c998500ae378fd06f9b5b7431b4763755a3b8f1f63ce192cf081bbe3c38033af14
z57e8c05e8efaa88b2aaf1ff8df3555aca494dabba0e53181e4dde5bd0175ed3d130927b336fe5f
z7a5e75b5eadabd6386cecd72d71f0c2446b7ece1bc394b4c5916ddeb95c9b8cc63cc718e67fc6b
z5aabc10f787ab632e93e2e982ba84b29b544ad3a730b70241b1756fbdb8aaba98e101d2016b283
ze6b8ad0c7db7ab323436e00530d86eaca640ee83d080b4775dc3b438fdc69535273cee0f834a58
z91488c3984a8aa2d9327369b6f9bdf14b6e758ea8ec994b001cc83ea2cfdc0874364226fcc516c
zf865f4e47a88d7d644495d7868bf4b4f7e7a9c0b578c0a40ca37d588299f253b5965b1c2cdc168
zf96c45b24a518dfc549b5b387996145c76df6e9a402e1ae7c727f38175e68eb06fa65c91710c6a
z3340af9ca918132d8949d62203ee7d83f2ac54511ec09d35eeae81cb6c19b17b97823fbf427e74
z5a8bf15b66e01ea1cdecfafec28b9f5bab6f25bc588ea5520debde148d769a67b79200b22a9fd6
z98205f948ab5887cd4f2b469f60f28b3395640a1e6207205f784173eaac0f2e69fe8f3ef871350
z121f1a2c7b38e41a8ef2194b5c41fbcbe65b7dcc3c19405b4788fafc1cd5d16b37e28bc1e0b4ae
za9f4360b9879c3fa93b386d842e7cd88445ebda794fd495cd422fb445b48968c0b9ecac2ada1d6
z45712810f079ded8f514f74c189b7ccf3d792741e41bd05875a556e64c80dbb342b35fac7acec1
z09d4500676fc211477080870e2301850eaa21eb582c1b3c381e37189b18d026d0669855bbb4159
z6d7090d60b8c7008ad57816131ae2d3c53c496828a3a79bbf9cc0beaa0cd14bef1981b4666e62a
zc827bd9bc9a554eef19341d40e5c977cf2d58d93b42924dd702f04f3169b09ce5ac3aea7d714d0
ze1de442f64b325e27d3ed7b182910198b24b014b5fdc1bac47816f9d9b08bb087be1117475b4f3
z4be68b1c303e54eb4dda92db8a61e749d62146094ae928207a736b8330546f3d3e4170c3e523e2
z83d2a85efcb25001d04a37912d57ad9687a29e5fac2c1e8f772d9bd44353d58790d3006264c1f9
zc5ec4395e926115cffe2589bb45ef44dd68e378619f61c40c34b43fa73d2c1f2f32a4c791cf1ce
zc254ee1e02d4e879a8569060f4721adf199697097ff44e5b5d87e38b72fce1eb162298a5ff05b2
z9aaebe062eeb3adee89fd757bd5e4f9c8ede9dfd19e90ebc4f22279fef9d266244d59fa3c17c3e
zeb5a9fcfb7182385d40c90ebb77cbb4e4dc67f793f050db7d75318a8505db8b69c8c3dae6a5455
ze7d8b605d887b7b966e2d7f7e3218c08d80ef722b3fec64503a85d60a8162dcf10b1135c8e8dcd
z986acb1c8a56c7729861b73e25e57e74d26e62eea99774e74a5f53f23060da6f8b4f2ade042b48
zef98d113642b372c6ccdeba28424f516461df3e810eb8bab24de8dea0d585ef2fc90ef888f66e7
z9a74e2cb0af6de92f02c68f1112ec6dedfc52ebe114c1d8b93385c01a33b309be2e5961b2dfdfd
z15ee17b62774848ed01066b578f14d8aa1688b4fd110926bfef89ddc8d495e6323b604341ab852
zae115cc5b7eec5f668a5741a863c5bb0e626e682a80747eb41784f48374450b8ec34c60be40c1c
z1e0910a3f637d4b11ff2a17eb3deb1bd03756f04f8729a1088e9c4c9aa5cc5f38f00455e39e521
z5067853f2a015d3deae69892cf6752b42c1c9b86c1bed8a1961539e89a587ece4339ce0806d20d
zaa3128290f1574dbaec1572e6dee992388fa3c8be585fd0c2bff8cea1772f131f7cece2629f1b3
z006bc165b6b85120f369fd30bc0073f3fab571fd54d8c82bf1f169dcdc76841d60adae86d126a8
zdee14a582039e6a47d8064e7945191e63ea5914be9ed705dd9b922cfdc6bda22e6848ed8ddd4f5
z819f441f90e1a64c0901a85dba4285644e93b4697f57ed3d42946c19e20c455c8137763fbc2b66
zf1c9b1109e1b13b8b3a327f556a821699f0fa0e6fb74d83cc1d11e41a12b4548c403acd230435b
zceb8a497a968ce152f3632a9526b809743c92713929fbb6527a712298a2e95258b4c12df1c3c73
z6c1e59ab80c3113b766149d3e7bcbc628304f4ba7cb0a24d4a61ef33a9d1bf9e788ba9d7f4f22d
z71ac38b8151f836c55dd08d52a62dd1849fbca7ec67a1107fbd38bd7ad9deb687c153f440027ef
z642cfea95b2d1ab8dee5a0e8c001310048416415b313d4c00ad2384f7d64e6d095d63702c682c9
z8a78e6dae72003ecb607faad414b4c5db6ffb4f71ead8ce54917d88273660216d8e900ab1b009d
ze645dfa5d6ea089779679f0e6f87a103e4b0fb1ffc4cda2b0c3611d6b787ce100fd9dbef62eb81
zed619f61d0b6967843ebe6e90f61c5ce1aac506d6fc18e535c90763207d132634f7e98306d62a0
z1b73f1e8dc4fc4e01b91e61b7842a6c3263e298812595f78ee34b7d24d74ca0f456dc23155ce9b
z6ec5ba09cf342423ce93bfc9af2f21472f95d312695f8a38ca02ecff4f2809fb3c60014d17d8e8
z2a088a1d6a6e6a89be8f9f8a56573f6ba79b532bcaef93a53772e8b4af36c07a0856ffe6869549
z0393c6ff0754614150f60f61394c8139f06ffe271462b63547929c87a749eb9869b1b710bdd2d8
ze6842c466c3b93abd851b900d848727702fcc59ea0856cc8b82166b9eec5f74d2bf0075d2f18d0
zb0b8d3cf04165c7498e0dee13ce054041638ee67449930ccefa8cc8e416da69a93cfa49deda114
zc16be0886172037c8e94a9efb247b65820f3fa1e90491dca25f3f57f48c06b846d5e6e016fa1cf
zf0b620c22bcffe34b5ef358126c559cc575132a54ccd2d0cabbbca208babce68f7d5364ceb042c
ze217994be5e91228037d68c146c84b6e0484ae0af9b8826365d2b747bb7ee728d25bd50574efba
z6c96e1ee7e1b8118d9d7525acaccb1f084faca377d2334110648ce53dd075685d1a06fcaa8fd7e
z47ecb765b3ea3a5be853a7dc239af6ae3f36d25a3bc7b496579dbb362d31d33bb0ba3545d9d85a
z83595e00846c62f87774d050e92d9d74b4a9a85706de5c721de418b2b1a045b2003ff013ab4711
z4886b32af26704b750bd11afd64bb615cf34a899fa8db43c9a3c004c8bf80c9320cbc50fa123ee
zb5ba9edc4cf77d7722747a4880ae9ef5724da60bd164317c42c77b58ef8c540c9a4539c27e4e10
z2e359341947840f3afca6ce0bd70994fece2fc445d723e81b2018e2fb4787f2b36de5992a562c8
z210883a4a1bc60c363ff97504293de27fbdff6e2815d0e60d291fc8a765810662d0e229a4c79cb
z1c994d6854e301c1553f1fe485c5992af5ca0f657ed43deae7069cdaad9ec344f0dfeb17d0483b
z1f79db2fd56b3fc233f06d4b55d9627a6878c46824770ec81604ec4374cd3310075e46a35f99e8
z70a7670e9a1de9c2555e2350587e05ebc2ecd171583034a2279d1d500e798746724d5cfe6b680f
zdd9f9b3425858334591226c532b9aa1cf1c3f9a268f88cceea8c6fbeaa037dd7461b6c183b3d73
z12b29df602a2057365f50fbff4d4be17a0a5b7965a3b0b37c0ff1d7403c07faf7b52c2976de632
ze0a60d40cd55f20ce46a3993cd95de82074989dfd8cd61fc13963d26f46aca15d6638294d0233a
zdbfcbf3fa3b203f9b3f32210b4f434152debe6f5b1c31f1fabf9d2b439d8617ccbd2622771046e
z2d8afc80f57bf6f770e92fc53f820dc58a98702aed53555e1a26af096da22360ef182fc5809815
z4b903e7669e28d3001fbc5fbd5f99a768da81336bab230a130a6ed078f20d90ca111dca0e13a77
zb01d9e652e23452d69c895c974495475c11e345a9e203123b45b822364bfd1cfa02402f90fd65d
zf57cb4753e67a33337784b8ce9751e154bd9f798a82dfb81d8b61ddaaf3966dbccb46318e19267
ze5dfeb89bb2805c96a902045140c086b215e565ccea1f390620c064fb9d31dbe101f7831189097
z66a17bef15eb450e553db9e6878389da27a6090f413a093204b017dd3c2b5ac3d01a32daa44f21
z2e95867565c773b7c1e35c95c54393c4540c6d86153049101d91ba6086c8c1df10a7a9699fb21e
zcc011422e01ed74acb3011f82d4843104c5ef0d8f7e0122a5cf9f59282455afcb84195f19f73ad
z6ff173706e24d68e940b750b46fe46e51d35691e672822395a40db643fd52b323e3ace68e52118
zcbd425d1a4c61d129526bad67356fc95a79a0acc803ba1386a2e48dba8a6e3fb6ac6a6f08ef595
z8fee4d2d8b645eff3ef19102e3cf72e3e041af816ffc31e25b4eae14d3ca5e4b9b626c88976aa8
z2c2ac0f07754a02437978e8e8a12a20e37b2ec09490b8dcc94f36fb006381f1a1f8544e132e0b2
zbc84a1481d4f5b6c1a1b7e5c5ad946e04154be1133ef128ff903d3ff5f69d40830df74a9a71567
zc0c2f81dd85176290c085679efb77935943c874c9ecc7a5444d4288b4cf3b229be72c14af63cd9
z70cddf640d291f0c872b5679a227aafac514e1440521995ab6593143581f2f91e991fdc91183df
z863c89bb015f89073bd3ae95659d5c6c96d59af98085ade252376488b28309edaa6eaa4f22d6a1
zf83f40d4886db014807b2c454a83d8457b9b6a971e703c8b0850d806549619ba694fe90654b02b
z2fd2d6dc809fcafc23c482b776dba8f56f720e3f5d09f3a406cce84982b9783158986bba992dc0
zf2a51ba563696743b1d020774c6dc1f3e870f72926f3de3b938928616fb16b298c49bf1f8fa7d9
zd832296fe93a47e4e2a6263e9260a708e593e582b4b2ad10432cb7b3fee85f2913f10a5eb33ae5
ze3b1c655933dd2d947371075e5e11bd097aa40ae5873107554cefb22827e114b8e2785123654c1
z37a0c469a03eaa3f37c27a62736dce1fe8a19dd72f7a1b681d656db805cd36f748336e11a846e6
z110b70813dcf11513b4e2970dfa9eff49b7bcfe8a8b4d148ec030a4285b2e913be7f9e9bce3f79
zbdcc80093139c7bc3d83ba32cfb994e19de5f193b3eb0931cedfdf3b75e3d01554654d5ab466d2
zaf547adfe330203a1bdcddf3d15e851c299b5e586a0fa9db3716b2013047ecf7a972420715f634
z92a7a1b25e2d316338adcca1703c679fd2bbe68073d83e012fbcd1dc7d54f1cce53abe21e2bf81
z65537d8deb525f9f31f93ccd556f3fd761d8b6a63f58cb9d29f938be18051d200bca6b80df0221
z86f4396fe0cb6338554b73a40f8d4c23afb7814af20047d4c8b9975972f0c4eedabbf1f8bc998a
z6dcd9d477355c99bf1a3a7bc76585c2345817d7c689dfd74e2828eb2d61e99dffa2ca8fde437ab
z0e6361949e7992e51b687751b7fe024b043be99d1108e94e078eaacdbd4a4c0a3dee19586db1f3
z226114d13a7546629955f139b039ab20edeccb43a244c60f468bba668b9a9c0db8ecba0331963a
z033ce4737245ce0fdff76975c4641edaeb39c4380856c896c62ec930b855396ba010d5130eca09
z890b5738eb2d62920110bb138d699c9d2ba058939963d4b5c2e44e10cda88d4fc47a34c465bf5b
z9da2276c745bb53524f23abfbb1bbeb51026f35ab6e537960dccc4309d356f0a85c9ba1cdfac6d
zb187ba7c1a47c8881406e61d06cbde54984c241479b57e5c28a9a95b64a2eb48e00415163cb204
zd48ca436cc5d9ca98b0516435f01e612b1c1f4a95570d4070377cf090564b067c200b1548de081
z16bfce5936493ad1f1422d56d26183a3841f8d099818867a6b248cfce7479d5baf183410215819
zb6d01f7b4884e401de78e1a3dc9bd256f7aa49c96ee8f1f788c0cfeca0e8f831268fa89e8e254f
zfb275dcaf45bf2daed80928130caf4b19ab4fe8b3ecbbf71579a8d73c989589e56559b216213b1
z38a57ed65516dc65b64d0b0b4e918cf0be073e0054525e062160e0c776fead193b7201f467e308
z81533c914c55a92bddd5637da17f519fcdc08c0b166ada00f5ce5f6af9a2426d8d705688caadc7
ze4aab1c13c507d4bbbca23ad7fdee7cc4034085981ed2249464446b3080a6d20ef9afa2c683615
z4651ec9501ab27697e42125b473f118be5933ff450ee8118da1f73e7ab57dc19b3d606e3f989ec
zc3e5c15667223d679a29587967b68c4c179f9ace45a6af32cee24ba5be4f9ee803ae7d52f4be97
zfef9e9c7bd18590f5acfbeb9e35abe70eff25f4937b1062c6e2edd480a36407917e9254fcf385e
z56581b484a8f455048da6ad78b39c69f28bd6de59b6211d0ee907545ed1d58b2b04886b5fe7dd2
z73da0f994c935e0f9dc27f68f83c832bfebd3408774f72dde60b981463f1da275f16ba879573a7
z0f26802e78141ff04e98e65e20badcf7dce34523651bf6d708062951d30daa93ccefd4d2c45caa
z1b306b5fb7c7505200121d8176dce6f80e07f98b7c2004e4a4b1385e71e4fbe0abe4687706eae3
z408e6d07985e37f9872a484498919f623a34bffa3964227209c14f3cc54e594604283048c701da
z6b85eda98718fc2aa3c143e11e479ec4f27bff8b74ab602aaede68054022bc1837cca4ee553488
z90e1b87b94e49ef03af0637341b1ffd4144028f1e9ca63501e3059c50c284ef345b0be864b3b9d
z65674166fa4ebbe942aa94f0f998807fd88b786da665f0a2c11cd24ed0419435a483de11add3a3
z6833e8c5412f0169334a1c478b3cb1520ad9c11ed09634b57058a463f9a568a8cdc6f8240975d8
z9de83a47bdfe7c300923efa0a4c145921f0bbcfe24d3952d1cee94e1101e23dc8227da10892a44
zc04d04b2f7fe9f4267f68908fba1c762c06a1d82fb769efa7680f8dac79f6a877ec1a146f3a69a
z1af8eaf1eb83a9052d21896936756bf5153e6deb05967e57b83ec086296aedeb4368af667bc200
z17132a65a93978f183371edae3e4be27a8272ba0f45a9db1d488eb2e129603985a5de611159947
zada279c27a5ddb5ff02b47dc37b37475d47e3ee56fbd11360fd1f0b0ac95e6355f4d5d6dd36921
z730a9fb14412681483c692aa1e0f28225c8b8c35c6b006434f8bacb1e13b896d3fce04f4368814
z0d195f5e0cda91187cbf2cea50c367d88ff535722dbea028122a158835f49cee3131b652b88d8d
z19632d619f71dccd6a94abcad416cf7a5b9c4e42bd53061d437eaf6411b6fe77845f255cc04801
za07a2df20e3a343ebbe76196cd3b9a67f51bd76a947ba377e5542754dd568f10f98a56522aa1fb
z6af06e7260708251363af050d69b9e942721b1fb14383317e12b708dbe2d5153da4280687b53e8
z172eeff046f794a57eb97efaf128fc65a365db4a77642dad95cda846b07fc08cca526f50591e2a
zadcc3e2e77f6ce0739b95505bc3675452ce5caf29fa4c82a8a54469d24b41691a6bda834de0003
zdc80a4e53afdf260081c65db0d1799ca9a5fe6747d7f37961dd096a9db1de41dcb8d5bef73bf53
z5bd80d173e91a31136bbfcc15e321beec5ed3eec3ef0fc0475d0359ba99ade59eae0c761e1a66d
zbc96052586ef5a908c926f752b9c2267a3b97be47450e5511da4c8c468ab6a13fb016cd3768b67
z1e6dbb213a8de98b466e2382ed11c92beb33973d855a5cb9324a17b9cd0a603c1c407d6aeaaa16
zf57135bf6073b2fb54aca1087fe39e0ad6c37e2a4e1c240073f4be4695331ba5213abac763b299
zfce62e40e574b90ad0fe93b5476e3cac00f1cb337586ca3626ab96e02beac9f3785cb56f07e81f
z2349f00c06b4b3b9cce501d4292e49b1a5dffe4961ebbaeb71e3166c938525afc3e79e40a22325
z420d60c644768537d4eb7262731a1c3c72b76c6fa62a956b8f644e417491eb9d6732ab961598b8
z1fe75347c5d84248ccaba7274d19d0c46b999274f25add068896ed7a67a1d1847d80c26bade9bf
z64752da0748c12a2af5f788d66ecde09bd5fe7b16c7a75c2e1512bae82e3591f48d0c30b7d9250
z9ac112c651b28364fece6d0448e7eacd4d02e7ed1b03530a49ed6a9c74e6743b3fa8528e035b2d
zd9162ae265e0709d62d9a03918c59cacd495483f77f1e915601c6128cadeecffd14fe3c7a8fa84
z2d4a3215d4b96d11601177c906378aaaae658d4e9c39b024c3dbd84445130d07faf15b55897f55
z4d8af8be90d45fd2003fe374d1f77908b9fb62ece67aafb9b9ad1337262ee4470c3dac74e9444c
zfc29e32e9d66b47133c924d5b7d8d9135c0be2db2b190c450200247ce5df049d072a8e195625bd
z22c6933e1f9de44208dd123bfdc0322c4b59940ea624afd26e1d7dd2beeac90897f0b0cdac3d52
za1724055ffe4e533802b6b714620ebbd1d4dc849fce0a888a290567d22066b7db42da006b48e02
z07ce486c0097c3c640e2170e1f995070c03358266d1b20bb05c28671eb8fdf3a51664d5fe74843
z10ceaed267724408ae1f6cb4f31130d5647c05e223f8cf5be9b6acd2d40d51d86d25c3ee7a79b4
z4509363c779dad0d71d07e5ed3f1dc573b6f6c0f733b22d392d1290f234136108b13716e406764
za5b6e5541bbc734fccb9be54ea13efad827021d3763f5830bdf678056e7b5eb6c609fac0903101
zadcd3c5a9d78c620f36ceead65a3cb13b9273d4177c166f46ca4efef6adbb930038de1a490ead2
z0adb2dffc73d30ec4ded95d7834b039fffc6de87d8eed96903b5fc148ce080931381d9d113f28b
za3d79c02000c243924cb3d9fa88c087f496ee9f30f3c94552d47d6fbdd8f58bbd7fdf35e2466ed
z27fd66b3e69d3bcc42643e4363532f1c0ba5dc4dd9e1eb176a7e1a4da62a4a825c68696a36f58a
z166a3df4d14c609077076466d3cadd1b32eb551b302037acafce73525994448c24b09c90cc49d8
zd09629271c5630a7e28c09acd447719f9487ffc0e6ebc92aec558b3da273bcd8d5ae27b044dac6
z9f350093dc8fe99019175fe0c0cc59730018ad5a3280d492d2fd44811f43a02c681dfce87f8dcb
z48f29041330076beadea6aa164d8b6333a40a083da61dd4b9c43915c2caf723d395909109c9d30
zeb6f8f623c5544424cb7b4c6121a68302eceac7a2f166bf93cdf173650500849e5d28469476913
z8a405e28c17768a2e2db308897abd38cc1c7fe25829721dfe2ceeda0deb95b825c842208849f62
z713491822635bac6a6226a63f98a16e236c1f2e4e1f5c0e75d34b430fab1f26d76590a825e883b
z8be17e1af5aed1ed314224c110b8baab0f2d2d7c2d26d6d11b41444fa9b4108944693cfbd11a2e
z9923408cd67ee1b5a67b94189205de3aba295b4b481281a89440daf83fc4878935f031db75c14b
z6cac8fe145375492760758f9a64620ae12f8d4aa1fb89c4bb06e6955231d1ea0d8576615f4a893
zec649ceb376e3ab4139b110ef8bd7950e0e495fafbfda8a4dd18e1ced6a42c02289c76db4ad907
z682e5b98a0e513b15eec6c7bb995dd3b63c7971bf17bc0f3e4d188f55a0fe9f66c2802414384cd
z0f707a6b31279c8babdd76b91fb5662c37095106da25d690e8e6b0c4b96c25db0f8ba78add3f28
zbd12ed31e19517ee5bf1accd6a753ab437fda3fec2c662dca0cee80cb807eedf12022a8fb2014a
z3f74e49f5e0b244c7a30c63c2ac6ee8aca504189fc8cb8ac46db9617cbc1f7541f7791923ba944
z2f4d13e67eb1d4e5001203eefb2d03cb4874e668ac7ddbb97a31beca5dad074be833583cfea115
z136d5eaae5bf48c3afbeb331a0b616b3f6cb02df75f8fb39d5dc498dcece23c12d03f28a466835
zd07bf9b3716b7635e4a5b02f19212dc8fa150b316688fba775879f0e984c0a5c801407caa752b7
zc0f1ae09887a4313298f3ba434ee77b7c11c69e0deba07bff770d6592900cf8a26e3b51eb3e749
zabf0ddc7ac58641e474f6f1e9c8a2f6af35afda8a77d483f1217a16df36dde607da3f571ce32cd
z3eec78690a43c4ce4e9a23fef93332d6a05ba089748801df5ad37d5f42bbb9f43aa8d4ae378a4b
z72b00a545a36fafada9774f01252cb6547783b0ce98519d09eb3da1b6381114500f446f044ef25
zbfff4645dab7788ee81667c339b28c99b4ff5b12e4c73f023f3f1be1b665b9910f054a1c01ed5b
z553de6833fbd2a2c5abe4f4520c1172f9db5768c5218ce680a127196e17be37f683e68e838e38b
zac07c444baddbb1073452d83e5b022af169a158c200e2e489170e91ccb98b360bac52a0a867cdd
z5611d97f7f4fb7466ff7f6db111f6191977ffa6688723a8820e4d966ae7dcb598dfc96728f26d3
zebf6cb4338b5ff859693df86f114653154a7ae8bb40ee0d12a27d5be1475439cf75fca59f41ac4
z357bbfabf79381bee5ecb74eaa7428ffb22afcb350e57bd42da112510afb1e1fc6cd62920f13a2
z4873670c9b6bdd5526f19b7790170c959808b11cb211a9c1b788a97ac3abb76ce36ec909fc6a58
z1509f140be79ee3b4a7833b10d23e2070f947c266db1bd11274172ff2e70d7e04380908fbf2fd4
z8d400f23b72ddc79471c8b6e101b6e2e38a95ccf04c421334c834b8a91334e5b3533534755b38f
z6ab8e258eed4260071a695876cd6745703df7d1882873f9aac20eac24ed66724e3d897a644ae12
z235662171c0f145b6fe3e269670b88dc36dc01bc5ad418ede81cd53ddd0e37edf0b76f2fcd3d7b
zf89604850f88080acc669287a9b7c105b960beec7c8d3d1195c9dbcd07f867e05234b6e749447b
zd939cc00e313964efdf1cbe173a56e4d02e2c68a145bd94d27fde6314e1f4068e6fdb7d80ec8e1
z7e2ed4c0bf1720036b348ae6c438fd76fb9ac0a669c5a56ee2506d6cf22025ec02e9be0025bd03
zb2c3687bd4b025f5899176d3a8ec269f802083b4e51e5cf8e2d3c1e6f96ab36907d6569334ae4a
z89424b5b29f41eb2471f9f7fe9cc511f33f3b94a2cb7978b487b3f8bc6d11f62152963427096d0
zcaeaa80c2b2f962c667008ae68160f6c08fe9d8aa3b027043c56c1cb5a9d0eac627b94d013eb42
z661d6f4840b220441050f2bd06c24e267f79be5a28c815f7f7c1a3e87101964773a025bffcc8c7
z243386015852ca15437a323a9e80c166c8e47b7eeef9443982b6a6b3ba0e812133c71f5de8b50c
z16a6b9d9a870810c4223e40babe2c360e4b2d54071f38bb7ecc9dae3b25054909885405fc6cc63
zf46cdeabb0bac3b5150b15366bf4cafdf3ab22acbcecea95e504a83ab59e1d6ae7be4a9c4e8fac
zc7e1e484fc60f2c73c59ce352016441d3d558cea2793abb599c0ae474c4721ad8b92d9ab03eb88
z7dfe389ad4923b80f196821ec81680f19aa5489e9374951701c512991b3a014fbda56f40808672
z49cffe6823dc06b35e722e846cbceb784abc9a8ebe1f16854fbe31738f52109a4f7086c9774277
zee488e1f829a76a1b70d20a502b1cc011374d6f03ef03510dfae6ce340733051a090d23981125b
z3367c024cd9137768eb1c0814d30c82e67e95b74fd2fc48d07a25ce7584e13df819e2ae3665cfa
z055568c6b05c91a7179ca52229266a6b153019b21c9a0db8810a4f9f9e0d2e21de880f57c14e83
zba827a194d8943ea6ae543c23e3b893e5e6eea070415439575a276cf812021b465424543130155
z6b7dbfe4f59126841a01ce184cee248bf5d53cca247db9a82d6666de9f85ef514e87570a66b4ea
z23c5b82158a2d4cb1e40955fcbf7d048019125fe0fe5fd122745a3c6caab58122e0f5fc0444b2c
z3065a489207420a6ce240efa415ad90d4784f3ca77bb6de14c1dc5155a766edfc0b94e46d5c671
z7a3b5ded45e58ebc2f45df82ec7428d4ce9aab466ab9d0fda9d5cf53946e7128289fa44e9e679a
zff810c57af46f648a77294697bac3a11c3f6061d13830256e88326f315ca2c9088bfd6ce62523f
z90a87fef13ebd90fa9c782762fdf4348fb6e7cc2eb7944871458331ffc771a35290e5187995eda
ze33c0cdc995a2346ee87debd7abbb9af95c988b025e37842c5f522aacff3acb2bcab1272779d6f
zfa5fcaed9017a8b600a761c40082fbb6b843664a50fc3245513ae0da92aa509a6c873bdd3a86c7
z52b62c9bd0b687c4eb614207bae4684c914c1c169f1e93984aed83a27f3f8d2f43d52da7952fdc
z36f60723463ff6bb000011cda2c3d443ddfdbba7de8785a15acbc94cd0c4d4e933f7436bc773c6
z9c9e39296520f59972710f4f0de2f029fbfe2d385d3b018e211cc1d69c8d725576a0f95be6fadd
zf6b93297236fe471e5f9132fd2b5473ae511f8e525cab05d4e0b95af1d76684414a775e79bd6ba
z3c8a9d8e4681476582900cfb98b97fb54b32f1f141a38fac7af043ef42784800736fe997e53561
z0ee6b6b6a09a39fa670879a60527e022886ca27e587ad5a3fd14a7961e037c4b368455eca5e565
z553c5eb7b3ea7e5c7b756fad4836a14fd548c0eebcca5e9ab5a9c652279ddc6ce36e92f5231651
z413f63cbabddb73684193f021b1b760cf7821cfbf71f4d4be2e3ac9a90639d82698d6e961c547d
z97f504f905231c2f44fdd4305609376993a7eae4edf822e2702edbf761d2ddd33522e35888cdbc
z00494eb0c2b8b8d597d7808b374dc84cb220df5121669cf1fb8fdc091ebd6144224e2c811e9c7f
zd56c646cb9c2306aa851c02b3201c26b379519c8a068eb6024d892f6e45aeeae597cf7effa1c9f
zc2cf38f468eb7b122c9a332b366e3ff8101af5cc71b6c417a474fb415d9f82e97682d17fdd0b25
zb58876f466516ec3d1decbd0f8c7ff4c6f7ce7cbb46620eb24e8bfd134ff9b9c388b89d4693731
z77d772adf814929cdd1ca6bae52a53126ad3c92de6f961e14e3a9ee8957d09cc196f1b7a8c7088
z28fcd96a4afc1157ec5807e84cf1de2210c178b5fded1fb9d06f2704f0f720ed90d2518e8a309d
zce75281c5e1264af0d798d261069998cd760ae7c0798aae2277b0d41b074301833de44f3cdb467
z1834e0607b5b39143af2093deb69c4d3c2e0e168eff3f6bd83e461b8131b22abdb6ff2a681ac5f
zb1dc0e9b42626383ef8f1993e7b273869bb06e8371502668508057f9381882af224d4e19451855
zeac563984645174e3aa9ff8044e2a28fa886f24ee85130b51d5162d54ad78283156644ec93d65c
z1ed31277b3c5dfc1bce53e4f2304e96e0b6ae03b5a9862374a6ba0b374e5df64642b80e3e121ea
z9764d28c428fa9a087d8472c4b6dcda1a70502378d994da5a74966cf6271fed641d7e3fd8ca2ab
zb4fe1efcbcc9c32c2adefa90ac5fd75aae32258062a16a3972c40f5cf88c3e6d282cd4cb8ef52d
z1acab6f9bc70d71108eda083f2b31934a65642eac1b0198e57812c0ae5efe55316204e3fecc123
zc24fa5ce73427c4e293a479df4eb740e1234bb0a935f0e9510887784b0170b06d2f0b250bded55
z42e47cd7b9a0e75356e30c48e4fea46cae76bde42564e8a72207f5c16a2e5f7b88a506221634b2
z107864583604ffc7e0a8f8c682af528360b678ef717834739939d650f6fee841e83c1730c27b50
zb9943b20480f2a93bc326d41baaf91f5235644dac034c36d100aa5113cd65dccf774197ab4be90
z353c6fe76588a3564bf47b8b9855871f2d0eb2b931c5ebfc04dcd217cc4f9aeb0bbf79129d2631
zf7f26a5b1d311457ee4ca1f93e917cd1e12a9b9a8968f9de2d75e92ff79f086a21ca90a0eea6c1
z95432da78632bd9191faa6d20b31329798e7101b0f3d08acd9c8d8e953109654225ee67e6eef1d
z512ef9adad8369eae7536e9715df0b580c51d5f7da685e99fbe611566d91feb12eee6ddcf2040a
z46c8e24297ab9808cec6d69ee561e37b6dc6da2ff6c8c98ddef167ffa062d7a72816f41627cb52
z8c9e2e38caa8ed209edafb97d7abcab5ea6702bbbbf52e54881c47082bdead025bc2b0f07c6072
z7dd69f24186e227facfe6db6f6b38b71814eb43b87d7b417cfdf672f22b13c5b20df2bb5b3db82
zd8b2d63f93120612b421dd307d96eee0ac54b01fdf58f55863597b270b05cdf40d263798e29ac0
zf3567b4454439ad57bc6ab4c405d7b5f8944495959c902f3b3a6e317af2af439985bc3ffbbe066
ze0dd586bd1149a79031535cfaa092fd020a6bbbc25d9577832600e096262339d9205128cd326f1
z52126710e2f7866edc46ece4266957f9e3006ff171525a100cacff115885f4f16c31813dab0cee
z7e674a7e57ff020b15db2e44ad5cdc10a55883094516cd8adbdaae9bae2276c2f7545fba58b6cf
zde4592092e890b4b416a4adeedba3d2bb76bffbc64d0c926f1f0b456c295d12084de055857d15a
z919507f117c2a5a7bb99263b8374b320f758b38ded0f244ced95e4de3ddadb694557a76dcf3b1b
z7ce6ce659c995d446547d9241e1b117fdf54c8d7353d1744870b33c67f99f09593ae0a2bb63b52
z49f0b6bbd6506640438abef4bf0deaf22a1f079b7118be7c6b1189a6447c4f7a9ea52d73868212
ze1eb3a871b1ed1878e4758133880bf5a551c7ae79ef677d65fae376fbf8170860f912562ea5d25
zd96c4d2c49e5aee76913a725f2776cac3d7146e398be4c152d4c9b39afc265b6ac5236dd597587
zc1c86625de256dab423c0825839b9e5255333acbe09442d49410bf072d2e47a8b09a4e6d23d7a5
zda3b4b738c4cd85d157c2c9ae7ac905d9b138f935fa98e09f0544b714b6b9d93a9fec46ab7743a
z198bdf5accdee70ddaacd93e5b3a4909d14b3c2e2e7b9120ac930df29b42337c156b57a31412d8
zcc79ebefeb0224f4c65d643ab1be77128fbb7826134d5d88b542e84f4d79cf6f0ee01ff636a5a3
z0ad53fd9008b52dbf53212fcf997b706bba69f47ec77761fb540d09b60d072326c5da91cf2ca13
z8d88e8231be73e98211eb2d43f5adad9ce4920e169ceca1cfeaab1d1e76bfbc808a862044eb34f
zc3e5939838cafb09c3b870171d24f70d84d378582464314850596a7bbcfd516e73b72ba3acfe09
zf93a0697224a4c5b04c4e9d140cf9fc557556c943807a9dbddccfebac7e031727034330b8d9e16
z510fd47e986931a9e00ae30de65b0650386075e5a06b2eda412fc9a32a28897b2d1c1297c8a298
z421b59e88282cd139529d3f5caf366cffc738d9a1b38f851c633e492da9c96d29c60a25d2c5014
zfac2aa5e081d646c8b1e0cab92043e2c6678407e042e3af97ee8e3511f2cbfad2bfece02cd0367
zd25d5d07a3aeb107ae9f51b6d093129235d90080bcc525f28c56b96ac1d6875d3d5d9dfdeb8248
z0c7233f48d09f9aebb344c43acd6acf0a5025e5818b2b03029ea8e149e2beb846c7d0142792cf5
ze9e742cba83d7cc860a314b2c929d14499ced828ee75396d808befd8039f12e8c493237ed0f351
zb6899d749690d21862c1604fd1651383abc85e99ed32af66da7b1eba291f4c332d93802fd8ccdc
zf8c61ec010eacb4f93397b810a1ae057309ecae3d0f659fd0e3088be4b400392eec56f5a22df7a
z9421b6eda324cdb350ac90abb7525dc6cf6e2ac7df241319746f2fb6668bc649b44bd07089f1b0
zea6ab970260df73558fc4244a47230fa22251488c042878d486cfaa4a9f7c8d6e7efe41a4909aa
z71901b62aabbe7e46e4cfd320d2c6a28f08ac807b65c3e59d1ae7c8913b113c3872e437c3fb822
z7732e300ad6cf16332672905b997b988fa8d6894bc1cadfae2af942e290a4b9c28d2dce14c334c
z895f4265c4dcae99c0d3ba4b846105665f0df7faff3a71cb01e1c7b154d2a93a379df242f3572d
zbd9f4732200302604880fec49d9765780e79f69e0bdf377e664db33af304de4d6e363db2ef8c4e
z34270584ccc68ca1ec3257158391b05ac15c325b90b13e6b6ab9aaa78018bc2bfbd52c3493960a
zd7c8022aa7da8f20c8df2bbabb93d19db1eabb1bb040195860b9c9c2529b2117d3b74e9135eaa1
zeb427e83c1b5971a1a0609acfcc8900cb985a362022bf5b447675f6a315bc76f465dbe826a356b
zc66071506666de400872dccd4c548f3347b71df0b389bcf6a8edc0c19f1e2b1208c1e1e96d89f8
zc3dcf2df7d1d6eb8c81442a396bdcdb607d4234c67374aad92edd8db52d625bbfdf08b2797d305
z3196a5b0569e8e50e89fae2527fe842198fb91b4671d9e970d498d3f05814c60b629d0d951f2ca
zaac40a45d6c3f230f26dcb93944df1d32600e8b433d04f3f42ba211669d832f22e54ba80b1b013
z350128fafbe197604d56b3eb89c3cb67357eea821011cbe468649873c8ca348c64e8083135cea1
z3c3476f47fe383417232491d84397f646fac57832b3def384841caebd0bfdcb815503253ac2499
z66370029e9e6c41ba4f20aa5a7f45b996dd477bb9e75eafc29216a1f5f321c6c9ec2515c589a82
z8ee5cdc73cb13376fe95f3e3d2fd79ee595fa2f96ff85fa24f0a1b5eca38f50bb3bd2faa881175
zc908f7f60b9db103f63b5ddc1912fa148e9fe47d3d20b31a7698fd6821db9b96e48840f88365fd
za5a6c5abd86d71c2bcbea61bb223ce65a16602dc293612d2b399921180e6266427b8e6867be64d
zd9291372310c616d6a96fa3d6a0135ca792333e3b0ba2168370551f3fdafc01a55dc47e71e9c16
z78cf5d101c1029471c45c6a447132393283b29d01087ab52ab756a3c09c403ac4ad6f968c25925
z40c906771f8f6dffbf52c02eabfb8dc040f1e034698dd6999dd7f40f0aa726c780f6f12537344b
z4b67b8aa59fd3952e4343fa0798e7b2c46790d8984fb19049e507f5b272afaa558b5ff12df1c7b
zb4e3d035d2ad061c51929c57a0b36222e142f8983e62a7f330e4d02b4fd6d02787a99c87863de7
ze876ebdfc7002b9b729a1025ea352f2fef842cafb66c190a4d10c02ca4b79578a9ea795ec124fd
z80bafaa92f959c640a157e92ab17dc7f7e973de5d291b555c172bd00f05bd36a6e0579290f26e1
z7d8d0888c8e9f13b8d58fe5ea9446d1bb255cb65a2fcbe7f4502122119aad70b2cd7c9b55e2f10
z2e0a3691c335d3f22595f6cce521b9f303a5a176c714720a666dbcb9b90a005c6c59d6a7b7333e
z3ea311327e67ab407bd72b76235599c5bfa5f06bd47b126dbef164e9c6147cc854530636540bb7
zfeb825b008c685acad88fe9d24a9f58206ef93b7307771d0f248275815d54de7726fe9a8970df0
zb78869da5bfecb6e3ebe72c6af2bc4390a879049574e2628d404208fb16865c8659561fc992c8f
z9d2d688213204c7951c2e191175a17fc39c7c7475a5c5d6fa1eebaf1d8f8ea4d32380e8b58c263
z225daa8fd5046315969e63df863d9182655259789e8d8796059c3ef24e49f6c7a9124dcd9aeee4
z7d7d0c5f54bf1fd9d9bee39c8e557ca6e5b1f7a0b7a595a2c9107458d479220f77131ad80898e9
z8f7a15d4f0c24ef133b0bf08f6dd8d3f2db3261433224a641520e3baec6a4c36008a5224a07d96
z9459549f55ad4b237bc8616745c9174e3db0c81a885343ea4d0047b6a0b062b07b7d5d741596a5
zbdcfc6234e2642562d9debfed1516a2963cb53c0156e9eb0ca3f13e67dd38f0f30c0708f705727
z90800653b6a78dab8a35f0eef91c11900a5b8447c453acf8d266cc46c7d014fff2d09a22c53a92
zb676d9554ddef3ee51988fa0a2bd573e63664aaf729f425a322f5282973c5d0ab2f14e3d0e8785
z8074d00a17131f2832ca4a8f657fedb9323ac234ccf404894604f97c2419be30bb8307191525c2
z925da9e9
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_value_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
