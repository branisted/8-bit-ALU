`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab30857016fc53a
za25afc8341302f0c829d94450c399b8ff9b0386c187cb854ee330605b7b59da379b1f26f488e1d
z36e675f0b1336408b3a1ad87d0723054f952fbefc8d5a33eaca6ef5be8f42bc59870a29a5cc9dd
z4fec09ce6e44cac279651402e7e1f590df88ce49ec26ab39f12b4a02855703c6f03b1e85c797d7
za357087d98e5b1f45502e45892e5823d6fa4b762932009620038c05d74efcea7c3fdb38901d620
z36515d0824367e48d1bc182335f158c262d396cada6b0ad58add4f945eee634c2dceadbfb5118e
z14969c29a743830a07124bfa78707f3952b96b0db7af7c9ff36f77137d8c490c4f79328328069e
zd7d5280e4f95742c9841340368b9764f0f80413adb175ecfbdf3c40716abca7b8cef6f7fe92ab9
z6bd2453f1aef7f7899c5365c5c83793cacc7795c269413f6cf0dabad14d40e9285afde8c01a47e
zb61893788ec5060288cabde8fb553f21b02eac61ab0b48ad3d54f4d1d76508b22f0c600861b5ce
zcb30ba708be817b1f50f59c0f6fce449203e7355c1be55b662fef3f92ba58243d81537761af8d6
ze27d7864d2dae99372b2b75bacdc0437a4f7e011d68c3487a89759e3625548fcc920ad06471ee7
z2d701aabf726859343208b0a543c73eeff8406febf277e3babff437ec820fb49d6b78e73bc2353
z884917487d35a6cd06d7d73ccff5f05355122888b886d1b7ae29679db6c9d2d7f218ac9728369e
z0ba3297b105b1781345d5dadc1077db50a0833d4730649f7637b2138ee147e4467e47d68c8e25b
z593a6bca87484aba5888b0d117862ed7c2676f9edaf1b7dff2a4c8c60dd9f44351e4f72dc5a0cc
z078e18bc1a3e16169dbe18fa92cf30976c736c34f1e53045f4ea0e07c779b0c89edd9128640419
za470c9548911d77ec74534902e23ed1fe0e26bb1c75a601bade4472cd66f6a9c1a514451027749
z3c93bf4c9c0335941b7fef7a1c7aedeae746dd2e714ffe233e9e081c98cb79e55bac3fb05f7c26
zced71ca7b5b51499355add111354f6456b1e98e25958d5c71dbb14058d120698d689d1f50a5605
za02ad7c57cbfc7c7db82fda688756bc64d7e0023dd49024f637f6c449375e0bfac80df91adf122
zf404ac492c6b75d7df921000659a850b755a85891c4128e6191a4d518976af372a779b7d8a9b8b
z0013eaff9247beda916c0bb4e0ea49ce8e9fbbe0d9e63237c715063ae268f5d8bb2b1f6dec0bf3
za0e3a465edca5bc93cd5be4879175db2100b0bbbd16557795d3dee8ee87a830b490d79f81310aa
zdda52bf79dab4a231976353cd0a46551df4bfb2a01e5c272700fb95f896ffc230a6555dfe8ecbf
z776162702794fc443fbe7651a5ca7fbf8d05a5e5309d9a1162ac6b89f2110fcf7b85ff85b1a8de
z13d31e038f801384c2cd5dfc8c7837395ef27a048f0b751dcd389f57fa1a1b39c7cd4b9aa87702
z8a951fd712f6d5d3b3be0e0510de2b0045fad1f1b8d2781a349f8aa32f6e671de94fd2ce56030b
z78d39f3b544bc9febc6e35e6649f0d656e61a57a35d36da8da51dbb0861fd53c2891e62d7a184a
z5e7d7a5ec135688b7f8b860f10cbf018aadf1e382b34b620ebb570311eff81235c83972dbad89a
z759d88c3e45075996649df88078ce4beb53b9cc07ba8e612c52d391b3c4a54f3cc0d12f9318a11
zcd6e7c0de7191f95276b2b78825ee9a0f06286a1fb3923238ba12002fc4a59ee7e88427e676c0f
z21d3afb0550a21ce51195f8b2c367b04bd490be197f95166ee3d624ec1b7ac280db8c59db795aa
zc8af9d3d52f3d939eeb0ac079dd7dba5c6fd011ed28e2f60b2faf88896663d03cf2aa8cedcf6c5
ze50cdf071dad163c3b1b947c14f4e7ccf8d1e14ab02e98e06a6df21398b795ee00b8866ef6d89e
zf772ccc0308845f51c2ab5e99a0d42d39bf23ead5842afc183d1016dee801463a09173edf75665
zc1de08db89bb184997707cf723c13751e65d8e5879778acc0585a5f6cb901e5695ebb14fc98183
z804696a0b88d95ce81c33a7edeff997c90a829dca42ed2336fcceebed25342500143bee4d58c50
zb9345bffd2fa417888a88bbbcdd1f0021bc686d5020391dd3906340ad00b786f1649b04bc4c476
zc97dfe0a92250063c00666d09bbda2309b2d7f87d2720190dca22120c2201c1cefdda6a9d17968
z5b6d7c7ae938c1c46ce22b6ac2fe7dc9317eac873d58e4faef3cafb134ec04a7ccc6799ad13ac0
z1fbc7b430b27a1881bfd26d0d9026402af951c80535a49caabb3970ab15e2b75b37efc53d0214e
zacacbb2a5b23cabea842190e22fdb74c8e252f6cce42f184877cc9712b903282be1d999c9cc0ac
z3d5075e490033947ff7a6a162d61aa71fba8d02f4ed23d007cfc46292e2daea23caed96926eab7
z124da6f503bb36bf2376de60e01f005377a56b40482b6c0ce27e250569d964de2e047fae7c44de
zce3d0e7e8741346aaba02c832851e3e84a30b922beb309497e6ef38f3fda6b175448a02143e311
ze0413e33530eb433580013b6e8cd4a3ee68a4a7544e3c7c4faf2c4108d7a19f41a5fe86a919516
zbd679f86ed3671418b56f6aee68db9913dbfbfacb5e536f01c5ae3803f8dcdfeced7b42ac77bbd
z70288d05319683c462f4f168225f388bca0872e4919f71297e17b8a04259088d4c9a347e20a2e5
zb993d6cc000a61d1f94c41e760f63611d830bdca37e149da05fd48f9f56ed2c2c1a2c0ec345140
z2aced68b6ebb6bcafd81abc278f08b9f3e3b7608b1c01cd89bb15147dd9e41545b5ab2b0a4f110
z822481460c3b0d525d912fdf79274e7086d9bcd5e1fd1d2e65cefe156fee090bb42514f130cd40
z6df9af2eef81f58b357c587de7b8b9d4a7fbef5b381059d2278e89fe6f722bde7871cde6bc0555
zc67240863578f2f1f3d57385d8cd83a5b63bcae9602509318b68e9933cd7d88cc9eefc76efb768
z59594916dd88f49f5c8a3e8ba9d9a2bfc0468f178a30352eb515b55b5842d7ccd94b4c23929dde
z1fcd69e635abf8e7ab1e79d9e24b0aa5f25633d7c8fbdbf0384e6438fccfcf5d2ae30789a660a7
z8b6385d250e5553a925783d5622db1919d341af327ef8ad914dee745f5cb37a3b6782c4ae4e7da
z6857cd550afaac8389bb3a2d1b492485b711cc0ee68e5162e25e0460dfab31135567d119885971
z52024bc1fb7b3f5eb91c2ccfff4fa836e7d08b4340f10997509a05804f450288737f4defd3bdfe
z9ad85c260dc10b1886427d10619f7a1d98441b218a55e26b45d6d5a3381bc8755e24593ff29ee6
z0077d5463b2a9473906fff5bcf8f42cabd354be2ea55a57fd4e34f3074d30ca52620362da0dbeb
z349e09d8ba56e4ff46c6e090d4c0c020aa18681d4d449b8a8331b8da661569278308f219d57f7a
z1cfedfee6e971057b59f7ae0cdc571d709daab94619fa09fa9ef804ba95daf5ce422a9b5c39c41
zbeefe559723271be59c23a8216d8d2666c3c5f1c796e1c604413603767f3fe63b55d584eae9b07
zc4b240a945224b0c7d952ac599af03c4b725c82d4f8bb776b809f114b4f77d860026962a58821f
zeb9858d91ec795716120bd224d6969a5fa671ecb62d8e9aac6c9e6ec58de6eca9918b4854c831b
z863b3bba4b9722b6e3a720e6ce2c4fcd7242a87b7621a0af648cc79bcaf1292a592061d2e33fdf
zef5564f5df8375ce8ecd1cd5ef59b6ac9dbafe5bd1ef177d3890de3b1323bd2cb08c2b20913036
z2a55262e86b80d1ac5b1575131cf939c59ee268d1fd5d4990e6bfdb3e70f681ab1fd364b218de9
z844553620fc92665351401dccc31e7682f54329238908a5b572cf57a99a41cf34a69dded7af652
z9d3a0e58bbbd388f436c6cab1115ae9972b254f6fb31529342197d0b8705e8082017ba6ba1ae84
z3d10f2362bf5f1c2e3d0750a0ccec1934b35754bfa531546910249af5c4adc5abde0ef52feb28e
z5d6d7d15d04633e4c283b26731d2fd378531028eccd97ba434c74e4ed80afee955a933410eaa1f
z9b263b2788865ce4e6fa531c1da62509b336d94ba1164267d188d83bc156ac55232c2894347e80
ze798dcdcd9a233a2aa002e32083fefce9c3b58dca56930a586f3532a712428efc3be5e63f57cb5
z888726a42d50b13bde88a09d01ceb43a9a1cfbdb00c3d975e6255e599373d06839d06fcfc55e7c
zcf27d0f356eaf88f23d53581e8853afe7fb22bdb129147177581a0394167e0da07a2179430219b
z965e51b3ce14bcf7ad81eda52780e83e9ad2983ed1f2d99db00fe2b72d72e853a841b6c0f8a985
z0408419f40fecda732d83a21db4acc7ac87ee5593ae828845de749a8e79a506053a53cd71818a3
z050cb2922a4ba8d3e1f7164c0152f18bd24d9ee7a030e8ad724d185c6705a74dcf8544e50d7850
za51e9dc48a275f2e28cdea1dd2be60cfa41042cd46d90528ab39743c7813c0ddbca181f758f8a6
z957b63baf233731c89e6b2c6d83c14eebd87546042ba6e40e7a2aec6f0b5e6e048504c5966b9d7
zb2982efc409c1b79ce52687b35f596c36e36c92142ffa21051f9d45245db6ea46c9c641d3e1a2c
zf8dcd9c3cd3b30fd80d4dec5eb561fd56d35394392a2cff21d8bc1110ac7ccc73a8f28a88df097
z992e24ef7de18ebcaf30b0d41d147b3d0af4f8511723b6ea8b9ed91232e32dea07ff4e27e0504c
z58392fdd79178ff48d5daecebf3bb0957195759bcc67e3de3fe77f9a83211aa4111402ade6325f
z390c2c178866c6dc738afbce5fcf8ce81d51e74f89a47c99a1db47b6550d1aab1768433afd9c2b
z22b9dd6f99708bbdb8c2591730c06b61e15e38cf53c6fe334889fa513565a9e3fe95c54da9bab9
z84be6ffffc3489fd6d64d3c3bd4e4d233edaf9e6acbb83272d4e5ae71ade43e9e93d623a6d2056
z436d7ceb4bc1fddfeeb766da774d7bb9558a3dacf0c5a8c55cbdf2b5e4fe99bc8db7c9346b462f
zedbb5db89497712da86adfd42d5f09e5750f1b0218ea55123c85e6bcb89788b6658c81ddeef8f8
z1b6d51f5db074b326f52b93504a721692b6d02d72e166f26ef0ed7adbb61c7c75254a4d6712432
z3017562bcd3978b623d1c2b84cab698834fd5d581468b26f8c5488e46f160b1d204bcdece11fb2
z41c126c7937ea2370643e61f80e708b4394b5f4d1c3bad96d7204919e2b304ef2a00b8059169de
za987de64268284790bed2ac88cc81b4d8d42225f0ba19df4d036b55ebbbdc9adfa2aa2aca4a4eb
zb859dd24d8c5610e04076ea891aad952977b62292f95eb02ff5d27f6d84befe60de434b86d69ea
z1b3e8c907516eb7349da1f9eea85ebd338dc720e8b794a619e38d895b692969ffe88fb553cc956
z3937f05e810c0bfda06c171ff41045cc604c287a9a95e0e4448c0ef73f65c0a49804606dbcff4f
zd3aad6d86657111a7929b6f7a9a642084450ac8296dd9a8ded2150a29ac40dde214a3e340281f4
z08fe1b916a037746e98b8c621e1dace2e8968f2ed4af40d8767be511546eaed26c649ae04b32ce
z5c8ef7a81d9361ccdb019bd374cf696367b8b01b560c88886876a9474040ce57ee9238c495644d
z73445202aec92f62737d2a273e691344451efec968c7302def3a861427df22349452eef6004ebe
zf37a85ac889e31b080465e4513858a50d1b9615b9789feefd97da51b297b3597047a7402884881
zeac40abdc846cebd262e8a659873790116d8026d7bc1c0a4679d83bb3a906567c006ff62a84de7
z8de578f6c60d297056cfed402aeeef6cd6dca891e021194b1263e53701ce28b4793e71f9b9fcc1
z2a8ef1de2b6a92f06cca3d1fd2cea54047485b6810d693e46412560d1ef0844d56b8ab5f3ce02a
z1d1b37a4e423caa59f974d6b37295af3e1a4de8bd703b75c7d03bd2cd0edf53a3465295a8fa986
z0cb6594081b883125ae36049b6de9368eee96cfe5944575412334a8e1fba6cf915c96dee8cc758
zcd0a55d053a5d0ea7dd8aa91d4d9e0c5cd7de5131a1d810201754bccd9296a8faa411667f17569
z974a20ee5654bade8ab04a4264cff63399706d66a65d5530cb522b58c8f855ea510fcf2aad5699
z69b638ab3ce8ac89bf557a2f32e8ffbf2b1694e504d407f023e8ba7a7b0e0f998f9f6a43503f27
z88f803cc3aad5ca9085d6131b3c2911b39879c3c81e3b736b9f6627a56f2425be4fa57b363bcbe
z6b952548cf92f4d3f65ca61bc9e165d5ce36c8685f7c90956ce7fefbfc3bd1e2e1ddfdf320afa0
zb9577a99bb264d0ec3c914fe14ad22f592ed1c8dd3f7ae3c4fdc84b82cc5729a3d868f575b9778
z6eb69f2e2b4d32abb255d516f11e0b2e31ac29b84e6ae2e71265014adfea13f199862253509f33
za5178805b16f99198576203d7ff72581e03b16e08fe0144ef9b9468b732084b1432eb4fc359309
z3a2af63d99c5c610de17295a8cc3e4be39808673667b6cf77d66de517096b3010f49c65210a360
zce4fd85df8a26e8fdf933ba24b75652bedff46e3858236b75ebe9c2ab21016fd79be6d5b17ee65
zab971ae76c0d04484ad63da918a409b1be9bd6b1ebe820e3556d6a6f21cb14df5951c120bb118e
zba2e8664a3eededa467282b7afa1996b3efdd48c6261956fe697bed84e85b66a4b35c0f88497e7
zc372877f81f428f97d84f6dcd8b21b6926cc6973d8f39a7a2eb8a0582f1b2e19f29f6781314b74
z772aa5775b20eb7a3000bcd68b8ee30aae2a22e78a0592e3323c80467e50d371f179342aea89bf
ze2b9b74cd293ae078711f56b0fc289bab01063a3da6ac62297168018bba21bbeef131d4d321e1b
z94a24f12455ff7c424a80de7593c78262e50a331cc8c4442e8a418b31c6f7634d6e3c7276aa1a8
z8bcdee181b180719866d68342a3a4de0359ddd54144eb423fb15643fcedf1e354804cf3ec526b2
zb74e953da54e536795f01df68dd5dafdf4768df739fc352bcd457844314188358784e6fb110faa
zf20c89d62426b1ef75689316b7a3277b0929a77426776a81d8a32440c67a7926abeb919f030402
z06d70ade63dd8ae9777bd1264fe3bc4b101db990fb48c07d4298f90ca2479e3503eab8c1949618
z1e8f6653f7eec210c73e0745997cab3253d76950135c03cace63c9c0ad4d7f4d4ba66a01350e95
z44c179f37c7e37d60530e65049f3823fd67b619f936a7a95c11ae773927d628db51a4f4e2b3843
z735e73d2138649c7c465061f66db2bf7ad3c7d9aad85877458f7f21a7d316f916ad3e680251b5a
z3c23445109092ad0ee525d7c8e8afd59f897696ed7e08c25a5a19495a64f91e60fe2f99329640b
z153c430fde334f44f72e166ecec559e3f0f84c64fd7afc7fb1c161bdcfbe897bd8a0ee4a94e606
z9c794af35ad59c10ce037acb6553e8a09249dc55b012f49eda3476498ad5943ab3baa132e9022b
z0851acfebd13d06a81e23159c2b08eeb9fd190a197bbe00929d7772025105d30b52be2656a33fb
zf66bdb857802fee3eddbc57519fc1583a594c7bc007511fa713aae2e452919115bda90b4ddf7c6
z94f3fe6223ba89289bbc611cab7db95ef187278343db4c176e4ea08c8291ff301dddc5724c226b
zb820e2ea623084f5969025a099ec967013946a01771f4b5371032cdf834574cde0cf62096a6ac0
zc79f1308ddf89dc2ad7847a509d7eb8c2e4ce78a7eb5715424eb450420d78b7e44517db46188ba
z160c210230620a723e65789d32faebb932a57c55c5e97f5848a822791c3933c30b52915836d467
z7c0b002af87b8191c4475ecf1a4bbfa6917819d8f7d245731f8bcb6f216635e17cd25932f96efa
z5f1b98f4f5465ab81fa32eb2362bda8ce7f414cd57775e02c0a867ea52da278316cc62f875bad0
zc12752f1ea3cdc0ac35122dc4dcf9c8002e7e6e695a51c6ea0a3c9168f8cecca8345af70acf6e6
z6b8dda6ca4b70741e844c593e05043a4cf72c18d3b71ba9263d5ae96f9a518652c5bd93eea4f92
zf5c7acbae4043471249de1040ac0ec6089ee3b9db9766c61c4824c54f679e1a6058c566913e6a6
zf588073eab0eb1e5b5155985813f7a507aae03b34ee01bfff6115de282772140c7e05c4b7eb299
z13fac8a39819912c05e6a4c3b6461f20cb05a8803207699040db8ababd124891728d8134a6e7fb
zccae7ff7b25b5fbd9cd0497419e06e5abf5a96a58625152b50bd153f6c398e05ec47631f6bb0d7
z76db04ae66b49c5637aebc5b242cd27114949538e231526e46951de63f2341158892d7beeb1cd8
z94bac4001234d24275e39eac04780e5e9e8eac57f08e294341c5622f6248ff0cb89a6e0b9c2540
z858dac54b1f341ea6f6d54703d896076a0faa9f087b5fff24c744704e936cc0659f07b1374cb3f
z04310ce90351b9846400ecc631bab92bb7ad81c7d3e96d948ed404d9a005d9278e3b4253e350bf
z00dff687c7b23915356d8ef0bbd95de802aedcc1b45ec82aef067fef41e5ea5b7e4cd48f812a43
z58c93440932410b93827707274d1302f3ac72c33b419c3395cc3ebb24b668702351235f40f32ec
z0fae04a2b1c020bd7c16fba3737eff85052d466fad090cd982402bd4aee9e87dc23f5cc7a27984
z91ac60b0dc0d26ef7608d5a5a2c88fc32286ff1999a29b1a6f7f3920357398b7746ab0cd12057f
z354496e90ac45edcd4884cfe3eabd86243cf08ebff9cb6ceaa79688a918d066f009111aa87ae94
za0e9ee8a44fe825a8aa8d25d41be5ddfdd651ad20b6475c4d5d314fdd3db63821fd3b116e40086
z180c00f4bf1e21072cb5aeee58e7132b48db8597fa9f79e7c4c57f54cab191831912b7cb83e14e
z8e7292db20a1bd3b828d715ddbfcf57f3c292d2bc1aa1c5d4454218c225a6591b533b1f50e3c10
z9d5fdc52abe64373c573303cd3d98008b566ae0145f9231b021b4c39655b095385c11c710e80e9
zd9cf89c3e70fe8cb6f1423097931150b58bde9be1b18c42ad527332f87ba4bd9b65c01540c7c4d
z226b5ddac5e82e1de272cec609b02c68582f5ee6b44635849d76c54d667b8ae43f4b64c749a71a
z96a16ea3e51be266c89de1254e97a4965854d7fcd30013df85770a9a32103937d31b6c8f4dfc6e
z1a6ca5db2fc5a9dffffe084395a3900e0b75037941c0888222fa9a8b37c5ac810be20d5c86537b
zf2e090007fc686c5fd321aa6a2673dff9311da015b79863515c4ac12992b92e8995f2077ca5b77
z0fadb41046036e10c6b14bd88a7019fd937492e7c2610dfeadfdc815ed28954b5cc337ebad6a76
zd1db9b7cd02fcc1a8dab031c982c085119c33998c585677ef0e08d015c7e7406142cb08a6b4958
z18576fc095af7d797ccad3071ec0d134d791f8611957587cb6177687cd70af5426ad1265fb103d
zc66561f2dd5e5403e0b4a1c6cce9b96b99639fe7c26e79a7781ecc53e6cf8bd94a7b686411314a
z280e574adfe78acd8270e50647c0a7b6755ea81e2da4f1c7aced3cea8aef340502b783b6ce3fc9
zbab57226fd1bfb6f47120ad5272c9004ee32542c83a0a6a72604e8e7db63608f8fd8b8582f3ca8
zfe467c011a8af84087084d5cbd1e35ccd3112acb903fc271beb4941aff93e597765ec5f94602aa
z2c2ed226fa90da135818dc57d3789541dec76bb30372c4a1149bee1223d100b0e3d52c1cc42c52
z70d8ee7d45f06b85e17275a68ef3169e38527479245b6b62ffe33df4c537a2c98ad85241cf9eb1
z7b7ee5a1caf7090ca1f280aca9fdaa1019e3dace2d7bcbf5fe55cd5dc7caa94020e71a2e6c439e
za98d65d170cc4481bd496684767f59380c24ae88bf3647c9958847c110b50b32d1b8d16d3b8dd7
z9c231457d69f04843e48076ffac10a9a4526d585da3758a20da9d37531f28d02945b7e6d524a62
z442a884215ade94fe0fe78f6cb4880fff950911fcadf43698253d7f51e7f3775a002cb4a226686
z6ce4a3daa951ff4f3d4dad986d6e2bde41299f68af5a89e28f94a671a0a09452fbe9f6d7079f73
zd8eb685774a0a485d98ccdc4362cdf72ebd9ba879be225daaa5d1e6a97a7d33b14298676afc649
z7df092fe9a396dbe648e900e7412faa1f292ff09f9948a289c0014aa5363e60ed6a5990cd632c1
z1a46871ee654eab0fb407813d9d980a95558e8f7695d207335984c5496f4e0145d3ebc20879aed
zc5401601bd812a150348165382b97152b6b4838e6659b4f99adf47a2b08e7ccc64ed0953b70ecb
za4498ddc8258eb1c1fc2e030a7f5f68e6ef76748a4471ec8a92cb97641e9f31ac3c87d376bc749
z4f23fbb4603e24e9440d124c589be31525144408fffdc16ccd9ee9f4c97dde2bf21051ddb982f4
z79172447f185cf40bf2c3b475ff4a4086fd00caca7d31fdaf7c268f3a98d1bba8faf778a7c5bfc
zdf37746ae01c1f036d1c2bb2301f97461a010c43ea723ba6e94e0ff64799d1dafe0aa7050dcfcb
zfe0c9a72c7c2524ad02d7a6c41e2d9519f27389a7d078911743a5bd7d72d7f5e9414fce3cf56a1
z3de603be0ff205370f91094524f5ae0e3f618e26864ce7f7a02b22ee93fea1e6f6e885d1d6047d
z62d167729a0779cc5af1b64f533d0b76ef1c5865060399068a8d263f0699c47469f4b862d87b6f
z07f915ee7df8847097621761b9a92cb0f5cd0f325dc88d051ef88d98a876b776157abe518fd4bf
zb08f353332de528ba0db29e99c1c166e1ce014f67b7809004a55dfa283f52891c27df985bf1bf8
zebfa62439a9f68564d3282445ebd1ffb314adb39a9eeac3aa9a07dc86b7c0ba2656bd476ef27a0
z7e7fcf1f5cfdb9ddbea090250099c73b1d5a5b8c1767df6042b0960bdf6c28fb025ffc77ce69c2
z0d3e25e5c1b1c8c497c2fd34e5be8e1933dd1edd1b610ba8277a7d5f07ce1d66e645f55c60d036
z603bfecd21ba14f0b37d8ddc95835651b659a552ee45ddeabd9fde79177d58edbf4dd608b84994
z178838701a61984c1db15a1e11852e03d6da10ee71113946d0dc720c357e8288c438284c7581e0
z35ef606dbf8f43212975f8aae5c851bb91f0df4aac3f2da78f7e809fb5ce1c42985bd3ac232068
zfba8e933ba78a84b18095dc05fe41e19288dee570d8515ec3c117f8ca54c0a6826c872d265f44d
z444c8b28315380f31aeba302db1d107777061ae36fe1fd09bdfb8c6091feb616266a7eff37d20c
z26e4dea1dc8ca88fd6e0af5f04e4b3cb706ac2466cba153af145f5c775e6d8116ffde05401fb8d
ze624d2dde598e13e99bb45c8432f3b2b4fc2955d05deaaae36123601babf3dbd25a9aad9499ea5
za9f1c76b48789c7b6dc52cf9c11092dd5978e11147895ef26f065dc55a642e00047bda0c6cdc48
zdce64eb98529f97233e732becc563b429ad14f689f9eae5ab6024af80c96144adf130ad2801a49
zdeaa4ae7a0eef897318e8704cf3b152b13e2786c0ea9cee723f973dac0e1732a39a75b0a250586
z2cb94d0fce7aeda469d5e863b720c498b286048600e41bef8249c70542b08dee27f3182b0c3e38
zaf4f21ecc1e424e04b2e9bf11fcf86a564f3d0706ee2f89fb00005f97377d7866efe918240e84c
zf18d51354d9a1572bd131da562c15a365b03011cf69a59834b39ab9dc2d37b685daaf8c9141116
zd963350d21c31c3b8118b0377e12cb5f7bf8d4d667793581193fcebdf8a240f934f4135bffb3be
z90ddba3e269211963e6549a1d2aac456b762e9fee9dd9f0fc47c8fcfad799909d7ae387755144f
zf71d8df6eb663237a1899dedcb0fa9675d7fe5a8dcc48c36fe7b8d84e394b4f0a858b9080ba617
z73fb84f3e304e06f68d367d98a2affd03638cf66dada4f27eddb7d1dc05a0c8f3c99b79b3cf800
z2c3d7e15bf6d0390e6a7297be625ab09e4c2cd4bd6a1f600f9afe9f1ec2ad69cb9678991121df6
zd69dedceb6b1022d7d75e84717aa9afbec50c6dfb05050f5884f597b754781237f628c512ad393
zc5c64e3234e46457b2338ec76b804d5858e3feddeb04697372e8024cbcc152c9fc4bbf85cec1f7
z8f0c9e71b424bada72d504edd5e2cc648098dfb042c5966f87f517dc88bd5b1f5d590d0a7a0e29
z24f67ff690502ad0c0f0757dd8a372e854245daa4fc24734fc12c25a6f553af052318ae8a90ab2
z6e1ef2e4d4216f402976533cf32655b78fe76510230282e3f97ff1e6c98a6c80254444d96d6ab7
z6838dc94ad25540d680019d2be2a878cf88d4ebafeb3e05c312d01af54f792f57ea0b2f786551d
z5e5ec0aeca18bcd25d9514c13313b12895c57bed965615f66484b7031785e9ad32015f2aed6913
zee0193746f4d39c089e2bd945830cf6ee632a6fb864c8373e9cde63d905d886eef4fe36a41a307
z8572b4170ecbebbd81614af8542d398c68aa4240646f710fa05417abc688daabf8e6eb2427aae9
zea9bdb31ac27db8f3494afb017ae25220d54502e403642781907066ab008bd56a08fd2334d6e7e
z05a214433674b423ef61b6408cf1a823ff4ae8dba0a50b9a62b10cd0abc67d2ea17268094693cb
zbb3f19c9d7211875d69ffe61704b3288c0c520cf99ade5b24b610ac38c2bbd63d4ef0d89650e18
zc3f8c084329d3ffc560981a5d0ea223f23e52ed2d898a8185e1ebb57acf2fdc1c3a09497d0c5e2
z1cf3908e96f8f4968107e43d5d88c4bceb7210ecf89e134e3877e3684fc5af1e3748f76003a04d
z5464e9dbe32cd996324aac670ae67120fd6efaa922bf5eb68a83b00bdae02d9708940f7130df90
z8cbd3854318ec46b5e53a556c1136bd21bd0610d6bea8aed0801713d3f9e2704b233a6724af69b
zee94d5d91105980be6c969524ab7997e3c3beecc265ba4248fc528d9ba80f919d79d198012fa50
zd04b2992ed15bde84500905c58fa343c09e3f1c9e033e776dd135cd06f523a0bc95ed2bb1c90c9
zb743af5f446114c5c8704d7b84b7c2fd222c6798c9eb7a0e553bed30430d263bde75ace22c4660
z00f4ab06ec6136f4e460f90d716a1f49cce1ed6d7f4ebd12d92c1eaf1443f329e6661ae58bc768
z6339d53ff53fc414a9b47fed680e3b09fac95b5870fb1833b981e44bd690f35b87bec5821af857
zfc9c77d712b22530a0bb7bdb73bc50ee4a4d3ec5fe90a3e0f9452766e9e4dba88905574400c18d
zdb4f136b016547fc75015557c4cff1702578852e844569274e6c081ff2c8932586473c6deabc6c
z11a9ff7b43e4540a9b0e6408834f2123b8412bde04532f1c21b5bba5b194bcff84467967bd49f0
z5ade7c58c8571e782f6db361c50ea4f6bacab34a0df64add65e4946d0d3fc624c0d175332dccb9
zc30f8f99a2bc3090db9ceed2954dd01612512952055f8c160aee7b7e1a881eea1654dd5a692724
z11529d2d9cc0bd2a88f916207273f4681833000853939c4e2526bba931d5fa5975ae756e01dc4c
zaca22049b891cae9c16763eb33d4c1f1f3861b997168c33c8990fa2324d8eaafc79b7eaa32619e
zfe054832a385a75f4cac7e02f1f6fd4599f1d2834697a73d9b0b9cfcfb966b8a87d669341ad72e
z7b8f1ac438a509a733ccc2fb9af6e3e388fa9d3f5b902bf25824fd34470b4c51c29f0df328ede0
z839ac0d808474769944e15b752ee32b3ebc426623a0fc1e695c4fb10c00339ec935a5840c95dda
zc435a601eaedb1de8ef2143a73f0cab13845cd907fb7d73c625104e98b782cb6e1b4cfc1f123d7
z674a2d1ec9e1dd8355b56dec46362e03f4b560df9d6cc60fa5f0463e4cea78699e2caf9fe4e174
zfefae0c78ad005d87fb16270d1e932e9ff865d54c174f4405237da90447e6d266044789856046a
z1823b64706c932b65e9e6cef4ea9d12becacbe0f66a83fa9a9ae6f0a07c9cc202712ee50ef03cf
za039e3ab5e9ad4aa2f6890f08158cc0fa36b44e2146680df58878fe8dcdd5bb823b503f627bd91
za9d3d93956283ce6f55891240f3876d450ce63d6cf719d73de81ce50e918fe7c09b86ac65b3742
ze5f35e085f302511d6203e5259ae7e5f120ab62f6a27b65ec49137303b959e9dd847dcb796fb15
z223ce125e519ddfc807ca899456ed57253a9e0e9071dc457becaeb30a3089aebb5e33d9c887ac5
zfa6050477738c2c437c23497d44e83db4a803cc6832006eddd865e00ecc8f7185b9d7906c2ea3e
zddaa3125d91179974ffe6df3e6a3754ef9533825d540d0d34e5257728fd9deb92baa92b39fe596
ze99b615b05fc858afeb7c0992e8e90a997705c2bf46abf6ace079df4356bcfeeda51362a934561
za5d45913f19e860f1b5e7f2e1d5f080c61b70af0e144fb74d759bc252bee4850fd202be1744d19
zb1170ff7254a3fe114b3754cffc44adf83083c28aede40868880391f3a22f7d3bfbbc20121b407
zc175664fc7f6b13330959f2dfb0f7fbc29caebe692666ad8752bbca79e33bc03a46dd8d463082c
zdbadfa2ea5abffe779dcecf9597f2d3c13b31155ed569b7d0c0e58f4305905140e434e5b94e19c
z3861c8b379ff11bc3f754b80cf3727f4fd084a6bd6d638303ba5786a7940e6409997849253f15f
zbd27515d2f0751fefdd0b297805d11eb9af660831d6907cac2c5daa4d6fb1b90d92db3f6821fa0
z561aa2c0b395658477788be605b15f8463b82614ccf3ec3d0343e9cd42cd3cae762a3595711640
z1339f5ac17543f5293a153111e080df1deb9ce19bcec442509cbc40cfc7c2d49e23b62d6a0ebd7
zeb95906d51da7a02b8326d9eec4c61ed87b1aaeb72985791ee17325745e0ad853e7cfc924a4cee
za013b05c6414cbb99e5b22d5eb4f190e1e96a6fe267f98dda0a8ad76749527642e58ec37cfa494
z7d1f7138d2bdb0af69863a1c5771686c43e62bf52d7bbed0932d7732f1adcaaf2ff88778911293
z1fb54918901c58d02ad69b949d97b253b038c25795d5fd679641cd57b72c2b6635560b457fb85f
z6c8147ed81bfe39ab103d19a2f169bd85a899c25c9e43e2ef589ccbbc4d4424fe22050c55f8918
z8cf9410a4826dd4de8f7b4b5b16ff61a9662d893cd8adb5ab44d0dba1ad3abefdeef6599df1f67
zca6af5b1df40ebcfd29373c2d48639c3ffab9a2ae27bb78802be3607417f82d3fe8878d22ff1ec
za1e7a506ab41e575c7ab47a263c2aefcd15142b1881d4fe8526882f542f4bc789f628f22e1c78d
zd7afe43cbc829c5f089d14b28e144b3135309f324e620d95a1f768386f61499c4cb87da2fd8624
zecc42c441f36b909af3e3c553136d67fb2b01b86192b1a5973c48355d5100fdd6c7d1624ac2756
z70776616ecbeb258b81c267d628f839fce005b7f64d706b879a2f8b2d059e1ff75f60345e621c2
zbed826e4d9bd9993b1d81631815eed4c4e4ede7d29b03038ef7e1185b2e39b0c622375e67c3a83
zbdeede4fdccfd7484cf7c8275532659459d6fd8da446c6b06c31ae33311a12b644bd957b2becb5
z31b4ad5209337fbb1e8ca8e85a0ba3f9f6d242d8a32f32059387a48e78743eb14b6e01c8952125
z2a143c4693c5d614a92fbf935cd1a44102d3aa263e6c80c49ef17bbfbe8d451d45fc22f1528fb9
zb8509cc3d9b9a0a5fff01e6f05f7c01dbf03b6a912cab87a41808916f068624dab5a393edebed3
z098139f7a6f6ae4369c1207f54d41d2194c10799e2988ce5fe5d8e06b0060839bb3baa08aa39b9
z84e467b23c6e6f34cfe740d71fe7b4fabecca5dd6ccb48b7f9fae7d42d1a779e2a05553a1f4578
z0c76e34143610df2c287f3c318c616344910845d5cfe451a10b7785e9be0b08b5a254a02809cfe
za7fa2dec44dfa81a6006c8d84c5e3943cd650657f025cb0d74370df508cfa8586a403355f9a615
ze75c8ab617b5db0110e720c9886bca2aa127655f638049ab652d7effd0a27b0b403c167dd62f42
zb9c697938593ec828db31b598f48fa4347313fae427243c8d7128ddaaeeb56a74b18ce52785ff6
z4ee20f8157cd914363d084b221feea2cbda0404ccdb9ccedc91552f98795403946234ace5082e1
z0da0ba76199078bd0e3125f19430ae58e419fd25618daf013ff294c72d8fd40cbd07ff404d3b93
z1a29052368c145502b91f4fe19e083f24b47ad6a207a2216e57a3841f4e3cd6df3fda57457bca1
zcd51e37528b4d17e00cab10689cdce7e248702a0f9d2536d772f1715ac04d89cc3f6469720cb2f
z8750d361fae0f74a29ef2ea278034bc8011524c65d5722010fe772a3084f2994638120497d849c
zced8554db338083e7da830a9609cedf2e28689d1eb4add66566da01af28b6200abddc26de9d655
z249993e9c69312b6185d0d1b2c861312344764d23ade4ec80738170d024ebbe5581603cc6d5509
z537fb104ab62a1e4e09ca00e90a5c92033e0172af21486bd8113dbf4038094e3ee5fa83ca3b6f7
z3da7257267f4392c3ffa5c7df849aa8ab740c6d8b5433a7d6559447f0f712e197521440e69e014
z39fb4ac76b00da22d2c64221e9cc183b796b11ecb90bde46cc7130577e06c2e06e03133f727973
zce05beffca03d19cdc939db95b85095c5c8b4bcc2d1dfd1e39cb360a16492d0afade3484162d62
z14bf82570039dbf2f52cd31c8c8c88929d3da03991f48b49f42c1fe689cb4eb97133d35d570103
za7975c1d3692c38f2e5e9ebcaeafc3a71ad8ae8812449d4103e7de72f88f0025a29b856225b07e
z7b937fbd9c3e83d1e92286ee2a67d7677440abf74deff54fce3fb85ecb1d9fe8a7b3da35b5e11b
z6f593bf5bcca589cb2f13fc0832ddce0979bce02b32c6d82e2c4bf314d8b019282023fa6fc566a
z3a4a47f0b9b4bac45247c4319e11ce8562f9078ea31aeab2e26166ba7044acca663ec5cee62763
zcfa4bd6a5444908d1627d4b4d1f4d6ea583b63166a04fbaf2f0a8f4e237769e6532d7bd6c54a83
z4512cad736a443c2f0fb2e24249493c706a7f2479ab1bf92de405d61d926ca4f14c727717bfd53
z589feb30b112fe0204fb9cdcdbfdf3eba9be45d2f84057a2b39f2d51f8a5890e06b6cd2bbb4a84
z66a70066993c3b648a26362d572db436d31445ae2cbe006dcd4428a3d45358c8b2e54dc3d2f7cc
z0adbf8815851cb006dcd7a96ac72ca163098f2ab95b8e497eff2cf68552dd8c8436bd9606cf129
z81ba0b18c16dbfcbd0b669ac9c274a8064cc20413a0d19a7788f6454fc82b1913a75f356be0b58
z77dbf50611b5a62d469378a1707bc547c92d8d9057727b7f79bf02d26ac9ac3f9c7bdf55833f91
zaa8a7d4e692b9bd27665d7bf6044531f660b3a57e2f7c3c6862a1767aa8caf56343ef7f43b5d0a
zfeeef784f12bb6a078ea2c7e8868b68c7d937a299c12ce7869255099d15beb0ddd479e69ef0945
z326240d7dad045bf11e9954e14bc5114712b0a8bfc7ba3bfb5f864dc501142bb10de65c74883f9
za61de3e20477766fe3cd7f758ed90421f09e3a75ef94ce6d6007ac090fb5007ef1e129ed5dfb3f
z379d7cece8e09a5f1df22823917fea7a200205bbc94392e562beca973e80e977efc3934cb66d9e
zf561f61ff3d5c1081236aa70b6dbe59a7dcf2ae3d88d1f90543d9d554c8fc09c8f20441a6f4db6
z9c57fc0cc9f4ff8b33d613d0b4e7e3d23cff49612644ec870e88dedf728dca5751a820eccc61b1
zb7861bb272457d2d4464b20ae085fa7ab49a0f069c6fd151664344919995f2fcc10773119ccf9b
z9051eacd1d907e60d842c370879db0f4f13c2f367af242ac3932694a1d38105f7e0e34dcf17c8d
z8df72d1566f21e97c7fb5bdc5bc09eda8945e760ac903de8d418743863a7842e4a6ab46e3bffeb
ze391aaf9170245267107f6972cceecefcb9cf26c88737d4a4097cc957fcbb69fff3a063ef1b9cf
zd5d148999335445b950903684bfdb9f5ab0d6d378d1d8098e3bef7d9b72dcfaceececf82b1f899
z1257128bf02c4c6ccbb3b7e8efea442db23e2c3c4eca787731e8ecfc8066b5d6c3e24a0271d0d6
z1d3b5464d87d4c0a313637271685e788d3447f7b91e69168336ec397ce77823c7c9df8457db0f5
z58ef984f508823480b3f6887765c64cc1d44736e512fcc571f2ba93dc5656ce671436ef704d0ae
z46ba09fb4a34ab988fab29fb17a4e5357780f58a941193b79ac95c91079b606dba30c376890f31
ze2d5c7334141a84b2d934c26fc22a132a7f17091fed4c820493ede3e3b7e018017e0d7c8f1080c
z4d1bd5a677947c92c66177b0b1b6f6801387ba674b58f15717723e8de6386a2e73ad3479f17b46
za08cd3135851ea5cc7478a393f04900221ed3932aa0b7f55755138a1895108e0dd55417e68cc10
z57c33db9d60d25dc1e0e4b51bd72aa7fa14b49e5a9786b4eb8115fccb34abebbd85ed8e7d510e8
z8116a423d34ef3485b903adcc682b66b62514db712ce8cc2ec580d5b6d5040410823615346e396
z651a10d384674a65e9eb27910b6986f6424cdc11db9c4919015fc1f4acd9e2b49fd3fe13c7d7d9
zac6cc5ff3d8e95ca702157f077260e8125a8ee693cfd21fc0880b6dd03a60f13ef07d3fa5d6617
z23e4c4cbc205731f824a1da3df7ad12c19f4ccaf323a66a11719c3bacae324113a9f216766e144
zd45a3586c26d5953c62df16d6ca3a99a19d549d655bc627bd85422c66545cead608b90aa9c7271
za80f40cae14d91ea0eaabab9537c6b1b60f78068696949be485075e3f5cae40349ddcc7d1bccfc
z75d124f93590f21cab120226cf2c9894115f96ec7e6e92bf6bb10d6f01eba1651b0ce6ef76255d
zf4b15491f7a75201a5ba2e9d2078593625ef779a76bebd15c0c8a2b05fab60aeb9cc8b6f11f699
zecb0c1427098e21b6ec217acbbe2ff7816fa88bec05de1f90dae8afdd8e2a382047c22cc1b3690
za762f61aa9786fdb40f52e1cd1562c1a0e02ffe43c5461855b598e5404dd8ab9991402d19631e3
z7c6b0c28105a47891013d7123a1ce74c9d066143aa9bc38f8753efb2fcb34b70fc4c053d19f64b
z0c4ecbaac558aac461655363be660f785fe4764235e65696e629a7ada97865ef5d546e4e5e4138
zaf372ef4517bc4e4c147fd08783a2d504f61bd3090c502842abb6d2d31feeb27512812ed2584dc
z3db4c5124914e63cf95579a0023bcb501aa139c36732b7d91df429d460c39574258ff0a24c9256
z9773d8486b8aaa455e7db518489f8a0140b85d2e27ab9e208ea8ffc588cd2835c8de73b54ffafa
zc22c2c00a96f97395e1b5e2832b70e8affbdc1c3a2df10e616d684abf86f79951751251e2b60e4
z8e89382e2bdec5d5aa960d0e661f7dcda3755f19ba33f3e3785ca6e26ad35e9da4e22c4343106b
z375b1cd1ad9a4b7e95905eec869eb9559a659e7332679a7f8ad60106546307f58a2b0b2283ae46
z5e236a2dde8e8690050a3e41009d96bc17efcf840b64a28affb5f94ec973b7f11ead08330ef90a
z57205735d79fdde6946aab57a484106df72e2ace6a3148c816ba92ac9949ad11e07700f7c68995
z72713e4aa9642c06f6fa43f6a50dd913070337eba91a6861dcb6e8620239af1b99f6e2ce5e1727
z3b3ab871e964684703703ee15d3a7ebfbad31969a8ee7a74c1ccd6c4f10b61f8919dfd88c4cd0d
zf26d3f86e2bc2ff1ffb159cd7fed9f1e3dace2633419ee2767d67a119475424449a5acec55b42f
z81d60f5fa92820a35ea93032905a29529f1ae5feb7df945f85849395d4ba52fa4c109130202375
z5b5ba024a288beb7f30d4b59842b7fedb2ccc0caf61bbd7aa8bae55b502f209541672795f7f814
z11321ab25e3c5eb7a65ee8e5ed62ca9d1df444781f6f65f628fb01d62244e67ab61bdf4c70d55d
z8e37233cfee197929e0d4962354a5dfb3068b401cf838fc44f980d33bbd2ffbde2238e26774574
zcbb137b4de4756213ac43e9d1f8fb85702c6e4827d560ab60521c03c7deec7e81cd3ef5c13998f
z5592c2fc090726777a1f90dd722d14d6071f117253106769e5fe05a1f2914996c4f841244874c9
zeffe332689c2b9e27273d4aa12dcbefe6220dcbaeb90b47955b5f0b830ac0550005c84194c4abf
zf0fd4f26c5e0e005792da4ed373f96fa2406bec4a9a6c9c5f7b35fc689f0712d8c8329d4b2ad8f
z31ecfec1076db8542731cb4ab1d6317205aec70311c0f226667e80644f46c3efe0f1efcb65e21f
zcdfc125abd96d3a9f421d98d67215171a47f95c2753c5cc8da4cfbeff84a4ac81692a8bae7a675
zc83593905bcb5f8127a99c1ac25889c4911d1f07c83a94d9c94b5931dcc0b86e3892efbc524108
z0e31e5c3c657b2dd857b412f1a5b90d7f5b9f965db4b589172ed753ff1a5ba834677343b3920fc
z3b5f1d3846850bf12944f522c71142456a47914beebcfea21341e31ba90a81ba6a0c9ddd7aa079
ze06e037cbb446d67f430bd5aac331c513c6a593018ef8eda07814e9937f3f41312d267c4b7f267
z129708513c479d90156ffd7dbc1eff2ebe2489830b5ae7dcdcd4269a91a79a099439bee1d93c22
zc49bc0bd93782f908440837a68aa7ac0e06211664ce93a4001689e1bac15583f531b49b94cf961
ze5cd3dfdb29f0a3a9f0d841092f33c3a4547f8145d6b5dc8424064f27e9b4e3ac61d307d7987ea
z55d2ac515d3d2b185c1ae3409039f27fc254a57bfa02c68f46e3426ddb02c9b713103ba4a59995
z34a83a5dd5d381345c8a2e48f2d4440f3f3990e0df809c93c0df6d84e90307809f007f9ca4a390
zf92dbd012fc3b237256805945d70df4d8f2897a1746f3f7b121eef1736006e7d37eab0787a281a
z0320916b540bdfa26437109ec10c2fab5074645f889c8a3d1c09051962dc7e4631cd32b322bedb
z653442e9e3ff3f27687976f84c060d4fc76af19122c75be94241ac8f99d78813557b7d85604154
zc6ebf9010903d9fb802f6ab5e6330421735ce72fd7eca0f609298b785b7f2478032187bb3850a0
z4841a06719d7728024aaeb13b8a0f1bf9216b39ee4a9bcfa5d642518d142fe40867029363c9f21
ze47fd5c306893cd71e1614d2065e4fb5ae5c43132a4a6ddb2d603ef30ad32409f6b2024ac630c3
z214d8b98cbad3a5a9cdfb97abefa8f6f0161cc4f59c6211a6c38e9123181874d4fe69536dd2c96
z32e52541653485c6cebadcc74f0a35f75caf234b1e91623ce9b4cf4b46b9500494e0dba74e3ff2
zb48cb293cf10eac0ea2882e8ebdfd2e2cebf9cf5a452fed2541802be0bf8f71b4661fe3d1d2ece
z0d4e954464c906f3976d380f14e6b9a3887259bbc395c964a8390d067378d9f463977d2a293629
zaef5ac159e4933ffb0ce661ef182f108a6c62f9e05c27b628f3f4b586367440a0a47082b97a106
z2de78a782555037645da6186e495edf62f3fe0c9d75e5a4f5b8dd1fee56b4c24518e72cb9033db
zdface858a97a60295319a7cb329d6887ad561640e67972d798559e134affc6679f2ddc39229b3f
z43ebd429b90f97a1f913c57b440d57e551a4a5584c7bcba86aae2e7a0b419c3ec140b1d8ad11e1
zc5cb6f254d4dc785f9543315b152038fc32d7e3a73b813706ac99106bafe821f0f072e6a7daec5
zf108e59668d909083280ad3dc6f7ecb79355f1fcb71bb7dc13ed8a51f5b5e95e0c71b1cbfa5d03
ze675d5cc9b753d219d2c8785d2b5a59a2282bf8b35c2ee0e78f75980e2b4156b73a9b58633262f
zac26979919879ccfd350d4186d7b80d6fbe57f5fcc535a597ec67cb797dfda8e93a9f47d0b23b4
z105b20c9f916e99bb0bc7ba81c628475868ed7529d8c9a79de919b020adfafad5b2ec504788983
z844e129866e0de8d7f9a4b5d09a80ccd410cf4c14c8256163f5e42bc9be06940591897a6492003
z3dbca5a39678f193939541202aafcf9db09149f7970e10ea16556b7735acaee03bb90f9fcd133f
z13bb547ea2d51eee7682bc2c1e73ebc43162253ed5186ee38b0892302be1f6cd2734058b0b494d
z02237ad8448c1e165c52a787d4be340ad163f4955be0f25752b888271af401ad4dd9d4401eb2f3
z0c18c7793c2897300af3e5cd2180bf140ac92327faee43c8e3507b339124d6fb1adc9b415161bd
z91786a01059e2ae0b29e5f66ac639e9f102304e8276b6b17f569d0f065270024fd269cea17d737
z49a6aa7ebb1f3836b3cf577728d9a8d81db8da8a1c1d184d6ff17f5706fe8699e76fcbd6d12de8
ze25e23696811bd6e4a4055adcc88368a86b43b4b82c9f232848b986cb6b97fccc6f455093df4b1
z39bb7b126b81aeb4714c04c7201b4e2456c6c2d21abdb398a1582d256d7f0b83c0ecb470bfdd7c
z2ee7bcc3ebecf99b96760c34815016859cca7dd71f54a27de936184581a3f4dca56e202a08d132
zb3cba15ee0389bb94b7002556f0a363e3918a8761a938d469e10748ea23a0c790f0c0ebde04b77
z0aa86f4c66e47447b41d586ecdcebe2239c1e7dbc95a324ddd2b6919dc31de8f8a202df116f204
zbdbae10267b8322c50415b43a803b645e80a8b3574825a1309807c7a7ab469567da1c36d4c8b45
z38f6aac8fbc2020e7ccd69a588c1a03c24cf32afa4a9a540d8826f0b394673be97d0bb7002ab4f
z3ac2bfe40bbe9484201b15bf7b983e6897974adaa79390bbfda95ffdb38224fd8818d3f7621cd7
ze8bf644ea5c3c5b9c91dc8c367441f3d29f7158fc7673ff8955bd3cd936fb1780a9f32a484cc9d
z33b6855fec21872ab26707e7ee12e57cb5c2067530c290f804001e080f3ebd317a5420294033d1
z7749d8e708a62c3108bf27c346d86b0b5237635ca628ad1fa55b69428c0d473bbf967d9a382ca1
z43c9ef3d3047023c505ad0862ed3b1d1a04ebaf88391131841bf10a14f578479c248ad914ede16
z5e8340a6787a14a8060498044b7e084a366c92014bc177bff1c313eaf46e9b4b316964535cfde9
zb2293039d528586a428a19b936158b56703835caebb5e775be2d39b2279eef7fd9c65c03d3d265
z6c8326ec198ab1952e06b77e34f63c90f0d96a6e07db2b57f802e62de99020c45302df4393cfc7
z8f6fdd6c423a79863c3a9bd7c1b9afe1af9e886bffd9eeb2558da92c562614c0acc0b7d413cbb2
z313abd0ccc3dac4b93123c51c36f58e9ca21afb3911d7e9b771c3b93bdd116c474453c11835660
z190cc5e7c7a4ca5c3aa9de9328327e9ae7cbb8a4d6fb8ee5a359f001e7bd1c36ac961ade0aabfd
z2ae3e09f6f78183160f054d1182c0941350fd9a7c3d1d1ae1c9fe25afc59e36ff9ddfd4370ab84
z1c0de143ad3d101938ad822e8580a30537ef968ba21dcd58442f9b8f786af15108ae82e1d8c1d1
zf089ee05f012523a74b1aabf2e32718867bf0df76097132e5ab69db83b7c71a0b49b532e885366
z628ae695435c7076f67f9f68f9df19a8f664b6db379090943e8cedd85a36e28a22d588c7bdd2ab
zfa08a252a286b0e24b27604a8684a3aad8000d1d7b48d32098f486a7ff8868fd10c0e75510a0a1
z24cb193bb6860be5242a7c81f2ea916d9dd81b981b74faacdf3770df8c02944b49557d9ce8357a
z325239f53e25aa4c0229304297518d78f4884da766d75f5719ff62e9b91d733fe55a08451f4d8e
z3cbc78d199a24a27e45e5cfbf6e4326f235f8648df923afd8271b9e1b42d9023e5e734f05b6770
zea70c301da8a3b8cafee612d3e7fd188197093a75427ed256a35ebd1b9efefce4dda4a37ef718d
z31bf81be48b77ddf9c9a2817c3c2e141db7222e69687ae4da1204bd8396c9981da69f7c6f17c3d
z366781ddbef9fb8f7bd8f1adf55b311821d8df30411bc229b58f949db7548a775fa5430df67076
z3ea3a7ce00f46c3f9a15d677fcf56b13d7a6c947700aad3a00ff568f0f0bd0e465952ebb45cdb1
z95c49e073180457895f2884720b2b5eb5a5cf6f832d112b1d3dca3f5cd6f119e3011d11aae7b04
za635eac109590ceab13b96c9b2db8da7c7ba0f998e745b6a8e4833f7fc7c1671dec3a559403038
zc17121c287027aeb88ddc1f18ef7cafe7c66539584f8b887c49d712ff794e74627432ecb2fbe70
zdbc4ab09379b30bcc8ec128b50a12dcdfd9567ec4cd5d92bf300c78f0a42d8633a9c5c57e0b242
z42595a3a8c2e3dc93d8d6cc6fce30bcbf1f929015c8a0d830906690772bc0fa85b2ef5d929f03b
zc14549f2368dbfb81c4bf3131959923bcf2a76e9172d3bf8746bcf0c3db89bf31526fae8b4c19b
z62488feb9506d01a6a374295b0ba398ff4857fe68f6b7eba71c711d2ae6f53c6c36346f76db5ca
zab1a585778065e9cdb3257c25f7116e7c438a443dacb7c02bbf556a427398a1e089e2ce16ee3d8
z4a6e091fb460e0a74f899ecb27c3d6bb6657e13519a8c20193e9055b8fb5452b185167d1ab3b4d
ze056bfae00ebb8f55653b6305a8b673caa9228ab74f48a31d82bc08ed0f1811b7a3e24fbd8e45e
z380c9830729ec25c5c4662a26795ab6939bae2b50c4e133947de918047e028d805f6a2315bfd18
z085eccc8a06d63a2a2d215b85e11853d12fbf0747dba6af7ebae87312e1095c0931bbfb2617bd5
z83e7fcd6e9b2d5bdfd2c233987fd7ffe71f1bd76f0afbb89953523ce93c67a520b98c7aca2618f
z3efed42827cb08293b313ebf1dfb393265dd9693e280b133051460f2e41ed2aec7570906f4f563
zcbfdef22f886545398378760329e0b9304fc956c55266e890556df0ea681996acd41fa69096062
z5269b682cf1138f5ea5cbe008873dac94341998ed5e2fef33cc305e6f14df9c10579e283a2aae1
z231ffbcdf1c900610c2a94ed7133012c2826e9287f6612e1bebb92f6686f9f6181cd58d96ea30c
z4d8e9734a55ed4a8cdc340f87420b5e2b43cacb5c9fe87155bdf0589b91a6c0b485382d155a561
z3f8f20d06db0c259acd3f2e442c2b447794ccfb6593981da7cae63651bc435d1bd1c831aecee6c
ze28d30ac87e9bb3580b6fc8f16ce012bbdb4b9fe341630597e658a0d087937fc97a93f3b93d126
ze8d89d622cc181a50a7b8ae4e917a3a3abb6a89c05ed4769f8e5e7d39e24474e0adb05c5f9c2af
z025a48e57cc49cde6bba08ee6980d8e98cbd71bc7ec77b7d04b561d8cff876dd6e06f88d02b3fa
zc52de748b534c3ca8e95f8c961dd1c837e87e964b11bcb11c1808bfae08f459c49bf763a07dc47
ze8a1ee1b70ef8638c014037a46197447807a1f0495ce934db29f75724fe75bdae95a6636381479
zba32b8a86aa7e0b836e51fd2d89c77923c84d0fa00bc80d3488a4cca953bb5a1309b76cc471f37
z8deefa07ab92cd7ff3e67625ac36f3ee2c6bebc03ec2fede93f779a449abf4eb0ff01861dab243
zb1eeb23e41a1c52ceeff02819458632f45498fccc5f56c2ebfff934138e49a3d876b7804779696
z9796988643c44f586df8993388241f6ce3462eaef34793541cb0a6d6cdf96395b98b13254a5b62
zc158369332a4bc805fd3662372f19f9567ac5d4908bb3c86bc9894f31b3cea7f028cbe84921cad
z181aac6d3f51bd0b6df0d8a8e43233644f9d56ab11738c41516ebb453ce852076d2a72dde6c773
zd45f2438bbf0b366b60515700b4697c25084fac11d91450077f15b5ea388b02f6938d63d8f561a
z1277c8ac9868ff605598f228824974aa31f05f245d26fbb017f8eabb8d1c2d608c3903d79e0d72
za6d426e91b9424f1661d568240fc8d05c6795d67bdc0476675029f01b72ec7fabd2f3a64a5b6f9
z39260dc0b30051ca7e5b857758577e7b12f8547d188f8002a502dc31978c0920e8a97792ef7e09
z8aa1b7fa43330a2657b00005e26607001922f43553f0e123c3e4f1e866af215a5da269a5e1e167
za745cbe67bd9324497008dd305fb25580d69499d1cdbed01183bab205f8d56832ca8a3c16dcdee
z9c2ef572c2d25e4aba906a5f53341a7f532728022a38d77b1944237981d915405e088fd5dca0ff
zbc4eff14f0eebb173abffe2551b2ba75d8f08ad7daea908c8e95c10b5bc493ae4bdf0817fee997
z6de832032e1137b27a565da645cca1a76d2abd2c44e7717c69083c750b3772134da76611fa2f02
z496f7049ae7b9ce59c7abf1d35ccb559c028e7a1164b00197dd1b7bb7d8a59b47ce6773ba7d893
zbecf7381a2a5dc5b7d1b1fe9b9fd239ca7f14994dd74c5b23cedea60f3a93f6d303e56ad07fa59
z21a4ed0fc3382c11f658c66028001f568796dbf4047157c6712779e148793308dd2ff23b29bfba
z08a486d2c1d40d41b5ed61d00d31c9966ab57263ac99288630d8d50ce310e6ae6fb580c7ac1915
z03ebdad290c236be644bc206eed636e3895535dff55b8de025f14ea9e9a3b9de0ded5634592421
z173860de49220b6d7fe109ea384fba9a4daea096756d1a392b74b1ad23342ea2c7a0f9733ed498
za63b939be0d288e59c9aa342142f92a0abd426454277b13553a04b22a3977fbeee147c9276766c
z285a08b4b44f6d1edc609cb26ff29eb07add57d755002c1968457274b5458e2752bd38bc01685c
z8361cccc3d10800718cc9823e8177f47e2e57e6f4f96f787e6c448360f91c9646a03f6dae043b3
z4357bf3b7f6adcfb72e3b9671abafba46ed45fdc035234bf2665114edb17e93b5f7daecd063017
zeb0542769c2fadb5a07f0bf8e2006a3ab2711e3f55c0e5758d9baa3586e94a35a5a3825aa774d3
z408d81b471173a9051db419f7a1172951f94d3686794452fd83b7be54bb1488630776283a0efba
z0b2d65946d1d5d5d83c7aa1ce13f99c5881d754638fd13bd76df2b8de5c12af30ee90deb70abe8
z43b4bd9c013b72e51f069613166e016fd4b9ec2fedf08dee516d34c148bda43877e5708ff4d6de
zcc15b4965f244c86ebb0a9e62a088aa7871bc2f10a79303d58eb20451c77b1934c690d1bae66e9
z3ad0e9c052f78e530067701560d7d3064a9893091247a148a785636bb7d25cd980a3a5b635a316
zbc675ae1a2a0aa858f0c329b6967e0d2e521487772092e1fd3d49f1853954f5a8504963187f74c
z717456fda3b4601f627a1dc5102f879555d45d98dbd77afa6bfca6e6e2eb89ef9594a5b3829f1d
zc4ec655125b7a98404cc564e250e9ff5d06f446729d8464a6b5d6807560b89d45c72051eaf355b
z8142978ece0acbe1a9007351b41e436ce734a9f8da173022bc815a469edc74d3aefecd01962f86
z16d76ab48cc5bcc7a54dcc12c6587b254b7a5e5be7d504d636ec0c650202d55ac4641a49058c28
zab511a4de127d37e2a4030b590ebdce72482fc51f1c35e3c536c9f7a644041c0940a4b5ea153dc
z0dd832d6ac7bccdb45222e74031225872e3e724156e04ff220d65c157fc8251701a6c9793afaa4
z73c0085f428cfc044abfd1b424a4d15317ddc9a5659c50aac691ceb618dc06e5c5ea982509547c
z5db84af02860d8df038fec29b4d47269757a728a89cbce10e74d700de3925d13955d7be3ed7461
zd99beb50866c9e7936b62befc33a7f356cd115da85fa1df41c982dad23749aeb845d330f7b650d
z341f08882e800ecf2db90b6efa7a9ff88d742479a9d78623aaec074bc15e1dcccc46065a55980c
z3fb061642af90b0a6a847727a6089b68f03a740ab0a235b14d01469746076fb05c982caf35ee73
z2cb640d7bd00f4c978410cbf3511eb325f3d116423b68564e94d5f197b8457dbb9f31371aa3ccd
zcefa250f11e0e5450b670ad5c7e707f0d4a871a276cad799aa30b3b56d15ee0721797e117054fa
z5326e832df76be8609e83ad3f2897f3163df08aa950be325be518dd041245c5eea135db2768ff4
z63576aa10bd3c0bc5deb6eac8c0b210563521bb086fdf3fcaed3adb15f6d496205ca2c70a10135
za24fa1011e7213c4cc93e0c7ee5e129189d3eae9385c52ebdabdf55e98d6f3ed46a9f9b80136e6
z2206417d3c64eb07270aa1e41d488e886015e0af668adcf16ca51069e6a63e5943929985a5ed92
za981c6c191bacb9445d18acf6588960c9312938a44f1705ed863885aa9af0c926279e6cd5ada0f
za0d04390c9e577285bf3584253835cc1cf00adf8aa0d6b35f9705942481c563816577d3a9bf378
z80c1106d0ff3e2ed94c356d6e76fc217f047cd6046276cb416d375e25b4b03ee6cc7e84353343b
z5fb9268279f960e80347c41a6751bdefe628a627e1e3d0d16254e38c60371537de0becee99079d
zb5e6322ad1b7f591581123e572e346a046ffdf35a88400f550700fc9914cbe9da684cb01a81f3f
z46f5add9eeb1c2cd8024189e9dde957a688d768f7913258f96feea1e4e3d25334fff9427ade84c
zbbf54939abd7bfbfbc39f1169926b6d78b6d7be029f0bf73e0971a6304c29087442d5bae155f1e
z6bc26953d760a9ef080ef913daf602f2e802fdbc4a2e4643f8f01e5ff41628c4b475a38612b9c3
z09db229ce83996660a1792a74ed1be501c6fa5d156515abe6c6038aa3471d18395fd8dec39567d
z90d3afb2dfb9de1d1d8bffc814537a591a15f3a97475aacb965f5237e72e62144320b065048fb0
zc0531ec439aa191d6eccfdef2eab8831b5e02eec72f09498d44dd9cf6785e4606861bd931471ac
z03e9be673a4ff44dad5d3ef1a94fa2ddc1ca8f8df11ef4a3b0395acb0c134aeaf9bad7515c0e03
z38aa2da85fa0f5d956ef278e132d0680ee5f2ec051494a0c2882abace03a987f75bfde6a37a77c
zc275ebd9a76199be5d31c0fac9eda363d15af730bc1cfd26ff590b4d82e4a4302abb7ea301bf9d
zadcabebe23fed53c299f8c49863a806471cf1ada2c53ed3d0b9e5e836f39cee1c2a778bd078836
zf42c4f6e267a36099a3aee9842f135e09e1647df4c47c27c54b586dbc0297a42a6d5260798ce25
z289be0f9554037d686c12272b8f47f31bbdf13b53e761f31ddf948c2375be51c045ccfce9ca971
zc9f339b67010d0b97afcb809947578affb993a3442700dcbad939d6bb9b551dff0d311a33d604c
zf46e38d2a8395662cf2da0662a1682c9d2e2fc6f08a40d960c1b598e897622aa47ca8db187df11
z49568ec38820243c9e3a71407caa4f4842527f89b03ade0b8a68f6018f5738d26e6dde84ff40ef
z8d6f23690155568c4b998090bd5520842c2b25fa91c255f0fa44def43c8e10862509ca325ebed9
ze462fcf012f04ea6729e55162a691ab6fed11cf8e72373189955ac19fee76202c5bf0cac5caac9
z08a4c846703459acc571fa139468ae72fcf77ac07575e161eb07057c3b48d53bf47ceee3f46262
z2327930107612de9df2a2461327755e8dd7ca0f0e08b823185456ba4aca5a4ab0be0553cda8ed1
z41745c5cb23b6abdd2a900fb242fce666b0c7cfad4fa2af1e7b7a569b3355c74b32c839f2aa594
z94a53992037cb42c7c65d28ddbf84dd896f29470b576669c008516b13c4f5d8843a22c54e427e2
z76d4190df610d0f607f07d0eb1d52a8a5d9bdfe6a60ee5a0e8f1592b735d00ed7daf4de6e9b826
z96fdd93713b6a79fd45d92fa84393da4c75224d80c15e49db6492d3a52d966d30b654c03972460
zebdc1601df5fc27c19a8df169aa25282173ba0cebd9fceb1252abf7b10bbdec9d27c081a0dcc7e
z984a7d2ee482d3ac344cabc797390843039634b62b7c5f87df642b0f5db961dc85ee47ac8f7e63
z783b9ff0dd823980839fbd7f6015aa86a1ee21c79d5adf2657b2653309ffba9c66fcd5538001d0
zf0c345c5a8105e2ceb0724bdc420868a10f488c67b9b68560d5982fe9f391c9414c3949a506716
z901eafd16b4ef2b35fbc194895ff32e28cd4fb012f2f5cd4125f61559b880aeb56db188f0409b4
z6a0cc7e1b56dbc0f3d47f1b2d1a6b9a3c48aee971bd9c9315276318db049b1f7d48781902c5ba3
ze06a0364bc4072cac1c82d83a857753cb81709a51178433c061e20a2a88f50e2c6c69752352cfc
z3c7b5efae7bcb01b997d7fa890f3337844969f63a0dda61cdc7ec198939fd6eea8b5696324af68
z50f5a9570e9190044ec40e628ca2e066db06956791a2fb32d4c44a42a4957a124e3203956cde7c
z2a454926d52f2e84d326f433d8031493599f3a4dd5526b407444828d699e8e6511c28fc4d73951
z45792b6165b2fd8f3bef7b07695d8ef3b144a3ce46a61eafbe5574b85adf65686a3824bc06dc0a
zb3ec531a35110251e4a715946a53d7ca49fb1e8a52b2a07a2aaac9127e95c5c47f6705f40ad05a
z8b859b5d94b4c0d95867d460ddc55a917b3dd6c4f373d3561eb1d84322cabe3d720b8bdb2a40b2
z2832f63cb84560fd166e56fa45a45feda8fb9685c8fe526d909211edbfabb813e64a3f3a1a4295
zc0df8236fd43f7a94e8e9ce4ff72d84746a2e942f0e162ef53207a0b763fa2d47855d353ee10bd
zc3dfcf33407f9f64330615bc445b42b78a11fda239f9d3c2839ffde4a717e7fa14acb93f9b320b
zc06642a7fec3ca5fc4a3bcde74e48dc4c3b65c4a28f05f8d732c8bd7a72385bc48ac0577fb6e40
zf5aace254a4c0d214864cc613343bc476bd7b57cfd33f4628de35bc86d1689c7a84cc0d2c1f727
zc28a6981cc87efe0914b4135822606058c6176431a0b72bbbbded7016f4fdf16d09d480dfaeffe
z7b24b8d14294072742bf09977629d83f020b24a2980a225af78a52cda8b005d1fe5171dacf477d
z97a91da40817f0bfb7cc31378ba0e20836612dceaa860ad2cc8ec822d32cf44941c27a4cbe1b3a
z40d37de2451e5c019e1bf29fa1b6e132b750fea478371aef6d549e6bafdbe15980a8aea40d4625
z90ecabf94499a333c1edaa29e1e0726c4a2437aee6f1011f33b40e0d79e8551f096782d6563010
z0a8764e59e4802b0a64542ab3756b591a679e3b24bd54414e044918f1e41443bea500fd7afc35b
z524a1d1da8003d5aff8403d07d7df954f03a7d935477794ab46c6743aa3e955075276b5dcdaf9d
zf6ffcae65cae1cdb4f16518bbcf5931e79b943e1f820a2556c8f4fe82fbaefe2feec631c2f4dc6
z8bc1022ec8515a6a67c7e0dfe739150e8158a779a9485da0fa65449de84be01914f2dcae2e06c0
z611f20c6c3ed5b0d042f5288fc188c86b9aa7954eeeb49419e67073565e051c3ffa6e163ee4d2f
z534713c27a4382dfcb8822abc53ac64317f9c98b3e8ba7a1607bc9ac042c47a1aa90817a6df9da
zc078792a53c6e55a3c097d96b8a5b20b6843d3d82812acb51d384a02b7c7a441d6d08139029490
zb9d136690168f892ae824fb6589fc8c6c9e3f17b370ad9527877989893cebed4db0d8d9c6e80a5
z3f619b643b8d12766d1a301230e0e64ec876e05d62deb6b98fcaf1f18185da94af31d9c7a16db3
z2632f266e98215bd889f856a62d20d37e0916c98ea9117b4b12d1967151a5aeb5c6e928eff374d
z784c2ef721ff93cece9f47f5059795146e6efa66e6b5819a869b5747dd230ea73c217b38cd4f28
z0edc340c912c2bfffab5621dba287f31f22b603a62f6db8f5bfca9f6dc0a02187f618f95ba52a0
z4133c6afcd544f36b6731e886fca931f27a67c6472b0d7b87b636d34b8664b3608dea69bbf4e06
zf9897beb0d85e79b5ff064df0ba7e9c80f1b97be71df8c69423ce5540c675e78c058b2cc6d0d1b
zbba480fadec82843e58c919ec78738bb51ebc73fc0bb6788ac2dfd8d4e426b1c6df881e02062a0
z67e83df81e7f30758b9baff7ec051050042235c1457fa5e7f7fe88dc0bc36acc7390a580ef9578
z5361b5449ba6f20e200dd2f55705120a0a623cb94e94e8d8797ee7c58309b3159f3eb2a7d68fac
z5ca66ae7627356a1a94296fc459cf8d63072c70335aa27a68f1429a6c967781fbd87c4125d1cd4
zedf86b9a8f4ebf84bd8403d98de592636f43e3ed9ff8493ff8e4eef9b1398cb7283097e9e0edef
z5894a3a5711db3a1002ac09a74ffc05bd1f77b1057d376d4afb2434c233b3898527f0ac8563fc5
zc366ba8acba42597526dfd3286d3aa21aa322e0cd7e27ab0a049552daec9ca8f7ec8c400edfbd2
zdb7b0b46e1847ffcd12a53d7fb999fa16fba593c6f733a4b2e1757ce4725c2fa78108f11bc253b
z90741ae12720ffe1d4c38390bac322c0d8c2b613fd83fd91398e91de367aef96dff5db3a3431ec
z7e1e3a9b4525c104e389d5ff24e2372300ef25d86815a4be5a3517f78c9634789c5107d342218d
z32a5a29e57a8b4e678724e476121f7bb8626e51fdcd115fea17c03624e93b1793a6f0cee6496a6
z4dca3fab2a2999ab88c3adf6b318b322804b25c15464d15b0d4d455f169deecb9f326fe06ecfad
z5dde23ce693bfbdb6d1fc272d79c2d6d29d57a605f0e4780c272f1ec23107100e1fc18785a425f
zec586c11ce53cd452c2319e091aef8f6ce158c5463ed6f4f20618e8e5a6c43ce2c61197a4341e8
z76ab2237550e30d0167d3e725a39f8bdf787447cdfcc52641528731e938183f0b52133c040ac49
z3da5d71c364ab7fa84b6cd3be85692a7c594720bb289832acc06e78dffa9acc22c2db1b6d2a137
zd239f63b57356464a155ce0986179dc5dcaf4b47a8a801728751b89409a869b4604f2a55042e9b
z98404027abccc7bf3c5886ef770f46702bf44ca6fe2fefb9dda902e736d9a913d3d069428b2e21
z8fe882e5d6fa9dba1c980dd1460f91471c53ea0ce8e88179b806d707dd403fc7ff1f309c178615
z0ee06085302743e18b789463c664b53804bb4e5ec27b464f26365d3e352d940c9a114e689dd05b
z25d9da37c1903d8b9d2cb4732926b4c085a4a5c85758372ae755308315e657d024048a48c6174a
z7a18f00ed99447c7340a8e5232eaaf1eafb05f6dbfaca83e8335273d306c19b2185758900b4610
z8488dbdd854984ca59057224bddeffb8a313e116b7aa55430b203592f621a4d2c4764867be2ff1
z0922e3548e7ca893d1731e37ae6c29e0156bfab0ded1fc3620e2f7ed58f56e235510bb6f8fb08b
z3315546158e8b9754aa7a397a2dd98293c7ae50eba15bcc2bf254ada8eca0a8004aee3fa4b6275
zb256185f67d987d1f097ac721c722a7682b9625cbbf5990af45157ed6adc01163f5d9ff94f7d8d
zb80e8bc3ed0c0679e0b1e4206126b742b7feeedbc58f1c4eac5da2ae9c91ab3c00bcf370bd9b70
zc36182ab679a3943e85ee85ba309936612c5b637af802063b7ea4d16563f832622959e4fb417ef
z23f6b04f7b6cfa064e1e231dc40fde93570ef176cf5bf105db459f012e0015524309dbaf8f6273
z6c77940c723687b6e6710ad5bf2a8baafb322305895a5cd87cc16e33aadaf93e780b4fe480e2a5
z4bf1041a4c249bf00a1ee6c57de5839fbc15d015d5e61618af3ded181512f598ce3f97f9a4c90d
za77a15ecd43d15c9c438f8c78d9c0780a85acac4cdf6019f6f2fc537816d1c4700601ccfa52a77
zd5b66ae4a75d967f7cf4895ad4809cd739239f66d3c02be1eeb57ed292d9ae43a3f609dd8e3f73
z433a2b231546d2d40ac7889fed9fbafcb825ac93560359fbe9af581ca847dc58a0e851e92fc427
z5d225923765802c5c929eeded7d994bcd5404a5fcabd3d3601c4ad1d4fef8358e9160a505f7fae
z641f1e35f4dc32cf34a91faeaa2c33e8b1af8e4361f150e75e689eadef45d4c49af9418a993db4
za084b7526037fbdfde58eb3914c83f654f4b823364daecdee10bf923c132db6c0d646df04a6b97
ze12a0dab055774393101913925c2d988aaf92c3f0aa60af523e19a575ab05bcfb82f665fa20292
z841599949d93f25c87df59a86fe7c4303994a39589efc498918bd9d466d980813356a9fd0c43d0
z57b42d6d610ac9c611448523ac749c9ec7e18695a603c0ec7d81fb5d52c044db3f76b830f84a44
z970e56337d220786a4fd4f0a58cf71a64e959c2b2364628b91ec734acba0f439bed652fd411437
zfab717ddd9027f8c12faba4fc1fd8d958e203496a2404fb44db6ff9c724bd1ee0242c479471fd0
z02231bca0cc5bb9cb1e960a3220bdd7e751f778770128b12260288154851fe79c226d2eb7654db
z079e8efdee0c8809fc8fde2a675586dd2f1d7e8c82943836fc27bc200a0dd1bdcd42d8adf3495f
z02266d5caf818d808c0d6af16e36d6e741453479b996adbc9d023e07f1d002caaa50b503165ca0
z602e76e2958677f947785b8875051a47c5e228e099d628e2c7000242d599c1b7dd3ba0c94c0808
z56adb587a95aded4282e4bf8c59186138e656c28117982bcefb681ef8ec1a320bd98bcdf329502
z1d56af1875bfe868d563d9ad2c38cf0590c8a55878a1fef47736a6ca71706a471d74f70400f3e9
z8d1a73c1619028290ac7044bab1ff39fe43b17e557c8d61b7cdd9d528abd5f2eaf39315fd9c462
z27060717f2ec1457d8ff529401e308eea475bc4c3c5a953ced2df543eceafa160abc39663c1e95
z7c2cde505e1ad5cf56bf5c3c0c50d7a7ab8c6242180458f6b9cb2b797594ff5cda04d0a0db4644
z0653b5987e929db8e79ee1aa3da6b12ebbc0ebc4ba2b16369238e26dc0d806bd1a117cba51326e
zdfd17d20004e145637f719af82f14b90cc9e166cd0fb804382c219f809d363dfbe35e6a17a7f02
z2f4d88f84888f049bc64115284d646e4710e43ac126dca07a2c06ed05e6c108d74874d31e6f283
z488f50624f6416ea9c5ae86e10e1bb058b9f05a2787681f08e6bcbd0a982105949d214a4b805c5
z76c15cecf8fb440b8a1d8bb95cb63989ba86d39ae241afc0ec6c648fcfd7486e8b39dc5ba46556
z0ba5cb8b7511832d5d3d98c457fe176e58ff78c6a535395af1e82ff285dea28a447bf5379af83f
z0cde0d0fbd00378aa57e9748e3230beb34ee6cb42c8ed476c748d1c6b3df3c86b1e31c2909f1eb
z98689eac22fd294c413db3fcc8c7e29703228060b7bde662dbb998087ac371f2cd0ccecc9a732c
z028204584d207b5c501b92ef6df9527ab21cfe3dd639370ad2bc93bc412db58df3f96dce8f07d5
zf98f886a1b54809ea4891cd2eda31084601b013c99a0bf980154573fccd4d6c0ed4ed8cb94596b
z77c874260a51c35c0daca0c98f5d116fae5d7e10a0c31f6d0369d585c66ecd77353fc7f47ad3e5
zbbb830c99c3b710ece3a9398539eaf70a397dad5fb9adbb5a1ba87206540aa22df1397d0e0f80b
z652a243fb2754699d2437bfec237af8373fd8827fb7355499dd9fe97f9890bb08bdcc92c507f39
z7ce5641e6ccecdbd2c5ca8bfe09bd927e48684b4b913cf135e62acf1f715c64cf374680c5ea02f
z912d4edec31cca1ced8f64ce2987e3e493a6252eacbca531a3edb1798f73e25481ce805ddba0bd
z222fb746bd0589d227c4fae1b129d52a88c0f57aeb82b7f717ca00145b00bf5578424e8ec0c5ad
z80c49c7a6011537cb0f57ec2fd965b9ddf80f675a6b60b6316ed7a74e664dd8c10cf28dc884d48
zf7d288f5b46f3289710c154ab7b1633181d53e16136df05c653e27003588d480e82691590659a3
z2607a2460c3da29196de35f54bfd2cf41a6f3b413d8a0f2817724a6d3383e85d819f2b11a4d366
zb590ba240a19674ad0246172f9078b723ab3a4fea48f4faab0576066b5d30b15d39be6a7e5b5fc
z65b26e31cbbb859c9bd98baf2af397fd00e708084cf62f9660d7d184bc8ee33d19cada608cf2ef
z0946aa01dfca5a346c4ada5c05f343a7361d40dfafd74c864b0e0868c06b974ce3f13acc234ed3
z45a795b4294690adf748db4c4300cb142af42cc3f232ffa0f57b88e5ef5857c34c85860644f583
z2a29ca01467f1d23f7451668830428376f2bdd1335f6ab0a42fc90746b27804e82aa0bd2df8257
z417c6329ec78df4b3d0d47714d4675ddc65974b4faf6ff124ca7021ffc1459170ea9bdd05c247a
z89f068b38b8e5b5444742c3c40b7e445136aeb181ebe1050b1e85c4f820b1c65c9e969545ac2d9
z1dc66da9f5fd6dc6918bdb6ebe1bb0df8a896b2e9b2e9424d014aa19c3001522949ce9b3338b61
z10aef979b4fa4a98d7b869be86bbd66ead4301d978e7d4b45bdef292615676e24ee0761919f545
z2051638e19704c131d73ba526b91bd35de39190c0825dddd5595164e0b2d5cfb0aa762ef7b5ed5
zc6085e8afc2f866bec9d5c9c4943a915243b7a315335b46bac060f85a368f69afd1b872336d7db
z26e40ece3426c0108a0f03a3ac0cbafcdef26f12c2944cbf33c46c6df9f4f96672403a2200a77a
zcaf05ea7ce83219684675e02bec2a1c756e4a2e9882fab0959b3b106cb815e9dcc7073d021f273
z53a9a153d481350ac2dabc08bde181f714b9006ed3d13ed46f643f6fac210926c50f8b6247fcab
ze241b90fe1dbd887ed4be38354e52f38d5ae43638b99aa0353914159d63075239dac443a1bbe55
zf1ff26b1edac2432d0e7d9963da262db1a2b81645db9ab7ed51fe18ec2b196ecdb7bacd99e1c2a
z87029f97dff1d2c9613011854e9f3b5f6cb512bee917b612a55234838eba93a79e99a1861bcd61
z520909b0070a9a0ece6bf314cdf4ced2b76555e6ae8920be9da51e8bd8e3058e21f9d9636c22c6
z0f9b998cd2a5794d3ac26be454b1612a52e06d7e1d777c0b5621ee344e52fa0fadbd47e8c8f555
z75d5025a90338efb0893e2730debcd84bdb41479caf3ee43b0dcb4bbeca2fbb6c34d8cdc28df88
zdc80e08dc5c51eab65b5aef666a1636710bf678c58a70136cab0c60282480cfd934cb5dc149e1a
zaa956e8d29a32d6518621c5e0f1f4b1c0132ee4f753eb548460d0ec74752ccc741da469bb7d7e8
z9d7ee059a34bd5fb947374a0993f56b6eb9a88bbe60907f70f26a56f88fa760a48f74c1f44e8e4
z958f6bab8d6a915078d0532b2beba07e48f2948ddf2e8a7b07ce50e42bc5b5fe49ffd81da2403d
z1025d4cc3a33af2e178d6d030e8857b4eed1308663a2847b1dffb3045f29850235267204205928
z9d3c4a3af1241a37b9785375e46ce3b6ea2f9cd7f1129fb4e5fcf746cd1098aacfac52c8fa97d0
zaee740ad29be89de75ff55c7bed24aa1fa0a1fa46f80bf84dd052d611b917763a28d36b8bcc8d7
zc843889c22e26082cd64b25eba6dd5ee66fb56651becb8a76a4cf2f0f5c0c9271890d0b1da7ce3
z959a7c02139ee6ece1260c75db10c6af653a0295a83f43f7e178e9ba76100f588675755471536f
z4aa49be1d734540b3042f7eb605558015d1d2fb4fcdbf3cf2cb6d9e10be0a664616ff039df7e37
z4199f87ea81921b0892d208f3ae330b0314db0dee5a422e6790926b48585af86ef258ab64e1962
z8623c96fa527f958e99666086328032d73f688abcbcaf00fbbf18fb9d42928c703467a5ecd19b3
zb993c9b3b52da80efa0f3202d7a8b3df24e4c1a9bb19be82fc22ca13df7abb9c61a10b41740b24
z41e939aaaaf81ec67b1fa361cb0de55c57410bf6925201dbcd1d4c0ca309d41792538b8599cfb3
zdad5d19bbef43a23aef0602831850631a724a66ee82b00c1c270c60fed3e7ba47142d6d4f69d36
zd56882207ee6e86cb127c3e5dc9eca08c85bb9a725939e681115ab4e209191d421b38355434199
z8ce5f087c8c9082c08051c972512783dd2a60ef3b28a8cd6c31e0b7084e1799aa49878a5c3491c
z46fbc37c1f76679b6b3ac39bbafeba54e282b68773cd673dc2843764a5403a5a6f17afb0a792a4
z0a044659d61b0c0e0358a8cecf1f174ec5092cf3c1558eb0ad1cfa09b113b9124a86edc3cc573a
z6a678e0cf38d3a814a22f74005a8882c7cc4e45bfbcbb25a30f08d3e1a359b56e8bbc3d66975d3
zb331d52166946b82da7a0efab70c56943edb9f783feb7f9116010621ed89d8d17bec7f9b0e0ddc
z65267935434d8515d7bd4bfb8509565d31649c26700b9ec8abd52d5598d95d9236f80147e7a100
z53b9ab439594bff6b5eed988706781cfa92026803358bab0539b80355042f8e7d65f3e33944d51
zb2ff8fbb9759c1d7fafb769e484dda8d75532ad314282882ad6a6fb3eaa6fc734a7fd6f5424ab6
z4b57fe91caa0a4dab0379637ff20b727b63cec9586c9bfcee507d9ac9c440ad9d05ddb85b39405
z81887a8b6ffb4e94458f583c129965ac511ba2fc7b0cd1dad08db665cd996c7481cffac1de559d
z134e07ccb1ac30c9059a3eb760b8da5a90418a84e69856b60d0d319504e5878d9aaa920d976194
zb263fbfcd21b29472c6e42a8e49fb67dd0229c7f89b4de7b6e237c33c1a11103bc8ff72cff9226
zb03a6d3c4add8b4519b36b18d107d9711e7afebfcc06c8029566bf2db4272ec6ac7776b0d77e1a
zfdaae1fcce5eb38cf9db31691c278afa65e66e83af25bc41aac02151a3021393180d0f02eeeac8
z7725c6c8728f0c44b87e6582f9377404a6c613b243f3dce38b1e83058034203b73e3b04195ebed
z1614b7878f4a5b2b74e8c01368301d1a536136749b81702bad566f0fd6ee3f53512ebf08d75794
z9e892706b3680737e110072d1335c1a3d4cb47fce0c10341831ff9b231ea1d3a92417b29106efb
z50b2ecba007d8824777e8ce635fef67fece7c3d404c950acf3907efd38910cbc2a33c74bea286f
zd6d38193635ecd4c4da95ca25ab5ed9a9133d754358967b5773254931126e63891dcc8ff4eb238
z5621374e77284bf416918aa00765df1be5ddfe921beb95e719a2d7412c9b1b37d5727c1aabbe99
zebb3dec76f9bd946b0abd6c951150f3eed445d95df5bdcb25d8a44ab9db91bc71f150df95f2c12
z44f9b763a22b9392eda6184dd6c82849bbb448dc09f33fcf2a499c2fcfe226e6ca2cccc68703dc
zd78df56696d3da4c052391c6574746e870866975644831b6703a6ddec129de10f9a26fcadd71af
z3ae7d2d39b14531e974e35652fae7c0cd86ebc2ab2eaaff485ab1827dc04b3ad99fdb13247b472
z7b7135b3ef0bcde0ea13ed2c19477679c003713d6672fed60767aeac8ce2de835d70b82e1d51b3
z98b3a8856f9bfe69997364b6df6b11493811d6c1243263b8796fc9713b52101070db8a609e8526
zf4dbcd0c6b468be23a4f318f013ed004c7cda308d91c77d58bddbd72068decc2c8b76ae2f67af6
zd0187f35e79bcdca0b7d329014c23297bf04fb26d413e62106bb6ff21a3822553a6a9b65260e34
z794a807297ba0b330c0597ab2f13e017f954ab9f7f9f8fd844694f9d0e1d7c63c3864e3ad5b1e5
zf044fa4acad20e7712dac8003e5c4ca09396f658a2e34c8b15a9a7dda2eedff0336b3d677d64e1
ze2ada0584ac76a1e76fd5a0e2374f6ec2a4d2a4dbee3900bbb704aa23c77df8d7aaed3852c60a4
ze992007351cdaf21d754edd0de9d55a2f01798cf9c343788c506055ac2f2b2f9627b33f92ca630
zbdaae03c7ba537aa05ac3c3f3c6d4d87a704de2258baccb1b02e231d32e08fcc9ed594d4699add
z3cad467535031001a70b504ae653edad9dec9dc87d8c25fe9b3e6a21f5d5b84468175a9d3f53ca
z441b2f549c7e219204be7b23dda4df2b20ae23bc77acd52af298587149337e4309419dc57296a9
z69c616a7adf08917e07c8f24f6070ce0e5b664303cdca962584d1dae453b3b2122f95b1fca5123
zeeaff81417009cc2e7187a8cb26ab3cf7c39c04bc5cf512c028f6be38db9ebade5195a4e9f5cd2
z2045d3cee83a197232cf69fe6ac88c4f33f837102cdabb26c665685455ce4770d63cf6571c3284
za5a3b7351208028d2aba2ed6086dca555f510d03bcb623474be2d110a583f65a242b57c820bb5b
z74ca51e7eabeba87e094171b8e193c946ec97f1ea73851b0413ce0941885086b625ef253117400
zab72115b1820f012c5e21ec3ab59ebf80dfc4f4fa7dd2d8c95886edd73b5965ca2a4630d447a35
z0feb0f438e29c80715a5b57cad294426ce342c3c927466fdea522cb4f09fd36b3fff3bc8219ba4
ze012a24081f687309239e2bcf58da5a886d715c21bb8d788cd0cbd3f215885b563a2aa45356b53
z59c957d87593f79dfff73548e019a0d31a7b235718f79faab330f87c2297cebff1037b05c70df7
z94a959dcbbd2a09310db85d44e350ebc0a7accc715aeed02f271580ade7464f32f58b68498eac7
z136481117c14e4b2843a103d4117373636e5cd6e366e43329a5145354757d350c5a1a2b15a325c
zab3438051e1c3bd23049096ba038f8ebf519376a96c3b64f0ad4e3a2734d1f266c33af7790b20e
z95811660c7f786059bab89630b4ce47a019ef3cf020ce5fc0bc8787d717b8f4a1dc154098ee362
z3dd0d6f19f7081ad29f9a1f39241a21978b4d831f0d776fb01377d38fd2c7300dab02d4b791bfb
z4fc29b36d344eda67fae92b2110d4d4a4afd76ba4b446a3f37c927acaf5117b710476002ebbbb2
z9d635e0a3d080b2ed5805c48388dc9808edcec0f61ddd69a95109f24162e4f4d2e251eb5fa600b
z9f094f85547ec72e3736dd6b82e67f186f3961966059feeb44c0517ac681fe756cd1609e93b452
zcec60abc8861e5888397760df9ad67f803534d31eabbd921e3d1df8c835f4a87ca453177d6aaba
z1602581bdb896543302d8f6d9d98e978045dc2567ab072350c7aab6481b52e5a4c3fbff5327d6a
zbd824d15b71eaeff283bdb79895d9e134a45c4f14e4b2365c5e05ddc44fa819708b3b38b2db5cf
z147ca82058039289ee86319ad3c8ee4ebdfc19581b00994c8c581e073c7740efa8c9f5962dd267
z24a7553e86f09ee62660730654f59f17726a3dbd3de95a77c88983bacefe35c2270e3e473f731c
z1c5d5790fbce6a79fdc8e6daaad30b5bbb7a3f2f1b1e5ff5402bfb13a1b77464eeaf6434be53b4
zd818793b8a95d8d127579f66eb9c5eb0610c1d92e1c5da3910a83f9a177efde80407d89c6aab90
z7a35c1c771e58b1a984aff2e03a308bdfe7e3eb4b9822b22e53848c96bc7d9ed30d75714937437
zf3d39fc2f1cb0c24fbb72aa07a68b1fd8a1db5ce868b51abaa1dbe11b9751964a5e7a97e2372d5
z50716a1f923aca4674ffadeba5e03e3846a5bf6651cdfff419605b792c061133f7be5a55f7ee70
z6764cc5e9cf6834c50d3d37c86f030ece043585059a7db82748ad4f0c48511112a11d0fa9b51c2
z109e40e8f3ef1beba6c5b7c946e5c8d1687a5cacb7282a16710425ad4b8e89032372230ca1eda5
z48d610a4f3b2cebfc9e7baa70c52203f1cc8bb2a256521ced1f1fef880b144c173af9c1147fa45
z7f13d2afc5e7b53511e54f6cef881c06dc82283239ae88527ceb790a25d5d7b19399fede1efcad
z98542f0c875d5dc5742baa3fdd8b28158d4fb8d976c97de35ccf6d9b6fb7a8c8efcf9558d1f6f4
z6846eb09c044b67caa220e3b1543949f002abdf3386c71be213def6463790a6cd76d50404b4cb8
zd9fca958bf5799e6e066a640ef808076e205544b52717ecc1cc2bbc5632e1f715133426cd73a19
z2f3cb2189048118b6a3651c46c4c00f5e14e57256794189456b3240968520f62dac42475c1f94a
ze7af1b9a5e99fba3369d1c0d145c4ed0b34701e4e87240fc69eec794e086e2e37a9a901e9225c2
zaee01a9928736bcbd5e417b25e62684d48a1cf9305f814044bf115cb6ab288f22ae60d5992b6f0
z52e5bd2df57d52404970f7a932897a5070048593e5f74c5c8a61a9ebd86e56cdaf245d86b9038e
z2e76a8afa6909b75cfd303ee1025ba37403687f45e7228e3cd7a0aab0a555ff1f4b7b216f78b2a
z7b7b1c9b599c9dc75f44d0061eaebe95c602ba86611cb400048963daeeec8d1ba9ab78b7f2859c
zb23ed9db04323b2eef669f15cd9d2c4c5deaf76eb1c952c18134209edcaa5f776a1d341f410384
zec17df9367a770c6f29d0d17d9379e81f1a59098b7fbb21ca6d1cdaa030cc0109be0dc4f9be6a2
z1c0b23b9530db006f9350017f111229a161f81dd179d2c582ebf95fe576f28005fe15c0f2ca640
zbbb1008e61bd33028a02199a0e92ef269dc6f5db1e7f3023e68f27d36bea1897ae5dfd5de317c1
z25ef48d1cd0827c359083ce09f69eca5c757ec1647f2c1892629b692c54a57b14b653c681b1932
z2bf6db15432a938e3b06bde86caf951e4a68c9c0a9abdd235a46249c274227000571c7afdbdaf7
za1e6c6b978bd5a9f5b3c62d356c6b4acf5a6983735be48959b8c229b4bd47b0b9a1105552479a5
z1a45eb7bf4bd71a30ef1795acde156f3901740a7b4667349deefd6ce82c648f35be3a65df9f17e
zd71b1a8f0a9c9c21d83122b9b3a1d8b96dba3d8af76c29f77cbc8ea2d95d73239391ae3dbb2393
z477706e5840a184756e52d72f463505fdddc01568ce90e99e261932211c0691af1e7b05411dd8e
z202a042b9e0265866fcac3d2ddbb617046e7f214dd11fad0fdb8ac4cc26d418fc3299b82eacacf
z893cd942fc432c9b29fc4fdea283cf43b1687cac259c2a38d973e534b29b1c6e19601ecb926585
z40e8c94ce9e6fcab2e09a80daf647eaf28ead4c65ba269e88fd81666224e470df28639fb508f6f
z17cffba2b41dab3791dffa42fcfc2fa7f35b1d8685b94356fcfa0782ee1ba14847902865e7730b
z8f2c95d748ce82582d1de1a6545c535ea11bea3939cc8ba48b12cfb65f96be143563ca0c6e7cdb
z9525d4cbf5ecf600208758c15f9f7c1225c7bfaccc4f73c3d6a42d8d0c40fbaee0b2846a8cc566
zd548aefd2761ec54ffcef96711fec649393d22a34df7af836d51b8ef17cc4af734b04b476fe41d
z8610ad0c79f1db6a4ad910141714bc85105829e1d407e59189aea01c625d96c433c43a06ea973c
z284918639072a4879e1707431dfb4547f8d416e8e23765b8f133c4c364ebcac87b7215bf39df15
z941b5073c25c484a59167688c13c2b3cc115f3e6392c5020cba0ace5ee645e43152e8cbc70cb3f
zdc9ccafe403be3b97f826c27b6625038d0d4f4d15e8b107403d526466542fd9bf51f16e5b13211
ze0b07a85026727f72131866889d26d932b61f4520b6d2d4f33365e236312b7ee7f3f6f3f8ab26a
z4fd1e35dcfe1e7876c8b7b926ed386aaabbfe263d5d488ab8b669b544ad7660bef57ce6222eb66
z914729ce1409c5aece8e310235afae6e47be06f1c5b66715323a44810b33291d4db10d25e8474b
z1ba1ca184a1abf3e69ab14c6a61b2af888a97d770420d3c8731d42221a648505737aad1028f982
z13f8cfb3443bc8a91330fafacd23dba2bc9281ef9bcd37216edbd4e505a4a4df9d33f3fddd7f48
zfa0f507a701f9a3994477b9b1cab86cd81b479b4bffe026bc75b08f6eb3e7c34b4547d03885091
za33d6b7ce912596d3ab08b7eece15cb592f7b3746aabe0e47869cb074725307289081f7c4d2dce
z83170f5ab2135b04dcb28052f2fb0997ad5abbde4798f49b6dd27ab094c2c7aff2756dcae1a92d
zab185cc6102f5459340ae61c8fb1ecbe9c3614d4b46d498fa7ac28bbe3dde6fed571619f18b428
z29476cc2ad8265ee67957c805bcc4be921b4f3a669551320fe076de74079724e047dec632442db
z2bcef4118d9c80a1b9ae2adca2f35923866b989bfee5ff151f16a791c8bfd67577456ca985705f
z3ee24f895a27c459547443a6b2ef22b685c2907a914e5cc6b07e67d5651b9e8f4b8112a4054fd8
z6a080bb0653589f1a666513382d116e54aecdb914acf2fabdf288ba654d6aa9d2ebb1a54b6e885
z839a91b88341d138cb3b5e08b348a19bcd31edbb41f1a0cb77141c752c41f07f0a111e8f95337a
zfc62eb1a147910f06055af824b85abf63dc782b58a79029e0c2511de994b7fefe5283cdff26499
za667e744a012a4cced7ee1d9efcc515fd07339ebfd0d63388f55457cde3070b2709e4f2491f576
z82a59a9319de459007f4ebcff93c874d349aecdc4b8cb886c8e65d97d07022cef9dbe61a61bc04
z2a870b07b2d317faa474196396cfc13b3901ed75bad46f9ffaaf5572859d701bb927b1c05a9ea5
zdc9e6b771a0ada5f76757817d707117e3108a76024c5dda85133fb21f9196d50c7ceab400726f7
z1de1a68244654e2c74e9429870d8298ac66f262d9b3e520e6af0499c7f94d9ce6d92f03bb1ee0f
z5da703e60e99b9f1ab61aec2cb825bff84cf24e54b5ec06780c6a3fe7a38d6804a0cd0d0279416
ze4ca86ae3a99ac7394f47090487516659c77e2678ad5e8f2b660d403d9a98d769229e39b9fbc67
z4a10742aff6c19d73565437b9649e48c810ddefa70f62fb4d6df765c29cb0ecb56911786d4112d
z439b9e6d669ba1bab3db8104690be465da649c0472102413b289baab893d3fc3e6a134ef86fa7f
z3bdc5b5130051beccb7f51f406beb66397e154c8144d64647ee55604a4977054b8444faf66a4a9
zb9aaebcda622e3ed090a66c3be9fe6dcc8508193c096e7ce8f708f585051d225dd50b25f3afee1
z43a8b622e088834b4d956f9a4d30bfd93fd75ce2019adb5c9626c940201d4eddd96073a71f97d3
z2d37536e31fca46f6236bd7647ceb34914903ee02df57741234ef2d05d57c170e1746a03805c3c
z8004c09da0073b66918c8c917104290012b0dd87f1a210682c43f0b10e0fe49049f35446786585
z52d56ecfd9379262de250d2b42eebdc9911269a7ed8edf0d082e4e9c46683455d6d8f80dac49d2
z0f0423b29c859e8c7cb72c99d305d3787730d2d04f8a8de9d9d2dee5f0fa85c960573c33c07dc3
z79c73a1e79b8b35b4df7fbfd010c26f0cda26830f7397b4d85c51073dc0cf420518a123dc6cd64
zcfc9297d0e239552bf21451e7a771810b61803e4b1f286bbfcd4ef4d7d35cc560fa4bf22968904
zb34711494915be458c1d83d23c52853b94e1853adc2eb4a68c564c7448c2756d24f5e64ffbf830
z5e7020575ffa646aa498a3e8900d390df4c439b6e83eca245790d7e4d723ffdb9ca01794f38dee
z4cfb6882514ea509944bc0b12a3c2e2e9b89687f85f3ea7829844311ff1b45dfc283bf00e967c5
z90b847c03c42c114894ac07290e968ec70acc98fcfb6becf629dd53cd9203105cb7dfe7b12bfac
za8c6611d9e75f9eee140d3ebf6e1f64d7079dbc8145a0c692ef2e6c75de30e1adbc1f28cd41134
zcbd04d6e23091353476e2f942d1972c2a0aee8f9bdfcd404d6ea8b76c26b8e545f22477f154e95
z71b006d07bae6c223793d6291deab2182862457dad7ee55b57a9fba26e4482e1a0fc84143daec1
z0edbe5ea99ef2781f0c15e68340e4f8e3ab773d60982d130bc6e5b7e2c7f444c383f359e3c02c0
z33d2a8f338912ef7fec0754b34f6f252aafd7b5f57eae04491915f02f8681c6c96a999d9db7d49
z8beb3cecad91eaae5ba32a0e6c9c81bc8d24dbe09a56bbd982646a0006d12039725252c802989b
z69896122cbb30f5e1df1d85952439b91c2b8a5b563e70528ffa070ac4dcf981eb94e06ae319799
zd8a10c13f8841e3aa2d527b3656126e34dabf5aec99f94303c6b1b07bbe81edfd576b4cbec6172
z32b4381e984b0777e7042130614206756a0dfeb895b6f0c0e14a35b5b67a6a45dd5b15996e11ef
zd92932edd0716cc90b87ea1e09d56ad5d4deeb9e50d10c6e31bccdbb7fc60da1b824d92770bfe2
z116af4abc7665c5cb0ea433ad24461d432362ba8b2b5006ed334a84942927b2f907ee6de0d0da4
z90dd73586593dd6ef4ebc989a23d417b7dff194558afe5c10ea2361ead4315d2fe733682a59f2d
za9de86c63fa52a31a8d33a9a882ffe461691b6dfc148c8b3cd237cc975f06a39ab65295c25f6b7
z867db2e0c952b2980638146ffc7c2d9e628eca28503f6db8b0250acf5bc567579d5285cfbb6cd0
z46a07ce46e4c900c51c518b49b500b32167a02e7a035ad5c97dcc7dea1d1efed2f9dc5f12ed668
za32afa01fd480a3d745e48c445ad43d3452df4f9b1e29a5e4b95cd7f5609f7e60c7ec47b2e6d87
z4fbad9b003c2ba8c8026c1e2c14360bbe5eb3e459863f34748343c44434052fbfb8b493ccd5c47
z5d46ecf86012c14439a14335d495da6edcad465168bbc4d1b158f1f618200581b8f13f6bdaf100
z8ba2d4f7e9a453d44d9b79892eb391b0e01471532c6265e432a39f1b1beb9f179aba06281da973
zcb260c597c1a16557453984c2fd51e26dc832b282e128ff148e4e3aa5785093f9bd2b449f95c73
z906ec5e07edb419dea2b4e39b7da4c43d8eb2c97786f1391a2e3eac8f49a779439a22751e75784
z9892b9c162a8076e854b4e394332a6164ccc82cc46d8299954e72cce9def10e5f500f15bfb3c59
z62e352d74139a69b9dd0a2026cca09fe8d960d67f672fb6c3930e2d1130a30039ddd4df45873e8
z98d06ba2c9526d44028fb8eb093e5e62a2eedfd87cd3ad5d2ab6e16caed668c964e971158b4a48
zfe1ac4193dae4efc2700512fa4b66f3b2658881e5137505551e7b71efcce5e97074f446bfd098d
z038b1329076c3462b8ed8363afea4311220852a144c03adf3f38ec91421110186c4e5825bc0aef
z014f95c3a910fcafdfef5ddca7c8f26a241bf407aabf432773fdb4aa6372b75cc1d1bc386145f2
ze2e6c0af1d0847fb0a4f0bffab6bd9d8b5caa9e63f189b499405287875ec30dffeb341db13964d
z887c2ca66ba1ee254d20fb733a6d8f57e0681c017c8c9cd72f046470cdee09cb439438d2d8b05d
zfc90347631c76f78d6587e0d3b5f3db17ee4b84de1769a0238aaa3186cb8be13be3165f4ab0e91
z1bc56b01caaed291445929cffd8958cba48c5b276be1931e5142c9f64368000cd7a37a22a4234e
zb5519c7242ae5ca7390f876018c21df63a33e95bf4fa8edb8d8bf0a7644925fc41158a773692d1
ze70fab511fcd8b2fc680ed51eb56f0e816c0a5b9f9d0dcca84d8c9b9408a6f407572d794eaa4d0
zae48dda69740ed5b6f8273dbd5ff66d2dd84712c53b2a8916a2c11caae32b9ff74fc859c9eef1b
zadc857da7de8fb9c5870da0d492ba7d04016d46fd7a41b9f0fd2af19f8d577007e4ce2ea89f8fd
z6a3866b9ee5f29b4759f55b316cf7422074296349b85e9f6e8b9f569bc6dfab0811d445fb62ce1
zf2489fb22f5b230a5b353077bdbee197b0d24607e0c47dbc0107b2a289cacea5c017e69fed1b5d
z11a3e6fd8f890739a51ce2b58c5e51f473d2951ec3c13c35d4cfef4a88a8cc1ffb2f328f99b232
za64fe938db3ad8f2cc15129fef48b34487510b7dcbae37f9afcdd6d79e0c8e4c8f578756fc6764
z51f9407f1516686672cb35eae904d65eb2ee59c03d480bc1ed1a2156adaca3c19daccc04c630a6
z21426892cd1f9c6eb0ee7e98d8ab1039a23dfb0c482035acbb6adab35031e52f5ed84e6975fc5c
z6e25d2f5872593d18c57dd2ff6154079e7d144f4dbbfd20b0e8e262228bfe87a770d7576470c70
z326080ef204ccea67c2c93488f5affb00ff095d95b10f17e2ebb678d85cabc2da50ed81d867baf
z5da3558d30f377f62657d7c7e8734ed892c769c172a3c972569f549eba533eb091ba081cc3640f
zc11f58aa5351f72d523312e0119af51316f72d1bddd3c11860cedc473d35a05a3031c74b86f6e7
z1628197e20261a9e33cc9cefc6eaa7b8d231a92d084c13358229781146a706f4cab60c47ba10e9
z06626ced50c1e4df9c24eb488f25581ef7fedb9378280bbe1912cd0ab39bedf852323c3831551f
z8b75cbe8032185d40260e43c300e5848b4ba57bbcd89edc93760785fb89ba6aebbd2157670e2df
za72792a8ecabf06bc3ecae552b79fc1a1e19b33d9089d4ad802a332076a7249e4cf627568b55e4
z09a1a8003ba0f0a21ee85de9029aebe1f5fe05e0ecd8f00995660a881c6de63bb221e8212cc082
z1962226815d68197d54790bb3ebc7070bb1f8c28fdf9d142c3cc09d29d4ca117b10c606f13c896
zcf442163dce98343a94af1131fc6412c93793a5cd885fbdd2db39be832976810795bdccba8d2d7
zb1d3e0488ddd94c2fd33b3f8ff7d2c99c2b64b3cb0bad1365e6231b5103bcfbfb2f476a621b4f0
z281acf64cba24d69d7d50cf7ca91dd59745e9722296b65b762b70088fd51210f8b2c9b3dbf885a
zd7e87eba49d11de0ba5d1dd3835f7637b6f4186f6e616480017d7c9c2753c3c8fb78b0c69b76cd
z8928536e7de4732b16b57b289dda1a5adab1c0e287f95b46463fceb81ef6df034875bbb70e2273
zb80e6f46f7d935782dc4fbfab88ba5e294015b8a81a1a7af662859dd8617fee6b6abe1095a1d77
z61abcb55ce0e26e9cc71d04dbe9f6b8d53f7c2825ba9b12239ef57c89878a5959ffb67f8f866c1
z4c52bf0cf04baecfa75e691e6efa8383ed7504ced0e1d3ede4b0924f181a22708ae4cb405eb327
zfee24ef927a63f7346511aca96f27e56e595a06018db7190b77a9a04d732fe6be611b41ef2df34
zf5489553299bd25b9cdff3bac5b45c54e684b34da45b5b496ec4d0b9c1b1bb96e70109ec285944
z1caa876e870e285a28ccc84ed77e0ab89f01c554c570a4dfb4e7487d919fc8dd62ba62e0c7f8ca
z2a65c2c09fe3a9ff149e015f6a1333d837bf900c1a88ae21e93c251de576792d47f57470eda4da
zcacea5e6388fb41f9606e8b32c8aa9de9bd5870c971721753e0f4b7917586ee70efd100ce4e5be
z6c2f053231d391246081fd964fd3dd9ab77ddf2c444a722385c660e42423fafdcfd4f4f3040e98
z60a404a8a7aabb2e4a68c2e1429df3e393bdf99a6fc00cd760ba729a8513862add102ba8d9407f
z83ddc6ab22484fba355ffcfde101052ec5afbb6261cf0ec5cfba5ea7abd04c48ff406da7a489e9
zd6c9d29d4fb96875ec10abd2552bf0ec81fc62999206605c4bdb7b67fcd152ff6524ad6f3d174d
z980a11d4247ba2cd4522f29a36d5d54247e2ea6373579c0b3da167a06f5e5c54e894e852b45cd6
zca73d7435702600f5728692a0261d534f14f7cc25a9de258db4a0647a7b68ec0285b8f5e575a9e
zdeebb26735a4a8905bff41892fa626cba22b4acca55e2bb4494d6264206722e16362901146cb48
ze0932d788c81bd0e83b90c9fbbaeb2c20069ebb34eefb7fb5e9cbfc5e24043ae0e2d069c2ca0b6
zda2e5f1e742e4b6ea08524f12546f0170e79fff7eb874e99fd9e1d45e2c481a0f7772474e1346e
z7ef80457a7591340aa6f544621777db371d5839e1715c34db61042addbbc76b714b1e21268b4e5
z2930ba5e1069acbe0b3159f25a8162c25db24d836966d3fbb941b89408e460b769cfd778db0196
z88889f5da85086e0ea664e7294193f419c3c41c29ee7ac4d41bd23da83ffc2becd83ff7ae95cc7
zb1b9675ac5572881b4fc0ddae3ef063556c0958750a4b7aa95c047d04302078405574fd56b616e
zc8d00f0abef3387550ffa2c1d8451fa185fa0222c439eb8cb4fd6d49edd4648d2a7be8227b19c3
zcdb187212742de78e0de89de52eb398e1316136eb125be6ce3883c643955b1b59e843776a3399b
zbb60f5b0c91aaf17afe3d922c0e1325f53fee7c98d15000a206a4f0d14907564e81bbf6ad6b075
z6a864605e8b2154c1de95783b895a62abbc3fbcc3f189042ca770d15bb03b14c1db4bb94be57c0
z2a430e93881accdc0aa5c2695027d871320918c715ee16f5858da83f7e773af4877f3770ace11e
z57dc124e3ff6963ebce7288c3a872c9f2977de12ad8ceaf3d741a3059a6dfadadf10508418e5ee
ze25a19579150861555acbdf7d8070d055f80f4fcb0c462f8b75f055a4f5e48fdfb818a54c77a5d
z0801c7e4efdc5b13cfa65fd5714088d40427af91ec394ddf83fff42bd2c742b9d0513c41cb31d2
ze6e32117c840813f80216220648c3474677b78a0f50a29e61895911aa16d6bab5b3ce180709485
z79f4d51e64d3585f5165d20fd6426ab03210f3f8b2ca0b36064a7fce4193d5b019fe8af543e607
zf65e43785790aadfc2dafc46884fa974b46822f85713247a7b2270c268609b62d9dbd4c3241e16
zba97fccd03c751ded9d28dba9a2a7363282b883070e995414d0a3a46d6af3709a56bee7c0d85c3
z77b56fd6c27e0ad12f21485f5e9c977684c0d9b1f0cf68e390fe1ef8e51f4360ff4bacc058ef44
zb60e9cf28a35291da8ecfc0edea42472603a625021ce2d06ed483bfaba17622939f52bacd536fa
z3e48293b98eea13ef43bc707b35b0d903b7354c2fbacad36a18a2195ea0597897f65ba47020ab3
z7cab6fe5d261364e428bb3ff19018ca17e7b2fd07f89a2309d9a8740e1662f3e98b816853af2af
zc2143d8ca96f9c538697b0e56b1563730f3a80b834acff8f154060b3ebe8a3856e5bd0bb5cfe2b
zd4ff05997ffe4010b33647e830656d322785c9f8be916745122fc4a02ec28e601399d82b883bc0
z008faef29eb7174813e42d686b63bfb08f3cde294e7843d4dbdf125531c40ecccd971031e8311d
zfc74462347be2ce239261bbed228e2c15415e5701ebd0a4338df775941deea6a9248e09af7853c
z8abeb12c411bd711cc131b7444f8f4392520a18c5e7987d4391feddf235671d798f45266c9ff5f
zd7721c1741d90d51b95504b6b0dc4fab5cef440f5de21d01aba6339ace2d3d1314e4773d686dbb
zcd53ae805cd6b90ffefadbbc3d32d3e6e50ab24ee4c8cfcaf7e45e53071770e7303d3990a8e5dd
z268bcc5cd15f1b6345ec1f15f622f8a53910ef1d6f9ececee34ff5ccb1cddbf0c6983ffe4f2606
zf5868052a33fcc9fad4080a753d610e298a90581b63a234b4e83326f86c5433be29b6f77f9308a
z1ace0de9945768d985269d28d66a846a30eef0f4d8354e30b691dd506eac67c2bcb155c4e912aa
zde633f69a47657c6c3ee01cfcec07c2c2650439cec4c2304b852ab570417d683f79cb623457e40
z6ca00f1a33eb49cab4a66cce4380819e4e28c02cf8515755c6eaed303e23deac8b2293242769dd
z63d3f0d27202ae6d898d1a672af0be3f9d40f0f5f44eaaa0c6e620de5de1462bef4a7ac9921b11
zd07f150e80e70dea6eb29a72aac150981aafd9f040a23ae85a8b7348a6537852c1b97bcfbdfb86
ze79c93ec66d249bd230ec6f429b08440b05c361a9f697fc972b7d2a288e9f72cbb88156d504437
z708e4178d01b2f05926cd85e6accce264009966224fca087851caa7f40bdcb88fed802cd36c702
z79cc406de311b9d05dbcdf703e5372e18181329335353c15c7896ada44c92e9a0f13847b3bd5f8
z599c0636a99f4d65d2c1660eb31727f75ce2fc9abb04e0ef666193cd96872eb795b2ecb41ae2a4
z288a7996dc3ea501a933d07425f4bfb32b92572422ea2595e27477706ae79702bfbd8b0c8f563c
z129bc55cd9a9a918af3770f2935aa3fd86672ad157037403924485d5a323afa291d11d06a86790
zd449d80167a88ff0104f551090614ed40d9cdeeb7d35efc91f6398d721f16a4ed27c9910a65ef4
za40fc2225cfdc730b80f83a6556c5f6d80228c62016cc742b680b3890bbbe17e8d4e6a06e8215e
z89b97d9527bdc75cea79d372f74a11f07b607919dccf0f4afb32be12fa7096c2edb7bd07576498
z5501e07a85aac175e04b7eb8c3bb46625fe7fa0086920a12b9dbdaf42e8b1340dc4c91f71ad3b3
z74d9abed0309433fc140c3a43888b09ddb24687123e5f1b7c378c365bbf5842394235db060eab9
zf7db89f6f9cc94ebbca1511b294f3f7dddcdf6e91a5f042dc877cf623636eea00b59d9cd93ba13
ze1f9d7c20c1c3661e62bc2f5879771a147c4d7e018f58f7d61fcb19d6b2e65e6482878fbfd95ae
z287ec8ee5e29bdd232e9a70046fef84228cc1ed504974ccaa4793df88f229baaa10a2523a3678e
z57b049bdaa4bb9360cfb69605c401d9ceb289f94f909d2407d00ad36f468d5d7415bd4871b19fb
z2cbd3f8ed52a08a7e6c9c5c1f191266b58f3d6a9ec9493c95a6082e8f0f77793e1d209687f5392
z5b47d64f997074120149b1ddf125139f59907261cd464c1c85468201ccaa73099634e5f631a99e
z8a8945fcf6ed654bd19648dfe6a6d68e3a7d7ce5b6694c2cd3097ecdb8b27d39982e54c5590217
zb09e04ff009c229467ff8ea155e345d195648515c0b0978a4d64dab499105d491eb62cd9bc022c
z20b3ff7ba5861452b763e24650431b035af40a097170c7bb6e18207fb8f1639461e369b96241a3
z1dfeccd8c157871d7b41e4a4708d20cee698f9aa581eb24d58f88c12ea04eee84927024949ff9e
z717263903a39326e5135f7ccff121118e034ca4a41dd539e0cbdeaba09008654667bcec5eafc08
z332a6c065973686670de1857023c92bdd4190266c7830c8b4a78ae1986cca6a58eb6ae3aeb5358
z588562dabbfd49ad2458e73514e0d4b2ae9b7375541fae89a848dcf90ba8f9181b61b6baf40c41
z79f17e58048f6aa01b1ee52ec9489dbc9613291f5f2cde44574dae587dedad1f9d4c35c9c1d0f7
zbe70beaa50bd80940591868183546db1803e17b7e5882d3e18c4eb46452d4e2d1817a8f0b1b209
z3ce131bdd8939089dfa81f9d74245714f55bc72bcc41df2bf70d6d0835008df9491f6b0e234228
z2ac01c863d6125096f96bd9bdb93fffa3bc43d0ecdbe96713785765cdea2b9ba848b3b803162dc
zf6c8ccc70c58ed928525d9c27a2f0fa667752fb3128649d6dafeffa075838489d34bd424a8585f
ze3a52c613814f141ad10637cb1e954c7823decaf5727a1b7b63190d38f41c595708dbb395a27d4
z9ecdca61cce27549088594219ebd47ea4b1dfd9d6c0cdb58a986ff5279e9497cbaf8f8c5aacc6e
z8df5415cad72e08df84ab70ea3d06043dffa831fcb5f8c3c90d63d88d18036ecada3f64464f4fc
zae71581439bf290f9f9fdc2c05af82264062dfb8f4f1d397b657acc6fb8dc466163b279c38bac1
zecd9ebcc21666c48e6f8d47faf312574963b15b09ce555446b16efa40e693bcf6c1cabf05a7b65
z4f888e3a055429cd5388b75062d056bc37b93c736c84bce10aa6f3426e7fde13552a40df22d6bc
zee8be05a292f00d74d2dddd0399e8b8e269894ebd432ca2844022ac846d4b8db5067413a0d7102
z1d231043cb925c2c6753c25fbba476bde885a5abfef924ab698b0218611155ebeb267f23e6c935
z003538bbd977b45f27de475dfcfff55a70e2e2769d409dd1c326eca1dae777d524c90a51a1caba
z6df8b09959199f08632ebf234289c90f374b7903df7d0019afabd9f0d383360e55301d366d3607
zc256fe518c1bed49981ebb5868ceb19bf2c45db265f11a6812522e3abf9ebf2bbe8724c5fd57ab
z09d63fe0672272dd330c0e3eff66f0cdfee449d92156e25c8a4a5a6ad6f9c23f3342ce7c367107
z988d64f7b8b900a3ab55eafd9eaeb41868fcc69b913f898a6091b7ab4e1c936cc4404ea913f647
z73df60970d167e078e90234d463ee19e8cf88f88476737f7faf41078e9d853dfb98cc3b92d11fa
ze5b4b04a596842093ced424b18388cf96b43634542b5304edfd855b1ec87d3a766d571e48cae6a
z6cd1430031c247f35e17b0e7f1538028d0708c2adf0de064791dbe3c37ed66ad079e4078d3eea6
z491e57c5174c216be5a3ced9fd3867fdfe1e061c2888b90fbb2b06345d4927016b71ecc3e2833b
z9ed68562bcc85eb904e25d88fd299f45bac2ef284a307ca7d9d2ff575db433a89402eb787abd05
z42889e504093779897e0b3f63f358e5e3b0f033d2754679d3859023f7fb7a583fdefba0c815efe
z0439ac759990dc5df37df38d993b9a41b1bbfbbbb0cafcdb5133bfc04c65451459f1d629911e1b
z7c27b96bf2aaf11da4a2ccdf1f55293f9bf8e2f466c0b3ac72a3e97441ba478e786e50400b091c
z3daa7bafc903a3e4d0cdfb979f4deff41bd2e5744edf93fccfb15f4d12e3771009dfa8f59a56dd
z567811048ec4773a95376c8dd2b28cbbed1ff01b8bd15768b1e32273f26e7d917069f0cb4355e2
z57d25c390eaeeb4b5bac317e2fcbdff19199f5c716dcd7cfeae8eb417f80db836dea8177a1aec6
z4d7573ab72d300eb55471bde687c5f7be2fbd4a3c977eb500b63895c818aa6dd89505892190b5a
zd36f49365b86f4258f4c254948a90eb4d0611b1ca47bb2d36799a7dca7aacf1f593f8e98183a0c
z2cb5eef613134a0c794b1dbac416078731b4474443ee5991d034e79c655152e51edd6b76b78557
za0829bed7b32d0b854724c286318b83c638373e84fdd0c7b47f4b8035b3a35db9f9f49dbc5c011
z02919e85cc1f04430448c2b57c7aeebd7d0a6f099d439299865a48de3dce38fe11824288347fd8
z07a7a8028242d1e0eeb344f5d03b2750929a3580a18a7c38d0079d4b33d304654fb3755dafc851
z8af056df3479d3ac838e7b8c697942ab0afe6c4cf354b6df4388cdcefca47b26de7acd4c64730c
z2e28eb1ae95e134d0bd7eba02bf394afe5827a4b9f347a0f9799e699a90b1fe14fbc9c3a0bed71
zb41869be4630b857082598fdc6dbd5cd2459df22bf6425e1987c87bbe3646f9a7b283979e428a8
zb1207d3d557b5d349743842d277b63394830326a2d98873ad0ea466dc11e5426afcd61dcc2edc4
z98455038f922de43e0424fedc0f97490d460f8696c0e53b3cf12f578e0deb7df2b9203d471d14c
zc0de5d86a79f8f977fb3ef3ffc2276176b6960fa86873145f1187e4e90d91979e778c8ea872dc9
zb42bc2cce494f9e933c76ec36fc1097ef5dac4790585def2f44b9479b75b329610844ecbe5b4ac
z983a85c2384483f187f6aaa2dac1debc3aa70f61cd48dae541421271f09f292835ffca49706483
zbf8c4140198d562630af46f3706df048971010535617816737bb38838947654b774eba1badc917
zb58eba6d31cf0bf68a8380b59f8e91c968c9e720f053ad4eeaac0f99fe95b1a36ec62356e7eaa5
z97a16e2f002d445b3e33c6d32f4944136a07ffc791e836ca4619b46973c27b522dee42c090adfb
zb3ae863102b382afde9a3f45a1f7baf8fff7326b770006a50941d29ce889b19098c5d0f66f5d76
z15171d6b40f280bc50243602343bc2d59526c14afbb244a1c02df9e3d9f02c62aaf0978b0a5384
z33db09cd59e82c5a93647b6aafd48726191a6ef75bdde5247071b48636a32b2cbe08df9492a60e
zc4ad46f1ef88815c002a6b4b6d81429b70850a3732adaabd32e766c6a59ec64e3c02810bfdd3ce
z81f8a00243180e37e7f19d9059179b4254c8567c8249c1d9c30ab138e7bfd98fc74aa12c897452
z551109ad477f6dd769f545e27f0f707a14955957a396b897bcf57a6a29dd31233808f2ad069da0
ze24d0df664f909266033bae346159904cd4d4b8b74028d07b28ccc8085fb63cba63eb09aa6df49
z574770fca22c1b41bd0f7dfa8a9c92965194d085a6eb8da99795998e34e1bf0cbd6f8351fbeeff
zae65300759247bb6d63dad3e3e5d0ad1bf00e93e09123430a529818a09e69a5c2b0cc0074ad848
z213573032ae902847c1dd7a597d943e31c283740fbc1c4f126a243041e6ff72a5c8ccd8a032030
z46ed9f9a6849f244f70a99d742876ac43fe3222e9cbac77b6f5aceaf467be6e5d99d5df22c1a75
z63f6e28f15ef7fe8e90f7863e3a3934f0286248ebf7faa320dffc111f9b3152758c6f0401c2da2
z6f30ef113e881598f64453fe206b4ca48acb3c307bf9d97295a18b9799f02e6a0b63d7e94ebd1f
z42b9001811e908890f91b931ec7777a7e988ccde679bc6e5976ffe55b49a34af0865bbe6bed749
zcc2e86f2ad764c7063a88cda2b289b8c224f8787e3a6c0fa20782590fa099eff65de6451953893
z4fc83d2c6639a1f2678eaf731f2fccdce3ad77a3b87634259cace00ebd7c55645fe08d887265c5
z3e777f30fb78fa9ce6019b62507ab348e30cbd3b969c8a29b4348b52ed7a38fae0f6ad1803f1d9
z29b6612024c19fa7a96419a34041995bf95f34b5b801b0a56a8cc4564d604fb3b66f38f0963b7c
z69548e2199a0c614a3109cf2788db45972042af9d76fecbb05b404faa07c5baeff11e2a09323ca
z2ff1165cb3902800e77114b20c94e1e204b46b8fa2f79463ad21ca4979ae57e956c1797792a6ea
z18e04e94305d38e87edf795dc15155d543a3312fef945e595f65f7dd11dd1429866529a55be011
zc48d3e0d1cb18fc8f8d76983fbdcb185c47630e015e1acb3728e7f6b7ddc8ff28c7e42f53bc2ee
z01b7d0c4ad76c356a621d8a6f141be21790f9679014a28cf36c435c04e2a81e5fe79572703bb1b
z309a3d33afd7c0f21d0a8be89132d8784fcf26707695ceb4eb4994a5b817bde9476db081c59b83
z4e944576bd5cbf9e8f7649150cd09de0018a4d7701fc8fa54bf70df3ec9fc928755d92e72df5a4
z15e52ba825077ff8c987ae4fe065b0400101aa00fb6f9d31637efa770eab9961b1fc224735b59c
z31f5746869a9b04363ecafa2fb0794eebc94dac7165dace4faa87255e4a9135d659a5d36c4a13d
z462cfd1f984d519ba16802281d4fa936016363def20d253adf8b1d36a96282a2a6af34e9165d05
z78091362ee6e961ee7da3e57e84c4e06f5a9bc353555f8248182fbca3381f83e6981dd64457ad8
zcc586f4fee13e4f77158dbb43431de9c66ea2110987392203910503bb70996401f101db947ae74
z1436d3e995d5a51fbdbcec5c74d5d5cbf0170dcb7fac9619a9d21a188e52922237e680d39b6e65
z9a1cfd6d0644fead940c9b2b8e19118c6fd7dc9433c1a4d1dcb43d835e629391ba84c55cc14dd7
z96f7f775e1c5cc86c1923834d35e6f05fc85d9f06a56cc35610e2b7a72d4de1bae85566f213c0b
z37b2444181dacf207a0e0ea8727d4810a1bf1f8562511b20650288e6a92cf52225d340afff7f7a
zfc995cb6ac67fac327505e73339dd91dd68a0e19ced0b3b501e85d30ffac351eccde3d33a07aef
za22155e20776317887b85ec6d9de9baa4692c27ebffb7d2c5c35b6f9fe6cb4d828c334a993369a
z92b2410c3b02d1e94e65227b9c123351a1de904057ca486f6b33ca6c1c85953200c63ee0238f37
zfe27d4f40fab5957a100bd3bad1063070644171dd05ef8b462a6098c7cf6d239b5ec1252eab449
zb4886489b6d7e0709b63f80020048cd228ea9c95a6d18b03079a7c222fece9ae7325fbda4a5bae
z8ca2b02e8ab615afcad8e7670a6400493ec2287855de515b094fc1808c84e595db35bb2a28884b
zc4d12800f3e2110eb164deb49eae4c3f660ea4823fb417f1679a9a7c14083a386547f26be31510
zc4795a9b1bf62cb687224ac26bc07217f9848737e5a35b4c37d7fb0c266cd6d8b0a494a9b0424a
zbc958910124c21c0e76d7eeb67bbe58ffbea7a38512eb793f0410c15162951a0dc914348d77fed
z46c43581f768e3947411e0b2a2e2c278a1465e1a11102349bba92c899c7fb518b52fca35a5c4b9
za4f636f25e05224b75fab4fc3fd05079ab0fb04cca7f62f34e38913a59350260dd6876882d85bd
z4c617e612ee60b224435b9aee0ac100fc4ae685e2bd5ed81bbb18d01970a67393d4b307c8e7873
z0da4dfc6ac14630e6070518b17b9be512ca1a14d3b1c09c6cf56eba02b3b897b0c7a00034652cb
ze403f426dbb4244931dc51468c21c58a90eb7107fc73fc58744a3fa9b66d72960cd6118ad00365
zd1077bf22c25179d22b6b2dcb6c5f639dd3fbe8f02b0fd1dd825e26b611b8e3e15c7a6973f8e64
zeff2163bf1590d327dac6a45693cfc1a982e701aa4ff84c6e8ea9b6e556d2ffdca9c9945533304
z688adbf01a1cd4b64b445c091a4751af654228b4b6e7d1f45e3389f8939370ebdf71e2ddfc6420
ze9356b7bb5cf1b117158b4adc6428d7ee55cabaf61c412062d384971023e79ef7a96ac29ce35bf
zde6eff9dcdc6198bd27559fe0bfa4b606cef69678e99193346b26341e93ccdea2a62389d67280e
z2010cf123f6b4e268ab5271c574699b6a2b23aabb36255665b492bb0401ad21dfdf3b540035545
z6aae5dcc2b3196180221e412264dfa99f1b03671cd2a2e0bd24b0df550c0555804dffaa0aca550
z64bd3336613a03c445062e7ed002259898ff74d71b7bdec1ff9ad03973c40831eceeff9d57843b
z1685ce98c7d9d04e57249def7934ab90d599128e2abf4924a4eafec3346de46ba9ace076d0deb8
z62217d6935674bc1a45f1a90095a5599584321a3df3751757808e1616096c5584c4639bdce95dc
z5c0f05665e08a0da43a177c578e60474e335aa4a69175cb02ee132433c6f911a5334d129805959
zace99c7e9cc30d9f5b39fa632b7d9f9beceb7229679ac92760909497d8df612113776048d2798c
z42a045f4251d2f5dbf8c442e3b8842cc114c8533693ffdfc8adf4316f0cd8961e25fb6f41ecf10
za2d32442b9950832ad6b021f08f205542461f25837089a8404823f60d656870052ac71903a7bf2
zd7e048a7cf441106e441cfd935e1ee6f0a7c1fbbb7ac80f1248485fbacedc7043b12a697ed2485
z5a708316680c50b76d857ca6aa27f0ea40f0337cdbc682982d0c2544a3a3ede88ac01fbc9f1a91
zeb6ae71b463b47c37b70ba1f66c2dabc792a355e7ef4492f2916cc9d55919eb52b3a98714ed134
z487cd1afc2f1c7dcf5e22da54781f8dd314792f62f6f21717ff3347087ec503cd48241f3c6f08b
zd51f3b903bc4e9bfea6bed84339a3b0f87e03e1b714584ec2072b80bf70f5db00d19542c91c6ad
z53cfe0670c6dc45f967cc43dee8966451d2f07551d7dcb760474b270763bf1715bcc40ba66475f
z8d7fd1b11d64c0698787698700f1572d0aabf1d6cf517f26a3fe273c2e7b39709cf25cfd265696
z5cce038912779e2d9507b8e275231bef6302166a9c04aa115c94e88d4fb47744583f05b15f9a91
z65d42e87b5d72f59d8e97e9bd61b8e4e1ccb769e08cf9be3276911464c78c963174d6225a79ea5
z50b56bb76044221742879b5ddb811aa73e4fa8d446eecfa50c2197c851d023973028b86e685d4b
z9cc92c7f31b9949be8bb452fc091838d416a47d84e80cb390d29c7186ee7f8d959fe57b7534226
z33fadd19a9729fa35cb4d557f50c2dacd6040b482c9324436476f976f571745f88b9fee1898004
zbb68dc6f7267fe8eb743772ce67fa4b4c98465856798b77840e25ec362c27682974ba5b1ec918e
zf74ed4291f9e2c809cf02c60a37931c702b8356943baf21bcda254f13ad74909bb52d22a9950f3
z279921041426121894a400e6cf3519307a7eb6ec7bb17574c2d1f6ed4d74e3e6431f1124d7f16e
z45ba42b08aa7f5c2c76a8f2ede1f2c058fb89ba4d2eae9e762c4ac11696cdd4b61628234d705dc
z7524caa89a12c961de24e242c6de6953e7e88a48f418cecc61c9b31d93700cc06975e4c0caede0
z17c4331c673648c0fcd36d992e384539e0a430b7fbf5f932551b6c82ee2f5b451518b98a506033
z1bc16825f524cae2a6642b733beee4fea29bfadec21cfe88ca741f8f1f5fcc98441fe1a52736e5
z7c96897a43856d50c2ce45800b7d86caadf1406e5bcdb59b0108b8fb9027ec06955b676a942879
z0af430fa6f1825383f17c19f2d452c0ffa7037e31567f1aebe6677928eba5ad26d3a1733394434
za148e0e2cb9db84ab568a168100303ca70ab1d73ce71819d5e62d817f6ac4797389b91826597bd
z1aec80e89bdd52b35a6685ab6ac826a196306346085f85de96c93d327075fef24f0d45a89f7f00
z2d3ab4ff7c8e830c56b2bc4b8d68dd75fc22b79c47732ed3eb6c2bace1d28bfcd7916f7b829e95
z688ae01995ddd782d1763083a3b02be68424062e18fb325bda53799afd6c1ddced009fd75b89a3
z52f503424af22b629e05db92e32fd9d5f6c5569ef75a2777645925c3ca0868536566c826b8ab51
z4a906edb5f497afdae2559479b8adb9b8ebbe5d6fbe5af047a7bf0f9393bc71eb55d1100df1e54
z10a2911ac234498a814954168bc3ae7f93dfd041e429455e4c77ab1d765e58f019820825030e6d
z7fde13cc648ce91480aa12f08e2e47478342914c6f2e269aecc019eaf654982354f0eb580e2a23
z1591c51e41850855bf2c84180ecfa0fb58caa619e61a1eeeeda670a1b6e7cff47aa1c288737db0
z4376a8f734971a0247bd9a81fdd783749106aaddb607528242b44697906e776254bcf484aff654
z7d3ace5800f2026b50aeaf3d0e635dac4fc77e651ba73fc091fd2537ca4e1f294749385826e1c2
z23323bd54a967a7343b1e1b447e4a18d5b0538e1153bebc3f2a953fa6b51c0dc50abb2bab8b951
zab839d8df8d3c1bc2d3f043484c66e241257754beba0d557106fcbb50a24a5780e9beeb6363f3d
zb5e818f6b0e312152e18719f557b09e2a95c7c47f487851834963f6cafbf9fe23e897d0906c2e9
zea86fd5dc3be0db059d11045261744b47b3ead51e541d1b4fd46baaf169527032893628b38f550
z4e2b3b9cfcfcb3c28ef2a7b5bf4209f0f6c24acdd218f6c2416fa597cb17c9c4e8fe68de3f7e3c
z09232955e1a1bb70e19de02b230cfd2e18d1a162b8d0e7bcd4c3693be5d0653044118000bc6208
z07bf315c28251649fc2c7ec90bd68f78984a489569db143beaa19b34579eb7af6e5bace5f0f8cc
z946057948593c7d192f75a0c62a38df2e9972ca8a4509203b03178fab34c83c96862878d872de2
z585abb7709233827b78fca51c5f7d9954a3fca10c8382d8a597baa5b28741beeb2889ed36d9cc0
ze7e5ef8e82936a84cf588e2ef9c2139ba999a76597b4d7fe76c39d391e8be9ad00438768a0cbe1
z115d3621d1b325a0adf149fc1c967cc0d2b11d6dacf229a31dc34a6f3d5d0c3b71f87ec8cf53e0
z33effc06a183314aea696d34fd443f385b22b80f100efb8b235680516ca70a105e820d463c4649
z72899b38ef6d42b8f112631e773c397df1bacdd0678183f14117666f55fb4c42f5250841c40fbd
z8e425affd777b27f02f20b8c953e99c66728a4b03881b87333bb02af6d67c609117d1e8b5b9bfc
z91ff9be7e8bcf54b55b8b933c56f81cdf3be2e39e5e4f626c4827016c2effcacbfed428f3b1148
z8b4560388ffa5acc4855116f53b20e3026174fe33dbfde5d86017f02814068c003f8e927a4b6fd
zda5f61c89d4d364e036f942a8261cd5cb1c2399e98cd603ac20b185a1dacf099be4aa0c07e92ec
z62d25c9142d2d7dbeb7dcdba9b6fac48076c834c68e47ec9d47d8a57009252c8ec4f65cea0f8e0
z48d19687eee14524bb7d52dd6b497928c1e561053ec983ffaa33946a429a92bc4b668395365cd3
z4ae76519bf4e02fce40d879e36a9e28fd1d4467a328f61f0ca782ac9005d207bbd60494041fe65
z1ccfd239c09fa787d39a3e6b44dbae81d9ee5596590ffbc9b6e10c4ce53c18b52a9bd37d5cfe7d
zedb6f96b16a7e61b370fa286edc06414fcfc3bfc0aa803d0c7196ff9b8221e3b46d859164a15d5
z39f42e180508581e24f92a6523b8031d86acffbf72fd1bfcfcc5b434503f4b7301f45ddc84c452
z966e2a5ded2a43954d6f75129a2b2c3cfaf491279ddec86d2b2883755f1139ed0ec9bd4e60ef38
z015518a2e037185e599389de7653883cc44e5a49755957e8f0bd431ccc04038b0cd284db08f24c
zd38b4d25ae55cc16d8ac9cf22ec1cac7fa448071dc81b2dbbd8bb5e2bf47723d11712ba257e3ad
zd5addbcf8a757e7f05e2bf11b2d9d52394a7cdaf76b5ba610e9446b9a07ca64bac9dd64e3d9d0c
zb8ac76166379177365381bd1c1d66b453acd2119f1201249d6b8922225d6242f31e8da41fd5a5c
z187eeea5838a4746ab0e990d60ee254fade77964ce41d94c44f97b9eb80562b8e3f09c834f1c80
z682fa714a429d08ff11387371e4c6dc26fd468f5952666dbcd3e9dafdef2c4bae08814e98dd2ef
zbb63c7f14fd823f69dcdd5ad7ce1dfba1fc818b40c08c58959943112215070634add63b932daec
z40d47e791b957dce9270730acc72860cf4e15788d05565e067dd04dbe228c02a2de77d5d77f522
zd1ff3661f6ceac6f942a38ee16e01561b49922b330d5538265c58ea50841b889d73ea8a58e7549
z167e5c5aea2302b52cb5d4a8edfab2aa334ca5660af0c8a0068842d90f3499c248f006aeba06cf
z787f0647f047daeaf15a465ff8f46dee52e218f949f16dc7d25f63f512145a8d9a8ebe2e7c4c6c
zd3a8daaedcf0ad24870b4daf0edf27971eafadd566b8fddd9957f995c1a6c77408600483c287cd
z4d02b24d9703a84a3aa97ca9f5c597ca8c8b93cde3cbbf77688a49ce9b1f1064c64e378778088a
za89bb03a99c6858ba286899355f0ac2212713d5c38bec52eaaebb821a97b15f495137bc30da7ab
za5abd09e2401f11d3db1b237f1c72fd6f710a99d87ed158d5ea2b3957b055f643324e3724087a6
za430f2c0ae756f2cb71a3f431ab18bc75e83b3aeefd07d58328f2e90133d21e9f93f05aa5c9ba5
z365125f289132676900dc18a6bfffd946d7f7fe49eaa6ac6066da4cc4e561897af2411cda4f93f
zeeaf38c7d7434484346de09055fd97dd2db4d35cbcbc33094bcd28d87a432d3a90b591e5ee7798
z889024b5c8e5bff3fb760e350e8f32ecc51bfb337d95f6794edac296d7eccd5a98141a01c2faf0
zb5432e8498de4fc840630e2ba75841062d2c382748d38d41c494aca658f49922535bc0ca213e33
z1c0cc3231e31340f091fa45a42cd9ed79fd8bb44da9799d9133824ceb2dbb1ac004a4bb7076494
z097aeeda94903668f1fe2a3ecee3e0abd68d5acfdaf0e7be5a3eaa4c4245805331eafd5701a56f
zb9dffc7c29fe2e743163ac238684cec80c42cfaf1711f7d2cd557c9ef6d82cc2ef1a84ce3cfae5
z050f59c2ca30dcad18ab4e9a7a3dd231584c33b6fd0cc08298a324a8a6b430ebf9ce567154ac53
za6216b29729f126a2ee53250f82d868e0d36165236a6e5363007317400bd674e3547c1343be51f
z4a73fd55de4413da62a53b93a7f553a973330521682cfd6d58e94e6284c546db81ffbcccacfa98
z040f5510af84c8a9540c206e3d7ef56e9a84263f96393082131673ba18429c673b16dcda1b9ec0
z56d1078d08b3a6eae67287d6ea73d289f7fd0d590e2f5ddda05a1593032d681c9c79cc590e9d59
z49d8dce3ae0f378a6639374f3ee83e0b6e8a495a720a16ef4df32c0a544932db8ab8485ea15cca
z4288a6442c587b73ea808f3e67940917e96fa9ce162b8aea7d5dd6de3704f098af3b654d657747
z17e4341c629518523f00eb0ac32037e7b616e15d4215d51e6f16f72eec95b9d22771994a731065
zdf6d1038b18c6d2b9aec61a864a3cad47f78ed9bcc1eb5845c0ec5b382a758ef6d37fe1a775dd0
z42f48aa90f299881bda0dd352eb3cce77536316ab1249ab27c97f885f732be68d6ae280bd10e31
z341edfa42f3cfdd28f8e8734d44090c4d38344ed72fbae50827efdbdea076250e19aca77e4e89b
z42f086dd01c06e4758d301ada5add1eb61bbd6171c6d0ad52a48cd76121aaaecccd2ae06886bbd
z9ed8fa97415a8965ebba149e733a7e341960e4418f4103f516bfeafa6cfe4abb0cbf5c63e8a77f
z6dc8b1ea08292a7d7752e44d20bbfbf9b7371fb3a12a0ce8eb78a61931c4d403f507a6deef3300
z21b3ff8aa1fea08b4699ab6dfa97253e3562ca53f97366e41d539fde4588f56bac774759571ebb
zbad78b0f36f95272f82e913ff20600d3b528947e2b752ebdf7411d20e62e420781815d5ab39a6b
z828fa9e1f01d82aedbe339712593d86ad6941bc54459ddec4c217c739ecc0a587c8fd1e9ef37d3
zb5c366ef0648222a062916a86dfb987bbb8546447fb18e487f9881d582fdf3a14d10f58cde02cc
zf994a84c12d031e99921c8bc9f82985b13e4678d5069752016697576e97056ce653b8a86b2620d
ze31609aca7218c70d3fd3497b727bb1f0a936aa2d62b2687052c2f6e87e0fac9de8671887bc09e
z3986d4c4cc461e9b51043d0820c7b71bf4bf8fd8085b32aaaf446c80aef93608b8ef124d123a0f
z23231a6aff07434038b7dfdc2dc4266a88bcf65765f021358cb9cb960cc12a8e554e0833ffdd18
z71befd75fefa9b516001d3ba1df3e97c07bced3bf79d4c8cdb1db5fb2d71ff0b83562cb50a79c8
zb2ea354cdad54deb66c6c745142ca28650b6fb573cc5cac7865fa7173b6ac9b7ad0ddf2a93524e
zcded802699454aed5e1418c05d2a9d8e2936cef96aa54bbb7b9acd7e23ad1c84a7ee4d75d5135e
z4ae8893a4422af4afa99518efb313e00a74a39823f5c32437e34f82b5e3837e28b99b888a663fe
z37d24322c57c7eaf3391a905f04a397538f95fdb0d68dde0c5c901349965759da5c1cefd711bc7
zde857b709540f92ff7c5315f8d6dd1debceac2738a323ff04b4d98d0a82ece1996f84877bbb776
z9945192fd6f8a9e9e8fc116a81509531144acfbee7e067a785ddb45182ae1435dde7f6a27eb200
zf09b93fbe35feaca1e6b956f081b7802f9fc476dacb338922af7fa5cc329b1d4f90349e353b062
z3491274af7ca9df78f5f83e6b60a2e82481f3e2b9d3f8164a26def0c2f9021e6c33ebe5f52f3cc
zb896b061d0be56c14525fd9d503b1740bb0bf6a7754e9b08210317946d2d3c805f6f2ab53562f9
zdb53fbf9d5ba623901a0449c3a0c1d72a5315952c7cf42b41fce45afcf147b234076dd73bbd809
zc69d40581e295d27380f060ef9fe4a477d15a827b9436023bc39b826b67877391fd88ad64873eb
zc5d35e11071c0d471df03ee3baadd4b4903fd047fb8b0872c198f120d2cc4d8cfb62219be244f7
zbd33ca0fa602df38a024c72c58230854ad17ce599b292ff17759f3fc937ee4845e5946745f37a5
zc644f58fba02cf32167da58b65ceb384f7cb0c5f699c7a3dcef2e22dc87ca3a36b38100b38a871
z6e7053b4cac207467aa0407272ab5502aad569aefc2c061c8428e2d265a47572d0ef69716cbc06
ze139e3ddb7ae7322e502d7944316da2e376536576ab61bbdb4e44a5d0c3e532e5485ce23efef80
z6083fce15e7146bb0918fa5a0c1b01e1a9563ee432d4c6015a1262a7beaecae82037a6367d3f54
zd542094b07b82ca91bf4977cb6804ab9c9d80e84c28f387801534818724140baef4a94cf0e8831
z179e4cca13c5475e390704fd301fcf9c49be8c2d15ae220bcb6aac25a87f17626df16c5e02745a
z6c192aebd043d24e0ef84cfe0cf97d883f2b69bf840e2d73079c1b15dd781430dec297d2fab190
z9cabd9f4c0963c05ea08f2a713f004194d2611c335d8b3dac1250f38a81cef37fb2c9f4d44adc3
zf86b9bfd5d2ad5f83ee3affcae0f4451ee3da46a29febf9f17cb289611daa5aa7bdb1d904b1574
z077d9adfee902276a72b56c2a1cf1780e8ead386265736853dec6182237d18bea0213113b1a34e
z546858e0bc4a099d289f3a8c75a09282a784cb451ed39fb877f233102021751228bc69a65f5b09
z3a6841c746955aeda9b44fde832ac14b1e3e1747fa6c1e634e6cd5a8db99c17f9c78f1e7bf42bd
z8fd9b40ab6e54b4630bf307aa361cd77e4d4ebe7341082dcc73af73948b4a04cef93faab0d5148
z57c1aff74a8984d9c16ebcb96f36187f1430790d7a16c620d6745ef0700c0a82ea02fa1073f3cb
zf6441579dbd2a7ab425465d6fe478b876512b0a977a00b0589f29bba87888d4935f157769d56d9
zde3fb599876926012594f01ac98f04f085bb984bc30faac96ed3a404a456f51e57d833fe86fb96
z81f45e8ac1b57b175770cad52f3c6f1686045353d6dd3107895fff49850909cbb04ded11668391
z9401d8f893e718fb842db5e2e7132b59f524be09a2ec1873c940e97dfd0e8390dc1bdaa32cb41d
zdf8a34c14dfeaa7808229787481dfaef577a2c7579859c92a8a36acf2a4c6fd2308dfd784acd9a
zcdf5e38873290579359cd7442b7be66124d59a7f931f98670e845af19d0a233463b390dc2f3ed3
z17d31728039975637f4c22b03a0e7342647f17c2f02a9224fa0f860e21add1bd04e8b8ee606c87
z6405999543854f12a93c811ea32baf59a3e8133697e4adb1c122e6602e839d5667952eab34f45a
z602b11c9269bedc49fd43ab0a608a0a44da5a7ee60f6985517e90579f2e70f46cc933c5ff4014b
zb3b10fe54a5482bc1bd91ba37414b07eac3fb039c92342e7d04f9cf56a47de1d3e23b14b86ccaf
z035903b5541b9e444c7c5c1f653b6104332ffecad84cb0128c7e677aa3bf9d18d1b714fca91837
z6bdf7143d8d33997cb2eb1883b67a6195b2d28af44067eec55e220f046d8116d40a0e79be3ca8a
z24d18af95f568294e379cc384f15f4a504eadb963afbe894202de4bd6aff3c73085e31cbf086d6
z66e836507b24dbdfa48201413cd84c953ad7800b448d81170a8e881120c034c21d21079b34c582
z1c626a86f3e2de70cdef7ff382c435b0da6bf26c8d4fe45ad9badffe9ab6de48ae49cd7db39b6c
ze7bbcc214f40338ad7cf648eab3294b64abd3d9d71de92b5eda8d3aef1015495c08cf29e02080c
ze4ab5b1371885f343d76dcfc364c743d3ad46ea3719cfb9b6a9b9bb0f965ac43caf84a7bcb7693
zbbdb8304161a98354de2f4dc823868439842175791a12c1bd6260017620a14fdff36be135c7bb7
zef9ac6095413eaca4cd2b7c7ee6d8ab77c0cc51e12f3b3786e7e76d2e401f8329fb4550e47bb0e
zb27a0c6e8e80c9ec83c693f368086a7e1af7df16f0289c62a9e6ecf2178c1df1dce882d5efa8c4
z6c6e1083b49103ec12e15e3f7e9422e91aabcba91dcb31744a8bc107b51935ee21bafbb9a41520
zb33efa04f7543bab42f025727d25e6569d64ab048a6454542135e62e24902e752d2f42d286a77c
z5622797ef3997c35eebdca8d0324ca26a36336fd750550bd893ecf5f59bc40eea81f83e51dfcc0
z92895c40a9f3976f1dfe44be732958b01ec2d7644c1df894fbee692aa40d79bf43fc88f07b9994
z14c39f7fee1220abf7a4b86dc7c0afa25672c252ac5e75dd2fc356b1b09cc15b184e26c0a85c1d
z3632a69dfcde61427d15c340faa101ff471442e2e459c260c5bcb2413cff9570d08a0d7405aa4b
z0121385436a566edf1b844145807e42aec896234e434177fc17238149337d669c96865fbd7ddb2
z92714697c04183c32fa56b326b42cf497bb0c91bc312abc543e991c26c7333a9a50e271fe9875d
zff48ba365703c3a862867c0ae157da8d423ac7de296ec2e85a7972a17ff739455c7a217384c9a0
zce1c2e70b3d8631d2a2723a7de55e59153f47a02254aed56a021a6e6360bc7f477e35a511fdf4d
zf013a6158f2a5baacacde77df7317f4efe2057f0027eaea96ed201da2e7e1fdf0f7bf37856bc5b
z3a0e847422236755167d7b51f5f94e4e2df87f078e65cc5fff8ce875318aa87f27bf4c7ec1d8d9
zc94e38db76ed110b136524838f8f5c63409ae312be43949e8160a650bc5e64fb2331130af11a37
zec86295e070293bf863a65c82c3fb83888e8f62d9a336e7b881e8fc6125bee64855c24e9a88d51
zc2b6453c3899eab2ab771288535bbb36ca4c36f99654cfd371ffab67e6318a4981d9a6ef0d590f
zfe3b3f5abc6eced2b3061c92831beabd26487431f411a22a386bbb04150d5895b550cf5e4167c2
z6c467582a6522947065804e017e5d146a71f31912b8a9bb85b4a324cc301fa140d81529bda1a4c
zafe5b61189e6c02d60241cc2b852cacad830ef5bbaef50417a185ad87fa0b3b535229a4711cd0c
z9dd937ef57f99df63b1ce792a9a01c78f1df4ec0956a4ae7ed550538580ab2c118783c2e3cc776
z602fa6cccd8f6f6952e75ee538c0818e4716e38fb65471f83b648f512153937cc6c4cf94e99d17
zad5b79cdf54fe99c4ebb8f679667e78a8745fb53d59b8991d044a99a10396f115d6235ff0a1ce9
z592e3ac0e875fec91081558baaafe7442d1d686026936ad8282c3e1e9f2fa9fb49b1655a1b2ab7
z423e6eb08502a6fe57ec781b06bb6d9f1844f5b5c4c3fe1c4eadd40506a4ada9f3d23fa17efc02
z9c8d85e6f61492bd5f323eef0daf05cdaa2d79b7f873dc0be764560483fefb04d598681148879b
z044573915a649f392e522051f927498835218c21b529f32710addc96e9904c6e90f20b67e5867d
z380564d53468ebf046b7ed545ab9903f3ed442649bf29181260e5b757dc34432237fd4721d5f8e
zba19878e5d8f49a9c86f8fb6391c3b322953fd421e59c631a1331cb57e3bb3fd5e701b2ff7fd8f
zbb3fffa23f66c76941631746efcb564762da1e60bff30f9ea946a2b8bdf4657d56e5ee0c46cd13
z5e1e00ceb0ec42762f1acfe7811b544a2a2be7e1e2e4fddd15c5fbb85b0002a5357ee6d1cabc5a
z23b2127b0a174ec9791f487fcd1ad0af5c61435bc9f11fd7d4177f7b5beb902f1efac9eb15d3e0
z1d47d0e60051ef50fbebf6f61680f5fbfd9250ce12817028641d86ac88d616de943689f4a8537f
z04fbf53671ab2bbef5cb27b5c5dfe71d1cb7d36f0da3f980f0f7b8543e253e57bc45f3e189a4fb
zd82dbcbfa80624dec9a0f319041305c915a66adaf55d6fca499caadd5cde0fcb9de3c963ffc72b
zcfd4373d702189a4058c9a956ac2bc7e55c2d5d24b34a1a637fb6affb316902de8071cfcd286e0
z651dbf68c047572c1fe6ed3bdcd3a9a1ca866b0e6eb4ae61d9daf72d058ed64ee845e725d914fe
za2eb60e364bab1810e80b27c4d2e2506370de0baa99d73060d48ead9ba491dcdb1bed1bddc7f90
z31edf94241c0b72fd89802605b485b1cb2458a7e0b57a1ef2f4cddc2c8ffbd61064d3b15295863
z088f98ac1d1489c38cafd2ca26b98ed80fd037832abd8d9e83bd9f331b795918ba5a86c9931bb4
zd43a3ab8f0e5a9075397c21438096f42d8c71c30843623cbd08efee32a7d2a3d29672cf277ac48
z4216f5f9833d968d9bf56b1b57b2e933ba167e3b724829376055f6d56f94fc790c82057a8b79b4
z208763290d0c2a99633d3e1350055864b0cf089af071d30010ce7202a1ac32c9e9a9c32a33d312
zc3027db38890d79ff39dbb6871e1641f0aa98d9c077d6245d7b09aa0b1c5ed868dbc4737c8c9be
zdee95f6beae033a0b48e2e43baa7272764143f066bb443b84a0f35cb82de9b779d2ea8038da8b4
zf731d829a3ee88b1ddb4641ec6918399d680de87747140a9bfeff66ffc0f16614758810055073b
za45ef07399fb47fd6a2fe1ed42a1ffb765cd1de282f6273f945d529e0c94fdd8ce6d42aff639f6
zb0e4f45c04c7d7c108984f7cbc4768145e7c8cd583822101ebe020a748a6ebeb193239c3fe23ae
ze9bb929983c926453f855823ef7edd5f3651e1f30545f7d60df1da7bd1f83d3a4f39305c0cc9cb
z2be37db5420ccf7a157f22c0e9a725f00c940919e90a01bb6345d7ea5b3585da0fcba8aa72a4dd
z6ae433f6d910d8de5973c83a5955f72adb150c2c4c71fc104f4e873a756acd7dbc7b042b1755bb
z84035b2b06a6676ae91cefee2d036a5395b6691fd7305aaf12e2baa17f1f295e3d921e4c3b3d42
z98a790a31ef7a11e85a48e550c54d6ffcf2e77be80e2689b4d972326a43d2416bac91760c9876d
zb40b5ec0beff7b3e6b0ab429c41ebca8265e57f23f560d80d01d64b52530de0416478aebd34826
z6b852212d0f8cf1ce28091eade85691a370dcb9009a5d1dbb00d560aac6738e476fdb6bc149e09
z59d67a9b2b74471220656ee6e83e1cd37075dce1b49aeef13a3158b89042aeb355acb19d4623a2
z3e0a42a111ee9f8b0c325c521b28f0f033a99ce0f0422bda0f1cc4ef054fe20d215c5106087aac
zed0ac65513e01255ae3c711165242048201d7467b9acdeff411d45c6d25a3d4369c4a33aae9f21
z77bb610636a126c758f065d324129b7593fd44f77a4b0d1016e48afc8c639d0be7abca2ebac9bc
z3147566b549654a3116de7878fa1411e01e070d41108ce239a9b45f5c54be468bda26db0cb6bed
z310c44320581adf89bb2a3e0a7d2defa7e818074881864a98d908efc074bc3c13e7556908c41da
z86f3834b1655a0a20e0e8fc1996cf1861cae286a209b80b10dbd9f8b7a078a1c159c6823c19b28
z5e4dcc85cbadf8fef75f04abc605fa7bc42aa88e4a94163afabe7832542f58d852dcf3775c176c
z3f524914ea15c0fa0f621db517cb6440762166211e35f2696ff98fcbb9bd2fb4dc6f4c0849753f
zae7aba4e833db6a4928403362a19fdbffa1023c4bca9fd908d923b2a4751b3f55a69bd4447c904
zb0709c08482c8ab2a587309b1836dd35c0522a0d9f69517d5cc61dc500e411d7e50afa27e49fb0
zded2332f707ac938bd365aeac28df62bbb7bf3eeb5732de988eede9a961b7cbea1cac480ef13d0
ze7b596167b640a26d3d95223f2593143f51b69cc9c85a3d970848cc4520f5c58d2f7d1ae7aac8d
z70a239a59a7302c407435aefdd6164693d829e2c57e16f0e060ee172d80cf827eacde5e04aaeac
z1ea79084a3dfe486e68c4dd3190b101704623d117e8c0cc4d67e6a6f2fa91cebfe098589bf58f7
z225aa3957689fd19699c15e6c7aec6a12e1cc26a8c3d39e1c98b0a43488637314a4f95455b8735
zc65e3fe1ada9b251d41720adbe1f8663c3f9c7dfd1eb79361701fb55a2c6dae1dc0caf41d7fb9f
z604901dcc829fe7963a974fde453c6c1d9e7b1fa93b2d6b48a62ef1fdaa8661adb80b89fd5d90e
z8676788d3b0fd27db9663279617980dd52a94c673c3d54fc2bb25f0057538712cdcf047048f1cf
zff999bf4a4c167f1f4798911b4aeccdec765c1a76e9e01187fa6e1a3d7cec92662b4bcf7709c67
z0a43da523e367766dbae02555dd367aa3970a0a5dffd7b9eb61f78b7e478f5fa15330ad4aee7d8
z1aed84a4f97807ded27d9312fb3b0ba0535e2cde6ce09b0101c4c0d2916538196122e76e7bc197
za1240c4db3a9d8d101e228af6d4965d71b80f074fcfcd58cb340998fb9899ac71997622a4ba995
z1f51c9774e3a5c86e52c528a3637b4a3e34bb9235e4d832740a2558edafd596fbb3125e9c9fce3
z4fd410c2d84e5fa8ebaefef818308d064f7178f6f86081d94208eadd15a78046d67df2723a834a
z498cab311911f7e41c57234963a127d6f063324bfe2f46b9d194215b2d3167838fb1d34e6df68a
zbebf6348e512e2e4b413051ac5f8523f9fb46843677c48c8a39c352418fcd9518c7da3c0b7411a
z3b5768b23363cba7c51dc3e574d90e20edb1c9431904e3253836beec22c003dcd0bda2aae6af81
zce53643c5893fb797922a789767c7da02456989d82b8803b0e0e50c2275ff7e04b4f53a042c788
zb4a31c033fb97a58254b508b575c1afede5ec80cfe05fd1de1d4725797784b7260b45e7862313d
z923cf0cf8e3fb715143301f5f5420362ed96fdf9badfb9771ea34a867ebe052fce3bff4b4dab68
z2d690f94c25208d064f8efaf252a3a5db7171ef58092f3aa9995a6315c13d715c9b8839010c294
z454fd41abddcd56148c264f64149be87be335ea8bb4687fd83849adc1589440b2def0ad7985f48
z5b4e3dc113c263940fb740562cfd5cdd3ba60e26145a4bfbcb765f16f3869927f53a9779c1a4e3
z7a9aa1bd74f99058728a5e989f47f173343f73489bc93da5c64aa2f80276062424bdc95c43a176
zb479b070e273daa2c7724a9732b63488ca7eed3a843657aa2f79a84977ce4570a4817ae8dd5140
z4f4b19cd49c7416d9e07f2e81fdebee0fb4d72a66b048580e580bbd5da4558f4a41bda331243fe
z036ff0f2e1920f9234bcf76198f5cbc7ebedb96f63b7f6b34661aca1c0327756567d0225175531
za712ecc7d73ef6baba244c8bf8a695d92d9847b7daa595ecb584488a9aa595d786d277d879c71e
z4c7e3c030e503b3089ac8ea7002bed714ded1ec5c698252a321038af3c5fcf57a6aa3c1291b712
z33dbf2039d15f66aaff5b1c17d6c9911859f981820fc17640c4e66f63be98c39085c8fd067cdbd
z90375642a153c559ff10763851bdb77db3ccc05f07aaf38dc9439af170100d9a879e96ce8313cd
z4979a2bfd45c36a26cc6e0c4c7564eed3526a1a87d11ae4ba549b467b3db10f5982f586247d2a2
z50aaaedc45e2ad282fdc2a4e22a2ae08334c649b8c02d4c8bda9235d19ffc8170147c76d40b308
z94e80efc2427df758b88572bd81267d83460167b35acd218cc31ae12ca4e25e68c2042e5e27f9e
z4d3de5ed333c04cbcac15fe70159bd2f3f4cfa7b002b52a031c3bb1307462bfcacfb9a67e120c4
z95bb143a6600b6ab68b89f7ccfa78bc5cbc276e981bf385f6fbf57d168a43d72ab8aedf734a054
z0d08d2f86a3c39f4841d5f7b966a44aec1b459332e11c8ef3e12132bccf5eafe2956c1f7dae59a
zd7b6e0c5f089af6ecc61cd4755112618acf73595471a1204e68aa1fbe2c8713bbd24796aa7d8b2
z2aac980aa407e1eb29b3489db71deab6c4b225248f593119d730572c64dfdb3beff52acb236818
zc3a44f63ebc277318869ba42e2652162712eb2c895e8f8e3416c930116dbf6694a7d54b2a488f4
zae9c89c8417172618080394334a2a24576292bee990139855cf88403407f7b741e0323e1296f92
ze54de1c14fe57aa99d57201ad07b4fb16b072b004e203478247d154376add6b2e21af2d349d41b
z01f6b31e86732a25768856e150512cc18609557474bfcd0f672d1fd361e2ec9763de26ee4e3230
z5ad892e736a78ee75b13cc233413c38424b7bca9da4efde49c9c48ce1ee9540dc9031852c275f9
z72b2e4d6b746f51a514f9c521b853c7b5ff59f8d2e4e457ed1d2a3611e1213fad138b95c278d02
z3fbd9512e384ea5b06f36093a920b7a7591a2d82cbb5b97237946c411ce42d661fe8087bf74f7b
z80821adaed964502cf4c074b3a0ced475c2ad15d88b6281a7878bfbdc4ba5a83847e0f5520234f
ze95d5443f5353bd36c4c891c3fa8f48a51241246309b7a0bc3c53b246fb2ad360a32fe2f08f226
z21d3cc25b2966dce775b013c29f9fcb3d86719dadd1758445256f7619ad68a76ad31d16943f095
z075e431a0b1da344bd82a80b9fa2d0cfb47b661598f111a1449aeb9ef87c504b54b2fb0cc7e9eb
zd678978cd644fe0ebb2116582c4579540101b4f1b1993d71bf617ed59aecea2ac5daa461f1fd75
z905f81271ef6657721dd007d2efa50d359ccd6d0da5ef831ff8bbfb48af501a7b7dc7d831a982c
z55b342e62aad3f94ffacc26dfa35bc353e837c84c8d9a53a67dde91410b3be7081b1c97d439ae6
zabf45f287a4234f273fc21e26240fbc3a58cbc2e7abe3d009c62e23e635cc7c66965efc7ef0c52
z315052dfc363b2472a7e15d276d609a4239d29719266aeeb56d35ac27dcc5c0688e79b2d368b81
z1e61a7486c053aeb7a4b5ce29f7ff8ecd94b37457337039356961ff2a9d18073addd933b16ebab
za73afbb1a15fd3d849ca86d8e164c49d540a330924b340cd4ca2a26ac9454cecad004ffbf293d0
za521db6c8f312fa0957b394afc248c1f9dcc806768ed4720412df928c88fac310af2b39fd05a06
z13514942a6d853686f84f8da0f1937bd099ff9f59ab26e1df4ea09c0eb428d1348377610c06472
z2835c069daae9d43657b3edda34d3fc47df34a72b1e83bab74eac23fbd5e453b93409d05f596e2
z94aabef3e2713b6971152db0ee46915212cf3faad29ff8df828fae4966ec2f2b8612562946e412
zf021af99b27f2fdb3d290dd84efd075acd7639cf79ac7b3e6f3a56f4260fb9f6a10909a9902930
zc59336ee114c2229f52463f2bb9cc5990828594b718849b37835d34a7b1de25b90f2d2577433ca
z69f3f817af545d1fdb4d9fbf498b9b493c760e1f1193627ddc511c67446e6c0ddafc8c3ee2bf6a
zf38bb075bccb34fe4b00982d00bdb20fd470df5a42f4c2186f778659eed5e2a5af27f6e52650d4
z9aca180a19796a33a001fc7307bf3a664939191438b38578c8d334924a2607b3248a27cbf29bf5
z19ef046d1b9c872071b6faf84806a541b7b780f199779b7964f3b41f956e470ee952307115af7e
z8df574924d72c6f21903205d98bdcdc148d66f5ad307d7ada30dbd903e4d403baa0cb6f554a058
ze006280f7ecff7ee3ad44cbabf68785eae4cf3d4f540cce7450772a4f73a2ec5e362c6fa56f675
z49100eef751a413c7bb2fa44e1b7edc567679b1506bd44bc371f8cb1228fb2d70487d88380ec23
z9574d97caf0b08e140fc4a9a981206a2db137c64e9ce47c0667056921c0f05c4325689ded3bc91
zd3d43e76dde0e4b4a0901fc0008f559163cacc7a60f82cdfcb809bbbff8d9a4c300b0c7130dbc5
z7b4e586af80b8c0e1fefe059d7ae8f094a87656f4eef8b39fbab99f6c79f9202d4ecd50430b409
zb4d898eac99c3dc5198977fa9bb2431eec56589a77e5acb2e50af388e17434e6ca063499e372ab
zdaeae19adf36fcd8bcc67c36a02a2c2bd952b5d0a3437f9e3b152e04c34361ade1d29a11e28c79
z0fc7663f15ec40c7af9a82b93c70b4b8964fa9153b4b24746a174ccd8f75134f192773971dcde4
z2a2c0ea4542deb8d9f05471b2c37b477a82bc634237f8de5e1a9c34ff00a298cdbded7a9631d86
z2898a589cfa4943a33a5161ff532878beb5ba22ca71e04cba87ce5e7529f61d68ef1bde3de0cf8
zc5e584090057b47c14667c34ff2fc4d4ceeb1cfd3399d232daa9b169eb8564e0f359516327823b
zebdfe6c319ceb45f04cbfabc62cd1c717a8e3024e1210aa457c22b6499be0044000dde5832b880
zad5d90b0519be2b215cae35d33893a2e68a973eb0b70e6c076335133361575533b89ee7718f72a
z1cf1ae38fc24c6f052b2dc3408bce1ea874e9637989e04725f42be5936663b17cf9d8aa025c5c8
z5eec8abb17f9fc358d1c96d9b0d02ddf2ead1815768d991016c2f3fb9ea0d9ed4d897c95380313
zbadbefc71f7d5d712e2b5f7402b803da8d0c37e4c7f514525262627c78830ebdaaf92ecc9ea307
z04ec36a2a624e3f356f66a12204983c54cf33e306d191d4fd0a16b09780b7a78875fa5cfc0cc8c
zea0133087b4cb1092efe1a222aad48fa1505d9b9f2a53272d499b8679f2a2f0adbe1eacac55b52
z082d5ad954f849609710e38e7f4d042cbf6c620c005a9219adfd1d1c8df3ecede49a4c29a4a331
z104268b054ac6316a51fa78d6c622720f0a9bbd2c4340a1bcaf3ea152784ce992bed2599e601ee
zf3525389c508ee0bc4083221f2c9e4677f81331c17573ee887928609c192bd23006b110e7e9f0b
z41c2320bab9f8649bbd7011b53a3137ee083521c78b642fa8b3c387402b887c7e088b97d2bb60f
z18ee489e4e9046bebfe971684e48480a128e1240b4c098100a46e10b151362a474f7b99058bdee
z705e3cf6b02f32ef2ae126010a5b36a4df95d2853ae08bca4a0064ce8cc48510ca7072302a9418
z3b74a73d630e98f1eff054ae9e2e702f945129f3cec677f5cee14e4b9f7adab9bfd2c489d769a4
zf0a3f7d6f2fb3d9636057574cc73e088a1c9eeea71a71044b73589efe8db5beb19988caba0daa5
z41eed4db72d2d64aa7cb9555acb95775c8234373af3ec87778de5bc314964c8aa65cac7ea18451
zab415882a59e519cff0bfb12c9b9cebb62041761ea7449a95e839eb2c08aeb3d699a23d7769bb5
zaecc19b41b2672364b8b3064453340816b687cb72fa00a4e50c3e22a8cef8e550983ff114c688c
zd34143a0b725a28449fcdb3421315bff5043ca1d026122f45be24c0d863191308fb73c25bdbc34
ze781fd9611d16107ee0ae8a06dcac322accadeee7aeab22abd3e5d8bb5e2e96b47cd785e06e381
z33ed3de57c71f64fdb597cacf4991b40fac133f1a34104b1c1b63b0b17664db0b5b343bbeb2865
z39b7f10be08cba5daad98d5c24e71e6fec6b52684407a9e588e154705958c89606920029f44623
z15ae213d35c6d747dd549d0349729fd429d3d9a74cd57231e1523fc6568ff140fdf26379272f97
z9c8579c84ef3b02e4d8000f2181032941dc3ab6718335e41641e98fd31acb6aa2856d0004e6927
ze5e4f42a47ff8bb340f8ff8dfa459a4de170f5fa55523e0b784161eeb685df797f93c63d837ed8
z8e3256e4692592c15a40f9fd197dc6de50f3227ae9ebd9c02536d92b3e301c28a40da596b40f2b
z0bd8c53aec8e25bc710cb5a1d21d8e0aa31b35db3ab17358ad6f7bad51ae58121de2ea8d63eb8f
zef4c8bffcab91238a59474ba4532291809c80a3c29c709ab92804009ffdd14c7674508bce53518
z969ddeac212df3a849a0f32776c9887978007a3cb674829d64abbf2f495cefbaf14404e815c96f
z26d1069247052c09605a364a672638576c438597bd6e88d349b49efe63977555595a90b0daf22f
z421b0e03a7e70813ee12b7c4df3fbf15f3333bebb616ef3733cf4ef67fd00f974a5288d1c1d89d
z8f5760f779d20721b547f04c695cd2484bce9f09156992f12fb16e69e6d69ab3c036ce667e2da2
ze44fd00fbac6c6e9c9a0b06f1a0c774695659c56b147c899302540ab955998d6a873e932419491
z7da8d9d61e3587c44276369b136b88d02c20d0a0133a11543bd553553055466eec4ce229dbfb32
z2579e7302e67dbd7c054396653679e15ea088a1eed5e56120821da762806a0613d55bcac7d1469
z52f5c13b7886fae90a446fcee61303edb5ce7c765c2caad49cad6be120a34ef67aac9f2574b1af
z2c87a2e972da4fb20ba4ff64528eaffd153639f3a866bbbe9e55ea29d4140d2192ef4e5cd5c11f
z2e740135f3c32681f7eab2c87fb8fe2e8de238bce4ee7b000264a691de16d06237629d2310c77f
zc55040a8ace7895e3eb2e267b44cfa8179b1b6edde9ad22e10b570b67d60053b229df953c2c013
z58387bc1a3736925cbea365389faf871af1b30a43882f2cefcb4296b31a7ebb991d646707c79b1
z855fa27a7991af9d89c263c864e3432ba7bed25548e671123f673ee5661b7d914cac120ff9909f
z99c73c5b7c33596920721ca3a7e16752f6d6c2da246c7cee0711811d9df7e630e07218c1b0129d
z56c5d74eeae514c034dc6fb817d94bea11f7905f51df095ba703ec8fd627a9dd48cefd0ede3cca
z5f4c601876a9e16cace3838456f06085df38d35d6b003f1c3ec47c79767e5d788182cd1da7e490
zd4bcf8e04883e438569302cee0eda982cbcaaae61091050114583996f51d5f3738a0eb459562cc
z5c88a6872c33c6a406bfdb208d9127d84d53b90ec6c36fa11bc4a3e494743429560317aa423c2f
z5db204c64b479a641d93e0b3fdc7a27ecf834722114a2b5779aaf7e05a282651b2513a8df48828
z523d9a62e7c379be763a00c9913d9aa8ab6f818b70a841bbfbe9d085b09a69ca43757a6b2a259f
zb3defdba47b3e05ed03f1ea7dec0c5239e999be8473bee55543f7e38bb053722a73451a4a1d913
z6d47c1204620bff812ac89de97d64e7af214a393806d3f83e9c1bffebf499459ad6ad3c28e58d2
zd234b8c82b85581dcab3f451715f5067b9ccb16c0c7921962eece084f6cae7acb0da611bd88091
z13af4a735fc025cd10cc628c5e5a7a40e2ebe1758d6b29e380bee57a5cd446340b2e50684fd7af
zab49bbed59859d9d5bba18f3a723dabac3fb88c4522211ebd0dcf2b246177bf0beb15159fabf13
z63d8d0f2e6732f7926ccd3d1cf7260754c23dc3cfe5acda3d61c8a6f97c3e1bb9a178e3e1f5d6d
z488c22428a0671adb085c72dc97c0d19c90cab792454e7c50db9f83e8396da82ab305420b20b47
zf3f4245a27c8ab4019afdc12972e66dd0c281c8613b7b8915bcc320610bdeead99a05d56508c88
z650195c57e6facb9bd91ffc34ee5981ad22493b49a7f25c9f0df50739d8f1b1a739b5796c75b4a
z56c4882122cd1ab330b22adf2d047143edaffd2e08ed459a4800a017847245887c0003f57e3daf
z349d9c1fe6c8b88148139a738cf8c20d59980b3f32a61c5afac112fc76ebda3f7cb2726edcc6d0
zcd625dc20faaa9c5bb363b8fac433333c872bb55c41318b191f3fa0268d7ef3fac4cafe82658b4
z95a11e50fb056fbebd1e3e7669a3d9d4ee6e4ce6fc5ce07395ab6cc0deec43c81dbe55440a285d
z9099604d33aa9967cdb805125b6148b8658b135ff720d50aa819d3c72dd1f994b214e10f24b1b2
ze9fce216144ccc2741282b7ce5ccd8c7236bb17db4c00e2294519d2731eb70f3a5f472bd366706
z3cd19dbe207570ece7b9fb7cdc31460eea50e8511516dab5507efce29f136487e15802b3ac1c92
zd417c17d5314e07f642912f6e0bdfe1d4c76f8e3bd06b3a101ef0b2b7825c4c8acdac9c7b58f32
z9a724bc765d05f9f66c87ed5a40eeae726de58b90a2cfdb9a926a6f852fc3ba558e2ae6e67fec9
z1437ea056cb2850bf6ab6dfe3b09b1fdf93b447f5ad7dfaa1a1837e5071a80b926ecaa1d452f6a
zd5b3878138fb3e77aa6a0dded4dc3e68348b8290cba5f6b4908b5c0e51b2b36557bf431ca3c495
z8f4de5778c7c771eba93245c935c91e517d3047f06a51b6b31162a50955378a09cfc96258f0966
z569650890005e40d97b35da48dff66eb22eef5b016a739c4cc7e1c772659929bb73f1d46f459c8
z7b020e347ff9f98675dde187d564461ebab0a5b890e044a62b29a8e934a1e99fb86f70b2302ffd
zeb4c42157af7e97c414f3dac4470a564e272ab53ba7a7ff78557aebf8e6edd66663ff5e27b2f9a
zb795a4ff8f5455f1983a167364b6a2a2f37715c4d9757a451f4f2c40da942240cfa9a75e3a4862
ze478c8553a77723b94a3ff1f1300c02fe8da7d63408df7d9c4ac7311b7bff78c7e06e0a6bb1c34
z6230e8b572ddd0a86dbbfa2170d4fa6d001b254c22112cf44a4eaca9b0188808418e582bac76c6
z16c7209a52a340fbad5c0352b101d0aed1e8701e29397c761a834f49d801f7bb2d19baee76b11c
zda0915e37fe7f3c79982e4a8c095a533b6e212383628ead626c8a68ab33ad059dce6905ad2ab17
z3b936a589166aeafe618dd7eca36f18eaa3d170d6620637b22e38d97b010a2e2da0e6593f025b0
z642d6a73dae0adf245266dc31d3064614035df99ecc117b16db5efefe7f7fac49231e972d1c1a5
zb2ec6fdd280e8344ed508932e00a3a1e95d96870adf902c4f218631aba7860313e7012982504c7
za6378353c3eb5fd72f96648b2e98f1f1bb00ae6924af19bef7a54c6626e04ad762b9c1b69e7af0
z648c6e6c6a78afb9eb9ed32bf3f7594e07c0a39433f0a29561195bcf125ca41d17a6da9b9a407e
z2c4675d9db2a3d8ec82851531afe198e4259280bf7d1e0410ddeab53de7fb0d9ce1a0f34259f08
z7117b5c8273a330c77cc7efc426c324622db50f61ce20a2241f5c93e3d340d111cd173e18c5041
z7f63b7d42408b6dc414e5bc4c6f76d240e68414a7052e5b32d28fb9fdc1fb395436f9a15fa13cc
z2f2845f7be737f1c6687eb4ef4777f28b0162e0ca0afdab8bbe0fcb716f27952f068c7f369ceac
z086bbe9fd9e451a13aa1576cc5f0c5310714afc78042fc43b06b82b17e6581c1889dc23941b7cb
z13187b75338b44bf546b714fea57d79a1231438a7416753bceb55ce0daece3c0157981ee9e0d66
z0babe0fa99ffe1575da28c934347ee91ce8444844a6cd180d81c107900b45d9d09f0e9e7425586
zdd38aafa7affe88279b527a6e49af3a00a2df77bddb758fd8324f9829f89df64ddcafb06c6ef3e
zd41b0605f9315f40384bf0b6d375cfb4d443b54a9b3ad6a45963ddb1088583e6d4f00aaef8aa97
ze2d2306dd48e6d9de5171c918e7d413ec814400218972e58522bfd8b748567c1aeef47a554a8f5
z1c9f810a7ea76772c9b74682db810d513280319bbfc2324a28b45900987f7a23c9ac1517317b0c
za05c5d8153f65b3d8e36622394be5462cfefda49731892cd280d2de4979502b5c6cf05413109cc
z91b99930f06c2e02c5a1fe0b860df83e10fddb40cd89b916ab9b81675e9be7cddbbab1fb257b5b
zccccb7657f9cad2bc4072c3cb628297581070d47a5abfaa465477e2df19e22045ba448a92809bd
z279530b36c709500ca58107b3e5b1da4ce08a4c9b9117681a0cd15b432faf35f91bca493c0cbde
zb76f9be7b047580b212c75ce3b8bf60ba628636972df4622b36fcf6a2daf7457c3991e2c5f2ca3
zab3953c777b25db3d6cfdb70456f170fa63382414068f32e25cd3354bb9191a6189840bd200d6f
z6e1630f7918992429aa951a7f0ec9ebcce3eb40ad33af46c19291adc7866c2608b84697a927b12
zedccfed12bfedf45af946764b8a7e74ddc7eabf4ff6ccba406d778d422bfed9e82695f660eb529
zda954fad25c45504824c9a8b6c18d6edeb407dd207e2931ef45bcbcc958c1056026dd850f065a3
zf6e5b9c8f93075752034ea85d72d8ec9aa44b78aff02c5d0c232759c799c080565a7c5d0d2f1c3
z976fe9f86fa2cf17624f0beb36eb3a03e888f463006369c4fe646e1c4a74bfc1bedbd8ba70e7be
zd93387fd82c1d445591eaeb38eabe4fc478fec14cd0b525e9468b2dc2b262a68854bcb959d5ef4
zccfd39ab96146eb6a84bdc27c958c85fdce35ac5f16ac5bbab5e3698c701fa9822c93a327f5aa4
z1ea92bed270e88bb22c9b58d5fff027f4a764de4851745ddd3e6bf81c65d99cd3afed6a33ddfae
z045bc218c6dc3170db9a847969a299aee1c1551d6c928857d7308a60302258a62357fdccd35b83
z32f184720126375531edde5873eb244ae95264ef83eae044b034c09df88412cf95c425c0181c80
zdf525fc6e4ee5157d3f1bb53b07f8f1f22483d0ad66309de035b44e5fcfb7506cf3893e0cd37a8
z1f28b2f529b378c44206445a5379168124e473392cf03dbd8bf8e81011a2fa7a30c80b9431c287
z112dc9d58e5282e65bfe0b6b28a91076a3a265a82a9c80c221afda00a39026f5dfc2b96d3787e8
zbce5b00a6fafefeed07c3ef86805e65560cd001a908fcd4e1a77551a179cab8c1d783d25b45af6
z0522a288ea5bf3dea810debec467f27947ef6d367331152f583df71497ebd8ed4bcf1b68e55fc5
ze0236e64c4239a1605a851cd2ee2500742b3cf6799a4f7571273446e14899b6951a216fe195407
z27c94c51c97ae1b3c796aed17d305ff36681a417de077b58d109ef617316e6c8f29216b59e8681
z53548a0f667ca62baff2ddce9c33811809495bc6c6fc707c8edf9ce21b3f028ab66ec16188862c
z8ff34fb2cb92ded0c28cf4b44821b567cfd2b584d7d2f851e58084ab5ebe24f544a37d94cd78ab
z92d347d1d29c70325123ef136ba207daf7f04aa78b7f3081d8a7d0cb1db767118c43053a25975b
z4d41e6649a30c1314de094fbde1c1c40be124330c26f63819b38e3c6255b5f6c9882cce4e73304
zc8d7825965a526785f68237c2f43e00283c004b9eefc4fc2315d0812b54c2a8782372b0344c16f
z8a8c00aae18c714b06260cd0103bc1e397b555af3720b1501539407432034eed6a73ddd0258c77
ze85174e689299043443a9a57a85df641741b08d099d7f6c55c9446d436067557a7078fc2efc931
z946e2603d34b2f160dd250d74c2f1a443aa4eb9449b85c7a5fe9e7987de18b547245d2899edcb9
z0df7e0ee16a9a268c33fe92e20dc908e8b220a5fe10f7ad6f77ee8cc657cb7ff6248e936ff6cbf
z1a9e61bdafebde7bb040a7252facf55e64fb2855ecaa5bf9fe7d5ced468b1c6be8a559be95d0a0
z788574b153bd22bdd2c4d83f1c7c0cdb056e9ac851c6c159452166ad1deb58507f8a04ecee4f85
z690af7daa8a61f0b9e50a26a65fea632addeca971a9aae38fca9d50ac8786a001dfcefb436e4d7
z569e747fff95db71956e4d9424e023196fa36b636844be864b9ff717b1c4e0323fb3eddd088e7c
zaffd275eb1e6dd2f6776371d4d785f9c54cfb60e323dbf28738f5b684bc9276c6c82b1fbbb6a07
z54610e906067dc8247b323c9d5f5616e3deb767ddedf7b1fb2cc346590cbe36a4fe93bea05006d
z3418f6022c604aa2377281cdd5f88c69efbe8b9924e73b313c8b890ff05b980f897654b269d767
za76bc982fc43b16f7df700d18b90c1c238f608ad5181694aa48c7a402efeedc79a275138d23ab4
z577b6a5d35e16ca7dce796bc5984a56978210c12dab73f2b4eed805df14b4f91a486cb0749e770
z62210232a884c5b47a126c723f8d4c917778baf0a7d600d1e3544ad6f3ad3a976207728eae4ac2
z1509f3e2f68f81c9a9bcb5557938770b2775ff69a24d43bfd61807670f48d312e7373490bd3311
zcb37f4ef7908580f078d49aea595e4f825b1c229688e4f59aebece8bfe8ac20843065a2b346764
z158113705648651dbfe65515b1ae4e506ff134fe430c5ed798a0fe7b748e60bc9b9a423d7a633f
zffafaf248073031e0442366f53d1f1a8bdd26ef907c82d3abb1e72c2d8804be939d630e6b9c73f
z802751d5d31e303d9977eb60f7ce342059e8322f9d2a2858d60a03094ae47d40d2f64296e040ed
zbf8f13fbcf4ab9f6f0ca1c3fb161c33c5e7fd8c107e6305d61be5822693c17d422517eb4023c20
zd0b6857544a44fc91b319ed6cb3e2ca8895323c3cbdb62f0796d03b7b11385ac0434d7a24c064b
za7a95b5b0a42208de6f8b048cdc210b63fae07097beab8c323ef2e2844c479056e0560d718a2dd
z0525bf8de2fc5ee4fee39196f5f15f3fe012a2811127327beb03b3f482bb6dd383fdc1ab8a21b1
zc6250270ba9acf5066214ed96449af6b5f9d88607393e955bb4197130e6e2739f3e036ca86b16a
z4dd8a70f44db86d64b2ab060a208ebcaf846ddfc3c5d7d09e2f001db99970612039ad457062faa
z88439705e6a382cdba743a022362851687397c41449872564604990d417dd36dced940c9872669
z31d583818e6643abc51d95fcca6d5f66e16ba494e0878303ce3a81789febd1bdeab565abf4b3b9
z882423b1f334c436888c45891fc6404859c1220d8b4714b05106bf8bea1ab51a0fb49c81b0b2c4
z8515aad4fb7f04ccd165242f5d002d68c10deec68f11da76a9c2345fb9eef9349bb9414633f539
ze61db8687d2db8ab05aea81293119a228b263ce49edc3fc158ca4698b9cd5ba94a51f9657c18c8
z26241f80c275072bbc172c646c70d4549e2d8c5b5f5cb336a49e3f882670090350ffa1d91ea6bf
z382a8ed410d1970c49dfc69a88a28dfe44771aca80fcb19b15cfbf35b525b392244be0c1127003
z7be755833a184ae6b0668d4807fb479fd1acdc46bb425ca1d4c8f5a2bb2398678507f3786df42d
z5f82c5c3aedbdbe109bb2fe12605ebf4123f105cd6f8be140100dbbf76c8fa7fc9f8db462db1aa
z15d22a13bd24eb84e479dfca3b067c2f3a46064ca7e1fad7923bfc55e4465ed4e1377d8e8e90a5
z619dc9e4597760f6b668bf8f39144b96a8c15c0add82bbe9b76ada371e4e2caad0920d2cf7dc04
z0289db8afb0bfb45486644a8e1508d89a0c96606b98b19506a80d87f063b60d26de15355e4d399
z1ce6dac9f72fa28b8cc736ccb11c51657f5433d9cac7760d56f333a45aff80ae65b95a3c93e51e
z290f44802365aeceb0237a23378877f0450c882688224fe7f8f8bc1cd99855debae52aaf8607f0
zab2f3e388df797b2588539110442a20303e8402524a7e45d4d8a0ea48f492d27216d2535af8207
z140dfc268cbdbb853d5124cc95ae78831060e5ab8a638915231b213fba0dc07e5fc08c92cc89bb
z1e46d22b0945e29f4603645d6849058cfc44a38405861bc4b97689ecbd50f82c9f1391f5787ca5
z099643f19c1ccb674c8f3d18f623bc64239ff66f10f7ee34c243aa87a88486418bc2fd12b304c6
zded1ff0414a28203fa112d241ab18a45a24e725edcb31b3e1071f2011c7e53054d2f8794ac61f3
zd7eaf1f6863c1089ad207123d110d0b9be85bf639f6b7afbf1c38e8310ec481463333438ee09c6
zff1e593d01e9fa3db79d6a66dc4fc0a7eb6af614b3afbe948dd9a221260b793497975933d2f2fe
z5a3f704cc56f43fdd116ee3e1d915bcc93cab2f17cded9caced8032e532c8d38523610f607dd99
zfd356946602abc079358fdfc33ccfd69589179f556a1e38417d7e89d4f7d7bbc6e096bd13d2a00
z2b7952fbe82a470ac420288b82532f35fa6fb3bf0952e67619e484f88d012c52c8eeb775567ef5
zec35cc6d326b413c377cab118ebeb3197e09ab2ce2f8f26ca4581193b883573b173fbb59732701
zcc22da374530814f6feee8d46fe162ed06faa508292a9876250a6da90c3b1ede0851624c4e042f
zc6e0fd87d182592418ba881136a6da3dfc7c410545f9c3b48cf5bd1f9fa6a2ea8827fb81b9343a
z0eab856eb52042e0c75e8352b2ae962200ea8ef6381f6553f5bb86923baf7903fbd269184542ce
zabef38c54b8be56b6081650d0871d647b01ae4b0c667d693c65e5da886f944a8c5632ad325c811
z67ed88761efc811e0c26e22268b8be89f3d13aa1c3f71644fff44967d758ddf22ad8de4fe8c0c4
z7be3411cee05aedf1ff64d75dd58f6e95d62dbc7b8bcb2944672f506ba4d780d01cb6666b5b47b
z6d4bee505179d01ae5ac26a4fddd8ff2c5305f2d6d51af8dba2c92a787058bab399d75d6aba35a
ze294148e37219d137c2ce20fd6f2bb01e377fb250a3ec167a3d9d904572f4a38101fe0eebf5f11
ze1a20ed91364c2c80d2316d929e16721b5ca0b4295d3ebd8092a57e69bf3fc260094ec040f54db
z9ef199afb1451124d5a3295f4a2a3585751c861e5173fac042fba869320edb8fff2cb3d6ecd814
z8274ac82316e7ce51e5e88cdbab7369126c2a7f22a577d20984165aeac97665d4d6e1b7d8bbb73
z0100b7e8ba583074625dfcb6dd28bb61e50ac6f1d1fb60f8e5f8e013a827f3c4bd03607a7e7941
z3b5009bbcebcd5c331e668880b91d2b3507a082cfe92af7d4c7226dce0d24d373a088408f7ac85
z43a4d4f50ba7bc5a1556dbd56c7cdc7901fd6afb6105313900a67652ac08ca665a03f9701881d2
z884a035cf2db4f599b6601b6a2ec4d7186d7343bd897905967ef77428b3cd0e082f422a0127684
zc5c0ffde998279b2aa2ec6c6fee1e01ffc317414f7d88793b3a0f3eeec59f17648b7a142e5d6b4
z8f5c291343e43396114b20c9d9ecd4ac222e726f1fa5dcc57072a8a2e2dff1e66180c5a2e0e9fb
z407091a008366278909c24ef4c8f60e8d0d6e8cb174fbdd4bcb4ed9b3991471fbce662c414d8e4
zb443335a495b34ead9ab3fa88c335a4d77a5b4d892bdcf2bc054ee992606fbdba706bdd599fbb7
zdeef32ad70440ef42ce8720b9e8e7ec8ceb8343825ff44b4390056d93e28f0e8e05450a06cb865
za21b1515f4fa657281d10408582dfdfbd34ed6e70db8f300175a0d6e95d842bc2fd08848365f90
zf4819812f91e0d7f5326cad20a0a80335f727ab6774c4f60174a913de3c80a1b012e3379200252
zaa5872b9d627e11767ba680b18ba2439a54abee67ebf9b21040a66ef39874085f88e0856e79b72
z596c3605d47a67c3801cba0bfe06975f1c62c729e1a08375d858cadbfc8f9731b110a2ee94dec1
z3ee21d7430b0910eaa4566ee60445cc2bd5d2afd8472ee3af008f5f09395fc7cd5c9c2b1d01e20
zeddfbabe55439fe0334ac43fdea843cb65e4154af5c7634251b99e6944847988493222c3f35205
zf3cc75ca921fcf9a8ecaef841e212ce43fe2f6faf24e13765cb12559f1e4851c4d835f61348311
zd23236d287cb219e3c2a1ccd82ae6294c70d083f05233602bc942f523ee2863b56a268c27f4098
z31ae592e897d42fb5d594d6646aacca675d0218b30f3e376e13dc974f554c81f99e60af8027443
z9c04f64214d8cd793d96487555454b974d616efe84cec985e96b9de335c99b3cf4e938e9f448a0
zde72c0cc0e0f72a9c132a901007af8e9d33a2bd9f1c6c671899e3b570efd5961e6a049d20af307
z1c3b3d184ce15bc5501ffe8f7875819f7910293746e2f0504b568c3734c456f51dc989a1693a3a
zd7eaf1cc3c075c5c4b81283dd262e28677a91e8532245d8e84faae75478b38b27a37c6035eef27
zf71976ce7da9fbcbde95c0d2ee9f2c6bd09e028c7578ba618bc6bfe552da6898a306a8de143f4e
z7d5f9d608de8a2bb0e686cd857fdbc764077a54286fa0496396179b046d096fda515d780325b9b
zc9de98e2edc5c41303d484d3d6bc8f8bc9e3e590aa48f3864f8cfbbbe3aa5748f87cab0511d308
zaaec25f2b9b8d0c011d633560820058bd7f6b2fd7821505dd93d2659b637594913e8b963d9f2e8
z54d9cb6fdfa3cb0a6686f7b1f1083ff00c775f5628224bc4f7f210bc56050125f1ba80afefd89d
zab7037ded2583eaacf6678410035cf2a03ba5f4a4b19eeef89777ac05852699dac48c024709899
zd157c23941add263e65ad5b34b4f1713d4f677a95c44afeb7506b86f14ace812c03bdbb7469125
z8cfd9244823124beed9e2025c1600ded6232be2b243a2d2082b217d794088a07971156706b67da
z0b82c171d46420fb5bd04960e80e6a58b71ccde9ce9ee2eaadbe4717915b1affb513b5e75d1cdc
z821ae7cc5815b2100ce8f7c6db12bc4d3c7fd6b35b2781cf51750ffe094f78baa6b680e4d2b026
ze2c742106a3462fcfd41362c280ab112fb2a7a04679c52d540656ea230b540093eff9bba4776e9
zdc66702859c7b2ea004cdd8f2d986dcd936d0ce16f053a9107fabc0b87d6c1ab1d694aed740097
z3f375a362e18c3798c5d937d6692993a22f3b4cbe047dae4d887bef9105ac9abd2617c5f9a916b
z0491c76bf3a05723f3c4db2723ea5b0b596c5cfc5778c0b0bb005c75edf933085752a9963ac2fe
z9f4c0fe7d4270b0b36c08a68303828cd3242baaee56d734caaa9bd1dadbf9bdca53564cc28bd9b
zaafce38f2241125fffed71e52c38e4b89ec00e3aeabcad89af7a215526dc059429e7aac2bcab66
z18cd14073bc77872b3eb4f5d416cb9cc684ffecf8cf128eed043dfa51af1a983524d4007e3b1bd
z6cf6f18302dfec3883b89b2afb834b781c282016c5eff6198f80b68b96007f15e352094f3370cf
z6d3abf3a5e13d5688613da830bbb86d29aef4aeaa5f7fa7840378eb5927b757f28adb94eab74d2
z0b877ee0463227ee152f914a0e3d61c9b9cfa06724fb0855733797043cf6969135d22c314ec343
zcabf9be6174fd78cda70f0a9e1cfc6d1c6a430ae0ec2d068474a160b957b10a0e91ac07d0d3c10
zac12f5144063a3f95a6c570bc5cb572bcf1672825ada5cdd42c3d677b529178fa2187cdda2e11c
z4b675294ef98a435c7f91287ac9b7139131a2c769b587f67a52645ab02048f9041769ebcccb965
z53125306e0265a81edbc8bd0cec8de59be32340fb015ff2e06802b2e6fbe303645b5b808549ec9
zd01f14b30e4436ec406aabef8f70298bd5c67d3992f108a59362a498ffe61f17315881582867db
z2d2e2169f4ba39eeee1da8399443f98e9fc3361ab44b3318200948fdbd0b73dadb9a95451d89b5
z343d4cd52622fe74d96aa3377b62e34ec3794d465655dbb0cc2474c4c71b315d33e622c311245b
zfbfecfdf48f38af999902c6786e0aa1604cafab2f42f35e0b06f132d9265a97fd33e59ef2e93c2
zf03882f56ce83eb043d89644bdf1f1bf9e6a296c8d5929a6e265f96b12715cc878cde9ff7e5483
zb54ae6b90ab0a0b98c480537195030f219ace6ea605c63f546bbb7186e610cbbbee063d8d84d9e
z6a415d1457ed5fc891116c1425e77ade998d4fd2e1dbc08a1bc61c7ffa2bf4d1b61ab9330b7720
zbf0a1b0ce7ce956a4ca3c31be9a3beed68190d6990eb9ac1116541b42e449d7a59280391c65df5
zb8d0e1b5cfc1a489e6bb5c8bc000eb4aeabab152c2e353ce71ec82773da9c077c674b0fabf829d
zdf5e1674f6291587b18e53e58b9aec379e1ee2075969e2c2c7be46bf09f8c7d30cc41b7a648a46
ze77eb4ee25a241bac7fc519c2cd1147727432825efbe9b3cd3345d678533d671a634e792b71ac3
zbe097ec6a1f3f6d7a3051f71f45b3a901990348fb10900a8e6378b8c5e02a51d94568585b125f9
z2dae7d0698303fcd9d2ca1d6b6e4d6819a71c9735bb969980e68facee995989d8f92652d142e1f
z476718441d490859fcfeb6810d345d88dc3f76205973deb6527ef1c780d7ac065a78cfe1812fb1
z12cd8897ab2d1b7159a87c3dff2c3fb3965d981af580458429e105f70700a0d486a1e2ec1c795d
zb240aedaa26ab52f53e9078e3821178c6ba3f6608a85ab89718195c5d6f81cfe06b4d7b5d44cd0
za75a7b5c46f13e5d7247d5dbbbcf8bcaaff66de3a2bf205e5b9b13336e65e4bcd47f1a78ba9242
z3dec95239327d8948796e1d69b0232497e5289d384ea51d55a1f0bf9c773c7ec6efc53978a0588
zb199778dc2fcf105ecb3cf2e524a476b00a61ba166ecf2f5066f7675a7580b015950488ee9a6eb
zc0c843e7732a1dc7465126042fe7341eda138ddd2d678568db2440493626dbe914cf06080ed7f4
z45ec0cc769bc28a7a58809d55e2e52a48631e3174467e44c280672bf9181390ac22a89e1c2ac39
zcbcc474f03e435760b990b2be02e297463e9b477d0bff1e04bca348dfcf11e97fe2787ddf71a36
ze8e8ba8d7cd3137db5376d4a3a75b8564dc9fd6a4bcf160dfa8048334411f7701d58bedcadc3e2
z29dce36ef468251052ef4d7d98b12631c1984f1e03e1513da9de99a711ea9835760e3148dae621
z4ebaea40bf5b24158547a08a8faf3a308bd3ac9ef159da09652d387911f924d5853f3462ca7ad6
z0c08ceca1a862a662c27affb645a783182ae2a343b88a99d5029bdffad4e2cf02cf336097a1b50
z014b032f223e09a1354e195944a8505941b83811c5f67a6e0d82c566e76bcc0b3b3eede7cc8050
z86e7ac1883c4b93f9c13d33adbcb52e04b76ecae4f2fefff015960da516a22f765dfbec207874e
za04d734a815b34e4fefbaa373a453840ba74a507a4b9ced08179403b314b5277a96f90610c0035
zdf6da54ede32a8e9f6c3f79f24d5f0de5ebad6b80a4ca1e1a22e167b92bd8fe4f09256410ec65a
z84335378c3e7e31c8f7c7d450ecda470cc1d848926232d3a26cd7d1670ede0a77288a00db74e8b
z536d3630215903a07d82b1bd733bdc81a0cdfa67a0524695153a7f18be3988880eb75db7a4aff9
zb32e77134c80cbbcc2d50422f16e2cabd980958dc04364e378c569eb97820c8281620c97962c60
z02fa70fc9f1358b6b84d85b882e5eb570312acdd2954adef0fab96fd617c6ce6e51db5ec74f2e6
zd6e20c18cbf35566139e4f2834ba63a57a1e7d0c2d9b436dce29489979cf9c6f08cda4afeb7db5
ze6aefcdf23d3f1d8b5d0028384134989d30237aee9b54699a1df11ad627083944a66e6ce34308e
z23e703cceb679a767abe2588399eb7a2e07b0b139c1a65071d2b4ff8f4141366eba06066fe821b
z7ec2c62b88bb0c95ac7a34bdd7838a161d61a716704785f08421ca4118b0aaa3f06f8847456216
z2a31332002b7a60a1f7395e64bd9d08a58004f781cb9f011bc4feef4df3a96168b4171fc923775
zea93e34836e276d3595f4148257503e4d014cf7b4995048731050700ec33add896d55918a4b34a
z5ae8985de85a4dabfe6dcdd254fd853e48afb9f70eb8ab2ebaf7b33abebe914cb5609430e2feba
zc58f86f2880ac3ce8475be9bc3bb127fcfbd7ef24054d312c02ee6be5e74c89e40847a0dd18b83
z5cedd82969ba3fd3f367ac2b24070a8790fbe7809d5eafb7cbca6321be519f3b7e8cd651739852
zddab84068e128fe1350d90f4286da7e006288b4273ab44d9373a147112ab4d3aec97d7e22d36b7
z497701daad21a78cffda0ae8b8490776836029b73c1e4d074308aa7e2b9fe9c75d71bccf2946fd
zcf8dfdca9646fd8335c821f85c83bec5d579a3f8c9315bb94f8e4f63425abd380dc0b5cb8f0a5d
zabf5eb43d9fad18c4fa48809dd4cc99b71401e3a3d891e565b5fc84f580aca7b1fdbe9ef250762
z26a5fa634fb5a0a339d2dcdb76aaf0d6e64ea002477974a8d1921f579220045eec38b2cb2602f7
z5d9cd69348c2bc552093452807135cd7d9380468526edc0215450d2e62503a7ab27451a9f9d6d7
zb9f6c7b2047fe81eb5abce72c56c3946912b85b0dea388a85e4db3ad2b5de844e1d4031d68ffbb
z488a357ebbf05de68ccac8a9f9cb556e079feecce1e5d952dacb49c0a2c1754c1f4e3681fa7fdf
z96ca0a9e9872102774df91c0b5f5680aee9ef8eaf93b6d0e967c8292a8461f014dd922fdcca21c
zd18964bea3cea3998e08b3047dae04a523aa0a1ed048f5f05545e811dbff576032f00a5adc6cba
zf5082ed9c0f28104c27b57601aae3f775302f85a59384a9f1a1ca53e3102f1fdafab6a0495bedf
z0d18ecca3766b3b870bfa618ad2718ebb5dc9251798d5a968e6dafb7d272658af42c1d959ab96f
z68fec93f4362c003915165d0ef2e2a3b9af8e77b65d28b9361674f3179a92aef4d8248a1150c8e
z77aa527aba02b1256bc3ce02f0042a216cf57016008d75c56ab48c780d1ad4aaf59cb6b1395c1a
zb22710259248639fa0f545877954a307c6aec0ee3ae12c4d2b9d15abe09dc03b6ee797e5157787
z041f17cb0e67a19eb85de3637fe044398017843de247c45c2e1bd28f136ca111ed43b9927a5ff1
z8aa13f9ca0271e79a63ec542169de5662aefe8b6db899fe433b39741e9ae8c1b2d23504993f659
z378f9aee91f3d3bc2eb641dc0552211b22407a37dd38fbc16165547d30d93799503adcf0d61e88
z46fd2adc0b93678a586fe8c58b9a5e53fb984aaac753b5494fdfb20b99af77977c4982c8e7ed7c
z8d58c6bd79d3bf7c6a533486394d63bd7e9115ab9510750c8f8a87ff982c20850d25dc0e76e644
z4c38bda3412d74c0882a5ca47c4bdbdf42f7d3f06eab80b952383fc03d12135f1556118065b9b7
z760055c0fc1d8f762023d362041ca6875e7fa9661989bc3be00e8753e3c56309fe50c0de4f78da
z25dcdae44f6543883ae71dcaefffe8bbd9389d50e6fd0f5f30b25336b55ec167811390d80ae11d
zd9757b301c3091c038a5ad6dd1c813ccb379ec64f14b968aa7f83a929759a9c3afd0062d077f8e
z70e3c801ef8e992994c7adddda9dbd487fb2352c0a13fc35638b8d557e3e236888e7e57017861b
z6844e9a46d3b8277a243eb4a85d86c392f9f23def48bd454c5c2135694b6821934cac635553f55
zcbcea6fe0d813fc7ac8f3bd99626c705c03f74f881ac88c9a54321feaaaa941212edfb7972f812
z06f18e387d22a3f4ad840dbc9f66b98ff30b27f66d8558bf413de5495ad4d51a8f40db79428293
z5192c294f923dc85846bf9bd0292e243d045f9a5c3434b00ecceec96bc0e7b792ac9686ebab3ca
zcb3f35d75c65ac952217de558eeeaf8141d3980ef653becb072d6b7d3eaadbb077d4c8c34b1532
z25000832f9d0a13b8e7585ca31fa21229c00b15841cb3f74554be1e72c696e76dae8d15b0b05a4
z286d8708ea932d8a4eb4ae854a6e127c2021e93c30cad0928d5db899f13d28ff1660419ad8d993
zac0203254bf278bf93905c6de21c8d517e0dd68a4d8e2cd815ecfc494f5aa4d43bb55447895c04
z8b59fc46c47805e492a194eeb58c711baff4d398098978438d4145217ce4ee28ec6d9dff8bafff
z52317a6dde464fa0e02ac33c29721f998c90af16d4c467ec3e87faa63ed0a92feb818096c341cd
z257925d63b0d07d64a6fb7c9750c6524a822231f1c1262d79b3b88ccac982b346410f89397d420
zd1359679b71a2b707a92c9241095e6dabf7e80bd99ffe77a647f13a8a97fd62aee70c23019509d
ze75b92a31bd0fda34c7bc2bdb69dc1ce1b5f9b1d5218fdd801fdbb53899d4256d327a0406a1804
z52938ef6b0faa23db5e8a41549da1ca6daf73d809528678e702e4f9863b471af75afca9950dc8b
zb3bdcf1e0baa351436d323f4215ed1276761b91235c62675df45d0e97e57d18d547b95d1ba08ad
z5e73865a6288d2cf73a6602e29e03236346db4bee598807a43225043da03ac60548f3b67a8f0b1
zf5f67b047a200eeb5b0dc6c87500fea89e4702f627980976bdd8b121718200e4dfebfd15b5e16c
z0035d8e357d75d5fcbd174232d99745ece58937c630e8177378fbfedf0e4134ee959a83e158022
za98fece1df51fafffe6b921847dec2e6b9fe9ac5e80fc85565263e9b08a06a854c4a19d126b555
zc43a790600c0866631d327574a7967bc8ab64fa1d6f4035a22db7595db8cb36b0ae9ae9d56c26f
zda01f202dcff77945441f554bad10ebf9558b2b5c442c2222364922194a626882b845cce6132ba
zb4fcb593487e3b15cfbbb138b88c2bb78c42a6541cabacfedbc106622892849c8b71717d7919fb
zf152ad36ca3a9ee009daf21ac5f9c5080eaa4b67cf5832f438b89b338ef9c7a55c379edf750af4
ze8186eb07a5919ba4aa3620a839ca48d974712367c7fb47d0ada172416c99db7927cee15466155
z4996b1cacaf5851fd7fed993555e71d5984c8327f550604e7843dbc5276b132a4231b486694b07
z90926919401944c9cdc01d64ec0ef4e57d9571432f0022d2919cae81d8f041a27adf795a7b53f2
z7fd2bc3160133e70b4d42b18be986cc96e1fb269658b6496fb756ddd4b838341d8592e7abbc1ef
z9e76c6ea7a4a8e432ccf56176f8659334560ef3d525d4f2cb05f673bedbf8fbc68b48f2310c4d3
z4be9a3291097b2bfebc3b6ea0cbe981001e390d0a6e61aeaf9a3fae3eadfd5e4b8d1f82e3132d3
zc44eb2b07db20d2fe793b8003ad9c3aeb920b0f8b361cb4fbdae3c277568129dc5d4b1d0ddc251
z7cbf2403e88624f1cbd9aef3238c1750aa2c94a5655052d1f2dae4de6b814533274ccf2156878b
zc9884aac45094d1356c7284c3167db07729c06b0c054a58e8dd561c9a55cdff58489ef99885d0a
z098b320521240fb7794d7b88a0010888d643926337c16507aeb78ec5184ffa2b8726d11547abec
z5a91973bd7357175633c5f08c48f7e2cca56420b1776095baa88c13250575486654c8bd9e1349b
zeec86b55ac0ce6a49db2b98aea0f8423a68d6c3b77f61c60bd805adeab69b6af912e0dade6e581
zfc275697d52bc312c8fd090a0e400960a9ee0823d77f8aede9b07f9e70e784c1b20ef5b4d27e18
z58c779fdf4cc5bf594a02d04f05df2b7f8631ed6ad760569c07fa3b3ae02a748fa95a68ecc1474
z1ffc9c6da02debee9e759ac38d915305bf791a68533d49f4ca8d8b7140ef5c5f87f8b079890364
zb9c88ca4e1a37a04e99689bee087ba8e77c7a70d4792f63071d9e36618039009ffc0bad19ab980
zc870bca43752c0edb9ef2de7b91099814dfdca81488f9cb846ac5872abff51726d00e145b2d333
zfda79ca4dff8504562321cf8c58babc81a2889d26c8e364a099043e7d99e1ef87d62151e44a15c
za92914f0fe5f029aae04b925842dd7323ec259e15d9f857b36f82ac2c6511ff2d67eddd5427294
z7f9489bf9a5d4c5e1833147213b797a5a48a4d9d102e2174759ef94ce7d5b062fc7a21d1811882
z2c7aa98c83b980073889727a61ecf57c774136e5c1304d4c43721a738292c856d26d323dc935e1
z3619a078b5eb43c7389758a7d70425d3ba49c1d97b3ae4165d6df20889e2611802397fab5f434b
z7efe0afbf9ab268179540ac6e319ab6d59db92701e25cfb7d13a4171973380780316cc2961bbce
ze0c180825a4a088e5dd700e6f35e5e99d20e0725243548b78481b5e8ecf1c68427c2aca95a3d61
zc3918eea73c849ac86439b886dab9fcb338473116063ea155966f6deb119c096788fa55201cbf0
zbb0a7b7b867bcb1ea3949e8908fdcd7d36d0e10a1874dfb65444b1dbbf89a8aa099e269aa05370
zc3f9ebe611fce9ccedddc0f7c166e5723512a6c8893f8a6e0de2b6fb5ff9391f582929d32d6d32
z4d0d4846ac86fead5d2e21a9f6f7b81ba527f17778fc4f56f2eb373ba9a3b810b14a3b14545869
zc5ebfe8a65f6499242aeb7d85d7c7071e10d444614db96323d3a9c3c47866082ce4e08583e1c3f
ze9d7926b706eda8aeeb5f752ccdc01b1f0aebda135ee3c0269f37918bcb98b68d5eec929acd828
z724ebdf6e83069fc7470a9125941047a6ab22e1b5572c14ff7baa0cb79fe18e006542c31de385a
z2cb5bbd56b221805249394e9bbcb1aeb2609a49d27b48027db52c31404050da2422e87ee59e30e
z80ecc813e320487f23aa13c4740544e650aa8641f1d6807484f19c6a41d3c0395a57176228f5fd
z6ab93d5811eaab398dd37ab79792375167450f6d78d28dad5a1600ad5069de71c367339ddefcd2
z758835e3e5b233b89d65e8795e474d511974ff7d0032fb4c4c9361984b6d6bc0bf15ce1a89e570
z4fa76f8238a449cf33b2313ca7efb359ce196752b9765a8587d0a78fac15da07f9522d892c3eb9
z332c1cda79169d96d00135a8bd3fc5eed85e55b7828e906bbbb6a7c5b1fa486ababea8d598969e
z0a6c45ff21e3e5b469639d6ded660faa52fb405d410d7c235eb5a94ea13bb41cd94e1ca6942860
zac9a01c0ea3a1c1ccfe4c57bc757a853474cd923a996d9996f43e23d30b8c95f9f4be8106416c4
z0840865e635894c2c1b9733c7377962b4fcb8e0f14f4eb903cfe13a22cfe27a5c560566177d9e6
z1744d0cfb1d441b0575068c1e38613a0dfb136efadf9b9a5175c2276fa950fa6a82d3f8649f3a5
z6458c89531051aac8bf26191c4f242f1209e00c3c58d38887ceb928371ec1b339a3db19734e15d
z84ac522b9488b0e7a2f23833b7e1719f2e1d67f28e366cbc316f31d6d01d728c88ceac11a4994b
zc5bf91b378b5887c78f39c47d1f1a42e3c0e692fa2628794be40ccdb8091f0712caa1fa3b036ec
zab4ef6f67535e1c99449821dcd3692864d5636241cebaace9558bcb8be3e04e437ee6651a69722
z41325db7dc5c9fae57e636fab30cbe3821959a9c94adb7daf11b74f67fba358cad7fd5fb95547f
zb9d6f5829c64e7e9cee64d09df69d1f72d34a3a129a64d1b35bf0a45173c696ebbacae0df1b8b5
zb1c8aad36a4734471eaed347f16650816d26f18cbbf99360517a4778b30a440d67d0da0d6c61ed
z56cb6d3fcd3730daf64a54ad085a91e104e5b341fe7e8c441b0a8f0cd9e50b3dac8bafa2fc3efc
zafd753855c56cb0010711eb794c491661b0cd6bf127074e431f850053e4bf7ce29eb277f9184cb
ze67b9e6eda05a3b6d71dded1b35f149130044a527da4d8c0aed2800a71e50f2e13ccc6bddbe106
z7dc3574f206a4f3cdda3f13fd111ceedf2a313bf5fa7fac7d01de076fec6c316ea17fcc80af97d
z860f8f6ea7a423bb0d4e67a7673eef3cfb92a23359dc71b1d8900acbe18eb8ec45d12d86b74bfc
z3933f58d0be057f6942f5a92e2136db505c31958ba7c88caf9c2efde73f26ffa12b8b482406251
z2562fc02ab481e143388117c90a5025824f9b70c6d8da3cc5cdd31ce2a61417d7c19956790b826
z04c7604a3d6be05a1aad28e6a99ca47642e25ac8f4b49b086072fe6824e805668582fd2d946ccc
z5b6bf102a5ab9e592eca02cbaa71b96a467ea5a71320979084ba55b55084588bf4537b608de4be
zd555d7f83078d5d3b3cbd45913879bf0206f3a4db9b3d4c0b40d7c5091402cc93fdc358988dfdb
z1d939f944219570198e815bb08960982c25d7fb6eeafe5b2cd98db83dbf2c5b7bac8400e7b3204
z68e124f95e0372a026ca3b29594f60eb0b98397bce5b6bf0a78c9fe8d206042158b1de0c189b60
z8301181fa6ca57aada43aa6bcda6933587bb55a08a76a8f57b9c03bdeed24a1231d6824567b7b5
za0c42ca60152dc872a2bfe95278d368010bd9cbc4ff58ddd2428ac74fae1aecd82b4c67491c200
zc8ee02aed832b00f43b4d1e513afab0374fea130dacb5c52cdd418ef95790d819e1aa8f9e557e1
z9367d5fb9d2696865b5eb4c069b1aac47350b8c405df38e34b1fd80bae2f6429f8f5cc60da99fa
z0e7c3e278fc8e93a3c8fa4ad408d8961c10de34360c8a6987349162041e2a8f24fb864ce9820db
ze9f27fc36ab076cb02cfeb26b1854135ddc5531dd2698a8ec0eebdb06ed01ceda16c68209356c2
z14d476ead8adccd471d9c8febd1346deb28ce49628a891d0ecbe9eea73e4901dd68edc4a1981ec
zd48ba5acab49d654a6e78097f431a1b1646bc280499bc9fd76e5566c1dd8928aa90600752c0738
z7f1243275878b880e8b44376a5bffc576b0607af11dc54e8fb93e85e18b33c881dc024fd820d2b
zf37d9e7120e81c4204239fb28c6d6f73c1d5d67a5e75b616844939306d5717e76739c60c32910a
zbe9c42fc948a08b4fb94843faa3e1154b3a4cb416753278c5a1163892aabd502dbd124d3779918
z9b42a3de6ca2caf7ef05f2d508529daa0a5dd95b2401de4a4ddb44de8e91a2d0c67ffa97bb0ad9
z11d1917e3ba333e96a81ece2355aad227a51d34de83c2dfff3eccd16ec7479babfc591097c0daa
z92463b0babe0fa2a48515fa7ec87f4d0f908b9a9b90cbe2d2f46df8816e957fd8322d4397dd8d5
z2a08732f58901c644a95d7997ab6a4f47dd0f825af96945c51e5f8996bb81439f90013f0c691a1
z5fb8578df24b7e05da2e3b35e7af3a499187beb806e000a59d8cfd7911068e72ebcc616ab96788
z1e2b951b82c1ce5bb3b796570de5f2d399a2c2acd40963e38cf69ce8b79f55a2f7863ce0767b89
zb0be6f69a444af1d8b3d790c17114919cfacaead36094adfe967d1a296b870b377011695b0898f
zfe2e76ecfe70ae184ced36ad9132544e0fb257376defa377176fda2e8d42c7f32851c903fea0eb
z18ffab2bab568b4f69e13214972f29bd1c2a2cf382223c789e08bba6bf03ac85b0982bdfd3227d
z1f0b988fb657aea34c1fa95e0afb3c7677cc3989aeaefe39764be4d3e218eb04dcfbb10398e624
z7ebe6ea9be29226c4508e0fec229d1f6bc0e566d5ff9a21c2f1fd99a0ea8d4c8b3451506142d3b
z3ab53bd753fa471a7a2f3402e464e16b557aa015cd52817e3bb1cd386b8fdd8961416d1a2da90d
zc97bc6cda0ebc46b6171000f809eb7e13943fcaf93c12a47bf7ee4e0e1f060cb76898993c0ae31
zfa51f52f696fecac3c7abbe174a898c404675b3f94098f6a83f0b93d1af73448890242349eb3fa
ze79c0c2cf5836729322b16e5a1cf20c9eb77353289d44ca8555c5de5590757b91b35c496f41b28
z5707cba1222ce79c138a9a842c2377a00fadd78e9a365bcea1836c2dce3f572f36568184d57e15
zf7c10cff77b08ddc7fdcb506214c9d163930273a4da230a4a747bfe0fa5d4240536881c1bc57cd
zcb7bdb243abf946195895f7dec24e933cba35e2af3a4c52fdea82c049f1d916a6cd64841f91d79
zafe43f10e600df3b3fbae75d25f3dac982e60394e08642e6ea3b2f638b8285847b95ea7006eb02
z08a96675da44e07eb23e2f4eb7863c2496d43ffede4b97349df4d942c2d18cc99c943251a3a223
z19f7e341e1c9cece3b41b8c861d7952e7bb2f5b0c3db807c476c196946b2c1c6b200dba63ef781
z167f28e2b6111c7e7974d006b6f8b6a5a1b7f4ae7fe2ddf9bff81d5fe00b18e135b63a04c469a8
z58e4f6f62cc82f8ee0d4ff2308e3007eb6158114670162ec582a6fe23c3ac053c71ac389a72d96
zeba7d2f4403c8d5bd06dc63654773b2d164c16f1f747bf43e7b57ebabad9e1f724413d41100052
z6184bc452c8138a24ce1b88260e33d6eb14e7416bf4a42095a4faf261e4e939c3fa9e90bfe158e
za34fa0c3207fb7bfb6521c764b60cdd382973867ad7cb39eeda680a6f546c0b621d9a67ca0962e
zc93b6f40b34cd621521e912573d43dae33e482aff80f5238df1640da2bf396242928a15420e3b3
zb1f5b7fc8da0adb35a7a9c53168a3cb8cac728a0591b95c5210584d1e774a2e565552b9abf765c
z49d8e8bba176aea7e0aa94af7e395572f442e8ecc84752f442a0683a634d8f40c16f14aa3bc866
z515dd6074f0389b2ba524b286db8e2807f87a793bea9810a292af27f30e3c9e0379900622b032b
zebbbcdadddd9f83741c54a990cae7e197651b297a466581a6505cc5adac9eb48f42313ce053e31
z3af67a83efe4472fd127f80bb4ada50260b7a1cd73f481f5f29aa3f046d6ef56bb8dad213bd316
z58c7d97883b210f61c2c1627ec9577b246d608fc431e6abaafe19648b43af8a13a00a1c8cbf202
zee055bd7a6ddf977a7585a7e9a8886f176c94325be0b59ab3fe058586055fd893e11f816ddfcbc
zd451ebe0cc7d01c238a86cde3f84eb9fcd3e4cbea86b82447d14a0fa5ebb3650196a92f769a0f1
z32caaa3f4e076672d0d91f357b2fa137d4205135024346ab133c19c78ef7efd75342f0ac0b989d
z65feb80c16e85f7d21ea18ecb27c2ba037cfe1ef202c6849d596939feb06d7cd9e3c9b49db4f72
zd1ad561e1fd566e4eeb4201be4ad8e3c79789f3d159ee6fae5d7b924de85af1cf4b8b5d78b7a1b
z82c18036b0841dac085da98414
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gigabit_ethernet_xaui_link_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
