`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc89607e51
z10be237a8e467b1652b13d902d77ade35c75f54af54a3a25edb5532d5f1dfed98cc3457cb305fc
zb8eaca599f16a4f92caadc3c4003e9e85b584e072fba51c103aef06f0d2d112ced5770ac12804e
zae87a68e263dfc3d344610321f6959f787c7217ef3b6512dbf4dfc7b803f1a05d09ced0639fd78
zcc21a5cb1439fe44e55f89053a508a7df930aa70f350c4f77b7565ccf58a5b7accaf1e7c4d26da
z1c7829762218192a83a8d00ca75a4c6a05b45585ebb64ca409fe7f998b743ae41906f99e78f7b0
zcf1408f020664a3f0060c723a750afd3be35752d5820b179e28f92d1228f738b4c3a4313f8057d
zdaaa51f5e79aedca1b88f43a2cb2427391daaae2da41721c8879a1966458943b1041c18ac5e164
zc7d88b6e69eeb772dde7a3f45da7fbade1d7267e5f17ad10e5e8f1a3426c9f56d4a947a7127896
z35e3ea90817a0ad7bdc3c0bb780d66219bb4bb370116e6b0543105782455079ba963c79f45ffaf
z0827c96dfdfaeed1eb7bc79ddbb3f7a19305adba2471c1234191158e75d7fd311c067be0a7d32b
z3d571250367f7efa4f675acf3787bdbc33e773bc629e3ad64b5d42a846674b144152a44b00294a
z6df3969a7fe73195bcd11be5ee408a04bdde2bdc0191ac0a1101991e819c1ae4a8d82b8b7d6d85
z839ad08f57ef99d692fcc3a335dfe379fa03217b633dbce44241e4bce46c8078d07d3c7deab872
z37f9217ebab03910adfd3d3515c77a1135dee97f83fd554190d9ffeb88f3f01ac4e800e162b5f2
z2d4bcc05ad8b35800515b7be35b7e482a2ed03754c448f2d7fb4040f39cd0ab174b2c537278230
z260cc91968ec21f15892e29e7da13eb9a9cdfa728364683ec87e380e41e2d2207293d74f99a96b
z4600c5f0946ba318e8c8b2f56034b0b396248ac03b6303e536a46830e00434c0bdc8d08064c681
zdd650d01f91ff7624d146d3a4f7631b4ce09cd4dec072cb0e1d0a44b79f4007dc4ce323f315c88
z07612ca35fa33830edd5f65bcf2012028af07cd3e9ffec645894bcc173be6433af097ed237e6bc
za2ac615dff423a439111425050687d5b05ba3bbdc6ccd6e9e7c6bc7ee4d1330279d34f4d6e45d4
zd4d5ae968e2514f4203206221c51bec4067552d641923e094702c2a85fada2639f2d1c22c118a6
z7bc8c40fe7d670d8c80797b06e143008ced8488220d0ca82c7510a0bfca5d5715232d22d35621b
z166e505af21843c97f9d8d9bf7d35f38fd8d4a16a481c83f7da42e3e89f560a11a8add506dd5a3
za32464be3aae437567f3d49bd1ebfe138a4c78b10c02bf7b4d9c9b62f1c9c1df53aadca5d83431
zb9dd831523fb27cf784d9e741731f40c7438e68f9ca41288fab9fa0c71c9c651408b8ef6ec1ab4
zbd7a7888254c417925ede48702caeb326a24f5cfa5b20800906122887142d4fe29dc533910e375
z24c7eec5bf04769cec9aedcb01525241834598d822953eae51ffc19f6c48bfad0afcbcd2e5c91d
zf2229d889edd134fa4beedacf7793d1a5cd089ecab4db4249e897f1e3a92448fa516aab23cf636
zd0936f70957443d75c113a7e4171be2c1bdc9eb03ad1a8de04d6aedad83372b63f7f081affa7bb
z00cca930a5fef4aae0017c636cc52047533e3243a820695fa18d338d0f3413b1cf53b8c509a5c2
z48e23e07742cc4502d61684c16b81a236f74344818dee5679071d3b1b721c9acecd26c43d2189e
zebab5cdf48fc3640310f04830f0b1f0b04a8c92063c8eb0bd472b362bbf0a3454780503632eb46
z72e9eabca76d128b5d4c7341db94b4fce738cb3436c20777ba51ed6a13f83a0c3d9406e27a4490
z441afaaa10ce90cfe17aa106c0098939096088cdac8776f6de3be048f6aefc99d4418afe0a14e6
ze4cb3cacb66f6c6c354888f272c1de8e87380b1774598b9df6874da831be411bf8be71a52e893a
z1235433489152e6d6d78889c0249e417d16657f3dac8139781d5852f3c7f5eda553488b0c81831
zbbd45b0112370ec5fcb9ea84f1c503f49865faf51a29d7484f43f8ff2d444ca56f1d830ce715e3
ze5f5a9b8aa4b9ed57a9c290fc08320285867f09df2ce076c9841227e9173924fafeb7dc08d99a9
z6ebe9700a4a41821cf0be55ac5785b4ba38308c33f08623f11872139fe86c4b6ad21724c2bfa22
z3eb52ca37bd6c8fbe8f9f3d2958bc9b0b4a2510269b1fcde9e40e0cfd381518df08a4f4624f62d
z63ea7141965b2d5757679fd534d1a3141b6a28cd18b7fc97bd03cbb04977bf62a17b13f6f2fc9c
z07f0297b22adc9a46f18ec14abcf67ce85184c4ce1ce49731ba71beebf535abfa8a7821e3e6e75
zce6efd9b750d606c57590e2b7a8adc572453cb596371665009941f34f106d60bb98d3412ec81ba
z39da6b2881572408dd8462e18a377905c027f13569bb16532e34de805eeaef5e1d0f24b2dc7e95
z999944ffa369441e38dca3e14d16557a9c78d08e7c8d10e2bc6c9faca7c71021932ac7827adad8
zdb22f7ee9e16f826f2b6df6c700d8941ea9896dde0ab0f519a3f54e73fcf96c2a6f4c2a0fbb583
z2b85fcd5c37cdca250abcfb0dac8678604c1e2550c799c588c5d53a242f3386e72ea25eda4dcd5
z68a94b4ac6250e5766346ac7f192df22fcb0ae1f92d18ea4a1e33daff9df9bcfc393beb97de5e6
ze7ffc468a65bb0da31655e6c13b4269c4360ab8a855ce03b571ba1beef4cbd5418051860345774
z588c39dfebca6f1981f707f1be57ce83b062e9f713a75693ffbabd6a7770a9b8dee914000e2dec
z8604afc700f67a6f583721ef5554e206b9456d0535871fa3d3b298db76ff1ad5d7a85c438005fe
z821412d2dea2962a218ff8ca5f5687f86a47380fbdae0a29ef6cb4660d2f8bce14e80312384a9a
zc52d4e80dffd15882ae9989a3383e6bfc57906397341db79042dd20ffb632b451d925932b133c7
zd873f2e9198f1ce3dfe9d5e7a5ff4c10fe7a3eb77ece61b0c2731f121640eca2a4886a8937931d
z4b27cb48fb3994d7af8799c3b3cb5b7a5f5225184104e60bf477d8ea5dc0436e23f00f39344508
z688f648fb7ca1827a5bc53f60f8777fe7dad2d21894d4efd5c3ad87269f4d253655cd9cd02e1cd
z5deed8d5d77cac4a0a3ad5d4a631728900d7b7125c74501185af428fdb148930b5c891399c2b31
zbede172e2dabf9199692c6ab953399798a13402baa7a1f3089b682ecdd0f462d9a0f9af0935606
z6fdb56e43f6bc10a46344853162c0b2fac3c056748a61dcae6c58e60cac4a17ed08eeb3ecac59b
z0797d1c7999e900b6219ba89c5d831e788bc41fbd16463eac86293c69b0e8a92ffbfa97ef96d75
z8d762aed24b94f9fb8094773597866447d2f59eb3e61018fe2d4678a79d5195b2db65563960596
za148da6c0a4e69f9dad1d186cb656f3502c5a871470405ee3e366ba79042c02d2502f5fc5d26a1
z749cd796bcf14a07fb908075f8faf3581b50c5f3bb31f11b6eb7bc540311d72b0599b8a69b8eca
z1264189dac40ff5c5a15aaf49addbe1b8541be400e737c7ea526c78615e072a535b4818b228a81
z38498469cf3c221df03d10d410e681c2bb95657b5b3a67437284886dd0a7d9019d59fab3979ad5
z51e8fba586d7b12e6fa746d277f7c7fcd6fbfec8e8167289a9e0374ed33c2e264e172627492dd4
z67ed380c5e1a7552599f4d758014372cc44fe923ff3323ae056194854caa1188b774be29aa85cb
z46ede0fd250f73d6de8b0ee482325fe50d45e136f0fc460b035f8f44a274640e89dd98ab3ab41b
zdfa1c7a7eed2fd00c075699ade98aba2f007df3957eeb307671aa019f2a29c8e8bf3f1679ceb90
zf3e49c46f6934791f6c3a285c279445f5fc6a2d39c8989a1a6e6d07fcd5151e1cdc8331432b439
zdf3a9ca53b1a80a70cda56c0f878150b73d2087bea6a1d10e4d6e0a3ec9e5524a4c61136660732
zd7f3f0a9d734013c0995b3e383b70694f618d5e631eac47d29be20ff8645d8eae1ad7957cc1de8
zdc5401dfcbecf03225f8daab95895b67b4da64cc86fb918c9e4dc6605ecf6dd2d10ded4335adfd
z7b92933389a802dd5b9c6f7d7dfc790151c4d12927de15cbb800be5f7b35335276a31ce8ad1c2b
zcab14db3bd58a4da72ddbc762a480d1489a40e0e03d32b865ea22126ed6a18c361e900743defaa
zd733f686923b61229d411e3ac7ddbbff00cbf7166716d167c7c434d0a7ffb56d4082b1f382f634
z094fbe9a6b13fb05d8e39cf783be849cf398f7fdf6bee433bfda2c171bfab419b0de54a86eaa66
zb2b26eda29d0c5fe15eb3e732aa796120b5b155865835241f5ed9c6889bb3d41171bde13592cb4
z2e3b84a2dbc0c80886f97bda84c10f6db1b1be018f73fa629c7610f6e101c0bb244d12f07d6cbf
z80433dd973ce55e7f40fba5649c40838a261c85c263c1d454321488114983c4046091e2eeb291c
zfaca8b5d97098f490bfbc0b0b07ae935b38ffaf6c91be3bb503b8bda573964efc7e53939806c56
z1ec369d4b853adea2a8ad6c14143bfe84cae68f5f775d8b803b39632bc99fbcb444eb7b12b0e0c
z4b736a1cac0c843b520497062f5cb62fcd0c65b8cebe5e3c984d25367bb3c54600f743cc035f28
z5f70dd4a695e0f5181ba3c3db5a8a13e891f17a119a5f49c1298a7fd6b96750e143a9d368bcad6
zf6e93a47f120139565d569f289dab11dd152dece536b59d48c239681a8c2270225be529d179e4c
z6cd5fd7199bd5bd165772a2663bfdf23474d3fc7a48257925bb98c8b9f83306c0779119dbb4fc0
zfa134dc5aa3e2135d2ac52592b6248de0a26efd6007832fda328821296c05f91b512a140b35a93
z5b8d2630f72bf4cea3c6f3482e8d9d3c73c43c4b86d13fba15542c7171679ab712036ad986f6b5
z742cb7f9877da5aabd5039ec446fe93018a7504c8c32300778616fb965f9ddef5ba3369be4c673
z4e5686485ab34487c95e473c19bb2c6c581ec568040318feef93a9ee0b673430328f3b278954ee
zfa3cb6dbcd2e7f78a090756e10680dcfb5ebcd5a5155018b83142109071435523e238011e5189c
z22ca3eb22decd66aeffa2bb73ac218af40a5f7b3ac0c6f32ce3b5fb3a76cdbb15c1ac79dd145fb
zb17c2f011fbae1b2bbad2bd24bf6f41b76962c25e98536c7301e10c4069f7555d2c14cca19ae09
z7884f0f0c9761dbac3a5da96b50bd7adb128c83c13f4adf12943e083ec1929a31fd14505adba78
ze12ee8a408d0183edf4e49f497eee5d6d53dd35869b7070fcec65c88b55064e3c10a11f0c12b7a
z068198ee62e11ef964e1c1acdc76832814b3e11efa0c23ecd63b2538a91bac1acfb586c9d420c2
z4dead05879f26684e321c5a0e6e63e9b359dcc28d41a546e7c17491d88965e0ba5166bb5d817b6
z061c8e4cd79915fac1a7f461203bc977b4c7cc8c6f4c1934676b26a57746f6dc2ba69e3ae66d53
z51c0c583d9869a4fe7876cfb4e83236ec86718eaaaced209c9b1908378652c48a394fb90af943c
z5baf1cf550418e37c090f83fba448d024713ced42c0380d375c2a9a9a533774d57d215299bb8cc
z6f48147cb0573e7f00be12f490d14372b2d6390af075014e8b1d085bce38fcaf48a0bd8ef03485
z237c8ff14848507f5d92602614fe2b7e47ad88829a78c9c667fb4690cc9d596a16706928b54bbd
z8629d7eb3ae7079518a5568803bc1eade22c1365f988ddd90e23b9557ad2b70069bcf763a790a9
z79e6a3239ba819fc9f3668a9890f642f0bcd17889f6a7617183fd03bf4c013856d032b5941fa3a
zd12886f12a540edc1e9c21cbee4b43ad693ad37eb860f87ca6fbe42608e7d616891721c745b3e0
zee3b1a6b919e20fd75dae0a2caa564c0598f2c2ee147a0bd9f0c0caf41da83f9e444a3534cb6fc
zd819c238c796bf794f16f3e3536cba23663ee3481a1287eef41651745ea2193530ab376a967a97
zd88b4789c649ea0df18b45fbbc22c3f85a92bc1e37e9b10cd48affedbded89086629c04d7c03d6
zf4d465568d8e09e40945c8f2020d7acc13b8c501dd08ed944a84050b22d2a0212c4a2f5a2792c7
z822b10511816f31c8e06e07e6e643eb3dd716d8080f04d1655cd8d72609f19062ab885627a71fb
z2dc99bb765e6f7857a8cdca241614e3156aa6686ec036ffc7be5c18339c9bfaae65da750057631
z22a53b4a9c8c3b0231cc8745cacbf32445c03d8096a8aceb7e32b38a34a6f90209b76378194028
zecc0693ee5cb1643f94ff6bf6c20d5f1ca0817b9ec562d023f5c224d060abd3deb8e9f09ce89e3
z1653be821545c9a4b0776dfdc19e10bc6fd25eaabc4e61aeb8d66e7d3183e181d3187337e2a375
ze4fc36d1d5ea0a8c3adf01dc275cf866dea25111be3636698573f974cc74dfd9fe41998ea81f96
z0df474310a42d30af0fd3ca17a4a7dcae49a3d36f28c92be4f009e957c817b4c8ad7a2de536d25
z90f8108fd7d753b569d95f4b7f223872b3458084a5afce37d3bb0f22846fce6432e804816259ac
z61e19adeda8af16f4d3ba112cf0770d724809e9efdea450b771f0518daa53ed57ec2bf6c3058f3
z30dbc17244cba2b78229c5da79f84a5962661d6b35ecd63f7be659bae7d0bcb8f4f5b2a4102fc6
z94cc291c620671e364cec0078beadcd9a996fe7a76caa92cef18470eeec845015729d543393f73
z4991897a458b30982ba7c2413c92edfe546aed3644db7127531295b11ddec456ef33d92c6079cb
z8b5ba45e73342c59261d4658173efc4e154e1a2f7feeb83bb2b4f773a2ac2856368a2881083d2f
zcbee9867a56e1e971703946ffed46719a624108325b5dcd13e4cbd30d66070afcd3f8ea99aa15d
z2bf136acc78ec8c4cebf1dc75cb03ff12ce090a17c7eb0ab4557581efd13dfa1b3f7c8ac6a6d23
z9365b39d5d4490280041f1a97d83218847b30b9a8ed2c31f559789a999378fa44a0880790dd7b2
zff28087c8c8803a27ab12a27de3693e57f71888e26d338040d33d6ede86b66673bd0d188dad3e3
z49202063f86a8209ebd9cdab6e3a8fe885ed87c84cf1415658528f9f31e258a39f018244636de2
za4c5a41dbd71ce40c24c502be9b5e75aad9bc6958ad7ec7b226b3445d35b69004beb43aa6f49e4
z645cad68ab4a25b55ce163c8366ea794199b7e9b494c609ac553165a1ecb5b28c5c523ff899289
zd2002c179cd254224c58b875d8a5a01aabe95424cd6ac4b5626c4cf75a22f46b3a9d9fb51a38cd
zc91674704e423be12b3066a8766acb66972065ef2e596ef659924cd7244e9ef7399ede227c4d22
z720ce41878f5c242e7e102a4f3d178a5dd452e88221e98e473660fa559a0e36630b65c75e25cfc
z6187e169a317b4e82298a27f83e763e36df0713ac30e878882c63464400ef9db2a115c951f201e
z5b7d7f32088b022236e5076e59554cb1ef962a07d1bcaedd91cb0b90ce7412dc20d07b354a7d64
z677d2cf4f61021f08fbae35986ccdfc4ed44e17252f20d476c31e21ef81d8107e5b873d7ae52a0
z35f821fc50ee8ea322060b53ce93347db587408ed7ea64294e7c601b0374d68322b7f08f17fb6c
z56059c8d47b614c8d6a72d718eca7cbdb5c656d897a1703fa0fb17d1dfe18b72457e479682e2cb
z163a80dfafc80cd49ba319772e885a47f32c45d5ae60f2845f25b6ced724077cdb3ed3e4c70083
z5b0cb1f4a59e62147c87302d0bee32157826eb3cb3e7a449ec11e21d68e0b10b09aca548ef9580
zd25c982a98222455a6c0a46e4cf99e5a5ddd5901aefed06ef3ddd50887107027453f967622560b
z4944528711dbcf3e45f80ea8cc0efe5cab02d81cc51da3979ccb50daf55fd56c6e2e5b6ee82be2
z7e5b9f5871125ea11551e52d5ec4403c39fcc102d5f9430793afb46ea25c26326150d275f846be
z35ede6037f4a5477c4130b352b53102e496e5a9bf7888728195494c88863c03df81398f5456a0c
z4de169f4d47b09fcbb118652e90cfd049d38aa10b6be783e38fb6f0afdbb57c57332f7a395bc1e
z33d831041340a22ce0cf4cb05c3a1fbee7acf79c9a354d1148b9b07a2050406be1c7e2d34b0c13
z6c68ba15554c8856404f338b6d731c9379a13dea6317d1592c4f0c7da9f5c6df2176cc96c87126
z762901ab222b9669f4d650e246615ecb34f6fb7437e86759c3fe51e6cc44ab02823f09a112a80e
z24e000281399acd71765963eb19910564f54ebdc9577cdaa0baf21c380a8365c9bb0880bf052ad
zabd53a262d86299ce4f4944aa098fabe9aa53333deb20ce304c39e046a2b26cce9bef13c63bbf9
z246f4afadfdccdd33172f83ba6fbc1b84dad4815ce030e49c96341e37a9d89a300fa02c172aadd
zc272428fd005ab0ee6d2d0b378a302e43e4f2029b90bbc83819d7f9f39c9c4581d6441064210ff
z7ed1606a24fb36df809dbc7497e462cbd17e83c4cd2599ccf72d997eb82fff5d65284067378093
z02020d26ef1bed306c7d9d17f4264955ff9389fb3aa98b1e9e9e86bd94cd7b4aa73850f7e4d4a8
z6d344581776c67cc3363c271bd6c561410a025fe46fde90c721b8d16b638c68fccfba354e9d8fe
z54b156b3450ddb467b4ea1cbe682e80843a24ba0f9fde4357fbf8ee59a0a25ad97cd98c8d27905
z06526c16bf001ee3d9dff9fc5cde74ba632f94014da32a732eab13ae049f11833b46de2a9d30c2
z02c35db50ffc9c99900737cc7fb8399ff0c97fd41a038fa16d4fb336410926302ae87a3ca2196e
zb298fd1315b0322fa78f5f46aa58272d06a84c78acc8187d03b5373bd6d2411d9d6b4ff10bb031
zc9201d577d93b931d5978a9a2ad6847e9638ab7b2e5ed4e96da6e234a48a167590ef6dc77142df
z7ee36d0f8f0da3c80c19be678b1e8edf457e5741deb279924fb5e2643405a2ca87a5a9df41defd
z741c05d3d265799a5aa0d3e7ca99b9740f31b0a2d4f2bd6124bc382eb2df9a0344cfacc5bbb4ea
z877a467476fabe5c3e84ab299448650a048bedea64575582d663f37570b28dd77e966c1af70a3d
z7f521868c64d72ce22f043e071734305ead48e6d052fbbb35c435d7e40fbd2899bcb7447493ecf
z3ea2fa775e67d7cf2bbae734611c26f731a407a56242810a72caa8eb084d59fcea7e4723440ef1
z07d93e8dcf337c6c45a7a82421bc27085a9488b7e08ad0a44f6c70e7d7c2ef97310e52cc01228c
z97940a3ad08cb515cc2d36163800c902c7697f84f8f38a2133f210d566805ff61af141c193485f
zfaefd508ec4450664466e957f02c0890045af0da11ce8040da1870bf0bcfa0bdc26c5a03a9b00f
z4471d525d010c9a41d5dace78eb4e8ca930df3b26643e91f5baf24f560005e05a34b46e14dbe50
zccafb59c123488b7e706c6cc199e74b85e044b54f8fed8be64579ad8d9febdf04fed75241db59c
zf98ff3290d83b348cc315f8b6cce24981ebc3a885baa20d481392f9b2d446e63e7cd4f5a6fa87c
z2c2af0a785539aa2b59d0ae86756bf04b684ab864f4b84c40f6c0233d4dcb4816dca5c3a6c780d
z879924b9b194db589fa94ca6c89d1fa4d6bc43e36f63f30428faefe8eedc692939a12d110cd019
z6f800463be01400c51c67e1c9f0d9b4b08b5c34308f18a321147d371d0ff075e54cf7e9b2d5ea3
z98d490f6364ad9b3dd6b1f6d5e3b7ac8a6460caf477f65bb3a158200377aea3fc2fe6bc67cc612
z2de622b4ca12be127dc838fbc9e9e500a42bde52139bb61e8d30c7cd974a6c15f91b5e57eda838
zb7ff37388e2fb64e00d4ec68297951ee170e2fb3119cd7edb54ab950ddaea953d94d7355ae3713
zbb9b8cb94e425da70761e82709e3f29580c9ead385565d9e81c209571922cf727df6681285d005
z11582d5bf78fe59e434cf001dcec6806f4e95d15db7e4f04696d24a44d1f39e27c84716328949a
z6cdf1f56e5c20d6d173efd7bff20b3ab3c6fa5e29becbf9242a64f21887e6c93b8a5ffc9a570a2
z64f9f0a66446153c0e8a97a7e3346fd02eb234ff700c0827e0ca937994fac91d248273a2eb16b7
zef2ea19435414da8a6a5371cd5aa27fbd6d16b12aefabcdc5c217e09afd52806b68fe84de17516
zfd4d148b12ec3371e670fa0801ab456de4173b6494c07063cd407f715459673e3b85eed73a4a76
zb8c16ae304d5019464fa2bd118f5cab3407d9c359da9732b03c9b2b5f14afc9fd984ee399a870b
z01a953173d6945a0eaebead25a37b23f21f0e62e4ca45ac90010e639695c6d879054cc447854b9
zefbdf54622cdc779deb9635dd3f7d465b6659e7d69391265e68cc06f86f0d29de916f224a2abe7
z4e666317bd6b5d8fcedd5f40d80a8141b8f783a050849202b5d23c92c4d91c8ce7efbcf3b08356
zabc5cd88583fa54be6dee46e995b74a626a16af851c2471889a42652671045a492fda80b53ede4
z83db2154a9569a0ad41ac833c74501f113da300bee74510346b81d0fe633b29ab85302cfeaaf4d
z1ce66f03cd3ae21f1f47630868a69ce549c7f1a5c615813c8014bbfc0d7e00c4c0eb2470f7d13a
z5b5a997e4c4adf47feb84e5ee640fa3392a56675ee1cc8ab77d5aebafbf12f3a0f1a1e58bc8aea
z5927b23b57b285044f73537b5e7551aa75d44bd30e5e377160c0a43870a659d2d7d976ccd7574c
zb096159aadafe5b6c05f930ea9263291979a4988bc2b2f4e94e29a012eaef2cc5b4e6d1a74f9b1
z3fc1ee4bf5129cb4ee5c99a7f99b626294f8618ed3ddb8aa16f9c27405d3ab69618251b06ac6cd
z3f6d024dfa5b7c69a753ce4a44e081ee1ef982d1ef576ca7af8646fe493bf4407475a223aa21bb
z4d899ea823823b18579b3c00279f1c4b08d84bc12d1b8ccfed391e4b809e03f4c1210ceb983a02
z53990b137bcf47b965d28771c65a486421b0637f1fbd7288554379148a77ee1343018fa3ae484d
z1eb08983c533b6112bb4715b300ddcbf6bd8086430c4b3f3d6e9f8bd3ae7ee99baa8ef7f4de1fe
zad2fe8aacc4840a992a5070216dc18e2d10828a7025b2166efd355979c67ebdd7c2df918be79b8
z57ab65fbd0d8ea2a68314e505290f64564d2abbee0220d42d5e4527ef57af0ae23cf6ebd39161d
z508c968a123b04811e0e766c8fc7d7dc6d1126ef7ba02115f119650efe3707e29082e3cc0a027d
zc2c82bef3c00e3e9e4b3e6afa3b333677bef24728fd45465a4d4e09f0c2a8f73fe8fac65d3164a
z10e4ef4ab5e5e0cf40771a98e1efc83f166b7f2842fe31a9be516129153aa394c0dc7b4536d62e
zfce09776fcd3855bfb285dc01bada324d075bfa8505a4af0f2642e457cbea6588b4ec21bbdc593
z220380217d7274781882d4db2a831b985967a1058865707c74af7cb8e19142e0c57781c512327d
ze02a096611bb4a28378997a380c8c6ecde6c7931b8904c3c59646bcaacfa62107f9673754c063f
z75ac259dfd181f32a856fa7a3aa5af3321085cb575b123bb3601cb812bb9c258ef92c750cda291
z2f8d1b2abd3fb1ed6aca0fdaf5b5e4843f342734352cf0ab0d801f18e3dce7fbdd3af2fb049ff1
ze24ae799f87ef07b1b8590c77f60884c354d1ef37edd13dbac877ff1533003212cd199992ba2fa
zefd3ab63ae806ec88b9b9328d39a90374726f8b336709296a12329298782de7f55e1f50f30ee5f
zb7a6f8de53c986dcf94a3be7cf2cd01af33f566f8250a2a3596a25b946c358135271994a203b39
zbed128f18efc9c73615798ffb212fd12825b6fc33ebc026e7d75f98b72bd8b8d1a9f619e8c36c3
z2298c1ce1db7c27d97c4cd843d31b88a2761b2e25878ff99e3cb2c98a27b5210ddf281965660c1
zb282e4cd89fad5623fe969c36c703d7125a3e84857a98b0445a66bee5c9129d6cf64a4112491d1
zf7c68e88b9a1268c85d540f13ca04d1367f23589e8ec517db27e0c07e1abf3b88e0f7d1de69ffc
zd24fd04a617a583cae1adda0e604b656632cb0364babc00d626c99e44a2a360c7311993baabd58
z3ff02f777bb74e26c7d90bf2bb1e3cf5187c42d947d55a6e15f61381031583b10d26c5ec6962fe
z6628aba89fac69999bc626f6285511c4100d7adc384abb5938f600277b9e2c8318b27ae1cbb658
z1a099e843348064df1a98d1816eea11f7928138722af097e6ed07e3b670c49ef9f732db2ae08ec
zbca2cff305a500d95ed38dfdc66b63d54a45e9386b95b561b942d090413126267fa50bfbb33bae
zed7e7c277dedac0de07d63b8082e54a1e89388f68a2375cef9feaf7f353db9d6f0a1b0ad3ca3f5
z05f26ed9c006333a4584a40040455274b617e2a64843e30e11a019c8a393e3a4731fb5a57f5fd3
z2ec9bf7d51c66aa5a1298520ebf31375e60325896d4d8f6db7b171059ea8815a5d0fc9b366f44b
z3b4664208d4507bafb91e70c4e06f39af2317584583c04abce4647d10eaee67ec932abef77485a
z9515b93dbbe5c0665a9ce03445cef57c662b0cec8fb7564aead61bccd1693a971baea84fa0d76c
zadc0564a1adbf2cde0a02ccd0079b5896296b8551cc2cec1d3f2cff477d80349ec84c6b7744753
z7f62ebe7c3de520bd5111a79e2761f779b8efa98d2164cd47c7fd3fbe1da9b3949446bf556df30
zba73d03f16efbf7d904d1a7e2d1dd315162564d3dfb6e3c3291ed2a2a80cb3e3c9f2f1b8c2a62b
z75d309d54d256685601fc3ac5cbcf643f8e909b95c107c6a0d06ae7a2e1b46d515ac32bb06b7c4
zc022b8c60c77c55d36680c1ac6886dae8eee8b70a1b91a45d1e30f965a899f989f538013eeb7c3
z7817a95a6214c2cd3e763cc21ef7d6b1054883a4dd4d2e70f83022836100e45a0594a021564021
zf19cef311969d955b94f604056d3bf38561e056d98e9623bb2d70eefe1e0f33f968602ff4bcd86
z349164e6b4af3017d954503f5e1926ea960f1a2e950419f0e846415c81890fc3acac932ba7c9e1
zad8c1e3662adb55cf7271dcf8fbb5c07ae7d4d154a5e2f2f21418f52833846a607df05dcaf6c7b
zbf80d46a006c048e36edcc8ad887fc3082a0f4ebc1dc2684a91f97de23e2c5e51da5684dec739e
z51787eb674683b7817062ab5494be399dd661b9abe83ef1edf6753fa8111bf7129e4942ece63a7
z271b009eea1fedfb4958f342e3bb47e28c4a7230b1bf91a2daca8837e2f3daa649be76bafdaa17
z8560ca7923c98e50bd89de1454794b65149cf3a683191aa46ac774faf6e03e055ed2079d68c6b1
zf8dec7ab8caaa23a01dea0516ff418125b320cbca03310d2b17b297083995c84cd9a556999529a
z3a61647446b6225dd95f74f98448141b94e9e25d2e850527a03278d213d1aff054abbf89e59016
zaf6c541c702bdc47c2f55a1a00455ec1b3f5ca3fbc37078c9805a789e4926b339b9e95b439fca8
zecd14b76216ad61602c816e0fa3c6a150d64c23bb21b339c2e797edef66b3e8bb5084aecfd8c60
z2e5b822a6ba9ec14591478960de7820eaf515724298be8d97bf0b22c5d7d0e4a6c94d17e453955
z1a632290031115eeba2083beb3d283c56a25d44828ba353da5a216c2dc0a5b81cb6ad09b244426
ze00313d5536a96561421130423ad213a1b6f6d07cda356a04637133c6e855647149c9c7950b937
zc7bf956b032018657f9581cdb9041aa008fa6647bf5d3264a192b6f3819f0d251a375fa63d0bea
z61b4ce69158d69dc95d1923f42fd533d507e2b9af0e194dfb36e4f6703a10bae26cca6e2102379
ze107886c6fafb747eecf531b59062df7f8dad3841340587e6232b818f69adaa0e2e0f56c32d5ab
z6125f3f2c01761454fe40cb91cef7fa439a112ab76328b39a54eae995f4dcc11a9023a5a721f70
zf1dd3908a57ff7e1df5403a562624fef1c9c2ad8fd80676f5c957bebcf0a5a48c8c1418d975e55
z9e774885c9422ac440a2bd12f3bb5a4403156b814a71788daaa88e0c48a893b1783abbf1ddcc1b
zd2ca831924b678e14b72edf9a5776945927021986c5e529776b995bae0b689cd9d06aa1d06e58c
z7c745586d40ed5758e8d2c9159b4f4f7321b233b44180112f2a6ba328f1d1c60c2a56a3725f466
z9de9feaea7f1a8ea7a834c25a0ad968106379751772d438585111dc8e9666756056df5ed00f75d
z99caab54f2c3e8f5ca8d2773d69df1803a518c252384eac9fdb8b9715ae28deab462f39c06582d
z4c37bd777350d3b6267a5b7882981090160d80193a863202b1406394b250e90b5f4e0084822449
zf59c94c5668dd97636d0ff40c39ee71c2423e93c7a5090b41634168ae918fa2e01d8c6120f7372
z1e79f30e06b1b534baae4e75e8ea6bbd3ac3f2a91929a2e028c458add9fc638bb83e35c02d25dc
z6cee14f24548831447db2c9d2f698b62a3356c900a9fd8442f5259b2b8bf8c9dd715a39171e146
zc9184b138363af55661b4344c2580a416c4c5c8e352f0dc0d64c4f0b93be0cbb8b8e4f8de88a73
zbabd387c9f790e7edde3b0c1a602687d6c2f1fadaa0b0149faf3cee19c2c4fbc765a4b69b4af6d
ze147953265eeb32d780326ba12b70c668969d75ff2b2ff93bca9d51e6f4c2d09d9800ee9d178b0
z1639f87c0ecf30988bf9f8863ac62945f416dbf3dcc4b6a30904cb793a87a0ffd0c290d3708643
zf545b2ebcf4798b870f350b8f7961c40626508d4b3b675e3d61c227a0d8f566959945e4b84e630
ze03037688cfef3e53f76aa171b64aea011408490e10928cd3a03db581383bc62fea23845f24d9a
zc16bc23a99a153e4e3710d5ef2eff5697d8aa0ce4381a54f52177257b1773e39f994a252b0e071
z3e699c6f31dae61610d8725f178d877234189e9e3bf22956674bf130aee6d01215b4ddb132bf06
z7c57b183ece8404de25606da63b1d56eccee7d4ce3b3528af598bcd4cc2c8a7eca86efcfda8945
z54c2b9c7e67ef5b6103491cb67a6468929dedd4d903d3274e046d4abd231075533506014e47ccc
z31eca48d58aa2f3495960752b531d590f81053bb3beffc8365bbababd6d1288eab6caf2d57e805
z1a02a781510130c1055cd7f580706c1421bc7333907ee32ab9be4f33bbc1ca2c3b4341a857c96a
z095ddafc8f0dff4c85e661de6bd6e90e43d5ac5a9fa4880015e38a2f2d7bbd3a03cab7863f8b46
z0d598040e517b0ffe2b2f3e6fadc515e8020fc0709cc752ff00ff5a6fa7f7e14db5c1a37a4235c
z7951a0972578f456c327fb3a2fcda7ea71735d539aab10a4bc35d396d8a8e54b83c3e2fb4fa6ce
zf07d6c061e8d002eff31840dc15abe636747d717d5701d15321ef7a236a5db88874449cea3f89a
z06cd59dd327646e94b4208477acac9d9216f8b34fd2a1d7d8417839c425b529890c1ece0bc8cf2
zb6b0b84decff28e7a97c8f67ae5510eaceb37c5e2acd60400b5e617b719d46a2a47de3591256cd
z93a78ff4d9cf9d42c84da73d2f22136a63d02e32ce68aa9935fbb8c9aae5dcc86cf3effc8a4b8a
z91cfdfda066fa84eced3603b883d2406e9e2cd6bdd12ec92426c04f293cdf9bd7cd407637e9bbd
z925a68e6955e9c8f3c726336815cee3e2d50659c80f1f87da46168110eb14eb2c1d3f3361d9d98
z2f08fac0ddd44d38a28f4652866b075bfacddba3a0c096c351d1815279faafe3d43a8de4babfef
zc4f317b8f8d44e301ffa8d860568360e6c338121ab53a534f7fb5c0a7e4f54269f8221129f81ee
z6c4fa86639660b268c75fcfaf9c90d2bba973181c81ec695b31cc670ee6fffde157b47c6cb5d69
zfd94ec7f974fdbd4fb279a04b3b7da280b3086957425ce2577f33a56956a364d88639b8dd64c70
zb1915cdb3a556fa84374144dc26186341677672418aa7bd58c1053d92c799013975726d0fcc317
z6c7d57244b1b7f4c05ac70a153be2396b0972537c09b6cbd7db957deb304f485a65ad1222664f4
zdb9c83d4ee5d9106769141d2760c08769cbdd029e1c574ebcbc79798a6ebf7d0e7ed57d8a64f91
zb41ee2eac1dc4bf3dd0df4d7fef0c2ba3fd84afd62e98714c2eb6a5f9e2c41a3070fa50f067f4b
z8b582e3bed82880820c144562c2f47055995b94121f60cfd63f66ed8ccf30276032a3a2c8ea9bd
z547c40f9795fde4d2dc9e35bfecae4d99f7505a61b1130675b34f1a27944b187bccc121ce6d03c
z2aee4c2fc4a8b6f9427410600a8ef0ac3038fd5a16cd5ff0c81a1ff6b18528ed7cadd8fa714b29
z2a35948cc1f7af0057346816f1c0e0f985488f6e12a4af222c838d938dce61f8b05351d906bc4d
ze612c17cdf8bdc3c13517035f981577eede7d2a9084735b586527506994ed5aab7d3d55e1d9b77
z08645f2938c6cf0b8f29e79272ed48996867b26aa4727eaaa6da17355883d4107e7b3961584eb7
zf117bbb0d038ba43fb2942c4aaa36f6de0d8d9df095715700e689e131f2e0c5e39635db64acb85
zd2f84b489de7bf84b4b6d7682d53ae7f017e66d44d0d8a4a7d1d61d20b5260477b4be4c7d57318
za0bc93b9f183f3a379079e62f24b0a4c440bb3e63525697a06ae6388b292f6b2c8e92373cabcec
zc40f3c35141000751b6732e46e5ab0b3bb9b553ec6753c546ba68ae6bda038dd5ad25f9b805413
z6f707bd667eefaa9861c590051189ccfd5b7e0e2a0474edaee684a7231138cddc8ef9e8429892d
z33f23e729be90ac76272746cf9918e739c64bec041321300186cce14dd0431dced5346f2b265cb
z28953b0b7fbb2caea26e72a7c372ba3f18db304f2f74d3a5adf58226cce86428136c14808a3ea4
z8628ef1f68f8274bbe2b2ffbb6905df1f5b951b5adeab9be6f3c2735faf83a037d1657908f21a8
z2da949224df0e840d938498894c593493c982b9105ba8cc9e5a425f93cc4a123ddd409027aa427
ze0661006e1532452a9c3d2948ae1f206c5e5c913e300e9b0c485d22b6e30ffe5f0b1c76470253f
z6ab17e859d23c83d9a5e77086c5a99f4eac41c691fa5b78645887ddb440aa957838638b6a440d9
z177a7fc64ad502c1749eaf5c176c0308bd669a428787765ca1e764fec33ccb157ca1654ad04756
zb27463f9d4683f5cf29cbece5fd5208d3e78311495e16976b1fb64dce9c91a21d0cbde905e865a
z6336a3fad5787272acce8659a4b02a3668ca94df8317e4e8f2d9b155aae9a2b40943a3f94523aa
z06e787391463fcf9a2e9bc8e86adeeae1a41f475f1c2c359730daaa6a78ba79775e5da033187a4
z1bb0ee1616ee5c474ab7eb97bfd4353027ca19da17930852a51ed65f6a6b3339fce24f18060cfd
z891da3228863dfc799524ea8224710390193d2df5d6451ec8b0494040279556c751bdb974b997f
z64b6ed85697570af2c3141db307bbe7078c3cfafc741a57782cb2b2fda1d2f76ef60fe72583b82
zbf29d29f732f42f982da618d4bf83f924628e06a9055cc3976f496ff029b058f281ad46bb54028
z6ff8025610fc833cf91ffe786480f3608a119b023edb93e7ee990957c17b91267dd58fcb58510e
z38e6f47eb2ea82ed6269f1756df522da4c75f3bd7bc62f1a698f8a1c55b2cf51c53c8da5732435
zddefde7cf2da527792406e2f2db541a4a94360f6c826764af277305279defe8bf1ca56954d8659
z0d578daa049866e94a0f5f4e73d945dd2070737a34c5b61bdf64aefa44d7150a554117599c4397
zfb72abd5ec2060c6ebb8bafb4c8469f770dfea09bbbb9c54ca812d1ecb245f0420b21771b2e9fe
z17d9b368378b8207f3f793935adb13ea4c1b2a91041481bbe15a37f01db0ce9651726ffb264f7f
zcfe2e20f58e19fe12ef1e495a8c2450694147d3838b9a2fc2ba017663187c5c4ffc7ddfe219251
z1f06162d93c1a2dd0c56c9848eec0f59121406e714cc9c9d7f291d1f983f7e4c056da92ff256bb
za1a4b5f43b5a87e2cac5ea86554b8f97d946c7f17ad935c10259810410c0c14d5aa74673cbf30c
z88f4304ecf75f15daa8707ab6c4db906fc03919fef46a0a244e4ace56ac29c8c3070e4869c4ad2
zcc51b49aede5835883227235ac6bbf4f5e9295b5133d8c7d83325de499f1bbe938620e7c62fe94
za955ed63565a77c7dead6cf176f343fe85211f7e3e6811f7189d30e45e4c78bb938e7d8eee44c6
za2fada91c5d1be3807fbca66e86ac9b2288ec0552602965650f0e5ce0b6b89bede8747f70b59f0
z583ba628e10871db7903296a33919ec1b099d31822e898a02cd59840195aecebf9019525cb2238
z7aa1fd0e4bb2ac733b6cd8ddcc778f4a9ff8a2c08ba9bdbb64b505a56e047f17c76e7224b557af
z204f3f2adfefd5e440e4536d0520e24a1548150f7e343aa518bdca51d6b26049bdbc9423c3b86a
zf59e4fa92f1f59fae36772594f6166f3593fca9fef0c3ec2fcac86c25d0299754cf20954a087f6
zdff0c1bf814b2c22c20267d28142158aa2f5305dcce02be7ea08feff485aa951fc5f961888108c
z551884ce2e9847aa9cd52a6a6f5a3953b0f8254f548a47a0869df0d5f1220007666089f50fa93f
zb74840462f90db3031abac3efd2c53a53b9dffb1fd8947b9d09f6d96aae5f82cdacdd4c45392cd
z7fbe7016b77b6bae8dd5589b9bbc17f3bf045dc20b6bcff1ca0e2d5d8202f6c9237d23a901be5a
z906369f208852f462eb0805e6d86599f11fdc3d41316bb4caa640fcb0e88ea083ca60b50328711
z074eb6816dd6d0463e5ddbb61ab509d7730c973758ccdc5d9970a0d3527abc71d8b209d3ac2e77
z7c682a62d5de50033c092d2911fc46a3e69f03d5fd3cf7b4c0efb5e3d7219cfc169892d3a790d2
z4d3eed28a5b621e8f7d918b35ce65f0832420c2ada386440e92d42472b26fdff366ff81f8f9bb5
zd46200e82522db9a8c71421100236754cc4f4bd88840927ed04340e9975b9a1b23d669ae7df99d
zc68adaadbb3049ec2e7a3a92991babc67cfc49564ba5a497abc70f908075c742648fb56e2909be
z59be98b3cedf60366ffa31a82db145237c5eeadd1c7151f3e663a8cc6fde321e35e44aedf2bd53
z3f2efc3762285104195489c1bd1eb1e924e65ecfae8d3a04e0ecb2cb92c6f35af9f5a570d3e215
z1fb95ba1b20dc3b31caa76fa5f8d942400f4d0e5d8a17d4ddbac3311dd05784862a822d26223f1
za5a1ce1b5e83eb7807e7d1f28671cf27bafd27590fc5bceab4c054e5a849217033526d90a7b870
zf6ebf284b2bbed10317af6e47c654e13a2e3d5724b9d627931d4ffaf4d97f3a52c97627aa9ac94
z1cbed79dd7681f16e4d206b6deb475afb1615e82e3f6d2b18f7bb2cd315a58e7a64668e9c961af
z9a3cc22e5600be7aef16603673d76327b026af018bc83acf51cfcc6269678aaaea2e0b6625b86f
z28dabfbb94e451c9e3e667dbbc314258964936490c8700d7aa8b9cba2023b5d65032dc50d72300
zfca7c27793cc8f06621c772be3b6969db7095e5e3e488abf1dcac66f1273548db69589233a671f
z58cddef6727bf0dd516f5368fcbbe0fb278e605c58a2cefe5eb921ab7d0d03ba64cb75ae0eea72
zde3fffe64c6dfe5c837748457f660368befdbb4fbfb294b66136b6da838b10327e0fe94692ca25
ze0c2c83641a226a5a1ee3e68efca657cfe4e4f92685eb30d41073aaa5e2d5b39fe8710ed1f6bf3
z26c217fe68ed1173d3ba0688bafcbbeebc82dbaf2dad153a576e98e156eed91969e87e12cb124c
z890d067b57a52df07a38748fb6c85438e1fe8d90a17600bad619ac3ec73e6352de893b91202e9a
z6eeb8e8984d692107c6da250c978676c6bbc5c252611ff5d6b028cbb82ba1cccc97049d6dd81bc
z12368df5374ad14fb44c127dd15389b5ccfeef1010c7a0b3e60c905a34fdd3aac75dc8c1c98a96
z1babc2c9015b602032ba5d658349ce0f40d9bd05d0315fd49fb8bc4c76a81ee2eed54bf266d6a7
z83c9ceeb7bc07fac4e4803780f498453f559c7e2bebc3f46c4fa4a7a2b63c832447fc636a36b03
z12b4801977c5efe8c155a04cb225e2c761a4d7f7f94bb91aaa06b346a3bc7ca01050adbf87784d
z653ccefa6634d8ba7680a8ea9b851dfe395d418d76ec109ea625a44dbb24583e36336838b4d1d0
z91620b085ea33630ed109a0fc22f133db2729859e2c9e6b3914ab55cff1045ad422707991ca399
z616807b31afe68845897d7273813be30d6e98bd2d29921a0c1720aafd5da65d7cb205d150ff7b8
z6d4ef9df703d58ee4eef16d270193bfe6cdaacf9230446b331b4f80bec16939367b3da93254f04
z67158c4915ea149e4799c4b1608a3252d767e3d14f555c312ab44eee0cab732401066b7330ef8e
z85daff644215f5c1d3efdb9d65d4fd9aecc4cc0d346436cbeb3b099fabb305357e8482e2b258d7
z3821e1d1af282a86efbf2da86fba11adb5706e44ae4bf0ca2da1275b141ce366bbe71feb72df8d
z2d5c239a162f49cb7a14a23f054982ad3294e4b37261ce9f3df120f748bc407d224b20bfb3fc36
z585ebefc5521a96ad1b8ab80602b5402c12dc8e5b29b996682e0a57e0be15c46f7a6de1d41c6e0
zc5ead16933fe81997f2d2af4f45707c74b31ec1e167acfe523ff0cfca9e0e8f6e71f14c3139df5
zc9eaaaa1e141b0cb6bd2cbdedb5c39f919cc61915e03aa01ae3f1780b8ba128948e1512b97fdd5
zcde871199e7a3c2347db4b7344813b2bf212f9f6d9d6798671bd5648020414a13b710c7716435a
zd716396268d4bbf1bc8b994fbcf265dc8ab4bac5d6e9286b311ed95f72345c8658c2411eb490e2
z98bd91a3a0074dd816b2551f3cc697f5d81cfb5b319962c341ff085869efd89f3f99a2844b3f53
zc864c84b89e900f94e55f4213f8c75ec2f48b290413dadfc7ce00700aa5bc2c869d2b0a555fb6f
zefbe05b8c99675ad9cf6bb727cf509b93c1a772925503b0b6064e1c23b2ed88c9990bd4b4a6d73
z1e2cf2dde51a4890478e35cea33c888d2ba50071ebbbcc16e87a7ad2d3683beadddfa41b2cfa03
z5538cecbaafd8a59b12e527da0e986c6b31cd6122f44813cea4bb145a5d3a7519aeccab0a862bb
z0bbbe2b5e55ad8b340d8040ad096b98b9d6c314e280526e50aa88137b86faf702437925458e6cb
z8574c4e4fa0580ad5d2c043879c9e88001dc38c735cef3b13fc54e8f7039c7495959629c2d2236
z7a33f4afa80ecd5e3f7f55e991219c482cdcbfef89e1bc30667ac770e13dcb9810e791c2353dc0
z9d66932e053524378e7af0df6604bf8fb893f8bd23c176d7cfc4114a713f87bc240c6d064ffd88
z8feb1693793b96d9baa5004581a751248683ab0db1d293854abe3399d4efc2d511d3b0bc69ec0b
z2af30c3bffd43506c190109d8b9203b7a6e7694604bccade69d9f0995d0282c58a79be89231e62
z1e108d15c03629e70032a86253d1ac50f75143c4b5d109f1c56c57d3e28def71726ce7d8888f66
zef7a1c43cc145df0df3e32202781cc0a3088b4cc67f8c7267c8b1235aff7aaed4eed5fd3eb37b1
z2964c6cfddee402ac35f668d2335b230338c8d3367ce0c6bd81e5686ca16f8536970c8c4985e62
z39f768d05ad82c5ecd0f2ebca1e495d6baaee85c95d70e964459efab93ebe23155708d010efa52
zde7f7d58c2d6e21fec830e9b98357d2b136997eecef47ab9e108455b6530e9a83f1cdd47de8e04
z480ed4191808d997935c137cc8b7ee31a4c93c9115cb92580313fdcf779316e3357eec4aaa9b53
z9000796a4e9e603ff4c5dcdfb843afd81858b865aded75ffd1a02ba722d6d2eafed30654844816
z6dcf8308e073f89759e910e567b0044164bbe12cb43bcc34c890750cfca208ef189808b165fef1
z4be683972bb3de35130a0fbd40d3f589cc2d306b322781deba2f1e369a35cbdd308baef29cf75e
zc38d7e82a27e2970fbe70b07a9b5bc0add68119dcf456b2486fef6ea42de1744b4cc67dca7ab7e
zd4d39d24238e9b357825c142486d0dbde1a0bf102adff653beaf3a3fa401c8deefa802b0aae2ec
zd1af1508b90570078d48ea037cafbb6c04a7357f21f6ad9cb782cae37a63da311160b53b346ef1
zfe6bd6b1e0dc241d396eb982dce7afaf3f4662ae0a2ba473048400725a7b7a5d7831845e856524
z6d86f8d5732594a2f757668aaea0aa8a85afa3b8130a245b981850ae24b2ae80737dfb99606b4d
z1355601293a8526e8c282f1d86e6a788900bed2fbf67eb263b10a3c26295b673d14380c60629be
zb7a4f5fe09d17b6af0bcf2d27f2433269bc93927851531d6b2c5956f928698ee012c3eeb1dab94
zbd443234f55e7f70edb54a3b1cf1dc3b56d1c44efc6a8fcae0fa2f7679113556cb668355a49c94
za1aa38783ae4a136c25169057cf5bac056245780ae0d85914617ce18e339a6e5e847581df73d1d
z4e100bb1eace177aba2aff355a9ad62e917c240c891d237bac77868ef52442b7537e17406ca9d6
zb00e281d9dfaa2402e3f8b96be2929aeff61ba693ece28e9f7c3eb75e3166785c57de31cae892e
zf6d5cd999caad50a56b75ef10a2a95e5d62aa3211d203c4aaf09dc68e895238729140ca9ee0990
z077a8590051cd90a84d506ce65a214d480666366ae367b23e17e270823bc67d064173145110a02
z9d6ba62debc6678212111276ada9e9baadf23a16eac186e9a46a25b6cb8557234d22b95001e20f
z7c0e8eb6b7f2a0396fe18b8f410f8c323374620a8853ab0fa3090e0f21ad2bcce80b0f441169c5
ze6bdccfda531c036fb018011f9a22a297c3eff7d736f5674105f3abb807d106e7aa673f6eb0b94
za5fdf3ba1d2856e28f46f0192803ae92d70595a0a26f1b0b67b3fd62100581760ea26a3333307b
ze477ba1685776c5f2da3bdb35f9c9de489b4c356de9f8dae1d59d41e99f1dc17af803baac2c8d4
z25c91c80bb1eb84571b1b1a0b316829ae668a47497106142c39d58441109fe4b6bf760a99d1b6e
zc7b9232d65d5e784c3508e68f122e187e95617e8b00812ef77c1f3d9111cae26dbe5622ece69d5
z6e1eedb2ccf3de9162967b5dee0dc20126f05a994e7849f73de3e7ecbac49fd8c9bf6db543871d
ze9eeeb642e2947e8f2ea144db620e8cdaef8848a6dfebab1d124743207d6ac0108e225fc452061
ze88d09bde41b6487abb55dc76841bd4bbb5cea07120d0b965e28275a3f51bf8643ed521f6dffaf
z726e9f83bc50341742d88a5abcf966e14f7ecafc3250d4dec5e69e9f4b383da86ef5236f7f5f1e
zc977f2f25aabca47163a0c3e19b67b67455a47d2c8f5531b02ecc120fe26eafd11e7f88d597266
z8d3d57c6b9afa298e96be55aec008447b31aa8556acd552c78544ce0195cd5c1f625c4f8f90f31
zad20c20dba63dd3b264f3dead76bb1dfe11338ab1fd17abbee9e778b747b9d87c93f00c0ed3956
z200e733edf798c3633f6a8facd67b3d4675dc29c66179399550cb8449f4b374bc4d09d2db33d7f
zb378f73cf3853f77afa1f195059afc95021686d7f772cb6904b1898f65aef05544500489e635ea
z597f1cb192b19e2712ea32534d8d75a6a216d61d26d8b0f0543b70546a91e84a7c4ceba6788fb3
z7b65cd650b6ed2aff82251beeda00bc2ef48c82574e1e06bd2f93caf5cdc8ef17a31e56bb71fc0
zb4a50aa9aa40842bbff854f7588932fb3aa520d6ce5089a668950bebfc495c43ccc813858f3003
zdca6c23c7d893743496c07b48352dc7392ec9ad05030da6fff268dec3afc533a0a6b6da0a50782
z65969a38e16e32a705f3e4becf1c1af2a547893ce73925005610ae1858394677ca6ab68405b798
z2d5c9b3fe042496ac282c3e868b37d4e8a615c218b168b41d14135d24cf5282bdceaa296b4eee2
z2cdd932eaf83651870ed55c5b2321bee0121321cf39ac146a68ffa091f263aa72527f4d6e7ca4f
z894b491ff08d2b7125303433a3e37d2ee6ef4bf428bc84cfbfe38d4d85cdeb2dda4252dffc89d6
zf35cad9a90620e9d46fab3b3ee05cbb7db10c62992b55bbbbcea328a466cba2a43ef726a5efa11
zcc54174cc648cdf7afc4f9a0da7466d8cbbba973015c74e27ae125ddae93d9f99bdb2c1cb697b0
zb47a99325da3d776f13232ab84abf5f248826d3b6cb89801cb07ce29198302d24a13a945d0d81b
zc438e038de4a7199728278c4a0223b267d049cfd687c7023f29eaf10a583d6660871501b5cb1ef
z34876e0d93ebc1997cbdd47bd3ceac88a0ce5ff4ee9ab603ab9c9542b492b1f8f0d62cdb205c82
za5944e33cc6b60fd074f58ca893d2805d681563c6b2c0ad5b18237ec390ce813e958a77d502af5
zb619197c8eb5f11111263893c02cd7235f70853eec1697963f9fc2745c8643421ad982a4c8174b
z1844799af2bc714460016bf521b8753595f51d8768451e9f14bf7ad910ffaf5bd20d7537a66a1e
z68bfd9e9def74aa70aaa6d9db1c5a2e82c4c7d388bfc610ee56ee3d94ef302bf023c604add53ae
za876873f0b776f84001c595dbc2f26b48257934bb782199779081c065b252833f2cbddb13be6d7
zfab9f9d2888d20bd59f2696cab8be876adb4ee78eb5ffaf79e903ec103bd7d2efb583ef1833bd0
z983d89af2060124477a0813efea5b42dbba94839db090d00848cc5839a4945f96fb08656ff60ce
z51d67a5d0f97de64c452928db1b93f5b9af60ba93d6dd5682ee20b73545e3fa4a1da9f5a29c9d3
z5d9f70527ac16ee5cf7af029a92f1c4ca2f4a68c9a62960f756e9d021608d6c50ab4fdba539bab
z576169d0fd67f61c389819f34358e297ad2815f31aa9f726e182e093068911aaf352c8af5a5f28
zdf64fc31a8d188eedfcbc4dd03a41f5597979ba01916a8758a3006355ff11cce5b6e25964059dc
z2e397dabe630ac06df13131838901712dadbd90b8fa569081b70fe7a4aa4785683a10a30ffe384
ze98b61e68b0e7f0631ef9eb27bc38a475503f8ed725c84fa7d7b317a89fcfaa84aed9c728b7cf1
z02ac6cf4b50cb5c6db4fb9b418648156b8d3645cf8b518b3eefd4f69961c84eb98da270960eaf8
z3c29e7a843889840ecbd3be3b11134bc4930ad738f9793f02c00e25f44ed505353751a3dc5d2c5
ze9bd2fb6795ac14deee3bd652dabaf9b530d2b8ca6fd9cd7672227aa3cce29642b82d2d07b16dc
zed4553191d299ae2fe75086d1b89938f97c448c3cf3d324eaca770b7ec845ea4238b19390ffca8
zf1cbbd99463d89a90ec7e237e97d7ea045ad1d04dd6ae57bbdbcbf28704b700bb52e2bbdf77557
zf6bc7509b57a8379b1ec8783a165e566270247cb144254fb52684660dd89f74e96dc845de1021f
zd7bd968d2514ac609a7224464bacd289ce4f157e791b8b6f62c479ba09f4c4996ab80451463e20
z38a576523a4d15b5c90e75988e075b8967a3fcd8823087c84317f1dfb697ef67928836264a5901
zcbf793063e31af9431217bf7f604c4d396e49c07f7ba44e214434757078927a7c4c29d39cf8d39
zd775d69dbb04d8b56f56b09e32de1cba9e12ef5679e39ac3ff199d4b90368a11c96fd4fe6d4e51
z6d38bb91559bd26102f5b170a6220229a62e3fee35781cb4776375ce339d04c5eed2a1627fbaca
z38936c967dc3751f069d49699515b2667b19a3ca0c324c7f613b514524e34da0bec35eee4dc82c
z76a270efed6f2a85128a46310135653b8eec10c60dd801752369869e0aaf950f3a4100c9d9bee4
zf468c128f8833ef0c0d8182cb5056a3368447a6314321378296b55b551ce1f8ca091270f7de961
z0ac036a4835869f3167163bf84e3e049d484441f5e845e9bdee118cc178ed0972663e8e15f2a45
zb03e5ef67f46ee4aa4468fdd6e5f96d78c47ba446216c998be4f485eec1c67bfbf0c2473ebc40e
zf1b370b869636013dc8a4ac9e45eb34f70fb1cc303650b8c386360dabc6c44ab8dee8d30def05f
z5a2dba4cc27c58f294356d183e01f8725bc4f60790e0586eaf2b948c699393dd96c8b0f36f0395
za75263972a4e020feaa0ccd33f237741ebe4976fd38957ebf9a704f9da224988eaa1ce522b7c06
z9e45e15870771006d0481620edb4f88ac30ac0078169348d0fce1dade8ebde4aaa613cae14c4ef
z5b1b2ef7bff7db0e871f632fe8e873dd8b930611606229421ad629a08fa617b9cfe487636fef6f
z039a7e86cb2a2fac71c948acbad7c6f2adec89d674e0cd75f9147d2fbabd84f9c2c75f4b2995c1
z2eb3d8b766997babbb608ad9e5baaabecb5f8bb2f10624bb82ce0a5da8b7c718e26e8680118f58
zc3ae9cb53cc28907044bd4245e782a51dea5ce897fe1895b5ffcad6038fd5cfb3d6c2ad0ccff19
z2ded3b3ac3fe8b72ebb6640374c1e8c991e89362a17715d2a1b9196504d41c623231760394f61b
z77ff8df54222a1b877452c2f5771ec9f03f744235507583e7fd2bfd2a21d3c6b96f89969b56881
z80b621ab11339f13d4601d852d747cf4dec98d23af9a8de3297b5da8913e6088289129bbe47c52
zbfa89779cb0a268a4e1bf91231d8548f021a4cf8fd333607d0d1a01ef2688065d24e15f2fa2b67
z1e35c4957fe388fb519b9669b7aa72dd61e83696bfdd65939fdb5679099b6bd94a7d36a95c7f0f
z7663ddbdb5b9bdff3029dd3d5ce7c6f01a713661378aec4a847ec47f8a99e646588352543fbedb
za0c89c857da34ecaecda6e1bf5c9da855887d984e4064504b132b0fecf4d29ddbdcd08909af82b
zbb049954187eaf78e2343624fc8946df15e3447d45b736567de8ebba60a88fbfca52cb97dfae51
zc41f4d15da5bb4e1c879c851ecb51f200f88a8bd4fe0699a5d739246af7ecaa2c99e0d67475400
zc810bfff2c5a1e96a57230f271adf48f90847de7e740d608c841a87f02e7f7439af43191c069f9
z40bb9939f5cd890cd3121891c0a56f831be88a1e0de1820774c96f82f3711d15bac1feec2dd66d
z1475dca1d516ffc435da57a795741be33074a60529756d889376eb534552481f845959f996262b
zf010f47d6517f58d3b8c528f86c35d78b2a22602e5dd69eb2cacf8716e4e4e186078773cab62cb
z0a0e0de9d8c2935d1a0c51fb5736f7068287dfa2f363ef2dba4d2ffad42f6aba3be3b6e7814c14
zd9bbb40cf7aee8a424a3b060d26a8d0c094666c5d825ca5be081cea751ef2f4d8e7009e53698c5
z14d8a7f64ba89c138c10883096dcb83656b2edb86c6cb7aedb4c5e94eff40f027094976ff86c8b
z29ba28e46055977202a6f0549202c676956239c19a60bf1d2fad43eb4ba3a421d5028a83875b7b
zf067a4ddcddc6d2ecfe9bf320305329ff6c37eefc5f01e01ca814a32566c04a4c02e11afc633d3
z839a07108cc22b9af7c9af5a763cb05d732a5aa46eed5e407232cf3cff8d453fe70243347f0a82
z395dd391537272f5bd6358f7ebb82b7fc20e8745789eef1f26b439110472a015eff147b6c57948
ze135717e67ab4697c949a727ce63b5b3893f8e36d17dcf2b10f79aff5fdde2e50f1b955c0a0e7f
z50da32439db3b7d750ad5d53bbe13613dd26b9cb26518066f156f103cdb7b03236a6373133f80f
z6f50b4bb816558223498faf428d8b890cec1ef0cea3b2daf685534698e010fa74650d792c0563d
z3e385397d61829a60011d857208819ba7b744be1c5c4b771d25e80826760e42e2db4e1de251578
z2e1558e693147e4cfcd5d007383883df0bc54551bebce21cbf43a41dcbd8a806e5247bc8e09aee
z22f3f6519a0a34ae23428fbde27409b292400545b5c9a74bc97741b653afbd832097a65d66153c
z612000f58d4eafcfcc009c39b4fe2d7d6b36ae65db0282eed0fea1092787f0bd4cd85a9c93d662
z431b858e058e95b35c6d46b97709b837a8c15c8a1aa9e34d99832826647df54894690e107aea09
za867fb1ad4407e1ff059492676c7d8f558f5ed05730425e67340479c6c7e860fb2d3c4deb8998a
z30fa6b032a3af9fb4b3b941e87c6ff7512898e6625659664f97a514ca30b4e8bfa35be1df5f30f
z009fb807d46e3cf81703769c8a4e08bbe0f9ec61197a9ecb873c790bce37b81e900a39f822d666
z4b8bb1c883f73295e06bbbbffdd6f0482ed1711771ed0b3f7cccbd1d16670b16a3dbabdfe2c061
ze6233cb9735138eb568c8222b94717d0a397a7a12eed544be84140ccb0149b5d10e56f15f9ffa3
z8587b43f5278b19644054b5a67eca369d94b1282d84e26b7c99680c0c6500a5259abb82c1fe2a0
zbb355ae213655bc58a7f9c40a50fff13a44d13bd8974f7a00f7786163e47b37e53412448127765
z9697b00e34c768cab55fb61ab44988854b2d3a14a65c6f735170766fbe60a974b150d135cf071f
z34c1cf1b99345939cbb2bc4164270e13514f416f57b8ce53e5a6016911880435f33291fff87bff
z47c4a5e238392416a91e6bf307384d0736bee126e7c5b325e5779cf5dc2f19afee000a17bb46bc
z9a21a1d1aecb7b79db84c90d938b2077c4fa25cd006a171a750f6a45125fecfcb98182017c772e
ze44c9f80afa4c7fd667bcbb21790421b3005525dca37cf2e3914bcc645f219c13b94f51fcca4eb
zee131e0ff22043ea30a06ceda219c6a719bd609481a761e120b23aba083867925bcc93a24d752d
zd06602371f696251f3eee3358328d3de357ac8f6fc2edb2868f6cbe01ac352bd6dfb273390e277
zb8148f20a613c378092c86f904ecb2688828c57c3c3d0756a308841277646d9856b75a285f209c
z7ef9e8851039abc39a4e0845a12aa329ba6de49ff5dc45eebab61a3a90c8f947dd9bf9d3973aba
zff619b11f7fb970e004bdcea38b13cf325cd0203fcef4f06bf3d0c16d899a45e0c968099a44069
z63f2b977ee3e43e08bbdad8df3aca61b35b272be069c4d6086530be4c0b241f3047d532df2446d
z9d5533eca6f1601d2544a3bebd26ccacf30228f1c3711ff46f298b76585e0e12e0b016dcd7cbb5
z3f5c0bcff841d83e7e5e947d818c0e8bf02fd6c7b1f46ce1ffbc2b989f4e2fa308f648d54d586e
z153a86e67dff5c280418767640853f452271d8bdd54864ccdccd75717e64319350227cfab49725
z0767bec2b75f43be8bcb1ba45259da52d1e60e8a06e489d62f001e370ff2421fff0a9e4e9cbeea
zec4e7250e5d8c5fbd647143acd691e5694debade4f37ddbd753dcdf0f31959010c29c1957aefe8
z20d973254e737fd76053cb591cc29138b97244126e99461cba714d95c6575ccebf340a916d48f2
za7bdc0147b756b4272e3457853e9cbe3c414a37b8287e1a9c266a24b0fb3aee855de3843ebdc4e
z6c94b29b45a82f7d78700e9d1fd1c2d5f8b183e8294f9afba990e40bd2153b71bc6cd4ddf8c69f
z797bd765241525b6f10c05943806c2296f8ef2614f257b5ee90dd78b9c4fbcadd7a15d9d034948
z521e05b5650a1b41ebd4da204470cf4156cd1ddfef48bb7c0c70d7dd8284f85a160d31b99dc5d4
zaf85a8b73c2a1fac8318b146fc2d51952c73ebd470da4e83ab1f75fb92843fbc724570cd9119ce
z81ad6d1b0bcd02c599b916a2323f78e284445c42edbd2d9c73d4b0cef921de3d50de1a534c5d9e
z9eaaddd13dce5dbf0b4f0f4c2075851ff2aa7a1bdc873fbf13cfd0a215fd2141fcef4d06f49644
za95018a585b1c659fc3f4d88da2598b152438330d9bb4ffff5c81ffea6d722e7710596623cb6aa
z6a980eb6941acae43829f4ba218757c6615690187172d7a7de15370f5daafa525be9508d5c5607
zde0bd352a4a5082edc3f156867ca6cd8cac9c0f9b40b6b69007769f31222339da2cfa87ee44634
z3a35e31886524420e0385b992d3ade5803f2ccf33c9508e9d23a5aae7a8860eee24c96e68b0f81
zf6969414f91f7edbc447b09113146f09badaf25213de04953d31dc91a4bb53e62c60c5c5b2f71f
zef6567160a7dae01f7c17045889e7ad4bb3b5d3facdffdcbd670957b936749a6530c09be0008a2
z3b1fb1820892891ca5335ba53d66b1bc93cff7f8c7e070f23ababd439b7dc748b839ba4f1905f9
z257971357f60cc8cc278e0d3bd507717c0da012b37c61daf24b43968185d508249595693a65804
z9edd30ccb5fa8305bd9a69f98d831d0bda7acc0f14d636dae51189b197ebc677a36fac8d111a5e
z7dc8fb5bb44385c57500ce555e14fbbb819bb440ec7b45abea5ebc09500335b621715671126e3a
zaa93d4fe99b3ca9bd0df4a21ac8ed0f334846951e4c35de715987ca723975b69a0c6ced1adc784
z3e0092679a4e93cb6acd37d9c72da25594a03acdf2709ed2b95a89aa7b033e29708daed8a91a58
zb7c7ea5eeb97c037edbbc2ed39b3de83e772e95dd6761d0e56fd8ab4be530dd26ebd9fb6124415
zf350ee1080c78f1da977853279ad8cd69abcdc781a3db262e7c15327f5c45643b2e0fddd2651e6
z7bd5aaa71d110cbb7a72ef488acbfa42517df036e52af1461bad3f9ccf70a8f2ece17ddeb9667a
z74d3c6f973c705c82ae484982d9473ea5e8096c6c521016e6462a2e3d9ad446dd923bc688f441e
z4b457c28d4e0ab223683ad94073e3079e3fc020befef3fc2a0773a8ddd7627d5b0429f5f1e0233
z5e5d08776e81ff8d785c40dbb8c4aa8aa2150c16f5210e4d06951db74314b776952e09fb4af8fb
zae133b46032f4541db7cc6d9c13b003e489ab54158424d64daf0fbbbf6c12e3b5c8106caebebac
z07fa8475a7f3daa1ae6666c1caf2a28e
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_assert_timer_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
