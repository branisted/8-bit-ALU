`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab30857016fc53a
za25afc8341302f0c829d94450c399b8ff9b0386c187cb854ee330605b7b59da379b1f26f488e1d
z36e675f0b1336408b3a1ad87d0723054f952fbefc8d5a33eaca6ef5be8f42bc59870a29a5cc9dd
z4fec09ce6e44cac279651402e7e1f590df88ce49ec26ab39f12b4a02855703c6f03b1e85c797d7
za357087d98e5b1f45502e45892e5823d6fa4b762932009620038c05d74efcea7c3fdb38901d620
z36515d0824367e48d1bc182335f158c262d396cada6b0ad58add4f945eee634c2dceadbfb5118e
z14969c29a743830a07124bfa78707f3952b96b0db7af7c9ff36f77137d8c490c4f79328328069e
zd7d5280e4f95742c9841340368b9764f0f80413adb175ecfbdf3c40716abca7b8cef6f7fe92ab9
z6bd2453f1aef7f7899c5365c5c83793cacc7795c269413f6cf0dabad14d40e9285afde8c01a47e
zb61893788ec5060288cabde8fb553f21b02eac61ab0b48ad3d54f4d1d76508b22f0c600861b5ce
zcb30ba708be817b1f50f59c0f6fce449203e7355c1be55b662fef3f92ba58243d81537761af8d6
ze27d7864d2dae99372b2b75bacdc0437a4f7e011d68c3487a89759e3625548fcc920ad06471ee7
z2d701aabf726859343208b0a543c73eeff8406febf277e3babff437ec820fb49d6b78e73bc2353
z884917487d35a6cd06d7d73ccff5f0292fb3df6f439aded7c8bc5dd0187f22a0fe1ead93318eb8
z8c6e90111edd2a748769a8d92e19030b0323140a1ef01d3a257fd16256b12b03810bb4a4e82398
z2704088d587398546935b6339280ed10cfe93a3a5b7a4f04e0a6f073f8fa718c2f9190d76f588f
ze9fdbb73c2c6c983be7680e758043939fdd6803162983f37193ecbd51d83a9df901bce5c960f7a
z91451ccc98f8cc68bcf6283cc3f9b8b51e819fc5551032ae29e144349e39be15f73760385f3b1e
zaa10d4c3c0da4b4b70a060755265bd43e18429556c824ff54bffceda07d93c93c945db5c21a789
ze8fbf98db4407fca8f361df1bfb254cd88cbcd56aecfc6fee807db8ad4a60f00d9f7ff17bff2c0
z77cb078b0154ee4577dd19692c01efbde3d7d63a11612f14e22938bd85f072db23bda55ccd466c
z5f40b0cff9c918d188bcd82bf8459bf9b373e72076bc38a2276ebaaa6151f611eb8412f55b9c98
zca31719ad32a0c5a52d9e787fd2bf3671a94f7bf22c26d3d8bea2df43bc9a30692762ff5e4f86a
z46f932edf61b09ac566aa5153f08bc292ffa186350c922714c3749f6f013aa9c955bbc875ab1a9
zc035d4e9336398732c02641cc754b8a201d54037f9b9a7a3fd4dd13f25055c83b0b2656901a3ef
z9218e764103ea255202b3902739a39bc67ef37fa204fb6c5f3ecbbe2b6e32048689e161a1e664d
z4d47b582fc6332933b23df52aa948081988bab1100d1974c647539c0bf6085d54d1dabedf9293a
zb51b9e5b9a56d6969046e39b914062276737536b01fef8006cc46c69967adaf6e8164f4f02a813
z287834e7ab9d12606be2a713b5860a18c7d3f8fc8658f8c62ab3cb0958a2a3c2db968bc9fed218
z44894a1d1fd303a5228b02470d2a84e6e8cfbc771120dc1a297e9c87c5f6d366e1664611e993ac
z187ad5cef57c4608ec9b6118a8218fd5acaae7e56d69acde7514a2f7a2fae5beca37611dc4cd10
z17ad6a7a37af3f74688442fe08d9683c64cb0e069ce137bc0f201b25c404a78d78a7ec45d6f453
za20f1d97b85a7e9e37266264509a3338fcabae693f12c0a8830331a75a0e23a84e438b5540693b
zca24086ef3ede7aaefedc073c8a94aca5bc514a458155de7a658458ce36b0cad615b11e1c85468
z562bedd7d747bdf75e5940b1ea62fc45f124b89c31ef26617befebac676d700db98939d2d29c95
z2fb48fd60374e4a445983294020789768f8967df867c175d930f477ea2fc7ad77253a465d307b3
z79a12ecebf998bb59f96c22c8a2ac5b89ffacf282949bd9fb8ee8c0028a2462b0edf4fbe951839
z8f82fd3c4a3227c0d2ffea519dad1a291b696836bbccdb6e3c41963d249252a50dc5fa2b9f433d
z70cc634b328cfd989d2baddd66c542adb795df7d35c436a05e3bb99e1f28c4b74740d6dcdcd374
ze5435cbef3f414e9129c52830e88d804d7a28559da5423dba4acf8d1098a5898fa9b60ad9d99e0
zc8324b1c3b431cce8ec600cbb62393de187f5a7b63b0341c6eb6bcc8e8fd2879cd27047bf410c6
z336b37c4f8ff8cbfd8767be3aede3e38e76c5e4ce80733e92bd72b1957cce41fda0c881d722c0b
z1394f0f4002706bedd40addfe2d90e696a02ba4e57d77beb0fba05df08d85305c076e9e5f891cd
z5773b5afd973a65cd20a321954dc90e6c697000f58feb83ed20d02e083aa57154a2b253d807511
zfb984f7f5f05c9b6a5cd8ead9fc3ac4ce35b9fb26d7b2086a4e5bb4736fd993a12d10c122601aa
z2bfa4d26ac7b64c0951b5cf83657467c06df377709f2d4719fdcf104f67432bff4f6ae512f1495
ze36251b187fe10da1558a96549cb0f0a5cba90f80ae75623feb41ded8c7271c55dc40355ee2d46
ze97e118e390bde24e986aa78f8ca21276f1897e931f46d8c6c4ed5baf7bf883db5d76eed0cc97f
z987ae9091ab3c4d416f7d361aef913ac3dfc38805416fdd8bde4479d0fba3cb45fd366ebfed923
z2ebcb2d6ae0d089b871a9cc3ce8fa51dcab47f15c7048e2dda3e010fbc20bd602add62528e6e19
z4902e589d2debce4d5967be7a188dc299010f9aa67a7bc1dda94676bcd962e47863d0105ad54b4
z6680d454c6bd8277f29530b2fb7f924c89824ac426ad99627a41360e5e4d22f7d56038d7a0aeeb
zffd710cb120effcbe361c634d494070f64bcc9c62746d7cb1928885bef35e7e0ecb5d70afc8cf7
z10b255d88e21e9ebcd83f07d960ea524ff6ff7c11165cb324113b4b15c1bd95e57ac5af8fe88dc
zdfb2423a712aee1e33714361599ce645a735e1778b6c5227f6f5e007e038afe153257bb8342cce
z5e21684191da3e46d90e94732b9bfd15e31c5b7219eeed88c5f93085aa2e5b134d493ed66f563b
z36f7c589618e538d47c6a2282e9b6e474ded3dff3b34fcc5520c4aabeb85660fdfc5f89584cf37
z943aefcd0da64cdaa338988155d70dbd0336df30a468cdfc608a3aa081c3853ac4d87ba12dc69e
z9150cca61818a164159f08fcbb79c6e828a72b60733e798cdccbcac3b18ef728a617154d45a9f7
zf350b37ae9742079f66bd87927b0a8775cbb296ac96ec27b279e81692544ed45b44fecbae5888a
z873d9b6ded06cd11ff04a328fe7d1b9a0e45439a1eb95a586592cc96318365690bd3012dbce20d
z6990ab452b5f9701a1b1603f8d1d66dfc0be9e1d7ab7e4211984ee707ff4f11f825627d3ce40f7
z92d2a647a1dad854c8b47985e57240c408528910889ecc79d5ce1862df69c336c17660bbda3a0e
zfe9cdde8acb1852313c1f55921957ece0645bd6abb6398bb080f51af0d4b6017f2e743763d9d44
zab7f4bc14a5c330882fb4d12b7e9f7e105fdcab587106212c0e8778059e7729ea31970b78eba73
za62ef7d375db2e697350b7cc0d4888cdc1919afc73859798d5e3142a5bdbf2a90543507b63ccb9
z46b823a4869c6f4facaaa7ca5cfb959cc48909920ba3156df02a1cedb6db7ff9817267723cdc41
zc563d9aac441c4d8452fa40cfdfd2a1b149abf62181c4b14532a135fe236d071aa2fed2b200ed1
z0c095c58a436c57ed8aa6c72205d47bc5fce12c9b3672ecc41404150d17e689ff813ad6bd710b6
z91cb4e02e16e2aab92c73ea0f070b7e01edc0cb6a2736047007bdb9a98373d88348b4a2d168356
z68a91e6e1d8b0472d79800c2989d2f7a97abde011c2d6fc9812c940aa957cb946f1b3f6e792c95
z2c630759af1288e1cd4d40a24763b3acce1396a8a440ce2a9cf1e7aaef04c2ec36ab3ab7cefe6d
zbe7a65bf921f252b7bcde655b257fbaed607c633c064595be7deb27bd179a56e50e9602ec3df10
z05f6fd0629eddb1ad7039b33e49516198de90bbadbc540e4169ae23533023fb6ab3b05e968c90c
z2ea9ad168317c8b3314b0acad0bc02d7fb77e9ea7f97d7c17120142240b98355c61cfe45b5d545
z3f3617da1aed13e5f5d4e766406781e757b7566b37cce5baeaabf2502ce97f655a1633d7c061c8
z02aa38e3325b356c9cd8666fd69b8f5c8f3cab815be2cffe336135359b1c0ae2772d573b3d37a6
z49a73b0c184e7674d0d2e7f693e27f7be8236593f79030ac9aaf5d45f4ccdfc2f1ba54764b992d
za09b38cde0525db7c5a633f4f4ef0836a3ed1e0dbd0099bf53db35fc0a7c206560437f12545651
z3f68badf1d4ef90c85c8b8eb1c11cc9ecf079ff09d1edc8161c0c3f98c4ea6bc12a7f3611e3f1f
z97dafbd842c90e2ef3f845224a61ee90f6581af0c25363bc074c8616ad239d2d5dcf98b05fed24
z31083b9ce6048627a9abbb4f59e3bdacebaa1a566246961e00eb738d9a7f26050a8ff96b39c7e8
z78f09c6c255010fc00734f9e20dc853f2c0fa7af024ba66bfef1f6dfa62fcb1ca80145c3391662
zac3dfc373ad8a7a96e6f25ac173d7af7ff6fc8ffb9717f60963dabf50b039d2f8564cf63b2fc28
z9f7391ba97f2b14dbf91c051d4dad9e2fd0bb6ab5ec0dccc0db8f314218bfb5ae18cf107fd017f
z1412eddd43de9a53ad31bd75d606df809a4b8c748b79afcf1af135bc3d69ac7007562d8c44e77d
z7c47421596bf7fa981712a5fda9e6acc9d61ee1b2dd27e6f526cbc1c20c6631ea4847a37b5b075
z02b7df4c4a1bd06e8200ef31d8bce3d304442c1e09d1db657de9afd79c402be555551afbd71cbe
z82a3524f23efdaf8e6f30c52c7a5e01d0eed23d08eb60783ba12090733d39ee42291e3afb8cc5c
z60850e5c93b7da559c20236bddf7ac75b02c57375e34089fe26b8ac1c1afb102187e3cf4f6bd8e
z7c976edc4f52955e00f4ab72acea95e8bad0502c6002db1baa583efdea46553fc04b65324a352b
z95feb1f9b5003a433740ed34bb99a79eeaeb95569772f82461a60e86010a45f59aa1cf4f601745
za985849b2cd609207dc6bb7b07500c547b57708e39039c8fd206964722b7de5545ef2e05bf51e6
z7139a193f7a1deb0f79788d7791674c733528c0d7a8b9e8013c3ec9a51d882997fa10950223a81
z0d0b275821a03bffea67d45e55e41979c1272c4b6c954f9eb0e9fc90a3a6eccbfe9dd6c6b5fffe
z9a42e06f82bfa0947b1df958e5925314d5d2f32b66619c2c2ca9c992781b4e43240fe9ef561cb7
z06ea22862635530fa7cac0fa7e3d11dc09269676fbdfa463d5accae7ae810f172076033904c041
z1260c393f69b2753cdc75d73fb5c901b39eeb00d2985bedd12580bdaf4be3a3c1b005612e90076
z13321f7eb92f4a88707a83c010158084be2512eafd217feec60f700de62d71332c2eba97ef6420
z89b0314ed71c82698d0d490dab09bba52c7cfc8c445997abe25a284aeeaacf328e6ea13018b558
z0912c04acf7247a92a959e6b3f60982a1ddf6d1745862d6cf73fc222ae766b34898d9c0c0ac1fc
z0ad99cc4975db45dcd708bb3705e2d7de5eea1e969ae42e34b84a59490961d190b851958dee3cc
z321f0d200c5584a47e991ec6855bf9a8e635d25152e8fa6bdb87aa68aaa29bc885f580f40b7f9e
z8aeea498dff735818cfe82c0d46418d662c6636e8ea8932be52482bccc270f7561570feefab731
za271283e558de8c3f6194f90e0110c53fe5b559f569b8e5895c88a2808c838245f237ae07c9c75
zfeed2b43f0209ee945cf2e0a9c4811d8ebfab7bbf004ff8546e28a581cd851ed7239e49ea78ed2
z316835b95be41ecd22fe21925f180460b31ae67652a561412363bed87c08ebebf7c4328b654051
z519c989a6285c23818e18fc78f146d6228cd54997f514c37805232e647687e74a422b2ff491cf3
zb4a62a7d16f8d02924c2cb19fdc2b0d095caca0d2cbed03cb9b3bd96c760ffa97ea6eee4259f35
zac15554a6f5fb4741a7c1a2d32ec54d47797fa0ed7e6ede591bdbc619d064c6a57ba993a214360
zc7249abe18cb5b5ce8f6ac2699962f13665e48cc3504d8cab586ec796c53b2f3c99b10181d31df
z6246b47fcf7d6c0d9d55748fd7c346204b0fdcc6b99b2d2c75f33fcb1da18587c79624acc65246
z43546740c3748eff8d65a5a727fd049a79e7e367f63283e526ce4ff257ff4353ef8f53de0c1fa8
z879bcd2b799b6cdc0fa789ec52ea3a1fc18e91b607a58ab40a1e394dab4fa373f04c4f45b703b4
z87ae85bf72962d587e209a4a0d319f634f07d4fc529dedb3f42aa7419848dd6fc093eec016e09f
z3dfd6be26b4cd78d9f614abc15b990faef90ee02e3fbce8c6de28ab063374f360fd799934b1294
zc612861c437ee3d9569111aaca742af7ccd20d9b9a1e762acaa14dbeea8a426f187ba1821f15ae
zf7c3f64beeda4b63ae5206d3c0fc7a5ee0336b280c6250b7e280010854c550571b25731d086903
z3970bccd6b82bbf0b20cf99642120e3fe1b03c1dda92305a50a9b590c31785e62b46c80ee3b045
z40d21e74419c1384d8cfc54038c931a4703e77f7cbfdc4c714346b70cc1bfb25c64071368bc34b
z63f7a689cfa7c9a8e7c600c9934d52c940f68132b6bb4bb698ac9bd1435d7530231fd73c969335
z283243080e361258684eba9fd37bd4587b8d112778cfcb8fc312ab7c54be1320b39a25811c97e8
z7a3c83d2f3a344f55d0195ad4747d47ef03a831aa9755c7f9833be17b52edf30ef2d44a5401f81
zf25930948166f07105cad354da4a70db4d251404c06792a70a7469e62455c5343e4537eb807377
z8eac972b22b752fa44243207aa733994f20b13e7635d0d46572759b6735bcd70c4877770044ae9
ze82921c259de6e798a3fb7a95b4988a658dbe2596a6f3d5c1cf669653d1fb8015322e634bc7d97
z087706e40e8f94861803eadf88caf3a5e23321058b92bd5f6968efb753be7380b7afb43cd0641b
zb117076e82ffc3e77232364a1e79d1cfc7b40b9862731ac66a2a5f90dca725bb681f3e92f52765
za88e8fc93ffb9f81c4349221c1bb7d4222971a07f1cc6e7e0a2c0dcc4264c13bc94f5f59e8ac6e
z4c99a6dca0d6caab4abf629a19e89e95f345cf018b3f330fc4820bce202d0a5dcf2fda1e2f2d4a
zdf73c4ef7ab39336b93512f01abcad1a68331924414b2caabb6e41fbc240eff088b06bef4f3961
z674feeb567b2a8509e91117f295a4e0918d6e91ae6515caeab3af8a0fb722e0099f57131dd4430
z8bf410517b8f6641e19d44d73dbd5a927165eba86496172fbd13940a2b487cdd00a6b8cc87088f
z142baaacfc0b3432af742a203d320fc55966e7a8a1794a74a5c67434dbb222d50712db28f7a05b
z9ce969ab5d3c907b615e71dbde1143d2e230c4675ee4bed1659445b9003f4098fc8ba99dffece1
ze7e3ae475db6dd550256a6fa753bb1c4a5ed84b656ae87d49d64750cd29170883805cdc56fbafc
z9990d822ff6394ed5c2af08edc1fa41b270f1afb86fab5932de4f11a59f2e88aeb8b96aff6b958
z92b465eee99009c86ce1b16d673d0e2f0d5549a54071b46999ca42520d25067b0f489b7d94b6e7
z333d637bfcd52272d8af3faffcd4f220a8d28d0a2c583c88f9bc66213c3f9e31a4870437331047
z5aa6660aeabdd9fd54afb4c966f3a0ddfdca9e7a82b1e08d1303c55cfcaf8e89af16e977c4c828
z0cf69adb586823c81ce4567eca649956163d4d0b6493f184bdfc71d6f400c87fae58a0d05bc51f
z7ae3cd7dc66dee438a2c9f009b1099c5a3bfdadacc98ab153986ff51a71f9a69e43bef6477ea6c
z27974030cccb86556fd568d52c2af93a2f02469b2898735f2a7ca20eb4673c4046c0aae652f530
z7a268bede0eda638151e964c09a4dd295134ffabce433a9cced0ab5ce517ebf91074a4879dace4
z9de913a60a4dcaa43c2f1a20e6db9e8c0529a7f6fc7e6348be7c9175157409ff48e0ac9ebcd8c3
z640343515cb56cd7060193e1a60d0be896cb19931872ce2b1260df23c201d94b3f3fbbf16fd5ef
z908b1b6684a8a3b0f7264edd9dd5aa41e9629b640225e5179c8bc9474c575803e55232354f8d3a
zdb8072d37fd1f7ffd085deff9da027ea2277959cf8c1c500b1f45fd61a26acee19d5ff95be5b18
zd154d80a7ab3acd4b1a74a7698c850dcba0cb464bc657f2aaf76d4fa5bb7e61f7cffd3e4bcc788
z895ebe7839708bf563405efda2d09bea790aaf924c8de9d0591c809ee475da88c5b34134187d17
z036fc41306ffefbf3a22af3b6544a59d4bed4d2b0f72854478b4bd4ed13ae108324b7717f9b81c
z63064df38bf76818d882169f2e98f5e9484ca1bc633aaf3e7c444d70afb35356c17e0607fc9efc
z69a38276e238501070d55e7c38434e023d4e72a23a210ea8d5c73a40a158ec068de463a09241ed
z5ddcb74604bee78c5ae2c33216afffefae8a0495c26ec18914093f2029794b41dc5a6d21904eb8
zfb924ccfc4e7a0182a45a781e71d7661801e3b28b63fbb8db30e6af6b370800fd392dd417c5b38
z26d3f908dcb579d913deb6599a98319a68ee78ad14ef2bc763374cc7165470c012ea2d38294343
ze9935ace627a6ff430f9ba4aabcf730497d8d591f5d11493bb1da46fd20819b4bf8d906f85601f
z05228ab1684b8676329acbf2d98c14e70ff84746f966e9e139649eaf134df5f2f48edcf6632a15
z7f26f6e44d70658928b4c27938f64b765e42d56ac8609c2c308514c4ae546196b925439d8da147
z5faf3dbc18916010fbc2946e1dca08f4d7be086fd4ba2becdffe5f5a36902f5ac3a8599246425a
z2e9998346f5dfe0dd1412749e373b0065e2905b68281b9a0043fa69a30d0c2b52df899efdb537f
z2d94a812d7f9a152ebb7a2dd9f7b771ccff61405252aa5878f2e3f9b10c5fa3d412652d68ecef6
z5ab071ac0d2cc13043bb866f5fd688a0e5815c6382953c886f8677731b4f4e5e7895688656a6d2
z456479f8335e7a41e9785bc9497216503cff95ba9f734d25f57608589742da05770ae592495e43
z62539ee81f23003f9a625b34bc1317858cf5c7dc384ad1ba2ca1d40264a5a724d273431947b962
zd0bd146456d01eec145b27721d3df8b0671dabf74d0f766feff3cc2420faaa35221fb77f20a5fe
zc07d68994f3c82329dd96d57fe63b43b9a7f50f7ee66d95fc41da0da670c76dcadd0c1865b75c5
z5f9f12036262749b7ece6b2ef2af5317a0b0a5191760f2ca356286f50fab0a56ef0f0d98027998
z3c2daf2b92c7334651f8e2b80d150167a06cf1c9c33685ed6b27588f6b4e21f0ed06457041ad4a
ze645f92d5d74624039fd694453182b1e142376e438cde21a6a5d5249f9bcd6d9c71ba3b7faea03
z32c48bbb5039f0b8cae6cc0e885244d0b1250c813a94c6e5770c26edc85ae3885b7ddb36369a59
z5626bc3e0f0c8e22d8dae071f64211f0251a2403edae4ccfd15dd94c60b8d86ae56670aba5deae
zbb836eb3196162bd29c7996594939a677efb6078c22d03f068a6cc2a2f3a9c9f070d596dcd3a89
zdf448c78d7c77e4ba78b4489bc6c290feb4626b2dbb1e3ae9d61d822dd66b69a8e1d8fc196b962
zd2df2d42e73d37743aac59988e240dacad89e3d07ab887018ae642cfee82deb6bfa5245a23a560
z700256d55620bde4c1d56d0f0a838a8063cdb66235318ee3af9a26dc7dbea4caceefd19f22e3a1
z6c6afbacaf54db3cb8c9b4a05fa19c700f56805d7f9176ff3a7d9235401a7bb56c02620b15b508
z6a101de16b4f701638c7f37e3654872ceaaf01479c794f23f1b1ec92de4be0265c5ae6e404c169
zbe7d6ae1ec953623c178f358d9665353e4d90f821df827c01420417a1cfefaa6935cca1f638731
z1aae71a0757920b5baace40bd82a23b10b4d5992fd590565f3845dfdc76f0164168c8615af46a2
z0d33208f7d38176a25448a7fd3175cc84f7d908c047f871082d7c4aa530204c8645d2502ca1271
z5cde06e11b1b1fed9285893dba98a728243ace43e0a2e7fa12cb92f13909f31da2b5558f753434
z68de58b1be64dbbfd74bd1a0fb5ce70fdbfb9c89b10152d2e32190f4bd0c63363bdd09213ad5bc
zb2382bef420852c1ef058124b3e9aca7ecea1ffe4704873ecb237d12dd9b7231ec0df781d2bdaa
z5206e4d1926d83b9b02b5b9fda450bfc64cc5504e749dc423725850b3533f151400120d04d732d
z56efe884d1d9a1eb3d3c4dd304652eaf7bbf1f8d60e5cedd15bb91579c3a7103f15c74db3608a9
z3e39861d688d28d307fe345a1d341d98be622a752b87d7a0e52d35948af7022a3ce2451c5087ae
z2d3ec1115a88c3b9673a4d6597a6c052dc15d53a0d3838bdb6e18d5a66efa0865fd507b3dbfa5e
za820e6fdaef219564940fde5e77af896f6c423fa02f461e8c9546b77c1e29f674011792192a79e
zd1049babd43e143f2338c5cf105c79f424edbb0a24e88368e8726d91b8f9baee456ea8f48d10d9
zdf263c805825f81327516476a89c44430f4a3356a6067404655001a58a9aa72e7a2159e22359f3
z7d1d52487b4b2bd34e9a8d1ececbf6e0d8ddce8fdb45e5c525fc1a15b740144fa0e8a43b156404
zd0f450af62df2df2201ad60e815c2097984afdb540becba7bf6a57b0359c2d76194be58dcf6250
z233ca56ed6ce9ec8bc90705d5938e3d30bb27164286d4279ceac6429d54f9b028b192960bdff0b
zf10b1edcf372a3dc772d60ac1207c76854e74496d072cbd8008cf3fdd27bb15e087f729d09e75a
zc5b4f13480825e789a389d5ea9a0678592ebdbc88bcfccba0b7a78dfccb76fd455c92f17c9d7d5
z97c8a7a69d32b30c783f57ab24a4491a0da4084a48c0c88cc519771fa4d5d8b8092b152f471c1b
zb354b1143c6f7db19c37a7d402bb553c039cd20af47d736f3bcccfa6c3a08db0180160d1bb57ac
ze6b29ca0f866f21a70315f0679a753fea0fe1044e51857539e9fe69752660a460241df5b4ea80c
z26197558669cf108f54ddc21bab14d7c68529607a96e51768f80cd82ea4f6c870f199c4f673de4
zf651687505a87c6eb942c5d6d8b9b3e54c9da39f62c244fd8018553702c1fbc82e1fdb3be18d7c
z3b2fdeb922c355970175d065a70c2e2101b252a350da9d59aeca68998234a32f209697e412b056
ze7b2a8faac5aa9cac7843f49842b67b954871f2341d49d9fb62ae678805be3c72b46784f535bbd
zd2c1bff03834418cd129276bf8befa1ff8665b64217c2729062effe81b8f1d7e71292dd24efd26
z5e7b0f72f181dc7455990fa40f2cd2de75a0949bd0b449ecb4b2e0bd51e4fc6f0e5c76818bcca3
z9ec8a2ca458d7b2fcd5041a6545617f6a3c2ac14051b64d6ba4041d6f3f5119d854b04be1b7864
z5dfb4966cb500d778350eefcdd39d1d0fa836983c17e980139047f66edfbbd27f38eaeef059306
z0471e0a346f0aed215f19f658a259d518604c6c3c46a8f6a42bdc70f00c6817b56da2da1255bc8
zcf2c82652c83bf0e904c41be9ec1a70cbcb6669c8757649171f992e186b04a3fa99c71dc803ef4
z084f03e2226ea11f85d21af96a0ce2f29a49e5958fd578bd7b764d40e6304bfec5944276063957
z0bd64be243ee8de434ec3768739141ea47d3d53445a98ecf4070a8fd7a51d6c30afbcea03e8352
z9aa38bfcfc71322472fbf9ea950b9b62422b7dfff9d772714898caa6059c8a466ae30039a235c4
z3ca9426be6cd85c29150ba221f00ead51af1a76f750d1fe307dadd52d778c2b8d0afaace15ec43
z24683faedc20af72475be819d8dc54e49b8ec2108f18ed9f0b4ebeb086ed412d192ed9bc876122
zf3ccb5e6e408a975c3ef9a4e5a2c362465db474d562aec90d67a8ca100463af163f4ea0e4efdb1
z632e0e718c81c7f04cc3de383b7cce579758f7f15da22a822dcfec9a51a2e4c096e31cda949534
z6025329c2249a452bef36ed356de8344d47dd3ee2eb420c245099c53ad7822c10ae1f564662162
z11c811a05a966394fee084936fde07663efd6fe9c774470f036c778767863ddc0e71dbbd7a1451
zb2f6077e102bb1c46600ee43e59eaad0aff5ca8befe43ef59c7d9e7c0b3002f5e2130048e7f960
z6d14f0c34e174e6ecd3df10005bf5d45db2676c6a7112cc3d0b8c24fff73d7829331666574e419
z5d6d7c204e6cf30f9efb6e727112c8d31af53e5edab5e5d42c6732631598e94363bd4aa1bcfe6f
z44b92299fc5f4872938b6f9e389741537a05231e3cae8738165af802685aa7eaecf82e4cc2a8d7
z4d33ed1fb87bad7874d023e242a4e0c5de9b7442d628053d12455eb79d9577adbbd7df6420022c
z31d641e8a2c2e5c1da77d97962cec36292dff2d58ae8d88c2e158458d8471d97c6b15e212caef0
z8576aa62a7ceb079c1e80bc26a6e37c87ada6ef07f85793f6b6439f8e432f92e2d917b060e17b9
za554488d2b5bed92208dad61e84e0e728e524a33a288a481ebda491934d2f29ea3be071999b221
ze33434e941e2365fe36db27f8ca8d2709e1bda913034e3c03c2ac9b2530491c219bec73add6940
z5f2d0656a19b803630fb46fdf3b6c120c6c7bb40bfc2dcfe7ff895dff9cdc14be9962e620a229c
z274b18102d88c84a5e06a609b039a0d92b3a22f9fba2dfc908c01d493e1a0c2f7991bcda50c0c7
z28046f193e7dac572bf07fa8d27e9aaf80eee3ef4f7762fde6d701b5011dc32176224efb423c93
z900010bc8093ff0996a393de400a40cd02a98e373ae97117b7c53b90b34e3998f39b695ab2edbd
zf98f95e8ed7200f2e4b139b999a1a6f042c55fc6f3afa3a39d46f87165f79caffbeb70a27d707a
z0ac82be7ce86e3f4faa1559297d4b083f73f0e2adfa2ebac0aa728ced952e2e9f96fb0fd0227e7
z5fd2a7b0863cde230e0739b0fe00134569b81c55e71847fee8df0b361bef8c4a503b081e5974a6
z33dc1916e46e38c61cc524e56b5f0f06563697a9475e4a4d76e1ce480326e3e7802f661c72d9d4
z8703324442991e2725b792d49ff14fac7a396f2763b67c456548f5d87df657591498f8f6794dea
ze2da1b36b508dd13071d6457feee603a3bdbdd1aec377f3a972bfd7db3a7381f6bd59b39be6ea5
z37c9be8a417f1796ed7ae15ad4a9cce5efb018f600165961e46a5ee48cb784961d24a2a231bc3b
zec2b3095fb0937ca43f06c0fb9bac1c1d2645a52b78850616e2a4223666800bdeb37ea1c646d1c
z2ed4b1c5932e0d8d63c7c12487d12a9480e95b408feda254f7389cdcc2f907455608d38f513515
z91df1a162d93375b3dfa8401de5f786fd4024fb3ff9870d45a901373d59d3c36bcedcce62a29d4
zf93b01bab81a2ff3ec872753b3f13f0dc9a2eeb529b3c597a5d88be026907747159f29094658f0
z8d2adbe816f81fa50bf88c563ea509bc92ac8071c59994f98035ff4078b08b9ecc0b9b0a14fd42
z9ee7557aa4996101fd14f07ce8ccf899aa86b5256636204f7722fff74007d070a4d9f76f51dfa4
za6665222b6618bf75c0b7ed040443d25fe490552e21d8d74ac228b62e5ecc56246dcf76812886b
z1d59224412cd28528e9c0145c434c54b776acb213e489cdca7e952a3af29d65da497baf4b58112
z0cce0614e2b006027e1b85c7256c89a996b2e63aa5be462b1342ea7b32e6555bc8ce6a7c2ceee8
zd57cc3bfdf468000ccc1917a4f33896e1b65cee971e86f8882e9ce346816c11b7b56856f63b8e9
z396a7e0cff7d75fc1c5e35aff3da1a0e1797089a54586f16c672a77287a389c07adceb67221ff5
z826ae6577d3046808956dce32e90cc98d3193eaea0a43835c570e9512f9cfacc29a11e738b1aad
z1588e01ec1c1909773fd5ea775274c71df36b049e15b9518706fbcab8b6ddaf5035aacce51fe23
z77e65266167bf55eb4772ffc3d5f644aec506372fe1cab47ce6bbc5e7a96df754ebbbc18a41738
z954e9074a08c56b312da7ab3a35b19727aeebc67033942248ed3bdd43baa1f96239a4129934ee0
zd0a22d4ad9b656c0a7096cc0389efb60d0c846a9334a37df7398b0c00722567d46c01f44846d99
zcd681c5a1054067bbb53785d662083f4c5188b63790326fcaee980e388f8ab1594669cea44630c
z9994fb5e5faaa29055765ce8f284f1cb3e08cab1bb8da65340ba20da77ea49988fa7d152a5b1d3
z68480f829b53073f8583bbf044a4763e0f5245ec44a351173f8492cca8a19dc37f45481a31700c
z445728b79f0c315327d4d78b6bf594c97d88b9649e5a1a7044ec2f4a2f62b0d003f3ca2a569c5b
z1d9b1e1751872e0a15e8a413e18ced4f502a3a2fd5c0862e8c0ea269d9d1e8641edcde778315f7
zc3cf5bc428e63d86aced966b7b656aab77dc34bbb5e9ca3152e9b2b21911623e6bbf32cc9ac0c9
z7ecd9ca6e021b51c3f6de13029de3b0c2e520f36169040bd70cec84b4ac7ca2868308b30e48229
zbb1c2f75d82535063447020f0ff798226d3730ac645bf35e28066edb3e4aaea363f0839d6f6cbc
zff74b18f78d63bbddb2adad1e8a30ef7e9e774fcbf2c1588981c8f64c48097cf1b734550b26bbd
z77f48e55b2307f51ea721afcef516dbb89714cb9cc750b9f1eeb248e1e66a1c1dfa8289dd3f15c
zfbee72ea146f5b04587b176d675c434162425fa070d34c489ac3675bca832ce876fce00f5e8bb6
zd7fa038fb6f6419c8b5d1f7284de2f114d57b43486da7d69c86710dba5ebcb2c5ea21c6803cc6b
ze2a25d8f48b3cb330b31c71fc68810ae5eadde097b5edcf7e8edad0c2231caa3da9ee235ae6bf3
z01dfa4b1e769e44dd2914a12bb6653a3fc83fcd71d31c190fa35d0b4982c9994fdc9b214e2de2c
z33b0fdcbcf7e79588b67047e7c5baa0a4e69cce49eb0d0ec101eeedd1f2c4652195049edc4eed7
zd1f994b75f918f4cf7491ab2dba006d8658cb28c4fa13b3308e7030a135a49fc3b6acb655ca1e6
z5d646e0453fff764e3a9e028063013e9cc839609831effd4f8979f537c9439e38180d4259b254c
zabf3a301d5c465ce5310afdf76a759aa9c07276cb0e5f5544d4ae8a620ca96b03cd16919f4cb31
z6c0be8966e777f7046fe3f922cf927a0d9076919c6afdfb77761c53e8553a34348e710c10a1a5d
z07e28aee3db707ffda5f1f829e449235fb0a3c37029d73b7672bb8325510da9818adfd4adb6ab5
z4913a30f2a49eeb66589654846885fa2b65f517448783fec95867c1b7fe542c525262799b7a597
z95bef2d9586624fc0b23be338aecc6d8213325170f6a1935ce7c44bf42e4a8ea280a27ffab6b5e
z701403d5b526ea400555df3843aecf381c544d579dfa72de9059328eb16e69f7a2fe55425832cb
ze27e8fda32aac027d936ae7e9a194561d068db3c9ea9525316951240c87d53072c8f7ebeea0553
zbe592646773d6f3fa8bb8a1fe815375eebb4c52b1c059411f89f3fbff866fcf73b89c4bc314db2
z3d82c161ae62275ecf9f10a13055a78005e3ab38a253c93481722f0258bfaf028d2cfc501af7b2
zfd1e4bb13bf1df8d220304e9320f2f407b4b9abc0f85b45c9255666371a226b1e9f40915d037ab
zc8a73d92b0204154597c16f621c33789c050d074a449b51d473b23eb7aaf66969a1bfeefbe5380
zd456baaaf9dd09a9b32fb0271e947cab9d473a9011c24882874fa060e15fff9babeec9f2c7452c
zd973d80f5e14e7140cef93c7f7be098c41723fce4a34810870e64cd56de8caae88f1932b548d57
z31d82c1af8aecafd5aa5ab34568dc9870c9cc4a88aa4881416a9a2c4bb900d0b72c22095ace48b
z93d01a33c143636bd7d730c2ac836bc40f3680b07d64823acab2ad4f2863c19fbfff6f8980b3a4
z9d8d0a5e8c03f335f4c874165130d2cb2209bb95166fc5128bc8065a9e58772f6bdcc5467dad82
z77bef6a4e1f0855140d2a3621f83868fe7364a6ba18df409a39047f3ad80f181dd2f6b1adc1df8
z058ef1348fb741878b6f364885ef5c5112352b9356651527826ba9656c9a5eefbda1ca7a45b66f
zdaeca1986545280566ade4c66fe1a8483b60cb3726e9718e0095aecec6b526e1c286f1542972da
z1205d050ac0503bfde76555a5b810cd748b8ede1dad732e42e12b25817eb3e81253f5263fc960b
z1a4e5383a0467f698c80ff6dc4142d8fdcfb9fbb001dbb16b6bb8c5206d68e7cca7fc6a6719913
z2cdd3506cb00d17e919fe6a0d63b76cbb7e49768e51b7aec66429f099f8b2d17c09a6a41bfd17b
zbe24d191cf7dc9e1b8a681ed918b9beede1496f01997a4f1999f1ed90543a858e87b35d617e452
zf68b17d2a61aa9dedcbe9f1f9e54666b475f826d0f6d17897eb1a04a04b041b50d5982803e18ed
z7d3cec7af220cb94b77446b566eb2f1c1c8e576f101ec250eb77cf6bd1e248a67df16d6afc55ac
z7e1789a6d6558ac2a51359c6336d29fc265f0cbef842af3a259f2a28e9c54b658f649d9ed21280
zb1879bfe77aad6c7637883c114165fe8e40789ccaa87b0ff11224688cf0ef2161a229f4d3738dd
z55667d47ceb58b2a253dffca01306ec4718da25aeb175dd2440c29fbdc05e94621f7bfebfd9296
z8b08cea979c5a8c5aa5acbd20ec768cba9dc7751d8597b2de5adb684561fa04fc5b8ebad972e45
zb94c39ea5644a8833abf08701c0645830da1ac6dc0362430e9f001ca2ddbbe7f07b7840f384e49
z7d4ffbdbb68174e16b2a701fffbe2e39d1c7afd10f3306d3617a4ee66dba83ad1ac6632301e17d
zf9a3dceac03b313663eaabe593ba1da9773a34b51346dffb57a7f06a7597ae9ecb8a2bc3f685ce
z37895bb3948277740eafd130fc8cd596d823c4e5bbd55ea70af5e686512b48c59afc9baba35852
z8f30d734485da59678d40d0985150a617c42ab5d7f67103a5c0ed89c83991057648a6545ae6827
z6fef3e50514f3db465997e436d38b4db9587838e3f35a09f7d96e5696b697150b0d2ef1ba4b2ab
z96c14990c6bcd743fe71237e7a09e90d551c7dde79a34b96c9c5bce6d95bcc6166f7aae599b1ca
z3bc5a671d973592f9fbca74138fcaa945f86385562a22e44ad058fe894cb99f60f7a3ebdb6fc4a
z76ca2a6936c25e7beeedc35c566201b50218cd404c39d5b5a417c780ec13403feb348678236a7e
z3f357ae687771d1e49a2e70c4f0d4123028ab67181c7f974f331b150e5a1342834f5d9f094a4c6
z2085774b7550f5485ed21ce6f45d7247f2a83431a338f53a8a8c2ddd4ed3d6a005f04c457fcdc3
z5d875ae718c9ac3a4a275e8058b053f8915342872e69f25c1ed29833538ff4322ad473b5e13edb
ze7706c523489f19ba11dfa49411a5c216704ca1b1da840b2f828eeb8d0dc99a9866db8e0762871
z9f8a654d601fab8d45b495e7e35d3214671165ee9c10d3fe8bb7bf8e056e96897135c52e58e012
z6310a23c50657a9c8e87574ca7c3446c025dfe794134789bf96e22236870c9b58784732c5ebe4b
z54fa8bfc9377a13381c60bf9680eb0f1d65fd0a55e640392e58fc01b3c651a1068ff99bac14822
z578a16a1340070452bbc41d9bf85611eac7f24a1299b9cb4aca8bfaee862fdc9f55418131d6452
z09e5ee5307ae822b716095a0175d03632b06358d027352184b2cb0349cf62a7ef22b8a3dd6aa6f
zab9acad356325cf488d94fd22c14756b97778a23691006c472e541b323884cd120b37b11058bc6
za5e74048350c2f7fea0f5aa4d67d7b388cf9aa0c56625de6c0311b8dde04509085f969273aa5dc
za008fe04cdf877b0f52a09bc1d8319b03f1e3d3a9ccc8f5820be4a03e1dd4a5e8fdba4eedfb371
z506c6736033cc253797777661f9ee1b4425738d179924ef8d8d9a9be640a33e46cd58faba4a817
z482394cfdde6d31b095b89182483257f30e8dc7d73276fded837459e2553335afdc5940c3677c8
z58073a9f1cbc227f0f97341ede88ee13711aec1266cb57fa23d5fc72e3102434bff50606a2db86
z443dc0b2447e8caf1e67a3e936852c9b9f46b635530a1ce3489cb06e6d714ddf8a47c7334b4642
z10f4b1d8f12944e925bbe0401ffa2915fe3cd1759e834d16a70816b45ef048eb61f7594494a59e
z79fb042ba35a4e551e27e30be596abde9eb69263a12555b05e44e868412b681c97798a2a26f384
z90af0ab7c902060973fc922d56235ee82a18c4481384b1684a30627322af4377d640be090ac094
z2f6afad3c68ce10feb25d17785c2467d93f8d97e2cc6cfe94c7f7a7ed44f3da2578c7f93f31468
z411f719ea8574d54fc6478328cb4f6cf28d9cb991153dab6cb928f74d480617bd8eb8d8ac7e488
z6adf5eff77e7cdac4f8ddb704955ea5e1e39c4842a8a1f9bc3adb1b3e5ad365f23b75a16ec130e
zb0711d7d792b3657b640d080cfab9e16f3112abf478c3be5bde28518431a67c9c6f38bf4841edb
z5c1137117cff131a7a4ff5e6741a1996582322c4837b6b325dfc147c7609bc2d33da1217eef156
z45dfff8a44a675c758bf40e5890aa5fe44e18348712803b700f65e2ee0e89e13a1246b544d8c3c
z0469d4b5b0370a4f2a415f15f949cdee12d70e1b004f80146a9899349d0d91287d182fc7e0dbee
zf4cd1f9aa559c6c55d51778eb9f214bea914c960e732d63a39d210923790ec63eb8dba388a16c2
z51f4c9f852f9b5e6a75ba5894be4d91d2a8ed7b1a4171cde094fb90b44d798ec9de859d61b1939
zbbb0a9bc4dca145f6d6fcb2960360d70297ce5e5b18145f3a317d74a5de727e70c4bcb8b7ba437
zd0d93cd07f536024f4372acbb8bfb4b61f2206ca10bfc9790d685ee1d1a216889fb3478e8745c2
z20f22ffd2159186f999de3af342c7079075b82584973be4399c91fdaa829a24219b66ebea30788
z8bc13c5ead6bf6d23996f396432a187c91d4a5c36ee7e89eaf0677c97ab8ef1a77df10a34a5e82
z58387a9e7a2c9f59d7629318489b226a85e9a98d59153c4617c9d4a3318002e9e2e35798f96d71
z5de17fcf460eb679e9676e88ef673123123d8df3b225eb09b831f27a883ad6ed80c55039bfe5a2
zee11bd15a7c94ebd0184d4d6ab090b345bb98a539942be3e17211440f12960a0760bc8339178ed
z918d59449a65c934f9636a68a1d030f2e372e1c4ebb2cd81d7012ec9f54ea767c8e6079295f2c9
ze6b76cc2517491fdec46bfa5dfc7076f9d2fcd051fd1df388b544250c2c69406331d85b96a644b
za00284b4ec2177df6a72d0e7ef5278a7d734ad9e9b06dddf0ceaccc8593ef8bf5450ea2b956e21
z85e53cc3931e84907a6669a1f947bd43fe8e7f3b372bcf72a098e1718a073899ffb6d9d5ebf535
zeaba219131a19ac9995aa47b84458fc670fbdae2627032cb9a81b1485a1bad54c2b65291a79ebe
ze80caaadc12c265e0c2b3937d7e83745862907ed8af72c28a15a62a9912ca06734e233ce696d5e
z63da8a8f440dcbe0c745331bc5c815ba8ed3231a5da10961afe2c2bf90096f1ecf6b3716a46ae2
z81ea4dac00c78342d1d7e1783e1d02a6ed5a49ed00b9f112ff00e995f726fe5e84cf17fc6fc002
z71116dfc7b607a8509715cb86e5768ff8a251d7425ca30343754e7ac8d65a8d4f1aa52d2294750
zda863d37e48a227d7c12c8adf16d027cd622cce5c0257a9dee50b21342e0600162012b3af395b8
zdf6bb1a7a8c60f05a7a74e2e2e94d35b664049e5a9a292c277332a8e878df7cab08cab827364d2
z141878c0f679cd9f7b0a7c5fd3fcfc9547e42ddd66c75abe360d1435285b859ade77e18b6ad90a
z434e1dc50c431875eba5c7dd18c5a5de6fd247c41a368519290a7d740337d36c9c71022faedba7
zd93b86a08fedea04efcaa13127bd833cea89ab7375aecda9e9acd566ac743c5271b844a8afcce1
z45f9e9994132303b4a46b73c5828ed71636867a77198f6841a3472bc1e3c09d8f7f861a6b89480
z8f3120908f4cf447b6790c7a9cf2edc72831fa6d98377503a659e2cbbe65a8727f48df805a928c
z82a5fc3a3e9cc22602c39b6abe24db70995547bd86b3921ceaad977a537cc587510fa392b61808
z3c849dec1946a22f78726eb2e5b7d4a5a86c619aafe9b60e37ef799c5c967cf15ee30aad2ae78a
z624343d5220d11306e20b355bffdb1f43a01c452f341d0a2601c2f3b8a2925a11577e98225a22a
z55dc90bd6a237a50da9b822cd2ae77f444065dc359de61611ce6cb56c5f06405f58625c0d3be7a
z8442d7882f7b1ca87e188a7a25120040553638d3f3bca825f2b5367757ff52ab8be897e766890f
ze3450fa2de51aec9e7600ceb725d86965601c2a897a01982561606a5a0b2c9248602d2b9436f48
z21fae71c28a5d9911ea6e980947fd08297603ac5bb156a5af1547b88d0f7b0e282707fa14ad933
zd2ceba3d428a05a710c4e01122cdd80702d6bfe190b816a49bd04d95dea25239c884543914dac9
z57ebd393b55f1f4bd5fec616285f6adc910af0e2663405f88842ad0c8b5fe171c14d04012c3593
z712f53f072d5e37738b13cd6df153cf404b5cb6ee97e132ca4c799dff5f3a8c01c390dba99e153
zac18f1896c0a6d7f592b590550c5916ff441cf071aa974f1f83c956e5d282bede787bb3baeb689
zc35bab15690ae88fb629cb7afe7558a5600c9e88217229e5625cf7f548ecf9e9287e260c58c426
z9c98fe5e82ecf20d3dbdaab26bc07b86c8862b00586c01023fb8b73d57944076e9acc1c24d5220
zec4d21fc728719f08ff50e009dbaa278f1f8eefa7391d34edf7fa4c218d67cd456031235bf7f56
z514679fe405e8d5c9f3b2e0c50258234ca646fce7a5510d5e714a9c0a84f9db632235ce30e2102
zeb8a458eeb23f6fbd784678ef0d18dbb8ddf839f358056469be6e8515d9e371ad545e73f7649ac
z165f7234b1556e888afc74990d11c504fb3830f8776e767c133d7cba294530394133b081412db6
zd01b5ed0b4d912a05956d5be9c4f2fd09973949f107b6caada7cc7b8a90617175a3f5192164228
zdfdbd39df1da25b7ecf69e6a1f6ef6b3984b8ea48f0c8a6b1123a4dfcd9b69e7d868f28dd76aef
zf0f298c70dba493fede770ef69763337593d3d06e25d73b76c85adac902794f79802b1b42a844d
z8759a24bae70262fc82efb75001a31c4d3c1892ac6be33d0ce3d46c8efa557b4897818f06cb38e
z41658557b23d809b442eb133a7c66363ef65da72b3e8be1fcc6ef9e269b54b86c224c4adf21e73
zb267312e519ded8367eddbe388db7d3d28b61c6df454ce220906d59277c0a7371fe1ce07fb6929
z5fe8a98bdcff8009108be580851e6c878f03680cd59f7089ee4a5c027ba7b3c8565613f0c68ca4
z32c4ecee6cf674b8a558395a79e61c2acffbd70d2bc644abacff040261f333b24091a2e285472c
z09f1ff9946346e8a5c4fc07dd98c87dcfed8dd1fa8c7aebaa821d8309c9abec09d5bc9c07f15fc
zfb9684514749c1db6bb15557bc16178acd0464e58dd4d0b53d9d3920
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gigabit_ethernet_gmii_link_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
