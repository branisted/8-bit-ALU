`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026251e18d0ab5f991ae6977f59097
zfd09fdab6b6409e7e0a1b9964ed96e3c6b19e365696040da73432c85429c758c1172aa36e7d4ae
z15f3667142a7ac89d952acd463bb3819f5c7d624ddcb2a025ccc36be408c039904aa5c76db930e
z528784e18481378e2497638f0cb57850622da56bc84fa996cdd058073fae8bd7f4c22ec641596c
ze86dc6e6ef940fca0e2124ff9774229749deb60a8c1c358f5d82e60684892dab5383fe63a556cf
zdb66397d055cacb01ee28d4f04a36dc3d722a435074a3225e6fd8f406ffc497dab3981ca6d2940
z656d8c97db2e5699175630397d53c14683ac087f39853388ef2921629d649a06b4b4a766d85aab
zebd355b007043898ae1f8002c023a26e58c44c262bfe6d1d60b1903ff1b56a082944c8d3b6ab0f
z30c3d4759ffaae3feb89e3fad854c227eb5801f21c6738fcc47225e19f1236fdb23c02261f1212
zf0413d4bc275f99903d4a137aae19cc3f1756419f525d5f1beeaa716d21579c797990c2ea30ac1
z522f7dff6c59ec66fe63444ab1c28e50b47cdf2f7c2e7721d1bd7708e50377616a0bdda34796c3
z2f6e6ff488b0ee9a10fe73f38030faa8bbab5453500b7eb083862ac2b24043eb06acff76a15664
z33ec7887d67c975f9a45bb60e829547bf7b13eb71ea95331823db3764bb73a5b8a5afd8af8581f
zc712ce227bcc564e0439e64c253f6dde10c95bdc348428e0f82904a2b6593c166df6a143f26ee1
ze06430f4ecd2dca75bbe883d45a049f1114d3ecda999102eb88be661ae1cab766965cc59127395
z926b5732bfa04fd632f4159d39a6c77b33f54f020ab20b51b2fd5c383c163f728fd1e9944ffcc0
zdb54138429e197b75c817922a46bb0fa749a1ffb831e09abec382e985d841aacac09568b0856c2
z6503ef7bf480f659594ad17754f8dbbe0ef9d365cc81cf6596beba11440ef18ce57b638a61461b
zffbbc543873404d3732cf97253b26210a0b854cccd065619db78ffc18184985057733110f6bc8b
zffbf6f3fb93da57a2dda6b762f1bd4b1e74e0e960f05448093ebdf9530f5cca24fb57d9f914f22
zd79063fb24d465b6a207b1e71a2cf26eb914e4ffdceef16407df383b4df0ba6aed81c5bc4bf4a6
zd4415bd5f1aed71b8fe3fa388785c87498a9d7c2303b80a45e2ca7b7757d164d3e7ebb239fc150
zd776f1c3a26b77118bf77993ca0c18835728ed686cdaac5e939c985cdb8378d32562add2aec0c1
z6ecb18a974d08ba9ffe4f9ced7ee8ae7dfd1778c20849e4110bcd8e012155cb9018c00beab2516
z90781004c416fe3fe6b7aaaaca9d5daab563901f3412546c021ada54ab07d45ca8e783a51026cb
zefff78f381b92a018d1a34494787145645fd6ec742856c55036229e6aeacdcea51565bbbad423c
z8722c12e73c872ab3498e16180c5701221a90d65abe3ae60ae0446d592d487159514906d7ba853
z3122144922b976e0b881497cac97ce68b2d1c1df86235f2d6293e656d406ac0cc580917b4b219f
z0fc971ab6feb54ab0c7779d5b70a671269911afb5b60f03cc4ba01dec74188cb42378b8132045d
z0c35225a745302eeae1ace93461d6428a5e63773e11a6eacfe58004bae75979f77974ef78a0ba7
zd57014d00dc3fd74ad89508c92d3a667569e7d8b38534bb6ecb484dc03ab880b172ab0c26cd92b
z5c1143042d5aee27252b36b09c1eeb9a0d463aa15d46551d3636c339bacbc5478ce5c9c17402da
z2b15dd84253b1996cd009ae97a12a8e1273a385f2083611407b8f02991ef6c1a0723b44f5fe2e2
z3e1174fb0dc1d23e6646b09e6905ab24ddc5b0e647a9e4429750dd5954f9408eb4a19be89cae44
z729a3a35f692bf4804c4fb3d90e40fba7eec98ee9c713bfa510dcb32128ca5c11fc89666c55659
ze14f2b1c1cc3d729f521ceb52d9ba1af71a2abfc1b9146ee7092d517ac3c21cf5370532369deee
z47aefbd920f87c72d2dd1811bb441ba7fcd0925607c3d2851eb0fb07074a69802266ee3ad3abc3
zbd562819bd1815b40b85e0bc07631fbf450916655f20696e6b6a2b4f1a8dd69b8f31536c33b88c
z7bb0bda2563e9eb8068b6c2a5b7550dcfd29b4da1f761995441aaaf81b898d9cb99f1bf8fa2675
z5f4dcb15298eeadc47ca372c220821e36759fb89ec55a25f930b40a6306ec29a7a8dccee0e131f
zc0ecc6e8f38b787427fca7d8e53124b770e24729b23ee61489e256392a814f225b6b2d8950c8d4
zae62f0c740dec00106e9cad1cff0d400a5f2492391db7ae76e28a884b72a7a74a960460e624b5c
zc6b541dbfe2e5ada30dd62625fb2b9c9a87e81755ea720e2b95538105239a2985107eb0cf40eb9
ze32ed6daf79ea3f3b585b7c39da175df59ad2fbf8ec33a3dbfc6d44118d9d0c0c655442046cb9a
z35f98f3396c64e10809ef7b06053a96210db64e4fafd9dbbcb3b4e2110aa353f81c8a5188256de
z391a6d21593a136bed4fc2db8dacbcfa36267f87993e81fc3f9605b633cdee52080c253776ea6e
z9e570bcd55a248493e8011d8a09c11e8c7495483389ec46bf6ec8eff053b194d7b0e4ed3dd17eb
z2749242de9fc646a04bef87729966a4e25d88753c5287f058e52ec77e679e672a0c16c5abc6adc
zc41a5428e38093264027397914bbafb531031f7804cec436c3d9d4a7448c926989a2b77fa54e87
z1f6a7f932e0ce3b00ba9d1b771d8aa230e437d7879839c87b95d0b0e16d0036978c98654cd453f
z7510c310906aa13a2f3bd28e0371392feeca39ee7c195c5fdb3cef9475bc5b8802839be0c608e8
z38c0bab625e339bca8d3e50b043dec0d369af3012cfa08af77ada242a156f7db3ba7957810da58
zd61ee5ad89ca2a47988b9dc5ef871d54393430d0718f36e98444545d28f90f3cfa956e6a45d28a
zf949cdc64a80907129be6ab7bfb999c031a71279aaf41edc479856f7c9510e3a1864483f9439a1
zd582e5edcfb584fd98a725d0ce270b3365d11f9ff07277c48f64ab0463a66302252f1fabb1a6c8
za0d0e3da75d18b23c230fb4f563f9e7460d231fba9cbbdbd5c073f22ad65099729ed52f897eb8b
zba55807757d295492c387e1ae080274c543d97a4f8ce46611262a0e3a215841fb8c59e7a7d094d
zd95ed525b9bf71200c0b1fdbec8b8d08526d3b2679d9cf78daf4384533760795fdb3873d644e8a
z82c60e2b71d148fda7c958d450205c47a0fade45b0f511ba041aa1781e9db21e16d8f6e6904d6e
z0d143fc7066210c7d1af3e0d270392c080f7b25f1a4b576987b0385e9155490af82170606d59d6
zadcc459c30039ef6b302b3733d029339450968bc77e21dcadea1155c7c3f3b87d6850c50c0bfee
z84baec01a78074970577d70038b589acac1a24415d793fe80e724aad23ecc708051cae383e15b4
zb0ec36262afa4eb192b55084699f8406501c42ade1d285f4674e141729343e2ae3d46a2f2ed1cb
z1b5660de2da3c8900043c33916bdbd6156c066b7bb940d1b6151206ce98c3face3228f5cd617b9
zf093b738759ee040cfe32847d77bc86d1d52dbc0405b891db2e14d73fbb446a98c64e62ee9a98e
z9ac793946493940c160610391cdbc977db8d98047132337b9351b915cdc2f8cc7eaa1b957a2d62
zf3fcf608b5cde5915ca6ba68af8e9e28296696c2a4dc658b06144dfee7ef4868f934fc63171f87
z4e5e7f717b2fa96640e9eaf7f64edad5d1da4c7d08bd0a7c59ba6e05acabecc264016e9e5da060
zec0a107a8a4eaa8a372c5222ded068ec68db7454b0bb5ee9cbcb6ad5a8f0bf4fe7b0338070d22e
zdfbbd0d5db03a5ace7b20672bf368e86af368e21f16aa6d9e4b0399d788195a15742cec1dc7ba2
zb265b51ad97140c07661e91799f6da39ca4dadc092b39301b1d043075bb206d6315072193aacbc
z36f453fc3d389e181e12e9ccb6f70db0e938a02b4455e1b565fe3856438ba6edd727cd1243beb2
ze22cb86481b80fede1347bf304b12e9827613062446db9553c398a40a8c4eab8c7213a6a11bd3d
z4532b441deb66af33dc7bc0c2364eb4b82cb860ac6d2aa61dd6eecd35f6860ab6a2e390d03999d
z69e0437242244a57baa1a72ffc639b8c9c55e100258345d0bcd9dfaa4ee7c2e05e21d4ecf95ea9
ze5cd186a310acf3cb5a82659590e698956b1b0ab19937157d9a8decc05e877c309b8ba085db7fc
z6110ada56f35795079807b0b854034a0754b55e226f37acfb384f4b1e34dec203684e2a0a26873
z17a9ba2f75956f808b35868a27ebcf0e66d815e60bd6c707af8051cb80f91283a5e542a6c0360f
z655acf7a9ce8694025c320b6f0fbad123ee315f712fe150a59d52b9f7bf2b5b25f3f45f11beac1
z1454a5f8d479aad407f710c20f5cc0a5ed761c77857a27cebccc3848767ba46dcfcad0d03d5bbf
zde73985536d5aaae8e9b23adaa06b34c2dc4a8eb0238a25eb07c73a2644bfaa1fa12c6ef754bf2
zda975dd9361b06ed337973cc3d56b67e08a84c577aeaab85957c7f1b217aa2e10f07c346d3534b
z046c858c5b3cb49eb2c968bab3143e4a5ad08710d2d63e362f406dbba49d95cd1e879f3a34d2e7
z32c7a0e6562e96c62d936eec0b61f27829dd73aef6b41b0bb23c739869a3d439051ce4c48bb512
z1d15e0bd0dd6f5eb86f6b8d86e58f16c408a7e837929c00a91b6bb3488ed542b90071ed0802019
z20dbfd5739b30bf1cf656dff2195aabb7d69f7014e9685cd81ea1b3c99e0fe979adac27abd927a
z2eabaecff46640c2fa7bcfed2e557f5b1b5b3006e9c2e2680521d7fb000ac198068ca5916b9ed0
zd9cff7a9afc17f3c7f59381cc9312af0adb22ee213c10d8a65c3762113ef1e6d10768149223808
ze7b3eeec9fe3e7bed6c24a18887fc1d13e2ff8fb966e1760c436c01689d1396657604f00cf3ed0
z278dce4aa2d4caa0e79bb0c765eb0ff594435dcae40fcae064bb9561e7d94d5016eea0ff2ce90f
z3b6284b57dede9874cfc27154bacc928b07264f80f15f973b8f9e3b8b373ec678ab49f0eedeb3d
zff02898576cf725d803ae96326f796b4cb79558cf905bd2c4de2413cd48afafa6fc3f3e1f4450d
zbe7db85b47168869f75ab42d548a2d69e2acf1c524eab5361fc2090aeaab66320e900c0f8a1130
z788854b463ce66fd0f57c5d78edd1f81df7bc0f898cf63e328bce12b81994bc792a7fe3656ed91
z5bfcc469bdbd10e6eed81c6e5bec382caa5246c567a73ec23240d554a32b2c654908f50b2f7470
z8b6083d4715503b4071dc6683ff7a81b9408f454599c3821fc81adeda871a866629382b98dc335
za1d800035f624b8e2a728eef013f37e9ffd408fdcd7802c00503ab8e0f287605db83de5d686db3
zcc398f44386ea7dcc4003294491cf9c6ac3e2a095151ba26e8a3a61591927c57bd1ef0378f6c42
zdafc93617d6bebc5b66b9596ee07d167ee5e133c5036776f0753e5cfa2c7f1e2e57e6af14149f0
zbb9280c361efafe045f8481039c5e58e2ec875fde15d5a6d66fa7f73450957b3e66151ffdddd65
zed9a5b5c9664a70020cd014b237723c4331b565a8c294cbea10e236defbdb9b54f022438c4d14b
z8fd0f4b6e5e7bb5e3225fb986b31ec99a311a64374cdd303ceb394889a930fb136be4a3ae74871
z57f3aa49a0ba220a502337637d88f52aaeb759ff26202faf65c52d52900b2f7669431fd2ad7590
zc585f8818eaf65a48956d03144cbaa414534b1a1717b7bb1f096f6944bbefba87723d0f55579fa
z121a33c3c9b509b1321d68cbd2ecd0661ef171a2c9b6c9ed020fc50511f290272f2aa4ea123a5a
z8424832d45589bcdff47363570ce28978aa41e94680a11e4f4e0a1c330362c46f1314f2885c406
z61ca624135277eda200098c6d250895f7ca81da811c50a5aa8aa20b135ab5bbf928dd2e57fa9de
z5e2179c1c445381b7246897e6ace637fc3f664421938ce09f7fb4a1538b2dd8122f77020e50522
z25e763c71406f5dc907e66edd0c2a769e35e7a8a034c4a2e9575bdd91c1b225862f4422092ebd0
za38db1e64c02e8b437265c08c9b13dbab3418aeffad9f2087dca500b2159c61e295d7a8450d8a2
zcb8f5593b843a577a2b0cfb287f49359a7a7707d3608460b5e902d8d0a28d6a3e370b96df3dfb2
zc97fcbfcb8a3b5dbbadf46c3f380fdc0ccb0eb84f8fa7a8e823a6d9951f13dba485d04c1fa195c
z485bad008464eddaad13b440d05257c19b0f264c30685b45fff648aa0de62cca451a318a3af26b
zf1f540fa956efc14c82528a3870da8a98de53c479d3523b3b3b6b99ded5d9e9f8a9f7e7379d21f
z0c356686224748d7e8a3bc0272104565260c3a0cd0b3b3141d45d6f3a37174cfa3fbd4527b17f4
z80f6530883e975551b59f00fb8da00c465461cb17e934a0ea39002001f019e2031970d1562f8aa
z71bcf4ef9551bba434d3ef3c9c02f26ac426b9e41ebfe36bf74d6f00e0beae08cbb07cbdc0c0a0
z7ed74011136092d937e07acf80337f9346cdcd769ce935328757d98240fc55fe44e505f417ec2b
z567d163c6337f5f983eca6ebaf79f4a2d22be92611d2258119a0e991580fb3a1b17a077a4c3b3d
z5676ea99779197b6506841241ccfd74fb0f3e1b219dcbc1b5db451dd658ada1b42210330721bcc
z6af300af9f3488ab519767aefe9f1231a2e376c9fccba8a3e95e688b7de4574444d71388995b28
z4f6fb6f07caee763d77e6e3d33d6d386ab47471455db564d273c5169ed94d3452eecaa56c230c0
z3742ff7a9a1e66c82d6682f684581a6d6d28b2276cf2bd0ae137caae82bee808f7f4144d37672a
z5f2d671abe214ebbc448348aad13a86eb7757fa252866826e1a512684efb03876e9db1e0f2ec71
z478e1122d6d2ab4179c4bfc443740beae54faee7e3d098d1021298047e4c8a345d1acdbf28b209
za95ee050c4df174f3c35131b23f911a69e48f424afe7ca888b086c7212b02b4ac45f9537c896c4
zc1b5ea1e739ba04f0e29a7e49e4f9678ea3c0e2aef8d20f102dadbc52a87cfa8a3f16dd25914ff
z3f76eeb34d44417076c25033ae12d0bbedbcc65e9783125efaed2683e1d943fadaba5af6ed6e7d
z0b64d16a030152eaec2d45254ba2771618a1f0ea94e4e958a3cce545e45d50cfe4ceb3edf93797
z4f79b0727ad2ef9aa4d27c477a0683115989da4205f9e7734aa702ba585b3ca577708d938b2a38
zffc49688a7ddd34cfab2edfa588c3bd419167cef1a38bdbdcb0b3ee566aef0a3a66306ac877bf3
za47d712e48ddafdfba81a12f3c61f4ff0f16501accafc3ff17a6fefdc7ff23a1e8d35b93a4e224
z82c777b00d228cf3949ec3286085717af422c456ce4262ce80dda5a1dad2d130ddbd6c31e24af6
z6f4aee24c229330a313c6f3da3ff9cdd3578ddfcdc59e7548ccfb6e81ea67ba23a128b2479612c
z075aceff74b878f48d51454616b2dac1d5756f55d6b3a14600589a71f97f8763734e101f2c7937
zecd20f2d34d2a330f73f936dc26743b8a89ad1838171390d7384d94546af18073f1b9fca7ddf76
zce44b4df8dd96c7eb4ea800c46d09b444f4fe93bd6f17c79701fa80b22c59f5cc847edc8d2556b
z4730112a5b194adbdaa0e07f558bfe07c09d59c9ccd933852007acf92bade74ec3b1748386b3ac
z28e97d72c3ee1dea5e62d72729864529180057f7a4eeef592b80b6b5626e8b74abb481067abb9e
z443e14ec64f3ef9a56b45fb17889f699f3bfb0fb958012cb37f4df932e203b69dd7c4da4247d49
z46992374d02da5d5957ac8b3885203c79a7a783c6c22af259a65f52d523a55610552bec27c388b
za34f87c1734e6f75e7fee48a6c6daea3f61f24618f905ea61e012b5734515769ff086273e3d14c
z6371faf0467d6640e3565991041b01990be8963426557674c50b51f3f201fc4749f9cefe4727f4
ze11448bfbf83533226d0dd71fe44cf750d6e8bb585d192e4cdcce3f833086107504c803d7e8749
zc1e5db81a3ef896ab4205cb2aa590bf37fcef07af5f4204261c1345d09f8ac3d7745656079e115
z56e5acb06da46de91de180fef041c323d81a0a4008a89ca8303128036d670bc79f908fcfcc1de5
zbfd22c66b2f7599c3fd9541a22d6ce1b8f0bff12f7c9a5f057ac9930c4c59302aec904c1884345
zd286e059eecbe22dcabc8cef45ff7cc06f4134e8aed4bb1969be5566852fe207dfa9fd92eedc7c
zccef5e0c17a1777033fc688d0791ac22e70f0f593e1ee07dc70107221ec6693260d807e06caee7
za502713794da5bdb12863ac1d17e9814d182868e726ed0aaf1514ddb8381dd2ff610615e518cf0
z45fb37600d661209b31d895c1e463a5f1beb06c655908f5c41f47334e3a1fb0d05fa183e0fdb21
z8451133d2473d69362019fcc7b7b3679bd77f85c33f9885e8b8a857cc4dac820cc73d55ce7b876
zb3bcdd506159fd98c1cfcb8e9363ac603eafe1c9aaf63ba7333a3eaf7d8a9928acf1bd0606e9f6
z821367347b7002c7e4dbb86bc860f98ada9c1fc8686a48dd1e5017ae422c565de341cd4f42e43d
za908118578abd67126305be76afe294a1be3a817434841b754d9a534a8b69b653c83f0dd3a4f69
z852653effc347aaaa5e1719bb7a0ef3821a6dee576dc890e10dad10b8c46bdd979f14f639156bb
z9c436ea42bf624faecf88bb6e2a29f398b70171a6e1957ebbae769fda652d26edb63c3f3599261
z2c208a8ed897f65c41b07232db98d97be56b1df673639a1084d69b51d675ae7632a667a7db63ec
z257afcfd7c2f3bf3a07bb83b783d371bb423137157d4f701c9a830437b0466838a59f9600f23bd
z22abf940b1a9f8ffc8ff01d62252b216ab6c23ff293edf9635e2efb41a3c24af182dc965e9fe59
zd8c2faa22ff91da73823711d8f08f38c63b7a54780e34f4231d2d5c9326d01ed2c3304a3b38df1
z3d56c01a1f57b56e94dcc417b4e81b20442727d91da5675cad66571cc124573ca62336f536e42f
z62c1067d7d10d811ad880155b49757b276ed295d03b248c5f9bbe9e66f0db6cd4005f719cf18fa
zc97e931e39fce02009c03e10289b3d39bc8b6acd42d962076c9af3d815fb92f20cbcdc8bf76ba0
z18a7f707fccd8cc838f20a0651720572fd127f8335901a4ecf2ea414a4295a1ca0385cda837cfb
z45c0f768771bce7d34a549add0d6cbbc26628e50c23c4f6086d12caab49ee43cf613cc54c96680
zfc6122a3d3e5f1feff5f71569b503d37c0cc9e7d3970bed947842d7b38a967bb5ab3279e75c6f7
z6c4cd7c7e0b3bb5d930ef9068e9aa02e72d127d3e6ca41911f37ff675177254454753b08363dc6
z57c93c466c3250e6fb287a10e6d61f07f1d549854389f7126795b009ac937424dc4ad5eef32c3c
z4f4b5404ec42dedda558749174a480e2aefb7a40ca2689329e6b2b72f0c315d941283a9351d248
zc998e91800d318adb39bf1563a93f46a61eab4654c87284f788b8d24a69659bc1006f73a1a4e77
ze2c50021014361d8fa3b63872e5c3f4ce63df745c6267c77aabb391472be46f49545152a1b295d
zdb43169fed022063ba406c8fc8e8281d64e21b72b6cb708fa4c364e14d1a449f79fa6aa7f62ea9
z218367151fc861643fee2d7c8626eb8f218547543546a6f94ba54bcfdf833d9c783fcaf23f520d
z5bc9aacd8285825211ae7daf861b38c421bd2295d7dd71ee385646aefab63c54956fa84c79aebb
z3002426e9307749f8f2722e983c0fd07107ac72067f72ffc06f3d41aa2bb71b484bf8ab74ba07d
z3aaf7e39282bfb20a7324483f7e92ed8cccf25a2435e0755bf5400f2be53ee45672f52b1b34fa2
z203e3286592bbfa889bc25a2f0635b9cf60f0738e60da8bd96a755aab121cbfdda7a0591cb8a3a
zb1715205b4e35d8e70c1be6354f721e56edb1efd0e8606f689d4621a69a92ae8a69af8ce4522f0
z68b3c4e26f2a728ce657e1389c3d599b6bcc4da04dd87938a4f932288812f7cfecaa6c5227b237
z76a9a305f5882da235ae05cd049c7560c2c6586d7c7dcb5e488fdb478913cf8d2bbe1476ac4b80
z3c66e8f05b0fa8c40c0a53b3a0d9850d0faaace018acd0cef0404156ca36996668f692538c5c01
z9142895cb92aeeaf1e26587801e1a1b9e97252479091cce12d50d9ebc99a66ac69b6973ada74f7
z902b04a56d6bbfddfaf1ae04be8fba5bcb537ae51ca9c18f7cee1667b375fcbc975c08e6910e2a
zbef2294f28da5be22018556f00ddc0c7ba48b3a144f4befcb7392e4fef8da1e791eea887e3883e
z3c801253243e51ffd1074b56d34e1748ae5114b63f514a8cec253dba1638566f13f85cb86784fc
zb5324b013ed9c029df0d4a7d32e154b46109f7028cfca20f4854cff90509d92fd771a9f5cecd2b
z7d740b6b080f20bd8871c3d0023cfb8cb9e541beccbd8d55e06948358a93e37bdc6cb305fecd35
z8ed8631395594c8b5247b17034c13850e41110657c2b280f96fb0ae2da9802b49f65142441af05
z4f611d148c7a162afa8f2657cd6f0def0e6ff4f8a5814131e9cc391ac479c6ee7269d3716494eb
z8bcf403ab1cb2abcbafea1669d88dd35d755cdd627775e0bde470a557325d64e251651a370a957
z46c8faa20d4b7e076a32c9d3979836425762b91c3d455fb13381741da575cfdbe67120cfeefa3c
zbcaea580b4efb5cce66c0b3c5f18f3dccdeea34f370fd5792bf21bc285a75791f92152c64b2dab
z452db2523ebd70e95df1c8a94ca4adb7cf499e5802f1bb0fca21f86b7e1dff11be6caffe624df0
zb5550a331f0aa13d5ccbe27edf047d8e24e6048899e2802251c27449cbe12ffb50883c2bc365a3
z90001f0b5d2e61141d21b6b91c99506a4b64423fd393847ad10731a28627131a068a9f1899b396
z553b2c0bfd210b94c2a8019fad51c5f1cf2c3c0d0aa23c3e49baaa3f2a8c6b71646f2af01f5893
zd73adf46e7a4c6c9762cf60d00a195887e593bc302cac2959cb6a765765f11cfad23083212a70e
zbd4ac25f8ef39a5bad7044927145689ab1984f02775874429f66ac3aa581813236eae0cfd8f22c
z301a45445a3d8eb80b5d7436e9e60b9be336a1c6531a25cd82f0540efaed1e8040e107f972cda3
z3ac5be33abf0cec1b96caca4ec58bcd247cecf11755196f7c3185ee06a6e806ef7684bd14faec4
z558f38f0f653febdb64a61f172b6af2d447926176c64f090f5d164420e691aa4d0fcba5f9d37ac
zc7c99f655f21fad609b3d94f1fa7c1f7d84408b0ab8184390a446a7a9db732cb8c72c9692b50e7
z56dd773fe677e40d6d160e4f28ea8ee9179cb247b3aa29c77a2ee863416fc70aac452dcd7f6702
z1001bdcd64ee584b5609d80b8c357afdd495ee7d51394c2580c3444f09fd611514979ef5856979
z319ae5e9a3adbb4da2fe02a26f8a692843deeab9b3ebae705480da636b949a5a6257f751ec88f2
z528926c5317e9f7719d65879b34233690c7cbccecc14a88fede3f8542bdcba88499d9d4b6980d7
z126ae65c7fcb7ff5193343bfd0b43a590a03128ecf9f183bc9df76f9c5363b83991a25f390d914
z02341c49b092e6858071cc0a65afa7ebd79f3fbda2f9d22407794a8835e898129592a8eced76e7
zdd855a0544cfbfa4da5033f24d1722599b612fe6eea824d1ae59532abc164542c922ec13c2509c
zde45cb0318cb0326a5ff8841b50f78cff1d111eaef6bde46172949d84171fe578c03b1fa6d1870
z90dff31ec68030328e2f3097f1753c1b69a82a7a3adc94accff2de50b538248023376eba38f08f
zae032ccc10d238ef07795006db0e03f44559d3d61767d07ab64246032b82e0052c6c7c9182923d
z2a7048c34611779eb46f1010c7354c755f6408b12323568a4afc30ef4e79c3d682844418f30d41
z79b79f02f0a456b17048dc615e9378c4e056bcd4e10a9667174d56d9e3767f19046afabfe048c5
zd36f556f113db15c27cfb87e908325e9420cf0713d4d544f22f0d5acefd745f136ef36bb96a69e
z4f50466b36bd7ab4ebff912608612f9b0c9f741af4e40a8bdb670df70f15c562c44535221787f2
z52bc29e2347fb51c2aa7f53b28122666c428493ddd8d0500f76013aeb2bc02a5c97c3c11800fe0
zfa96348dc47c92279afecfa3719e9710eb1cb006452427d7cf0d3b541be32f0172e28a122facf9
z0fd1123af308e1307cc82c41f02e2b935dc0b78f5b70ed26f7ce26f9efc6018c446c341ff62e4e
z173a5661d458eef18a87b4f3c15bf938fa8413a0981ec59f06ba25c16c2e76bcc0b9f4c511fdd6
za8255c01992d815284f1dedc74dba35848f195d9e459a2a15e8ab8d51b7c96ac896115b544f5fd
zd813a5ba7142976a32304dd14839fc3ad6377efbdb0192f763d90e0d5a8645eb13cb260716e98a
z70b77fc2593e342fdbc43b88a42c1d81c191493d623e794af74bcce0448c4ddb09b3abb4376a58
z117ddac89f5ded870e6755e31d23d6a4706f7f8895ba0ccd0e7de6bdb88f002127c9d69e9a0803
z8b95036e662ecebc78aba628b89c6b762566b8202ed656604bea99e2689ad3d3fd7e3ceb5bd960
zeb4e0c0fc99a7022f6b5835395dbbf7093b65665ea3feb6e5fc37fbb3bed7d7eb232edb71ccbf1
z576785b7379dcf5d6c1c2ac8b33a1b2b3e4e812e598e146768d226f36df8c750ffd515faeb5a8e
z519469528bb5e2e808ceb5942ff5e5ade12f2559e05b73b163438ea6525c63d3939e4092b043a7
z1ed93b63a428b617e5dd1409924bac532f7fd958ee5d4cdad9c74be95028a8e25af7cbb55ff503
z98cfd01a79bcc8c222fc7fdbab569b5755d0d8ba7a18e2c525bd449a4a9e3404d38cc1722f048a
ze01bcb6e450d1c190127ec0d826c6016a059eda7e90ff27513040e2465cfb88535ca7a9f237278
z3034edf514629a3cb45e3baa2550eef5d208c905790a6190bff8734c846c0733e061468876c47b
ze60eeec8943ae7c9cca1f37c85f41c7b4a27831c349bdf4caec95a3f3897e53067d012d23dd9d8
zb82692942ce24229a9b3fb0dd371a9b02c3f3a5a67e6361f03c2786642e16499a321a2767d6b32
z9b8ca045703da4981ce6196ea938fe79fc7f4864469ed6b08ef273c4ad09f9b2868646e0e2076f
za96f90b0081599851348a825e71f35889676a139110d2eefb57a4ebbafce60833d1bb7294266b9
z43f9a365281e1ce0cffd6244f78e1ca14dbf7862538b0a9c4d2f32ae6b72bf061314fc05700899
z7a51b53f1741742ae60700362b90f7014c2ee6074ccaeced702a02fccb4ed4022b7b5be692b3de
za5c74ed0cf62c48a053645b12457fd950b00ab797dbb5ec07e45159d5c787c40a9821e31b032a5
z81f8b2e925adf439ce512f0d4a59225fe8a18d3722d74d9f36d997cd00c638f696719011851f9e
zeefb1bb6940d5f79f881d9fdfaa52145cab9ad454f33340f722c569ad6519dd2e31d0bcfe937eb
z9d7a5bb54e6a84abd5c55c692108aa7f8085b16858de3aaf423033d9e6f396be37c01b126fc2c2
za58c55fb79bc6e9673c57e99f15988bbd3d249bd57bcfeca63fb4ce76821bc4a483420d2f9473e
zb429ab2d1cbf1e0603c492d8871c0ed20c4002671a50f8de78b931ec4e718721e1a37ac9e0018d
z08faa83d652c34ce122379075b4843cd45be301f8e48ef16aec4119bc884c47acdb8c2cb73447f
zca3437382a65345d687cad1278e4fdd17164ff556e0c6115bc10d0e89575ccb9586467b9afb95e
zfb8ccebad8543d1a5c99dcd7029b4f361a7cabcd211949ad49755f2cfb1fd5b99e2e7bdf031cdb
za9af540a432e6df232f77072b5a1fce8c699b3c4753350e0759283de4ccc291098442634a28329
z4191b93774c6de57a5956aeb0cb50088e5c3339421858f86cdb7a133314fb2a908eae52d86d459
zc9804cefbd50760683432c6c3686f3bd9067b2fce8c4edbf11706aaf248fcda0038ef5368682b0
z22f70cba78516787e34ab11b78bfc1dd633a3acb774a54e050cf8b44551abcc513848d0309072d
z250037b6f16c11e118678bf384170d74524192945171c5c816940c8d04acf3df08b98cee014b9e
zf920b35aed3da9f66fc1b0c41257e6366017297ea95e0f2f0a21a07cff418a9ddeba06544644d0
zf2d5484458965ea1ee9d6bdcfe722fc6a6bdaffe3cbb8099f53e791122152fb132a01afa1fb07d
z0364171b606a333627b9444fdbeb7137319e03ca8fe87a15e0d90e7fc2169d7c4abfc92d422b76
z6c60aec025321ff80d94b9843ad907a2a648ee3abc4440749d66ffb1a11bb0536d55170543a45a
z4bf760a60c1920d8b9c0771a9433744cdd46524f6cd68f4588783cdd5d5b036e306830e28bb5e1
z2f1603a110b8ab5cb6ef976b283ce83b6c2515ff5ac3ac32986f9af59a83083346965207ce7925
zed9610d4df5ba36a0ddb0ec6dc1113014156ce40c0f68d950f7d21a494b31abd618cc435ea1b57
zacc1dc221a8b1d7e5a2ef1bb0fcd8563f998574947527c1a89a7fa7412cd86af5e374c07a4341f
zb79a0f355c86166860d7cd2baecc28542079e4bb7ae9c74ed4dc9b8497d7aa1043a7ed4da3924b
z1dc0eaec07f19d43499c79ca4564ad46813e30a537b9c020f1bd0109991f89695051dcf9cf5854
z811f5a711089e9f4f3549ea52ac361725e306380368fd2c3e1e8adc7a70e836b1bc6380955cf23
z5da64ddc4ec6736fb688e2362993e7997a8750b72f2cd5378622b2e1ef9149cea5bd7b03e86d19
zd218a7279cdf2b877989c1f7ac9629ca466b49bd40f11bd1e18331c4cecf8bee653576d506f9f7
zbcdb406efc6baef41f0ab47d8d93b99a24af17343e32adabdf3931a9c741e08b7dd212afe8f0db
z5ee68a2714218f3e051e04b8b135377f3e6575862bc14e936310b7bc282bb5a7504a6ccc26b415
za4c84fab6581e59e065a961c786fad0a54b3d69c8df88bd02e12a21b9f3676d5aa9e852df07e01
z6c5fa1f7859c3ec2fa1c1d305e60b38520eabe9ca7f179e4b65246bcfc389f237bcfbc56b74d3b
z5f8ac932f3bd1dc5d0a3661d4c59ed0b86d87043f1d33553c38b2fe425381f821a636b461e5a71
z6a795a500c0d008866066efac5524e36c5fcbd78e0b102cc47dcf2ee596035d4cef0753e2369b2
z93ab9919a6ab0d88e1e46d83a5de7d8417d43ebf0e2b37540cb95d7c95703d15d1d51f9571f0e7
z996394a9cadbe3a92987014db6b4217dcf4be8ae1b77a0cdbc0e0e8be6602945544fb2157a9ea9
z6f72c25474767b8056cb6af1efe0aedf17bd5d04be80180c56e282388808197518dd552e83fc1b
z75c51b2d8c5c5c93da70cba652660a75c16061a890ce6ceaa2c233ffe4a300ef56829e872716c6
z6b0ef5fc49290f6272da9e45c96a6179f4af06d13f4af83d8e6ae263eaf69d29afe748c8de8833
z08c50633b3de2acbdbfbb1e77b500467343d46c56f964b3daa8b91a6d996a866af0de71b5ff105
z41d4cc5daada0f98c41d51d94337eedb5f2638fb663c0e608cff00f2b4c14630189e2d21f6775f
z6cc3ca4c330973ea0c41990684dff322c99cd84625345342c9bdee3920385c9a52c80b7cd808f1
z62bbe429904b8879eca0ee5cd0a98773cedf86035faeeaa8c5a1082c501bda737ad05b318de63a
z3d224b053e81d992e4d6d9bd1d88314bb59dacac2391e6ad2036f5fd2f6dfc6501e89983bc0049
z5937c05c33c390f83a2d4a8470291d00c42c1f4e3791d0809af3d41837c6d43ec5d2c96dccdd29
z66f2a5c10c87e9fd1adb8e3f07fcf39215c6d5769c95bd794735b709b2503393720655817db4ec
z3fc0f0327e49588a23cb76082e0fb9fa7ab6085f397c1fcbb3528f718d4a60645da2a54bb192c9
zb46eb9afe90d1d2a7fb150e3b8c284c129add53a6f99ff6ffe99f389a5c60fe163be1a859b8c88
ze91a23337edf8246b3d035fb8e1123c6221b349cdb40d7617e878f0d705ee8316c1dc204d98ee5
z505e29aac9e07b438dd1853ea214e34275d404efbdb0166aca7bbba0b0dbb90e4b5d014f6831ff
z774779f88fb676f661adeb548f84f0e5d4c4ef2e4d684b431444b51025ed0fc1805661e4eb255c
z21aa3bffdce98de076637c1bc0ac05ee70e5a7caf5ed769b1417805d62d4a1ae80a071c57148c0
zb8ddf7a661aca1374d307c620491d41d771a9d8a350588a6b7926eb6454f1b66b4b0ea1413cbff
z3561dc60e815216389622656fa1cff1b49881d3902b4efe8dd18c1deeeb7067595327ddefe8c88
zf4328f72d4f91d448bd03eada596091bdbe5661beba95bdf5a5d80aa61d89f43106b0bfc04dde8
zf93cd5a484e489b9172402ab565fcff724c4e02ca2af5493ed52120ea704a90563aa938eb3ae9b
z2f0479e6424f79122512319f7ba8fa2e7e06538edc47b941255f7637afecbb87c8e14d8830ade9
zee50ebd6cf147ebf0dffbac422c5f15b725177a4fc03d6b0fb02abc35f59f6d20d33a9aa09828e
zf97b6d2a2234f94f2f9c48648ca5dfa94688986820e7876c261878fd7631edb9c8d56af3c75c5f
z1ba6e72cf0e00d9ddfc2e3b61c553cea3529517d3d972b77c3ac819518a80da9385c315dae7928
z0ddbe658d438e9ee6559ff3a76b1e5cedc78bd8037a16fcf37e8c300112eff3dad1a5a974f06f9
z48ed22c2e2474fa00a7409877e703b832a4c018448ca8d58ef6620b61ffd8734277e1cf2aec0d0
z4f1e559402279ebf26cc3948872bf6dafd4b104ec04b1c952beebb21d467982be74acd25332a68
zbcd096f96e79ee359185b12dafae022199c4e133a359e940b9dc8cc523f521de91ea0a46799264
zed765a48e633d89d7df495f3360bd07eac166aa9a8eee3355ca4f93e6500fa1309e69ca7dbe59e
z1960411c4737a0cd475f342f923388c8e6f5c2334fe10deaa211b756d682ff3880941e13cc8bb1
zb2b372684bc21b307c47386a0a25a30bb1f4411484f8520007268ccc7933fb02e17fd10735c366
z78015d262a519f816d64e583721656b686e494ec97ad5d95ff567e57d7147ba09e0320e48c751e
z9ed71d24b7acfd11b53c1e02f073fbb689d756d5fd3a5db0c91bd78bcbcc3f195e48f5dc0c7a97
z56c0b90589ef3762735c41fca4cbee85445a3d7e9c6a9dac55a5b1d0b41a35317f3a366eb2b1b4
ze2422332a68a8503bbd687e8b3fbc5af54fe1246a93e87453bb9986b2769993219edb8a606924f
z857cdb70d4beee296ef2a492609cd87875a4fe6362e9e5d5695213bf6a42e12f22ef15623f3a8f
z951447228b8e682ca6dcef8d38bbb54f3566366d4b1d65d57ca8195c5db775eb95fd1ecf5b2f2b
z76e9e755a86d53d4a9431ce574780d074a961c17af44af50ef4f7d2e3f445e25c628a2b76e1562
z883d1cb7087a475e75e6c1340d4d5f60be92e16da754a29064d99d55489b2622e7b5fe89a3c18e
z1b40158d9fd629c70d57e7356bf3987bce34c9d99afc5b414dca7bb4fb67878c788d56241c2e1b
z31dd4b403159c13c8d6544d5fea294ef3f9aa7eab08043d3ec8876904c67e289a98951d1fad697
ze42e0c52920b6d3a427c6f1c70027ea77a9a4b87740532ff6352e29bbb4fc31caf90445403272f
z121531295deba47569742a3ed4bbfe89233eea0b373fc7035330709aa72d1b3ff34be930fa4168
z874465d980593dfb5a0ad40d06553b93f57530108ac5443085d261af65a28b28ef033283f7e59b
z2305f02e227be5f515ef4d5d976f50d626f840347ca97482aa3b9a7f4b3088946d4e4e792b7133
z6f682a8f5afa526e6ab3003f7a5aae5992d06847a9cd27448c664ed6875788da15776ebd47c35f
z61255113eb7ec8cb96db88345be08a19997e12d267dec8f03519f3fa0f060f882570969d907f04
zcf3f286b31b96fcf853293eca90b5c9bfec7d7a81d833e50642c24e3c1a9a728da01afe112192a
zc2fa4c767322230ad8585eb87497bb2c0edf8acd88458cad7df0270f0eba95f850e83a41728ab2
z72d27fe4d5faeda1487557866c90dae4efb6fc95b6289fa22b280774ad0b0947fd27dc7cf90189
zf48ba3f4a70f975cd2e39ebe99777b705dee4cd6d19c4746d88d0e34daf719370845942a6dcfce
z09974fce0e84a2a9a77ac5ad774c23638afa38c8b56f6dcc3528f7d6c735673a0bd5e8cb48a0c2
z1b2f83455535c7764b4d907dea4edde66b0b60fcb93e787a9ff55a21945f020929b5d526a0256a
zf4a6376ba1206a42b979fef4ff20dee4969f094e44de1f286c55bef3ce084beaca2148411eb9a7
za684d08db53b94c33cebfa06cd00622efacb69367d151427425010d67b13f26870633511f21bd3
zf64d650d29ac7b616a9e947963cfe9dc7ffae1d0338c5fcb2e87eaee278febffb915af769ae600
zf386aa6ddee38c67847f514c86c121cf4a0804514b88a41fb46e79829474358727013ab3b8ef39
z715a50d58b99abb80dbc34c219ba516220aa8c8e3bbe2503fa5faa8879af6729852d182ae7e7e2
z570ddb856782fc24840209f68f79c6d4af3852f500fe8efb8662f636e6efdedd9c5105ad7b7399
zb2bb5aa1360c156b254ea1d4b66cef84669f4816e40b98b33579bdbdf3a45634d7608d717f3336
z14e0cc22620aaeae0719f7a76f2a93b4fd6f7b83c6781cc0297a98b6d1f19039eb8e524fb444cb
zb249f406943293aedd8a5210cd9aea478608560ed9e3d2addf9d6513a15e16113e80c1de15bb60
z770e9d1400221cf25f8f13e6d30207f505b5458cd397f8234b130c791785c533f44ca9aa6efb76
z2693803e8f9aa9ca302a419fb642790d384a4228897e7e1356330b7b4a8c29927a071f27eda2f7
z515bd3099191ba03a10dbc7e88d1a11de89cd0769aaa9d7c1d4d5e9d8b55e2f7097a6feac6809f
zb917928cb915d7b6db132245ce903d6fb4057a896b221660b85a1e30a6c674d97fdccc6e633cb6
zff1002827e7ab7f7301a96b8a6b3a30610ad91a1e827848090e509551018169682bb033a8c4a7e
z210314f137ad7a60c405ec35c290caabc3730bc56f76d0a73abca4fbd8be937162b4039e4f82c2
zbb8eca3158d38e3c74ab2ac43346bd40e860da2325044e1dbaf3d3c855d89f747cf3bb729c3a2b
zb3c791a724ef14e43d815f0b87065a4d8701af38e5d3f94b25d594db32a43e8c62028d0e0a6359
zb1bee1aff90a195dbd99924d81967cf9fac0f84aebe6ff47a3c4d9560d6ca4393819c615c0c937
za46850890bd44f837a667c1bb40e8936bedf14b6fb0c0e80591e459236a3974da7dae3a6bde8d3
zb535de46dba3ea10c5a75b2223ccee0d7083175c998f4bbe44940bb09dbc25301a74620df6acf3
zc7bf8edf88b89c0cd71ce2dd5e351fa2eb7f839be65293b9ede71e3c148115986dc64f2ea4004d
z42c3cf043f56101bb5ca3ca8753ae77c076a9c88d40ef033ed7751a92f90e14ea282080f82b849
z193bbd023d9a65472a652860265ee571ace704285cb0bf2fd099e9441a5c982656ccbc51160255
z3a51ba87d373e552a8940dd350514f6611d0e22792d449ea4c84b135a00fad4d34b01fbe26787e
z1c45ab51dcdc7fd28772331a3cf66c3b9dd4e94d98743df9d31fcacda50e4254fdb630f8ab669d
z4bd3a33a83e0226c83ebd25c09b0922ed5fdea5803030e12592137062e18fa415d6d9816f41ce6
zc56cea0ab015efe1e57a283917bdb338a57d80d52ddf330519f784a6352c0470c5ffcf13b4ce06
z0b825c29e1754e383d8e51a46a3dbe1be33acfa176e29f0edf70cd0da1c5c2468a7a94c97f7d3b
z162171dd2268d970da2abf909bc99e6b641e3326b8c41c9c211d72979404bdf65bbe578c683d98
z5b6c7dd02b1e19392189e58f5fc8494a7c2c82f4b35a50c942eeadbbe1f0c56b90c2b8397580c5
z27c7a0c860e9f7e06dfe5bc0f0088d4b461c0cb8125ad3716edcb0de9c3c0b1b6d4de17ff11720
z91716a2ab93d08fecc74259402c407be78193df5bb6dfcc12cfb378091094ce983eb638f0dcb14
z13d82669262081ab01eee3b1562d536ae81ad5e12d3407645c23034c6ce77bfe2083cfe8832fbf
z2f4bd1610986d5a692e40c5edec929dc6a7f13a25167fd7b0dbdda48c7d091cac7fedf4cce58f2
z55428c36a49347b427ba70020fd346fb3c45724e5901561627d20ea24efae5c21da6bf6f23b1fb
zb882d3d3e321feab61c61012ba636ae5146bf80ce59cb55486c88650c694e04431108bcbc501c2
zefda63d11fa1b11ffd3c583dc79f18fdd66c84a7eee214cafcd38f0f02fd1b55bda974414f44a5
zb789b08746de75dd39ee2026586332fd712ed3fc793bf92caac6e9879b081e08d16ad45dc3533d
z383efe5d2ec3d606c06df81be277fdfbe6775b4f1a19b2347f74dcceccf4f0172ed38029f89162
ze3b1c9203d77d6e358cb19953edf5c00075745fd87f368df73313a4a161a6c08b2bc31a1d964c0
z3498193d7f854d94b80d63b8f5f594bcc71bac8dd051f7bbf212ddbca2ef05bb8bff93207d97bc
z5aae2c2ac2adf531e5b983bc68d54daa8c1b698af638f5e5eb928f313ca85fb7bdd898fa141d53
z0fa176a69c7288991446576b328c3c729f4eae025a28057d08432c6dea31770e98259c2d03a5eb
z4fd15d50923e967d9f566f785e865a381bd677e5ccf99138fc6c6f623845560d4d7e3cfe5e7b1d
z9299f788ee74b66ea0c1ed6f73909f3e8ebfa81f13d1da0c39837c10295eabefb42a5259bbdef6
z5d03be5a7f0e8d1c89e576a179bf1c45816c0aaf8ac86739166803482fa3c0633a7be4a42f658a
z251a39492169f919201dde58fb955567efd3638b29ceedf4a12f4d283cc7d27970c5e7a5fd937b
zcecd71793791f63fce5618ad62846c02765c994c06350ce69635e4bcc64f46f77f07d97a4ad8c7
z4bc7e20a74fbea7a179e4858391a0e97b336dfff42c56f363f97d8ec4a304e45b819840277d85a
z1b00abb1d1bb3b7c13c69dfca4807c6e9c4deee846767c9ef61f320e2c58208ae8cedd38937102
zc38d1b5a47dc01d132d98e9dffd6a6b405a2478110ea21996c93eded8ac73be783efe65e41e22f
zf8dc8dbb1f9e24816a89becf8b572e77ab1e9826a0be08c59a11c2ebb324eb6d91120dd44d625e
z115dbe635a951d1ca5c8751263921e55cc41a75242a081bb7491542ae54ccce4adf1de64e3695a
z12ec30bfa41ad34552c4dd59c953d4736d15c1ed708044db99c2af9a542e865ee5b1ffa7a29e6f
zbffe31a1378de38d0e48a6ce2a605b982ae668826758175702f75bbcf1d59b2f20fdfca01c4c61
zaa685e5afce51a1b64206d672efccef7a53847404155cdaca4e80a17a70b1c4b56e295161a601a
z5ded53c094b87ae10338db37efaa34f8976485f17e34cd4fb12cb05bd5ed2eb8d5e9e0fc40b18d
z67114d30ad5adecf99bdc3387fb5b4088a6601960f39e56ca0306a75c9f2d75af4784d93c169c3
zf385cb16d63b6e63b37b7c988230862b8f61c4ce525056eb208a485b1947c1848932937fe2439e
z63014a785ffd60231c80a857089bba73de35ef4cd75c4c311da881cc1f297d1289c2c46d41f8e8
z13af63ed5d9818e28c4208437c62b665f819c0b04df5a95cab34cdc660068189474e8a768b025a
z00c2269526baa688af30dcd739d90bc359f9a1dcaec0ed6f51e26ccb956b23bd058167e951cf08
z4666985bb53206f0cb805849ed1038336d23aa36f02c4cc04f2ab70ea2a3227a72356ff4271bbc
za51a47742cd2bde40c7b64e0884b0306060c6f3d5185fddd9230f00122a0ff2f10d62bdad7310e
z3d8c37a43b306d0bda3fab5a2fe035455eb571a41960d50d54d75c91c15376b665aee83c7b84bf
zfb6fab914ff1a6e9e0e4bc9a68b4665dddf57ec6761c498ee89b399c96f979ded248771dcd3023
z09a8633a324e1b2661ec30246924b756a287518f3ec875bd0e932c17773cc25c36f5fe54846193
zac3d3eee4058aa613f88e522761070d025440742fb17848a5744ed5d8711fdc64e6738ae63ca29
z0cf8be81945560560b5afd9779ff607d2247dc6a7d0ce53a62b78b59fb70f4622654f3bcaed340
z45830c07f79d75cb4e43fff3c1178625090b79ce5eb6632e176fe510366e063a1bb07f0951bcde
zd08fa62a8c4df29fd3bbf3d810e70e6b83c4f0ad717eb3255f94309f1c131e91104e2803861498
z876a994bdcbeef605029950265f9e87a8b7815b22054986aaf2ca260e368c5f0b18b63880717f2
z6ce97de256aaa8610756583f66d4fdd4b6373caeec9b02cf1ed3cc256b4ee8929bf9a34fd5c99d
ze5104205139ca6a662a7d7a2a508e3b843b88843e834ff455b5a6dd0a4ad21b7dcab506be8b8e3
z23aa3e582de7321e2d0c94d34ad1fd4c73c9e2b15a6a7149d03a833a8d6eb92f3bdf968b447b4c
z55f4e219784e67335daeb52491ab5ae3c35c00ca8e5db4a5958e3b487e4b19d8852b5b38e4d282
z459c66169553434a68aa25c042a1fd2f70fc19e83bf86eee6878106f0d531c6d448fdd328410d3
z52e80bcac3247c27ccde87ee15c009cf97aeb481a3df43e6367f5e3b67d0cee724fdba70c6dbf3
z7c980cbd4348db0e8e30555abdc57113684215a5873edff635eacdf60f7c4176b4836c1ebad957
z01590fbb4f0c07d34dde7a03b9d24cbfaccc89d831cd7cf4b04bed21c71c3e5a31c2db7902ef5d
zba164155284b8b02269ae1a7c7ac62eeaed4f822f3b72ad82caf40bba46833f3e8a1ae1ff287db
z66e0bf48fd05e709d8c166a46b4cfbe9b3a3fd4f2b2e44fcdc512b30c5ec9faa22e4f0cc71bbbc
zdea9043dc1efd9fea254749d97c0020cef0d49cbf7f44e80928ca6d295ee4b6985c70008ca8e6d
z05c99088e26da13dc15f2cd3fd5658279c0b2be4e849887d5f7cbec5984be3a15094adc5917715
za69a8f7b01c1e0e8340b12183dac0cc7c75f72a79ddc1b223f120451f4d8554bb2b7eaa0a037e7
z36a3bf8bc5949f0ff47b0580f2ab7c84f69955d9ab2b8668a99f5f0aa12eb86f6c33ced9345370
zabfeae3074f0459fc264c9228283177cd70e5ab6005cf57709230fba9121e9c921bac161a7ef97
zf6fd8e3d2103cd85d5c0853f9cb08a51d50542ea0913ee79b1ed85a305c4abc4b88b873f8c4a4b
z4038dd16a2a9008ffa29644784c6ed4bbf954fc76e14ab375d4ef7bebf5e4108ac60a3b5253b35
zd134771af18e5799514fe7a6ac7944c5d615081d80dca1f3568092f0124f25b2136be29eb77819
z54716ca7415f4f2b7d3bb6e7c7a485369fa3c2da1f9cf28cdedef587b9e1d5bcffc372df7ed9b2
z96ed6488df59d246b19115d4ff3072a43f949ba36ec629e4235b51fa19b9ac88722d1bb402c71d
zbc7a7117f7af30212352673c0769143bef0974ff4f95dc60907a86b67a348472b2ba0af8a776f5
z4fe177826c7d5c78685a74c296db84037b430e8a3c6312c1d581153c965af3a3ee0c1c7fb5b6d3
zfc96d054ade7b550a147594d905a8117883bac0274f3513c75e3605c535d5014b712a79ea6ce24
zd0cd8ae7ba6bd9b628a83fc57a8b1d5b972e5fe50c7d7259f13fb6529602be2b84a0a7dc10e9fe
zed6eab6f9912739bcdc7fac829a0a2bb370e786c1ed873a5850c3c350c0f7fd5942f365d997a42
z87d1a016ee902f251d396b4476394f7fc7ff89d9b261a4b0736fe951dd3596adee166394be558f
z9e90ba848f3ad76f9e3995679f276ff64525af3605cc181cd7489401ab105dc58a0586a1c643aa
zd438191ff2588fe52f338327653b4ea0290d34f28e6b05b73e46056644935f4f7fc9b47ca7e49b
z8d33144e6eec24f846db491174e0fc801d08c6d3b514fd7393083cf5d987c353a13b1375bbd0de
zce354fcc903b2bdc1c18436113f6010f0bf921186184c630f0fb50a986754cf87560750be50a37
zed43607a7f5266a68dfaec438158eb464f276b81555e438c9a613421f456b9949c1b13252076e4
z51933a4fba0783404fb9ba0762c5e9f617282876ea92a6ffaf3496f7a9b448f3b00108eefde96a
zc44542af3037e97dfba91b534b762fbb325d456f0e84a4b0b7c2a1c98fbfb8146ee6d116ee8d38
z151b6cff4a71d5bd132382bddc57af6ab5872c81724de309deb9a5446bb6bfaf38498b638eca14
zd6890a92f3a060225ade86d48353398a63d6a8e49f84415c184da16e8878b87c695b39f3457022
zab6c1393cd6d0c60162ff757bdece1bae2861f54e39f4d93bdd37e31da1150489abbe5530f4c95
ze1053f38be2d3a0934b3eddda46d10a3ceb00bc988c82f7f9f97ffcb5560e0a26e58b4c3b033ec
zc08fa379f2141b3a00dea72dfeccd2338f6eb76b15fa2212b915e17e5e7e825080fd2ea1a633a9
zd155e7a13d5ba22dc6fa2913f66f9caab062d754c1f190f7274a048253d45ffa1318ba53c41add
z2d2b623718ad7cb65b24224a2e320065760f7acca2ae84c88084dfc9e140d8283336733e8bab2a
zfe2d54adda2125c19bf8334cc74ac7c15059ae8b4580026f86c0d4d49792d023e30271e187290d
z15813e3a944e2a7fe2a9acac85c5bacec7ba4b6f70ae1a2b20c46a202ff53e70c3426e0e68a5b5
zf7985827f8f7ebba775a299daea216018e6e99899101a5a53921dab2ea3c85bd71f4af4409ecf3
zcab70e9d1cf265efad34cc74329a1a1c5ab01d761bd57b8dcb3099599db6be6549dbd0b3fe2b91
ze327d6b5c3b5f8f5041f0b2bc492dcb1f2eea70b6e972203004919e3a9789c19f9067cdccdf004
zd5af7e6fc41604c052cef3089f1683bfce60a0d15864ce4982b4d3089be860b9e602c85ea0235f
zfe0c92c6912ea52267cfddbfd04aa825c92bdfeb06b750ab12d78619f0553fae0da6b9c3627b27
z501c2a23d099c791837e76b6f63d0ed47ceae92ad05d7021667ccc32165f663a6484139a288aa1
z76ffda212eba8c26e459cdf6d8b8f8083781fcdd8ac636f7fcd80c1d687934eff30260159e9407
ze51021dd15476d01624f0232abb4030a8637568d9fa5b907aac5ffe0270896e517c30d13312eb6
zf589e3734b9eb9b68dbc2334148ae577835015bbfb0ee42bb78945f787cd2822cd10253f9fb471
z371d9d1fd06f8e95b0b59acffc13934b1f486f4233fdbe551ab836375596c37a778842b4278570
z405609d9a1fd2eef1399b09b4d10aeef5eb61dfc8854dad99af90f41194743b7876a5ba5124d8c
zc79acd4f21e08ed681dd4a8624a50fe2a3e658c91c3502d7b5995cdfb9930b99b577057a6c79ae
z5f8c117beff4bceed8444b0335959803a06d63345d451d71b0dc31a872bffcf2c43d59fe617806
z6a74ea309d90f4d67f5c55a940a49bb73fe6b00fde524e071a529c6901065d524fab4b7dca297a
z8d3f920863eb7588ea289f2a20c507cbed2069d42cf195c9d71e46471ac3c21a085d26896357b8
zdaeedc10e30481a93e1449a59573c929a2007a770c5e9845e0eeae3435774adfc78c103bb9097e
za6b3934884245a3fdb2cd3bc9d39e46fd8e1e6a57e838930b6044a5ce4eeaa4b481b0d0b6fcc34
z536f9ea979ee73df1239353a5e5c1cf240e4a8ae869f8aac767b94386510d550596521be0272cd
z2519a3916f0ff792cbfefec42c947212b6a0abab8f6070738deeef2a8e8f8d9edeb2b2d6ee9970
z4c31a321c2b8e6f02695f7ca7ecb3e27b33e7dba4678c13a5f16246c7f2848dd02f371eb2bda4d
z783a2380a0a5c0b15c60a50c94b4e316291c2ce96e657aea8b88e1e016a1ed547e00613340b4d3
z57f5b70f9c4f48a338f56e09a89ce6cd90f458aae807aa44b2962d4362ac56778565928950cbb8
zc6bb195d45073cf69b02286aefaffa0aed570cb423e0a63fc3f4f779950b975fd40d32f32fd3cf
z133307e3c05b8f7c70f29d7d87056942f672f1b60b5ae1169b9372727acb17e019608f998b961f
ze4175d8fcb40ce93ee52822c2bce33c201bf3d22cc417d8d3eb504f6c407da00ee8f0fefbcaa5f
z0380d6365a027458593b218bfb3be34018cdb22712ed68449bbdd042c82c056ebd9e53b84d85c6
zfed7a170dad9ded95da4c73bf54619af7b5e1cb53d32acd12eb36176f344fffd5ba764aa425b44
z80b2e6b36d2f107abd83b187049f0b66e95f7ab0ef06292b4590bab38fa376733c83da67056b69
z9705479297b4d49640a835b07b750d9ce5d6dcb57f0ec5d4c14a222aa12a4012b9a02d08455636
zb7ac275f17a802e8a01ae3bd337230ba4d5768afe7955ad41d0302f4e77f72a6f49b0a0ef812fa
z8def55f838daaf1400a9dd5cbb88fa4364f670d81d92a36a915c6235d3b8c7d72979ea37da22c1
z8c283dc0121dcac55a88bcceceec2d0ab7c3eda00d1c5aecb7e90f0b181aeb076f5ae24a3751b4
zdeceaa9479642db47e09a3fb12fb20cfe6b587e50f217a0f2d98e1cd847f6eeaaf4cbf99356d9c
z92696a68d37f82eb085d0799944ee648231f6cf1f24692fbe7d58c90ea8e13e4e56208fc6fe338
zc71ca45c48a1a9b5911b1ef6292e5725ad1a6be785d39966f25f8b23e464f1ac5cd6fd99836d05
z4ab40f35972a94672b1e2f8aee2878815e6f528b291e1bcefebafed5fe0bd060b2443be2c323ab
za5749ed53d9096090e32ff8602ba3d95f3d8d10c62f229f5968e125bc6aa92cdafeff6a1dff867
zfe7903732512f8b5265e7407319abf5b9fefec703190b2878d97eb0c78e5d86820231a3157d11f
zd01e49066f44f6040cbca5fe50c9ba453dabb10b5b8386cf6f703b9346a2b72583aa7d37d13670
ze3e37d9b40e3febb0382d1c076bb4bba54fb581579da4d3d177bd25a77bf89fdd703b052381874
z42a3e4c88dff34acaefd2eee57ebe5e9d15e20dc24b5166651aa1ec00992d9c27109d63bc02f3d
zad59fcf24be4d8b6212c4bf2a3469b23da45c57f51b4b918c61e7a67ade392024ac9ab167e8822
zf3450c087e689dd2067be651d02fb5c206cf27c5bfc27b45615741911c52d4bcf1b28710a941fa
zd0a786f9f226c445c10a455911d9905b94a9177afd6cdbb9b20c870c1167055bb5c51269f85fbd
z0a65ac15eb1c11a7a8453ef1b8adb857a511b65bd0cac4f08e3757d83d6e0b153fb306328ef76e
z759cc132b79be9e551771057ff2fdbd45abdc5c61f8b0ec6cbb373dbac6ed2f3226654a837abce
zdace6001caef4b0358fe6e1152a51b32ecc02b6a9f535ec21e4d1320d93481d8b4b97028b968ad
zbdf6b8452887a5b6aa0bcfeff5e365ac12ca82345c2fde557b9f7fcb191d70038d5c0f5dff7d6b
z64dfb9abfe5889853375d4ef3b3e5d7dbb25aebe69c136b5f38db7eccce8e69ca556a4bdeac0c7
zc28d2816a124b79f446c52f9d9055acb9e475b5aa43964025ae55c1a64ff574f93b7ffd4ea21db
z641a2533bc952e062ce2ba1e404f27a767b6c9a8679d53e26f0bb092138a33fb520c7b7edf1849
z9342ccfc88896ac3a754b40a2f1008e7d4cc891652bcddf015158027f8358b70d5761e1d487d7c
z7dfae0eac353e7e7fb1f9e3de7e2d79068620885e01e262c1b18bfb6d1e8569480076d5fbb5a75
z412209aa292887694bb2e0d1335fbc86794fb82f75d3c6f69299046c1b189f6227e4291e7eab61
z11af1c58d48000cc5245541262c94f59a4054ccd9beb0737c2f831003b631c8df8b03f61303411
z8163a701c3c5823177959e5ae1abe4c5836aa5dbb592397cfc9c07f7deaa2ed43218932636c5c0
zcc925a46b2896cf004dd7866a6574fffc9320465e14bd7df1ff7f23216391d6e87ffae87e62645
za71a89054086354fba4156665a5ba87294b79730c36acf87b62bdd70d674e907e63fae13bedc20
z1dfcb2eeaa0ecb68100417772c04677197900e0bce981a3f4feaad45114bd85cf1198022216aa1
zb9eb8060401758aa8a28ea0228e322762dacd6a9a51e64c00b3cc7fd40af08504576cf89672ae9
z85e15d6367aa72ddd50c528eda271977e68c16a42143a3da90f070e96c979aa7b8f1f9ee71c78f
z6a6d7a908aeeb80e03f1ebc1ed52be535992e394d0e6bbf9a201375f94a02d1b315e20055161bb
z0ffb38f24961b0f01e35a28bacafbb6b6867dc13a76bff199210bd4e52be95305943fd9dc8e131
zf3d2f487dd38b325b54b8076781b0a0ac2c35089ba8018821606df3f55ca71c34a1d28ecfbce99
z0552d43b91ff278dd77bf5129f96fc93131858789813f42dff5d7946d3817dd0fb61d185b2a4dd
zbbd77b75e5740f0a6e644845346db1eb8516814ad504b74f77cacb9a94040c712ef6f2aedbe119
zeca1d978319c93680dac059db70d656db14a0d711b87aa1421a161bf6d08e45c48560c98a6ec47
z63440a684775e5214bfb731a8b6a60fba3506db5ad8895c308144e8c16e81169d2658556555c6b
z71291200e6d44fe7f49ba2e04a7b57531da5e11743484b32be98781e58831b3dcfcb6d0b178a1f
zee4754b61ff7c4c033220e714b82118a30fdc9788623f03a7a2779767eb3549fcbbda952abee29
z524d93b85460339863180ba54a84ea4a7a5032b5e59e86bd8259e6a2bb97c664caa543ade6872e
zf7353a6ac6c7f510aa63bca059105a23987ea3630eab1f777281a8418c65be391c2e06be012e53
zcf7b72fd7d4c6615f092767429b7dff3d731b76512cff1ba47037a19e8ce2177c24b293f0948fc
zbd10ec4abe2efac215f4b40179a41a9a23a6ee5ae6d89b5195c17cd45c991376c4f88825cea3d0
z4a0ef736a7fb088f46e8c20d828e44c2889eefa577fd36a875683c5de4265d639018fc6a6188aa
z9da8bf5c3c58b92201cd4c27f67d5e23a48fa7097af8178d4593b29b3a35f8a13abce655fdb7d3
z0338250ceb8137834952ed4d11273421b9f68d2ef74be5b1b330ae419280ed955f5dd1c45bf3fd
zc9c5786ddbb1540f4487dd35d9dbbe31422985c7808092bffbdcf666aa7fc397ee87433af5b47c
za2be334d3e59c3ef7c7a4c0b6a3d9c7ba119170c6864446a142a3cddda286ae587f5ba19ce9466
z3ddbb19ef8781bdd58e265911a613199b29a843bab356e2453ec3568f7e3891a4baafc9adc836d
z2d1805cc57ae519454b2e0bc1c65478662e3cc3b57a37de11258a65f082f07e237e22632c8e166
z1235290a5f79b368164f46ae81a84b65d5d7f53a6c1077537e04e6b8b5d79223db192afce9a6ca
z3dcb0341468ff206981e5b0de9dc80edf6ec945e40e9dc2fefb8d072e70619f01099e0dc86fdcc
ze8995ad234c0bdc67e4c07bb5e71a9da058bffcd83563e0a0ff8aab6a43101960937a85771abc2
z416a37836fe6325f6a8e83587d1dc3b925443762c44783c09f178386216b59d4ac1328f79cd158
zd28ad148a5a9be6bb0a7f3cf0a343e2fb8cf667e87492955324e260b75cc2ab0efd0aacf274f34
z3e3f6079dd1f5ac28b756865b6ac85834f555d59d20ffb0704b3a94c65ed11d152f919ed2a8099
z3328d50ece6dcd955e0b525b9a250b82edeeed1ac591ce709011a34b6a680a126496a8d7e7483a
z90a94d2f7b1f09b66371fb04f76ef11f2779db22303f5dabd20395a349d1c1a09b9666183b5a17
z5eae352a15699cb8f13c1b0d9b94e66bea499ec17cace954ea6b23bf4385eaaca12f62c700f4b9
z2b61b8222ee6f8c8fac187e7c13f8449a2a15ddecd21ff1f0327617c74e1f29c61119b2b356a1d
z695d9623c326185afbccf34da2b5e8f91ee4f0bb4263a51fe5106e8fcb20a089246c9325d2f002
ze689ae3d24c2a1dc92ff2bfe1aca787b93d90326d4b2968790d725b7cdf4c0
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_state_transition_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
