// Accellera Standard V2.2 Open Verification Library (OVL).
// Accellera Copyright (c) 2005-2008. All rights reserved.

`include "std_ovl_defines.h"

`module ovl_bits (clock, reset, enable, test_expr, fire);

  parameter severity_level = `OVL_SEVERITY_DEFAULT;
  parameter min            = 1;
  parameter max            = 1;
  parameter width          = 1;
  parameter asserted       = 1;
  parameter property_type  = `OVL_PROPERTY_DEFAULT;
  parameter msg            = `OVL_MSG_DEFAULT;
  parameter coverage_level = `OVL_COVER_DEFAULT;

  parameter clock_edge     = `OVL_CLOCK_EDGE_DEFAULT;
  parameter reset_polarity = `OVL_RESET_POLARITY_DEFAULT;
  parameter gating_type    = `OVL_GATING_TYPE_DEFAULT;

  input                            clock, reset, enable;
  input  [width-1:0]               test_expr;
  output [`OVL_FIRE_WIDTH-1 : 0]   fire;

  // Parameters that should not be edited
  parameter assert_name = "OVL_BITS";

  `include "std_ovl_reset.h"
  `include "std_ovl_clock.h"
  `include "std_ovl_cover.h"
  `include "std_ovl_task.h"
  `include "std_ovl_init.h"

`ifdef OVL_SYNTHESIS
`else
  // Sanity Checks
  initial begin
    if ((max > 0) && (min > max)) begin
       ovl_error_t(`OVL_FIRE_2STATE,"Illegal parameter values set where min > max");
    end
  end
`endif

`ifdef OVL_SVA
  `include "./sva05/ovl_bits_logic.sv"
  assign fire = {`OVL_FIRE_WIDTH{1'b0}}; // Tied low in V2.2
`endif

`endmodule // ovl_bits
