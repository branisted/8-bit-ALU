`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262ac56ccafe221d4824992a69d8a
z0056c786d54cd57e5ac49b6b8aa4fb7a6065bae21c146cc6f3a280ec9ff5fb2462d8759413581b
z93e05d192976492891eda0fca2f3ec4b5ec9a3861c90250c47bb2fbaec1ec83cfd5ee7ecb80525
zdddcbb6c783031a964477c94c2f1feb714f221d070ae59db13890ab42f6439a11c7132097f548b
zd0566d90979468eb425dcdf7edc2634488ab3209ba42f72a386c5010eb81b3b07deaa410644433
zbff0c8605d35fbbf8acadb2851a661d9537feec5a5de5206584aebbca7f4fe199a2a8c5f56ffbc
z977ba939756adca046f9f2cc0827beb18261e660ea6a308bfb159ea78bebec8c6560db90737e71
z1f609f9280be9eb705846ec8be7399c5399d77f815e203d0f0641e14b3ca2e41deeefdc9cfd5ef
za04bf0b14c2164fbac4483366f7d8ba22d21202810361a89e3a17f6c89e982127ca87481b8a547
z3b8432ca5df86d5f70ae3cfd33fc2fa54f2f2c7b569eefc39936b43831c81b0144d63ae3a350a9
z92d309e07d27102b61dc09fd3c869963aaacc3c642307db2d5769a0e2bbf647768d58b097db084
z9f840e1ad8dc80e194c2d0e9d7d2efaa6f6d368977771080a5b1a3cfdeb111c4cff8f4a06e2307
z773fa1cd515097b4b0285049bc92e098fa9dab02e9ed7812da028f5a0256df1c84cff05e858957
z2c93f77fcf26f5c76d8ec7f8c10ea83e4a0dbf5596da604dda8d1b5c66c2acbc3dcbfc18fdb6c9
z2d516b41bcb60e99249f6e61d41aa45395c66d1894115caff43c1eba8fd6c96d59c723a46cb915
z901ab9d1341eeeb0c040d9d7fbc22f0d5d1ecfcc2478e752674941753a3b05cb732ae292d2d8e6
z4be139d6a05c2fb0c2387a8cdc8ccdba2676496545c8473a3c8ceac1229e6a272e1050c4bffba4
zdc615c3564238f1d65cbf72e6b97a3d149dcfd7c6e0a52552a9c256b3f20aa7740f3de773a7f90
zefdc86b3be4e0e720229baa02a3d4372865d86987b5bc0d0a249cb30b21bc67d8924806623220a
z3336438753a1da837917a5f5806cf7e9eaef38f7b71f6089a0dfc66b4d7dc9159866e66e432e89
z61a1d1123ebe1fd77c769d010795fc54713115faaaf0273957d071b9ce91ac4fa2fa0856eecc7a
z703c9ddbcf840a507db8a23dc5ea3c78138d63d8abefd45db46b11d02e85e7169595bcc6b99afb
z3fd9fad632698e87ac17dd8ea0690a5b513c72a0eefa01bab38fbdd3d9adf1ffcbe8e3974ad3cd
zf90b40426d8b8b62f3c88a4d5342ac5b22df6cb8d0f057360bf84cfc31cbabfaed0df8f38a2f14
zc9c03750281f3c82e7304daf888eff0b884fd48364e035426949fa7613b53b933562cd705370b3
z145fc1544c0f0562f84afaffd68363d5612a20811d05ae6b62a0210f2d73c5a533c623429c64e3
zd3eb3db61c8aa7fb0e25aa113d08958a11a003b2f17428b314f2eb66f5bc49d6e438bcf3fa72d3
ze24dfee56e895d9e84a7597cfe277e199d1317c28b5642374efeebc59a21d15fd0b6169bca34e1
z80d64d14dcb3e1a69b3aecff553e01f32bf293cae407d4b963396b4639c571ef4b9667a99e33be
zcab59f6d261f7dced65d0c14477148e5004a160f6bc8ca3a9fbdf674da443c4e6d75df9ecc6117
zad4f706dd494a0812eaf4d1167901c5955674c90e3d089f1da1e4e7e0409179eedf6b1f798e4f0
z7ded5446f6cc16ffe87699ce272c88dc684ed98436573ec3f9e5af0bd3187b04e59defcd9f7c63
zf9a319aaaa572daad97728aac90c2a16761bc41cf83987dcc9d802309e0360156a912aaabd7d60
zda61f5dca9539024babb86f7874857418c1ad59d3b745bd426947ec12d39cf53f7d1a2a58b66cc
zf1d86f03f087d2b40b00c944fb37f2187d618dc262bec9a0fdd84ce136ae24981cc4eb7203ddfc
z515547cad5250a4c5d6e0676c5ec1359b1b32d4cb3bb6e03080ffbfa233c4ac9bdfc40a2908136
z0f47b7ea30c4e249d43440854fc3a7baa040ccca8f291f495f86717143e9aa127edf6eb19b839c
ze6b85e8d82ce4efcee37d469dee7d176b164128bc3f4730ed262226355cea4e2fada7a2477b0c5
z689b5b349a16fb1f6b80411dab0fedd96d62537555b02f3d6752e9f5ac694f8834a809eb6b53a3
z3f87ba90e0aeffd5018a825a512595ec176126d453eafdd01d26de5e720c6b484d44578d8739cd
z1958a8589c34e21f71c713d297c4b25414fae620cdd0c016c0ff1de8e376cb00cb007293031497
za32e96f1dd6baa552268eb5fa140eb25b8ecd0525f071513cde76a5c7b6525fe9df70ab9f3614e
z89c9bd6849d7251f01c2d7a9b7050823e4e82e289137e484e245abc24de997be29a732fe8bdcd6
z906fb9f8219ddd7fc0808f5a3ba1ede6cf649d653d1c77c69226c79e55e9012deb4b714b319dea
z371c4d238761cd42495e9cc86412f1234adb036c10662abbb10ad0c7cae117985e699344695dd7
z6d199c54e2c0ae4e72458b9063a962990a275dd797a73e416451de09292bcae7eb1dfffecf9e71
ze0b170cec8093a4315eddf62d06dea5073e17b6e770ccf662a3d8eb5d2a5689b71c8171705ee10
z5fd1f9aaf5834baa2f780657288fced13e1511cb054128431c7761c96e4b75b3ed8d8d9ef6f780
z440d3f12a7ca1118bb46fc8c568f7b1acf525c8579a21275719e0491556140890adbcb5610d040
z46a2a505d32004e7f4debe4ed373259d3d75ffa999d85338459daad92245ee54d1698be10aaca8
z03112e2188a8354cf431647ec8cc70d55cf8c2fbf2f3e0e31fae4a176b855f7c3a0124aca8f1ba
z11bb17d2dd2b6cfc4055f64685e743a53911ba3c37529c2bf44723b8e3fc106bf0de7898fc348e
z2fd35647f984dca75c43163c2249f12b20d8232afbb310502e301ab8f7bbf880a5fad2123b9304
ze78415a8cf485aaed1ae9a86cf78e373651844127de1da65c1b2eeff5ac34b9fdba0d55018e7a3
z3c6c461b1d47fcb810390418a865f8534a96a8d7585883206674ea2925517bbb9aa4aeeabdfbfc
zaf84f1fdfdfaead208f314cc55f3a2830d617dffdc053099312b6bb7b1de2d1f150a6122a1c59b
z830d5881780ed5036b5ae54ab8dce441c58f5c68e02aea1ad10f201080fa8aec612d05efa1f40a
zdfcf2a7c8ee9e3a47c24f3dfdb299b3ff50a4d6f889b6ac090f19bd9ae306f467e1c139e6be599
z0cbc8469aa51a73b096be983a06ca3680677e0af85b1aa88e659b8d7a2a674b18a683435398dcf
z607cebc27a2d333d05501cac7a5749e749c2a6a0656cd3c8ae3c5c7cf36c715faf99df1a509c22
z9da5ec1cc0268f56c10ef57d24c88420195b7bf5c7be41fe789aa95c5dde8a5026320e80db9fd5
zd920116cff869ebcf52d5a611f178005d22a86d1ec942224ce1e8db69888e1dccb703cb1977a95
z92fbf064f94b7631fe1d938326123058d08aa7b1ef7ecd0992f977745b527539ca3355a9396633
z4f94faf6b92863e8c50535cceab2b0f289d392cb5b15d1471271e38ef16ae00f01f04c92405063
z3093d4bc7bab7d67503dbd971488af9120662c7da386678c6e6a9d00d644a7fed70dcc9ce7ddba
zd9d90c7f7eb80fe0a575fbac953fcb93c7c11003de78307725dac732cf5c0b16c3833c8a6bad50
zca96d597cdf4d74ce29d1d43ae657cfb938b7508c6ecfb2510fec6456e143210d4655dfcb1626e
zdb7fdf135df0facfc9a52b8ca9571cb2b229ee46fb71bfe381cfcae38cf8f23390cef89c532032
zbd36ed262105f013e3760869906f8b4b87e8438053fc3b15f7f88adb9d99a40b65895c6ccb0f8b
zc0d900ee4e9e7744696be79d59552d3b3949a3bb0c523416e0a9437a7ce21e70d0d0dbe8dea08c
z85ae9765f6193c037a9d7d3d5dffc58e3bf0b2e7cfe4cd4f1801c02d58cff1f5e47d840e0e7701
z6a482a22c273e21fc74fa9fd7a0f4ef86695a70762a0f1d4efd87211c4ff7d9485526444a52af9
z29aa0e88f7baf42146c5ae9c0e81204dbcd66b30656f3eb6f649579baf9d6aeec1cfe6f014a1bb
zf3fabd019a86a0df19acc900947f576e5a9bc437a0fb971064007c15b90967554a1ba85fb12cb4
z1aed8e055b022e73365af1513296daff1072587718267f68279f5c63a7b7a9b4576137cb74622d
z3f751cb62417ae80f948d7a533304d1a1ab017f122c8bef105a158812dee167806993d887d7c6a
z5e5a6f4cc95c6b4e7ebe62de737d57fc53157ccf76958d75e4e9d760482155367e6ba15d9f6be0
z5029a9662a829f0863f03e21302e3410a9c91a55a0bf098c85864590aacedc950809e7854bb58a
z365652635f123cdd441072f4b68564fbcbcc1b711e2208970d8ff95e567820d0795f7001194fa3
ze5d17fe84191dc167c524770cebaf156e18d8deba207173cc8f8e780e9fc34e2244e0535b3cd30
zb32fc0ef3ec9b54e6f13a0e574d4c18de620a2b52d150c58059934548354a22507324469aa2d0b
ze164c877d44e880de8699196fd5a80730dd96ae45b3b6416230d50520a1a0910eaf15c0b1d95c6
z8e78c45e70566e01e41315b9f3174294e4b5f0f91d87ad70710581506dceac6ed958e6f78ddb45
zada5ec684fc03ec22ee01026fb2e3d39726ffb4965a7a845a2ab2f17668bccd4f9a3555767ff38
z0689e2f6dd57c9c3474856d734ac5224152210e64cb7525430dc40a8ba5c5cdda2391e1fa72835
z85e38ed634e31d1d48b3a46a2088c42a15831c22eb3362f248fa7762add0f162b89649fad4a6e4
z1e074469a84311a5aded893ed97951ba6a441b77ff9535094a9892cbabbf811a09e47267cfa581
zd1cd9ca8aa221aa92ea60dc8b169703c2f05021dcca649bf4d7422fe94119d972dfc3d52d3b13a
z25e6bae5a51443a4d62b528db2c970bbf77dcd0d2312822da14157b48dc238bb9acca9d16d17ed
zaa8006a87c4b76576f220cc0bff4174815c5a1893331265c96de33e53a67960b0b180a49c0f853
z0ba02af9be044a1950d7950c7109a4882148dbe70251f09259e9c8b6b6ccc6388099fcaaa49d31
z51cc0dc8ea9379651ed44df7c3a15aa1a4e8bc55049d5454afe5d418f2359f93d0593b0861e99f
z6935ade89aa26eb0603f572830a434fc3830260d569a20f14e204b7a263d1eaa53f5c0dc464752
z8b773aebd08ce3a05102f511b42cbbe15ed43fc5d4200da532b50175c78eb7cbda15d5e098a7ec
zaa21c47ffb4c3370371119c925b6d2e1bbd3c2d00d319a4639363838b40b789f2c6957c1694c05
z0f9867c969ea4be9521acbdfc953f2960a577ea707f8e20f64f714d2e5e9d74f7d7b6055f349ca
z4263aebfba0ca47c2a3f0038d1b3a2c3b0e2f0292900ac1108f7b5aded399d777a3b31c9acff0f
zf348cc68d98a26279a959c12e6e2c657f726dd5a5cc4d155fe75803f98ddd00a08ceeec7ea1659
z0732baf002af171ca64fe545e7ec8cfb51f9d053b6548fbc7d1d81934f9b7a7ad380fe6c956a20
zee7cbc958483a3e10104570b7ddbf9f2f23a55be82515bcc484c7974f8d6617911ae878d34c282
z7a7dd04f00b966c3b71598954f92543056cc4f0f49c0185aedee9623adb67d7984c1932cdcfae7
z893c297889421c7a55a81bdb5484a44a0bc35aa57960b4e42a60d99ecbf77ed7ae3a115f8b22fe
z118baa351eabaec3f9b4c8c7f0b65dda7347eab05b2450a326e02526397f524d8fa6687504b89e
zbb83185d1c1ac9c24be8738973e58d5efa59f907fdc4bcbc185a6416837da76ef2aa9a26569856
z37dea2d32f7a5552869746c2ec13c40d6094cb6cf6ac0d62de36a0beb1e48a723d6637757182fe
z0a8e0f3d18f409cf8761155d7177fdc6e5b2e15ee7d3555b8a209216fc0e07a9df98a4e6c2e668
zdfcc14da60c053a431ea3898d6a4483e31e4d43fdea94ca5cb4288466be9afffefac580538356f
zc4ea8b01f4d5a6648c21bebefc7dacacc2a010d63a6781a36203ccd210504db5bd52f270f80634
zd41d1a1c6e1dccf473504e233239cf7d3e0c63a8619aea5d0b080f4d5576105282526b386393e8
z69420b1526d8b3dc16b7731404f116b2d9f0f2089de3907eb54411bb813f2ebf8febe01686c865
z5e46a99946359f8d8a4b6ce52d4803eddfefa321a6f5f9442cac616bd1baee7f98b4802390e434
z1680681a271e74ebe83588944be6e00725ae741a206fcc72c21302fa512a5d93c37e65d4014861
z20254436b1d059b3bc91ffb140339f216f79abec40c3d2fccb80503586be179371c446eb80061d
zb001507faaea91ed55c89f0c2b78071112f926ccefef629e6b20a85b06ef570482c8e11650f58a
zdfe626e7f3dfe8750224947316252ef59858a3651f7b90e6dc0805bde76d3cd739f6118ae49aaf
z6788baa32590aaadf5b13a56c2933b4aa2992be2b344262f8d8f8f2afa94b3e316ad2bb8f5fb23
z63c068a9af8278d8905e39cddd356a331ea7e212ffd0cbca6ed3fd876d8bb8c92a4105656d9632
z19116cc5fb424584dc83dbe07a262e3b25b92897757e4bd3ca5f55e03b5e20fcc862ab2297e308
zfa5c64d4fde646cadd5818d5ca89e9091d90f8d8d86c7544cad1576b0633684c1202808f259e5b
z55ffb6a8ef3a9662be1ca1d06ce1c04b96cea2f6c6246a6c9b5ae1615911de48165bdb8a47503f
zd7babf214762cd38aa6e579a403906d6cbecf62d6d72d11cb0c319c28953e3460380c716465264
z4ae89fea4f1edeabf489d70d45c56904a23058
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_same_bit_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
