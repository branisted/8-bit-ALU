`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699166942afea5fb71013544a379d857e14685a03b77f81ac
z296de8f163f6909d2cea8160366dcd1069a4ec7b3eafe2a3ca97cb83086a74bd9bd0fdac0291af
ze44ecbc1f91d60b48acdd3afca719670e39357f5448e977180eb5cfab3de63dff72cea566f1646
z0120c08938d14dd8a38e1ee382ccf375cdfe4d19c75b0ed7c629c009781b4c8941f40c232e5f43
z17b5146380d9fd3edeb219b83674d2b7a1edb607f41678cde95cb4b47d46df23a7fd46ae218b37
z0989f0ea404f34e59583bc532b4a5e4407bd70c0de32180526897537c1b3224a441fc88708169a
z00155d21c0df2df5f465101c77bc93ab00803a4ee64bc17033a6405a312763e105117b518d5594
zb11b72507d9a6b005514b8b6a15fddee1b21a04a517c72efad33b87a1f2b9456ba6eca4fd6a23f
z539122fe8615670ce4e20bc6a14eb2879d240e20a895946048d9091cfd13c6911629d8f4c21684
zad62f70f250bd7deb0d6f359daf6e4a6d84087684f3c28a718783b43f040717f11f23555680682
zca7a224b3608699ad680981b35fbd4a767892ddfc4508fc7ab58af7ca1dd43542edce52216d2c8
z9168a4e192babad85b34d9739353ac4dee29ccbc8a204441bd447f1cc60a09a939e4fe53d66be8
z44b73bc0d951f02124da0d2a6a44eac4c1cce5bc3780ab2a8a4564711dd46acb375da42a8f73cb
z7be9c655909357183550acbfde5e3847260331afc908d95aff58de325ca9d3258a2a0a32c1e7b1
zb41ca01c1b0664ba10eb1ac386dd269cc930227d2c6b211157a028660679535a53671c88dda26a
zbc971d50243fde0f73d8692216e4ecf74b896f19a68f9b2ca3aca5b55ba05bd5457183d6ed7ff8
zf560e42a5cb123c0f5ebccad242f1c7c4c4cd3b147d0cb212042457f25ea567466af2a63edc1fa
zb2e7425b666e6945d6a3efea85ac48b9b8dfce3f01827efe3409fb9e53b9040a382f20c662a800
z23f49381cb580176461ab83bf783ac594b5a239ce1c57d27db1146cf6e74475b84e4574a032401
z9b23aabfb517a7803e6c8c07d3744a273a17bcca0a72c7c80446e55d832019bf74953a41a05e48
zef12029e6e2e2895503b27a9466abff3a2ab1a14bcc00cc8c97a42132ff4c2b4374bc750b52374
z30a95eeb30eaf219c75e55c53cdf52b7997f9e9ca77d3cec2deade8e9f8222fe96fc6d341dc63c
z0abf7f50cb7ba123a74c56e448f382d801ed9b042b4308133f0801c60f592333e2b50088274095
z1585090c6bef2b06a48043bd2ffa48af97e969c1aa9bf702301b0b6a168f572d30405bb59db93e
z2170b9ba923b0ebfec5e22f7cc7398b821e93376b4db18df6cef161374a579d798b9cefc6f254b
zefc54e3b575395d04e34f530dd81bbd6ada3685b3e903ab411f8d03747f8b9b3e03acbdf1951af
zf07856043821be7ef3d469a792f980da4dc6c4df1e2f58f04c12c54812c6bb4bb322e1386b6b9b
z1ea1dd0d639eb27e42ceced01500522bf5344c20f2045cb5d597502ef3eca8791369bc88719dbf
z8d59663670a88a7fae7c11c320333d17ab9755118a27aa4472f0b44a9d250273d31d8be81c81c6
z0ed25392190f632ad453754607ce2b52bdae928aaec574354bf91433d20b26cddda845ffb8d543
z813ae4489d21de26d560258a2a35e2349a92078593a7c44bdea15a98de57a8104c8c557127eb23
z1ce048c4be028e0b41b8190576bbd9fb17aa61e6182ecf40a2abf5280148846fedd7f4ee231969
z73afab30f0ef45ab1ee078d50d1780baebb90faf573641a0f1b91fdd7f5e0feb39305fed565e83
z059d1e8295b888d433655408ad5763634bcb494b3856dffa9f70f0cb2908bfe2232fde65b75dd2
za8aff3ece12216841834e35a832d39c443d866506a980a94faf5ca6d0336bfc5e9c31faed512c4
z7ce65b2ae724ac1958200a6ffb411add6667bc4b8f50157f000991e770a2e18bccffa308bd754a
z4205cf5b28f509c4e33e1dc080907006465f6d178e2596bead5f34a8384d134bfd29ebb0762a6d
zdbff6d61ffd2f11ba8af6fdc11c62b7a0487e4aa0ec1052ee8be8ccf046e267c1e3663ca8ef6db
z46a6efe0dd2520fb6e2f19c896d1a81ed7638acc24cb9ca1548e565fdf248878deda969eec93a8
z0ba1efe8dda686b1a7fd28fe06d0769e18827957d303a3677a349f625730c70404b10ebda98895
zb5565a75f6517f9744b4218ff4796db0a3214df7f66e365d916a43688e3dc3cbe5c7f88d72ba30
zbb3946c478b76db0a38b60b4e332b327291f32c5edadebe2bcab9b1d75d3cb4488e72f64fd8869
z598b48e6fdb2c8709ae95471043958a831a86758dd06b57ed3785a0f1d0ca8f53786bacf1e2f50
z74444532eb1e9156a65d2f867155e246c70c2b6f51edcbee2805a8fa6eacfa4195ce0a525652df
z51a867b71faf99ac1764b6fe34381d92e52addd708855411247baece83b5c7af312dec109f76d3
z84ea0b68620e60d1685ba86eefc8fc55cc8f8cec4ed4c0b096447430addd107a7b44a9fb853a77
z2e68b1363c6552f20ced28d37a2b161acf81266a5fb05b0b9f65f3a41cdf1244942a751639be1b
z30c46999ef2ef7a858a20fa02a53246ddf9a03707e743b8a73bcca618a32f38e745f4510b68776
z421bf00396ba4b83f9082936c1daddf1903ef42c74b0bca7e8588adbc1f3211524a7e711491c66
zb30f29cb818d549d5d5ae83184ce489b8f91e882fed3ce8dc6288c9472365f90865f4c18c042fa
zab5ac792d5bee96c2107ea69972a0e8b2fa8a568e100c9af59d3fe8c9906d86b28c50f2b97071f
za3f0af16ba72b2a7a57cdf1ca9028daa5a55dbe202f26b204b44b34a395f8938fd4b7c7a86863e
z5432a824f11e2ee1fa6f12cc3d6020912f0ea6f0f7d003f212186c7d7f70f60d5386823dfd9df2
z824b18405bfd65fd301f8efcb57b1956d28af7bf4f2d9eb01770be06da37c65d49f68671ba8568
zef350af8314279782fc1c8d55785082b013df95d67cde40d9a72ede46d0f5868f98594206662b9
z16d2e5f3668e50b7277b8392c6e7e5f571500bb7576f52430a0d91e2b66cb625ae1fa59d19eceb
zeffbccdb06009bf191714d21720a90a98a5834ecb8812d2edbc9760a4a196d057ac17255b65dc1
z82e1c4502584fc82b8c0f5de00de9fc83d36a8f4890053458eb38e110b3c9f407077d67517684e
za42d464fbcee8697ca93b97b344d4e82a3d9b3f615e8edaa74b21d2983e26746fda154ce88c755
z2565156316e86a4b5596a00faf0b848af68bb36162d72544198be02fd141d2b3161f3b58d5f4a8
zd731d07dde3a274c57f504738f7c5cdddf93eadb2b91137f261d37adc01e31bfbe08b355f53306
z729582e5c2386e08f8a80ba1ed2baea9394131c8c3b66163a7d5d574a250f4fdcb6f3c87a3bf12
zbd19203b64a4b415baa5ba1bdb909df8dba50a8679532393f8c5fd47da197de4b711e396915e8d
z2535ceae2346a4aefa516e24e992185e92ac34f2f3e285894494ab5ce05b0208ce366ff50cee32
ze55e2894d30a38cadb30eda119d28187fd15f428d8fa6283f7a9ac4555b7fdf6ad91ea7a86a581
zed44e8b7dc5103f9c92ad9d56b071124158295c993748d0917687f6f0156c8c62e922ce99e8732
z6bf00faad67a9316ef2fcf794f111954dd82e87c19665ac09c736d0ad01c29fed1bdb392b70015
z78d91b8b5b6c5b4618c8bca21ab193515ba29afc909b78f18a19412b56e1d868d415b3c1d08ff7
ze2c09a05854b285999a24d4ca1160f864d7972272f9ec3151d589c464cc4266ae027425984517e
zeec2cbd0dbca863fd55780bfcaa9bc2c7d8d5f3c976f6868cb4f6d9c39ab0d2853bc9740a19ebd
zceb219e49be7378c2e890bacb6e74d2d323cb62ad7fab8e3c83d835330ca6e6e9533c02c35b47d
z3cd08b4f9856ccaec101e2b3eddf3a54a9885c9da217b5edadb708d9feda6fb6d3fccd9e69bab6
zb2c906720c4d4aaf841cbb946bc57abe8c78fafb3764803428021665fee98d29d61538a3faa937
zbbe16f6f0ed8553cb4cf39671852298b8721309681ea03d9fe0097959637e8716af669dcbc0a2d
zd90dbef05527e3bb21a22e05a47f44ea22878ea6049c80919d66a6b1f3368daba6c6161f6276bf
z2b6cd7e330d10b30a737c08f15afee045d4ded1d3f058cabe32bd174599b40ea75e643359cf629
z2a14f2a3e21890855819d0d8d56b671b8641acdbffaa4d8dfd6431c70c3e3aefd8645539af8902
z88216195c702e49250ff8ba20c4a59c20b93196f971dfe9bdcbd14c17e7ffeda966aa30e929d7e
z01ea19245444f5ea5616f701c955f1f4825a3e940553add58b6bb6b28048d5e81feb77f9d72fde
z07f0d27cfbaa0afb2475e18af0e738ce3fcfadba8db66f923120104f4a0fc919c247b91bbb9267
z1f64cdf2209001e06e350006f33dec4bdd43b8fbfe05afe9e19c244500a970f04b53d0d18dbff3
zfe1a8d2fdc7df48592a1ae3d7d35413ec03e1cbffc8528c92183c8ce0dfc6487918979894c4580
zaf951967d4e8ed59228e0aa60ca8484919840a049bc4f4c3ace5b709fd6a7bbbbd0a9b0c5f1f56
z79efe406831f28873c726e61b13f9c7b18240f833bc56f0681ecd8e624f82093cc0e5fe97c8342
zdc8075ea7617d8790399e43b3220d0a94316c4963c00282b19b35c6c43cba804547f1978817d4c
zab0d45a663bc3bd8fa3f6ce4708b6ca6583a3014fe8fbe2cc169a2054052fccbc64a00ee48416d
z773a9da8e71edd6448c2089afb04a9b2585ea782c26db9849a0dda2f9baa0f057a37f9e42d9a07
za4f65f5b0dd81ee531275032d1a41983df72aeee65143afa73ab7e2c2de1813d2198199256af49
z41e9ccf5cbc57391e7eded94b358f1a715e334d7022d621e690bc106bc21ce1759b40bea1fbc3f
zf4effd3268dd512a7e98ebbf7e6101b25ffc6ab73363447260ecf576664b5101c454c00620d44d
zfa876e10196021c07da4974e9051c3a315f3b9a9d5436f9e1bf48ff948bedaf1723cab94dd36e9
z8ea8deb9e8a60759781fd62138743ff0615d535c2c1523171bd92065e610d70230d13d8537e520
za2339c47da413907be829e263d3876e67da2e1a134d5b0d9a5ec3765786ea5d614917c30570ae3
z2b6c27e776aaf2025dfb960f89be7d66f82bf11289d26442947e589021232bdc7954a042f6c646
zdd1c3995e006b88754feccce351b0a9b3850410de9981b2add15b63d2be59b9d0a39748330d3d0
ze598be1e6c506733b0134328f90ce71c8f962c92b63f4203c7c982b772fcb2b02f2d4acb6993a8
zbfc199962f6f3f53758165cc339b8a41a0591eb375f1bd19bde0fb5fe2f61265645418b1767cb4
z4caa05d29ca37a32676e659043177ac6cb2384b42382ac43c2bb852331b0a7586d293be7a5142b
zde049b2dc510c4025d77699153a85c213933980645e71d4cde35a85bc10ad2c937a7c4f08934c0
z94b2c9967c0dad57fef88908c2aff6a5194580674ef9e5fab6add50b51ef6b509bbef2f65da825
z70706b36e8621e0d6f6a6063db9d4283c5f20ba5606a3e93f91618bec4bf7020cef741a84cfa7d
z52b0da89959951e02fd621bfab2a547618949259af39de9f74dbe7dea939bd0dfa37737dade8c5
z01b239ce594ec82e5d97a1dca1e82ec2cdfffd0bc4a2c3f8fac192c1ebfd651c6e1c394889b51e
z0288dc788e8599cc9e1ebc15aa3735c9d2068e3a448dd7e548d928e9ac04c9badb5819ce762fc7
zcef13723fc6a60309235149687007de1f1ac1afcef1970cf29122c65afbe6a009d49999803dfe3
ze2573b772928894e56a88695b10cf756d85b8b932f3c8d95e6bda8cfc2cf652bcc407bdc6ccb5a
z7def53b81bad41a5313b8690b7d6b969f35833c8c44adc75963e08f4e31dd3dc96ed46ab49cf5f
z20b9957da2e26a55d8c87436bbf23a228931e8ef8acf0e1ca46b27be475038a1da8f8498616bbe
ze9c2d956c12196c78b5bc3c76dd57a20347c06291397d342f401bc8e08cc5dbf0c00d31e132d8e
zf3d86448d930d29b1f0b2a2b1197b4f84fab736d1037fb570cb5c13ac10f87a0067a086c9e002b
zc32ee80fd963e2b1f2c70e3367ed4a1ae0ec0c5555bbfc33c20af40acc68f64386f1535c7308de
z837879feb5ca4ca1d1eaecf156414cd730596803f826854f2611f3bc0fbb3f25d146d3fc099a8d
z034eb412a02b42307ef18cde697be369d0641f47c2e30ba85127cfc29bcf81ecd5b49671b9e548
zc86b7f032cd7bef2cad464d70f391804e95243aa2bfd0eae2f3391db3a0caced01c32cdf3ecc06
z19dfe2124b5fe677089523176315f06235fee356b64fc6996b92eb09b7f5b3b3924b77ecff416e
z33a954b68cdac757e5c5245ab6ecbdebc32b3cd35b303c6c0e619a9b18406511fe036821483d76
z1fc463613f8138f91186d3c90e0a5e793f18c943befe43c5e2b6fe8c94436b759d11d097d26739
z21fa2213a538eee6944742b9ffe1c240e5aca86ebdde018e23a622253e6f9b9e9111ae18bcbe0e
z65878557a49ce4bb8fb82b636de8d132c5cb25f0e530512ce00308332c5cea6db4668ce865844c
z4de9afb09ee037c52c7a5142695a46d008c9e438e0b86c54d0ab4afcd1d7e4622f8464029406cd
z31748085fe286a77cd054d81e3eed75d4dddb006d5c458371880b05265ae9986d96cc3ad816a01
z5f648323bf86ee669f06081ad45c34899c3aa239aed695c66c2ab4191abb07075f68d9a9633a74
zbf27cb11da07ce82e87322c7bb8d4fb747d2128e1c7fdc2dc815581c6e725b3d8536b5251154fa
zc96e9605864f487315fc586de601ecc40a020160c50bf7def791b7895e292f45ad0e24edfb20f5
zecfaac449924a9d525d2bc3b36e76ad61a0df8541744e52baca45aa6ecf686803c190eec75b25f
z5d4a74f9a702b6363837cdda1fd6c5811bce3178574648ac467f9bd36d2affc86ad6a4338a9e1f
zcd21dcff7d8de8fb2f3cf141efa637a97d312f0e85ab8a01fa0ca1224c861a1e9a1efeb133d29b
z21823cf05822b98a5505f7d85df2a002f82bb246f3111fb328d5642c5e66c452c111fbc49076f6
z9fdb2c91bc1e5bdb8993da3076aeef437e400e34f3d57be39388af30a783b19de94a11a5152f80
z162a3751be8b6318a8809530d47f2a0a4e452992acf0ea70772f8eb80ba0589e3b4756acee1a97
z548e04d17d45d95fbb7928638d3680bde151a2a348ecb387b81a177ef94dc2687ac0b5ba7aecce
zfbbe258ff88b8191c755239d92650174cdd5a13b9db40942756501845e5b7e6747e98b88637688
z770f9d0aebb16a89be283e64957f49d2a65874c3f121f6789452b4a9a1a61b2c9241ce88f493bb
z54ca9ec19bf6c5bf52a44128b9ea28639886a4a21576dccd9e8a33e94f6be33d26f7f6bd7f2100
zfdce0392643687a88df72cc3d5d6f796cac85465b25bed13b80c6ed9d714ef138c33e4447657a4
z1c815083e1bbb0718b8b3bd3bed4c302dda7cbc6b13615ed7c5e345126d1a0fb729379e57093ce
zea0ab7443fa9948fb30afcdd0a12bb308159b9ac081de9c858ea404714a58b0a711d8cf574659e
z5fc2785cbce140f47af97fdcaf1414c467a9664727b7878781d5c6480e21a322cb4cedd987a69a
ze33b0aedc339ba71cf263febd843a1f259db41f41256878b628fdb603a6abab0198ba68c883fd1
z838e5a98dbcf051e7f53dcd1fdba7f3e96f4cecbd3c43276dabc18be71f6d5db9e8f28402b91b1
zdc7d2940f73630b2a96bf1aa97d506087ce11fdd271f7f6692e0510cc8e4d7bc2157b7ea4952b6
z1abc1514f10e2fd187a491364eb2e03cf497a94df5dca8dbcc83b260618768004ab8c7cfe1788d
zcec80423617a708fbf54a82f52377aec384826bb42405ff85804a34c1d257ad79f20985716f2b8
zf89f9f930128f0e2d0cae1b85f5142acb9e310ff686bc9e9635f4d5f9e00bd9b25c6f1504f811c
z5644c814554f02e7184307ffbbc8260860eaded70e9a85ab5de64c7f37b59cc85317935fab94bc
z082a3fa51f019fbafcc8e3d37df245c872a4b6a85227a96c58a01ce47cabb1b10320e06b6f811e
z0d826f24e2a96d77e3ba4b7090aa60d75da6825cca1fcfdd9cbecb21bad8177eb881130e95d359
zfebfcb213ed9fb222fe7ed0463b4fde74a8fa8c041d4c40b6911877b34cf62d178bf4b9b87dfba
z29b0da29d2b99c2f1b5ca4474384399ab1aa49214a781e562d3f80906837d8aabb30a929a4dea1
z87c81ceb50a92931a6d390ac666c2e5b75e6ad3920258e5abfd71e3084d6b931ccb25f8ffc59d0
z316ea8f5862fc3eb94125cd0d125b07a06b73b9b58675abb375c46c9a2f5f36314544ab456d4e8
z5b5fd43c4f8eae453bf7963cea8854bcdd594d7a4bc70f5442b55f84047447ddf777d93ef82888
z7bc45e1a1f7bc422ef2b604c0f94f661b695558a6ca836b41d6d09d203db5f0f50adad38bb1b62
z999b03f132e759f0855b907dc36458eef466b7d7ab8999768c237832249c6b1e6e3a499ed89dfc
z0ed1bbb963e68a8d4e8d938d957890f63f5b339e0b80a70557b298bce00681f633502c8a63ab0d
zfed0ea77ce30067bbc3812157a5cec73067a49d4c37e16292e464759d4fa87616325e379f39451
z89a5a0a4c9776dd5f517c32feb963670b076ed53cfc588c566db29c7955d059fd4791d237fdf42
z21316bb6a59091015a9de7f0e30754d6abab6f03e9673dbaa99df867a7b2d981ab230c0ff2d7ac
z6805555b9112dae7bf3853416c4768416b1448870a1b10b374299d56d50e9b136b5558012ed4f2
zc666c0c364b5fe3d102df3e86eb6172ba738b54638c75bab042c98ada75abec0ea406b9f84591f
zc6df92a06cf36b314c17380605810d49216d5609b1abf049ce7cc07369f1b1ce943c229c60902b
zac43ff15e15b7515f6bd44e9a9cb22e58d8e509bec194e55ae3379fbae203556163c169a43a5c6
z2f229e0a415c8e5dd640fe7e98075ec6084988027ce541dce70d48b08a3700456004e839cf4361
z0dda5d481fa0b1bee70f15e98893150c5a3b2a345f8309ad7abdfb2d3b8da121f1f88013788abc
za03ac798f8d703e23c57cd4343bce345c632c7710f8b39885d1e20355c2175dd97abba4d62c248
zebad2f297e4ede258076ad4d0dde19479a9e157bdde5ae2f3777f00000d7277709d3c4fe4a6eb8
za972e4a21fc52d68e490d1ba3b5f21cbc5c929599887e2517ffa340758eea519fd6829a9c63890
z95973e5f6dacfc8a7e370e256af528dc0a74ef6ee6b2b11b270641c40e1d9e85ade15408cc2b58
zf5fe66fcc4e155050602d6101edc49214f4b93db4be0e3a6a8492359ced5f3b9aee8db7c4fd141
zf03885a213dc642717d542dadb4cdeeddf5ba96468126a0de7abbfaedf56cfba7db4221768ba08
z5e0cd83467673eb7d2a8a2361c237b9d383b6616416819b68083659ce58617b180bc80f3dbcc77
ze8ef4f11c570f49be32b6bf87c37a481a1598c0d94f3c18a7d4eb6a1e622b5cecd77ffe076729c
z700098765a185d4095bd58d8f2ce9859188b94838155c34aa26e07328b03f1e91033d2e3b26415
za95dd15f36412e4822883f1218c2cd53e9b506c3d43ee374860e313802eb10b3a844d8d965f1cb
z1c9e5d35f97688824ee1a10d0eec7caf5d4d3d5eec8f99b2a7213fc5b18a335f2a3b6ebc7b54c7
zc90317da5ce840ee1b6f7eeea5a6c02274f50434e7d444f7eaceab202094360161809a7f3171aa
z85f1376ec6b61731bde7d6cd68124f6c66c5bf31b2a8937d1a1ad9da49fed700d9625a03e5e992
ze9d4263f9a228df7cd72cca2de0982e6665403a37294c1f0ea5f0f615e2cffbfaee4762e861b1f
z3959978235dae36a88f62de9d7f8b404a8cbcd6e503442b08ef372bda71c259117666d3f8fc838
z084527cf79708d29c56f165785506747d5ca61341ee28ae0a870f8dabb9d34442ac750249af8e6
za9d3ce5ea262df80f64808a57d2b848890f0b5c42604640ef4077b72b20b9bd92748c2a9c2b61a
za9e66f8fe0e9fee384846faaa9fa999b9fb43637e0bd1a31b1c0d1eda51c822449c5a35ca05c7f
z10dd9d09b5b1e0e79737e1a67c042e5c2d940754a23a6158bf8bd3d8397b49f6192eb923799425
z2eb2e1bf51c8c561a54ff8791805edb49f1289056b9a5096c4b7c373f7f6db0f0748b1c6df657c
zbfac4ed947c2844e7d5d1fde9c1e05ff05a1ce331379fa4f7386ca0b2edcf10bb7c98c111e9a5c
ze48059aa2962550e27570b14a08ac1cab2f146664d5b756f45750da123ad794ac951cfb6eb04ff
z82a374bb7d0537f3d8eea8f80524219dfb1dad5659de04fd600a09ce764a7cbbf62df8aa103e9a
z1bfb5c47e82c873d78b33daea12879618799387a45a8571bee74d0cd7ff53ea26b2a4fada8790a
z8790cc4f35d840fdea089caab0782e47c48e4915bf39f83e14783fa4d198111a1e9e29463a7adc
z106e6f9dcb8620d3b34268ed91a51a91e5b6b8b01f482af6e7da364f90c8c5fdc7af86d407a793
z2bf2e558940e24417bc8d1ed5972419251f77e0a3deddfc6881305214ade44c8acb2b69bcb4ed5
z08bc75b74b1f8e1c21965f0e5b55d65bbb50da58f63d14992ec89f38560a3217f553261d0724fd
z528f2f18b3c6aef0e947d39c90b6be57791089dc8db218f7734f72079ae1f2c379c3af214b024f
z454b49408b34fa34182f4be75920fc9e001deef880b0014a04fff3e2bdc0a6e86d837a2c9bcab1
z44f249e5e8706f488c14ce1fb65b61e7d13a09f4512c63c9f63f2d490f394d4466eb49c09cb76a
z33d15f98d7c05490405d0d2e03089f24408d9a1f989881b0fe89e6c6a44504d8772e3595280887
z375c0cf1b33614ac516a113cba472070ce225a60f5c3dbcaa9d03f663fb05f6488c43fc47c894b
z7dfdff5715db5d40582ab08bdc04a383a8e3736e3bc03b3434be2a1e897862cc2b71a67566b7c7
z7f897a2a6b8d339aee163b9e6f2c0e3f117aeea8b8761f17a9a114ed9dd017fdf2fcde0e9f33b3
z49f150981863e299dc1d1dc858539c883660a319a76ea7076b3986e6ed42a53e178e7df5a7b6e5
zd74e5b1148d157112a8323b77a3ad7912ba8e7f2b6f9a53798fd08addbbe08ae90f95d6a50d414
zc4b26ec71091e134c5ce8d9dfd997dfd2c92422a2f589b8a863a3d1cbbfa4efee08bf67830e9ec
ze30319eb978f65b6e299b4821482f9b65af67e67d8f1dd0304665bbd130b4e9af274fdeebca47c
zdb5deaefc98bec9316423287840fb963f19d0c4e992f33c9bad49236cfab14bb6d105a9760fa58
zd1e56287c58ccc4ccd7d4d291eb3ec146dc174a870f6975856ffbcffecc0aafb708309e5cea49f
z109676d041c7546acda0728388fbf21682eae3c6324c30bb18ca0c1b506e8214cb3cea3986f825
zfca04313be2d663da8e2b086c0e7c418be98c2459dab97c11dcd88a5505387421aee8340a31807
z5219b4e399b2b9267011a623b5a253e7e799466cee4bce61c68e93dbbbede84ad2589e8b4f9568
z71afceab2d020ff68cba97ab8d2a7b8aa89c8b83746e320701ebcf680c9e5de56072e3d02d9d6b
z3ae4de9da17e555e2618693d209bb0a1f6498dbb49183ac4ca0299699e720273e0cdf7317a3fc6
z3bc5040f758c31d0a7cad9a7bccabae7fbe6ed9a255a7cace6866b663b5fa28425626c5f564e90
zc6bdbc199aa2039102522a965dee31887e9056e81bde4dd270b69d6745e44a77cf8ccd79b85bdc
z067046874834d6eccab42850ecb7dd009f10e2e57b827f2cdc454fb9434009df076809f6083f7d
zf2c5c52572a1146090ff4d3e63a48e90f415dbd9afd7ad09c9b13b7ead5a4d307ba90de0131237
zc5d46628bf34b34efdd3d1ffaff57bebee0a03c72a7727ea6c3045cdfa074a5e8a1fe5d6d007a4
z58eadea380bf5791c24dce6820743b26be7a5f9afb24c7832e2be6edce4fdb0827dd4d961a192f
z6c324e0aa566dd83e84fbb82c3ae2fc374075dc30b2b634cae6d49f045c7e6cd449d1200d348ef
zc16c9ab88e4595e57f039851dfbafe9429a4374e93947a5bb280fdcbccc6facb578b106424c4af
z79bce76315537acab384aef0a0be84b1a9fbfcf27fc52780fe0cf7e6c30768ed8531517b1721c6
zf83e60a7e3a6320ab8aa9d58ce124923ad71c697414488b7605509cd49edbf98e845942bd08c62
z9a9ec25e0356cba061abcf871404bc4f60efb8237b0cc7c795ac6a4236b25c6737b95cc5dadaf6
z631b7ba86662b44d85209aa1ddb43c80477ea03669b654ac6b22d2ec86e6ef19ea19769512050e
z92c31da57989c0ad004e5e941c9c0a57d4edc3f572952cba4bf95163aa8522e5986ac46a4ce70f
zc2402845312589b696459406815c9b0c0f5c7c142c8714a321a9e4235a030dc7a4e73b1c873d69
z63a1a522de85adc19abe07c55ecaffc4a2546e3410a9ffa49a5dabe2c8c545a3785d7502a98fcf
z97ad1db753bb07715bb289c6f3c75ffd283227b753a3c15e876789401ebd4950969ec7b339e84b
z7123301b9241006d67533f2e431403f21a86d5ac2b722abe60e28558a0c18c61fba59cfcbabdbc
za0723b6f0a6f9f8b2be514040da1ad4a01ceb01c50218e6a40c11860a3e6a6595f2b3710531671
zc94601d4c34f2fc0763a3e60eeadc92197c9c7b8f431760b932ebdda1f72eb205377fbf44fb9f5
z61ca0d3453b9f45c22889fd12f26658fdd79bbcba6ad78913503a2dd48d110aadae6cc24548b57
z736aa357194cb5116506dcfc0bd42de682e247a3bfdaad00ffd59c858d7794c53d3bc7249ca99a
z374415282219967071d3191f20d27f74f084b618ea2def8b088b8688fe05b46f9bb8a56dbc06ad
zbe8a63c1bbf6bda8e368c2d899990f2a60f748eda9df376a3cd43f5b50e3a83666402af8fa97e0
zbe7c61c4bad95c05eaf42eb670724994310cab6ae2568990eba9933a7d84a7fbf59992791a75e7
z3bab39fa030744d51f1bb5703e502cd4ceb2f7ff6cfe8fd5a19b907b4e650fff9e00e18a2f5edb
z0c315b6edd3137ab8b1079f191a5059c38becc76eac145ef18e6c59ea53c83dddb00e208ab6f91
z6ea3e6f4ca8bd8d9ced714aa1490771d24be9519573e8073db6fdac110bd2c82d70afc57054282
z1ce4dc19e1e321044df6fe56ebe58c170ffe4069708e81e049f950cdae7050658b53f1c098b3ec
z0957dc86178de776243fe4107e319934414d8e50cfb3192f5511211548765d870d2e1f5088d0ef
zc4e559fb071a84253b731725f31d08bb24384d33f24fd714e6f4c2610a6d3532dcfb27ff46bdeb
zfd34712eadbaa8e5d08a87faddee7248f904ea1450c5f51bc89737d0645dd7b5d9a5f5f745a24a
zd199cf664c83b562b9a2fb0c3df54124867081e3d220ef2cb03893edff65f0b6ec648977348fda
z1cc5318605f054c03aaaebde35a4b20e8cad9ab7585bb9095ce42209c4914c5dcfef000d5c2b0e
zf89d54d20f53af11877ab269403cd51d0f02ccc8d4b1949287ea662c3e7f5a824e5350515fd63c
zf09e43e26e075a334e889e1ad4eef7e3c76a8b412205661b102948f0ab8a6cb1672d5987063611
z7b86d8f7a6b9fa2a61e72f38891ebd91e13ce7693be17396ddac07d820ef04c9e28f5f39f0f212
z6f14f60ecc22d5b2d698e6236e45cb0215314f8cf279fce21a2d8802039b95b2ebbb6dcca336a3
z903a70fb7d37e3c5aaf59c7d342b8c7ca4bb705ae26d3772ab90ebc575fbfe21110efada042a65
z8ebfff4f3c52635b4d62da785c1d0cd104c7209c165b8d986f82a714de97c1f8b15838369f35b6
z60fe4f4b4c2b74179525f942b1df19bfe89667dbb48870c32142439cdf15f3e8a8047888d56040
z492828218ed2219b985e30e7ea751c2de8ad5d4ed1fa0cbe33da89abdcb892dd010641173fd3f9
z420593b4fde23ee14ce895319d1a215421afa750cd7f973cf616d1729365c02a38fadcba10a651
z3c1d2b0c9925cc2e7c42027933d34d4c26853b45659a677ef681f4cb1bcfec0c391ba730778bdc
z1240a16d20626725f8fd5856f030cde98cf86cc3449e510c04d29e6ce2641ecf5643fb9d023598
z1aa88087aa33b11ad1fb8578768902eaf9b254f5ba438d5e1c85f4dfa69e6205f2d04fbadede3a
z0466cc57ef6a86faaabcbd4edfb2cf0530cfa224aa234da9e5462ab53ec2d07483bbd0e22d160c
zb94b37e14e0e827c5ae3bf0c03be24c9b40de2d34d45b1359315a65e47102ff64996cfa13eaab3
zcb9e61293400d5991eea3fd557bd92f0dd6ccc2763b5298e5a39ffa91a52c65194cdfea717bc11
z5c64f82fccd9fb729629d46ed24cd5cda9c1f38aa720aa8768a55268442d1d5fd470b6a0625f63
zbf7a49e9ec3773b1893eba03d290266e7f4bcd83ea59ea8cede5a6df91f7e3b1995e05213a4ab9
z058ce46bbbb425ba9129315dc09c86346d0e9479f256c699b2f6e407724f33aca9af96abd9868d
zd3401d648d4e12d80b51d4e74457c7bf6ea4dea25961430b5601aa72a7fa747b45ad4232a2d799
zad47c2157600cee079df16c4b0992f95752248307c9f34ec909248239f890de6303254d4912703
z192be7f248b113a8e65d7c94826c013ce18a1bd1859e6ad3509fea1dfa88a42d8238e64205834e
z5a85cd050c37502f4fc08349d81b7bad7d7eb741adf7bfb0768b3ee4af15877c3bcb111ea82878
z5bf5f8c79e88c5cc4e790e3d7b0b057ef9e2cbba598a97176aa01a73c5e3e28830390143827c4f
zf442bb4970777fc96e238619793e2f5c093aa16df2cc3ff2cdbc9c132c2e9b46a0e66c4eb09366
zfd73f8320f0e33c30bc01882fe2580b147ac8b642114d0ce326e003b775353b3e948891f864c44
z2f60d7a9421a401801930795356f060fc1a66196ad36321f99bdcfbc843f150b413dd5d960c11e
z720d89b7f45a4a5f913f238f3786e11afb57ce07188cc57df1d06948ea1c56aecb657f8dcb8b2f
z27d4b6c4b4bd7b3de76c85cec64c09716978aae36b38d8d7909696f0ffd2a52202d196bf782c46
zbf27973fdd81fba5ed0103b912b86b271bbb9bb62e95f01ea5d0be36288fe81e7f0826a21a6c9c
z0c71ead5470d536d114854303e7f4ffbdbebe775278dac810c175723b19ca3f72fcb236f8a3ea2
z55e1e02f4b411a7132af52534735dcd3c3f76505d47c6c8ab9006a30e879b274446c15cf0a0f09
z55c25bb6a405d8500db12ec74e3f0431e531e80325a2de71261010f2ec3e39b50f26f2bdefbba0
zdc48174cd910db4c47ce092435c8a2c006168816c57b5489451515d5e4d195d3235a437779a6ad
zb57676477de654310ed273f2d03d80b6b6dfd9d7277592e35db94e9bede68fc38a15a010121dd0
zf684e5c811cdaa4223b9b30abfda573be225b908e689d211c1cc3e4b7338e4926018ad9c30bae8
z296f884917f1ad99ba11417255b324e3fa23d8a32b76ec39fa337d12281d2169ac28ba42e0b4d6
z939faa2c95c44f2322f61736baf39cc611b5f39348e0225ce5847632c4b2ee137060fee01d5f68
ze31295f90d247676e08af57438aaa62e0572aa935ee06f8b295f67af60e2547f03965f6498e4cd
z653ba27e737a627aa1c5ff88cbe9e354b8022900cd2fbe0948fdf7b1d32de1187b752c424ecbec
z1a633612854ab18972daf26e715db2bcb4ffaaab269572fbf9d3da588b91ae71a82c30f3206ab3
zf5ca68d12e762d4feaa76262c70027b72cbfc825d631f8b5bfc64341e190cf43c8e720ff36fc24
z7050bfeb35ea28c0fb0a7f2998849259cb88767db73347c313e0c47b524723fe3119e8a55e9156
z77cc4e1c360ef00a81ceeb5ad8fe0364fed4ec5940eedcb6ee174784661fd370da4da4838064de
z11d24365df7f232ad79fad2af564e88692715e6e811688d8a890e47967e564a983b0c10e7ce0e3
zb0e9c5b96438f296105de63527ab105164b9cf85dd2e50790f50c061c9fa1f4ce90f22a3cc8c20
z88f5b71c075038a66ed402956961977d3638936db080cede95b132f23b6fde6fb9bfeaad663445
z9d99905a7b758913b0f9ad262ee3f429bf760119c55a1ecc485d2be8673b2d9aaf6e878510b466
zf7cd3affa51d700718da5de683b058e280642d814430f23e144f390256d2b1274613be0d9932e9
ze70bc1f7afe9355c9efa4cd834f6babe72e309ec8f649895dbbe11c8c26b97f3ba007e9620ff7e
zf991bf7e23a9089c6e94983e4eeed3b666ead4a40e042016e556eaf648fc14db9f5906d37d18a3
zed3ba220ac3ec925e26fa79b227f11292556a677836a602434eb95d1c61da6d87cf5d966600971
z01c4559900a64a5b5317f2701acd616efdc343ccbdf47b1a6c69338beda81218121035036449d7
zbf17cbd32595b4c3d38672d7a5fe510407ef12fc9e67c72b04320f9ecafa3e7b28849cf3721afd
z4dd917c7d05c2774f4c8706e4f2fe1ba16156665b3a1f0840cf68ac394b4d2b75683a26265e5af
z56abe8f0f97f16ca232c4a4a7dac152be73e0ed7d7a40e46dbd39f30c0ba20eee50398cd8e159f
zc0b0281b6e25acee644d1767b8e0ac3d978a7db2f1f47a6d4edcce90c6166c4d4e418393406e1e
z78dec81b8f9ade93fa013587a0c155b368c767e70971c61948b771b32d8bfa6387e5ed7d3e21a4
z599181acf5c0a9e8fe2955c7de7839b952a69f7a16694a05846d0f6f5ec84d01cbb1d7f9b5d1d4
zfe580d25479ce929a014b07c7a609dd8b397b56ec3135128e25e287eefce2b052e81f7618ed052
z4b8a13f84fecdf9ac3d7c7b2fd8b69b1e936ad608c46d99186479b8406d17dd6fc8438a9c9a1d7
zcb5898ffd30a5c079824335d3290b8c0d70d21c739838779e92174132d8ba5166191898984103c
z7cab9c5a6dd1c6215f31a88659ac30c69e0f6304dd8e715861dd0ee2846daa2a0e86ec24fd3264
z01c093c5ceeb9bc5cd003442ef2c47024e4cc4b24b478e457b6d3e64fe5fb9cbfcc50556314330
z73a0581a5189e3e18a2bcbfd234e11551638bcd4259d42adeddd622caa415e1cc9b076e6372134
z7638e27d033ae8028988327f9593adece541c22aa6458236bcbc1987a1df155724e2e798d2416c
z4ea5587187c2c2563e7249c42a4cbdd6f2110c9c24db919d9071d1ec133ab82646eafea01418b9
z0737ef40a8d74fc0cfd194e737ff66fcfb5a3c48bb3426c80a1d22ac0a4eb505bb861d69ae659d
z30cae882a6d76ecba4219ea74a0014771b5fc81e11cef4a81fc537f10ba4b51638133ed890291e
z165ebdfe47ca70efe703ebf26443785fa2b6977f4dc6c117b794d68aef37e035e1c00d5cff1cc9
zd991a7c0ea9fcb58be68621ee0ad8efdd13cac74de3e7ba734c899aae10b6d1175faedb392290c
zb35e745f2e5f226e4932eb686f8d0110083809b3019581e62fecf2982a6303724f2070637b295f
z776dd9d1a0fab607aa51455fb51aba92b06ae3f70ccf9bd9c7330755482cac256fb61abc329d97
z48eedb78ef0091cd3765cb83e394fb8f5d367770278edf61525674dff5faeb662ef5f9864322dd
za4846aadd97b6e19742e1b8e2bdd0a5847dac54bdee7422e6e69bd7b2dc2b5ff32c61e6fad5d5e
zb83ddb229587953c23c5e16fe508810f11f43085403352a8f32cf0a00c3a06cfa82e75a8da4eb0
z865a0762f36e8e4732078baea1a8a9b3aaecb0b6ebd629eff2c9dd428d98cb7b737dba0822e299
z2593dbb25be650bd4e5a95a7fe8cef339d8be68582ef7bc3ae7ff0880e9dc84fd53272ac983db1
zb11d0d674eba203ea6f62fca492e0775eff888c621562c15094e212177ec53044478ed14e73bb0
z7953dc9abdd97816f1a8fd16966c6d804bb01c7e5c364d67aaf2959db21b889a804baa3412657a
z42a10de23d5539376832f82464654d85a37d700b63e776491998f10954553bda737271ceb0cfdf
z8a0296edb254e498db7cbc8e709f68e1fff39dbbba16fdf8ffd1e4637621d3ab7f9bb6af76626c
za2fa6908bdf5a6dfb271876db3d7635e8ebe4ea9cbb57a9cce9ecbbf401abea75a5602ae17853d
zab26cf8a08c94c801e9d2ce4277aac138ed8ce5912ea86486ad71450692ddb4b875a58fe16fec6
z050049705d67d92ac87a614a6cb1a2311a6068f722c0521e35c004554ecb29bd823fca6ed36144
z9e7abf0b956b465d7cbef3222082b824bcfa476e1136cb5630366b770113c0b247a9da70a5186b
zd2517c327588135f12ab9fb3473c1ce02226976ecf32db8188383046012061441d6602c6774694
z9d383c63096a2021967cf66caab30ca10aeaf5247f9b22cfacaf77cc38029bccebe0e61cff94fa
zfb4d1951071526b67a6f0eb0974d4aedcd0548c0973782af3d0b251c3c04272009a90f9f6bccb3
zb4aed090e9158de8efbd5edd505474c7f34bafb3335c84644c5d86e24dc4e80926c34f328c217d
zb92aea699aee9d0554814257d1318dd6496f3db77c51a6dbd26c74638662ad831d05c867523bbe
z0a4127948136367a78c98db0b587140fa26625c2bc7dfa4bee810d6c56c3fd9bc554ec6c7dd98f
z9048ebd264eea690629b6aef6552fd091a8175bbf38d4d0bbb306571da4f91bdb076e10b6341d5
zcbadce6f73d4aa60f84c75fa1f7bb666a0dac5b11082b91a83d0d7d68e84e58b5506967ed708b6
z5370c6fe08bf101dde3c5f44c07bb99f09c2e92aa717db23fda243c075fd31c6d5a99efa87b953
z5b96d69efa124f3ccfadaba28bf7eecda77f7437ebd8b4f5a6bf59878627bef974478c96c3adf2
z026ae064662ee88ab812fda7b33b4ac982e543b97877806cb494add66dacc3af452b2e6a0b3d97
zf76c7785fb07a6912492bf0ed4cad496dfaa1f89b6c3590d6fc78b12931855ebf3e015bb173a0a
z1ffcdab729d31987c2f84e23ce0206c72fcffef939bcd5d91b4ec06a8b68382eff21f243f9fa26
zd9166cb2d0c4cbae09d665923057cc08e87369b216ae3d155f598092d52fec98f17c4f0c640d2e
z08aa6ee6a76f687b1ea513d5c9cd641417ca6c3d29364a907b4ea90ca238445ecf476910f9d00a
z5b18559398db02a28492d6f0935838ae1ee002549d688f7f3e5e606b68fda10ee076c8ad80c8e2
z20ea0fa400435cf91f7dfe17da56b6c5fb285be4c8b1bd0ebbca9082609cb8cb357235e93ee79b
z6bd051f39b55c67507763985ef2175c3cec49b5eee3a8df23f6cde1c4abba82dffe6ecf6ccbac7
z84a0403ab2399db1fe3685500d3408c160f10103dd1f22698b731736da5e79e1ed221f80e7a433
z321807721deaf0da28336707ec9166f125ec60b3b8a7dba8ad5e4de3773b2f083541e788ab0f3f
z916026871c234f7ba33f3c3c8650b6dac6110d7a83f05e316aa9016fa7017f38334b0d7bb25183
zdee08736483a589557101d968ae50b2ddf169c85e880327d3f55185c829926a4d72ce2bbf44919
z22dba53934d9f051cbc96f95ea3a4f2c99bf7f8f3dd42e320650b74faddec2a07a4f7fbf81624b
z4999aff3ab88cd03d9759d49acbcef313a1ad4e8feec358524ba170fdc47e061545925271783c8
zbade047d9a59e8f0b9a66668ffeb223e61a79c45313b798fc1150cffb157650319b54c1e76a3ae
zc36650d391b8c78294147e3dbeafbdd9a04319e11ce5a6cdeae3c940227fb2346ac363d0d33fbe
z0a3362811553ce98f6b448dfb5aeeabb2dbc6e2b62aa94b5abcb4ff2617e08652eac1620584759
zb8d24d48e2cb875c819e24cbeda1fc7e619cadf01e024ca0afd2bfad632c8279a9b1635a2dde48
z051910fcc2e7ca5ee303e5eb821fb6dc3bb1f3052d3c1a60d8078a01a43dc5de01db40d2291e30
z1d155048671830f0d0ca31cc2b15e479ef5863762591c7ad3dab3fb00c7ff48e40e9c6f01cb30b
zf60cec6d7389b2d961fcdfe8e5ab2a485c88251be365902554985b4079632f6ca574fc876ed2a7
zc7b36df0159aaf8ce48d5f77395937453e56afe0b7f6e846ba5498f7ee4c03b0fdd765d9be1338
zf86d6adcc25179b46a592ad59f3395fdd5ae82848b32b2c850b59fc14ecfa4b63c8a1a7feb1815
zb529b302a3695f3c58b879716c03d14f577ff7710bcb727e67042e16162c0776158221d4a5374d
z769fbeebece46a5eff9bcde87c1afa9d2a14943d7ae2cd3eebd152f24f3077b58b24f7c1ed600e
zb98db36d058c62ac70b36a0a78da425cbd296d942919922cc43c135874dd1b21e785835c3641fe
ze48c85039d7c9cb607dc60488c8cf420e53b4fbbb7e6756a41bd9607aa530d8812b22c1dd2ca8a
zcde92fa704652561c9bd05447eb06e9117060492024c880896537248d4ac454168e4746108474c
z271cab34bc5cb4f1d41bc3fb4bc26671b0eba4197be7e8059f0342f660d318e531a2f54f538eab
z560d5072eeb98707ab955622791ca500d3f01c9435c8cfa28ca20ac87924ae45e6334a6cbd667a
z2f4092af73ad23ecd8e0680d193a03cfb852856fb8021e73a4b6ffbcdad31115c0cb2043d36ca6
z2a5788772623aec2955d20c0ea014ece1fa38bbf0685494f4c8783a9358427162fa3f90504c377
z73e35a1f5521ff49aa3eafd40d7fbde48aba51cc15750f1202cdf668c7352b0e46ed9efd85e70e
ze5668234388a6a8de1bc42bd401e1f24dcb049c560e2b3f8902944acb9d57f94ae30683d1d85bf
zfb810dc8f68996dd3d47c7f5492ec254b43fc2978290681d0147c68457e1f261f91766ba481147
zd47373feb44f2e7464594488d061d728ca3d6b67352bd161857b2ad58ef1ac062d0d9861cbdac6
z3754e8b43462f35481eb91ef929a2210146ec07020e8ed85cf5f33c3789b00f912bd1cbac238a0
z9d6c97fd645fba784a9360f62719514d00d4aa42175cafe97e086bc1d94c2bad658aabb1a791bf
z4a36f1b1bb9c109ad1a5b79c4234884e3d0cce4c2d24065381cad37119566ef87035852b9bad32
z21176df14a5e7c58879dea55681d045a8dab741437db4f31096fb962983ee1e26ee88e7505f7f7
zd51a2485c8f1b2760ef0d443ea464340dda04733173e6ef943ea87e396ac6003ffc85d3b791558
z0cdffe7056bc1670a9be5dd3bc63f6a85d0824fc2cacc9f6fa3d5ed9220f44a49be89cb887560d
z278b32ba66ee831b2cf39ba549d17df4f3f618f7218844f8904539d3d6a509680b4c1aecf528c8
zcd7d9a03d9bc7745a859249a714eda3f710d310d21987a1187ac8384629b32874488cfe734cc63
zee53bcf65c89212e397e6b1fcf8cd21d526a3ebdd54e19e24b73844edf2d4f4d912ccd449fd404
zcb98a6e4376b25759b29a80323a9ade8df97f758efb82ee528f50c4591999ea47b09d13a89df54
zef8149895ed67c7736430bb0d1501bdc176840422106fe15e99f7c72472b1cb98c201334067534
z6d71755a59f010b0121a360393624a382b1d101cd679b8f73e13f0f503fa122414d35b812883a7
zb4d9f7695818f49ab9c4f85722a3a254a0e9fccbcbe16477b3425a9711d6c80a8236e04c6675a6
z30ace9c31c73ecf0e459e38c9d4dc215db8304449953dc11bc95a9a77f40eb50f4526eaab809bd
z760f704072b9f6340fe5d6add36c9a71ca65eeb6cf2abe8147495ad8afc5a63360a2aacb6940c0
z415dfd5a02961bcdd0109a20d94fc9b11bffd31202d2e22bd1f371622c26e70ebace8fa746c62f
z0b6e5a9ea0e61a16343107ec8fe6ac6ec6c6669b2a5e2802d2519fa62f60b3568d5d0893a347d5
z616cd159ae1e20fb71d1246e41c86fda17781faf6f3c2fa41de016fd7eb5ccd07fbb046f46a61e
zb9219b640b8dac4d89384ff37ca26de1550b9cc089f36df94de61cef8a625480485a56d9ab9ebf
zde6d0a13a96e41f16f567b71449c80bb021d3d7c623dd1238dcbc6c3e6a6a288edae3ba137f215
z161a151b1437584186ec2b6d9b3d7b809bfe6a6b14706ee3eb725c3b34933469f381eb78338cf4
z5b51d7529d16e49953e279a17c8a4e163925bfdce8ec1851baa6f8cc15ebd3039d4412fe8ff853
za9a8c1e52b2edd4a075a9ce00d1b2df40c46fb89a95f7d582e1d6838d1af305c0889c3786c6a7a
zd2111ec9808476e7841a3813bab0a2198beab6dc0e38600298043f9e992ad47b1b952138938687
z947ad8c5aebf151c75e65e8b4e8a4fff922cceb9d4efedb6ad43253b57a958a65195e1c0fb35e8
z827e9a64325c5ae55d18febd8713c4050e1a039500c0c75c97bbafdf237895a8eb8ec99ed0e4bc
z4b19f253abf9bc9ac822059a3b1a71a0dac2918b1677f4f2ce8d5ec1a700d789e55aa7c3bfe1dc
ze852510d521fc869fc4217774ee150dfc18121caacb5fcd048ea53281aa3693f28b8311b93c1c6
z243ec5a5fd61ed40b516dc06e6727b30c6820999d2b39ed68de94153364cd6eeef00871b2239e0
zdc11de8f37f146150754230e569694de18d80530a37e89f00e670343a857cf56d8b70b9d09338d
z339b5648980d98dfd95a3d90e92ff3746c8ea3ad9971b8ea1e4de83f1d647a6113769d6bba830b
z3707d692c421f293e7853683256e530fa62f91448f3e52997414553d480ca0e30e4cd017d3c602
ze631be1e8c63079ab909938184d1afcfb4b26b438bf4e8e62c5fed0c03a40c6940cd0d62884543
zf2b261fc7aa68643cb49c365a6e9ce9746843dae639e5616
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gigabit_ethernet_mii_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
