library verilog;
use verilog.vl_types.all;
entity tb_alu_top is
end tb_alu_top;
