`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d5e386fdf9e2cb5152bcb6b17c5fb03279eb4bb766
z695f5d89e36663627cbc4150f70e4430e6e040faa587833e5d25d897058d3c2d050032c2fd2012
z958cf66b328b38f4ea6f084efe3f3777b3258b2594ba068d3a85e5ff19ea2240661a8784a10595
z814eb5a1b06596ea02a5e03dd660a072af25defd4ade83cbfb343849bdb069fe74a806d4a0dfb9
z1646fe7a492674cd7313c2495c716bcf3ab9a1b464fb6772a9eb762f57b382238961a44e20dc15
z7e103d803b28d872da8fd82e2c041bd020c7027707d1fb43c9b3fbf938dbd6b702a88c2753ddf3
zd33b98bbbd4ea307ec9e4b1420e259dac5b2462cccf2ef82174003bb8c6627c0ba0b43ab82987c
zb36e2cdfb91bb2990df17a0d1fcb1bb98736cd7f89fb200abfe4a833f906144dee57d8884a2e1b
z5217714811aaa8446e3e577af4896a1047103e0cb0f20d115064aebc488e5cfc0806cb059060f3
z86568d14b54778b2f10d702f4ec10fb8585d822b817903c62f96e7b809f501c241bbfbe3fc37ca
z32509e1bcf6aa92dc8c551687747bfe8bbd55c60a8d14c42da4041fa796ebd7a9bf163bbe072ec
z310ce4d4fa970f1eeb6a0fd735a80f14a37e52dfc1ad541fdd4f070ca16835d9ef4c5d54da13f0
zb12190ce1c5c4f15ca979090cc7aeb369b896f2490ebd6994c5741c59a4899b4187a9fc1264a07
z435f0bc112a5218021f0bbef713c4feb70f557a2d70bb240885aa41121403ab7b6a09b0effa5e8
z4e6c3128c74f938cfa3965f0cd8fec88675306f053076b00d3d5db0776a4a5bcea21905131a74b
z6d81f3d64e7412a007351f82e6b6689e1879a350b8bfa498365e4e6d8f290b3b0aebd65109ab2d
z7a6c69d918327f1e98e9daf5a0baa69ec4f985bf516260784065cbed19950c4c5bf265f659c4d9
zb3974fd14ab11fc11088a1276094f088af5b0c732d406372125ec81810b7a9da70211969882190
z2a9df0f80ea91bc3c4ff17109b0236d55d0120046284cfdaeaccec26724bfb74106d0a8f6310ed
z52e6430565ba85456916ae44f5d4d44f6edf76d1854c50ff1f766f5ab3a85e741365aea40c42ae
z9a7e0f93f5f6926ad3a0f454dd908fd746881664a1d88a12742081cb0a2f1cadd69fa095f6c9b7
z081ae68d4c2d667321deee5182765c15d9a8494779178e151f1aedd50a8b8059f85ab9dba24d67
zac1090cca3bb6d9b647b81010618929e361b97f54e942cec20f92f0cf41118e8dfb1c12dd16306
zb566202e1420cd22c046cf8976b7eaabc2dea284b7df442017dff8369a1897e6ccf81716996869
z4abd8350e9dd15fac56f6c81d01e2d2df59688aaa7eb6d5bec9ef7a33471d7c788076dbc956b99
zd2e9bef68cde838cf0ac164ea2676f5379bc9889fb38cb51cd407dec14cfb24855d81891b45479
ze4a98c80e160fa519c712d65d78b42f61209e2cc62a625473379a522868a05cfef278ad2876c6f
zc853cbe6ca565875dd546b36a948b255cdd6a984a61b40a899d9d036825b85c842a8d05f38a30d
zeaae849b868256073be938d982a2f2adde0e490b9728184a32129a22365eac878af26478ad0b48
z8e4bcfa9dd6415fb9f6a5ecae5d6d0bef7df13196c554ed2b1fc193ba8c8328bbb10b3278e597e
z92e64b9cc041bd6f9bcedd473d1bef5fa56628677860819bacd69b6cf57571911925d9418f67ee
zc1e437b3def7b9a4981a6818451db0384ab8061e725d2cd25c96faa76529c953004aadcc16fa30
zeace7e28a0b629eb8e422ee5fbeb9456169cd0fc0f6a33a00921a6460e6afbbdab0d4ade76e68a
za7e2e32e504d35e0c3ef492916f2c70c170fa9dfd6be5043a3a4a22620c8419096b662df8ce984
zf95cb49536f8a8e6422e36ea5d663a61cfeaf63c0d00f89bd91c0b90c5d78a7eacfefad3096429
z3c9f004f3fdb6f5a0445fbd1334931302d8a02d5fb198cb577e622cdd16d03a7f00c2dd5cc8213
zb1938ee9e98abf291c4e950ddf68555edc3e72b1ef83da43e1b7795e0baf8de05b6cb69271f886
zdbfa00c35d419968bba35632d25d4b34038fe63a9c8127e0cee715a8ab33443f65aebf31993134
zb198862814debeb381a69afa0a994c576fa815e6e9ea1e147c825a5edc9752607f94e746ec3f74
zfb3bc3a9ee18d54c50b2af85b5c5e2bf6224c41ee7000b6b67321d29d422b9202a42562115c9c5
zd0b17c0dab28b91f35dce8ccc6b301b03031ed93e882fc65559c88aa77cae6dda03677a899f547
z85f34b749793755e4ce8580f02ba498d0a452542ea5ca761308bcbd960031a5c1d2f67bd743f8e
zae274d7041c5c3a39144c35e618bb672049817e20a133a844c2b9de86e2d30a132cb60120221a7
za5233fc9bb506304fc20af19bdc27c1c97f24fa4896c0c5b12ea930fd12ed50cba61f51f9dd86b
z268cf28c0b7ad7fba2889243e76a6c30e08c776123e1f2ba0f5dc52242e67f9a56bd68adcec561
z184f04f0d1fbf153e2e8c5d1a53ef703c564829baf0e9b4d21c1e83102244baab1a1139cbc04b8
zfb41f421ef5f7ecdaf152fdea0ed694c70e9503eb27f01c768d6402eef8f3c7f28839988c090de
z655d1d8eb13abe1dcaddf6cca72238f2853e91fe8c8baec6dff921eda2612441534d36c8b12a54
za4a9d49d6b5e60ac586da33db930c964becc3b2059428ee34af097ee3e6135c054808e49259a95
z17e58dfe64aa7d170021dd9b141ed9624b9cb3ae158544d89f59cc80b1ffe5796af0906577a242
zeb6b0a1c80f5901f3ad38ab19a9f476e6d80acf66fa69025f5fc38341afdf25fa10cce96e1f403
z637b1fbd1ed5d10c8db571c237823d12971de7b17577245b66b950c91c77f3dbe9d77998e62f4a
z26afba45fe54436b206db90b37d5639452533be8723e0e58e6a8e1d9ce6204f02489993ddc9aa2
z173f46c2f52826a3a6dcfb3079770cba9943d61adb775965dcec9d196ad600427d72de8966f8df
z2dd5e58e63730e0c58aede233a1ed30cd2e00b9d4378fee8ce94f14a25d5757c946a5d01af345b
z1d8c3362e344649811427def8e0a1ce35bcfa46fc5469828bb3a2a6a835e70657d63c8c6db53f3
zd0a2292477ec805cbb49bf6ca9df109f4c1a50a49490981f3eebd603d2133de1d89b5f42d14d32
z34c095d588e3bf4ae9268bef9e46a33131534ed156c9f0eff8339cafd95052486580d97624fd95
zb34ce69d56c937bf5e536944cb203b4fc76e2a7258e62667dca57d0dc167f24b4e94ac55377645
z297d74d38a2a1d7c02b805eef75ce71355777fce2724b2e83da7c94d847d3a45c1da41d5d54421
zc58f39dd536080e61b29022080b78261b845e25424a58692029a79ccb1c67b0d34a30b18b40fad
z6400a4b46f265717f595a1ff1930f4dc6f95d1506b4ca241c7340187270658db6d693570f61f4f
z386ee9ca42424251f1474e005c09da0cfbc2147dd9d5b95dc5ac0d9868433bd6e8f88f68188243
z5e265fc6765f712bbbb06646134115ee036ece3843a25c3c1e3a40ec79081c0954557ff76170d9
ze53238d364449f4f54acd76fec4dc32d5daa1623591c29b15c0f1a3f6e53412f722527342259d3
zb27ee00ae46a9cdfd9959c909647a954bf3e3eafe6239650460bb82eb7af6f66ec095936c57de4
z22afe7a9042ed1da9bb2accfbc53b1f7be404e0506b5ca0a8839191f758355ff2020a2df988623
z64b3e83b7d47180cdb80e925b197e1233e796507754792aea906fb2e2d1f651c7af79178d7d910
z3d0d9f9dd1012f451cd0626496906bd972497ad847052e18571b4efd54fac135400dcc23aa90e6
zd1bb2c05d69d4a87b375dd9c6c31f01f77c1cbc84dfe787bde87615db66893566a7cc26cfdbca4
z981178c8d31b490180a5266b0db7426cef62172083e827aef45a6c479563eb503c2b203ade8e23
z9e1d1c61d01ce5d8baaef92aff091f3a63976bfca893d7242e07711586aacf3968c5bcfeb05ec9
zd30dba591bf0e3b475f877afb1860d6cb5a40a06d9d5545e38786fad1b7af41d434adf125a03b8
zc3fda5d81b4d6c4c81c0b1a2cec42d02c90ebd2237ad3c536b1f6d58e17d09ecac5a4ad6c2b415
z12233d392dd167ddc8259245b2738f61abd42c31930b9cdc01dcf8aa989e0400782ed79ed9fd30
zb3354ade8293b4a5fbb61517e58f1b7e8a6ed22e4b783550ba39642ca0b8278a32559e0f985a1a
za2204377ed7c61fa592aa8b50d5f3afc8c25b3b7e735209f2775965fb0d6ba2b896c3659984338
z84b1d76b3346873fd495794545458f460b87323394bce62bac77a460efdaaabfdb7be9e74b3929
z5b0a91fb0ba4ee1c73d97ee0a600ea6fd68e2c0633e06c4e0c51a38b59cc5dec7daf3b2487ffe8
zed837095b5a4e6a33467ae49c22ec071b95e28f3b5bc9295ac81de827a32cbe0382220214d1ab7
z14ee4d78ce1a7e1ba260313e4249c2b6efa59e7ce205676dbcd8847e1bcf55163158a092bb46d3
z1478c7e3f9a3276ffbce5033595a3ef74880e7052835fdaa2401615eff85e8109cc9ae9d1a8441
zf5fc85e2851f37712aa67f410d177b1cb7cd7774bfc78bd1dbc4b597a3a0a358d4f75b2c607ed4
z635c79cd4db427c382f8becdee5aef144f10f08d710ae3fa8307831ae37b1cf5af2f3b60c82add
z4f98c53bcd77342ff1c96b591599ee6d19ebd60833f243bf221cddda37379aa5e7180cf42a9ad2
zccb48c4ec7388102f1ae18e09a1dcaf221f67b49646ec79790637c1d8d0f7b38aa2f964c892ddc
z9e78fdbbfdfa9ead340030310d0587b839b91424670a52d2499c4c3d996bffaaa62aa9e711d6ae
z54b9d1f0dcc545332b70eedb0619db447c70d8596b44dca3abe41a04340d12bc2b14fdc1934790
z2e1147e4fada79c05f7fa6a5717a079a67a82b6605c5b3889f2913ce29d78af342af53da4bf5fa
zea6030caa79284efe72325c0f0cf27fc7e1e504214dc17df226317704506061f877acd2eb937a2
z914aa708a213118380fd4fdb36054d05be15548bc45bede79cd6a6b0f5aa8075d54b5065aa7a1d
z8c0035e1d510b7b5354f5c95b5dc6e8f01f197413c71a873fb026d6568dd892f022939ef3bae45
z8bcd4de9eaacb3bf74b4aa1765ce6cade24c8847fb6a49b8c78a819685f5f5ba5ea39370c9a3a4
z47b9ec316dea139317219f57fbfe22310e0c456d0ffafb36fad702ffee27523508d689ffc134f0
z9caa357addfc062d41ad42c5aa03977b08a4c15150a0d8e256b0063e63945f3c4072c203c89630
z149e761566ab336ba58f0fcfeccf049b7cbaf07e65c511c84c67b3205bbff1bf2e6df28f6d17d9
zb9287d2271f5ee49ff9b7672718337d4e0564db45a353680287f29849c136e5bb41b8c02f39631
z61c60bf8b5f42a34777d7b92d0ae95f5bf02e5916921f2672b02992833e901c888c28119479ed1
zdae66ee51122a0b826feacde0036ef8f3f10e8d093c0a8f20dbaea6aa2da5845e21df17b87a24f
z73dbb2127f39277c041e8df7d33672028b8c7b8df63d2c2166ac14f3893e073c2c31511be5b840
ze54c8299ff3a4d453a20aafdbf6b0e49c140c43b7b875a24db3002e366f232dbf90b9d509aa6ee
z162bc8e3f10969eb99f848e5c77e6749304ba67e3196464259ecdf9793b193598e95b5ed631a6f
zf737b6ccf9e339ad6c27ab0fd4a11e0f489d60b2646edc79bc842f9fa002898adc0015ff4aaacf
z78e3c8cb663821cc10ea76e59df991974bd5fe17bc5f6cfbae39ed0398595dff222090f18e5559
z53fa1f7b707212b5a7f20fe5b195590d1d372924c46ec205138a1bbf175f1d727c7e6f7f1f60d7
zfbeb939635120071fdcaadcd9ff3146ed716d2f2c9a3d8262323bf19d39830c79f3daeff039ecc
z2cb8796ecf80ae902678465ec6fcc5c8bb012256c312ee78dd9b7b0848c8f1ecd61043c9297693
ze8d3f034d231f7b89c3b9f20a0f2a4db53a5e7b8428539d3d6ab95f0a96ea2bcc5da65befc3c02
z2e5d976c19573f9b0f3149a5b5cccdf202dbfcb988c2f42fde2a5db6435f985591297e99dca797
z10d967704778ab1827b1964afbc209f15282f8f77e397dbee65b07300d6fffe1f0a9471974ec12
z3345204df2c5a0c1ee0ed15ca2fa519387ac76a5303685034df75d37e98d099de84b2f279b96bf
z9d56d9564efbc5b376690e040faee22b2cdb09b5f0b52b1fd86bb5f2b31553f94dd97760030780
za62891986b6c06e69e9de3a088c06b0e5b7f1d9381a2f06c46e0567c9d25cefa2c3fbf5ee3db13
z14077ec379761244c1c10dd663c7bbab48d9baee88909369c50cc312fa53bb6fd2e675d302457a
z556c3f812fbbfbb40bd347a58fb4013175b2d28f4f94faa93f5fb3b9dcd86d203b51fe49ec19fe
z8e313feaa6bf98218aaad38b8168312ae531c8700f01d2b8b5ecb6dccebe2df0441ee69923f01e
zff35b629156a5ebfc37dc3352fc23192820157880563bbd9a6c27a31fe3f45238afc64929be50b
zbc8b23de361c63280da335fb299c400998113afb440512621b4c74e89bbd1079a6c251a7fb6fdb
z4d013646be63cc9fab072bca15b773ea7885f91120def0d118683a454274addd06248207295038
z0cf9cba2d533e7e0c39ad09f586f1008c3cb2f3fb55f1d2725934488e338915b7708787e8e579d
z79160184c75cf4efb1c974fcac301d6bc995d07ff81e4d4290660fef26fc58ce14614b9717a1dc
z03522d85b1f5531ec8b4f8e28d5dc5e7b87800a63cdb9dada3ae16af3fc7e766be7b26e17512c3
z97e9ca8a34823e6f7756c6169ea1b192aa03f503f0d4a083d548419cf5337f23a02a62671aef67
z12b7743f2b02b0d8d1e55340096b6de8231c9bb260bf1eae3276e3b8dc8d10d75128499b0749c0
z5a24a9dbe631dd9f6524d3e4b02b35c32ed9ecb53a029ea8b488cda54a9396dd0677707b2f4da8
zd8795737d1581b1cea0a11e3fb7717f11754f15cd9a0c950ac332c87f67dc848cb5519976325ac
z930e2444650dd2f6f94d80e7af6f2dbe702cd5c41469051bd61017237428ebaeeb10a72bedb74a
ze974cd91478a86225d7bd8b305cad4caf64924110f669b5ca3aa
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_same_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
