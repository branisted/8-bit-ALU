`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc6039eead
z7d07817cbebcef2e23b1e790fe833185ea823248656f1b9f541b526005ce77793c3bf75bc31386
zd1c797cfbe346b8d30cac8eec15958a28f5d44aefaf1736c246ab55c9222405df0b9c4a173f981
zae2fef42a3a96ee8abf5553ff93a3f9612ef59a9d47f6253c53f6e03083c421fe768d7bd462ca7
za039ada6bea612acc17150a1f3cfe5db7e34bdb0218850979c0340904609b15fb0df159b926561
zf9454bd76859adaad6d36d415c947a257b7e47049ef1701e6ce64e7dc6fceae25bcfa96cbde8fe
z2646b5588196a9ed57ec110795144ed71f5cb9a13b84908a19f9b265f2870f499f80a5b819fb96
zfaa7e7041409c3dd1521faf012c8b215bd25c36ceeb5c5b018f67088faa5bb99239cf304d6f1f6
zaae1734ca4cb01b62efab7a2d0dae23db30c12a21472da13979dd5d339a3b0d656f19866f22d69
z2c431c56758974458076793c4d0fc70452c7610ee42a2a7a3f24c0ac030b57ddfd36b844df2b5b
z03e92792d2a04fee5805c60ef35ffca5090f93489e88c2b6220e9b5f54110323e9db48076fa504
z13e69e09af0f0b99d3f3170be21a0003378b65b860e3a54c8adb980c219d028ea1d3cf962ef53a
zd43477596575a3ca9eac7ea7f111b754d3852575bbbb6c968be1a78d627a01d684f9a942d47f84
z00c38617328d2efaf3ec0f6fe289b1540d9cf270e8685bda5768690c287ff4fc7c81dc3aa47965
z4302e44542c9249838501d97e4658856e682e4da5ed5e3cd5bf1ac1866964a92b40646db5ed5be
zaf21c2e7a4174283d5acc90be700f5d502b751dd3fd2111951892fe63fcc417a2c10aa95faeee1
z19d024c219aaedd6e479c29b394e73155a0c11098cf44cb4c38a00874d9a6597e440edd2ce33ea
zb5ea535606786148db6037ac2547326c35e70468ec0645c27358d3b57f0e201a9da231153101d1
za7de3a59aa01883f2023d8cfb7a52fbc23db6a2c04e5c5a7ac65447573192ca8a1c65848f2be1d
z688b851f18434e5d01fc7c89d1549b42839209ffc11f99cfa8f6f8a349c12563428419c9ee7043
za2ed0e57de77c5aa3abccfd892f499efef36020f2cfb8fc3261870c55a2901261804ad55a9dec7
z4f6b3a415fb2de07109e76604031889e683fbd6476ea05fc55a160e0302c35c5bc8c30c5e830ed
z62c0fc8ce5383bbad4b8097f63e5a1488093f60ed8754c5d77a55704a64584a9ef94581241a23e
z5271eba6eed89ac9cbe399d6550147ab8570d06f3ac0e7b10802bdcafc4c5999b69d55434c414c
z5923a4cedf6272bb0eef7cb13685b566bf4c9e7f23b82658b90376fd4ff679e75893962292c01b
z4a19318154ed06dae18bcfc772eddc12bcbf1304f355613d5e74c9df1e904e935c3a3956c4b969
zd8013531489e94189c8306e7d02978cd5f135ec0698586f557b9ccfb63b0219acd112b16a5e768
z325e5b7a1ce77299ca22844259ba9ed714d966b522365cd2edb7944bfaa45b881500d96a46f241
z74e26bbca2d94f532a6321a7f429808d4778fb70559466a48c4a4c968780d00728e2b198f44a6b
z5b3c23a55eff1bba12a3c19eeb255871c3a054ab3dbd3d14b9718153281835cb8e05add54d4ea7
zbf6a7feb623c297612388b6934eeda4a5bf99d3da12e35825135819d4120375da7708835a84b78
z4aff2037e43ac75196f8fc5db0418f4bc1ba5e701bcbf31192e79f90edfe3a705c8fb1deb15f15
z312937d3689e58a92ab2e7180c4d8de2dcfbaa5f6df6a29f36ab253d414310c1799bdb5075f43c
z7593354d63417caea6b84608aad695d248e665e5eb863af35ce352c08f572ab9c28cff28644d0c
z71c3b060e6863f33fe2a1971191a54e49acb3ecbc13aace6a30468abfc86299cac966f038e1dd1
z5d1726389edeb38c88a4b65cd6c547e822e1585dd0c9a5d8e35d6d52f435d4ed923615baf4e703
zc6856597fc04f11e41a6cd8e0b1bcda837ef4e1a08b7ecb626750c08b0f56c66d6e5059be6acd8
z962318f84e464d98864dd48520344ae2a07fbf479036421fc61a24979be0c0fa35313965f6b8d6
z6a29dd4230b356a5f7f3d23d0e91b3821fc2eae1c4eb695b4f4ebbbe6e79bd8c7cd645524b9117
z23de10e33cf595b0f5fe79c7689692508c81fbb3ef14a2e8709e79dddf810c6fbc5af8fcacd880
zf2bc4117e3c6a509f29c039ee9fa91d14c8020158e7f185cddc725a6eccba4e108d269f9a6ccb7
z67826c9a91bc0086f5a1fe3f36e416b1e214efc96d304e6629212a87017ed381d240ed2a4b7349
zeeee2137dbea294aed7b3bc70920acbbbb59ffc2cdf0de346aef634a66dce6d5b35148531162dc
zfcaf15bb647637a2f77339f126785f9dccbc061f9b6d57fa7260faf645680b471ab286a0bdb09a
zb76d892e3f44a83cddf2a192c4f76c7db3faa862722f0ea9ecedd5795b94397b5b175c5e729c48
z4ebc2759c3e58359c176677bb9470a1e490825b48d8d5c532844332b83414469a2a730d7e0e67c
zd03c476ed255c6aca0e549e0518c56404d40cd20f6c39e04c7890693663bc2a67049e65db66dbc
z9506443b7f4006a81f75f841a029b298ac554ad96cdf22319d98c9d51f3f84b9cbd2541b4201a3
z90c76b3e427eeb7f2efc50c4d34121fe9832021db71184e0692ec6d5ebc78acc549810b9ec725a
z636c0bf248e279f35a3abf66c6a6ca07df6cc60914c47d6536903d98d8ea8461faf82b4302c38c
zd17a740f07f41d81224a8ed8c33afb15aff2c08624119c35e1eda453bf1a87b8964346d4d16aa8
zde0bf3fec901da7f548c94a9ab0f596ce8e69d1701086d52a074fd5ba146571d6efa1395acb0d1
z1c6cb3bcd878107842a831b04bebd5e1829b214c1b9ceb79e5222143b6a8b969a0f7e8e8aa0531
zfe5c630513fdef3de521d36bdcaee95de9e50f638909e807bddc0f8e14a6361d41cbf2759260c6
z360c8101db47518cfe24a9775200a43f72d63fde9e04447dca8588b224983213140c100bb95a67
zd8c4cee8bc2d65ba724ef20610e777ec8179899ee003bee0c90e7f875f4d1f930205dc04b58bd8
zb358638d925c850adf507ef6fa572a715f79c10e51a3824b0fc24092bd2f98c9d37d41c273dc22
zc2dedbb7fda411a9ff6dfc4b1dd987edea26c01bffc165c0ff1e4253d8b4cf126de5063926d07b
z68a8e7170f4d62b10d7f93dc7118305889b82b1703eda003b46c4d25e4865d21b9b19c2816739e
zb874b09ab1329b0686af1ef9505d75c93278afa95a01e8598ddb0368d42e45854c30ffb7b32166
zcd73a3da564379c6845bfda53a93b59045e40f90f1c0453f854d8ac731427510b982af9089c0f9
z5c10fc8cd345624e01a1d16549d2c34a8bc0999c179dff55ecee18542e7e4305eefc080394dc6e
za1f924fee55854b5da3cbf94b6f046b7987cc70f5b0654877f6cf3447af3258efc9095644b91b4
zdd77392ff16f22dfa10209972ac5175299c9cbda34176fb71a867cae8a270650ab82df5a355692
za56a2bff5609502343967a6d7bd4e339790ad60c1b4280e402164c56cf2ce3c65a4d023e6fc4cd
z30d24b835152e7481499629876eee5cb6c4658ce3d1c6fcf1ef7386446d7e85c13b31b98ab3100
zf887276780515c2c25503b70ab97bbe702acf55c0d8c612ab5d109056b5895803657027f7c328b
z1bf2cbd12af810ac98e6d24e0c63facafbfa06e53b4632a9a644c8a6556e210a0081e834395d42
z5d92dfdf0c4c42f66b2410cdedace1073ddafdf9b18650d7d6c98800c333451852176bddaaed3b
z2c1e39736e2cca401a9dd385b1c1fa4fc77d747a82bb0be66a66c2acfa1b700badbd41c719eaa9
zca321198698d24584a7f2bcddbc2bf28a5fdeb9269261603007a7dff460b3faef8c78e165c9972
za72d0ce73451ebe0422bb74ebe45ac649fa4639f24bf042ee0843f5f5e33958dafb242fdcc00a0
z2bd8dd15cbc7a45ae245a679284bd8a3eb485cf6b465bf7d70f1693e2ca6d35677c53c17926866
z6d1bd60e2639996ca1259d026735e92207c7291e5c2b2b38425d671fe9913bfaae228fb07b41cf
zad3ebeb590809f23b05e76b546fe945eeec3968575427fbf049fe03e9f9e9b9dc267b43622f7ef
z4ed1f8f035a0cca777889640ef2694142dc367d7b217265b98739b7fe7f530c95230d8f36f5164
zbc6976039b5ed9bf654bf8012f85a172d0c39cdd157420e7471d405bbd8d8df081b88e6116b313
z81cfd2eee7e62e27c3f392e4a535fb73cf5d421e0456601fbbd397e296fa91c928b3e7bf9a140a
z33ed5bac5c00475f444e831df2d085e0a8c98f26455b0fbc99c44796dda450ec35266ed06f6349
za9c49fb4737f92b2f7928533d18f231a01f554900f008f4b072a02e60e6f0789ce6a98026f8bb2
z785e0479bfef64db301d9ea3010a3657731fc7ac890997ea9faa20dfe3a89b43cf33f3eb5cd2a0
z1fdc3d592626d87863e30d5b4acb7d9efb3032bb53df6572366f3a57a420d742cf871efdbae0f3
zd3b6daa2ce9734ae7ce79cdb1df27b725381e7195e401efb4fc19d8181b3892f62b21da2dc5ae6
z64ec949d81b242954d969bd206fcf113c1474e90cbd3f93535fde79922e6162fd3d24ea003af6c
zdaaa589536dc14d4e54da54cd45b28cb59fdfb48440dc1f1446ccae369de41bb8369246ab5e309
zb2c31d39b2d4472f165570b1afa351faf2c9e2c51df33822a8fa5615d06a83c524d99add1192cd
z9683f58b8f56c7720c4d8dae78987c1ff4c4ffe3723e9a37345903ff480a4dae22ccec10fdc9c1
z5bd0ca39d73361d2b2353e91a353015118a33c2a7b65710f99cfbad8d654cfd3a13597cc7e029d
zdf62d2e7a6580208cc39749fa7ed1a27216d1c66b36eccbcfb5b54848fd2fceb98f061a38c2a17
z82cd12f60456064c559920d4fc24b0c200e16002c8c6be8f3d0d46b5c0babfce39c61b5db816cb
z8a034fbea01af80b6438de823fc786b1d14770cccbe6b38c73819330ad0751d3f46c404e8b913e
z38eb4dd7017a391e966a165e80f09fa86ead9c62e3bc7325ad712700a98fe0ee49731107487e49
z54844d85bb5a4f1828bc93c162580ba3a50f8f5563e24b27a7d0b890614f70edf88f27ad8379eb
zb1bccbe3e318a8ca2d99249eab6c297b47e62d5d6618ccb4451179c3ee52288d5aa429dac15b2d
z3b3f80fc5ead5424017a71fc9a70e53301d3f0133d654bafc6783064ddd0a4b5d6ef815eade264
zcccc3684b3ebe12663778b005fc4e3e103021374d9b03989dc660484110180a952eee91ce58a0a
z0ea3f9049b3ea9ae609d6604024d1be48030e82b1c9e1cdc8a7139739bfcde3788433dab7b92e9
z0f0da90f66dda16c19fac803e4a5a065354f3a250dd27ef1b656f4677057d6855c074c20583153
z8c955a0c82b48ac6142770e2e43ba738a1f43771294f5e94f7159fe2939317e768482e765f7c5f
zbfd9404ca90f529ab5ecb49140fcfd6f69500cbb30c2428ef979f99b85a27a0558cdfd7e803e7e
zcc5cabaf99bd512517c32f915cbced285b93252a8f41b9c6b9778275d06b8e19e678b9820ceffd
z4ecb247b3f118fc1fffc5055f1722bf81156378802111cc001b93cabe17f01065439dc6c155b55
z68b43f4fc3734ff0f802bdb83d18dd5da06cad40ce78a5777d0796c9b48298fd57b7b8a28a65bc
zf19383f0043fd0b65279fe07a63c5c9bb12e029566cc031094ca5d59dcd8337008d384339f4e51
z3e53bb69828483ef721b8b241641b9ffcf881efa1ec62cecd9e3fe2024aa29e118b3cc0053867a
zb9728c15b991bffab6c9cb8a94745720ebee0603453d64686fe09817b820332d98648615436ff0
z6da04319bd5fcb12077257884f2352666a8f864dabebc033eb693f8ef0b749dde1df6ac8f02636
z5db5fb1bcd68f8d4820989d8b4f0efde6af76c28043b462f3fc1e7186f5f7d9f6e28aa88dee97f
zcc1ad439bb7a7b1a39a3aa1cf33f097b1571767ec83950850fd1b688e588ecc1a26293ee78347f
z32e0f1fbb12ecfe3f981af72673ffebeda17457ad6ef9c9792546d8351a1ce1c5d06c0d7170f46
z4995bc482aa4ab737268bc814ada0c88fef8022e73541e83396666e130f3d7bc9e861dbd6c25b4
z77ec85c5e75e0b7f39149a2ebcb6fa1074865c6aa6a16e94626ebc3ad10fee4db091822005ab13
z24231ef626fbedce69293cadaa7ab1505c8dbd0b1288361da459e0d850187a41579bd08dcad494
z18376d2ae1d78c96b57308f79597787b9744ee438eea4a3441e3b0c53fa2a87ddaaf2121ffed89
zae656963f13f62046d61f89fe14c4e94b388a9d877fc44683a95efbcfe3f645d3e348ece9a755c
ze1e3aac07d414cccff89dfb1cb5dc132c9a60d4fe148f279f42acf9842d6a0926d0be70b98012f
z36a4e6ff9fe32915632320849c253915edfc0b20dd7e0c512d91d08ea524fe1c5241ad12305ce0
z5804e4184a17fd3b166e03db480570ea7fd465a5effc5354dcb4f17898d9e129f8d2bd70db93b1
z1b7e7a0b3b60471d0ea488a326033159daeb8a5890a9d16a0ba931e7d084d6937ebf11b5bfc0a8
z53cde808615ef420b8951d332ad4364bd597a0a2b6a3f5c584680ab51f097fa67a559e762bf716
za546455af47c385851bafbb2e1c5598b0980801114377f1db136fa1db6966e15c49f93445d7804
z4dca4822ad6ab10980d8a7c8dbc3405b231c633fe6fc55cfd4d4f7f03c1e8b257106c63d9b9606
z59cb3190ed4cf6c888bf2bfb0e06037f0b86bfce2dc6e56aab5a96fe6fdba62e8f31cc61d053ce
z0f1ff777460cfb73d79db20487d99d6d42f2b63f11cad1f94bbd20fa830dea64dc0ec9e69081a5
z97bc0377d86810f8f60c5b3bb946ac7b24618e9e6ac1c27be9431eb4ff6cc3988011e86837c837
z21ae4372c2943fca9e58a15ffc0bd29028ae1716752e915e10ab63ceb60932957253f85a2b9491
z4ab3aee9117ebe990973a301523e8242b88d034ee22be911ec1052194476868b4cf2db0cc907b0
z015d5ce0558126800e32ec84a61eb409e6da546dac8adf1f89d1ab8ef88bb1e12fd170fd53bcb1
za20c36d8e26e90ff59a5ab2cc1268572f0ca42ca6096a71a6190ac3192e0d0fce586ef70a8d6fd
z3491dac308a52b151381f56d282c756b716845ff0cc16cc5a7f7f8f960edba84dd2fa2be879adc
z1c0300909507f790706731686e861a4991239a6ff4babe11994cc9ce2edb25816bcae80b8dd7c6
z9f4eab7ea45c19b2fd6639bd93ea3248f3167b88a6945f0822e0b7fd372b1dda3250d46ae12312
z163437f053a12bf2bd8c19ba62bdfc18fc56e10d13259b04c6a85dc9519450dd0606c985b4ed34
zb5bdd09b9445f160db61a98eafe991dac4249137de5c107c7d3d9d607d759ff8f47c943be40b45
ze3cc13908b69c2604019253d480a8cb5359b4dd9556f52b0dd2e3f80ee137ded5cecef9c3126c8
z2cbceb003f310b2de7fc9dd3d722abd3807654f1c4b14d5ef096284c306aea4318a0052c530bf2
z6a993769389829bdc7b5f62fb1c3c635c3663739fbb25e750a380e370751abb0a3c37323eb0b84
zc3241655b3ffa219024156eea5f00bf5e9d772763f8f4906d7ce807a316a937ebaec3cc8956d7f
zf65e629e595b27118a15960735e5eec09ce75355e4471d7ce609cc41d668eca5ecde0fdd133635
z07843fb63bb09205a542b599239337bf8ad1799c73a34a6e08c61d69751bdfa0e1a2dd106f957e
z32812f073c76e305c54fac73d3f86090d25902b895859f318b9d60b2bdf381639bfc7a8cd30a59
z375a7752128cd5ac4159abd07b767f411e96f9c67c623be2b1df2dd03c6bbf773fae9c75ffe0f1
za995800a844690d185bbac3eaa02375706cdacccbabc7f872b3457ba44abdcee7c241762ecae29
zd4bd9889b50308b243d96906a00486e9df2d02b85d3ac1a46901d0f9f4209909e6a3da466c44ff
zc596d940b9b390e8280880960f44b77cecb1c546c0c5df9ac3319f8beec57619af47102ba1fc31
z38f653a232fe4c05b58e600f432414f79d8c32c5f58547157190f84d3d718be84aeb5c3bef5f3b
zd83e92463f9943f30f21fb181e5f1d10126705f5c120eb8ce706924b363ac53928f2eafa0feadd
z4a80f017ed5fc96cae988cd5ec68867a32874b819b4fd2178995142e3c0ad68e68b53092661230
z8a431ac1db1e544b9a122e8258087c956e021b6f9666f0138a51245f712a10b0ec4f122d3c9d35
zebd16172883ce97147e8f3820fddd311f631cc4fb11aa6f844de70b988b63ba826a22b889c89d3
zfbbcd4d7a0502783d25abe24b339d7387d81b054c1426dddb33033991e3f863773f094ea7eb8bc
zd45736257e40d9fe12ec4b0a40460309a085fac973b031bfd099777a0137c4077e11273e4ff6c2
zb2ad13442efe67cc81d5f2b840e384589ea7a5da0a214b47c6369a7790043db1430708f6ba66bb
z62247244c4a5cd38069de4c5c282d3d399d186a52add5362bbf5607a08e53c653cdfc48b2f808a
zfba2f4d9bf528d3495fcb4ce68f253de1d88748c92b880dcf78897eb83a89af4640cc26673b612
z64256abb209e407332aae8336b7f884a8edd0ad0028c8ebca90ce49bdec1ba89e9321e57904804
z224ddc74283fe8b3f68974c694bd2b5de57b44305b8daa1611646dec0090c6c134a8563df28862
z18821e0a75a6f0d75b20465b740cbaefe3a38f70b2ee943f2bebc0f8865bb4b22ad85e63f38437
z9adabd1804d9d5a656c0f83607482813d836651caf878273bc475eace738a390bb5e52a22a1dc0
z4b1bb8e53ffffa8519eb43ae58939f7a5c7f2f8d516aabe44c21759211ae2988755a227fe27974
z50155b2e47f817ec713ce2817970f8295d7e7101bba5be8265a7dfe99d356914d63f3c556bca2c
zc3eeeb5c880ba885369bed2ad5cf2f6c6805ccca8e987dcb325312581de682809ad7c68b8f0546
zf53ef69e14244f0cce810e00081a5a6f7c6bceda66595fb4a1ced19ed1594dca757358e4699bdf
zf971e4f3215648eb1b21ad776e3e06d298d1c64888002adec54e4535a660e93cae4cc8bcc373a2
zc32e9b676ae3552688e068b11ec2c8386a0eac34195dfcd25fa88763c3bc66a7c374bca9f83c07
zaba24969c4d4013370dc8e1661e0ab0532cb582c34ef2c6464c4a988ee10e7cfb47762de698876
z854bf322e21e2b95269cee27c097c1bf8fe7e0fcd5376e607fc0af3181405d484c965272b11ae3
z07c6a9e19029c41ccfeb16cfb1ffaafe553c1424a33e72476433c748d7905b881720f3372da69e
z569844ff41972417038c6e5789f1b88bc065382fb7832b5c30b835b3ad8651c2fb23428b590a5e
z00fb85c6308edd25de76da18484a665dee2f860b59b5ceccdb1a4eaf54e1dfff0ae378a465d803
z377a7adb324beb961c0b71b9ef3953038eb2574b11b0a010f0762e254772ac38a23e85864c10d6
z33b8ecf6997483f2ebe6edb3bb529564fd73fc38a876f2b03cccd06645860c79f7e4f4b8661c8c
zf7ab4704d36f83daca75e14c1154f0fc934f05ad04644230639047fc18625b0f767ff2d2634a70
z3a3a62681160bbcc99fc3da6c77934aeec8eb2f5bcf35099cdc61d1d1078a08dfe66395328ed8b
z246f25bcd8e863b68096924ac3154c7bc91f73079d8455e113cdf057136410e24aeb1c2feefb74
z5f2371e31a0190fc95df7dcbf30eb3f0eb55237629e1199c0ec09db198efd0357eebd25fd3b5c7
z825bbacc3b696aaa5221d95033abf98004f8e21b09db4a43f6d3433c2afaa5e6f6873a690cadee
z4663f4e31550cb919bf47e7850ce2b9f028a54a9ef78837a7a38d31c4b07c70d939958804a8190
z350213e7de936fa28f75067691c31458678169b6350c4b7ba1bf97424ea6a925cef0654410ca98
zfa2c4452cf65979e18759ab3a592f4ecc7d02ded3fa7f4a687a5181fdae9d55ee913b632ab37a1
z5863a3512803cbcd718ef43768c7bf0c6c3b5f7f98bfab553a8202ebd3a80056d5fdc4946ec1f9
z811c009b4ed629b611beeadbdae4e0c53d331317a5fd009278a43be51f7b103e6c1ae45171e0b6
z5949256b03585d96e61800ba3fbb1f570756fd7e019987c49e519b97afcd72772fe67552ae2d8a
z2aef6b9c88273b57a46b8295a564e9ca5b67abbbcea638bb13f865293ffc803eaae0ccdef8bea7
z1cf5e5c2754289bc5227f53caaaa769db26eb2f12d821ab1920fde8102d57a08c656e543ea84ac
zd85bd923c7e7a5a3094b44cbafa14fac3fd60e5a519c4170c164d5d43085eb7120b8d808eae995
z6595c3473edc8c4e492bf19bc53662e7fe0070a47c96e735a5bf1edf1501e29908650606d18bdc
z8674731bf52b215a48266161cc4eab18a56c901da9778176d7a2c89cfb66aa648cabd3a696dc5a
z07d58663cb761ab821883cca19d7998fcc6b31edf8771d8bcf08e83f5ae2eeed3273b9b1ecf01d
z4f8fe490045e253630d1ef3deeff02de69808224c676d49d9030a8a947007d55afc9ead674496a
zbd478717cc1ef031bda3f09bf4ab3346f2aee9f4088a62964807beacb2c54436de5225106471d8
z89908e86cac723682e2c272fc47d55aeabf1f73367a381d94f71c36436cdf0080df94d3022fc43
z70677adbde0186d80ab1de1d3a5ed98ed0218fb5d1666356b98e68afdbfed3b28f4b12a6487c61
z014a91e1b41090d2f1e9046f0df4584e56904b9e2842d41a4472329a445f852e75e6791352c6f4
z26a45b4a33a9abb14b6ca9954477214cc45e83bc9b3b8a7db08ffbdb2ce71fabab33b7574d6a12
z57541080cfede1af62bb1fdb3aee04931326c0026529032bf75240daec0062f29cc5933127cbc5
zbc6d16c253a5c11bc5f8c6c6ba4981a6922bc8c2e0b1055d161e635a49e2928fa163ceedfe6091
z71b2e20a3c9846491da09b0658b3e32d4eb7005215477f901ae23ca4dcbd3c23962ea963a8733b
zf72cb1aaa0dcf8474dfde471a9ef5685386b3deeb256dcfee947d2103137fc58ad5066134d4ab1
zc938e98437fbdcacd986fca046fe9707966319d1f9b2db1b7e2066de07f944ceb52bac743d0afb
z189a91f13c2dcbe5e99542592124c9107ddef6f354f17a5f8a3995522c54eb4062eb43de4c5bc8
z8d5ffdfa6fedf4e952f3e78804e7ebc70dec41f368d5024e078eb14a2641cf25a794dfc4b074eb
z7efee85f5527ea04b74c9c3f1594a83c6948d34a2c8cda934ba07dd6c41dfff18a68265e5bbe53
z8c58b85c81552b7964d3da62acfcce757c10a6ff8217b3201b150ffef3b2dfe4c04d410cfeb39d
zab251e89d4fd24b2a86325e773d7a44a42e03aaac884b23504c22f856b4984d65427b09f1e6fa5
z56290db8b730867ea49579779e68b0432f6c9729060fcc4fbc7334f845219221e85c2fbcc38c3e
z07d9f72fbe70e8e8d6f2dc5fc93fc6dfe379a666bc41991d878fba1e250b3acf7beb7349c3e5ce
z00e963b81a65053be3c0dfbd74f159c014d5c81a3da1d58b02130ceb9e6dfc22bd1306d5caf9f8
z9bc04412cd6a0f73a9cf54667a74d0416ff45035fefeafb06479a2dca58d00b0340687c01cb9b8
zaae56598d5bd6757fa56d13f831338d6619f96f06ac0b85196ce2cce465e0c2b76d8e249bdb009
z09fa0ea218ab1e4bf7ec901016717d0c24eb4d623892dbae1362d21ec078b3ff932cbb09d9a9a6
z175f6663723abf40eeeecaf5e737babe308bb79ef4c32772aab6ba7addb3b4e08deec09a59981d
z4a93276a0ea2ba0d9978c0d46801affd206b29d50412398483f8f0018813c9ab60e979a13585c4
z25d23ec4a53e0a3350c6e5fc19b814c08a76a09c75510699ab0fb18d4f7219f41e7ca96f3c3a7a
z8aa4d6bb42704abf6e7f4d2215914fac25d7d1af13d8fdeb10fdd17a7c190630c73ac62288545f
zf8c0fc2743b8416eb9a5aae03ae6b5c558b4030c7cab1a1ff885dba6642e2869f6aab06dacb3a4
zd9cc832bbf641c5e0e7154f1d6d89f2eb73c69bccb4c66e0e22420cef938e2f2dc9f41b75969ef
z32c02127f5addb7a8e5590d162786f9626d6e057668182fb20e418a9b33e573890311d4bf1b767
zdba3b174aa9477c8e70ba1669d79c9e3afa669b25c2e81071978fd7e630fa18a8cf5bb940e72bb
z2a2dba97f43cb881c7c04dfe85cae854fe95b6f463caa58e791be355861472f21f3b947c0a63e0
zb88c66bc65c8b563fcd1b61a2119c8aa3972486d8145b005e748987ffc5d9a1b18131e124a851a
z2f70082027a64d8d56dc890eafd404446490c4f932e390507ec307bcc663e2cb1e7d61766ae0a1
zb6748a83bf4619f36844e182831c26204a10f0b9eba5ec47862a2b7b7ed2f8216d2cc65062d6f4
ze854503fe45361f40d025283093b4ad809e9c94adf9917cb8a104387326af6c2eb23be28178b7f
zc48decf749b21c0f313178358fd1534795b9369710333067949896d0c819e3c5d868d89574e5d2
z186c7b1f92c9dd944da01cc406b6b21d58d3d5000a637196e72a04c9613818836b7b3c02eac3c0
zcba35c763e368db825577dcc7eaa58c247c12fc217ad1904e100af1b351d3399fa4d3aafe021f7
zb2af48344705efd6733a3cf2054c150c346852ac4afa1028148ad42feba9b533a8293898a508d0
z0e4c9fc9f7c89471e30d177abfbd4a7e082f44bd60f6596260e2702f064e6406851242086f0013
z71c82ba96a9e8c3d88694d9f7ce834b01b826c6ea01b6fb0cde00a35d62febd8ff7447afedeb6b
zc5621e6258f289638ad9697cf1f887695d8b951b29ec2a1e525dc09002952148a1935dc1b0c96c
zdcc2a4260285ad42d87ec7233473efc16e6a7cd1505aa2ebc81f506a1c4d72cf9c17554ee6c502
z010207a1dc7e62b2143b7948b6c9931cb9bc5aec5b10663fcc07c9cc15e8a405c240aafbaccede
z71dc8e82059314fc5d89954d31474727a854ee83e969d5aba3b4637c427af5a97470076522203b
za3bc38cc25de8288be9fbfb9aecedd2ac01109b9167f6f7ee7f3762940e00599a85819f958de84
z42c039b87bcabcc5b04ce02c8bc254686ed53993345cd9234a7a4f8b8d9d7a21a5c8b0268a7abe
ze817d341a2a3d0740477288cff1a5a1aa711979aa98b8ec14a9ff5d869bdf0681050046971b4db
z7728aec34c5d07edc90bf9ccdfebc78de34db2d18b6cfd547c6636565ed1a1e3da725eb023413c
z077672bfad4ed91a6d6329a24c3c8b34c0e82e02da303b59502226c23f1deeaaae5291ce87fcd2
zb6ab778a986a0245246a329bd5a661edba2e18f738fabe5f130f3ca64db2849583fb277aaef502
z12c06e95c380ac533e0caf968795b0b7415bd0be7f88de6ae2f4da52ef6d041621bbec95681b3e
z4f6f30dd942b52fcbe3c145619bb5c8358e6c440eae9f5a1b5c99f8f17ad2e481eb695fb647eae
zfe9df6ce6a453174f4c1eb0b30a7f05d11a80febf20934b30da5f5889fee18890057c8edb4fb4a
z6a7455688066b8d5f7c3e1dd5c9924dfdce9c95ab5b81dd2b385750e67daab52880f42dcc0ba21
z13bb766d0e1684c0bf7bfc01eef718863c7b35fbe0a1ec5ffabe79645aa518b81c7519b68e838c
ze95b3f5d013e7a4a65cca8bffd3e7f0fb7654bc02e64f3b9c4feb61b9c2b89301d4f6578019902
zf2d0e140c5865bee250dc4218ae5407a17924cab8eb3c71213a922187d6368688a56bdbb16d0f2
z913a2baede82aebf449149b99051a9f106af997b9473d9a42fa3129c450033b9c90bf1b8cbcb60
z271e15528dc45cb5780bb41e1506110dcf7acaf05db676605b8ad6b3e9a95ce3efe9dc42404c50
z3906ee58e7bc3aad25177b56f4862ad991771e212d9c815295d2f73a1bf1f47eb980fbacb6b09d
z7155d98a154e1c45c69e0ea6092d89db3db93f448017536d20d284c2cb3865ff6f1e34e8da7a76
z6466eee98bdfcf164dca3dd35dd4878fc16e90bfab46dc7786738b620b3f4cff7db350e9f86306
z0e82c513f5dbb5d2fc2dbd9adadae30cca7754e5eca0859a830ba8a395088a3aef6332e26f5a92
z753cac862f85004e32c2f8616872c4f4697196322c7c23872daa603cd47d1a55d87f77476c58bc
z6ddccb606f7c9f9e0822134b7c658a9f87d7439bf1d2461313c3ac0f51f1e27ae491650d69aa1c
z2e740a8dff1b5ca4790ec4483d29dfdb8acf5fb586622884333784a5c05a66d782c2e9acc1b63d
z19cd48587838897985649004c0e0f0caa9db0aced34aa3e5d5c19c35398ee281dbe4bd6857aa9a
z3357c21f4afb974b32014bf7232da7716af9185310916a96a8717d8a9bb05b426dabccd512984f
z83b546305072a7e2846e58bc1266b74e9e56da548bb5aa544214afce763a1bcedcc585387849a4
zde2c81b2bc4c43e37c0911c5fa150635019c0a7357179037a26c9981673ceef63504cc32711842
z8bbecbf1a454cad8825e198569188318bd56bd2a4f1352e90688f209eb7ba38d92cf3afb06b243
z6d39651ab4b601c62f460d9ee87552106308565537562072873513c95eb67212d6ae3858414082
z097e16e8f7e1574e30c6eca376fcd53a93eecc1b34016ac3d1ccf80136b9a9e86bf6c1104d4b27
ze99d6ce55d63db7d3d078ada532bdb40de7e06507b4824e11f39ca086e8e18bd1e5a3b4843ca90
z6979c4e7c714f9937a22376a0b49b97b49308895d62a1f15d7d76f5831871cea6efb50a127a31a
z99a4e758a29b9c8222d1f2ded7923c782d5ae4454cfdc2bede6d6f599dc00a066806bd9680caf0
zbe62ea7076549ec553f1180f259b8faa4f90e56c41197daefe5b19daded90d930ebf0e58ae1b4b
za54d6fda0c05322f5f2cf46edef77782ff5affead41b27bb8f5a87af237282a2d9effb002e0648
zab871b7d23f9dad174035c8693f47ca1a07925e7a0aa33fef32cd4c819718894e1bbdf13ea2962
z86b59dcf7a135b960cb4e3e007a6c9c9727ce2cb0273b02ca47c519cb7af499156367a1692e7e1
z7a60b59c52294c6e69e69005da7910d54c99bf38ff3246ca6e49971efd2f38e5227135b36d70f6
z70b20f139d5adaebea1d98f25825bbe809242d3dde2c82a69c84189cb63b32ef2aabfc09844227
zeccb61fd405436caaedaca5ac4010373fd1a5c04728fc8848c8b7b205a63fc1cdded76b495d6d8
z2be0d14a001665732b958323e2788ff70ece303c2e76881c1f6b0f753fefef6d0ca7ea59eeb68e
zfaa2457e543fe72f7b2347f7a1766ec6777372488bb801a557784001980d56f74351fc60884060
ze4a5f565161edc6aa614e03dc5733bbbaa861ab86660d9bfa49e251880b5f48540ad4e3e7cf5d7
zccf0e71f5debbf43f024d751899eb68d889e7fc9741c474f4ad7b1b1cf4aeaa46ddd3ebeab5c2f
z1e8a4d04d9c79b58612bc058ba5fb544280f5aea9f522ef7eb8018c27e48cd526074932a540e49
z4def0f001034a8fc74d3641e15af28f65dda90df0705b0675d0599149cdca47e62dd91f76cf48a
za31545a3001e434ddd5fb5e8490d6a1262e28d632956a01a5254e5aa63c702c0b444101c74520e
z7dfceb3e647719af156fd510af6f7a2d5a28e13e87ff594be0bc7d72e6a2ed51faed615e5f4b4e
z11c025728bded5ced61653b719266c235dc97b60bb171dc7b271be59fde8e8dd05117bedc26c09
zc640ea13a6910d20422f4f14aaf77cd727b1ab4bc86e1dc48524871a0f54c376cb0a235db46c73
zba5ca1040d57bb3e9e3de640819c71def6699ef7ddc00dd83c2b99d0278c7808f5e9b1a997b154
z0647185e879a786f6009c106e79fd2c1b000ff4ab00bd23b247ce139795c9a1261f48763e9015b
z0d082dd29dd7955851597f0ece1dd920d2e48adddae8d955084c01e48621caab02159c745dba7c
zac00fbd5c3fb0c95fac46213c59a11fd8d454e4ef9c35a8377aa8ddd00ff654a7c82bec5841cac
zdcdac7ca1bcbe151df7bfc6c634802f0951428504b0ecb3f793fbb8175d2bca52a1762a957035a
z9a5e20465589cd47a0d80bb35b4aeed48f1d9d75ad79cf968c4e4958c1e9eefe0e20baa7417fdc
z5f813278e4066e959cb5a6e5ca7c1f048cd6c47779d4bce61f5452280635bc1ce3fa6d9aa1b753
z35750771abac168bed4cdf2f950623f57978fa49067dd2db5091decb15305646b273381c4a2600
zea993656fc43ea4adba1c299e3cfc8edfe9402b4948da19058a3881d804140b03471d61a46909f
z825f0b1ff44ec6f91a696d99f872fe14ed9c41eaeb098264fbf76edf76cefcea4611034f5a65b5
z4b249fd2dc404b8fef30cba7e135d950e48e1a40ce646325f6cf37e18b4cc260d0bef9269c23b4
zc2b4d0fc2bf3500c9326898d1ee38c4201747fccb6be009ad779b6b90583ebcd6d65ba73b8ca3a
z61fc98e0ec81f1aee7c9218000f666d323d6df72f1ff1b9148c7cf5490f4e2616284554569452d
ze979ff0f9122e3aa894e43609a13cc59027ec42ced16a8d8c250a3cc99e51a28cd3beaf4afd502
z1d2e8c1a7e7c88348ef2841fda68d7cb7cc5b3a5c5a3b5ce6bb79d6458407c3111216aa45feba2
zb12d0d59aa0d44bb117447cf200c9013f3ec55e9f3c2a97504cdf77ea3bc91f27f988a6502a290
za3f9104686ead157fb1e4619b79c37d5c012d9a895036f547bdbd58d9a05261c008d73f5027392
zc78d44796418b44a515871bfc81495d62c65ef54c33a89178883073ef9cd80575ead3c4e02c86b
z89233b2b7e2827388a77380e5d5a4ebbe320fbdfd879e94746d409faa8a0a54f091ea517f32d42
z3627fd4200c0919540951bb9b3985a56207ce207dd48b05198fc3322ebf2f8d94bc1164fe4812c
z2c9132524ee4f262c949823c82a424b261eadceb34356897335f638b24e8ad1922da14631aa06a
z685e13c1e66904aaa833d8ece1e0756336086bb3da1eec1a71e2b81089545fb2028483f4d2fdea
z6cb5997188248f11d7c795b64fbcf3219b2358f8675590fa32ee357697754c0fdfc3f34000b998
z35316096b35d1c81eb66ad80d88995ad7352d73c2adb6115339d4f23fd62b17be53db7d5b995c0
z137b11d3c0505164cafc49219f01b413a191d80fcd09c1d4f2c162a947c46a2ea8a7a4da57a11c
z4f742c8105c2af6b351bb3d1e5a6b1ddba34ec7c27482a9cd1fe46b4f99601f1f5ee696df08ae2
ze92529651c9e546150d5bf8a7241919309d32c28eadd4a253c4f1b434f63ab85e209d096af3556
zc599eb01deb585d0e1368ef25389e190a3d146af565051bfe68465ae815a747848e09d48e38dca
z2eacd20f50e4a3082430b777cd0815726ed246f522e7b7def9fc3dfea9a917b964e5a763525a98
z51d3aeb435e044e9ed95790d291aa4d5f0a3aa95fa70bd16c6584cc62c53d1d35e81d5bc55ad53
z43f22501027a0777694229b423b9cebd3a3b4c02291f298dc1efdf03210156479a7669cff39499
zeb4fadfbd8657edb5f5980235a676cca000e2aa5b1bb87d0f40f7bd2974bf77caa10176ac26bc0
z8ac21c2eadc1b82dcecd7b9ba8bbcd15779d5dccb93835ded68919e4c7f7495082011dd457bf32
z376c32e26aa33b58e910d02b68a533885d2bd3302ec2c5f9b71ba44788e952303cdfb8b6a1c453
za6af7500dcd3c0f4536c27ed393e50cdfc3dbba640628b8507568a0460badcbf22069891612673
z3a84b1addc69a8654afd2d17a01bcfa648dde864488036e647e54b3cb2e601917e3d582f40ed4e
z1b5df3ec86962c3f6f18e4b88fbc67674abd34d84f8d54ee92a645eafd6d10c14cc86faa997d28
zd3007af1f1195fdafc512895d3d959373daddaddf7050aca12842863a46f1a85b3b94d78c02b7b
z76e49d4fe450b5d7e6360b6591d933ae1045077932bbcaaa2741ad12ff34c2b1a78cb918855b24
z5dbb98bcca66a21f8d2828406f6350c762179055ddf8144ae3e0e942abfb4ad5cec940bb9730b6
zddb5397657aa368b293b6cc093c18f77388259afa3ed3c38345fcdf01cb900bd0edf471fd1ff76
z7ec2228eb955806153f59bbf766d1f18a69e83619de90940dde8e9c3de6c971874b158b74a5b78
zb2b8c5156b06d0fff902294ddfc8fa32e95969613e2b3f48d142228fb6f87f28c6292750e01e6d
ze433eba859ece2640b13f11b00cd88b2cc694c70a682aa69aab7db27c954b8fd7ff937b6387af4
za8198ec4ebbd3165b1689d7bd67ebc3997cfc5307644d8cc239547c651c6c7b49a976162c133c4
z71fb80651afd413dd41e279c28255d4c4f0e88e77ab81d985361eed6705e231cbca6cd5b67d65e
zd7480c78b88bd8856cb5de6cd635ce5c424ad46e76b02ac0d2fa9908d6df45160729f07bbcecf8
z6c0fdf79569aaf13cacada9a142ca6cb637ddcabfea43dcbc3d479a134cb115cd5baf462f441f6
z72e577b44756a84cba081ce3718dc1dec152a1eec56575ff4fa0e647d7aa0a5f9e2ed84251e8c3
z2e28e7d79d1810202389f694b2f347bd72cbe8bb69b972a0eaf4c5b63ff29a2cdd21cac0c47ac1
zcbc223693e3447dd4d10f3734e69f5198603595500062c5c67fe697f1e2f8434c5bdf3707ce497
z26fede46ca0caa11f1fd593aa08eb22ca621e0a0be5a2305b08c24ca58e3640bb9c8d8c84774c2
z55ccdbc991478a935ae5d4ec6278009ac2c150de4377b7014e215e3d52c9689a0aeb30e783b2b9
z8a9d4c8ce77e707c6677d873851ea890f50a1292e348032434f9a7b4c9c09b676a2076c58f4e04
z5ba43c3ef810803ed4343ff802410bd598cd4677452006a0b640763a7e6c2ab7351c86c0d9d916
zeff066c772bbff782ad4804aef3752441d6490da1617c5d9ea5a1fc5c5be9b1fe321139dfe2012
z05af93d2898b7abdfec5341dd72ab91596a528a136b9b1d26cdf97bb6a5e225c596a78cb04c111
zc02bb20059a80a00a515d80bf8ca5a3eefc7d668aaebfb9c54f738e86d8bd1adc821a0b460a2c4
zda02fcb819bcdaa6065ad601d1d5ac364bdff99421795f051c6e72d486edf9910f81089069c74a
z6e0171f29731b1ae1349732209f383cecce07718dacb60da76870703d0b33b8d3a667057ef81e5
z3a4fd0bf839fcd197e3578bcf6b44c1d2e7ed99bc461286008905cec71e98d5520fc566cac9de4
zc064ce3661250236cd68c178c211391898bead247068f2bf78d947182496504ba0827d98825877
zf354d764e317522f4f96ce76a5de0ecf6f5bd3f8008a936cf24ea16c26b1db782037cbf13260ba
zd0e7837b69cf60c40fe80926ec2765a8bdeea53afa27347f9ab94380b2e17b479fa6e61f0eccfc
z4793cb74090aa719d70f11e81d6a31eb2c41e3e29279a62eca4c2775d280c208df25f2ca405f8e
zc4fb94e94f8305478b9bd157625d53c9aa785bbebac6911767b6d2d3073fb3e2084148638d0437
zcd0eedb470307588d28f0961ff6cadff8c0edc5f9408fc2caaecdb666bc4f26179640448fe40df
zb68fa1e78bc1f430eeeacda315d63fd54cdaa8f7b999828540a017fb71a151f5e156fe5a5670a2
z5a63338c88e550d76e0ee56b9207c03c2d3102a2ff37d780f5e16e313b71d27d270d752cc8b8c4
za8f244a8247c04670e22313ce1b21af556b5acb825356ad891ff3ac6fcdee182336546af1f4c3b
zeb866f192042cd4d4587ee1c2ba0abab6c2f8e699d6b381e27bd05d13683867f21a55bad5f6d3a
z89d66d805125beb2785dedc2701e577986289aed23f98d61f69bcb618c96b6e403c9a9c9b8675a
zadbd1fb83a9d2379b8b874ac2a7f0959c72328fab12c10c493706294e92ef75b0b33adf40a6a43
zb51c65d2c077aa0b0f13afea6ff65a0cbc8d7b03e509af3e47cbd46bead880e2d496e91f3481b1
zcdcf24c93d6fb554ed1922153ba84121e2b0b0aca4bdba557818295145028bd67dc7eea4e31d53
z3340137eb01c380bd767799c591de275a62054a516010f6fbb113f09393dc6da53c9bc9aa89f7c
z31bd6784fda90fa264078e266058079946cac3b2d7fc44c729b895897f5000771dbfa59dfb5b83
z6456124993e982d00b33c5bcdb00678c3a083df10cb4eb6cefbc26b7daa4a3d6154a2a36bfe38e
z381898ab432454b2a43b069d049f18ff5e4aa05293b252ffb4d63cfec83b0f4f894fef114a7e44
z39ebe51e223c9d3d8ea310c937b1f805b182fcf544f20e5980e3f844067ef12d47aa14240933a7
z1adc28292e2e72a368ae89906c63b1edb644b76e93d7a8a9261be4008809e2723a8abe6241fa4b
zd4c316b6816a295832a3847128cac5268289f23699a282fa12c3be7260440e827b6ac2acb6547c
z0372986c2da1fbb8f60d01b633e93293a33b5d8af08321cd7203dd71209eff47d9a6cc7b85487d
z51139e0a16ad5932ee6c3fd3a8ca8ad2f0ddafa09292262fa79c2d078559c02fd6c8a045cbfc09
z174658143050244182c0bd801ec6936b62ae4a37722e545d257a61f2c1c5e8b9e91f486d7ae34b
z012dc3e5daac71a9efdc9bcc6559018787f121d8e99e60ec18039c7a9616156a0638d1f263b0d5
z9bdfa55a00e7e691becf3de7a4d020fd44b5da3f800d76d7a115feba03493e9aac1749916a2161
z7f40605016aca7b14531970c681a7868c74cfadf7de7a733788552595701b69c50987c07f61881
zccf5f79d39e5acba67b1e1e928857b97ffab6f7a0419232f14b9c36bf56a076cd6ef3eb6ff218b
z49b74c476826ac93e32d042683db0331e7891323140df77bc6d979c87c4769e640ae4dd041c3c2
z69fd07fb87300fa5556814b4b07189f08ebfb727748fdf3b6cc1304ff1a5b95a1f094364901190
z7722486ddbc5f6ab6e5f4811f6d2bda59b03a4b10236cfdafc38cfc91b56a12937703eac36cf32
z5dcadfb91f74222f6bffbc89ab1e72c5d89b094eef054da1000c3f38eda3ae78a74ffce836eba5
z94b649f7e7dcde3dfb8033d96fa33048ce11bf60b812964ddf3e65feb5b3af50488844971d219b
zddbab859092255bcd36c100082f6cd0f2eae4216347f93d5201e77978f282323141f4b738db5b6
zffc08cd36ab5e760df37aa1be91b141ff30fc4a64557d240013a623d167a4a074016195795ccd2
zc15ddb474b9687d4fa23404f211d6989fcf88a0b3f4d58c3ad68fed53e9c1339fc55aa4253e235
z8458e7857876cd49fac6342b96bafa2cf30658763f8b8212d1ddd81e4d4e75bde79a000c0f51e1
z3afe7d7e2773fdeaf0594749796b7e9b9ad189c729a2527df4acaa2b86d17e0ae92955eac9e0fd
z05525ebb24896bd47e737ea39b765f206169ecf2feaa8d5c4f219802bfa7874f2240a71e9b8bec
z99a6f97889ee0926539740b35bd49dd08e8a0efc4fa44046e95ff365c80920a192abba4ef8be52
zce3c68e30de94fb93674db871cc634a0d7730aa72cad9d6769cc0d6f8addf903c1f2fafb676b14
z86b80acbb8ed079426171e8c74e30dd27bcc5fc313e33cbe20642b4b64ccc9b7212d9f9e1cad23
z5493169f8135cee659532949d54c4a9c2d6f078419a99712bd0b89651d7906b53cd13ac8e11cb9
z4cc3495ab5ff4000080a9da8cccebccc44c413facca91543234c47f3b7ab1f3c31506b0a23da34
z2cdf6b94a425dbaf0dcfd1e52aed61f7423e6de4e4992ad60306c8383c671f87e15be6c88ee6d0
za5f9dbf6f4b8fa39fa78beed256ce3607f321a6faad26d8206dc545f4a69e35c87168db997ed48
zf1e996d81d9916fd74f50c47b935a0b59d5a7988249840dc3a3d854081dffe34fa0b643460587f
zf8092e6dd508c1c83456522cdab38a19f98099a960c9dc620a1472d9116b803773d383ba6f2af6
za14d69c65619b02c5caccfcb3964cbc59b1f77d1d1536130832c661b91112093fab90d4bd2221c
zf022d0d2471ab7c752c53c57566507474fabf32bbf1e5f41591587f4d0acaa4007fed2f0ed2598
z5555a471b898f72899702add9d6e9d6079dc3a82fe531157651604bbc63b0285838052286c09fb
zb0c74ca464ae50f3d66292174dde32e3c0ab0f86a1f0f7ebc39eb370ee4bf29d780badd2cc9adb
za849d322394a822348a3e1bdda1ce7bfb482d6e464d86b4ca80e90ff377ed559ca710d70329c62
zea732dd33f9699f814883122855cd945f2910ce8397be3d0ab36bfc1a19efba7fa3d357b062fa5
zf0a851a303fa8dac488df986384e492238cc18428c1ab557bed4707203cf01eca9a57e51cdb36d
z1a5fb83ce8117b30ba943158ab8327aba34e2cfac1965986597fdc25a83942c67b66bb322212c9
z1330c6d3c62536c75985f22813055cc459022f903c3e42348d0a2ae3c1d93fc77694304fb22948
z4179d3ed42c98536587bd8ca0dbf986fee24b3e7da0a65f0765fe3f1269c658880818d1cf6479e
zd69749a258b787bfe207ff9f7708e2a455503e077765a1a9184e1833a9431ea7617d2412c038a5
z1a1e9c6a0128a3194dd65d5d41388e35e6733c69bc14c9a749855297befc4ab39d2688b3e464a9
zbb66ed78397dbb4628eaa36fe0dec475a3dfff6909695de527121eb4d708b16fbe6fdcf08ec79f
zb6766b5eaa62938cfe355f1dd35a0778ca915e6326fda4cb6a2e68332edce81602e3972af3839a
ze0c2b7354ee35928258c4da2abd22a9d2958ca38f3c5e055fed42aa4b22614cb5fa1e5cde4ef24
z05a8750db7a65cafff8fdb63c1854140b4afee5382b1a60b7bbe956bd9ccc1b54ccd094e558190
z9e60d18af419714f916f02cecc64bcc1406f5cdc987c363ebb5f726a0e8739d0b0f4b6e8fb05d2
z417475abe9104403535541f1351d5bb1e4109783a0ef465004339898e361ba4043538ac18baeac
zad025913f208e534e3db54fdd10341cf2f3f8a58ae943af008967c977fe038c71d7619dd02d09b
zebec91313b9c1816b334e6c8ff9c16f47c59dd509feabf2eb1548ab5b787534fa231e4a0916af0
zff564b3988a81af48a8a37ba98ab963f67d2241d45b501511e8bc5525fdc4552cd62a7e4efee46
z0c456f7c7370ad3dd34c288d4996102cfc4c751d9acf1232c2ad8d5a18b865e7bca1958c9c13ea
z07d65c2e10a58a276be8ab82fc98f8764f6154ba397a80fbb7d652c4883c166aa6665401b72520
z8eefff6c77f979fc34f091c663672e4fa99d4b1c666ff5988931516375e676dff49f3630ecdcce
z4e588fb97d642c8abbe73563a6c5896d6b949d0d952485661373054a637f3e6cc9f67660ccfe52
zc7905d1bed24977a1d61f900da858427ee570621fb49cf538363a1ac500deb3467681a2f7ef3d7
z529428a5437215096f70d965c8e0dd307dede697b1c893aadf987c0ac3fa07e215ce1312884c55
z4e209e4bfcd12f885b05056586d5cbe31eba44cb3926c196eb9ca5d4ccadbbd5984e68a1aebf9e
zccd5c207017c5ac3813f82b38dcc149932d9aedaa636ba76b5eaee787a9a5f781957ba364d8800
z213a133169a376a9d57927d70b7a37ba7a563c1849b39743664abe440a0d9f7de7b061bb94b934
za131220f8bb7a7bd33b998dc88d881003ca45e07fd49cba8edd25059d4a8be2617c99aa90b37c1
za944b64b752bfc609e6e380dde5f36948e1a82f68db711f4d5d727497347037f5dd62e4ef9cd54
z83fcbe8f71f8e9ffb9345546842a179bc13a47267fe2eb6d9de6400158757a741ba44d97f19a8c
zd128eeca8e5a7d332485f2107637c181df2ff6a8eaf0c0541cafe9418a79cae034abd4ad0db86a
zfa663fdc94f42c02c02848ba5aeecf323f72d56b831fbf3843939ce23969d7556ee1c74ab20b16
z3bec31c3e44df507c032c382a91bc5e2593ef378392aac95ef2fe9e4200265160f740f1e17e5a8
z82e1e717502ddac71270adb276d51541089b2c4498ee2732ff818768dddac1586b9c490d893d55
ze193019a44252c2a9d234f0fc2b83b7a1382eb8b5cf2ceef5ab51b7e2253572555abcc3f62528b
z28f173441342488ab6de6d06be98994c784614ad84771bf48efc6558031bafa7259fa5bf8b0bf3
zd5399d0b3faccdbace28e703da09605978be82546e866340ef3d8f0fa6e942386403108d590c84
z04cfbce94a6c44c5476b74a948137248c9b588415133f223662432815548aebe533dabc8e142e9
zb5b5c7174a48ce1cc8a94b15a0e64a1f6c7695eb77d2109929dcb19c3140ec7ef839fab70a4567
zc1deb8e2f14b19e7a2571ae18627580bc305ec9fbd5002a1a0e80f20008ce34aca92365655a72c
zb60965580555664c69a4a38a0407bf4ea3b5230c8e8fb5f9be44bbadf896edd4422227c6f2e3ca
z40a29e10246676345332f8aec4da3ae83ebb64e30e71f9f745d4f67f34a61c357b4d2663006e00
z66e9c59d4d899e628787a52cf07ba8f72f8cc3e313e1fcbb53b91bd8401e70228f9c517661d6d8
zbf01639040a1e0a408c0280d63421bfe1e22d449e71fb8ae7ff7cb01a3840586b547eb7f9b1524
z0677cc56e14cf183f2f2fd828196b7548dd1e3337d773ca5ad74e910200da12938b67493d77d4c
zd7db2adddc7c9bceb9032816b3a23e03da5d6523e77b6f92d4615c3d8085989b0a58f0050ed2b7
z5b5bc2d4fdae2df01b9c1b27aeed8d9aac4937986c1250bb12f55c017c3d63a59cfe417dc74ef0
z3c9ca3a43b957c2573360fd12bd352a3b6e7bf46f60c7caa6e0903e531f9152c2a11c451137f07
z7e6857d5ba25f806be88420a232987404409d8c1e2642bf39063298d9acf5a8cfebb18ce78119b
z29f7f1eab233c18806205461ad99ddb4bddba99a4a1fc796af10689b23e9b057620555c07da455
z7910a53bf981acbbabf1fb655252799c534a8ddf88c0f84955fc924a5ca8131c269fe325713bf8
z62950c64244f65e4dac917a2af7b8ee45c326abae36ee5e72c159301366155c8969cfc4b84eeff
zc9826c4de374f7fc09caa592980284b8916812b7a8f0c09f31f25590696ad8fef426c37bd1a046
zd5c2ef79b273d25572d1b4026a8efe727e7406a3b09e192c4c5f096419e63a7854dede50b2e6c6
ze53310a6cb0a323600ad07b5f6aa10afe406779caf7a047c4b98d6d6e51e59929bfd59fbeeadfa
z5191dd90c9f4625531468a0e126045e29d8d0dd01eeca9997baea1402bbcd32669deec7ff1cc95
z471b402a902f527102a5665b5482821647d21638966581dc970fb1eed46e8ccd06132dff068851
z95403ba5363754ab4eb9319af640b422f142490598808cd9c8297c6ef3759d9cdbfd862062f0fa
z20f2af1134924078f23914a096d62bd34485bd1419b91d1fb312b38301e3cfe908273be14992c5
z9b9848712821fd16ccfb3931184e977cc13924af8a34aa76d8a2cd2f1a10c3cdca86b612772fc5
z35372848e4415465cdd09a1f1a0a43745244b659e205b54678b7e5a0b001d9f6cc7bc76a10a612
zbb87707e1627ebbcb1be28c443647e66faf18fd6cff6e3725f18e7baf260aa96c22fee3505be0f
z6ec12d23dd38ca03f3158ea1864c4b66b8a51aa78ff933d6884ec777bc285ad705c9cc1c1aa085
z129c9d5d699d8f33fdf1da58fd39bc0e25d9481ea4333fbbc32935034540d64435446db5b56f58
z38d8d0b92c90796e19d02acfb9731449640db9b02521476106d2cf3c64563e04aa77c13a682fdb
z708b17adcb36c425f8831a9a06007c65a3e32be95474df10d384fafcc56841e7917062bd91ae7e
z9681a6f69532deccfd684b2ec96ad0e3779e8da40363c4bff2b511264325ccbe5fb6d064327db6
z912be44860ef9a0f04028b3ef254823d3d0d6418fe5bcdd38885889fbd8c5faa1097fcb77ad458
z054d032dd02ef26843079fa52ba319fbff96e4a3218871ce3ddcd1f19184cfe74add890f03c7c3
z571526a722d8a77e05874d4b4b6a07b4fb7438ca6c80498e2661f29f2c52b18cb7f34c668eea7a
z63fe1ef44e3d105574aec1ac17626f08675ea04ae70710c72091126e7ef48573b948fd5ee1f477
za66e3749acc341a3db6c8c317a947a54c5940bb055e535a0e6965a11b4806911be0bf82a0adbd8
z4689f6c478077a8213bfa854d4c131a12b3e68a157944b94b1cecc91f34779b229215b61ebdc00
z1e819f3771bdb5b6d4eee1bfe46b1bf94ed536d545142bbc1b3d8c969edc7fff8ecaae3a89a214
z1880a2a861f3d5651aa848038afa2babf405a63c05456cdd24e2c359c498e2dfd12a6ca5661734
zd2db9389b2532c9d163ceb2554402f386d881b86f867ce1dc7ec2f9047979bd55493e00c349bea
zc04cdb9c3322a302ac868581bbdb19099eb9f3fe872215642f894cdeaf44e2d2d5b4c9c3e5f8e4
z5ced8114cd398d781405b50d12b260ec4a940da9ae8d3817bae8e236cc8c2165fce3e32a61d2da
z29d3332121a5617a9faae1ca26f9b36b23c1fb5b1e466c447293420fa12a93204a75fc6bc23596
z850728442deca79b54579ab79d90a64d99fa3f5a6f3bda792189d53d50c3be2ac3c427020ec449
z189c4980cb286e8bc78b6b39d1e1d41b41676d53f1bb2f8085d30757e122543d6edd6abbed3e5e
z21a51d2d50e2f8a1103ac578c6d99703afd55f12f281baf31a271c520b80fe3f389ec7b61de4f0
z2ed7f0b2393ca0d71632e25d7ed955938192dc499ce1633277601c6fb26ba9d446350a60ceb667
z4d7df9ba19dde2a3387d14cc338f6f20ead382a555b8f2e923602ab3484261088e79b85f128480
z8222927aa492ecaa461db3dea00319fb3a929d5ae77806b9a95c32c2a74742c47c898266224dec
z6d0c8d32aa5ab3d297048e76a929c9c25f9e6f3eef820aea4bfb263e46842028f545283fd3faa2
zdca034618461e20abcdb1ad8ae31ed112b4365e182b625714fe58dca3bfcfe958f2b21687222d6
z2903464033edb1dc168b95ad58d3bcf49465bd9ddc27fb6b53b8def3986d38de85aaee001ccd8e
zf030d6b18bafc30f36393c97a50709cab511efbe84ee87b71b4a0e409dab3213992532686fcdc5
z7e922e01e181eef87e7b46417c95fa8376bd1823b4f64a3396b836132f06da381d5c0217b3996b
z89d4342193428e87d8b723e04e4c9d762e77bf250019724a6631aa947d24ad2db9bb869d90d319
ze688f276a8414c32c9802c61d263dffb1bbb02e04e2c16f3bb41b3ec2ef4365cf609131f19fffd
zb11462299ef10347cdd18e15dcf2849d32ddc936df67fdaa0a9c2a4e6c31e37fdfbbfb6068ec8b
z69ed77b9f8736606570dd13944ad2d6844fe0418bdaa1be931dec8f16d9f347def0269e9473f58
z7c79c7779168fe8cafc6290666186f9201bbbfc3d628431f5035d70f93b9ba337eb18c8b6555d8
z385819372fabfee5fa71169777bd608aaf39c770d2ea9f0839c2afcbdd84742bbcb93d5dcf15c9
z759cc1dfbe8b98e27522ecfe53073869e4a9fa18f09ff271386ee01061e694e6c07528bbc49b8b
z21cdc317c0bd1363e3fc8e40cbd32ebb72b0ba3868bb197b455e491da0b81d8f5c41debb33951e
z4fa384f55860a98dd373b9b37460b95d89f898fe289b23b41ad6fa0e65ad7bb291e65d1ef716c9
zdedfeb094448cc32f1f2805cfa923dad1681183b5bd6515cd09ff10de29b1dd21a5b00a51f6e64
z6b534397bc79e0bf2dab492c535f0668d9a8b133117e06f2e17b8d7837806673120005866e87f0
z9e448f5b27775ad8d48bfa80004391d852b38acf511743cd8d2edf772bfd44d0acc7616cfea14c
zc438b75abd2c83b24ba0bb81c286ed378e10a23946e8f06b63a2d24c5303d317de3970d25f6aac
z375f936c6b2ca48c9fabe510dc8c79ce425cd7709700304ceae187677846ff553b6ff9ddf0a72b
zedf75e12c9f0e1ea7edc985a7f3194bad0aa8d485dd8bb6719fb7bd1dc6a34d1ef00edd23812e9
z8176cf48f2447b7386224c8430eea9c9151cc37fdd0c5ab4b3ee71b2bdac10d115db4acab956fd
ze79015a8ad5d6a0a63a713c4259b37419b970f3111b2dfe373ef4ef89f0e9b567fdc4bddd03bc9
z6b53b4e305a60c11d32213c49be59ce22094e354f34d5b987e2350df181075fb0d6e4e2a32cffd
z987cde7fbb287addd5db2f3807cf7bd79970dc0409abf89fb05ebfaa5ff7c4f55c4cf220f3db39
z1068524c2c2183188a7131a4072cb816a2c7e388a3cde0d6a0a856c04172bb108d563b2da36d3c
zbc35813f9b0e6918e23fa437801e58050f1d438799f34ccf4405fb4fac06a32f3131e4d3bddaa1
zffaf6f0294e3d29e35b88ab9117d95f56e3f2d243c5cf65ccff006f9e2d099eb34c9f7e7d19071
z7d6a3bc9613f40c8c7956ed94fbd5e70ada6599f2b73db7d62f2c6e090bfbda722ac41d3f00b16
z6286b57e994f8a59c7b14e10b49c91efbea71f0bbe81e5361c915f5688d84e39c057293f9bd98e
z9cae9b80d245a1a60b9e883a02ccea2123671ea369a3d8e31226938766a185f53390852c94f1e1
z78a85a28b9ffd322175f4daaa1d747222f47c465df9461d0167954d36b4bdd74526a18bc3f2a3f
zb09ae06c2180d024ef4a500f51108a03f222b64b8dfd2db18733b9afbf63a6cbc57dedb26abbef
zbe5d89192fa50098b317029b5beef19f5a0f595871dbe359a2d4fe00100a2c9c9d846c8a401d3f
zb7bdaf384ae022628f9571163a00d26b2602e1c78303e7781feb6d50acb4ef2900b7cbe68e3cf7
z9ad2052ac17a0cdce607240731c651ff8fbbfb51114b2aaf8f7cb333faa6c615cbed627cc9c2b2
zc796f52ebcfcff009112334d5ab8210bb67c8c8cbc8045ead54cd9a00eaf941a9046fbfedef2fc
z911e107929c69cc2fe51dfa84bfaaa7bc142a3123d69bde14e1d86b9ed666a843301cf105e85c7
zca64bbb32b64f91bb7389a0c30d133223686f08a4ee56573e5d32a06334b2f9d3bdd99490dec57
z0abbcb757babc3c7e1e3a45a62f122dfd5d52f100948221aa6e611f11c5c212f16f8801c68ed90
z565dd3b7fd7603fcf2456a5c2111c63976ae9e164557f3afd1353680baa72ffe6e3eb7c32ed186
z212c74672be5c5ff56ac1b5d8ca246de319cd079fb9f33f588c385fd92fc036ec9532423960c76
z07647ed1a612f60dbea5bc7527a9f8d9c5b92f7d83de304f8b761002a09a755a1dd8987cb665b0
zd1cc9bc40398b3ea7d77971825b07592d1dca76f98a57ee7c1ad5abc3f1fef97c27c70b626800a
z3a6024c6e26d0d164137456ae77d8bbc890e239aa7618fe75d503b5274a53b938dda8e5949acc6
z9578f2b76c2f97f11fd2e5eb36e48f0cd102e40bc616eeecd640887076f4e2fed2718815de5db0
zff7cebfe8a28e26a2131c771d87758487ba606924f3132cfd19d055cd92c4db29e4efbdbdea230
z0a89d65f8999bc13b32a18c3cd0df0442c27e49622f3cb9410ac3122d9cc32b9a22b010106c6b7
z506918aaa1d93a67c0f02c635454afa86f65a9f94619fa2897f389b6a2d7f4e2933e49eeda9e6f
z96f37c6c7d72b604fe8f0f3b687fe41e478852222da01dc58aa5567fb715ad38b4a9c6869aea03
za6dd022a975907ad87d574130c29400108b93f0471afa3b5c20ef236028c81f91514e3a6195057
z7bf473ed0dfc7ba29298486b4e690670367d58d463b944dd8cff8fd066d28125eacacf7893b01e
zab75c8914989649ee54279cb67d7c7e5490f1de94a253cdf7968836e3c10185cce173b030e5076
zcac4e3795298f46ae25f7cd82314208deccea7bd8a0caff41dabddda427453ae1f9f58bc7afebe
z10a1f2eaa3b47dfbe2e8d3167340c085057b2c22629bf8a3da0b6c59f8e3202041a119842dff9d
zcd2f1e95ebc0f5ab54f3a70fc77c90142c6fbf5696c032f831b638918ed22738bb4a53425cb7a9
zb6e0e6c653ae79a5bcb0b6b45d49488d155fbc29191ea1e966fd82811b8f3d10830d000bc39225
zb119bda1bed14b26aebf0e05a3a5db9db2960c3273ace1f533a55978ba1fea1b76dcb214c0a86d
z71825b533fafb17927972cbc05353f8a5d8f172edcda3d680251d9282c2a67a21c8a09d317f28e
z45a1c3f78fb0aa35d7ddc82ee93a72a243bc7b4d6ac02570946b51afbe159514db88160c84d150
ze935175134d8e1c2dc02253614edec084b7a1f45c26ca78f0a75d6eadd47e1e305552d5dfb587a
z470d4381fed0131422c4a0f99512693aad5f07a3325262315de2cb76276a9f1ecd39fa33dc0b6b
z7d0a902d5235c6db371318b96601efc7a350040f00c2b495592ab252c4f6c8a7cf6914cb3acda6
z0523b25a49c5837d818b213c9c94ada42db0b288e42fab419ad741b63843d58a1cecf5c688d094
zf3494f0f8797c7ce39f571bbc95b56c8e4610296a8c326532f7ac0b2d5562b95b9cc0164894506
zd15e0912a7da0e448957312ad457c4a4b69f0d4a37f7ecd073e36c465b57460d0d4ef602e9e146
zf8c5358ddf0c7b927f9ff9214f2bec7bad49bab7e0293c7c4bb47aaf5291c4a6cf60fd8d551b45
zcbf15273e5fa7321caacfeb2e1ffa4103cdee44a31d303421eb1ce8ef3272f328fb4eeaa448f03
zc64456ad4a57b991716c1baa7ca11fc4211c0eee41409d32b35be10f420bfff85c266c8bff4726
z62e69bc375ad5dd359fbe92b7f03050e2ad919567836b83d7799d00be449df47ca58ce6cf80e08
zf6b647c1eea670377eebdaec4f56e09be687fa331b645a1255144c2cfb5fdb49af5a8be97c7ab4
z10a30729c5e9f5269c3ba536562d2b0f9be01ee304a8bcdbf971c92056ffcbfd3f9a535a6d05a5
zc0bae0d0ccfae74af9323f68c63e0dded660907a959dfa66ac5b376f2527c072f945ebe595164c
zf8e03bf2d442366d45040acf2dfdd1086df7ee19fd1e40023a7dca024d429e4135f79e972c4a12
zea1892953f3d2831348d24fd1ec2bcd43e8924a32627105020f7fc6c2488f55d02a269896d0b30
z4ff29a00b496391018b77d830ac1e3b2865d8c030ac893988eac03c8e87237f637beaaf746d140
zcc8b17c2e510adab90c8680c38bbd3a3ab046bf97ae5ec9c5a9c6291edcd790b898c6f99f93337
z478c08b2214184e22cc5644df1328075d97fd27f146a9aa824c2537b6bfbfa369cf38a3aa264ce
z9b6c0b3b8662a3ff9bee09a1ef5a589f13d2046d48a37990284a83880e9a520770090ba56fddda
z39f7c9dad7acc05004e192cec5fd1381c90c91ca8651d432d5ec25be2cb7338a0529484acb7d37
z679d2c9af27d2717c513974ceb4cdfaa714590120f3a9b18ba469f3a9649123a13596d05cf42f6
zdb87ac1a782fb76be5d75b0ff8dd041d359449117c07343b2f55553075cfcea5ddf655702e3ef4
zf744456deee20365854115743662bf0ee2aae78bbe1005911a50b047f1e47ec0366d6232a7cecb
zc8be3936d5236b14fd457c92d753c0dbeeb03e7b80803021f3c6d672cdbdb2b7a78b015a2c7025
zc53b6e912b5b6f2a8400df5574dcede6b3f0585d1b702dd51b1709df85dc2cf77a1faf4fb1fc00
z4d9dbd0198802b00f9e919d8027969c47a74e9030d5117d38d311b360471095ffa31f7c4b81bf7
zb8d17bd6d9bc9532ed7a329ee139a6366ad97fb20c2b826e69c1e072c04c58459889d8d2e9f8a3
z7fdd4c6c15bb79564f5af5c961d2da65f03de6c2db3b75cef14557bd160ece316a8c391547a347
z4a720a131a99c4f5a1e1bfb9b54adabfa82c8a525bd76005272ec74424d26ef2de1994945bea8d
zf8f38a2528367bcdb7c1216f4c562cda7d6edabeefb08a89f347b5eb6afa2189306f200a9180bf
zfecbc2b7b1819b8ce5a1ee7f0531bcd70f597585186552f5f9e5c7ac10e1e300d1b1e951af6278
z7f30048b68fec137b442db6fcdc0fa19333814895fddb59daf7fbeaddbbb583d9db3a2dc93c2fe
zbbff56a7521152d053aa6991a33d21837f962e1c772b62c9ff2a29b00fb7e47829e96222d0f02e
z18dca47bcb895df452a42356ac2ce1dc6ef8377c96296bd06e987aa657fc09f2092a66751f09db
zc13e0a9638d18cdfb9df43ef634b1d1789ddd5c5937d51b3221d520827118ffb797f695adf81e0
z6d37982618698698572774078cf62de354957076ff5a71fd175e3c2cdd0ef50ef66ead08968b53
zb79eac8bee31a9143e4674819c5a5a73fcbf05de206b7f33b4d10b0557a66d0933eda1d0ae2b1f
z2f6661fdef255cdb102ea903c50ceb79d8fa028b7ac3998af8c91762d9b5ec7663224ebcc71f98
z583102bfbf72b365f18edbd5ff579af18681c44c9a6bff204fea07b46d63ab3d27d63a0654dbbf
z265ef04ab5465547059c169b4a4aaaac034b1b36bb9778a9aca2b1a6e0a31ed605ddb7f832cb4a
z4b3e23094f420d3075d6e4d8d5fcb8cded159afe95abd2e34a745c2ef177f97b900abc8dabcea7
z7172211c483915641f99df07d0dae6c6dd62a5d052ed21ae04797f8d192e503a76cb48c10dba5b
zf66dd133b3897155e7930a4b61595a08dd67cf9e57fdaf173651e526137de925c480d5ded4b855
zbd1282fb0d61bb8d021dae0f13e9d18286632a86af39f8e1b9d5068300be600755de8d0dc3f9ea
z2512c0d9ed070e0d34e995c51b154d94defff24c674e4711dd6b0e7a4152cd373d698b6ebca235
z81a17033dbb5f608bcefe9ba3deb640b4e548cd509c0c1b50456df75ad9568970a18e239c998d9
z924785c0d7a686e1e7dabfd9b947130a4e7206d7b02c9e034193385b52d0375994e619850a0b03
za5504f4f4c1cc7239188fb04d0fe422d689b6d8ca85c7179cb26e8f7dac7eef4f9791d1c2cf24a
ze148d18a69f9d5432d1eaf20ce154a6984498e315f37ff6c1f1caf6fd1aee7ddc263a4ce9a9f95
z27c29c4a94f7a5110890674f84745f951225bc053d243f8c5a63bfb3c1350ead9c98f3d6cfae67
z5e9919998270165a69a197f176bab999e36f63aa090dc6e4d5263f8e86b4f92d0337e98bbdc1a7
zb47979b96ed520bf87dde38e1e08e4bf2518e010f934b2597a1280a40bf0e24c48abeac3a8ad0f
z6844cad41ad45d0a473be1a9073e8a53bfca4971b4cb0855c0357c56e85d5cae2d43e6741c606d
z53a8ae20bb415c625d931e7a6fe12429b60701b7e9811b887fa30102535267c16ad0bb325bee57
z164bb3b5a9b0ed25623333f7e8277660b73ff9c826f392ffeba8e1335973b34b02118e5e1e37db
zacccaab60d01cecf820d381ebda72e4e888076e949373d1d67b20c3c431ba840bddff27498dde0
ze6220480d4f4e9480e79d83b62d75f748c54f4583684d4919f6f8569f0014141c6917e65cc1632
z315cea54801eb15c52147424174120cdcc6f17c31ac081b8d6644013bae5afadcb5338b3e6c4c0
ze6a4b676a3cb1b0a17a8909bf8ecf40f8ac27f6b357d780437d9976484f9445aa53158891fb3d6
z95cf4b01d25f5ebc989c00b28a17197b187c839f770ac3818d950712117ac676d46de4cc4cdbd4
z0f85e17c84e67105cdec90c40cbd60c3e8c907c0a53751936ff35d9a731ca737fad0af0942e54e
z9d23a69d11884f267266c9d8303b904285ed6562c0fa9cbd8089fec138fc0df72598ccff6c9fb5
z2cf21abf38f32fd116074e00dd154764d0361fe17e6dcc860eb431086bf0f0156e3a17e555e808
z4f50e64512f74a9f7e4f484bce3cd6fa34a4cb2ae1f52c4c8881a0e7f02bf6cae30a3917fa01ef
zd1f07827901c31e3d88303ccc57f8ef24662113da76ca897ce3b190433e2704961b1168ac3037e
zed89623b8e83c51ff8b85cc8b9fba84698cffed2df975a45f83f04ed86318b957d231ebf64f65f
z67727cea591f83cddd0b97e600e3a5d6643cdb56510075a9321513def41a8c91c35a89a5b54680
zbfed3c15ca8c815be4fa544a5e75983792f3fc59484ba0da635dea6e869458b9828e12829bd82d
z676c19a5bd1a8e94789060b4b2bb044d329e242e7e9c52def77474f0b99f6be9acc610a10ce5e2
z2a6ec0cadab39766370a992b12dc8cfae6468693ac536883cfa85aad8c383a3812cad7ddefb84d
zb458a176693ec45367d3765168f3c2678a4abc78127e5c46abe489a8757c89bbaa408c367db737
z7798b58eb92d7b0843990496aec96719e993fc613a48cd372dc5d5688bbff5228d1849da44d0fa
z17643567fff8f2ddfbb897ed9e95398819da9b8226e5f7bfd0025724d2df2b1a02665033d77a6b
z650161b4a21b7539df93ad4cc7ef8906e1f88215cf9f9418dea9b84b08b9a3eed37776da06212e
ze51495a16a4c654df17cd5fba6db30a62a506dd1203b81ee023a1fe830ba637f38cc469e9a6ddb
za06c299d0d3433ae47f29da113e9bcc15624b39b0017de88dee1e9a96938d9617576e6b2eb5d63
za5749dc9167ee0f54bd6b9aaa2a070f8d395db3a961fa8e0ff72683be975bc139e0837fac10919
z28722bf3fb0679cc895793f5352d071728f106bc8c08573abd821c77a7341ef5b8affbe2e15f16
z9fc5d9c5b5df8e1a349cec249a2fe9a6a6032e5fac7122405b6b1affbef56e799c84a752e95458
z67800b15ad4f2a497a2c72590b4783efd5cbaf19ab1984817bf1cacb0ca15da177ff411a69595f
z35109d02ca77e43476ccf8419a0db5cb5038b180a89dcce5626c814cc691cffb33661f843b5521
z984b05ed759d366f33bc6db63ec844a25d61c9abc5bb61bb1e9535f4006ce722a06399fd0bc3c7
zde814eee5df412e37a6d4930d13461b2c4d355fbd1432c8e83c064a8c41bf7df771d3afdf3aa79
z1e00ce4e4544349531b708e188f76fd32477ceee4e355c0fe5dab837c9192286471302df9737e7
z5ecf5f5fa4ad2fe0537aafe822acd8c377db846a3eeb7468c40f447480dee322e2de236f65d411
z97b8a633b3129e065066a41840716f1d81c91a4a11c6333cbafc63cd3f8eec859d64d603233c68
z553396a5badf4e9295948b277a4eebed6f2f11e29f6958c3f4b6d5c0c02d744dfd6c3a30f57ef0
z218561fbfb1db8bbbda125f98a0006fe56ffa7493078fc109c6dc404dac1be9f50a8c8c048a1fb
zfdef1f00122c085eeb81339b92e21c1fd55a51b6c8884f8ae3b977f40f0f426acc3a7fba57bc92
z36feb4ccd6477f5e781d77912550d8d634ee3335308909a7c78799473b90c6e7af76c67f46949c
z935cb68fca25ca3ee5c2642c9e71c80f7e4fa0d8046ceaefadcbb28d2efaad21c07d232a79ffea
z0368cab47c9212664dca4d51bf7f21348e1d52689ac07a84d02ad954714c5c059568dd51089bdf
z63cfbb2886eb8359fc61da4daad92e5fa60354a56c7093518290ef31fb9e3e878b78bcac1a651b
z99727e173d1ff7e291adfd0a39a152ead66335c08cdff0e1d1eab0781e4df4771ed3a2e7564037
z0655fc89f61606d9c3eb4a542dd14b28c2320ee11517767058977e2b764ab74b41e5a442fc04bb
za65ce55f797bfa93e4262c29e39fcfe9dac9a4ef6e0b6f7748b773f4386d57ef82ffa00e22b997
za2be2e3590395b59f4aa13e798a6f07c1fa81b7a774def9d4ff6026b7290376652b598b84f201f
z32b389de7a6a0ab0e982ba94eca71dec84523de9a21f2042d5bed638a5d616bc1a5ebd2db0d58e
z5d198a0df9c14274271b3849aedff5cd6e72849eed59685720d31648bba4641ce6637738489a2c
z10fcbcfedbf384b75bbf1de42c20f5f4869594a36c7258c4cae1006fba586a7bf6f26f2faf8581
z8294acd3d4bf4036b2f67b2becc0fc7d08c6c0f389cdeb9ac056d8f3f0413922fb9e602cb722e5
z17c4447bc5196d6c653e709095cf2c15c2c7fb7582ddcadda3b70ad070f24d00f5bdf5a2df5a7f
zd9a7d37f01a3b693b6376dc365dfb790777a526b3832437bb1e1ae97e3187c074151752e407d23
z30f202b791591c0e61ecb3f0f5b73cdf3109bee43b78c94aa3590338adfdfc2490e2763c9b1341
zfc649f80fc4c6534b4cda43ca212e6d3cb2c912fd061eecb61194bf0a2cff34e4c8819dd613543
z1040d27f1185592b7abc5b699d4e34af51f40ecb3e1656f67a67c4f96acadf245faab0071b91d0
z7e126209d7c98dde44867411abf2a44db4a2846b349a27ce463e46ddb6e0144cc5d9b8dc83956b
zdaeb081988f0aa808646a3909e78243eb5a0bf0d0385fde4c6757e3540d4877a8b340e6cda58b1
z9482ad9ebbca077661816ff849095cc8b6dfee67fd0a0afb7ebb7038168f14222c2acdad573790
z5808b7426d17d81e6c43f7d4afdc69147f21755f245f4f497a0c12a2d8e5c05c7ab2a4dc740028
z98806776d50990a098880f2016df2def89348bd7646b3693b554dd3c3651cb52f578f3adcae636
z291930bd19f82466c26488c07736f8eeaed7f8a8163a51de8d4a1253022f318d85ff8c86419ecb
ze80dd371341ebee2803aeaa023dcf64ca0da4b056722f0a36ce0bf20edfc3921f90d0e865d3cff
z7e3a6b3b9d402bf6c78a05b83afbddb6963bb977f2ba5c30deb67c1e8af8cb88a187c65326c788
z7d1f84e66da579eff25e41c203feb45a2dc553cb69f330766262282674c663c2fe7dda3c3c5977
z4e601731998cf8e62ef8cbc8aafc9b6b2d437dc2dee12151b354cb47074eb3248062ea69e432fd
z414c2bc5cd296e72fd086fd34f9d08216cbfbf76099ed3fdbe6210b41bde89a3e25dbae477b4b4
ze71666d39b389b058339d69a89a15ae75f6c316a0c18aa62dd6876b8cd13b3bc1ad0a1d627b5e0
z78441d200a7ec587809968e50efe683a08200d50edccd19bc09e36afc6e8895599b9a76864c412
z215d23c11429b183eb81ddf7014135711fba22382d93885a0def84d6c9558c48a0e7679267c043
zf2e87e1a1819e5d9564d4eeba9c68c7564f4a77506b99b1991ac67709146244c1489e772beaebe
z378ec6b216a3365983dba9260b6621e6cc15162be4e5c96b5960f8b732c5b7e543dbb56d079462
zbb787515447d1f2f5bfab00c3651725d87ae5b710ab22bc5455c2e783c9fb3c67b6d1d0515fb60
ze88c5c9ad530fde5533f323c99fda63b0992856f29d8bdefab168152e0a271194629e9b8262140
z12d7df6b62485f305045704a97c58d36faa52bac4213baf6158b1aec88c885048c6ae98a7b6aaa
zb6eb9e9b5897b18c3bd2d43136a33e3a6c4436abad478ffb5e0e553c63888cb389460033d65d91
z1dafd425c2fa1b96d0a5952d279c2edb2039718f522e356082e7cc40e2b03ffc9299b1c1ee85fa
zfe77bddfc28635cf092ecbcc5675c4b517beba38c9be999e5000c3d846c2099b5216a4e99837f4
z3e17230e1bfd3c2575919dd0c1d568321364fb19c4ccbad6b7b689d82c336e9cbac6fa6d120b9e
zdb34b3b315fcbd2be68c86dae83b8968603c6a740e3815bc00c37c1447db21097b6512f840029e
zc088b5f6a051dbc88ea782c5a6321e32a119ee3e9b81d3a3de767c333e870efc6fda19eae85df8
z57484f4da59d45a0f81f6704ef52bbe1fa0d0b221fde17fcdcc54497579072a919819d38afbdbc
z92660bf4d767bd45ed3c35f80c43e0e52dbb9e6c27361dc98638759e8607f625458c0fb112c3be
z5e8299248e5ceccb792f7a20f09cdc89490e2e1184ca8f9a2700cf1fcda9e98728199994fb43b2
z58dd2b447efceab8462bf60a8709e9b23bdd155bd3f91732eaa108911e177a88d4d80dbeda785d
z02175077729aad90a48acc6f8790e679b363506a65c3dcb20502a6c5445d5d344e08a4235bc78d
z49217720055e79ad71e5839a9ae02f5ebe0ff57050cf677d1aa694b6ae887683add14d473caaf3
z0292783766d1e2c36c9e306f9410bac1af80bd9ae4de4a32299c4ce74c11b9a9a746046fb555bd
z555f5349a53fecd84578ec3dd229fcb618bd49a889aff12fbffd5086729cd160ddc2e404f9876b
za8e7ff5232bf1565a5005ff64bb92e883e22f209fd7cf49832dd9b77376b5b5552ec09cc392ae7
z206f6ee07bbf2fbe1cb28eac2975bd90593c45d0ad33e60f649b442592d568eaecb3073a8ec1f5
zd21920976e6479f7715f229baf59c5ae579dad80bf3ce06ca09f57267e4b87d1733b7389935720
z5514539f11c5c7e220544c64aa065d73f5359ff955298883b7866375d7aacce1e5258a035a6861
z6e1cc61cdd1957781272106d048ed18224a03d76eb57b39b3d425083c55d166ac916d7ef5c3821
z8d878bced35b64e8ac4d765fdca945e2e39ea678516a44cc44728875399cda388a86af89379d73
z63f105a6a2832dc7589115cafaf931a8f1b96b1436d044d78e0adebef2920c9c0295a165d8aab7
z1b21a31d7e090cb448ab8a8858d9e61c5cbd5ee74fab55e5bd9dd066daea738595cbcb32b90ad4
za3ed39ba2dddf2a26542c11e51b507ef557ffcd1708d6b44ead3a38fbac62b4642bade3ee259c9
z08574e3a425043ff158335f559b20912ec3f9059d096106d82b2c5bac12dd9bb83ee47fc5f20ca
z87f06b698eeb3193d11745fc953f3d74f5993c8a2cba680036cc630420b7776e991c692a6e4323
z00e8982abadddc77cd2f829f4519641fd6de5dcb9e5cc8aca8b73aa1431a567b89e876ead4d7d1
z31d315f077b41e1833f8f7fc696c61703a3fb234840cfbf48f9838c78ff062272a7657c70c2e5e
z4f4863c9e783c4cab3b8c29a2f7da0ad95a30044679a80a854485773755a429beec468410e4572
z94f867cbd1bca72865e5de42c4844d9f8bc1591e96832fdedad42e6399f0478aa24d479367b61e
z39ac2f4aeb200c866cfa5201c1ac134eeb1e9ec32bd2a4a907eb59b69867f7dc61c9fbe2fe8de3
z1d2df4df7e8f53617ffb0505e112e0f3eaa3a8860f94aaf97244fba591015c2761f9ed1374cab8
z5ff60d61396c4110d0693de614d93efee0a0006e5fe5c439a575a7d75d828b06fca6f7d67529ad
z85029b13dbb84a3840c9912c37ac48052f86b963d910ddfeeed7fa10818447f59894e2017ebb2a
z35cf7172e7ec9ecdd88183bf7400ca2ed49bea8f9d95613230323fecfbd612e6bf89f5aef6598a
z3d68d64dac0fe31b9be714a2d3211eebf7cbd5f58f4b9ba7000b3b94f1a8d11090f15214789e27
zfe078483ff4aeb26c3e0769d1af9b9afd70b83c8b1db37913abe88af76443773a4b1d07dd05f0a
z3c46f6ed867a816e27f0bdfbb72c6d1687e3c7e7d3d1077d7c7158eca93cfed455b3e7327bcc76
z0d84fbf3bc0701245faf07a641426362752ebe093f111b1c275696760c23de52493c754cc509cd
z39e51008e90c22d4dff89a5bb758dfa641ca00e6ba34f0f1d4cb3e57fba16d408066f9797fc5fb
ze098b950f78d8084950a6465032b8ad9b98e05fa44b0ccf68e4a8db6b31ec60335ba5d31425af8
z537ef2c66c6db47f12d4eccdf1495971a7025f264f3fd7425126bb93de41396ee6a8410379dfe1
zdf0f15f7623e6fadbe290c8f88c914358b3479c7c98c52f858cd7919b7127eb85695d7698dca61
z306b4eef8ca518a0de0b588adf2df66c3946e6cdfb8582651248266fa8694f6fb738cda3ed5840
zf53a48ef132c279a23fe122c78b0214257348903f485c0c136f4bd1501f241baf264f3c47b431e
zc801408b1532a14075d9e01b850af24ae3766335fd958c55a1edd8e9a4ec98fa23bbc4a22f02f5
ze94be334e8efefc1907bb7d100a6382025eb053e083fa4854fdaeaeb3e0032e516f424ee1f3ba3
z1e6130b7acdc162f08103d0406e6245077038b566b44647cf9ec547712621713bbf219828061d6
za1c9c42b6ce4f6a1c6e0d30f65d358114354fdcc42bfb4f952a8afc9bc16cd4bc21368f8cf8158
z20521bd6a382b914da4690c7ceda44a0a7141740e80bb4a45831357f51a4216e0b013f80754bf2
z58b6eeb1629b676b7c4f4214e67f487d15eff8eb01a788bb5adda5eb7ab0e984bdf64d4d40419b
z6a4d099672c788987f5c4b96a93023fec73275e9beb94936ff9353236b0f17306501b42d4089f8
z2f978b133aebc58d0ab5afcd53eade71570473c3da06692163f42589b06dc2d11a5f51cfc20027
z2f1b226e45cba4bf1dd5d52be201157acffb8e4a09e53128d4ccb7eb1bb5415016366052097ccf
zd1fd02aa5ae247230d61aaa695a26439fc35ab90a5bac260b4026604f6538ca4633721802802a1
z985c4365a20cb173505de8199e88766b7fffa63a53e19d78c0fac6f20fcb453b69213932290d8e
zcac0a707c855a27c6f0f21f48d366bd956502d90bad2aed94f50a8f6d210ddcf60ab47356351b2
z13f6889ea73839af46adc37b2cd0282da4a113cda2646f80e98740667e38d90a683c8338458276
ze6d16f494cbc84deb093ce58a3b9278d2550d4498e3103ed2693278cf6c835e1732f1648d2e1ca
z92e0022b9f06f57221c39759731a20cca679458dfcc7ee05e207c9e277d51af212c48d92c79336
z6b280462480b3a323e2ba52e5cd984f60ff6c5b1ec093ea5ef6156cd7141dca8f573667bf81446
z5fe29e93907967240171a16a682c76afd6f401e20bbce648e2d9ca302a0529c62c2c122e7c9cb7
z39a042a132ad460dd655ac5a80fcee1c26097e2fe9a9cb000aea934eab88cf37dcdd7321f38756
z69287620687c2092162b29109967770ab238a08b47ae261d1d68ea9d5f506f9c679c268459e028
z51081dce26206fb4f7ae26e14d608262f16d819a3a14280369c53369ee2853371c626844061fa2
z2583db835889c3086bad17baa20cf6ae4d1fc5aae8c20b62809df1abc931d2d29db11cfbf0c241
zc8dba5702600cbef9cbaff919a2b855d2e5348df4f46a378cb1a7fc8172da72ed36f787f51d996
z8f67a0102fb20bea3c54f37e9e328ee3f1d7c79845ab2e1281581fda71c6ab16e31995df37ab0a
z4b7d7c594118ccd1a6e569a595056b99fb9ac698fb37175486fd04c08ab0bab66d3602b3bbf464
zd0011406aca8904fbb407b0389bead02ab6d54e9ad44c11469ec5d33663bb3bfe5310e5006b838
z0d5bcf0efd70b1955fcad057162ea3b2d20c636dea5ef54fa2ff5cd77218d49a9656f84d9ee436
zb7ae51702aa428d84eb57a6ce9fedd3133b8373583f587172a8b2e6af077fe8f66390cd54291ec
z5fb48f3cc88595495e7e09a70643d6ff44e2634713c0f0f8df5d9ee92e6d0ae5237537603db022
ze5d2a4c6d33ffcf1943b322ecb96c21fb95464766ecaae4fdf3a84c6e97fefe3b95fffeb2cdeff
za4e7c3c84a2921884d4d02e4bc71238e9e9ff01de142b17d22470779470930f05d218ae14eccee
z231dcc6bd84d6e1f54dc3553bca7cbe0ef34c56b04921ae81f5e934a95e6750ff06c321e165525
z8e4444fee5eb57232ebecac1ce43bc8e184180216ba0bb55f0582bc0f64e711b042f495a087b88
zea376695f6dd81bf255c57ada1156fad4e2cb4bda1749ac040396f9f64c47c47c4d38d6fcc0205
z0c4afecc5dfa0701ee1750dd5d05723a533d02f0410d9706483a3e3ef748102e4a9ced3fa89498
z6e93c86e82b83a1f3d773135676e1cbabea06b0dde96d449863876d256ffc1f3cc9b474e68a565
z684a1782f1c5f3a25e53163e6d9bec51b3f82e893d98a74693657414e37f4e9c838edcb017a6bc
z7923ba6af7b1bd2b0f82880c5792e1471fbedffa4e5414a26123b2e4f9b13ad62c84a1958e024c
z0da569164a1862179c87350784ea4c86ee20af0e0eca2507ecce44431119400abff894f72cb0c4
zdc795504a5e457750d6d13a79c741c6c40339e63c9dfb626c2501586d641a4050cd0543cdf063c
z557691c163332f81c893612727f352f7f5ade95acecc3a9682658dc89c01e5864c4ddeca101b6a
ze3942404aef5e0d3296e3a1e928c65bfb6237f4ee555c80ff1e757d75aaf5c03c3cd8db4dc1ddf
zaa7bb0ada947fabc262710453eeec6003c381b6b1b1695c3b3b6cbf33ef4559e38c89569658b8d
z0ce15bf01ea48c5a6e6f47943faef59891c83f0f4538981bbe61225420c5c1e5409936c6be581c
za8996cc4970c20acaf0a31b56e32dfd67d97ce4aa5c9852434deb3216df6465363aa4b6cb5babd
z442c7fcd81b0ebd50f9848f4ea02291f4360588921e14ede682573cf704b1f48c0cc97a394391b
z4f892a1b9e78f0e1bacbd1fd94ea41dd4709743d253757d8e6a8ac5c3c7900e3b29870113e4879
zea150fc44a39f683010375bbbc410512e0f1f47131ab5e452881e2918f596d0371edb4478ae4f3
zc7b52a9a0403c6e1efbbb56dfd7375c24933a5591c3e0195b88d787e8c7cc3726e100727ca01c7
z0ccd3ec5fb20ccdc3e4d9c80760a2c664fe1b2555bcb2fdf76c84e916f15041e918b304b208e7a
zdfbc58708bfc7ab705870fb8c1f84c424318dda506f6f7fd855fe5b131a86bd1faa5ce7fe2ee0b
z91b79e5c51625ee2fe0e67456c5c1e3a034d8c86a192cfa93d9b213396b6a87d4c45f4900e1f0f
ze8b4ffa05aed1f3fbb1166a491c12133bfc259e38d2fd655d5ff24582f60bd8bc26a02ac134b4e
zb40ae300c1f69f9b3bff17d05e94839752d3b5832db9f51b70e85bfafe2c88462553b1503c8f03
z6a876d0d2595316c54a318e68c127d2aee43ae1c33b481f99ad84d22eb3a312964f58356ed0f48
z66503477a6009f00e99cf8f0670199918c7d1ce26b8fb181f1f0d1c0f8a644132068bb4c033fd6
zdfe8b1427a83ef288d0b122a105a4df39dd2656ecb35e83c8f2251ed078aa93d55c0ed197501d3
zbd87641c7debf0b44fa9ea4da2e46715a91554a087fa45a2106fbdf0c33e3156e4e6895fad09d3
z79cb0ca3e52bf866e2ee9180d727abc8556011effd8c63f82b5bd86abb82bd688e5819ed6aeea4
z7cdda8d8a26f830c87a67752fd256e4fa24693a37cefb9f64649ae6ad4118814aceca7de9041e1
z16dc48c0bea372a68ad51c0095f3a5ef76b8d32a73f50320024d52e6f98b9e3d8d2b611c3887a6
z671aef09e701a173261a6bc69915cc5c63a393360eb8b9b6fbe846c11e04a31ad5503c6a980604
za5219780b47ff6e9f2e66da91294471b1a17eefb3cb8bf3a24be85652460dd557f4c5ef2ad80cd
z2e329eb5308e5f4aa4a12191ecc14ee14ca968288fa6a9f7a765a31f94d6f6ebde53c53c1dc34f
z01233343d26af4f3e7154352fec185dd42df3cdf262afb3d53bf45f4a7776c219bb0f694a26910
z18d3983e93628966bb7d739684832d059a7380ff6017a3f548323e94f63f5a6629e7c9f68c4a68
ze269e0d4c1f7c5b08ca2fd0333c91c661942e8c17ec8b5b790c8304701a4448a3914da7d388589
z36a351c86f049194f05f7cdc5a6b4da68c1b17062518f0afdaa9969cf051174b23fd343fd575ca
zb92137025b6195382fc492706b136db053e03f414e5a3aea7db11b8c4408e04b6b7a4cde8a4c00
z0daf85845362849a460e6e77aaa65c59c48f1e5326b4b6f42f69e0f2b76137b3cfffc3c6a80a08
z3e01226bc1d207f1cd1641ae14dfdc1a6745a2f9c5db2801bcbdbe3ee2c98756d8ec10e7f7a2c8
z74f2bf1ffed7507f98944c115aaed5c3e6d24912541ca4a70d03c9d318ec61714e8bb25ebf12ee
zd4dd58fb1ff107a4b997779b6a48305eae137e78f1a338186aad287f7dc06043d0c6728d76bd83
z6ea73e58d876cfcdfd0360f9a5f1511c09806af4025dc9cfed6f96e54662fe37ddc811a9218cc1
z1be5e25fac3f56a633d50d45d02b1f8233a1de8db3864914cdc48d47e53baa080861109dd0dc1e
z218886ff1d447b09b9bf601d1608aad4f10a862c2de2c607a4bb8c1625425258e95c9fe1150d22
z18d1177fa7abf4ce1456d6853087b13a34ede47b193a62a75947caa696019bc0063fd9d4f82c7c
ze8ba2c8cb3b2f09e1aa84988f5fa124242c0b7d621d1f3ec369dbd4e914d40ee5a36faf1351747
ze266942780b440d6ac6d9acf97728e004267dcb9906a2f4d0bb876a632c4aded1e9f5f8e251fd3
zc812e9703758a068dd9698d81441d724fcaf54c34178887d79627bd72111ab3267d14c5f0b219d
z8644f57152a10031e29b8c740add02bd608ae188f4479ba3965b09c712b40192534f6f3f2e3172
zf5930c817d82cd0e2407e14fd8dfd21ce236b260f63d1054e6c7627690afc1040cf8daeb5f0709
zed21f507cb037fa56a10085af7575ac08616e76f8b11e005be13e8cb793db72a0c2d06d6213a39
z325f451d1ffe0b7c7134408af121207d31d8e227e80f32f9ed941d408dcc091231eb79da6d88eb
zc8880a1713f2c98c55b34a27327d63d9841e3d746dcac9259987f5ef5570498f69b1198a17143f
zbc09a8ccbf4701f6ca5e86f2c4968ee0d2276603e299c435ff16a80a298cc618cace9c0e88f8a7
zc8f1ae7ee250f569a71723120a8efcdf0bb129d79f14c1fd26b45fb6c097c61bf6b28b66eb92f8
ze1e8b56758c55ca813edcf05314f43158e55f5bf8a9e28c3b6db17ac8b6ec656f2bf4982cf09e3
z298edca2960926610eb3004e661c6344fa3e0a12f92c811ec6b37b80451a0ba2b665fd1ab58b0f
z5a8f813350cbfbe61dc6d12f48dcb578f2495e1b1122c580c0bd95f222b998e9013f07deed35fa
z34c8aec8616f138a386b0e345ef4c089017d61e08dd8bdf4a8768a8aa344b1a64d728d1f49856f
zfc8009c677ade1353ac39b336af9ad2499bea054a8a5ab322a382fc429c6b81d9cf8b15b222e66
z76b461a56fae74797280c4284a1e9a6e81b656ea69802f5d2a8efc014576a6f0bb89ddc804e0d3
z1e1d3912ebb6bb8185addd28c551b3cf21609f3a118943c5273325817e145ca861fa9f58c6207f
z5a429dc5cde14bb24c9569b003fa4ad8f6a1531889da374ab46a4f64cc7176a938fe802e3905c7
z7b8133ceec8fe57a9cf3864ddb0c73f5f224a87d0671af56cb918fb481ff2ea94ed93d659027aa
z5d9934b3d56e3450d1b2f25d92d09735f54879eae4bac97136aab4802d5ee36e57e71ebab6f8ca
zca3bd930034699f3b91ef5f80ca6f035a7c7305ed166e51942ad8b7f408c52ae8ebee596057371
zcdc627a5226ffa5bf69d4459bc97f821db7a2c7117f31ac0aa26e0ea4f25b5792a75c3c91e188b
z131fd0574bf80517b5d971a3dae84ccf9254fda4be7810480ec3ae83af1c039d323ea6f3b03caf
z5586a75141019d26f0268f09b410f8fd2b70e956aa4e014fadf9eb6b76fd2cc5e8692dfdf4e50e
z59473063d9d88a543d88f787be2e2c46c3e1e41ddcd80f143da10af1fbcac03418d1864d511a78
z20980a329855756f3499e09f94697940730836377bd44005f7e58ec1e7ca3df08c2e112d7ca022
z89a459658505dc25d4a5dbf0e0fc904d6aa1fbb05c0134f0a28cc6631b34643b383cc3369777ed
z1827b60b2ae4304451db67e481db1eb828624e5edf2b5787d30d729f56bd47e13b8ca5af4bbb9b
z6e70999e1bd2368b698e2b5becf23916dd899c6e8dcff7dfa16001b373bd7348e385c4dc953a1f
zaa8a333c099624d65b7988ed67b00cfdeeaecec08b034057a30fc6ba837e98440810e52a761bcc
z934e32edd37eec249bbf2be5b2ce71d32dbbe77c9c0bef10a06ba3fad4f5f365d8cf137c3768d3
zc8d78ba05220df24a319bf00937e2166ef46b244f134a23db2a5ccd44f4aaa66b7fafd759c5b6d
z0aa87c3312912921c134ce0ea6677e546abbc41e151eab7a79c85f982e105b7e4376099daefca0
zede735a6f615d62355bf2027754dbd49debb67cb5d26b75c2a1afda3322858432f5384c8cc7ce7
zabeae9347fc52e9243bfa3933da66d2d106b5647b4158e1ca3c560e57ca320a89d57024205b22e
z221d811ce003a0af2d9afc05a73a45980ec86fdb9365fe817fbcf6aaad27e7b293ba95f6553bf9
z6d2cca4314e0f29dffbf1adf5ef9f770a5b21589ecd9c88defa09bd877ad35afe5a12ce05368d3
zf63729bcfa11245c6e61929f52ceaff5becb6ba0d5d47366e048d0aa013992b8e3dc41e38ff1c2
z677677c2cf2c7e297c6848577597a38be84fd31197d3fe2c1a3d952144d78c2bc887ac4f4ccf57
z0ed816049d6ca5bcdbe0e236c2228aab9f8e5b910d2abb64e714ccca18b21c6cc07a6dd80d732d
zca73f51fe624b3088f7c5be9bd6af68a0bfd93f7c8822894e4db239c4d2511fdb1e0df7631907f
zca5a33ae547e258ca13425347ad528cd7ba70ef2bf5ff42bc60849559c65d09dea1625e00ab056
z6f8955d34a5608f7e326d4972376e54a9caa60ccc6b9cdf437291d2bc5b8ecc19a95b5e2aa4f35
zb29f43406dc36462bfde88b59458e175930933a7e8c8234096dd98d7299bebcf3ddf850d46851c
z6c061d0ce437e237cf258ce5aa61d4061efa3160b20a07d70d8cbd052ee414fcdc2f9a53d8d29f
z375fa7bf3b8184faf9381184266c35b83f314c6095caac46a00e00319316d48d45058dafc8c0b0
z8c58183a2bf6ec20792046e2cc49c21ca8d8f2e8cb6c5096b6792fb7e91978e3583b0aa246a087
z42c06c7de8969e337b415964b4fc24b6cc96c2d39a18cddef19968f320fd95b0296c1016414dd4
za9c779f86a5ed450d0eae632df90e1e2ea40a92097d7bf9aed3c7881ddf0cc959a192a2f3dd082
z613f77a9173e1d6f7169177a993aa71aaaf5246bb4ff534be6fe71243fff5d3305e386d66b72bb
zfa9114e5d28e316d505cb90f2e20394542b166c6cd03e9f8bc3068326277816b5cafcbdf5a206c
z9b975c313aac6b41d0afd213fcd80223dd7e1d7edeb18fb7687f0977851f1e30b091bf394daf3a
za5edc97528198f7c26e631111d58028aea7c8f43b30798ea97e42a50d430ff5843c2a1eccc543d
z22df7ab65d30514f3068691bdd613f81044af35c1394b13e05da940767a0723bc38dbd44f596f9
zd9c0ffff8335e7407e0b7fbd19d3e3428f2d2b9a2bf4fc733ba4c1792a910f3f0ad96c3a71884f
z4df843f9ca72f1765cce3dc7ebfc8b87c05433a2e7fb02dea9f5cdc8cce401404de77a6c6fe997
zb2263372ab835cbf0c4d25dc7e6847cf6365fd33d01419e0fe6aac488c33f9d8c058d7e5d048dc
zfba782cc06817fbe74433d7014e4beda3c18499e501f61ddbf6cdedc7fa7de77cfd21a91a90524
z77a1cf2fc8d810fa548fb747116cc63101822fb6c1bf1611c99952f90d7192effd8b7d29b5e0a8
z8e9bd7e75a4c5ad221131fa62e4a219542342e8c9fe0414af4acd9f4aa4e0325526929ec9abaed
z7991f2b14bd8db16fdece7f7ce06e32a01b61b075c215de25995f70e22b098882994451d5a93c1
zdcdbcc93c471dd777c81ab3d5bf1baf79d9f41bd2af9171c41cfaca704f1241d72f7ce5c41a68c
z452825969cc8b3090f14749bd2ba2a675eb5eade75aa55c4b44150221f29a5152640c3df53ab37
zf2dc9ebb6a9679fb0e6305c2e0f3cf2d2e920a24209f45124f204ae0be3bcc6db7077be7c73262
z0949cef8b92212b8f2b281a0f5532349297d2cf2c33ba64c6abd6875a810a719d7ac0a9465f23d
z579bf88092d455cea0e19f4bac7d8222fab63ad3a72ba46be107f4f2cc3c8df16cddfa84134de5
z85c21c330f9ff2b5de54d125fe0355e54dde454f6f65ac156067eff868d379ec3b5af38c081fa0
z607a31e627fa41d5608da6eb11418d90651c2da1f72568b19d282212d7fe0e02dd8295a626523b
z4d4922a1443042d6325f05447364bf2ac66bf8af1e16f87a7486883613d6814b411d558d60a42d
z88733f5c97cddcf50e945a4afe36be05cf8da699efb2a30d428a0f8c917858d1d1b7fb5b267075
z0f04848663323d265a87ebc618c64ad6bcacea9ce8e969bf1d80c43498a5ac4133e732323537e0
z2f1eec440bc26e21aa1d906a7b59e8b8213cdfc8949dd9db11a5e356eb9e0d4193c034dad84eec
z7a480039aecb2c6c4dfa822ba6834d9b4433779430ceac02d54718ac20a62eea4d7e82babfa1ba
z7701d40d5ca50d81d47ec11fccbf0df52d8ef312789252a76881877c63910633e0d071f0cab63e
zfc6b171593292f380592f6b75b61b286d921db76e52747324b8d35ef3ea0ac687d2f7111377bd3
za77166bc8b7b7fd7478af17eb810cd4507cd98c78f00e6aa0fd17eae6228a614a4164b5e707cf8
z6011ef255185661517593e54e652db8667d37644c868cabe01b6587f89a4c933588168505754cd
zcbcbecb411fe2b5bfe0b11930a7cd8b5f92978b1c7053253585153475b60cabaf08c96776202b1
zce9314317113b8321081f3338c10410e59d95c154902c3f1f98cdc1638c348a6e5d7e34da4449b
z895d32f0c128fb3233b63bb359f7199af42a8475933d29720c89547a2dd583c76bbdb724cb70d3
z8730d0747e021e73ac2cf36b8c1fccd5a3cb3cfa53d2e73ac85674babf9c90bb34745a4c3b732e
z92c1f83ffe19c9b0bc9a7a3d060d9f49fc816765e61f825fe0459d4a8ff21eb0a44794f2a43038
z7f5b80340a247a896d8b9048d129088177fe4d15541ae3f2281c9be5543c0981ae4830d4f839ff
z86fcc06757ab1e0bbc3fc7f736b4c1f6ea971921320c7618433389ac0f4dcb0212d8619c993c53
z1165e43ca07ef6c57ad6a2a137db0f60673f321b0d0114594be0312e0e230e863d86ba3e028da8
z465d58f4eb83fa96e673424c79bf88d68049aab2b5e2ee09010e1adc5efeb8f30b86d007317e45
ze19ccce6492e6c215eae41ca46a23cb3c4662c43218779b025eb39cb2180e617c03eb9c2a08521
z29b2f605de8646e4c139ba0d3a24ffa8367e9defe1c7240bd5114b6ab953ec5289a6706163ebdb
z699f1b08f1fd3c219e436902e13471a9f6c439376e7b10651aafb5f7e34f27ac5a49bb944316d9
zbed1eee1e7829c430246a405da7f6a94422c546bccb587fc59f199579243dbb21f29184517d435
zf2657a52f2e8ae50f1b0725a8afdd17586083600a97d2385defbd21d3137c6d9e6a70e9f3d9e65
zde264df2ec29833ca5e1ef1936e38d8c7c88427b6799eeb6a593637d105ce99de4fc29bc714566
z0ad5a949617a7f26dfaecf1f15cba60b8cc16edd3c41cc3c050d83a6ccabedbb2b951501b23c4f
z896146255aba773042f79a4d179b1e5e357f52c416034a6ce44249d7505f1866442536d97b5e58
z09be0598607c10944f6f3112737a53b6f3707ce1babf3a1335a3c2762da21d74e69c2964a56f41
z2f79ebf1944823c17ffd30890f7c633f297fedfc2238582f96ec4a6626542f6d50375f1ce8c7c3
z2fd25366511c4a90ac09d2f6d5934c7969d0d43e68d6ae2020ca3406fea4db544b6cfc044cf309
zfa9f30d2d570fa335b70a02f0b1d274dcbde353b430e2eb0ad2152bbb318b01731dd64c423c50e
zed8447d93ac7951fdea75cc3c4aa62179682a3e413a03c42b838bebc56dcab0aa8a356964fdb26
za2eabf047d344726bc7b31cf0d62380572ce329d3d0d6ea9280bd4074f35b71e51bc1c7fdc22c6
zf073a7e9c315d61d03f8c174a91e4aa1660260d9308954be9e9b2b3d74ec50dfcd96b691693e58
z77911e70f6b4a6e594dfac5d1d62baaaa9b0bbc60a8a92dddb036b0ea91645ecab50d0b8507fa8
z4b254e32685830aa6645cf077821edad3540c0439cae269c4bb51c04d3f673422a76d63622bc8f
ze76337b6be2d3ca385147b6ac7f98717a1ae27fa62889e9239108d688412056a53f9e6224cfe3b
zc9cdfb84c5fd38def45c153813e8eca2eab76dcbe9ea93ab2abafd77d17911fa2463bd81f67559
z79c1703f9a98b2370b3d784a38b216e643b4c7a0cfa326e79626dd796b7bdda8672b54075f25af
z25d56b2631c1de9bdec59519ee0b12a8bed4dc7348c798e8e296aee0b97f80752cf9626683c54a
z46b952052f78fa2387647f78a11cc60d471c6cbe6c3d469299e7dc96fa80963e6127a0b7490fb5
z5008224cfa5c2a4f5d95961757647f28e995429b6655e7bbade6e5c1a94183ea5e23b54c68ecee
zc76ca2462e148f88577a8b58f94ff8e03463cceb7ae16a4416f7043d23b4efc9c0c47b70190f53
z7f546d6e101fe22b27f2087aedfaca49c13d8a3ad3e6c050bb13094641a7e63bf3185c00dda6d1
zbbb12cb466b98033a3109d931023812aca2d1560c570990ac732e6d8e4909dbbbba3f2d8ebefaa
zd83d2fefd3aa9f45564f2d61732ae6fb062d3de97db91cf9e73208cb18959d8f3654f726f929fc
zfd98c80c930e3538ebdf9d1e11bc30f79806d1f6129f5776053143102ad631711abf75c70ecbd8
zc1da7fe5c399fee67a72130e3d1660defb4c4e7d67e9c4f814ff6b84a23c56dd282159a6c1a571
zaf764d967bd0f56a4a38199fde10a28957e93e75217973746f971a4028d43e84e97ef93a5bc0f9
z53a813615a3cdc96babfa61c8bd01c33cd4d12289f941f6923c85df79e50e10e7a04fe20ae1ae9
z92364661cfe46fc4a2d6c349087ea24235f7325a404177b0dceb21f124d33c59be0f4dfa9d60e3
z877869158781d3766d5b7d57436cdbaf2079f09969df039965fe9911528b19938dd1df19ae8bdb
zb73bff836939e42885dfa7aa605b916a1525d5ef943401f84d8305729d745e2f60c71993d772a5
z1fbe5ea78e66ff90bf527c4e1134994cb33f62d9ef402d3f092ebccea91f8a3c0639bdffca7879
zbb2a04a1f1f426992fe0fb33f00a3181561343f8d327fd08931145bfcec639fccafdb022787c52
z26e56bf24fe0b3f43af02fffa4399d3eaec43a39df7c9647759b31da6885f97770bbc7420f1a11
z443ac45a76f29470964d4f2916cae8b3fb1e4f746d3470f2251f03ef10672cf00964c7cf410691
z7cbacd5d6e10bbe2ca645c761479aa0b396feef660a74b6ee7df638c4337d55b41fba180845cea
zf020a9a522a0833d6ff9351a48a3dff208a7f318fa4c0933296e27abd82faa2a42c8306e122b00
z7f4c47c56970f01d0226f8f9325887bbc68dc83ae317e246df9bc66a08cf940c93d07acb8c400c
ze31940b97f7ea94cae605351b1e5c37b2ad57a237a212fa461daa12f1946d7ab781869b074c1b4
zdaa7ed28a0c2883e2bae594e0153f2515f703203296c8f0150ab3e0664814096585602b7e8a6be
z7bd5d5f1db428fc3b2800941deebb05192cdf79157c55a74ea7a1f78eb6d3650dff56f52e419ae
z5f2d8dce4951004b0b17b70a9381810048b566dee9307f1ff8844bb39af2f1c4b77226d7a75268
zdb66f31a104333b16ab13e88eb3e957ad31de2f6935239b05f1ae6663f523722b5c7e7e74fbf3f
z39cc14783839dbfb73870163e4a0480853f3e1de8795fe25255ba01ea115d71001c16d51b47770
z153250af39b380c99a9999770c1a1bdd557b729f84da8ec8977f1dde75c758c825af5874cf79bb
z286a293d657dd4416c1ebccd1037d5d283b90fcdd1da258d90beaed2e1340167fe279caddc9ca4
z60bd6e93f739a0f7a1a6abe32abb7d668281146152c064383fe5da17e9ba1e1b03d4504982f3a6
zabfbea55f78b3ae9076f6916fc6784c9a34a5626e1bd4b192ea4e01a068a66704d728824091d2a
z3c4b409330bcdac54e08eb58ffd8084964b156b1e71f75ca62ac64df76adcaebb8134dedf2847c
z44f0d70266d151701f2e1d4077f5c7ac7d8ab0714f3ef6db6f7400ad37
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_parallel_to_serial_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
