`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab30857016fc53a
za25afc8341302f0c829d94450c399b8ff9b0386c187cb854ee330605b7b59da379b1f26f488e1d
z36e675f0b1336408b3a1ad87d0723054f952fbefc8d5a33eaca6ef5be8f42bc59870a29a5cc9dd
z4fec09ce6e44cac279651402e7e1f590df88ce49ec26ab39f12b4a02855703c6f03b1e85c797d7
za357087d98e5b1f45502e45892e5823d6fa4b762932009620038c05d74efcea7c3fdb38901d620
z36515d0824367e48d1bc182335f158c262d396cada6b0ad58add4f945eee634c2dceadbfb5118e
z14969c29a743830a07124bfa78707f3952b96b0db7af7c9ff36f77137d8c490c4f79328328069e
zd7d5280e4f95742c9841340368b9764f0f80413adb175ecfbdf3c40716abca7b8cef6f7fe92ab9
z6bd2453f1aef7f7899c5365c5c83793cacc7795c269413f6cf0dabad14d40e9285afde8c01a47e
zb61893788ec5060288cabde8fb553f21b02eac61ab0b48ad3d54f4d1d76508b22f0c600861b5ce
zcb30ba708be817b1f50f59c0f6fce449203e7355c1be55b662fef3f92ba58243d81537761af8d6
ze27d7864d2dae99372b2b75bacdc0437a4f7e011d68c3487a89759e3625548fcc920ad06471ee7
z2d701aabf726859343208b0a543c73eeff8406febf277e3babff437ec820fb49d6b78e73bc2353
z884917487d35a6cd06d7d73ccff5f0292fb3df6f439aded7c8bc5dd0187f22a0fe1ead93318eb8
z8c6e90111edd2a748769a8d92e19030b0323140a1ef01d3a257fd16256b12b03810bb4a4e82398
z2704088d587398546935b6339280ed10cfe93a3a5b7a4f04e0a6f073f8fa718c2f9190d76f588f
ze9fdbb73c2c6c983be7680e758043939fdd6803162983f37193ecbd51d83a9df901bce5c960f7a
z91451ccc98f8cc68bcf6283cc3f9b8b51e819fc5551032ae29e1442c4035c513e9c7b3b80943fe
z301a7c5fa2100ff52aed78938b3539056756c8be0eccb0271945748387ba5d649a64d900992ace
z2a404851521534f0875ce7edd0edd7b65a1912cb89b858f7af5e01b6c3475d5f27c6e38a8429f2
z304d3ecc5b845a240e6a0fe770fd3b222f205391f40af7bca99509434f6b7b1f7e2fd3fd1f8222
zceb6cbb08d53413f951d31a677658a198ffc7474b69211370a5977f22ad28ce06079e8d0b5d6ea
za811d9e821674fcbf7ebb1c7d8e230b92ea3f8f6320794237b222dc4f17a9a83c961dce15d8a86
zca99b1c76ac7e4fd5950bf8ab5a4c7fa73109b98b2d68efa15a620aeed0af4d81ab0255fc6261b
z95d52fadb5df4bc32af36eaa7ccbdfccf4e37a4962cb8efb08059dcc490a07554280940710c8a5
zb7694e7af6bc9a87db732fce9a43741168f16e1763c1a387651b1a9c3cb670b03ade7fd65e9c05
zc40f3adc906159a05c1bb22853318cddc7d3498e190852139f067fe384d3e9f8f8bb0b22414671
z85a82a0ae266e96a6dca3729dfdf3447bdedcaef943045de1379271c848ffbd75b4de1b8405baf
z3fbe93570a541ade8602b39e5c063c3fc3bca0c059f291f6e2557cb19ae16e0de9b6d6637ec5be
z9111b35421eae4f8b8544d47b576f8845b0de8c2733a7d42c257f2c5a0fc163f2976c455532775
z102143bf9b495763d37ebee81e3d2ef1ed8769226a76ecd2ec67079d15b4b6642009fcac3bcdcd
z232ccf7aaedc0b1da4ac7e056a54fc1135b79684629bf2a932c80c42e25da5655ed0dc9242aace
z9683fcb7614f6774b71b289ef6cbbda65b89feb9b51a6aec00697b833ef817c4d2721d4d9bf003
z6e06d5b89378cc5d5dc4b27712f486972ec733541f1b34786a2a4df8a8c5fbb24f8184b54815e0
z3084196cf39b52c06b3efdf3f08bbfbc09d66a9cfea807acca7b7c185772036377fff3fdd3ea45
zb34a4b8226f83ab0a5f2dd9f586c5f533993bebd3e2d7453939a76572622dfaaa9f04433107d9d
z823c76026144377d82d5204a4a1b2aab2c516b8e669ab263cea43da66076ec39ae7f668487cb4c
ze8110ce1af8d7e06d783c46441e78f7590b6ec08ca58531cc64b2985966c8a5e85bcd84fddab73
zfd1b387440b80e5d69bd1c64da4be437056bd9ab9b7efe1d8c6f660f61d3a1d354e2722fcdf427
zaf43219196715116beef2282bb73aaafdcbb4312874c88a77abaa114c443278b74fb2c07a68a09
zbd03b9105cc3057632340118507978f114dd673d9a59f3cf55d5380ed98aea7743c488b2cd61ee
zb9ce2713391f2eb6e1e1954241489381bec1578523c0b0ec373cc564d1ceecea1b8e192cb420b2
z4696ccfdf18f4215f22137bd808a567e91af764540f45d751c4809a83071bea7fe365f421f9d4b
z2c124c17b95a38d19af5c36ab58880e2d27650c10f6445cbfdc947dbfaf1557812ca17ed58dc34
zc57311795c43b007d034501899628c461fd20ff17dee026930a153e1bf7199418ad89cc210f6fb
z35f617ac13f3b42e0fe464d3d643e8370e717b12952ecb5d10931426ea195457415fc8307f8a65
zb1074e8223204b0f837e756da6cd49f9ef46a34beb56a2a7cc6b78e8831ec4a64a2d9305c06a7c
z157e5f8bf80412aa974870b0e10a1e84920a473e342c7947ec8685230d9f9f3c92dd28107c90da
z9b94e7e5d01f446fe4a97a72cd00da234a46a4e76c6f998bfb1626ea4e22b087c84ab8b2364a5a
z11a28f7afcd6351e9387ec6fe58c0ba5ba791e31e547b895049ffccdbff768749f3f58a4a7b221
zf6169247b0e7f1fad400b47cbe9f3c2336cb8a130b458fa6edcafd3a417e8e4310f2dfe4c26328
z0f93b58a06c73763292fc562abd99a61d7a5520bd4cb261c04ff4af11ff74741d958b047c651d3
zacfe6aebde1736fce0c9101cebd620807f2d2c8d76849ddee4bbc3f4b8417b32c1eaee7c297b61
z28e64574419422e27794b9ae960c325b260e7885b182b8c940a27e48eac01fe8c7ac85dd773e7f
ze27958c1c7f76aa39c15c4b38617c021e740be3fe45f6c317bab3b29b679757da533e282fc9f77
z55eb3cda65326e791b9e63eac086c50402ee929c7142c2754edc882d2777db1febaa46acb39058
zf5c24b743d5ea37b1c0f87ed3a38cdecd9af51fecf5c4f533b6ac70142bd567665d43c4fe0f84f
zb8da7af11bc13fd3a29c79ba895b25ca2e0068822750eadbda05b6b11e9c8ca234d92e25fcb253
zde8e4034a89a663e7736067ef7160800a01b6c537bf661d9af57b2b79cc084871720a27cdc3e99
zde5938d915c99f48395309465560ca399f3848f5984ea11bcc6dbfe2e9587cae3dbd290e82bf7e
z533b166d49c1de5f88492b4748f64473bc4ca34bf73aec7f8e80eccaf601d96216d6e23e24b692
zbfdb7fcfdc3b97f4cb9aafa32339f02928dc9a41e7cfaad7eec2681ce3db28068e3ad7fbdc09f5
z5cc62109b22205f23477624a3d274f120143c90240ae056b30ed56228addb0f504baa2a4c55a4e
z280704166699c05e6659358cf7934befd1bafd1d5ca232c1bbbe7b9a10ef3e613b3aa3170c28b1
zf4b49edbe5d910ff2c732465ff0405bf6f4aad426e34bf9fcc9b8038678a054defd85f86b81ff6
z8c397881af36a1d4c88d8543ff03597f1f090b1e06b4ca0fae61e1d3081723291c0da4f5b95ee7
z37964142de2386baf2d142878b45d9ac2868369ee0022286ab5f3b9c526dc867c49e74b528919d
zf6dbd69f1c20efa7f7d667f2955e0f5131a0f32e4ddc68e4d8d90e1f6cae1a2d1f6a5f8f7dca3f
z4cb4849c8a1b4d60ed05b49414510d3c4fb2343c7e627254070ab3f5e2803dfe8dd023ebadce8d
zd080f43b7b9bb9e9a1c001720a7f28b967e40b5db3f12de459ad5b56482166a4c2f8c1ee8b993d
zce3902bda30124b925bfa1f27206a5c8157058484394ef360eee4556aadd6e31a73df050c6109f
ze0aa349a31ebe1b95dfb26391001ae8616c54bc26fa466774236f865d78d34e7d2553a516f0a06
za885f26dad65b0361b973c227e6d76da08db58e88d050e89a1df228bc43b608c4c33cbbae94b08
z602c01e9f9fb3a090933f2b31c72df95e1865d4b8f5b3c0a224cff58d589804beb88b34661c50f
z84c72694198a723cdec21b4312ffc371f22a1624dfb52b989c9cc4686c9012590b2ec0a353ef3c
z99f45a2a23bd4ce115ff8f180e906d89a62b0897675a1789a0d3556d024185c4f63a21c34805f5
ze051446867001398096314fea5315caf82ec8740e62a9e88e9df52ff5897cfdfca6051b0d5be2e
z97749ba5e3da4fadc0f838d3a62c094ef0c91c1ec9de497bdbd7b40221eddedb0ca5c083440aa3
z23c36bee67c4e3c89914f5dbf39175a67251e3c4d66c139fd916241cc27eb1ef1080669f5e2597
z8878a01d56b58a2cc5c4070a0c90d778c3855bb9cabe991598eb025d384cba5c512e4037a0110a
z8577a44ec06f5be23979da0e6fae87a1a0be80fcaed434fd467581dbbe7e20fa656d06de6a1da2
z85781270a2958a40dfde8aa1da5f3b056b0514d5b4d9a842aff66fff12ccde2854f1ec4c1d239b
z709035f8beae8ca64cc5979ca7d25b7867463e5b0e22722507f08248bd23ccf99b03b1cdd5d803
z05cad7047f754c5fdfc028f1c4fcec149dca2b7978b80294efb8b5ab6ede62ad7be18e6fe5b8a6
zfdcf08b9dfda88e0eeedb0737cf7056f7f9aceae6aad6bdd1e36e46dd613328947674e1600ca27
z339eb9d7540b81f5891ddee74c7fdc6d8691e26a7cacf2d01877783ee683cd29211a09c2c2cecc
zf0af9379c7cee6d31fbf82c74762d21e7121fdc45634e7905c77c4705ea19dd5267d0e6c3eff9a
z6f8129bcadf0efa2c8c58318a8717d9461fbb2fc56fd9bf21091b533fe41de15108e27fe058272
z3854ffe6a5679633150314954587eaaf1229de2de5b61ca078879e7fb5bd318096d17d4a6f40ea
z1bbd4df8cffe0e40d033fa0dae8b93872da8fdc546c587123cb49446442f4d17021f52c9d2f70d
ze10bd95c5b4cf80421c932fd183258df2b7a18ed4b6adc1ba298b7349ba9a536afedd42752228e
z6492eef01642baba466e17a7f31b79219d8838e11583b34a62b31647bcdc48bf8d431b9c14bd60
z50bda9b53258998d77d40c82050777affdcf3c0537907836c8fda0544dd69973466fdd4960620f
zb50d9812a71f571f8c68cef78311080c7357543ba15a86724f67c2bdf651c126424bc7739af325
z8ffc4907f3dc3d8a7f21382cb2df3d9ed8467a7a8abab9dde675d84cc66e7b7e53e1700c9c50b4
zf2526f7f250be0a2ce4928273ee53d5620f507cfb52430750368d3da86ec2aeda541561e1cf874
zebb7b34483fa23c47af28a8ee98f730d8faa4ec795f931b0855dc11e9defcda9736dfdcdb1672a
z0c753541651d5b0b58af523feb7dfaf4178518f7429ef10c89106a29500c034e5295c87034bc4e
zb07338b5ae112f0683ab64dbe1da13486d192959c544c6dd5fbc4311133d56145db1f29ca7a3d0
z580ecba385d80ce1d98bd4053ef7c6473303cf24100ebb7c2c3d4757021fbbd7818edd12d6c28e
z7fb04a04b5eacbad256715f4a424c59ba7629e810cc6805e6279ea6eae426a2d50f9c4fcfd00e5
zcfcd1d9190629ba0c047fafb9cd1fe912e5b12ccecd412a0d2909331893c70b60e3cd026f161ae
z22d0ecf63d0223db3ddd555086f872881081767ef1d1b596e6590435aba0d37645e387636c644e
z270d2f2b882aa45a357ff5fe933e79ce6e55f0a6de5cb07120aab6aff4690f27b00322cf248d21
zea2c8ee7fc9000db079c0fb24b82586f1e7d5ef65e365c6ca9375875b6943bf29a9a694faed77b
z02cca6cb00ba8a7da672b3d0076fc4e6aa2ecb96ea34159fc7a646c9ab058116ef68ac085ac2ca
ze9c3cdfcc73bf60d9b23b577cd2ad972630e0842795b731b6a1e871f721194432c80fcad995b0e
z8d909fcec81a41b645da69faced3c44bc6379f1a19efc2afbb782d6d2caeec4eb11e37ca0316d2
z2345a0a0a5f005bb47e8cf17baf517e7e71007fbd3f3893fa81d64c7da2060a7b2b69e197a65a0
z8d62c7db8127fda79ac7119f1e82187a4fcf7b35e9b155ec275a5722cffbd678888616d1f9fef5
z59ca531e33945fdbeef8716a2339707514cfa87960df06a969b26e3f12b47d792d226731264beb
zffe32e294977840eb18d92a1b07ebf797d1b82373ffe4cafb4abeb4f8d72b0e144fe73b5fdd0dd
zf4b455aac8cd921f8e9ba744c00671ef44ab0f83eac49197ee2b93889ff2785a310853433b8b3a
z15a84d09e60fde32cc97fb85327f000fca5d2b82d824c4370c39b99bea5f0a0b629e2a46bebc4e
z660db38f9c76ff49efbf8d7559085ed8d10d06b2429b5921f03f90c73128079d0d75b27fe213db
z37006ed6f80612fcda06ec1c6fe520073ee5c17a207571e258e43f36d50f531786f4cb308e7495
z6006732837429aff6ffeef6b1ffe76673eb284156c41ed5bf1b8b3334045698918e00238e771a2
z0ab03b972862c71ddd2aab250c9bf52c41fb36e2f84ead2e2d5c201dd79ab5197f99ed31181423
z30c2b939bacf3aaaa5e200f0a97f66e3dc5269d2935675b67ffb6cf1bb0e6aa376353ba8290c8b
z249c3a6eb0df92f25ca5a313764dbf2ad5c98d9080c9240e5948e607b19c423756b41c49d400f1
zf1ef191a9400465275e1272dc46c17a25eb75f22349eeaf9b842e397b2595ccef2c2a418a1a6c6
z3740da965c3d7f9cab7ecb3bd387f977457d4ff4f9c80acadba7672ee93d7c8d406d7844401251
za7e622a893bb3902d3f3341bcb7fc572ac408d454a8d34e3539adfb24c3b22972a32e879ca8f04
zf724a0adac8a80b2ffebcfb7d3fc0c0a9f07eda450d2d7e6f1df3eb0a3df4dd0dc842999e45cc6
z95c8c7aa686990059e3e9f6b6216c8593b4683d7a40a78f382184d6f64db344938e46ab6f7b481
zad046baf79a0f31a29400fee3afc6c916566d135cbaa76522d985651ae548d417e7e5530f677ad
z9622788e047901ae012a1713583d34f9ca00a5328045eda56febd59b7041cf1139376105a76737
zab44683fa0c3d74861cb92743c7776ee30471bf00e600fb8612a2291bddf0089640b5300ac2cb7
zc9eb2bb3958c72810c87f470b08bc291bcb501f36fa69b7633ffe239e6684d1babd1e3361c87aa
z613f31ec051bb694f706421e76b4d878b186e8b1ef210ffebdcf78375745572462ec9189991075
z31edad59894a2ef5cbef14fa96ed0258bc19a29a8b5d3168cab8814b248c55ca67801f4f63f4cd
zd74bed8b07d633cf0b9296683ddfbe541a146578a38c592dffb6f0194dfc4241e0cd7aac2c01fc
zae851ffd028650f93bdb15068acaf502f800fb837050c495d65ca8e02dc7e89e342665cc630444
zf9ffc1750d12428cf16a79e69c5b130abb01e25cab3ea014ec77f7119b8ac5571af1704f4e8f8a
ze9bcaabfb7ff2c4fd490eeda9e3e22843155ca0d88a04f56d358d60c2cebb488711f764e7bf12f
z43ff43b9acf229f00112a61808380cd7014d269e8442c0d3abb1149b17dfb574361f48e74ccb27
z643c882cd8066689688dd60a067fa2eb029c7b72b3b43c8d6987b04839a3e7db66b0ebd3b8bd6f
zef62429a49b8bc53aa92a193e29c01e130f633c1510e92e85ceaee8b7fbc32bc1a5bc22f1e9020
zddcbdf9728d31a505f798df6be106fc5bff1583d659e651a570267dcf65c385cdd2c3aa8c7b4a9
z269a939a601bed1c38bd9f96f0a757599c2cb4b036ce22460edadb3ac40c1b4a971fd236eb6e36
zf1c3c5154d3f8a43b1cd06cf1fe6d5780e5b12d7368fbd7e5434ca5e35e5d69aed2a1457a20a4d
zf92785587819398420f8be16ca861294b29134069ee036a4c71e75d2a73865d431bab7aed1d788
zab0d21e1fa3744c90c51351fc0b6cdf208ec03cdbd5158fd03200d0b88fddfcf248d366cf36540
za2657f2c52a2be72e432585b8c30bb73611b94263f2fbd4c5775cafd84c4b8874e65c5abdf9ad0
z8bd42a75ddfac41672ee331d213afa04429f7d4fb1a6dde617e0660c11567c084386dc591ac880
z4c8f94e35b02d771525b552e24df1a035e4690643855cdedcb544f91bc6acbf027cddd1058a89d
zbd2be4460976e2efb500fb2518db0bd9096a39e119b128ae828dbe7ccc567252044cf9e1454d93
zce1a60bdf41e052e2848af8dabe697e75a1a2ab54ff6d97d33d25736382e96ce4622a7c50a1c68
z06245f7ca8cf2443bc02cab7775f3ae744aa1e2113332ad00450d801b1aaaebb05432ea413404f
z22774165c23423feea89c3889c3f359e42da6ec4c03d85ba9ad8dce1bc9bd627aea038c1a7a693
z29a3638e545a4da5cdd65432fab9813ba366c775cc36ee1e20853955f6159d05443cafb65b274b
zd139b60682457a711ddd69638b24063c4119ecbbf2b274fb929cab476d6afa477f8d4a426da13e
z2061ec4b53ec8143358e2346d049d4b8ed072ce2dccf8e53c5711db7aa17349ec2f5ad494e9a15
ze76bcbf27ef201a94d310b08c49322c7339fa5b500155389b2d646aaf319fce25370df55cd0533
z9372a29bebb0ce6173a3054ec372fac732582ff29df86ec36331e5f7817d0076130e40159d614a
z655ae9ca66c51b71f354b3f669e8c6ca654e0720d035337b9f1acb107a51ad1ff4a6c8ad36b8e6
z04f11f87417b15c1332b38e40b54cf29fa7ac0a839f71eba8cdad0f2999ccad922a59a055772cd
zffd161b5fbc00104cb280da6bdc70e29e2332286c337829f51ae12cbeb51eeb23acf5fbf96d295
z91469678664cbbe7f6f05798b8517185a646078e705690897b96d156ddb94a18b0144690fd99b4
z6266463357755d6bb0c2ded98d8bb777f39a27f3e9dd78aeda4eb125e841d9698135dd16442500
z0ae0460b0a9d604ab56f34939ec8c32d0c36b9f4f58c1ad02ae347d0d561b80ca2469bc3e25c04
z3fd9b823af2d91acc2a693b07998e8628041f5e66671edcc163be5e73c28843b5d5b711cf267e1
z613ab629e7941b6a6e7c664be6334a4d3073e9c3081dbcd17844b4f3926ca2f1fb6a82ad51a500
zc888327ad9f33206da75bda944a460d49f634430b7ec1dec47edccfd3829f39f5b748a8b03e454
ze8c655ed4648cf551b15c18760ce6b3713b8dabd06450f0798ada99fca89374747ee2523a46b8a
ze571641de03141ae0ed39ccebf0617bc30b6ca15eaa37076f734325a5e97a156f469eec0a2ad9f
z30da1fa6cdb72cc2aa765c9ed7c58e91a0e4b5e3f1ee174c4e10c9b96903aef63d25792e3e4722
z2ec9b549d350c857b4a00fca959de59636a903809c210eb80d862836ab050fe92f2b06db4aa2c6
z8a212d3a45a7d227ca8c77ea2b73aaa9f970621e5eba4bbaf94c0b8b907f58ae8f586fc62d7314
z6c19d532c72da5e933cd18cde7ea78d736601bee0f7347e53e53cdbc22e0a1f7e1ed55e22bb01f
z40084e1feff1d9b3b8442f67c1c760053ee274d9a29133052aff59def45ea45bbba8886ef1934d
ze250012086f551f2db29430dd2bdbaaac91cd1ed8dc945e2a7eaa3c55e9ec97c04ee7741f5724f
z902cb26805ecc15fadd89602bbfea6365e45ce4a58faec662a4c8aeb771b4be96e35d139ca9c03
z53a930a678fe655f2d411e5079bcd118c9695f28951ff0991c89eb4de1f302b1050514b2e443f9
z1eb007297933bbbafec32d8be5fc73dfa3efc0734169d60f97836ecb8ed731069eb98c4a050c7f
z477c67901bfa10aef770a5e9aadc39b592390654325793334693c9a1724eaf4359f18b62cbe48e
z9c7a82d93a9d557f4bc95eb653bd4817c1007e8b481c4c509f96e8fd3131b9d317de72986b4ec6
z08596eb9c33142243f81a05b9bbe98aec71058d5a90cead91ebcc6e6714bea82d56e717d94cad3
z9d088a3f8afb17c09c1023335df3f70bf6de76db2f620c999c4196eee9b79b36cfb7b3ebdfd7c4
zda45b78752d8440578eafdb09b0ba05a3c080f552b7fa6f7f4b6f7cee81390fe434e28f4a2677f
z4b4b88aa21fe9e7df8a63a0e07abb3af2a737784a42bfcb777c8ae2c4890417882aadc7c32d98f
z2df1c789bfb31da47c6c21ac468d20aa1bf35e8c7ea547aa52a702a63e062457989eab1cc84d78
zd9458cd62b9ac1fa4825b60465ddc4497f37897f3ca26a405416b7975437369b9daf5c0052ac66
zb1bed967de9b1e7c5266e98ae40414619fd8d7c5e794e00b122550491f13d0d66bd131e49bba5c
zb90bbc2901f8c6289e4276a81261fb1baa9c96ae5bd86aee2556b44faa64a93dd03fc67b8a19c9
zf7fbcf5e0920dab4e1f94adb77c297b7ba6dc0ed499662c7dc3180ff6947ffc143db8b5efc91bd
z2bef713edd6838a0f1bc342a4a50bc4af03ee04a1a51efcfa29741735565796d0f87bcc0bb1a61
z24d613781c425dcc163b596ca502fefbb5bacd33eb1248b18d8713f8efcef7746335969e91abff
za339164c9c24253234b2d3682db66f082eb4b7f5b20f74d93f8f8926dec02d981f1d341aef5a60
zdf8d52d36fab3158e7d24c6bab6f015a9eb07b16dbd62c5f4a1e4eafe4b4e9494984de5bbc6e29
z3eb14704948d249714d3ae633377e506a8ae4d79edb09d1cf1fd6dd909697a50f80d81cb496aba
z6ca939c0297b57d4c13d5f2bfd25e23f54ee2d24753f31acee7ec30a85d0357948d648584fe75a
zc1a40449e721bae078b5aea2b9e7344b4ca5d1f156567496a559728fb94f5cb1bb8adf2baa26dc
z869b312ca6fe11ce934521e1f650c31e415ae6166b40645607514d73931d414c173fb9330d4545
zbc976b168ee7a3e5de6eba814e7047c64c54304717167c7be23ea129d61cb96d4562b48d6963da
z96ac35fa7865743c2fd0dcd0bd4fea3ee64f130832f79ab0cbec009515548df7437ef01900a605
z1e18b760fa3fcde0a85c36af3a1392fdff1286496190b76a4cd509f3223ac58ef952954d6309d1
z11a546616bcc1ac0a949de49118c156d791370fa66d96a03dce143efd45a6be49865be84f586bf
zb8144fe9f202e7c08228805afc3cb87521877bc38a06eb4399b5853eb26d716257aeb2bd957c13
z94231fc06bd1700c76fcf74956d10550fc1fe962d94af7a8404ec84862e6cb9873aeeb34d44df5
z6e3fd5a43e7ffbf2f20cec7022f1c741decaa1aa7764e96f158aced16bd2e6905e97c5541bb077
za878ba15def33e5c0bb65469cd24192907eab90e3f93b37e4b34298251f73157c2988c653c3b53
z7a621bc3d8882253ecadb2356fb5c616add20a423abb4b00153b77e7f23b7c3a64af0bdc3f62a4
z06d35d41c4113581a1fcc47703092092bd31efcdfe040e70fa6bc08461cceee56dd4c834f8509a
zfde3d3862f1fe824088adbae256a5aca688a9d34c9e77b76c96becac8a5e293660718e44e13d55
z7a9c4071b67881168697c18933a614992b83cd0ce04b934e4b6e71483f545e32229c5fad52e710
z951e3a6d955b5b56da300b563a2c6b724f26812af156f9100f962418e3ba5e8368531ad9accf5a
zab7a941c61337659b3ba278e0b3f964e710a103d180ba1fdd740f98fa2f88c48714be38172f540
za4d1698ca9b7d0c0eb83c21e91b6951872a55af0ae921036468ea68d914554085928648d1929a9
zb36636d4d267c8e22848141dce0a89481338d28b1e2424a36ed7b70e4d2ff1cd20e88dea0cb3c1
zad0f3abe69745d83b62cdec4fa698580bbdeffd3ae7ff9b2df0319f57ec340667f6b80525b87c5
z934a64150238407e9a5a3655caa16e642bab71274afc88a176264ff3a112556dd39d260705d059
zcfb6a760a820fad607de9e998ae982fbaafbf60912bdb773f027967af772e5fed6ec25649936a2
zedb9d93b11f4abe359ed55cd679e3a865cc99996871242fc31dcdf800abad863354feb26d0847c
z8c2fe01b65df7ec656c372583f609e406e95341cdec22ca770508f7fd65de780bf57548df544f4
z91c639ec479a4d4ab42605a88d15de0ce3b4b5d7b4d94a6f9eec60635fdd9876627831e3f7c665
z1b982dbda12db34d5b213e35f3a2d18648c8bb1914bfe6b9eadf37f0908abb9d2a8337bd4fafc6
z9be8d95511205f59e141dcef8c9013d39746355abe784bc97157bff56c234aa360488c441ec253
z555dabc8dea6347ec9fee829d9995d46981f5cf830e06f396abc7ad9efd72096d0e1ca0cd83924
z9386488436b1fcb6968b721ab0d866bda7081cf7124ca052033a6eb6a9429dd4828a898c011ea1
zeedbaf14cab0f0608e49e238cf0f5e5c4b77894fcd10602d1c40305400cec2f17ef612c7b69ba8
z61d24c3b5a53853f762cc6c76ffb174027291e83d84302241f8ab20be83db11a3556957e2f57ed
z430afd9001e149fbb2eeee49b5848510590f717a88fae9836d923665e97703d675237a2606cab6
zf289be8cbaf56314954dd1e770176865dfa78908684551b190a02ccd8d44f415947c12048d4799
za52d1f71ca84132f6f5a14cebc5e4af695de77ae69b32862f6a1ca49fbd45035f253dd11ef77e4
z632689774790010cc68ca7e0a543cdda2bd97d5d98e71021d87bd331e99e63073ffa3f8f6ad5a7
zda2c4280c7c092ac56433cb61342269f4c4c3ae58019453bca38e1288c57f44ebbec601ae46416
z6416daba3d84aa353ce51ea70fec39cb903f231a1079bad6213049251c5cfe6ab675f87bf0ba6f
z55566c3621f49efd80ba34193d91a77afe710d1d27bc136644a148b7515da1b9cd32aecf70222d
zd93184f408fb33a958b1bd9ea460a7972af22df236cca15464a31bb3c24d6144837ed9973c3711
zdc6a7146affe96133966dc0b77d3f7b8a18c2d44958aff721b210c64f29c1b021ffa39cf00689e
z845e65d4519bc94feed824dc1b0146e23a12ef56babaafcef200bad541aeb52feb678626a3e65a
z19bc144a52d9fe8ec08649f753290adb186db659d8b7d8dc9b86b9b04a447370ab13cf8ff0a9a9
z0e1c34208792a757b0edd68ac1ef0526297c0e2a34bb0f79d476e352f77045b3d8ae486606a8e5
zf37d3fa23b930e4ad6a51ecda1b8f2bdec709afa0ff2634c508377cb952d8d5dd9cdbac4d52693
za46cb43dbf52c3944f62cd92b515c5d4558a32fb2b67ddedc572584b6231892912d918e910a232
z1a8e748b3aa401db7400b7002cbe0a4141d027782968231004bb4bbce9b858ba0237e0935752b5
z73209eb10c6600f2769dc5d735839ac781ab7426c1935566bc53eef6bd372eceae52093d0c8322
z921d690be21df36ef0e1a47b4e3905ce20b798556e83916f37e91e4fb729cd8d5cc2d35ecab5fc
z7b2c135cdbbc7bc09a3f57ed0525e45cc89ffd76a2365b5050baa3900b7a17e5ff79f97771f46c
z629e997cced4c43fc9e18f6c8bfd407ba526246835943754991b7d79bc42799e0b30a2c197afd4
zdddc6686647d4b1ac3a4c94d089cb1d3ef8e997a3cc20deb7c7b0f0bd681409a93207d46e28671
z125b736c9211871043509abd4363ccba3b5ecfc97d07b1c48f0a528d3adaa0c1c18868e738e7c3
z5a315c7943d720fec34a9033da54b5ffb83fe734e65bdad623a017adf82a399cef9dcdf7603c09
z125785743c6df9b61964eba48d25398e029fb40bfac2a1fd939909bfc49923a0a24c794688a919
z622b06d72d3f8da367279ea783c80667791d3edcc7b08ab60802a902eea9a67ba6276ed0eca18f
z8c4044e4e3ddffc7b40932f54f6f077e3e70e90318d8b77903957c655c06517b3b35701c49a8f9
z25d54c6a0e4d770bcf3344cc52af2379a9a3d4ac965f41986e3c88a59b76efacd34836a9c79589
z3b3acc803858ddf0a4ee0579468a2176945cf50dccc6b289917e2e57020b7c06a38c0ca3ec0600
z49ed51ed3fedf095f3c6c2e2c69adc49e138f279c74db6c2020c76e22466520aaf050a0b370dda
z34fce19dc604b6c4739b6a1ed652a3d85f182be7a5c7818796f556092296fc90c12b91e43d345d
zed2ace9dd3557928881522ab05dcd60724c5fe08ac6eb3a3023ae3cadb7e355989c806a2f9a4f5
zfad66cdf472907243f322351f5b7bcf1f8f57764389658036a43e8fc9919261dafbbe9ec918e90
zcca5597fa57c770f0fbb542e5e8e86efbefa00ec3e66e686ccee4f766930a6474341ada8edc5fb
z6acbaa398bb0e116ee23fb9b8ef05e2b2a28f14500586331f048b4914bd296a73e1d1a3aaed40f
z580c137601cc85b9d29d7b72de21c7245870d7401270edae96f0038856ff014f7b77991a63adb1
zac2b1ac37cd6e2b2075a17993def8427c5a25631e2424ed696c81512d7164b46281b2b9822e21d
z37ee3edc564723bf75e69b3087fad737d5774002a1acca6f75876ed9614874c1a91ba6dff1d581
zc0181e3e8659c5b38cd4d98626e46d6c91898b9886c439db0af3cac247b5ab4209a166d6120c5a
z901b60374c7d5f50b966e6f9f3c0a28406e58964cc519973a5e9f91cd47aaf6af1a638b07c9883
z2049062dc03375f53ad5da02086c6f7df973f7d88c02dedb6b5d51f37d96de3a6b4dc07aeccf10
zb6e423b912d36e4acd633dd045c43627d20952e03ebda13466cd7cfd92ae7608211b012882eb92
z006263adf36df29afb2072af1d7350211b7b81d580ce291ef5146c4b5dccec5c0e4b0d81475fd8
z94ed8fa7d4bc9b752c164ba98b334f2dd29e6a69241b4a6f9f4ec1820b745eaf0216f1fe362568
zb07338c77302a2d3963c444c09b654e0e6b28c11ffb7fd2785472081f1aa8695bdec9fc5be9d37
zc5d9db79e6aef649918649a557f15273369372e1d144f627aac44479c82fa6cb3ab3a2ad0b7db4
z7010988a71f7667776ffa53d2227ebf562f48a42fee3632f754799ce0ff8651257681cd18c7a0c
z21113706a4f085b70a6b87afdaeb31e2c0e72aa2f00e0f897b7d402e1452354900a999101ec1e4
zcbd8aba336eb457069e23506a07dbc54aef62049e8234f1b019bf6482824c02eddae9eec8d54f5
z7adb8a234ba7086babd7f37624814dc2000a9e8f1aaacf6033b9fa2e008a9d8023b5617c439da4
z98cc2fb3d47bd6dc30e3d30af71d9b96189a35fb0c6c1e9bc805c2f6af9ea22bad394cb4f82291
zf2163d30bd6b6bf1d2b5f1e3d6cc6c747fbc4dd5304e97f9b77c8a50258ac32499e5e101ab650b
zd2829bfec9d910ae25d6bc84af9ce2285a189c0e4fa4dd90d1775b20641bb90c7ae2fc28793866
zff81af16ff819cabdb7c16300e5a68416b7aeb572e25226efcdd6f2d112883916c67789713519b
z044721394d6b1d059a380b8f627c70787186e10cd73009c443f83cc2c1782aaf44384358df4897
z1ce7ef72ff5339c6482243cb411cf11025f4f39ed61f3f5d964fed9b58f50387fb8655f302cd64
z5877c45ed8409cf58186a69a8716fd6eca5f36c3e2fe5eb11de3809b96faf20ea08cbf027233d4
zb1e4b9494b2e2b69453296fc7e14c2ea6b397ba61c21bbfa8889ec6277fecde2ba8d32454e7878
z3afaede9431c25756e23f999770dda6c78395a739951a948639fd902a5236fc4bcd2a109aaeb88
zf68b006d2c25e1a89c51aff056d35067f38d7e6f24090239c88b64cf2916a2921a322293d30b36
z8da5656bb0fc6bf0f8b9a0ba8a9735bcd000622d4489a32a47b7f84be6069b1b7f33615b27bc47
z3bd8dc915fe78f30f462196067c10695e168d404acaf5b15f4c964c1d7ec9fbdd68eccb0fd8f6d
z10addd4bc9dc89b2864daede8cb785019b76769014f1063ffe4980fae371aa5393f3b2fe499887
z035197ff52b047705c7f0ccc090db11545a323c97ac3a58baec0d923d5f46c41d5e91a6b22a294
za3bff74adb791baf1103f93e58ed4ef1feb1ab7c9d38fef728b160b00af2fea00748928b2f24b8
z389bc48e99be8ff30e96cbd4f22e7fabb85db9cc3b7e6852a96cb6b26b04a5124470bb11584a71
zd2a459b191d17ba58a3a6f7b76521c1a62e3190a0676c3410861a4b433d58eac76af8eb04e9fa2
z24437ee34b26143f181145a98e97d39d2dcf53da4d349a280df9860e396d7da4ee061a834d58af
zd836b3dcfbe8282faf23f776f3046454b657b1a9d7a89c64b70882c1704d1716f6935067ffd280
zcecf9b8fa71a37312deb985f498e708862daf7de513eee5ee2de36a61186d2a0ab829829f24ba6
z8413fd2cd1accdfbb6c6c89066042d6aa41dcc683732613dfb5adfd016228c6bf9c6970c0a1f46
z96451e91aa6cc9af366642d92fb8cdd33f189779829984c480961e318661239209216a3f38d360
zc29fa2e169ffdb0f671f4a5a9e1ac9f172f559c1a54da6ac162b1a6adc94410304ec5adafe5713
z6cc71064050765bafa6162f8988ee3fd3debc8c9475a20aa6fb5594a71399f77a0735eeb66e443
z02cad2d48be0ced316241e9361ae5b498d1ff9799896ca657aedc8eb5e864a2402e1c77c9a0c94
zdb0a9fe4c7a87d1351b04190ec3fc457a7aa9e381009a12e2821c6e35de6e6f1584239506f00c5
z2d2bad3e9e6604cf0f20588f43e8cd3605682eb76f3eec833078d2cb9cf1564ac238afd8311168
z4f1e9bf9736cc364826a040b1fe5b5fce806ea523803687e7c54a4e51c46b7666b67de9bfd1151
z9e2a56bde2a8af83fa0fea57f06c9b3de5785dfea8e927d8ae7c7a3044bae825ed8a5d99a4e4f7
z23119ea223dd15e657ab8189ef67900da4cbfaab71c16a03ca869e4c5738e048df13e4832dd1fd
z24aa493dc70c95bfe002eca7a9e6ca999a69b26314841617c7ac0a37847c06c7de7a782544f369
z6cfff00a5fef448da8552efdeef62a2c7adf9b560993a930c18e61707db989259ef4baded4afc5
zc0f584c10260719007ab416b3d438c571bbc5072070c2f29d283d2e4ee134f17a358dcbc13fafa
z454f35afb807b659b7b121befd802b68da8306d82beae559bfc182d9d12a7fa0514f21730ba4b4
za8897a050da5fa360e8014222908b2f0641087826c4d6b7b1b3f93147d884d8f3e21db055824ca
z5e35e683f3d94369d19c25ecb6634f18bf9d68e9a0198d6f6e7b4e32f0bcb1606ea3a0713c4f22
z817bb460e848d51e21839c482be67902fbdde163b22688a2fd571d53bdd72a31e4f1f8df237240
zfb0ee17186545836ebe3f4263dbe49e9500c03eaf1e8dbf49afdbf1343fa62f9fc5579356d0f89
z32663f42a6c6f281356187f1dcab0112dba1111fa437c6ab6aa680bb7c83e537457c00cbe1f474
za928f299042b967c2213d0876c9878fcba541e52f301113720859ac73b87209cadd7b2719e4a6c
z0731acef7fea1dfd43a720e5868b31296815d1ae5f7fb778b754dfad5231f256c0499222e941c3
z9a6ea8a953054e555ab3d72170b7932e05890164337c9c386efb38f389db4ef68c008f770c3ecf
zba1b84c330dc330c468f255687f3ab455d897b18f89cc69ac587026b672af7db9d1ac5357b9955
z4a5739c22198166262b94dd16648b6503acf8d0cffbb63be4291423e0eeb8950fb475b73a121a5
z618b3df48b24fe0b066303e7da4ca644fc5924194a568087e04c9d9924abd35583943e2b44f7c3
z671ea597c9c970d88b64f9bbca9c4affd584969e19572bfeffcf1cf87cc5db45f062176f696255
z65d5e9b8c075a6521061bccae97ae6b318e7de166a159350bc9b72bbea07bbae732481f10ba8de
za3dc5338d7d52c4734ab151a506d849ac0f184a6318ce95bb88627333a972a1e10174d9000deef
zeb98cb8a6c5d236f63265ba12b99a24e6af8e41345265dc5f477725608ce0bd367c0c4c840a237
zcbf5ebbaa5125257696ae1b07fd10b2ebec6bdd96b7c3b848c84636c81fc98e70596b191ebb82d
z6d50142c5348d08b8c8cb62d4d1a9b6efcccd12543c85b92e08bf1da525b88953f8c5027babb00
zcba95f87d848fbacd2325c8ccdcf35fea97d6c168b3726e038877137d1a5eb01da4a30eae7fe6e
z64229b226c34a0acda8e236fac2dc688aa4c3164beddc4e8b7fff959a30023c0e4c940e844b477
zfd916b0029db3c516e70ede8634492491fdc6805ab4a29fb8d7075d6771ebc3da1987a6af75ac6
zd45f7d1e15d1129eecdd95da795c27453fd3dc458f9424da699b39cefafb7232cd676751a4d1a8
z665a9e6ac1f93ffbec9b43bca5a17316d7499506415691c9f7e2920428ba1c182ef220964f1054
ze6c5e6de45f4e54f9f9c4346d7967001b413a7303c856502be9dc2201f4bda066a98a31314489d
zee47483dc58ef7f1c05d93d1040a304dd80377600cff6aaacca0aa6e26a4a569d9ad4633f49d7f
z340ee44c1672f89523c5c3d424320028c2b0b3fd183bb9a7571ca713a9e58e43da7b0206aea574
z3b3f28b741c0557f15057e89ce704665e1e56f07ed453c697a7edcdd59f1463cc8ee843ef7c8e3
z04c2aa06ef54e94b62a4bfe9f5f5bd674419f4ca167ea0858c972752fa0463afdeccdcced5ae76
z59566869f45bf7a89a4d672132a7c22390e2903fac2f8b02f0a14ad367eb52decd8b77feaa72fd
z57098d014688c0730a01acfc3d8f09e18150c0111a3191fde907d9bc58e6cd467128a714088ac7
z94019b6c66dd9ece400e9b421615a162973340e3462eb1cb7355bb28a228b12b287ca56b12d4b3
z7d636e12dd3148900f7ab43ead68bfea0b0f249be93e771d0e7e52f22298082f1145e8e932650e
z39211552502dcbde8210079eda463698b3a9789bbe5f008087cce6c71e8b7f21fd4bf4c7d7f729
z64ff24993ac495849b16fe1c7638acebbc19a875be18611846bb364f6b0266014195f9298a9092
ze8e114e468a37c1e69d1ddb3ac9d111b8dbadca60001ef9f77a1f468db5fab24bdbde223fb67e8
z3d4bb3609f6c9687605d4ee52dcddc19281fa96bab284244519535c759dc00763b864edc6cf1e2
zfcb6ecceb4427e360d146d78e5616d799bbd32281afc267901e240c15b89ffec5758b251130b85
z5cf48305ce1d05266a551b5416708bb9201ab7e90e3edacdcae2777717cdce3e381b3438cfacff
zf87c00fb586bfc86f72de588719b90b673e7d07f88eda5ec8816f2619e0df4d26da34f0e6ce2a3
z4e8665ca61dd67d01b4a102f7819fdd046ef578153fa647a4ccd2766efb0dc70f8ecea724d433e
z1863bef485bec1c56a68c48ae274c383b98d83a5fe0e7614318ff4267718bc5e5952f2586e3c8c
z9f53059367bf63658e77b333b7a08ea2ece339cc6afeb3b718db999d808dafde5f531dce986672
zaa08440eedec265bd276ac7e61721cecbecce2df70d0b8d8d8fbc32de2d2df3d72f831a15a654c
zd7b15fc4edf6262a05396e9eb548726e65bd302eb2439802cc530f8fe89ebafbae580c4462bc32
z1b7b737a05a637836ce31f651eb0c865fea442623e7c61bd246402a438b113c33e68b2b648ab3b
z358f34c9fc15ae8659c7f39ed944dcf80c50a995f433e6be8710f685fa7bd23a89c996895d0680
z80b0f6a9dd385ae0658e7dd468654ba8d8d71738ce185842f0aa73ec41841a88d8cc00faedf95b
z143edbe76ae11a84370ff04f4b3e3395e494b7528613d5f9a97531df8b8b031f06271034fa59b5
zac448dced8cde3daaea27c974ec3d8fe88bf2c42e7245360de3c3397abca2f8ec3c775d461d8ed
zfcd16cfd99dad8ab6d18931b61240cc6c266f1dc9a101a205b20f428c086bd4369a23180bfabdc
zc2ba75ba1587af3459ed0e403d241356925d66ecc1730ccdfb8ae0f2d5ae041931634a08472f75
z28e8a85bc796db8bb3bf2d1f8413f5cde2812d686614c63973b56b7aaa4d6b73a383ad03e94c0f
z9fcd0bf42d15e47458be20d42502e811e642eea5569d8b4edf28d06b057dc98eaa85591ee674c6
z8d18657a77a0b41b498a8b17703507575128f967fca54587c6e31742f80985daa39ed9ad75e8e9
zfbd3592fbcf89504058f514e63fa0f6c4c9de23b7170329f3e5d76cb3bd8284b5ee1886aafff0f
z7a4b20e4729943d64aaf00c975feb905a4c5009e80b9f382d77dac3f92cd3b604438c2df7621a5
zd250834f1a39682851f3931d0db59dd63a2c8cb7653b55f83c48e0b6253ac733157da7e477cdc0
za83e0035448502ba6d52791df366eb18debaa5d998eff2c12b481b5000f50d09d6c9f6111fc470
za4201a5b801ee7c0e61b11d8ea2c87441852bf48144cb66c15ed84c385ec708faed00070907f33
z91f840d2ceb24c79c965fe1bf641c5d83abbe0e8ff399506794b95f68a3e2df7a96519d7748025
z0bbe11b0cae934df4c06e007c7a4d5cf37c37adaaf3d9a3af41c1a0305349458449cb7b0944b41
zc89b66636202b17f53903c0588b58aac4e794aebd6ce56bc11e258153645fc0c8fcc1fab0bc121
z9f815c9c5fe18027e4c3d5ed96ffa877bafa05b696d291a27e3068909bba8b7903fe448af82e7a
z7087c61da626579635b7e3c9ca4a92d08d411d8f0a2fad8fb84d68b13b2243eba8cd231548c709
zbcec18fe656962b26660acfcd37947766980d99a42045f0844faa65603a6d300a978085ca471bc
z9fbbe39b4519fc1bf5dc75c09155c2cbedb881971cf87aeea67920527008553fdc8f10a5dca48a
z644a8d64df1f243590e34cff550553804ef9b268c58c904d0adf17f9e0cc531cb4037c2a244d0e
z9738825208606a9fe350db521eda57050a83430e1a27ea0c824dc08f0f7396b4e58ac0c57dc454
z3a35b029a9f16b64a590305b048a7677cb740bd7d62707adb285da759a4e9c13568a04ddce8616
z5f222ffc989ca62feb6fa83cdb634cae788849e63c75c35a8e18c7d190fea201acbaf57039f6a5
z7ca86690d475ee140faca6eb600fa0e5259e93b957c63e810a5fbb843926e03354df355594bf39
z995cade7d5cde60b4848a5f3c4a5230e27019262ed2bdf98b72121e13131c9e56445948ca74f0a
z9325376e22968ab26b92636953b74c6177a65302d30581e257ebcebe7beb39f2254fcb1d484191
z1f1fa85966a3289f1e0f566833766ef3c5c209b8a197b11a1ec7205a24961df7ff4f6ec6870f25
z985b666da6b9b94454e791f58481985079e9c983fc3bd00e2d36e1601372abe399938ca0d189d2
z883e1b105441e496d8889eb64d964f79a7bdea62efa2e7ac65245892d6099edb54fa540ab197f5
zd9dc9e1dd992cea19dedd8abcb6b772a10b4ca36ce4ff9973c3887520081a47e15b0cc55288355
z225895a940c3272d0c782a81b80b3a89aea902f61e7f06b3074d9b1b9073cbfcccf6eb6ac261f9
z145cef6dcd5a5822e348bfb9c43581a94c66c1c25d14d3f1664b0ad7af77b3617f02f1e4ad9ffc
z8c4243e6e899ebf9c15263771b171952ccd622e8dcad17413ff80b6852326519bd83198f1053e5
zf12f072d94659cea88a032fc091aaed378431338b6d7088c41fad8348a07742b8bb674a95b33b4
z06394de7fbfa77e669412a6dec458cba12317702b9311fcaeb3a929e8f5e70b05b448307e59d70
z905dacbd9f8a5a61a103db11f9ce9aef18946267974b736c6883674fdd758a37b89a3904f55a82
z39fa002cbeb35f04df76342402cefc97e3955d453460ad37c5ebb6b68d52c0b5a16ef0e964c38e
z87f71b4b230f615b14f36088e77c277f6f8fe051ecda11791a07493990da422bdc44f505654f41
z87223506942e52e0b36ef3c5f5791090680518399d956814388a7f985bca04d8c2ef47e1fa5a0c
z4c3a3d6fbfc877698ae3d38c2a56d12ff0d7e4e9140b0d35046e7d9fec7ae8a984101d5516c21f
zd1ec87ae572461a75d929cbe1430ba4272d91b09c9e00452cfb9bad81c258022a5f13cf1d26b16
z1dbfa153bf255a7391bd8f17efd89d6e47f38cdec8466a540e3a95819fe642c13f6c12ec316932
z21c14e291c0f0cbb7ca400ebbd82625e2913bb403904f8125b587fa0f80c18b7c411e174884fc8
z05649667674fdbffdd31ffda79e354eae89a03afff5138d58164454c3f2e7b45d974d6efccca1b
z2c3ae2dfb2957228c6073afcf68ef07aa9f7033d25e7006a3fb31b62f4f88a469109d6248340c4
zea4b43a40df575986f8f1cc964e6b9d740000d66ee57aba232f789167f74c3f506a77b05146193
za22885f67212146b3c68562f83ce3c8fbae39fe3a9473226f089a48efdfd2cc657a73353bae112
zef52a7ce56d8cdc72585f5dc903eccec84179ca84ad33f8f6606ce1e08c74c9d980c328290e97e
z7560acea8c66fda16f65bae4063e016e87c3af7f4a18149cc15d554e9834661b144f37e6ec5dbf
zd8f341d0ef0a1d1b54814787b002fb9b73e2519c391d9b1f9171ee60383584f016c077234b6d5c
z84fd130be115b935f7b26c36791707d0730be426203d63f5b18f65894f79a29f3e0918497337f3
z4c3314110f389718e3662b6bd7738bde36d83e15311a5015dedbaf03d339916b3bf533d6b2df44
zb8276d50184c3b62dc3fd97a222ea09551cb4abb66c7259a60653c7887680d3581fd3381be9b11
zb38f72c0a3e346052d45b849d2f4ac0638f074f253cf8993afd2acca4c6ee079369eb601cd20d0
zee3ef4a4c812c15145ebaeba4e045fed92e283bf7d0b4ca0592a14cadf107c56e631aee239d831
zc7db3787a472652be58aef10e110ca5331a9c3780d205f0e692ef91c82467768625cc7b3219eb1
zd01af5521a860656b5b37ddc7d2751ba0cc729a8a5cef64a89fd16593a2954807c64590c051096
za403a37055db0b51ebdbbc9be0c19291c811423398e81b20644a93aa18c9b3b7d63222ca27a558
zd400a964e97b295783a82e961cb5eab682368a1fb4791f21076409dff2cd7c98c9ae56ffa880bb
z035da5c6d4dc0ae8af78cd8942970edac41ca4ab24f0e336175b3ee42070743a6ee1afd03510c0
z7647081edb074970cedb21494f2fcb482ba26c6bbc6e800345514baba7695927e200933bce88dc
z5fff278da1ab2e85618b2dced1d2440b143d4eb1c521f1dc9cdc6f9f44229113aef2cccabb3487
z2987ff4868ecadd8308c30bdb4fa8fb6c6c65be6d8a0a9da0163cbf5d49171ed875bd78e4f9e4a
za16fbf874b4b589823ecf20f1a4efd0f2446c05853be2a9e7c3c4dd3a7a49cf6d6fe7819d3b294
z6733ff7fce5d0b982d46edf329e4afda35c863b47dae6bbad69ff5f960564c8a1525020e23d979
za09d906981302a67c06cdf993645006aac7b688b9f329aece13361dd3c4160cc658d2115c26dd1
z8f2297a8b91540b48ad7808d9bf4c3494a93b163868291791bff1d8ce163d0e18ad32af05d0661
z405ef89828e8adfbe0c5c4aba89c2415a50626f659efc98849000e75e3badba1c87a76a9f3d8b8
zd60537dfaa3101bb534c4dd2915a31ceb106307db9b7a804ad6640c08cf18792ba110ba458fb9b
ze632a54ee252b7fc30ea675235794b2937c5fb043e265c2b8c18e8bcc84c259b260d32519828c6
z41c2694958c995b503570125725becc140378c3c6efa67c6e5b334f768d5f265ca2c4190821387
z106b4922f589f4d2ee222038bc040281bc3836daa99df7fdb671319e842ef7fcd743f3a217fae9
zc4b229eb3669e72827d3cbbdb350d47180eb97454407c82fd90dc0603033b691877d87cafe8840
z94d8bb69f31ad4a13ed3fe617bb54f08d534a9d1c80f40ec9f365dbcfa030deedb41a93a6823b5
zf391f147a05d6d7675b7e5060efc763530c84303328adeb772e5243ca1c89d224aa5e76c7f3bc5
zeac2352bbf7e05f8250edac0d0d5a465c5460e6290134b1b8109d268d1ccb86c010a1de4f1099f
z96cb72029aeb80516fafa457aeeb0e4ad8731ee5fb188a926e619bdd7abe4543dcbdd586889703
z854c279d6811f70c6ed1944c92dd73f359e0528557c90efdbb23e1d4d3ed593634c2b3ce9bc6dc
ze3cd75480250b550c94fea057bc5bf27d50b98500a7206cc7d2979ff2742f75345f338474a7e54
z51b68b7818341970d93d7017c43b23423f2ec970150f43096c9b51896344f0415ba58e4306e4c4
z9058d2ca7edecb9f6fdad854c7ea3b9276c7c3c0cfc2b1757154ad3e8eafd93f87930982207ebd
z1b10024bddb9c42248aecbea116f3e9b9d954d3762c71ab07ac77aae55e8c40855523570e01eb3
z22ff3765c5722568e35f4a295cb51c5006c5364f068cb20903c1b39b2e37b93f3e5a66e07cbfb8
z36123665658eb27b56e2158ee017a412d6b3ae854a65ea496d8e2905b55ebfcd1908abf90a2769
z1933fe992cc9a4baaffd8b2d16a46edefd7398764538c05c1b544863b69e9fbfb17933a13c8a96
ze23e4425c12993a7d725dea493591a577dfe41a1e1745f9444cbf28705457a77ee937096eb54b6
z639323c643a234df24cf069ce39c605903408fcd236e71d04a72c728de46cdff5f69afbf4d6687
zc931cbb3aa0bd547ecb825455ecef6e70232474866477b708f759799e57a291ffe89e17637551e
z2e52911d6bb93cd2fad0cb47734c5f751a192544f29827d0cea9b1de8472b459719c6125f500a0
zb78a18633efe3070bffd008c3c449171c97b9a66b477146955d309ade6a525336b0400f9128340
zb8aa87daa7d7c32fa56feb1c4c6338a1b0f63c5f49607786ada615674a014203d80cfcab3b715c
zbae764062207839b68287ec87592f58a72021cede45e46e307c37e5962364d6340a122e1da007e
z3a16bb815802622a699d8d111cab3605a401636381338e84d7220d9c8805ccf4547de2aaaa25d8
z71d9c1c9babc350cc39afb78c289427095ed3fca04880d4e97e2f1b40c0054e23e2ede0d7b4b32
z0a61359d9472ca798785c26cc7293cd371e072133b6bfed000bd89e2c3935077324cccabdd3954
z6712fe779869e86a0e21805484971cc900d3362a9275428cddfe4edfbc77c92d83e932c10fd4fc
zd70e738d4f2a70b24937ffdc764f05dd86a895fa2ac85d788f23320512eb2bda22f73a3978de43
zfbaa3f33ca5bdaaf34d9881c2a3ea814ebb081982a708c8a5d76a319cef231be553a11ad3386cf
z346dff5e12770fbce9d60f16c2873065b7721f1fb4ad0ffa4dbb8031680259626c136bccfb19fe
z2b03145fe95f524317e4b56fb198426010bc6d9b5e3afd5ab0523983e06f96a121cae3cef43fd7
z478575e854a76de51107946f3c0380e74d6e17c3cce88aed64971abc99e46b39011d1fd2d4881a
z18923aaf4051e8a4899b9a6789ce9121fc85022200f2ae5e951459e178da9f42e5704a27b6ecac
z5eea8085373a1551250cf80677bc98e368f9227c6db270d4e95cd8779e880e978dfd0a6f13c48b
zde9aff5d59da2a8f361d8e07dccebf864d227640d4b3fe680df14b17db95be0e5cb8f1f8dbfe2a
z8e021e6ff7e5a2e8062b3fd977ed577bbbff141f7ea5c87353a73839d34130482a7db86e3badf3
z28bd2805eba10c42d891d3f3b45afed93494931b680aac47531fb7d8e9975d1602ffd7ea6c39a5
z3a2e24e3577ade2db06f43b63d18d71b2c7d06b091e7bcabcc9401fc73b423d4ed04cc165df617
za8ce09dd802ba5eeb5826d5ec31e80f27e03883dfa9920827ed14fc20853d7c8143604eac6995b
z4ad506817df6d7b7738a12f2e6548e2d296ac82c6ca90e336e75d3d9a323b2fe4e31789c00013e
z06c9bce58891066e30aeaedd36487e618a9c045b31b8d3f7121ebe4c014c2e8f8357d88ea996a5
z95fb9a595a2bf404d427944ec9090a99111d52a007376803461c62397ed106f9757c969ca60ea4
zdfc0c1882da5d9018f2ea0c9940aece7f7ddc4c97824753d5d1b3e2b624c5b4aeea6c2f557a964
z787e05683cb557c95c2c183dfc828f7997fb91a751f640ab14af6f277824192d21566a0d48e08e
zf7895ccdf4497c4aa0678408ceb932a6f1c7a4583b51d16b2a0bdc947799ccf953eb3619725799
z2811bfc56556c03706d340ffbe69a4ce9133871d63b90e3f85c056bede1889a05c77b99a43d0d7
z2f8836b846a3cd41704fbc71f29456cb107027433e3d975bcfef8b67ec239ca2bbdc08556dabf5
z8a6cc2f06f799467abc9d052155b87df7a5460ba66a942b304ebe3075bbbc024aa73ccb07c1cd8
z1122b980ec91507e3d7e37bf466d8e8369545354f2720799e7f953ffe779d5c769d84360db0b8f
ze1a0721f1dfc42f5bfb6d2f850725f324389978dae0d6984cc89108cb7ab5375fb489a0dfbb4dc
zc2856f223ad87372c370c62ab2b0480938047dc219e5060664849ad8dcda6834ed4d20c8a2c03b
zfd8e5576436c76267d7ccd4ba6008353434a6b95ab8346c60e8dbe519b7e135ee51d5b6e1624a5
z57432f9c4bfa7da80192a83890b30686f562549089f162e3810d1ff76f274e629c0d6ff44f08bb
z9c86964a12d9ee9eff40251e8ed4d9a5410e7622bc1299534dc07076ce16dedc71e00778cf2cf7
zb5fc3d01cf595ec7ff03c79dab9370efb84fe775ecad99eb1448e8b96c1378498cdd0718b807cf
z9d65aae7dba07bd86309db6b0fbc45fe5670d6cfdb26e0b561190a222a13e9cd5afdc256001059
z1de397c1082b5745be730a223c35ab080e4220377f52c4b9c57ed0149fd57983fc9b3612aa2193
z3842a50f29f7bea5fdd8f0ada9a7f002308e4ad6021fbb491558286dbdc8af1f9597faa9bcdc3f
z6aec4c13f58e9b119b0edfbe576472e5e6e9d6ad0b1b150ff55f26222521da25e1110ff2fcc187
z2c3e348807961a1b6882417afb1dda999545627d39da0c2d924bba0868d7d639a2def79f3efbe9
za7fba10662255b8301a6952cd444feee3de6fdecc98269c8cf4150ceaf600fc71d3376b565e580
z606cc3ebfdd01bd384f49028ce54a5cd39577f9ce8264459bca30cc7905102dc8ee50c23756153
z487035fe2413ecd931f99fd90f10ae279c001510145f609c4c41a20632c6f45e20624114c1b760
zfb932d325fe414667cd9cc12820aea95003cff76e42246d2904ef173d50d77efe891c3c4edb1d9
z91f2ec766fb22fc15ddcbde218e9bf0ffa14cef008d312344bd78cd60d45c764adac177032be8c
z08ae07aebfbe356e709df51481e9729d4297f8f64682e96889788daeba9211f3402e0fefb18005
zb1ff47c2680c94b8f504cc3c68925bdbaf6832bcd02b0d78bab5d989840ee6431eb02fdcc77b83
z0adbad4b8a89b25efc40947c5ac9a661d5bd0de2a9ff2b3c30a8101765ad59c3c9f2fdd462a997
z9703d087775c2f66b5f97fed7e0427baf04990fe03c6dae594563e24a61227dd4ea1c34205fd13
zd228df9121c3459580c982cf060c10d8b1964ed0fa52cbbbcf384bde16ba1688ef9a1363cd6c9d
z144528117fc73f418050f70ab598327edd95037546db122f50120f2103773fb010e9ca4a3c0bd3
zdde732ba2288de30a96130659f9f8f3d881d3ce51bf9d8670baf2edb79ee2f22c46d00a99694af
zd6f542403745748ab7bc82dc1ed7d393b580b95dfcc46c2e028584db8c3b2dc418884789b3021c
ze16b111570e8d4613e854d3e1c3821ae77857c5eed9ed4786afdc07a7cc82b4be8510930eb49fb
z30190b2e2f32591e6e2e26ab909043a9a7dd559dd296aa36a96aaa95bba9d16b5d42ebbf0f38c1
z19d881fe4cb367b067b35f0335abbfa856ab5ee70442907e7e0c165f28995a542fcf840d09ee60
z55986803a055034e7a358f34a3264c2a12240b9567bfd6be1c16db6048278444cea7e50797b41b
z18198a4e86d6b4f1466f901d0c480f066df054532d0f0a6fad4a50008b2aa2651ddb9673d52514
zec07c92f4f7c9246466950e364944d9a9ccc074598da00e48ebe67dc6dd1284a19d6f8ceddb424
za539df96bf31a1f94771dae4a619076dd17fb9e22d9f38494bb877569d717c32e3af16527cfc67
zfe3320e2478c003a9d5ecad39355c2414bd42d30435a615c6c213e68aa5d0131f1c109fad841b8
za56693f666c2d2037dcf1ce02e06790f1088479bf436176766448be95f27609b3b3fc49c2659cb
zac078291526b372e5306bf82fb5bb1c4aac0010f66e443ccd69c42d4c22e6feebc4882d5eb9d23
zeed1fdd3928f1b8073380742e413aa2f1bdd6a010c1da5e7395c6f992e61931aa9dfd399f52b16
zf579033f2b3c990776567f40307388bfdf63e4ce3903a7433d7c1b28dee814c2705c364eabb89c
z207a74400f800aa936e79b279edcccaa9aec47b5ad9ebf6a117c412496a1613c66c829e12731f0
z27e2ebc2c0d3d11bf6ef7e8108ed4cbb26d69f0749f73a0c648927a63e53fcd4501a42a95fd294
z34da9ff9c8d6e6141f66785ce486028fcedcf871c5513f5048f7d14697ef14623ea69e42b97606
zb74c5ff0c35eb948f1eee8b485273a98be5744d0209b6674f14e26736f7d2d6fc8a88acbe2bb44
z313f134d017f7a9b3d6fb6981d0ce3d63396bbd54a3acaecacc74114a10db3c51b96e62d1d3ec9
z1402f7899ab09aabc24ba99cf467c0b0847178bc5965d5f3e6d6139716f6d14fe3dcc28a202591
z52ee8389fba137b22d113d1cb788797fc285d4d7c3f251f202fb218eed3138cdd8795feb4b0ca1
z1eb03d5abf99968592c5db4b01436c0a86d7e663f909c68320e755cf0dcd087f472a3bc5b34278
zd62b2e9bdda808151881b9488304f52f2e476739f99c6120b37d9a0c4177b9d362fa632ca61b12
z0471153da8e7741a9b9da602450a17a0d2612d37e1460b3b0b854597b6e59c0d785085a3d003f6
z27f1058e823e45b4398422544d986aa40b3f9ba19e452b1db2a65c15e7c1d31db4d2b8f72dac29
z5431a0f77de7135bc7f9ed5d764495986c1d618c06a956d3443c2ef2ba9cbb2c64642537ebdd1d
z2a5d1d1e85391500d51a5e0b7fa559cff3002ec79cd24b644b198a6b0cae7e7a92d51e9d6014ae
z37341d25b4e46041c4479a5cf5b39dba3b53f718269c252c8c4f7aeef5455acc2f2ca019af1b51
z594edc8d3a84cbfdf1e62dce202349846cafc92b632f8c73ec476d0368db81b4b51ba7adbba8cd
z0922b6eec9f70eb7549faf87d06da9dc2cacf87a9a5f7e819c755597eedf028f00b6e2f21f94db
zad886a71e51cba82a96ad5d13a2a13d384d967a469e2aca9e397efb98a76045d5824fdad917176
z59b710593ecb3dc03bad38ac313c2e035c97394111c8a26469df3d9d8f734a3d8e454f2fda55b7
z267ac0d62a02669c76456c820a1c2453914c65e152551e080eafa162b7d41611f1ef0b864e42ba
z67e955fb0823cf13b64e5fe3ed506b38ac8afad6acb60930ff8c8d8b4947e459faa980bec3acc9
zce17dde179d5cbbfa3a82f6f86b96f44a567c698d85c97ae1cdcde850f7d443d55203feee9c261
zf6ebf3b7b466787929da041d9be2634eeeaa9251217445623ec97685c12fcbbadcd6019c48c238
zb5e976a06a9e5ffdf86c46ab860314681582bcaf7655c638b6549d3042d0fdf476d36dd64edeb5
zc8cb9dc8810260dd8d20607e0381e46eebdd0ccc39ec7dfb45d60aef9d427c26e022abf8353e09
z2c90770d4510b80789039bbfd52ccd5fb78b697097556ca46437f0450cce42690269c56c0609bb
zc2cf01fcf252de7c89ca1a5ce5c92934fb2ce818af9d9368326451ea35baad20fa146d49b722b8
z231674685236a40a6d38e9a79d95e01da80211a34498a68f258b68f491d239698b1cf8eb630bad
zadac47f98581c9f6aadae5d08f1f20f64e61060b43d3c6fe42345f903a9fb884d2fe2239fc12e7
z7ffd5a7285375fa721aad3b3dee066d0305625edf582e313ab27bd5c1e6de2b9bf29a6e3f4df26
z6c45512311db2ec652fe92b49be659f1d12d61610e4e047622cda117de4856f25f89dac74a931d
zb110569a7139f9e486a4f1acfe6f72c10ab47f8da770cfd6518d92838f46a47227777f8fb70a48
zeef34c975d7e35e47b8fe9baec489c135e22c07218b2993c39e3068cb13e928dd345e96114a1aa
z290262ed880997ead02ceac7d17ade542b3a4a9bb45abc14351194dff8ee41523fd7767e2c2167
z6c41a6af7533e72c1e7e598d4cf98d4db799ef530ee4080bd922d2716753a6f8ed642c81151b6f
zd749b37c102bc62cafff0eb505364ec5e5143f3d2640a84aac0e9866f467df01ca68b858d65a4b
z4fdb133d2f35df070d22b6a6029c864c5757e56a48464f017d598ac4484cc87e976f641b3ca587
z1cff03566caf05bb59c353891aa62564b579d2c6f9cc64e629acd5c1f042098a611eaffd99c423
z4e96621696ec0fdf7afe26b62d8353ac233af6c7fdbc02fab58990dfefb8e02595313f86618f87
z2e4d70bfa187c946a0942467aeb236a5aed2a0802291f04e815daa41540b78c517a5a2e9934036
z6b2cefa8192f1f7d31d5db19dde6f4f374393bb020b3559c494e3f577e92de20e828159e0d3eaf
z571acfca9808b5485d7649194efd2c1b0dd60d4925aa407ed58d2264936627a12946f760268258
zb445800c7b0cd3e31bc451111247226594a422eaa8615f6ebdf60f01f8c9a1ddf0ef77e0b57747
z4963aa362366133e82aba55edb97bb833f72fc3a9057d04812d41b4d096ba1f4ee62768ed5befd
z6b5a227519f3203001fbf88678f912081a6fdef78b1df3cd8d7f907e536115156a003433f6d36d
z89d9c25a36099c5c985985d6ea56d5e71e614381cb9c4f736267a608bdc0f29f09f0266141aa8e
z3d1dc4fa8d944d5ab16ae495160054bb083b145e04bb8efb6de1a3bd690c76bc507e32247760f5
z39209993fb97eb45e1483e802a4bdc850761c1f8930155e2da935512a399834de19213c6073712
zb326d3970eb96df773e62f0be2c55cbe333d9a732dad1d68da3e9e9b59ffc078e965e42dfcdc2a
z2f089acf2abcdcf2a9c30d569783541f9ec8a83372557525b520c2f88d7a85c51d498f93c25709
z50a87f0e824f589ba7bd33f0faff3d6c930fc8097b2c3686db45e925aaec2a8627e198f19f92aa
z07d1c2c9c203d7394cb451cbafb3710a0911a6400542cdc0b892871740bc33e2188b704a954ddc
zcdaac026201ba3920cc6f38741240a2b3acf40bfa7d6d787036339e68df11a49b412efc0c934d5
z5f71711a74db146ce36136968454d87d2b13a70fc9948cee02ed9b77993818cc245be5eef39d14
zdb6f3694ef9856787dd2d9b17ad06eb3760094d26f115f8e6619fed60ee70db7c2245be1aefe33
zb5f4969288bf2c7d9ac6a25f5cafb6349c1e66afd82da356457aaf14aedd01071e5dc909cd2055
z55fbe5737a739d471a47efce745eb46eb3416bdc7b94c8c56aefe571cac5d6b220aa087c3509e9
zba8c4c23abaad36137c2c928667a4be45132f5ab881590c95e137582b793cd56d3475729f76cc3
z873b8337f9e1e4f204f5efa0333664f8c80d2c4471138204c8535fc036030f05c71ab66a048b87
zf41275dc73dbde037583b52ec79cec15846e2f6e329ed9aab963f30eea9af06a7daeedc5272b08
z107124114832bce6e5183f99bc9e71a874687b4474f2bf221750f01a0304add787a238b5908826
z2e94f2edf368953634a435a725ea202a90e035a639aa8f35bc33cae8ef5603b2f8e26cc745e90a
z4820138bc60cd1218c8c507e42b84c1e32e1f9292636de6e1b0dbacf69debb264f422ec917fa6f
zf7794ac7b8b5d977ce45587247864dd4735e653f6c58dea8c6f06dbeb406c2f2f76cb949c45197
zc8740237050c17e0a5fe093f1969efc409514f32163fc800a922f5ca3764d98a205b88a1718ccf
z1df7a0cd1521a462d6032686976274cf0b73a14c11578f62d2a5dc5530708b93e2c671ebf5fd41
zc5644461d1cd0ae3c665c99721950680d7c546f51d9e954ca9165a39f71caf6fb7cfb46c896242
z58705faa21876e641a48ead431d58a4b0900a7a75b04f6b594f29a37e7b2badd5aaa965dfd802b
z3ac722ee1af8f3968f8db85272236c86809ba96ad4b991451be14a3948b8fed63216f9b3c5b09c
z3eb789731867672d6b775161f2b148a48b16ff4f9d35934141e9c62264e75e2bd0efe5bc2dfd44
zf6ea919b849d2c530bbfd09e4e59765822c7791231a8f5a16eda80304d3826bc4ca384b1f44074
z8158db722b24fa71e2627ced47566e65959eaf6b252dfd9f84c7ebe165e4f1bd949b5e77f983f1
z4d366f27ee484c8dc3e61a8bbf91b819a7989f14a401e6283a9d5286edd7280d9502ddf35dff74
zbff66134d3958c6daaea0eb2ff2b894adaabd0dd3841f194e5b48a43f6f598e95c8240e20d871f
z9ad16f7435828c1751efcc91e53525147bba82816cb6b1b0f9d1f826ed64f36707f202476ea5aa
z1c9ddee21eba91a98ce9e706868d396e27af3f6d78623565a58e7e60d84a7a730af5fa41b46063
z3f8d71e19e1c641b3d23eef1ee6dd2b863bb77299b61a0db10204a24fb4dd348088192ed626b4f
z196f7d6feee72084edc8dc9249f756d729d9237154542fc1d94adb647eaead3dc3baeb695ce47a
z8c377bea4427f0ba09047966dfc6be1204092109102d96ac7825ee24d3c7a74dba5a570b6aedc1
z56b2de4e7be4159c44ab7b1794d7c53787d830ce8c785e7ed63e7cded2f0bb4d7a1b5ed6e79813
z963d34b1bce2dbfe6533109179fde0645874f0b5057f05a65f7d5695d0e36c92ace87180eba09e
z63bc62180cf7f43bab7023cd292ba2585bc61749a1b388488f9887a7d28a5555f547629243bf5d
zf1a3083ff3cebc4804cfdd4f8cc3620059d10ddf6205df67d082cd48541e67a9ea7c8a1a768b78
zec910c63eb6f933241a120ff8032ea19c6c620a965ee69fbd68b2f9794d00cbbec66691d188cb4
z4c58cacb2e1b9aa262a434091a9aba433ccb2046246c99e57d835ad54420014defb6a033c88ec9
z67338c3176d702a847dc1ec6586d95701aa8ad3c19503e080ae8fa9dee4a99109c5f4f4382224b
za2124b776a880afa345918053aeffb3fc29525411f81fa26d04a23be2d99a826c6350d782b8488
zb8e9a8e89167681c91347aae45b70dd2db63041b7efd5508fda04a9230e4a1a01749c69f02da9d
z8fba91bea4fca8d18473e7c4d3e4a7229b34153ea4e7a73a9c2758439614b9ed9b824d45543482
z17b164b96ab61899c2b8bc9530911433657085a8d4d6e6f2661109f0a99cd22f066db170c6e212
z7296a1fb45113c12c9eac7a9d1dc6d4feddb72ad88044970fe2d901d3d9dbe123d91b32268a356
z3ec77de825d1e973f044c942d8c08d0e3f193c56a13c7dfa86c2d3682bc05a516d7876e0e97269
z026ce50a523ab7cd965563a1ca1a71476910c553483a66001d2e3ea6a4b2f8c81349be6d996bf5
z9850f9a4860f50ba3c8ebd8b3f8ad5ca882dd90488c87736bd5ff9e55a6d2e983fe519c85162dd
zdf6aab0c37798a1f5b937faef0e3ea82a25f89c79433cd80af8824e28973e92069fd093c05daef
z4aa02e44d50fba9fd36238289e4940563054420e98ce65d3de2667f5cf815fc3e4a29b0a46bfb3
z44821511da8eb368a2ee93f9310ced0685d73aba4a1cdeb2f1d2071b4e8226ca715602a4a3b631
zd998f8f2d0f59ef893d04202daf3ad69d59ad13571823f040850b18065a9e047bd98ef790d94bc
z332f39bcf8196c9c4e9bf089fe48249ecc8a0c1cac18ea785a69aa003f8b4c89be14d8493a5ea0
z87215391ca189ea081d932b39b0635f349ed01be70377db40c87a2fdce591c4aabb745ae22699c
z7b35b95a2c49c4b8bee415aed62281d229f799ef88f0119b0e7a186cd346b1a9543dcc82d45f26
z39a2c9da22a95953300161f37c5eef00d9af6eedb505c9a0858daf49e517dd9f83b0c39d8924f1
z74a4577595b3557e3afceb10250af6acf2991dbfe3dc0b8160d41398f525cd20a282dd90cef8d5
za2fc337f2a4a41ea30e794b65a737b60b5d861019538db673524f91cc796cc0ec76139ee8af2a3
zd8e0f02c18bf10fe9d62742bb7d72c46a0f57dd10f4c4feba7d3b3a27e34536fb45d305bbce2dc
z56d943e9d67e15e6567239a334a527f92c09ecf399fc8fbb51603348ee41945e2790850372c299
z1ae9bef4072b4ebfd3c890fbeaa680cf467d2b00930b202f433020c378625ee760b370dfe396f5
zb4132836dc5b64810b27b37ace326c21448990c55f212e6bcbfd68f4bb3a0face2cf23133e2045
z1361da9d7994869f46cc6809a952fafb4fb85069d3f68c353db387685803f64c4195c05d4b731a
z256fc99b649d31670c5edc87521c0abad1a3f6ea2c8bd721d3c242d49df6c8eb25e8cc69c1d688
za0fc6cdec0a32b3a4b3f4359a95eaae595d8dfc0e6d20b0796f0267bc2903cb4db1bd3b1c9292a
za5d0270f6397952f4fedab0d0b795dce876b2c4a553bdb9442a1d68ecc527cf2cfe615a6748aa9
zd6fe20a940a5c85aff9e0c90aac1ef742b76b702eb3e0bd8316e66df2df22fba95b885fa2fc423
zc34298d5b32710cfc8edb9cc278df779473ee2cbd4d23781658a6d2073290692bbda866cc82287
zd5ae06e6d1e1975a887c9f96df47bb0dd0b1aa998d5c47afc06154c03e3d6cb3b92c5301320108
zaba2bec6a62ced9daacb95494cf1f00b991662979d8de2af655c751782d183ff99d937ae2fa821
z1db3f22a3937bf2b400155dc92b88064c0863fe7275d77773a0a82d76db39ce169a171f0d5d041
z017fd1dd15e42e9e026f56154465929db6829e8e142aa06c776eb5719b5d023aac4462997a62fc
zbb9511fdbe8e69f4b62a6d263b077a18ae0c373f9bcda7bc971b0902d15e8f554743c657cc7739
z583e5bd63695490ad09dd082a3850c00516fbbfc047ec9caf686e50eeff49b0853edd46c3bcef2
z54a2e91dbc01f1139e7906c84f2bc2b952ebe21a23d3c2104d5b499dc0b7fe809862f1f55119d6
z42eb57710cd0b1aa0887b549eec8c0713d0579f2ec4a016dec46bde41412656d662ad97493ebc9
z30cb468ece2134f05e0cb1ec5b5ccca350f36f5af6e1613c183d20388777dc4a523ed40204ff0a
z5efc10d4c0cb3e74a190c37bb6df9ba473e1fba240e9641568d70150ac287bd484bddb3a1089b9
z9953629e2ab4c8d101e35a1f7c45533e2606163a63cb8d8e2f4dc229ce8fde21c8d26b19b09d75
z461285038d72c77cab878b19bf4de4c0a41a56dfff04e1669b26a6729ceaeb4598a59b50c6d05d
z866a6fa33741f5560df9f99354ac9300255782a8b81915c7f02c635d15b8ebad6ea6b29161760f
zbd5733c49e62c020e1b2020e19d0b0f134d20483bb170e47d6c2facc891d29ed448099fd948c5a
zfbdfb6f521f35b5723fe18ecf9840d6277e3d14b96a66fc63b2cf43c892d1bf81579235d1fbefe
zc1470fa1030072275b53f05dc06f0425c8f4f5a03e1b9e07861fef3c08cb71ac65c696da0a0991
z8f2cec0bdc3bf887b65ce3b9cf7815f0c47388e067af3d0c5c087ac6d8d98ca3cdc87022e8cc09
z27246667678884abd6e468e0195e267051ee1840851889363d3eb24ae19424d7922445a92b2dfb
z630096273461e8e7b47cbb7b00930dba0d2100350cbb49a053c75c2ce44786ef9f5e7150f3d175
z63df831bd1b9b2832c6f712a385f6400985b97e8930872b68738339d1e268ae0217f07ca1ecfcd
z79977628c8b8acf5daa05fe77c07c97acdf095c7e39f252ec3f8946bad1cd3d7b72160c133ae8b
z33fa83f6fa99a783a72bea86eca5bc88c4438bfe43a9293ab09dcf551ea914b6f5b821c877c745
z18f6233876b3938eaafd847a446445ff4c53a202db132a70a761b1407b5a6830d2db70e8a43bae
zf0d3d9e597e057eaa7a07f92eb3a3953f7ef8c49ce9e3d98ea0a62e066c6171a04dc147e4ae61d
z3497e2bdb196721c30feca33d6ef1516bf938b4acc0b6375354ea5b15324f2d06fea44edfc4fb0
z9779e0a8919cebf335c86232925317e75197b865a98ee0cd78ad2d0d2b5f9b923fb07d5df30d48
z2832aaff0a5d33897997de33dcb459cd5cdc1d01daae67f3c51d6290c9244a4dfc2cf94b6a87d7
z66d42f03c26543e7de19914b19aa674532e97ad189c1986ace5e1744009369eef3dfb685b681df
z31c1daca9d58e241f58e37111bc5580ed8673a08749f42c27615e525513924ec942bebec74fe01
z06812576421ee9aa56e52ecc395c58d8a780a8845727076b714b607b0efd6185d9c5a4ed8fc23d
z83621ddee646a0be562f857b91849d6c5a56bcef03aca7138add78cc67ed29402dab6981b80419
z2fafc2b87595bd9ed736bb0339076eac159a5a847faf8fcc38f7097763084caa7af3e116ad2840
z52c26d184d78b87690e3832eae6c0728e2550f865d7ac7a36abd167818b7dc49e9489853dcc548
zdd54dcf3906150e695c61620fe4a60e97e90c19901a347678935bab5605698a7f06043b53fd8d0
zce886030522b6c6c6b45b54dacb6a62d535828d3351e5dcdafd107653625c1f47b517870c5a6c6
zbca5efa4101a97d0767b07e81727c480d7737de8a279d0946625392054491e7f4f99cc62f7f955
za9a32bce634d1ca960cbbff72f5a8414371d022638cd1918f46f391e2533368807cbf6aa2e43a8
zbebe6c5d871222a2eea70e5b0348049a21b0545e347c46874a913b1db86c583526bc3b5d084c46
z60d67fe309310c971a45431735f5a947171926dfdccd5ff8d7f68eb3ed94abffdd74703d7527ca
z9f70e880ec8b277ce43e1821e65696ddb6a46c7cdb3d135873d28f2c308c39fdeaa962595aaf0b
z9f06733bb1c6d2b327bbfa3b1a6532d8944d9890f85ef0f559b50d35b8968b118868ab420d777c
z053d2caaf3c4f495e2d895b96118fcdd364d4b80ef885701bc193e975281d2926e3abc559614d1
zaa5d0ebde5ff5fb58bffe5d02b9d43fc6d3e86c99eee2698f5c3cfd0401602441a62a01f380ccf
z04db9578342dfff0a1b3ad27580e32ea51c52cab8054f2b8f8ed3a96dac5f7c23165ea52257019
z4cfca88eb12f69e6eef7534483adf8a4e21ae5410c52cb25f91afaac4fd48f19d6dcb0dc151146
zc8425f2ea06b7fccd559304f9af1b6d5766ae70d71fc4202fe31e21012bca6f2f738f1b79d828d
z261d7edb79698c8cdd941ad6f094395ffcc79db92125190c7c29d95296749eab9635295aadf1b4
z7103e5083cd6f1f91dc5cfc1819151421d61aea08f98dd1ac4f675191336ba6c2271e8ab96b6fb
z9e7c6c047d268cce5ae6f5f75005ad21f1f722556fba40d3ac2d0ed9508cb69d22ca94936bde35
z25e3202b671c6d1ffbac4fde0759dab7a2980a3f2e3ecc38aeb36fee20cf692d71db0459774a0c
zfbea6b216e9148537ad85b4bae60eafc166cffbce90039ce749f738c242684db958ca60cddd302
zb56fd68642815c346a814c848b2cf1c54d5b82f8d615d6d738f3142c28fbec66460f31fcc2cf5d
z59db1b079e6e38c29ad16c53e38a411c28d0bafc92e1fddce6d2a0fff233b4fbad6c14ee0fa932
z30c5554c3e7c8bce2031db921d2334b40fd6c10e23f51d845d910958c94ddfea260a6ef37138a0
z63fbd37fc2a6f85565fe2f26046a5ee8efe1cee61951c54caad04ea350354bde2a33bdbb95e514
z7051713cb0ba2e4b9a4458359c313995a155144d97e2b56f5870c1dae79ec93588a61afd0fdc05
z3c682cfdb13db5160d37502cea66c60fa6cad000cfd30e437e416ce536b4998ddb4df4c93de3da
z3180c4a79b9ab0d4137010973ac8c421c77a24a695d69405e52868ba18fc53544ca56329cb4fd6
z65708a19ef2be1fd9599fa0e1aba5271670897cf362b68db43ccd5142c1aa7a64b83093fb0f239
z56c125976547efe91dea80dc9d4bc49865a612ec906b24853d017cc5e69ac4f98654e745064ac8
ze98ad5a6fff3bf983a6db3609efefaed1ce5a4146734f264d4fb0b0e05b76dd7ec271ab2ee8447
z0213dd89ffe154572b4c223d955b30ccb3923909782ada4c34a4bc5fc599e6932764b1c70ef793
ze6d7c64de24668576d147af17191f78b071506e25e8215d7c56fc23c40a6c075157222659741fc
z9675af88fcf488a538371997817a28972ed052e560e8cb681dca7d55aedd03c5b7bd0b2e7e4812
z33c0a1d4d110ad9ee7e080914f8a7f36706aec5c89de901e4b7db423ba199e133aa8e4025bd17b
z464a54c096712acc46e2b7ee06f8e3634c67e39c021d5d5998580ddbfa6e16af864f33e826e2ca
zcd58ef8d300bac14fefb27e737e39d022cf3dbe933abc6d95f128b4ad16580d3ee0ed5600a5bd8
zcb28a159a9480276897c581bffacc79193f87400aa4af4c8754fe0d40574c9c116e1c05de2802d
z22473b2a074693b5d5b959edb7b6d2d1676424f70c9858f96f43a7b21898fe4f81f006bd5a1d8f
z7d5bae3200e87e463106b9b5f00fbae42f2117fab08624e35fbea3374fcfa6df85c3452b1cd0bf
zbfa43a4090badada9492f179297d4e69ff09e95309e691436695362f5e70e365c046172f177a34
zdf95d0ade7dda356f4f6c86b7aae122e49d0aeb1d839756bd1e76f80b4637f12793b2acde2b488
z6a9aa8d7989ff07eb9e5d65705c8df14f24f41badd6bb798260aff603af63711ec8679229e7dda
zdfbc3555df9fff0d78203e8510b25aa2f6b5c97252a340e87e3664ad97e157a8d931e38b85a6f4
za52275ee846a07713a807a89e81a10ca948103e186c2126e1056598f5863eab79dd87ef7c6e3eb
z7f2218c9711a68bfe51feb64ad64dc26c39677ba6ad6d211ec78e09797aae7d870eaf2a2475481
zbd7d0806651ba7188988ec3f3b1b6134d6cc99bc6c9c45021cadf44541911f271cf815c3be4a43
z36a04b709d997ff5cb7ccfcb299e54f0563fc026d831fec0153a70b993f9abdf158bce614383d1
z842604fcc387647583ddeabee0667366469ed3705fa389603e6be6c6dd07a97cb21b20bd3b1388
z366fe6bd04d341fafc0725e1ad10dd917fb3fc3511dc48e4df206771f711a2aa29f1825f828233
zef6c9829ccd91c830c157e041095ed7d6f1f1bde7ee869e864d0296b8dff557ced43cdd74ad086
zd851dfbe1b23a9a301252cb083496e609c62005ee53accbf42a8315e1c35670027376044833893
zecca6b542de6406c1fc12f2103859fd14a808fcf36f15202a6c1d9edd3dbab52cd6045c26ff6ea
z7794f1024e611b14fc2d62b347da5dacc411c59e63e52eea41b7e816b69aec54c0ebe0cd772ae9
z4dba5f0e99b53c9506f8dca62527824478ad25d9b483e9642553052f43dbe89f61dc72a7fc2b2c
z47437da1ae61258faa9b70f1ad2e00c8bca583cb8be53c18349fae03af8a3cc573d62c34eafbf4
z71b3e052cd5241123aaac9dbaa46cbd4f65eefe2c35b3e3db3189c3267b58ec6472a45ab51f490
z1c2ffa0dce84773f694dcac163539f255616865815d8b28c55954fd9c1749f2ea36086938c6241
z672dfcff670c026372d9100572499115610624a83af066501165fd74921a30a9d292b114b2f132
z56eb51a3c1248e5d0b104b86802c0d1a2064cf762c043d41dfa25cd1d0c5d03db2c05aed60b68a
zb6b4f9c6c1009081d75d39ef1cbdb724c13045d270c7ca64f1940d90cdc6f121f095ebe5d558c4
z449fa3c6d99e6e94d44083bc9924c9644d23bf4519f672d07f6f4cc0cb5907e1c3d0eaa3cac721
z4889dee0550c9745ad3ed988470cfb7e8249b527afbe18bc4dc0d19c5ca05bbb271df3d1f94fca
z95b556851dc7d71006def748da42f5dea94b474039c0b7206eef1d6d2e57598f1590d2802c57fa
z01d6091ad93a425bbddfd34c3e81cae9038493cb3f8cad6bee5c272401f490489cfab306fe1b90
z17c919a60ec825728f20b0d6d8764ad7107dd1feed14773b69eaa0b54f4efe13c44bc5c33c45b7
zacd6c06a818836059cae022d8179eaede666ba7ae54e4cd80bb2f61929fd5fcfe5c8b1c1dcb064
z23acb9822fc805d6a335054babb003746887c85baa6ec182430ed23adcdadc40e290d84e41bb16
z88d1813e2716fc34ff92e91730a2adb0ee220157568c8c0df39622aaa368b2f4bc4806eb3d6464
z393e9c9616f2c0b19be3a00837201f0103a06d81d08eaca8f267f59e2761a926b12b0fc3dd11f6
zda7eb739d99e6ee2571e9490d8eb52a5fb117298753f70915e98a8f5c9c346328f1a2851983be5
z0071dafadbd674d7a89002532f777d6907f27318fbe0b5ea2480c93b940e27992f4d2e5fd559e4
z901c56185d708e2bb0e13297eb3ce3632197dc7729160534f157437c6d115ac0d6557ddcc0ef2c
z834275009bbc3f1e9aa4235a00d83dc03cb6168143ddf8ca210c27ef211692dac98b41da165b7c
z0b1873ca95ad5ac26f975b94d1efbd9c3ba1d12b9ed8c94caef168bfb2e8d9047d88fcc164ae2d
z5c22b50229546d2246603e412afbddd6cc27b513a183c294c858a07066968111773cbfcc389f1a
z70754a50609537e3ba355729026cd03363d5c1cb195a6a75554d628fe5a4b7ce56cccee22f00fd
zfb21f1b2af4054c682e957d5d35c2c3ea89924e59bfffeec7024b92fd8ab06c422937c73313266
zea08cefb23b2b3b5f9ff3adb324955b7a3b151fd643779749493609bd3d96b46ae2d2d5b54bd84
z188bc80b6b288928958d21051449fbf4458fc21dd9d0b192b5370831e589b94271754395664270
z223c7175727a74fab6df1f757c2dd05a3fe8be6722d1c0c8364ed72ec0e5186450fce588c8e443
z2003c953a8a169ba67a6a4b499f6f99914b9ade685fde9dcf1ca826744162142b4d240c62ba2d0
z368ca1cfc9d287f9137d1a2398f81cee9d299feba0487e62b689f5227a8351ea6c70d2e23a87b6
z9d7be0db02ae8933a0522090aaa3843e5c730be3807869fd853dbf2aed26a2a51c4fa8d3ee05f2
zc658a3d343bbdb7ea687948fb6382fb014b96ac65623fe3be19188dd7afc33b897089d2d8043eb
z32cfd3e142f075e103db930db098312c4e9f9b6d5a7a108b73764ab446ba674a2e433d269284e4
zd56fce232494f0a8fd9ca220a0438b3b382d69c74bea9fe54e6b76106529d63cf2c73735d9a711
z6394cddc7c2d71e541ec691417bf1796c72f8f9ebad00f7e6489486b0dfa5e3344ffc9cf422bf2
z9e8d2e5cf96dc53652b97d62a8e086d6f93e4428375df9d84d488bf161a2f59c1eb20adf774931
z39fb6cd7e489d7f628f01f9a3de3360dda62dfc6c8412a5d3b4b25743a0a6f24ccbc3316e45fce
zf3611a5584e4e47d8b8209c3baf0c25424cea41a5e8077df4db95b59cd0ae9305dc0c2c50c6d86
z51b714e618c5112cc376eab4a012a44d97a85c25359ebf4352d5968c1ec33591367dc8ef6b2ded
zbdb7afc68eb1d3e91ba4580416aa6089c3bfbd6f830af3fc49d6513e03246b548f6aa58f246aa1
z62f1bf13ddd7afa80a1231b5d7c90c769051bc5a1035617d2f22430b8b62418d219a37e0f65900
zfa16c6707f70608e4b75e112914ff460ddd78a2b9707f7c2726b5c98bcc8ffa2afe2507bf5aea0
z5383f9b4ab781bb25359faa6f753f778c340f5fbebaf87a760d8d86856a19f52eb2a7d55afb436
z4ed65e2ea3350a1c20156f2f909d9d98e9c941bed872bb047c1253b67295431463f65690b07870
zef7ee08c0410901954cf14638a7c88f57362670be122beb43f82356bb7ba1542e1b8a4b0cfbdfc
z6f71ff8d80032ff2b0f29bbf6a1cfe21dc152e0f799069570642d2425556ff1801c94c69ad192b
zb85e1885ab2672171bb61b2d02c685fae870e9367860e15d816387bd2cd5ce902785bad7b686ee
zcccc9070c0938241e9d5111fcd9c1a1704550a8c56d65762fe0f80236893dce7b20aa76b0814dc
z7b33c0ef56b2465df906cdd56e07176d9a9bde22e00fb9a2410fbb0d93448a52e8b48f06ba84f0
z4175c5c878e0d8eb89978d73f91afd6185c7c330401d7e6ab97bce621b1eea85c765a5a6280a41
z811ad4fc7b037c96dda00681798cb4b44f604527bbd7fd0dd999762ceb0eca08f2270e2dcef950
za9082cfaab2e918bbe13aaed969effea5fa0ead0f68ba8698d3bbc0d2624732fc75ba106e00617
z67b9c23b3a58d24b422ef7fe61eb42284205714a2c80088442dc53555d7b202000b229a7f62921
z29949eccc274c7c4ebed76888bb13d8d39331d5f8e14d47f0179c682928ef323e8ca88cdf3f9e6
za629e17c7ffa390c8a7ff9d1d1de4ec387b6e69426c799770f1bca5a3643400ac213fe004120e0
z4acaef05f2878d7bb3e1f7114a26646e59bf6325c9a967d76ce1eeb2534184fac863e3e8352a8b
z77a2a555b7610cc6f3c3c19fda21184fac87dc899ba776ef12fa16838bdf950397c88b1a2af373
zed2f46f5235c5b651cc265f3249bccd769b84a435322e8b7888e0153856a33fbf82635cef0bfd8
z9edc06f70bd983fb11f5afe4ba3bee9b6cf8bf5e2a695986608c1888f2acbf96c6698e73cf0b3d
z33cfe292cbb4a8e607fe8496392d7c5b97354fc37e43d710e28457ad1d7201c446bec1644e7cdc
zab15d2cecc6d29cc163354a051416a1cd54b205e4b1dc516d4585f2790622c753178c6e583368b
zb60c990fe8ea2b149390be7e78bf3f7f95966b5fdd2a8fec2b6d69b3b4ac8a60d2b13fe08fb3bf
zcef7a335e2688fc12c6eeffc433cb147f6e45642bfacc615a3268d70f7e2967ce6f6264447edd7
z032fce1a7cde43b021fea706b1653181b72c3968527bbd6911bb54d6b227ca3b6b1966922887d6
z217991aa5cab61a4bfc4d3505438244c90622a9901ea8f79d64fc07c3d9077b3a80d3d8b917d13
zc14192f909df3ed88a9d1364729cfcb67551796fe8a092021a449fe21abf74f76607c91f8e8873
ze026263047279d04a8bb4043478d42fa1ae95b2963df2b783cbe4797ab928a18591b0a6c51f1b2
z9aa7d1476566d3b0d56830c290920a204ea0990f4c8ff57877b466c68b882a4cf7877dcdaa32a9
zc20234d103f8b92800fe3fe838368209b06799f0846478551eefdc3a59d4b01bc9f1b5aa28ad7a
zfd6a89cf7934e69585aaf4091688cf7cc47acdd25f9cf2dfef5e4faacb3deb05f28de39ba441c2
zd3e83a2a87568bbc75ba66c3b0eff675ae7066e732c9852ccd0707605ec4048602938ebc086a36
zdae2c57e13673ddd37748ad47f185034143048bfcd60f92c3aa3e83cacb6b83a510d35ea685dfc
z0fabd364e90c4f083a166797c948ac223eeb8f99dee39dcb3b46604ffcbcf77b3e98efb0ebbcf0
z97a0e51b8f404efae1bdc9b75ef1b59365d3085d196e5c0bec0fcd2b052b0d07b231cb39274aaf
z7cf398d9b9b5e20d2e91244d7dd68be61ffd7429431880e24d71a29f6c7d9656c50aa7d5d29ef4
z3afdc1a4504c5dc4b025c8ae203bb4aa58ee5ca821bdad08e1323414c85f6590129599507f03c4
zc9c7b2c0fac732bdc50f31e070cc00e24f1fa4cbe38001dca8fb415dfc9d9841c8828bf2fe410c
ze3428726f421aa891efca5b4b9942b25868c4b842c8cda4150ca20c978c8219353695a1da73bf7
zc960dadbc6a7765df42ccdd92dd952d09260de43db2eaa53235981b038ec96eced158bf1421e74
zcd408492676769978ee0e84747b570b0484ea9677ec013d236962da4311b765c9ad7aeddcfdb3a
z71cbc8faddda0a14cc3d6babb05ac8333c693112c625ad07808845632ce2f85b0838ecabb239f1
z66d693ba02d7c5a4a12325753a5cbe80f1bcd48b2b8b4e2d5350d53f528b4595051a95d3506861
z706c232e941fc9db04a5e5b5b0d682fd465d9130496964c570befeb4c9e9b0f007b744057439ca
zfff76fca14ae38c290e94a11b26b498aa546a8007f2f498cd8e202c46c8d483603fb3605edd2f1
z70d080589f147f3e471e2d5df802679cb1225492114f539e74b22aaf9d7c4803b5d64f9d65aee0
zc03419c55dd9953183b55f60bc99ffad38270549a271c60add330c583a75c70b232a5a8a1cc44c
z27e2cf6f60406c567796cc73a4e52d7c9d0f47706d55f06fa15cd21e068ea05b1adbcfb1c680b9
z79403306bae6fb51580df750608873aa3283ca0f2bd2f23520778e2b8051aa5f787f2de76550e5
z59cadc163fe52f5bffd09dd4bede7ccab9f24f557082bdf9a67f7d7ddc0727b82baac1562ff7c7
z21d0b45ae3afe95d8f07fe09ca25e2558d95b9f841429500c814efc01ad85fd1253570b08e0a70
z652be1a271ea8c91df5b62f98ff86a1c8aef8e22011ff2223213ac145dd2b026d8fb2e0189c436
z4fc66b8bb2271975bfa53b6795547cefff252b56b76b1c4bdcbc1b05fa3eba64d699f98a03a5ae
zbb849b84a1505e72e5429818722619e1ef0dafd01d5a664775c260b60241461fcadc9147a459b0
z5e20266264cf72cd1e137d44643fc95533655d61a6e328459689aa8d70b3b7f0e1d71eceb299f3
z15f4920c3f37361c43ec65edd19bf64e266913dccd661dbccff76ff38994d17b2500e719d23b0f
z9bf2cdee2fdd7afabc07d24f1f9d8ea4b9f9439df4cac009088af01c6080d5eb1ba63571d05f19
zbac6e9c7007df663e08af6d5eae3ee4400940305a70280148b3facb2460b820dca781b5d4dfb94
z790578b70f74ce95ceb77a4a1bdcf078d0237caf28a311a4bc9b9db30b9baf3eb66878e399ba36
zb86671880b09aa1cdf15cc8d56c434a273dff553891a4362754413d174f962996978c99f69a922
z2c76e26c70e2bdd55b631c696d6a14117b67f51d5780181e6633b66e55f9bf2a34408eac364d65
z59e9fdcfb9292b78683d52713403bacf5bd8ef9e7e0decfd60229f80081cd53bf4a73fc9de3ccc
zb21f68068f6737a3a4908e2b90fefb4b5bf49eea478c36d386ee2076c0ba8b4cfdc38775a7e495
z13b18b5a0becf9ed0a3d74df5d9109f76ab41bd96fe79a9a4d22d71b18a60285428932bd7eee13
zb90d54c16f10f0697bdfaed084650e29b5394ee2f2f600ff101ae1066fdb7c8aafa555fb98af35
zefe277c1d52648e31d9482761f7eda6d607c32c88f50d80763cd5e8f1e77b96679caceda514912
zf6fa646c5032fca8f083ebd950112661560d4d4bca10d7a1dcc2728e0e5ff84b5b1405ac2eecfa
zb98d9da827e79e165c5dbd48f2d5ca197db2344f3744f301ee422caf6155038a977d53b019fdb9
z4d757b592413fe065cd3f584a7ba62ca073a0e036a7142470e36fbdcb38625ac57d1f6d49ff892
zb4344bfb8f93b0accbd7289f7bc67fe2ef34f9b0f3d0664bae8694f1a282ae15ca526969cb6418
zcbf879168be68f3a03fa3f0b37ce0519f8e33809f0e8ef610b6fbee3bcaa7b22ebe3c7481805b6
zb9bfc42651f847c6a79f268330214be44d35fa1864844418f28bd8bbe2fa3b2eada93fb9ca4160
z1ae8e88738f605ab4ba3ccfffde31e456c41ed6fa099ebb0111e8128f469c2ff1303af6c3063e8
z5963f8dd33b4875c543397f888b9b64518b3dbf59179201357e2ca7bebb543ddee16f2bcc0341a
z0a65d21a7bf0d9e8d9acec8e3a83645a065c954845328f917639ba0c9249346417589e0b03e9c8
zdd991bbfdedba5a374a3f1999890536f50b2cb2ec7a92f9dc41612c679d4e74f9d506b9d5b38c7
z0e25814622b1259262905721ee9298c4126b4fa01383eb34d58566b0e1acd3253857c2f31fe135
z0aca6c856acfe380e513478e7922de92ba0eca97abf461bc10d166e3f77cce669082d15b14d48d
zd4a9b7378eac7c270004d67ead53f2852d03b070b0d7a2638038974ebef72f746638540920314f
z77c3ef0b7530c144be16fa6c27894185f5fb4d21acd054bbb5387265df10100e1e03d74fdfab90
zfea394c74acd0cac8b8e439f31533697c6a476afff7f3049886edfbdaf49a705c247584fd2368e
z95858dc6f07e5a40a489eb7a85edcee2d69138482073360bc4bab08cb247792bfde3320a962bd5
zbca4b4b314e50b504d36e762f9e94249d7031b3cd45228ff93a9e5d7250929dc9953a82283bda5
z9254d2adeca959a2d7dd7e95512abc990afda1004a25912094291bd8b2585925ac4dfd12713f92
zd4d6dcc7c1c9f3fa0db649069b00eeb7747d7a397c9389dfe7c889749826d15536efb867df15f8
z73c7c363690750d933fc73099f6f468f656afce7db4153e2c9245dbf04c7be4b1c5820a84b9690
zd4d0b27a96ce662607ae637e70e3bf8fab2abc492a28c8664056195ff80178695be58c1ac30774
z44e1cf2c1f6b1bea33c03af17a2f814c6847e5d88a0551c07999ea0b7700289da63ceb88956f5b
z491726e28205ed3ddc31c9bd40a88eee84f52fac4581532c913039493fea722450011b7d7c9a5f
zfd8a5ce0dcf6f828a0509d203ec333eaf6e2a2708ae12d4b5d40a5cf57d72322f521fe6cf919e4
z5a08aaa5ddf807b9efbb1a2ca60ffb5e050e1079028b25e9558e1bc2b51ef8ed0cf5e696f057be
z2f54df75e70db1f4c4d8f4a0809bd23846bf4a1fa1906e42084f859ca8858ec0def1e3f5f00fe3
za762a6aaa93ada76b4456dd5bfae428755a750424e8eeb6e1b8c6202895ea435ce806590ef16f6
z39d8f4c65215364d8a538cd56c022f0fd30b6ec3cdf50ea02c07c9fde9d71b57a91fbac21809dd
ze4d11c226cd815ad34e6c1b139fb22a2000e7604ec6215490597e4c26e5d29176ace01683ad311
ze584dc759af1c3dac09cfa25accf6acf35905f7347730b2de1bc4ca35b45cc0961edd937fcf148
z95cc9a290569d2f81b27425d2a382197c79991b9070f1f6542e681a9b4ee1de8ab97a9235c6cd1
z55c5ac151fef61f3e59865cfe38ba821e7e7615d8a5448e73653b31f27684fddd43806a30721e1
z3c09057707bd907d3d756da5a4ee82c48600e7dc69db71fc6e557868415c97c68ae99f31cd86b7
za3c43593cea07902f4568849d75a277bd274ac10abc45e87c97a0a4c34dfbfb55cbeca04e1902a
z76eb7c429297b62421c7f806053b9e5c3311dfe5852ce44aaeb38a7c4cf33f05836f4286588cf0
ze97515420351a040d9d0a254d06be6bd29c22e9ec7175ebb7e43ccb6360e38fb1ef22b8acc00e4
z4ad5b3613755e7c1c280711f470eed36a3f52634805d3cb9b42c8b1015a7fe4fdcc03da80e57e3
z7d5d8fda5fe0ce93bbfdedd0cd165f63a392dd0c12eec711b921e7a8f8c8affb3955c49f772168
z28f3db309cf697c6b29156111c9c1d0e977b98bd3c213b528a91f04c1df7eab399ba68b4c6f017
zbd54dc405a7708fbb44fbd59d3b691f2abdd64b292baa8832be10fbde039d7af1c68b90b7e171f
z4e3dab3092d9dbb217c94745128f520c6e95399f07fbe8f1cf68dea1d2bbbe01f3c31c9a92a678
z78736a4083a43866f671cbf63473f0c1ed6ef8d1d74bd87ebc2949c3d2a60202ab438f5b61b8e2
zd025fc34690b1af4e442e2ff038768d2e9bd943cc74d0e0ee06549f3bc55ccd96626afb25e0e68
z61ee0fb1e5d2764f70ab6dfff7810af8bad271bbfe4c81b3c3ff73b5cbeb71a4e66c347793e4b4
zeb0191c1adc2ebf3a6665d8126b39236b06c350329a2902a815ea0d8ecf3acb9edef2d5e982761
z86f2d1d14480993d34de29f2ac5397e2f7f8a00df6a6cf0a008ddc1de643822322814740a87208
zadf9c9a408dfa5dcb321025bbe0e83b3d7b145e4c0c7719a5eac677fb518fe4b965812843ca3e7
zd79141fda0398a5ab048ccba27095079ee50b67d10b540be852db39b3de3ea589966775c5264b6
zcae90d86e7a868b3107e313d17d9de506d39808e0514a6cdda0c6d326797b85af5715925ae7ab4
zdf79eb1a97055142e76b877763b667fc5d8d4b80f424e041d63c6de61f2c2851e97a680b265642
z7728a6929e7539d1df7d00298c44adf6f709e9c26f6066c06583199eca995c2e663e5d78e6777d
z8c4c4ea2eba6ed7c44a98585b788dc061340141dc4691e10c065a66034cadc1b6b40bfb6151264
zc39708e0a6b1993eca81944c4e00df0a8c8fbd4c70faf6008177ed1e344878d09e200325140bed
zd0c77af89d0d7be4f78bd8f933eb9f42652861bfcea54ca9923790ccea05784baf9903fb29c1d4
z503491739d0df997f4ab7073d0ba9816d1c109acdaa1da391035a03ac2eb00a0d4ee64c7cc15ee
zafdaaefb5efaf25c8376b07c7cd1217b3be63c8a79bee0f60b671fa0ea8b39f6fbc137bad77cab
z950086e202614f7e6ffe1df8da44b2e2bc2a29f50b13ad74bbdc51e9bb3facb874b09e43aa34fd
z55dda786400dcff8e6b71fe77c1bf1b7b4092ec7445cb98d824ca820174f8476f4eb2bee2bfbd5
z7b91f79cb0561b94eaa79d15516c0fd934e17b7fc4c442fc02730b6b7d9d98c96e48a6804d0b6b
z7b1d973cb8ec590e3e7cad82e4faca510442cce2130fcbf58a8d1fb8766916b484ee5b4c61c73e
z7ea43bd1e83ad47495e7d4f69582bd6491f24089788e72b88c7658dc83a635d058d01cae0c88cc
z1626ccbf5528d2184a748ca903287a639fd3e1e89ed3243b0de0d4107e1eead07f9fe361b500a3
z4a75f86ac29c1bed9d452854ae8017f264b5625e54186a14a9ea77b5898b8fbac1fa573255d7e4
z0c998367c0e32ee812c95247d9420eddbf439bfe6caa9683694869eb0faa7fc099ce4d2cc3b312
zca8c79037f3f7d5cf7203f163047088c50009f9bcee65b843670e81227e06254a9afa9d9ebc873
z65d83f78a92453135dc510b5ffdb875fcede274cf86f1350946a8970ca798bca4fce0cbd5805c9
z3f82fcf9db1ab57b9ac36a3b280216727443817613d7fe5136f57dfa31216e66a284180aa70b44
z2be8af79c768b3ac96f1d70c4aceec6e9c50960b822cc850290788b7c3eb4238b867a28a1e9a9b
z755cc7081e9dec4034582176da6229d01d83785dcd9867a71a0eafff0564c5879b656283f670c7
z3be5ece90ac682c21e39d71e4e7b586372a6f1deff38f5330c183903abf809ade057eab1740230
zde659f04559689f000a13abe846802fb25fdfab30020418465b287591417399e2b7d7a7a04f646
z2d28cf0cf9748087ce22315a1409b9538ca05a6de3be28b44b6a3214fbd0d6afbb1ef7d8a2d88f
zbe2ec99f601fe639736ae2ceafc3b073bce7543ae7cfca44af78357fbc767752b0e965e103c404
z427b5d0ef9ad7c26745cc0b7593c0ed78a147dce4121048c51cb8d3d96f530687c2da1024162a6
z25b672f1627dd72840f56f7eba674f0c492470f41d11b704a2ebca9b88d0a9a70e25629496164d
ze67dcceffa2b3636d0075c723938735cac9c19c41c2a5d9e54a16ba4d95d46f84ba0f225301c13
zc976e3679fcf2d119f938b4cc3d24f6a67d84ce34dce511869fc800c7c2a043e4dc536a15aa032
zd97996564d8c238069a5068fca8eaeb5091686736466a3d45b87e2978a1cef91e65c6e320ab0f4
zd60dd1a45941d1acfeb8af1c1a6f70b9c51b07efbd01a3670dbb02ed2c1fd3d21fd25d53870dde
z80bc4d24fb3d8343a245a19d7ca62ed79cdf8188f29bf59ae0477f3a07c60c4044ae87c5725d20
zf5d12d6637c4eb818f3af6c55e6ee220e641b44e21650e44ba5fda04e5b748addbbff2c8fc1e4f
zc908b1476b1fc4497532b87a1db087c06e036016c960604aeb5ff5ec4427a2acd0db0a7a1799d9
zaa497baee3a12abc0735e55c970abe8d25ca3f4923c4a5f24017d572f946cbf9f1dd47cf155c99
z9610c12e3d21ea17a2a904645ed5aef08bd29f47c10ba9570bcf4ea0f8a51dd68406df34b0a244
z90d90ef20404ea95cd5dcb24da4f7ad787ca995396914af0ae75fce5b0ce438931c55308bfa03f
z28eb8aa8bfdcae31c6671c87c6788222bec8e3fe68ea3301626bec8d9d594d305527f12e261787
zd0e84ea3976fe41e89c15840be6e3aeebe1b1a458ecdde2ac9e5fdaa55933a22d0427d8d068ae7
z26b1872d9e85cdc0d2b58cb1967ee9d27b975cc3d5c5528e33a5416fbfe7f35dd4f97cb264757e
z73ee45b3ce9c623850648641fccf5a2908c2c6e889c833603c667f157d1dfa433f930308311ade
z73e9cc577bc79c721d04e72fd9d9405a4777b8f9dd7cf18069fe291bd6327b3d20d121bb9e986b
z9cdadcde30e5e7c3e1c64f8dba3ea8f7fc2a5b7ca0f6a61c44aa0d09e178bfb2b61d90b03dc3eb
z7f4ac25d754756043a396b1e140b6f1855805b985a4d5061c2b61241722a632cc750991b5d9ec8
z0d20a151e984a979b364b83f2e16f38317f52c6d46bf6c251fc4189084b0cac674d4a556863b03
z510ec2654c486652443ab1c8dabd4aef45e16e307b010d1d3d2aaf0885e44e917c927cf5a0ab66
z0164fd12651ef6112bff6dfe6367df9e1a7ff9ed992119a1cf1d79ad8af971905cfc1c6d2c1357
zc3a88b35bd351be9c03935edc950faee4bdd34bf17b2e08a6d7709343f49309647c0c4263626fa
z9c343a616371c50e4e54a88148a658f1cabeb57b866e5a5c05821ba82d4b14914f098ac39fa4cd
zf129b7778945de083a492a8f9ac3e730841f95d0c4ecd8ebb3375d644c8b2f2db39a1ed008e3fc
zaa9a366e5cb45e237cffb484793f4948381732d51570b6d70a477081b2ada38cfeeaf4fe1c0564
zd3e9d17d5966ab28ae58e225373a4ff5a7785d25ef0993ad5a485d5e9eda360d8d736bb4f7ae07
zc6f3a317f7a86f39d2295f6432b62be9a12ffa0e0e8bbd02804340c83a54be6e1f7ae3d088042d
zd45f2a7b92296159ed08f17131d27d3e62c9505ba6ae42f7d8ab65d199cee6453c1329232c75af
zeeb4d293a9c8cda7e5e6a6f6d02d97f76fcb753bfd63a2dd11119ed7b83c41d5726a2d34372e08
zb72d45c6eec72ca71b729f48e665a171672488d6c891ab1c795c9bdb96bdb2ba9fef58d23969b5
z70f602ec5a40385436378f2355372e436161c70cc3e39ea93b9f7751c67a4183661bbe3abfc88d
z738e33ebb56dad69051d5747bdce5541a1e4c86c3f996c74f29ac68101358c14e57a1085bf4191
z42be1c37b69c79e72d8c141bdccabfc327c51acd22e83a8b9ec60d423654fe2e2f825e4406aa65
zf9cd52dd975010b34873ac663f8ac26ed62b9d48f7ab13b1a126f12bc88977fb95c264673b5cae
zcb061e40c17f65ef6b5874375e8f51ba169e45a86afa9936383b13db259af9abaee3c88c3ce93f
z986f384d6ed86424506e8b384bb04fa49ae362478d9324cb361d29443673bc80e9d750e404982d
z8d539c3b9c011d75499f4f76fc6e6c61b8fae6b0ae6e6db1566a95567d96ab7520ff84bfca4607
zafd5b67573f38c4f542c2fa63a7d7181f9597886c025ae969789ddaf869499d1dd68726e7660fe
z8580c2f89fcc982d70592eec615a62bc2fec72e36e6c992645198ff1bbdfc639676ba199c22c0f
z2131b02936f05c89a507ba65f567aeca01539b0c2157a8d9eb237b7804c86f237f20024f100b10
zf801c611d4b99a6bef540cc9c6cfe25ba1f7878f5ef3f3b458516c162cf4824b6d18a6cc453814
z20fb47f39e34d0a9c324f2a3d35122b599ec50c07606ca90e2be681aa2a63e9e321070c5bac183
z39039beb030717b51e2476631e11071c78541e498e9b829a28309df0c3461f84a4b5d3196595ae
z36c5af6f46a63a00b7e9bc0c80d3da34625be15c2fc678205f8abfb3fe70b87442098545cff108
zeafeeb7cbc9fbf253c090c28f3784c7745c5aa89a5a5d4579a61203d4a3b516e913a7f9891aafd
z3fdc795507d9de4194d3cf8a68a87462abfc546df57f46cf8d1e86f9ce09bbf26cd03fc5dd9a6c
z4be801dafb4e51e663980b8be5544e3311adc4a66a53968abf8710301242eec227f204491d6095
z96bb6e07a305cd0dca19a47dcd0ff7d7240ced9c43ea9d8187474d9865be537ef9c8b103cb9ac2
zd04155cd49bdf513a3dd8cc8f8f35bfaa47150feed34bd09791dc7015d6569c8bd1ad543204110
z6177d6654dad213e73007f361c1d356781baef5fa99b75b0c989ea46cac020b2e89ea353864370
z63a359dbcf83c4039415aea797b5704f2a04bcadbadfa3d1ed57d86c0e9ba38659d1801d3df3ef
z6aeb685d3f465f4cf94ac0eaf75622224ec870553d88a1ae9cc7f0678aa06b7bf642afe43bbb05
z5a493bbdd332b2788a9b74b809b6b0e29babb3b604aa35c3bb6d686426a0edd8216aa88c674257
za568aec910b8828e1d9b34ea390eb63d4d9a2c2b211b7af08386111626013b73ef6f3085009a36
zcc39b97eb7f0ddbd1a624d36dbc8c30a2d0866c285a0e2469b98c1131a38c81c5b5f2c791c1377
z1668500efe12829a80f608f98154d22bf707b86da5a3355ed6f2d3a9b0ffe53cd23be1d0f214c6
z7dc0c2c45c3a810a25a9598bfa207717b909ce7f90b710a2ee6a54729657113eece298bf0cc6f7
z211274afc548738842175c963d2b45895e667e0d4f2010bec7084519c5e025176172bb3239ce31
z22be6bdc3bc75c27c693244fe9fec3bd6deac8657aa4d87b57687651f314ad01dd741638fbd743
z46be700844d1c32c6794f69d4b8e6f73ad59c3e464f151638736a7e461e9396114701d0d1466d2
z8048a3618414138825cd69cd94ba9c51260eb97383904adcf169fa5928fdc15a846c540585abff
z4ed4d47a5bbe2c62ed35bf7b7df8a33e3e9d6b6ee06864ac6162ce63f52012b5cf8c6d79e1aefc
z1660b5f61e38ff0611def60791861a9a76d174e0e76e8d7100fb1a2a0c69b17bc06131565fdfb9
z445436282f40bac8ae0f4bad71ada428f509da3ed663b83a960e40a9bc9a4c151b0bfe75c61bd3
z14586552b9b68e673b69aefec13d042a6b2edad03e06fceab05b917f037443ed2396b571bb2bd9
z3756fb733c951a7f27066ca4dba97a3e703bbadf6f476938eee0c90ff66935ad5a27b2481dc8a2
z09b2b892929151360e7d5bb8f042f319d15fade11389c8c99e84056bd2bc815ad846e119a8d6c4
z57b612a6881675feb960f2c80858fc0a5b31fdf2dd224a898f37c9095af00219df18efb1c08114
z4c0c3972e9fdf06df6924cf97a7bdf57a16b2740f326821bf6cb07fac6f96571de6a3d488deb89
zd183e7a7225d9b6b365390d2742bcc606522bae4390fbe2a2903200f28db49ed76a3a1a31e4bdc
z8fdb30ef1fb9346a3b92bcf78563019d830511070926b1ee828c9220d7a1caa00114283d9b38b6
z684667a6693ab888a5f4042347eacf091365c2d132520e65651c6566fc07ad23ed991277512d43
z9a4872feaf7a869e176df89ef714d7504aa49165b778de87de0d830d07e3435cf88d1e659df7ad
z6b7e12543ce138f7093ae12f5cf5d000b478711fdab3bd548b0cd90d9fec9c30a5f8684ac36a31
z59253b0e99576c101c78e650230f9b900dc30a656be723fba7e711e231ff2745ad09b167f3484d
zfb574290fdcb78e397bcbc08685a2309ce61385fd5e8b60e420cefcbcf26757ec2a3ef800d214b
zbce7e5b3664f13bb9ddd160035893da81b687d3f2808c30ba67c1dc911ae285ed0bbced009fb50
ze55fd695f7cee6123cbb0054c2472de7f70281cdcb701d6355e542bafd5478eac7b0d5171c1e2b
z02d762db10f81e467a390551aaabb6a12a89c5ed49f1f751193039058d4e069644b829553ff923
zcdb102036c72e2dcab15c300d57a91f21cb742770f99f35fda4a8060875bd2df0ac28c141c721a
zda85b4975fe977ac6f4e223d4ea492c12a6088b49fdf30574e8a316cdb9f0d458c2a7154671039
z76d52aae23da853ed5852b9d21d4490a55882e92a5eafb58aac2a56fe9304e30aa177e10f60a00
z7187e70fec3949b4b99f0abe8b587553d14be23155afa7544d99c16a31da20f9f26a8a7d531b36
ze93b780f2487170e142d282070fc2e2d204a86d8713c0fc51e8ff69877300521d76ca0fd232445
zfc5b6b5a2683008251f5d41460e7b1f7b65dc89394a26d3bec93a8179ee3c992b419190df470a6
zc147a577b1b088febb8f676688bab422ca011431ea1338a2081c7c6cf8c412cedd1a738f6f265f
z6fcc59970477e317fded2b184af70753c8ccd704cebd8fb100f094905b5eac04a37a958b778ad3
zc29e9fdc29a99c30a1dc8959c7879a115d73855d19e6468c074596c076ac9bb77331145de2c879
z22001681270aab9e8167d12008486102eeccc3533b962992580abbef47baf92be856daef7ec8eb
zcffa69909dc9c0f9a8df039e7dd73219e0c2194a8277f42ab7e48c3371c547cbc695d1947de9f8
zca3de4726813c1aad5b78f1d25d7eacd5bc93cd376f1963327805c9fe8e845c76f632e6194c371
z2e05c612cd13887332a77eccfdd9989528639286a95eb0d9a7a0c493fc4fd197bc20f109aca30e
zfb1b5dfba879cd1076c23180abbb0332dab5243cc44606af66cca84062412d14729383c468cb03
za34d94b038cea466549be22585b36f1937d08d5cebd5b7125e84c69c10fdd0eff51dd2c2cbc146
z4bfa77859045fa256f8fae7aa3c944964d30dbfbd4e18c32b469d7cb7ab6d8cd1fe18944367b7f
zc2bbc6e8851bc679abf229908aa096fc25a66aa38175cb96e73e2d8e8edd243097b0d76fb9f7f0
zba2c309c3a47478d62522e814bfc88f28b0a7d0709b23a260caf93ef00e9d49844d43a764eafb2
z691e256f197926988ea6e0c9f26a8afee913508343424ad529a41d2528af619844aaba527aae67
zc1c99cb03cbb3bba43a4e68688f0e13ba969b703119b7fb6e39e6a690b85a23f1134d5b4e817ee
z57bee95d375c3b3bdf7272b2de63e587da6024b541f5c3fcdc972bfed1844adb755543ee9a3058
z54f8dad31046c6d08b791fcd63a9127b8b5cf41eecee0a7b2e37326f6ffb75f883ec454e768aa9
zf41fc73492fef023280c8a8bb113992b9643ae743c10e2a0fbf35d5f0b0d4d6b8a5f8e99af3aab
z19fae134a0687497cb018a75e95956e449f34a614944cc65028a3ab7cd3872760a3f9ef1b04d38
zf07d2af1e96468194259c19b4697cf760480a7dfbb308904e2120612bf244725bb0c500d0e472a
z6eab11a9e78679c5a48c744191cc9f1e84879bf628522d5980a5a324d3bb72a37dc5225ce7041f
z39b17df8027f292d4543c912c293aa2478755c0cc317954d0498f51de916a14ea3b698cc7906e8
z479d65e065219cb15bf0fd1dc330db1e5130838a7a57f673d07fdf229734376bda4869d736b13c
z74cf208e473c0fcf20aa6c2a39ba68b261d76826fded0f8b543917a8b50d3aec1f03640c8d8c1a
z70ebf98043f037969998910edc5bc65acc840724d5678df46e3768a5e22723dd5cf20b6400c367
z69c3a52a6e8a613b34301c8cdcb5463e9a483ae1f44c2e35be70a6b6cb143b166f25783e7d568e
zcf062e1d3162d6cf049e76239ef96fb71cdf778151a22a8dc364bc6f1f7e4f18bdadd19eae60ac
z5c92ee0747eac1846566f85d3d441a8e3af4ffc92e0721d20db0b59bcceb662dc3640af72f6f5f
z295180c5e21614a80af539d9e22f41ceb7c1b1db45c126f8648e4bc96ee669a1a83305cdccd44c
z797376ec91bf66385713742ddc03ccdf7a41b66424f5b2ccedda288f4484813cd0d2e9ec28ab7c
z1f2c571f4afc1354449fca18a5d103e2c2c5c2e241d47b456e82b0e274acb0c9480d28157774ff
zded94db62dd4afb8b7a0cb9a8d7e076fbd7fbd8fc23bc44bf68f0cb5596076053f236bec59d75f
z9f82079b1b1e0b3fa998d3494edaba117df77eee2d4d9dbbc4838dedba1bcaee7ecdaed0b9a98b
z0df86a7899e14769e49cd7be737eeca97031ae85558ee5afe559d6a353fd029dc39bbf15ab46e9
z12dfea47412c4b17836e3ddef26a76d4bfd0cd1e4554a73beed99b6c0d8a509768e7c15b4d36be
ze99c03b471ae8867146f9076599aeb3a0a08684d701d6748605cc1a434282d7a46554597ba127e
z54041b25591997e453fc623730cf1b62965e57da40f26d3e28b4544589bec3342b160f356da571
z82c628a76f751fa52d89c3fcccef442a1879ed4cd39fae0ed029b9843fccbacb2f7223eac7bf46
z4980dbab7b223cad958aa5a7b985bad0c5548a6251d1a399bd93a59a996408e91dd7933676300b
z85b4f33d02c25eed9ea8566899ed981004b7188b63f2eca7517f08728ad90780251e0821fbb3b8
zc96372d39aa4c2d28805c9304853c5e84450eb7289ab47f34c7e230323ad19d746fe68f85cc4a5
z221b8b56983088b62c08052259b78f1581b65fb3ac05229586fd71ffda302f353c2c28fe353d81
z02bf12497a6c7408746f174f94f51709450bc6b3463b6eda2a2c0ac3e3e9a850b78fbfe8cfd90f
z8bda6e64bc49b332f972434ddc79fd78746815e876099a7db931ff02bab365aa4f772c146d3328
za35fe94dc3e04cc68044e0a9b0db6f57e0cb4bd46ff7b9ca78dd09659c5a52ed40781ac0dc2e4f
z7e4f2e993741deb3a2718cbe93c3ae5a35740f21587615a5303ccdcceb92a7b2f794db054866c5
ze72f617cea5b0db1bb051939a9bef1fed85fc6343dbe990f4104dc53dfd806d054523aa82fed32
z3bf9e9499f252d9bb2f2db08c091f5166a8dcdeb47ac57cc288bf47eaadb005860f91f68cb2521
z386f6cc6851569b9348c30059adad81b58e8c0ce73a56a6f88707591aaf92d96811e1242456e9b
z017a6dee85f47ab1983a5a640a658360099f116534198d988570da78e308a456436f43c9576a7d
zab6165c5e8556e0e15867f6bf7c4908063b5e72656dc8689c08ebac469bdcb268c6b0b0879ddac
z092be54a3876c138b7d7554a02acad58268675ac5705e91b6a932f63cc3fbbb1f2766064b08688
z16d21a9d32c37d69833465b2010f9a064930508c3fa1e400898798696cee0b7044e3b60c7d4ba9
z1e0aa60f1192e43b37321bc4b40cf33300ea5787b4966450908f01a470485c7d7cad7654d0c2fe
z91b2ce24df912005c9b2fc78210842bae3e33814fbd2e324d1f8ec0bbeb9bfad190d5bab75c8de
zf74572b842c02cbec74c452478751e47483540bb8d44e6e1112f691aea30cebbbe45d2e483f200
z6fe641806ad12f243b8c1bdff71d29cca4a7926f9adeae4e8477ab0e37fdf244fe53ffbb9c2a7c
za73ffc4659fe44c3b79a4792d84d2db51b4135668be26c8d879b7966f75f2baee61b4e36c21c32
zfacda34cb3412deefad25570703bc5a6899438f8461d60b36aac43b904705daaff28d573d7713f
za976e8239f43a24d952ae953e9b97a445d864140f3c180d7667707d42281a2777d4f2fc8c35b68
z4ed1b754927ab1dafc38429fa5ab0cdbf1861210f8788d14a22f0efc350d24b41752dce6b03a55
z639e50ae0beed198d70c53cba88de7a91a700d78ed876c519077359a887dfccb60c7e3df262484
zf8421f670dc02064c6e8d5537a721f05afaaf4a897bdac5dac3e60f85c8d00920e4fba9fea69aa
z24543826bc40f6a28f3eadf52b1e9a0044f5a11545cb08aa76033311bc54225f348851a780a3d9
z1fbbd8bff5709edcada3d075c590e0f90f420ae8e57d9f2cca5be6d7fd467382c2250cf8367113
z8f8bf1f62a123c247f8d5b7ace2f1c87b8f7dec3c2bc8831c39de95bec5f1b9a89ff6b5cbfdc0e
zf72f51c5bfd651ac4254c799e2489691f57fd72d5c99bd1a39dc3f4463b8451b336c474aafa2a3
z44daff95f5d836bcc23d79e675cd041e5e70c1014a28ce1e62a0da6f47aff6436b48b9105e2bb2
z52f1105974e0fa82c39ddb27097e3a9690e917723372741766e74f4e921e6b861a3162071d3536
z5df7736a57a0bb0a6dfb57586b70c77d205ddec9f23437eaa9c64c6d2282e31f5d08
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gigabit_ethernet_64b_66b_decode.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
