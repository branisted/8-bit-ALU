library verilog;
use verilog.vl_types.all;
entity mti_debug is
end mti_debug;
