`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1bc235c2ceff4f6e3b1ebe72fceb7af9adc96a
z694b4bad7241bfbe775016041d7caaa74d9c0e7b507ce89e8b01980415bfa35a8e346f54c548f9
zda8767c02ea87d27eb7a843f4cada7dc3b575fb5cede69da7a4701b2d725c73f1f7375e85a74e2
zdeae70c30f1127407402c955b283d7b9512dbb3cc85aff97f613d57a4efe57b3c092e5ccc5b6dc
zd01018bef01fcb6b6afd138be37349905063433d6fc88423f78d0a5cd8c325dc906237be6d3673
zb87d9fada90e2c892651aecfcd04caae277f299df76d77ce870132e5e40888bd3b3b1b6bc6e799
z48a23782b89d176bd848937c64ea2b6938c5a6c2c52409c3721f00cb676ae49dbce756d647186a
z2d5ecb2321a08bb462a97b513b2f2f7e1913c836666420a662f742f4dd090636a3381f28becec1
z1708d87f1f0a00e76b7fab8e82c4b58a7479b0d3618edbc64d306b42be8b9498e21a252a9f7760
z4ddccf620c22105b64d3442eeae29848475b6321275c60da85fcc15cdfce58c0be67611b4ad217
z85faa32f1a391d7896ecd2d6a476653f33c744e342ca0bee6222cd817d247928bb48ab87008585
zf4c934887ffb02320d1f5e9901371c546d07491c6dc0560188ddf7660969a0521bcf06899960a2
z846b97706440dae0671d4d93134b115147c7d3bfbfec814d2c532f2bc7b5a866f7796e878f79fb
z6352953b57e9db9e47653b1e11547331dc0137729d159986fd727762f733f71a51abb4c40cde6b
z54c31b12df4f712a2c305b789f9c8c8d46984771a07097977cf132585a196985bb181add954404
z36bded7d75961463e3e276ac2e2008c390d0d00fad22ac8caab98e40b05c933281c5564459e8af
z8f9aec18240d5d36f086223b5e95222f73bd924274934a787a3175a67677b85f713dff1bedb855
z960c8dc7ff24d866221fc620d14d288d5566aaefad917b6aa9ba4910366ffdfdbcb49a0161b60d
z71c4abbe05562942e7c4a09a9dff28c943ef7c6c1e6de5057a705620dbfd1899a77a946861a2a3
za5258b51f50b15e1e9d1ba5773de6452b231c03b1e4ee03b38af5571c17b694de542838ca07ceb
zd73b049d682c025de3028ea70149c459fd5fe8c1534fd2073fdb5b708ca80de4fe0c24327d7ebe
ze6f5ac9fe2a7d3915ef17479b49e00d476bdc85cae1e1c7b0b7fc872fcdf985a836855c52c6337
z753d70c0046642b17b1004cef2598fc48dda8dc428fa2961de13495007ee5aa14104e778359466
zed993b1ca5d5d91f1c91a832e66da662129c06cb923667066504505d5a62665d284c9ea33fb58b
z2477a57131bc88465ae49002e3a2077d80fc4ad438a952fb10d7859d6580dadef38473619c0c60
z4488020621dd5dfa9cd73770e2ebb616ba7eba5e8ac434cfff5f7f27dbd9905c1c8b3a661cb1bf
za821c2f3f1afab9aae7f62b759c53f1389a5aa085f88f9283cfe4a10649d4196c851da4320cca0
z09965c93affbf8c487be9f4f854b119204a0dd14feb056de691598efdd65b5bd2cc86cd23bf668
z4c888bf8c824a326528b7191d2be28381c6739ee127eddfa50dbe45b766205ac45b962c8ece8b7
z54f61dab50d0fe48de3a131de077275ede28e65654a11a62c7dcb8d18860e6213dbc6d0ad07552
z0275cef6917654f5979d02fff9415e2524fbaa98e6d1cd1d28570f1b2fbf7bbd32f7d466cc3f3e
z73d9512d1129816bf29fcbff6e5508795fe6a320e999f74076fa20ebd70ed9d4c602a20f88a40c
z4b5f34a0967bd3d7947fb410b5208f1119234a83009a53c24c55270153fec89789a02c01cac15a
z028014740bc45b836e1a539f21e0ffb50ef4ddf22725ef069cf13344e188c30bde00b3d49c27af
zd2c433327745af3d6389bb9dbc7ab102c46df7439c9d84c107389b85a611b85e0ac43f13f52741
z4ba9d9306141074c2d4fd44e7c0015fd8d1698434796b11e7149eeb10c665cc4b6f42679ff7ec9
z6b6d307da20a2635fa14a368a472b5107ecfc94ebed16d8e9030b241d838d0fb352394c0c7af3c
ze3bc25b4826ff20ed4200bc80a94e1bc339de8d5cc1ef43b7603f20d2ae586890f629c2c049754
z598403c78a069b69dee27298656cc31ff2b34cf867561a2527328e852da739f9bb126276292920
ze3b2e4daab448c369c7ebe0efbbf0b2ed20ca7309a780727f4de9552723680f4f13bd5e2a378ab
zc2b4b5ea11cb48b27cc583d3296d112167103a8859657582566c14b40bb1aa61abbd6a876ecedc
z6a829ecddc9c32ccbecad05361fd8341cd62194f545f80ffd497bcf2b7b857fbf5e1d968998d13
z6ff3d8edd1884763990524453b8822a6240ca26511cab7cb7db719b383c34c510bf28267d723e1
z223de55ba13331686a2bed93c409b1a2122761aae8a35d4735b644b9d1a9954cfa5519d61d83b8
z8908877c098f2575dc59748e185ecf7d395bd29b0b0303b683d7aea441c06e6429fdbca6d47576
z51a18b86f6a8174ca75f4a1a0ea1abb7a7b5937a7073826284b31e5ec933a33598f5e3b3691c2b
z1d6580dd167d3f3c985a2655d3c50542c6b064d87fa1627430face914bf4ad2e8480cee0fa43e7
z2b1db67299ddca31d62d42ed24777810563717533e660a5d2bc8386a43cf025e046f79e09893cf
z267f9bfbe188d88cfaba1e2b843a5ccca4952a6465df2a3be338f234ded9dc8d6533c61fde8d85
z349bc725fbc246484081a493efafbc2e527fad73ded74063cebbc7ca523112d01e7db46a787c6f
z7d9b34f4f8741d11ff03236f526a7fde909336a81d14d38e68b39459cbe85000b42c6c4b543ca3
z5cc7afa1d5353677323078ba6913b0772c8be221733bc79a65998e66be75f1e8681886776eb12b
zc1f62daa4f62545d11f5036701997308f6f31e99d9983368824e6947e7ab68db1c85568c61e305
z70abebdeb7670e49cd495ad6b7f41d2e90c380de471e7822b56984644490dec97bd445fc0d83e2
z03ef9f5f41a4ba4ae8c6b77952e968cc8e7920350579d85cba4d256e275462e7c282666c9886bb
z9ed23b912a018f973f187471976493447b0aadde97f3435cdcfdf68924e98a223cdd5a1c2b8d59
zf246dcb4b08da12a73c53ea7adee2346f908f4eb3b732d67150f7b859a0e656aeb6d428e3d9091
z8e3f406b9a5e9a9e66947bf35008bb49871261404203eb51819ed8b52c077bd914a895a6ebaa84
z7e7a9d9afa0a3307e9b329e33ef393019b0b752316cff4dd67fe4c6bf54f4b5763f5c0618c977f
z1cd309678a0062c51b9d10298a2cbb643ad7500fe20adcab32c2ea3e9f53aadedecf7b477a5505
zb916def6693cb3a3b64c753e24d556e9274ee15f7116feffce533ef5770e499e60bd37ee21ba47
z2810b0d60fcec31bbb3c6b505cb6373d8901497e86185824e09a270be7c4438bdc65fc93afc7dd
zdfb557a5d2ac761da8125c9ad3758613c7362918b81c85373e355746543d0d39739985e216aa93
zab943f311021c8d00f5e2d2607394fc30976b4bb0fbab86db4f5b62fb32ebef49944799a9ba202
z45dface9f0ed3130fc9ddfbb4df9d7ce3e15328284f8f05c2b61f450b2c32f2e960d944150e3c2
z3207a4bf47e1d5f327716a887e750fcecbc282c52f0c075b137b2b140213e1fdb36175ab0046f4
z3351491a3ecaee1ba8c9f5bd2ece0de76825d3e936dbf58d8cc7bfbd76e3d4de0f2b8789be7c9e
zca74b72cc644f9b8761af97d7a6d87095128582e356bd79ae64131365dba7a89f23f4ef80ff80a
za6fa70b1550a84ed206d0e071082b53509572b42cbe5b8c22dd3920c9e3735751ec40b9f58e143
z32c103f742b41801c9a913995b0a6f37d09d144ab6debadcd6b4eeecfc27f0e8fafa62674ea999
za14a69e1b2ec7ea3f1b413f6145ad39be52f320f74db7e9bd9e38bcf2301ffede3bd446af0a32b
z36127381fd16467606c73d31caa1654857f0f88c7082b88c9c6c3208ddfc5468c4065465c2cd46
z7257f422f5b3859379e68ab2a08d0c2e9706e0b5cac896ac2229b51e5fae239662ae3f5a025f2c
z919e2f1b7239ca40adeec19b653a6fc109f66318b4ad7a338e717a42bd70c6d70cd1b33b43928e
z87b25b392e0d68dc3322dc92901c57b2df0ceacc437d96a81d1b735ee4b6fade6fdea1eb07da48
z8b6e9dee5dd1f1629cedbc9e2f84af3fb7a44b2722922e7415ec8738cedb740faaadea904932ce
zaa95e22b2d412608f3dbffa9b7fdccb4e05dc44963388f3aeb725c777b0ae294609e6f1e30dc8f
zf6b65d499aaac5ede92110ae10339c32f80c7ae9cba457a0dad4281997a0142582625095359a29
z4bb9cb8cc05fb2155d52bb2a64182f9fd9af2a1cac7e319e0aed804afab5e35698bea3805f7b07
zec8c656b8265d28c44585280fc868925d831b05eaba34206702b0e89da8e85319253a93d9a9c35
za730f511b3b1cb533c644be45ebf23c4ca3639b7fbefed6ea3a86abbece6d9bf5964484ee45a31
z97b961eb5a7bf550fe90778c3c4c4d93fdd94811b37a309f770c3bd036da190ba91f821ab69e13
zaa25978ba9121bcaaa2f9d3681e9a8f87e8367847948ed79bd03d0d88cd2fab915a8d38771adf4
zc21dc6fec43a62e5fc42970537934b414bd7a1d8a93da3ec732ace6bdccce8fc659833abccf26b
zba1ad0efc7ef1be07a8da6d13140bdcdc603c2e87ab7d4a92b2c0df7264a323c76fc2e345cf382
z9cc8babdd50f2d9350aa83502ffba9c4e10fdfebd3e3821a4233dd6a409f7b4d9c5dfc07c5493a
zc602070a445c0781faea4477dffeccd2f5bf50c71a683a7c31e593c15dcc0969e1c9a89585893e
z3c8eef6bd6fef84c29dbb3bfd2a67870f8e3dcdb147c460140e77de6be69a1a4cf1f01bee85507
z23547a19e4eef0a9500fa7ffde6c41dd100b80d90c1a9ca40604a4fdb068c17198c5cd62934ee1
z76e9de550c726ef2a97f18e51c87e2017209c711ab335a8cac46deb4fc03fcf84dfad54f80e516
z988e90974615c6c3d2be759bc1d0b2ef6956411e0afc868a4fbee5ffa5de7ef9b3efdd86ef328f
z310911578ec5bd0b7a3c9aa6e868386fe0213380642c9a697cae082199b142549c480c34f9933a
za2169d6bfc4a9d87844abe95ddfb53776ea7c66281e36844f0a9a189867326de92922de2bfd424
za9097b43865ac7ec377d33f7a8281238734d26f627e9d5ad2f30e3ff74676e54a6cb94e2357736
zecf941df0be823b53027e16f3722ccf9595b6eb3904d8254a702bcd91057492392d43c981ab66d
zc990a320e9e2b31b849f3548265aa24bbfafcfd7664bd79af18c294dfa0516c63d579de28259fc
z8485bf17a095ae6b3f30a64b731e8955a498123bfc1006e4fa22f2c5f6d5c74386b49259b0b5fe
zbbccaa40c4becf8865deecc2e6c66ab72f535dd4e32c3b7349fa8105ef68e80045e9fad4734184
z0ba84e7ab229c56a2bbda829cfb9347fee6632c216cc955d55095ec23345ca30284bc32be76e0f
z862f0ad8879dc00a9e18004deddb4c801384d57c5802c45a780050061a5bf01961531f51670db0
zcc92ad8de2095c875eef424c1ece59b0c79095900791730942d57b13b4d89afd5d6bd7fa6e5bba
zd32554ab0f797362c78a4dc52f2845ac6b0999a3b4446c46048e8a3f2d2686492b0f4d3f7acda1
zf5191c927b797f17cc517dfcab3d8865ce9888925aa204c355411870f4c517ee7da1d67c4412ae
z6a869cac74cd4423f529f4140c4ef244b2b024cb2495d0666dc06cc893fe9b33aae56127cc92fa
zef70bedbf6924653c394ccaa7e6df99a86ec9bee54c7f59d37099ae11fa1c0aac233d3a9cf1f44
z2941b2eca3ba290f548b2e567f2e91497ef3d6b580b7c1a49098c1cb31578df03d6b1f0fd21b3a
zb647d203196c2b271dcb8365d8ba626850ddae0c08120d38b43b1d536aef66058b29cb9cdb41e7
z8f791b4fff261d63a7f4b32c193330193673231151ee79c8e42b7e8e838a19030d583299d583f4
zdb29a989b6bf1fae2d2222268695e2a74a4e27c58c43f47f2ae831c4e9fb55c0171ffc051ee278
zd1f1410ec6e580b0a71b6f14cddaf1b3830867bdc09c541a196aefa98242e35bfc13cbab075c2d
z480e7fcd24759692078bbd2a5c7d723d81f6c437905d5389c3b5ac3e70c4d39a22451b4ff7055d
zfa8305b376eb51b6caf5e58c4f62be7e116398389d9a5630381a56c9b7294da5fe8dc69d3d5baa
zeb8a07bcb819bad75f1b72d0b8604776668d1b357e0089c0d6db2c269bc0e07402e62a06271322
z3e68931003bd2a29578ce84443c458ffa9f86c1106be21265de0e135a1a139fc0d3d304ca500ba
z116c679e1c5955a8359f2f313fb8a730b7c8cbcefb2560326a6392c8bf70deedb03c74ceb48493
z5d5080334725927b7aacaf85de1d5d7d8c8261c48fabaccf32fa4d128b27d4f3e07554f0bdcbd8
zab05d4c8e8faccb463826ff400e567a4fce9cdaf43e2f8a5352825ff4276f5f448672e82c42414
z7253645163d26c7d82e4a0a1e5e47dd59a4cac6b927976202beadd75207d5f1b86c3c92a383f28
zbf931e765fedccf8a1b0c825b483ddab62d3d4462400f04040ba77e6364ad3467d59d42d0ba3ab
z3f197bb997f2c08799fd992042d4269ba57ec9d8521718268c10ea0e2250a4271081b4fd2b1ee4
z14aafd3ca43defbfe213ade759ad6cbed152216ccaf5e72af307da71ecfed13effda66540114d4
z72a8a7c8c011190840e48124ecaef1d99a0ce2164aa90eed1bc8652761bdaa2b4e94dd607f97d9
zd40c9aedb5b603f36784a1d1fd3cb1e187e860d7f24fa6295083cb96edc60fb3fade523f243b8e
zc2970d3ea88ba0a726126134a77aa93c77427585572a0c3068c26603494810482c97610bd8ba45
zc79233418d82999474431a3073cd0c5f0332997b8ee6d85f13a35ed53f3af81743ac490959fa8e
zb97157952e402c03d61ecce7dbdc3801fc19500e93ac204cdb40381f987fde66a0027e69c8c6ac
z054f70219f37ef54d0e2d2342d7d2bc4590488eef6399bdaee3b4c1fbde43199f3682ea7cffc7e
z740983ce683c8ca474316d0027127d63f7535ff83c784e08c3a124bd6171ff89096bcceaf33be8
z95f3c860f41082dd90dd658f9565d88081f895692636051e9e2b7f2630f2beeafa62a0b5ce78d9
zeb9e273fd22b1d05a218ba3bf6029f238d94055c0d7c4553c30d8ab40ac4711657160b8f5f441c
zb532bbf7ea6293100e8010dd66d4f0e9648e17011bd415eb16019542e5dc3bf64bc31db7ae2f7b
z62dc76360a7be51d86015d98082da2dbcbe681625706ef2ad3a82b82f6e2dcf994415948c2948f
z29a29fc9ab5e12b938aa9af0f0a54955b58020af786bbe2ee9b1b3027e92ac512899dba9fd821b
ze30570268e23e8e92da2704989c9a25164f51e9fea9682eb7269814dac30fb084366576d28b62a
z6d6fe1a040582a58459138f9c8942a39b4dc5d35f9a95acf464e99af099813090977a7e523dc86
z70849a642dea35863a30ff531d70369933c23ae796c766e6bbc4e7f5fbc49a3211e59efb828a52
z75dac95ef9d1e218c6ffb11e7abf54a6e8a8faa1cbdc6d6467a8d1f6f9ab0e1315f0e0181b1c4c
z9a7f91922adcaaddd519d49ee491d4bbec8ef7d8436acb33c12db2fc3659ec529c2b7c54a6154e
z0ec74098d47d7d85b2e4440c60bcbd38c20b02ecc3d96258670ddad4cb3bf45bad81092cf1cbdf
z36e99748a5a198f45bd8c874f8ec023a3b440be5d8767c9f04b79e4b592e10b7dcfbc67a27b0ef
ze7ee66873d34d072ccb9471833e7214ab72499e241411de71f6d5721c99dfdf81c04423f4d674f
zaf854498e707ab324d2bacd6ef6381c33cd1f6fc3e4d53e6142d5500709d6848bb5bcacc341e77
ze8ba8887a68261d245cb30955d82a84374d78b01c842c3b67e4455f406b16e19fc19fda328ffd9
zf6a8e22c1ff7d2ba9c46f67614dbb9add087bddddb28c4967d54a203d64a57695cf51ff33f65db
z8d98fccd3cf3c882fa5b8d4fe406a86deb98e3f23b443bed445c314b48e80a2b2fb6cb45732be6
zbcadc42219c11c8be1d387e9646a83daf18be4bda364d7d3297b50e1a09eda9112400f86c07917
z6f46e9fde8987017d7e3f7d8cac97e495a023b0aa53128a59579b3adb2d6b74db2d3e9dcf161ff
z05364660d7c18d625a8d61d1a1dc43c71f094d654cce52e835a3c14145b9599a2c72e3919ad935
z7f750f4941658d42590784f05fcd1880b255cf6b93f18cbba1ccc7e403ed0efbd1a3df20e53cc9
zfa2bdc8543d7459d6e2a716a2e2b03c57a401fdcea247f97161dbf0a54090aa33fb8adf0b89a42
z0b04a8879f7d1fabea1ed6e2e428382d6941d7063b195787a3072f4ebf41a76aaaaf5f7d5b4d53
z3a312132c1ff68005e17ff8dab5fe92a91ead767e81cfb958242aa912fd6251551250becd626b9
ze52a54b2be99783a039ae11b62c6f9aa972d179eb6ead6f0618424a17ca69faf37153e56da88cf
zab4c0f01071b9ce0c32938683341f48ed1d3f7ad534e8e47d8d34f677e1a872d8ba78eda6a49ca
z0963a43088acef7f7c82a7314f56681f9a38149c92a7ae40641dbe4f7a22c005690fdd02183b33
z224ec7b01bcdeb52e1b85b5138be530884fdee164592e5a652064fe23cca34595a3e791ecb0d1e
z1f88b5565aa13c5cafdf156aa26a0504df047ec560462cabb0d87c479f14ca2e2644bcb1d74370
zffe9ae0362ac0406cbdb263eb5c9f6f95023c8ee5d61decb2cf1600767cd8e4a62af22fad238ff
z7a412dbbe2b766459ce36becba60f58d6ade31901a985ed3dc176caaea1c97fb5d1b0a20148f46
zfc46b900a79ce7ee52e441fc480c514f31e2ca40aee2afb001679a9741b6de2e7a0584b4f774a9
zdf899a293daa8cbab8596379285bffb7fef8c0b7789fe5fc9a28edc9533bb7ac36ece8d8dcd27d
z0d60a14f0d8bfd1b5c9c3917c91ff5694ef80d525083c98612799c76b37cb415700d398d417f98
z212e117c167f18e1e3913f0a744256a9c7713ad6cc64c923013057761fc0ee07781fd86b474f58
zfb1faa5aae4d79f9f4b370028863325ea2d50662d8f833fff42de64e5a2eeccfd6dc172c8eb3cc
zb789fa665307e9ed14cc5cc45b6fde4f8ae695d271edd193731c63593d098b1045a98d3971f449
z3c515d380f5245a0b4d7b6409d0437a5f3e14f8a02bcaa794d4c5eec4b1b38d69f893c235ce95d
z5ffa293306bc6ca8e28d21c066411834cc599cc83be7698d8fb747c5a215f08aa1b046bf845452
z3d584087e134abaf7a486c339d340db151d31085ea9b7799e312c2a40ce2a7c9e4e539937fe80f
z4f53c7fa843c60716d842fbba1b1d67633dd94e6a2dc4ce7eaa9d8a358e2ff8f42357463fd1924
z2abaea4882c4dae9aa0e6757a0ac64422af3115aa1be81d2cf00ac8f5ac44047dbb318e63a990b
z3cbd8a46c880457cc7456b17b5aaedda074d92b9f71ad3f811e38c06b819e9fa5ae180e37589a7
za7c63cb4c8a2508f1bc31c987d44da444a47a8ac674883a6fe80a98bd68c4a3a9c56924f6a90d7
z188bf1033a6714eb7b874e1e85146cacdbd434b82274d93e581d461f7c013837091e2ed9b57225
zb92fd42b86d804f4c661bdea12d851e9e176e4223dcc1f024cc7036aa023942ec2c93274379a16
z92feac3856cac0e6fac3939a541464c51bf17722760e2b60ac48cba7e4c3004fd73262140d92ef
z268744441fe17be78d9963e9395ddad81d7d2311b02af23af8c7fa95d9d6dac4356d28ad31fdee
zd47c646a31e077b37842329026644808134eaedb321c24e93186449d1425010366214318a4596a
zc8236a60d9f6f125773fb845e59d15986483c65cf298a7cd10309ad8cd1c31342973de91edf53e
z62e1a64f296f146d8d7391da626616b93297eb73bedebaa396761802223cd6e74c407a0926f00e
z7b72334f2a628f7a73d8d773b9c68167beb11ddcf21071e48dfbff4f4e372730537b1d950fe2ec
z7ef19641fda9893b1faa629a49729b8209d0c14e08b20fb195d6b1b1874776db9ffc37d19f9f98
z68a3c506894701c8ea49411ad304e6b44529888d9772142cb4bf622ee6f0fddf1a4d5a06491580
z0a34a1da123e4e411e70aaa11fd375db163a8b7954aa7dafbda6327756942a951d40ff5a63778d
zbb4994f5a290a0b261c6192d27fb5ebb4c8b062ca91731ec286c0171f0c43b9185cfef8b48867f
z03671b76a12251186cc542251d92081075b94c7e9250b1b654d4cf287c24166eee1c6751eac7f4
zb50afc677ed2470cf3d6d46fee8dfb199463b1ab65bf85f372e8f3e0e35c26815d7d77433cefcd
zd77f270232db87edfe61a9653d726350ed81733813c3d329f0f27cc30d2df2bd7899e80b773921
z513166e923b703bcda17952af59b1fc6d7c3b87bd098586a752ec39189498de333533f9cea4aa5
z818b30994e8938c9bcfc186b77fa19f1dbc6bd2f6ea7f3d57e36c008fc299a2bdd9b8fb4aa866f
zdbce1849bda1f1fa3e7668193cd1b8f78fa42709cccb56a0035920a6ff06975e9e42abfce7fbf7
z9d82eacb0e0b2821fadf556b4582a25ea3adf9823903b7867c1c2cad25f12e0ef17ca475192eeb
z53c51ba10eb050f8660e9d2076531b5e71486b7f64ac52559d1e55cadc318463ff28195db63b00
zf38211d2e11d627b1328f2b2701cba1b125994316bb85b54a5c901bad5427461b765d67547ff50
z984d70965a82197aa5d1ad0a6275912f886f5e21b6b1fff12b9a7d6aaef2bfb9a6d02ca4ff9f70
z0532ae79b73f06a5370b5f187ad95890a8e18bddae93bad5b0eab27d5d362c78a8d543ab1507fc
z684017e55b18dfde1391514f1f5eb434ac0827b936bd9bbf169fe4bd9d6a99c9fad96bbe1436f0
z673a478d2f9809c106ec791869be8b672bfc638392a19789c40e8d4ea5293fe3a409fc1faa9a3c
z022022dc87a49bd45521893fa2aa53332259eaeb17032c88a7f9d5cdefc86e496dec379d908a0c
z9978d293891d161794d067660159aa852deb2d584d22e209a7880eb5fe7a87ecfa10df8d6dfdd8
z7afc70316b66f8f33ed2c3d1eccd4f91ccd6a06c58b530145e4b72413157bc2b741e74fb05a859
z10c1fc65759b9aed78bc90b043a4d10adf052fbb98c1be91d08fd3223b9bbf611a1266e3eeaed0
z16f0de8a482b128fe4412fc666636c1252d5a20aef137b329bec09cae1f4c3ae297ebd3d4ed141
ze1c2751e47a9473d8c0b86b08e742d571d5d8b451fc6fc2edcf321494431654bdc8cce734bccbe
z45b98714fe80f6a6fe38b6228eb2af4f9ef4299d2ea19cccf00564ef7a7c4262a48c14d8705f5a
z0bfa6dbd1468c12c6e3809e1b1a396aa6ad654a3f64c8ef1597556d8923a365723fa391052dfec
zf248ec909707532dd00f66ae78fd79399b6180d295436ef07ab93df097dc092690eb68531584a6
za216c572ab712e286bbc66f9a74a7eac2c340ad044c1377a5d447abb06efadd34c49f7fdcf0c29
z80028c305cf5e2b2d00ba6c0a9375162e6deac9c00027e4dc741f985ac8dc5e28dfbb3fa146211
z51c5347a87987c95eb2bc61e1ba771ee1ba78f0a7cf096c908cd184515212131a12cf54887ffdd
zce7dd7e9605e30dc57686dab43868c694f7a9d9fac2bfd4468749f73cfec9f1eefc11f56f3d4a0
z95f31210041791ecf882ecb8caf28621724d0c90137935337e4d931ef7899b07e2b24cf16eb6c6
z68b39fa16f97294744de513610a56358ad5b53eb9247e0bfa4d09a93a712c3c56d1022e275a49f
ze4f33d77c65983775d593bf24280415f751663c9ef3bf615909d9843a3d339b887e817da93dec9
zfd1fe8f1e1bc16eb870f3be91cd43ef851103278c29a1733536e640bf8e813f20f7b8b16e4aa2c
zfbd3e301a3f270c20febdae6560822d78a7aa465b28b50feb9b42ceba69a9ab259f772c8e18e9b
zb7288685135eb49d2292b88c71c0dc27eb0c4552b9a0c13a9d7f5b790a5e069b26d0613f052849
z144d9ef93a4520162b9dc79e7f1f9d4b6b17cce28fb080ecdd6da995a71a39caed89d532a29a31
zb8e37526b14887bd4ccbae5ecf23b1285ec3f0f28c531791c3de8fdbf979bf570644b3d47e522a
zc98dc0b44558a65d0f3b2deb72fcfd62c1ff32569d21d89f64b76f2c08ad5f21da8c9b58dcbdbe
z81fb0b2304f2f61c4dcb2c0034f3e3728f67526e28cad5356ce7f3f1c0ab4f90de62e06c09861a
z60ac0b6a4cd6e733f84412e07a408d023e688c95b18944ff78827a90cbe7c28718d1060d190258
z48fe8054d8130be7a7cb64547669d51f137081935f9c70b2b8ed7049aa1b4743e6bac4866cae44
za38bf1732e3b52e76f3d145464308b1593f466db291ca1437f505d962558538953d648fa101aed
z3413785337bfb451a2a05311afc4cf72854ab052e5b64db2bcda809cd6865df7f19bef4f488cee
zf5b98d7c812988bf0205ad92770e37c32828a05b5ae69c8dda402d3fef7291a9f49b80a0718595
zce722e8c85dbab0d40c9b4a5ee2709a95e05eec55ec6ac7b88d0429ff5290a8c13afdbed813415
z08e9ad7749ab9a540ffe9f0239c1c3dcf57aeeeb7ea3acc101a1b98caa4cb2abffbbecde8d473c
z1f8cfa83462e1bcc5aed56b4af579c03fecff419e324394956b831310053db7946ab4740133f13
z3eb8b3befe29c9a9c5ad2b67deb5b1ed793e96d337bed380f124594e4f7b715daa8d5983f2ef2f
z65558c2b75496c7d8771ba0d666cae0883e6f14c350f922c88c86d77fa8e5c33781eba6b46a72d
z8f49cf32860f4156f262d312cd93bc216d1b077c38f29818b21074a6b08d0727698715292b6ff1
z2769c56e959eab337327fc2478da3395aef876f7cd7f817494d50d5dc309c318011d92764a3fc0
zd25a6098fde6533d0575b9afc8e00a0a6f9b40baca9291994709b09631565ff6e9c4c6841f5239
zf47f0c176ddf02fc292ddf408ca9f0602fd47f404eca2c982c246ba014f6a177e7b575bc070b03
z0669dafddafaa0de1e119d86ecb642602558d2d0950592023cf4ffd30c8a0be74b7ec6d7b45284
z85599c87a15a653bf54b03b18196680d1f4ce8572fdb2a5d0804760a6a766307a317f27aafc1a1
zd81fac65a5a348c02b0f2e4346a924a9ded53619b36fba1229b2320f351ee5837f635e7a379d89
zbe8dbe5764c517658f358d1c763c43cd84982f9ece285888db25efea3e246c88fb80097a89e6a7
z7713ada1ad4c70f0ba8403b177508531adf91b40350722b95c947636905fc485a9562d710630cb
zac7e4116af92e8222d647cda7cc2dad3c13aece85ea6cad04886b89b37c29309386b6ec12dff3d
ze0be334876dbeb0e6a606006f822a63d68d1e559c0ce2249df1b81ac32c68afd0f8d76e0c53c6a
zefd77d5e3aa475a89ad867c1845f857a240a1dd18f04bbdcb656b81d5c838354ae3190ae832e4d
z5bd068f387a162c25a54a6f0636aa8019e7e06831fef7862b3c54981275f88470cbc7c13060ac2
za96fe4b799a08b779add171ad04d8e4c38a612ca54b936209322e6ce5395b5b8cb7b09117addc1
zea7257d82ac06f4f60e11be4ee4aa8dc65f1788f1ee23e9417660c86e873562aea89e0a10d80f7
zc4f5c391a89e2b83f415a33a773282d8aa5f9f6ec58ca95413ae83cc31a1f35fda96173330e260
z4e65af68b9455176bacd5a3d5cd0a555a14da5486e191b8126410d270bfd60529fbfa298993edb
z89079fe44269031b88cf13351d72fdb8197f78807654558d2119fe0714263e6ab63816af2e7be5
z6ab8f31f677f6823964ac00ff2fba90b3be65fe920a0b8b0b71df507667c5f349418f0d0909b44
z5f3596c1411a7402bd41bfe4484516116331fdfb55d73060a9a70a17bceef2f35f33316be05cc4
z8a3dcc81551e06cfcc4ee61bf4044acf8159fed2b09a78d5d11cb3d7b3634f13275d6c040f8266
z3019500412abd64558ba5e3d9bccd5133b56839e4d2a500529ab234c7f89dbda41f2ccd211e428
z7463b7e37cecdead9cbe6fb4295bf6353a61ec8fe20d1cad4f15553158b641a553c214737ebb9d
zdb9f8ab8c0c43bc845e4e48b91d959ebb0ef156567e3bfe024f48c4d1d7b09f05f38b097a5f1c4
za6abb40e42b472bc7741a97d7ed72884b62f020033cebff973a03b1ea805ffb558ee39578ba04f
z94807705f5235d350a72ee578db0a2541eb2566403ddbdddf9cae5b41d04541dbf8bdc5fa0c3e6
zdb8c2875e298bfa48736c7b5a941a13da998e6293ac6783f2da500d8ceeafdc9b3092db49a04d9
zb747b154e9c9262cea135f262f8492b0f537223889c276430207f9eefd0dbb90b7beb845d72e50
z29eeb19b182aebc5d5ad6064b703abfebc8eed1bd6f59c8642d411ddc4801e1339feb1db0c1cd8
za441b7ea24686b97d955e6f964beb2d96959418d353666bdcdcfa8bc9ad649d2c8d871fd31cccf
z46621d03792ece07b09dc0310a5a14320b528a84b53d2e5907e8b22d19ca8583a9556e4c99767b
z3c027687c0868ef7b28a3e169897f261e40b8b2046f338415bfd3d4744f13cecbe1cc03eabc3db
z5c8261f70d081636c2f87d07b4fe488a8e65d9e504986b31c941a531d04b93efb479f45a1c5a96
z6acdd7e1eafb81be4f43a40defb80db3edf8f35000a457715d7612cf9612eda37c6dd6b04e301b
z595f540cc86d978c2f2bed55f90f055216bf8e752520a4a6ff58792c59d8b4f1d31376ff51c819
ze0917fc57990ef3b0a9e49076c6d630f2acba60d4601c19a721f4b6b8f9cbb7124b75f12b12f32
z31a88dddf7d834685ab5393239350d099d8d44cf41e5c3a259acfebcc66ab1461b7777b45b0909
zb88ac4b55b60118a5ff5fa9a20ced728c808c3da6ee48a207078dc40d64792cfe0f927631ee393
z3bef843216407841402a8f6bf6b4b57ea57d02f7a15c69542779e6c7d82ae6174d20390ffeb83a
ze6dfc0d2677811ee0b9e4a97bd6333a27e3093e8aefb3a1761dfa5d2d43fc1f6fb504af595f1de
zef0f3590122afd68fe63e98bd298e20c75ab9cf4317ffa3a6a7d2ea93ae52b40e909d98f7474f1
zbf4e281d7a7a43397967dd8d2e05666b95288cf710607ed6569609337f7d74fb3c526408c12e78
z2637b16c890594f82a829c8a92ccf58377d49c02e224a80889c2831733ae4cc28565c208c8a751
z618412bd1a171b9d5926228baccfb380abcb69bc727c9251a4e4cd305ae42b3c7eae008709b392
za14eb6c7ce5199eb97a2dcfc9cf81b8b915978fd5acd9fb3d36d76793b65f35b5756b67d1b0955
zea38704671004fb0b96db1218e1625b6872c2e4d12fc078b986e613b02af9c4ad8c180a06dda50
zc187d4077c0ecd814a424e16099aa7ca8d48024c2cfded22c63d06a18f02959c500aabd01e309b
z48c2190df93784c5089280124f612b8f4a3bfaaaf736c707c99164dfc96d73dca54ba8e4acee43
za2f760e9400ae705f9bc9611db0a9b73758d38706f6a3d18b3cf91209e1ffa361117934096fa2c
ze45c15e099d50d7e6309f2a8700a2d597497de5ede473686474df7121cb993e87e30d3882ba153
zebaf303b409028964a95ff4220ea9b8cedfea540c94b8db1370caede0bcb98744a3fae9b2ee129
zc1f1e4cce82cb9264dccdbbeed3445a69e29fb365fb2e7b05572b6acfff4b4b5e6389a8a75a716
zb91e77298e23eb3a4396c57ee1aaecefee6785e42daec296fac1a404691ec1fa7f05839eb56d8b
zf6411e3cb4bdc26708f5a97dcb15ce59de342b3732262b5bcfce4989dcdefc4f9e40a00344274c
zc5f05c38efe8e68064773eb84aedf942c124a5477f53252941de8b7f2291ba7290861b65509745
za474072d7f35a853f7527061fe63df5e6fab61d453cea8f4a68ae5f8e6f2a5f755b35ed79ca611
zf3abd39675e78694e9486096a1de4b9581ce5f3d0df6e8066da674c23ccb3fac4f08615ddd21ba
zbde7906eecdf1ee55755941d2f4e801d1b26cb13ee7f6c027543cc44efd4a48174abd1277eda0b
z6c9d5f95d4d16c8a863727c2ab6add7b49d9af0ef1da9caf89e902b65c4ecfff4f1272a23f78b8
z9ceb19a112abade9a25aaa54b3c04f71110532212095abb9b0e4165cf3397df98eb13cebb7cc74
z154e010f72fa8fde1a18d69f1bbd3a3ceb9fe9b60f9b461c8ec5b360e2339a0aecab14a7b3656d
zb17fd818d45eb3f86b84fab0081b63fc923d75a6a13d5f0631566a5ab15c9c70c57ab4887cf540
z986ac8f593c8ccc8e5b415c25366a990a3a37d6997f00269c5c35d3ba5ce7f49cb9860b0687a42
z41ebc7b099554e4268821a2bceb70aae51872c890ac72e200d9ba6e68932174a61ea75eed7e743
z3920f7af7e4328ca44081538373ff0363901ca0bd8da98abcd61780285dad44d87c47bfe824838
z36e599e3c2c75add89dd3f92b8f5d5b04bcd604531d8848b3327d5f772b1faa4ed07b298c29b3e
zd872c9d4fe0da0ce0bbcaa616306e51b357c458a0acaa5aceeac6042a715671abbf428bb1c2bff
z782d5c478002de15bf7d4e1b6156f0d99cc6202c50f3f4a33872cb708e8c2c14e939ea90ab6e6d
z1f048c139406c6a53358a08d66c97dd11d6fb1b99b667c56c3613169eef654059d814a565e13b5
z0b4e02475939bfca9ac768230bb22dbe1d6aae3a84e99cc2f45d0a63a7cac126480cf208f39b9f
zfb45eb31b754799fd17219694d9c056eed52f25692ce1cb90dbe5e9b907bed8f9791ea4bc75524
z674985057fd10d266dc187bc30c2e9b7848b871ae3ce008f10766608b43498405b74bd4ed26ced
z0f3db5b317edbad2aa6ce4c840c1e9fbb84dc8da9896aa86f2959a1b539352eb4c8af06963758c
z998b8b73d1879f1911133221b0fc406196b2173bdcd687fe6d0a8c1be77af3d2fbfc07e9365b30
z2f14e29d29c4271244db8f4e295775a8635af015b889e8759dc51a95dc548e5b1396c635654ef4
za3f82921376b4993cdea80a644973f5a6d7a1ecb8912641d8eb50bfba226f74fa57daf043438cf
z6b598273956e2709337df09afcaffa685a0ad340e6d931c90879be874f5ff0429442d4f45b0ad5
z58c414330a8da6b33bd67f09e7250e82b235720d2c3e9ca96666737dfaf1c92cc230b3b5b7aa79
z72b22fcc62d069414d71054d67e6ad82c20f087bc154aea56f6d0b4cb6b7df0451b2a0a121912e
ze9a013a8ade6b26b16894e341ced659f184cf41b585d34b0afedd6929004a0183f14ef2fda5c74
z5c6664d07a19cf2644666f67c27a81e66b169eca2656d9deb4caaa35205f2404851114fbeeca40
z831f9a2a53c3e228ac0c8a95b1a92aa9f0d398833a9cbfa19ff23d5a5a42facc6a5251cea6bca0
z6d6f2b5da26d9d7f917b7524234c3cbb9ce9869fd35a07d8b0ea99b251ddfd43c9e46b003f21c1
z58e36260cadbbe3f6ea2bd3767156d82cd01111a020157326065f0d75c8c0936a23abc65abc457
z7380885d590dd74f8166dae04ef27696efbc4162aaec39fe295cb4ebb774e588a056f937a76115
zb4a3c4bb49faadae1000fb10eba461055f0340ff3865f4e55b5d2344d86b2521ed5f126de29318
zcd657d4a56fa8be851d30b1099e8a5e7fd2a17e2d2c831bb025f02092af62b5eecd9670b8da624
z8560ccddcd136155de1c4c95eadea42bce64b35572e7741aae248520655df4b803086733e7cb02
z7c6600e1a2e89b6fe05221125936474363b5ddcc47a27d3d2a797640e331df9baf276f7dc88dd4
zce3f00e149ce8c7599da4ed4e50f7f7a9534e80f1e797cba568e5b41fa7fd34f584fcbaa40584b
z0e1312cc06af61d8ac93ad5542b1dc29353a28a6eca73999f4ae26a715b524bb0051cd8ee6437a
zbcf20a1518320bc300132e7ede991dc21385a85d491b24dd9047944f92db0d25e36bf305abf30e
z49d2b9d958339a8f7883436a2bac91247face47616d5928ba296ba2e8c835eb6922676dd0a8cef
z89fa3cb4999c4c3332fdd3d3371e201cd6389e2f4fff1ee9c61e50dd4fade58577e9fba886ee8f
z7baffac711611bc6d006eb1807f424a135c238b18b47a64fb6dfb791a9b5fd3177f11dc62ede39
zbc96ebbb7aa65015e0f05f63e78afee28ca4b304366f423c9de678ae1bd15a723af28e79cbea29
z698dd60c946c964034d4067c50f1d836b632ac393eb6a61aadee8dc6da7a4c0f4536605ccd3b1f
zf550afd8874cd206746e417d76d18ad9fea69572d17d4b690734515f48094b9d4796d6fc915d60
zcf9d906f9fa0c0ed3301b8d8070f59bce17f8b81dbdcc4b512b7d96011941be30936f9e6063033
z2ce11a59fde02f027ea04779a8b3293208027ed337af1bbd6fc31d51cfc439c5c5e12feb981700
zf79792ef6c60beb2177611200bc480bd7a6665ad92cf6c5fd3fb598a6a958322b5281f9a45cc95
z4155f3a053f911e8bff8d9b983ff002425f015122c6890d051a6488e1a3cd18ef18c69c10e0889
zbbaa7ff446d0862bcb55923091f344e7652fa44d3bfd82071be8e123727f7205b4ca733791ce3a
ze882f3e3806a9c4d4ac69cd5f3f372ba5a519a6a6136f78c8320be98a4ca8a20aada0f85c91601
z9fa5fae1960aeec2a21ab9829e04f54c253171b92c3e45993f978b215131db7553569639cce6a3
za98837951a5bb696960108b51d3839d908b86c82c012b423adf7e140e344c4a073d0f928bafbc6
z612cde53fb69738bf2ac5212a5392f4848e3986779a8b3ccff9657a826ba71a2e062beaaeb24af
z2d209f81eae9649b15e467582e20913b70f273cb72f85df7d968de3e10344a0470eb74c0073b2f
zf44ca66e6e63c66c2e3c2fa0603ef135c30f2976807e3d19ae4f84edab0b31e635f5d931ae06ca
za8b64757f7a7d0201bbf9565099402f96075b933846950068df26b204d502f6ee2ab1499102e7a
z430d6a7c088e107ce6df116edddebef39edda6bf2f12c895937871569f73f747bd55f017c6769c
z8f128c73f0ddcb5db0774f2c97a6bedb601605246a224370841389d0528026f4ae63b6b1354f2e
z45a0cbe24b8918c44a057a0533f1519de46caa77dc87c1c9f25d7391a5275126479ff0428df7ba
z78fa24f37cb5117106def17bbfe8bc8d6d6234f5cebc7c16781fd3971f0684b587584c9d002e3d
za25d2df02392f8b6bba72d7bbf75a06993ad3a2544a33dc5106dd492bfea4d25a609c4ac5ee7c0
zba4e01a65dcf6b903de7023ea34aecc63f3769c245793a492f553064a7b1a448a6fc28838442e5
zddea60fe42a2b92a34dab2398b11d7e54d85d03f78a38e29d21099be5cb3f3ea04e902a0ea70f8
zea2bdc82cb9a6eaec0c09f4e7caa4fd08a4b794eadea73c2e7c0f9f1e5d5fe63c2388c7b3178d0
zca23b7da0488636581fc971b9b9618a456fddcbf8d4ead361f745b728856e5aa4f096b07dc18db
za22d7fa959341b4b07833f8331a74d8beb54eb72d33d458c977ca0c56c21ca7b331aef28ccb40d
zbe68968e10ea7344c3a2135f3eca96c6e2fbd8732f83d6b80b982b482921374db9979c1a6e00b6
ze30c987b71d52a73f8cb2009333e327f8b295e3b0113ab47e1e66577ae8035ea1ce3422ee48796
z13ab91f27614026b4721b60968c4eeebbe24b0a3242b7e41b644e29338a770fd42f180474b7f93
zfb1b03e23ded9c500eb26fc2cd0603cfe3d78729de3a2695dd170e63bd8005fddc8292b86ca101
z50d729349fb5f1a144b22fd3f1579259301298195a3aab5fc69ff246e2a78e7b982ad3cf973ff9
z1a5519230c5f8c2e2720ed923a15ceca161a35ba8d543c348e509b14a582e743ca52b13c0745e6
z3b89a1b51ea2a685fa7cb362b676deffd1db7e555eabedc0431cd6505c873b36b318a88980fd48
zcc5630171d7a1d3c8abf49074f056666b767ee688e02ee14d5057105f34f8b0214737e5b9ab0bd
zc0dc23a6f2f029ac30de6ae64e54c3eb3edecda56c8952dbc5b0680141188b322cb3ef5bcc34e9
zc3d478495843e1f314b347833a3ae2ec830eaa2b4c5ade8dc152359ba08fbfebab4ae6328df2d2
ze6977a04f542dee847688a4b443c1320cba7b070f25e6703e24a661fa477abeefb00ecb62c7ff9
zfe49a9e3dcda9cdcd5663b36d0db127b749e9e63fba61806ed8adfb8a8e5836d3b264ae6633154
ze4a1a61a3d2b454dc92555c76c8426f131b1e49053b049eb6d28ec2089f3b332b0b035d15a218a
z2ef309ed67915130027f2026dbcdd3c8e1506d9a820fff3ed3a10bcf9d77c553266163e1627ebe
z79dd5a986a70e2e615ad00bc0495afbf9b97b6001fee721ca5eb8d10ea3ba8728d258f744987de
zb1f84bbb2848a4d2368c04ece2e36ced4384b01d1fd4016b83d9d4929d337c4eed681691cfe325
z021871f11789bd7a43236ab095fb59abb93732f08617773b52c07d10e9f742e090346d71203b2c
z373951ca244c72da498518ca441704f46745b8408348b25498e687a0750d5cfda8c9197ef5a20a
z7992028655b1e9f4ab2ecae721002ef282d975bd71c67b37303c90856a85cfcd1647788fc57b0a
zc9a461a9b80d257ca01c46e32a6769b82af8d5551645ccf7a35aa93d054a66e7e86bf2246e9a2b
z7afdc65f1e7df43690f6d0bd61320a2c76c6c163a352d7d9a4501069f9335837bd6e8a9307530b
z080a7ffbeace334c6b585965c7c53d7e901baf67401a524a19f82e07326012d79fa59c83972e50
zdea30bd24afb8b558150de5e5a7fb52872dc49cff86a7d5be7ab7962ae147665ce3efe773fbd18
z6c5dd4b82ae6f6fb176f1b1f42d16a9010f3d07a41d52396c692b1b0b1f38ffd59e102b4c9c2bb
zaaf82033f6f5836b3448febbd5437cbe0176e5b8b6d56101826d3422b5bdcc0d3fb885f8a0e8be
z6d69451a719348b77672db244321a02f0bf609b43b4a149b52be24a9fcf28a0f974b126078e129
z06172b844ed6910c785fe8f0d8a74ab00c4a3fea58478a661476f12a88b3c62e41a110879de4fc
z6897f9421e53ac170025908f3ab50dc1c4db2e9df8829f4e56dede7e1ded650f25c92a1fb4895c
zf320799caf660009d013e0f0d06d541e216914df0523368098af7159fe1f7aa36ca3631c263d7b
zd639f2725795fc6ad0f4deb0956e703c9e52052d0e0ee02827e03840cdd3b7ed87f529b04aba67
zb6e8d67759bf47a1eb84df6423173880e6407c55be1e5e7d609b84937898dc2d7aed4511a60c58
zeada18db4d1f6f758ed916b597335cc200bb364c5312aa3a9378fea445c40bc0eed8855c5c8565
z184af31977ec493ab77f18c0869faf8fdf5973de513ff0aee7ac342040c44f294c4f3bce25daed
zb39568d8fb0aae2e7d30975e18cda712c21f86e63cd811375f7962c6ad4d203361bea544a0bc39
z860bb4787529460d244d0188c71bac9964394b843ef1a38a5c523c2026128c58f49fb300a44aab
z341452cc6486bc3036f256f3aa0207d2d7edba0b4786d61378db805012f9e7ec955f7332418579
z5407bd112c766d0839a5ad8853804c8d6291a581eea0b34a2c34308fe5f7fb14740fa2ec58292f
zcf2f80a7af114d956a128dd5a97a6307c41bb1236a6414c5a02d8da7c6b62cb40865bdc1cced5e
zb875dac6c0bb4983199a155c34d6a30ea55c7e06063e0078c7dd3a0e586fd4303d36132f98db93
za44f5112ec5fcd35200a65dfe3461b729556cf3ff1a0179163a15d76ece21bd82ead7bba161b6f
zb603f3ad569f5abfa68aac9437344f9824a64c411aa15ce222829de75f64cb747c60fe4358f7d3
z0ec250a53510c276674e90de98f7f1f78ab20478ffa71526e8a36429fa62f2c4a1e3080b29e8f2
z88575ddb51cc9fcdf344cacf5d540b73e37f4e6df62de654c704aa090a77868fe2b226bff8f90a
zd30504f7074f051c210b90719fac8da6d8bb7d887645518ac04ec1f08f22662282fe29db363cf4
z89efdb9d2128000c98eaf80603ee5f2d1f535d53e3c7dae5276b585f34c6c8709e122bee3edb86
z93bae72a11a5eb2aa9a0f5f4fba1271cd913659a0af682ee9c1513a214e7829207c99b252f65e4
zbc2b639a4243fa9665cb2dc155980f4c001435a5056c38b2da0ec05a6e8955741bceb40d1679a0
z450f8176ae7727661e90b58fc9f26ed8309cde3054bff3012e56c1856167c33c69843b45231eb6
z4ce4100c2090a2896a78e350e607e3268152c05f70bc427681b2603c7b2dee72cc52071d1e83fc
zd2c00b3ba04c7b965438a38d0f921236baec82b6edc1729b2b4783c85eb8eb5aef55f079af6794
ze4ccbc3b75d46a42be70b5beee4788bfb1a1884333cf8d7e1dd2708d3a2704e88dd3d76bcdde2b
z670d72f90677ef19795fd128498c155e64fdd11c56dd2b1bfe60b26172845efed43a728947c644
z0cc4d092be3b3cc28c77c5b6e6ba5896098623173f857b2d8aaa82bcff49a10ad6e109076c56da
z8caf03e7c98cb681febc02c28f9b90958232bb44d81422b0938aa415d1de2b1cd61eb4d14b80fa
z9bfb168605f6341a30f0b5637f6d835eaa34457efe6025c85622d6e54bfd8d7cc76eb9d607e48f
z0d1dedd812add0f55ae7927d1b99c93d33d41e5412ab570dd5d8b4b75c9022c81e7755297b7ba2
z37f9c751c61614278d3693b5c1cc1a43963720f03f9dd4109cf85d875050538298365a1a5bfb91
z1110a44f1d316c34391e7c1d10d0ad4d48f9db45ee8d02f9be76deb3335820250e1db01db883e1
z0c66fccac07055c8276309d18e99a5d9c323ad70934e2444e45cd27de19a42a410ed0f5153a742
z69cd2c2feb17416ed46e2adc2e1d38c1a76ec9303d6915fadbc567b2987083959c557705003ee3
zecbea1be1028d7fe243538f10d7c8a88c12b3c2ec668c05167a35e9742a85d00f70de3ffbdba4a
z502c7964c68f4ba62b7a05225d57b77e954ec5da3a2482046e0436b14e4bbc46d237b3b43ed39a
z8f47702ca077736077e4a401f43dd79efe22b6d6ca96825b9d057c79c31c0952a076c89c7d2a6a
z5dba166cb2933948689dec7ac833057a930f2ccf9140c2e2a397dde7715315ece38083eb733bb4
ze07c0b881edcc7daf99578bb4a0c3cc99f4d96c175b21d19df13f997429f569a0bb4d7e37b5965
zf255deef4a108ad3937c11e4d0e1d561da369602ffe49343e31c911b38b01173a0955c5b2fbfd6
zc978eaf24edd85d260ef6fd9805d82ede9aa1190247816861d3d1be39032178e752cff3469c11c
zc5c7df2931b511d8a1b36704ed8a6a47d009532a41b4b2b6b31631597d15da287e5e5ba8de0ebb
za01d31eb5ef16f9339afe80ff61abe3c26e0babab7673e2298a2b482e892aec815637f7660b025
zc3b885eb64b50586caff94109e8f2fd0b8c57ea8d9bc658b286799534cbf5692dc402d635159c3
z7d0cbbd9b2396dbbe7c4f585672feb8a29a93f0126f778e7b8b7dc95bd481e09575dc570e16658
z2e14c73ff846c8f34d3fa15d5baa27e8832bf2ad5623fdf750494199094e0e230728f443f9ee98
z0344305621990416e467d69b3da87bed732320d462e0cf40174b7c13dfe35027643c3400871722
z91a3b51d3e8614979ec6bf2e4d92e1a57bc8fcaeb32947be114331c073e89e64c570be4a4b0a30
z13587f8569319630e73814fd321d758c927755f952de16b17aef56897860139f44b8e8126e40d5
zf6aed554d444be0240292ff4d7a6b6d80c6f5266cee7c7375837cf63f8754b69daae6df6ab3f6d
z7b2848044e42075998474b4d3adaccb6e6023e6947dcbc2fd8127444b4ae5032fdf4f882eef651
z9e7c94758f311889dd1adf2297d24d0b2f3f15a69b73bd92716dda448038777bb65203ca6de7b7
z912f71bf7ff04815a0305203bd45e61b2b4c4a7c6bcf8d49bdd41d3afba857c80c53c4c57f8ed2
z3b57609e8f46240621e4e46baf2623531452002da4260b3236f2f8ce19575f2402afa5d5a6d91f
z5704b3f092611e409e120b3cbe9f20f718714ef247f6fb3ba59b1217e47e91f5537e7289ee3823
z77ae088862aaaa1d134301c9672d14903e46817904a78d241fe5f5b50e3e2d788faebed695da13
za4e16d501330c3cfc521ff0fdb8f6941f7d841a1db3aaa626b993e76f9710f4aff0d7ef266afc6
z029136e636099b3d0de0da99533bf577c6c28190e6cde13723e27cbb6d12c5f005ac1956dc534b
z617822d2b86baec4b56d231f3659d86fd4b8e7584856afabe75987403eed598e28feb767c2745d
zc21535fa87f900615510b8830db19442e66fcd450b3b0945b69c236a8f6a363779e34966d7e150
ze8f5bfe63407506403286d861d3d7081ab7a773f8dde2e1e4cc6818c9263cf545c2ed121b1f905
ze04636b7039954aeb77ae10473f7c19ee0b2971a9408eff2c2d3c340d4c73f4c1e2b60362eb687
z5bb1f047becd0613cc5940d3718e53e28961a835ddee8709573d1486d22b0aa9072387d58527fd
z76dd657af0038fac2de9e1d2b084789acfcacfb21fa7f65c80236f8d86f67cd9b37e898cdc8aa7
ze200dc6972f4088c22ed301e5f0922612a8672c201187bf9fc2226fee6630f0c301ce0b780288d
z15e4a65f5723cf7b817621ddd1ad43cd0e3bb1a2f8c347c0a4b428912e538ab2cf64cb71f8f1e7
z617d6f5fa0533fa7096cecc58477537506a6ed1c39549d5fef552d1b1a368bb77ae2b683999c98
z5ce50bd13fb1b95d0b21ff1025e9d5089678007c5da0c1dca89c2763939c65eba506ec84cd98bf
z0b5294e02fca90b2eced0d1225381f3a13f006f137e31eaf7144474b3e6445ec972890d8fce155
z5a0144314f74580565ebc24f04e311faf31eda761ee20cd89511d63d83582be172bff57f54cf98
z9241af9120d7ec47c877331e97a58fb6727c4f5db89f22378b14c72de21f64b5f37e6686b371bf
z6fe6039f57510aa773a93d795216018ce65bf51812a17669482f03e1b46aa5cc42c1b8066fe459
zab13d6070620f997e746c8522312fa4d2f057ea5e42a0a71e9358da643890c5e7d284f320ef5d7
z1ad933b21e476cf0d057715135c6627d1ca80b7dffcb9e78f40514056e6b410a3e90af7064ac70
z1497a63535ed1d122c65d5b90335e75b48c78c2cea8953b8f7da46ae54c267b8462b730ef747a2
z4a725b55133508cd2dd2cd488476474ebf0b7e89481c31a8382a8ba2efcd8d563de3ffdd2b5e32
z008368e2632dfdf2ee07b2be86ba829b237bc75824c64950aa81eba62b4c924cc8e8c9d7f9fe9e
zc66b31c5cc86c3571e36afbda30e346030ebd2007986f64ae39828b3bd5672be258611d086d92e
zb63ea4e2916a41dd68201e8a3b18f28a817b21bddd01ba39998a11caa174c9382713152812f44c
z1342b7e202800fff05eb4633b048cfe5c1dc508620fb3edb4eed6ce8e2fd527ab213221ef99d12
z508ccf8294496445aba146b375640f377786adecbfde354713f637ca9346cb3f054840a06c440a
zc035a51f472789477a64f377d6d746e6814bedf12fdee8a5faca5b1c086a309e2b05a598ac2060
z91b638ec619d95ff093aa797d12cf942fa1762c56523018eb3fc6d3810f68b14e9851cda2d05c7
z88c7d7c1344537e6fd29d180941c1e0c2087c58c3bbe706233713f25e5b1aecce4d17e221f1942
z31adfacabcf261ac7ac20f5305066ed58ecedcb5efe0ccb795ce1b050f3d9824018787e4c722f8
ze3d131a50d9c758ce26827f3b6b41ed5f659075c391ef494cf37c8b78e02ba85f4f86141e35ae4
z0adc9e9f09622e58967716bd89e97a8b4b158d4348987ec9d0aee5451bfd3fd2d22207a3278f27
zb7f8a168000e2a64bcbb5690c5ed04251267121c9d4eb1ded38f104bb9c44a52adbba6758dc090
z1eda77e4ea96d4c44017afab4034c79e04e801bb3096caa0f1c21598d29c17fc96a3fe4c6e2f54
z0985fe394bdb529a6e77930bd3bcc36c33708dbc18279efdd43a32bfdf1062cc37ff94da2e8203
z26e2ffefdbf47338a2bfcb16001181165c6ad826231ab30c24c760bf0c5a9de3bf0045a31a6f29
ze453d94282ff2e907ef7960475c987488498a6c79a1c6c26aef96d42acff48248e4646426b88f6
z65ac41aa7952a2a20dfee2c0773bcb3f89a516ec6e494b43f201308a7627a7292840484e2aff21
zf53e8b928f408005a58da809c95a7c40e1ac54c36daf25652b97aa40515e4bfaa9c689a3d6e60b
z9d93dd7a2851563eb65ddff0305e3d13b70aa3285defbff127dfe6a0cdd8bde8d8bd939c2c9bf3
z7fa3530d90349e9f2f6a68718a54e1046bbf81f6c919330dc0e887fb17fee6f4e430b02034b155
z01ee1e9e16e62ee3b218c135b65c4176416854c84abb0e3e05df3241772270c7e561e17eae8335
z3f8c355767da5673d0a337a6e760881ebdf2a333fec9fc424ef32be8a560af336fbb7b956cfe5b
z032af7073b4da8674dd70bc5df78303bc9ab030d9d8e8b623d168bfde5b1d3c833f61f7323c0f5
z1a74c2321230293e46b125c8c34f12c40ba27beeea0a1e8c0632a9be1a31ea6571f4308bdd23fb
z03ea04c3e1e9f65e8c3111d4e2775898ec5d3b3bfc9982731e837c20d46eab19c5daf9e5231f22
zf06cbe1b7799cd2fb53b516fc80f46714b144846613825dc029de0b491da91f8cba1977f53e4d7
z512ae4dea6d6d69226c22a674478d3442271232be24f57cb5653af413f22166bcee7bfd5d76eb1
z43de8a516cc1c235f792727c15ce193f020932f0f83014b16764d3b714e91590af549cb23a9a48
z966cc1977f81929be985506f4641120877d2ebf42442d606f493a3eef2b38e0e22f86e4beb4f96
zed2fb7ebb988779ae7849b752484d443a7448b4d4f3c235c299e1b6cc49c4c4463ed7a86bcb644
zf993842fa8dc9a3f91fd1f99228c1260867317a71e1293f7b8927a74898521aef8a2e0be21fb54
zb092facb197ba2f0a1264e9c4cc0be1ead030d2313e58145eff3f6daaf240e794096957591bcd5
z757e2f49c2f719c1fd7d6c69d3d6597b6095d57b71ee5e3424e0532041d73d58bce1d6fcd5a2ec
z9a9c2eefa5c46c00d3bb9873be2e31843ea3c2600ab838566be54b4a66c4ec378a7b7da2bbfbce
z6ee37f0981a56f185132482f125458e3e0e700001dd7040931ed5e44d1764ef7b25ad9057a07f1
zaf35328e56a7949c04e3564306af519d449280df9b57ab453d314925cbac711534495495c99f71
z0b469cb47e873ebe236db71be5f7f9177252f281f578c69789e1ed39a3af1e859b30e8a1bcf8d5
z63ba5a9cd8951fbee779c595ca2d82020b751a5ccf6aefbbf91f1fcd316e45f14147da7ba0d3c5
z6ae924635666888d6f785d93978ed3b05e8022fa068162426cf465f9041a9a51caed59d4c98139
zd4d55a3f9f1ee83249f5010e7b21cad3f638026937116552d9ca785a72cfd6d9db6e1706d82a30
zb1afbe6c907555e46f88ecc94411c7f7b9e2fe1fd3990fa3be82e4909a47c2b56858a3383b86b9
z422dc78df24112f711929acef233aec771434e274c2ab919581d43f12f724ab95ff07c13c6934d
z77c49f2dd5caa76acd0077914787d9d2caa0d8aef5685a9c88c7d28240e0dbaab434798a0de5fa
z74d54db7a6e64c4fa500d92d4cc8e5533e3795c8dbb713128bf20931c894781afc8d04992b3483
z617ba93d2203a6352d04d9a51b4125359d5779db00fd0f11ef8f07f92f2fe58116f0479e838d60
z37d8fca55ab1d12355d69a03103710019dacaaf210a14498fecf943312739acdde8b4a8b822600
z06b2d62476ae228c0e88504c0ce6e345368ccc1f0e3b9969a8ddd24d8a1fee3e41dff9af7cffa5
z0a6df911f893bb6732cd3ebc5d7e0d4885352e02aada6be654f0893d57652172795f10a52acebd
zd92a29eb49c66ec4c554acd22be0db7b72ba45de90754ca1f4a7d3e762e3fb9bb213d6f20a3b83
z678760724ca751dbb057c2dffcd106575555f9da12a3fb6673b2c728cbc344c90d34cb4662da77
z1c7c4afda879b13520f97d91500d4b1fd243c49c15599adf20f1045e5c2a665f38af7f05efe314
zc8636f24b0842398d10f3dc685425c8a0b2089ec0b55fc2611b5f18867ebaab24ac93cd3d8c1ea
zc423f73652a21fdc481735c909d46cf5a418fcfe86357e0d2a92054e2d956af92e4a1f7d7b9ef1
zc7b0df0cb85cc83ee1f8d9cba7cf2d68c1d3679eeade0dd03a229b26e237eb6b8f2b19f5475ba3
z57f833c7df74e1e577f82d71faf44ce300915ab933e03f6abea43edc83b0c25ae138942f0ee5e8
zd8484431c55f5b0e69bc04a17089277ea4b3b3eb0f69ac6eff00c6ef4fe3e62377acec6e4dbc86
zfbc8e22d54147b4ef456041cd65e70305cf9c34b8174c10c6bfc7a390491412539a21c8733fde2
z1bd81c348ec8df041ed122441a6b624c2b1f7bba0f71e3180b745242f2b7c671cf6c97c49b98a4
z605f08edc5971842e8e798fe6a1f06de38e5e4fea5f970eb5e94b6ac1a6fe8d1a766fd2699f0b5
z8b2ea695164f0587573a89b08b4c9dd40e224049acb197882ff7a155aba2ffa7a205220cc6a5ee
z31fd344db1f075744ea858e9e19fd5a04e4f6b56b203764e971df66157275fde96afd273ec37c4
z14a62d90e52f5aa1f5c562b34fbad19bb60b3242832f44d26b9fc9293540359243a3c9f6bc3284
z23e5b6f076d4eb33027ed43a6421ae3084eb3385e0945037b46b062f46545ce525a0ad3801fc05
z4e94d0ccc8e75bcd381b3eddb72d5689e3fc0250cbf8f97eec03ccd55a43e197c89a41387f7765
z1edc1ce094ea3d8be8ecb8b08cb1a82993e5f86ff353009582d14224c7d6b205d0300392f56552
zb35c4ff71491f6a67cc0fe2233cebd8ca0c75b3e5ef31f202d85271527b716e307d4d1cc6d9347
z84855f622bc92726c1a99c78c84d72a39bf0fe71f3e721170fbf66106a002ceabd6a5e0c7778b3
zeba3d30c404d697422a9121d81ff3a4272565c0cfc7c7f4c829b69e6c136f497058ee8ec33ac67
z075ad452646e7dc8e7a776482ae5aff5cf5eccd861540d8c835efbe50357328e658107bf0d722a
z7d5699f8d034337ecc9a6a6a40538af5538fd92ad75810c0b345531e8521fd882265a296871c14
z21e7f3374c69303c3adb2a975676cc3d52ce2566994d76a27e518cdc5b59c589797ad4575935f3
z02c21c6185c65ec5baf87f93b7ea3426ec5baee4858752f1e9d22bb014131415a708c233b01b65
z69aab287da97855b7c1f81ca1fc36f8a3e79b8af7d4442c3908d2b4d26edfa106cf5f0f8dfe0ba
zb46a836e441182f8afd96cb86e29fe74d2d4c34dfd28c0eb870e6d036b7f904e66cc70a5ff0a58
z0e6c9883372cdbefa36779c1aaf8596169a776da0c1fb1affd3a480122e71bab53cbc714adb6f0
zff9e150b53071d376e8b40ea5c39409910796aad40e13bd9edcd89edb8a9a66c885d7710159b47
zae5683704b242c1781df3998de852ff025e99d74be8af74b451e626ef120eda5a5fadb755bafdc
z035d9f6c1b45bae20184ace1ffc539b52ae5ab54d2a693dd9591c8c6d081ad68a7c7eaeb28c6ac
zcf7add644d2506b844c3d9963f90729904d5295a90955fed03da943e92586641553336495919f2
z397d3fc93fad3808ecb6727fd960d0a459cfd052b4144c4ebb727153644ab3425e61133d50ab1d
z1e88639fdb0228751ce23ce820814eed5285ba615811b9cefdb222e2b373177e37ab5216b1c49f
z785d4eaebec9c9a429a8415bce29e9867721c55eb239aa9ed92c9581e3c00089a32f76eeebc2da
z8bb5b0158ce9a7dc1083b2d1fe6d341a91f67cc401aee47e8c3ce3f41b9da861db71c69d421f35
zeae9d0ae07eddf096ec0277a1d36b45507cb9efa7a414ba2383a485780eacce883e419b63e2a5b
z2162255cfc2f4b396d5c52dc2f3e114ea5417a2c6e5df09f488529f248c1dbf5a4c4c3396d2d86
z01f39999c3936f59737c8355c7de11b390852aa75d2193c7cd7acd3632a12c2c20dc55bb0872f8
z9b37490d98b9849b8e4015a386c198a01c298594ef7277d62c5c50c7fc4f03e3a08a103e8f1cd2
z30dc6bfa67402bc58f02f3a0c5249023c52ed8dcf7d3c316a7c2a81e2e85c229488f87f9318187
z702bfa69e00bd3fcb37b6bbaea951a00db6f12b03c3c8d2c215b8a89512a48c9938112bd37acaf
z29d0995479e242d604091b2ec364c3c5292bf347847c327fade36e8745b81a81417ce192019907
z175ce6d98693460ca421e93cba038384cd2c0b02f105d0d9ca8789c65d9a2fa43fcf4456a939da
zf146cd10461e58cd9e259da0a02a5f1d30e262e0c8ee20cc812d01842be7e28c1c88d939c8271e
z8f06562b122e95bb0d4cba4b71f49b9bcace27e2dc4565ccd94e7a0526bf5db554cfdd015bc6c8
zb1bc557d07339ebf87f037cb5e16a7b12a55ecd7c05159638b5ba7baed3b4e414de46cfa932ea1
z3a99d0315ac0214f2419893ee5e751b36f99d0656f1fc68cf4ec963a891e1b38644e7e1ccd469e
z06c4dbaf12c7bc7f01014b2dca543c3cc36f70cd5c2f6fe76be0027d57209983012213b9bc3d82
z79641a32268ffbd1deae75efc084af0fe8611dc658f47ada8e43b5e2dca7ac4c171d32dd35a685
zd4842b0fb1606ef961f41213422f80d417ab6e7403f1000a7b011bca9010853d645c7de365720f
z5b2f4a1b1cb9ba607d230f88c5aca6a04d353a3adc6852235a6838c546ce8e885883f16d012156
zc2c50fb3c1c46c48ed7dd6ec533d740b4db1f8c987d6bc2ccacb798c14421ab4699853b9dcd82e
z4c8f5eabd788831f5d555e5fbab93567d0a6bdea8715305500184fb8b58359c1fc6cf68235f358
zc5a9771626404ed216268ac0336d7588c0264f06f9083bd3fa5076e7daecbb189ad27f30f2adac
z4102f1d69c91e2c1a866ff792564b1ed68e2eb590773008419b2bda95ff6eb3e4f761ff177679d
z11f2382d9808d0232d858a1498c54b9d7b0edc030c876dbb48222663f51092b25f2cd01af034c5
z20d43eeb4c325acc1b9a011e80da54448334e8eec96c54eaa98af0c711b3af760b54e2058a089c
zcfed655e7868cddf2bc8624eb689a5ad9ee296ed9b8dcb90f71dae8b2ae2d32a0674c90b536070
z5a3118c49dea5d8630e4f797e11e97204bcaecb35680434aa797db53e784ec63237e23647ba5b0
z65addef9cc18b570d208975fab529b1400f821456ddd4fa10156b552ca9dca78e2dbcefdcbd999
zcaa3582cddb8f0dd787281a1b1eb274cca3a72be508319d8b33194d55fb53c5e62477a5448ff16
z3209c1919a38b53d4119abbfe09d5298bb25236de70296110cd25d2eddd57f58951ccd9d2cc874
z52f861f5d1be8baff0e8095b1ac6867e6d95377feb3caabf27167a254f5befd7ec6b1abd6a56de
z60211ddd7b88e2f5242f3172137adb39946742c41fa8df034fce89fbf035a292ab8f99a33fd6ce
z1c9248ec7dafee7eba59490715be2b41fbd63fb4e21d2a5f0e1f5aecb2bed8d333f38d6ef08b53
zfe3f71b820319cab0bcb0d0a6b89ee7fcde7103b99b64101cdd9115954e8aaa55f3ed9445af993
zf8031ea1eda3110d5cb8df57db65f8304a73de4d5ea081ccb2cb27ab421952f1fa1e5b4c9b78af
z6d7883f3bd9ae72844cdedcf5d020e67a20b8c7395d495b3b711c13c436ea01d74b05aecf54a34
z69b4ae23b2086e7d8ab381680ef1f0a24f1985618bd76d93a5e28a25d123b3bfe561e4bf5e8604
zb1df4a1d5daecd8452280711f49839f59c6c57b5c65b228c7cf12c8ea28d478c0c2c0c35d03932
z50e8201b502977b747945a54295fbcdf9114d285331151d8cadd0825ed1021400ab3d6ea3c9ea2
z7f0e0dc9f893e45be6ba2ed7993054062ff00b4da0876ef7445d4444f9b209bd0d3f3e19fb8810
z2519369d330b0e1a3e63f9e692f5059044c5364f7c9c0e9ad63d8e0c0293c38da4778df54d67b8
z2d151f8f399a28c1e35b30ae5e90854a3e851a14e0a15690a5b715cb99b43e731bfea44d3b474d
z7c710d8dd089006134598f98d0297e8038b9ce5e154484d39233f6b26929647f66caf6a7f27aad
za2e12115292eccc9be7e6cd813edb084042a17dd2b12e3fc4d68bffe18eb6b9ad994e88292aae6
zb460d210d9364068bd542e0e37b6deafeae4a4624cd6e82bc576dfe8e97bace1274124e9967e65
z2ae0d2c99d28fb7e90d0621a73f155cba1a86bbb44ea3acb7797e26e52113c4ba2721290d7929d
zef88e47db161fb4a447dee8c639be272a87c9922c527d2af2ad7673a4230288a7366e28576e3fc
z6544a835dc5abe451c7dc873d1da928d7c90c3aa7488971f11e124eca9bbe98134fda702c0b334
z2312c57515dc904e1f651a1be368bbf830aef04c139f129dbe3a0d31aabbe5fe99c2d0867f2980
zcd66f3f8e10905c7007a07d93df3b2231a1d6795ba3e134ad1f6af243a981742d0c40525945023
z61a04197a4937ca84455baed8e7b5c65b6dac45651f631eb135e6ffd6a888f4dfde8b279355f6b
z11b69ba66032f453e2207166b79acb7f2b46ed6284f217f33281edd9a0344fb09a086a9e7d883e
za23c9397016de4f50989db2d35a91bc5c860018192db906601b0496282c71bd7fba9609252a19c
zc1d132365d1bc8452191c907d44d6876d441c4017e1b8447c720a65438005493e35f6b8561efd1
z238fe46cc8bddfe854bbf6c5e9d5cad98ef23dd113ab058c2f5075fd5bccf87b3896f110801e48
zc52fb00a297088b2f882a360c79f07187fd6bf8a96244af8d4f8f942bd4bb6a329b8172e473950
zef4bdebaf5c8be3f362453ce6e7451cd94edeabbf2621cb47661172c76d5d4f7d179d024a27401
z8060095942d22a013f696ae0c662670f376157db8d1f60674090328bbaee25f548fe3cc25e912a
z0f5514e2b183040e3e216c2741696536b354fbbb0dd1b9034406303592fa904795e0a48d8cf240
z0bdc24001122f98ea12c2c3ad4a1e7248b9ee6bb44c4862d3f6279b8cb0b863e1068ec6aecc69e
z9abae627a3d05a0cef9dd6a229894d1b49aab7a2ef9d500201e4ff0c2793188ac2a7386a31ea5c
z5a2a189ee03374d4c98eaa72aedf64b4e51f2853e506db68e37a07400049d39224c652540abf86
zdb6053af2a371c4f8e9785c76c267b4b55dd45b2bf20b23e986621ee6c2c9f28907c755755f013
z086253d4d11e23b45bbcbd3bb85701d76d566242a89ec104fb740b14524b8fff56ce0bdfb60df5
zdec44c22595f713a640b1f4a36a5e204eee1aa52b1b6e58251048fc8bbc504ba3935ef0880c921
zbfb8f3e4146e390662411ca6e8d5e0dea4f6d11e87f096b690171151fc78e114892d488a2c2283
zbf10b40d2f05941fe77d4d409176a9afcbad892e72e36a999aa195fe162644df9b68fc07694e53
za491305a3810034ea4b09e8e5a81114635edf8e6238977d1a0cf5abd27e019ad54154a4cf06dd3
z9a7e13af5c1137e634deb5ee0cf8da51174bd3e35922807e0142bab4a5c0f2bf074b6b80ea8357
z8d250e4b516326424d29812e887e83ad3f0659bc7ec62fcc1ab0609d1808abf81d8b6e5bca3d2c
zbbe00a073f4dd45eabc3cb582f8757fdd4d18769968e2f57265a58cdee1476bfa71cdaa97c734c
z7e734785c3c130b1fa84aac66996246d76ef236991163f81cb6703e630dc4d6f05618cc3aefb76
zaf6c38365aac870343a3d0d118894465a74f95e259ca8f32a26bab006e7fd66d564bcf7e418cc5
z1c8756727b67dcc77180cdbb52c73b8fe03739f04cc5ea51a2b610d46096202e2574e43fddacaf
z36e3438d0914d7d3127a7141da6b0bc1db08cef2d51b45fdf90c57acb40ee119896d92ce25a207
z6fad144b6fa7d35cbb1b6558905e0588bdd3eea75c373020d1af5476b868115902140e83410351
z30435e72827a2f48d8beac9d62eebdb4a94a28bee180196db1c0533aa8dfb97dbe1dfe7061dd04
ze2dc0a357e194a6b52b4523f5c272e3462debf2f8309cdcaff504e96a8d28d2d2d60ad648b7e45
z2e6a22736e23dff24d97198bd3211d3d3a80f56712b38616b84a55c083a3047590c524208a4bc6
ze0e8130298370560b30f059e036ed433ca3e337bf2c00dd45dd28c3096dd6ac56389ae337d5a9e
z7da60d2c640fc2d1e67f01169e69205f384f8a71576a470b24dc122ff85ac4bc2d3fd3980e3ed8
z31d23c5a1090b91c0f8bc790d1cdd76a1310f0047bdc1d60509eeebc2c5dfe211fe9254cde17fd
zd7f4ec83552f70de6d1f5610ae6cfcda0c5fec157dc60d95686add3ede92568219099a000b6317
z91f86886bed5364782bdbc66143c082e3162d54f122fe294489a135d320757145267237bb619f0
z8e9f62b057811e7ae9d99dd236e199fedd3db55de6ea1e1cc67812d3c5d5e24c9ec4dcd6e9083e
zcaaa90d5cbd42adad05a675bb7cb48c65f21dda07b29fad2d5dc2fcf2e53793a1805cc54bfe4c2
z1189c10a36ec569b03b043ef46038bc2b1e23c076157cd0369ca0cdb7380125be2f28cb9c980bb
z631734dd78cdf8d4239448e1e4cc75e05561f604c65389b6350f679ef3693b917e16710f253e51
zbd8a0fc1a4967c0aaa8444a5a1766de851cf8c87de49cd3565f5e41b41886276c3b415021cba75
zdcd91a22b7523bee7c9bded217e08f392a1af8bfaf50d0df30047307ffb31a3b67790538d592c0
z787c4c51ebc40327b4854664b9bfe3d6a4d538164bd4d3c731a65b8a72168ef8dd4640763c9527
zd621a296231ed7b41141b59a3247fa3140d0c53daf9790d5271dd376e8751fd292746eb1d18fba
z9e7b13201323e4ebda0341093cb981fadd4d2d89f5f6685de6e26b9ff67c41cefbd63474c6cfed
z16079553fd9e265f49efb378c665cc69002049ef6b178618df4b67342e4a9378cf017e341a86d2
zd7b6081cccc145342feab0bf5d2dc79319e486e4ed193233e45ef057b15026feaa709648fac515
z9e5ca4bb670a1371b3b3ed20a3ac97a9a2603a413b6e72881d34e6799a1e95193b7df12c4bf150
z714424e71b66702751d95fca1b8c27121df3d15bdf651bcccaab9ab322c3eefdb592babe472644
zcb12ff09c278f1bc74e79fd3a1e4f2cd7841f8211719eee5265f2a2a6629878556d656ae10688c
z22310befb1de45d30376b4904ae660bef7c3bec762dc076942445dadb4888cbfa6098e924d6a5f
z42b377b8b85040b261cf5593e80cf491bb6ef14c77b443a803eeabe17cbd1681aed718e285dd6f
z35a5285cbee129b288bf65a44dec35c0d933506c7245018418628f3092dd0e570806edd9221e4e
z25c7f3f54ad782d1879b67dd91286e9eec759df9ac067b1d65fa7dd0797a6b600837cc5ac06df3
za99ed2fe3c6269283b3b0b4b5cbd6519c8c1e09f26aac59c78a718b9251dfd823542ce227a6d46
zac0a92596bd430b7de774a74295ea0ce0bd5d76437ecbebb541d49095132b18c73d8c09c7c1f27
z9476a7f67425192527c265a71d646df77a7bfafccd205ac8d8a85e5da98f7e9d3384bff242afc1
z343e3ac72a46cf68ec501aaedc863455aa235983f3d4898b1611587b70388c09df327beff2f407
zb9eab7fcede26bde796593bb0580534af85796a0fb5146d41332294a83ba88bc2b8ddba77cecc2
z68814e826c76a5ac5d00bb2511e71ea69ed002167f0be47701b74d5840621f568840a42029afdf
z0ea0cc0409290c747b9fd07b737501829d8f97a381d04c89caf9a638f205a77d10e9a790255406
z5a97fb8889984915d7c883d5505a9cda841daa2a2dd6ba6947e9cd171a264a906f4c73a992fd82
z4be822e20100b85e357dd2761435a39d003afb85d5cb5d11ad8882ca86a40298370ef030ccf337
zd57fdefd17de2e7c687a72037564e096e0fd3c7c067aab99ffc84546ef4beb865ff4f459ba3f84
z3115b8988098b08aad1b03b34c9fc175ea31a5b43b043ad5bfe226c7482d5674dae54e5d119cd4
za7901afc538f1313d20c4a4b2d3d6a46c5d04035982a41c9338eea3583823dce252c64558a0eb7
zc34a87441f90815d587763adcc5d352567a91f0143a92e0dd2f4086c52ccddf7d64bb89ea73fbd
z7cb1887c0455e6ae3d60533a86b400f7e4d1098c88fa122deabf046431a574ba6fbbc2e8c70e4e
z70ad9e44daaa6851763f9991f2b473da4da39287594544f0defdc220e31e318e5338d69d315f46
za83fbdc622a299b9374b4a0faed3493d12ac29707e22afa8b6eae63d7e2408ca6896579bff3b03
zeef4340f1a27995f74e4b5ab9f483a7735bc008bcd96dc285cbbdf685650fad643b5c061c845ef
z0237bdbd8626307ac5861832649f50c248df04bbb1104647eb1589fc6e0ba461e0bf87c6adfa34
z118aec28920c4cebe2430e8fb341d8335b5452d6cdc4e59d508a84536c9479fbe9cdd3c1b038f8
zca0d928c3619a93787a6b2c860976abd47f5745855336e6ebf0e32f688547b0e769659928c3c0f
z74f1cc0b76a9cc0c762e753bd930d2498978ecbf46f91b144edec5d7953638ae97cc32abbdeb85
z17b8853895a56fea0bf996ee00ac6a6a6f643f9b3ae935feb7dfc0a3513c8fd0c82b9ac61da8d2
z16ea2b1ba4bbf93e729094426a930ae15e1fafe8d9c638bc6046edbc0406313587b662157fd365
z9bc054efc4dcc2d8093c5046d4eed65a77bdc2c581c47b517f5b6018588c776875926ed8cbdc35
z7adcac353ca0e3d1b9c4963794298bf40f3c2acd37983935c02d3fc41839acdbdcfa8c487acca8
z4c50b995f5ca2ffb6f42ea3f4c18523a3afb237af299a43a2bdc28b1f8c690a0661ded8ae59e76
z852711a349a22d421a94184a57fd6a0d9e41da1eeacf43549164948886d7c79e5f9a25dbad72a2
zee14114cd8bc2bd6ea895aa1cf8100e77cf76eca7c82b434f377a114d72620b0a01425d6965e9d
z35a3bdfb268475be1903d61f7282f3605f763747d4bf35b97e45c989fdabd8ba52e8de60a9cb48
z63442ad560b04cca3c964ad83ca8233f8c280336bef8ff4309bbf609a04a4d05aec072efdfdace
z8f2689859cccc37af053756bede4b7f14056a09cd5bbc3f142a1f2eea6c521c28b3a478b776784
z66dc45206735120786f482377cc1b23b2bbf65a0812c009ac0965832bab03a4d8e194a129bfd0f
z5cf0b72b949f0f01800b7c1de65465fcfc1baca8fe70e70331e1fdd2f9e2dcd0f30030b1b3c748
zf57116644f7b945bac8da5610b343907dbb577a26a19460ec1cbfe713d9d2e07c9bb063243a601
z830b3967437cb383a70cede29293319551671fa5b586232ab3a457e0f9cb7a74d2eb3b77d39c06
zfa76752498983bbeed74fa4dedcd0cfc9c0b926dbf57425e8971c96ceb46530b71f73b13b371f7
z1a9d331bb11af6c0d9487f888fe4ef9035cadc34421b4194492dbdfd8777753877ee71303526f7
z6bcd639340fb9d09d8abb9f7ae4d873f25db85cd4a80076e4d3e15734f93d7faec8b70630d33c8
z3009967e2fa0036bb253bbe6182b2077d601f3e76f0e5d7ca449d48956821e19a63d1bc63d0993
z22064345b65bf0dd1a12c5f61697eb08ec7c51a8133bd222c6a4ee718581c9fa87fcc31e91dd6c
zbbf7e7fb9b393d8bce92f1d6643fb20189097a633e95b1ae72388c63e40ea747631d0c574123af
z6a61ce0fc3f4e9d764380370913316b7d84d3b43afd9cb0e8542e27ca4e397a6952002c0f942f1
z989736ea65413eba8d45a1ee473e8cfbbc5c9f22dbf96039b95f46fe64c7e344bed695ebcc2123
z6f090daf60bf3781dc1ebbec1a0fe32e78f99e44659fa1a4d5922be6e7acb32e29395d43506549
zb5c705728b714f92b0f5b01c1245fa92498c9617a805b09655528b50dd1ace6dca5c202ad678c0
zfac390d6480295fb50f6d9b5f3dca73cbcfcaa93ee96253f16f876ea4f3d8d570f699d2f6462ca
z400f531564804a75958067011e3d3c2149f575899c75cda4117b9f76c640e7778c3a65d8bb4ade
z009de5cd0ce172db10f528f6cbdb3ec6529efc909482a0612381821b8d84bbece624e82d20249d
z8694053f406e1fae62d36696926a35e069cc39c7b6096aa0f3e73f13eb4b7ddc7bcf13aed49bcd
z2ba5180c14c5e3e7757dcaee6e01497c1d5dce357f09d709f2e73c4388313d0634269fe06686d7
ze7f6ad3eeda1e829fc889522918be581a66ef6b936336510724212761739558014fe39b8608a39
za0685cd9ccf2cd2b729c8c176b4035da234b55edfd1e655cdc59bce24c9a749e2bca99cf771db2
z3a656dd82e2bed581c89f99ad7f3e1a301e7cbf643f262f50c2c5012645446da999745ea18f6c4
z6b5c0ea2a80ade8c30bb7afd8c0b782cad1fd2f7a12a35b0a23abafb21abc69a5a058df8da0246
z751d6034f696091995eff8d8865790b50b49ecdbbbcc8954a1a8b6c7bb403d38bd38faeb2248d6
zae26545b196e6982a0c26c91cf8cbf5c577b7b5a4da3023419b4527fe51a8e9acb271469ad8f33
z4d1174a7429d5cb4efa7a9bcb0f77b7bdb93c5753835bdd67353fc4edf11f01bf00077d4d03db6
zcfa7ee636cb6906a615a63dbfd2332bb41316251c3a42e50a5ea4241739e2ce8da9f42d347647c
z2cc2a4b362e60fb8e9b6736ac304ed3980f2cc046cdade8e0fcc0d72ca37bf1ccc3339493d55d7
z722cc734db9a314fd169646dfc0232314b4b7aa6b6138074ac6eb82c3f2a17857f89f8c59b4356
z3762c468a767fa314895edec4bd04fc4c9196341094e4435255c2dde5eb36295c3e0e6b2c7c0a3
z8edac9e94fdceba87b0b19aad5bb83a6a1852c16d0b62f4b6aa5405c7321309b7e56fda64de907
zfcbab56ddebd90f20ee6a199bbc3317c72ad5e3f9d8f4b924980e4996f8186ddc844af05b7dc60
z54442a5317e1b4b89ed3ee58ce86fe10919aec927b65551679b65cd2727421f4413be22eba03d3
z51db0c7a5e9c39b1ca607e90a249467e4842217a9e29bee06a2f03ae39fe925a792e4fecb7aa9d
za28746485489f91c78e3bcbf93dca506ec8b73882c97e24115c9c6bfba6aa22f15ac8de1ef4104
zf7631f1be4375bdcd864ff068401b8652b1b726866e5df5040ca35131a4b9f3f9a203bd42dcabf
z026c971c6954b8ca27df226822f5e4d5bd377e6082f2fecc4ffa15125125fbc7fbf493659777cb
z022a99f0536f55a30f60cd47a4c7651470a89b4377bccf8cd517f36562811258bed1f534fdb6de
z2f841b345c03003dc0ba27e3d8a2d31b4a3669ec27faf0901cca5b82eee1f77b7ba3878c372d4e
z8bf9042e2554302630625bb665eeac192c44b9461f299489b1cf302eabb2fc2bfaca8965f976be
zc5e4e982f40509fe417586babbc9499ebea8c61b072c45fc86217d5730067f09f817a244780249
zc3b5555475bce84dd286fa48887d5af37c1c628a22bb0bfb031fc0581910d39abb08284733255e
z3cc570f927aa574b6725367719fd9d63d125046d6f12e3c486437cefdb4fe45344e8db2716703b
z74fc8474004d8dfb6f14836b43baefffa090db6ff88b1b0f0f1abb5276da13e28554587081fb18
zfc62b9f67385292c060b842dbc31ee8f30433de77d667a49c6f85b9a73e6037106ea9528893cc4
z04d83f76a9b80ad53c71e58e057c9dbc89dbd23e64d69bfb6033e0ca942eef64ac45fe8a4f846a
z21b8c3e011a0ff787de24f6c97380328ee7301a1bcee81a5119237f1c4948edb05ad1cf5fcb320
za1f37df4ca3196e7b24e32d9f410259ab8020e7c3c79d3439aa64fa94a6a1e743f0c9eaf46d19b
z40a84dca0d1dbe030e682af8b0de61e2fb67d5116142a536b58998fafa15a5c226a492b364126a
z1eaf1e4962f7b07cb958ad0e8932e9ca67ee0c8e22fae6ea001e4ed00c5e286ea4fad92cf14b8c
z15ef4505ce7bdedecd598b6e3e26fb2282f5077d872681f7e55e976dd6083055dc9ba8f082fc92
zdf523acd3e83d47fd9ce20c503ddcc5e319b106d00492c9e2c093638f8589557ac4e709c7ffacc
za5a18e1ef44fca7c9fde822707e009a924100170b4c56d7abef98fd19b7ebb7f6b3697c3453f19
zc49518045b400917bc8caae80d9d532bcea1c19bcb988cb8b0687f834cb016ead590c5faaf9dec
z483e8e221a169ebcd68e007cbc6471e07de54ea3ef965167bd5f445c9b9be8cc8218d559427013
zded1a6872b1ed25828899a837c02115b286940bb9d28b523195b9dd93a6b99364a0fa4219abacc
za7545c9512b5db1d4b81ea7b4cd7f8c342f96a28dac2f60f63e5a84b372188d571d4e93e0ee9da
z45c169878d593a4b9fed4b26e76b332bde00b19a6a86f9cfac094bcf5918aff56a9f500645c220
z2f1dc2fcfd80ba3e7dff86d1666c9634313efc5a86d2175bfa1724f7ddbbbc6a2a65355f03eee5
z4ced01f9d16b70058792f9c9b4d4cdad5d86bdf90bcef3a895a2fd88041586345a1a741a8d166b
zd90e41a1b9592039de705c3f008ef46bfbbecba990a7b14f2f03cb4054f5affde4575069f3d4c5
zfa6383e198d470493aced45fd9ab0dc95273a1ceece4b1562fce2cb950f905dfb1543e7a861308
zcaec9ff91503972b4c896cff60600060dec5732b31965f322f482edd96c446eb7fd4844088f74e
z07b12f6f5a48750ee784ef7d2355b6fa11e04cae17688ec055b6155869597d13efb1522cad102b
zc85dce3a533500fefd2a2b4d25973500170836e8e0014a3f760bdb24356e9cde343adfd0e432b9
z3ec2fe8028e67b8b2f301881db63c79f272f38c6bbe044e3951cd373883396b778fe9a76ce2209
zd54bd6175c4e0b978f04ddd984140bc809d15c742786e9cd7bbb4879ab34f4c066dcd8592ab456
z51d5d9bd503c797fa6a314bda8226b727e9f359209b8f0f64104253db0c443a5a817b9bc427ce7
z86077c6c995538d68100acfcaa8cbf278fc15b7ec385eaeec39a5238bd887cd8234f95f06e7eb7
zed5dac04d13b4a49552c81cba1e4790296fcc1411395312659334b8ac6f568db14c529b1f74c69
z3a3fd50cda80df5a412f068df4c4ab16b3c0eaa25be9512033d185168ad5bb05de18dfddd62298
z018578d92e08dc6a185708c6580d7d497bc9adae7ad75384886304e9940ce7dfaea4c2529a03fc
z1c96ef5a3f03cf39f754cf1291b83008f50cf4b1d0ed9d8899c89fac5ea2d8ff411c281cbd548f
z789a99f2af523f1528ff0f83c5fc2d8ef55475a0657d2ade5599a8877f732f1f1a298d9e4caa34
z1f60113ade3782fda2ec901f1c88eaad0d62a5e7f588e23fefbd2f305912e267bd9ec2a22c4377
z923fee97f2f4c40e0778a04bc5168b6c01026a6585208e862ddba356d88e1f6ef039813204c7ea
z183957e67e1101739b99ee72202c28a012e53123228d28ddfbca0b7a71b577c4d9f4ebc2ba1e9f
z706a01e89d6ad23af84b8c57e9cc15569dac87d9a069a4b4302ea9cbd83bdc148116358b3a04c5
z36a27e35d5c3b54a31965a2748987cf388aa92e529b32a18274a50d91b9301eb1354b3777c90e0
z7403065397f37471d51daa1ac3f510f46946b72f59243534d3c20a116ceb94a4f2f74bc8899d32
z056b11c5c297127d74862182d148445f393bf5e89705d09084eddd52225d540a0f36b19cc20f85
ze75e01833c73cbcc381d0adeb790666239d6f70aeee7160b69002feba6d5d2232923abefac1e95
z1565d9833939b1ec4567b216f76bdc7b9e21e79c6d2ccebba7ce6acc7cd6f29ec158ad3cfa5eb5
z05cdd8508a8b250946211a15dfa1efb7e76ca56cbf2fe7df9d288f958cb6429ffdff8840e57691
z7cedf6deb09d50229e163c26969553301edf854c82517ba0d3d9cf546cb4745929be289b4bfd3f
z1d18b7e2bfa41ade0e2fd2a023ff536eec339d8215996108963d17d9352597abd8444e079ca576
zcaec5067ca7f8ceee5bc728dfe058a3e0c39cd5b472687ebed700695ea1e8371fd89c6c1a7863a
z6dfc4f8b694e7f2fb6cd6012d703a2004c676e8cdb728b5599a2e098689cd208b6c47d7def15e7
z88097d3c3ff178909223972bed189f9f6a54ac159059fc62284ab9474ef2240c7376fa2e9e938a
zbee15cdfbcc58fcce42af42f8784350cfe1595011ccff4fccb97a3ae38fec9b73167aecb902656
zc3d9676e8325684b2e8b6b8a1286d161dd8a54db42991b5413889194aba25f21eaef0a1a41496e
z0e90b0a946fb909f60692c078032f51a412d7617ee6630b159ba514d09942655f4b45962742f8e
zaa00ad61b8e96f11a632012ac81688fc96b2100e03feaa2ac61cfef59fd4358cc9a8f0c9d9ebd7
z956befba76eb76b9debd5035fd871483d895249698c74d31681b4a1f01085b51b0dc5b66f2933e
z81adecfc9328340db394406a0f146b163e008ef345fcb3a28053aa7fe1071895eec259faf5b721
z88f92a5114ed56fd293f1043022a040b73763bd9f4060053b47b84f528ad06f53ddc1fd9c7d4ba
z061051549cbc5d62f6b89d23d5a6a8182b27a52f33e41c249f9c987c87803ac4623520dca508c4
ze66bfb06d55e09c06a594408f0a8dbeacee8f37f90b70c90648a5ba481d2d08dbba607c205ac76
z8881b8249101a285a037bd7e6506e7bb0bb61151f5db893ea696eb837952ce9dc21c4937661d1f
z92576aa7978335a2b4382d151b086971f1720a7825deea42e2b54d67cd9bb462b6c916a47f33c2
z2477d324a6a82898479d73700dd0bede75ca8eeeaa9609c37f211ec88df45950f986a85eb16e6a
z6de186f1c494fc874416e048bfb9e30da7fbf01ce21ae903bc2c0775f5ee86a2db03c4de950429
zc660396271191cde463c3aebbf940ed2be5ae9dce4ac9a1d73538a60e902601363c08c518a21c2
z3731595d450216b4b024bf4d77f639444fc8156ca9bc436b9eddb88dc8040db7befb57cd85bb6d
z06442bfa6a2619ba17cd07de187b2f45cdad23529aa770c0dafbc70f1e49eeda8e084ae7617005
zbb4629dd367d94dbf2948f13b4f9d6f34724f96bad026b040e325f384a69e0b4552593b3b51fe7
zb479371d7ca55ef94e55f9c5fd3d2385259de742326ac9e77cf4632fe4bedba9eb246b7334d0c7
z7cdb11bb50eccde17c02850732633950211d12041b9a55a259332d108ba4cf0bf4d25ee4ae3053
z5b9f956e31f27620777437c1be8add692fcb9a17dc9be9c138bb1c4b23532c855d76c32b48d73d
z4868fdbffefd1cec466648aa5fd850a8f8ac3d044a5a10300182adc8345ff1d569641d27cde6a7
z3c482c61a2fb8cbe25dac59e1cb463f5dcddc04a86df13f31993e131c1df4ee7770388c743342b
z376c97bba09c3733dad5cdf3e83eb6c9936e4ac16bafd5fa8f1a10f8ccdb05b72f9c01db216549
zc2ae9a6e1e81711b47ed5d1dadc4bf31f6d2689ef682a4385f891c15eb920e1bfdd84c1d5c0f65
z46bb9ad3aa1119e70481bcf4d295c68db10c7f8ff6c95b5c915b8d084a55379133d9816fe48487
z431501f8382f9e05560206a43424093a5725b1b558b890254e197e90abff8265d16619df4c24e2
z604629dbbdb09b64db5f9f6cefd6deb5df93fe20bb948cf88d968e8d7e85affeff2ced57f055ed
z79f3ae9f4041e55af451303ff7f4a4eb0bc67c87647d0937c6af110a8744a8b43d1001d9cb8d48
zc93a7170f8c259563b8e783951cd31f8698ee3627453aaa8e4330413cae3ccfc4277172089b472
ze04f0d1f906715c6acdef2b9064f319f3eca11145fd30fba4426f4edf1a8c32e821656f62383a1
zeec53b104c83b4d4fd9c8dd32e0b5522fe06c37f52e6e886335bdee00df533439b42ba82371af3
z68462ca1280ffdecc80d4f0a19821878445d62f218c12ef2ed94dc0eb9ecf9265535c027991ffe
zd35b47e36108c622036fb2441ab1ad6c72bbd83bdf56789fa96ed136b20cac9125fd838a39f987
zce7cf7dc301bf57d4e69fd71aeb3fc5401d7265ce80619895501e57d396f4ba2c629e064738247
z6522a595763b650cc1b02d91b8073c2105b1dfe54835940488dc67a2d5810d748027b6c5bb41e8
zaf4f8a2567a6c8c4e7fc5fae4760b4af0445a12bdbf0bc74143cfd26d1f8583c9f75560222b048
zf62fa436f77a63657743137aef8b3d989e8de0e6b6c16f79f04baea310d11d84632edf2d641ed2
z572c6d4e22dbb31e3a34d58ee8112dd044c978b724bb08cc350ad14e433bb68cc4df134db2f278
zbcd2eb2d94f1943707164c179cb9db3144b173f151a41baa34377b43be64bb8e08f92611d51ec7
z8c43d616410efe974063c16444dd56eee967ccf278a8aa7b0170f4fad9cdc7bd3879bc0e9ae1ba
z2ed2247c6de6a920d75927b441de78d3227a37f8276b969283b7a965ece4cea197151634c523ee
z083c513c688789261b6b909acd083054fc88f5ec2b92a5703e4f53306b64ca8ea7f7c9e6eed04a
z6da3efca56fc943dff85f2e51bd81dee3d3fe60c4d904e82ca8bf7901b7d20d04a8364a4758b27
zc9059cd7e217dddedee1188fbe9f385ade093579ab457a237a709e30077e9ac4c3766edff4f62d
z99ee79d1ee08c9ccef952a323e03191df4ed1849cda6bdbabf8740e5c94398425c6388a90b4105
zd2f5b940d89ae03d9ca795fe48080636184141a2bef7c3b42b77b35e3df68c017b81893110919d
z2a298b8682924dc447ff907090b8091f5e2ea15cbd2071bf85bc745124312fc993b61b42ff3987
z074a22f03021c02d3bc08b5cd33bf71fd7c93ce410cd6e65a39e34e3aed76f667d208f8d71b7b5
z0f83e51f5bd59c7a7102dcd984b0648d6b299a11148edb12e13e6ec6de938ca8220f1273a4cbb9
zbcd07c719eff4db0543f129a72edf90d143164716a83eeba85be3272ff82ae182fdadde9e9eba6
zf6fa98bac0b0143acc5984c95c8a06f08c41601f0dc36f2f34d3d4f1c646b227874fa8623d2760
zd8a24e18ac5df6f5311e55057186be420f1eae29b9e17deceed933c78bed1643be52ef5878fe84
z5bb2b38110e32ac611fc788d5d5d06fec84815c5d3db8575b17f563d546fcff4824329f9145eba
zd8f132827c4bdd326f0331998bdcd81610b3de594e396fcdc75324e8b1d15cd0576af192df61dd
zc60fcf7cf2d521b347a76d5ea2bead196dcc2215c0de2be94a7363f23ed670548827beec081a5f
z02269421c5def2738a27d661f82ac7b649dc116782ce8696ab90e0c56b4d68f797ce5c26d3a1d2
z07bd667cdb6c2965ef99a3b7df06cebb024834e0f9d8d332c9276be82bac0efb5455cafc9a91d8
za47f41598a0177baf5fa55eaf7647f166e55d7fce5ba3e31426520c2e6b3586749e2ae86a13f45
z0898614f493274c31b95dbf4c0a515ad13fae00b3ad332e9b785e150a2ce7caa6c410be83393a1
zdf5d221ca44d1a5a1afab7dd825e94af6441823d695fb2959da1bc441be206769412690e99c469
z86d5001635003ed4b2edd1c91cbe7a733119c1b67b3e06832889d8c8a036ce5079d518f6b176ce
z1e43677085d0313714f82f8be3cae807bb324b914c30ca69e63db7416b0ce44c17650c694851ec
z007f094d638178c8dba7c881d0450c70ac508f21e6c3bb53e66e6d682852a2dfe716716423c948
z820d467013e30382f7b3bec8e555614efd94b06c42fb20650d6a1aef63959536a21a9351e66fd7
ze6a7fc427bd306d45d2b3e3bcd1e69ca41a15b54b40d63eb67d7f5f95702db810e369e5c21d9e5
z94ba9756709fd30694dc024c40d9357bac0e38c78c1f460f7f9d129a52def80d911914cc5a1b2d
z65a1a87fb2b3efec9b005f7d04054d1aa2030bf8b3c1355baac96737cecb2a9d0bc662005cc1a6
zb811dc8701784a1f9a77ebeb965d01b7c4fe7920063f2caccb74c466227f0e3efdbc3a9b966b3b
z235b7fd84b8e9b1d552db878d97fa2dc6c055429e38d2f022fba1bf14dedb521346e5f2bb1cc19
z57ad1d6b3320f8db57dac7d3442d42d100dfaaea314b05b9977669e0d2b03449af8f62d7856c6a
z5dcf1d3086736397a651e95e7c4f8c0198cc071b782c6c539e5a103847b358463020c91a7d96f9
z0f5dbc5261d1f1d4df305472c424659323b98e987bda2f800443b54020ceaec074035cbb8e69ea
z7ade0d30d73eeb5c3766c3f7e042e5a6c86301149d126f1abfa60b198044ea8333c9dcbee9cac5
z20edaead990b750fd9f1dbcd2fa70a702ea9d314e5f0472da4d7cc4bc6c85edf38e0d228e57921
z201335182129aada591b7c8482728a4ae70fa15eb9c3aaf3958ed7ed8aefae051f49336cdd7c92
z63d167c952c00670e163222bafdde3fa9a26fd496d5530babebc36814cff8f98fc7e08cbf01ee0
zbf3395e704bf8ade1363b3d46a901279de45b88f902006633edeffa1c1ea8b517a2ad569fadd76
zc6bcbb941daeb84de23b99f8a7228397ce057991f6ea896ce354616a27b21acc457624eadf60e2
z0f6a1982e24f5d26323687a8bae66adc0ca2b61183c0606a7c99aff3d2dd6b6a441801ef5357cd
z44a89feee2709d7fd94cd19a33e6111b7528d0b34a7db249dcb8f6c735589d1e56557a1cb12709
z5944f953c686a6539b6b6066b24ee958dcc84540e02a211b6823644264573988386f4d9be18598
z3749213117ea1cee9942dca73c6f14581fc60d5070b7863db08f986da771cfb4ddb4fa174f8a39
zdc58227b263afbf6e7d3e027eed4214199add80aaef59c8220f596b97f8f9cc384c3955ec82d6e
z7a83c15b4e65cbdeb1df953afb53bea6a71d0f27424a07ccf8488e84ad09310bd81103433286f1
zef266809206b21662c4d8052050f22c1e3c3a0bafb213a213e8f5eb885f92e79454643869f4462
z2428fdbc9cf0724877c9f6ab87b06775d7e12c171b5e1a617535c836aeabdf6fb0d35ae13a040a
z3ac5fa4a6bec0e8c9e948978c671d06a08aa80bcbd095415b5beab520a03a539e087c44f44559a
z11c2ca63c8ea45a84916ab9f79dc26bf91191f39b5745a8e323724edd9f4a74328ad39834d4f57
z08493ebffd64436d0bbcbe226b841338089d663c77f46e8f77f92a3a1b8064cefecff4cfed3d26
zeaaabb8f76ea83876f073b0571a355fafa94d48f36e030e6d131253c62a88172a31e4d8fe5164a
zfeaab1958a55f64c4290b6153e9b33f10e3238b2a61623adc3aad9737d1f66534aeeb36e9a8726
z1c2dedb8f3de21e0e0d34eb9d0578a56508c2334e0575e2a56929328dd86329708dc4994da8a8b
z7f503ad63edba534ed09299617d819ccd8a1ff385623e6974ae4c4a185c79b5fdf0899a8446154
z6bc32feb87d4ed8b79bcc7d765aba09e23e9cc2e18a776fc69e109ce8fa80ea069f19d0b6906eb
zdb282df2611259febb5acf3a2f5402a3c6c6ca85dd426dc13add60a3f876a81a5994f677872d29
zcbdc0a9939405096d4320b69d90bfaee6f6cc8fa3b2a1c4e430fe73463cbe0c002bdaba1c71269
z3fc61cc416e1d4c0cf6056cd200e71a109a74bc2d58728764639d78620c499a21b318486b0ac05
z139e1a036937ee0e842f6f990505e675228df9a303bb49d17cd2e435ecf33f7d9118bc2e2abb25
z3c1f06e163a429814767dd77dee1a2766e951899092634d81c6b171e68243232f555d458f6c182
z7a5ae1da2ca2eee25ca220f4e5669c03835a659b455ec0fdc15fe95bce7605a870ec29db1aa95f
z3eba52710a55160846c346dd842247e8a1ea9a86d5f60721aad1971abed4ee9965c3ef83b96ad6
zb262cc2251e4ef4245a64409d506ebc420d6a8e0bfa7c1a79101817e330301dfb127975a0e20be
zc6113cd8876c23751552447a76dcccb19a2a6bbdb3b5fe5c354b431db91066ff29e7ebacdbb43e
z293d249af16414e275ad1646c293654069ed4a013fd9e078f9ee8913873d321e2369fffb338d3d
z7d4b691ac3489f918d853f129b85f997d990fa6a955154516c73d16b118a9b656622fafc0aad1f
z94250138261377c64a97d2eb42113cbdcda36588c1a924010e5a2731207eb695c06c84d7a03dfc
z18fb7ec0d8482f2fc6b009c01c09ed9b3ab797f98fca87afa71a81bb93aea01c95217d90909c7d
z57818942abebfef153cc3bcce571a04748ce4edf00074f7e4df18aaffe02cd169e025b747fca49
zf6e099c6122d7e988f9687c4b772e3d8cfc1196137b7a9482b0614ecc6df4a4771989483b36b4b
z8fc37df522db2c2ca147e1486be6e97a0693e0e1b0f8c73400d4f761b174130fb6144f0bf022b2
z9700b2cb31e2eae3b54d058da0d6bc28ac14c618e18230ec25def6c2c4dbf0a2def6d146bcd264
z7d0c3e0670672dc728fe7703a9cf2b001ab87239f9ed87c87982a131648d14cf2c4290ad15092c
z27f62b165e1ea7c6094e141bf85adfd0691525f1aecaba33304bd43f2756ff96ad391a6af42543
zeda8eeaaf838e6ba1c3986ae215e421440d4f92b83035fb2bb0f13d557960176d8b3c9fd6e9967
z5d54d12b8ac80bf4bd1b473f658cb34f374300d95c73676654a082f84301bbdc40515c295ff826
z648b1c18d7d4ac10f7d969da3763ec7a937c0e63078f867a222ee4a488f1fbfbb83139a7cb8822
z9f8628f9a21a11a1437d43569331fb0b4a459eeb4b8f0aafa7cdf8f0986b752f0d78a00930107d
z705d195f4078031217bd1e82d2c277343cfa70eb097a3f1dacb9ad8161e574635e3f337ad59155
z31e02ac63b31fb4b606d092cb3c81d28e72f32e1142ce472d6bd6d85bfce47262cbb7b66a5bc35
z7f98f60dda1104bf6f66af19c43fa474bbee0175e96a515b4a9d661010639aff2a077ac2b0304b
z6dd3b6438e0cacde121d44043d37471ff940be3bd930325e6a1aa36e346c49ded59756a77d4888
z955ef2bed70e5e8ab93b86e4268e8df002b7258fdc391782206ab0a83d86402a99f55d19e839dd
z217a6b7665b538aaf0c8ed76b1089c30b5bd69cf0d7669f30dcfe89924d54ac1d5b1c092443a07
z796b260afcfdc915a0b18a512fe72d348ceecf833618d44d3a8e61b8739d14b2a135d7ff0bd2e5
z836f7b7775864a96c3ef5921dffecd5a5da9ea5832f71078f9e869409f47c624c94aff6e6a621b
z2a7e68d8196f6923b74d348d0508ff4a542e08a20c92e7d7b7ec4a9e1f65e17f7cd51f1a122f8f
zf77250ac511d981e518a31b3cef4963c7850ffeb2c87c42002e6b3c9716c401d4321edd5404884
zc807d553e5e32c5a030f00c3bb32319f48420c9b38589f3b8a4701c872c051aa75d02fdbfb9fdd
z30722602a658fe3c020444a6dc1e78390bfd9424b2e33c7093836bd39634d59be252720d08ab8a
z5ebbebeed8c1f2121ae9a43498504fa577e30c558ca0daa5fe8ca0377d52bdf99dcc02922a1f88
za6961d44db837bf8c766e6c8ba8eb6005fe8c49c12526ec54151371b7fe62863f257e960a758a6
z0be93053e111a549295391541aae7c9f5dc63de0cd86770d66b2acef08fffaafe89ccef78212b1
z3839ecf5a7f2c0b6b5e75056715fb08600af8b34c790887a3fbeed312f8cf405b7040be1574535
zb2051dc42ac9e2f4f474dfa4e69a113a7f39a8b26883daf8f891bfbee70aba2cb01ee23f6f8ce9
z1c57d273be5351eb571eff1baa9fc3d162a4c38e1b18d3a9effd3286b7474f42dceab2e8bd28c8
zd9c2fcdb6736fad21324e33ba74ae7cfb6f545c2b971e8813dce76f20b22051908815344dca455
zb8d6e8676fe084c995264ddc3a2f7d5d627fbbd02e612528e931ebd2237b2a631cb091243d3ca5
z698abfd603f720363b3900293b0c60f782c23dc0b7534ecf10effbff0e117cd6ae5d5c73fdd806
zafa352c23c75e5485e0f75042d2ed0ee2b8c038c2c3fb09813ea5e3201c142543e57964ed3cf88
z97f3d666f30963e7199c5b1ce3ab82832b5f7688d535272498e3717c3d1f48c58e52ea1526aef0
z3597cc4e34a63431c97a0c600b7509efea218f86eec2f0afa0c4df6091d2689f538bcdf9399003
z7cb6d2c00bb0e73ef70b50d5ab97c1206d76e6670b7cac3393c9ce0e130eb7186ae680f0810d8f
zb5c6f986f18ac465b43cf54338795877754002d56e5dc45d69e399d8aeac69e74866d91be23a56
z378c2a500f424765b18efbebbc80e0dd6e7a32b5c0159c6284eec911d6ee903f50cbdb47ff25b4
z58a13e50127d0af7d2150ac39b1d95a6d5b7538a39dd28aa909d8f27ba830c964675e93e9ae0f7
z809e76b436f0cdb34b699b9106498adfc2cf65f55539cbb3685f4dcca53efc6ecd12804ea61bce
zfdf1e4c34b1252269b6faeccc47536f0dd891587924359ae3b5575db4a42f257b49ea7bc6c5975
zbd62f0e72ea9f4fa9bea36669bad0389f5533f7762e578dc30a96dee9b48a2835d5cc8ffa45972
z6d0f31eb7350d834e9a0dad67b4c5c2b06f76be0c9aa1b49e45e486fc1e7f844083e5bd3942399
zb24c561f8daf6c3a3bb2bb503f453aa64f2fa3d0cac7aa9232052f6870c260e7d5d7a1eb821348
zf222c06fb8d0d14f25be923fdb70b0aa385d1e30de057db81c34c428f8d1e3c68aa3f2625fc8fa
zf8ea4982bcbf5ba0771d54ba93d6b440e3b70c0511f9a0a3097eb914b44ae31a5311c76e7b1cda
z8b580b47251b38d39bb6bf071bc42656b18d750b54403cb6c04e725c7208094981751421c6fbc4
zab104b336d5f29c63fa3160944578e5c2a69d61c66121355bdc4563f7ecb2862c54084b7f46759
z09c5b3e0204bbeaaa80fe68de9dcd77b1472e0493afcbaf36c4618c2d07b3bcdca33a423643ffc
z257496a3b7b9e85811edf1b4ce7decfdecec957bbce7bf0457a9d5c8efccf34efcad707f6db3a1
zb58b514f87a3bbfd140c164bbd1f4a8a8f82d1b57a319045de53bb617be28dc35b451e702d491b
z3e9f1163a5d2d12590ddd2780f2229d108051b83ba692e3650664553d5aaed94e073c76ed89cd6
z65581243424c840c0a15c329aee51b26be730ad7b0db9095344101463ba1ae1d9ac8b2d058a4ec
z2fcd3b46dd0662128448f47248578fb0060b111d9543a411247f05657bfb497799fe22ff3809b6
z11de6ecac1f8ca22fe1f472c3b8e91447745b28460dfd9b68c429a37eb340791e26166a16f4373
z07c333d8ee0ace24ef7327f2972502bcdc04896b3de4c5d8d12c9e75b83628c13ae08c70d9078a
z9f58f37981b2510002dd3f666b439525173969ca0341ca3a14ffbcdf737d7ea0019ba85e4711b5
zfbd80947f3f23cfaa7e0fc0b6918ef43fc139f7b1429f58ed23a209f9a38bf48af60c70b7fc629
z595270099b272e82eb74b40af47a186ea327d62e1b307af0504214ade0de8041c8bf73b96a1539
z694f3b3fe7b2ed6fa14897da24037fcbd934e2e97bb44d72291a12d4ba3802d39d713de7d3fc43
z2be8524cbe454730df2f74238f7718b975abf1e8c5c223926d6dda9917e0cda92bf697ba996b61
z95d41eafcc918f83421689e2e17ec5ee32f026e508caa53874fa2b44ed2f183a4ac0919e370c20
za82aefb84441f13229c8683a3ba595cdf21d94290ea16bb5ec360cbe4f9df91455dbee05737c91
zd4ef51308f45a1a47ee5b8cd2bf6949f2681e154d2673cf6c1fe6a70170daddae5703eb1a979ac
z58e505914209eb7046a18070098e52d5dc674ba03393284ec661a4e4a4f69689ad8bd3dca053f3
z4afb6aa008650b0a53d581213e3b88facef2cd1e3b725346a3df8af25466fbd4d6c056e0c9e000
zbd34c192c7adebbe2fa72762909ae12ed9bb02b69b0e923271f71a1eff486af367297f4158b1b8
z9b674cee18a36a84235698a92a99afebda0ef2eaed091a3142cfbc62fb6f55b14167b4c9877563
z18bebcdba2a1b427e8b0311eaec42cf9b7f4d4c08cb521b445f1e8a80c11a2f5c58b153f59cc7f
z6367d9d8d68caf696407ba5a6ad8fbc18a82a4e45601d42f44ba8e74752e1fc3a64b7914502fa2
z91d9b0803294ccf34f38b322ee941319f98e068227265e59693b258a3aaec128e1d74cba2bd301
zcd17cb0eee1b879afd06235be23db6118561686a2b63cb57caa98b27a081b9248322dc47356d60
z89a11a636a935f47c08be48286e24cc7c3f95c46c1f4c936cd77f454291ddd65f261dcf83a7b5d
z84339077d408da6bddeb8d15bf3b829e3b30052c5332cac94520eb31342cde0b5e8146149a267f
z5ad9e796f41a07997b3e028f547fce27486de9803eb5dbfedadd2288be6970c20ac451bc3b185b
z8586d982b0e6bc8b2a766ac6e9fbbd24d910c1604814ccb6ae1e8c57e357601c98f01105adaf51
zbf6729f1f929053d0f978da7081732292505ce12f1d99e326270770c9e6ae1c5e47d7e851aa4ad
z9701afbf3d04df48115e0bcef38022b239edcf801d61dc64ebe86adb67601dab18e8e290b0f3e4
z10aa03dce99301065e049b5b6830ee7a5ec621baae9f8756db4b8d1d814d38a37c4e27ca99ada9
z95f7e0ac9a128a00f2ab02f669d64621cc8ec15028ac28d0f1f5c2c1927702e34d1e9afe3d0b38
z29723c834f5b39a04724a607818d42eaeceff1c008d684b0a0cde447eaadf47e56e4749084504e
zf5b46bf9a68721edf0f0d985b67e2b52705838fe3c0a0acb636961333d0192036408aa08c3bdb4
za652ae2bacf45da8b35ba9c65796ccbd14515611ac18ba114a90fe8e272973801da3dd8887705c
z7d6b9fba468e6ec7d0d41f0d1af31cbb1f023df06525b23f74784f9932d75cd2f348929d5fd946
zac85cd667e4712669bf94519e82c93779143da873422d3c1279f57d3cd541bf9cf9c5e2824fe01
z37027f743e54487c5b0c4ba64bc20651e5cdebe20562d102113aa40e1d42b170ca59e2c5c75f08
zc143d40c8a934188dc426896fa01f2a056e9a388fa74a043abefe3753187ee74f84e96e5169e35
z4d88f99ca988c361e1616854b3aa610442d14a7ecb1845213f9e88fa6206874e70de9a0539e620
z0ecf29636bfca9a7eb5efbc43a62bb530f62c3d88d8273e75063804487cf7594881abed96be37a
z58b308d22e4545dc020d8ad868bed78ae544a34742281639f59f376ad73502523c24b284ca1f95
z1bfc4e46d8c76dfdab81c79c1ded5d86b37729d02ac7927d67f0433691657134fdb1ab759f3bc2
zd850615703b67015f2b02a70a2bd2d93d4460bb35d6239cfe2b33f298a76007e225be6b5fcb129
z12aae6e5e60dd4487e469466dbad1fff6aaf4ffdea58f3f6da75d99961e5dd15bd3a96f0500820
z80628962c9aeea965947cba340010b42719e43517800983db6b1f3b928b1793b9f952fb1faf0b7
ze9330622e8163a97675e0fd20fb00cfb8f6cc332c7d0431c9a490d3b477c44dcb936526220dca1
z905e75ff69f2750c6fc738d47f39695df5e6127180c14882bed03e60bd952afe82feba54a5e3e4
z6953de610e5a4e55b81ac683728006e401210b011cf375212734e51a04d2fb45a7d26c904443fc
z94b854bd8be145c90e6f01c81b7fbafd979f75b4ca2bcaf916d85e580dec177cccc34c2fcd7683
z9abc33c8613bc1d2cac4364a676bd23689323ddc5fcb52d766290fcddd6e9e3142879603b262f5
z99fcac812492431a2b4e1e8ec1957e3fd7cc980d703d53284121b54b615b111414459c3f926bbd
z2b538da8b2e6841e1b30fe543bde8ab78cfb594845bec17babf1ab55266d8fdec7f3d52d2753a5
zc011864b857e6b3d27afcb451f59df66e559164945d4e6d3df8f333de372623024784d47f0d6a4
zaadaf7093a3db93334ec10b454cc53387c0000557b2b5db8550b3eb8ec4da403284cf25f908c3c
ze089f8f0509c4f943e27c0dcaad02d8c85e6324b5e14efb7391279659fcb8909f1cdc12ebd2adc
z31862814ec023e94b58a3d55e163029e75484d0faf489cce92a99ded90d93fa2e8d53265617806
za381812deec18c90aada869a674c7a242c47e52bb94fb1ecfc07de0002527a5104c940c5d2e3c8
zc0681d5bcade79ebbe593db71cd890211f61b4a51ae453731466c7070c0ec5197cfaa357ef170e
z6dbeda4bfff2fbd81b7706cd3fdbf41ab7dcedfea5d64e3ec6e744b2c18fd68b5eb25b38e22b0a
z8fbe70ceec7eccbec447af8380a1c14b2d394495b1a132ceb98267b65eca92c9ff1203748907f7
z78dbc92d6b138bc8195da0d29d1c6fbaa06c7fbb40c6ba2337c80871e081006de943e85b697579
z90e4f2bfef82b9e2eaf0e8b2cbaf95a8d42fc94d15bbda44a545badda0c863f65bada6b21fb8dd
z8d14989be9e9df48b2540bd54825778ba0f62a1a263194fe108bb361e94264039f675a0e380f96
zc13fcd34d370370d7212ca62cabfb2bfdbd94797c0e357ac27418b3631a08ac687ef0e486ee07e
z8fadd5cd60211e5905917ade30bdab4138a02b3b87f29eb1bf91f9cad1a95fd2bf915d1a96445a
z07edef6dd77e0b2f43e8ffb4c8ee676b724374d364839985fe42477bb4ff078b21140a674a51d4
zb5fb1f73d1f58e2d83417c0451828e260791e4fc01894fd335cc65d3e9e25333a35147aafdb339
z65f7cdffab7a7e5ef4b8c026d892de3b4d76d82be5ff1d1682e0dcab427b5a6ec2d5b245a9defe
zd361cf539ece18e8bc46550ee541d0497e1977cf39c9583b76ad758245636a748fb81fb7d16f8a
zfe8fe8e0dea628f1198fdf5470e1729afc1989f7566c55e60b28b7d2b8ebe3b470faf6e13af111
zd8ae0037b5b3d772ee73003ac1b3eec9214f45042798cb3f066c0b975dc0363826f715c1836d4a
za5fc507ad0b392feba8b3111477e7525b5fc84b95f2a93ebf6325918d3fd9accd924ececa3ab6a
zc3202bb1296d3a00bce35c5ea7c052c2595ced27725d3daab1f0b453f7b2d51298572842b998bc
z306dc2c86e4b455d39641b803875d662f2086e3d212f4c56516b8780c424f08f3feadc5c375c03
z7f547e556323a0aa98887a6f211344483189919f97ded351381d7733c1fad9e65c5cbc65a38897
z391a9c857bfcb335de58ee941960202052b3f740d439738a01e12d06347d96f111541ec040ed4a
zedfc3d92d8b9bebc072b13dded1994ece28bec35cf76732c33a55551bed21b0f44f8e75d1dd6ff
z69c452a54c0b3a8e1786adeb0bc54d88444be9b23a3faabe252a0d0f6f4aa1d572c23246d8c6fe
z4b83416d3ec12f0770fae89fc2c133af51f32caed21c42ebdbd14bae5f73784f1f4c0b07e5195d
z10407c51dcbe9584951ece14daee9f63417f2d0675acb6bf801415d32e317050c94a4310ec0945
z6e43fae523ca0b729024cc117465e57622b1d8a896e930f0c1ad5fbeca9e2f1029cc989e0bdcbe
z64081ffffcc9271adf4a83d6d5fe547a32a35195e1f0f1f3a4c3be739482dacda8bec9a62c8087
zcad3115d292e5c32278713e89b309c0282286a2724b756aa986660872bcaefd8339b144292ac99
zb5971de004d4a21b3f2fd72ff728bce3ce535746857daeb1d192ea64c3ef083fea68e1db94973c
zdf89f501c1f0788a664dba9ab0d36144b087767a4cc0b767bc8f956d1e9f671ce1b15de2396318
z59008226ac3d441b09b9873c1025b4fb8b8f65d9ccc23e8f09a26b5032c0ec8999e09ede13353d
zbdf906e5b203bf85fc634b92b1afabb04f1a73d9c0a153d4b5a58d182fc3459d19ecbd44ce2d0f
z40b63db96cd3f441a12aeeba6c62522a0a8b4034d094ee396d0f198e4cd367a892fbaf67adb287
ze0ae53f7d07f597fbb76492636dbfbb61860431f28cb472f7388d9144c74768c5832dc9033595e
zb25aa5de91014749945993bd624d25f0912f3c327f9e048694aeb33772d79bb45469273f77ea1c
z1f49690ee9c1dff4ae0ee667a3169beaef2cff2d4e5c0426b94d1cc3aa8977e18f2ba796b4c0b0
z6bfb2bb87e3c556d5574dd44eb5a0eecfb41348be40391ce5017396b009413f0030b2c6211312b
z44a260d6ac3fe0849cc7eba98eaa162965a9808297099d135f2787363390eab3a9fe5e24e631a7
zc2f4377e5d9e5b6fdd5ca6c633b61a908809fd3381d7a0f91bd82bb43ed53c35b4c85362d8184f
z773fc5c7daa5b0f35645d51356c979d7927efc44271344bfba3fe20f99e12a4e238d7f76538a92
z41693a77c52134662fe9af7091aafb544e1816126b7a92fd931dc81e238f969ac022eebe78dbce
z8f950446aa365ab8ebbb3143f207d9a9ab6fac43701815228d547e734519b04b20c41eeadc1e99
zf15b584a99468569939bcf0b4503c3d5157fdedaead65959d161f64eecf27fdff136c445983c9d
ze96d5ab9836b32840fff6446a22f06ec4313fec5729834ea66a82f3bb3f6fb2aa58856e5efce27
z9a409e0f8cf0d0d9b224505e3594609d57b76ac08a83116ef3657c692ec581abf19c8fac9c0814
z290df945c3486b90f672cba84d4d2de85a1ff82505f04965116faf2863798923cc7b8fcfdadac5
zeb010e2cc5f618663b35a82e9fbc10cc722643d16da9613efecdb57a0cb1f88e202f84572b93e5
z661abd87c9908cf1f059df903ef60709707964c7ccfb88dafaf595fe208cbb48b901a798fdb72b
za3366dfdc5eb3d030d747646d88ddd7091cf4f703375660cf890eb5730fb82ca4e659a1a45253c
zb578b173b9993fab81b6e385e1537f434cf69a0182bd9e1e2b2ffb915a7e322effdfded4285034
zf3944c9a89eae33c9060fa24c7d433198a2fee214dbf917862c6cb929189ea59768ed935ee1c08
z7f8bd81a0a74f13a7f23db43cdd13a7ab89764280d929582843ebd7254de5301894d3ce29c5c2e
zd1b6de0f418c87162748ebfafb03efcd36e4018dbe3d931ba8d5a78ec66cffc25f8c052fb08098
zb6d2afaac71d6a2be759257781116d508a1dd6abce8bf0e92f977dc571ffd9aabd16928baa1f99
z8a8949e9231937163af4f2262c065d15d198c8560aad3cfa35eaab4b8bd67d3a74bbcac5190f20
z1f1bbbbdea13d354abef98d1a3e29c6365b0b3d01eaf4eb8ec6c36b4522c8549f6a789ada1ef30
zdf01cdd48df643d6c56ce9b75c8872135cf446390b0a07e578738c5645dc54216a75d5fc79d843
z054bd9bcd316808b1a809aa881a0d558a89448ba5339381a889a9dcc62d95138809bc0b7781c8d
zb02b1749484b4931c817975cb2c6c61708e1387f20dc5e3f4286239736619047957d9911bef424
z292aef20a97c92ca1646e9379179873a2c9cafc6850b2370761f4b9e98bb5799080b5d69c6ed6c
ze28c8a44a1dbbbaaaf7e1ab3030e7841ea3d196fd3d2962a070a181e338f181e21f65808ca4ad4
z88f0f2974bd9e4df0b411b9275399cdf156502ad05af6c4770d9e73c68b3175b9d5283f2beba09
zc96e8029b39219554d7bba0c85308ab31c8d12df2572b51813c014aa31133186d425483dbdddbe
zb17f160a160f3afb2725a08987fcdaaf49eac417e2cebc4ee520aac9bb45a8f765375a72364fd5
zeb9cb709c1bf684d09776f8f739b06128b2275aab8e8ed6ccec5285d783b6ddf7ebdddbfd386cf
zdcbc9a3322593a98eca1ad4be0657e3a1fa1462477c431aca356e3a110f2b78dd532a8b682f500
z3db3ef3d14e17e2f79eb3be0aee22e2fa7ecfc062cea9a9f483111620264c487a2b4777e224fb6
z0ba025a2437e5face3108170e671086745bb048d1a9662102e988a3da48f42188610ae0a48b5fb
z6d6d8bfc5e7adf5329d7b52c2de3ed48c40167b5ec077ec216716e6e24008393baa56108db9c26
zf033416e683863ffce8d332eb7f2507ce17838454266484bf0da0d191b879d87f80cf71c21c6a5
zff07132940133306e26bab981340699f47949b2daddf45e94f3d32c721da94e1f1ba87662ca07b
zd9e443f17ccf0281cb6bfe8f15ec4a18f8c3e0f3e3e0b588f78842f703c73c562320f4e41d7cfb
zdbf1a37be2c1860ba789f84688c8dcbdad1e7701bd76c17cdd096e9a6102254798a2db20fd542d
zba8f116ccde229ecd9cc2ebae208f2185e390e1940abecdc0c904ab835b189bbc7ba1ac4e16615
zf3afca45b24b9c469e3f29682d4f8c54e5252dc2d1bbe7431e6aca2a124167e3001d6640d39877
z4e558c1b3b675e8abea7387da4dd2f42013553e2038d87550bfc869685bdc241227f2293359911
z36c1b164a6b2e979843c18ce0474164c0a6d94b6711fcfd15c86f3cb9bfa27959bbb29d0dd8d28
z1421d191712e9cb8aadf00b68fc756ddbe18516ef3277ffab7c7ff6c6569a04f5643f8ee699a4d
z28c56927ac8c29eca136547d9dbc9ec30bc930db19e1ad74022ec9adc40655bac29b5d7bf56df1
zf08b15d701a28a4f8c45619c6a8892c47dc82e30f3d39404f880291fcb34ab58450acd99e59c7d
za47d75f8cebcd980705189153aba81379c64cdae5234ff42395ebf51601e2770da0fbc3ae53cdb
z937de360b69e8881372cb281c361c4fe6728a953d315971923f91926427819618e7c0ea2df26eb
zb75f60223bd1a34322577f67a7bf0cd6ba68d8def8e47b5a0d1c58d90541032a8675f7ffd316c5
zc1bc49869d49f3aaa03e5bf5155f2344499692ad30a32f8a0c83d8907687c2368e72fd9ba631b5
zf58af96d6b7fe7ac10eb57c4f755877015e28286231deb30eaa91f99e8ba107608c08a92345d49
z4f449c893b0adf3c96d2877a93de0a03ac3c66404b07a9b1a2d503a8d02fe3b146edebc61fdb3c
z72020bc32534aec0a08db3e9645eb394bbc4664bb2946b206d9880b683034ce059856279a883d4
z53e00cc58876dec9b6757656112f3cf5869913478a71a3610c25b91c279be700b1ce9395f99c6b
ze2e43e634f1919b586d7a26fb099c6491b55d3738b292e5550d78b7434da5db7baefcd5f012aba
zbbfda04c1c6d9b0778e6cb7ab54c4c17e8247a4f94603812170b37c927ffc7491756ec2ee8b421
ze0f8e85b5efe27a1be41bceb7148dd3584d1cb0f4491149795f5c0169db5c5f653ac799d34fceb
z36728ba79556da1b76d46bebb6c8a1898efd064ad4384c561554b052f84de526811bf082c2665c
z4d72cbb135c9b834924c902f01141c425f088f81e44d92f67df50ff89cd6c796857c2106ef9c6d
z973c8fdb679928bc7ba562781c0431fc91e89c882c3eb64ceeae46a19a78015eb72f938aa3728c
zb15670ccede439fbc69d211c42ce68da482ca81ce86840258a6ba35f094ee391310f9783105300
zcb67c89a05c807ab623ad915407426330e4b5c948a0c64bd440638845c225219d8aa2de5d32338
ze85a5e8ad14774d436a838236d614dab50a410e8b3c4c633dc3a7d45222d72461f259d816331fc
z57b7251a75260167504f779c54d11c7df02cdc8b17d6d46a28d23b8da21a310c711748713f356f
z9feebd3ca3f4efb38265bbfed0465eb232d4500465f60bead4ae61b2c66b8984ba2041ae40026b
zd93ba41e692b88dd0ce7f4824479efdbc33204e09a7ee430b15da657b53daf2d6fd7e2e92b2eee
zc410521cda99a94d43ef7f7cb87562c07c5c546760404f2190d6b329b86dffd7f4f914ac316ccf
zc47914fe02e10f0422637ed3def2b4d8e91e09bc434bb35f967d11cd892c78ffbd0404f25da23e
z706ba9cefc1ccf7c032888a87cf25d4f91ac7a0471f7c3208077f2ae21c2a75c848fe6554ffe20
zf695b61f43675ae9e95bbc86b020d0114076b26ab755f6ecc7d59f0db82bb8a47294df0d5bb926
z3df28a3d8fa782d660b1171b75eaee77985daedb47e8f7e4062a31f59d9e5c05bd91355baf97ba
z0d015d486f56be62c0f78110421e88e078d4387d9103421ac7031097ae0ee199f8f4dc89e97d3e
z885a9491348c176624856df6f7bf8095ee0c771edfd5c5bd83f37d2a79594be335eba28d342dcb
z94d1ec279f1a4d47a34948108afe4c9e2dbfd679ea2c797b9c18c4aa9e2bdc8d1db88338e4788d
zb859235119bdb8f38bae6c90c5845ce4fa2b5b978f7de00bbc2cda12514b2c175692287274e754
zab534ad25fd4425691c91f4e2df17811ef9e43c340904d30315a8f0923e87832099bb15a015c8e
z7c75d57ad5e8ffaafdb5661322fc3901db320ad9dc2da58f7b0a150c51927672da7ad890796382
z63887a71c76dd3aae3766291e0083b8fbe9ea164065fbfbca2bb230ce6f832d58d3a4b160c58ac
z9c78195d8b165b064905d5a6a8266108e9631d00ddaafbafea3faeb1d8935a87f7f395adef5491
z2e5505d79e388b99caf72a89631586e67e9cc2e9c90004a174e1edd8c14811ccf3ac8aa99f1d85
ze63c30ddf42f990cc0561c5f514491189d7f976eea98de4b4e0e7f4498ff2070b0d52c17257ab8
z314e0dd0e0a75503f3acfe560ea502dbafd8d9247d8937427e4eaabb1f75cb65ad4bf1751a4db5
z36dd3b31ec1527442457fe1a0ec8561ad96de5ab56ad2e81f87298e9001ad147250b458b340703
zae5fa0f8397289e1370b67225f3754b2bfbd54442ae961ba79923467336babe8d699c9f71295b3
zeb419a8fd058ccdea4d6ed2f6d983587c35c412dde84885644413711b8a10915ae9621823f1d66
z140bcd18ad27ad88951e34719016ba4488e56f99d0e6ee4d32a1861d8df94041c2840dd2dae9a9
z9f86a3699526a59adc486b0ea439082e0733f7c4d495660f91938e6e3e6aed6c48efd409fa16b8
z6cadd75776a292da84a50cc3bbdecb176a5ca25a110e37e1253b5eefdba0f972de073c8fa5c5a3
z3a6eb9904f8ea453af7f9bf7d4c7a06fe23ea3551c01a08ef712180c6ef786ebdcacbea65f5ee3
ze85564027f5f61d658bdecdbb01d4ce0068e73b0e9fd8f7a2a89db5f020d78ed49dbab04299838
z6e9f8733b362f279ff01e5d1d69d1cd07f06077f6cc8a95b853859edc79a95e561514648d0e687
z830dc3852d2e769f5ddeb743806e41a35ad9607f31fd263c014aa0af7884bd60668ae9494ce8f7
z19da1447d5e7f28208b6e38d1ae4382568065595af5cab5410260546eea88e231cf5ed644a05dc
z17f21b68c04f14fb7fe1a6c27ae0aa1af454ce5c81331aae42746cfab1db8dffb1569cd510128c
zdffa3e9e1ea28a0a972e4a0adccba289c8b708f420681ece0344f4cf85970c494e3dd3a951a934
z449bf2b3512752628d97111f28f230bebaa59301d4becb1f30c643d695913beb4d332eacd3f03e
z91652c9bc0e92a2423074e476dc7de6bca15856ea5117a0f8820b95fbac74a3f59299ccba05247
zf98952affd610efeb174f3ed37bcb28cdc7f7dc3cce3ae0e35d754b39b44bb10a4fd67e92a0cea
zfb2960eec6c0d080b7a46afd3912d2b5adfd45e4137042e5d8e222471dc5f1357335c12799ccf6
zc7d162a8727d84dc951dd8b0b35e2934b4fddf2d4553bce501f7d20965c30ce2ae3cfce6d9fec0
zb556c47e0de33c1ec284533829bd04e0ccdc05b12452d589a76d394c3c394a725e5ed689668370
z8471935cb9b4ac80355b7cb155f941b2ff871811e2676928d79c47a005688e789711df46662428
z0c7f50d48cb93aab9bb5e8dc5f6c9e0429bce59b99231c76cfa628254185b11e1812d0f2dc9b6a
z467034aa32c6804598d08d5ae682081ffd52e1ec7a1106a0da4202a6ad3a957caf27b59d8f9ca1
z04356b7eeef0c738a41ec8cb7640811d877a7cc6c09df4b39f7920a9137bf393469121340cbb86
z6fcf237118e005dda1edb903a6f698e9d1e47013d00449938635d03b89616a60748da164a0a51e
z5148cb547f1bd8da531c4158ec300f64c37069db15b6a0669857adad32e61a41c3e45def85b01f
z182397c2efd4ec343a8826b63f17053a328b76f1ba402c61edc2f6a02395d472a0c4e55c769bd8
zf8103c3b9dc9866cb0c925a5fb580b1531d802c92f0ce0e934d9bc9b8a32effe3ccbe44198efa8
z34edb370dd369745f31b87d9318ea9524a686efd5cbb7bd8a0325ee3bf7213b372688148227cab
z31beaeb5fa1273624e59173af0002aaf900191493030386176ccefd19c8e89fe80473271af9082
z5dbf9205c13d2b01b8395a81caa1eeb05fe3f8c218e2917727165e943a9568402bcc65d50d8e37
z2012319ee5e53cb73f5909af8ca41f136a83b012684cc72b7fee36d30260b9652ea3122b7c653f
zc78f75827c2043458f5ce563b995e111cd4105326ab3b31dbb2fb2e88aac40509fb552380fa1cc
z046a96373a038200080b88c7bb7dc09f6869a993ddf4acb9bbe30e032010a7e8d44e00d3f71e4d
zb620e1cec6e22ec2d9e8f9160b75abc929aadff8cc55ae43c714afdf823cdc0c86cbd5b2c85b0b
z2ca3ba190b300d745700c36efb25160e573704ea0a7593c1edd8fda405d1cb5eae750dab66819c
z379d7d068e11bdf6b2f63ba1a5c0b69a5246a025a97215220a44c65b47b1f03a466083e1163bef
zf0f2a1d9f9f38fb28df1b67c133f636b5f8fc2f1e6fe0a3ed435b0411aaf36496bbb4d29ce99e1
z69b3169641b1a3321742aff77ec7346cc0bb1f2eba4a1523530afdf965d213975cfed074f73e94
z0fd279c4f89bb6c8b25fd59a7f11d542187f7fb185375361f56cc7e01db411deac654b5163f474
zf710d29c1d291192d3af1a33e347607f93d2ca53046cd7f654fa7b12967ccaa02b4b9502d83208
z74be3dae995c675ce03df0a8d31dcba4232861c08f9a324e159c41e59d11578d367d071ceb2cbb
z02728f3902b888757ac9af071e04bff4af84aef69d98dd13ba5c53be1a533f302455fdf97fe40c
z6e2143989b06895ab8de6ee505e8056d1a206115b4b59f43c5afc139cf24fb40ae81159a2d116a
z8b0d587848297dfbd1410360667ceba8e5d0749986c8873fae7b05dcdf79502e456be615b2bdad
z333fd4dfb4f6dbac4f41e9bf5920e6081b94f6310d5c10fd60d41e35e4727d49f4c2a3fbe51533
zfb874f89b55efa4e79fe78283b9f491cdfe64cbda99256b6823e1af7f3b559c70a07cdcf43d786
z609b1f69d571721c860c525f8050eb93cf4fcd669d4e968edb76065a9d01eb81ec19715217826b
zbb1b9924483a22e0ef8cf43577cb15afbc5f2445a5606978b18f0f966a96c156956f8b850af1d4
za38065261213666813f4de548fa955caec9009db919184af0f216dc305adb3338cf9da8a785252
zc8281f7c5588fe73d1f08569b2106fa62ccf00af6a9a9bdaaac40ebb15e1791805b583b75b765d
zcda3c27805c56b159a2598bec4b116522f04bd545e60c9bf70da3959c8ba90d5f5d1b2d4d34839
zb05fd54492b14e52a391a85e6fbd1df832b9ed42e9010e100dc596ec3796d89654806d43cb7883
z78009f991cc07e0af19fb1a889c0bce1c60a0f27e4e4a7db56c526f4400a8f2930b611dd6041f3
zc51a44c1859e723a0d770169095f0b85be6525db34ab2ef1f9297d969b8df6cfe0eeda14bb4f0f
zd00aad2eb261286da977936d5d45594d1e42232be480f61ba2b792648198a1b3782c8174f839a2
z58fc52761e109ee1fc3d7b6e5b4b88a11c6dddea73b3bc5b106f0cc03d465d28eb92a264df9786
zfa5ee389b9d769c2f480a5acfa3bad7695ce245edb29f0c46da03717cb996946b5e1aba8cf35a1
zc4c07b09769c146af919b04de36c9c6ba2f95e3e2a52a1b484ffb5ff1809087dba8f37752bfb14
z28ecedb8ba8c28b33683a0954183ee9567600890055bde872c036ffdeb08c9b2ce21a41a39ebd0
z4594e0e48d52e93cb03c74f9aa6c8f3c9590924fa06e3bc01fece98c14d876144ada4c4a50745b
zf8960c9ea43927c1ccd363a1e10708f6f426be347bf02e62f3c63db8ce7c5511553152fa29047d
z4c992edb5b7e8b2aebf35f719733af3146543b984b18b38eade26a30f6ed5a4635e2d01f78d73c
z3b60b56b5a5a31bbc1a84eb0e7b0516d6cd8e7e60ba95b56d15b6b685332a114d04de928a2bea7
z70b5986cccd505dc35374f0ddfe2dd680aac8f244c08dad264901353ad1990fda156f3c3d0154a
za077759394da3c7bff6763bcd41d9a350a03a06e386e407737630c80ab76a41220226fe20388e8
z71d1dede65f37be5b185c0887493b6d3360be42131d05215d462e5103141aeae9c204da02517f4
z466219be59a3081b3ba63cacadd11150b3015b8c3cc7b1fcf9f2d2bd71cc6fb08bae7272500c4d
z72aa6703810adea18014e553892f6d85480d97cb3cd695ad983b930b4232c5d48e95f3ebe5b26d
z2d29d320eb5bcf1c6bfcb9ad57eaf598e1dd00a899a43360f31dd9dac2c741474844064029570b
zda8e78c73b734d9c8b367c73e9773c3785f0a4debb9bd2fef018ec2f767fc27730da1ca56c00c3
zd9c84c0784f4feceb07d4868b09eb193d78c8bad984ad9bbd4f76253b0c02279e08df297af98c5
z6d677bb266018d036bb199884d2041616b7ff777bc24850778f1a0348247a97c67dec567539652
z39445c1de4dffc4e3acd10bc4d9467c307b924cfb7371bedf93dfd42dd3e8678d30f8db1f7f037
zd3eb84195f692ee4e89f455099494b324a8d1cce1f795565461e7de73ccbb58dd4cc97acad846b
z1045993d791fa9f354bade970c62f7ac09dcdf7ebbc0e9e1d38c594a0e3c6f6b17695679b79bb7
z8c9eae9467163e51125dfb4d1b00d58ce9ddccfbabb5169b44cd3a03aa9172e7b8e33357200dc2
z9e76ceb83f390589a33fb9beede54ee8e86ce2123b42baf0adfdf77b4f6a095a7ace452bb770c4
z32264e238378e374b6a91607bdff13626f60ba93de275c7b727c2162117f230a083ee9ae123db0
z912088130725c0ee842c2d1b77f82e8cbef501ec4b3404ba34df33da0f9a75c9c4991aa988c112
ze15f02ddb8a8226b3f56e8de613cb16a7156aa56e1e96de5c6f29f18eb6fe9eb5bd529af5249d7
z8e558663fb23420e9e1883fa83fbde28659865e4337573a7599da711a8f1ff7e3c527c7c711f49
ze5d2141e1e76d1b2f365a521222fe6e72e35b45e0639b66c45803cc2b7b3b4641181af31c7c6cd
zd4c5984d5af81750cc95dee4a24d3e9185beda94391d140bf29105ac1d549827ebbf6269cfd073
zb77f242d92ec4f4acaa30fd99c8e974005b20153e1c8c25fbfeab365a884a40e49bbaaf5ca8ea2
zd1188dfe907a7b8ea38603ce2cbb7d3ef59df368d6c0311f1faf22af0cc44af1daea6b290a780a
z59b756dfde6982701d02f03c55d02092cf1ff61d51a1e14785142a30c1276f9c07be2e172c3ed5
z1b475f2b917a1e2dec36402c303874f3bd9d294a0f0f57b56c5956a7b962415672c62aa953e9d2
z4608b2b79244893d867782359842cf8c3f6c42c129bf38010d27bdcf2fad5a14ba94372945fc5d
z21a960961d7db70f09ce2c1cf3d9119533eb1ac709be15af399b55d708b51cd412588970ed4ec4
z693f6f3ff77c7bf1deddb656450115d433263f8df019facf34d51b612a1754795ef64ab0c1c47b
z579460bd6b47d9c5d2522988dc6b14ee6531a432a1f71943e0a8626b77b871d0d06189c84670aa
zb22685bf4bbc6b1d2dad0bb72b8c7366eef822f8ee1e20ed68b0a2c0516b860f01bd28676e38a9
zefc65e784ea6049785e0c0289b5229dd30b7c684a7648674704df354e34e604bd5064882ccb38e
z9b9c7e0a6f83a4cedde0287cf95322b3d8a2fd89aa3b01e523cd756cf505ae6b976228e0b2b7f7
z6a2991f50e1736a1196ffa2db6195c9b6a8e05db1829f52f3dc47fe6ec11710640302c902e1b21
zbf4a93874bd0d6aa1778210ea2f90e0672e33c3d28df0c341abbc2f244761f649cec8bbc97bffd
za4043165d1a1d6aafdfc9188caa72e6c051b1fda149775f3722059736ab62de04baf09b854c75e
zda90a1d41aed6a1f30bb65e21714ed4050f59550d6729729fcfb5d85064cc4dce79a1f129c4f70
z05b1811a3a764b75805673fe7997496c95b74a4eacb20d9dc51c29daf070bca37ebe5c733ba670
za09152503cc779fbbc379b931278bed2dce4c1fd2ca0f1318d04306e40bb10a64cd54f0e07b66a
z212977936e663c70127708123e8b2c2a6f6fc7cbd348dac3a8957775296a025d3fa86688926624
z3bd4350ccb1e5d450b1b0ec12eabe9ea6797a6c0daca0fa2e917061693c7a85143097e3d8ba858
z390daf32107cd046cc8125cd56c094a13f1bec3f3951fe990392b4d095f7c46935b282c92dfd17
z4bbb233b838bf309f8e45c7b2386ca6f8881220f027e4c4fe5f765808a18b31ff36e655b2240de
z6161ebb029b0da1ad0af309cb4cf7712360e04f1ac0f4e0c959441599df9be846ecb6064dc3f42
z4ce0eb42a159ba686bcd19f36ef0507d07b1d655892e52ffff38a283fabb792c3c233e4818e641
zf3ac3257ef86eadb967309683b89ef2ca782db452d706a0f6cb8f19d23e2d3fe762a4913068d99
z136458235898f0837a952bb4e3d6e2baa45f57eeda5a36137d40f05cf62bd2f27d6a487169317e
z432b7ae46638ad7510a4ebbb18aa6c2a49f68d810fcb99710ea7988375c6bfac5c349d17826327
z6c2c8570be28f3e950332242770ca8264d877154326b27ffbc1311eed4feee488e1d963d936d34
z37df54fe2afdaf9c444550aed59236631a27f53b0d5250453f6ffca92277c571fe95e68d9acd2f
zd3e4b87db912c8f74c1ea007b4709f9cd05200b0a198b1f53cc048310ba7299e22247f7e8b077d
z6f8e3a366920a17e9d726535bb273a3e0fc4ca37bc7ed5e470e1713193fa537a3856b59a037ffb
z490dbe7164ce7b9837e1e537ad2a828ca98b3ede119dbe8653b870595f5ccf233b5ab4807efe91
zc688a24e4df72446d13011f77123517585fd8a3068586d3f562ef9ecbbd76d470e2f5473f54416
zba27805284dd8ff9f252b3491401d6679a5c1984330ead9e31e7b0be1de23fbd9e0b4bee9885be
z775eefd460f7aeaf08af0d8691b336434331093b5cd8aae1628694b7eb56de35993a6e922a58a0
zb0aa1634875352ba421924bfd55fa12642548f40037719927ed6983d2ec21e6dd5dd10da20e166
z7cb8ed4f549c0a0b2b331d8697a77dd700024c1141c3e1d14e641aad793e93bf1c49b9c0035c85
z14154c48b0042701f49994d82617ebb19a369a376be9958bb652295eb034d71e1d35f783a245ea
zf72a538fabdec1cbb8ff1ef38f5c4c7adcc177187e4d37634a7506cd642703dbf4140515547c49
zedfda9914ddc060099006c04ec139099f6740410ac33627c9c655595687cbd30f91767f93a6bc3
zbcfc8df1d340287c768a5d78888f8b012c51f0171cfb8866976bd01eb8237e9188c1b414eb9a3a
ze67fc4ff717f9508a7afaf8f2cdb758761f860fca099c018e9af7c6110b2b0451205b47f126720
ze121923ad7b0010dfd5879de22ae6514e16e405f9051254ac34d95f0f865f942c8564287d66dec
zb8dd17fd590a0d85d48e1e9da66ccba8a1055998937c6c0bfa26d727fc93ad4024c5828587ceca
z26467002e16631db31a889d02418ed7bc3f1a8512f44b7aeed1e87ed31f4b704e2baa03d9df00d
z884d5709562234aae967405c45d410076c6138c8f8a3baa60080546cefe7566f295d029b198af6
ze1042c8edafa89c592f16d8b871ef302ca9de591c3310c42835eb32a1a4b4168d81817ff9acd4d
z4af104cc2f8f351e92c1fe9c29ee64d25f53dc0c6053e505b21af42151093b952879bf88a19a27
zc00eb52755ba7b7b8191416fdd27b4b5a0a9dee4e36ba965d2ed88c6291b91b6924794b08d6a48
zc6fa1348ce7544cbcc399eda5bdaa837a710b6d3a6dd55e828ccd15f59babe336077638037f2bb
zee4df4129baf7d33a977311d08085da46d91dda1109a740006a6fd15627bc145cc0814b1d4c185
z3fcb656c4799b69046ddd0f72c6a144c00912ec439eb90bce25a1ed569839bb419e530aa4170fb
za4a1ed209327eb82042d62804220c8f0c2939f838c67a9991fbf38ec9ccafca1d9206b6e3c2560
z82e3262e9f4b7bd352b6ca65c283a860c7bacb7971be2eb364d48b19155b96b0850675c57cb91a
zf629439ba5f1bbddc09584307c75e1cf49abc854a3f01998dc951921c4e4ad26761434b41039d7
z83927aaa93b6e325ed0731ceab41bd5e07f193dee7eb733ac706e494c72a96ce686267f51bf095
z911430c523dc521d7691d648a2efb91790d5bb37d3834981d0b0250af8d2d8f25defde01e8e410
z375b543b376930a915c6bae55a2ca300b2bbd520bae5f0492e6380a0fc456fd477cd262f6a46f6
z593def0656eeea9f78b23635611a8d11bdbbcdfdd7de979ac77fef2f0505a3c1e2b264324e7eed
z500a3b3a4dd72caf7314635ba1504cf4258b314163906d7353b3645453e9976c30dc3be675afcf
z4e93ef4e2be2c884c4bb071fee77a6691f9fb865c161f6f8a77ccee882a1d460425e0f4f0496db
zb1f7216256c94a883471fbb4f2188b674fe96574d37e6199081c1431f8aa4311642c259a3d0251
z7d2a5bb798e539c918b01d05ed1cbf2f6df6dcaa9f90cb210d1c7404f59c67e3ede3ef1fac82c7
z41f1e44e156f41122b489028805b6bc3a860e4869f124e74067f15e1392111b161c50a5bb7433b
z487b5175e4b136361ac7a270b8b42f65a2602fc68aec8acd24e8efe92e11ade8729b5662449e78
zffb4ce9ea5c9c4fc58b2077d54579babe683004e9ac946b1091cfb9cd42894736479d9d76e6f75
z71d4c6f74974adadef2786bb3552aa565722b0f7f83af60f505dd15418d34c4998fd6c1095398e
z1344b178d0aa1af7bedcd2d49b590016967998b5ef2a408afd0a1eb70924041d35c8e7ca1399e9
z9593bdfef416fd99aae947b2dc95fecc3ab9e74bed7e1445e318fb8af7d55d3241a1996d00f96f
z819bf7ab043d6104e188e5a5be0e10a1bdc230760805232df81cd21b1babe9d9717f917c1ac6fc
z5e779abd918e75f00cd21c94439833a7a27df204e6840c002a60bae649c967f2aec4544302b0d5
zae9311c7733e0c1839a7b99deeda278dc0642bc1f2f8720f18da0cee138015ed5bb5a6da2471e7
za5a36527c3fd28bf3ded6d495b887f7cac8a46ac5251054558dc67737ee515bbc597388e0410fd
zd76b13c7366fe702e613ec46de1f68754797eda93e0c8631b1f275b586c41c7a50ba54482c5c6e
z13b6a4489cd80b8ed65085694e63e0308e62797f9b927b8b9e6deeadd054bc56f9761e2826cbce
z901a5cb06d4f93a9cf3afba3983da540f61415e6e8bff65d07043e3d42c2ed5ccae5a8e3e1ce87
zf048fc193293d3788367012b378f1a1d4a34d7c20cae1af907530a597e5c46a229a54a9681c6b3
z0334a4d978f88b813cf469666ec3f9ba4b1b663c98c89262b8e8202afd99786270144a5df268c1
z87e907777e8ab49e20e2e4e6df332b54df6da16b46503b04ba98abfe2df26a05ec91e26e14fef0
z9a795cd94cfb850704747207cdfe726a62736d744b6b6b139e43127bfd583a339e06b0098ee675
zc6c8057d9f21d607b72fb97480910271fa529c1f77052b5f4f5a8642be31a1eae00595516327ff
zaedcebd8f9e1841f8c8da883642c86b21df9c583e0d762984011a7e3ff40b2e7fd2018a143f7d7
zc649db074a888a097a734428b285ba5d1551294e7069f95ca23564f9ca39bb53decef6a9390c79
z99e4bc177a8c83f7c6d940c94db6bcbc44285e9dd27efab4dc6ce51c019d5bb28b4f9fe3ed818b
zcb9fcc4b68f442dc3984d672b5dd1213377d33bf74f95c74949f698f93b98e3778cff67afecf1d
z67cba75803f3e8fb9fda84db8ccf18d9004096aa13308613207ccbd8fd418b4cd1e7ad54bf25d8
ze6e98eb0d5a1fa766d728b373cf8837fbed1910f0c932ea065a453dc3e12a21cc685d5b5e687ba
z2df2e6078c973119aa1d869e7cc0d11c69fb99e6de290137492edeef1cf4e54d7a550397096d3a
z33f3b0ecec4282a7ea8cca491fedce17e9518be6583c8e341fa3d3ec34621e44d3c9d06fef2aa7
z11dea6232a2c2afca3de8721b8dd4c0d810cf6cd2500e17f55f2beb57caad7c78c7c62d6825235
zfbb561a6db6f6a6057d80d3937f3bc10cf96ca28c5dcdca0c4145202ef740be8fe71b5eac0458e
z7d765fc2b273d3386c61c4d1e69a527c2c437afd0dbd2e093ffe1831a8d63c880c7f8edd6fa9f3
z191071e76577be29676abb8318fff984bc94c4cfef462178babbfca442feb1ca3770dc1cc512fc
z5b546cbca1d7cc769ba74fc08deeeeda87d0006767530e46d171b952241b01f1f4fe06dc2a114c
zb29cb023b9a157383809edf5f34df492e01d55a38992ba6deab9ab69fab294d75c3552e3e55dbe
z9e3649e798878e303cdd31d1a5b837e4d6211ddc929fa7af91024ce5d2039f66dd8234d413ef6b
z8ad088cf68ef713d64eb9a9dfe781e45d4ea1962abd70246c52b823c039595255e56352e78ecae
z23f976cdd478777f3d1ed1376c46339e18cf87c9df1cf847037831c02cbeea11cc7b41f52057f3
z4231d3562e43e96f39c2f74e4043d199f6b98ccdf556a1fc6aab762900c95b4e14cf7262fbb363
zcf687df24ef4ac755a41e8d4b1fb83ea25e6dfde3b396677d586083bd8398966882c8a0891dbe7
zd952bdfbc455a37af6c2fd269d1e93c0f3df7d43956268c8c0ac529f5db65744e7ae1a082e7ae5
z1f63290fb6182ed5001e48cb560e51b99109f1ab46fdfe326eef073d279b031d1ab4a48c2b586b
z6a95eec6d4510a14ac8d70c9535d06147cc736f9928bea5215ad20de4e552f9b7cf38eba7def87
z0241e2030981b7c06a718e2748eddc97e62e1230a7754eea227876a27adc7577defb8c9e99e3ca
zbfe3478c5304c4f4c81e6f506cfcb538b2afc93b4b63138d2e4c9c6c257ed54136dbfa5c979339
z755be27e275f79577a65d22f86e046cc0d38aee3795bfb4b35f78ce3c3badcba4e38b0fc928cf2
zb62ce3f038fccf9fce60397629c53f849f6859a310dc18977f9f82b6a3e4e255e02bcb38402cbb
zd2ea47ab7bca04f16ca495671d6bcaf9b31e788e81c29ca1423583e1950973e372a1d561372113
z59a0c7659860a165ee50f7ac8b6878ba753e2eacabb48005bf105b5aed09ea3961ba70ad7cf707
z871e69a138b09fa9194a2371505e0902262036425314a2ec1864176e731f06820eaa16b326fb35
z6cebfd04292637e4b614269a5e5abf4d8630b25295aecadaaa1d6f69d257a84552a08e59a76791
z786603142cac0d27fa34cca08c3076d4987cbb84393d10205cef252e2fe49775eb6529ddec4e1e
z7ad146597519d21a34920a4b8d84e64a126a912f3cef3ad95dc40856b7c8bfa9a75f517eb96a4b
z01e497a04a46e8a493d00ffdf139a18525ded18445e84b353b534c7c2c0f867858b899ebe6550d
z6283fa7aa25dfcf11751ca319c3836edc85cdcda7e2c8b922ff024111066532abdfc10a762a945
zf228e7adce45f06b9295855dffed9186d29ac4207eb7b01faf65dd80131b11ed157c4d98773eab
z3155ee9ec073d000ebe8fbcfca9ffd42f57ced76996cd4a5f4c1ff5c9d4b16699cf02c56d1cdf0
z82216aa0b581c4c47f0b31dfd31eed6671744673ebcf20b95a8022fe249cfa6597162e7cf515b1
zfb6014f72655c3bc060f2f94dfa2e00171085718a968bbb6c74efc7928da73573d57757fb1ebd8
z754ed24c02b81ec75ee71ad78eb01f85f8ac2bdd31eb04ca06109b5d7718f4590a1c5143c41084
z4c7978d8773c416a40208495d962693b762ecff9a55fd58b0fb4d544e79adf09b152a65fa9d63f
z2d0154470cb14796cb7892d6c750b5b5870603b7c52fc385a1c85ed8a99894a9fd4727403dc018
zc5a450d396127f24f99c982dd52438b5fcaec7be800077f2eb68ba0181bd0f51f09160d682197f
z3951485439de2c2c39750641d281a3582364329c21ef9183520caad35ed804e96385d845fea98a
zd8606ca608af844cecbf5466c6639c02cd73b58c5129692a3303d494b41e75bd10ab41ab4b0aed
zc41e1f57303b708125bac21edab388d08a393f094a3b9a22b289e6d42393486f943695627e0b61
z7591b1542df3e7cb1c31c96051396dd4349e9b1af0d0ac0f9c173ef9b793af7882cc88efeaf192
ze81c67f091a82b0ba05679ff00466cac49e8a1453f63edaf93cf28822484ce8b7f884b88084b1c
z18e2dc6bac87611014e36c02ec6c50529f62321183997040114c948cf99518d942ed6aa981ee7e
zf280b0c00f038e7d5051ef93d9292e9c53d128463adce362ad9809a54267ead6d927bd441fc9fc
z3541d74efebfc1aff229ba0cb47a11e869711d52f88b5d54b15208efc89469f133732dd9c661a7
z6f94dfedf57d8368f28fac594060b3a75120d802e1744542255d220c0c350f50412a7f087475c4
z04d1c28a85ee4cafd644b53cd0011d0fc4604fedf3da6f59f14eeed1474bcf488bf45806b5fd8f
z6d5735bfeb9a3e7c6b343a773bea771e8fc43d173c3e9848ea1b62a9cc228482299704da903354
zb0ec1ac2f49e144154f087bb07cd603b196c5cc184f61824a1776c3e4e489ebf58759918a8b81e
zacbc60c00116a634fe99cc4c79a96b59ba6156df9e2c3d9417a333b58461342d795bb1d07372d8
z6527ee9c2f98ca2a8d275dacb001d2d181fd13e817352aebec33d8541aec3d8654f88809fe31a2
z9df42cb83bb6bef08cd6f713b8e484f55d66dac78255b07449ef642bf09bc257766902c2b5f067
zc04e82b75190176f6dafa7210c31e50c9e9555c738df5b966eb3f2358da874aa3da5143a2ca21b
z47ebff9045919bbbe156bbff6296b95ee9439f4c57b425d9c09688abf9e1ec83b72f4130c8d216
z8a77db8d2ce60c44777aa2f988738969cb211714ae9d7b110f0ecd6d1837d7ceb1569d663b552b
z17aaf7aec5097bb8f4a3a4141d12c09807b5e93925d18fca6e8b25f027d97f8ff8c373b8b47b87
zbdcdb6dece11a5c5421dee368f4e01ed9bc481550fc6549b37a972ccb649c7c3443c7c7a4202c6
z5f0128ba04cc2b709e68d79bee244f521940b56a4181b9514d7e21e6cd42e2ec60a5ca667fe288
zefe0233214043feaa60fb845d90196e2d60c02c632ac06c6ffcc2b8144282ff57c2291919ad210
z23c75f47d70a101bfefb4ea94d6ef9389b2d79adea1d241be470d2ad3b0bdd57f42437e01fce33
zee894c2ea53058bf559225d438c65fdfbb2499115634a85f7365463d50d5d77cedb5ec6d2ee0e9
zc0171eabb5fa25a7d52bc60cc07a745a06d1a5d05b6c7ab829815d482c5a0ced65250fea3358f9
zd2e3214e1e18f05719cb2ec08bf1cdb1f277e8f7d596b50bae99dfbd817007e177825fb355a125
z5f3c5ca918f532d6343c8c2faea59b435af2b29d09a1e4ea84ea05152a3b7f65db378a0923e215
zea1146f6c56a106bcb504350f262a361bc40b7141eea4a6616e49948e0ae8e108e99d17eb72b4d
zded314d88c7e692471bb94376600fec65b7b7683170bc6990665badad0b014cd6c6e99bdb789c4
zc2fae73baeac7890424f645a41069ddcf91107881f0ce81aac9bdeb06f4ee38259a34fe25bdadd
zda756dbac2a924faea412fd12ce4c6213d6fcdbc535e76dc61d3eab3f36fb619fe30842e03c4ea
zde9e69195d2ef6e0a006ab0f18ac41d7b58d49d1b1e2d9f808f6bc22c276f50c433fc1f366bfc5
zcec821634a727165bd1e59234cfc73e8d010d85ab2319cda135d2abf3ac9b5ae038695edeeb3a9
z7e1b66fdb9c220016ca32fb6f60bbba6e8a0b42d6c11d33cb7d7a74f7b440e2931823c97845d92
zc51f4fc16b6f1c410962afc05e78012bddb9f22e6ba009cc3564bdb712892efd8c83379c44ab4c
z54d4a9d2f238725129937d41aa2649b7eef378745ca452e4340343f2065e2dc91f7789ce5df976
ze097310e5205dcf46a08f1245e0394f0fce3b29f46e45cf54a03d630c9060a6d936f1a4d91a65e
ze2230f5bf06f101881c097299c23abd40a51e2d7c4a7616bdbc4fc114c03aae323bb345b5c9e16
z48f06e03efea7d8692b06e8c28d2f877436d1e466c594ac6eb63017560b5fde3cba18bb94bbc8c
z310c98e45a169c1afd6a85e0e477982b070d39bbdc04bd9dc8c3faa9b872222e05635f01f4bc88
z0bceca74b282ddce9ee67f4fabc47f1e2ecc4f7a58cb404ece61b5438e0634b9631f55b2dc6a55
z1fb02566f5dcf13adaf8ec0b52b048f0efa4135fb3234a84dd71ef45b55cb61353ddb463d17a8e
z2126088716b29bacae5cca579323df339c02ed794fee8a745488303ecd1a6754c9182670651499
z90bae7a56f4bf8e94dc1ad34d7e0573662c10417bb733a8d5100247b69dd93d42fe88e24ac0cd4
z0e70bfdc910d2448f15c5606aebf4b0db0208e356bcbad8d34a0439e5c2944b3c149a94d6f3283
za0fbd0a4ce2d6ee74cd97f02cd702fd64019f0ec1c68c153e37183493b3d546c1dc186fb5871ef
zc67fcdabb953422cb0e6b6fb16a5ccbc39f7e8413ee8b02c114593db0069486aad42046e71a2ec
za282e7282193a0d76c6e290b26332c5dcea52cfc390f3a0d2607f4cc2f10698f51a3230904196a
z5cdc076c89fa7fae834dda1a33b40a6ba64c0d2c8a5409aba0763f34bf396fae217d7499a1375a
z4d76111465ee26b935b6656d0dc46c83f898452bd5d405db3b7ebb29133f5fcc116899dca10d2c
z78b1e2fede87b93ae518b9e0ae219e4d45e00bb91de059d1520a16418d89597e16f72ee6324fac
z7b7e0865795d797501be944b8e6ca14b8e4dc2ef89603f0d3bd433f56f6a39e78c0110e0de2b8c
z0b09b286d395fc63ab2848f161d57588d107dafa82fb3979aaf8fc1664a2d73b4d0b5ca5a11c69
z74bfdafa57186b4a77c107f86326dcb45735605ae3e38e654816e3d5b701add284fafb6f79fafd
zd1535add3597d2141fb065dfc9f4ff234495327ab78a89d61e1d0cc44815cb9709d544bd6ef050
zbff7380cb3c3d65dfd7ef06d06d526fdd869e7ad49ebd33237b8ed9f4aed610bdf0064874adfab
z5ed01f6335a84f8809803a607e8efc386692eea1bfbc7f93e5e02aa3c4426e33d6f90b1b0ddd08
zfc6116e9c076a2cab7f605a9f33aba6f0c65865809c720bbf10c5835581d827ec9fa6030b99980
zbd1c286830670e1670d5b59a03463eee153be0f5eb4faa7684f9e0dfc72a1e3cbff82b4d467833
z1635e609fca5008d80404fc92df8580e6542c48b100f451b406cdf94748797ae44669fec980463
z1084dd1eb6620d32357590110f7b97eb78b6e397f7d43761f704ab6fadda73687aab5744d2e2ad
zbacadfd04b67394021751a1f9a95b4af9306d624b4d319cc60cd773d165a8de6008bc4568eab7d
zd0c0d6830fd508a817f289836e9e2d4d5684da4c13f1a25a77935d0011a2ce8ebb18c594d8684c
zb566ee11482580d2956c17bcabf42c4c24d03e6406892d9db0fa5ee4b5e15e844a1a8618f14431
z8ab8d4b5e31fe3dbbb94132481d1969d5b2e0b0d96cb7c43f9f49171bb897110b2244dbf69ed47
zd3a628b08ef2e72a9cbb3e76ec8b5c76ffb0592eb1adfcef20be2d6684d2a9ccedd615a47869cd
z51224f5cf3bebed8333cd71a94239e109c37689c59d7df983d1bddbca949985a96d604ae4b4d7b
z755c618c4682230d7de78a6d190e946e6ee8c34dfa2bf341741773d78eb7b4ea2fd38fc20af720
z5063468566cb89cae2829f6463aaaf49136fffb419529af9a425b928b274fbc73f197f5bd6397e
z9bc74c73c0f5de4fecd59d8f4f7cb35cb5188c4d99571a1f66bce383a68b287302fa6cc511ae0b
ze16e7e76017629f4b2887475cfc6c5d43d20d57256bb8215cf38b790221eb544b10e2bd5251467
z909b3012fa9cc15d4ef6067bf1c97d2312a3fa6e31f68edcf79e93463a5ad1ae3e90275fd835fc
z703e6521bec19906c99b8a94a41e3ad3180941dbd683ee6df01690277a593a80b6a6e94c216c50
ze816270d34fa06b196041ab6255a66b479966aee67799f26587061b42ccb45a259aa6aabac432d
zc2b2c08417da584894c8aa4cfcdcbf4e241b33505d661dc7ef1cc20093a58ee6a4acbc78e7cc17
zfa09047cb3dde037f1d84da2783f480cd6744d68cfe7999e66759d80443a7eec01f5a5dcf69cad
z87269b6aef5e39371cbf7f7dd409868b673e6994b56d52a9054665abf0cab39b010cd82d7f84d6
z5de2de450f6ca618aac5158c794d2e9d229e7458ee6d76836c3047c9b2428b5db4b2fbb2d7d9b9
z7271f1b65c1eab56ddf256e41289eda9c6225f1f956689850e46786699fe0eef986ced378cb008
z172d7b5a25fb4ce3d88310c149ca61587f8aa5f39b186c22881d037ed5ec31c3969d60969e570c
ze686b8e15b1e84640957e31ed2ab904ad683c58a1a33f2d7d759cdc3e4762657d7a9cf796f92a0
z72d6ea7eb927898af3c4a287a5b363ecb0028d6f40d5c6cdb5e9fc36cd6ba2de3b75ece5393290
z1cb23cc237302d7171af76feb89ccff7304c6539075b81464f2da95e1de1df7f1699c30f6d6d65
z826f7098802d1b51b37297f2b949dbd7871f359d662926474bafd76886d712f2f0155f7230f5a6
z546ffca6840083300c60699cf20aef16b8e51b051e888f07b30d5d42bfeeafdde2dfbf0011624e
z0802283e9218a0224117c428cf4b64c424d0574c4ca30090d695ed504d1b3ae86f6e8519822086
z36413589b12568ce0f285beefdb9058f0683b6ed16067e4c6fccad5c1681f53f59ef5088a95628
z62411bf18786d2e50733e39f1e51af12b6607477beac5a4d7f3671197e6e34a720e2af9d848e13
zef311197cd3f3843544e24ebe782cc7401811460077b1877487dd603f6ea1d2b1acbaed513c5e5
zd00d47f499530e5aa62bbf6c19eebd97dccbda261da48776c09baa4f21bf693d7e9b2a6bf5b870
z055ba9656155dcb984a79caa63b9515041755808f3b2d46e1331a34b4cad6fd34636c923ae42ab
zab52c43ba7da4f43562f2afdfe1121aa7b420035590bebdfee620bad68c586b709bcab2643751f
zdf2719473f6c6012169e38cab620a63f8f519181512dc50a977d4d91d8f125f8f15e8f67a272ca
z299284adaa7c3e85c677f35cc5d5ae9131bd74bda35795eaeab6dbed0edac537be70b749ac3d12
z4b5e6d60b8863033cf1f45d501a1fd4e46b120c6395d8e5be58b97e0e79731b248420c6e547d1b
ze5b061b9b53999559b6d0785c7d116e3227e6b947942ee52448eb71adcbd2e44025602ddfb520c
z0cc9f759b649208da29b8debb5b76febc430a61fd5caa44d0643af2a0980f1145927ed46e15895
z95b7582daf8aec910d40ea385944d2a460b9a7dec2a04e75e332f1c229a368c839ff47137e9403
zbc32dcde1ab7d12cfb7a9668eae42bf8a194f8eb0d73bedb41e0851a4db9c2575a4a347f1a34ea
z826a57b5e7ec4b153b48624d5f8ee287602fa94389b8da39f23846f02ed5160bd0fbb5ca813219
z8e6f2ec1a6b98889e289e86a5440dd28738d956b7c0d13f1fcdb6bde81bf0ebb28717ad1d05684
z2a17e10d2657f73cda018becee6fabf78e85d3aba5bc31f3d2881829aaca185545b024e2dbb4aa
z2cc57788bed0968cdb10f9f00cdb3e653d732611a1b8570ca88d9845b336e0724a097ce49c8961
zc3fcc91f11c1ee67b1dafb463aeaf8e7615f1bb980bd4d710cd0d54aa78a701003dd22df554867
z5b7a0c8f6020245701578fbcce464bf6be062ed7f34e00ac3dd6573c91b3fccb7a0860acec8eb8
z27383dffb2f3dc8ddafcdfebdafc139daa80bd5a814c189ff162b6d01e7ad44f15f322739a9325
z6d6d64bfcab39c93750ce115554ed8681d0357f2aa2bb50b654a1f1c1711319b38c3c2ef2b9b63
z50cae50b0f60e7dcbb2da4220950b8d1a28a63bb6195ae317a89f869cb520a902aebe7a758da8f
z8237acae696a0d64e03da18e39b932546d2a99acfbce8bac6652b9efa90140e8607c278935c2a6
z9af6a525e440f2eb91f6e45e362b18318f481bcce44e88a70924040b0160886146e0c53d21fd64
ze7644df96495f50e3cb3d352e377ba76957d8488325bbe78000096f9ee1f1b7a1cb34eb3ca5b5c
z83a0ab17e5bde957410a7e104cbec889ceec32ff018c2c2664ff4f5bb3d2af0a9919a974852804
z4d4207d22b85359c347f5c54881ea48754ccae4211358bea5c792440cc9cd92a68922254ecc63e
z1fe488bd00a4829a0c5ed61d607c54a97b9dfc5a75d8cc224c0b5b7c51c73a5881796c98c63b8f
ze4782e2bed482a2dc299a63d3f391ceea34894dedd01b4224f0e8ecfdac60306782cc9ba4c406b
z909032bcb9de841b4115d877e0e1cd26f5c9e9de7c2f7afde3b1adbab7946131c994a441c9547e
z4607ae6ee98bc512872f6caa0632bff664f1f3c5b4130b8df88525f0202568fa28bdfc5d3b693a
z2b992dafe89d7c3e6fad6769e56fc5664af6be4705ce8379aa085d3fef55a2991e065661fc0a34
za74b3bf5a61c3cee3376a3d9456205a930318844c151e1e101de21344d5f03833802333e05b22d
z37758bf3cdc6588e726bfd9fe8d1e926c720c9666e771d8a49c079bde76b42a87565884a5cd18b
zabbd7c7f24356a3bb35db9da2c72e9cfbd31ac36648af9ba37cebea3cecf5d0be45f97c2ae9de0
z14b3997bda79e5f291740fe555e4367a5a8371ce798eae412f3893dfe4fcde9e73f0c1f33e19fc
z497e799396198f2b94a44bb4eff2f7cf92cdd888c81e79c9abdc696ea8c5c248646c5bc381b8b6
za6e64f226aebf017f7f42411f39dff11603db603ed5e771455e993ccaea7b1fa38374485761285
zb4ef44c128844f4707d3b94ee2676df3a4207fe1f77878fdd436cb9af4ab31b19d390c844d50dd
zf8e7e75ed1f3e07103bba21ef5af60b98f1f304f9b8c9c1c542097675d2d53147a7b565888ac8d
ze951e818f4ba3c88ad24a8ebdade45b9cad8aba0a9041163bcc01effd1de91304d1ae8b4638b39
z42c183f847f7814d41401b812b2753c3d9bad8a80da230a64e7d6271124a9e7acf04c280b86a82
z7214a676d7ede62895ba77fc8698a89ab750c81619e07339e5281576ae53fbbaa1efb0e3fbdbad
z9c3c0fdd513fa3b145487f5c78d2e9b03d37dd4a940cf77b8ebdc139f9204a04f2f28b95a699bc
z03730e820833784d54c236feb190ae67f69dd49ec3d11a4f640c28636d4add7b2c8c9e698d502f
zb4898cb1c6198aedf92439677348e90c54162d2770b00da87cd0275b271a2e549abddc305c473c
zf5f114b5a85b1a2d35c318fade197dc27021b55a7f720746be8c57bf721c9acab497645cf4b093
z739d2af24fa95b42beb3e0ee9b116fa36ab65edd11543aee76945312cffcbf0c46a9265baae1d0
z8e1f6c944515ae0640fdab50dff30faacea351b357ffe896588f12d39cb519d0dc4cb1eb06521d
ze0e70a395acd0e67974066f45f9551d0688311d0f0dcc58a1483fd11ae5aef9e363edf81e933b4
zbe249d85f86252fff6914b73d91e91a0ebcda16497b11ea42eedf0559fe98b18471e4533832c11
zaf3e400bea6b234d4ffd8b7a277f2c4aa110d51c790cf750ebe05d37b3bd2c9875940d51b83c11
z2cbcf73f86cec3898b9a7ef1e93dba020f14d030a993fa57ec49aacda3dfd6362b3b5676643546
ze8be716f58e8c8d92d7c4c662d46a7f1e22cbdd7dd223e8972c8e3b455435b03896db3c554957e
z962a635f2406aea73707ff6001d7e378265f4a4737d8cfd9252152c79dfc13032ace0611b45b32
zeacfeefda27fe26b20eb16c1c87ae31944d1811ac2ef6ddcca5553864162d991dd3a476c9c21bb
z79b8db16c08ba945be971b5e8d313ede91112c20fc11c978e0c21e74e2c825ea5c26ff8cd5bdcc
ze19d95ba57cd83b2d19e7453f3e8555fbb728730fd3faa0cc4f8cdb6c81ab4b6bd8370afebabad
ze1b88c16f6cbf12d3a1ec6b6d16ccbb5f19e74530d645d5dc64d9cc57f6ef8312958cb2550f05a
ze39f89d75c29791e0ac4cd2cde184103fdff663a681420239f495028f0477081ca1ce94f5c0a82
zddf603ad2f9c23d1ca64af44a48e0d5175aee79f5dcbb4a596f48c890d50fa279b16cf5b960e8c
zcb5293701f0162633257fe7ccf468e1b052cc18c77e4bed128d1e2c2465a997680d4625ed070ba
zb2efa70b4607d09efe015c4b9c498c12d3c56e5288968347233fa33e03f6ec7268430c6865432e
zd41999c469bc21da74ed122cc1a943e4f311fa0f2b8d773a07e784b7e9149972d053c923f58c45
z458ac3d49cdf9317d4b23dd27879cff5d8647e84b9856f5ef05ef0310c0b9d34141abc4cd5e57e
z1bc32560f847eee68befb232b9be304fba85ea2be12324937d0a38b95f4a25ccf7483754930223
zc44c01b94a4cece9f8d0fbc672971716b5d51dda7fa21a52ff0039f3b0d7f3d584e074d02d19e4
z7ee5765628117fe914402238017fb0fb63214e76acaabefb5c43b6480b3db70cddee7e6e3bf8ad
z3763beab314c910425b70dee2fd1079d8d7c875bce1a8b58a71723ed71d689f265e2d0382454f4
z3d9e555f09c5040cc899089e6b40b22d6020c471cde8235fc6051f945bdd9464d50bd97a3eef4c
zfff0fc91f67c24ed4c8c78e09e938cb7e5844c8a23f91c382d1785f0fd0f25b8c21bd522337bfc
z28a959b0227359cfc7fedbca61eeb9aefad4796723355278219b72dd5a922c318232bb5e6358bd
z3aca5f1828b73473dbb9bbcef84bd7f7343575f92168632858146bc13ce4babf897a78b52976f4
z6e46016ac3010cff1e761e12cee6849c2d799edf19c9229ba6b3cb04d5e1ef7ab74eb37c516b0e
z32881954db4d6197430b1a8bd3cd03c2605bd538d108d928753ff61d7997c3292dfd3c6422da89
z84a993967a155b861e45a4a31d6d00de73954e38134bd25be3b5dc6734e13c2eaee37a413ae997
z002cb386df2d7b74bbb125ca9be3348663ea448141a9cca41bd19ab4e676a8cecff8caa9aa146a
zd0190f0266c7c0e69a027c47bf5670fc9a87e52af0705e725b3cc25bed282006afb64888c3d65c
z7e631c5f0ba431b105268c88b19b54a0de9c5398df3f63af6340a90e24e45027143e087019efa5
za3ac42e702434edf2dbbfb1967fbfe3bb8c91ce9b7047aee2d7908c24bd408f7f44ae01ede5991
zc31ab0ab933787e7763b4c7e9323500afe646ab41f5665ae8cd5b93f6c80de654141cccc7406f6
z0804a4fde911350b9c9ec17c3fb2eb6c3e918c24e1567038c5f3088c1a3805bf9dcc31e184fc60
z332b4dc50fc018d1ff72a2cf7f302683840f7e6119319787ae41a209a77e886a1b31a3915bd7fa
z05c161c6ea6bffb84e3c7b33bcc212a8dd6c23fb18945349e23a5b646e3a22f1e2d55b8caa7a84
zf314ebe170a27e6e7206991b83f72efda4043f9679779317323ca0d93ff9bf4c9d763fcb40ba17
z0d1e4cd45d8cdf48d3404c13c7a261239e2e78b1182f5e5d64e591448b738ad3c69ce2fa6cb625
z212b043b2d26c1ccf2fec89a89191dd90f87d22db25e323fd0dd57d34fbd549197ac887f3af80c
z84dee335377a0450256f381d18bac22575341f3cb19f926ba608b7dd2bc5bf150b484fb9e51444
zc864bb2520ca5f81b0478d091a3b7988150190831a3c94429b4e54f1bfae2928c8742aa7543055
ze78d17e06cc7532d10c9a849e064ebcd4ca2d025906fe723ffe2e34a07343989642cad8b706a42
ze180c97423b564261ab1e778fc4391fb6871fcf88193bb6049752c3c25b7f6a378818cda3b2739
ze9b4c608d78d00b0e5e58a8a352d2a1778b3029ed5f8ca42de8a5c1bf6a165c73779723d3516a4
z09b36b19dc468aa36b7249d2fab6babab0cbf0ab3dce66481b21d0e3da3986c9df44f0ca467626
z5f3768ceb3aa20f3f6b249f88a5c3f6747420f6e7d363e07e091b7dee9b307319ea3a2f80e7a86
z0325708b1c66a56ddcb3702b272b96a89eefee7c4b98c428add1634843f089cb766fcd1b8ba52b
z0c051cb04691a6d2801700f66a14c806a8e80a3713c72cb9b90bc927cb143d30c6e11acc1a7ba7
z6bf806054b50e2eb596e7e218a88f68795be87a061daa78d19fa53a30fabf829a2218679e3b364
z3ae5903875bc7d8e568684d26b93ec1832e883b8e0808a79037ce58dc7cce38439059e835fbfde
z7647c42db115008a84340b18c3bb336d311ad7b18052d5bc954f4ac5dac84208c3a1f6e7fe147b
zfb2319360942b9a3cc6475e327078ec90cb91181edbac0eb98ad0693b02cc8e58e381113186e90
zf7fad306f664b2075c71e906c27feed9ab099d711c6c8f165cfc045328cbd6d1cf47c0bbfb54f2
zaabda66ff31352e0db7423c386f5d78a67624682884a662988dbcb681a1a32eecbb93b97fa6396
z84cabf9f472b83f0938b1fca57e13d3759d7a3b9c8e9cf3bca91e07ef338c0fc721eede30080a6
z94c2ad278799f5abfec66de6cfa9fdeb7baed1c4be96231252afc1dfbc574cd259130685a48235
zc015a79065cd8269f5b5f1d2f2fb90dba987fbc2c1f0bade81a7471be47f705508ee150f646bb7
zff8bab80a2f62051c0808b99de74b263ccf06c22805f40aaa01b377ddc130a5779e1d7948567bc
z74c41f1308d3b283040bbc93696c906f21e5f9d75f1d1c3f43d1f8d64730137827204e791077ec
zcc55c3eb4974dd5356fbf9f0a70f7f592f4c3a74c38ae70661a817e2e8d62e62da33780e590fe4
z52a5a79b301d00ea6266d0c3707934ced274696ca2bc0b1f31abd48dd00b0169ee54025afa4d31
z46de88a4f9c320860e91bfb04040c15daaa16441e6e5ff375083f41b79ceddf7938cce12ff0886
z5326ffa5732662be4d55e9dd1fef968c6d761f9cdd2bcfa37aa1c8b08b5eaae54f7c3340f5a870
z7b7f14e05296bc362b0feb69d89f5264e7e8b4ab031142342ff7e46e4279f3ba4b50afd122bf16
z1438acdf27fb8377b2786a6b7b3f1c878ca77e11f43c124796b80ae136c9485567e83877670879
z55fde32c4c1c2f3351a5a45ad4122df871de3817ef497e29b4327d30a249a1ac2ed7f849312d9e
za8a826c9a27beb51cdd4930c26856971e68c3d5eae2feaf2e1c88c25949934da15b2904c13989f
zcc926c127037000430c6925046038df7929b62c1bdb4289bea03383bcb2cd166db02eadf577917
z67a34aa195ba6b03213e60fd3fbdb74285f63091a55894f2418244186d7c9baa0db0f96c162bc9
z350c87832484bff831ea8df52f29ef79ba5bea1ce5909638f8133baf99e45a00e85c660e854b1b
ze9c19694a18b8820720d10ef01f06082c6c498ebf82a9195572ea76aaf3760d92d4909228ff816
z8efd5998fb76cb120eea0b786571f87cf89e01b23fb92df7e1bea1babc0b0f1ec3cb875de15cf1
zf710d0bef8fec295c84675ddf6516ed65e77168b7cb9cd9be17440be21da82543fc1a9a7390111
zddc85334e5552ba043202338ae1686b1012e03dec4b8799279cc334f933eadbab22e7b92d6e739
zc8e6045651abbac6d1fab1ffbc4fa43bf5d587b68eab248c52227b91bcfdd84983df5d0a9a7c74
zd10b48bd2824067c710301fdb8a56b7b96441ca01f3d7671a6560ea444b4d0d8672d0d514b61d0
z5862028cfa0077388e46a1cb2384c678d33e9d5c83d890728abde139a0a41ca9e42d05052b5d5f
z4194feaf5c8379606b7a524cda8d41e6c4fa0fd389066314d6a75ee3aff46d6afcab57e3d150c0
z3bc838aaf4f69997237c4fcfca2f6da8d945a9451ca194dab689ac92f96bc6dbadc4119009a934
z75f35628b402fbed336dd6ae9a64302574337c057db9a19147d4a4249def354c022c160e911cca
z18a92fbb82c5046b052bda0a63e22230653817452fc339e114ea513f7ae11bbd2e6cdb2d4946c4
zcbc8f511340320c75c51ef049693c56248bf64c54769284633ac4a1b9e6c34cd4f6f1b5ae6e0e7
zd614fc436136b4f8230000deca3d0312027f3a529907fc2a3e6f5fe0842d706117a240a59c6c88
z5f11ff923b3e2b77f220362f203dd26363df47ccb7c9aa6d949591d71722a262514fa26cf27d4e
z66d75f0a8870447e5eedc677e88b8f3ab8661bff916eeba8211c0ecc9201cbfacbd2a1b14d5159
z16359b71b498712e07774cbb7458e5dd5d8eb85b8fb534a6d25956678ac528fed15b65e6a63c67
zc70e25207b6a6077f8795a64877e6155f42a4af0ef2ff072f117eaeb31da4b8a0d9d45be2dffa7
zafc8395935d366494946f8700220b9596849c4497be506bdd3b9af12a1bea5e176b2bedca7559b
z1df6c99c6e4e422c6e52fd32ac34ada181f5a847d23c6b72d97c6abe9d4f6328c55cc9c395ead7
ze700a618b3f4a03ae169497fc6805b3a1aad7672397f223e3cdb26460eb421a4106fcb25b5cd24
z47b5858d48d73cf8c3d3a6587d13366c543bdcdd0a98cb9a42dba68448f3058517b40ac452f6a1
z0a4345c08320e1c8652bf793a8b0b540ccc761cb8d37b0c0bda8d1e8cf8cfa670c5651a241a725
ze22830cb2b2c50901eba174b4a1cb0c808ee81290faef2d635158b9cc5abe27861d835a64a5874
z8b4fedfd673056caf0a7a53b9e5fa73ddab1afd86ef3a83f331428b72b0b9d0035f86dcad12944
z445a699828bd0060e52f9be1853ebaa43ff43f4973c05ca9eec1b9f829b3974e9b7094254a7d22
z6756bc588bda89939b449d2f1f1ab27fa6a95e0bdd3628415655920027c02f3a2ee0bf4d9b2796
z5cb6c46ff5e02544bc9c481514e3a192ab66f7345fbab8d210c119ce3a7e3c1fb93cf059908f0f
z09f5d062e508ee1994cc3d12a1f8cfa556bd59a56a9310bbce4e8f2d2a56fcafa4212d93971d96
zc309e887b2710efb9f70835f83cc645348aee6f2b4bbb01a108cc4cfc5f929fc794a03d545c8be
z1d80827f0e0c0dd07c3193f12db77bd1f7f11d0d78a7bf46819859144cf8cadbe4efa10302bb99
z3645cd35444c65362adff4e93470863100683e72a17e02b8aadcb15a6b4f74963b70c8e9052dc3
z7a1205e9e04c7ce13162ee2140a13823c57afbb819734de093ac8f3dbcd714f988c482984dcd90
z7ed8e886bbb60094c4ba05d53c804baf2b8a9a699c08a38f5ae2b212d86398624e6325cad66fe6
z8b326559ce19bf5f6248a54f8b70ed68f4e6cb687eb1e2e071df0ac7567c57912db39bc4d539f5
z42a72c43d3da8c6638e8798f2c3a836a4c502b683dfdf5baf32adb6a04564742603a1f6d896229
zbabd77ee4d33c3efa564a3bae93abe7d9d77183deb5dae17ac82b36c15c650083362fd2c7c6758
zf1aa0f2d09a07c1c68157fd5dcd10ce334f681d47480c092f474fb0a05e79ff11d3854b640c9a7
z8b6920ba82ee4cd68d803e1fd29b8a35cc6a4f79e6446f0ddf2f7db800907e2ee75e194a7169b8
zefce5743fe280e46d394628b9d82c0c402a778e0403776e2f1e5594cc4597f0c151c783f87915d
zc61d27d37cc308bf3aa79960da3b19067657b9699c4ce7dbe86ae4404620950fc8b00f2ea4b7d4
zaac61801a025362403a24f6f11b88515dff707b58ef6f7bea7fc7f3d3182c946d738b38961262c
zd9a0f8c009917b9a420d582c929858ab50349ed7a6ca89fcf2b14adf3647333e23f10409ed1182
z4b5fa8da8bf4e7870f696b119326a5551d59dec7f0e3eac230eaa405a079e994e8356df17d471c
ze2d2a2fbccee73d7f4f83fe85a3dca6c61f69a92417f0de3c089993f5bb1de08f2dddd1399f21c
z0de5743f22237a1b06f14da44b8e71a07fc675a8ed1f169a1e83c1095040a0f951a0a4756ae89f
z204e0c96ca0c505c3adb6c9ccdad179c7d7a66d89044070c3f5e17adc5d9a9a492bd1c409fc471
z65aa1bee63d86304e6afc92886e30fd3b0ce3661a35374c49994bbe6f3777ad5d27ab7f55c2bb5
zf7be767c76bbe3f74d1eabd4415d3f32f1d207ffc45fadb16cc9226eb76072ee02d727937ce4f0
zb020263ff0e7462deadbfe85a4cbd9c534f5442f8e2c788a2860d89b30d8e311d46ddf84ada924
z5fd70b03a5430495fe996fbe006435520ca3398c48035f13a1a027bb39a48c5b426de03a41e4d7
zfb0f800a34f8b3bd2c89bb46476cbafe55867ae30ee736c54dfd4dbe276774c710368971742318
z9eac0a7f8ec80ab734de0761d7608ccc68aefe72fd0a89aa4515338ebd2463ad58f849b7a5ddac
z65cb17fca4f6eeffe872ccaab4ff5256c258d94127e5c69f59b31fd4c3f580cfea6cf2b63d37c5
z74fec114563e7b78cfdee7a997ce8b3ebac9a59807ae2f08e41300b23ecc10e5fdc0b80b3d86e5
z5538cc4514465500d9cde7d4e1b59a588a96429e3292a296dda46019e0eec2fc720002b49c40dc
z54338f9354dead354909ec6d3dd37ee7a6e25ab2f2a03e5e6313681aec8c594abc5ca51688be7d
zb9a7d531fc9c34a3097d6891abd8e55ea9529679bd729adea1ef44356e4d724dc70783e2ad6ab6
z5b43ba96bd3e52942c003911de3442bfb210e20662f8663e4dbf1435369df2922362c9db5a109b
z80c0fe46e1cce7203be2d53b2dbe9460191ddab7664b238b6cb031e6f73ea5aafab47f9a29a21a
ze34795a3876e5446b58e0c0ac9fd5142e10784a85c93ccd2c9d929aa537fad649a01da097cd89e
z72d76d30668b8671bd5ec64e74a2c65b62d33615c64807a72a1d39c3974ed74130f838a29ac9c3
z1b173d219127b126bc7084c164accb791ddfda68a2a6f0268b403958e9bf82ceb345a39d3330f1
zd20d1bb66f0739b4e853218629473643ebb2500c641748c8bb81f73e440f04d849e4352dd40559
z0f0ead3f299617cb5eb0d7f11b289db0778f0122e386a7852a60a49522589ee9dcf6ae85fbe1cd
z113ce031eee0998c4b59c3971a96e8b65c2ce02fa21cdfafa4f0ee3ebd328989588ddb19d58e91
z43da8d2107437cbc34d454702eed5f1be2a37797660724c3d0bece104fef7104395a2427620aaa
z4c6cd4270067bf2c5cc3586c425a05ea629c34399fc28f1d35bd99b9346965624112f55dcab2dc
z5192a107a9487ff64392f5cc1c84f468f1b51f60032ca886be2358ff6225f7282371a3ac41219d
zcbbe11d242543e2a9889289b9b47caa9d1dac1fedbc0756b9284a475dff73c5d3c7472b66a0d00
z033bd514a9d5775b0e0f9a6ae3380513b0db39faa65da934890278b2680b790f19109a72b07d8d
zd3a0e1639f8f337921de0df641197795c574fa2312431300e1708ed32c975e252199ea09ffd640
z92817fed6a6d4b60f40bccc46300fc76aadc8f4b7afe9e25081899aa80411fee925ec1c54b9a0c
z9578a0230135144c426877ba76e84203c840070f5ba7b7dc8a8eefd0b5692721724609fe4093f2
zbd2d3dab1e7265143bbd108c421b40e1880254abd9f5c4caff864072d93145b0fc4019579538f1
z7e8d9cfcdae0f0fcc05a451c45f2fd94841148817fe786dbb38f10470d602e5132311e59154135
z24a1ea1599d2e09ab082f353e89bfcde011049712371fe44733ec670e9665d4d67d36904ddf357
zf2a217a39068272bd1282b80e83b847fdc7f6c4fc6a4bcd71857974f91a7daa4b287e0abc152cb
z8d05e2b5f56ca7f0198ca707d1d6b9a5e89ad5d832a3c48aac4acdb85f6cc4f5f7ceb1535cf9d1
z7c9b1a425eba4f79e4bd4369f548ea21bf1a9aa37a071d6a0250d5033e278ca3f2a8ab39ec3a2b
z76196aae5b5e60d80e7715b26672b002491619e6804c208d1e5d82b74a4debd75c98c807840a01
ze82899d650cf2d36081a8d8150751df36256cadde230902f4d1e916c8970bc3186eed48b9ecb38
z5e168c52263f3c1e86a13661dc6f9088cb1f302e4aa5b74857f77f65bdf335ec65f1954297ac75
z1f053bb290d82b120f3d88427110fa821574e01bb1194ccc8ac259f3f76d855cc083621acc7ea6
z46aa6eb8eb9beca7852f8e33897f99e2692a1eb6261a7a8d2e57344a125f81d758d7ca7e7c9f42
zb9055b1ff64738deceda58cf504a939aca33ddb96a9e9d3ed3a1dff8e2d52ff20799ecac182f19
zd2a352b532541209de5c29d6973178a8a31bde5d086cfc118cd89651aafc1910ad2304bee9abaa
za36130eecefa38c0c4d61242ee21aca3a13721333bbe6d0be865cb67f95eb8034d68878a27ad1e
z3e37b0a92f230d4d2eee2393afec026b6782c21a78f7e7a61fae19d85a184191b1d4dfdb742f35
z0cdc8ab829c0f64d94fefc457afc372af830c1e2b729b250db2557b28ab344345d99cb322d6be2
zef236a5d081072787ad70949a338896ab1b942c43e1ab5e81edb257eb3ceb2479289260fff94b0
zf6023bb0d90f8435f362fa4931bac474a931612338b2e664a8d0f0b0c2f888c42b6b011bda8712
z2f4e86d726d839c787f8e6c02ddc4ed9b7ab754af102e8cb7af3628411b57ce6423a9f1eab9410
z0d98b70e4f34e1d9115dc2cba6f88a4db01bf399845833ee33060ed45d2eeebaa919761ca98671
z9a0df155657923d71c6f9e25457b56f2bb1a8f6c90447b1e10e97f5fd11109ea1d03f22ce83a71
z6c69a581cad46a54efc8586c8c59e81f67a14b054f349b9c15a2536ec1ba798eb18db614801ebd
z2c5d99f6184645274ca1bffe4fcd3f8cc55bbef96020f2d4f84e3ff35587a432a99eca22b201e5
z9e8f475a4b9fe54deb768d5e116ec955903fe821835852ab8996f6792a3d9d0fa3361846704f60
zcd9e9460d310bf13efac02b7aa138e6dd35dafe92c2a66a23af6d3305075bed3f811d14fde1a0e
zcfebba6bea03b4972281f8d07ed3454a2e69004f54ff4616a4bf718f6b260ced6403ccf37a843f
z9cb8ebad7671265852a0d2e331f000f5ff30a4d7867ce1dda33267ef8ef3646f9414300bf08781
z4a7ee577a3a4dd14d09d2d6d27b1ae3ac3420fa9b6d26daf09f12e069ac5dde3960c314af33ee9
zc1ec141470953315cda2413a1415d0e9ce6c4cfa3d1dbf4cdbafa08e4be6402300c9d0f465240d
z21e1204aab36b8aba63421704ae8f8665e465dc0de8ee99380a6aeb140492516ada3ac6990cc5c
zafbf1240813201e046a5e2781e36327bd7ea2a6577210ebf521684afcfcff2d173c9df25a1eb07
zc263b318d9300f830fb9572ebdb22ea3853d10a3ffd547965d350a81671bc24443c97fa065efab
z305e89298b7c4dd8e248c8c0818cd7a2c35f04fa4c4b673b929cd8a1c8df9128a103823c7950bf
ze252716b2af3087262c9633807097389fa16f58c76310987d019f4d6a87143c9d931fe3c6b6a42
z2b4422899112e7bba6d60701bce1ae3fe02be641b58fdb813c07d3a3687614ad6ffb4235f24919
z252fbad9451cf113b3db22101452c3a47f64182e0b51a055b753b9158908cdb921859c54c88405
z0d67793452a9d7d86656a95cbb69b13f28f1f3b86e3512987d475ef991cb6fc062a40934440b67
z852b6200cf4c32a096ecc0408c00fcd12f091930784da63f7f602ac8292abedb238b241b442048
z7719c18c0f2e2d51a8f7cfe421e90f001fccd9a256c3e2a58bc59a29ab1d624a55d99b9109e93e
z1d84bbf2062a20da3c73debcc4593a548f8aa70bf2fd3e993c5c3a184d438e4c0b3c67a490874e
zd0f33ce233dffa485159fd4ee97dfa992d94ab9523abd844043eecce55f01004e1a16fd3c77607
z4bb568d208f59f8a565f8541e2661e1bf8d4f77a2b4a5c5b2e04079d21e40165d29d23bacdd5f4
z1b1683be54a83be0bb784cd75a013cf1b47dce34c5c86d7549add22dea6bab8c2c221686959d3b
z3f5aa0fc98d45e314b7dd6d7cc8dd49bcb09def24526702a50584baec2ac5b320cc43badb7be36
zdda7cfebef23e70396635a4f133fd3be70a96c773bf9395b831732a785fd55e963e97bce8316de
z592933e87e54b89df2fa0f7c2402a19ce85d0803bc495f89cf00fe86669135ba6726647e0f3077
z545bb783bdf5da486559ab3afe0f8e791c92b1c300c892d3e452f4cda23a7c94312be80ed7fc88
zd199f744336a051dd7c7e057df46d62ba0cfe34789b9eae3470c41a178b7a0c42475f2fac9b052
z6a15d048a927d6ec6c5cdebc7b832c273f3060fb342755baa2c22a494c5f08d34b1cd0caa96203
z948fc4df195a2c831c94b04aa9bd7a1b9d33bfb4199cf865c075edf4d0b64e4bc237b2f88270a1
zc282a28a6a3ecd8b93465eedc0e50d0ff788d1613d4edbdf92a9e5a924bb3b5588fc26c4324126
z587175bbed971579cd752a757810f3f5c0a98e9d12031f7af0810b9bb7d275431259efcdd2e061
zf938f94d7f457688146278a3edcf3b8cbc6f671ebca2e59a76bc23bce1f466f8b14bde266f33ce
z0da23e5542f332760017026d7fed3428776a2205aef350b47a4db204cbd104dbba67e14a859047
z708c51fa2b9d3b1da4b267497f96785805f9cefd95a27b29c30988f9f18ec03c6fd10204b81f61
za6bbc9d348e213eab518cc0f51b23978c4c72582d65a8de831d5fcf3bc0b858bc49fc38a520fe9
zf0538100c148553fa6da823fba48e95414877692b293cb2ff31ee4c57301ee0316c0a29cc34274
z50e48de750e4053cdb9e130cdadd330f9d3fc657086badc6a1bf7dc5b1d235d858ebd00a907dfd
z4a00f979e4ed686dca06b1b1cbeefbc6b4efbf1c4be045a27bf4cbd2a1d920dd3155ae22190007
zf9118c9e7b95f27620f934fbc35a4cdfd4847d79ef7e9cbf093de49d1ed9d1a257dc1293544182
z7424f1b5a8347ff459a370ca440741fb90235b2c4a963e3606a355d08cd83fb66d17fe4ad2ad21
z8f109692c17723fc2d90f99314c9231ec055ba7454ea503241a7ce6593e9639498bebd7e9525b9
zb0401bf10731808b9720fa5043f691fd4541b07767ff6667d95a0f653bf3cdbdaed9ae41854198
zf92725eda821267102e2582dcad8ca73c47ae4ec4454de2896d1d121ef31bcd751c6e5ef58c829
z4aeeb9d825936475ad8ca704c74c7948861d82c61f52a4162917d43269cf2a40305d1d33b7c108
zad1cc2619f4810693a50e410a35a5a3731e2e6c0baff3ccc106d5b6a4898cbf31952ac05fcbe0e
z6de6d2958910595723a7d2806003003d8fca9d1608062d26c527b99cd7f7bfff75f34d67fc41db
z85652cc47b99d16ae8f26a481d9ffd6201d35f452fa50d7b2b03de7a8b11da8feded879e785d9d
zf6135da8368d7e52f630882b6d0282d226a02b46a03e784185541a12c3d544edf0bfb8aecc8460
z7076018f1b76f2846ae8bc211f94c5652c0b9f64b1f4e80d693ad0f8b691361aff72e65cd3e086
z1435e27026cbd88db74e64f3ccf4c38adff88cda74fb828d743e308e81a68b52d28a7a421b7ce0
zf6897e1911ea2d960c99bf7a2199b0ff1ad46b8abd287f7b0540215d74ffe3e7f5b88e8e5651f8
z372e773bc8a18c4c75c906867f1508a355b23fed7411906873238af284925c38efd9e4c40958bd
zb04c749782fcd640dc2462e908a9e08fb01640b38dbe1da6e6394491adb1eb315e6d8bce99b2e0
z21ea16e52a31cf7c2b42d8672522e631e7dba640ac2e39f4a125c24c44f37b2835eeb8b3f86ce9
z4a3aa11529e1de891ff2bb0a19247abaedf0e9cd6e20b20c205e88e19312cb058d480664dc4e31
z345f198ed02ed7510f99946db5a74a0173fc08f805df03cf9b5d40b5e98cfe3eee7fd998858818
z4410648f822dc81dbff4a9345a879af17af5e7f32aa4168656999c2ab004d076821dbdcb2aacaf
z6ad308e585a6305a4d81348574e07920025f7042ea372f766bbb36b5c3f7ee0b4da54c6c7876cd
ze6719d060032b2110a53fe660d820e5e4efcca8fa1005b663e83181767644bf234aba8ce6761b8
zf639014fa36aa109c4ac42130a72f5adc2e2ccc4e949ed691566e881fbd6fd7f04644c4209834a
z5438fc84b8a26b79deb2eed2e02b5dda3641a3b586c6fd58ed159fee2f78fdd38738d8f13aad63
za3999da04a21baeba168f896595290a91193920d86496616695cbbf1bb055c281bd61299348cbf
z7a7eef182cc365e31b36c0ee6c4d0b8242fd9c354afa30426b84dc835065de3ffdfb2cdf82b547
z0455f9d15baf7fb14fc0103744259b9a139185e170ddda2a2df3df938ce494af8b357209f214a5
z74b487574b8306c85e43b6ce0d02a7795d7485320e2e7bee6a7cf9973d09ca48cbeac2209c70f0
z7383e352290492bc071fc70b21ef281f71fae821302123cb2db2c449043c5860969da721877c4b
z35d1e43e18d70b19710f1975c430f14bcfbc92afca03c00d399fbcdb3ed48de0d794e000ee2a2e
zad1cfc1048537ddcd808473f57512e076d4ed16cc9ac1f61df713e9a4a8194352447c7f9f11180
z7bfae2bfcae1f2da8aeee81bc333ebea2aec5a41f65ea11c090864ad89f372bb9ddf3485a0c920
zbdffed163d2f92b489ac6d98cc774a835f709e390cca77c37c8ab1f4091bacf47124e9dbaa3812
z63884f2fff7278d8ab82d5613eaa401c5a1f1c822bf1fbc130107f5623686c2d849ca6c628c5aa
z4db95e5635e90d0c9c4e90a27eb667bc1fe27df4634b1986ea510eea6716f7230f9eb6cb256913
za5408d452ef5725b31523b41ade6756bd3a95d064531a31796480f8b421e7db260aa7da966c254
z691cf9478fbbae89fb89bc32de08cbadca104a2ac9c21516e237e37c50dcf7bdc85eb6360b4497
z8d35caf689cbdf73eb55fda4ea92f55cb136f3cc0ec0e5e2dfbd11cd326b3624d186fb44787e27
zc7cef225750c34867d6439c5335f3c7d0329ad42b7bfae6e83ed82d1af3bbadf515019eb7da5dc
z40b47edbd7b2f650d930811d88376d53206ee0034c78f5df8c72d9298b94ef784eace04e35a6c8
z5e56f698a99ab76001c7d9cc8869f0015651e2f8aca301ce2bf630e69dd7a55f67f1249360974b
zb10bd43db70f9b7451d4d4387279b86e42c979ddb5924c18ec9a47ef6b81250994ea24e22f1bf5
zff391ed4335bb65a3f57555601abd1331bbeff32696f62fe614a7cf979937fc846d71f4eaf1228
z3c10ab0976511790e45d0e22baef25a61559014cd0efe79cf48c8d99a668331704fad5278ef26d
za85ece74b82a01d405fc19ee332451385041d00403bfcb407cb605d91cd37f7d123428b3b72c2d
z3f8a9370b9401cd8f86b9f58c6e4a4b33b874c1a7eb9381efbdd014185ca6c96474a7eec8fe79d
zb3cebb354e346f2e0de7839bb2fee0b2d240c68738f6a22f7ad581c7f3def2daa2631f99034cc6
z6636e8d7906c2d75dccada341dae18ade659c952606a951a975fd384a18278367402913122ea8f
z47f8e9214784c4266fccd0b13ca3e68c3223883ab8a7dc6762940d66ead6cc9fd1707c4a444419
zd9c33e87942beafae7231365de38509ecfbcc020c778f31103b2182f07910a98f7513ebc668408
z6194cdebbe6e8eb6d1f16cfe07368ab29ab9c9058b0e3d361f520f77c76fb79c0bf1295bc75619
z8ba206c99897d3d0eb1f60e621eb9e0f0a063d819f35c2ba1f38c662d8de37e004c0574cc285d8
z484bc522babbf9fa69036cabdc6f74bcabcb6846f64443828233716ab8adaf4a152f186690d955
zcf384ff408d7894cec23728e07c5d38a87b6066bb0faf3dc5dff4a29d5c4292a4e121cf89fe568
z2cf69695362e225098ea9fa32aca76f48e8d399d59115fb07846ff9ef6f8f0b7263a9c1ced2ef8
z5ace99f548fae2effc88d404f2f33ab009e31b15b6ebbd84f7bf63ca8020c3be4db02da52d8efd
z7ea340a580e52e361ef86e5ae8ed94c52151ebc1d094221354a568b67f6d34d875ec82bdc8092b
z10323fd5516b366838a74c709778446f1e368760c88c442dbdb3999c6a634042b1a9850909dade
zce73403f0599eb4a07a7d1eacf96798e067d3950bc28653fe6f01c6f44c998dc7932ce4db2344a
z2513692310c5c8fde09e37756de74d0583115705ccc25e3fc1fd180fcf4ee2abb42fb095be34e1
z4251a49711154bcda596a1aec46aa5580fb4c6903ca09a090de300ff6fc99cb5847affe5c88eb7
zedb591f0108c29b1be6bbf39515c532b429c43313dae35134170a99886a1a71cd9cd7a5cf6ab75
zfe88acc5bd02bf6aff1967435b92a4b35eb717a9b2dc89b3dcc14990993adc0dc838dbf910345e
zbf47563a0a7af09bf735c090bd006df39a5725e157f8ecf1b0e1ad646f2f301c629bf9a4092536
z14a43d5960804ec6c3cb6eec755d2fa75adeb0af703320ae2aaeced7cd506144101550c870e07e
ze9e0d96a7f542ac0e2a188a10a6ce1d5aca6cb2712b83f6b7c130fc64476e8df088b3a1944535e
zffc9e22eccb75272743f82a4c44bd997f6a7e9fc3267075983cbfbeb502062d2651d215e5b8711
z2c9d81bbc8b94b2b309dc1a42da474528f07747fc09d9677bc7fc194b7703879d32ec7b99c7dcd
z68c7617c725a32024ed89ec1398f4cbac2f81007d59c87b2f2be350d4a1ed28c12ca6cfe70b01a
zed83e8593ae322baeedcb3b1b81f557992645a8716522e4b3551d2f01930b62647b0dc5bd9739d
z55789c6de92fe02e8748570806cf9e875c7357516e99f3ad7e668b58fa161f3e8a058dbc1adfd6
z2f00669f018392804fd45a38d2affc16ec22cf75c4a602607f3c1f38a83cef9594f669175e7c0e
z523b99c8747d992631bb42f2fb2e5c407cc77dfc22e87c7e48ce5cc9cd28e5194569b754bfd329
z994c5f7795f675d951ec3ddceb6e895fc2ade62fc4f631361fc9f6aae297fd0c8ea8d7432cfa2c
ze3eaf167fc0d4c0b50fdd0983194d041e6df82e69b20ec52cb19c84aba8e0042e213006b2a15da
z77260de33bbce06f876a8c5a6251d360a02abdc835a6cdb58afa28dca962f483f5b12cd9ff8614
z954e029d030a515c0864d36faad5fd218607da811cfead597c8f792aa4cc5b6a46c2bf6cb1d12a
zab1b411412981a539ac4d3f71272ee0774787745a618204790321372bda66b4b75d0de91f6a092
za0bd95d148bde7368721bcce693b855545f6773958eea789a07386e2d454a00c98343efbdedc0e
z49f15cd5ab55f6c3a457f4cbe5c108ab3faddc097ea2241f035be3b28dfe3fb97e8da4a556be06
zf6889192c31405d1bc827a1551e818afddec9fe5eed6b349daea40f625e22e92f519593b76931c
z8711c70343a3ef3c5df455bc110b3d32bb0bbbb48bec2360b1de134975cc0407c91afbc6ba9585
zdf1762d3070ca6c3351e29377f20c225e7998f8f934a441a5f226113c16aa1de75898ed23bebf5
zc2815c9efd10cab784f5f970d86b432fbaefc8c0a5ae7bc94685696e6da72e6403149412f9708e
zea1acb851b588a77ab6c8794a35fa84d8344c6e23513e2ceb68f4f8dd09ba83909557eb5ccfe2e
zd25aa9567b6dd5cf83dd5815e7d057e078cdfbb2ddc5e9d0eb141b22e7f4433a8eeb5af7aa811b
z2d77beec4c02306cd3ec92f0150b06dff52a2f2b1e15a5bf6f6295b47275c4da27efbad24902db
zb31459ecccccf509601d37c0181af532613510bb8ad63905d641921ff5e5d52c3a19512d8152be
z102d7ab0474dc283a6949fcc6f8eb7b2bd346b4c28d645e2a9320a8ce2edce7f45c5fe72b255ca
z0576ce0465822f299a6fc543dcdf96bade5c021b8758085528785072a9c17aad6797eac040469c
za240b3f058fae5ca3405a15304a92b09bbbce88292ee2cfe9166ce7cf35de491586dc44c2cffc5
z89ec36e25a61a8dfe9467e62cb61bce683dd927315ce136d7fb0df6517d2f51eaef754884e789f
z8d753f4eb0c798ed7631c7497b91fea9e26b88eb66ceddfc236cc5cbaf6fd7145125829644d03b
z12f1719c56c8348983ad5ad23627541a65116e775f0725e36ee0ca3c0dd571663ca2fc702a49ec
zc5bc117266944bea846cdf3bf83a80c587bfba880248576c80f25ce12eee76e6be83ef985c4140
z290bc4f7c6cbe6698329044760957b7ac29f82000a70ffc9af88ebc405987b13a356036787995f
z96fa326e32b3bc30d61dcf1e8d33431d1d484060e52ad6216fe335cd59d7ba7c589e9723661bae
z09abdffc094adc89eefad77e5bd3220b276e6dbe31a34f977a7b899a503d19f31b288139c357ea
zdb0fca07fc9faa44f0a428e48a6abea33975bf0beac46cd84af9dc8afa41c5b305e7e0569c873c
zb8b69ba227042b21a6caa490a43ccbdcce6964ae2b21261baaf0fa5219bc45d05b92a47984fa8e
z5667731ece84de9207c9f808b27eba721f2cf90563471674f1eaa4576ecc8ef253470d744b6f2e
z977991ae3e3442abc2132ed18a860f3d24d8c2a1441994b6d8213997d829d817ecba8fe87dbd3b
zeadc88dabbb3db4ee2e4b5b83bdb6d7841193ac261ca86ef4a1cff45fcedefef998af7c26e724a
ze04b066c32967c3703f464f72a6c767da5a99f2ff8f220dac6b7e4db209fd274d9b7fe40cff5c8
za95555e7809bed7cf5d4e98d3d6192e3cc257b980c2a1216116cd4e57d4a8c9bb6f7490fd80daa
z4149a4bdc32a76b100cdb6d72b8dd5a9066b8845f094f9b522f9198cbfd04e9d59c719acbb3811
zc60060489e92b163fc60746a60d510ae67d5b26da53ec901552b8ab2faea6d48ffff0ed30ff75e
ze71df0ef8872cde518ba2ad999b5b3ca3617fbfb8328085b02ac7e4b3a495746cfa303fbb9ef11
z405f9e4d7b70f89220716ec4b63e9eff0b2aced7a9d66b5bf63a3169cee62ff15f78b9cbeb2ffa
z67a97cc3cdd95ce2e1f203823e859d3759d9e794ebfc8394563cd55926c15d57fcf3a189026c15
z8d626342aa8874f63d69976807b164d7ab220d69c28066ab7deeeeda48645fb07688b18b000635
z4707ab7c60824edd524d809db4d4d4791930efb332379f4af2d0f40e1c71963e7222e81e474bd5
z00a17bddc27709324725f3cd85bd9e29400c8b754c644696f580891054b17565481db6d852cedf
zaa9b2c412bf80f6bb72623b89f7dc0da5c009d427f1175a35ec05eaf7fe243afb3748101fc1abf
zadaa00e071c0193f72a2631a3d450fbfb8f154d38fe6cffd33ed3f3ffa81bcf03f515a87536854
zb0064943b1e9710af49e437d90d3e7944bd91ff9e4d9f91c6f6c4f3b966ab42f69dd1fa403c874
z1160f3261dcf6b9a7c978daec53efcea4e68c4cd400ded23f0f2e2b0398bd555787be84a02c04c
z520da33044ff9bc21549aafa0a1ed2d2db1deec3532224042148bfd7b085346a66ffc4d6f42eea
z8a6303fc9bab4ff96be4b3c89648edc3cbda72affa3eb652a10268252430848462e911e5aef865
z545a1b59588b1ae54271d9274761c8d9ccb9cff1a9851d45b311f462a36f5373969208e1a5751e
z3865e4f0fe60c4b662d3e1cab908827d46d0f3ff25cc1ec79794b971f3b292113b0781161560a2
z32a1d1395e2dcf3df73061bf10d283b5a4cc608c1202c9f6d73d19a908a96ff2a182b52085c2af
z9c4c93116de5c3daabb6aba548fa1f79f46939bf54f77b5afdfcd0d5d28bbd7754c139c711d5c5
zfc5cfca60ec0e643ffd193b6215bf8fb7c4019cd3a817254b377b03adc7e675115fcdfb111ad48
zb339b3593ed9274b6446a146424ae37596c781a0ea2c57f26411b1f78a1de8f74357c54a6aa7a4
zd8997dcbedb1af9b4d03cc80747b72ccc48e36e5dc55c9eee239a1ef635275c6a3c8c472b7dc8d
z73cf4c02cb01a3bbfb77ddb176076c13b526383155c232f10a0c4c80dcadcb28c00ec45cba178d
z248170bfb037f6a7097e5d012303b3d5a96407a08dc2a7901da7509a0c2e99dbf6a3e0b365146f
z9cf79fba91628c3299325ae518f3e60b5348b8eded16a411937ec2e7abed900f1c56f355515b4b
z2f0bdb16f7ce8766025b384e1729a03b77947fadd75ced133d6f8c039bf7545954f874d1fe7859
z510664c0159d2c3679a3ab5263d488e6c0b850f8380b15fa05fe33eb30951122508a1c417db01f
z761e4019454147cabc675e84db3f07fe3ebfed49cecbdb84f2d6ea880fe54ba68b384bc85228b8
z965c1a945692e09e1f86d7ab2971316e82fe2d3609dbee69f8940dee6d7943372530138d5cbc32
za48b1ec5ee5a36289ba741ee4a7c5e90567b83110538c094b3e5b37cc7538e987ba78d75085e8f
z46969d58619031654b236d84e186dbe4927775d162cf608152295362a716490b8f4bc0c78b7183
za635900c83b26fb6d8ebdf2b80783b9268c0e2954ee83a514be434f068c5c678d5da7de443f935
z22a9cef16acb7d461801ac509982115fb73bb2531454a537324edfd4e6a97a13c4b61b74e2088b
z74d6cd86355ece9a6967fbc3cb077c965e91c9f7b6ff59cca476b5f14046488b1218474ca6f18d
ze32ef1cf398fafa97d2c8074c161601d55ed7764486a6acdb9c9187e46ce5be6842601f12f07a8
z8a11ab86b2401fc893c535ed6a305f65729e67ef04387859e087def3c2031e8cd1c498e6e32ede
z3ec6b82498df812279c243dff5e245767d0abe3a91fbe776d1435335a6c7e26a671038fca750d4
z0eca4990064d1ec7630f1e89ca74745361c16084f700d9a84ab0581135b7b025f3d0b344587016
z9d5ed1751d836c505636fe166b50ee9893e9120892a7a4670485b8b8a1b7d7ee9fb39492f6ad43
z024dc4367055876ead822c0c13204308a0d67522cb900b1dcc393cd6b8c0c55f66975697421df8
z898a232abc48d83e706093c609c005005ccd383122671b30306b57e88be635a5086521f4228d9d
z2f47eb91a3776f169738156a8d7685b60de26984a4ef940fc02d2cacae0cca95d679716808af93
z084cb0e56a69c5cfd6e1eaa04dbf78b482bc82a4344641ff74da718750ffd25379925d19bb495d
zda9b7ebac55798dd8c137b904b4f94db42dfe59c1ce31c7010262eecbcb7a3ed073841b0665bbc
zfb92f256d1aae8eacf2e0fc325896080db560939979dccd9a2cffb64e302b6894f8c1e7d987c48
z49e1b2d0958134769e7ffb111e45ceabb250ad2379bc6ef03f71eb6bc7503f5dfe2344fabc473f
ze80c0a4694adf8dbfb860275d31041e78cf4863abe8ca066ee010cf111f292611c9d5d456957b8
z59685058c8e1a7316f7f3ef337ce7973d2f9e1cc2aad94e57622628cc230c15acbe39f8d08de21
z07f2ba051adc95af87470ff9438db7ba6b350ef017afe418a31f62d439bc59890f3240a3f5d680
z50e4321d1ad68cacf39255ca86c6f4ff32a08798630d7d99b70cd633a0232a711f3dc8b03c7f16
zdb01e0258e76bfe7927d5b55f289b1ae88a5aacc1ab918225283bcf5bedc61adbc6bd51425720e
zb79e7c547d1faf5c1fd3cb257d4a120f8631786660939327465a3c3c880207e0b722af6870f2c0
z5e2e893f183a89332375ca79c1ae95411fa0d350b9078658ed12b75c0a4d642ce2994410c3a234
zc2cd3cd35b1b104f13b1c3a45632522ff8ea7dff0399ff6493f35214fb810ebf31f990bbb9d875
zb4ed9afc31a637e9d48993861a9347c7bfa202b828f157dc05c89e118c5c7fd81b130e116d9ae8
z105900033f8b48f4b7a5359ace4909e2133ea32c16180c99fc3124dba37afb33e935f2478359ef
z22dbea2475094afa3230bb99c67fc000fd590e29ca5fc5dab857903a84e4ae5457d57ad6e7dc39
z2c2c7b939adf016e4462921a3068e9bba44b39bc812f98af2a4e360371f45255185dafd8eec926
zf098575f96f0417d2ce20383b5891754acb32917dfc20bb29d73c7d4c3a8bc3e7d22eb3b2b543d
ze06866b592195b169a90df80688ae6358981216c5877698cf9d81996babe568c44d30e0aa12f12
zec174199c3db924e994f5692cea573ce6f5ca252f89e7fdc1cf03175813fb4082e0032068f152b
z3f665647fb69cb3a96ca0f4961ef4dd97bcdcc1d3dc5439e8bf7665e430f2ab582292a05f29446
z387753b9657aca63c28e28fc2835025b4de4e2c78cb2976b2400337692c56c4e772d0bf5084aa9
zab8310f4c5c4602c9f50e2196f575ddc19cc2464e5970c5a651ca06eae495f8db26feb0c421b6a
z3c5132fc7a1ff67c00ee1f034d9373aaddaabde80d3a2e64d001bfc3d378483419795f52c969e6
z6dc91ef00efe23ee51fbd812bdd5f5c14aa222cbb6c10dfa4bfa96a0aa906e7030d69347dbda90
z3064c5969b790e1852ef29f252bb9b3d4d994a4d76da47f480e0e1033befa92cb20122e953732b
z6d7034a2caa7b8cf301123621b7e3525e4d84f006d7d1a558d4212bc7393080e3159cd901286a5
zb883e5674a96cd052874eab049ef7eacdcd58b9b4ade6c01d60da6b3db24a973b7a8f34541a61d
za28edab818e8df731d6a40ec19e7097545e173929cd63073b420c89addbd0cd3af5e45fab4a69c
zf755353c0979bac86f007df0766678d7f94c4f6735d314409de617423c1b69dd98651310b776ed
zf13549a78353265f4c0fac9ca1d439b7348f3717cce2b0bbeda9b7c0a2b428d3971b9da407a576
z51fcbd15dd7d6618f7603ae5c5a1fc907ed30f7a5a7ff70a450c69ecd49d01407fe97aa9a0bde9
zedc3543862bd66098f19bfb453b240fa5883868c87403690103b6773d2245d836a13113984813b
z892a37da55bc7af111a379a40645bdd489938631f4b7bb4a16a33d8b606f729dc46adf2f9e31e4
z79f43567700a724404fcb43a2fe94c862b2d6134eaf80ea954ea9174f3c6be5b9b6ef51de919e3
z6e35a95e59f207dc9e2b23a9c7beb7bf7b976532c1ae5e057f870dfa140b45d80d7a16230c2522
ze18e2fc3eafef0711d16a16960cb55cc6ec57d89bfb3efbfed4a1fc2675ab1e5eff827f6a9bc58
zf2edb47010045e1f38eb36f3fb4fce5909f42f60fac7d2c7820d75d8faca6828436351b93b3f7b
z068ba222234fa6ffcc2d8a5f436abfc7272a4d2689004b5a88b4d8d3fb274d03919fed36af2846
ze59882f1afb85fa34687aedca18fc36462efb60534853efe588da2adc141050d257a81208b1f5b
zb032548be2e7c36dd205e2a4e890c89b00c5786099dfc312399ee859e8c6c93c6338485be2ffb4
z57e563580fd7512d04362292f3771de8a03b4a47f39b013fa8bc51eb45f7fc0eac353c39d03708
zb819779eb6dbf1670bfa04b38608b5fe5e39408000c213e7af0b9a9d3585ab3c7acb83d31bf71b
z9c44f9236a6787b3789761fd5246334981a0d399362af918553c6fcfd81af2889be530a93a0315
z3f193be2b93dd7697c35d1449160ea2b5e33dc6f6a07c73f033b7c8bba657d5c98cb3b4e60d8a5
zbe49a30debbad4afd99df1e049b84567ce3461966b6a2c549b0f4e323d73c3fac4abc1b64a36a3
z679a78f390122a7d7f59d43713f155a27371d2e9b2587b8bf44212d3e7d423fdd93d81d0a1bc1d
z92386b2b1616a460389a338e3528321c04bcffdea4394c8f7f8ebf75b0600ab077560121db167f
za347df69a0a87778a8793fba68b3d825b063e447626ac1238a74f51be1670dae12cfdd4642f3da
z0b12a7df016dd04425c5b1ed908f1b7a17b52c9c22ea111da7f944a0a64b41be7d627dc28ed3fc
za29181914fb07c73d4675ff95b1732dee53852924858f604bde23bfb637848bba1f5bb1ad6a640
z164342b8756edee5294e115b435f73cb09293f377cd774e052f19636c399ebd05aab38949d385c
zeaf90e498aa042f4dd5a0306a70076b615efaa3a08fada1ea2d32f75026a0c57ed6fe6abc1800e
z9779c6482a8c7f404bffa0861f7ac9b92b89ecb15fb11fa46b6f50c3dc2c114e9d126ea172edcd
zfd5ce5e4723f3cca5e98df4f5033df178e49cd82259bddfa76c7a342bfbc6fb099292564c87e5c
z93f31698057b5754b3163f38734985e00ce872076c42a5bd82810a1446019a41354f60b077b189
z0009644bc982f4d6b5702cd8716eb4dfcbf6e0e45ef25ba6b6164c4de4af61fe2dfda78598fb10
ze2a247337131b2436deb8518311a9e3fd93f31a8e36fb0d9e2026a23ac3d46002ae82bfdbcd3db
z8ad83a138e51f6d4723b032b474dad59ba41b757bda380616ac18b9bd894f61292e6c448013708
z4d455286609b477e584a868dc45963ae321480673df0d24713928445f9eee777139996a25c3df1
z41b72572dee2d4eac188995a059102f3eb504e3f485a67724e7b3a9f8e76d3468961fa26dbf506
ze17df8a42b4fcf3dbcc136955b006b17e1720383d5526fb089dd3ad5ce368b9bbf786c1252b566
zecc4c3ebf2774db94c493931a8da1b8cc94c41c1ec0055f4e7798c8c33c5eacd7a03f6035d2a33
z9a93cb7a7a28bf602be97b7f79f3e02a64300e71f67c47f1a3caaf49ce2bdfe87eaf66116c2e29
zdb903131ff06e1201ddebb9055661697adfe048b67b1cbe867e2668f61e1267d4664f0826d03f0
z6daba0a6873716d7b095780d2af154f1a3f1d9975197b6bf4329afa23c0b47e4866b1f03a71b23
z9911d8205604027a7616ef25138f7bb90d8106eb45e02980a5b18052517984de314aa1f63b57c0
zcc95dbf1107c78d958a18ee3a45ace0027825b8b05b121b03cd5c039441b109f9782d9ce1572ce
zeffc010b2d0b9016fc980bf29d5763636f38a81e9ff1d147b63b700bb64dba464d29aded2c2a5b
z31da15169348d8de915da6e99403d4519bbf284d3cb0c8a5669ef028d4fffae5b63f8a7478d69b
z72c75b5707266d515b04ec51bdcb50ad85175d2c33bcb77a0129b5a4b9c2329994ac083299f7eb
z1c6868f4aa5281b5d91a70ccd3ed66bdf5d8d2788b4b71cec9c8c39eebff5a64d8a1c9006913d0
zd19bd53ba325db003beceb6a6b9217e158549ddab3b3803fe27d62b9bb60dc8d235316a431b024
z8d1c314b1e42de8c75d686f758615ba4a86e723b495a442bf226d7a58d89e07acd1854d4036cab
zb23102c974bcf0602e6368e99ea877f0cb4f09a0b9fbe93f662e5f510876edaa6a4586250dca9f
zfc06e19bdda9196bb34be1b2ecb2f5b09d2994eb4455d5eb25022539554b74e3a9d919c094a114
z194dd9fc6f2435fa40b0f99136f7bbb9780ff1bd52ca3dfd34b4d2771f55572ab218b85d395ced
zc6f4358c3c7b320e83d4ae363e5e86253896f46f87fb803f5b7eed62480d65807779682d5ef5cc
z9f107039620f0d59b51b409646e973ebbe51d12a7ad2d193d732c21ba49eb2f42984ddee932fb8
zf158fe622567287e970842e9aa485228df208a333924c39221be43e6e8f7969405a23c8d44bd08
z81d16c7f36eaad8c6067a0c2417ea98744d94b7027018df3ef3f3a7a7f29d71003f3e64b9004f5
zb4d853e819a56e417b32b65c5bfce8594a715b56818d1c402667203d1c3e2e9efff016d587efaa
z76366b809be79655b9f60ff2b4572e0171d2e0ec5255b39383202d9292d1de15786e3df1c2c5e3
z1b5375958142b6ec62e7e0dc95dad92b39413cd4d6adcae593a7ba40890c627b2b02ab958fc311
z70af28a60e17a8bdd882411208bde546efc2cab7727b68695e0bb7cc50727c67728f129870be26
z17b0ec1399a1c511aa3932efdacc406b9d87c8832ea94ff7c90fa7886e7a3b1ed206bb4e2dbf31
z390782e434d03c08c66e12acca302538b56cbd52e9a3f3f4d45f6e8b3d1eddeeb7d5cc179f1532
z737b1c935507790ab47e12255f9ceafe022bfaa0c765db865bcb5905bc84263baa2af130ea5cbd
z0ce486128063ea9d46ba96e42054c94e97efde3fb4b6b2461bf86f666e17c2663227632021d8c2
z83437de026e01a337bd17b42878a926339047a5e48c4d977ff992be69a8329b215119dd8d1ed57
za0b9f68bcaed239beff0cd65cc44180a20e21f283abf2d61b8634b6550f1059270f16f33b84f1a
z0f0dca7da27f1bc32d42fab835e809db16820b4cedbeda60f4bfac4179c108733db9ed962fde30
z45cb0431a76c93a4fb44efc5ed1f5ec5de13b112d312e54dc63d3e73dd3de2a21cb5325b505391
zf9f03f1f4627f889020a5c02e63bd709de4891fb751b863ef8153007842cc35ddbc2892fe8109e
zb1bd2743b9f5702e21393b05dcf4f09a45971749cbf76840c918ec309ff580477b6efc30e95c47
zc4da0dcabb86a9876fb87c6dc91de1d7541c903868cdc06ed933e018d4fee34a2ede6401b4389d
z15de7835a62d74ce35810e811150bd7297da729466e84a4947b915bb210e629296781d561e6530
z62154f36f6d05e5673bf1027199d9473f5a06126197eff53519c4f9a42467627dca57bf52533a1
z6cae62f4dc9cfb32df5453331fb5651fea93c00f4872f3867c739738cd1c31b55f73a747be242b
za1e32c2b6410bc90f5481701381ae9d6f88ebfa81f9948b7778d050cf884d27ffbce84fb83629d
z80ee3020679198861b1cfec94144bbcac36d8214ebaff66c5638d71d93add5878a824ca92b7a3d
z17443006a77d00880b515c591ab0d473215191ed0283563cb2308d8fbde18a914f82c6cc8bd201
zbde744ccb3bd5de07dc80004d858769c8bb20842371cde8b2cf5a4f948a0a212b6a6c0698a436b
zf129ebaa0c9f335fac00b637ac02f9bb65360712a9130fe54ac2151cccc6112e12f7061ea324bb
zde6b3406aee952f6fdd1e46218fdbe23f65728512d93495a83f9c8caf287eaa425e9f67aa7effe
z7bb5e0ac6f3018d4582d8450ed5c25bf86ffaf596d0f83ee21148e57bf644db0f8f09428f8fa49
z2e63b6e7879b160dd11d81bf17b747f765b659f53815d33b6bb8fa14508ab89d02f2c5827621cd
zbca94c55885121cb8c0d2574edae3e1c1f62dea8bcd7bc27ef11faa6629294a0c076864043d3c6
z1410f8b1ea428a3941a92a88ced775c61442d1bfd14240d2611eea09181d0d3f5b7da4d7ebb0a3
z09ee5f02e133ca7fd78378798fbd4b03528fdd025bdb8375477e9072904f628350ea7175d5076c
z531adfbe0606820deabe4c7e43f27e3c3c841d149599c5aa0ab167414a84b5e18762f3901065ec
zca78205da53ca77a5150e68fc7013a9c7c313d2922d126ab1dcab5599d64c638f5fefadafa7346
z178dc4471d0fd5cdab58a7256714110d15d5d141e3a5bdc9b9521aff11a72c08450bf74642311c
zfc2929158b2c111c7deafd8e456b57437bdf3fd39feb08356b1ff4200cc9a0a3cefadecb1bba4e
z32f7eecd0aad537ed367dd4ae38e6be69031b05dc86de814ee8954582404d82558d85b1694bfbc
za23617f504c7767da057041ff6eeb626bcf145f7dc25647e48b9e4613319177453bfbfbace72d6
z51bf89256439de0e58230f85f674cf1a0294eb3db0312d06949cb81e98c667bd370ffb55c1e964
z925ea749142f0efee0d6f4dc3cc29a49ada73ce72c6f837a7ffaf767c0ea5b5511d2dd83deb08a
z6e08ded72aa2bd3bcb8bede461f535ac67be3b885c5dc2436405dfc6cc486b0ba2659f2df78451
ze0418b80ead832cfebad24e6ffc00a755355fbdff05674478897fa9227c342058ada46bc720e95
z06291b60816d3f2c2e9989e7d7bfbf7bcd2be9f9334b163afc239e9bdfdfb974c344e42538d758
z40e0968e35825da27c20b9020bca4ec048aa1178d2d80afbb910fb13c18f1a8d6b5c8cecdde118
z754414a85885783181a05e432aa5a146c6a262b524344045fad5e254c60d362f148d192004c22c
zc2e1b7bff611f14bd8fe867273a29a2f9166f2a317dc476376ce3c161b62e2d8bd1fa13ab3201d
zdbed0d680b1f73afb3dfa8f221d9bc8b32b6776a82084da97f6ee11115a4d7e5d7bff3f64e49a1
z948f3e348f302af8ccb6249692426c6aec82f82b7572ca4fb5a4e4539a8fd76840301e1a902875
ze5f5c2518a30cd30b106ba282c0f40252a8fa290f25b067187945a6087558fef87ef96351ed4de
zf1e8c151827dbaa8089f3dc4dc012c92d5185a635db4d79831a292d89653617d47d8076429438e
z044e3bf019c2884c27d7816361014d75842bbd555fba1850b9bb46d1b6408fdbf63e0e36846b0e
zdae6d7ba89b418a992ce734baed21cfb11c4a14bda3fa9de241308d4fd5ea9447e213531414271
z08de72258f980010c28d2920c89dd7c0f39047e282cfcb30e417018ecaa9afa7b60c47f9118582
z1ac4bd35f9aa968c324e810bedf2a4faecf4fece5afe82897407765e8adbc9148b5952bccc89b4
z0a9b1c0be61f978d44874afd346867c85497c06e7098088d05aea1f9a03d134f045eb82f4779e5
z5394c75649e5864f0f4c49b419b6a54b2e6e94d805df6df758662dcdedc2f8be7c8f40d085573f
z53b878e275111e1d3f1071fcb4ef6dc64dd55729fabdd387cf6ccc25b9ffbda5d4b0348186aaf5
z19372dcf76e3e662184cb527c845f5a18859e9150ae6111b3e2e451a0c9cd526e235ff69bfff0b
z8026896c4d05604958bf465b79f87efb3140aaadadbd4a781f69fc6a9ea7b39a279acb7339a420
z2b2d6d9fd5d0f0e2039438b951ea50c4bf9ea6007407ce156fbaff18ba6cf11bff66c8dd894e31
z51bd0549b19c04d5f052cb7d5d674c91458a2b3bb78ce0ecafb763457b53510edc5064aed01e59
z689ad249617e6ad5b3fdba8cb0831e64d3600a09fe433332336691c4d6f60a7d76177a9db4d4e9
z264fd88e669af318f321e6ded0325b18bc7c40021cc0892e4c5a286dbdf63760e80e676a868d20
z716be5e9d45c991582cbdfe129e7a43979e8cc0ce66b9f9f3a39e5ae4655dc231d1c6a7546c5d7
z34b45c1e2e8c26bd1674ff987fe95de3d405bb8fc2a8a3f3175f6fbd0857cd1a347893dc663139
z611f42dc17fe6268e71c2aee10a9e0099960af4b31d6d4c90f1ef914b1a7aa64fc598dbe349aa5
z348eb872e7a203777bf95d847d8b0891900f7ca4f780bf0e6a8a048f2d96137e0cbb015b60c145
z03a3af71922d7b9b258f2d7c45061f8c9dfbe32ff9f8609b5e305382ebdea0c9524601c8bcbfa8
zc33b0c08eb71a5575da3cb05d4999643271b34208ba11108eac1b69de2e75907ce5d28e7c98268
zf05c3b6ce79db3f7c70b5ea04f44e164f3912214481df3acf32eb3835fde30d649038b113c28a5
z605757dbdf731e492f6be7438469fa2231908c7b8da923d2521f15018226754b7d201e9bb46429
z5df942feea84120528e8d44fff1446ea9dd453868acc980b07cd80f376404e6a4e1c01d133dcee
z3083c22c0ba4d62f796e7434f6f26c27ee1e49a26d52eae256492e08a792b7371c41d4bbece5ac
z55683814373d608e5d51d36e26d9e0962a1ddf23833322222c412922e1b5d0e8cc40d284bf488d
zddc8189484dbaa7d5a5d94e9a551ccbf6b342a5636c8bcbfeacaa854db03be41d1d6ae33916980
zdd5104486da3143295b1fd3b21392de0b5434fdfd01135584cb4721cee13bb5eebd30c47d678ca
z2b1baacb2c4cabeb16304b864df9bd462c6be48857c36979f3a2159445d35e52cb5917ed49515c
z7df832180b1c3cdeeba37d6cb3a15a9b7d067149053fbf1857f2073b27067bd98f299493fd0065
z735570f580b87e1e42f145fe7d3fb2e6b58c06ced65f632bfd5ee1d740a9dcab7401899868f5bb
zb4f7cdc9db4cb177b353da6f0d6748e75d39c0334ed39515e3dcc80e677d64da8a8b7b3aba83a0
za190f45d42c92e42627fdb2901fa12be3187c2dfd20b60913bf31a3d0ccd579b47722d65bcbc77
z2fd46eeed6a3357372eddf484e1b93ece22971daddd3b2f2530ab809711c8f51a0e1457bda12cd
z12c7d58ecefc96231bc68e816bc810cb47c8b3699858d274b7b0fed9cb9ec2ff5dce1806c98579
za7a7e92231eb1a4cbbda9c94dabf22661750fbc30e8526bdecf6ff2289cac84fb2045419db3fa7
z33422eed7314871a1f1fadda53b41eb6073a4b0bf463355cce0e951e07614e94802b5f13dc827e
z628dfe0d62ce0ad82637e553ad44a93209b323d4619a119b0be57ea2f8445208443fada379137f
z635dd44cf0fa1de64ecea021e761923670a813475b14a154ced746490605a898c5fbceae21ab37
z41a8242306742c3fc3af8fb04de95f96c057331f8b444041c622d682791612ec7972cf7b60ef53
zb3f18c71114f80c9bbaa24156c4887a6cb530225c3f4228b3d8054a7de47eea14cbbb1c4d0f375
z48fa2dd26bc015eeab555e2347cdddbca9974429c318dd254ebf3b49c1957b92a295f00e46a8ad
z5f191f1872029310b9c62107cdad4f0f1b0aebe33f5dd0d2280e0dc36418cc5d7aebf67427bcf0
zdb5f5fe7188a554c7eeb00c1f9dcc943997c01a16b93555f572cbf8ba39fb96b6b965ed37cf7eb
za423f04cec7e980a62a6e5c3f4e2bcf49dd3cf2bdfed9db7ee778d6daee57bc5c9e845a4da992d
z2b0fc8b73d1ac8eff6de949ca5b46cefc3321c470c5b34c5970fc47825a9882cabfddc5e61ac71
z06c3d109e2ab20466f8d85656b888b2c84aaabdf0582104ef11d2d20b9f67f7e0df6fa7f21bbfc
z3ed075b88c0b266b41f65e0a3867559e5283b15f0ab3d6f2cfe1b70af4891fe7bfc398842edcc2
z8861ab93f9915818c2a26457392d57c7155a406e9d1c0f4e4a7aeb007f926e0050238c2cccf503
ze95e82b99c0162da43a96a774e1669eaff17bf4b44923c29d353accf37888c0f54c7931c6fdd1a
z9903732a88c70a5812316212592388b3bd7c59017515f320a9e00524f850563603075e9dfb7ff7
z037d656f7324ad172ff3868a0747d43d2e4ea919435bb9dc2b4870e5629ae1daeb5ac4594cdf72
z62df67967ddda58fc8c4fcd88fd66f1e213e4947e69beaf073383628056ec391cea084d303a0a5
zee6a01bb98a9213338fbe1ae12f85b790358bb936218307ef7304e29046cf6152f9d23f2f2a9ae
zd60fe05724b3ff860c898296aafd9d730a7966a8f5d514d8346837cb6dd6b876e868db5a6896f0
z36feefad321a9f64d8dc5d839c402ec89b9145dd8b351621fce816e03439ff8e74c345dcead232
z020e00cc2210be49c452ed499472379950fe295d2987b232ae16d63c75823ba6bb22bc3abe9900
z2234f1c947679b52a496bee981ba6281d34878c67f4d0b42625659cac28010321a3c95340dee55
z3465803183028798f667044c3e9f2f9a286fce5a5fccc98d03145fd50724e6fb9de4f390cf12ef
z04726f29ce13fdf7030f86653f00ea608d1f56b65644ee75c778479c6760fa51277cfbfc6cf8d3
z3134718a7582697cd74de51b9d99cf03aba65acf718bf9ba292b0295b65ba43e7d04340a8685fa
z2f3a27d16f1bfab30efc06b21bbaf45c09e6158246b07269a9f6008d8b315712ce869f1ff2681d
zcc5e9c09354b8882bbc9f22899462c32e16f7ee40bd70baff5975d96921fa83ccca5f7de8ddd03
z7e0fa6aacbf3a4a4f6eae2966dcb7e6472922e8aaf0c54d46c88908916d9ace52a77d1f5e610d0
ze29132f8ae01fb147278fc5a1fc7d08e7069a5d4fd7690a8036c045e4bff67f8ee424be2f737d6
zcfe24a9acbca5ea401f2805b4db271bb03e8f860fa928e2e9aece859d41a1e9b30e5d5d97d93f8
z6cfabdff9b99552add31c382100809950be0f332a8152ce4b390e5a1ca78a62118456f5982fe28
zecf0d0c0a1968155b348fb7a5d710b5be134db044c2ef6b3d24a853b19f45dd61cee94ecb380be
z9e3461034f2bbf0aec16ccdfcc24f3c5b2aef85b88fd6de403d308736e11846eb8b0f159f5f5dd
z91612b8d585237b59ea3175106e4fbfdf600c001f7f7f52e47d46d097353c8db7830e8a49559e7
z79c89af278602264b0f76c0e6379a214f31f3cfd0063c55e081e0831785fe77431c6f65e766491
zd912e36f7ca174cc4707fe763183274bbaa5416a24eb40f8455c50a54a6fbe79799d5ec20b31a9
zb604632b14221e2511132d142292b4b48a916ae33d03273e5f61339e91049a23a8f55da4e3d9ec
z31300f8f27275d34f7764dba49976211401386d1d580627da348de1037c107811ee3805295b3ea
z355967143daeddc93a21ef0fd0af8479664fe3cd9478ab007884aafd537431b01ed053827b88ea
z0bc363599b2e758735fe99373dd856fc1128f4ec37b5d9154d2058a0cf118636ad443cd152c5e1
ze9c725438dfa37994704662e9b21c9ec46e5d454462b92a24095e25d64e7fd034df213a3db9f4f
z5c80a174e985a332d83de73f00c4a447b2b1da7a0dc2f8118623e7cbf71a647f282997361d642d
z511da85ad738ffc3744f1891249b76ba8bd184ffe16e776683b7e35fbb917b13ae1ee2fd7b9793
za2d62370b599080609865a8664d7d4ee22830a8538122064370c2dc1f5a002b3ad2fe649958b80
z664d70e6898513195cced617d1292497f55577a4cfebffa0264768907ae3102dc11e128c161086
z3456ff814100289b076cb61b675196826ae90236880ede0b331a1fbc774c932c7edbb2f4b152a6
z0f483d07d265e222d69acc108fc52693d1632d1d967c3aef4123494cd55391d534a4a923e9e670
z3a8c6ecfb0751e8fb68ed90ee4048c3f4fcd2cea126c519d2a7d4eb36f38b5477f3e0fdc77ff3f
zb4003c3f1b0bd9fe0a614e36ee9008c1961750745089f599658a91b9327cde95104cceda584241
z29c521d4df88c73b13a9312bfd97fc47141280f9b5d35f056aa0c7715affa353ae0ddd11a7526a
z71098ef0e0ca02aab4217b2a73f1be9c7b8121996abf9d90f900e10021f61be9f53831d838767b
z4b55588fd4a1834f5fd35d7200c7937a54a8330a3ff98318ee48c9b0b681fd1b33d7eb6769e597
z35bc17afede86326bac118deb23ddb63f481cbf8e8a06bba1b08f8b938998d65cb6319f48e7613
zf0b8a19aabad07111bc74519795231a50c19798089fa46f4a44f9757ed715dc30db9e7823ff20a
z77f4d246cf9898e12af5a9eb1e983482a658cd8715b2eab8d4dca13d9c30ed5cea4f5a2b6d3d47
z854320e59b6e4ffcfe1679e0c09af65826097d47ee4b3ec21d6251f5ce5bfdbcd2079113d2111a
z7d22d98935f801a11112c075bfbcebad275fb78ca64bb949f0968a2c112f4ba1a97c21ad7cd6ec
za4cc2b91bc35eb82c3fe9295c42761b32644ade099b1db8f0aea5060322caf567498fe88382e0a
z4900fd5d188de07665a85184a81934b786b68b9575bad6ba646b1769002ba2dcb18e0b69ee5a52
z8373bd46d379c6aac62cf15a138d47a3ab1f5f5dced8ad16957eb5a22bb915a0ff0043a1b02f69
z0f1370fc8ebfb6fab56cae6cd13e13ea20311cd9afd104d5b6389e4bd3375078199039275a084e
z72f1517e6ecf839e639976dcd64fa2c309f78ab182a3f087db224675d1b947c78a91871d9df04d
z0db98f7af9a9fe7b4769d32ea8dffe153044c15013f26414dfb595977225ff91d1e32e6bd38c51
z3aafb2cdc7c6425f6825428ff227f13f7a1de916ebfa7235532175d2cc8eeb9e25f606451f8cd5
z530d732c74c5ba4408122a54f45821f623369f7336eb6ebcdb5f5dcd4ff8d4ad66e412f3e8eac0
z90743c608e9798491dc6b7eae4e29d225f7c40ea3516745f4e5e2bc1b1012fc1edc2aa98976eeb
z6b3d56a54aa79a7d9b09db1aea329542d5318d768d926ebecc24fcadaf9c973711f9afa1de5a51
z35975182917db34bc927f636f45dd525eb6eb0a025ab9c736d4e9a492ada9e50113e0b0856b6a5
zdd2addf86b117fbb8f5f8d86a68dfcd1bd36a1bac8cf1a539d5cecc5e583eb57c553c75953070b
z5e0d933a9b9e06b09f9da2b73ea46feecd2f21bc827b91c1e557140880e9028b9b1986d18568ac
ze1c9d87c386b023efd3a887d50515619aeb3bd4b8767a2fcd4dcbd0a2ee7fd42bf83b1e634d967
zf991b7383e6f43599c4658c73bcaa27f5804c2f95c5a694ff6a13e40e9c385180852a97164561f
z3cd843e7a2fb761f438e31f09bd84bcf1a030ea3a7c93ab539d53f508564570467faf36c04d29e
ze6bd3ec4f5c18fc94d40be57ef68d976cd4c5187f501ebf03536a50b2eccebd37cd06bacd650a8
z6b55e87eb1c9153006eccf33a90d4dfe8aa35c900b87b91bd6d978926d746922dfb62624198ffd
z32f4dbdd4f288a61f88e95e120bff6db846703313734a4ea8af8b3e2bdaf8289e88715e646cfa4
zbd059e57e104bce90ad43fbb4b6f4490cb3d92d35f52075ccbb982f564066ebccc2046e2c10671
z2a3a7a89481df3707a86c513eb8a9dbb0c76e586f086187124199830383fa355435454142d9186
zecb8d7c48ae43c5ace8e3866f6166a607023b72c3f3c3bab029fe52e8d44fc740bcc9888306736
z80b789758bcc0d6bc143a7be088ed4279914435c532603758f398839e49ceb0fdbaa237f3b50f2
z38a838d33583dc327744fc8d5ea6d1aacef37cc1bac4a23bc35d2fe5e49fa8c725b4da0b70ff51
zbb1988aab755948f0031ad4df60ba47877c1b34624d7577249804e92e66c570ab179d5ff5e61a5
z82e16813bb839911e63ce39f46a4a546afc4ce2ca8d9b910b704885316d8e9102789b55a958b3e
z48f241b0a0c7b46e7fa32d3d4738a6ce15f05282f17d63553cb0ad9df45cf3d65540b137f7439a
z92619ef4799f294cf4b40db7445a55265620f399c44c35a8f7dc419bf9f450612e195f963884cb
zd917ab0077599903df648b333613755d65ed9d9523992b45b03e8683f1fe843bd6cd9559586ec4
zfcc56919dd3c141070851eec20c652dd7f486309920244ce19dc21e578f138a6256c2104b3f9e5
ze7b765442fe8af9bc986637b72c45b307addc26afc49e392b75f97b38fe2e062caea203fa19023
z4e4b909fb218d25b4f86f7b0727d2ce5e06aa346b31c987b66da16b29574772467d39b9c1a100d
z6e512cd5ca314e8a3170e80ead71dd02e1805e0b8e8e036f63615e2a0aa9907f5c5092718d0a82
zea0a57ff56a118050e6ff5a5e6ad67d488bbea88d31e5c2f56f8aa95c9c8be3c674ee091ae01af
zaee80155a754fa25d779c6896466534312956fc0753bceae6de6092424a2316d45a5636540059f
z2160cff5a540a9bf9a0a9d433c13abf65dbb3d71ae02ef24f7adcd5d79e7ccd5ef4549b162f0ed
z6e6c9997aa0703bd34077311c0a4c8454677695ce750013813fc36c7330fad5aab6dc2534d7dfd
z0c21c378ef80d8a33e39f3c82ebefaa9630f8ef6004f267fb91f383b744a62602769b171c71f70
zb98b41ddee70b772c2468448021c2f75cdd81001080f6d5a7b313b832ee93afc9c0cfdba36b971
ze2ff679fb205c62e902ffb601d5aa22dc30a4c97451d8b4e973abe46568527e17d50c419c25cce
z92768fb7b5fefc8ab6b9ebfb7cd5f5616d6557937c8ebb4fd137d302cea157be6d203709b5bd87
z47a14886429de7bfdb4195c61019842d53435332caf52fb564bbb1b2f7f92a0e90fffc8c3c1b51
z6a3601b957bbf20ed8267dcfe512bc7d5e2bb7be06da140cab109e690b97361ce27bd10fa175a1
z05b038231c9d2e51a8eba5ef56b6f9bd085542e89c9184f0a8468c2721355f1a13378df81fdc04
z25688fae2c2f0c863df85b7249d22a59f8b740d268e3decc764cdeac9e03b9fc0ac6475dc8843c
z2a3596a428ee987830080ccf489c98b2d64bd24ce23b3712534deb97382fffdc09ef6a05331427
z86a68b0d7a40c84a359f2de763f53a58d5cf78f45f85941fb881a1ba71ad9104522288424efb0a
zd4b75a71b4d52e9f611ff04f44f72c61365c6f6812b9bbcb70270ff7dffdb22c180438a30673fa
z3fe53829ec8b60536796a4fc9487e2275ba351032884e67d6f94a52c74e21a217847f60353f144
z1b8a6b16da68f18a3e71e3ee759e117c3a056610a95d0423d1dc8067312742b0fea0ad2f51781a
z557a318616b3c0230515c8897152e1bfc44d10b920e452dd40730fcbc58480c81d82059eddf1c4
z67ef30e7d672fb3df2de3a8f943c325adda126e620ec82e528002cdbbccf8caa326052dd46ae95
z9dfe02b08c732d4bcfc9c9dd492270c37eeba4192b61d561a428bf0ca1520633e33f5cbcfd2359
z6938e221aea0549779751068aad6b88f62ff75adf31bc341b85ab93b07548a5732b0461bec1331
zcce1861479a1fa12b52ac76a0d5c9e29461305e1f17cc3c0566ca7d2efc0a6bd7d372bb230d53f
z2f4c21ab1e79db713f8690c6b9ff354e18f1af839f2fa7595b1fe906b7d9a45c7aff1dbb33a02d
z749cdec33ac9ab395942881ba5e8ffe8b54e6db1b9ba5040c0349ae4384443e968114633820b39
zf8efb35ea4e9c04bc9df507d8cf4fdccce88c53a1843abe26ed92bcc7a37e6c00f049dd6ae52f7
zea118e6b1e1ea2811390ae915513cfa2e6e41d9418465687c5adab981a10db7557d0f0dc179b45
z01321805c96ef73e67f06a9332577cf824bea3907f24d81392c6a66c060c572ef472c8acb59a49
za6f4b8ab7629c9b6a148055f2d6c5286b28b8a32a18a59a73a73f3046f6bc087fefd571139a65a
zf84e66be37133015411750b530247cc9240f142b529d6446d7cdd79bebbef0ef92f70a25967c70
z7fe3a21f11ba58205f98d92a97270b0194598cc6a8c76919cc70188ef5959bb3f54898e4b43121
z77479ad23987f587ee5dcb64a197973df0569892618e8bb388066e1d58fe458cf5d48ffd502066
z62c40e62c87837a050f297a6ade70d8e3a640e93fa02d0a5880295366940d022b7caf7cbc8b44f
z577388628e02d4a5ddeea7f5fcfe52c9d021d878822fff29d3337e255df852c682d16e2f7e95da
zce438ce88e0186cfda174c46317ab1b00d23fe0104d2cb061c4f4a3962f3a7dd0dabd87532e8cb
zf40d6bba869bd0e2d9ac1516003d3f38fa14500b84566332646dd6a4e5a910b24ab81420c27283
z4d74cc59d4667f90f9ecb47b0d0b29a558e3204be714bd1d60e8ce70cad87bf64eb27c60548c97
z39e1a18c50176fb62a506d1b6101e248472e83a10ff44988a92858585403b3a11664ef86f83640
za66b1ab42c4ae16a458374187e2412e05a833363a615263aff1a7a9979e36025f2c0dfd3eb52a6
z2e96a66f3b2806408590f2fbcf7f60ebef68e12dab4adaae0194c1c964f7a952278f4beeaa114a
z3329f03067a95c823f98add337b795f65666391e7f8eeabd0e360bcc4dbda64d7f7861ea723054
z135954a1ebcc957a47cfdd42fa6fb15e9bf74e7f166aeb9892be3c9a4e804a17d7c2a7eb81fbdb
z391572b2e6962e1c8dc8a07122a10cd4b336d3f2f7c684cc42e0f1d6a75f0d14a68ebad9ac2d18
zf0b47ff5b073a1bd92a969a15c379e6c8276de940b71328b69d17f6908072d8354eab4f3612b6d
z8af1f4a2df6530d5db6c2a038c1abbf0f5139ce879bb3ef76d3b21e3137e4b779609aded55ac38
zb4d723686e775b0222292ddced2a0e40895154b88910c5043700e988f1ce6c46f97f556c1a63d8
z8b675f339e7a59eb7a0bbe8adb347b61395759103713d3929023a5e017df000f65608541d3db2f
z6e1bb0ecb406b4641166ad7fa77addb2b4491190a48396a7bc637a3b4bd28ec3e11071d1ff3f83
z8cd466ec6f3eb0c4f417eeb98d604acede53e118c6386432035881cd78dabddab35ec4f710a72c
z6525ca103b8d03068b1678b5d6e028f9ef3b629d93ff948f6f8bf5205ab1860e29968ac74cefdd
z803834bb22e950f43ddaae3b67f80100b6d09b85931a0927aeb033953ce0b04435e10c7cae4fca
z897103d73ae23eb3cd3068827b80bfc4cbf715b8e6d0a9c277077df5e00a91c75cde86488113f9
z7963758136a7d83d1e820d130e513e2e79cea08366058b819e8bc273e03cc78b2756b56f24be9b
z8b432d5b014309021303a40ee48fedfa2da1acefd7e2cbd5c357877dc5e9c462779735cc5e1cf1
z86353b1910d6bbc0d80413e74abe36278862c6a219bbd8bf3914fbaa9538884fec7966821adf39
zb29c5664f6cd4b448dc6b9c767fc2a0acbde8dd6800adffe6f54aab40392b569e255d99385e611
zbd8ab3497774e34e1fb06d0741133262990e9c94d9efce47adaace93859c565836c54f813fe433
z917178662b339743df8d9c510b67fca79a11dce6d5d847ef2446a32b803b06dd3d351e143028bc
z0a649da8015746ee0a0fcd5cfc0c313811d7cf5b433d93ef1052e5324c56ec294b7c991a6b21f6
zd5a729d8ecc95becb6f44a1a139594aacbd7f0c88a211b366ae803580ce740735d3c3e5d7713c3
za1e8b2d876b3b1080e818a9cfa5420a84d7586c4b1f9b716b8ac17e9bf093dec491877bbdcb0ab
z910d2729e45121a2849376a8205dcf17d598541ba6323f6594cd40818f5f93a02bc99b3d36dd41
zf7ac3f45c23fb0d13c55f84fab59160811f6a25c4f1580f313161a497bc02e329b2e07e44c7fa9
z77f81602e81f138447f3ab9d8cb35991f0fed5f14790dd98270d28ba8013407f55254417ef012b
z595a4e99d33eed6fd8031cb2484e936d3c568fe90c5e736412b2027789dea2bd4dd3be53a29c16
z014b22c481a98e000683c4c15dc0dd4e020fbc73c9442bc2be7ae892251d0d2c994114beea6f01
zbe05b5785116abae05b3ff96bc2b06bd138ec496e1cc9ceb598a0f35ff1df99efac812b9601666
z67cfc86395253950994119175641e14f91869917a24c36572b2022b9980f299ee04fec0beb601d
zad1909596afe64b62bfa217d81478c1f6dbcfc9a1d65d1829ec709cf1b9b86c2f94839f1f502b5
z9ddf65bb569b61bdbae285a887a128788ce2d325381e8df540603685d072387dccecf9d339b573
z56a711da3d20cb3ec67021bc1f63b78035a4ba2afe18c68aa94e8506c4c4882a869f94c7f2035b
z73af6f42207d0384ed642c475da1a1f2f1b692dd729bb45c9d05603c4ef3dac357eb8675833345
zbf7319770c3f0059929b6c786d81f392a31b8020b47fd1f1cbf218118f15efb781182ee3d609d7
zd73d47be703cfe8260f082345eb81a73a9030171bf8ef31ab7230b1af9c5ba2cfe5f46b612aad3
zc9aa5b5a01dcc6213d44fbbee20e8a78d68aad7c185d0c11918dd27a6cba9bad59fc25a7d82b74
z541c319687e85569d6e4248844c0bbfe71bbc926e5127b1deb455b5bc8e2d3afab222ad5761dd3
zdf696c8e79dbf5b9f1fb4417294707539c77a6f7920ab8d5ea0b049799c1efb48807096b1f2009
z57c8f95dad8a6cea513c8c062c65a1661bece452ede6bd317160fa970a79bd6ca79760e2fde803
z635cd5c75176874968c897e02b2e8e11b0d3855a802128b1b15e6af450fd0a2d587f8a53f07c75
z59d637ce1bca160129ec3fd279be9f461d9f74b319bdc8df50ce478eb7fed86b29e86bd75b9478
za972a181093f12ed0af363996dcd53cd9a7b4383a3ed46058d52a70f4641b87d6ca307a51839d7
z4137a6ce998921a3249c6aaf79a310a279c87bb68071a3d8f7733e134db0292ab5253798efa50c
z0eeae22d8d7052961fcb263c51ac893634327ef73913b99ab79e8e7b76c741027bf280a8a07421
z05e86ca7f0fe90e0c949579b0c7377bdee3cf8bd2afc04fa59796a752a211a4f9e71ecb2425e0d
z036e4beef2242c68cfeda3ae4602b6116a520059c7b06fbbee6acbd93c06128ccf3855dfdb2fc6
z5237dde7570dcde50c841904a687b9d3eda845db0ab015f9ecf32af97ba7296deff6dbd9311da5
z954fe0565d5b2d232f3c0878dd157898533202c5f160908a7a15881751cb9bdedc9004a660c77e
zbc14a58449842aca451eecb4ca4cc16d5966ecd44d99da691cc1c666d6d03c2e2b39cf55dd9f27
z464507c6a7f9eac3b3de86923a8d82aa1b0627216256afef11d961dd65cdb9a5c101ef2f159f0c
za3cd647d80002bcb47fbf3fcf4efb5500b3e9911df849eab545b79a55802ae562c8a390e91412f
zc09f7ba8376003794ed8907d6a4026b1525cfc17c10f7f90c9c9fa5fe3c27b51b805fe8a557cbc
z8519cca5866981853bad9a77391b85da6d0f5ee9c6dfeb53a0035bc4e970189f28edc2c57105bb
z7cc321240e4b3499567c6200279912dc37c34a0983a556d1f70c5d8a92dd034dcff91f178c9704
ze4ec27ff171696604b15f5e20181b78838b6facc57c1de51daff7359397e23fc05af4fd203ec0c
za54fe58cbe8d0999939a4ed08bfd57c913686fe42c3641de37d6f53846136fef4c92c921fb4908
z182f097fbfb4acc9d9af33cdcc75dd41f2b216622db42551cc9d436b3e86231535e73721eb4598
z2cffb06bfdec04c21f84162b70811d18300ca7293035f4e227375619ec6c5aedd043b932a811ee
zd66bd4fcc10c8a84cea6c1f899adbc81e0fa3dc5100ec8e5396460a6b4f92473c037acf6b07e75
zdf57850e117ad7efa402e830dec3008879f0c32bf6282a15793508c6df3771b2aac0a6f6e691f1
z11a74284cfece302d689a8e995ca07c6fa98727923a23ee624eda82f06dcd00764efb581a2324a
z5687582cc234ea014628707261e1f9c38a78057f06fd2707fed92108f39e0313e51c92c3db77a2
z849ce34b9a1c87ef42b6a7f1ca4749f8f55ac01b5cc1488f4e61f0888eb2d0c12ee94e9afa0860
z9a753ab6ae94a251c1a43a152f403c72170db5d0d834f24a4ff04a9c185f4e9ea9a7b7e71afafe
z2d1521f7b830057148cc4ba63cf09a9fabe9feb9011cefdce06edbef56dce75ff5de130e723754
z03301793d72f8f82e667dd3b8c1882f18e46ebb537c4cb844d3df8251be47b4b2395ee17561f01
zd0384064bded6ac3a51afaf03a0b4585ae461dc65c2f35ac41ab93b5cb09d808620e2fef176c6e
zd5588cc99d93f7d5b5975214492b2084ee27cb4d2b4a8cd208cab0c866db17cf273d3f57020a95
z16a8609f4c1ae25b8c4fd8e29eb058af81f935dc970fa73d77638638c8766a0348106c0aadbbac
z3e5ff87b00826d5b57f68bb22f19b33bfa17a448a5fd85ef937bb028f8474502265d69d18a58e0
z496c7bfd801f3b6bde36f131336c217e8b68abffd28fb40db8d277d5c6ee77233976c5b863feac
z2550a08266cc44436a000b1b52c98efb17a6064735074616a08e71e3dc4c81511347a9eeb136f5
z0f729cd7358ed59b117b3a443b9d7103ce5e82f15334fdc0c954dfc1cb56267975814641390e2a
z8e59ec44b8cf3d24035dd1d3f2051742dd9c3add78acc4bd987cdfb38d2e64a141adc684708a8b
za75aa0e0af9a11c6878bee8249feed2129638895a016e707055a147c89ea4f8955130d31160012
zee952495021c5c5d6fe8cf3ecc8c740ad91fd67d1e0b79a2190d7a141e159ff6760bb263bfdafc
z60c73c7def6e867d5eb2f66d437a6a58643968b7d5ab585e5c75114261204f7fafcae86ecbf2a4
z8629c1abca17166511e0ded4206045c46cf960b7c37fabf87a082e178b2a023e0004eab920fa26
z23273f21707ca4c5a2c6c48e58b98c3ada02a742866f56bface9b4976d5b91662aeaa2a5bbfd03
z000de656ae6cb50c9011a8f164a99a56950620c84f6893ef58bcbd3f1c3f5530b1e733abda1089
z93c2d217d05ac3ceebaeb092720ede5e13d8c4ee2ab516ff3e6082b971d5dedd8f8406262c8068
zfd34571bb5988b9d0b93a834ee243b9a33bec4deffeac282e3b0bdf7210e49f1d6d2118bf65cec
zc6292742ffb99beb3f30d70ac8ab8fce22e7c9e6f5b8ed0a35028093d6b10949f2a3967bdcd0e3
z8e9dc202004cf49ef3ff48b8eab112307003fe1c095ad622fb851faeb8ff8fcf04d815f6a242f4
z518011368e9246b48848a433931c4591dcb91ccffb98344a74830bb511e1ca62a8b6e3877eb95b
zeb72411fdaf5eea4cdcec8e5272380913b1a671ee3139b0c04d7cb1846bd3a830fdaeb47946b28
z545d0150517aa00842177be7c4cec452a84f72448af9b6a2335ec08c4fdd391613cc7af7d8c5ad
ze5b2315cd10e53ed509ff962665d49a0fe9514a32d53024b9acbd471b896aaa19d3747eb386bbd
zb70cc81047e5bb20c1391c00944a008da5779bc6b37c37d6270bbba5000b17b7a49e38ca944c76
z5c344281d35b2800c0811dd2ee2c035570ece5383b9290a5664b260f49522819ccf81928632305
z3e3d8ed555b68f837606aaa6017e96d111d29e68996d672ddba2b605bda37da314ddcbb5710501
z4abe8cc6178b970fbf79d35aff09341c37210312fcb432668c7bccab6c70f17303bf28546601b8
zb2e405b448861af3259e377002c0ac09b71a74098a58a7aacb7aaf570a28ddbae208bfd7009f96
z7f5288a310b17e2f723e3da209942e449b565ee12f52b2fcb91f2fff28b3ea2817adffaea9838b
ze9398a2619c8f46c8f73eb588f7dbbd1a3b430d895f16643086109a3f2ae760071b978bca770c7
zd165fdf76261b5cc13247a27173cdf9cfffbcc651a7f80e425e1fc65ec37af859a465579eec0a4
z12dfe891b7f3cba21c7ce89de10e9de251187a79d552b80cc347159d7aaa8bba63900a1e934d2b
z92e26f397a7230217467570a928cef71cb09770bd5c4234a75f7efa36046f4499923442da263f1
z3e2c00e7bed03858105c177f986d83eeb8a1ebfa4bde68d27ceb6f6a0a0303bf49e89b7605a9cf
z54da1e7c554cc525dfc9892bcf74636b1c398f2ade3271ff2ceb1dd941e78e5bfbbbf3e02f29d4
z6ffba49beb245df87f679c4e42cc40880b4738daab382932adadbd8c2eaf38273078f6551633f2
zb1cf0738349a0f8611afa21fa972fb03875d3772b143a381622d98c5e41bcaf52f2bc3ed707e42
zc14e9d220b477a556e4910637a1b66eb331a1868992ad9faea7a93344f37afc611eeca1e27c3a7
z03c20a0266fbadc9107842a1acf5d591be703f6eed3a8341261528ee2669cb3207f4e862d86072
zb10412f30900d506e9727220a4f01b41a10f349a73635affe082ce5cf5f84a4a85d8f6dc6fc2c5
za87360c6bed5531883106296e992eb022708f07cde18ba70ce02722815a574e117e21ef60bd600
z33f9a8004ab9be10ee7f79cee09d1ed5f9c72c52d368c161ab6a1261ccd40faf961da3f218f308
zbbfcf53fc4b227f819ef8fcc705cceee10915c8f441e6b9f85e07e54ea108d178dffec81104477
z0ef2a2fe8658cbf369f47db850e63171a2c9c7b2a4d3ad53910d6742e4f9fdf58ff4b658684313
z2256eb51ffb12fb460387da10217eaccf321b43a143bef11d1625286f68edfc6b2d3b6fc53f26b
zc507f9334af50c862cbf07a9bfe295af85500d60f3bc95c71357c8c3567761076e8b85c9f23ca7
z9a0b0bdb6a9b4ab869cd3d649c86145de8609cfbe642a35b7130f80db0b39d41d44b1869b17a2f
z8cf41c650a51fa0bc247bea1b011e255017f300f3e16c35521e76ca05f15bb8a70d5f105a0caac
z04fdaa092d4bde58487e3ccdc1e3473c46a12a7c530b7da797caa026d0c35a504a7f0813509cb2
ze1c1af0c5cc8666839ec4587b2c2bbef8f30331a83a0fc6eca8201be19a20fa322dff300e82630
ze29733e2e0ea57eccb2a5e3a0317c3ca738a5367585dd0137e32dd8bb97fe5a8650cfb9840a0cc
zb5d05e3566e270b48fbb5454ebee2ca02525d2a2824fd847896e63557afa2a9bd8ad3a2f84a24a
zb2444ba41476d520b256ad6dfa964f7e232d18868c024ea0f497cec9d5a1572484a0ea1133d4d0
z4963433948c6e21c178c0c8548ddd11738fd2cdb58447b36d400f5f236255ec09d55b75238a762
z0b9a10c03d17044d416c407ef6be97604fb412c6266bec7f0bbad56d27ef222eac417d8baef8a4
z6dc7e2c85208da780db80af1e9d3c24730c4f5ae211147f3c4fcf9f8cad4840031447f753fa7d1
ze74197a1cc8669b2d02fb049d5ee2023dd33109d6c551c4e91a2a6528262dc6c85811bb0953c2e
zd9f4d6338721750d92b2b21b73b0b8efdfab54b865e826f931dd1fef314cae056e993ff45618ae
zecb090c5c26d148419ab4c1fb11fc13d35a0a225dc91920797e7251e31388b762f985b4550367e
z9043b159b2b88273944ca10eb90de37408bf6faa3ec5af39ab5e91814c68890bb7bf272450ede5
z9f9e02479b2a1433361e0987b129bee07f50135007506a4973838c0115abe85f78a692f05948b5
z1960816d35730c3a279c59376a3df50845b7e56136f34f12f90a5fb9d8363ef0b0940541dde79a
z62be241ac2c70475ce13491f4b5d89885058daa284e243d13ee19585372862a75dad47e37a9717
zf734ac2e6f965f84624a906714d8ee8c6c1b5dc394a040c975d52cfd0b8b9920d3d2d1fadad99d
z5748e7cda423f589a504dd5e7ff404b4958e6c75bde49f59f3619a83a4fb7458a9283d483e4f6e
z1b6de1a0e4265e331fdee2a5e33407d98a23e895d2aab5a8d8404cafa86ea79eb23e163ff5f502
zc3225ce73f3155a9f31f94d1b94a1cb83081bc96e0ca0946f0c272ab68d89787a64cc4301567ba
z0f894f0b91aab5f819e10b9bbf4bf8e9a0484087b1298c8f7e11e7d6b774b2d38ae911ea7a05ec
z9e8a2c5e48a3d2586fc4b88327271d340168c206cdbee44b5b52cb851c546d3e942318daeba87c
z9b85575f29d9ec26186b992b0237754cd67fdf6b8629a019322024a7110b7133b9f2b8f089525b
z72d3a1660632825ba098f61ddd86171e0cb49f6c22caeea87d61079e03ac489190227e0605f17b
z380d5bf28af1c87dd0ec28ea1fbe32d9abac96063e704f10c008663847247ea6968c1b5e9ff403
z5f4f09cbc59adee8b2055dadfc6b1944d59d237ad8f791b0d3ef2e14f8e3d55aca25a4c3cb6b0e
z1aa3306497217916df507e1292b182324c850d83d580a1c4c8fc485b7748196fb092833d6bc557
zb356647fed28346f3a3a17929a73845c376e27c66a462a4910775e78b9732945151759d5dd8f33
z0e4db614771a6a9e92e14fd7e785ef1afc5db3c0b9914267ef7a2faa375cde78643531db8ea8ca
zc8dbbed879556ff42ba10f3a74dcc41e11af10615e2e905b5f2658c874b1a09a9cc18a70d6fe4c
z7affe89d778c624e7ebcee8528f83d9fb341ecfe9faa592bfd730359f9a2a548d89eaf0948db70
z18170353ed13094d81fcc9017eed0a824ccb992ab7b857e7d1e7eb81268b153a381f3e7e284242
z2f5b5ae372cc1e463b85e3a3d635cec471ac78d17b87d23030916588a5cdb6346ee0f51be84a03
z918b7c82b2160ebb72680281dd36f3d84bbfc34a6d7a23d6745d4e5752729397b7d5218f1450ae
z2c0d4fbec3781a86fa65e52c7bc8f5bbef6784b782cb0b6924fbbcba81b0c9ceaf45890535f47f
zed5ea8a7a1d353158d43085b5d0b69ae70f6ad209cce20cc28d5b3e6c9281bdace0ce6986a825c
z561f2bfcce3398512fb25a3ec66c7529f74d5a3534348fd07e57804134152748689319272a9afb
ze0eca0e0b93e8d23da4a4c810621374e9ffd7df45e575d6d4caa99f3b7912532a4cff32aed99c6
z66b234e97b13a8732cd5f7d59bba5ad7c721edd06f902f32b9db941935b8ecd1fa268d1aa24df8
zee1edc320ae83e1813b768a747b7511e7b475bcdf4879706c58b1866e1e23fd913af0dfe4a9bd9
z3d57b50133b7e1e4299f3934d260a003f136d2738feef730411ff1cf82d071264560305047203c
z6d7ae3f520458d1ffef2597a802d1459f0ea3b3cd14c3b18703ee9c0a114bea8f37b98465bbab5
z62c84aa69122d79c883c83d74d6d8f05500bab38c9ce4ac0dcb5259fe5d0ee1bead7a9b2aa358b
zf687893ec6fd0ee5f4093c362206389664233752d4a37d796bf798446abef83845947ec9d43723
z4552371b01a9b4411187410d69bc264aed8201087967693ab9c9a341c9c0adb116762bb1da49f2
z52f3f24dc7ad9997fc6e7146cfe7564bc67189e924692b424c861a4be6ea34df049f714ff6fd3c
z48a25d67e5805e91b51e0b66dcaf25d55e3a3dcec6c619b6cf872d9255045939ec827796f6bd33
z082c35107970fb47cd63cf0a51e22b44e1b6032e70ecf879fff07094362f9224dca78f65c88dc3
zbe8deb916c8d22dab43de52b1561da29fc3f27de0fe94a7956c6080aadc0d00c16168ef2bb7568
ze3d2c66038345b0107c69a671037d248d198ed720a429066fbe56b138c3fd7927d9b6a49c67f7a
zc998e73dda2fd349746a991e5673c6cb88b416d89bb361002e8e433e3c401db961120c7febc3dd
zc7871ba23f2df4a07dd24cb63db5694dfe89fa16b45cd3104a37c7cdd45ea066678fccf4693f5f
z98ba0554821691d8c7c95236b069456acde7b9ed5d2eea05a4bf1a46a427dfb28d648b60f1e6e6
z3abc64e0d8a07ca9214f409c94e6773a1817f9d70d78e13c82538e0a563356d7f4e84574a33a23
z22ad25b729bfb4f719081ce559e6090616c67086a3d5ee4502082d79e6d023c7cf69c49afc762d
z779bd76c729a8c7dee29d52df2222af22bbbf880c68c27dd5ecaef559df0b588468f342022c3be
zcfbb683af550cdd6659f5fbb1636907af072ac94208ed5c11897ea6cb63aac6d59963daec192c8
zd8e784d7f72727f425eb50c28ddc8c3f0afb79cd8975b95f5c0209117a7bd7c8b0ac5ea23ad1ab
z362d32404aaea5fece8debc85aff54f3395369a061720ed0decf9c44c05b261dae2c5d069f3e6c
z81f948f0856935a73e50b5d17f4bc7501bec8d7a3e9968318c137dc9db87a2ce9740a52971dad6
z9935afc1687859ef520c26dbefea0fa4d6c5c3e74f4e93bab50699b0887298fd90df152239c9f8
zff5df1f30826911b07cf8613da92dd2f0aed0deafa4b66c8fd1235588b300ebb1aac07e4550373
zd8c06e8893bbe31ebf125799b4c8f7670e2ffd1adcd734b2ddf02897958ce1854ecaa18fcfca21
z24bb30b30bb44d4295d376640e4d6faf1c032aa56598007844d8fd34d7d8d8755e15d2996fa420
zfaccce8652056b14f033d3f4bd944e9f1c382189cbec13fedacc15dc9fe0632385fb0216b4a7a8
z3a997926fb6aad8a67d3d38670c9a8a00d44b5c1289234f915a4035ed5638c865cc98278e89891
z6d07102701a0654456cf4fc802710e13d8c81dfa8c7f14800f2429f48ebc50e307cfd764d82d1f
z6658b2eb8eef5682b1bca1f846ce36f1bbeeb46f3aa3b9ee5a0420851299232cae339fa23a102e
z2efd0c2542d8343f522244e7eb1ef1ae3a7e20df04e540d10e695756b854d7b26813dd965569b9
z84ecf6b54aaec4906a5ba9842b2af92e446a17b612e463c9d5ad3514733cb02fb314e147eb2ba0
z1e6934e1fd1c4a81833afad6fa4f147862fef29c46118adbb319a9d2229e98143164cffc85635d
z02e6ef51288c492a9777347f9d6b49714234f8df89276c48f39a36fb9c32df5fd5ceb596634e48
zd968ab3c1d43d67ae817c8e2aa8d4a9fab02a97128b6344f952d957c8fcf83d87376441fe378e8
zbd564b91278753334712fca85159433eed3d55bf8259ad5fab53c1bbee0155edc81b451550fd6b
z4e4b7a0ec933ad7524c2863f5019b9aae2fdab98e1ed428b0be79edc034bdd20a84ca47962b091
zd09d1742563cf2c575f2469cdaff25c779f5a9f386a01d12c22ed943c1f6376b8662de0e8974db
z1eada75e5431cb4eefa4c838737a13c36549fd55e04db7104ea0965da634dafaf1c5a06287a6e7
z5412995e3d311cc2ab1cb2ddb34ce0e37c88787562f7ab46d0add41ee8eb2ad0c2ab67e2d0468c
z09050d437e492c91cc065e7e7824c8e987d1581e76e7d5e8829a60766cc3617e301c866bcbbddf
ze6a31dd519b36ce3e5ccb6c6bff95ee7f8c6a8416b72ec27ee3adca9ef2fded88630ba1847628e
z63c50c6b87c5a9a8922b9bf43a3e5ea155c79b7a7b6d7aff14524ed71ff4fc7f810f1943d37c8f
z66ecae6d4b1f7d0f70888af7d4a442b04f743fddefcd5b8093f24cca6dbc1b1d98b79a79289b6e
zad945ade96c2cf752f147ee17b9311f81a11ca84d5290922436a07d316dd6fb76b0e6821c9472a
zf443cc22472538809df5d9481cf7460edca17d210f9f621effe993aeb2ef9417035b010bd5639b
zecfd0cd66d64d87da449e38465edc8954839e09dd3fef667370c89b1b3f0f967eb8a02a3335045
zd3d490d62d2360ae2e6cbbf3832d62eaf2990cd706f94306f4e9c39a3a1c4e3e20b4b884ff65c2
ze23f0958082923ca63bc2ad1936c0f11891b9d520dbe220cfc65b71b0a422560d0085afd048907
zcbd265ec365e0f23219a1709ffad21c2d68bbf78039f6e021d20c1c591bd1f2209816a6bb960e8
z4d8ca6e9a2e7d706197fccf9cc15b35458bb267023e84ad20e657203f7c27d7399e7d112cf374a
z5aba159a9940bbfaeb86b4fca1c38465d1c0df588b469a0d7194fff49362652e0707808c8ee7b3
z31a53465847b1dccbfe2d1a2ce006b4db601b074dbf986b754b4a344c603f7bf76b47b59d225b6
zf9efe4330f466adae086c5c44de6b883438c9a0aa6c27769f15347dac546b8b3a87b28806d3973
zd1016bda4f3546fa028af45fa2606357db9179093579a2d39d72a1103c3859c6f77f9984b93a5f
zf94492060e1d9fc098e44edf29fe3fae4e22e15b1859252842b44f5588095285a0f8f15cb55497
zfd8348d80266f0cc4d4013fdfd0c48e82db40d9f009c3b00ad6d548ca5dac2d2092aef44314c49
zddc4fa52aba1ff14801d20721274b2736e1f1769284267a31eb57f8bbb4737a0455e6c01d1a810
ze13ba2389ab854a6859337997b600809d532934814568d2f932c7cd32fe8a3ff9f42cfe5620a6e
ze2965a33ed43f45f6b42b9da983646ef3626aa4e7af9acab987e7612714e638afb9579eb5c37bf
ze06a36ddb2ab1d40abb4e44c05463992f2f7e77fed23e050f0db17c43370f5f91888348bcc067c
z59ca4c0617b577ad6e6c4a3dae33e180fd03bdd8522d465265f33c78fec92ded113c4eeb4109f6
zf5e2b803c95e9f3e67cdefadaf737af8df24a5c4d42bac0595f384b45326ea39b9db461cd28ed4
z6b50ab0f0e0950f3b0c26b5d8891a86bd71c2f5e040b83f1f89051d6cbc8186db4255736d94d72
z0024fbb4d1bc4de8c9c591ab0e65f9895cab69295fc48ef99225d4438b79845c39876079fc2267
z3e84a2055058ee5df52d9cf8bc74d49dd7e86b88d6e77e6f7a633c465a75041bddd198467f68c7
z0ed0f82bbe77919dddaeab9780e0dea62bc01695ea19f0ddc600497fa1284313f00ab2d35ce792
z131efde79118bb826ff9c0b9da0257b72d278c7fc4ce5911711a60357d7055b50298d549bccc78
z55ebf4b47f6238a494103703ad0489f8ee04ba899c5f81e543645b3e082beb8322c32cd7cc1e07
z156fe593f54c2984d9ca74d322448f20b874c99bfb5d6b5df619f82cab486435ff4285543f35cd
zac6f215d2db2898415244eacf88f46ab96166abf40e0376145ba3963300077de05116429d75ea6
z60214b0930d8ce882dc643d8bb65192cbf9770895dfd1a956eace352ef72b6664a6862accdd5a7
zdcf8f172a49064256ef13d1fe47b89bdf71dafebf87920c96289c64c53a54522b011e338eff72a
zccccedad61a38ab021939f8e32f3dc1ba86359c4919dfb7ad9abb9491aac044517e360f982a0ff
z22d5db8ff008186e4fa6be44724fc3944b39c0674a8806d07d901ee8cb8f9231b2b948604bfedb
z0e1bc59e694417c2d876dd08b8644818698fe6130ff17a9f7fc5592614d4e6fb5dc7cdcc873b9d
zad19cddd3576bb72f5e058c5c0b1063ff6acd252de37a7690228b8a40ac590d4d1c8b7a6b10482
zd43ac5c539c455357501496eab423bf6b876adf3f0966f0f8ba2653b15d85182c810d789161c1b
z5af5d7b8d0fd06493b886217fe8510623a7b9d2a34401b428fb380dc63f88f2ca99b8bb4cbaf45
zb2a950815d3034fcf05fe2aded8edbd4c969d7d70efc04120aab6b49c496f46bd74ba07eb36798
z59e1b3898b6c7dfe7f7dcfeb316dc7e00540399e6d4ddb8255a95191ce5f1f9c747a9e45b98f68
zf7740f9f56d5d92f590db1642ffa959a1bce63c3bdae261aa06051d5ce8dbdd61db3faec6a9bfd
z738d6974d4c302a7147260cb72872a9145843c2e20eb3e56361856bcdd2e76a816488607018c37
zf3a43716278d7706cfe3f522a4b44bd40cb9cd9e7f176e5fb38e1d01c554ec4920cdaf026e85be
za70c9b8d666888397df3d2d08c86f9c3240e819b3fb6ff296725eeac24c9cf2e9c8a7641290c71
za68a9b9dfd3a20fe4927dc26675175ca23348b811922a8dd1e700cf37a9cff30855f0d13384ad6
z3831eb62a69945975739a6f636610f9eaf2e35c00a210e0e067d7ad9d655c47b62f5b839edbdef
z0d2903477d45d5aafe6f0777100851c69ae9ceb66f26996204f6db0f2259e75eb83f26d0470b8e
zdf243c46e627a91c79bda138375ba9a0ccd1e99853667ca87b7e68c5d052c82fec4cf011ae8caf
z5410f96673b4bf1ee4b98d2073ff71c7391943c4b0d7ce30f782b8abfeb2371a0899a2a8a46afd
z41cb2c7bf878aed62afdd034cece5ed87ed5fe59cce36a437bc3de39412430272712f2285e93a8
za1b8c150a70fe281c517d7c7329334e00ff1941df72e55847ef247bf7f5c8293d024756f454d7f
z6df36b9cf8d5c5d64748b081a0d4e2550476e82c8b434803ae686be134daef9d92774475dff474
z64cdf60b1a21edec63e6db37c3ad976010553290361198b3b8e2b2e8c8148416d57420159a5fbe
zeb16cadeae2a941a44f49d44121b44ea93a5e2f08cd9c07f5f39db3b3cb34cf77d50d6adb8ae8f
z0440e72465ff56df1ade4b206903b2c05c01c6e969f0ca46bedbf4c26b4a6397d41943c455e0d2
zc0835185167a8b6237b7d8cbf0f71d4d210c1369782c87a9abee5f779f5efbccfbc0eb377a75b1
zadf8091cb41f9a52cd44d1c69b985443fa647e09a8be82edfe29395c2ee117974a4e02140e3aae
z0bc26c974807a231c5accfa4e9276121710b0d51a7367d08c87bbea8a476eb273e6e870f5850ac
z4f860398b652b0e237660e61a024967e4d6a0c35009413345ba0e6f2970af0920a1a095fc88768
z1a9a296af40c6ef48f55fea682fa742f0f73c17bad4af8ee2fc2156f5afa3ac7a1eb03ce1e252e
z657b9291c0c028b30e6b1b6c989aa96cc3b34829435af2189633b867660156436eb0f61f0017f6
zbb6f47abea474e15ac811751569993ebfcb3d15e16a12ab745538bda34411c495e2fb9e34576a6
z027b416f550bd44e024f6994b15fead0c1a4f85c44f20959cbf38ef2b4f1b9a705fcdcae4f3678
zc123ddfc89a037d5b66726b8bcfd7da3ba530c901519d435cadb9f63a518864b31036c7cb72a12
ze43c03efad79fbbbb4e8cf08326dc6b51cb99232e7c2714b281adef17ecf9249e4506d6ea3581d
z595a9a169c597d9edbc22aa6a0e00602b3f2b004db98bcbb9831890e2a38df9a2990895e995b70
z2556813028393947cf559d060bac8a1f64ecae3964437ad36ff6369954b072f3e2f0a2b6bab350
zeeb3147c70f60f0d18df3f9ccc949a5f3e5a282d0bc5529316e8e2ab5195ff0f7bc5ff485baf73
za52d541154998e1c15d9600f1eb911d2b2c4b9ec0e7b5b71e66fce570aeb95be1e0de69756cb22
z2a9a418856ff2241c897aa4212da8dcbdb31c852b429bff3d50b4d7e37449b79de677fe642860e
zcf8d1e9558e598cad0e1b0de0a255fd25b04d0a0fda60da4ec6b2bee4f764372b6e9ab84198820
za6a4e9c4ea7db02ced4c186f032ee958394c8daa596e719e4fa9a80c976ec2f5cc88dfc0be7dbb
zdf8b45e5f3dd9d483f734d54856c1c89572f68ee2d56d7b77bd1abc56b40f31037481d3cc5ec89
zee042603a44583cee4396c6e7a3dd1765a9fea994c8717f1b3487fbebcc24b6a6aa6d924a2688b
z8dc5299a2de98020a517152141081257c463262f1900c55aa1e025b576e5c05ccb34c5eb2ee0cd
zdc893aa565ef247b4efa75c754ca8f6b15d99dea9f41003c2650edfbc0adebd21075bccf89ddaa
zdd2b0fe699caa7bbb59d07ffbdac9912246df949f420ace34fa7067431251f85fea638e573d8e5
z3b4a074538f3a91c1057aac554aa3a4a8c52921ec1a28f4648cf00b3916324965b12fdf45d8dbf
zac0a4e26088d7c7aec0b38f7996881f0af1a06efa6658222b5e638bc8a11923c8b36be34f747fb
z0858189ac8267fefaaa88958596421aa5585a6570d639cc3b599926b5d2041c4cee2d7cf71cdce
z43d36c6849f99b2db6c142a2b1f7c8c4c10691efc78d71213f2a54235f78a10f059e33638ffca2
zb5a12743960082e50a05e6c3186e9c49fa17439ecf97ebbc977660fa41ab58bd5c4fe6d29268d5
z0e80ae2d0623c5ce9c8d97b6a26a14cee5ea25fbb4cdd8e1262bdb5fc19920f3b5ec5a4050e5e7
z3e84198fa8039847232fada3c5c5efcc5236b33e7a730f95a5e2a3c8252df63bbba0d9f1445eb8
z0655dce4cbccbff2ad97c18ec160382ee781923ed32349ba590706727414cd250d52819a0376cb
z5d8103c5b8471eca2b0d5f229ed6abc84781ed718873376f2f4a2cfab7b18b7664d1347134ba2b
z079a7a437fcac8af984fe22859204a8c996231b42b04347011cd2f8d512223ba2c6412447845e8
z3e45426d63a874703d6eea8285904bb7c28ea275acde83d0dc86d225dbfc757addfc9f6936798f
zf1d63e4008e6ee059e6a89bc88aadec3ce3a1c7267e10a6022712bccad446fbd9d9667c936655f
zd48a2b5a496fb010cb6e97eedd50c2cf4f7863cc6eb5b1fd87a1bf369d274e1ccb6fcf881e4c0b
z98f588ad2214de883b5ef7392c32858f167a5f089824920116fb684d6e1c794026b40b7bba5450
z6eb0a28c7313e8fd8aabd5f751d32f7b959d63b70e2fab1baf8a6aab5c9f806118cdf1cb7e14ed
z80b372c200b433e1f13bf7a925b6bdf8f7abf9a5229b0d85376596526cd724f5d015a84b1b14d3
zcca560baaf4fe70a6240e39c1990fcc8a0e0949ded9cee364bee15cfa55c9b7b54092016fd6382
z8910e78b5cbb6192a6cfa9f0f5605b1aa4d0c4475da445967fa2bdecd1c5572a64f76e991999c5
zd6e168ccdbec34fc0ae7973a8b8d43f7f23b5eb47b71aa91184cd587b5fc14b4bd2adfe169f942
zd32accca79b93b5b66c7b41f7d73a2686666faecf1116b4f8cccecd5d6ea464c9be75f4bfb3a6b
ze9bb8e96c06a0c7502dbd01489c23370b197f7aa024fc2d8fa747f395a803acca5a579949208f6
z4d89383f8be3506d4f4dbe8be4519e1ae8b9ba99a3acb90e8d80d3d5099fbc74633eebad8afbef
zd49ffa78cc0422199462dcdc1db5fb0d092067faca48f03c4dd4fce003b1f2e1e202af04a6c854
zfeac3c2f835b6bd204b23d622fafb2707b59bdda80b0692a00d1f93d8852be8ceb058608d80f29
zdd2c779c65d876e663fd1af1ff24ff7551bcbdb15de10333537bd30825e419a8bc27ff3f9afe9b
z7f8cb7f78bb024ab2d6487b75b4b842d523a0e7e7099a95af59b5f945fc87d4aa3428649b710c1
zd97c002b390482089285afed54cc1fa7a0c4aa78dca37fe5981af60d2280d1aceaacdafb6cb536
z87dd32ccfee323805fba9914f82d157eea89e1c7c268e9861f757bf1e4b39d00d83554fb611526
z094fbac5a5f1deee8c94f7b1890e84c18f1168b09d4f216b88ee8d1e32ad893c3c0098686844d7
zdac35f89e369e0f77cfa4c4d4f4d08ac093093c4063fdca9d1e3235f250c322f3fb0ad0366dada
zcd097a2d9e01dc4e20a1a3924bbb015c348d9f8d525699dea51012c54ede2f76c95e9cd2172d14
zc44ec6679f4f82679df02ff606aea4b1cbc7e171d952a9548c3e787952083faeba11063027f0a4
z85324ce8b42625917fc762f9b17c627dbeec955e06e6e1ad4255627558780480f24d94ec49b263
zceb94304fd8920286757075ce23116b63db320927200307dc9a2f985dcdc377efe153309a4db10
z1b4c7a176daef3e3272e83af3404f839a79dbb8c55b873d1a9d9e0d5c7637b658fc5999d2b01a9
zf6f274fb949e44246be9c48d8e9f6e2011470b8de4b1316ad64161125b281d676614702fda4eb6
z8175a5a6c0e2c4cc74070934fbd07f41db2b44192d7ce14c698fb4f18fca4e7ae93590eb85b09f
zbccb211059f62fbc57b28837e5d061783cef5a22622d4168bc04345fd3f1fb4311cb4d3904837c
zee1e1a03d8e761ac69b2b5ef0e79bf99f9f2d5f09c142fe6ec336e3a4f655d4c9a3657907bcf1e
z7a03db6c06430cca374c982a84b7ce02c12935c23ccff716559a66cef4bcc6c6118e3abcd15d90
z19b5717fd13af091339ecf6f2e49d0eb1830a50bbcfbf2d31857401b193949f95dbb78bb963c57
z7cffed94e716ec558b396a1eb8d062f333b4b6a0b11e523c932c4e3d0e1888c0a60dec010e0655
zaeb1ad0d5b19df95c176e3738b74314e665a4e551944ae0904c6a4e6e34f3912c074545e379098
z925a507f5aeafb8413aa68f30fae6dcba03c07e3f7687a6c3079db759ca56b5fbfa07358f43f3a
zbb56a10ba6d7b6c90def0997b04266625b0bb8bb0c396ecbd273eea765e632fba9eb76082ae15e
z6719bb167b98da6a55d8e92711da97bf0b6837465f12f21dd3aef75b6ad2900d6069970460b724
zf228125c07e5a97a5cef58e8755e0c8e278df9c68b509edd2db5a20e3885674a7165aaa1ecf246
z2119bca360dacd11e5995a95453c2af11e2be20e3f3610e55fe5b3fe1c0bfaa7c886d9feee9f44
z7ab46bd52618311b88e7249138bfdc34ddfabad53bf00c60c23aa6fdc78ef83b170bcdd0459fbf
zf5ed6bad8a00a840e65a5e49241e9399097b639440f79d6b211181a344093c146b298641860ac3
z6c0ebcccd72f01bb25e1a7838cb2ea7981a72dfbcab33b351646b69453869511e71d04f27b32b6
zf9e10bb223ef0b337744b8ed676d958a220760f7b77f55fe65911209a8d4b23d012fe3b3123bb9
z03e424d69db8ff292e57a7fecf52488e4b07bb659acb990619dee90e0e89906d14453cd33559ba
za26f6b7020981e838e7386fa01d93cdb64a0d99068b1e7f3010ed85ebd259b9e1784ae4816f9b9
zab733804e8455568b876342e4470e6c61df61e59f45a4e5d99179b083cfe5357100dbe8a4d1e36
zc9ec8f3bcc301d7dbaf0021e35199d8c9d726bcf1a267c2f8caad6ea433633faa1866d601469db
zdac139feddf07b608da17500daf7b1a3fb07f243493def8efeeeb58b7b3c8c42dce40d9cf04e31
z59c1d28cb330954737a7dacfbb1a2d8dadb3791def7258f0ed4b1660b1cb088ae39d182a5ed53e
zcfef76cf4b79d3d7b695b1f5d7dd80f76294b3939dda45f39c4198931272a0699d20f8518239ad
z182f572490bc025e91a38230845f6f46e62204c682b12d1dbd4a5a2df26566058a1ef02d5fd4e8
z73e2cf2a4b6a598b6579de53e1371b7f81a633f5f75a27d3e496f2c1f5b26919a1e5ccee99fa90
z97077e523ff36eaf1b7c2cd2f4e730a9ae150a0acea1a707edbf7c0b6073c7c59dfeef6afb19b7
zfda95c2686010c20a02a9041b0b0725f8816457689bc9d14d775677b1abfa0f98c14c1d7fc147f
z91336f53d2905b3a461f090b991be198c24ea033ad4b3d453270103e554856dc75236259d1e688
z1827fa143fe9d8733a0487d8903da2691060a70d2241c5677273e754d45498d8969c14ab2a051a
z34b0e95c468b2b87c37906df7ff4280b0fc411a67d495adf32237b66e3f5a603599dd152dae76a
z6d00d34a4641da7e144921d9ff8d76b0a9151cf28679dff894998f46ac1d014f1cef9dc3f1c030
z8ff74ca91ffb2e1a6f941cabbfdc37d90c8896036e18cc576ce6d66563ae306a822ec8027e9f59
zf08044d88feba30935748ee6024fb39449fcbf43daf453f4d56f77bb3e9ef32919117db28a9c0a
zb410524be4180a485ccdc9fe37384c8d7fdef4553a38afd037811a1ca52cbfffe95eff1c2aff12
z79e19634f25da88f439c61053f0812071fbb571331f90797545e560aaf13daa77b2176763a61b3
zc8a002777140b2860913b789e0a4ae156913571f8755a53fdb2eb64b82f2946034f92608642ad1
ze4488c017654ce546242789cda7f581d0299848d3726a2c822f39d384b3fd94ef3d51d2626b715
zd6e2f9d4520d39203528610fb7b435d1aad2e4ea4f7c8ad157ab378a093f27c1a859f62a978489
z94ba2a692e47554301f9ea8f9bd1e79ceb1630cf96ca93e3085cad602140ab6d9f19c44220c579
z21135e3ff8b9e4a42aad493ad3a045caf8c4b89cbea52d8979925a55407b2c788acc2e96e3dab0
zb62d6fcc195de1d9307fdf8ae84d2085450313439d464a366e1eabecd9eb86e72cdb9d8f54dd6e
z17a0b453944f3ed5bebe48421a035dd46a9cbd96d43593ff692cecd4dd809f4fdd23d94410d61e
zd24e0b5bfbfc6bb58b2828c8be71ec3673e7ad46e676cde1a4c9b909c3800702d851306b9074fe
z76fc130bc7fd57b692042365df218c889eb2ca18d929aa898a90ff1aa9f14d3bd9b66164e68ef0
z1bf75705a8e9272689e2f4c7e3620eb05cc0ef102120abdc9a7d0031a733260982147c41094a39
z7d53f4b8b40cb3c537dd8d48d4b881cf277534e782300b1537f7552154d61dad6f618942a656b1
za4107707cb5d666b775b192a064df7b02cafaa08998277a27660a4bab7176e5cc3d4b771b3d3cc
zc115fb091c07240197486238b6fd2c9567c3e7d15fd2aeadd9a373e2724aeb01f048fce4067ee7
z4e2260e1db995c664e2a27aa03a58c44e938a0e3033722810110b0223a161634c32793944c57de
z5b09d94b1673d2089a2a928bbccbe5837ed4ad15bf89e46e00b9e6c51de72d604de10641e61a5c
z67f7d45d713b3c6b54eb083f91c6742cee76b74797b098cc9dc2e5cbe0bda377c22a32ee641049
zf1e37332def9f5ca5be2e239dc2c183fbda6e8c514e539eb708563c940759043088d76a7bfe4c8
z1a5faea7c1407097ce733f8ae8e3d8eceae71c994eb06f57941ac6d09489ac9e10d2a503ac7eee
za248b2e3382bcab2ab7eca2cb9275cae48b62d4a4fdb15b194d7f72dba28fd5cda83b2bd0b75d1
zc89ad1fb967ba77a8972ea3f55f1442514dcb372170e50f7de3406108576ac6ba2641a7d4a163b
zcd5c6cd15a2fc23df8a15b1d07b889757f54a25583ab24cec6e39477eb2e7147242f73e820a49a
ze758e279bcab04b60ba4b15526a1b59cd0f9bed53dc01ede44105c7056112e9db06e1b0ae3bce5
z1fd7a155e73f727db5745acc6fca2cf3d9d99f452e6f279433c4b6495918045af204fc27cd5459
z26f2abf23f4df0550b8ea77cf50e6ce94e584ad0601746ef5a2a2d61d172a5f869d9d260f44fae
z4ff776750c5c3859d07d8124e69cb702efab9cf1419dc53bdfdbe1e618dfeee14a79cd4f93035c
z844288c73cfac056461aaa316ec4d456fe4cc3f17ecc18f1eb1e6d8409e99236e4b7f40e5581c7
z36a1a27c6b5c75fb59bc6a727928a4ebb531ec1e3e16f35a36d63046bbac174c8b5710f6b49ceb
zc4abf2638e91cb19aea21cb87b49b3d2b14fd83443cfa86f0430a448832f536e3000cc000fed0b
z3f79067ceeb8529cf86bce17dec05b10c244717f22a7872514e641de27a7403b4ca1d8a84222d9
zb2dc9bf9faafa560ccd6e004ede57aaafcf32ec16d3db42a46941620ff38f15b9b84369433da8c
z4bb1107b775d79d64ef48a3f0b47e81ad0183210c5d11a1a9700f48bd0b45a15d0bafb42830169
z43fc6583a331102f2d79fe60155eb7ff539964b363b1d635eb618337d4d5dab4c284806b612c3c
zfaaafbdd5b46dda795a649c2354d4db1fdc5f52bdc5ba5b243f21f1e248f6f08deea1293153a74
zbff6d44a258a4835b8728e035f1a5d88a77f263decb9a41e8ad2db39ddf83d430cd609af3250a4
z691402d290e69b08066a07af29a590867180562e335fd7a3e978fe0b285da8238a0aa69f1b20a1
zaa38c98bae3e76fd3ed973f9848a0b272bb076c8f113580825a48e3f9442d1613e2cd2ec952861
z9b6c09a841c32d815a8aaf31bb26d1095fb701811c75b19529580487c986888a44e5b8e03e6c65
z7749dc4766986ebe15afa48223b65c220178fb940dacb73ff1c35fca056f80dde13eb731be9c5f
zb98216cdfc675b3cfac5675e77fd7d2b03483788005a39bf83feced0587b6d5f49cdc52239a2c4
z8272628bc6f8db713071ce1d44e9247a9cc441e56228bcde5b29d2895d3059e6f57db646b8d2c6
zd58ef998fdc83a7e2f3e204dc9177a9dbbb16511f07228440928bc7ea5b12efa7b33dc42878f57
z1ed57bedb0bd12f31981455410eb59049ed71e7c35ce66a5489786daf6f5b1ec0af5c47087748a
z08dfcf1d2fe7abb766a6be3c642bd3f540c28c8b0ff70f339d32271ec232ea495139af686a5399
zea73a2cc69ad25d37581e0f92069cc280f8954e5851abfe0bb82701f747131c596bc35b2da56c0
zc11c1dee4c14df820dd41a097a41390b621f901e5f02025ed9cef70d2f024b74f08db199c07abe
z3996e0f6bb3553d5225a344c6526cd6a2e8ea1c743df05b7e20b1e736dd4eb5bc96a23410d7349
zadec44d3d1dce65e4582177e8fc89c03e85d73d49a22c4fba918277f8d5ee355f3b310af8caa3c
zed9da062b75e81a48b605a32e81a0aafccdf2bc0aa506d6f04a3e3c7d545f069d95329a3546ef5
z7b2fca6ed97c2269d76be45ecbb23227490a9453ba120e6f7dae17ed5e0f841841eb585183d6f2
z6e88936d6f6e4e7e67df9d7012da9e6ef96b183971ec8a49d47a8316330cb01cd62376e28852de
z79bd714d50afec49f91813047253d6bd398258f9e12add236acae4caf09d05ec7dc4d8c9d441ab
z12ca2631cfc9f1b1f4c20f28a993d214c3eb1ec73676dcd35206e4950aa830feb52716c467f53b
z988cfc7fdd46ff3f2a272586856ad47deb633dfe19cbd1a3282976ec105725a9f141bc714aaf10
zc6bc4c5546b7adb37781d4dbf71bb0ac784342405e6233a848ed46792be81c19c4d6d24498c06c
z750159f2d809fa22b03b2098a22d7eb76c9039b12b52f5127ff9834f3186fa3f4a3d95133d2c6f
z8c52a5ad5ee16e6bebb227b1d473d666b9fca0ad6706a697151300398316a3447da4a091f05058
ze0ac51cea4b1848dae61fd55a4c3aaedc83afc499f992d051c932f84751155d3a978a23446038e
z9b3c09b16fb4ea35d4c874d3a975369f419c5a74fdb3f741f94d12240ed91ebb8d99824adb6b0c
z7db3c9539bc66388d5957f4b4acbb32cc400178f9b3c43e574bf421e67467a330f544c4d3d6b67
z063665187540b642c97b2436d16d114f3769190ad5f4e51f8c01c8d8fbdf3d38295efa26ff6c61
z8b62aa2c78aa7ae482ab0a7042faa9dc12a499200e09fa8e1b8d38f7746a6645459978e3aec610
z5146ac4ddce7a575f768e9b609b4d1e8df00736bfe1189e98cfd3b693e4b78d26d72b741b38d78
zc9abeebdfc78c12f123aacf13ead428a272547e304f9d5d979277bf505b9e7ec54a4327e579697
zfde1661bec131b8759ca5c643550728c3aa72c757bf27d53fb272bb09d8b1f60664f83d7959f81
z98efc377ffc4137a1f028fd024e7d2828f793ef4249ed919593737d2ec6d4f03e4e75c823a73b8
z04e1b712b0a30c5dc0da55e5cb455909b94926c9c3e66bb8a89129eb0ab8bf71491ef4f03e7fd4
z8dc7509effddfa3ebea8892b06ed0682ce4597cc20b71cd65edd987bae9d3be1cc15eb3e4dcf0e
z573c3c23edf93eedd91f66fc8eccb14550763768da305b33d1960fc77edeb73f33903ddc015ada
z915b6ee11fa98d092511f501bc3b01494aece4ff5bb17090ccdfe871114846f05a986bea8ae570
zc5c0ab0842df8216f31913e363568364070307533703d416d3236c7dfb3ce58d14ea45546a4836
zef7f317b7e2e5351918f925cc8dc874a9327f46eb8e04d031a24db6387e266515a978885e0bc10
z52b361813d2e769c0287664ee1ddcd67b09b6af003a3b94d2e48b147a906ae8460beaee09d28ec
za0a585cb2faad4085dde6ab575c9b5039109b28e020626a1360cd065d405f22e46b04d459e5070
zceef7f0e0cce98105d9b2c87fee1c5dd46c2c1b9d41f3d70c61574da0cddafc355015e760b542b
z365889a50e0f723a30631c1f990867e56cd599c9f651b6d6ca99b8d12c0316507a76c272f2df6b
z63b8185a4c9aa05081d590faf5ee9f36589a1ede9b03a8a273682c583affbec550179f6eab4aa5
z668c54d7b44ca1346e3c27b048e05201081d712ae030f515f11b5574bb41543806c674110d719e
z8c920b324f7f638effd5b6acb72856dcdc5536bbfefc68616fb6a23a917cd5390bee05f231ea13
ze80c213ab438c549751a281ffe23165e2f1cb55a3dfa988bb626ca9a907b209a7fa43efa51c80a
z18f2fc89cf73b7ee382394d8bc9b1e36434707a2ab7629e2dc4a3a3ffd5336f9a08c5cc29b61f1
ze62c2af1081ed6684e375f9fb0c687f5a1e288688476c14509bd0efb764d819d172cff138eddb4
z402c1f8c617af626255efaae2c35867adeeda0330fe67b2a715946349649e76705a0e04393c61a
zcd1915608f5a2480c923e31166b25f50c2b1f6c74b0f53694cc782bb615c53eba80c8e7c0223b4
z1432a51d9037b8b805e6904d60ee498765a0450efb6d2d1c70915bd4eeea36833bd112ea706c5b
z479de89ab27ca6e431d8c460b23a9adb7a4a95144943d399124b0156f2f132cf24cc6c7ef0bbdd
z85e1ccf35dd1c5ec6c483d2d67a10f4bb2e5a495b82080137e267c0f01af952dac04f3345bffa0
zee093c70866be1cdd40b72efb766288cbc3ffef76ee95207970d6752aec35612786dd5558c485e
z838d453d8f766bd67eb37405f1ec9ddd189d9b878f53180efa63759f7e665a868aac5ae86db0c0
z6fea63b8539f99ddcdf2ac188b43cae6591f17844f106dfbcd21cbd49edf43de9efc51c34d8144
z0113593db3f29a49314b6ff715d11b570d264f6a75d43df1652fd52b2aab2890d85cdc56afab28
zc3d61a146ba86b4b1285b638d3d72df1d69f50533940c7ac7ed6b363eda7e30cc5abe5bb451fa6
zd0a3e51dfc3a784ba421106208dbb3b6eae0d8ee1e798e0302b90dac9b94cc6cdb66a5569fe1b8
z14fd8bd12a90215b9d1ddea170b482ac3a7e6d349aacd1dc8500c1fc6af2df25175768ed1d79f2
z6c72c5b2bcf2c8c517b304af7415870dc99f0d5598a0a38cf48076c0a4eacce6a51c0a438769e6
zbff2bd79bb5b92855b7548f97cdbe503c930021e7e17eae1e2ff049833ab818ead576ee128b655
ze0fb99912da1e69fba92b58bfdab18da00a82f236b5dc8dbfcbb657f0e9ea5ba29f4dc98b574be
z7221a1b4c7fa190d20feed8be4ca2ef166c129f59bb4f0ad70ca32c20ea08ae9a423a5366fc8ea
zb4775f4e12c4c720acf957045544eabf5d7645319e64c68d8c05d6e95f13ea49649537b3339cc5
zd3b9d1da65f87bd06da26f05a613081045ef2956656b65d92374a510d33fefbe0fe4c1df8fa7d9
zcbaa935cc9c651fc3787ad343c8d23e179d4695af749b483616515ffa6079f239467db5b2c8a2b
ze0e354d4b8094fafdbe098d630257caca45b11984f0985960652c869f91076a52197bd62420899
zbc84f74cbdfca89999c731581d23fd17e298b196aff984c0096af24f4d5fb8cc9422b172d8b698
zda7a8800f42fb6bf49dd68951d463b93409c958170770b41c832ded4cd941966d0894da7e1c2d8
zc9371fca24c4faef2b6218cdf2f2de2118db3066ef5638d3ec8e941714391ee60670a378033666
z42a0c831c2d4ddf315d53b0c0bc232d53aa45c033f2d942d5cada8651cea5af25b3f3b4f009713
z5a5f8273b390aec258f6c42338b42839e46927387e5aeb1163fabeeb1ab7a52565148e3cedd2f8
zafcac6af5aa347c736e92117b4370c4b7b0daf1f7a23c7d2f1a77a725fbb5b4fb6c83848a86a6c
z737063ef01574daf6cc65850a8fb9e188b32ead2032418194d151b068fb9947f91e9dfcaca999a
z4b0cd9518f57803e60b6deb6449c38d4403a60e6f63b091491cebd956dbe8849a993029ca6728b
z2c1cad29c74f326ab078968524352d4035006644aa446a28941a99571c53cb1489edb92fd4633b
z4176bc82793dc40fcbf66b0a7b6c6c5bb3c4de253752870e247422edc733f17d4af1d4113bc287
z0f5df6538e43ba925c512b53b78e337e06457226284c18529fd146d6735258218602d979f754eb
za3847f875a87b12a9c1c939d8ac0230cbfe0798fc896f8dbecdcbb276647e8f2f90092182c94e1
z9b9c0ecdceb6d0529989f3c178dbc14ef78dd6190b408d6764331bdfe4fbc48c5f5e3344d2f0bc
zee7a85f376090716198bec6504f9091c3209569863926e68dfdf1b7064f0b08cdf7cce92e99315
z7b39ad13c2f6f0e2166a496259d9e38c600bb6601874a4ab918cf082f06408300a3822cbd13396
z0b6558e723e3e807707f8dfa865a88a17d5926f1dcdde4afe279f565597d6c94d875a42a3ee017
z5eab164103813d21b540fa3ff8d1a9811026a21c83e4912cabb6d3085964c954ac76151ea54ed3
zc53358b17b2619bb6f546a6cd9bd6e56a533440d99de2b882a8b8c620429fc6816f81e7bad5011
z96dbd69c9c5c65c0fe56b0a3c72097a2620418134d78bd2975847397de7f841d922936af576c55
z53c0c299044a6c1d90486b880ddf0027ed48e52e0873a3cfdee0c2f69282e6fd5be7337e066066
z6d86543e62ecee3e7124e488e13918538dc43956bb69b2eab404f70bfe810ec33c565d5c87da94
zf5647de020a698f0a91e94d4153e4cb7757a060cd5bea6e8404a0f3b1cdaf5a593b0558924dba5
z3ed5e76315702bbe28cd37491b09506d13c5f4620b169ed51499c0f40f878d167319ea0d4622cf
ze31f2364e27cfd1486da9d2257296badf46305a38216b09468df1d365554970594fb503978472b
ze798a5ed637046899821d33006349c7f72a5a39759428a0dde899bd56e65b85c3c1d350cb9c29e
zc0808816a3e9c3049b99adbf986417bab132f79fb90624ba0942cf9475d95a1bc3f4638d35aea4
zf84ac8aa6abcfb658bd14d41a637a0cc2e43c734582046e46655b0dcea09887a0ea63f21445f15
ze1a399c318ff96d544ff2dbf6bace0006c19cfdcb5a7358d7b80abf5b63da8ae36cdaa2a4f0fc7
z9b92ff8062bb44d441b93016c7cd660b94da3f22581e3121a1f59acb47a3fcc1a77077c5175f96
z2eeee65c1b987e9e346399449ecf4327de595a9e0de3f7a0ee1e8c3cc91fd9b4692b01afe76c7a
z05575f36f5eddb03790bdecc4b7af9beb5b2835e320bcf613f155b07b34b133cd369ba565f4a80
zc46747ad6ef66e4806e6a979095edb306b56e99096ceb6a29f68cf4aeeefc2122603c0b5b9f3fa
z21be1e02345cb84ddba3745fa9a0afeb19ada712820fbd408286d5d113fbf622b946c89c7c0d14
zb0c46e73d5258701375ca7ffa07a02a68c5812c0d4e078f54d551e10ecbefd5dd42c551f561fc9
za440da094d40e0e156c66a42586336d490ce01cfd09c7cbd122c25f53e9dd82fd7c562ba420393
z972cd841fec9f6e0f0d1f13825a21ae38b560a4e5bd3d034a8323c7366a2dc53774bf40912e562
z5ca82c3dd3e1273b9b2ec6257f5db34171b06d930682a58f35388d49439ad389cad95a2b65c2e7
zbf51058e18a335a51b9ebf654c6642b5b73b6767d894f5511358564cb15394387e3693bbcee799
zc5ef1496b5ff5bfeb4c16a58ae129aa7886bc029c4691220081feb27244a0ba6f317758586397f
z383e8b9a43f800f650d49c326bab8dc206f0bbde29723f17f5f7a5941c46eb5a1cade2f643327f
zd370df7f301620b513b0a9f29feb437759f65c5cdc2520c861c3e8ea7ff598533e92acca5bcf37
zeddd32b2ac7e825493a963270ceff84b01eca8c16b011b0498ed9069901074292a87c3c96cdcf6
z0e33b0074e7e422e2430c42432ce7908c36b9348f11b7fb4d8ed4cc2c2ba764a1b5a44b42f47ac
zb9f784583473928affb46a810238b262a2677df79791776f519b66b457ed44ad9a7e1063035f1e
zd82b38e8220c642801608f82bc10205e08f7649728b2471f71d333dd65059a54c128e5ce000242
zfcbbc27f1e43eebfc863f187b9cb2d95f33900f6723f855abe7996697af9ba60773015f2ff37cb
z670a1b23aab329b94f02b47ee2a3871e6d210a2f0839005cafb6937a48c3f1fd005d6ea284be42
z6cdca12bfa37423c128e76ab82bb455bfbc3737add0d8d15d15c8f26a315e43bd12e0a00d52e4e
z379498a824ca28c852b37d235e8dae16315b5c1c38ed07213ffed5596e920e12a636c73f381f16
zbfc1444ba5a82eff37ba7d644f7a4f636827088ddf6e0ecdda77facb8e12c1dd3fa723b6212c0d
z809541b80c43cfe7e01d112211d6120cf45ad7c285289dc5e238f3fda07619a3ea4018f6fad4a8
z81a7923ec7367066e6a192c88ad65378f38842a0d3971d7dfc44c99f14c55b3e8eb3ce52f490c1
zdc2a920c0d2d96d3c95054a43f1052f033daa3f067dc1183f9598675de2b089beda9cb4ab28514
zfc477738746b90e6db5fa311cc72cd8a23c15d1fbc195eb001812b2554ce4df450cc591fb3be50
z109763e627f6a2ea1c48471b9e5e7f20af8b547ec4d7c42681ced024ab3448e4e717020deca3df
z0d2b0610512de67ac697e062fdd35369acb682fdb2e85ddf01dc17de3217eb487830d7b66861e1
z4a040e169f948a8f51fa701c86f6a225ce939a52c44a75412defb0b693d6e69a3bca1a793e7773
z02bd49852be8d91d383e460f044fd87fead7b0c8a6c7cea2df97b52e091806609b89d6c20f3c25
z1180891c19623783d4fbf037d8f2a1f2ec86270cb460e62cfd255ddb33761f218d367c83ff00dc
zb6b3b2cd0dba4795e50343e4eee5ad22d2271018997a192adfdc8a1add3817fa7a5c73378270af
zae4854829f5aedc5cdd51d1be1be1e4ec737a847fe9ec7184747524d844cabe9a7e68428f04ae1
z4db19db60a598ba95075eea0c71257932d90c2eecece9e523e3b6ac1d0be369f07e2332db754ec
z6e1f0d2a2574115b966d0ce27d53b70ab28bf237fe38aaa0d7b285c7d241edfbca2908d6c2a0de
z390c6a87f7de576470d2cd973c8c6dd015c06b741cdd7c38085105274eec137a18b11f79c31004
z5b476390cbe3ed0c2a016e7b81b6ab49d9707dbcd57a710fb1bf775b0c4b9d096b3d30eb53f8a4
zf79e6014aeb3256ea6da98791babeff92d82c28c9dc1d36add179dcd19a628d39f656aafc8a02f
z451a588d2e03f22ac0f81ec255df7d32c4a2f56a00e7e8663a663b6fd2c735b502839fef473f75
z7eed918b40292b6d8bb24f3c0e47270e36045ad30beabb8f0c340c4e5ce7883569e80e5525afc3
z5afc9b1f15f12013ef93b76ee4cd2f58a71e1e639b2cbc99839d6ec711b8d2f421e67fc77097b1
za41154e7b6c7774214f9d229170f51677d2b53d7e63385505e87d0753b6bac3d07ec8d31d86b88
z3d1ee74431b649df499604c4dbc6e6d54987b14fbbd22d99726917c822e5c78e2e6eb01ef58797
z860f2f15de079e64162963bd0cb16bf4f821e00332d4f19cc79766e8118c05c67fb9550c9dc8ed
z55664d267ca129f91b0bb770f77f3afd3327901d6cce9ca1817217f352621105dc3bad06326fa3
z0662ed7874c9153715b311089bd8575d6ed5082a8cf011b251062fbd243aad32c5731fdaa411cc
z7dc75c0d4fe940830bd3ca9234f8f6d3bba89126c9abe55937e967434b6a0292702ecabd52fd99
z70ed24c462e3b277ce6969c4abb5fb7283bd73152ad0b2a4f2a274e343f89b4c7919d3de31574e
z8185fb0fd38e4e6bbb6e2afb5712c85ad7d6bfd0e7c97bdc3b36a244fa6b4b95523bfa2b67b7cc
z73c65dc0a1979a89dc8f5a235a63812d8ac51ce377968b3244a3fe6bb59e606ef2f741f52629e6
ze49f9e5f28aea49453fa5b4f67db4f5c5c6ddc3d82300fef434c16134bf3d9b32c8e85a59a9c7c
zff28be8788713103107f5d0e4ab16d2fe600ae9e375c5cc8628c5d3430ed1d756846929e73a5bb
zf1df34c76530d195a1923050eb4c85b5e62f4bd1a0ed28e8c79492ed510f1993b946c47fec567b
za932dbd18867849e7c4e5dd265be8edf2ed87f48bc7c56400145ba1edb469cc2db2faedd21fba5
z1039d23f1862f279ed3f89e2de00e6af49d349ebaf7f37d8a12902dbbfe451a4642437c07319e7
zf9ec609e17d253aecbf090e63dc4923223035f131be6603ece997122dcecd158793140f14aaf67
z817a8de1fb274c0f1d7e433d1478d4c5d5000141d6315e749dbe9fb18cf57417091a1456e78f76
zd33627945675cc0a3076fc933c3b92271a23a695df797b18ee9752cc58d29f7af7fbf208204490
zecb35cb02dd6f821c2cd7f64617645fa5888f92a26a6d8a956d31a16981cf6638f03b29f9648f7
za9d7394eedf7faffe880efa0df19103ad5630babe513f7874e53e0c142d5fddad9c82e2d902f9b
zf735c3f19dd5405922837450bfc6f250e5291a21cae8a183b4bfbd2363f111af382be2c5281bc7
z2f48389b93611f9b7d39d870ad1e2dae0e66644586b9849fd90405f58cb540f07496ccbb9d72af
z4903c5fc7e4b2528de19e8d96b851421d309f2063d452ebf1a379ed57dd5bc5fd685ec5b7a2cb9
zdb747d6debb0d70d7eb03fa3d11e435aac9aa6a680bbfc2646928c869d29af0a0e5936229087ed
zc97422ab247f1d3e3e9dd5cc18713762d1a0052e2b1d0ab486da5851e0e904e04441dcf7c9bf11
z582d69e25e7b0501532a89c2af69fefd1f79c988e47978966699dd624e6b5ca4d6f26bc4752210
z77b6adf8e82de382d9f2c96282f82b0835d3a621b618c5502cacc124a5e2092d1092d8af35fac4
z955092004e0c32b660aca43135aa93449c255e7f6c9fd9509bfff61a0e9baa55890cff41d02ceb
z0fe974224c4e47d2a9f4d5b7f0b7c8e4d7e88d18c529ff88656e6ae23cfcd13676d79c67d6c2d7
z27afcc8c4d156802fdfc2dfd42c464f5b69b25122348c263f1edd343c1ada2b3edbd6345fed7f8
z684b0644ba16c52d4b4cf904056421512033e8972eb6d1192c283571ab0069f67c5fe6b96bba98
z2f540c36c6e1a52e8013da89011089d4cadba4e442977669055faa2bd8e16ec65f19490601b1a3
z1003e2e2d0ed041934a4dbfa6b7059eee916614ca805c98555568cabd4f078984a64fd2597c4ad
z70cc8df0a32fb55efb1d04988cd4903bee42385dc8062ac4a9512ab58c303ab60e8deb98f0aa14
zbca7ed91b730d0c4009fa949d0a33473aac1416ab802351ff76966e6d5e588cf4ef911e507f7cd
zaf133bb403492c7726e695e6369f1507a9fb2e0b58ee113cb8a5bc2ccad41e83ea44c4c6043bd8
zd1d51a2dee97bc9ef9d3fab77fd532dd08a1c20a00d9e5468ddb5f25cc86316f3b33352ad1c696
z1e68257d4c7a341906eca5beb59785b2c3962d9e3c7cd351f091ea2f1354ed89381b5c5e231c7d
z7670a0b4b2d193570a43e8c88be0a86123d844739e20847982540edcf9d08a143236d34b711469
z6fc2f96e6f31c5c1e3f382dc87d36b2774eaee1016a01343fe853265a59b5c6df44aa2448d3cc6
za626fe24b8539abd797a339b99934df3bd47d8e1a27214c6a7bd24e81a7717b2978b4c3ed41e9a
z5fc208ae6181f320ed945cabde8a0f823f5c71ffb3bbaafce55decd45f15a89e8c913c81988d18
z4f4adcac740b0a7a7762b1661fec8c36c55b89275c20458a728aba2d2a796e59fe1f01a2f3d1e8
zd73cb1b9cb26e3544219c2a21ef1cd9fd577002b784da0bfdf4b4d9fc84af0fe95290090e1a1a9
z24be28f774c81bb2cfdc115197f3b5208c7fbad7f278f67e50a46a8d92d4a496965a3ee10b9e01
z5a17b1a9f5807d1ca77c20c71fca018e40495dca435620951db53aa7c4c0e6e380724ec34e5b24
z8574ed5fb166470ca53610cddb399a308f71a7625088496cc1e8ce4f6474c39ca00c218940427e
zb1131bb0b69096ca1777cbaa2a5fefdd02aa0c6db8b97cca90b14a7ef7e68f545b62f2712d5fc0
z0def508c59edfc1bcc797028fcd5f9d44d9f8aa6c381ff3f9f9cb7cd863489659144fb4db6265b
z04f058020a539c71390d684c87a0e276a9c28c7e99bacff1ba24747a313d7d9ac77ac48cae7310
z324f7cf2f35a0832e0249e035ccbbe31254c9d10a5a518c18f0cbbd58e07c836ac3b8d212f122a
z54abf228865cb43c7c0d33bf48116e23672256c297533a0355c5e2d389370f39e259136a645b06
z77cd7899221aa0f3ad10aeff89f4d9774eceb42d8ab97f0625a9a681e2246e9bd4c51bffdc6b9d
z5ca48c864a4d825d4399fee243ebd6aa9d27b6d6752e653efd127d6e9575b8d1fb92bcac3b1b94
zd578a68e22650a4fd1f1ba53b102dd1cb2dfbcc1002e80b12ce1e4be1087a9cdac18e10b8d1b27
zd8049ebc9848255906ed643b7ef3d6ad1907002949e9e15af18693cfedc7f11f53532889038e06
z141f7e2acc9382f19f4e1bfdb05fea4f1be54bf121c304a4880b83b314262ba20eb64e6a1df5ce
z987358c0485e0e0a95757a923ac0e66660283773e461f5bf0d01f5afb8ba38fae8deebac42b15b
z487ea021a8eee009f6d23a1a6082db14aaa192b189c9ceca79ecfe9889dee16ec00585b986e9dd
zbf8ee9dc12d5728cbec641499994096fbf069b4df41eba38fdebf29b366c79a2854ca5cfaac345
zd6c3805528e9579c94531afa31daaae237d5db6ca61a7801c516bcdb6670a9f649b0e1cd1d7a6d
z8a68b6b857c89cb4f2d2e7bf6a60c3a286d4d76921d384672e828d3412aef5f9ae2ebee040e616
z48bb8f2f1446d36116e32c4b6abe8d83243c82a49b7913b86caadb9af89164736dbfb2fb82a1bb
z78330e0df0300b9681b64bec199b037c287e815fe5de2561007f44d76f52dd333e72ad7cb4195c
zdbfa55b874aeee6b5bf989e1b3c160367d045529f2d00aacfc6aaf80a862f5277ef3bdee16998f
zf79331f9b30543a172953ad4a9e3365ef02f4f78a64993d38fc7e3f95b3eca284c22b29e581694
zee8b75444a662d52f45005a5f3517d89d4d15107f4343edbe162d885242d49aaeddba133ce2a83
z74b106c5b4dd42a87561ec9fc1aa1e1937fc20d80b167ebc196e150840adf1f138c23c92be8dac
zefc9f095190636236b7a1caef1ee2f4bf710e0575bc8d30cb95416658b72d1190dea2cd3df4c2a
zbfb9fc365f747bde7a70aeb4b1973f8719a356b73da39890da28b534bbed33bc203da67ec69a18
z7e9d7b0cbc0cc669eff4349c47e8d51c0d9811d088d21c05db35cf0de82871fc5f683ac772dc9e
z83e21ec12669b0c1227f12e370907a39c048ca0bac13598f91dfeade36f211eb86efadb990d243
z9499a56113176ed0e25c3fa176be6c0872ce38d2e9a6e6b17449a9d47d178cc4472c9b1d78a2e9
zdcffc8b5453904ade41079a7e71cf29e08fe7e07ef7c8fff47989ce93eb9416c3e50ff8aa81564
zb4842951ea67b5bfc4f7c9a1a5d9eb4f3a02028dbd013006a45f680e179a6fcec3a029c7fdf5d8
za88790da29d7ba1ba5d40865d7d9d8c48d303c71a85be4900e57a58e28ba810c34d40acd27f4c8
z16e626b16633acfbcd432891160e5646ca6fdf2b6e02ff248a582b9def90703b710d699590c35e
z6ef38c78e5e80e21d06f58df17abacfa5848a52ea63dcf7de2e033a1dcc30e2c6c88fc634e32c3
zda1c564ec6b45ebbecf1fc8c2aaecebd27e5dbb2305f2c0935e9189da52977692e18757393f874
zfa1538eb013837923194220621d89e054fb7c11eb262d78d762585f37d5c2d2cc92277ccefcc78
z5179c3e834b03cc7efb178fd82c457cef219a6c8966a599bec855a4a98af22537bb4d2542cc88a
z3665ea99a29b4d55e86eddcc8da053f67664dadd99425f78319eaee1faabc61c3dfd530572507e
z5945fb7fa216232891808caa9b220633b37c40f14e97c57736cd89582a2b697de9dca4c6fc2d7d
z1826011458eae09e4ade66d9b47caf22ba7477c2264d4677c147dbf77d71edd8871d7b04bcd36a
z81847867adec4b24afae37bce56c51f0dd6890de934d94d1d6f345c826f3a2e5003a8af8eae39d
z2ee38ffe9e0dc042e68107e9b1f17e802d203431d5204e0eed9818794b31c2f58b44db57991666
z4562a31c9cba9a8fbf64c71c4b56a4442ee0fa1114cf24770a84c6fa1bac1c63eae94a0a98a845
z8e452bd744b7cbd0be5b6370463f3bdc7a5fda0ae12d5429eec71d1d837af19ed92468c4da36d5
zfc2078e7f278d83a6168a8c488da585f9d47da21e6d5fa0740ccc65d30f8b7f3b6a2e81dd96ffc
z54d4ca3e066773afe2b99354b0d2204cdc5cfdd2f3ee99ce69b20a660268079458f97ab5765751
z488606a858dee386224e8752e02cc3f68f119b71b5799cb55cad400c2d8302560aadf79fa0bfe3
zdc058de392108f5bc09da43c65c39126c3c8f1e8a0d2379cfdc6c7de100a349843c0d60597dce8
zd03ecfa6f9de49d9976f20f21fb84756fbceb3aea9c6503e7e94128a3e047b779330e07b62ac05
ze0923023898d8317f9f1fac1402908dcd698f894f6172b95183a26d0024e8beaea07edf0d7a333
zf0b9e4102a9956e95a1c002419d6366733d269bf9494c41f3a084ed25550148921fb73682ae36b
z267e6428cc957c951372f479fae9ee65b43d0dabeaa108aebb6a339e093ff80a05b0748abe0f92
ze4c0864a202fede4535a9a3d252c0ed2803f4676954612975306421d6fc80297fbf9ff05558bac
za7cc1d5850bd1096dec236ece745d1b92bbabaa2b91e7956d3bf7fbec12c81ffab5bb8bc3e4891
z6f4c515814f4516293ccd3215c47718d87635d4fdc9941be53482b5034c986a99d8400081c2115
z4f873b6fea25c2428fb0f49d9d47db1d19b48974bc09aa8d68afe7156205149ff54048a730bcb0
z47848039f5e76e86be82fb7716740d2f6cb8bb2fb451703469dace0900547b2e2d2108a397c554
z462bb65e864517f91e43178446ca9f5ab2a6bc393b7facbbd294645ff8f672be78f3e550cf620a
zd5572e96fcd1a943c1707a846c01551c7240f0efb6f52efd10b8e484bb8e1f181fcf3c64edb401
zf353585376d991a54ab2ff8a6ee5e5b50124a7efbfd7b5f720674b9927c1a360c7cd9b711f4c73
zbeb07e3e75d85aaaa13aa1f0850c71e54ad1a30cceb79d05780766f6f7a584fcf5fcdd2fe57e57
z3c5615f00f61d4cd0738a5af3b38c1c1876a8982ded5d51494b5cf7e1bf7e0637278f64f1a0bc2
zaeabe80c7df05e6caa3160b0788545eb91c88f79ea36cf27ba6f1779d00c84e1c570304881cb09
z116859aef98dd6c3777bfd03a0479109ce55334aa12d1c300eb8b22fbb3c6f663bf4248c88efd2
z969349216dac618e37c2b0b1efa2684a41990400db6ca2876386d8d4ac2151132bb255c979c5d2
zb4bedb7ecc4f6e93a0f6c38e23f52b8ce90954fe9110f95e7b69d6d8f6c25d1c8f20cb477011dc
zd1509f17e09a3d55fa631ba93698257410446fced1fb1992c9d2d9107d6589dd16750c7c846444
z978b0da6d9c94f8de3eef0d900abf773d3571f880c3be32d022ee3f9d437945e92952cb2badad8
ze17443e7edee2e0a07cf15b927c770b20144c173a059cc8baa09958dfb45ad22a2f384778830fe
z43b27ba3bd75a1e37e339e8555ce2d75e3fa88e54c8154336ade439538395381ff769331653d2e
z2036efbcacfc0f10bee2e3a83a13e385cf63b18a64bc5cc9f84fd71aca1b54980b946e6806acc0
z0dd6bebcfcd7ef1c4ed93bb6870140a319872c5d36084a61a4975231d21d96eb7a3b5c6de59ddf
z09dc40842c1fffae06685c5b1084841d3c4c6eef1292dcdb4ffcf711f207c7a61c4b0ae5bb3d18
zc19117147013e397b9100c224e811c8d1e7e6c0d2be3536dc3a3b286d3dd21d4c8cee9eb921a2a
zdb4eddcad631b5976b474513d985361c19bebef5abd8bd870858295b7d9a1a289542fe1d50d3ce
z130f5f98e57a847d3d5f21891a1025625c5221f6bf6a4d361c6229dcaa01d4d80724eb2459c960
zd62283cab07e08fcb39082a221651ce3971adc8693f0b3b034d1e632eed7a2e0093aab69bf20cd
z3ee78f7c3e7b9e231270c188e1c26c1f86e3d0fc964482cb8c4812d08c48d9945bde622c6a6842
z13299b770be948425a4fdc9d6902aca37d6312e3bb28db72846e0d11f65730cd9386a6ac2e037b
z29202fa495f5fa969081dfdb81f7b08b3083cddbca2a35555ee2d0e645947349ed6e9eb0874b17
zb1e1c460a519a46d5419cfbb1b1146cc7b57e314be61f0d5ecee8142db7014768defc27e9ff837
zb3d59c332a38c28c50f5d73b323a45a3e8ce546185c9510f4d5fb298ee16ca615efa69a837dffb
zbf91f5d0af9a6f81845f04993a97483aec8c5c0d81333d5a7e884e3dff8945ba572dba62ac155c
z9fe09191eb8d7d9240cca944e9947a5228bb2dc4f93d5d8ca1e89781c8b02e82e0903d6c86067b
z1b2b10cfd2440814c373c98bdf6f3787af976224cf45600754b659ee7ab1d4d6fc3f9ae4124bfb
z0a8d11bf58db86df555364f9760af739f2b6a7ade1cbe3f04d406dfd700ea8ed57462f378caab1
zd5061df5d0aa8d56ab15b9d201e6bd050c604aa9dd670e2a7e98e76bedbde3f1366f4cfe6fd7dd
zb44d618ca47f39d19969923608d43dd427738465bb54ba91755c48ed3205946d521b14d5ccbff7
zb37f910b6dedebf648c1fd51ce005c91ca3b6a462cdf10bc1a7bfb09ea815f9be48d655321701c
z2c27f121f872ba854a2289f93edee2a3a7556f1230f6b3c9705a30a37f3e1b8411fc42e1303c69
z70c414e632693dccb0387725c56fb53110f34470ba408a726a3bbd015887249d45079ec9c99d07
z0122a5df49294ca1c6d8dfadc5461e9c44f642a9d012916af058ce7dc57f12ea6726f8f585c0b9
z0c6622b2daa1725860229cc313869d49c16ca0508d503429e834b731c8c3432dc3110697dd3113
ze50c3910250b607e58914bd9c0108f828a86e53937b030879f3b51c7c65909ebad6f31ec8093ff
zfd963d623f4062b53ff38115f31ae74a17502f1f5b831630597fc22f3c1827e53b0ea6ac97e430
zc17e2fa5cc69932d03ebee22a529820f8195ea237fe8771d3eb39e718ad5cdbf3748b509d46219
z9f1da801f326762bc982b0bedabfef223c5ff7bd39c9bd33b6b29cfb881840e8e1d2ed4b77e5bb
z617cbfe1546638e2f62fe62e3ad086547e3565e1e71a37a7a10b04b03f46ba4007cb2704ec8ac0
z33afbefe7f47309f194466893d0268a33874ad684d7e8e93dd12d2687b5994a1b6f2597b1ad298
zdcba0cf57164b29c8d01fb56f756b5d27edb863b3eb2861e1cad441e1b4b1f7f0e00daf2d4135d
z737144ee3006dca19c0002e04c8697c77a7b7a681d1737a7bb2250e27ddbeef56bfa7d57afbac9
zfa2447a69364019e2ef2403b5292d46011e7ee39eb57bb4fb7df3557033644a5f56411e9ac5aae
z6491974efdbe0a5490521ec90ad86b968f1df041fd72cfdd7bd054befc6b988c6432940f4e1a3f
z88901d63eedc9a51134a0170d29338cefa8a96e74aa7ce28342328c8a909bf6d31773aa1f6ddcb
z0eb8fe6f221751c47a51b687317d4d6e50d872dda8052eac606f3a1562d595f0c7873de5149357
z244cdd8665b620cd659e2dc193848c7cef9a9f2ca45570716d29fdb9ff016fbe49de096f9898e7
zc13540e54394a428ee58f1e120429b74c7a7134cc0027b680f2bb161f7787327837ece9bb700bc
z49e10fee66f36c9e0f44449c7812add6e37a4e57bdb3d992f5eeb8d79e768d938a98f6a0a1085f
zee337e31e7a055e33999dc5fba0da821e8c846196e9d550cf3749d8c4b81e8238f4bddb663f349
z16e167126ffa87256f09744d6ccd75825a9d95eb709b7af62d5363c798afe42c3a2b1fffc3aefd
z18924213c88768feb42612170de78d1e409d7439598a62f4a4254294f192eb2a50d2369c140cb1
z67af67274c22af5417481d9c18884a9b64520096f06d84063a16d736fb75c7e5315377af038724
z9fa602d744223946932fdc580c1d0a05d68eb5536b888cf3245e7f70c33cf355f3fce6a3cef579
z1acdc18131cd33f91864cf5816d96a1f0df5b12bbaf1a37a5829eb2ac3538ba3b70d5545489b4e
z5a3cb5f9b35c02c106883b75580e09494ea75b7e7bab727b03fa1f6f75655e5d373a1fbd2bdb7c
z5c3b1e1e44e4e4572d59fe07f48fcfb3220eca9aaa7510b83b7e6baaaea779279e5818d87b8a2a
za5f82ed5e4a75992700d8a573240ada47851ec483af5fe78c8da60e73e19c09a6e35867bbd1b80
zb37c7e8d7d2305174744137b7bec7ec94faf42d6ebeae75be188e21ae0bb009eaf944cb3fb0103
z1cddc74d743ff363b3d262dcd76335859cb9cb53cb94fef7934d6eec495dc25af03a02e508b240
zf3a7f18f20cd0f89032fc0477546a4a05ec94bb311a63e01a17df21abe9b9d0985a386a707c39b
z9b5f140f830c1d10650802ce79b1e7113a50004c10d27263cc1e147e66d7e2c0f7ff6b0c0a8590
z12a929be926b8a63ff747ebf2c52754ac54e75834af5421b0fcf3363946a8df65940d3f0a8b8b6
zdab3fdc28f7e9f95a58d6de4a1583052a8363606bd50bb57aed51ba58dfffbaeafd08a596163d0
z6c74b7e223ddf1cf7126e7f420847fe1bd11b54c2dd7a4864b49a865071d3948156ab7a6fe4530
zb7ae357d0385bbdb85052b134fed09e1a5d3dc35acc5c49a7d68fa19afb470816ee9e4e5de8c89
z70fb25fec1948a71b82cf6a3fa3fd5fb07b5dd2f26d5dae8822560f9c766c51c14eb5a4e2857aa
zce5ddc5e735f17de73c153251e2f00300b72ff22101834e6292b8d41d377c03bcdfc77e44d2ad1
z5994e306a160ca36e603aecdb5efab0c54303ec5cedf00ee9e0f0d030ee8a142eafb94fc8ace69
zc354dcb76b3a1ebcb2ca9bd3c7d020df2b941417e6b498fe0053391f52cdcb97287fbb2d9834d6
zbc20e697d64190c1e3f9479d952982161f628f530669d0bbc18de4716b5a0e8f3cb8e9083c7e50
ze745ed13308e8edf20004c4670f465850b92f1ad34b744fed7def178d2a752762e5a6e68d50d62
zbdfa397534f00632228b7881cb644ce018236663ffd899eacb329c3901e06da69daec0638ee3ab
z6e1471aa32aa1ea3ca4ea023fffb4cdd6f116f4cc564561452eb61cf3d7443a2e7a1ef25e6d1de
z06d32ca527c326a43bd2918046fb6250705bf12d6f55956073d36e380746a370a525b085235a0e
z6e5d6f5514b7514c5b15280df81a49fba876ab97c2c6809dc20cc17a0d073f88a618905ece5ed9
z7c3b54f272542440227270a6a623e0fe1470d4168360c30e346abfc621ac3e447f81bb020ecfe0
z435c6fe205b8c704dddfa1e49960607ff27242c7dd2c76599b4349b3414ec2bb1d3fa15208ec3e
za4efabf87527480f4267fb095d054c0158d3b3b9ad5140b78d106d81fdac2059febc76feb430df
zfd2deb48223f21271f909c98782d5150b0035d620377a471275b60c25dca5415d1ca711d9eaac8
z462e75a771d69fc838bdd0da67fe037dbb2854779b2f31acc39e826b5fcf42b5808705ae8f4b50
zc82a61c235940999fcd2de2d5b31229194ee8094e37569e6d2c9b759ce0d66c311fd58ae0782dd
z976b85f5babcb26d889e6d345c08b2bbc289a66275c4c247e829c6837545e5624dfb71fdd0cec7
z943f69e94e4efa2c03e60f850258091543700fb646f89ac89b8b151b3e999f4765bb7aae151993
z6743beb5b82e6954868f6cbe49cc0e7e827c1e6b06beecdc1578c7b78e90d721549781a96ab456
zafc7cbd597e25b255e9b23b7e702a28a7e95269ab5eb62cba620c6e87bd23d85c4052d88558938
zfdde8c783132318b5746473b3433036af20d55902d9a8c66944a287163ef04b7f20b6eca3690a6
z05bc00cbd54bb62796b24636b835ce03d905444d98bd7e725ebda75f9d62744709ae1cf22c8c6f
z02e5f64b1d73475399f123eb3faf5f9091e85515e1d34f7b1f0e4a77f0050c5ba108525d2aa5ef
zf9d8607aa770814398dc9e5ca9e53c7ad8274a6527bee43d10e0d2e986699749540148450eb9c5
z3a4004239d97a872087ba7d7d8e8b3a2b57f1fb2d504ca984330765c82e6797e68de1fe75dd35f
z32787c91fa84b29ced143d17f4413200287a6fa6894e6fe013a8b004c912894150ffb21e3bdfa2
z7b2867ccfc20e1c9362323bf3e37af4b1947b6adc9d17684f536ef83257dfb89b0deabd3258887
z7d4634c495d24facbbed790fa7976d12078515b39a0ab5021d273ded671ce16f5a6db371746cd2
z6c186d312d0ea56740179119ea428857b9126f2988664a4ca0cfd02c2bc17eb8b07a7ba56483d4
za51a7d9d877c35195b634041c452640a9e8dd97ad61ec9dffa01b7de2d2257f24f087623b63aba
z8f195ec57c70f771abe7e5fb36ddea08c9a506b752483c24298163b49b251951863cd186725291
ze132c520cafcf18ed06afcf5d0f91a1768691e5d4378047fdec02df56eb870affb19feda1e2e52
zf6aface925827ff269a34d19857de5a3acfe971a4b0e746bf1ba563e58e9fcacddfea8af6d8273
zc0cbbbf20404b9cea6966a0b66af78abcab6695473f67993832abd85ba68e7a7be712d0ecf5a1b
za778b1eea1c19eb47bd007865976637c279b39df8a34b4e2653fb079d9a94400fdea499b7ca71a
z7fecfcf8d19ae4a1391912fe81857153fb92e89fd7466bb4d0f309cdb8974526324434fa889e99
z29aea15d192ca6868d711b4bebb61f9c9372d1718f60267a5d42ce82effe73a8427010737ae0df
zeca0246c0f7b0734f5c67c28a7fa3976fc8a9673ce3c552346d616a02d99d6d6be3d37eb35cecf
z54727358149956f4290c05faa39c8390922d1a4a69cd63fb6da77eb0960a189bff592193fd22cd
z09503e2a199a320d16c0b83cf6c49556aa19f3579d0e82ec9e06d4f579eda98bb2bfe5f1cc42e5
z73de3be91f7cd80a8cfed8be9e4a48d214b3ccc433c4af24e7f1177dc00e87bb64de45753a95b8
z970c2fad1ceadace64d80532bf7cb2c0545a7d7e06340d6a190c7857bd98273ec6ec5d9262bcaf
zae10a54713fd220b6adee9296d96411e0735569e68d688f0461030d67409a6c5f2524f4ced2f15
z62be2bbd85a92eb2af1e47663ac359f89b24525e8973d55c0c395b5e5f2e44872a5b7d22c00690
z7ab43148677676a55e4e6c0312bee235a13e41603ae4720bafd80ee8e26a31247fde8c4e19f726
z0a79dc7e40fb83decd6f75b5dd66164d94f07fb0eef4f815c31486495f50a02c78f0303a09ee70
z50a4fa40153ae1583f333e0e76128a744be15b67965a711b1b0eadaaa35eb1afe5b7dbbfc020dd
z1a500e20f07398338a2cbc65dcdf86dd4b8433b95bc1eb2ec634246d3f38d5b1eb25a564508e8f
zaf143fd04d527def97ba962e012a8de5024400035c5971f61c391ee3df2aac0d5c9e52c050ff2e
z39263c7b6b596d7b0133545b08b452a7ed51b0ac7561fc931d5f2fdc34ec7434b18aed1a831c4e
zb19650a8fdf9ef64b3e1cb8de65dc210298bdcfc43bb4423a6f411950f219154ab244abc205395
z39249c3ac45e40fbf0c695ead3a5465ba5ae19f4c1845bc0d9f0c24accdb48b4a6f44b81a22cac
z33fd8315a24f016b0aec4dcd552883948ee8e78a376664ffd025051afaab85e53b628a478d6720
za21f7a95969bd01c8bba9bd4089c2517110b164700c17d67393f1509deadebf906f5d9191bdef8
zd7e3cf0e33a15bdc840850a0f0101843d52596740b58ff42b28067fd682e2b170dde1fab1476a8
z9264188cc43719ef25caf052fc09f8ed263bb1a5f32c357232d15497d63e07db0084a984334b6d
z0be0f95be9e658351ef5046c4db2ed2d1479242324a2cca136c68d2c772d08bfaac075017074ca
z29426345ef5b7af9fd7c3fe4b280d82c263d038335928ee32998988770544982ceb02553ebf6b7
ze59b421320bef2ce9929adccfa1e507406258738472ea36a49853706c547f13603c68aee9995ff
z5fefedff61382657eb5d12e6668712e979167d61b765cb8304f68b81bc6e4991ffc3147b3fc4d8
zeb4273def9141f558840a37952dd7d7e20ec86e514f8bb889c64c1c4496f8c3303c53d44ea337e
z83b05ce98b76e4013b6c189a2cda20503076417949174d03e65d93169ef251804a49e85472152e
zd22dd80a6fe42ad67b046a561fe307f6e237f37000b18950a6ca4e14d77354de496b24f5ec4394
z5d6257ffaa972edcb7f376664485773eeec605853d80731ddb9c13dc9206471b699cbff23137d0
zfd3c7321805800db325e3aa8170dee2e55f5598f2f40b5dce23c6cab79f10115b305313053bae8
z073484ff491c29de6f4a55733f3b996e4ce3dc388a8c413dda2e8b52c563e816789bf0b7718c84
zd246c4eed6591d966baa66ff53dca9afde1ddc4327709f88216c84449d216955612fc74cbd64e9
z966468c94e5ba5d635f3eeb774d717693dad1cee483b3e4a477b0bf1690c523af236d125364675
ze0e8d745d6cf46df06cbdb6b956170f80d3d046b0b9d350e3fe3c9212e2e2decbf0e05622693fc
z9e9062a43ec106967c0abe22632116cca48693af618c69ac2a94d0b54b557286f2458d0333f490
zcf64e6c9cdafc5db127f9e64b85caa13d2ec11a0f3e4579ebe79766db36f5d92eae032250624e0
z6dfa996b5906981b74b7b3d1d15cb754938df14d53bf6966dba4fc7171d65b5f496bcaf17e84cc
za2b0233a40314f74d50fa3b693ff04768fe024bc05c386015a90e5d4aa51ebe8bf42d52dce6812
zb4e1bf1242f1be203196308da4bed0c36d0d1281b4831d424a57fdd1b388077d10179fff9c62d1
z99c9cdec973188ec20d458a326091f888384c213875842887faef38f321ccf117f2061fb122292
z325af7f0a52d2fd129036b2a28a5561fc0cb774e0c86d1b249868f9289c89e485eb356832d1533
zeeefcfa4c6b067161b1b73364ffd5166b838f628a2ec2196666e7a08874ad238a11dc7a7f6c658
z7defab891958c8e077cf20cda30175817454f7b97a797754ddd9e15631b3210358fe78483fc4f6
zc088b121815b0edbb764b08931688c57ecb4113eaa040ce9c65eb2b9dfe0979246fe7e10278723
z32a18389f0c24de5ac37d25de15e24a63b5dd95435a22ea577144ae3108616206a9e8fb86e5333
z9ad2d64f97c6ba87a68fb59e5f7a5c8b71a82409de0af046f7fcdee1daf4a6866bb2d2e0e148fd
zef9cb4db327213363fa4a19083d70bf2aa9b69afbc1b92a76821543b4ed79976cb260363e95cbf
zb07f75ddd148ecb8c1418117e00cd899652436b68d515a655fe488da34565005e20370ef59074d
z8648e607f5fa23722359b06c4bf55d543776a46051e2131428454951415fe5c3908d74ec91d4f6
z79aedc1dbdbdfe3235a17abab567e8c80385646790401d6979802c0e7ba89c850facf75f9cfc8a
z008b551fb45b603f64105d99b220fccb7fbbb9eb3a71177d5c12d1f663e635df6757b22654e99e
z97c81c274b6263bad399e388a3432118868b36d37a733444303cb4025ad21ee78a1f195896f3aa
z8cef0ab601ef239557b86a328444576c8536df07be6dad61bd6e63427d05a13882b16aad8cccf6
z56216e1e2acab5fefa61ccbfe7284fcf4926698b3c73e14f67734678068d80eda1b9538cf609bc
za68833361dc0e437321f228d334af2c6618a0bda657a9d042d4e2e8e1a80df1e8045972603bac3
za88b695d3913a6a41fa22dd960cd1226e8c8045ed5220ed9f28eeb3d976ca089df218d91a9cb1c
ze58d0267d5772471feb29c64a10bcee1e572bb7e90ca092592019668b70ad8bea6f6c87723a1f6
zf784131b0c2bbda5b820f03660689e538a892058de5a818feb30917c11b33df5654cfdffffa43c
z2272575be383861c4d77c7ba412ea79f04e5af9eb6d71a3817502a5937fdd656cbacec361780f5
z8913efc9686164f179243484209191c6442fd81a65cdb2100161fc999a65d9e778b3cb756caf6b
z0c7c5eae073b4288afb5ff8deb9b9780927f0f488bd12956b8291fa8dd27b04f14e19c636e9216
z80d3bbed073a000e629675d0ab966166c8b08fbc27101d2089c2e2d2b7dea04848d6ac949b86d6
z4a5114223ab92603b3aae2e4ac23a11fc11fcd1ecd66af2b142456f75e534e076fbce0352a0a69
zccd9ab28d853a11151026a3ee25d95b4898148a70e9d9e9997f1d6e37a1984bd04c4a04a149929
zcecddcaf98297a4a5adb350844f48ccf84a32ae5541425eab1e78c5bbb867bb6f76bd45784de54
z5ed265fd4b8adff30628d7867730a059de0c72d92b1df5cbc82cff91c0052e02d9238a30fae398
za16bbdd1d1514e7e6de739e8fa1e4232f8f7f7204c133933229593e46f103f2e8a2520eea96586
z0cad586843a57451d2d53e7916516f955482d8f992308789cad72df5350761b39cb33fc7128f6f
z9375bf0205cdc5f18bfee9de783ad55096b1e3bb54b86ca8136e87fc77ffaf516e7b34c36b7c80
zb347b33661c85ba44715dbb5f2366d87644771f74d2bef54b57f45a427b1c14b75d7624824c3b0
z53e38d85205d522e0c51c16f36366f08d76403d4c61edcee3795fdab32e490065b0a6551b0de66
z8fc213976fe5d854af97c179df53f406450e84682e1caa3c8caabf07c2a5cc11d9c6b46eb92fef
z4c2e439acba5c29298c9745fa160a07ce26e508bef5d58b727f626942244e7d7f655b9c31d5d90
za66bbd6d3a18aceef5a2ee54df621175ab502af058cb0fc2f092830553d2dcf58bb11dab9c7e7a
z744246c94df2b73b4a668c6effad460e290e4fe2a13433f4ea4f90e6c51a5255df8541628c1355
z1fcc3c99e62e54e8000ad03b02c7905d9caf7ee5eebec28230fb0faa12f0cabf70470ba8af786d
zeec5006edbce71d83f4447a9a44179c68c7614ccdd9ba6abc3e8557487665150fbdff0bf3b37ac
zc2aecaebe1c0dd7440b28a4e7302b60c8d65f1e9725582d3d64bd6e25d438e842a31c6fe9acae8
za9fa9ee539dc5f38a020205be5851324bc7afc686d37d07c851e5a8677f0942033287fb5323913
z7e12435cf676c8cb7dbbde7d7e6bb5671923b5cdd7eb79d4947a5a53644a71393ead24c74c7edb
z32ccf357d532b2981956f925ccfa9637526958527818d5ba57a18cca9f7664890a6906b049247b
zb720dd02e30d20c881de1086d58f0a57ddee8dd7f55a568de1122e8c620830e766fe882bf724a9
z8916773edc1d0b28cf702302de5f7ffa248e8a2e6dfc3afe45ae7ee27f9a57d42ae16ab0058314
z06a5fed3b7dc107f93ef160a74e8c6a83b99c17557fae7182105d3abea81ed3b23b9081542136a
z8252865d89d304997e3c4b086e5913b344f7d3637f63aba854d37d9b79672468b7b0d28845565c
zd02212bb5adbc8f5126287768937045461c27cf60be079adc7304d9c1481a3e85cdb60955d02c8
z1f5f1f161351d92714cc0866cf3dafbc69b3351d33749b0b9797a7c6c985a6f8c3dd907c2416eb
z6e15fa5ab394aeffe3ae174f848310c17e5ae7739cebc0755faa665e93e53de1c0054ac558fe2d
zff020ae03e2a307682ba83f81ff61ba360b4871a98dbd9b7dee1b5dd3925430b62df2258e3028f
zc638bf0532bce01fd412beee901aa4e3061653867bfab49adcc19b9ea3beaae7425d707ab6b5ba
z3720ae873417b6e0273415167edbc8457471cc55cec182322f744e90c632953284ce62fe3748a8
zb19b709fcc41ac5de18a947086e4abc9554d5cf079ec8b2dd68f11ff67fc280b628ee54788f999
z3c45fc26cb599ff6193ee876cd9ea32e6f1e6a46aac0a7cd4c4aaca80114f9223eccc87f7a175b
ze18e267b2e89ed3f2b1899fe4b4295178c7006248f3d135e73ca995144b0e1501a534154053dc9
zb2708cd19aedae19d4d581b88a3475a4314c43d7ca481a0581f0dc77fcd0b0bfad56f3fa43233c
z11e6e3add6ac9f803b004ed32bf2dd29dd1a65daa02ad74a39039ba8c4203255977286f23a909b
z1eb1bd9525d1c0f8da8d93698d2b754898db0060d7ed83257398130e317df3917ab76e82313af0
z0c24011f118e1bbcde0264f0686de641798efc5e92b21d6dec089b52052c69b3c41a746c4e18eb
z528b7875c7d6af025d5acfcb954f67bae133458bc5455b436ae3989c9c72e7985285bfa5bcdaa5
z033e548e1c980687b6fccbdd670867140311a5a47c7818582871c3c00bd8c5500eba0927d7a378
zab6d5f3c81c68a4a4e9c0f6321326bf814b465dd62e992eaafa2c50d1216f0e3ec3092a7469046
z3cf3f63afecdaf3dd8dfd56192657f4c3dc0b1f5ff5e02a78ac8c8ee80314b976b6c3a2f204ed1
z259679b622a4bfd2b93f830bef2f853c0bf2627979c5be8ea336d66954aefee983daa07aafd156
z632a56842e40ce835a85b045960844608ed86d3d4049e9aa64db4e3722f8b6f0ab1f015c45ff61
zbf7eff8a5f618a6ca4b45f2b1c2900f849e1700779116499c4d48a83794e5643d0cecd028572e9
z1fa32b2f150f6fdebd54baf54769dd66f62bf898313b64b8194b71c7bf7718c1aae690fb6a59ae
z95ca58b972381ae4b7558a98daf33eaf661c3c793f6f7c8e8bf9e8157c60954481cc942c24f049
zb9758d84fd18b43bd00c49724f3dba4f3b44aee620a377dceaab6428f7f8fbdc09f3696a984aaf
z24020a5958101844848659d18ab9fe15cddabca53425a739a75f60c7c7450b17be879a308cd5d2
z99a7e08c22b2ec08e442721631651f54ed6cfd138f1650388b34c0cca19d20831d8832e865398d
z82a869213a6dbb9158f97f783b632e5fb88aef5f6a96419c8d0e67e4214fb41f6eecebdb41556f
zf3be18b596d12369424e940d5374ebf565f44c5267c138b4f1dfb92fad534d2eaecaad7202ddc2
zb2d08184e3f5235f7cc1de119193134a84045c37bb7b5e910944c8b8edd16faf2e71b526bcb914
z0f296f8df28feeef17f114a4383feaed17ef666fa379f82315f2ed322b67835dbcafe71c85edef
z64895edc951bff9100f5690477f69dca4484f1c02b39a31b509046b05a8f7c5e60042f98156834
zf10bcb3c2d2619bbec5133b11f99b64100151330bcd5556ecb86b00ecd6b5524ce6f81d149d5ea
z2bd4013b8a0d6e2b3594d8cdfa584552dfc7786b31a4a17ac1a124500057ed90bb318cb641fcc8
z904a1f8b292ef365105277c50f84855c9afafca4087481c6928e9dc7881afe929df2dbd160eddd
zdfd0aedfc6e02bf0d0a25b1a68859df5361058756131eb15c38b022a4aa3baece832e89f802f6e
z99a83c5d4dfb21e4d97917389951079857d583cf24271a64682ca2d6c6b62dfca23dbcad2faa34
zdc2b539dd07e7df85a3a02a941944f2cfacc4beb51cfc0cd9ee56ff8644e97ef1cdd7214c881eb
z917cd63db55bf8e9e3c6d1ae43f532575208044024b813a409397fefc6030283d96e16c80d8539
zcffdfc027f1260a5b06a13056d8bd3ebbce33e93fd3f8381deedf10e6e11749e0e3654e34d85ed
z47fab12010bfb7a1962fe9344556b44d7cf027393fd9a26af581bca6b1e2ae3b26458d8c2232ae
z7dab54be743fab99f510eacdd072d1becac4a2021b1bc2bdd294a57f22f4abfda8d01a475ec918
z5bf54b3cf5c53fbac7fd66094946ed1bf17b8c7e2aafc4f90b85b6e9a7ece3581e62c2ba43f725
z2fcb15d09df95e382c0660f54813444d320c42eaea02f3c2d76fb319652507e8ff853cd345d2ff
z4e90e2cd6f584bffe8da604b6ce030cc818d641e1aeb1ae105558cfd2a9f97050f576c7d8580fa
zd307d2b7bfed80e436bcb90a4c65b9ff14e38b919a5c0f7f5f07721e79cb38551c825a9c066f08
z8c43655c67a02dff08adbb15029cda14cdae06526e9382bd789963647efeb85eae417f0d5aecad
za9d29d6ae3290e5bb8b25cd67aae68edfaae7832ef2230213c0f7c56b2f1ebaf0c410f7fb04d1a
zf79f780d7ac0410f0720d0d05013878eef760bfb4edf0ebb0b9161a2a44530daf45a76959da2ad
z9de454fbe6ddbdd631876b955212c309cf91a5c1609830e7a8ff8c4db5c9aec4192bb761ab2598
z091c0718dabfe81b67b5a505ef9d90f5842c24a14f289f9b3a168f4a09fe6d66f18368782b2fe2
za6141e256bdd78d0d3f4fab600a82dd5ea36e0e6efd99e5fc4b6be55a119867df2142def73ee4b
zfba5bc33bbbcba887c63123c420aafbf9070c056cbbfa3a411c0c35a54257994e68248fdef1303
z93d5b0daa39f6e356186b9402a587586d24d8bc5a5cefbb55e406e24b9bd91eb138f1e0a09bafb
zf423f714ee45adc84f8f6e0cfd62e59e5b1e8bbb5474b1ab780c7137eed831f0b6100465079884
zca9cde6bcc3347834c8e13c83ec2c93e4c7b88bc0bc62eaf8d245add226b72b868400a2a3080c5
z6354b76cf6d48a030d28f483c9a79bcd11019c60e391b69347aa50372746932f83a856de4787d3
z90e3c0baf7c373d5fa5c955402ea782f61f372b0738adac8d5aa0c62c87fe9b988a58087cc2d8e
zfea757f3c5ad6be546c4c05a56a6cd4ed4c1f5656cbd7950a0d761702d1ea823456ba1554ac638
z4420ae49cd26195c5b32d86cc26aba486eae9a4cc579e6bbeaeeb7411bb0024cb5810548960837
z49a6cc10c83156f2492329a88c1d84ea86f91c84e15083bcbcb39512f9e6a8efc312d44ce4374a
zdb2dc7f2150c1f76c4e275f9f8a202f1a2f7b4a594afdf006151dc383f59b4af58fffa6d6fe4f7
z8a4ef0c2d16224babd34cc47e8ba3c69a8703254206eb47fb7a61e3f4bc157f8744d0e45356cc8
z21a94d2206240a9985f2498785c7c9eea181d31cba02b130f5aeef443f8f4202c19759ce2ec740
zef0d007d2c1d2cf43e63d8cefb3428bc51350e7245b7efc3fd1f54ae3586b4f08a423cb18a7c8f
zed6aeed062a9d56dce79cacfab7f070111ca994bfd5735232296d07e05646f48bdfb69165985f6
z5c4f98e1a9d65a8797a49a6b74dae3fb04ab61314e306d70aff516b5e9d1583744c8d78c40f5d7
z0558d067e9b9e26f9a9fef8073ea4a78f1749244ec57fefd7f6501c27a2b1063202d370f3317d6
zc6587c8773810815209316e79a61a3ff35c72e388a23b12ef1b0c96180c52561434624bae47090
z3be7a11ba0dc4bdf9097048ee9df5ed8dd5aab72e679ffdfcbb4ed7989483de3da7ce8de53fe3a
z1f813a44f28c51b01c6803b11592daa6a89d2328cca929d00089b9a586d19e11fdb878aff17ee8
z86a59ff2f55cb79e784157f871f3c6c130ea0c15d7dabc87e08c9c62380ede1c462801aad3d24c
z95d4fca18d736a04548cdd4eecf38a6a84fd6a14d3b56ae06e0d12c417799b636d33ca728340cb
z9857a3d2338e9944da95e989b90fc29599e91308ba3710d7e9a7c7c3632469940378e292a79c2e
zb0e1bbc03b192dd4578812dd16619f8a2138044d5c280ef674ac581931fa37f98dcc244c71e0dd
ze00a72b08097787484ba1ebcd5276c7d98f35a0b5ddbab0bf39202bb8402a957396c5c12f6aab4
z20c9e4a4a3d2fc461ce15b326aec865ae110113140e41194579a04043181e443eaf050eb223152
z625a0f7e402519f5f5750529f832147ab434cd8fb9aa23dbf597968147e2ad97276c0c3caefba2
z3616fc571ad91f29014f9e4941ff5e3ca5ce60321a5bba3e4a8c9ed1a791119e9809107800bb5c
zd98ece843a365d158d81d06342bb170b19a32de141476cf07105b9ef5c1be03c04f062d5cd2f66
za322fe9249a1fea7d34f6399bff831b9a97b3564afe4ec8fab526e042fda7019d1f878c90f5fe6
ze19b326abae533556841887b1da854f3c305a11bafece7c4feeb07a73c1da61643f1b96e500ab3
z701e0d8a977b29320f7658a03ffb4226c0ec2ef34e2948d5d35dcc88ee0a56650aec784f9eb217
z1a37d0fb6ecc51959e97d8ad5c1d60e6b969901e3aa80af11378378107d095c88c91cf72fee958
z98a0e8056ab9f0f2ca0298c182f58729c9b110e67071121bb99a44ea57dbbebd1a5e9394f16043
zca3bb711205c3e69e5748e13c040c04f57f3e81d3d55b788a83625e5a21f1efba874420c67efcb
z8eaf84cb0a651d679de8c6b41435466a5776dc5e3c150b78b0c1259308aa9ee6ee7868f4492150
z301515de80d1a9884e430c1e44ff5c813e8932d74eac6c932035775c05e72d4e68ea40e9633246
z38e07152c97716baa3cb3b1407802e53edc180c5419b866a649db1400124ac2e99019b99e1644e
ze7e041c66cd5d63c8d8f17b8c490c3879bdec60835656205772df96804c7f9ad608ee49ac6403a
z686e8f15eecb6ae489db2ff07f62a6f63f266da8dda50eb0d53cfca2684a5cc5ca84406b940ade
zf769ee1b0568c5501d7da6b050f42b1e6f2d994dd0fe5e6c125e60e9f5f284cb60099db9af1426
zc82f832cde1f30286fe20c4f48674f7c837280efa0eeaf4d4e95c7fd479c105c00349a590e4875
z120f4a0dc9356956c53f3edc80dcdb077c9a34c142902c30b5f39a6c468f90846897f909e401b7
z9d7b6afc2e119f613bfba9c548bda677a151a56d994f1f82ead43bd407f2081e7f5dbed04125f7
z054e26c70c73bf4e76798a98797bacae7bb78e8208c90a610bac732e1f64eb3d8884725acd52a5
zb9321ac0a5261891b91a6bedb5e834e2fbece81184af3c16a34064d0a3ce365790202d19eb6e91
z523b27aa88e5723657efba11ca9ba09893e5b45d448814f0a6b766c8747e5bbb36b90d653cf2b7
z9d7c024d0abb227a17f9fcaaba32221e0a98dc8fa837c7ecbdc91c7318b97d6df2cbdf11f740dc
zb459ac4149e0bdbdb07374df2cffd4debef2740544700793e910136c2f1616652c79850bc07773
z1609fadd97e18027cd1793bfe9f664eec1a87d31a48655d0eecb28460dcbfbf77784b8fab8ebc4
z9b2dbcc02e49f78bdc1c0ce142488a93c37a68829c279d63f86806394ecabca9795b009665cbd5
zd2a8e9f4108018988d6bb2687f7d8f47ed5546a9c72328bcbca1927d501c8515f19e38c23bef5c
z406e5ff89cfb1395ce081d7d8a0a27079a5e1797eb998e40350d860fe620cf479c08a8c2c68ae0
zf8b886e9d594c1a2201b312a77752915e9d032e18ce4e1e39d4aab282585900cd5771e2b85f489
z72e2befb8619a0eeeb8734ea91bc564fd69219ecc4b14171e9271f22522c8a3b6dcfd0aa73a8ca
z9a72d19108c08274daf4aa17ed11ce998463e7d31a538550b5e5cbd65ed19f26a3f311edb8e9f8
za75531d0403cb39678ac90e66015f5855a6d655f198a2310ace40db80ba6e5acd1f1649a67799b
z93d57ac75beb4e6af3ceadd7fae5788f1e63d389872f1d758fe9c20c8952bfae94a68b631b8336
z991c316f0a5348d3ae4bf9a75623c497ce151abeb1351b42cd23fcd2532ce0ea14b8fb5b09a0fe
z4d9fe8294befa03447ee794130f9c0746e72f1373a51fafa26a5b07658909e1301a9870654b597
zfc447c74bebe0103955503964e40b94541f01b054dfc234510367ce0c012c277d69b133633a8d9
z00b842b171544962aa50705b086fafa00c3fecf5de4f5aaba8b8c1d0f38a6a28014a7d0199b2a3
za1e716617109a0c979985cc2a045dce79a09f1596e77a0d0c6328bedaa56f2f657731aed8b38dd
z03605521844ae98641e80ca0a081802837e6e2d6c06f84a30c6c7fb029772f967c1983191d6999
z3aff91408954d2b7c19cfa51dfed6bda5d0dec0b0c588b4c7d787c2f2f08303f573378239fb261
zdda7fa704e0875126091b897bc02bfab65fb466ced1effd9d62d8dc700eb397091534c257b5902
zde32f44a332fed3687eeea9cc9cca44f11003ba49a0669037b40d917f47e89b5904aa919566469
z23689eb3d7844299d7121e86640308c37b89ed21f75d348c208808f3d928af877f69a58bd402b6
z5213bebda88e40c07578a806a30b78ebd5840be65937ad3e5be5374e79b639c5badfc0fc0c5b70
z6c1993655fb54915e5a8f82bbd873264ee45fc0776500b0c8dce8bd026f356034d3c6bdf340dc7
z2c817ff4b25d90fe04773dcceec83c24abd23da665025874a8150c04a0b9f7199a8db18ad567a7
z9539e37a0e2b10436c27ccd085fe9a049edaa8f6493cd19074949fb5b07314546ca29cb983bfd2
z0bca37e4fcdd97821f84e96a9c11b08ac0356b0938939aa12b708219ebfad71758503fd154925f
z6677421c40dde92e2bc9e1e7a7715773d2eba59b48ec1b87a36518a4cec7c674a822750f95a386
zfb036d2e3eb324c96513f83e7483275245d691f394de3c9445b400d9dacc3384c1623005c98286
z49ec629a107fd1befc35bb2b8d6bb2a05b1824052855504a57bbdb8105038e5249f05f2d9f5619
zecf1274b2a639632db0efae001ac768004991a10155681e8a419be7b46b51823ecfe686a17d142
z06ff1904a62564eff2414e41d7a4f5e85214ff702d90d0bc8259397d4a5cb9e1ff944e94447d08
zc69b39906efabe2b4e22b46e23849be9f96ccf2c1cd2738eac7488708dd98b79ac10932a93275c
z5fc55a57f9a707d736f9cefb981b8acd65c6f951cddf1fa93a0da41afc984f9754d80cedca25e2
z33c16efa43289245f3f6f340135b70fef289085a70510ae8e792c05ae18ebb5efde06f5c0acd5c
ze9935b76d524d232ac438834e394c1322a1e4761df37360fb6b1cbc73e94ad82942a121fab8789
z14731d22e5a05b811d0b7fe1da9360be9b7572f7633ae39c2439480653598aae15c408ec4d78e4
z4df3f64bca135816f8156abf0dd3bb62c13a06384f573e0bda8344be241f24ed3263df32567647
z6a35be9f78ba10e30efaedc712761e885b34460a0eb95d01811bd1bf085c740dbcfda25fe55b80
z4349ac9027fd05609128e40fc82c0a41c46d77729b6500c6bf57152a31f0f105ddee8d857689b0
zfacfc7118d04a12da598f36a8c2007756876ecca28a527385625361a243d872a82b24e2ba45ea4
z5ce4138bc56b3505993fd0d84e596e4b5c5feee4fc8e951ca73f83586496151ed08b25091afb56
z0fb844f483e545ec4a77a359b5c6da174359410e31dc78289d7dc76faafe62806344db7c15b19b
z18e6f754b55574939fd4be9cfe979d97665c49afd4529949c22c5eee21795491baa2c5cd552071
z5fa40aff187836f6136926d63ef41526dcc092bd116bb608d8cb0dd30683161b6dd9a378276892
z6e302294633a2a9b46f490760b406e373c503299c3b1a192865523d591a48ac5ce0d7173d23d0f
zddd0953abddfca67f37328a99126eb1d42dd0ec43adc04960dd1c71165aad00532ef1e4d9763ca
ze51e58bf0eeb5ba7569f8bf32e4f41d64689bf167baf6b5a68f9d55ce2c0688808b7ddaa27efdd
zc088c98479b5d37754809794ec5834ba2ea80b16cd9c19a40185f53dfb496eb4822e02fe0ab3b6
z76e64880a8ed5fc3a3265b65555f9309323a1567544ab7e7aae48c4961a349a008725da0ae59bd
zac894608b71019ef759b271a3df2b9a2a164d95d6b821c139cba34ae854e05a6a84e1f523eac28
z2b0d5e40263a45cbb0946a1b0053417b3790388a0a3875eb318cd74a7032b70c007efc7be4c315
ze7528537720fc98098dfa699b02f8d4c9c6578e973b5779753b2c91dbdce3c212fb0bfca32f967
za552a6a81a563ee13e703881f6c6688df338be00cb7642041b0c4de3c750296415bc4166d732c3
z63ec5f91e4e4efad04cb9c22984c2470eff3162b638edc848adf1bb0f5347c240a8e79f4444d60
zbd5a68302bd01da703138071f53133dc942fbbdb71e9efbe40be421ab0fc43aa311e71a6f7767e
z0073d80826ce7556d6f3745c554e99ee14a6de647201410a157114e15c95881ad6fc6835408070
z976f91d335658a1b34b5a56c5996b20442fdb17deeca10bcae33568d0c646b32381e65e4f2fb18
z77d7e299cbe962b845b9b7f33189acde7384bfab0f0f460eccc16595a2573cc0df7a793123664e
za843b5d2f7970ed7b9b680dc9f4ac4732011cc8efac627ce428c40e4e7a2fd7122b452dfbb8e7d
z93bb63e8756d725f9ae6d76edd0e7aae64bdb3f61359abb7fa9328d72bdc9016e7e2525f5b724a
z6f5968f28582a1c5c5d0264d346f882c2ef52280dd933f3a114cf72e8fa6791e44cc7713201dfb
zf72a8d6287eaaa7896695f396c35d5adad30bbe9301b09130111244ba2b43bd2ef4201b8a2458c
z9c5672ffeae5b854290ed7f3dfde5a0bf5c00847b5a9d8736cf382fd7f78d9dc2d472ea49bc59f
zdaf9217e62ea51413a322bd33e0ce94d89a1874dbcaa1aa4791efe757809be627fbc0355d3bc90
zac6502261e70da8319abf44ebef5bc113e56793af8e44ddb6051896c7784a4b70a83e44fa92a51
z97e3faf42455064e91f3c1ab6ee8301d4615ee54b0ad5b16e8ef449b37c4b65380cf5529cf51fd
z77af5b513dd91d8ae57d27c2b3a98b0fb5b563e8ab11bf1379130f09d2147f1c4765f9e6b7ae97
zb3f5ff3a805cd0e2d7c7d28842d838fae7b6444491cfea88040cf00967f2313ebe3f62c14c9624
z1ca740aa3918c27a68371db6805c9b44c74cb8670fdc6bc22c64d2c5af588c0360d0f9e0c5f796
zbe2f1eb6fd69a415ace1846149bcfa3da99889497b87dc2a7791226907736393ecd490284d9d2a
zabe7f38ebd9df14d84361f2964ae7ea737457df96b198dc75e0b34b1c070b3cc5dccfb68507286
zef79ca918fb7826a170401ea75a66d2b6b4cfcdfa07c2874162d4afa78bf6e1210850de8464be4
z399c49e6578dab478198f426676e339848321a2b5696c7dbf75c530236c84f6b2d523009ec3622
z657fc29e7d2b6050b41da8f82efec41b59d639659e9833b460bea0eed881c669f4b2508a061dc8
za5ebffbf17874faa65015771941a61259235e267aa98e46bcd72711d5c4ff476c91c4123e27c6d
z96ae0104c4629190e26ea4fdc7c4bcc31d2beb15315fc2d36849ab7dfaaa4bb4694444919dab35
z057226341c2b2e1c5821ac75d32023b15c01caa21bb71e9d4c34c0f89100b28667f854e48d49bb
z641f9bde3fe10e2a9359dd1b4487effe64142e8ea68c6b2426124b3645cdf85039c93ed04184da
z2f54c3678e6016b8ec594285649733ac71bcf12010efd5196c33e868480334b887f42be5a2667b
z59927040c3a004a33ed3796cfd4a5a6be881575025147d199a6a748d8121c94e5754aa1a8df611
zea21365a2585b0fdf5ee14607e62c7a9f9bdb3dd308f13123088126e6f9bd09a52cb3eefe54aa8
z701e4b8ad95ea8003956f356fb3b13954a786af07cdb6facdf55ef340c13051b1c21945ec5a4ff
z9b462707bead6574a0496272240ffe09d81772f4d9efa58085a760690eaa5efdaf594dc2aceb0b
z11b2afc4d8db91bce896666d3083c280e17bbaa4f90ffc927319259ee7b1612c281b0b6ef4a67c
zb2443e2e995322fdd6f6937b5a73881d0784c1733719a7a04dcf640357821035a9ceff2c5490a0
z8104a64d6beedcd6ecf8f5b7ffb9297c6a8291cc1906ceefca2ec0c24790b56945b3312e7ca0be
z045fadee7e79d46cea34a912344abf2cb796b5b58b7e6f81609161ccfdc16e46e07af093eb5b71
z84ad703e4ddd87a3725442ede4a0064b40c7ffab9ba7fbfffdab1047a7f28c1f43bad1c31c711c
zb335efa626bd903db4b6cb16c7412ece7cf847052f41552a74bc67cf35ae73f7301a74528beca0
ze319eabe9c647a95fcbff7f0d375b5f747686163f82317e86126cea9a8061f4ec3f56dae322ff2
z95345b32e3bb99bf3cbc0e3d6d380a8f74ffb3341c175f72231919d9113d232342454277eef49d
z2b4ba94be3e65a577aab856729fc80a57992cd79f6a463486dcbdb48d1ccf9cceb6ef7fde3985d
z6673bfe348f7849a8a496831a4eec38f8b277fe703d4b259a51fb08f0d37a39d845eb8e01f1685
zf7aa0f8b64bc12b4a538229e5b4c7386a187e5f8e81a66b0f07811b34494d38516926547cfaa2e
z5db71064e802cf9ef11d0e3e598264ce920ef5a18fc2b387a5340456e3dafb7d3e728db334f0d0
z913ce52335d7bc5a525d7ce7bdf1ef1e076d8a8b4cdb32ed2cd71903db47414acc437d1a2dc135
z672d275f95bbbff8786bb21ca6223f31ecc677b008f18e3e8b468f12b3d2720504a7b00d08d8c8
za323727762c33dc6d79a589ad81686e908e57d8b4d712cae40023206b9999c55f3759821beb1ca
z8558a964a707525cfd2b2a312b1af78e1ba9e77c40172f48de43f2e20d456a91002c1fd08011fc
zc66988f0e26bca5ca67af5ece19f45aac12df860d0a051f0328392d88c1b5692cdfc5ee450144d
zf027b766ec3254b37ecb00b0471941caab907bafb01a7357d4233b047590c058de877e221bf178
zb9a8ec6e01739a1682c07c0df4a61cb9e440dcfc17731c8ee12343af680b160c0185544189a25a
z0f285e7bf00176c170e6d419de68e2c59004d57cc234deb70a1c49a2b78761d216e8732589110f
za118d4e2c4c98221ddb8ae03a9153385258bb13a8ef19da24242e23b4a9afa9558401e79e54628
z17fe4e597cf2925bbf6d36fb9edfb7ebc5d4639eb2d16751b68d43f1bba5e28ccf1abc66a190c1
z8ed36cd845bca245d095061a4865d618b64c8a760c752b435fb92971daabfb32e43413e9797020
z2bc49e321772c401a54c6d10ff5cf92abe1dc437fa02632f4e45792f3ff2910f99116fe067dd00
z190b418702d77f2ffe077bb8669302d26a8721d2e0a6ffa4486e9204779eaff3638f9eea2ea31e
zff202b4ec5f0142feee133d20de6a561154823b0296f93267ea93fdf9e60b49191edefaf03b266
zc6ef9bfc279af7c1df1b744aa03fdaca602f3ff7233721799336f07c9656912ef1331bdcf7fbbf
zc0450d6dbfc0afb33da196f431b8ffb7bd68913332ac98b1d29af55062d6b8124259675fdf315f
zd3bcfea853d477b4b109d5c4f4c560ad5b49dab52fab3ce8b5764e4e4db97122fbb9a982de4c74
z2dbbdb2a6ad8580cf400d44cda58d02c1308a00daf479098a92fe337b56ba1176033ae869c5e61
z40495b375a92246ef2281884c249664b1bbb6256882535ba1e92c801bb6cf78fe90ced780bd1c5
zac58597f16fcc0f17b396b0071d9cf22f7f1c4cf0d88af210f390ebadf94f5b8869d942bc974e3
zdcac381d4c2dff2df2c3b450e98e29816e0059ab438a204656e653f61affc787408a1e3648c658
ze65afe6e811f42b911d8dcba8f593cade5b8bb0bf8d7f71b8b0b4a5660526b455729db77216a2b
z18b7d0c9749b41acc1d6684af667214a734ecb591d6e2206cbedbbbd8a8db852ed0fbe284a1176
z27270396f6a7acf79d49bac360b2489620b22839d95b03e00fbadcd0497084ddea4c1e77028e85
z3440f9f108fe70290c36914379407e3858b37aed0c23bb980c85e58df555730b9ecc2c2835a97f
z14cccff9b02c8124709c5d5d5c85136a43818b627229f5efefb8f15eef5b4be83ed9b8e6abf3b5
z90fd80e5a459413f8f14d45d9503ed1699e8e5e829561da2d09f0968ce9d2fa79f858e3281cb63
z2f1e66be6ae644ddc8ae314471240d5a5ff787227e4e1f92515d73aef760c595935c175b1e2f0a
zfa5149ed11716089b834f3d0e59db46ce93c5ace6dc39cc5f135dd53513623f505dd668277c729
zbef14811c086dea35cf06e2a016dc14b8795329d92486892f959208fba7cd2d9b17a25975dc4d7
zc0f72322ebddd13ee58a22ee1843c60cc47cc664979ccc655f43717ac1064e755ec99766243084
z72ad45c77f79e0a2c6bc5dff36f853e31f7c8b4dbbe2b4780715317c9cc3e5bafe638689e08dcf
zc4db9a909df07f53a3da99f78bf0be0ff74e71eb1481b22fdb1fe7cc0a67efc3ef3c5d33c8bc1f
z10fe514a5554b79c387c69d3f7384a39ce99497cb39746877e211b859c08e7e58732a3e9fd2850
z216d764bac6dc46600c276e43fb57dedca02da0217469e7cd7161170454d939287033f227dbbc5
z9483d239bd7e3009d739cb295c4d2e9d04fdb9a96eed0174dcf3797cd67684db10c96474a3c07f
zf5de6ba06ed42f3bd33913f0dd225a282ddc29044761144a2d3e3f37e5bb9967500a4702682346
z9da5be61dcb14caf70f3a1dff0182b09748a59719557f2ede4942bb4058b0050559e3902a394c3
za8c4164b215856ea56cbd1db9762964c230ebb5e4477b71ed400a526a86419bdd0e2d3e05744a6
z7c2322ffc4a80c287f60e1e990c41fb9af77fdd8ec19cb17cae9a1821039dcf378a06c932fde1e
z2bb2527151d9d752aa645992ab4f2bcd38c0c8777a43563b0a65fd4d2fccbff15f7d3f98ad4f5b
z09e1e4376b67404904839702ef049ec66a9350207657f7df23932198d9b05e927de308143df487
z9998163c1907a2036c24879b08b7b8eea27d1f02c81cf558f7f4a5b4fd3735b1ef66e1c56028ef
zb78d8e5efa2fdbbaacb17ed33667e257160b6ac7d61cd70cd57f5ad090844612b391a4cc6edb1b
zc191989f9c15f5cc3abb6e4829672335dc71f084f8298de029fcf4d97c8b15e91afbdba0989353
z730159f84188a036990bb2ae3a5ba2c716ca108f791af7c696aa634381c16bdffceab2ea8d5f61
z4b2692501a243849f62f2cf627e31368cb6efc95fa9eb2960b88b3ab267974bb12b2ba8720c194
z69b1bdde00c6e911bb186f261300d89b680eeb5bd55d583a9d14da9080ac08eab0a960525e056c
zf1b5089e70973b8b18df1c764b719338020a058a27ffeb4bef81e225105b34402b36cb2630d9f1
z7a2e9be1c1fad45e154c80137744079719320966914272a256e08cd805cb1f01faa474591c7c45
z4b1ad40e887b8a5241727e1b0f9e03e035befdb8755fa3e669792b40d633915113045e5731df39
zca2b767e168f05c9212e8e86fb3a9655c351c9fb2fc6edc22773bf75c64bf117b73683da7bd8d6
zbf62965aad0d68b3a7f60d698676f89f3d6c3f0382a500f081a9d2c084b79cbfd8a660d808dbb6
zf45e05df7a421d4b2a081ffd14a4f00ff2f42ada1cb4495c9b59899d5f56b78d79f49c8dd4563a
zfe87deb202a92e047befcd959712e200efe2729c2d6389ca0e8c2d1dade287245d6bdfdf311c74
z557c6a14791c7601c1b14a236f72b4a5d89b1f5b5b702076aa8e77920ae093b4f8b421d0299403
z7130d671cfc6b943ca1816149975ad4558fbf217ee90464f14c321abcf537a8420c46e5c7da0f2
z4765a1dbd05ecbe0b9d36fac1c03a795de9ef26112fca13c46f9b7179c24076bf1085a58986832
z38d9a2164c6d5e9de5b0aeea97490a2b4a8c4aacb87a562fe1ffc8e105a7120f18ab860e0b6dc6
z5460056d07c6d1284bacbe2554efb3033bec12a713570bab44d858d5be3cdc9013ea4c33967cd8
zbc2f6e6206c014488667c3d76d849e09a1d6fcd38894a882ac08de2acccf50b5ca997d90b63ec6
z5cdf57a1436f09e5ee6aac8c751d778119ffb10b39fbd55935c949c4dc35f0cec44da79633d0d1
z338e3dc8a5cb86568a20bde81975bfe53b8ad9bfce37b0e52a70fc9b87499f22eb4fa64804337e
z8975d8462e10186bd18b1f34f1fdb8c683b33a5a0f48741e21a907c121bad47c3460831cc01a6a
z99ec0965f84e449c2fe87d1e8a49384deb8280310c09d50fb77ba75197d728523f095d69d704c4
zd14abb2f47b1f3a1ff0a70d80e44e57298105c1926c1bdb3c0895753d969d2096506949e32faaf
z85a457a0ec3670b01f65ec1e1a8b3bd5bee01434ee230a7d88f17f3f6fa9fdbaac5b48baff1aa0
zd90292176cca5e11d47aab05c26f6cf1efb10b01a47c86f4bdb52c5c4ef1675441fe486ec3df01
z02988fc0ece96e36d250f063d6d38b86e63f37ad214d256d250cec4063ea6c5250cac06b8b3940
z173068063a3c2bac5d433c981ec1d09656cb06ac2dd294dffb72ab7e41d9a8c89c64020cd146c1
zeee4af22232ba9eb0b6f893acce01e0003c081edf5ba54b9373dcae128a3e6d742ebe130e339a1
z38598c443b7cf1743742a6e4f5408d1cd657ceb898e1e93a3dd79364efd3676927288f03c626d3
ze0917d3f7230c0781396fc344f27934522087a22562f4ba819d82f5347e2750c45dcef2ed25cf6
z688b6d370fbcd01088fb775afb5c877cd805f633e4d1c15bca7744fddef593cec59ec3ef4df8e2
zc360d45966671ee465a86ba8fe04563d0d3956feffa47ba0be38d29b2ea1b4deaacccc1a1f213d
zd1d26bf86d6eb4d8a89653fe64ab475c5efd1b986d2546b8cd04e6364eda38ff77eb0daaa519ac
z92be925daeccd5f4a8f8ccc8c569b62f5d99712257b3a17d3993edb570f387b0b7792285a02e84
za3ac4146999f40225ed86c74c3176c3847d077cd82754377c9c2b5072782653257fa2f29861ed2
z898cefccceeaa555b418680884ecb723d810054d81dcb9db51a6ff1524eb73d27feb5d8027525d
zc38d3dda40bdb13f61a23cd3b4d9b76f78dfc88cd9deae9aad88a2bc538c1b844a1d821c566a69
zf10396e0159a38527f7520f0d0d69844d0eb3ed991e90fd3c61810011a58f40da9a87e5fd0840c
zc607080c148fb41b4a6706c7f9780a7aa585c5e9ac7a6c770dbad7b2c65366ca3e4447f630f287
z54818fdfcd76aa550b4cc4f3f5b444d1f55b22026091cf48e95f9389258ac92b4abd0dc0619fc5
z112c0432565edb9ae83629c0e2b05543bc36f0fe8dbbbe6edfa3eb4d9ee46d3632358099b1f08d
zdba307d7df28db2918356d2e7c1b62df02fe2df8868b9c59bc127b717d184c0e8b9cffbd584da6
z245bd45acb03b505975e2c942d1fd3716a800d0ce1ec9da74b255e951522ba26663da7c63ccac5
zfc09f7880155b27a1fb8a0c110a4a55e27725fe26bf4d57284ea6be4a3b5f2867b1be25b19cd49
zd27a1c33db8439632c85018a79aa4eeb1d3f3b5e1f6878843489329b7f96866f2b889cd5471bb2
z61c679465d25dc22f0f8afde8337660d14dd1afbe0dec4074551171e060159ef37c2957a7792b0
z234bec4224b3b36a2488c5736f90c2dbd3f7f6034ccd7dc0b44b43abb3ab7ee16e0e95db823ebb
zaf02fc0c078f874213cfdef44d345298971580c7dd07ad3e9010e105ec4b2624cbe82f26a53885
zf2a46dad97054ef3d534ab0b0768d6912f303fae7d211ff34c2c4efcec6d7eb8ac41f8605ded1b
z7952d02cf875681119ba9e4c6311f0986358727d4b099a516a26db34a0d221378c16c9693b3427
z3a671f9af2202ac398e8871908291b3e7f407342743f8dc24c8302d6e183f41980943eb96ebb31
z16704f2a5e50a0e743d2a1e16dc42b911ac411f15b4025aa16957c87106e62d5c2e7574d834e1d
z940b0ab7075be57261d7765e627c3c1e76352a2e24d06cc9998627b93beeb91aeeccf404e5359f
zeb68df15664bd8f9de76ea1ccd833a8984e0fc62284d90cf4354a6c3d5859fcbf0fd96d97b4206
z711bda5d824e984e2a0f6447a018b6ccc24acb456de82c5fec6a709f808e079990510f590a8ad9
z8057a2cd42dbcfc8d2fc0dd282bc217716f3fce0b9481485e2afa39845cc479d6e6f9b821d7859
z3dc704564a4290876bafb8acd4766a30a65dc7f421ca3cc8c00aca489204eedfbfcae17e0e321c
z2659c5b5a6b6ff48d619a027dbc0af33a1c9ba404141d34e0fe1742344d1bb7d9beaf17b64473b
z83187687c50e24c3e6c6643da485115a9a4c89f2431a07fa9e702a29a9acbda93f5e2504ffa145
z1048e8b16f96bf0a6b8b9b0dec2726a122a027d1978a02852e40f9926abb35a1b6b5e82d8eeccc
ze8b29cff34d9965d3698c22b5a14319fe6a7721eed02c10eb68ae6f839d027bbb00169bbddbd2e
z54eb90aa0e3f24660efdf53eeba49d9b8cefaaf5c10759533810a9bd8d2a991dd6b159d6aae5d7
zee38fb7f43ac75b889bb4426bfa80f2fa48548644180cef7eb0a10a95365b3207e65f7a20db638
z7d3e2eaad3b3e29a668ebc332453a1a7a7eaf01e360d9dbc13ef401d771941959e1e552aba2e3f
zfb773c4615fbad2429cc2246d073676887a08f46e893ea6b4a9c54f378fac014e297cc3a2bf7f3
zce1d5aac739289d73bcf6dddce5e9dd7c9e31cfd5d8a44bf1ed5f015dc1d9c242d92b4f9a6dbd7
z2f821e3f975241279dc1f72eeacc8e2f7283e7467c6205fb62beaa4cad28d46f7d5317a393cc17
z7fcd3866a776e0e381c896cf7513aa3617e2f8dfc76bfbc663d90b948fded40e5f628ee3e9304e
ze87e6fedd2e570ee58dddf339af46d21f65ae70423b38182dcfdd2b9bab65e37fe92f07ec1ce45
z1a64838ab3352a11756f24bf7b8919883403d5755438f212ae9e46e64774cfa34487f3804835ad
zdb6ccd64c17f68f1a61e01b2e58e0d1072ed21b6b71b8bf57b794c56d42e70319a13078027b719
z1d876d25a4e8d9a883a6b0acecbc46eda3926f87286caa416e99ca495fb4f934976be17b723849
z0f092aef4ce76e43d5a2199d2859a3d503aa4f533ad13ffd97cb8320531df6de2a4c5a94246849
z39505e0d8616c9870692656a3ae9549d27ac9fa6dcedd8ad5268b25d4f63d5f94155c7840f2d65
z7ff40449a60ddb1a2fc74e33086edd1967a833049abad398bf7103ed62fc1751165370b7102d0e
z09c2cf85d26fd9d8bec50a33f8058b86419cea8293b7b8c8a5b1a3fd61305e1c93388efcc23d54
z83182f3456315dd4d3b7996e1beba8c9b25802b13a42dc7b09c71260df2e7104f5010512d05c82
zf470ee4a042917a77eb2ecadbe77db3ee8d5d17ef70dd0964c9520c6e8a698ca9df6102bfe614d
z4766b6ef671bf5439415da116288ad3207a0bf5015e6ab44ca652d23b5919bd83ddd8af02fc191
z3501552593ead92d613298e635d5ffaacc87f976fc28568a9a1ef6666f1d0bad86c1ebbc3d76fc
z9d6fc3293f97bfb540d5cdaeec1f6dc1c854377ec9eaf00f9bdd1e2d352db8a3406cc6ff423ff8
zd67545de8949affe4620e0feffe9d553d86a9bbce045accdcb8b4015f6dbc1baa138855037c6ee
z36718a4f39515f0f63d77b7c9bc6f18debefff276125c0506eb26dc7cbad90f49df61967b73290
zf9db84b464235f8d33b448c389949329bf907cb9cff5646abc2364451b2e13ed913d768d8175e7
z7a6adf55629bcd41546b5b65f55dbb5c56da9e1714173c654e11b3517c11634f32011563eb7450
z08498f3ae860fae2c2dea37641118d9e832c3bcef352713c160990908acbb9f427b890451984c7
z48f3d0b86dc256f36f17cc513ec7e41d6e2a48e15f97409eecd6ff60b9b79680c8070b8885577c
z02e4c5848cc1311dbf744e287502a4500d586e91415933487ebada7c0e5ddd4364e538e532b88f
z04a9497329ba04f05191ce8af2bc6dd0b6b63d99facf4e246884ebf182c4ebe13b798df9d9f595
z0eb70b2e6f824a34b36b3afc4cfc856351b3f469cfd0e13fdf0244a5257c125d0c25c2c523a20f
zfeec033b666e00904575e3bf0cc0c357b10b8061e7b110762456235115f971a5d16eabb3209834
ze39faf3950a410ac07fb060ac030571a44e4ba566787159c0ee8cc07399a2491afa55822585a5d
z3549bc5c731708d73fc8dd31484a5b468af74ccc7496c9907fdd8683e4b9757fbb067946037830
z5fcff1aed7c4be8e76917fff3f99251211923e4a0382b0db025166d1515bf9e8a356eb5688ca39
z591fb5d6c35fcb979566de99d43122c9b3d492ef3282940d26946ab1181f5f43dca3b34536da32
zc1a2b2ef2756bad3ae25e3a514083f11347b46a6b02f4c25d4767808236a255b50778dcac9b64e
z6299c567165cfc4188a7aad29a9ee73fa29d6311c9aca1463d2c273f88a9e022ee3370d30ac108
ze276f7e1de7315df758bad4f87648d4d2284cd66fc89d41653f067768cf4aace347af417f9cbd5
z53e7e0446e0945e7d7b954c885a67cd962f0d37d200f92cc0cd56e2b985a9c8529a88e490c3e5a
zaf26c58286b08a701d1a6999b41fafab88b309b2dda68cef0b803776f8dd4a9f21c4c71c884e57
za8c4070e46a81d76e4d14af60a38dd8c2b55cc2d12638e581c5485ddea31631bf9bec4a0dd4f7a
z351fe43ab46b24da29d3a4c649879e60a23486655402e23cff45868cfbee42a926c50013bb75e3
ze17deb0eddf96225030a30f6c9c6ceb849bc60869ebda9b03ef805bbe432e5551ec5dd3c67e3f9
z0a37d81c2dc065278a4c88b0bf2da542269e8f46161c64e5013e124ec6ee7f50790641c2e809d2
z19dc1d3dac3d4432a8b0b19ac69eb243a988612f58caf331e45ab02ec28d95df83bd2176cb8e32
z5dd486b5b5534d9f88d4f6ecd6614a591b35cfe5e879dc26f6e2a22c8959a256badfde4025e82f
zd0413c3d4f094d92e968a3291426bbbffda8ceb80b420dd2e913addf0e73a2864bcfd9c0f51544
zbb24c453b9b1ffcbcc30755831062409544fd64b741048a76ced1f538ae80b66f17895299bc545
ze4ec529ee99d31bd8912e33fb653801e2d2a4e46b0592bcfb1db686623e279742ac07d40b26aae
z6b5a30a0eb72aac43f93cd3579c26de81be6c6b28966d7abce3f8a5381cd187e722e1b818071e5
z3cf30639a950c0d75975362891b687a58b0774c34879311d0969acbbdc831053dce18adb8a4b13
zf24efae0881af7d8d1decf44136867e255cf5b3d808c73d7f0612de417bc685011d8e9d31e064b
z9350ff27a82e6ba9483a51612cff81c7772967986f67888d7398f0f73c3c0d2dbec33d85c0f1ed
z352eb1566e73e59f83ec0d135699b8b9210a36ab91aa5482b18d5c98066f3078038968575fd12e
z88ee03bacb8a383c4b8088838f001df2ba89018dab1e38aeb17800101297fa6b84994efac00b6f
za6e592c462f3e00a8039238d552e494e477b612f866f2602b9df142a8d069bff3c6edda2e45337
z71374a201cb319f3e9961c2dc982d79bdc49aef43691cc7c56fde611cf68ff221647b2f6729d81
zb920fbd79f16d64e24f959bf7e1698f3cf8c27de0b53c89467ab116063aa9ffc479e920e9d4f18
z9e8bc86fed61a9c88a2320e7365f2c499bcede3d8dd10b2b1701726564cd14e8bd2746533cf24c
z123c21cfd078d5e827ce7414d263b88557d898eaacd332ab007edb8b13eaa24f20a9828babb5e3
z7177170bcf3ca040b0cba64b4795f014625fdc3900c559880ab257f1a97ce421c45fe6e6c0e25c
z4ea9c40294aa5a6beff0ae2e0b7b416b0be94c73a86deba9558275a0daa31b6e61f0b91c091012
z716c6f53377f1ba5f11df19cdb39e1d1376eb23ea257f2d565a6f0155e0ec21f8635d6005e41b7
zea9b8238b1c1672277b593490f30e3e947fbb87b04d8be707aeabe6b3c261565a01dbf0374d15b
z992225463611c763a081b8ef882c567954e347b37e1f2a5807cd7af7055e0f816044d9c554748e
z98b553d18adc5bef432491f213c38ed35ff8709a717646f3d8c83accb4e9b04048f233877a4ca0
z4c83449603b041fda06da699e2ec37e65eeafaaa2d056ffcb6f852529767c11b2319cfb4f84a5f
z2bf1627782522f902f676731956f3a24f6c3a2724a591b980a8fabc16ee67eb81b375fd794e8c0
z5e288c0bc9a71c6451b98c8094e16ca3482dcbbb7e80008959ed0d8ff9e75f1c1ecd4240af4261
z58eb3f672435b345bf16cf2ad375cba4316b8af2382c39bebbae2a4de1325084e797fc6fd6d9b6
z630abc714c61c5d44db127806b3f3dd56ac45f96ce835a7dd4f057204297e1d84ac2e6de06f9ee
z7083764b4aaacc2f817a09baed3aaf6113c054f388be90cb0ec52554261a68674265653d136e2d
z05b493f7efb30bb7bc490bf95d357d9e58a318f346f338e499fd8565931127d8f3f6aae7fa7792
z0d0e6a5be262a360db84c13d0062ce1880a5308d86f87a596965d3d20a5489d79455e8d74622bb
zd20cba99007c856c6aec50f27af7e435927cb141012c25b8f246aef6294efd610a2c918809b833
zf50164a2f8981f4bfb3c3330b1d8415c4c6e00af8c1018ce3253f808f1d97649eed1895331dedf
z8278eb926b74599ea78a23ea823911dfe4860d2f8a435ee467873c62e61bb9bd30aa5db58e24ca
zb88fbaf26be686690f245bf7970daec5e17d00a7ff762edd4fcb93d14ced479c50b3566e489216
zfd74282971d9767ead0502f2ab0187f028be53e6d4cebf6a1da01037d57ec71f2648835a3c70ff
z7892cbf0edd9a2e43c403db35289d36b607009a4b100b537205a7b6e503412981c15f88017ed19
zbe90d89efecf58ba8ccebc615432aae858d12352429ee01f67654feb8ec8ad2427a9896ba41157
z3f07e3582b942babda08e42b4b2fb12514a1d3796057019aef61851cda763385faba97029d63ab
z19ad02f9b14601ac6c47486f9ab576633616d3426ba852ab523207b50baf783958b78fe0147880
za29c624f7de1346d808ddade9d448268c832440b7c42bf9f44898d2cf24fb1f6b56830f0773e4c
z29c5ed0917f57cbe6ff491ab0e36e83c537487d7bbd689e7bdb39661ef65862633686d8d405433
z7ba6d459b2c7dc2837d0ad7b3c36cdd0eee51ef44078219674f097862220b4402a5922e05d5efc
z3cc930632132bbe2468e7d53e2aee46675db28fd11420483855402f8635f9a90be162f93b9bd51
z43ced83a12db5e41187823d979d72d68a7ab1fbd9713ba5533b15a0d329ed5c1b17ec4e9bce61e
za7564c66c3f1849c11bab7c81826ae7ece89146034cf2b4425c576f8a62c7965aa1df040732eeb
z92c273a29a3b1e22a51bb275023f085b628c66e13195a1d2772551c1910008898f73d2e715c486
z8c6be88d7f28117fc18d5156d4964351da899704bb41eb7611021502c7c31629f76d02a6501a41
zba27f212e673e5f0b35664bdaf0bfcc0551e41032ae706bc92afcc208eea0b2460e7382913c74a
z96a0088c9d0d65f915d1956851997956b7da272558456c9e5cd0c6477eea8120febb0c8503bf5c
z98c8a1bcf5a72179ad2ac4bd7216ca531e7dd7d66d7bec4bdda57f57fbac5c347762144d2fa580
z511c95a50565ea39b9b62f08b12219d9ce70e66340547d7d3e810456b51e6b6a36b3514cb11a62
zdffbb757f121660d8710d1bc215c9733f9eaa1ab7fe2046666a77debaaba0fa202c11922248979
z57ea577f173680da6d959b4cf96166162b1e7b0f001caac1b292f863218e4aa7d7291028e2efb8
zbfb03d907390715a39f8f5dfc45b8ea508f53f9f9545a24e21cb694ef74fd4c38c647ccac62d77
z7a94d94f45476a7b5e34706c5f1511048c1a0406107b1941739a37aa6de9dd0b43a9e4e3da7916
zab3bf473549e9519516686442f08090c85e943870c3a3583aef624eda88f48f3abc52eefb712ee
ze0eac0f4ae7a366443b1c211437a5b17b1b7f7edd670da27e6676872d7238fa0999bdff7c5ed40
zfc1397e7a6f3cbd5adc1a4de42a36039e1441c4af3f9a214ea253321af890f559743c105258b2e
zc4b8c64e27bba3d321d24007ce5397c4ad81bf4a3c632debe7a597c77cba649dd7de8d9c7d5719
z5d0ccc90814b8c1fa091468f4461f59394c1ee9a483f9582435600bc30157595a1b6e2b02c67a7
zab2f7e7553f7ca7e54125c776924b76bbd959d36d7cefeec7d01ea6f218a038c865772e9f02118
z245f37490056b11a37aed7a4436d220a7aa371f7dab7889774a71d159749f31932c4d72726be5c
z4ff83eb5bcb7a1118179b1b384ee34400dbefa804e2e3540069cde6e28f5c1be47c420296e28c9
zeb58028fc791b06e2fbb741213559938ce14f8a2fa3ad249a6099417ca5341b37d77bc9e1567f9
z80834d07a6031bed63bf0913e9ff366e5e54a7631599b54308d3177b7518cff29f1ca0ed92072d
z62f33bf697077e3851d2c64ddb1aa8ba4b22f33a8c0a9358bcde570f68f7bb68d003cd7b125481
zce37b92b360d05586dcacc7f4a61f39fda60707fa9111a58acd19acf9aefea00a9f48b7f2fcc1a
zd4d16e69a2166c77e2369fdc437adfdbb0f6453a2061efbc82f16ea21769ff9d8238d6db917556
zc22a103b6dca9e807d1876cb4c2d519b876763f7e86758520bde12e2f2a62a7159db3f09a141e3
zcb7d757681555d438d1a2e45ee985dfc7278e8ef1ceaff0417562a64958e4377ec3fb77bbd0549
z0fcd2ff40de0a4d2e88e4e5ac4a303cd09d9588d6151b42386076ab3d008c2cb90fb0b8724a9b2
z54fd5871da6b240354e0f8ee58fb4eae5a436375138c51e71fd640b5ac662c42615cde8b79d245
zcdfb19df75c3e723a0a6719f4aaab56fa148cddb88d4b83e0c1b77f796ca81a05ea0e8e3060d2f
z3ab7d189507a81cb8b3da00ca559d5dc73d064cd358861313eabbcfc2b3bbd7663e442856b51aa
zee3967dbdd1eb296ebf9f3998ef010610d1ead7e3d27b2535f3d5ba50db4fb709d7929d2317be5
ze69599a8b9982e6ea2aa10964f0ab3e5721b850d539745ce48f164016e3fb4883da0d21e469e4b
z33161d99caa7d2ec128532823bc6bb0f3a0dd79a0d51c5df7ced121b24d9300b52ed9bd0a1fa7f
zb8368a13f616522d8c6fd98e090996d1fa9cf70dfe431f48b7a69388ca0767eddbc096257f40e8
z8400d9e36f6b1075410b1118a3b6ffb2ff4dcd82eadc5edc4eeda6ef7d3a8040c9918fb15e15ad
z0d65c0e36c7542a30e19fe8570ffc7fcd90d09905ab24e786cb9678979bdc38ed23400b70bc135
zb5712afe2e848165d2072c95fe34267a0a9d4074f5faa665e8642d794619a87d71751bda5a4f6c
z8cf6e22504762a9243e17133f6ffcf2a4825f7556084071d566bbd872280b39c2d92e827c7989e
z30a48f4a6f0378cf4a23c4c434c1c9e4f97e36427053dc65aa491b15aa3f6c4b2113192392ba9f
z9bd71da49b5b73e913ca9c3cba85eace1c06eb83efb4cda802ae4c52399d12989fde72091549ff
zac56791fd96e4a4692f5aab9a58cac7e632f5efed7ae91efb8bda0b38523652d9c20402356ecf7
z498a3da9266a532aa69c58a61afd24dfc6d59599022d56593a71b471acb094778f85bfec2beb8a
z9e07b52223f8ae1840cd9d406a3ac70892f1e635d2160dd5baa57138479d6db6a54d3919a8bf91
z10f681124128434f6bbd31fae4479a3528f5632e8705eff13948aca780e16d2e4ae5cc54b22435
z87e60f4f2bf1a1760b4edf22d0d12b3010db7a81549ad13031c5eb2cf1ee82f9edc269a5f07356
z52abdd7d473509df680893d483dccb8ab5e39fd428f6c2135dc1ef527c21d6da09306913ac6d45
ze9421099fb16dc5d27077b64b6a91fbec310a91d537b4cd0e292cc0c22bd2b98111f87baea1906
zfec53a5f149ad01355c24ac50a38901d4471565c093113488aca965c4d0aa27e14cafed6efd979
z4c5f62e2f2d09fb6cf32019be8ba0fccef0ad43364130d88c2420614ecc2991919d0c5a30cc901
z3046814fe5638bf765b258cd6e394c7d4b072572a9ec3cf723fe1776f665e20bab0a0f079b36e8
zd68f3e88bf63a0a3cffdec0bea35f6a013cfd83f4bb0afd39dba9b61f69ab99aca7df52cb70fef
z6a4350341ce4de5b2a5c4a4920e378f4e58dfdc9abd6d74de728c5e7d3be1f7c8068a8e10da50d
zc7631617bd822f3077dad53489c583414b78ca7af64f320f429ff222b8cc32720287e9959273ed
z555bd55b44d9f44bcbe17ec9ea5dd17f2bb7d44ace4760e30da5da105c20e3a814e003d8c7b789
z0879c5dbd6ae9e1050774ae5459b11909b6e1260ed5828e7c07dc91c1f07ad84f046f271d45359
zc516e7494f3f0e8319e38a4fbeb833d83ea962652857f6b4db32c0faa4e5131c6368df4189daa3
z1994221d1c0194bd9cdf94227e77581573096e912bbd896861c9a071ff9774c28bad20ac75578e
z9f168801d53cbbd3707182e78175cabbbc9a97feb9723e022766b56cc80578ec8b10deac6744fe
zc7ba5f378df8f53c484463e18a68df970e87d416924fff7f8f9c9d1c0a1ad49b03a18639c60f66
zb615a9f92e1ad2172f9704dd38d78e7eb5a94c45a3a0f4d0ac4ed139d61c3f9a5e06679ff00993
zcccad438c6a9be33673da8d814f2cc8d88ef1e618e2637c9ca81d1f94683f9b469e2e9047b2891
zcc0947d5a02a5ec09a50c5f267a0ab90c9669e700b8a420acaebd8537deeb0d9c65634d7c4082b
z0d9b5573b019c9ca3778e61eddc0c742e0e90e4cd670739f1f1134993f7b251aad7538c5f2b925
z7173f5fe5b8720459610d4052b6f0e857035e1bfdbbfd4c3f2e405dbbc6a81e6f392ad59db24fe
zfd175fca6d5b22b3c58666e66cd8a65e16b0e6fa084684266462e69862255392beb1445ec672cc
z1d43a7e5cd42cda66adea28c5c95ac1bf6f74d998afd4565e30b6f01f2f48e8f1e30617d6fc28f
z932a1c3735d19300afe158748f170ad70cc107d90be68b4dafd048c9e7a7d4b4d04679e4eb35c9
z97d4e16d0d1ef1e4af8c7135f06216f2e7e38ce966c04582e5b61a8d3ba6afa7549fa33bc25b30
z9102e5cd303568d430a5ef7e13b06f54cb1deb9941fa278397cf238c76d5debc85a47ef41cfbcd
z0c97c235925488d37b85c5ab491f8489358fe0f78128d113591002ea567e21d892b6122ee964ee
z139a6fb1f9397a79cd4192e4806e1c5085affcadc4fcca1d16dd696d7283ea823b8a4176188c47
z217b583a10f91496c3ef0564f33226ba21c31530285b4a937a8b35c55fefc1035ed5227b875df7
zcdc81947ddd4451af3e05a18df4ef54bcacfb7934efc35246d6b4a357308ea134bf0e3c6aa88e4
z0d27288e9735abe31b7b46950e9e333355764c89a70161ba7a9c1a965e20a46e075b8aaba2efd0
zdba21bd6d5ce95e46e75c669603b5cf6c1d611d5e46673212f11f53e9ac39f4ded0720f9272d67
z8cc3c3a2a339c2105c4e92a866d42d44062ae73f519a3ddc1f48f611c1f6cc96b1fb6600dd21ce
z9b4dec0ed10809938b04a2ec0c161a71267ab390562ffc8267c8c96a2156890b3040084333a50b
z49348d9ebb59df963ef8c33de284ef17735638fa8181265ea6ef3ad85fbfdddaa880abbaaafe36
z2bd4e806bb563cfadcd51bd1f8bce8f58800aff6c9909f5562c8a09ce7d54e403bed18282f0b8e
z2a6ac5181fdb8bb4f802847b7c6827a38aac32487c27759db89a698744cdef1aab4fcc99acfc6f
zb65f07025c74b8acaa864d7c4d61d5a84b2903104d15440ce93d423efddc993c5d8169e925b199
z94bc72e27718e19dcac035563e03f4365480cc82beb8db21d42eb0a08f058cddcf3d656f014707
zcc9d4eadffeee4be2126a837431e28dbb173fe66d26d36929d601a2be1bb00efc7016a31d840cb
zb74224862c38178eea6497a7d1649e8725964e696e5851a13f3e53f6cedd0ea6a2caf9a78e1ed9
z0cbf733ed27f3bb1c880921b093f1f4e02af044649c26130ecc7a6174c27b418c6a9dd64cb327e
zb400b32730ef57d4b026ebea24340aebc4669b1552f8c2869fc82110e1ca53ecc3d7d65ce44d87
z6e7c0b225072f1bc077900ee1dd2aa888e3289947e74479d4bf8ca5b98a815afbfad88c041389f
z16cca8fa976471215613ee3fdd5eb7da558d66621326b6d6edfd134b60d9918a3ff227310070f1
z9b2000ffbfbfddb6da113e68b3b11f64b7c867725c297b579d3b79fa7407a827952a2748a7285d
zd1b0904fafb1b6b238b96819627adf6efeb4d256a3dcf66f21496b491cfe4f0b35a23feae44a95
z034bb4ca8fb60ab01500b1adce3ea9f765e019f0086bea5dc72d940b2aa153afb245db15ff1796
z3348da76b4b8314073e39296500bf5261282671acaff50271c5db6980a2e80b9cb3b877b104acd
z5cd359754a4a3862a1fbcafdc0b6cfea896ead81aa489482e9ecf28a68c1177417daf1ec0ba64c
ze89c4c2261f1fc17c12f0efb7a069905cb65f6404e979f0faf3b98188a7d6a907a9ba62b1f86f7
z93ff8286a857c6b000f32d78c349f7bfa63ba4b9f14fa280b94ab154ea36510d99478170c839b4
z55844066a8a955f874a3f7032cba2612a0616d7f2a24b1cca7afbe32cd66601bbc07329cf4e106
z0d34f0b8f3ee7ac585c2f587b23719d8e7a07e0005427789e1ef1c8744e20e33d6123ae90c7a9b
z552687f158d6824f5d0fb87e2c457ee0d011edbabe71a4715ed015f1fb237b1f994b0762e6d5a5
za3d0d1a7a0b6618e8f83bc72de05f9f14857a3f66a3a573a8be477d6e4b1a1d035ad9ce8e96753
zc4fa0fd9f6a4cb11047dc7237dbb1ca1177796da73fb1e55f4290c09f7171b708304baf0f434f1
z068f38847b98ed218704a836c4728da389dba58c7878b59683c704802e02f6d34a14f5556401d6
z110b1f75a2204e4e7592b3dacf8adb356abe52b82621e4e6490b2d096f90e54b30688ec088ef0b
z88f26321325935356c4e1c148d06e8361b7811a5eb692a534cbea1b423eb145672bf853e4996f8
z418f7fabc8664dedadc5fcf523bd791c0e25db5b2598388530525bc731c17c09eb87464e2233e0
z004c71b6bedd18bf79e208035a6106b8d4f18fafbaf4ef6d405d1b55f92717ee71c2748e892668
z13ddfd74aa0b011f0048209320eba65630c029976b692d4149ccfa0c27ab18d024f3820ba11152
z89eff2dd677095eaadd5526dff91bb3eea4ae99bb7b76968c5f3c44b0a0cd8c3688c2c8468d100
z457b9c15ac9981000e8688611801ab1bc4bff3167fd329973801b69c99f5584bc589615c285b3f
z6e2804d19cc10a522fa1a884057c46590c2894d388f0c342c60da925a7757c38f7f1ea0d558f83
z9d7240f71a38194c4db211e3d423f34150271a14ffb12c0eea43bafe7e1087a327e39200d2bf9c
z360e997890d21f86154b028b98a5a4171a028c8ac143bbe7c3815a9ad5daf7cf27f511c549cad9
z8052fc1a43d16a343e5580c5f12d49f32f84b7ab441fa0fd7d80180173ef7d9a6a5ae5b81c357b
z9a15b64264817bc7e28ea8138f5b14a40eaa3fd74ca751d430ac6568fea5ccdd1cf952d1d5f4a6
z1b44ef36428f80d1d6c13bea6ef6edfb6cfd994f802e45bac134bcf3379d3e4dbc2d385622099c
z9ccc956ef95f06f1c8f0ca25be4b9e6fc7d021d2fda2f59a9d82d669c0ed1979ea4c243d612573
zf7a52d6728c05f37fef98966d5a73318e1fe2cddb512076a6a87be5770aed4d9590de3531b8991
z961ca1fff6674a45e0367dc19b230fe5f65a22eadfd32d2adcea7e2aca01cb50e4f3931393172c
z27cc6bc9f157f50c2500046663574310c3d1a967229f5821f598d4e3910ec43581b10a207ca2a2
ze5d86c2bd2a2c0fc95a4d8432478b8df43ee2d3d381270ff4d51fd5fa4cd7bb015f2d9ff17d112
z691d58561905e95a77dcf7333e9bcd9849a1e07e05b55b8e9786c26471961e4feae7da01b8bef5
z92c13aac9103995fc1c8057e56728e13b7ad8e1b073b005efeed09c7a8d66fa300923dc068f1bc
z55749faf1142dffde4fb068b82730f412c972c7a8f9f36217c4cf6b85860b965d243dfc3623c8b
z13ed4b1287d63be98474f4dadbb52f0f47d61c2451708f77a0b6802cfbe7c7221552fa93e0ddab
zcf198644c578977bcd6b3bc04786f40f0b4b9f7c370bd00be174a9647674ba1a9b00eb328860b2
z582434c3130d19702af1f1399a32782c1bdc6683df9c3a56c85d2f11b8ef711a6932674b21ccf8
z42f471682e425c59f0b6ef4abe0549dc4f50e67f1ae7401b520da76e85b3733da45a7a29ff4768
z61e62ea7333e30ce8c8c5c503a477fa225cb19c31ae2e6e3f9031f0b6da12060ddb24abb663be7
z87a0351414a9973d5a172209ef5b23b852071f832fe2c83ecddda8b95e6639b2173629c5116e88
z0684cd206b6fab3dbc10ac63f3e3455f230d60e18b70171d19ed6da5c71d2f4a0f1069c12f9b4e
z19a0a393a2641113546961c1e14e12013aa98bcd65ae9d957004166567ad25ef201ac8b81e7004
z101834c3b5d044b0595c9253dfdd7fd26a9b271beaf954cc8b2d106b738b0f5c95260515d31610
z6dbbaa3f194867591193f62f2d672d1922d5843a695d8ad2f78ed675e4dd3557bd46fdf9826619
zb67888c6c15376f22d896bc4a2609410d2bab78aa74bf463b70d56996efbe66d537a53a1e1d06c
z2e8d9dd5fc2ef57222ce0ec1207f441f8a2dd507b1e31ebf499336451b84a4f95971751d69f81e
z44766511ec47303407444ecd5f4fe0b7c68d738617e70c711c9251bd387c1b4ea5bfaf1d71e5e2
z66b925f8a4f52bfeca7d4928ac2da29f5b141943b1146fd56a102ab1102226448334679fd801be
z97c58ed7174c69c4b4b13efba4d694d782f890a39f896d31c989baf95a4376a452f57d7745ba75
zf38a46ede3af2c258917a051eb0af3d9ad40437fd414f33d6ad18d9224e1d1c4f4ea3d73c1a964
z378dca84efb25a678171287ea321f92004a4eda0291b6a0bc61c562d541785c76ef3ad5892ea2a
zc723073f3a3dbd700bbe0aec30416edea3555495c48f0ed96dcf7cb757165cf93e7384eee3fcb5
za018a1a3676029135ace89f8baed56460a45e6f602397f0beecd679cc501685e8321add15d4874
z06e187a9d47eb2c18e2c36c397722d8cb0810677210ff13f8e2406c351810a867d6a1ddd431df2
z5ce6fa720df7b06567936bc36e0d033f09b2735cd577ba3712f87255fed4559b0701cf1923705b
zc45815e17086b4ffee08d9161c1973bf8af45cad6156d1cfa5c2a1688644e4f155a0b7e2984139
zea28f761e904ded58831ab6347b12da108c9e5b3b1223b694f3b5098fe625f7622834dd6c498f2
za8e240449c4cdfeeca301063a0b472d99fd881c3f519a7f7ae717515eca7f19c2821dd5dc7a9cf
z9759c049625e59e6deca973cd203c81ee40789138a768a20a145812a5e40cd4f46a421d4fceeac
z62902e5a394289564677d17968acc945448a57317014d6737ea4bd731d234753448c43fd346a41
zeb2ca2f0f0952846f5313f381cb0957c0c0871eeeff8e08161023ab2ebbbd5e01ba5fd78154df6
z0abf99b72c6dca7658429218ba57c4b231cb470fc5a44f45aefd6ed5b9a0c9405c8772f615fdcd
z7be5b52a617c5500d9ed74f02559719c20cbc48a9fc8e1069ab9365fe00b478d0a9dcb2ecd780e
z1a473c4a058aa2b70fb457c360c8cbf01fa2f4183a9fa9748b691234862dfd2cb13e25dd6649f5
zf9ccccbf0907d61aa3e4a6ba8b62a1bb5f00e756a47bfa9c09937c0061fb373d55d100d4d53bf7
z46d3811cf2031fa0bbe7e2769650e5d4a0d3a0d73fd71ec46596c4cbd9d71ea1d00d77ffc7bf3a
za670879053e9fc589db41ffa2e61d8a3b5fc6dc58dfc576ca7547051a9695f0fe95267c4bc2fe2
z8cb26710f020e7899f3d4336f403e586f9802efb5f12087de65411ecb3afd4b0c668920c9c7eea
z64bfe5b67ae49a26427cd6353f4b731d3cca6c393831ef7878cf845d4a2fef94c17f97706b327c
zaf6599c0222f3f7a47abd0bf297d49c5bbdcc1e45a19b583ec8fe8ff7d33904101bf35df877348
ze0838ac39468cce35f730d2d532ea370e0296048eda6aab82e6c7e5545e466e69b1f6be9b55ff4
z2ddd657dce2a834c0f8cad0d94a65ac9a0b7810604e186944b8f3c428e176d2327f3a05ab8dc31
zf50c429b7b8adafa7b69710c819ed69bd8a8da1e632a42a86b865287899671ad8a8b8371c48e71
zc1f0e0edf809abfa00225ca9485ded46b4d366606d36c1a8cff5fe3bf80706bc6a7a12adc6f12e
z75da063578b6b85b687198f9ee0a90e3c3f563d32d88bb20988b6ae40237d128cc1a07bb27f0b0
ze1e0f1404b5a9729c2ea4318ba3e735dd8e7750ccb00c66ac0c20545b2d30ad4b59d9cb723bad4
z56fc35ee6b3254b2a348bc83a620a2becda36532935faa4503cf9bb364ad19307b028f8fb5099c
z40918bc516a2a43db352bd2cc410e5a1ec2d7299a74ea61cb69c60eb17f0352f99520a1e62b6df
ze5957ae354be341742ed280c8b7331b8cbb72cd5103e18b4cd9547ba7ad9bf68291eb00f0f92fa
z7f5b9c185bc69c684077c83212529e62bcdbde330255bde5835e6edd1b6a93d0a63a3573a7f1ab
z4d5fbae21403d5abc8f5a9f345220a4b7705a8cffb2160bc7c84840a0c2be30b79dadc34561b0e
z7198ebb4a2f5bfa629ea8e5878a09e8907c81b4411ac67b12d0e04909833cb0457dd56ba119c66
zb179c1f6c0f9976d5ec185661e529b423bbc87f0e43974f1dee2126317a896b7b098b3c4fd68ff
zc1e18b63336919f0812182570ab1ff62c422092fc19262215f5f03fee927764ee8ca9de6c87def
ze879f72f309b69df0b06887aa9f84c4e3abc623a8d95ea35d1fe0c8884fb1d23a61e5c2fa5f6e8
z850c7ab2434441919648548bab885dfe243e311d9e638226418cb554e138283f2a1ffe9f7f6a2f
z173bf4b234c1980e49d696f128d26622204031694bc723d2545a829c8bc01ef5259053bf35df7d
zeaa2de1b6ab3dce94ae30c94fd8836f9df1c61b4a4eae961f19791c6045c9db144a7166926e1ba
zdd331c80a80f263970c704db4a960d8c028a8351c7460b94c8b6daea3523e2250667ab3d892087
z2a3ccae1cba5a8efc78efba5c74cd8e9a4101939ae05da12ae3c462f5093833b006a216761d639
z78d77ad20ff91ee76bb7caf88cd104ff0b92f594428d0df48cc6177d3f5359587515926d682353
z5d16ddc8b6d28d71b3d6d9b70a8b1e92256d5213318f0941506af711353addc53c5e8422c414f8
ze78e197618493a82ff922397591fd69d1f29707437036d4c0a14f94c2d0302909edf996fa530c2
za5fb0e78a70bbeec9f6f666622e677d4b4ed96056bfe2009049f6f278f390fdcb8c6954163f8f1
z71975d9297af166290032e4a21792434bece339d1169b95da6e43440cab43a62b31a1ee40792ca
z1d6f35fb858a88fa148d68976b3c4ca9260968deda808b32b94c2906e3a1a5d6a8a5231eb0656a
za2cce6fb833ebd98b9c09ce4b9d8b82bc0b49acf5fbde7084ce63761dd25fde5aa3a0e44562e5e
zcd6f8ce87ac75befdf872e60761b06d94ea3c512e9ced74122358a6af4a7ed2e60b2dfda337851
zb365a58e7df30681636645f4cae2c18c32a663f9ce1a95614e2dab57fed2ba3e1c0fd3d49d54ea
zc1ba55fbb049d8d969e4155c6be8376f153ce5ba19d48e22c57c241fb797a3cc29860bc7e07d62
zce8ebb36aca238588bc659bdfdc3f36c7008a6ec8164bef02f7e05c3bdc5b161ac316c43c275fd
z762356a3b935fa104fda7a618d6e9cf36bd0d0d7aba0fd47ddc4c0f46721f8ccf094592e74566c
zadbb602c37ed630a290b2bd66c8922c8643321d42e1b7bfdbad0f69407e31a7efdca555f163280
z18e9faefd6d2d848128bd07ea7c6bb60d150eb4e05c2bbb92c100e3f27b452f2c291f18ca4d93d
z598debc7c80c556d884ba627bcfac486af2b204e95eaeb8cefaf3ae7e46e8e5384cb2594bbb0bb
z4e2f6c96a260e8bf5e072d2ebd3e3b1c2ef4213d6408ca11f64f6714aa23c0fd445a808499a0e4
zc231ad4c4124728afe123ff5655844be513a7ec60892a72f7d6bf1d4014ac5b84e3f13e8acc800
zb1433f3242dbf7b8ebf8ff774a9c95583c16a05fd7fa0d105bacfe7f170c102dcebac3d75ee1f6
zff4a96203054093535ae5d569e365e44e207ec05256133eb00d24696434a313d8774ae3c972ae2
zd6ff96dce526b9358af64915b13acd421123abd636c5d358b1eb4242115d3af4ad07dccd18c9e1
ze55bbb8a239f19deeabd723487ef0ec7b7bd86a2e0059c437e14018db01cd94e7fdc8a26aa445d
zfdada49e20c2cca95e4e9dee1959962bfd13bbdada061dabcf17ae925e00114b8fc91146bbd747
zf192d1c57c2cc577586784e50242b8caa8939001b4f06116184b6778e97f7735f71a8d8f302ae3
z9439d80934048601d0aeb8e917287cca053da8b2eb9608d037e88da8ae4e67221125a9dc0fbadf
ze25b660ad6827e47eba55a31abcff6b2fd43fe6930260c069cc82c4fb6c121e43c836202b80975
z3dc7713488a8f5f6c24a66e66e95823c4dbd1c1e2dcc41316f27b8668c7a2471a362bca9bdf7bd
ze4907dba8870bf6e5d5159f9453f390852809e7d3d532c62e821245a5f659e56cd6241e6bc441a
z1c051f19cb065400a07e63de107e14f8df3feee3898684fd446e4dc142a4a191b592beef597b8c
ze78cc386594cf4cc0eb280cda0feae05f320b55b36b9822cf481f9a7a1993e0645b61f8d04519e
zd83d91a338234b82cab649bb1a95042256c79d73f12a119c9d79e31d6eafd411f51c4c80de95b0
z0880e5f675532cd4c52e32333f0ce3f8f5cb2cc64021c6a15ee67c9d21bbe1f7a83503a572aafe
zfe889d4889c1a9056410ab16bbed16deaa01fc6b434671106eb5f95b5dd0c020e2cb4982148a09
zf0eec32cb27cdc98bf30356f5766937c03b8637d1a491c089ab809b18192f5544d3f4e3f7868a9
z0f43600c05f30944f18f99fe45760da42962482f11593098c3f1982092de7dea86668cccd017af
z62e6d14b67163502fbbc96bebe30e145392f43a378ff54228269e6f3bc83426f8fa066c6dab202
z50b4d038ac41fa38addf59d64137198231a07afdb1655b531ab91bd09fe5c023f37ed42f422e18
z0145db3b32529c514c1b871b64eaf1ef2d498cd9800197309254d0ae1fcefae62e583ba32f0344
z273690e1a2456d229feac0d744501f15edac5451add6ddf3f50d4f9573d075ae3c6c98fee9f507
ze18fa4187a8c8a8a94428cd8d23a4b05c4fc05dbbac3c55232341e7158735aed76f1dd2fa3dfa5
z9943159683652c60eef86f005e5f6b036a03b54e3cd058afbccbab2e101b9d8856b59c310ddad2
z85fabadee1e8e366eeb48d3be4ac6796af4d25adc9aa0aecaab1d73c77cff3130ed3d8404103d9
zd2c5fa734f11556118e7ed8d43c7973f6a8b0723f40a94ec5e2be0fc440cc0289280e1a4669a33
z88bc5b0fbcadd74129843c7e67be4ad5da72bf24446f9807462d8b2683b256458e212deec824d0
zc3c0fbadcf49514096b43185cf2cec57d6a50fbe91a562f7c2c5e2e1a10c5b720a25f3a453d537
z173e195bf5f2b19f23f928f3e7e6f6fd25aa25f8a1e4f191ebe191660acf8003512b21ccd788c0
z2e5507e3e0a8a4019d060c1144daa25e0149cad82fd8c7cb457d8232b221f6d24a228ee09c0b79
zb762516b62de66acaaddc35d2f9940ec724622d6cb6400e73b1abd0dd25063684ad549dab924c4
z08bb7595c21fac7bdaddbee7111b5b8caddc2cc089825333ac2b5d2c170944e6b440d093a0ed1c
zc4a85b3d1c5851a5a493502d023178bd04dd138dbc22f521f93e636e3166be01b2e7df125d6e56
z586ef8332fe053c407887ee4d40e6a9ec47711591dafcd4321b2977c0481dc41b6fe879037aaa0
zd3a3e50c4db9138e019a8b136d8d1c18d605f452f8379be2e23d88d74a4216bd5ed97aad090849
z79339f6315a893c59f4dbe4ab6d111aed42ca0020056285b6f5cf5603c43914c2079ba2ebfb793
zb33d50e0097b8bb8735c679a971b356f416fe72c5940351db306c83786e7b584e2f118654e3565
z3db6838c18ed51df6c23a4f76307983f1056cd2fd11cf1f7a3b19e896fd011cecdb1507bef70ba
za659b837df98f08e4759ca0b9dbe8cec8a860dca23727437acd079a84c641dd74effb3a06a9ce2
za7dea04c007cda6fbe2bcf2e56b44b44a46aff6038f7d12ab83c481360b153702cad3580e3d153
zf37888a88578894d2624e4f121c4a14e4402b277aee0e3de775ad777e17a4d7f5d0b652ae9cd3b
z76d3fa0a781d7213b13d197237a607cc4587c6d6912da8db220d1cf6c74474657e1d79d9482e7c
zfe598ffe1c5b159472354d53ce5e3353b22117f32648256e3008a9e6233a175fec7d8693b2af1b
z21997797a5dd080681bf7ab107e8a37be43e6ec76a04d04540d1686ab250c3532fce1e7a4aab62
z7ec0f9d52a2aec320e80a8c00921e703535fb6de10092b6f763dcff2ad39b90389b99322cc2d34
z970664aab8c39e9679dd7114a8e99151fe48530b9cf3b0c9f5ceba3f0751c8e9f4f8f4ce1ebe70
z99af9986d1eafe162f4c0f0e044fc22a117e417cdae546a9f209a6bd078e90185ede1a93ffc027
z72e2dd0a7ba28b54070da872378e1260f42ccbca760e2688c42905596bc166177c1c7327d72daa
z6f6f95441a6581c4df7f8855d6dd74ef421d7b7184dae6363e7d4d947c1f63b79b55e9e5bfa648
z69b7c8b5196df8ad936db249a8d658074e9d5c4dbec3403a15b536e7efadf045c607309a429260
zf0b9e6c545e199acfa2df7dbd85e151d4233c328983f9ded788d2eb2fc6d0e21d0c653bdff30f0
z4db3838ed8f820602357bc8120dec6847963831033c88481460c2b8d8ff5d7362c8e02715d581f
z62de38f9662151994cf1e8843a85fb6a5012aece5388933493a4a0309daf4879c37ed47e23e38e
z808ad8041a79e7a5a42aa0976a674e2e9685d718f1cccd4c549940bdd56629f6689d5c87bd377b
z5d6be9ed89577c170be14f681adfe158b464604039a054720fae16451dddefe79c5fd4460bea54
zc20562415f3126e14b09e86589abfc514593cdf93c0a0df9e31476747f61941e8894e43860b432
z0cd9650dd331f6b867ddbe7e487dea755fa4989bdf2d2b982cef4e3ffdcee5a24e0cac0469a533
zde27c4fbaea7e44494a9eba8cb029b5fea5c10c7e9ff62d307a3e2ef83ea40c903a65e8d22edf2
z2fd586148662d0426eadf9ddb497f407044178030439f0993089ad2205df6717520eca7b47a524
z4215ecffb99023928ff51e1e99f893d0a4f0f57358000c61d667f0d25bb28f940a826c3ca41a09
z783fe3e7f43f2886ab6ed451b5dd36f8d68ba272aeb085a6f874cde2f65817baab3d2fba285abf
zaa83d38711dda8cfac7f8c133ac3a086258179e4fac5df3ce5e6e05a4fe7d68a436fac54191361
zac8cb2b7a55427c90e7594079efcd873f5c249263b1b3fb6164cb8fca30613c67eeac51785b89f
z63a2312bae45f797f6542f427a1f8dc4878ecc3a03bc4b5d0422f3a2e823900ba573a5b4082b7e
z9f7199666dfbf8395ae477e15aa7a5a2eb19f802f0a4f406d06100bf264a651197a1b0edf9e833
z60405d3f30f1e557437df6197cb085fb16f3dd0f1b20fccb3101bfd54290007933b7d03dab69fb
zf19c4f79cf24ee23e8254896da1bff70e906df3dcf377b409e03d30f66128f1685f02170ee92a6
zd5cbf70eadeb508206b28a5d4b9a37ca164ff750b1998a3c52517b74ceba6a93fb5b6116b7ea9d
z1fd3759411a15d93ef782b732b3d7d22f2bdd742743f7ac06ccf20f0b4dd1e1587aeb324d6e19a
z1ee17a765bfb920df2f35e82cd3b48a469e3b7a013d6277350b5a2a8be36e712e435c550b25542
zc91ff65adf968d25586d06914ea5574637e9bb30ca1f7879b0afb8083023aed4b1d01720a51c53
z07921bdf7a4e1deb4811d7a8f364c78a70b87997bffdfbe193960ab86e5e23790290f4f57e5d84
z00948f76817bdb7603df6672aba85bbc29aace4d52cc565475bbc6ca3b6bb78e30f9151791c2a5
zde61effa9d1bd0b08969b2a9ca5dd916542f16796dc141cbe06e03c35958492ff97d9bdfbb6060
z69d3bb291da528fc1822ab123932effffe69f7fb6b21ea7ad1152703fd4d1396f790611ef002a2
z6324584eab5cae157f8563903c6b23594e874cc4cc156ac11d8756cf246c5ba9edb85cb1a8f2ec
z8a385ced4db6b7d73c9194e809d9e613542bcdcaf8af6ccf6b6843b6ee0f409c8fd68a8e51c83e
z507439f0555371857eaf0f7a67567a0cabe77b65e73ac138fe8e21cdffe5992605d9bf7908282e
z51df3b2fb1f3183e023bb80052b0324e6fad5639dbd3a9d136fc2e29edc40b4e14a8d0469b4163
z8e8611d3c5b722cb7f22348334f2b1c2af6781b3cc0744ffe36d707e40eb3262f4aba5db3c1efc
z7eb5dd4ff18be4d74db49e872fa65dffe2e3314f27c1fba1ccf22e7672d5bdae87a8f96f7ad31a
zd9195a622f28c2070d302fe52e057febadf06147fcab94096b45ea6ccb6db9ee5bb4250450294b
zd22169791cb6abb1fd64aadf48775fdcae131bd2ed5354bee4cedf4b148bf2ea7f1eda504ec19d
zfbf5520dcd59e9e87525863eeac37ccd815f2052930e329cb84ce11d9377b6b070ebd21445fbfe
zb8cdc3aa8cf333355bd948d69f6aac87b77e92571d109f786c157e4d71ff00538808f48c5d3a29
z325771385fe8fc11c64c386c274c3ecc5d2aec07a9ee57224a74e293e1801f842ae03f137144a7
zb2044de42608f8cf9df6c1e32f107d6aaa34b2ae285719d7094fb7d1e4c88ce4a49320dd3fc9ab
zb0ee52f039f1f916205b514835e23a656c5ed49649e6265642bfa9cc517fb94f5a3c3f95bdd132
zd666bae45250c4a7b70aa61331081605e330653e7b9964482814cfd21f3f82af335d9458cd0a46
zb676eb0c1ffaa9888be15277c6bacd635b779d34d118ddf7922b015dbedc873f4192957d976cf7
z4a46839f5d51c9f54f398ef713c6f99325fd8808e0564f046389d4effaa471eb42e5f65d4fd3bd
z0d4f40978eee218b153ca0ee201533fa5b132d58bb98ddde67a49ee5aca7ef9dd66dbed9df059e
z73ab69161d15abe5458d38497edefd16a690e4d416f42149e0f10b9733fd2420c7068a62c3084c
zfdd2c5cbe7cc3db0856e4cafa87bcc330105f2f148ada558464a696d534ea46269432e22c39230
z1e075777db8817ecaba573bb224419eab20b6a6fee8bdcf5f34920f206c5631c86c67d08b62b59
z7e2555694471e007bd51ac0fc310f1dc51f3b00322743cbbfa069e404b34cc7063cd13abcc5fc4
zd475e9ba32813aae28e63141dfdbaa53e7c7a73f729bc4350ff6fdbf9063f050b019ae8d78d36b
z16a731a1bb77d2d2fa062d9ac85f9b8511c090c57482614c06f04d7cab4cb1696ca2411d699c9b
z8979928feb4c935c79c63c7775921e52d6c0bfeaa2a9183d1d9f340efaa498a0cf33990d9453b9
z1e4be853154aaed2159082d2ac9370c76d64ac9425aad808e9a176177c20f1b40d5f54d31daf5a
z608a8fa9409e4daaa655e706bc9f40a2ca61c570404fc7ca35da390d0cfa0bc3aef1c2432a15c4
z92bab1bb4842b3439d5738f6eca7fa2f39d42981cc07fc9267f9b5a50622a4ca35ddd669a1a4c7
z951678adef4ab110113cda17d926dc6ba4bbe859c6c22d34f06657f6fd4a447193dbbb908cbf62
z9dda46468996e6354e8b91c756a4dd7efa5bc7250dd5d625586f86ad77f7faf69c99e48be19af4
z075a7c66a5817c656d3be515e2fcd231411c8da1ed60378103164630737c7547addf63cd569705
z70a09adbddc95103bd7403757f8fb4db1467ef2f69aea4df94e904fb80e183fc00b7d24bd06728
z31997758d029b258375b888f14c8b8a7b8e7c23d9acaf78e5a85da0465863b74c736bf4eed738e
z568bfba22df98db035914c94541e01e01963e3094ac0b3d809e849908c2903ae008cc773124933
ze8453fe31d728c6ce6ab1f64bf92b59c070e1c9b328a20534ef0f66db2975466fba707d3ca1686
z4ff7915cb8fcc2b7a35ea88977887b5d933ea9c5f3a3527e76d20d09e95d7ac50c97146aed6b5c
z18214351737a5b61e01661c6600a2852209ae95d97aebcf350ec65584418186c4a59ffd0930ee5
z688813be67cca46102c8397c4a4c7f13a28ef952110b2c7ca57e094fda20a912b4d8b2d763d46c
zcb8b40c044e02f16d84908997c54de64dfeb5222aad30063df506bf321fabbef7de9a6256d7fe6
z3908b69fe0756ed77cdfea9826d5bc427bc41524254ee8f7af8bc9b745ef7855c1c6b26fc21829
z3ae5897797a96895112b88cd3ee14aac6ca05dadd4de6a47eee5d23c70fc3e9f8e9870609d7272
z2de5fb63505ceaea85a91e524a8f47bd6cbfdfaa5ee247fb0fad30ba148b2fba7bb9c5ad7bc99f
z6dd21d637d1d330997e0d6a9587a6349171495421edb9174ac46efbeb7e068ecb0e66e0191102e
z7e108e9ee7b68883e03804fcb1d3c644d3d0b5f6db69406590ae772516b517dc3c2784c0f71a88
z98d625df535c91f304576cfc42454d99f55e76252d94c743db9e2ea8e85a2dba713c0654b1adaa
z2f7bb28dd01a85d5b95169553080de83b0c99430e418acc58bc0a1e8a9221484132b686ffe5c64
z65b6d5020b6054aba8c364bfb083719972e093951ea91510fbd2184a03de9305dbe98b6618a721
z2905615838ca071724039871fba10ba08d01038516729200dd0d0c6f919ee59c6a21cadbb07189
z458964e96a2f82d9c018a70e866725c72dee24130a46d2f335b6d2d39300c29be2d2bac4d75c52
zc5487be2ad6da78d718ae4765100385ec2792057deb92e1ced4712aa10339e039704a5ce7db11e
zd68ec57f1261ea862441af2d875418f6ba8d080b063935c850be52d1315254a3c1b682dfab8cc2
z9f18614f5eeb8367d390b31891710a969d9beac44498df502d69e56ab5ea4be62b8cf1bf7bdaf9
z0fd6ea638594f49127cbc710c7c8bec3a644f3e42d9bb305681e0ff467fbf2c882af86406e7cbf
zc7c280ecf3d20509b6c23764b8a5629d8153fd3e0986f08de50acbd2da116484df06f1d778056b
z7ac376e5d7f6dc45606dd876d559823a0474790fb141c1dfa8f4f26ef7a241f6fe32aaef047dc4
z7a27495ae7c45ea2b137f00873d88b7f26a33fea16bb7e98d121083894e8015e387f7ec25732e5
zeb12b15c3d7a6d5cf6368ba0656a7e67b0eb12a04a7d2ebc30e37676970b6e73dc1914aa34ad14
z3635c123bc6cbb7cc9269774c53e4a180fa5acba8b91b5f19e94de98a89ec28810fb6cee427afd
zfee7d55244f2433772cdb78bbf488134cb6d815f24b4aff6aab0857a7dd00b6fe7e27256c0fbc2
z96d1da05f5ff66f71ae49c412b6fec7e6df766f3217e6c9bd7e0f4e347a1843f702b357f4029cf
z59ca4adebb5f0f8f3db4da1cfcce2cfb08d32a0ed927dc57e550be192d72433e7039465b22e07c
zf52a1dc21bfa4521a642506004a758672d8ddc94548fd1519d6a1845e8ca905d08507ffb621ba2
z161051d7e05b4cb14a9b7d36cb8ca45a195f13f49586d12f97e11bd4773cb0aa3615286cfb678e
z96b86713a20badd779a4e14a976889c30b21a6db1cb980c59f4ea118ae7ed4e00cde65619273f1
z1916dd7bd35323ead8e4cbfee3b7106021c96d0da89c1ca83c44e260e550ce94722b842b829fd8
z0309572bc66302cd5fce7eb346306460f9d32311d9e9619ff9e627d6a86d53ac9cfcd1ddc9559d
z3b12d4f914d6247fdbbb544fb5adb0a60137962fc44cb416f29a68f49e23fbb8aed7119d6deb20
zdec8d493c5190ab5b603ae6a6e4824ab7220d4f3eacd68ba54424968753b7a512a00cd23fa81ce
z68f7eb04519cc47be1d890d7c8a3a0c1300679619f103547bdde3af9d8b66b5346c42db972d482
zdf0233d439356e65beb9421778c1312b1be21b021718b82a16f51dd2d005b5b70d92895f05d8ba
z36914a721eabe9762ec8b4340ede80512a87a276c4552c0603507c9814f5f1897ac48f4db8fa85
z7d74e12f727512964c14f25447e7893364de80f4bf0c1487b8b7bbff8b6a64a939e5cc3b9b8088
z10503da15a53238e4287ea4ae390bb784805df140cd8d82dd144781de115711eec2aa87d69ce89
zb3ea0f1e260615e09bc914f68f446737c749fa89f3b1987f23772391c3b0af0a55431297987bf0
z166f55941f66de89ea03245c2649491e90c18422bef0bbf814f6c6f742fc908c83d8e8a6f933c9
zb3f2f4f5095ce03c0da04c6d2bbec5ddbd046248f79ab70d5729df829bd7316f9be9f476f4856d
z728134f65648237fe7d163b1df15a242b256d3a25f760decd2c4d5c34159afcdaf5afc77b21a6b
zd989da6448c7c063fc8e4e282f8052cf2b4d42643679638e739edfde25f9311d863d3bb392ef69
zaebbb232864ed4d20eb4c56631f4b515e3b130decc0a1784704dfff097e219125ab4c029b092ed
z3ecd223ad964a68a3793f40ee24e1d6fe88a6230579e6e082b77686db620ecbac82eb983b177fc
z575d4649531e304946146049c4bbd004d9fbaca13bdbefb8c263012bb5fbfa887892059f4d90a0
z0332ced4218f45054f85abad2bad39cbfa24033d4087e6241e89bd45b3abc0ebfa6f3b338a5518
zef47386fe3f45ac24f3ff86e7eda76c9b6dbfc890aeb83f337cced1d38483f2242efbb9afb2cba
z0c7dc73ea705fd64fea9904dc2ac1070e5949ecccd8e3bd306c52e7fb791162856701c8aefdb05
z50953f4498a16974213fbc8f71b6b40d9dddaa0615a83e341b4b0e8780349bdd5a3cc394898610
z81a0b58b874f4b32fb16c5d751647777284d16d26358d7c1089b0f999e66580af1d690ee1942e2
z3f5a95354a10558432828a6c6f37fd3e4b48ec3346102f3d4da82eac3a7ca1aeb24fdf5fcae655
z8c823db686e58599d29dfc53e5c98b1cbfb67bf9306ca4c159b29b63dc3e50594de7d9b02edaf1
z285b3728b15d6da48c5140d8d58bd68279952a610e6aa3b72af548b2340e073b148614e196ab0b
ze9f535545cfc30f40dff4a3dc6c2eb2cf2a89005d2b507b53e92fa4b750ffcdfd312134d010bf7
z96450a244c9abbdd8ece54118bc108e9ede8449bab8297b85fad400e7bcdaf87219b9f58acfc19
z7de951bd9729ea988073e2fb5b3cd6cadfe5ac8dd9e441742792b5a06491043e028dafc62168df
z2c9fd5bd4be35b452dd2c8258afc43d0efc14ca1b5cb9f0c92e8d8acfdfa1fa7f6c6e16031bb56
z380431f71d3573c758037505842d5ad62d7658c52422e794044e5f4cee150594bc217e49d56712
z4550a656f8ab55c4ab85be89917eb038e6d47244c85fb799bef45876a52344ffa1ab5f2f96de87
z37c0be9e49ec239e2845484b889250db87daca4c69efd45eab39ba5e8a90a4a29c41bc47dffea9
zd24e97b4d9db09a470701041a4d091d32db85490922e6f78e41e7fdfacb6b355f7a36a64d2de20
z99ef224cb98944ebeca73c72863571b74e06d56007c1a69f241e6f8b0c6aaaebae803e48cca818
ze06c70d858726534debf66e4c78613a9bde2b0ac4ed8fa85a55ceb815fb3a9e4806411e0f6d236
zf9b3c6c8e779546e84e89ffd016a9e3fb4d70d839fc977230940987a15259bba9469d169d1f20b
zbb2cf0f5d955248bdf40873c7d6dc03ff72cc63a6096ce09fb3ed87cb996230dcaf72a122bbc72
z7f54f701b9dc4ccd94baa2123ac4687644f152e673876ac4fe98477c4b58964b027bf3761afa24
z2336348bbd22ed862d4e8353b08685b44299398c1d2c2938f1450c471ba527a66d858d4736868d
z88dcb02dc6a4babb63267de0e7c6216e0e38bf309fec28c4f3239fd1fafd40536961bfc3f302d0
z220865961f52076fd2e030a1969722a3b04789b85e390efe086dce97ed3fea4ec17b4d065af605
zdb27fc5c5168bdb3de27d812e949835f9d4b8b3b810e91c79e70381fad67c1b4d05c070b2ad857
z3c8f1ea0009bba656451e99d5e3c648e468d82442ffd71d95454f8ae11a8d81a12c028838b77cc
z84639f326b227118eee668d04a22a063274af99a09da03875da8395f835c05d5cb62e89aef0098
z0c0d753eb623d2f2a8ebfc557dbc1d4ad2c1d23e0a0a273f64251338704a2d3a375adb11a8a43f
z907d61df4e4928ec72e8714c398682d2160fe0f5e1dcf888fe11e34ae0542c4e1473f6abfe612d
zf8543b7789693488f1bd16383a2b011b2337ce28a86f30ab5aeea9560d22bd57799785bd9da4ec
z332dfb787a2eaeeca763a8f2f923d9144eeff21b4f9c792ab18f8e8f8e8d064d5082e6d945953f
zd9602df3005d580216af494fe0e6581af20abd0b81733b69d1ac3b1662d28e646d992f97d9f547
z96ee0eff9133ac87a6a92ae6b45d8e8b48f9ff108c17d7fca2d9a80d2df4264fa694f8f5340835
z7330e78d3a8ac487aca9a43f587dc56b2da6e4374d34eefaf1235106d6c881e886cd07411bf284
z3b3e5b1f299a7fd97465163d3d106e36a05bb65bcc51541ae980c615a4ed25c39297971f3a4cf7
z9a3def0d81d451bdee8cfb85fa8160e6d3710b372a6d4ab794665f32bffe6dad8206b79604465f
z3f4515aef2ea24c67f2b101c989a74bb468fa58393c3bc839b2265617b031f99abe9717a1cb6b6
zcf173b443b57f1eec4d567efa2d2677be14101e859765917669e34849e8fd22dcd0924563e735d
z10af73e24de9abc81adf2949a6e513614894de64aa16ff62b540ad2d68f9e79d171cd8c3347f6a
zf8523a8d26fb87317d6ac4ef80de99f303d3beb1b290d9ebe252567b71094dbe2569ab155da080
z7cb1551e8092aa814388b8fa5ed68e65b497693a60b84a0cf1c827c1fa0ff82a9c3bc6c57a9e96
ze3154b38bb2a3231dd1e93cf5d96279661022dad271bf7ec6ffc53df593982790b8e0eb2124ba8
zf04615072290e68ca6a2640085593facb9e5edd2274fa4a39230f4421a618473fd5b48bacec6ba
zdab58abdb4caeb7ed2948aaba89cdd64fdd0804bf8f0b1870fe7ced583674f7257d5628c113d4e
zb1057d90179b3d795c6c972581047a424d0c08b1a1a54ee356d868e255cf6db024aa74ea29e34c
zb3a67327b7c65d1435cba317fd72dbf4f58dd7eb4aa470102fa5e92d607c0d0053ec93c1ab8420
zffbcd4efa642326894bc69000972774e27df668b2c0549a141d068d0616a25c86df4521e0fc168
za6d6a03abd2beaed2e674411d14773ee8e49d5d7b5978aef769fa97e2038fad6e029e355120fa9
z88b0abd670897389f27f99f3e9db025cf4936d70a83a9209f45b53c0262b9b768ca9d60fd260b1
z9628cf21a01c0ff0cb28963cf65f7f37af52e8e98f1cb7d36d45c8b049d498d7a59e06b93919cb
zb1f6888a615bd871e3d0454ba256e90d07a48b4cc78389ce772c2c174a23aa90106b37681b60b6
z0508d91fec22f9a29cb018cb8ae24051150bf59fddacbe72724ab2b75d56ba2a12db6a501184f8
za3bfbd95b3bc65a66c5dce882e3607c3411d00bdd6a4c82e731ec6e7d179b81a261c2a893971ac
zd57246bbf6bdd9ccfa97644ece253d65064129c296cfb312ef0cd4392bc68c2d2057faccb2596a
zc21356157675062f3ba4b0d473338a82f669762c8760ac062c568383395e5c15129d7844b9c2ba
z33155a638697e60e6c61d45eb4fe3334366d25e3a40eb3a5edf68c4c3457e991d2c5c8fab4d8dc
z37d210d76c91001070d7c4171538b6ce4baa7d77cc102073b2943ea7eb7721da804c001d945a81
z468fadc9c3f0823f54fd0fe308be8f106803dbe9bb1c94590defc171a727ed977325900253435b
z70ebbacbf2a25ae79ad8ce12d08771103f445557671acc52d876e469e6ca73c38f776ca05fbd26
z42195fb4aa7b3f636d38ce9052f0f13162e6ef19740b26a49e5c84c213f53517f9ab68d7ff4bfd
zbc88398d651c5901fcffb4a4a6077bac889d109c6b8b5f166f776c95a7cf2ff0508154bf2cd0fd
z5ce39a1a366a4181b73c281a48695bb2f9a092e9c08fdc18eb5cdceae52c40f2de6ec7dbda9dce
z95d63bdab6fd2c8cc8fbdc6868bd7a8caae9b702b193757b6b9fc04e4a70bbbd19e57c6757a35e
z611122608cf9d0d7c5c8bc04428c4ea778fcb6298a50db77f2de78d60f0ce50c92978574dd7cfa
z7e247fece828a4011d805fc7aa9b2e717cda8ee516b36aa34ae18f46618a2e00fe6f337dfb8d8b
z4fce7704dcc5e9716d7bece6265660b2fb24f959165068ac0144bdeda658095adf77ca58715eb3
z1f6bf84883765bcc8e8de106de63e0bfaf6e6486ad8e6d67c79b40f8a5c3ebb7004c2d9ac71d51
z8821693f84a29045ac6f27ce5fe2af1759500d315fc010ab32f7e1a582ad310054c1140bee8433
z1434d612d99a8f1a330e8b5529c0ad348589e41660fa666aab01016fd7ddd806a322a0a011e58e
zb52ae44422e01ea8a5bffa26c359e29176d86f6bb6c2a8ba900c5a40cc8d0f1aac9b8161430aa6
z3283b87cd6a05a96985087e9c8a8f1f43dd322262044c19c4f7c8d099622d0775801f2d47dc8de
z70a482450be436f923268d9057fbd69517ed77918657ced9904d19896da55cda17b2fa822c7c93
zbbebb7c938331421592234c28d26c1b8dd45901dd5aea1ac5983eed722e5d94d54050a451d33f1
zba0ebd3825bf38f0bfb24bac8adeb8fa74efcc3bba58e2326c7721cba3008ef62e883a2669544d
za2f99fbc82be6cf47183a83c768208c64c6141d8dc26d0cd430629e1f68bc9f90bbf044abc0269
z1ddfef9015c2367c7616303006dfd174f26ef662d9c9b77b3b80672934260841217be7ebf199aa
z459e025a85a566bdc891812f153c5b0116b73c597e2433a05ad1b8d08950f3d7f6bc71f5cf5b07
zf4fba3782eb36b096c86bb0bb0b0687792bdc203c786258e30d3cb73a8b47b8a996a58b3b8190a
zb23474c55dbb6a4c201e42b06484efa6966a8dc0687f59932bd52fafed55bc6e98e71682d2b69e
zf08f01b0c8179056467252648e18c1af8baae4dc3aad7d083fbb5ad0ce4dbe4fe5ebdd23a2904c
z88357a83cd63d6623a5a2e81a71f1a3180b553b53fee843d9bab05e5882310aeb6843ccdd84f5d
z6a17832d0d34368337c95af3b9e4862deadaff2094db11c499b6357c4c772c3148c33dfa6505bf
z28c88f0557b6d9cca14da85a266cf40ce00ccc8b413d50c884aba2007f72df2129612e8905438f
z5e28e2202db6682c9884b7ba6b6da3f04daec28e4dba87a32db0f0e95804f22ab8200b474c24e4
z93d432ca21385bf10fd5efc7bfd15c9621dc038d303631b9c850c10db55ce068305837bc6f065c
z5b6e6ab75219ba079d8ec7aa8cc6d01280356d0005d041f7e7958a067e62016a09cc0028af1136
zfc8fd5e48c3feb8c325b76834d199eb095749347a4f4ea7babc863a2a76fc2612789cbe7cf803a
z14107f7ce7c0da7bc0c79ac6961a9c02187c6639c5f7d4c200b6206ea4c248f246f49807b7d1a5
za940f99f7acffd5d2bee61a68a7e93f8065d0efa369a1b289422295c7bf3926722f09f847edfba
z81551c391f14984fb40ea8aad350900fd3e649cb4ae0ec4b64cbf9b0fa9923795162ef62d12184
z7cc4f4f461a4bef5f6699c90e64c607e7411e69dabc78c00d762cb7760f4e9d32d083ed897ad85
z1f535ee2dd4ed4e35b321b229b3acf5df8ce3f00ede098cbea1a6b9495bc3483ff52aac92b9574
z3b48e871ec7263021d8bd78cdd5f429f825aa72a936a0d0900d3d010e81007a0ceff84aa7846bb
z7fabd6fc4ad8c23dbe7f63de8b50bbbb3c37f6371f0a8842ea5c886d0b494f79c7c276d809fe95
za4ede99d55d8215270171090181e12fc23419caf386d22e0c14c7a7b9e941054b6e1fe7e90dd7e
z6544f1572503e14132d2ceab14ea134716babdd1421e3e65d7461dca26caa4b62f5634e6bf3781
za722f06ca853abb5c264a9b938f9ffd402315a5995627289d2ba58a482db1579d6d5b6465f3e5b
ze458406cc993f3f52ef53fc62586566344d51dabbdecdcd7a97be42b12509f128ead798d2692fb
z08d014b611b80e90680fa0a19c3529ca97ba961f41e0929a22507586a4872dc77a22a97122c011
z96389975f3ff1b962a36a258a7b7a334a799c1900c77d2b4009c169929af610a557a5c6ba6099e
zbdfd1d2a9bee175aad86edb2e1428b3c7517b24fcd38790f53ba917eebfca5de9068c59b089249
z0db8049e3a08b2d1d4b97812146645f57133a88e5916346773c33ea93d1f139db7bf4d62f356c2
ze8224b71dcdb68f5a857b9e2d10607fe59e8c5779c2d0764c0c32ec39166eaf80442090dd5d4dd
za548400c8e2e8c769c7b0f21cc009c41321a8c0ee560d99e5e6c71f0c0ebab1bc63bb67c058f24
z62971da6c90251b974e2fcbbd35947e3b007788c1a9e80c16bc7bfb582725bd599171ed04e98c6
z7d191951b4bb97913674baa2d1a4c74431fa594bbe782a8c1f45c9d50db60b54730769cc6a0f81
zfda3500f8b9716d7824425bc77cdb642149c4433c4b476bbb5b73796bfefcdda5973926161f249
zcd2414edbe8bf47d614dd39474f39b2fbc2c4d5b646966dd8c85cc8398bb8b6121cb82a70e6ad6
z7ad3e80296bf26dd5a9c34495b59ed9e1bf7aeea21f895de5b17723fcf0637787c9849b3ff4c3a
z84cbf2d4dcde286f1c9434f17469c76d0342da24ef25f9548755c9552a761cc09a0646db9b57d2
z0cfe9108d37651cfee449206456618f19ab08853b4224a76f0f0d78766b4b8a5a8b93203038e35
z400ac936c8c2974e552f9b57fbac475b65d0968119049d378895bf1dbcf99184bf4ad8e3612865
ze529692ea099c6301195c1dccdc41666bc3394bb036839c9caae80d143247db64fac5068ba5b05
z287ca91adaaa010f1cea9e0b487f247a9f975f4148509190582ec0d979b561f32ebebee07bb2df
z3c028cf1f18605a0ff95defdbc40407815e53f8d5b33f568fb9c3548f27f664b74f06150dc669c
zd8884d0cc44338a56894f0c3564693fa9382e90f157401aff33788841042e13c72a202cf007484
z384ba361736fd09ea7036d49eb30585ed19abd750364d08cb5f2798168ff7f8a824b9d1d7a4e5b
z1d7a52d7561f0d8ccae3486fd03e9245fc64bf0f32b5a1442e81ac2be52d0e92d2a9a048ad9dd3
z71a909910dfc70d5075febc932596093ba6b4a2d06cda9952f392b97eb65fb8e50be0bf8d5093c
z936d294a69736de18c312329c90d2fab37b06ebcbb6b2c4e5c929916344ee99b0dd36fa62058bd
z4e2aa3159f36e499f7b502a6f685a1c8d1e0566695d13f4080dd11a8e2d9e0721300b61a95faa8
zf0a6410d5d27d2f50a5c4726f00a600053e9ce61e1654edb81b50da03c6104a472d96237601f62
za9701180a4d2726a4bdf350c8ffaef7a1bc3b0e9c0651d2a63dddaa98e9bf283ccaa4aed4b8134
z0ce45d2eabd719d87bed1cc93abbca08f9eef85789e8320d31cf70e4197a754e07bb9c5f1206f3
ze47942beeb49b5c91363cbf6134a2a8bd7da9e041bb652201b7c767b6902ce3a08a07abf756f38
z5fe25cb1d532cc3bcf1e0507d04aeff54c6de92d564511d2d8c6462260bdaecac6bea5e6d8d65e
z804c3edcae529dea5b45829d97570cdb46801a810083dd0701ec3958e9dda0f3c03edead22fa0b
z9da5e93b413af5b098716f2cc6cf4a8d51ad53fc60f684882668f96261faa40d573e0d777ab444
z46285a5840a396d7967303c9f732f51e2a673858f1731750fc7cb8659355b898ca879e64a7ac3b
z78dde3710e9458d7d59ccac79a6b1402506435faace85464d05ae68c774ac02867f99d0f238358
ze11f1347788ef6fb0c1a40b69543d61a8114694f4cdba75d9f2622e313ab069d8b4a252a755d70
z79f33a4571a615f3344f2bd599040775d8d9b21108f00b629ea499cb6f30c4043c69fbe3c4d01a
zec734a8e706941ee2f231c4009be1d533defd304d59630578c748fa288ff1eab5f487990943e67
z61faa96d16c9b345bd741d0350ee5a4a96756ea8a55fd6cd903ac6a619c07067f0c5f1decb872b
z3e9118e4ccee69804c5b36c0fc2de4888e05caf98b6aa0a9673cbac4d9ee71946a068c0540a422
z885c1b49f9960f49b1a82aa0c692108e934fdada732f057cfbbfb015a0c12a1c0601cd5cb0c5ad
ze716e2080413189fa0010e781f8f27da0871e09229cffd35281fc9937099d32ffc5505c69e72c3
z090dec2171e76d324df13f0257e9c0d3205b0906a5b229e9557cad58f6922434164f697dc674bf
z8fc921c4fcdcfdd289f0626c9b170be664636c54958e39caed0db34380d033b3a3706e2047aa61
z09a8a84b83b998a582f15235b59447bc983c13b31c20f9b6b25b272c5200b0115e0e23cf511dcf
z9e822a8892a3292e5b6ce1311b016d7592de8e5b551b57059274b75713cd426679ac930dc40a31
zd5b144c36a5b58f84c1158b698e033e50bc1daa68bf0883f2d586d06976c02350372f02eac4b9a
za9e28bcf79d3e87e3bd5f20b674bb8ddb83fe9951ec350cff002f28b77dccf382c668a2f206364
z5b86373d1cc780de71b145116cc611eb3fa61c18b7eb287f88c484aa5d0376dc38624b04fc7c5c
z14463cdd8d685dbd84c2435f6717342b49178e1633fb6b44fb3d9c418663dce64c45c31daf86b2
z145a62b3fe2b806e53feb9e51a303efc38e6635342451d700bcabcee285cf547b9d5b870b4688e
zc34c2c563c6496637742ae1e2f91e04e6ce4ef2ba749a08af9a86ea5974716512938b287b44a35
z2441dfb4590d2d566b9581990e8ee3dcc0805ce10041e76c11909477d857e9c980126481323343
zab120b36c1a104d3d22327197696566283e876d1bf84105c487b20ba943554ac4aa3aa2aaf0adf
z94656028a86277a5de8e46bb65b63d7c61f866df752d042805bd3aa6cec8343e29530f60c804c1
z4169e8fc89f9edab3bb6ca96c734c1ff1d6ce165e43d2892681f531aeb006f80ae47d27f71a622
z4aa11b6f9d6ee3c7c0e17ba84579ff4d1c7cd2705b7efa62b564298e26b7dbf82c682e334e73bf
z0331d3deb2b485b5e0a8c778bceeee06c8fd65c8ac38a292a8eb02d250dadcdb1235747ce6f88a
z336b1a78c22a520bb9465e73e9182f0e8de85509701f607fedf76d17fc168be3be23825546d239
zec6ff811b5436a1f06f7f79eebad7232d2dc12640b824575f22ba0a38857a2768249d44cc363e9
z93305639e3c33a86d943ee3f25cdcbda714fae674574b9b2b1033758631cf49cfac7234ebec009
zf2834a92ece59efc1f1a3047858e3ec97574aa19e0c3dcc89526d8dcf054597dd8f65ff118d075
z9b4b7c3d8be7267e501afec6669f0f4fa6688dea283389621511844c957eb9cdda961686eb3644
z0465155b7b758b129a34e283a5c6d777cb2847f11081e5e2a2623e2a4498ed32bc7d70bb433c62
z633e2bc2e45689b96f81e92556ca2e091b918ecb96526678f3853efe10ded332079fc3af0840b7
z69417ae4570cbe1fd6918cf9e0329d33d66e2a7300240c70e9fe12c58c582c132713b8234e700d
zda33ff1aaf4dff35e2ab711ae97ca91795ac87657b535daff6dfd72a23ae7fd42f29b3985b96f5
zfaaf542194f4c18358d9ace4868639a4e33a295751c9f167622a42e0ecc02f471ae5daf7bfae12
z0d6f80afe40748642907367a68c2ece73a14175f1e7d232444f5c20072ed1762e7e8446c34e960
zbcfb0e95dfb719577eaef33a0ea32fa067c88e6d418f948b1ea51b50edcf31b3241a54d741749d
z6eefe7d4d3d9566c3eb178c342457e3ebdb2081062446247065b6ab1df06fe87b82b4f8eddcde3
z43b124d560b2c5b50a3e4bfebd12e9f9946cf8d9e774f717d8a24256eaecf6fe611de3b6be712c
ze6eebdac043344e5a5904d407f3efbff6a6b87ff224c272b33f57aa802c2adc920dee6294f588c
z06b4999beb01fdebb68093b9a2024bca869f525e8d801e490d545488be6f50852c9496a8d70a92
zeab23c572846db534613b51fcdb9d5f3a1e6335ee3bc2b3c13a957eeef9c159572e91ffd4838d1
z8ffef27449fcf226a7843ab859aadd808e7e525409f8e45f9a96ef80bc4c5760b63a894444ceb7
zcbc9d6463d0ff88d709a7a3c49d16d8f7a929478cd42f1f6a55b76e6d63039db1363b496a9004b
z4abeaf28539111b4288500749c3d29697c7ae0343cd42c7ec9ac94410fc7e95b4c9b0e3a0f5e39
z902ab1da27214a58d1e5004d52ae3bd0ca3f317a795e89e54247fd3f07adb0f5ab12fcaa33c94a
z092cd912c86b05e985f5668a54c4f20425616223294c6dac852c37edee0a983baf64912055fef4
zb3988eeb0077c10b5e02b1815aada9b03702e669355a8d347eb5d23854cf20105fe35f7d61e3a3
z51ce70aaa13b0670d32f1bd80c2635d4e4eff6b36830c093a66f8f718a113fed6137964eb7c2f9
z172fc7576e2b48e6bdf48d1f7845689b1a10d9d3e97a31003b0facea34a3f95ccc84b3c86f964c
zb43e6c608c63a84c9961bab2db72d232690afc979236ce39f096a263b568f4fbd029caf1cc127d
zf40157caddb6ea39b48d3a5693dbc16b6c5311e07d75dfe768514bbf69d600794368b3b493e11b
zd4d081fc7b36d9cc4d61b58e0def4b1cb65307f8cf321cc370ee5630e7d2f854b190eb0c8a0ac1
z790926123ff45ecda49cb4bd74d7042b6978183baa07424e0790984845d9fd1dd857ee96d1fc5e
z8276bb22ccf18a38ece79e50f52ff78306fabfab8d882f677cf38b2c34e3c6053656091453cb14
z45b104ee8105ca2ac8e80a282ee8bfb3f1a911bfb87651201bdd139ef1007906dd257f0436acb5
z75376d0a9bb5d13d3e0c7b6737da172cdffa51e0138d31d87cd6a62a1dc0842469cb47ab6140a8
zdeca2dce0f15ef3e3628a8e954c3a955b424e576824c6ee7515a67bf108a6938a0e3623d372f9b
z63daca4da0fbc450a41366ec6a1130505704ffe66c6323497ad9bfefdecd5191bd9607e3579f3e
zb6025cfe3ee6a4df26bff85b5098af63b6ada8b65433c706480163dbd76676dddc7fed7ffc442c
zbdf372f33858dee01df12877aa47e233fc335dce1bff071a0017e3210d025bb3be52efbaa42c28
z638b4ba496bc0e9fc7755ebe0d42e249acadc1e771ab98272c3e31e2bd23bbb51bb42705aa8990
zda99e3e9934f21af66f7b51686d52f261786819062d5c09b7bab3264a933eaaf79697920940be4
ze07bd7daf31c440fba462473aba6b23580dbc8d13b255d049abfb17090de6996c86519f5ef8b7d
z56f5a92832a153eb363f2936226fce5752385d871d824a4c7d4d1620a9253ca507d9baf4d1245e
zc09a27a8166fadb45a7d0802d5fb8b3eb81e8480a40b73bf27fee4d0c31f1f6a673de66a52b3b7
z94a0f37ee0ddce3150bea9cdbd5f62204e97e65632d4876f8bc23fab7bf4981b8d9f24660292d1
z6fee5f3abe31cce29f5243038b026204cb7f1b607b59eef189589e6d34d8de4a4eed6f414b433f
z26b03d3133861be568490d2a08c5c959e05f72fcdf57240df3c99d9fb2cb88cc946e378eb7af53
z78b21448911dfe8fc9f7e1cd5f49c07363ac5860eba0dd63206e69435f4d198af384adb0a42445
z1d13d2c0be59d9a5aa3c45c7fdb5099a435a3552dd727fa41e0ab90c73f98cef6bf31b9c4613c0
z6ce34fef2d718e8e47833a976f1607670004e9981bf8200324db81884d6eb3d72edca352462339
z847c5d7af857e42a552a7982e39f56679817093dde5233993b1e662ca839b1952e1be5f86d478b
z330afc11f19019f42218840f313b52de5c3635379f572c07c163e0114a061e1af22c305881e182
zf4817c91c1519d103999b4f055a33f399bc83153f8dc3e11defb99571afcaada42230e4aa27883
z229c254460b4b5addd38106cddb5a6e8f9563bcf5729e8420af2ee3b0093acaf6e02044132dccb
z86acfb0a5c79f8191d822863c7b049617898c1fa7a04695f17241a066c81dcea87fee28a080acb
z2cdee9ce3936874eed7de0347a0e29fe33b39079890d9a52292c61e2831e09cd946dc4aea3d6b4
zaef869bbafa5d09739652dacdba5e34f8e9903c2bdcc28f1c5c6705d36f861c52611ab0169b6ba
z816bfb61ad159fdf7169e7db8e9c71fc21b62349e128d4599d712aed6abd72a8ff697b5d425f83
zc9a69fb0846270f6e1174c6e11fe6da96f69facd336d3b0b945f2391034f18f94b6fd7cb61fb90
z8584418e7a715849ca32097235a1a874394dee0ada0af375fb0479ad7afef7a1983c8a944d5ccc
z9682c564d0b46e8e6945bcc5ba06b967997dc276720bf8c1ee025adb0298b48c455164d78e4ae0
zd4f0fdbf6bcafbb5d85f74ff157f317af56d247217c1879b8913a7573ad04e80ec41bbeb4503d9
zdc68308abedcbc101b7dd466824cc1eb518f86cadbc3faa6d781a05e436fdaf33cc11672dcdc9d
za2112ba8e9b79824acf718a319df4c81d0139a76d4f45c6f746f49e741cd1f36242a8c8f8f4e5e
zf4a11c5b2e5f04ac473803ed340121136ad6068c478c5dc246237cca8c02b21fda597114c76ed0
za7639778dd2e4b23462ec22883d57d655925d1b5aa40eb74fdb2b3a86e80d8a4c9f11d5e7424fc
z9e2fdbf8aef13ff36d638f6a537fdb1c18d07f4753fd04426db696cc2982e5a4cdc964a05417ee
ze1a803531a338189088f31bd9ef3d38df9344764a725bc435141cc82b899286e8cce2375f6f8bb
zee81b3362d84da42b1f1e23c08853e488f55e3381f220d648178d7ff2727c5f3376d4e45aaad5e
z09dcbfa30b9c8b0829d7fa25b83f0a694aec076b6585666294e6f4a843fc6e3b43a45c9e7d80c4
zb8a9bd8c0a6ddf97f6523e5322bed7cd3e47bb463b5e79e394463b5abd09ca05ffc4d7f35b00d3
z48ea41e675ec307695a7b058f49591ed529020a82cd425e5ed516eca73a6bf020ee314bc7596be
z88ec2cc9af84341846c7e7df8fc90024118e6b267efae801d0e18a04512f8ad236a56b7ffb16fd
zba81947e4ea061c6a8bef7234c661e560910db54f621940982beb1a77277368f7bd4dc7aaea789
zdec21d39cb87d88019d74e2a1a2fbc567b02eb2522d791228fa9100f678648dd4dbcde9abc008a
zbb3262eec41a8b1b9105774ecc9cccc9ecbb24911bcd9034395834f22a197c932e66be39dd170d
z5dcd05bacdb140ddcf08023136f0df4198591ea5dcecf743a786bce05aeeb006a4433f072a712a
ze1b111fb90acec2dcb53e0064db25149463a44d0e7475a1374718963deaaca02513e1df8b4e40f
zc2f6e5f15e83a68769cde13560c95e773dade3087d5ad8fd3c465ca7a62ff46fec80a68d3f502c
zd9f7ecf1187bf6e705bb8e97d00875270928fccf967337cb6167dad8e380231e5e942b02882564
z2b81454d3f37505d6d14d0ee93f8a121adc2822b82ebd676fddbfd221835e7f21ce06251421336
z76bdb9d37b2f7bbf622a345edc90922f5581deb255525bf0d4a0502575bde97ef92ea0f4b326ac
z0162a1248cbbb0a09ee780001dea89af7a00f9dbdfae781719c37ad6da85b1786fea94b4584001
za5345a48acda49621a3edaa0ac90ac6346ded73c9b84f0bc2b6ddf41c66dab531224d1c6a9a2a2
zee16bc91599cd404e99887d21f7862198c81452ad0d2685e35bd070a2815b254cb45f607f8c157
zdfc986cd7f4691c8cee1d5d35e95d16cdeadcbac84eceaa5dc79b8994beefd2ff85ac68038d465
z89612cdf006930b39c7a8b0e3f192bc36ff59b68c89d3718ed7b6c938159b8b894ad98581ea7a9
za2ff7cd0b8e3b06c47022b5edbd22652f25062c243f62e20bda5fe3705f878453a1c17e8568375
zca13ecc841f044ee71a6815607f93adacf633423545a1577efbf389f63c703ebadbb2db1dd9907
za6e69d81d6bf2e8d2634c7b37f622af7bf1b10a44c72b7e00fbd56b3b4e0d6b77d188d562cf8ef
zb63112b9dc5818af1dd8e5367af802ade88e1bb6286e4d0d6725db05ec52ab9931bab32ebb28a1
za2ed500ea0cf54cb38bc9c4b3aacf00068f2cdc057dbfccd81ed18f4b7b6ef7f16527388c8c857
zf7c1c9085f4f46e29f1c1ba57554016ab630a5de248968ba8ae1619493836fc484e818f7ab2376
za0f3ce15842cb36f4bbf62572fea1803f1c28894f4553329137745b787e1d6e48aafb19d73a3ae
z47f1ba8a509fef90a76c032d81a2418c7e65e5701a149b3d24e34d4da02b0b9b2ba8bbc03382c6
z5be474f7e7ecaf0411a965a4d9b5075b570cdc1f758f23ac2a64a004c886fe8066d1a1430ed501
zd8d684c13119a0e0c170742abc04b3ad6f53afe384c4206d248c50d8348779423b62ef767498c4
z878cc0e019221c0900a8c595063a534b56cd3203379d501a8e211a3f15fb68837633b3f78ee540
z89415580614b7963fcedd81e602157a5cd5b5e691403576bfc0a33422a025d3bfd4e09cb20008b
z1d7a274dc2fa99e3411ed0b07d0b69d30c4c74507052dbec9449de4c3beb930950875f6f7e4566
z44227753bb807b9da5e20453295fb5b8f8f6d5612f923e3218c641a174a6702e8ee1c02d6974c7
z1982fcecbe4c79c9dd796a61eec5178220c44d77c6bee710a3e4eceb7da40e4d61da7a8423067a
z22c1ba5ce1c3bacc78d6d986262d45f051b782e1f46653c8f7861e291875a49ef88e51e8d469e6
z13b373a24c52ff3492f1b4580cf3dabfc09d486db5136a0ebd91254c7a648bd650368d12334fda
z31aa357645f075d720a5785b7685f2ea37a4316bff7bba3109b7e03acbc8276782c24431e06835
zb1527196f05e99757876ad7751f9ccc1e095cfc9fae254eeec33f678a74d6c0d37397abde498fc
z56c7bc36da18489ccca05f796cce5898800aeb7273006d8a6d51f7d0d651ff1dcfe4e7703b36af
z7f2dfa00afe0b618ac1347389a52bc8e1c796d9248c69f1349a6444a37186d859a58cbbed44593
zd68f97277215581bafdbbca613c8094f6dd4a9542a82c80063469baa2c38090ad50652c4b5f9c2
z6198eff479a1502a4e87f3074383112de2ba744325f2bdb42c492642eabb563dfff9cb5f6b388f
z18047e97aa5a7eeff7860f799a6a7ab0e41e25b13b320ec646a14e141a8f1be03dd3ab2e1b2d11
zcb88050e88419d329d9cc4c8d7f13efd21d73dbeddf175a3aed05122406baf64405a2603429c3c
zd6f5b98cb23ca228a2fc7245113eb18a7634c334914ab1b9c19c124e1ab42b2d3f5b0b717d0e43
zdd4658b43bc4ce7cec5a3a4f353a4a213f29ffe27b820fe91cdf26806b392f120647251e09f4bf
z4cc28cf7a40d93e4dd0c0ff28c1af8d4f72bb5b5ae1c4e0d897fb3548eb10b93c3969a13479792
zedd4fd1d5d6a65589b93ae1526e0e3df71ba0ea6b5c8c0e9bc5505e9f02f93fb77ed1456fd969d
z9a0b11544be6562516ed5d1726d7352460c6177eb9bda4ac127c16a4bdd80ac28f258566c4999a
ze9f0f187394681bb629cfea525ac44570e30249cc669d7b673463afa25d841322e25c0e7cea3d8
z2a4d3aeae7757ff1df48f620523c101e91139b0c3182d0d27530ac38cc86693ab608285db68eff
z6f2e76785ad8d3f98ac0598182a8da1848b6f3b1ec2f2ed466c13e6515513e0c1c8ba22e94ef30
z942eb323ff3b092d8e28e9cebce444550872c1b238eb98c8d7da56128f354932469576f9635982
ze95b8d6fba07c7291db012bb77c0023984f483dd8a6124cb2023996f71d65926c0deb7f2a20988
z16e0a37e312f1b243afe04494b9b3e6c2828da9296cc4a52e972eaebc425b5eafbeb1d00b81e20
z5831131e0940175b9cb142abfdcd3ca81585ccf515bcd568e7eeb8c072bf4186d951677edbb221
zd2b20f8a70fb0593db63c869cf1632bba6ee0586633cf39526745a37d4b192b1a57d9da39c5dc2
z5cf4b0ed19d0a968a2c1f7e8918d92dc41e26413b1823fa3c637cd1068eae39a6b701479e1e3b4
z1d6e6ec5415baf87df637dc19caec3aa5e56ec46f27b10263d97450625965392ccf75ae812c814
zefc5354794d54e38073b881359e4e8699cd89ad59fdbaac52948600af83318c439fcba1c08fda0
z2513f772eec9b740922edcff0e3e35e2b7803cdfd659e66c346a83d5c4e8381757f486eba84833
z463fc6038d15a0ef9dd266d2305cf9cb08c6d6ed1111cb527a46821510353020d7f179333ecf09
z067d46be682a1d08e511e48d5a1495c504b0d0e841bb323496a93a7f768005519612aaf1f150fd
z8cdcd775a3cc0ec2c682bffa634971760aeca272493a05fd478b9f58b9aae4350516330e2d1e20
z3fa613e9bcae3616bc3e7d99f90aa90ffd0755c267dc8e5cd168d120788caef3eaab4cfc48b339
z7c807326c7becbc23f92921d52a3f23eacf003146383b9ac93b2169f6918443fd804fdf6875e95
z434f75248f1cf73fdb35de838115fefe26bb3daffc98ae8d10d22e3a44a32237c1366feb573ec8
z3e261edcc88778b821f85b4cfa7dee865b179e8d83c3e442fdcf975c5726239f693509416ca3f5
z6debc3c4d1cfc5110035827230495b3aa2eb24ec31e7607158e916aaa7b005f3ad8b8382fcbf6c
z5c2f543d9bb00332ee67723bd790f396d3519885d8c4a62779ddb3c02b1146574e802d6fae8c64
z7f3685e22b718ae43a4e37a5fdc44b66e62c8fdfc58ecbe4e65190d4a842ae6ea95e3730424826
z2db670b4a68e7c5bfd2738664a6a8ab3a052a8863b338447db89e1f37efdf5888a03ad3cfcb1d7
z77dd31d07c3f918197aeda4ae27e9e573f99a59aa2ee571beb9f52617991c7b26fc743d3298016
z33a6a7a9d82bdf7170b8b8a855f4b015bf62ead065594dd8728c33fac593bbb5eca70fc98565a1
z433107d5cdac4b04a0441952edc90e9e15e4f85893943047ca2a9e2d763804d72fd6094ac3d0c0
ze103dc117389f3b6d8cf17bcc991929456869d1e9612bdaba852e6835eba2468585e2e4c381bc9
z4a257b9599adcaf93b08c9015586ef305c546cebf1c793eca0ace1d222c06ac3a8f7acfbb30ab1
zd10b4035cdfb0e312db42bcda156110c07d690f9631e850c3e6d3dadab6502f8750b0ad593b515
zb4a55001f02e0d222cdf6c7a06785661048700a8a8633a17edbe01f96ef616c90230c06ea0e8b2
ze4c39abea46d25eea70e760968cde62500d44f537d435d1d7891dd71a2af0bc0cd7f07fdcc4ffb
z457b845041c589bc706c60aa33d015f4889f4c8528812cfc6c58b8e5ca1b972262dc275ed2b760
z525605ce1eab0839ebb65048689e1253bb4bb08fe6ada961e7af842f273df130049b1470ae9c64
z7c179f5dc8f4fb98723f8b3687ce4b1c8f1bafc78393619dfd5d4b16222309b03862f6dab781f6
z4ac9e6f6f2d7563249398ec237696c4b5e9f4e5b932c839aeffa99ff84372b3071b5e243ed7eed
zf5a664fc16cd3cf37f82799b4b64222fb5c540918db7f1540764df59cd4eaa861c7203ef8712ce
z70779dcb99af8c9b8a6883ac1fa66d6667d261a6c450c32247f5fb1834dc01372c867ba7a355dc
z90a3e34c18f1bd761fb28649c79e893ed87137079e6b1ac2b5173ea3d5949db45e8afb8131c4c1
z72c2934e42e0769163a2de6dc0e0fbc2c1129fd5be82c2e53a65675a08893e2b0926bc221e22d0
z1b5d4aa50bca85488caa844f585265706ca02bf22607be526956b7776afefa7f6a20056c3eb4c3
zd0236b36928d6c01aa8b59146bcb52b48792761090e4a94f5dd020720a6e3ce5dc31e5461b23e7
z1e976412d8a1cbb4ebfbca3cd7a5b645f1f7245abc6df3a807df2740b8aa29572a4c87a78ef4d8
zeaaa5b4d49fad48b87c05068f20f440373b9f11754e28a13239341a2d31f3947a4b137a00c92ec
zd3614cbf1174d67034d6f9820f2d8840da57b60052abb84b358396e53e028826ee13c83e3be8d9
z74a4dc7b91f914822da43c7338939071918cf5ddb698257b26d120c382cf4705feb56057204a21
z1dcaaddd3128c36f12954ed7f11e5611793c34ac29c638ff3a6ab2b0c6a15b3db8e70c7eb3e330
z276b2222e978c8167b6f0e5468cc0b8e8d80509ec02ef61f35d01efaf254f35d2e332cf6fe3510
z01d253f257c25a5056048c17b04366f87f744f3377de27ef4440b75bc1017aa5aaf7ad836b1e75
z6e3b4b944fad32a6c1c6cb8a1087f2f2120f686cb1e750e4657ec53c5890dfa8d2ddcc0bf0fc59
z60cdaf5f4a4ef3e374753238a293ff970489475736ad96e326539f9e14d12bad7ecf064ecd8e22
z3aa7816f7bd8bd77fbb1aa5d0e8a5351fdf2b8b453e235af638942f1cd2740b23c150f34c7f9bc
z733ce633e627e711425f8d37d6aca5183e4620d5e037201c69dd5c10bc0094914913056b0f2fc3
z376379da54aa044f95f7cfd223f5d20d80b585ec76b5cd450d04cf5a1eab7ca451282d727eae84
z3b8fd3ac7b80472517efa31694c473e970555a149d9ac6b676af0b6936c66ef843ce1de3df4dca
z39b07df314cd621a78c8a5bdf198e63437e3b33a240a7e8fe16f5ded32f4665c1f07af51e1f30b
z4abd8c5be865814630275fd976bd025def7a1f9f628eafd9eb0f98be4a10419c66ffbc53ef3ad5
z33ade0335a2858f923a2ac785b10166fd602b1cb30a4de37c49de76e8d0238d72c1907c55d8ae6
zf3a1065542cb92eb915e10744ddcc18c58b02ca19936fb860ce26b1c1c73c4692a0c5c6b241bfc
z37bd265af9ef1043ef937b44c8c1e21dee250380ef0d517a49d6fd1d5f2b7a1bdffbe2ae8d48fe
zf9207a3559af50ab57b49a9ac0d8e390b9d1df470625a75b07ab2b5294b008401dbf43985e7b82
z75f5006c632b17c8dc7854b1957792a3043fec066a8ff276a19932d8858d4872372ffb859422f3
z964cc8fa76a54902e8a0bfbbe4f30c9e5ba90cb0fc3b35f3596dcba9e69a1b1b887563b38f869a
zf5faa8e788d1646ccfbed42633b9c9e97b6d1975ae1063c3dfa061dec37f0ebfa2c4a09bfb91d9
z5f568e88f5819e3a4ba94273e7f709d6999b6d15cad3bc1168f5dd76db3b67d4c9a4468c2d2c6c
zc745fb28fcb959b1fa2e0f7eedca8bb9ee8f26cda4b0177231c090c5dc66889e00bc33e1c790fe
zb9b87e5738ef2a4f4d9910cc57135b4d6a1e0e0db9d5afaca8bdee5cd7a22c94e4f440324cd7ca
z5e579de658b1637cfd1b811b265bac9f6334b864580f4eaf8ceb29fd2ab736711f51a24f76449b
z517f420bfc2f897c84e474b4b53d1ca2393b218aa9f0a27d3039406d736fe7486d2d447d8cb8a6
z58f44d5f4e47f7bf6783bd6d2ba22c1585fc71237d44e726cdd6efb71ab71627e21c69f280f297
zd41439e35d2df67703d47c419a04fb23b7df9b6ba262de75fc1efd73a0a5465a0b35eb8445a9ba
z485f76fe72358642bf47e6532290a0a2f389e0a0307a491f6062b418419576186ee309e977e225
ze33ad6c73c6daab6d5263b64069ad76f49e2d936176d568553f5e32ed70aa8689606fb92f2a8c9
ze2afee7db3c1bc65a0a04101f5d775345b919f2b52cf5660676fac648512314fe17d9ce53cf0e2
z68d72732fe7fb84e34ab7b4548e01c9d9efa31340a5d784c31916165df7a76234bd8d9896231b4
z145ff255a4d8c68db43a2376beeef2f644541a1cf4d47aedb34b073db36d5436b093c8caebae50
z4cba8bfffa44f836ab09bfed59d47959f6bf91993b934e2c1b1344769d723a0fdfef780915e94b
z895e1f3842ccad54610f92082aaaffb2d994cffd0b2069603e7fd7c5702c0b9176e53c486f84f2
zd0e13f07e792c5e2a8ddae4ae464fe3322dacafd819f8508950c84f654fe64074bf1766586811f
z87edb84493d0fd8e06ccf482ada2b5526bcd1cda194504967ac1ad4da0d5e9034f7a2f2e3d4b9f
zf7ff5f41e821f4847adbe5042d79a60e6166559b1f16e290190fab794a5ccfee23460a60bb7202
z7807a244397cc5c09234b0b025ed1f7472bc68ea891367ccb3671900baa0c13f8182af470c1304
z4ee78a737f58da2aadd8675105b3a774055fb6352725edf909e5a30227f9674ba8bc8a183f7aa0
z8717ef77bc58274e06bb0ba805ea22bcae7d9076cf8be3b0211678f8aeca0c362855f2654caf20
z6d68aa53ba8f40c4a5c92100293494c846bd53d4a6e67fd39229e19fbbdd2502537d21865a9ef4
z5df30bb5b571471dd1398fd327f3ca6158f362253f07281647ac4857989db4194dd81c2944eb73
zd2a323a1d9b20277b16035f99ebd1c98a9e78357e5cfbf76b6e86542bbe7aee729b3f336173383
z1dcf038e13fa1f0bc5f4dd5798f6e091eb96940abaabbcbec653a899976bdf1277af53cd51fc87
z055d54f6ffd2355967fcfab19289b14a63ecd555a70194a87a5ab1fb153d0d8ac978e0aa5eb336
z25980daa896c3491d2902c8cd5967d27afb86f1c76579c854c19001950eac8c2cf74c5b9565d3c
z2b534a327d8afa1687aac9a174a8175ca23d863d8a160dbe66677ad057d6097fe092b27c6ec2f6
zae8968ae90ad6554be592ad007f592e0b37d7aaaab161c4701b0111c8c126923cbf4a775da164c
zc76a5784001c8b93920077caf4b270bd610d9450d4f0ca893576f887368dc7bd05f0225d1e7b72
zbbf328e14be6f359f23d2e8e7be3a3df68c8c8bfb70bb86db876bc1d94c123b72aa7f8cbbd3e0d
z1a51253f1817ee5847d2c49d7561c3aca48be027881f755a2c3491e6507776e4eb8a7008bf1338
z43f81b17ce880865e96c30cc8122508ef267d0a9603bd5e8fa274d41b1c32f5d2f7d7cb95b07c9
z470fc0b5782a6e5e74660eddc6262062408a90ca5f1e8e92a8ee63855a777de6c762e5d1ebd8a3
zdf34aba9a5aa6c5905431a0a323559d281e14be3623379d087f6e81a571b6e10a02cc98c225f33
zc0cf975df18d54a09b1c1b1bdacf448124447736125e844f6fa903aa74e122b3a1d549663f4c94
zc07dc955f66c6ca37e24c537f530f1eda9b9bfe49017d14f4e8d3838f7bdaccbd79ac488b10476
z395c4896bbcaab6b1a948ce627e898ca3009838b57ec83f932eecabb5ac90029d457386e282547
z3038d8b27c41c1ef12f6bb3778f3aefa543006da55c788a27b182a065a7dd2d8600b1d3a31e36f
ze248f8e89d37cd1350f176e93b0d13f1dd9e0a8e3bedecc18ecaddde1aec0ecc5b4b73fda28208
zedcd4ebaca6ee96ce48f94a65eb49569fd4f539d0c9943b8663e906520db5dd44d595df7b06564
z47886d8628c606509c123e541288694680bb4015cbed20773c38a5ba2439eb464cb70e1159ff80
zad10fb2649165b14ecc0130147201c719c51c14e92e81a7362fe57af5ae89cbf771969eea66abb
z6617256850e6744182399ee3a3faa380b5c836bd20e37bb7733d549364a229fdfa4dc26dca85ca
z28d4a77cc2e08b911bac83a45e5cfcb9485043e71f351709a0afe6367d38f96aba14acdc0756d5
z68dd5187d512b8778645b81a5a78a9de73607e37db7b851dccef644937056a9bf73b9f9313c932
z3b6cedc8332a877ff5824cf3bb986969d49ff019c77ac5e3bb9dbe3002162fb78349fbbdfe19dd
z3a69976fdf529f864c691f1e295caa42f1e9a6f9555c941127de33b4e54bd66138e9b2d2271358
za74f99fc658b73ccf3fe8aed36ec1669de7ce36cdda7c689ab78bdbdef2d9ff75c4ba8937ddde5
z4e9067cda77c7d7cb555ae274cc6940e2b3281b3450b2e8aba49077e68713c6fd1e8c8b7084484
z278d5a565ffed2d897ebc52dc1b5e7c11e025084d464bf3ab7ae78d57c5f7cdc54411c5a4da25e
z4b59118a331bfdb407a07050244c913fbcc03d9d57b1cf2d55700eb923f217be1b4e9314422530
z56e728be585d0a88126cf8ae53c0285ff65e9b5684881e369150795be6616b372fbe0de3effb88
zae2cba54287926856808fa4cc26a60d43114c4db8d011d1e9e29c2748fab86e1b0a9b8dbfe4338
z3e3e08f3ef97f26393584d2ca2bcf0cb7b32379139d8e11517a18b579afe051378e0eb5790924e
zd97e5f1c355102e1672556149e0469d53234bd5548d1ba04d0be7bf637274b2d14ac58bb2e63a4
zcd23e0e98646362d50812f1481b92d63d6cf664588f087210c538290e419252056276d09f275d1
z3e9ccfc6c6defc2c75ac771b4415490b9ecb63229338ead832733fbb73e0ec0a2449561f886db2
z8bda2ff81c4059bc9a9221200a33323d28c7c7712d6969fbffea291ac577d4b31457f4417c0541
zd07f3a71b2a0b03bc30affed9c9b7c7d5294d589ae3bbaabbf76efaddeed0544d92f4eb3c330c1
z9a4ff9b0d44f61162fd74941ea2672f542e8ebfdc7764cdcfeea172c370e163dd54c849404724f
z9a0ea810341ac15bfda9ba234dace2635dd0efadca747ef11c83f6dfb962930805e14d421e3ee1
z02c6cc4d7af7d3003efadcd57af58e68a8c8c03eb98af7a9d9f67d25639661b6eb07f9d793a092
z5645770ce3ab4972c54823872d4eb2da18b03a96d05c62fe96c188402f7349aa8ea51db94d1f96
z9dfb71a40b03657991bc06e36650198bf61c800378ce3611bbd1e0a39a41d24c7643e37521ee2e
zccb0193e19efc4c471f856d566336a919e9049b8807e6ff89325c76a0e34a2356ba595f8fd191d
zaa4c069c49eb0b5e04e5cc095ddd2ce25fff0ef1999cfe44f54134915302bfe54640bbb1cc1498
zc332f34beb6126ba45db6c99adc0d58e6882a743f03268f1351590e2af4c5d5e5b0f096fa90eed
zda63764f63517c527f791dc55caf50a4819becd435f08a286b4a4d09678bed68c604298678d585
z8df60e8aded257673490cc779075b55ffb33c874e5f52b2ac3839607b6efab2f9ff1cf721ce96a
z7ec6c7aeba7f860876fa814847fe491407bd90590355a5e7b2e7bb1f24603032dbd70bc4060c9f
zf0359afcd8e2693503c111bb52848cc3d79fc82e41a735681a76fe3ef18cf3abc4ff2ddb7cf9b1
zf1a31c7335f1e2062e17ee7cf6d7a2622942ea4474cda0cb4b785a514fe50b11f2ebd9c954f206
z3ad706d022f16c908adfb86f1cafe84292c6bdd879a979bf3139ab6ed9d2171254f9d96ecd15c6
z2efde4b820934a92efbd0a4115bca899e66bc91649ea84c173dadde2bcdac5380f59475cff4076
z03a8eb62a831fab731a485dd6d432d4d8e5ca4658f85d1cb0ff96908f05c05335c0ca37495e1e2
z7bdaa0a112942f7f670b4999442cabd07d6721a45f6ac13ca44286d4a184d9874608792491414e
zcb8fe7763a018a0c01741fc96f713c690575586b0a7e1ab250e8cf235773a39f4b81ae51b66c4e
zf30e43316205fb9c06c3c66889729a5a8cda8b516f296d7959ba58ee798201bdb2d9eb64d85d54
z3a5558d725fb1cf6d20995b471ee2f6f6b11e08f44a5fc8611612a799ab887aac5f3e7e108c8c8
zae98b6c1d1e13625e8e5e901f409ee49d5152a71d606ba96edc0239eeb3a2c6a5b14a46bf66fb5
za5543483db2fca70454db857f5c8ce660db56e7bc74bb837c5f24df87de149f280ff435723a251
z18fb70e4cb539a09d1b3bad6452fde478ec4947f2dff6655d7abc7ca876329185427fb5b8ac2c9
z09aca4a1bc6d6bb5dd4e33f017af3089aac1af664d9c19e4d7f173ee0cd8500efac2ef4cb421c7
z700d85177aba1415e3efb883085ebf8d223b4407fceacaee40de48d0424b0654ba5e631d203dc5
z78a230e6b43d0ab4fbec7306a39b4427af75e3522f62b7753c04379df20001e7bb946f2660a3dc
z82990a29b8d162f822f0a38aa7d260270a027c500e03f91e1a45b85909b96cd61732df2c880344
z543bfdb7d08e52883c6f87034363bb4c38256e1d492d85d9db042a78327e18a2ed49eaac3fde23
za9f65019e38f2ca3baca7e909e14857a124341d1f31327fb973e7c484e01fa2fcd8353f61365ea
z9f9690cdd87483f1bdfcef2558287af8f9a69daf86f771de0ed1ec1cf49ceacb65c4316ab75fa6
zae51f3cedbbe15e76257cd23d520b8dfb96ee2178f16d2f441ddee4be2bb437497c974d44bede2
z7b7b1b312797717603dee62bb55bc0a48386315d3c23fec3ed23f4fec09d6371ecc8a5917ce4b8
z43f4767482a6c3a64c267e0ee8e990ee75ac5f49012664b612a42fee409f80d9b9bfd3fede0a3c
z6a791b9fe8bbde23a65ad50e5f561ad55cd58103b0de8929000636e431f94eb7979b9d67549f06
zd1045b485534903ad45e2440c07cc879ce61c6f16f6b23856d9fdc9b65689a96d40117754b9614
zd249dbc998726aa28a7aef25eb9935b60b7cbb0389bdb60c7d23f5f9be621c810bd9f7d1457022
z3c186edca5500f1bda0055026e687ea947efa76e4ae7c36427053efe467f635125f3d31d95b749
z27824a553994f4cf2e3a09c93424cdfda363ad99e94b662807165d85642d5073dbc69dba4d09cf
z9dc7b525a6414c6e3fd3e8d91013b5f614fd6442af373cf44ab2d27ae7b1dccffa591c25854e23
z697b7f2fcb5fa1fb74bc50e1dbab67a2b2986196d38e25750afe7a803dd0494ef3891d5e0e17a2
zf1c82de45100542931044284c579bbcf8d0df23f743fb25caafc50c517c2eb33384c21655e987d
zc207690ad484962ae2d53920df4db4a1e4f6b9c0ee00d0a162a3c83e5197c0a4c99de25ee56378
zf3865dd677125a1ee09f404000480fa074ff6dce9e1d98e3f38d4bb628b2c6a537f679bbba4e26
z2083b015830c2416ea9be48317f6bbc9276eb08cc319494d70d062b84e919441d403ee481e51b3
z24a0949967146c2c812413c3bafe3c23d7569ed7cb660b439e82061658aeef74f26ad5e042198b
z09374000e95e5fa79b630a71b021d5774ebba431110a6763ebc302d40385350efe5412e8e4186f
z00bb256894a118b4ba9396e384c1c78cad743bed7c50ce3c43aea1822e209fad3207e056c735a2
z82e3315094f14902fc66e8d3e0b896f725f91f89544a592447dbc852df7fecfed936cbeb8bdcd8
z487df3d6ccdb3032e878a8b10d164a110c80cf51a603aa6e6d767c01ded112b03086bb113ae5df
zff8449251118b64152007fa732aa801f7b81ce00b0f09874ad6b68f0d9967367c50d61a3cb07d5
z77bf364a27d04ef385f858128e4ed353f09d644286cc3140c63ddeed1d6184e908b1426820dd88
z3d2098f77ba384b59955ebac2b41d506866724c972eda3defd2a2cbf0352d54f02568c24a747b1
z52be6ba1514898ff4ab2fcb0e3a4ef177e0618de463556eb1a6968ecd67a393086180e12de3bcc
zda79442f3bf7d60c5917cc9fea8d49d8945459890134959c9999eea1ae19982504429469afeba7
z6d61cbb5ff587f6f6d4f81dc1aae8c94c0e41d66765ce9d8d308ea7360960a24006ed7fc7390de
z5305c10dd74128fe0358d8fd2bb3f64aaa465a6f41fd686e8dc9f36adbdf0d8439d9a6261189c8
z46ac5f6161690d6eefeb7be44805ce9ffa602cbb1b6dd04010eb5e9befd557898001c72e7f96e2
zbe344172fa308a76d5856aa1435d960bda9073c62a17a55e5a44bc1f460367f021642bd856f763
z7570b0f01df5b0ecc3a5fe1e7312e5fbfdd5ba41428238cb06bc6e817e5ae9af801b9bdc21cd1d
z02d9680225b7812debcd14a88374896eb26ef7e087959f8044deb2cae816654b250606fe561a1f
zc119b2a1c0deb4ead79735821eed7c5befa3ba6ddd43186ceedbd471c31e4186d5d1c9238f767e
zd1541f1171a660421a8dcc69138afe753a1d84e366179911d3229db2467a8cc567ea92737c2559
z62f1c29ba7ed73908060e2c8972b6677c9cfdb10d3efc6f61c808828b5a3c8240776a7fd1c49e1
z51a3730804e46ab062aef87a1a307b7ec2272477d881fe802639d5a83dd1d33452a35b064f16d6
zab76ea6ac9716a9d0aded090eed43c10af214fdf9fea140ddd925794eac550234df7e974ba126f
z7cff396075d60e7af8b2148dabd7f0afd1a43a9b679ff9e761b9d672d7a0be0b422f546546ac3d
zfdb1297ff10c1cba81d7031884de5f9194f5e16065e5ccadefe52956756f4506914bf0f1f6bffe
z3398a55f288fb7685c61cd128b12afbf88783f11cd8e8350da6c1c070490614f15e868c445ab4c
zf50faa0400bb6c2978a4df9ba4413d24674c7697bbb4ac1b9330a46b663cf81fbb169a9001d7ba
z45dc8f37a7c6781fff6d2fb9b08f813c3b32b6e49f06899fa287a02ec025a43845f3740246e9b5
z4542f5d22d7999def0a9ad769b175af3f346fac40e42ec8fbc11b26f9bba544820e1f9957725ae
zd5d45befd867b6f901c0c0d5bcd24ae0df87eec58fe268a2908d99010cf97f94abcd6419ee7a0e
z67fba587ca26d2c1413786da9d3a79bb0843983f02c3e68d090338dcad28d869c720f110a0cc4f
z4c834f30898f597c7da616e0c33d3b374ef923853546965ca20e002abad0b5b09cb18f8a9dee65
zf8a04ad590bf3de96276d36ac343a6253a54f730445bb9ebabe3ba88bddfaf40766a0f10566a80
z0eef6a072c98830515fe685c35d833008826ecc4efd9e8113aaa4ef16a643c96ec41c5763c6f60
z51897cba181cdf8cdfb13104de1f2e763423bc0d73af4621ce433248fab8463eca075ee847c35e
z9a7fcd83b048ea2db13617ef06fff6d75b7470d6961163d677f990ac5efa04d81b51ffb2449d14
zdb0a675e62bad1b5fc251b49e0cd19f3b3809af9f3312482fd782b18f459b7536c7a892dbd29e7
ze80f05b4594ccb958da276da8c3462d3902b0e3428ffabed41008f6ad5261d6e79e9ed180f4419
z59b75abe62ff16e9afed95d14144984957436bcb40beac5c301c4e98f95fdbdc01329d7c77ccf3
zc4d8ed571201de09f5d98b9a1a25fa2f6d2563ef517473c1f8eb1cc9c9935d50d4140980eb8811
zabbb2cd5095dc55a3d8fd6d70fdb620b33b2062d3cb45e44430671d9f70ad63995f270e0a5dd0f
z80323a67c84f2f613aa74587a8e0074bb6c78483a91ea10006d9b0ab3d6f026c74577686892e56
z7ac8309dab82980a3015f58bfd5c702c62eeccd6aa3a35179eac11a5661ff4618b184a21aa4dba
z2e4d41d6cae7efd5f1a370284be4b3e0259843242f475dcad7c8d6afbf2d835424786b44195606
zf469ebff9249686a6ab084a1c15d67c5251f07a360daaa412dbd425f67520d5d05cc6f38d41e3b
z4fd40007012aefdf4069b6ee4fef379ccbb97fd81cad09e77d659275152861cf07dfb78b293786
zc5002fd60642acb580fdc0af51eec760bb3f0f359ddce7c5fb5e445fbd7f07f22108e2c061c3be
zacfd68fdf51bccd7b59625c0b679e2773bc6e0495a165e519664d107b157cf1c53c63c87dc7a46
z29c69029d7b0122165294b0477c76aaf3074f6156ff4e5ac29703e25b473cb27693a1371bd1ec8
za1794c9794e61cb1cafbc1becf1d774064f01e7913f2c98e0d09c938dfee0a80bb50519bce4da7
z597d0194ae299e83b478335cecefad4ba41833fe74974f37a0d6d289bbe51f6c4e66afbe9596e1
z9dfbfa2f953cb3f9cb160a381efb5dd7d4f46e459ba9deac8c2cd8886369978ae7d262aac7d643
z623277390ea3f52726634e457f6671de67e626510a687e230d5fdb3afeaf76a20a81a01d5c2f4e
za53a2b1656f45a03081d5a3af799b9dd460663665e6e7b777bc2094a6556b30bb93ec30181d050
z19f6a7f3c0b3cdb0fc34789e60ae64dcbdfe5be746ec01150b4e71f8f7b91098924ea9f78ebb9d
z852359017170071c4c70a08426f5ed20afc1d57743ef3cc4c55b5d79982320cc53193c74bc4bcc
zb758f63df166e77706d16d91092dc12f3d47aa2006b0080d1a016bfbac6384fd45b0fabd546063
z970ab68476af2f68c06552d518b46b0727e007638a5e4abc8e560ecd3b593ac8a533d38fb88649
zab0aacf14c8eca645f9d941288b1225139aac942ff993c9b153204e60610c57a43724621923fd0
zd5239da33bbe5555b6a072a3a74f4a16647810a0b3c67b61a42d6b79944036d949cb71cfacdb3e
zd77a9f7edc9eb1b6f9a9b9d3d5c3ebe081b14598cbe93211bb3ff6ac3cf36a362c60188028098d
z63477c482bf237610ce6423171676e0ca88731d53fbf3a2b3e2e7fcfe4631b48039228a9eee279
zbe9a68a9796a54992933d35560d874ee82da1f7ff7d13257c628e21dbac7363c765aa73ad07796
z9a428358bdb3bcc55e4a1d9936a4ec2d49bf8531d47a46a7e40a055acee2b38c4e9c469d0d3188
z8f489eef59f21934d802fdae4bf0683074ab1f46d2c3e71cf87473852dc933b49c65d82203f84e
zfaf415a6bab630f9cef5ae2f7138bb00e32975c94e6224b6e74a08381f1068cde5496ada3a947d
z75df649430035aba6186233d5112cf34651e2caeb20f50299db65b773c687b9a47093e59be56f0
z52841b29d10ded13f9334a69712b520225910ff5f9fd5c953d5ff93dfc216e3b12862bbea0d3a9
z91081864098fbd5af437d8d198ff2de32ea100631ce2ba5a89d5039a3f69374a30a9d155f6dcde
z7f2d689accd13b171e95462ce30ac702e44edbf062cf3e0c1d231fde0c6b31213b433ba24865d2
zedc3e9a3d08b8fad7cf56e30497f95396f54f808f0d4c4600479dd6401fb38870ae55d96b866d9
z7492cfd5145c238a16923d9224d43c3e79f81506744dee0da95f7444c04e469adec5e67f55509a
z4bf9d1fe91f1500d98a3831842c96c3bf3215fa8320b9bf0d7e1c74c7fc20f731a3443c542900a
z4668a9ae1e34dda65a18ce4ef5dfd59b6927180d81bd8f5f966b045898eecddcf919516909923b
z17fc218cecfa217a27768ce1eb8fa941e7914391afbbd9b082295a4ccfacbbb879d6671b6649d0
zec1b061ab7cc341e3818e3a25c954a7a7236c8ccb68c2770bada0b4912d6c8b3610d5ac32510d6
zaf36f6909be42cbe66c93c0b49c66bced798e751141681b3007f1db7ebb0f36f096c14a64ddab1
z37b8e966408b1bbcb387a736e5983dd5b1f5b8dbea1a0992e719f3c71002e07a7f60ffc4a9a095
z0222c8143098b4941b5f21fa506b73745bda78a47d0de7581e289f87c7465de0b80df2afb212d8
z68bd2d6d014c0d1f2e38a089330e187f577e8956accaf59e32646ff1aec608458da0efe4c99c29
z323644e5ee2cf328ce21e81ca754e21af5dd4968c109baddc8da06049f5817cd8ef7bca345b302
z70e1f58d36bc911760072100c44534edf6ac69f736bfddf3b14a94314049bcf9f84b69bcd6d32d
z1e5022d54da040461a29e4ef185028ba1d390a0f71d6d7e9894b20eeeb9bdc95397d048e7754f9
z669646c71d553083051297fa819554cb285f1690d22f939d8d4b0ad73a2117aa6127a5437baaa5
z2cf3a84d9821f115449debf518db82c9f645789cebeebf1d1c657d7bce3418a2ac7e6648f09a31
z59a9d5cbc5a739a6a8ffa507626fbade83c5b045895fc8f0a25308f34a6b9a350b39a0c0aa3842
zfbb564385d4bc2258caacba5eac0c8dfff88ab29be173aec88226947b259459e07082c1b010803
z57fb824a8085616caea2dc2a63a0c7b03a8968eaf18e068f8f9a763612fc1f974591169c860a53
z0a3f9d4b60f4b48ef110386e0a1b697f6ef9da3daf4a4046b14c2e79f7286143c4d31aad581a80
zadb30eb9928e3ab93efd8e4c0b4cecb433f4a0e2b4599d9b3e83ce694c14ef57b8aaffd5a6d80d
z00bf46145ae6a2648914a4c9ca9758f68947f3187f20f7ab2f98a2b628a5b6a9ca129d04a917ff
z1bd4c698d042ce665d3629ed7ca60926726ee56b12e02e6df1d53d1f6ec1d6019fedb30f73786c
z229d9c31dc961077fc922f46511800b5a167a78639b5ed38d69874c961fa8671d89d0e4f6a96a7
zf4250f2bbc0f1cbf063c4033d53cc5d1a32fbc5ae5056cf34e2326b0f1ad9f20dbd62709863210
zda81ca857cc4032019a60ced339f8745d02e8ec9f9926a11c89cd17b2697d3400ebcb41df84a2a
zd8ae33a2b6fb27841f39e6085a81962aebce6b209503625677427eaa7d1437e96f0b1c990fccf9
z0d47aeb8d690b00850107a064fc6b00d53f730241565826508d3b55abb7eadf588f7d97ec23e29
z152571eec49e76d5696b3cf4f50bcbe03713a11f4a4480290ed2d661f2f1ba8d37b1929be7ab84
z848e53f583af267ed1e8287e7cdf2c4b944bd13e86c3851fe62fb3aa5ca0f05882f7709a1a7017
z826ad0f5598e3217aa8a10af6659ee94c0d6dcae36984bfb2cb09902493e61d559c67a68eef438
z852f4aadf1bbcede996306bdf426a3d7037f8702e364c9ffe65a680e4464e23f168ad1432cc50c
z74b4b52538c04b87b5bb2460d18d85aca4ded1d6685841319f08038759915e3897a66bacb39437
zc8dc65b6d7d2fb1796b0a086e3823264ecf58357dbf6fdfe3ddab0fe733703c8503141c4ab407b
z79cea162859f9c904f0c68eb1e1b57e5ad1c062d0f3a9b74d2cb65a376b2ceb26831743a82836a
z98517bf78e96eda6e27febad7e967ce1e914c1466d73b07bebd0a4ffd9b1ef1207788731a19c40
zca56eea6c1d28ce892939100de8ff37425454a95aaaaef083162259516311029337b3d7b4478f9
z1dafe5fc2d7139ae400625903fa79eb366de6c6af529051ac3c4c07b44f5eb805078f33980c001
z64b8e9ed85d5929e2d9308a73691a8909a2074d652679f44d1c2c2334d5a4533d185f45f1ca45b
zab231351b61073021e81cd9ce4db3f5b6134af5ded7ca4ba3fd6a75d4935f82adf194288efb96e
z642ab99bfd84e795a894d9f27d1327ace91babe35345c65a0c99633c8b533ad6bc81144cab88b0
zf564aca83bdb493e9b3c9c7c280f5b63dab72826b68e49553fe7b8a97da62305e8ea90a1587245
z4d01e51e4eda39e875ba0577005a3328c810550153d0c60b2707f9d5e7b22b46809f43fff1077d
ze0be67a181767fbba40b6b9e82a59fd8040252fa0f8ebbcf9ef1d962946970d8b2637b92fb3128
z3f44bf77e8b95fd11b6c5f62caae4ad64943348a2cf825e49095a07daec6ae750a3a7cb369b454
zd5080b524d191e4d1a4a151d2d56b63a572460e5302f51dd6d820b06309f2bfc3144e7d2f176a8
z4482be4bd383d1c938670959c4f2af17e8f7f9a7610d313a03c0d4312ca7cdf0212bae28b45ece
z0a0bf5dabde7e71bc601f118177773322ba5e240de65f3aff1c1024d8102eeac5bd182ce4e0e51
z7c64c88b48e4da20a0a3dbae78e136003ceec5677940ffd02d6a4136f91d1ed3ae96ac2cf4817d
z97b400724796ea457195cd11b51a4882f7e94c45998fe0889b26771884da704a48afe7fe802a2c
z2774d83955b2cb6316ef20a3eb26139f4ed950a2eeffb621aa6d3a1cd7687c0624801faadf0c4b
z28f147de15481470551ec3f0a00a23e5f7e1ef86ba98d2ae0709e9d80eb61e4dfba606e707e77e
zf60e8e3dbef3fca2c5503abd496f4a9f06a02adad681b2aa50b57cffd6261035ed459ce9edbc2e
z496a26f27cb04e8e471ebcb8e3dd3d900a280d574da5fe081e749471862db3fc2272c327d65436
zc1e33b2b767ed8f8b923fbbd10637031f41c2583ec756624410affcb9739432ef11b6a2537a999
z339366caebb4137bbaafa8f39f989dae738eb5222e313af1498f401c11f6672bd607b25b3f9b69
z33cfa66f7a0b17b34ea9cf81274ce2f83afd4d7879d271fea2fcf5b58fa6b01f5629cba87c35a7
z0d95074fe5064d0aedab58cff9da6e0b26cbbeb70867ff54df4a2bc5d2d6709509ba297b4b1d12
z3237be1192ea275d1a4ec1708f3eaecfa841d2503f92a4b83acc24ae18e8ae1403a35db7751ad8
z27a0acf2366153e12f7c118c64d4dad7d2178a0bb2590df8f267b9a420b2e9187ca62c593fa787
z13d26d3d65a757b0aaffb44311ac381d4cb3975a29e1b3fafe509c763eec850fff70e14e6deccf
z559aea2c649a57c9ad871bf7267c62745b7f5dff0f59bb1be90008f37ed08c778280dab3411adf
zd974df806452f43d1c276934224d24760dda82416c206dee3e10fc486d8056fd3108095b73587a
z7a9dec7f125535b459d6f7f744bbecd6f928b4dd8beb391fe95a06322956dc707aec773b44ca55
z6242e5c047788283ebcff9afa562755359b9dda2db6a7ef4b033d8e47af4525cbce8dc077e19ad
zca903cde0801801c225e4895a6eeb4e8451822a3ca2bf7b2d04236a243166bdad026b40370f8dd
z0cab9170420cae3a630035f5d3d108f233fac80e1cb18c5df86d481afafe086422f1bd9423cea8
z2a4916c764e581f4a618a48d77a411c0490ed8a1c1c238a4ffed4c6ed455d92efd925948f9fe83
z61552d451f4561557c11346b76360fff13f55438f7a5a62107cc859467ab7c3b125633b763d49d
z5d92cda4a42ba758b461107b7c85e2d107e4d8314629dd18ba20950900ee2eed4196e850a99487
z7a1b6f3abdf60065a55085883a76cd717ecff7f6b34974d498339380a2560af8fdb95ff4110447
za0f221b5c2710365c9a8a0628e00dc907ceba57936666a2e950f0c596b5795b1f01850bd138fc3
z219d65de73106feb6ca6b1c55c315042d86ef57becf52890621df68c4d0e0401e3d9c5287c4b30
zb53eb5f679a40dee85572db7da01aede9e5595347d68eb462064763b3348b96181c1ed64ddbf46
zfac870e972815e149bfb01293b5f0d3dab9d753f995879caa92bc9d1b8a9458a5f65cbbc96167c
z587ec722437a294a9640b9a7e18c789db291cb6646c7023223a115c5136a2241a2b171fb91ee79
z713b96131bf82af29e294075910693fa4e360a8702e655a802124b0d4b147f1595be04b420b734
z11b4de513524cae5a1918ab5d240b76b1a7a197f5aa9ed52a430aab5ccb564bfb7646f7e1cb2c7
z284ed85b10cf15c00ebd1e4215b3038cded22f55a1d84cff82f1d6ff53463cfdf5e04e918af2bc
zf4b28a814eb42db5ec592811a1fb17012c43e0f7dc9bb93862233d02c3dfa2fdbcce2d36b2863f
zfdb34fe029cd685a0efe6184bb3440fe5b4a9a9468aebf63fd31e762258bdb214d6277c395948a
z15297b061e1c7e15d6c65bbe67393ba5f404f6a30ce08771066b0e102a2465df7e6f738d46d5d5
za0587c7fa5605570ffcbe3c438b400cceaae5cae077f55bde407ef350ac7d4f78a9437f97cebeb
zd842c09334c72414f53c07d0a44028c3115e58145764e504abf53818c9e8143da106d28c7a0c87
zf0e3c25a80f86491f4ab330d022ffa9b2d42ffcd167db44ae8dd02e48e88816a31cecd389e3c55
zda7a99cef0fb6b2af85af67bae1452214fe2956fe68318fcfd5e14cc1de7e9adb7f9888c8d1e8a
z506633fc6c5595012fd774a69d9bdac990e710393dc49ec6b22765dc696eaa65c170706842db65
z066aa93584d06fb4554cb31a715bafd300c312c10c4e914fce0d7d83c6f4c70ac1ffbd952b3cf6
zd3f8e77a232409250b7ee178888cceca02812cd818d0c9098626532fe2f41997db68d255a5c370
zd12c35e8b82df092b499109ec2b60b071a2cad7c6c04aaa205de8bc298df3685e9509907853d34
zcefad18e9c8a5939982299700ec094d27cac8e44609ed7c1b1b9eeae31717b67bcce642434260b
zaf83cd994102f0115b7a79f00774fe69072271f6fe9350904e694e619ef319ebf804c22bc37e1d
zcb84632013250d77ae35f108f1f4270b1e9dab9d475a7750a3716315870fda92e8be046365dc05
z5a7e79ef8908433b0c7d137a1ba7f6a1aedbf55692ff7a24dba6655beaa9da622a102eea7923b9
zdd32f706e98d342d9033bbf07f33253398741b0d5e5be237c24b0ebb09bafde68294ab250016d1
zee071d6f1f46a5a8e1897b0d8364c82231948ab902873d4fcdaee6c304d6c74543999da1fa656e
z1c0867d84d15ae2ea8d9324899ba05f0621196f9dac19333b1426e1161aa56ef73c2abbf20bbed
z7d4b598c61f9076928f8140d2e50af89d5321429af6532a359b713b7bba22dda34f8c6d3e7857e
z2eb93bdee2b922fde9dffd90e8ed4aeccb061b8b332485d8a0418de14581429f1791d7967599a8
z8f1c5be97a316bb20ef912b70a89ea88431adc54070797fd4df5034c8216234d7fca86f794be86
ze4f1d74989e78fa677d2db9c9dfd04d92cf1e6253b499685602de86f3e88ba752b6ee8a3388db4
z4f93864eb4bfc70efde464a8ee5990f0a8061e95195155a2815acf873a995c8f8e5a17dd96ce80
z5865fddd6c61200d0b2a3524c737d3468ba7a021a55896548193ef0801aa97bc3fa06c8dd99cf3
ze8c006453248feef7e553deebf32a4ff3e02b554d0d85790281ab187ffe19101a28cd433a7f3ee
z0c127c91a89ed98f01a87a8f48d8e43bc3a5edefdd55d302b0a5dbb331901f27915371a7c80a6c
z9fde2f203a5505958920454249b7a94bb0114c3fb7bb8b05a97b7102bfbf111a6c8007648a0511
zff2353230a16f8724a61e28305175e17b1c436d2ddbc642595bc04a4bb4f20e01fc186977f4e04
z38f1693e0aba4265d49f83c02b006d20e48c2a963e25e6131e9e527f19052242ceb578d674a6a4
z1bd1502ef7d13a47983a9afa750aac8185a98d82ea30e5ceb26815ca69feaee13f82cdf4169357
zbf9e5988d309f30c7adaa6dbd36bec72ffd525f398704fd1f2f47aab16ccf2895c46e982341216
z76e0dee426aef663d688c5031b7a19a75e9298ca84b6f048dc8fe5d78227a2b6118f8a86af078a
ze1bdb44b5ac28f83b26f851d8c24df31b7fa44bd8b6e5e98b1faa149bad3a5480914e9f5c587e2
zbd49fb84abdaa884ae79509c92c6df4c3e99517e0d040bc05e9097ba67938bed65ada8def24142
z4413d2bc442d2476e5849eb4f3a1a33877783ac52901d8610f7a94dc5639525ac594ebd2fe0d68
z09684092834faf0e14d764d7cc0743ade4aae5d905d61232d2216e61b708ef338521a39377e65c
z1974527ec34de67b8234d2197991c021ac69ebc5b96d50c790fff9d1b57b4984bd35603f307c06
zaf47921755539a34354601eae340b6bcb8c526674a6e038cb36b3dc8c769eebb595fe8543fc17e
z8ea103037d3d6a945231b2380d96a73e37cd792926a381e9c7da8a8e0e041147462613a3ec9c2d
zf5dcd036ef02059c85d633a1f171a0e5a5298f633a7a6f5a470154e6f81481e610452e7f5f085b
za790acfbb9cfb56f207c572a1eeb3b9bd2d37eeb4dd10192e8a63ad866d1d4fd546dcbe1b929ea
z4cc2fcbe443e61b3790267652afcb7b26b3670e6845903f942c10a17c5e44c9712075979b38dee
zf19fb4474bf4baf0e63cb95653d6799109ac8af16c0aee675af6d704a05ecc9a1fc521bb9442be
zf7e2011ba02b831bad1cfc9442ee87aafdb921ff6594cc1ab1a726fd1d18f2f86b000b75e22303
z8540ad4ac2266a40d6a45227834eed007726eed0ff40de1ff13f1449a8796809de24745c873c3f
z0f56c5e5c33793a80a6df244eb2538441c2aeb40df4a1b284b58493adc7a4ec4e4746988f06fb5
zaaca160a355572101951b2ebf866d0e19245a93143457a288f6c820603f80b8ed64a20165f1e5f
zb32ed45ea58add506f55951024b2f1440c97d1d64c3fc3d32ae26b4eb466c2bb3945b35aa00c32
z51cac151e1f58448661c5e8bad9a9510aeed83c1b393141b5707351ba40c05db6018c9ec259393
z1e1487ea70522c1166ab5e94297754e8bfb8793076bc45232bd3fa573cfd4e5f33137e2f4b7b73
za043ad7068c970f54557204d1f8a5aa51b77903444d63a7bfd993f0c6182c71d0a9314fe9d4325
z84c94bea9cdb26883adeeb7fe659b0a29f4103fc7d6e990f50e19a6bdda490e77c0f50e562f6ec
z3037a4dda12d09d27e4d644cf612f7ecc464bf5a68ad3065569439986aba9e1ac84eb60b7d75b7
z23e64899448530fbdfc5cde82722e41e54939fad1021ebb24b6caa83d23f983663415c9400207f
z86b163f44a254a0aae401c5b4c44a026e56d3f6a1f4d4af501be9ed0b900061092bcb31fce79bd
z018c47a098e1a4a308970533a4471926f79af2545ecbf0520e1f86104c28fd86e50f9ea4a175b4
zf7f392e51de54c897051161a949867ecedb4f2748a52f97f07444bef26ec427bbb183502782757
z72e17aeca538e59feb46bdbf6cb3694a535c6a3faba2fb4818a10e3f5f8ccdfacaea13c098077f
z68282df5a67e66b6391558b9480d4e9726ae23f3bd5463031e610aa39aed45ef3c6d10768eb6f4
z5b6816561dd9f899db5b13b128f6983befdafa2593ae5e144fa7a2543a910fae1f2fb86e11ac88
ze5509a91ab543efd6228ae7174be7c1e745a3e328ca09c7276dd38bfd0f4c3c984c2e08e4caf8c
z37132c5b1ff8da4dc7480d212b6b5634c8cf4b9a55fb0034daedabc1f0be9ce9902f82a9756727
z6625fc2e7048cdc191c9a74a937a7990e32ad2b9fb0be053784cb5a2c02ac108559eff55be6b0a
z1eca60585b89f90f04f83e2ec94391fc9a90b5ad07c5be9bc44e63d2341f6f0df49bc82a070e86
z2c4c845a0239306d040098436c041ef98d4267a3556946b2671d13c25bd27c72a74f65574dc291
z6eaca93d808e3c43d45b512160179ab19540dd60894ee2cf84911e01304a8a86ccc9cece56018d
z3266f39f4c403e5c16807ee2a86a550474c0bddd66295d54144341abbf5c6eb9929bbf30bb7652
zb253eec4afdf0ed951ce6909e5cca79a7056ea0362982c0601bc5364786ff754414554cc2d7cfa
zd5712330880f063924c41890f13e99574665e54905c94f055e7c646c7f5c2ddbf8f9cfc36d5dbb
z11a56953ac2a02b41db60999b3bd254ea244e559e3560fa0dd0c99677e4ceb20eaadb615cb4ace
z053601f0a9adce57f00a5c33be0369982e87ea3e5c702f34aae07206e651da5c165a0f1da9da5c
z5cbe93d197c205443aa70148bad0982b36bcf69f3d862302a0454bb948e081df3d230d0e58ddff
z75062108859aad0eae3c8be0f3a61d2e426ff82bebb3d981107526056e5956f9bad1f30a7fef4b
zc80c6667894f9023331b12b337d2a0a8e4b0a9b6dcbbffd9938d11308ee6d3d82c501d01437904
z3e19b204ea59564736f6994426dc67587f89ca6df86762e18abf04ec340fe36c142fad81d2d3c5
z9dc3792a6ab555716c19b92fff732e7ede809811e80becb42fefee3015fab59f44d8187055b910
z54a540c07d97b09e7292a34857ba16d8d453a72544981b76fef91343d6db7d7419167495d6341d
z926474c2244593a7da38c3b39676cbe72c71ae71b3e8a341d54c651b96d492c2d1ecf36e4a8e7f
zb344d50746f25b3f8c30b76149ef92fffd791f2d325640e960a6037ad3e44d4e431483532357fb
z5a43796e8ccbd0026dda0bb28ab56e190f157ab37eb68f53383ffb9008adbbf191a9bf4cdf9625
za2525b52eef32f1486c4d3838177ebcd204a3db55cef3fb8acef951482783df07ddfc6d0e330c8
z0abb092b4f2904e757cdebf3fef5b074cd06a79b1ef5d0015eb209136979967b6670f0a106ef66
z4263ea6f54ac926a0249faabbd34d534f3ad0673a2170ceefea6e6b19cdd5615d7ce98989754ab
z97d80b8f3679925ce3b1a8c210d4e0687ca5f8cb726d8beb702dd2778320c6c10fc413300e9fa7
zddc662d4c4336cb77d0809e5b2c426acd50b5650261127d2b480c9735c76ce71262079aed36a1b
zf4239e611b8f18ab600df9466078b5c5757beb6d26365fcfb4d20d1dedf383f5baf31c6f1b1a26
z9b602e333ca4ad6f13392a41957e8156de6ed5b54bd280a9e7a0d618fd7a3a0df81c850117ab60
zecaef98a80845220825f92311f55397bab221e0b3b49c7948f7a0c7c7d16b7828eae5f25e97129
z8117abacedfbd5f43bb748a7f9e11728dec7f8992ec8ca4ca5002af8444eb97e57e37b92ef80e4
zbcc01edbf89aaa794cee9e83463d8f8d07dbcd6360e967b727ddfd56cf1f79bfcfb58423e0ca46
z725c9b2407098b030e50fb3322876a415f999a04e5cd81c75c5ec0be36ec2635010852fe45b568
z90aeeb50b158e167d5b3ad08c4b53e8355ef0808676a73b96869eefe28ca3113b9084689551647
zeed81f1a34af59fd50671f3717f0d5c0bd4ce4315caa32d147b192e32c92510e8ecb12d301744e
z20a9c06c64ad6fb33356e0009fbae714b11eaf93077afbb681160944e462117b957ebc45cd0f68
z8757406e1a294eb64ff99d415d86a05e81f90a7afe3eba02050115e3cd56caefc5edcedbda7b6c
z02fe24510fe32ad1563052144610be753b92c953a934267f50046722a601f9a8206774e36769eb
ze0fa1bca68a160c729df256fe2c8ffd0c36d409ed09beeafb2e4d8bb4cb6c10051694fec900d3b
z4685f21c83a60243c32aa4dfa1a5cded392db2749b56ad76966cea2c6e61ff02984b19e505506b
zdd26d664d544226c118d533aa3d530cd4ac0b60798fb27ef711c8ee548d930e23378ef30192fc1
z4eac02f5627559a2307f154ee23d7166bedb63d5eb7a92955dfa4be746f6f4a77f5506badda1da
z84679f74034b647195a20123343d0ab04709716c5245a92255d9ce1746cc53f3ca553af0895e08
zef901fca5f006ed1a351574c273e705ed8d5d20e84339c592751787fed9fdca1cd0834dfd8f47c
z00fcb424fdfa615f81bc02bd4d60ed5762ba4e9686c7d74e478960e50d9ff6a9bf61afd669ee7a
z448e17c2ae6547dfc795d665d72d70ea926a3779cbb2a056098d0b87fe2463725b7e6fa51606ac
zbd4ec371b71350f7fe2f3e07359410e491a2a7de98b8f43117a39510ca134beaa3a575200245a6
z37157149c07a517ecb8b196d9c4d6ac4787c62e1af5cd95e119a065578e7db8660c5adb3ad399c
zfc9c01f1409fb1f06a02250f74d9ccff1acc0d105448213f625be087ad02f6938b7e81632369c3
zcf9a04225116ca648990549a2dc9d2c3b490b225bebb58f7d50cb37c78864cc42a7f72ab952f2a
z425a128220919f8914a24a26735e8ddb0a5f0dd2d326d0dfd52ca3c340396a0282e747ffd0fbbb
zf0fea81d5e3c7c583166013747bab5fb5f6d46015d87ec0a5328e515bd183f43c76145818de177
z921463e62e8be823717b3148b88f76b72ab281fdbf839056a7a6780b7514d0de37abc46c62a7f3
z9b3d47f1f1730b5c33c8e0dd158f37eddb521f1308a80a5987a16682b3db505df3bdf1efef23a3
z28eaf691db58bf962c1f7e7aef9fe8d268e97adbb071a724f1a9e29185161fc99bc06ef88ecbae
z4314b0934947f07dd02db4873f01791382e170dc306a76596d3c536e1b491b0d54ba9fdd59f107
z222ec0aab98b703e02bc02158d9f5a08ec09bd99e5b2a99d3f7c083369e248de8cb773318a8e0e
zc39194eac4a9b2699ee37361eea4a9be9311029c39b61f5c5e6c9b430aa075dc0c883f6c6dda86
z9b17643d9c3b325bf30f505bd46592795bd0e3e4df52040effe824cab424bccc631089a0388387
z53df332303e60e9139c024dda135d3dec88ddf5a372165fa24cfa9c26626e90f0288ac9523954f
z8f90ec31968da57f67a018258cd6b653ed176928aff7b1b86705b6fa498d2e8c46238e0bd1dfb8
z3da17d5c6ce4ec33f38e079c88aad3603ca9e4c60b0195b174c201b0fc4b81a345de9b85117488
za8a3f92835d92b1ce672f54fba0277bbf323194a2057334838c70590b159da8198793e6d28a2fc
zd9ce1c7e0c3bc617689baca66150b2dec4ac441c67bbc2ecf65e90d2d7a2167f7e16be615cd3e9
z924fc84d41d246cdb6482e951734a65798c8cb340790bbc77bbe1fcd465a7fe334ef434edc9ee8
zf5d8bce4cd312ef8c0f0503b4484e772c59b378800ac2bffbdefe905f33ed313e7cea32e91c5b4
z192e88cf750b296d2effef649d70757c4636b1917006037138013f323b55575271a711394d399e
z3e20883c3bd92118c20ef3eda37165e085a3dd1c33387dfcc7503423446ade101076908a10e2ba
zc069c41a1ecaf7f08758e472e6c624c394cf1bbf2d771df517faa2eb5995365d27a18f50ff2da4
z8a37653740449b7b6f8e2c654e2bc831d1fb15a707a2a7354132b2586f318a1784aebbf9b44f8a
zac10cb235a0336a86b713ab2dc322a410d1b756f7ec19368855d5c138a21a22cb2990ab5d7433d
z679163b3bc0d60576d714342e98da7cdc64c0e437e2ea84d3c117f958dc6a980399950b184805c
z7de4e48b9225da594800a5b38d4efafbecc172751073dc5c047843fa0c4b412bc3116f5ac2f37e
z429c6dc8f84213e395aa9e7193dba1501285bffd66a1c71e9be0f286ee95b34116a70151865fce
zd329c44d9991cd0c8e0163f3f64949fe6b50b15f47b47360ec780c9c0bae094c897030bba61f0a
z836e17d8e72964028b5382b955782bb67555b9dd8b47244b470451b9419fb1ee6b12edaba53f59
z860e439f48891f8430b36ccc5b2b770c34ca7de1e29d36ec6f1dd03d5ccd346339b6d849b054c5
z7c7d37e9fc178a46512f29c2ef871c9d6f080f7076ce3ead27afe41cb89dc4be6775cc260fe19b
z536b2fdd4e1a7628dd6f9f29e18285121ec4d92f642d00d09da801d444535a3bf549d03cc65fb1
z3d6e5196a1b3bdde461a3891c84c8c9e5d4973c0f5fc5cdfcbba2f1b45fd51395b035eeab3742e
z2dbe143993326c8013a022c68c01214f2bc2e9601894e394ab09bdad3acd44a951f068f9e86b4f
zd50c20454ebaed53fc74c60167c183fa959fd814e14c0867988e78797ba91b9ef217a1006ea3c1
z8afae979a46635b3216a7317d32a2278c3b81efea4bd9bcb2fad5ebfcf807a25f6ed5bf224c525
z62ee5177f3dd87fed30f4807e0f56f34bac2fa8579fa0b8ae186ccf5c85b5c09d4b6e324c472a0
z3777a366ee9588b2f48c0f9ce7cfdfa76d470bdfeeedcc7975596ec21090e5fda80c815f13ada2
zf68a4a723c0a085fe7601422ba66426dc8add93d4717c1f57b8f197b12e9aa80989c8a785bbee6
z8bc64442d0ac9b82931d8d42e70bc996c98a46d2f6434d5521cf59171a091fe102aad367faf4a2
z8d2c21d4784d08f9fe558d72cca9dd95e343dda9e2f140cd74add14e1b214571eb49690cd77036
z5f1012297256db7d229b4c787d774e32f658b230a86f248696912c82173918344af374c4541962
zabcb86a42e8aebf09aa064595e0a8eee832456d76fb865659bd632cc85183353b28663f61511cf
zf122272458504e3b15d251400a8c506c8e8bd9cd5d11d417da8ae65097c97a3e61734a5e008eb4
ze7de9c799729b5c27d18b634cde9e96ace01dbb2475c8281e1b168245398923cfb9230ad344dd5
z23bdc60fabe2b4c36d8f8026d5c0e0992f9e7da486d98d6b08be0098acdd86c32cd5da31be6813
z1f30d96df3d5230a4463ee354ad4df4241d0fa8683cf50e24a7bdf9b7427f0668e9a86e317cb81
z841b61d405dede4703b2c3a697412958c22bbe6a58e26b6e92ea4d31185b0a452a3b61111ebdf8
z1ec0e2476e058b287df3172ed71b97ca41589bccd7ebb06bac3085d36117544eb5ff16ace4f007
z040461d0e20560d318c8bc5d7b26544c77fd8c2f479efb13b920f6372a9cc6299ca77b1fead4e9
z3ef193dc201908cd56c8df95dd8770f73c1c380e1c2a965b1268749b57310cee05c5012b844fa9
z494887dfa0c002fbb9d48c808b80e8521368353c3a201409ca33be5be9376dd53615d98b779d5a
z86eb0ccb66085637c2440a7d7948f1b4def9fc0ccae79fd87570270f150dd933044863eade412a
z874d93c1017edfb9a82a4fcac0bebe84760dacd8b724472c6c41d09371ebce82ced1b3688f876c
z817c31ce15a8abf94621a40280e9a540670b77e7fae3a3b52c93681013ba1be0a411483f228679
z1ad2e16cbef48eef46ec6fe40871de6f42f05cf879a91de57d8224efc0bf9410b408442e8dd8ca
z66336b46c9305672fbdc58082a305ca54b08c11a770c9ad43629047ae769691b5f6121c7d1d13d
z03b79661cf69f72dcab7e1a77e6ef1743b8ed6e3da3a7c90a4ac85f778c8c49aeac574390c2d6f
zeec8f80126399c62a12d21f6a6093ea9b3f18456cd95c3b9a43d6aa4dd3b5dbf1a616df335d38d
z8b475b4b4fc397b163e216469031198796153b6734425802bdc02a44cc7b1d89a812e9441fe873
z46bbf610ce7c50d12c5d3e20b54b5fd581fbb31c4fee57de2650cbc446430bde261358c7a382ec
z4a1bd93e4dfbe29b2224e28d225a823e584afcaa4cba72105dd67b97111efd84ff95dd20433f1d
zc0c65801fe29f1f8677a2716f6c97370ab80de63f5a40fd9580e5b6333ff3baa8b7cc370455730
ze2b158c956071e4b1359007f56428b8af6c5e6171d33b5e298e1c303db37d08bde32a2cdb0c642
zffe4062f8403f2750d1402b65b298de26f276d60e202761c875ae198fd5e642fcb29d776a88729
z52417f6a0e7820ed316d876ba9cbabcebe285346e33a0ba35d80805c2319ecb8bcd600de968942
z6f4452c9448d592b4551e9cea2863ef830db8412590904425aeafeb0d6d5191eefb1bd7027629a
z99c4b1ac0f12ee8b452571a4c8f971f9121bd4abbb507d3623af091bfc35aa45f9bb22889a00f9
z61dc95f4f10ba3b507490c56c10d0e5285cbf3363acd5ffddc5b902c060925e2c2e94a8325e387
z83a761955d0fbcc41197c389ab0e853e4071a5941aa91eed35cf5938f1de49d75daccda1a6a114
z56ed0aa281744fa2bcc4c5d30fc5997818584c841f9b3afee315dc15ad8eddf2b32947bd33be6a
z651b157c1d346fff8e1e4ba83724fb7cba63407512ff4ee7d689e19c17284bd31dcfab1e2830e8
z10284c361aec7b54c5027bec80c223a37527cbcd14efb5a555e05e306bcb68c35bc451347ce17f
zdc54715c36aa5861a365f7ba6239c98a9789d29761632e41a14c9bbd8ea5998c02be084fb13ebd
zd4526e2e2806d5e71e4506158284e2ee4c644efaeed3042134dffc59e96c74bc9cc7c358aedf83
z8725515a6471672a2e5eebe9510444a36b0236189ce0b488ebf7c499d45521fa5b3c670ebd4852
z11995a619f9aa2ef349782943ec9305124ce784f20b19dbadddb5740b2617fbb57c85d6dab34b0
z444cbe16e1ef91144d5970d083a63e0291fe4f382d7f07fafffd7af68561307fe7c3e409c59487
z54c48ded7b0b3ef29fee78604df3fb796b5ece88bb6df2fa9ce1d5422a06cae9cce987e4efdb82
z2fedf0b0dbf6682c479412e72c9c699715e75c77d1d7a0308bd364faed39317e95a0c3d6ea96fc
z473266fea0255956c1a3c4877d5b5ad18be432a232d787ad34633484dbfea51ff0c4779127dc5a
z09f50a9a29dd1a87672227eaaacfd2e770c3a98dbe023bf0d0cdbead139220c89d1207c63646df
z87a5fccb02a80701c630d186de274637cd1bedda7e089c8b6bc358e55e5ad5ef3b768e093f2d83
z43ea587d10ce775e8791a3b3dd5b7f195e47eb72a404498391a80f7482a5f6cc4ccd35a2ff445f
ze51e9fd6e347d2a257f60a49967e853dd31f86daae74d3e1b8ea69d5b4fb02b94c5a19cbff05ff
z984feea9e71275a32edc43955ea123f780d41c1f934654b7515846a07c932bc59b26126c3e201e
z37cf5bc33a2ab24512fc562b0a43aadfdbd88cfabdabc787df6cf7c84dbece4e62ee90032dfd67
zc208f1ce9ea29b29f9cea4f0780ab7148e2ccc09098c62b316692ebdfeb261df454e92eca6e36e
z0ee7806468d378d5e2f61f2adabcf3deb556699f9b86425b0008bd85417227752dbd32a9e4658a
z73ad86678197da0498609fe6a75e7d6fddf566bdfd4491169e736b2e97230931a04cf2711e6d66
z2b6c07cc00e597837d038625ed6a258e0ad5936425bc3571c6e13fe1206803a15d9e94d44e0f7c
z89295aa8e2dd958a6040c92fe99c745b68a015bfa223dbb488cfd18bdb45ba7b1ad40141ef1ee1
z82892a579c262f67998d2c7c9be78f35c62eeb196a287534f22b559257154bb7e47c158b8fb285
z0d326506e344fdbd1473ebb20e9b8c36ff6d78117e9b8f6539769941914e76f487705be48add7c
zaaa5ae6fe37c3e162a1e81c0105f00164e259b08f61070458cf6ddd4f436c27d0953145e7c461d
ze7b89affd1dec330d75fd1da5eea9f044d749a08770e93e6382f69a04d7976bc225c428816d5b9
zacfd0bc4f826d00da90edb10058848e8a21add435564cf51d1f430ee83070b8576d201534b4661
z987e8cccd45d291e7d6bd67f75f5c087b24e49083bcebdaaaaddc92454fe9541f40128d0a645e9
z961306890bcb6d261bcf6d20c4dc4768be89fafcef30d63c9922b8219a1bf95ace22deb74ff4e3
z305f55d0cc4c8c38e60c45c4eb8cb00efd7e63b56c5e27d361189c14f41da3b24f0d00d45bbbcb
zfa8c9871b7be3f1441bb20472a0372fb71ca4a873aa574c212bbdd071a68bda7e96126b75bcbd7
zaca2c432ce5cb5fff3e99024a2089389010721f8280b3c3a182e4d30175ae17a888d7510bd5d77
zc2be758606eb371c213a7cb66b4d205cf61d4b3a292165c5af8802f43b17f4a33d90c37497fef0
zde9dd1c3fc15131517ff4f39dff8caf76f29452ef6301a825c3ecca793903adc3160648039b7fd
z2717c90b522e7c7c0f337b800e8651655313412bbe15ec1ab41369f6e7477d658cb68e5033db6a
zeb3537a9006dd069860cac5c78e9eb086e502fc4bc3dda325bc34441170e4785287b80646d0ad0
z2caab5ef8fa7ca56430a4d1d26f663402ed446a79adf81d0d4a26ffb957faaa82c6bce4590fd64
z137dda8f8b1ba383b7f5d185f336e64ad0e2a09dee299f0c6b7e1fd0aa7bd74c69d74b027e7ea6
za9d8ca1f9f4604870969d4c6539993cb90a4df821dda611a6d45d06a3f5e590e24184587568faf
z910633326ca2e7b9c87f23f2a5f84ca327403fae4427cc8ac99819217a4534176eaf0bfb5c459d
z5fced5e26fc0617487426ae8848d4cea886b88ab6c8c64cc16b3c3e27c29f9cd6f85255de31812
zc36f748f509a80c87f9b2f7e5042aff278d664d5520def8eb15ac2dcde9bb7210947c24edc940b
z81bf0f5e35502de93049dd629f247a13f6ce91787a9380382317f2f92e74f22a8fe127824a0453
zcca86c45cc81c9d61a4d73ea4d9f441508b3b2b913981eccc46b766e62a033b4c46035030c9cab
zc617a6b5ea7eb8a0c9b7e6e1fe643e5387253f517d23b64b3c7353a40ed22af9efb8b3b883d397
z6daf44c02e54a58731141c6156c7e4fcc689d3244f1df9533b16032af699595ee424b9236b0220
zf330d44fff711cf24f7969d70ff9a6b52e6288e6100117a67c458657ec36ff6468a66f24b7f4a1
z6ef5bb3497dafb6e9095398206787aa9c6b7a36c6ab1fd4b4ce352c946d71212b6008e4159287d
zc4793487633d98befdf39e3dd6fcdd9a5111a8854b1e7a780b7a42690e28f48e938651d480e67b
z73a1c6817854f3303ec2713e8f7614a09e3586152009d9f8cda3a450b0d3e0267f91410c2854a6
z317f7408ad559901673e54039661ce8174419adc07c0d9b992e9986d2492989c29424b37c42a76
z70d9849dbb59414dc38bcb1fe16ccc0ee0bed4a6f239049fdee90c93984725cfd556c2a48f2297
z6c9e2cf4d430f856e981c1c6722bce0dfe20559b33577aabaa77c8d69a5bebf867165ddebd3abc
z4cdf19f80bdfda50993fff364f70c9179d69acdcf173aacf84b316c61cecec523f53d872011b17
zf70708387f847a438ab4c47b5bb314acfe386a8d075e556d9cb5c8094ad45b1ad236599a45bfb3
z944235adc0ebe722b5ed179512a88434eb5cbf08744ded7e6bbf7122b34b911e811f37243dcf05
z9649ce1737c04896d33cdfd01141919eadd8434d37a361cb1d24abc96df2d4895c0ad000e419b3
ze71e052ce71719bbd08fe696154a817d2afad60281a288d02dcb8e0d9817074ae695e102cfd014
za500dc1daa9e10a8f950e48c01c86570189219de6e898aa127d716e525b1d728665c1cb180469c
z8326b12eb56cfb43e914e615b2c73392aed9bd62a682db0c79aa4dbbc5ab3ba45156243230540c
zdffdd5be64180161cc5720c9cc6de3d0f5ca92ff47f3dc03f5ddb54d724918b2196674213bc507
zc83f9b8ccdb3c2abce2a5d9fa638e5e111b42c61d80fbdedea561e659f32e255ad36eea24fee7f
z454b358d931d35b59b81cb2d4a1763f1b847321a8b7c3af2ab3db95fac9128ee638e15af0d679b
z3fd1ffdd7291c2ec424f78d1968c5924900e398a834bad4505ea430cdc6c6f4db4af6b4da7da42
zbcef8b97d5e119c201b307e60cc803a392b99edb56a18758b1aab687d24fc7333e1e850d801327
z7e72f7177c49f23bc7c518852fbb0d1349cd190155f5003e3b92c4fc896d5df56d4a01119cc805
zf3d308ee81520aff4c133087ce71c472eefd8906169da29db7236cc020bedf60758a62bde22021
zb5a8c5ee480f9afd476956de5bc267a1f406a3533cbdf6c5d872e9b7c7fc7872aa29a220c8d7f3
za3e685d2bad308259f36bac3ae65a06c128c7629786345100d84811262b57805579b2c050a1ee9
z2bdcfccd65e3700a5d920176c51ca21ae0aad1963529382d2f282471937a8c63b0a34e51142bc7
z6bd8b6a72eaf353c23d9d985d0696154a61dd9aea488034c5eb265aa4275ce2048c3c83639ab92
zfdd4217c55035e76245355707e27e6347c31a8c662333348fbea5574fd74c55b82735ccb8e160a
za2770facbb8107573274468d94cae3c4722dd32ac51bfb943bb2954ae09b81191a464f48fc8c1a
za4d725dadb5d927c89db8fa4fb85715d0b57990a9d664b082a6928ff47dc8e20a2deea165f0f73
za1909da83494e60b44a84857e7e34c8829d269992c569b89934445a8055b57b7b4a4fd980105a8
z8d0fab439cf5e240b75f4b7f3bab228fb37104487ece5792b877c0d71dcdf9e916fa2aa4f76de5
z6d08733645c6a630b03c935f45038cb751d58dd10d26cf38bb5ba53a5ec203e8b05cd8b1d91bb0
ze26f358db14f01d528f3b4656ddc3594c42be64901285c4a6d2e048e5cc74a54a9588c0df7c9f6
z901ed266b0ad3ba029471ef7d2e9fd06affedba5010a07f1a46bc2f7cb36ad840fa940d5e96fb3
z4872c5c79bf41b849d27601a96dc0ac453ab45885c189e6296474b64ad755243194f58bd5943e2
z6f2f62997e15b75c0518c64888fda27a0842dac02b08af3b36c28b301af8d662d5bace6dabccd0
z895d7cdbec75dd094d8df8aa5f66738a7650415fcf807f002adeb77b786b727d658175c61bcb2e
zd12cadf1fa05b90465d44535035d9ac64711009305be3716af42d4287c6b896b0c07c56a1de9f7
z9961fcdd94a0331a7659d872dcae504c74a3d2f85cd47a783e375b6b2facd5197828951eccf82a
z151a5dd682b40654f354cec18b7bd7f77e151886a513b51e8588c1c686a97b3c83303d7fbee77c
z121464c617c753b5c2012ac3217ef25740b4db2b16d11d45f5a3006b416c6a2db7911291d75fd3
z808b865bf5209cbe5997b8f4982e6908451eb04b09fe6d6cf7aa2d4962ff1804fe09dc36ecb273
z03d87d18614bc8424ead758788ea6285842fe4a3f6aa7be8e88cfcd3202c15d77a8cd41df59bb6
z4cfa6a665ec12f911e7b896f13d366b3338dbca0ecbdf6247d5b4ed43592cff98d2ee3024148f1
zc17d6aed773b8a1e3881a3cb8eb6cc1cbb51e1d9f49e865d598f57a95591f7eea13ee83b0cb0db
zb27a269a7b87e8027b4fd0dcb0cb67b52292faecf96248d5f58f70142bbb2129a6927c7b376afb
z834357fb536bbbd2de8c66a7c7e49493bc5426884d72223301e7726b7693d6880700c9c84058ea
z394cb364b3928c2ea0637646cfccf5d6305a4eb79fa899afe6ccc5dd31db9127f8a7b838033183
z0ce9d2b63445966ea8cf65a7f7817eb59cf801e62235d18b5b5ce1f1a2b69211bf2b8c7286e5b3
z1e7d8b09c5c61ffd8246fe69dc314b8316b1d24dca90b894b91119ba2f22cf562cbf4fdcd791c3
z25e4a6fefaba6873fbacec9d86792b2e5dbec82517de353fac56621a0cea5d0c4ecd1a22153887
z63619e60a3bd75e4150829f32935acb946ca44abb41bc4ba5bb5b6f0b636d61b148c6fdde069f6
zbcee1694ffca72b012784c956eeb7c337594c4b7b80b44efc2418a6393ce3a29287540cec478e2
zd17497aac9d219ea7e8a6ff25b2102b82ce7924662252c3130cdf393f33628924b776537931daa
z14f287447f24754df5ef386a174b238ed2f086c42d8dd2e7297ae9a78f4aa5510d966a02194e32
ze67c1abdfd253022fbccf25ef9fa5df3b5f9bd9017e4d99123a813569b84e669b9aeffef2c1bd6
zd981179abc93653535d7ebad818bda0ed40bad825663202666c7e43b23ec9d98d4900c286c738f
z26fb7e938b6a40c2f96d100d951355817e9dd74a5c23a0632c94cc5de1f5bec6f8cd2d13bb4b09
z2aaa9f2ddcfb533f3eddf562145e3a4de309d95a8a14598c281cb4b0223acd02b312d8f48286f8
za259cea9a2c86d74bfa1781b5b5297d29fdc0cbe11178a4f0560c96d708e4a52e12cb8c5b0e85f
zbb922f4a320a435ebe61eb9ff59410c5d5acb2c67df83cbc80790c66fa1a7873364fa08b30e704
z007a7631fe88a8b0e4f995893b1c1d77049b4974f55262b82a3bc56b737461a086eaf026d0ea17
z78a928c278a7eef981744b0c193d9b23ce0a6edca888315f7b64b3f022fbe27c599c11453f21d7
zd85da4144411b537a37510cb67d045ed3f746a0f464786ba2b760ae6b24d6ba6f17385a66ec9df
ze9a0333228f541e362990d5e0c19151b2f7b39e528c6fc33ef73a0f791bbe5b15e769d369f1271
z696c41513714f24ec22aa4cfb3219c0b130788822b1c081baf17409c87be01578c512409b9c86d
zae4a090d320a7c33142f40b1ab89e33d49802a6a0f2f907ba8837f7e4c770988c39481ac3f3d27
z07773abaab565d41120fffcb6f340117f6f28585d96994d1dc0752edb2b6dfe76e489a0335ece3
z0270fc7d3a735d17df3ec6c450f211b39499c49b3c1dd2d932f288b389b3cb8011b7ec880b55da
zea9dc44cd2a5332513423abd2879f99e53ed515b47368ff6781277d716706a2a066ea4bf1da004
z6c2a8209cda5812262911e22417b5f2e23d6f1b808490898b22b397768887f583451cdb91b4350
z60a84e48c5ef4288c1e390814e87201c5df316a8e86e54629adf15150eb7c259cbe4e9375c4bbb
zf35227269e278ad7c7ff246cc1704df26076050c2ff161f1eab10568f64149829c298decab8130
zdd60c3240610e8df48514541db564416cd3f1a29040d48a51276595a04d09e6a453559ae20b1bc
zb1673472911af07862e55069dd3273670bbee60750803849b90708b1a0366d0fa500aac06830be
zcdf42c3244a55093003c521cb591bdd49953c71713f6139cfcde5537558ce2d97095e6165737b0
z9e9b3ff7ed9fabf23685daa3ecf9a030a554099faa1608ab843fe12501bdb8dcb86022302f612c
z33fc0e74b767a363e99ed4241876ad26a003fec3b8456e1d86321e530df57f6e07416386835a54
ze2ffcf9bc438bff8954105042b1023ba8c51759e9127c0d9dbeb5d7851ac67e07b5e3a2eb666c6
zf7e8be64102a909c2c98fbaa42b69097b07e3dd65326608ad4c998921f816b3b9ecf5d78d37318
z9b8ab6cd769f602d1751e1102e3fa08f993e5b7e1a9d5f2493108274c11850bad8aafb35579540
z14a62e0cbea57a57e8b7f94bf5e26253c22b37fecc97db8eff8c9159ade854c77d41208a12156c
z4dc4ca6ce5cc9113ed8f542b6d3d717969b198d0ca0e0c46401d12d7d288fe4318174cffcf48ee
zc1e2145fdad3a3df2c19301a3ca8388635a9874b7b234064f8c4bf493784482711748bd0eb0da0
ze752e6c3c23c374dbd473aff8b97d0c7dd611d983602b019532ed25fec377389705e9ea6d76b7d
zb651c5dd9e69d8cfc76ff32d111dd2037467501608bdfd37f8ad2e8c263047020c2d1b34e4d749
zc5d4c7e5a0fb694df76c9969644476f6859df66b328898f379ad72b60f6dd0fa713f7a08ce9c3b
z1ebd12c99560a17c884007230ab3bb4caec06d6ed47685ffcfaf898522815533158d8c740eb8ac
z562175c0fc28afd6abd85004ace15ab9d645e4c95a682cc9fe89e55882ace358da32beb819f9c3
z6cb1b15258b577e6fcacf92e203efbb860cc4429dc893b0716e1bdb5e0382ce3f4046aef324f31
zb5490bb017385dd037b3980a5ed2264670bf6b3c23f372a4c6a97d67e8462a4cfc29a206ad54f9
z236c40509937afe6eb637a2c107590d87adb75e104c3bb4d4672bf7456b94bb2d7bd21bc40df6e
zdfa464da9e6422f8aaa708511835230efc969924c56ff5e652f880bf19b3462d50862e5a9a83d3
za8ddc4f1ce90090a78d3e9dcbf6a8795c186077d0d4fb1caf9109610fb2d7051bc1e91189404fb
z313ad5093f79a27ca091e397a4db86d3bb2aaf1a41b241d3839af3114a93c094d98ea26d1b901b
zc0572e0a68fd78ee38a20d83078396f4a6c774f4c6919ed3dc3c8a2bbcf6eb6e0a36695e868c15
z7ae6b4d8633190aa03b2bbc3d99d1ac08a47d2aefe38a4a42ae303f9a5493a01aa3b149c4543f2
zf3a0f8eefd4455d0a0c8035f8639df4d94f95608bddef239930300aff4d28bc9761f93cfe8a7b3
z186f07566d2677690a9a85241302875d6d9b540c4587204bb054975ac6fa4f723ebb19117ce19e
zc769057b4ed1c0292c0a16ff3ff3cfbd6bc5263bc497bfcf57c60bb816d01d4f6c03aad34bebe5
ze2a06f297fe89d9d79f0de2f751122aadbb9952aefbb22433998ee817e0e39456072eb66ad8779
z853f67d9db8e6c112eda5048e8b1d75dba7680d745b20c6031ac5ec186ddfbbde7523385170f6c
zda12c94716dfe83219c36fec73909576db99e647a20561a977b09ed4897f1dfb76d31ea16797a6
zaf9b99b43b7820c9a2ae3863dcaa9dd39fc71a968167d765c5126ce1d55e24b283c683e1f7fd08
zd8eb2b9b2c4ece534dd3e7f71e1f0a709af97df6bb84de14f9f96e188a123368851e0cde961dd8
z18e109efa67da86d3d1365e1fbd02555dc963e42a051d6af7391affeaa4d9bac2bfb542566e551
zf918ef85e55f187587104b9c93ee8a90bce4f9831eb816a22aaa48b4ccd7c475832984b0c97bde
z33174ba8bb115787e610ecb9603e92f4a970eb81e1df7f694402cef02e0324d78947ab663309e3
z3916cca6bbc047798658d6cd176be7a6b8477a74ab9b2ed822fad061efb0226b6e644d4620cf82
z8fd953420dc6f7411c53c709d3cfc59c109f36d978f2f263cdd5518a8096b5545b56e88cca3957
z9a7546b47c3525ccfb4d5638d11c3580f321890497103dce1f124f88a875d36154df3441b37fbb
zd3505eebaae9d9ccadeef19820a1ffd1e6694b9c94c11405c0506870a7cee01d6e279b147251ce
zf5fda623ae7f7358934ada1f5177ece9f5d8b97803654b572305e1bbb306ef79f8be88dbdaae64
zd8677b9ac044c73f2521c1bb2981466747ba02d496c7f1bf8b1d3c700c999f3dc6c6ce361572af
zf47be618ff40e94e3896e0e8bdacd2c6b1d41a61fb161b4a22fe1123c6dde842ba80cd6347d2b5
z5d398777507a7aa1cfed0528006f615dbc650ac6f70e87f9059f739e42a580f51f9c6253c9d6ad
z7ccc3e066851f19c6fd53e4373e09aaa2b614b1a724bc704e99ff094ce2d26eaf5da6f9e8b7034
z14b0c38a44779e537ef61e6db5aaaa88e2bc510439bc17684803a55ecee25a7e98084303d1bb4c
z9869b8d324b1b043bd6a22e6e2c87e867a108c2c28c3f7a5a07c23553a34b408d92018991ca2bc
z109b4b05041a0fde41a6a7adc29acfc36fc88b1da696773d669d5d62dbefc4fca1d3e3f93f8979
z16fcb9557d0ba453033672182ea3158ec6e9bd233dfde29212d881cff130b3d8beb09ff144af82
z13c79feb76aa3cccea88009f039386c5eded6155cbbf261ecbc7fa688f0d4aa2b26e85e3c572b8
z3c1b11222e8dd80b68f36b75c9f3b752ad606dac5000eaa509c9fa972c6f6743b43aae84ba1811
z5e5a7db2f2da707f80681473d595bccbeb8630c2c2455db458b08388cd34f07da45994ba26b182
z4171d998ce5b4055c5c705eb1e9d08167e8628509ad86a95e1c21f0dcb764581a830bf49a7207a
zc60c4f241aa68780fae58c2c64be1336061ce4e2900df7b09c40b8bbb180d89b59cbee5f5ee88b
zc7ea25cfa2dbfdcdcf29f2f20f1acbf3e7d8b0e3f097a7c137f3fc3f8c989d961f6aa062450190
z1e0d06ea4f1c2884cfa68a15c2a16328be5e2f50395172141ac7d98272f918627d0cf6b7413799
zcb89699aae6ad7137225ad5e4de05750901826bdafcdfd5a7c4cdc1903efe3dc0dc56d53f9c574
z455a1f8293363a5f50b724bb5b08a156be5262430f55f0dcac242b4a5f9986d2ed621a6b9895f3
z55b2afffbc9cb5a70f93e00bdaede254d835787b4d0b62dcd0ae32737def03b5281d60b08abd15
z2257360e5e62f29f8406ba9ae2ff186e6ca5f98af3ecfe0ee5e40201a1fece0b99f54ba22bec5e
z6a49297158404baa8ed97a59175be64319c07f3a2909f04e5bda3ebf7d08df21f59a2e03bda427
zde4f433ee895c972969d6d2a351c43502ead50d4a630021e3cc00b9291aefce9318bdf52748b89
z5aa525fd6d03154870b1eb1fc84d703616f4a7d5343807e14fbc94383411fd64104e84ee6b8fbc
z92e28b9fcd352a3178bb84dd5fd734c646b8cf5f148962e2c48444ffafb9ab4692ed6902baa4ba
z9020e727d9e2352d34c5eb7fafccd9a6359b56ba64a184e0454e91b482626e31e569cf11495df8
zce1eb4e48be96594432961ef169c6d8fbc2960d4b7bbf1af6c8f638db32a0631ff965c97cce77b
z807424872f0eafdc21be30933ebee835890b128b3f3a4b5992aeff99a270ff6a3ac31f715d9304
z16a94afa02e124aae4fd28cf33d2bf7ae233c079f46bfd8964dcb32086bdea89c6a9f05f1d8da9
zdc4d1784f9789fe9d3902bcf55dba6a6d8867c097bf3412c4bc9116d5915fdb28c584bd78af58e
z3fc24d14ce602b4060a529a515a5884e9f1f0b576859e5fbf4607134d65cc55d1253ab1f5d3406
z1e82ef29e3b63fc96bbe2ecdc3aa720b5a95c020cc21ce5e2a708e967a7a3939ea59d42ec07b61
z89b876eeba4eb4c4c2cb81ab32c8f5b1f222c8703d922991c792b990624b0fdb078393df98296d
z5f81111a01c0b654d47a8a2d15577f4a4ee713c889bd7edfe6d0884bccc3329ec477d9f6b3433a
zb44545e4cc9cb0a037d2cedd07ef1c3d416c409efcebc7cf1d2356291c6c122d898d61eff099ee
z2c407fede0fef4cb50bb377138086a39f64dcf7ab1e12aed32deee9d083a2ef08b434ee2713088
z95058c90b41552452a90aec4af8b7dcfe6cc4f32426e756ae39fa4064b781e335192b5431371f6
z7ad085317d678ab3b06b8142aa8b23114bf23d6d3c60b23e993bfc93181e156b2a82b0ae74d4bc
zcd23760badc6b18640e0e39d1426a7c30dd002006649ccde3f12dbd04f4e845fe19f1a32b34c42
z061c36ab3c680754849f981f40b96400492d305885ebe1209705f534f2e5497e5ed0dcc1a2c4d9
z9198f5fd61f05ccad886f9e6ffa3cc5c54adbf48507e82e0e77655c702078b57078c4efbc66446
z2a7fe0e7b18e7a528449b777fb69ba29bc47df9d80a8b53114c60a9edd655008967313266e0b7e
z04c514728d3c6c478ea49acaae21c99fd1a29d019cdf00808a51ba830040e72cdcee8fa53f4793
z0348e5e1e49c930505d59b2caeb3be0cc6ca36a80345a03be2b3661b64b8e203b4026ea3c2f8b7
z771b2e75d96359c16265da5f22bda9b1d6179caf3ae4fad46fc34ddbb31de49da61944ce085a03
z574a40eb05856ead7ab30b641f53a697b7af68217e86ec6763a74bf86f2529a38edaf8a4c19068
z2e8a8f5816d461ef50443e71afcafa3fa88c1a7bba7b5cb1bc28636d8f5c0399d2848010efe988
zad3f389b5a3e11176cfcb3dd19f4beabe8a4b40e7fb70e7f5270a9f954a585265e2f49810bcac7
z7597a7212a0c521724f17a229a1d6c841fb869eebf7f3fbd14a614e8f202d6e7837741fed8974e
z251107de93816b3d7a5ce33d2eda2c7b54566c9582cdcf6019f385d62e4e129f1712ae0fa99e4d
zd3e54ff78110b9de84246e7293c3ca1f4a97eb969142acf14144092859c69e8978356b6a1f2935
z9271da4fb7909ddabc1bcc8f6345d5b20bb2d5088153852d2af8cac5e80708f8096af0351a0006
z27ebdf0b397ddc0a827b48c1b72a6ab83119d6acd1c384e699e9b9573021ccf2af81280ee7d832
zf6f3ad3ea117ff8746e19193601a1a38f591f9aae8f8a7ae6c3db7d51e5afa78fe00220efe5e24
z545a6b6a59eed4698e1d959470a2fb006347d696b384134f0cc2aa654dad46ef0b8463ab11fb84
zfafe2ea5f6d9efd7521227f0e6f31a4fc0c6fae5b9ad83df16648049eccf69a175538c22adea49
z42e326168b286288b8b9ddc3f33794a18a8f0d5294933b73e3aa9d8bde05cb7ab15e00794f27e3
z3761e445c4838af9f0491ff86458757654eb44e9ec9a7a126fdac8329a9d6c64924228c39c8341
z5e7fd9b316fe174bed2cfcd3fd7915b29721cd8bd13c0ff1064b7671f0aa3b0f2054cfa8c38dea
z87aebb0b0d901b5707d09d6955de9e702d5d3bb19f35367fcdd19fc2a661f767482332e095830b
zb1a36620809271419ca07788b0a9eb149e4645566a0c409ee5d10d4bbe674fb8e1ccf2867c40c7
z54996f727f33020ce5808e03686b4e113291cc9d81929ca92ce2d1497fae5f634e35ce9b70f5c1
zfd7b265d5b04f9983db21a47f1fd4b763d81285dd692b4d4c6f4c8f9e32fb4823f809edeb1792d
z501c7977ccba9ae01a9473639d65afa6dc5880c197f5768f7f16beda57da1c3183b6393c945c4c
z56fcbe60ff683e6ae03df86559754556cbb4dd4984dd2da356156e605573105b257380788668a5
z3cbfd2d63d905f848fe3594fc4d605d2e79f3f9cb7b60744d4e90b947a0264631f1dd044c1cc00
z78e3e1fbb5ed91c1827ff0b49ad159445c1d0e92bf7b84c4d4f5587cb6ec2acc27cefdcb357bbf
z8b503a0165b9887e9b774991ceb6c623c1b2e1781c00f15bfdc5259ca7916703d57a6060286b57
z1f847521ad0918ce565493554fa8e37341a41cf4863b52f25e2360d1f191251137a78fad2fa2ec
z81a72b2d2d60c014be9ee28cad348b18f0f84ad550d33e7cb7e74c159bb001b0c93c9f4e17383e
z54751f25e8943a07dd14d0749414d2df07621c2694fa8064246f1dd40c5e41ba84b4c937601db6
z4ec25e481b5357ff927159417ee39859135fb0b50d34deff235759ed66b91a6d634a73e890b738
ze67d07e598186b08491ab4cbf5658a6f095f8cd484da89d402632e38e074a2758f1ea354c52a47
za666553f3667e0660a1e7f9282bdb51a1ee72919e1c85aca4c1037330d4297d9e43040452074f6
z0ed3bbde1145361cdac5d4b001334bf40bfc592176af914d2f9791e58bd95c5496028c9c4205eb
z0020b0b54d611945c6b37ee8a6b1294c06f0c848daa0b27d8caf1cbf93016cf709afed924949f3
z063dbaf2fd6ea260188ad3597f20e0c30b394f45b91395901254fe9a1462e6901f87f61212f379
z3f3d859d26a93c6c8bdb0d7ec6b79b7421c23e2ed97fbcdf63152b0b3aaede471096e01a22b6df
z731e5f42ad7c5cbd04120b78fa5bbbadc190cf5e1d77d12d2df65b209bca8d1ed88defaeb6615f
zbbababe37b498edfd557594d5c3ce9d3a3a3d7f90090a46b7915d04bbbc4ea9e128528aba50e4d
z9dc6e5cd91d9e4f0612864f112fda9dd3004d255ff604933dd5348aa81b6c5f6b670616f87fb5b
z7acd1e003c5207f1a29c49df7d3cc2aeab33e4524bef8efffa54913e97b7dc71a1e28a032fc9e2
z423da9caaf30a4b12091b14273225509b2ba9d030786733a98b6ab3815751153ced78f66533c6e
zb82c38dde2fc0ef81619c2c8c79246f888b593077166ef16e8d8c01067e15d58ecfa99184427b0
zde6b2bf643b82858848a3631ebf516e71e2db704ecefbec838d99c67f145659f3552a92db22e92
z79368777806d9acd2a39b289be93a60d41b3c3d5a0e95ff8aed6f2cd454e20f7097c8725145ffd
z40b221c9d92d0d87f6b435ef5a088145dfe3d3ade35258c354c922ecddc7a76e9943f5b61dee31
zbf553e3302c5cf4e06d955b1bb798256b4ea3bd0796514520e0b0104b8b285add7699d35e0736e
zcbae39e6bfe42c8b0b2817df572b611d7aae8367d45078b6db2c881742ecce6d96aca9db691c2d
z54f258c8fbec753daf642fded5c58e76d0fa86f02b1c783f3b0d2d53078faa7c65a7679b10b286
zb6a8b483b4f8c18059ee8206c2313be052afdf7a6e207c2b50c2f609582d59f45026d35b734c30
z6518ead4f14db204eb786f71eb1664b56acb305b1984bd2008693e2128f6fab7e502fd1aade337
zb2f2a60f71d87e0a7b187195303720810ba04305ecd6200d92a1920b46dc5267dff9b2563a57d4
ze118de1488e9bd30b8de5d82adcd1c0120e20d11ab713b9c0bae2c3d0c5ec860004fee89c19e8c
z2062c2c9e9dd76f4d873759330fbf89fcf64fee02d88d122663870bd030a1649f26b3a41c745ad
zf2688af8ad104d83714f74ae7b9d967df6804d147bc4cb45eb0391247c07c9c64beaf7af56af3e
zb504696425b4b418c9a291d323ce23a16b7ab10a4d27315d45a3e9e5e0a151052bde4f5dc4210f
z59ec82222f5ef80897beb438cd391e8b028e69ce432dd8fdf8dcdfa3d27021a373fb1cc62f134e
z03af49756edce03af56780232c63c555bf75053876912e22761392fcd066144d544ad767d0f297
z161503ac8afd05383a03e04457521f0ee0e7511d2512351c8999befb39cd939451fc45024e72c4
z36ac799273ef5f5016652e94730f16d9fc78a311a532eca0417f8f0e70b5688d47031f230f56f1
z0eff4c688a3f4490ca465f8e48cdee973858f1622e2985401208804f63f0c2d456e89a0849be4a
zf239ae2f08f0cac15c71d1c37f8f9d8465bafedb5ec22bc9b2395e907d9fed828eb3da0e4d468b
z480364b4fb4ef833176a9ea07fa1050a5773a06b1db4b3da34e1bce9ccfc6074c4c39576e43d43
zc2e4ea9db640c671718a02df6c06ae6c4930ba852ce75bf3f852128b3bc41b6fbf675db7ebbaf4
z05093420f1bce6482b46184e743ca6331a8e9edede277316910b38c79c7675b8e6da6d0bd9bb15
ze2d75ad30ea0e2084e91b619a8ff58fe2d8d817955d7f88988a6b8533922a7820768c264f7952d
z1477d0381b2bd995fac0619c93f002623f30774454bc598275205e25c4421607050c68b418efe5
z39dc4dff457ed55047bc61dc82a47fc7cf216d065dc6e20773b186d48aeee62c17b01f71b0baf5
zf07b9c119bbea3a7ccc3f44c03d051876c28afda4c7ffcda509b0033e2a671b9f28ff5a56f87cd
zb056213619d6d16546d176a13a866e6cf06bb01fd0dbbf7b48b75ddf402e9744abed88b029b33f
z70f4cc16dd3cb4021b339135286cebecb416610325a02af494048c3ec08b87984c32b43d1fe3b4
zd0de7e6e207e9b5c9341b8d03266a129a707f4ef96397c5b49b66f79a73ea7a577873eaa284fab
z1708799ad7c3f1d41e38a3b28543e861d8309f89ec7d5ed493ecec286322301b76b4e2e01c3f8a
z13690a11b20ac9898d1c10a5517592e4d57b4885908003b5a6158e905312d79d63200292ffb0bf
zd0efa667673e7b4bf85f4e5ea17c10e135ee4bb2c6cfbe4cd03f16ab355307b71bc77a1f6d4a1a
zfc8f36bf0c833c2cfb98481bf1f7098e603f57e51af124a927d2d4062f4dbb15c47c6caefdfd3f
zab93db3b2071cde34270e3b07f613f1a01f37426652a56db309fbed8ef12d2eb3e62e8cd8fe4ac
z5442dc915f01a4f22c8ab3e14f37835f011015bd3047d98936b3abc1a56f0a86d22333a5f1dafe
z010583fa416321a87191e565ffb2bfedd84a57a31a753ae3ed717ea38ba485b533ca5face83565
z2585a15f7fbb6a65eb3e0245e3e3b437e047e598db25e5777911d4472a2528cae12d353e767829
z63a4e06d8ebf2b8e18ce34355a654ee8e3dde48d64fca55e4bc3fc0a0a1e794aaaf13f86cda905
z5f2ac30a6de4b1398a880dd24825e908117230930ab40092f4d569a73656350f6c8b68ef2fea91
z58db5aaf4ff8307a011883ecb7a0a15f1f6f4b5580a4495ed193f79bee4765c63d51b2bd76181c
z8efaa8cd99fa5b45e44a68cdf7f8dac79d2077b3bd2f7a1e95936b23eee9c6835d9b985f87f7e6
z18d2a8d2c441146d9b63b7619a7c51c6f25200fca9dfd1504f2728125ebf0801726ca317e5b913
ze8a139085e308abe171bb6acbbe7b41fb03867732c2f51c2ab0d5cdcc3104da68316cd02609e66
zaf459d5a1520be8c30fb1c3351d79224246b9928bccc59ecfcb758af04ace8698214943f557d9a
z534a2c122ab6583e4447fd7a30561a47697cd89ef2273c0bf4b3641898aa520da12a7f4df5ec90
z5077d6c66e78b100badfe6a37162ce120398ee8f3007f95336bef24bcf1e29a728ef94953823e9
z9b8ac095341d278ff2d1e10993f65c79667f81cf787568e6f5c1f5f46486cec50b4b820a750c79
z4a691cbe266cdaff43836b1ead3e27adce8f4f9ea6b3a52ba7e6c5fdc7f1c5d3a3c33aa933ce7f
zd960214e265b25a94d33f19b36716f9b46b30b10c91ed6ce98ce6026dd2cfd05cad0caecab3739
z647a681855719c7cc358a2a674af2c332d4cec7b3bec016511e5172b1e1c74f7ea91b6fbc68436
z4f5f1ce0a5bccdb880536930388d7d91dbc8cbd0f485e5c10b31be2a8052004ced5c7701f64acc
z0dafa70675740c90740f5c5e96960a1736806b50d3c0a58e5b5dbba3f280b1e83ff2d74f8ceed9
z19a142382c7c12176354059ada5d27e8e62f06e1e459d2e3f8cf52335ff641a4e4b2fcc2d6e36a
zd3eb84deb7bd883868ccba9022cbc187c35d0cd7c517c801836d4967748d5bf85c03e583747eb0
z7f48df17bee8158a50434bf6f54b6b05656d9c52881f68c7dbda491662fb39036b950d3ecad90c
zf0ed5b64da6206c46b776b75d972265b0b3cecb50ff858e8e01b05a95b7cfad1a20450774ca0cd
zd6c58b59d7db56e900907f51134c04fc1371e9e8ecec3e286c6e9e3a7de9bda784ab77dbd16335
zd53f40b59c12c544a561f9daf63617d11c2ca392326b5eb6e1ade55527b3787dc42ac0e7588bb7
z05d699688ae0e800aa938b2693d6031ac24db1d70845aa67ad0f12ea1c7571d34d523e1d283b1b
zb147ca86d54674dc6de8276bb5fbb22b4640a80d649105c9b6924fead5b931dbc44738944c07e5
ze056f626bf0d9ee13586c906c519b21fc585c0e4423e56a153b6d3037ca80be276b88766d8d544
z37ac157ca01e6f7de48d061effca5940e767686ad9f3fdd094f58ca44478dc0047fc4e0f6404eb
z7bf27d2578fe501139fa2ff90d5866ee8d2a459a2a42c74381cb1de28abb4e7c33b869cb5eb685
z22eaa5302ccaa02250e45e4d28bbedb2f6225ef9eb5b73a398b09828515e40fef5353f6e7a3de7
z668c828684cbb268141b499f32227380126a5f75eae8f84fce985fcf1eab55656b9b84530c419d
z1c8eb056e1a3d7372e23ed855a194ec4f4bb1d85c36075697d6fc134c67ff77203d59f1346c83b
zc3b36c377fbf401acd84106cdc557fd00031b238368d239db8c0cade80cc3de54f21688d26a05a
z2fc9304ea1739a81eacdd1c2c30d96caffcefeed98cdd0d0ed2da79683daf89ff6ccf2835211dd
z12637e73a061acf24eaa5c8a6ad9c24716ea7dff7cb4b80001455c9a13a3f2a5fb6e7c6a685ef9
z9e423dda8b898a00215fa490a3c9dd6681c2095721ec0df437c493763c326836b265b3b3602059
zde221b164e548efb9fdd72e9dc9cfb6edaf38469aaf397979b658a63c84e7a0743a7e9b6086d91
zbee1f66683736c6f835da4727091b7cbf526232214234fd97f11ed8587da4fe98e0c905122a253
zbcf99de8332a06cc008f5414652bad46de3b54f473f425e7d69a9249d5257a52362c2b84ac8fe0
z1ee79afb12c8bf15a74e94eebf015c2786e92245e2fed53110d92c5aaed785d2aa5a4292d970ce
z1ef88f3ad1789af2d78d83715bb6cad7cde40a3ffa83f557bae187929e2c5934abf2708b4d743f
zd05f77e8b8b0baaacc29780a517f845846006bf763329c35114ca75391f5c7ce229807bd6a6912
z9131e0ba98c0010d8c478c7b8451cf770c8f125571fb26e643dd7b8bf5897806d833657204fb78
zacdc0daea00fda7004f3517096365c83bb35baee288a2933fef0402f80422aa820d2be69fd7472
zdf29f22a46d906f4d296d00ed24a6263519610ac1decb688d9a4c7f528a1d392b7dce45cb894ee
zcc86a30196b2b9a0d0d0679e3957730d36261fa6756ce655fae8ed56bde112b24797cfabdf7952
z429166d7d7439f25d6a21b9a9030f43f331734788f3879ca322bce22643872c387da9c7f67d042
z53e1430c029fcc54c0f2358c9659388b01ee24286c210d59c2ec9ee1839f2e5fc3c90ab82e84ef
zfbf2f27bc4a44e5323197f9a32530a5d2eab29d925120c89e9d77365deeccd7ba17d8224a5362c
z7d14958040fa04309f3a0a48fceb44fa2056f5ca9cc64cb50780afd8b3c20dd516399ee00b74df
z8cb43ffea0bacfc85f02725a2b6bd257efffa48644569a5c384d125ddff60c6793cff6ed603cee
zfdc5fab9b008118ccf800ede9e3425ba4888e79eb2a4efc05fb5ad2955d33f593cf0a51d8d1cbf
z81c7c22ac364e2ad2490e4215452f8ecb1cfc45b18226dcbb733fa60d74b8690c5314f9f91a13e
zb87c3865a9196688f6ef7f0074199a47a7adfafd20fcd548287d85fffa4d03ceed5d894a9c34b9
zf971ea00efcf89cfa32cd1c873f38c6a1313d558f117ba22cb287de0ce022f562b24f187e57726
z2d9e8ee0aa5cffd11cd977dfe7b531275516ff9c22d1f9d1f6ac98384704176d737d24f360713d
z65777d7fe2e5c9c74b4c8737c501284c170ea08a65e942a65ea2de64d64408dcd91f4e602342cc
z474a4031dca6a663f4546e3e6f231c1ff39a9c9ed376553ee4157225cc9d45b6cd0554a3252c2f
z5028d62bf504f1325bffaa656a4e8f8440964dd630815dbea70a02291bb69b1fa8a8a07ddb2016
za6968a53dd2b63a83c6a1f2cb2803224603c64d0e95e75a30f63414dcd5b8778c76f309915e224
z9229eefb87a821ae8174baf65cb14e8da4f2cbe61c1469212febd8aed82edd0da7fff550c8bb70
zc850a7cbb7bf176507053aae0347abded988380b20f6c4befe25855aa692fed8a3a210ed72fe9c
z9764cd9b8910e7ce58fdcd5f435e1a4d472a83655e8cb89ce94321439b4826800ab5c3a9a6e7ec
z3e9830557d2c6b05c87ecb86196e51c763286c51e5c66516bb9729e3a00070333c475705a9725b
zc6de28cd36eb1afce34e9981ec2910d6ff69481e682de35660139d52ede5c0aa353f9011da0fdc
zc75a8e212633b87ecff9ed3fa3b4c986cd11909195fa337741241895caebcac335124c9b41b7a5
z951637d362d2d71f6cfb77f70a914169cf8508e4cdb224a20da9476ad626215d5a05ef0accef5b
z0a8083a614a2bb98adb37c67a0bcccc7461a7c0e871c578d6a9daf07baa7aa887721909d45b11f
zc935ec1b0cc38178a52b1d618c6e1ac1f73e7ee2f80533714bf8286f975be5e1a1ad5da893c175
z2b3c9f280f85b48bdb7c9aa0b021237c0b9110c09063414cbbb5334ef9f9a2cd2bd42432dcbf3e
zb1e772e49637d1d8abc787256bea7e908ed2216208a7026f83093b5d09ade27c21355b1ff54cd3
z3d1d51e2bc133f9f7f9f39f188a1f7a89198dcaa57e8772bb1e5b0474b1deeded517adbf40fab5
zd9907340a05b06b50fc39af7bd387a1aa4f9c9abdb7db0ab3a61109d396313fc0238d8d2c212ec
zaa498e8a7549db8636890f550b7bb4616d26aa28fc68cbef3114c2bc55d0842f0c261a0b741608
z1d9657a427a7b88e013ef069150742ae85fada816b450673820257d84d978b2716f4b27e3a67a0
z6419c192655706d6c32cd5841d13748fd91c548142c33679eee03c6f2f1174bf84fd4efe6b0968
z9be21abf56edb2ce41be8ada8b64d55fefcde42c02249b6beadcf5dd2a8e71939c896e8686ba11
z4b3665e1fdcfc8d5155252503bdbb64eba7e4864cd8ed4f3478a779476be149448a50e7f8166a7
zb74e52c59ef4c07f49d36e4d01348c04d00663df8133ec1574589d1808513729a40167199fe370
z8e58ad4708b016b4e0d31e717acccc1d8cbec50058a5796f62daaf5f6191de9462ad63f2a9fb83
z3aaf99cc63ebadecb2d2b8106f9b2e76a37e904d2266c2125036a9d1bbf2075c69d2c5546670a9
z90d4794f9acb89a2b0793f6d8380f53baac7773f404327067b3a11b6ffde440e3e2cc4b66d544f
zc4f8de533762bab1f293b81a7a5d3548df4acfcecf5629acb3f82a9f9389938c0629ace03cd487
zd6c44862c8fb95ee16d1ef518fa35d03437bad7e80fef0ba59cbdc03da381b9b77a74e155b376a
z415568ce5ef39c00c56227a2ca8307050cedcfdcbb66939f52fdc67cd8fd68fb56e169166e69cf
ze750c9a41a0856a79665bcc999e9ff72172fb2d294a5132796fcb7116e4ae06d2f7b7961de9426
zaf488895f3d926acf83585aee5ba2bb10c16c16f85244f45bf9431722dbf1f7db75575aa36b208
z695de622906580b908cc232fb96b0e310d9aeb95f76a6cfc6b787ccf1fb5bd1bdd07105ec4b50f
z2f3cacbe2a2a3f467553c7cf941efb80eb48f2fe8fa67393e8926b517202fa34fcc11ccef8441f
z0ca1a7824c07ed5ee5f7bafce37f69cfb8608ba64366188496e81e33cd7a02850ad349dfaa30e3
z1dc13f6de79eb15a988221337e89045f95a3af9f25ffe822a211eabb28da5af6509d2829440702
z7f211975dd659b4239d3367fed90264d00a8966c63bec7826c5839ad91d68c7c45900bf01f8e5f
z06603c77deb3774f63c73b675d1a958dcf51064cc9a92fbb7217b32ff5f45cb3b1c78ddff930df
z9bace1a0647b6687279584e81c0f1e6ad1149b0136725703b3c217153bc8dde180fff9d350a0fd
z11911d5770490c4ae7d7b7b133e9e61c8addf1d12d4d15eac2d308f801dabead1be6c78d72c0c7
z8bcf0f1e88fe1405137b126b841d4cf2a1118e11a8cf237af5533207e74beb448643e751f2572e
zd251bab165c70103c4c92b1b6f7445665b2af328fa086a781bbd1fa2202d70c1b3c1bc1a220e43
z19d0a5bfb143bb966875e79127ea78701f0fb51d6bbfa994950c365f01fd6ef054042e581bcb16
z3a612bc987dddbb7a0422d04c1ec3a679817830772503bb4e71badcde5d5c7b06a5d3c05cc01a2
z822f96d2de3364bbc8b1b70b97f84db817b7dc029fcf86e219e6fe66b964159cb67e78a7661e71
z42e4fa97a3de07c5c6aa673e4708adb30a9d90f77187b60229248aae3d5c1f90cc05b03bc3f2b5
z11ccf157d85b153f7ff46af42626b83b0067c6b458b4da7e432647fb2ed78cb661e892445472b5
ze8d51e850def717519ea2014ebe4443b9e6a2175251088c7e49923c180e0452ae5d35b006824e9
z9ba82080d5b6130643a738c6123b76b32fe05b40a791abe098f9c8dd72417c970c10cae4e85934
z1fecff82717655dba590ec8e2a739cb32da5763021e684bcbf98316a6fc3f1540967afefa45df6
z1e319dd55f348da3f9656e54f8dfdd505f0b7a3f288f6402ebfca9826b8a9a7bfe8eab66c79d40
zd4bdbcb6407aa4508c219a762152e14753163a1fd0c4ba013d5963c366ac09054dab05bec5ec92
z8909acaa73fdad2561745d96b1db9920fd699d13704b0743544108b2058926261b0cc47ba413ea
z89ecf2f719cffc2d833cd9803d80780bc79fb06158f3ff12fe684a913817ac222314f4b246b217
z8195cf524e89c3b851a357d0d9dca9a2d0baf02ba55f5a456165da24f38957bef03dec57eb13a9
zf07a133e0fe96cd732468c947e0200abcead7a33ac9e05d99442ad8b94744a3a4eb2a0a0eda1f7
zf46bab0ca74eb8461ba2efa9d14566e6a578c6dbf62d70d00ef54f35e2a181a3475fc72d8e8efe
z9c5936fac3ccd720a81fcf3dcdaebabcf9dc4fcaa15595e037c7b40ed9a9146f287b0a95db1321
z331c15879563c5aebc84986ed25e59592ff3c1f36acf7445e7efa101a8c24fbe99e1bc99e8f473
zcefece1f839049453e8ef7b494fc8964b6ef7842854e6c5b110f348f988e4ef6ee8ced4a4900ed
zd3a3589bca032d71e28369a827d424ff46c8f667fcece7ed8724bed824ed900d2043cade68f9e6
zd910cc3a9c2f99d281a3b8f94dd6581608cdd1967d6f43702ca8fd7f8c1efc97ce1a476280766f
zeedec837ab11e18807ba95c0f128031f316a718b06de9160bf4f3328e2ae826c204ebebca17444
zbe0460013287bb0d57c288749c237d5dfc9ae8ae257ed9f84a76208fa7a3a584347adefaac1c6a
zde1bd5993d364729daaa0479053c9e4cd28cc4f993c3cd1822c5d10006a3d32a4372be93b5f329
z13fd15efe27836faf7b896be101e5706127073305a1bea5363124af7ca337d34a754b0e7ad346a
z49a2ecaa85298b2e2aa62c18acbef35c4606445a41e5dbd0f3da224423bb25034f5ba6a017debe
z306b58f5f2ee58c92b92efdaa6e4763a46dcfc549923e6df2ed64fa1a7221fead0f4e7ac7f4431
z15463438d9adc5e2029f702449fc8ef232903ad8f826f45a288b0894f6a6f5a417c869320e16df
zf65efca67ed207368f8b808911a8149d019b802f6ceb1a7ef1533d2793752a4499de1b6a9f56a5
z263c19dfdcdd8d07f5d812b3f619d31a7443e47decede21a5a821e8f696c81fd7d7dc4b24fff5f
zd5bcd8cb9e48066c92a44bc9899187a30e6c7ec21a51d23f1b0c9dd9bad4b1811b5fcbc01b3472
zcde937760a64488f5b57e8db6df580058845ab892a55be195e1f1a797460687de38f022fba0af7
z5d3a402a1e9026483ff7f4caf1fb09292aa90d47d1bbf49447a9dab04fe7b258a36a39af569ee4
z717dfccae7b9fc43f070a0c9b9e8da4ba3eb2519c8051fa319f1a5a5a5c45d73b4780734532f43
zee1f949e621d9d2c71cca6194f4484f808f47f96cff79d3585672730fb82f8c0f9612c97e1bc49
z65a623ab73837244e63d1034495c5ed6f58b2454293e42988066f7ff6dbe5a39ede9e8cb1f6d3c
z2cadf5c17e62faa8ca0d74f132d7270f2b5f46649f3fe3cd53f859eed540754d9c0d79ff5649dd
zd401dc16d2d11f39bb49a69014edd36fbc0338b99417e11c414455a297586876692183d6944646
z5d1bc825d4dc1df79a33305d28b6e6ba3fafabdb5b62e3c64c9656be628997f61a96ec50c1adc9
z57e2d6d1a5e92bb43e54a380787c610a09fb68bc0a7879515d384eb02ad97d96dc8a3501d3460f
zf9c3920a7713d7d64eaa261ba36d2983e95f8cccc782968a0bfa260f903c34e07007ef0cdd4436
z31c2136a11abbad69fa88e189812531068abab068001a93d376c7e865d802dc35a2fbe9c6bc786
zdf33e26466e184cb854642325edf23ad9b2070cfb5346c367c922251da1dd94c88e16b535a7e38
zf8db0b5eeeec10954ab6864b9ea71baf5738772a96c532bee586e029f67d3c9057dbf3e7e635db
z4dcf957e5cc6705a7b55b2fd81fe4c958c0bf2d53ad1b95be823f869fb61be5d93e25d36126d24
zbaa477689e68cbb539404bd6aecdfb5a462d1227f54c4e45cf9074a8ca5f5d7d2290d96ed17847
zc99b452c27ccb5269c74452764e65f29b3cfdc5bd3cfa3596eae5c4372a736db69ba2ec793f267
z7711f85084a3adaef1226ff983d6efc2bd660ea0c2bcfd7ea9d6552f0cde29082c07b755966e34
z33165112e2e6e070304816174642c43ee0cf976da269242f1dbe5f611ad03f9daa121fc1fc6d07
z8ec26da8edbefc15c33d98a57a219e7f63cd6689c4366c159b9ee15914ee01bf0bf0d143696edc
zb7d55d11dcb4fc964a629168ff1027b001512545e6310af1bce4de0cbfbf8ee12b2a93eec4ad11
za1dac5b70b3d4259078933ef74fcdb64fcacdc435eccc4706e997179e185cbd9652712b814ee91
z4de11977212a25c812f38fb60d9e7b5b8b28ef449880ef3eda89f787be3a35c0975251c8eb382a
z10f03d93a2b67e5ddc9bde146498e4fd2ad4af34d046c2e2bef02fa7321072b5b8abb6d1d80464
zfd8f412e909d23ccc2f8b4144ce6430f4af113745485f22bbccd9f180d5c1654076fff5c16c38d
z891ec1318eed153e0bd5934ec6349dc7d01c68dc574fc971cc3c1a0893675aa29a9e0170a44de9
z74fa526f22f9e0cb082290dcb5c9a4d8a78cd4926e2c9a6e04b5e2ee2c77baabaa7ea813fcf1fa
z9a00115e9e20f16ff58f8814a84549b0f9ea3af446224f97e15e90cc759ddd8a40d4bffb59657d
ze2ef04efe7a3afaf200f9c3172b5de706d85e290bc66a03032114625f615fcc463fb1320177ade
z57c28eab81f7a1591f4a4a45979a384beab272f26a176808b39e5e158f15f51ff8f18e3c16fb3e
z5f9eaa43507d1603fcec3e25a05dd63f0e75d3c3dbfb80816ead53230f6ba9340d58a4142265cf
zde13524410e694a355e1839cb1217979b9b14cdece5b25ebb1d256ad3bb142e724d7831d3b5ea3
z532c6a38a6cb55f03d3bbf0312162c8e4151c242de8a6beed1d2293ff2a1bd4804b50c7e7a9f8b
z770716ff2c600abfb379aa66b430e3b8e8147b294811773a6342a290adbf98445cb9406f6023cb
za6577a9b17a318ae2016e433fd92b8efd62ecb1472ddb49609599dc64c7d40688cf59a05a997aa
ze9418066ca3d2f7d6ed3a71da749e5751924ccebc3323aa66d9f3437b7464f9d5a1ad71b843c73
z0ca0be2ef1a4a8b189fabaacf0c59ed1eb87c37f0a4149d5f88ed8890f548460686bdef19f817b
zd98a855602093bdf84b35d691d037667833b61212e06a3a9bdfed78e8db23ac195c3f543910d40
zc342bf4bf89721618029ce73851a5be5a4c098243a6f9d1995e833002c34ee3b8c063f2f02f9f8
z999c31183d10e0364b6804bafe73d6036121d82b5e46bca758e46e203bcaf224948f138e03bcb8
zf1b7bf6cf0075c420d104b3aa0b87c91b474a7ae4106502192e21dcafedfc5350a7a5512405828
zbccf494187457d9dc58c4d23df3554b5682e010cca4e703ad56899f921890adc103ecc15998550
z17dcaf01bbdc9538106e6ad55d6b952ab4ae47c6ca90162fe56e8376536c3399a82632ebae0c36
z94650335a700af9aadbf504f7de554374b611d74a47a2bf16a7a5b26f3658df2617824d46d75d5
zf458c1d4ab67b712daf95adb560ea27cbcf94d13aa59b945b61354c35a6c0f8e8ace1fd21a1995
z3a5bb8edc40eea3c420fc38e73cf95076510cfd8c519fda2c8bd0a4caabede5f4644be1f332e9e
z5d6fbe6f75808925d2c7b01b8659d98e158632b7695fe534d818942dfc4a54c1cde62fc8a23186
zc31ef3f6bcc3bffa78c1d92f62ed2a109dc297de0f3d64f0605a6acb5a1c5534f5a8567d252672
z5a18c57d24fb5bcbfdd714ed6e97019ff45cfec11fe963a5dfc046a583726a5eb6bace2f37f2c8
zfd7c57221f2a338c6059d6788a421b19e213ecf0af7df4d92e144f566b740daed44252ae37d0f9
z8c70b0e14184e9ffe744d7e419f5877276bc062a9c776be7955758eb32401a5fcb7533a4b0dbfb
z4c91ca64150fe17e9ec1ba5716c4e283a131ebdb4da777bb0ed5d808db8b1bb1abc8b0f7d88173
z9b4222c6050062ed116c4ed86f09ab9a9c4c65ebbcb37f8177f5e336cdefcec95accf3219a7da1
z5af8c7e7ab5aa53ba95d096c2c29661c306375e6c1cfee914e50ca3f3e779a1c3006993769fcf4
z899364a1790dce6eb91489cea1ed4b0da34bc037df7b112b341ef94af201d96328af9df8bb2cdb
z57fec913a4906e57081f4f5588f28821f6efba6025a0b8058a7a84953e23fe953bc1b79ef4b3d8
z2177fb9f8e12632a8b9aa6a36ba8e61879d50eb70c4a796cbee773019290faa8fde49c6c817a41
zcf705a1d5e641e3f6593f922f624fa3daa29d0743b594d4f3d2a1036921c63fafd505fef4b0562
z1e844824b90d03e840447ebdde99f542b9f6940f85ed429fe8c7b9f8ae29ff0ca7f9e344222752
zeaaf47b868c4f5cc889de2e1a21b1ecddb9d2ad137239beadaadfa4e45e291b543c734c258a256
z6584ecd342a3b3f87715089891fe2c9c9073a7f56e09c53df7e430a3f0b181ff525e4488e28b9e
z9e5a004806b5fc1ee936a33a02103254c7585b662fab30b44dff63e05cf9229fd5d69b7b160737
z93e2923bf43133317239f9a80668b543979e95636fa1d7249207dd21d46d3c3c195d75fe49e2ed
z928d80c74c97faf5535df21a386cccebcea6a38023845766c439623ce905def00465a7ea8cb097
ze7f2bdedaaa36a2e33cb63e1e09b1fe0f75543d71b2f68b3bd43007130db65473af0644a5e8cad
z504b0da7e599e981e5433a6353a3f63f0552ac442c7d158273af6f231af96dcfc38e000525972f
z8c3e90ea52296be504990b9a1a01687b1d5d3b389120c3ed7751aa20e838ee61b35d384fe30c3e
z765dc1aceb729804ca4c87166742ccdcdefd85477bfc85230f0f100242dcf3ff2b203ddedfbe4c
z9cd03e59655cd286ec11d7d7546a5c44dab45527f53f3f6639dc7c07327db1fb5bda924914f723
zdfb314d8f2e8763cff05d2bb2dcf883973c83db91b25713d91a325a2feb8bae013ae8ca06a57c3
z6f442d3174f76fdf42ff15961ed45761d2fc41405aa70b433bd88b568934ef41f17bbd775ee6bf
za66ad6b40915fab2621f9b53bc2ea6fa689475c7a5ae488aa537615f4fa4f8e501a1fd173e7605
z8e3793c796c631e9a018680a78ec96116fd23dec5f9f2cb76bdf081bf01b4675910ff060a25c3f
z5381c7c14c068c5caf559ff0d3b9a09f7c2613cedcf19259c20ab8875ae4a180950c3787bd919c
z4742854469c77a623d8d07aa5a8151b26ab959289a667bfe1446360a31d16fc38334eb06842f97
z6dc9708aee866d002ab2e45a3b8c3d2868cccff4b8a5b664a98af9fa12f67e622e13965ef87f1c
zd43e67b801f2d6986ee7ab51835e71dce6bf93d078c3cf967373eed40b9df467757ba25cfaa2e5
z7c5e0712bb9fa4a94e3c229c001d1ba6763426d0153d5ec557d1bb50e79e77cd815498eed536c7
z4e4555cd1f999a60a35f8e9d94672e8de2740c4ce10967c99ab272ce09c847d396b38a0dad4ac3
z9ebb1bcce1e6d51e11f6936849a4bcdad802a8b5cbe73c253b729831c2cea7d0aa8012520c408c
z28217760632ff6eb9dfcee7a0c7ff27dc5f2a8389bb18be03574842261fd8b97b407e7a6e54fb1
z7051622f7b60a17d7861fa6dd0393324d25a8e460b0ad236e84302495a4dd36ae4094ce2c40db3
z828edafa563f2c2fffa8146edf32d542f8c3dbeffc1c676806d596798c5148c9fd2de625eb4189
z3aea184456e6f7f2aaa1b3f8ead9b66bed560de4fa5ad185f461611c4aee22643234ef6657fb9c
zfca16770e79dcdf054f4f569fd8de6f6057954059d2e816beceb0f7f89696ba3fca7347bde5941
z377b5cdc6591d55486e3998c8ea2d9100ea784e75d5cee76d3cef33de7f3bfcee97c4c73997dc3
z308bb595ea6df95dbe2e07bcf883c63cff14d3b74da5b2392aba78c67670a1ec9ada509f0c263d
zcc2780b56c52aab54070454110df17fe00afa96a837e512919c281031e9ac9ad50c996b6e52ccf
z7275ac92fa359e9bbcbeb49c2d8c73cb021e1da71ce34a109e3d6ac26149d7b681dac82d3fd14d
z480c07067d552c5afdb3222513b552e1e4d543e3782c242b053df5d3d01418530b9350909c8965
ze74a560c87c5740fd62d68f9ca304cbc73f397569a2fa284dffe67a49104b6954c0014a795ce62
z205d4e00d3174fec25951af60495210f065379bbc4d9a4f0282481bf4d0c2ddac99f8fd0a1138c
za274e77820936716730b69335ddb0f10877f564baecf73cb74911c176c4826076d7f0ddd119590
zdf24a0838c28f32a1a4b3bb7fadf3e710f149c108813f91d3c283ad85cd3d72d3ef1c1e54c801f
z66db5532f1639873e4969937c4bcab5e36142afc212fe3dba5ca38a298eb4f3acd7d64e8320319
z62eb491784a0cb9ce4e11a3273008accd87a2ee333f75cd0e96b9b4295909de23b425f28d83c5d
z73d0be33fa958a8b0ed6963bf82256aaa7706085ad69506d9d5b98e321d78e03583b0c595798c4
zbe312cedfc568666c82a2e27d4448a8848bd0439358b5ada46e9935f50183e862cdb3b3c717d5b
zee765d688235b8fddaacc774f95ae0caceb113ad069f30e7a44933ad2398c086f568473441d812
z1ce6a3914542f7eda1d528fb89ec8bf512dd7ce0607f03f1ae5f17663dfa703895916a4b834f04
z43c44b5a8ba4975dd10853bd33f9cc1531e1c34562804e2e2cf6a48af0abaddf5ae349fd7ba186
z3b1555a489d01dbf230e61631209283c8ae3d27f7ef3567336b12ff3710a803fc52f632f0b8be2
z24a21302fc9f519978a7520c27381a200ffe3c1b7114d2782409badfd8310be5e3b2c5190932a0
zeb26d7488d1afa6a27bd292d895f5aad5804e133017468c08471d9f4b54c00839fe87a54b1c0e7
z780ed4f7b574c63dae2193f14e33148cac11d8f5694ce3575c97240ce013f97ece3ec0f02a76cf
z8c29653e0ffc889542fcdfb3125a8ca5f11f6156211f1f99d9a0cd34051aa705367dbd08718414
zba3bb72eb4cc4fd3ab83c5534ad0ef29fe7fbc7d71d9f09c95aebe804d7699407e4d7564a75dfe
zf5e182e7371a256011b19a4dc294deb8ec083bf2377dcca9afb3ffec7e6b183d666b43e92e4d61
z49c43c1f91e0acbb37873fb64eb3f8a36f5c661f79ba62011eb23bacdf8916e7885a2751a41d3e
z6e458ddbbe93b0b0bb7a1681c29035ebf790f0eeec7cfb259e62dc8b1e9bd0365fba143c86a4d6
z22977b50b275952e18e72a73803ecaee2fd06372833bee8ce1d5cdaa08c20dc688c81f0a752027
za71646c9dca2e7e90646ba3cda33b8798337b1d245accfebd376495a256db3000e9ee3fb30843e
zce85a6cf0a4304ffe88c3804aeafd9d357a31b76727199d71667c9de38460465f5eac0f6acaf1f
z2904a9311ed4c462598455656967b25e6746c401413fe69155b7ad66835b11242506975d7350ee
z55ff5c062692ebe9ec01d6ac4a56e50a53488b21483530b06fe65e8eac08edc94a0f258f5e93b0
zf3e54978d7005c00681064985cabacc3774016ee3b4c44ae6b572a40b1f0b3d5b87ee2ff545e96
z450fb056cdec8e6a2a0d9569eb13fe0d99a664f4aa25527eca9bf26349bee8fe766c81b41794cd
z4cef1143e4935472c65becdcb4c11557f05be0e3fa7fb591aebdcd5394d004b85dfdfd486524ff
z484206d47911ebcea308d8dfa3436c5782ecc33257a7ae785be2dbef7ce7e8f4c4c23aaf45f427
z8d652d9fca3113c12102e4599760c6cb349defcf65594a49f3d88fb6f2c3800b9141ea7e35221b
z7c5969703965a1f3c39054dbf94b9670205c38b90e31554d2f4242524115a28062947ec1055a24
zffddb9fc2174795930d07ba53dab1f584b9afe7c9c1a3c7b55da3ae8f1f7d7e3acd8597d9ebd1a
z32135b2ed67cae397881b38145cff84a0b027c3e5d9e5dbeae87b14c09fc2a60d8212fd84c4937
z667985caa350c2bb03906ea621b5a669ff4677e91ad9ee72ac4740b55e54cc3893ede89e17c481
zdf1dc7185af6d0dafee7f8d3599e65155024f8dc3ae6894b601a3ab5e3c5c0ee2fbd5ef63ae7ee
z35450310114d7537f13e111b231c67ff4efeb3615ff37bd2c0ef6b394f554165c528a368a19c47
zf37c6ef649bde6e451b9d832022a3aed9adc596ce8bef660db3ec7be74dac4282b2552b0aec809
zbd1ad7b353786ab885ba887cf200149db48e540c7272f92079b8235d8074fe19e5f15e9b2f9368
zfee94762e14e246a5e41f2c0981bfbcebd74fe9f23771d232754e0c5d88214077e6150d00cedd7
z58903e8333b09e5936c142e08537753aecc4b2f9f25bf219bd64e05b1ad12a20495d13e9947013
z521aec3c2f939d256d1b0c7e30d638e06a2fcc8890e3625517e3e4088098c57142e53133434271
z63c1f93f7a4aada214968581dc9f29773280a83c2d3b550eb202e0b9fdabc91f3fcb77d207e418
z70f0377c4860fab5f7eb1ff51f02da86b8c109015da4be6e50f5cbfd3e98dea43f283bb209e923
z62fc32812bcf75e1bb77b1fc46e12961e8626b3331099a9eb7a55cae0290ea941cfca07e3dcaac
zfc3d7e870825bb5b38f10928ea5b543cd0b69539db7d373427be218b0e9498287756f3319c6d9f
z410d22e414342f0f7f6f02f7adb159bda8be788c525fc72aba7f77bf42b39626aa3714fbdb7848
zac2ec787a1a2bec308afe21a1fc81c6349757fae773c1328f6a14dee193a08b09e737a17c27285
z4b0320f643bea22bfc3287dcc58f08cf61c5b917f73f76a7cfa4d15a8f2640eea0e0c4ed4963e6
z5574b1fe1f116a78e0e80c4df325b777c9e7c0a4e081fb798642dc1a1ad5758a947d0f3a85fb0b
z2d3eb73767f0126773be465099a703e1bf7eed4135bd7eaff0f177be923914765da643d10adcad
zf28ba4edc632ad83e54e916faa7d091ee4655dfb3a6a750414002a14c595d5841f7c9b8ea1bffc
zb8e85d7067dfb165dc1e837bb5cebfa6ff9d01fb543bef10ddad47a020e592e0f051e2213856cb
ze9f9488b522d534f108f2b9f211db8fab2cfebdfd09468f32de621f15c60762b7db4adb7c6d533
z11e6ebe76c96676663f6195060d12fa790647d1981fd2c8e176c4359c369357a04a772ee6106de
z3c9910249f0b1ab7dc2b67a5c8f59ffb116237e5744fc2ba1b7bd7f602c7edc23d281886de3a1f
z84ec00c13aba0a83187c668d50079b319500827ad0ea4de4f36a9bb65d33eb0ac4df50f822411a
z31f08ef4998fdd6c01f5b55bd6299fce4dfcaaf18a195b94b2330b93c5137dab7c93d0e9c212d9
z8358ac162d99afae0d7068fba017e12b20ba0e50222d1f4dde9ab86e9a8930092dc90f6ab80c84
zfee5231f24633a4675eca0c8c6319a1ef21c487a2c62a36faa12fa1625ae9abaa8bee0f5333773
z76c440991bd095ff69acfa1adbcaff365854db64b309f89f036f95e9d8da07a71f981b38f26a73
zb85d7f1462548f84d2205dba0eb9ef839340bfa9140bb2baf0d631840297682978a0710795fead
z3b5349648803de00880632f00f9018a7aefcd3c01ff867af4fb7549e3165bf95ff179e7a6d51d2
zeb280c2bb45c38d9d0abb6d95672cf9c9d2d873a6ea926c08fd6ecd2f98e853f9ebb26bd98b5c1
z4d0dd04ad5963dcc6e8b3f26fc2c05e22862ca311c4d06d57dffc20338440dd2cc48518857cad8
z5f8416baeb2be43f1f0e6987fbbb024b1fa4b08fe48f504cb1ec9f133e91678f29008b1813c267
z78726e663da248a08de179d438e5a63812246dcd80b25a6dab89c87f111925e2ab6c58ff9f4da6
z78973a18f23c6c20751f53f4e10b24c416e879c82cd160fedae0caee2c7a999f01399f306be200
z5d129977a4f173bd55f68e0fa017000d952d9b325a3833eeadfa03d2efa31f0f6a6e45d6403965
z38e03e59e71e231567cb87c5cacd668b5a94682c57e0a088cf08d922b72885ee60163688f827b6
z04936af345ccd50edba0613fcc8047aaaaa42664d135245b7d7009d3f1fe38720e8d9021366be3
z110513e4ff0949d14e2134832c9b5d546c15c8ef94191188488878bf7455b2120753a7ea0107c3
zf7dd198138e249c2b55a09180bd89f04cb82e035fa44e6fd8710a8a4663cea1d089989f3f7c889
z49d6a2a966c6eb27701987d1aa7500ed617534c87591a1892ad1d70268675cc718063519c19d18
z93bee52e19104f8b3f965c994f5a18405ae62eac89b415668b6dfe4a5d9f40bd851c32214f923f
z1b66f432e89c41a19fa19ae8176f3acc124f83d69acab4df8812fed75ed1b515c5c0f0b874200c
z26bd14b03a4796a99f096db30205a205a2e192604f1c4e6236890af0c95b0b2292b17f5573e9a0
za9c50afc8bbde267689f14835ae314816d148664e3d5fe08a890b2df682a973bfe480c2b32aced
zbb17f07865be93b1918680b01bf8bdfc104d45fb0e6c0dbd8056a36edb0b84366f89708601007b
z6a64f5b33f0790c65bbcba6467890e84dfffd731b67101a79489dcd3a4166280c2c368aaa0aa7f
z74a821d7e70cd384ac88a1599622e3d0bcc9c36bedbb5ade9e88ed22137af2da16b36db011abfe
zc62ef5e707cc564bff8a0da7acb67bb9f2d4d3efe130ce4cbff8be46260e161ccb03242b55b77d
z67cb3cf04f249212fa194cabdac58946e8d33340b79aee7e60a2d283e2cb55625e86f87007eab2
z1e7d49db56daf810e1a9e9ccfb779fe08b9053e6439afa72bc537d4604fa48da1c8ff6b120349b
z8b27da26c2e181e1c4da11ed46c20e5be5f2dbfde4c621ec113766e39588044269051ed9e18aa7
zc74cf345b7fa2e579c2c61d576ea8ab4a758e335fdc262e510ba24a425d3cdf6ebc139e942a11c
z7b756fa10e794b7429c8b41ae5872f85c1686c37a405c5fbf41e26ead2c0f9744ed20127e63ab7
zcab1953ee24ac74b11aacfb9da4377d160fcf6f8947c311fd415510ab0279355411101bf406b2d
z4ef051ed0ea1b657a55349fa084f483ddfbcd2aecaac161b7506817d6cfd7571fe0d7332d399a4
z2e63699547c6501f9d954494d2a3754955933c1ecf83b260902c6f144d00baee33b6099799e692
z8b3f5e8600fe657eefc95bfd66aaaf0c04737cb36c5c2d6a06ff7693f63361e85ada2c01cb1296
z7cabdc149ada1f34a5a1aa8997d74c4aa081e29fc50db9210628c6a2e337f52a6e0bffa5b6d4ac
z89e312988b12423b4747460a6f1d6f439cd1122a5192023a9e53df0e154f1e643d207816988ab1
ze7c93caeee43e6680688278d59a71708c794ca9df628848a9277e9a79f7562263fd4c1b6897737
z222dfbf9906422b85daf9640c298f2eb9e30c145ecf9dedf6e1f82d55a2eb61dc4be263ca10ccc
z77e4b58f001898257e55bec62f0ba30ef4fa98821ac19fc87dfcd260049e2c318a3799bbb31c01
zd616849b5a0f8d3b892caa3eb4e626f34554ef7ea08585b1ebfb3b39fdb1fffc8a694b1e1416e1
z22f74291a3a318b88776b841d516cda34e5f3435da57b84c330d7c731d7cf114b677c207f05b87
z6ea6ca3bbe16104fc191792c3f6b26eaebf3759626ebd2b9b11d7858447154ae7804c4d380e248
zeb2bd31ebd3e6c0a0b0f8c41539788c2faa896daa335539da33785091fef6816705e104bfb4228
zbfea7e3d79b532add48943395fa0d46e8fefb0c31ab2141a06c10fe5c2473102dfeeb24cb61b01
z3d6034ecca6f9d21795048bd37a72ccee7cbd261968addd874df8fc501f4e84897f5779419c935
zf8ceb0c860f3fc3e2f8f860bd46582b9be0ded1a5dc195e6a256bd924595741d39574fc3d8648d
za30448e2eeab39aa33223b339baf2791242720604b3ec4d742ffeb458645f5d77a27863ff23b5f
ze19162d93419c20024b1e7e5fdc62878e21c88cc00a43a802a6be32ec06922d674b8d0f0a02e12
zfc5d43a591a0102692d862f9c2a874a3479c1cdcebb5ee51f6c9af91d4e939593d753a6447ea69
z3f91a1ec7fe19cbf145b7809b0ad7df9cd2c41a57edccdc632489462526309a541dbc5afc01f10
za8266d0ed9cfc327285142db68c6719bc155250ea802feb69ade539ef08a3e437a17c67309f9fb
zc8cbdc846744b32c8f62f6bc997382a6591cfe4433c454d295de4a32c5f1ad5a56e1d9a96b5644
z16a41cb8cd18df68cecf06c119a2e0e8988e1d548804d84cda039d097b3bec76fd7fb97e80c023
z9837c39cabb60e45856720aaf569affb58a8703ceabc9ba4be8185e572868d36a2d0ff81107eea
z3ff3b1e5f4b6e0b820ac67f1be7a489b5af2d521ab262fc4e147137350ca0c9d11ddb245b340a4
z8b8c22d8eab97b7770d66eb856d5584fd65d7d71995bd0408c1580c644478e556a1b6df99d4987
z0cca4963695222f209f8181198cf66fc2e2b7abc375f729dc9656cafcd56e5a4b65faf78df8f99
z933d128d95353b41a84c08ab836f9499821370db6f7255a8f7825eb556e7ccdcbda832fbe03b10
zce2a8e777cdc5be397b37c390bc11666b8d0235f1ab3c1c82b0e474a797908eccdda44d4c6aefc
zd1b3ad33b00e25bcee12d4706f57bd883817fd8f6056c802606d7d8d76674cc4e817a445f56039
z32df36ea9f4b574d10f2029534dab57398684ae5ff7acbf366f1cfdb90ef3dbdc9beec23c0c09a
z9333d068b87ed6674f8ca2b17f9257ebd20270e1e2fc03648dfd1b4ec624bcfc576b3bb65160e3
z3602e6aa8eed40f5b1fc059a9ee4a91835f725c45a6b14fc1e7f6aa88220fd8906d7da6a7e83a2
z589aeb8c4ea89a551334e248c6187b48afc47b8a688c95fb927fd68871a1a6a50f502c25e35dc6
z36b4db293a14a51b323ef84f34421efb177a04d5b87b6b0237fe95d784dfe0e51afc52f35b010b
zae18d634508d5e498bea271d467d765cbaf23f9fa372c05b6bc98d29899907e7c1bfaef76e1ffa
z2c61a18d3f9f914077c5e9794764c0233d59dcf6895cc51f09cd56f3cc2d0c50b8aa34f03d516b
zcd5dc49cce35b9d591b2b989b6a88751895aa47d0ddf7a559790275a3ff7d3c9007cf7a661ce57
zb16715d51c7aeebece68cd7a459d6d1f240f9a00ca0964c77f810ca5fdadc6b45244839dfc2b88
zcd49681832b220ce18c89573c7838a9dc356a3a25a90e0fe9a5595e38f409e2ff1fad1fc170f0e
z9fba58977c228531009027bf763572b69f1787cc90f12792103fc2ffaf0c33cb27145ca119fdbe
z9f38a1481ae8da2b50fdbf392ce9efe0796604e9775b306d12d7adb6610c4df660332ba2b27b67
z49a45474ef8a4bd6713fa2d9113fab0e0efd19b3817a01481eac56cfbef2f8c26be2fc1ed635fc
z847085a8c976c998c3e29d6a864c91d24b4583e1191f0227dec6ac4095d90c239c80ec4e1b3182
z46695d5c28ddc6c2a5ca4e4b9384ccb214496676d4dece855bbee305d1d80ad4256219fde618fa
ze034e3b68749b1ba9626080923c410c612a8797b7ed06f0720b33398e58b2e372144e3ebf8fe12
z4696df17f5a58d64819ace1db88b5215a66a5ffe85180e0ea6af6a828ca0ded81d215ef1679568
z5733af74dca88f953d3bd5eb7d68e9a8cee90e9b4384c4273d7d9a6f75b437823701b5467cd73b
za7c4e230988b174ff9c3d98497abdbfae8471a27265e2d95297632114221ef540ab2ed0e85ecdd
zcab767ac82aee04f8393b85768dc39cff259444df19f98a7d9f8118746f3da064bc580767207f7
z70eaae5b7807b6574a505de47a5b4fed08274b7dc6435afb0c9a5cf5f4e820eac22e8509c142a0
z3e26311c133655bb99b935178e12bcbb84cb04d7dbe08ecf9711c5e9f59ece2aa75d5e9783cebe
z98c128fcaca0d6661bdf606d805004a584031f5ae2fc4748b5cc64173db5c95ce6985993b3fa39
z9905640904a626c0fd5ca51bec3f4d3be95814f5014e4864d8ff3673a29788fce72345c94043f8
z4baab47a7cd7817cd97669ee6c87452b8cf1d5a9f23bdbe384393dfc51cb5da6fa117e1602af32
zb59060e3eb6710c429563428a005cb24284cac9e00db8b9e94072352a15ec7d103a1d96d177d88
zf1fa5f9550498bb0a822d275cc496e3c25c9012cf0e09fce6da0f5d6591f146a6321274f3737d8
zc2993ace30666a11e06bbf3e5e6b34964e641cdf15f68703fd541afca5dc4de556042e2b4bba24
zacc43da4797126489f3f5147739feccc2ea438d492e530af4a54c324155bf96396315d99d9111f
zc021e745e78270855844de8f011be3efc2a01e84672a903fcfca7f0d1d3d0558dbe3470799ad27
z0e90a76eba0499d67b49ded87c6e9367166806b2b6bd0f14474da6d93d4c70ab5162482f6ad43d
z7ae861bedb9affd4c27802e84261ec3ad00f21fb0304e8ea84a4468038e0feba4703784855c9e1
z8630dcaded7764aec0c177e9991642e9230ce81b936d3660f0fff9bf75a02c58e4d865dccd231d
z12a235e99c2b59b7c8b219d2b3a6cbc811b94b7af0ab7531b958fd4346b68268f2472c443e5afc
z2a1686d365420f5d63c7f879c0e184c5e568fba92a6b496bc8b34d43ac4c6ed64a96c97d32983f
zdd69c12cb4b261ab827f856b37e2cfab0d704d083ba14fe37c4ba81563a99e944892479e802934
zc7a27f1e7d5bb25451cfbfb94af416b6c6d8f756d0f656c92c73115618d33b7dc2233ff17f0bb3
zb18ae0fb8d5c5da98460f964711bec7bb813d5ba12e12c31f8d796f831a80c7ba1cfe975b1482c
zd04bae9ddc5aee5929070e66cf56680308f77fb237265cbde23ff9264646cecb3e98382d6047e7
z2720e95b8e861eef35dbf74fd85f05bfc82b1b08c3b40e1fb4c123e44bd2fa4c826f1e68ce02e0
z42bc5f43a18783046911bc314d7bcdb1a652a4414efe98a7ab1e7cafc0bc59b384399026ddc339
z0aa632f4a61bdcc2efc8fe329bfe32b689a305723e09f6536253620f2a1d43821624fea2a79e74
z4fca56e4e0c5d64304711f8ac14f930ebd4ce5e9c8e20781609bb87b04e5b883c3e0aabf9678ef
zdc294ca54262659df1a1e2a2d4274331d043cc31c5cb0dde0509ae745beff5252d81b570933f3f
z7e5c4b567e472afc50fa402453ef1d5838143352fc1c8b84ba988b0fc7a94ed6855afbdca70236
zed35f23974dbb34d92a18f4425cc65cd70520823631a2bb688440c9e363893db67bd9973dafa53
z3ed4c81fd12937f2cc8985a8577aa4d3a218aa343004bc268be5e9549e8e73218fbe5166a44d8d
z19805ad5e57cf3bc50b93db4bdcb9f6f079c807ab749be7db53c1d321e3bf2767bad4ef7e2964f
zc7316936d1885f48c32cecff3d48da49862ee943527923ba58a48e5f3b112e5c5d241fc0226c3b
z109daaf8093fe24c729507f425cb13e58f2e94f2a9c9c1a2e062ad970ee51f9ba9e5133c08caf0
za2d601f781fd0f864d997b9b9339eebab5b35f77886046509e7921d5c2579c27173f3e0a4800a2
zfc3d717e144b0ff9218a03c4f166cd2e27e9f54468fb15567c1e432a12914d6699210dbe446a6f
z3e9808e4613b95780996bab6f056f19f16a3b3598b11b0244121021fe2cd02de206f893b3b2e68
zc5c4ed1d069041ff955faf879ef6a3a90fa3e41e5092ca2b4e131401824f48203bb3194bf5eed9
zdcdad7f93377812bdb537d861fcdb0205f91aab2d5cbc3aab84504096c113d237ee70926cbd35c
z80ce2b2813193afd2ce550ca6287e9ed20679b5a598743b9754392b2212a807f8bab6bbaf1ff6b
ze441bd6090b82dac6601a45f1329e330e1c9c88f1a57a917d701c8bf98374ab217db98acef59f5
z3bb88ea11f6934344caf1049a90ea2f334c2ce7bb9a0eb1a30136c6239face1d9aff82768cebcd
z424158a38866c9169cf39b39a828f285ff6c2a0a698cbcb05179675083e6141fc44f20e156292e
ze7f8caf0ea8374ee059a6800046f419f10cbebf9f658c3d97c71c8cd8953a3f3732afb029998b0
z3237be5e6c5a975342cf77867d1ebc524a0930e484af8f86a9aa03716dcba00ff06dee5658ccc5
z904b7231c8b3bc1a0181176797adbe81b07aa1529e0ce9322a66e01b3cd2dab8546fa724c06aef
z9956e6a1f5fed8e8fbd352bb2cb8f002f4e23a7d57f1572dfb2cd4593a85a726bc26b560b38897
z34be9b4f5bf825db34f00aeed355a08b08fce50cd6c19bf5a69d2a0dc5af89f3c197a8cf4e3eba
z9e33fc51046c25ab52a739f82cd126e24b8b1b9c5344edd393b7a60e78f3a86c0dfa7a3bdebf53
z7ed96a640f64136954df348bdf9ad8b89eaf2dbc6b5b5074468037a4decfc751434a1462e1fef5
z83ff765539786c51e1c237a889a072a1a6c8186fe9421482dace210e4b9e75bd07c55458407ee2
z19a85bdf4b303423500d5efab47d6b219ffefb8906538428c6baad458e511275b7ee29fe0a3dd1
z8178815979fbd36106dd3f7d77c6483e3038204868c6c5c03f79072c6252360b0c8e80c0b5d5de
zba35616f38f54d8f920bf11f29b719958b5e16eaa0be506b67baaaa4b037461c4c35adcc74f4a2
zc9303f368a24f50c92b85c8c7df3381dbaf8aa8c55db4c46ac9404a32a9abe6beea4299c2116fa
z43f07b6a0f7ecb597b537c4cf710258fde5b64d75ad3fa2af3bc93060dca79bc76e873f9cd26ee
z0944e9294a7aba1bb7d55bf141bcec6482215e73bd6d67d6feff15e696a35e529f699283070121
zee5c0728098dd4ec54f4617523746012ff18aff313d79537c1798c3326bf1d7018e904cadc384a
zb02ab5311cc99059234197e8806b05dac0e8529d43ba171548f2eef0fe29a1879eb75ba582c032
z120f3ff6bba5d7cb8531377cd639b63cfbe4076fd2d8d02360a4e5973626f8ca81cde5289ee0c3
z8e55f5b5ddaffe11eb061c83c620b24924a3dee70acaf3e2cc228a635c037966fa7c2fa12ce03b
z95c585cac20e32c6a7da42b87bfcbd33e20c33549446867ae0d893b4a59cf86dbb0d000d176d1d
z72ab988256b3a73eac5dc7b15fc1a4db054e5efe765bbb05d4b5119ea348a30d9e0fd8b77c7d3b
za7be2cb0ed27f216596f7953ec88734e7e0d8defd8a6e24bc98d4fb4fcf6f107e18b7c7dd234ab
z9bb8684bda091fc4de4d9fc192d89bd7dd2c2cc1952f7bdf013308398b1d4c3abfe85df001e89f
z090bc12e65b1ebbf2713e6b40b5415bbe581524d8c35d557661e2542207b563a59cd43d8c2e4fd
zd37f8874d0cb655e211e6f5061abcb28a46c049ddfa419166e4abd38f08ac351159cf9e6ac059f
ze29ec219ffed5d62ee767d39fb7954aea1308bffe62cf42ada07fa77687488ef0a23acb14bd215
z85f9390a6918b461dcae1997877a6e3175f68249ed14b1fc945d3c8e5e434316c356a566e93b5e
zf9082297d893afcc27945bcbbf749a976b0229f558346c086dd6fd41f55128e6b75dfc384df30c
z13f2e775068e42b1e66b78041da756e2f6f158dbe9142d92e3c67aaa933bf9bf62c37d6cfce60d
zd7d7e7f88f8e43c02868c1a6eccc25e1ff5c520b5da3f5492e074f4206d240c5cd6f083beb7a65
zd994162bbcfd903d7a7b236a7ae018f4e55b8617368f813ace8c037bdc4627ae95213f96e95f82
zb7bc1fd65b2b06ffb85e0c5260c1e1b8eba1775d4718e6d9f0e22c45c4a58f8fad6e6d965e6970
z49178d989be48409d64a7b3e51d817316992263fd9ebfaefb4681188cc3097ec91d370425a2472
z063a8cabfbb211c0753fa38ff24e7af76e901b76df31ff5234605092b3a29d1678b460c710edd9
z259152d69064ed70f2cc9c4288e4589f76a35bd762e53227479c283322fbaea523c7a605338076
z18be9a897ee1a3c4a2d29bf9ec3f468ee4a11428b552b2c89dc9c4f3676a805f744108187d21e4
zfc73161a45af61cdc04846fdcd5da148ab240a64382d70bebaccc85f87ab10236ec29bd10717ab
zddbb69f6b5de5f1e6df7ebba24d812f7454498e26d9eaa9f2624d95704a1c04ea75785ca17874d
z6c8f510a26b546d46520c1a29bcd6e329491276b2766ea05498029f71018e4c85b672db8e81930
z304d34b043456a8e8d7e9dc0f9c66efbea353c738e2eeeef24aaef69215d7284ba1c85db9fb490
z79ed5ca4e438307cf63eae8626997a226e2cae388fd9459e89181a94b1cf0d9783716fd96dd879
z4eb31ca076694c55b111883e9b983abf53a2b2b21aca4627c7a3fece05f4b862546321bcc66918
z8a45889f3263bcfd815cff3d7ae8f17c3dd827e821b900b016ac1384941edfa31db67d2d9eb581
zdedaf780378ca1031273c3bb0b254421df00f8cea7ab41e1223079335603863c49ee31af764365
zf14584436a34cf15b4dae2d0e34791ad624f4dd9c71bd5caa0bf860d26a2279e703b0816016c8a
ze7255ff59646f6e1302dd23fa8942e482d516c8eb7eca5bb6d8db9eb878dabe8141691e66c83dc
zce37c5c12fa419fe4f6c44d80ad4c0fafef429de6c785f35165ec24c34778a2abf62f1300f91d2
z8f3fadb37fa5ea899fbab4630b1a55651c254ce6113634ad2b0afe99b013471fa5dfb9ea7955de
zd969471c670d70f3463e196a50986cf57d177715e915723fc6f724e8595289cbaf608bdc2290b0
z66f3d539f46f5629cd1cac73aeaff0ece2c64ec925c3f4ab85e5f8de644dca42600e4a8a7a4bd7
z3082fab85d13a1f2f101a1bc6b48945e1812ece748ad820ebd4cfd0e3740b01c9749661a96f004
za8d17e3ed45811fe0d0f3d6338d44b0b700551e75d663e5d651488128f00f619e25766d0e1e92e
zf60c715d9cebab32b4525cfd347035865d2a523fb6b02c07db7959d2b7fc2d96c59f5c21aa6bbb
z9759d47a88d30b8eaa45e8a822300c877416abc3909112517ca87337411f463cb1afdddeba6955
zc3322b227b8cd5d778ea8f5a1accc7633032c56689f5b475616528c03c561aa23891c89b499fba
z8cac5430403394c9883725c78f55df6b2edb8f79870aa9999c45c3e74998f7fc1f34899935fc70
z366dea97f8749ab995d8bf9af0fc116f0f330be4303c2b00ccd12e904863db3cdfd6bfdb107f48
ze5a6f1625c0ee4cd75cf57f117f4f689980f10f0013bfbca580b63f833b199ba6998165199ab6e
z677e8f6ca5574f572f517a73a09cca4fe2b3566dee88e56fae297ca61bae6618c8d9b0a9063ccc
z4b8ae1a911eaff64c5dd5f77f2bf086db7f88502a2c556ddbd173957d6579e8ac0d4e5054670f7
ze24e7d8c6d08cdf4353eb739829164f5818e111189ad7f9187a6794a7e74c61952c6d9b7f162a8
z04724fba82e6569fb581230ff48c80001250bcb18b83b61c766e235ca93dfc3367a04b119044fe
z87e1d88f8bc9182bf1ff6b791a001c4c2ddcb05cc701393427188b9a838ecbbc4ca90a08ef553e
zc52b79d7156b4d18722c29b2bcb59f71deb23cf5f48ec296e5730e2e041f271bf361a1d337de3b
z4937fd11c1f28179d88ea6b330ee07e91ad92ac1d1574d4d332391d75daf27c840a83ffcd104e7
z9d69b2ba0755859d55b630a372473f7d69cdc6e1115e4d4f8db5448f49e64acf56df0604e41f34
zdb48a64850683f5512e4d3cbaeb0a64d3537c5a747922fc828252cf65a2e2a37fc4504178aad97
z048493f235aabd4d61851b1e33819f04043816234cf7bddf20db4c1b6ec3a4c587bb183028dcd9
z17e17293fba56d01b23e44fbccb8037b3e945689ca63f370e2a1505f650acc604272c2faadd44c
zec421e83ecc7c09e36c9d454d171fadac020a0bbe4de8a02bdeb0eb2b47e63a947901a3ac40e5d
z451b56e9fede1ff9e4f7262a908165e7f82c6ede2b47c897d11bcb7321edb1bc60b3f5795feed9
z452f22ffdd9d2b48da04fb1fce00b05cbf2513b21e417a1699669fbf2ea92069e2068912754215
za895fe8903297f439c67366abde685be9ed803b3d2410ca7acce8d9d6b2fcd17f050195aec77f1
z853fe8621744f8e8e3281a13081049171f82af696c42c260e242c9c72b459e10db6f78ec9adeec
za275618339ea868ce6e1b372da77a5949b785ecc31142ca2f5e714d90f12600ec48d0397169840
z830290465d94d729d7c2fde318821bdf77df67874bb3c483c0f314a35fa214078fe1f24f944810
zb27cddd42b40bb1c6ad9f6ca65a6d01b1fb47078a2e86e857c54d9721bb9e45aacc8d44de4f0d4
zc9e22fb7391eaab4d6c99541eb7ca61ae1623bc20fce1e906d37c6ad7b81fa24c25c0ad05752fa
zdce32e2342f78c5e8475845a0e0478f04e75b9c805b0b7d80f10ed83805e8a39ca4d6b3f588ca4
z171144a2fcaf82021b53c7d3596892e8c0ab5df1e90d1eaa7cb5ea9281f91a33b0225f0cddb60c
zf9e39a09bd4ac53dfa9a9d8404f685257e8f25045b76b76f932fdd8fb781b2379bed12783789eb
zdbc85eb53551219646118180aea1c1562fc9100a18d458432d819f1a639778c0540a8bb44d1668
ze3a7aff42fe8f802d5731488ae3c9cce0955e3cf9d2ad85f07f427ae6b0a5962eeeffd26879de1
z9d0ab260a5f9c7fb0d3e9aa1c4b5fbbaa5cd877b8c35372f147aba66b5ed90f69aec2909dd0264
z00231a6eda226a40c351936a9e5e3416de30e8e186c89b089ebe4d95a6746681fe8810df992701
z79de4f576aebe9e5fc818ecf3db7a90365103a020f10a7931f439eebe5c31dee2b5a6e49c5744e
z1035e3fa14152cdbe05f93bc6f7487b81058b9392c36bd999e776bc8a952c39b3cf4066421afbf
z6cbb40183a740663e64556ae3cf935a29bb581703fd77bff68c862d2df58da9c0971b7b4556e4c
z575fbb309df47806ebf60b30d1ea72efd7c2028d4f43067fba57b86dca056285f76c0a6990270d
ze4f7872ba38a9f43e76a5104183a795962597068a6cbf51bb730ec158b03cd273b4736f2c274d1
z543bf9562ab412f58fce287d98ece51c1df02879830214d15dcabab3a2e2c4b551c95b3bd04c34
z23e5c7ccf011a7f894efbc58440dd700cdc3e8fd1e112d82bc515d534d7991b9b2b928f9432bff
zb1abb45867b839f356e4f612c2e634c1de8542403bd945044b14fdcfe6d6bc53269851cd8a6581
z4c65d48424df9ce77b4205b92d128a20c2d3189542ab8a12370cc815b06b9f2778b60e5491add0
z282450774cc682ca5764adce4ff02f35abc7ac50eeb034d0b3776479691f0313d3025e495ccfed
zb10140b2e4684adee0ca1042601fd1b39ac391170a18e2a0a36d4b9b5df4027e90646159dee16a
z98ec2b30372a66f24b2c288ca9ccb12b7314360959add61418ea78d0739b78b1d4455dce21cf7b
zee6bc3216f40b610c3b0d86f20ca1eb640fc3fffd7f93c6c10f15e8cea4359a3ea226fd5fb43bd
zaec105cbec6d89d9ccc2d2971bb199aba0d42bb237b9531a21ca7203607b44ba2fd26a550ba15f
z04d5faab3bf77ad71535ca2fd915b4e3b617e381f0893abdc018e9621f37b1a5b5cb14061ba238
z11292d53cb884c8245afd0e83166ef7ca86e44a2a23bddfbfc196f6a46c012a591b493a6fad1b8
zbf7ee02454a7c363683d66aa5bb1f95174c56e51c75abc889febc0506b17016c586893cb4c6b94
zb1a762eedf151e471c682bd5364c987e25d51a059b14027ba916d79c63ab0496d16e05e25c9cc1
z530f2297077f8e8e134d4532afb1524f82f9933a0aeb36b2ec167878307a34f7c4dfab80fc49e2
z7642f7af9359b7e417375a8d441543e05820187cb6319639f486137a1fe2501312ed38f18246b6
z187a189efb46f8091d4bf18ecf57ebe29b5d474e131a3fc60871cb87ba2b450b6f89b8513de45a
z28d7530d3b8d9b55ac9d80c2f839777882082412d3b5c0ddf02bf83cfb6c3c6403e04db8c7e99e
z8bb63395e51804607383c1ce4f5fcd9bffba7cf3543970bedbe6dda4f2525c5a9f39c3c5985e89
ze81099195d36e10cca94fcf6f7f817fdc1a2e5b540b58471a4a9b25abbb637da2a9a59f1ff9b9f
z845df3c59382f41441c2d977290cefbaacbba44e98009068f2ff5ef9290666ec7e8bd07fac9427
zef54bd333d1bc056566f8e07b38f94cb858ef058bc1ea74c7dff02a2ae9ec80861b745ee0d997b
z09d388694b605fdb33995d05105cd2bdce9d98b936a06970ca34ec26e8b3cff00a937428ac9581
zefdea6bd39faa061871b621314635f21312b0f735a19a90ed76dc869c24d0bdf9fe1bd349e21aa
z3b1ce5650d9b7dc0ad634020583c3390435c132689440d53409f8c906ecc9781cb15da0604963d
ze869414e41fa8ea938b66755136e3ff2df80885aa4b168a7ef6b73bd5d4c6120560e3546a41083
zffcb926a547995df1025d5a23d16d388873ba8dc87f9b277736105338707c8e45bc537939c2d14
z201b09df9b1b4ae471378574b81d58ceaeda9e5900c545bd9d3f145205a5ae7ddc4ac75f4d32ef
z1dec1f68773cd3ed8cd22691570de161ddf0a1c71dcd7a8c3f114bca9a81da1a5550f33ef00346
z8be81bfa807842f27ca53a3dea297cc0963af0ab328485b635426c972a4c4295935616bc3973a1
z72f3f1e9f88305d6189691359a167884681d0e3f0a21be21e74e1f2a210d337151cbe373abc0ee
z6fb8d7cc29e2453b84fa792c248857ae68eac4677e4f08340837be298500bb49048ed106558136
z1c86a0119f2fe8b0370312452797eb32b451af229578f1a0c9300f09bb73cdc1af495f9c451ae9
z7fa43eb514b77634fc2f630bdcc64e262836a4f8905b6d4cc2f7597af421e71d8d220ee40c21de
z45a4a36beb84e180bfe70a7060e51e7f848d29f0520b53241322e21606a409bfbb8bd641c61a18
z4f7800360f85d3271fb78f8134bce5dbcea74cec2cf964b68bcb400a540f757b844c76ad69a5e0
zc3bb0e8b131be8948b57a3c85e57bbc5684f8663cfe13170ea9ad2e123fdf43c601917b00d54ce
zf00e9d5a29f41741e732212ddcfe091bb5b4fbbffa36e6c92e87f421c882d9511412795b029a7b
zdfabb30c0f5a0cfada067188476b415d53948be93ebf587b2cf900a8bae511503229afacb3d9e0
z4cdcba652f4094d2cd5cfdc278dc3f5c834ed59712f57b6d5968224c5ac4dbe2b44ed826d68951
zebf2b010d78db1d6bdaebc25ee52ec4c6bc16c28dbf22fa0f650a815a5e3fa34423e208f0b43d6
z0a1f979fa033acadab27a86db9e78d648814a58e794a1f379475b7400e94f235243b5653112172
z10f26b483a5540692339d33b4ca9ea79610e6a16d31770e27546ccb9ed24b6deaa5e4ae75f5340
z8b4e7d88a4954676c62c60173ea0c2c90aac210336cc475cae0a0104d367abcd567e93b2a592b4
z485605e5c49f4d51b984a7d5d4784226c39236c48fd7b096054ace01136c4093a504e86aceab81
z3677e33f2698b9608bf5e76b7f4c13acdfa560e93422a76a3b6d50e5d4019038156f0756b195db
z6917d8a4d14c088c5ad84376a430098bf3b2c7b034df7982aef2232110f68abc7fb51831cb537b
z33ed78565642d73e601d3072aacb6e6ac355d74f1b344e5398ddb4ce417ef0d7854c96f5cb457f
z1f759a65daf1be6ee999992b03fb1898afa136f2a4470482e9e194d64347a72b6528a0a63fa6dc
zd1de3500ab79dad88f0cd5fa77e3059ed438ec182a29def1c72ce70b78a77357a9152ed0e8fd12
z9ccdff6b3257f13fdb452a50786101c70885086690ac3383f7d707285042e4455bad9a443d26f4
ze5807e9cab3ee83e02ed10e9cbc23e16eb435d3eba0f1fe7b20b1407073196963cf80aa624eda0
z56517f8a149ff61eb22759597b534f7860578ea9ed1b7fa770259cb4fc28352cb8ced1181857fb
zddf23292ec4c0b56e9a1d0f86e48f54ac53068e49c03d0f31e471dc479c314008269689a91ea2a
z2c98c5ace0df1495f86fa4fecc576555c355141416f8eb342470b5f591c4f8f793036b07529133
z552a1747d8c034d2204388e1cc095d50337d1b7684b34d71f97586aeb3d8aef639bdc69db5c150
z19e58aedf54f9d7fc76ca43715a0be25d1611fae8e2da2f673a4e2bcc1d7976decf1236df12e72
zec6f4192daa11184cb01fde03bd5e16179bf55ea78375ffa48f05dd4603d205e2df5e6e34544a4
zdb5b991071d7a4e7880fdb1ff922f88f80fde79c50db8d33e78ca669305845a1097c110af7829d
zcd58bdccf48c14e6c8f066e04a41a8ce11e3725dbd09b56f2e3ba33f9ba1b485d4eb3460b23710
z8577e925847e9667bf951d56e036c0093bfd4d5ceef10f71debba85a3ec13bd30c20dd8726399c
zb97c2e3b79edd65ee3475fef0eec5f71ce5dd89f247f62b45784aa7fd7a21387828af692b72640
zf7ffa1c8679329ad0dd9b0a99c1e2bb74fe9a5be54b9e5b365a966ac9ac2911d9b2ac605cbaf6c
z780d1c24a73380af514b1e90fdc931134968283525fc3be3965f3ae729a5de97aba7daab618d78
z3d6765a08cc59b6321ee8b0dbe25c824e8ef1ddb4679bcc25d632f89d458692099edeab8ed07a7
z332762a6efcd1e82f55a54e275d1454643a544b91de19517faeb033dfd3b8197443dbad284efb1
z14acbccc250a1ccd4d93e3612118eaf39df122e44b9cb20a6525c2157d98cdabd41fc0be26a310
zb7aa8a36e8356bd494fad65a0609d4a91a914735dd863ba1559d2f42a977bd9c8d483fc479ee2b
zc3d5db9f1515e7820278af070fb8a7474766915aa7329ad00147aa13c6a371feea3b1a66f2e18d
zf12d08afb1086db26dd9f940b78124cf53e890dd89f664f3d27e792abccb4003f32c583c169ad7
z7d2a33cd488ea735bf3c77aa62268a478ef8875c32b95e9157894c3fd0cf8c29f1c9e5d20980af
ze9c18aeb036e38fb8fb98f8734ed4b144b076d29c7bed26517afedfe2bfcbdc7ed5388ab2bc047
z73f39673691689a7a102c6c88f263bbb8112468dd91227cdc6ffc773f18db9b8176f3c4df9aedf
z9b1703b282241948edca2d8b1be354e39322486bcd5e7d0dc6f74dff36f1aaf544d6d3881f3d2c
z9af3fe9ccf7a0632378eb67a3fb62fe424777d1108d6c03c63c4ec064319ec6149ac0198f550ad
z81af4497f7a739bfd026984b5d3fd40827676ab6d3f80dc9c828cd981be010df94af1bdcd095cd
z67e2ad02b91217a6eeac6358fff7e852458cfed8f68800a3e29aeb906f5ec4e8e3d54830759334
zb8069dddcba1b6acf8b8d7fafb9da993fc2882bcf03530f9a567139e51703218d80651c1bc0798
z3499e67fd95bd2a2c080d87b8e2d85e33a20dac3c8a15489a6c3cc0358d0ce1bdd890739930ee0
z2100e2bd72888a28187b509253eedf82a9aae60beb1b4b2545812616618be34664a13462641ebc
z563dd409b990842491adb7a49a1f32fc4fefb370cdc9136819f1f4cc1d25e8e270d66b5a2a5f83
z5ec4e3795257bfff94e43402cbb0e3e8c71dc8c42756e526c0670524fdb77b0d181302478ecd26
zdd33de6395c81dcedc9d280264b36d840f0c39d44be262d486d3f8eb3a6f9ce95882d4354c1595
za98a0f54d34f32fe40d7b77cf833fa5810b11f3754d299fe898e347066d39c1693dd4ece2422ac
z63b21b349f46a4ce10a87a5fcd0f3d9aa93d0e1d972b0c2fd8def6c8823c1e8091b85b53e97d37
zc9bc85248d3fed7e739d676754b81e917bfd6989020104a26ded033b4f2bec9869a03d9c44d9bc
za2e90c54f2739eddc2401e7ce66f01ea34174e05b2193682a5e798d72bfb660d7854a4563a3382
z278a81884922c3500a5422944106d5af34d4aafc188f508f7f4a2fcc41d2b7a65c5e397442d692
zbc17a5a972ed5742a8798e62c268f21373a555648d3e8a16919665451520e6730c6ca268decd93
z0736a78872e2d0fa8313b33fed288c30fa6342182ad14784eead85bad80329ac31f4476a412487
z448b21d99b0c6a16b0639211e4119cb344b16291019cae4d815e1bcc7e92cdd80f3e9dc2513570
z8eb23f3cc5117e80ca67f0fff5e358bac1a7523721f661e06bcab20e20f109ed0bba95be58203c
zed24bbe7d9b311305c44bf1abe82319cfdc094cf9d615cdc9c78eaeb2ef08d87e687975acacf5c
zd8d42da4cdbae0c03c566fd9a0c6f7cd6d2c41101a43bba7ddefd99cf9b1efdfa8c59b16cffc39
z525002b0140e5634bb748e43d1c5595e60362ee133ab7648161266dede8a8a13ea31d86c2dc1b6
z1ad8e2af1a9db38584c97aedd32b3427d2a0a01120ff959324c9e91b76c851619295d5b7bc028c
z4d38df69dbd941b6c88f463b8ea7286b7c0e16a0654beb329cf23f209101e06d9e6c82a744bf70
ze030b04638858f399feded90f8f8a4001108d94da1dafa9b8b1da15d8d822751ad328690eeac5d
z57c4882f16312656509d9dde26f34ef5c7eb27b365efe6fd3506e406f3f33ff8860c8220f2d76d
zfc091bb44b500411fb16f3ca8eee394c132dcc4e4a08d51a7f7485f0a82f58b2d9095dfe2bae91
z4429f98d046439e06e685ce12a68aac4d8ec20fc028e9da9cfe77f98a48d942e96c244f1572ea4
z9bc6d7fe1e48708521d357a1a89817f2e65ced2c5fe0607e35d4e66db6e77b9a4e2b38062491af
zb7937d3123acca5992bd5531c67633e90316ca291315a3aefba2c24baacdcf2833114fe7507b4c
zedc1f9211c78a3aeab9392997e4459bcf7b766cd9cff7776481549d112d2d38815d719aaeef1f7
z3e61e356a306035edf963e04110ad8640fab57e2ce8106d0973eadb4d5d1c2e041b817bfd9a9dc
z4b8987819474264b58282951b0076377dffccda4e7555c949ed56269af0a83e0f347ecbde96679
z6da9237f86154145febca5f600bbd15ce15aa19550f831d47581a93606163783c0c91de03b2788
z55a525ecbbe8e056b421ad9cc6c9d2b4b48a6056d42927d8d0fad06049c5def53e501c68418588
z254ff101432990c3e23809825fbff4cfe9d4e4bba290ae7964f7a59a158110f973ca5e492cb2af
zdf5370f49e86297968027f3b95f1490a4ffdf6feecbd007240880f32ede1e2b88bb5b91b434753
z20a24a6ac266a1695a2e3dca2c2f7530555ce49872078a59a0155b6b62a85e4965dfa80a51304b
z0b564eb597387aa73819f012274bd79bdbedae574953ae80b591185cdabb9fc9a39ddd1b108be3
z066ff6832fcb16e9186dd6939ce72319840fd9824fde3e40d08c595ac582a5b8bddeaebbb2cdf0
z92f143c9e436f41d6c3dc1c532bfcd5aa1b1f509f2658ff3f324853a877a75fd0f5df56729b51b
z84147b4a448af847696bd5322074f7894a2199447693f9e72412b4625a46eb6c28d77f4aedbebe
z023fa635160f39fdd61036a5d161ac3c06ea764ef6f01d32286fedfb377b966ec2f0c87a8508a4
z39ab078a8bab3c5d2babeed0f893017cd6859de93ab8539d36027d4e501da2678f3e804bbc44b3
z10848722e188c73cf891e3dc543c6ac68cc47805678323cb722ff2726f6db0d7e4e065a684b7e9
za513532220b95c4307a4711304b599945e777aae3ad7100de1b4f93df320a1d4b7b876af64e1bf
zdd34007aa19ce2de3dd33ec360dc27e350c2199b48d23f39073dbee15d8dd852a5ea0e52eed402
z8ed34057785dfecf75d840f4e770fea24657d9006336d307a9feac196d9e3f52b21560f0bb5829
z727084fa88c63f20cf5ba5d1238fc6bdaefcaa1a15bb5406401eb15bf067cee0eae58ddfd39328
zea94bee541d9c04b5a35961fc58248dfdc15cc7e7fd12bebd502613eb11e564e5060ce9fcbed76
z58c918ea780d3518d23243c2a4d65d8eeb15845f7245fb3eed433a332dbb7d10ea4c62468e947c
za596f61b374bb60bb90744f2e23532b4d0151557c0be45ddef2af7a38a060bb42e7d5ba5795b85
z7dcff181fd380d93b82e277a9ac088b22f37ad187ed9db21898080a0cb572a52560030990c8dd7
z72d672e9f5b33c01cc00f07b3356b560da64632d9ee141caba9ead72e023dc144ff84b3575fe8a
zffa470b4453145e351824ac436344c542b972e083b160a15deb2e3f07f692b40e1f02fe304a048
z2c542fac200408560b272fdef237a9c3b6792d5475ebecd4a98e624ed0e6ca464b5e7a18f51d5d
z75e83852c0ad4eecc6efa61645975e840656fbb60799711a1125651b53d7baa729fb24c8392190
z6bd1f87fd3b7664ee7fe86fb9793b20ddd05f68037dcada5402fec0e860286eb83b0a4dc630205
zfb765581c80be585ce082ab43a1b49be9934b63253a837a3268b292d01a88ed7edfc6df954c3f4
z91b643e15f808cc986258d37ece8462bf99cebcbd3bf0b77278cb0fc736b8f4ebde93b529a6f32
zfab7d0510315eaa57b297f9678769ed3a82ff5d6ebca2c5b5ce8da618f834443067ea71484e3d7
z28e371bad014caac179b940225018900381b93bb6db6116291975ca6f03abd5a152f4bb30c4b7e
z75c8ddea20f1644482ed66772f21bd5fef21c7e6b0766701a6fb47b44bd9fa8f9f2a3fff88ada1
z9fd9bb5e96aca12f89b7a0ab3741727b39a39053bc9bd84d425b19745c63e5101f960d1e50389c
z3db43a2bb250665678bb706d3089ffc478374e623da7de31fa15721c1025611c5b6999a64dfa64
zf7644ff6105c2bf7490e98a6f4fe1034aa4cc7f7ee23069e9b5dc9cfecc744d8802afc4bebc356
z7a96c81a7a1714fc0dc5104c7b1c5d08c0e81f0b8b6348e6576cd03dee15f6ff3efc23608faa7f
za80241daf743d00e718fa81a926eb144e603e645d5d937868931b823efcc501ba2e330e2e7e128
z2e5883fd8d33b7a87d8ba9211d30ad489e37a90d0d126e3c0699c6e4eaf7e55acc39bc50b424ef
z61ae60c3886c78d6a4725fcfa10207ccd4e63f3cbfae297b676f79ab1020b006d411a76908d6d6
zc1fc4ff17150386d09abf1d7d51ee231a261600b4fc2c13113de5a15ccbbbead9496e4e2a797f4
z43246a5ea9635be4b6edf459547ad13530d2a0b3e8f7c7ef14b45a3ec78796ad34acbfcadebf22
z812154b12cee33113fbc3c5d40c4daf1e4d2f98aa1b562ffe8e39049fed60ea11b565cbb6f8d31
z427648d204d665081f8c0fbe2df304c500ee84691d9ef03f67009faa19bce88cc2dc7dd45b749b
zbf35df8c977dc49175ffd4496573a740adf2180d290554db16c338a6056a1ee4c2e91106969763
z0cb767e3a4b2843db78f07a195fb4a2a14431c1f753dd56052eb7a41fc9de0e46fd3fd643ac0c4
zaed655d1c2d22945947ab64938fd3d06045bfd994cc68e9d6fd9e9f5e15bccdc33c4fed515d337
zfde71a7a290f85118427c8dd7abbccc6612c14b02b795df721080bb9a2c67b65340fec166e6149
z70e3653e00714ac1808498df3d18a18c1c81883649f7cf6580d4c7fa48e7e8c840a4b761962272
z552012c7b58df83b057c6d0bacde4108fd99839b3dd42173cbfb309ba450c4248fe7eacd9db5ba
z39d26b2936e89aafdf37df4e520603dcc02ee0cc73685c9e538ca62b664ef30b0c377f77d2fefd
z771e0f2c8d8c3838759a4f3fcb6092ae65f037576ed2df9073146893112fc71ad406f176352467
z00ffbce8ee5f90120a9d340c391957b9d03a7e301423ed669d4853e006dcf878afabab80645adb
zc42c56513d695540975142a23b9af32fd2c9dc4380f1120dedc2457e7cb6f9e491c35bd3fb7a3f
z0ceaf4211a589e33f8653f6be3aaa1e0eb863009962009ad999e896e46893eea1740077b6fc708
z8df3bbf5e53946b11eebf92876aa8985c2598ad7c5212ea219e5a2d2d358b571854010e40cc3d2
z4757948136b26e51b6100b338cd6ff1dc0f7ed5ce889dceb573a92cf6b60c4613c7c823e293ce5
z551166447284ad7a7d208070132ec0445421c48687d25642d587c7caa3b71aa71328168dd0a631
z4771854952914d9323dc8bf763378f839a07cc54048d6d61a6e9fb5139da02d27c502161d59b99
z48dcb8f7c024a7a65cfb0980fcc69ff5917605b2e3163624f941bbad6ba1a7069cd32e0c932baf
zf18ed039dd0a0ba15161102729d58169ad091798183189245ff2979c2ae6a68c4a08bb8ef5f640
zbc4fd90350619a4069fabd262039b17a2747137e5d4e631703bad6e96741d2d759b02d17b845c4
z44432eddc541a15cd9dcde4c4fd00896e2c0d134f86e69a2c960dc8594ea5036f1345ea601b307
z822948e5d098c55af449f3739be0a3255e31bb97d6056e20f62bddf747b41d42876c0ad6dc982d
z4a8023c541552bedfc3d8f5ca2f6349035632d3f6288fc886a9d10805dcc72b32234091e02d32f
zdff95d09753561ce8f5a7c2b520ab0ad82bf1f57e363956902f3e9730c2f9dd051879034e54029
zfb71dcec4120db05a2373ecc4f80391c43bd86be117c999ac859504438d52b69f32ed05a9d2919
z02aade11827a5997e0753b1d7f5bc146ba638c22c10daa4aec182400e8d8638d637af87557fe2a
z7d036e7c44c59947d5fc11521871cf452d19e0ec5aedce30f48360750212215c7cbc9523ecdeb0
zfbf9ba4030b23ce3a89d5c2358bf4f155c92b54d7f1b25477652d07c738e24422db8522f1254b8
zea544329c623a2f9ae7f14d57df6a55ca6d2978e7e724cfd4663b7ad7041f3260f2dcb7e45d829
zabab9170b7bb98223a7124b20295748b3ccb1f5c7ec32bb17eaa7d77286655020182d31b293b05
zea9b2f962a7ba5fb65ad5b065156c652ce67df58d034142fef05388b4f46b7e82c27abd6864b1d
z062d06d2f07347d135975d3c36451b35c33374bf983d79a4311f6921a05e8bb78712bc7c6c586c
z58b544768a9772ab745583fa15792d40e97ad8669f397006655ca6df0d4135a89633862e683f71
z4cfdd910e3f442f4ddf29b131424eac78d87a65ef5a7ca558638f272147a6cfd5dcc48dd6d8d60
z271469126fa89644689ece45c2a22ccf5ae0ec0381a5498e184bd1ee4e87787fbd4bae923c0f3f
z6952ac414a9c136ef0bb4533744c6b971141609e0cf3f8cc51dc6a73b4de8684ceaea0e37a1b93
zcc907128dd4ef84650f766c62e754b64ef8b0eae5e8959a1ee0132f9365f44ed802ec28eca844a
z1d54796aa0fd296c06f739846b99a778a6ff41b4af02e473e7b7c8c8fa514e5c459dc5eefea76f
z464ec0d3c8dd944c9ba714a532c46b913756ad073f2464765cc31cf872a7a6c9f8d8b4aee405a8
z3d3b5e504790e934519e501cbda5a5744cd24b0617e5bbc40087218bbfc29dab9fee58aaf6fa49
z00e771bfb7532c90a155e3e16b3e66124a6454876599c20e69c4e06d25a1fc6cdeb2887c166ca3
zbcc3a908e102b18186ae7b03cc186ef98056c6cc8ecad4764ebf833e3ea432015d579ac1a4464b
z57b86585d0e70a3af95ff9dc153a27fdb35491d246d53cc092df3bc95af78f6f16fdc40dc702a5
z38ff34fb515c4a979bec5b57cb84b0e3c08d20523598937fbeb0d91fd4bea611342dbc8615bb4b
ze5e159233d320241f78fcbb11d08a32e97703828e3b589d9c4ae6234ad94ec176b19a1396f700e
z8a242a9c45db49f566e6cfec5d4c692c8a00e844e401c3eddf1235018160bc30dc469522b87c50
zc1db0207cc7af2673f61059a456494ff5318c95da6850e68b4a2b991fb31ba1829c2268d00d8bc
z43ee01a52c2ea89ee9157fa3443490cb45f8a36864f7d4e6934eb2b2cbdf07b1622573edbd2f93
zd961db1be37fc5e2871a7b0ca6771e7e74ce1985a1a0b2f3352c8ed8ceb90376b1b448d0cc131b
zf21f9e22121615f4963d968200060958aa88f07c705d1c891aec340e8877146bc5c4552cee1870
z94da734252f35c3ff8e6068e65b9abf4ef68abf79694e6048c4e9e256d0805892113768cb205c1
z021109da94c5894490c272a45dc13259601bcea9ee45f52b7bc6fe1fb3438c65e4a66fdd33556e
zf09df1ff552bec37969ff1795b6236000db37ebdcf1309c1b58fd4f0bcc7528752d496db6bd8b6
z365a214742ff274a92bee1fd9421603de1202a49980ff05dc49fc379d49ff3b11836d2dd5121a1
z3d538856ec2083459574b296c801ee112d6b5f3c2e3b751519f1b1b901e678f9805fd6dd672026
z25fd5faa9207ef3cfc29a656031992e509e5c68418b72e6a4bc6b092c9600b27df18ddc0efb5ae
z48d769eccf8091bec24bd39dc04c767c0d3aaa22075fd3cd2eb541c1bd38e92619424c68a79a2a
z6d1b06519db53ec6838d4f4a329dfbc5288f23a22296c094e05ccea69fef71d7c9a28ff0c0d67c
z2225f36fcfa51c629ab56c6442515966f81f89c7c59b2a14427dbefdca940a76df0555f9b0d02b
z3c0a8d7d953e8887b8db1a5350e85176705223a51c72401dc07851f9003e730dba2b1da95bf581
z3e2b85eff7f7906b568cda9a7b24af0b43dabc13410a42d9eb5a2aaa4d003f568e7692dad459be
z5b1ec1cad2b704e7ea76a72aa0a3222c5ab03010120e411b2bd57bad8563d661b5b17d97e0ba67
zf335070fa62820139199b91c423aecaa4beb094a6f01582049e57bf842f8e61b2a2eca08c42b59
zf5297c36edb6e022a6bfeceb49dd441980edd2df25b672f968188ebf2a99099a9277581441f317
z7a44ffea589f4ed735d3e6b311aa8d70ae7c0aa4ab895e7b6cf19e1f8da4d493487b2168c9c20c
zcde6668722b6e8e4a660a20906a43012015710f488e687b8022f2dced7427833ea9abfedd91348
z99eaab5a526f8a7c00acf5d5c2b0631586d66136bca7a03b82b2ad8ed4030ef05a740abb4d4262
z5019ae5e089ba4864c3920b7cdcaf3fded0bcfdcb017a826a19d35bea3763c79a8a397fbf94172
z22a2809067a93c5d2412e4a212d3dd351b8dd5cbb0b7e88331bfa98099f1094958988f665e9d20
z78f56c9f75a1f45c27e6edc54cad298de263cee1f608009a88c13f8e80e2527215da00412af385
z6af86ce14b253da5a917d6359b81adc0a5f4a41522505bd997a1c8f8994966590daba922d76a57
zf04076665845aac9f374c9e8a948887d32193baaced33f755177e29bc901dc002cb09cfd1d63b7
z94dccd6b4562508ca7e022f89e6c2af6d2d022865afe66466ea3c3561ba399f70877882977239e
z6661a1c999602c3664986160f49c1ab3fdbb87adbf8fa523be9d07301221a30134069c6b0e0db7
z6cf6ec0a9b20e9a6a659e4dff37cd2649fc6155115d9748aaa6788bcb962b5695f07f8f8a2e8b8
z0357fa5a15930aba10ba5f51fcbf110829df074087da66496461baa52262231fdc69173ce3d1c2
z90fab1054d8e588a2ebc76a0ddaa1e4223c3979ad7abb87c7f738fb2c7fd73173265cf16bcd358
z8fa928420368c0a5f69366dbb47d8eee54eb34adc200867bfa3ea3bac0ff29c72410d43245c206
za01a97e449f6ae84fb692a1bf03f3720dc65f0c3bbd74fc55ea0d0ddd4287c6dfda86c0fac1a3b
zc6cb6e6da43483d192b92a89a4eaa5dc5ea898529e52a03e1d5409ec6796b6dc08cc3c0ed16a3e
z56b5dc57e30b477da57ffb811885f1dbc77906bfcd8fdc792d731555c48173bba8c5fcbfe259a7
zbb87136769ad4f0d9d3d7245ad8d858b1545b227cd17914b508506f9675cc798221a6a725f6c75
z3088f4587bef2e9709bcf3788965abc797f89edbb3a38f0544eb53078380e9ff3cf9b53bfa3f79
zf8add4167e20788013af73289865cacf01ffa421b4e72c96978609f0462a5c5d28b02bb87fdb05
z12cb0263b3672ac0dfe67df21592a1c4118fcc881f2ff372b62a86d6aa561f4f672c102c815568
z6091fb52a1d1e710f81211db67373ee47460b3ac40ee960145b274d9e98015be6147f21283ca27
z8e18bdac0d3517ae14211026443edf96598c46cf496ff31efacb576c2a2d0278687b9e8ffac3e8
ze136a7d58ab1629fbb545faa207adc09702b49884852f3615b125671760fde652bcc205d47f816
zc43d9b38c3476e574964f034de62261514b16ca1fe7208e97e4b8208c5f8b7035f65a4d7be0451
z3e2490a2283ca57c3697f5b86d8aa7ed39f1aa06e138caf81394bc98968c1ea02036c9fa823ce4
z79f236414081d7df72ea9cfbb5fb57c7614518bcbd022495fca16380cfb7a0906c0a505e093df8
z068b6580e998c1822f6a0cd93a9ee4c8cea81785b6eee23c4190ea8d2d34d55fee7c7eab94542a
zd294ab53bb775f5e6fff0844f8ef8623d29ff335300ae8e57b5a1093dc35059e120ebc1a55a4de
zff91134dee1071e39554927a8ea6df952c026c259ff0c9504cb9e3ee9a5d37eef33052fcb027e9
zeae31d14f271535d8a92d06a21ca7cc9c2a9c719366a208a90b778b1c156a5ccdc59e2be0e19ac
z6661aa9c32e5fb74a36646ec09fb1b680eb1090359c9d2836eede968be280b9bd4a931c7ab9ed8
zddd9a05c5b413ca481bf8af436375dd4214d961ccd68c781752037d943e6e6f94a032fff2ab172
zf0ac2fa339b46670f69ee29b3ec5cb1a2cda5e9479e416767e2c5c6d9a117c40017a086581ae8e
z5aadfe8bdd5f4bba6a13c51ed91d66f2a39131388ce67bce87bb553ff1073878b3f087d870bd2e
zdc747b8545779187102c450777e8dc891f415849aebefa897821f0d302c98b9d4008ad1f7ee061
ze1455b7d524f724a1bc19c77faf1dd813c19709cb2f805ad23e38941c39661760f1c151e7b7624
z9a8c940d7cbca62ffe28055423bfffe622e544642df049eb0869ccbe59c70eb17ed9fc97fb87b7
z2f145568124be7cff229004958f1a9a17da922ef7341b14b24ca466753fd3ccd8524386b2b3e86
z36039ec17175cda83afbb81ebdf620bc8d2834216d053c1f46631ca2ae1ecd650ab009ef5320a5
zadae9099ebda3a1429595b8f9dcbfb93add4aa9906591d3f01182787d804246b4704a90d0c200a
z581f815f2521171fb06972e5c66e584832bdd593c9e8ea4470371d080cadf82ee83a49ae173565
z3e7fbd39f28c203651fb02ed9fb8df318dcad14ae788557c839d37e0628ca3ef5f999deb3a53e4
zb0438e226d1fe88fdea7f0ee01f763d53edbfef42a3d0f8b4c4c6d9e3ac7a958944e2189a75b9a
z736ec3bd2d202e553b9e07065e0c146eb2c452b193771af6d1061b0a3ea7ea908131100969cb2e
z82f23e1cf4e8faf7eafc513bbcda7b1197f0c9f5a154135ab97ec4814edbd20d03e358ec8daeb7
z993a21c3cb8c9a0f30602c3752693ed21bf1eba17ca7604761e0f2f8f3cf81682cb930b6bae733
zffacadf92482bc3aa494d839515b694dc6b8f2bced35f61e6b0f9d848aed45c3968de61d4baf7b
z2ba074325e85c9b5905586235fe1f2cb6aad6d8434eb4cccada56c39a1dca8eb040f495391213d
ze7c2441df5aa56f99519a07c35f0428a10cf7c5a7b655dbd8f6c8d5da3aaa4b5a15c5d5fc503d2
z7785a5da3eacd4956b63ca8e39d414e63b582a7098dac1638e17bb4785f7cc1669ad12ae6c7469
z4ebe8d25033c5eb096e630481a38dcbbc5955ef369e8ef4c07d911a37b2207fd7c2f25180cb7bb
zd237502d77614e8fe962bcfd6dc53e5e17536aa6dd450432d5d6474fcebf2353d72eb2e08d5e1b
zfa82d3b17e1437a4b5ebf02964e36e0d85780d7a9b8a94ff7d2e3b2dfcd2f3f1bca433769aa790
za59a4a904ed354747b5c95590294a83b745a04a8a3d9a634156b11d4d94a05ec21904c465bd539
z5d87b114cd2a667c1642347e28740854c4cd10b943fff946c8042055a7c4b49c4c8a5f0b08e30e
zbe1548e14d69d85b46e0cd3cff48ff37915f7527b4ff3baed4e78fed165c3fe588b07fb4f42dfc
z3be6aa56a77c7c4283655ddbb369700d3957cbdc6334f8c1729702ff95651f1f1b610b279fa1dc
z3794f84ec15253d2be3c5d1b5d11478bcbc61c5e993b7b10d3766bed9384182c59172a466339f0
za530778ac5d12cb80e9db837126b2deb204a9818bfa321c64f8a1ed7077f6a3919abdc410f214b
z98ba7d4cb6701ec2cbe88102ba3fb3b39bbb49b1bbac1fb3c07bba3990539fedb3e7d14abfe0c2
zbe3680b299708288abacf0891be0df020e725a8ce85fbbca9939557cf34da346cecd9984e20a08
z11e4aadc954a8a5af6c913d4fb95e05dfe51e2b1a73adc3a7ad059759e1241643b48ed7e7772ec
zaa98f8c20ad727486a9f6e1258cda9b03bf0a3528cc5d40828ca169729dea6f0d6e17b2609a117
zb4fdbf0f51d3391536ee699745ed47bc37f02ba450bc839f748bef5634907c3d51da6665f13b89
z79f320f1a19b88a41d4596901b0f185ee926570b57edaf43983aa785d65a38ac65c80fab072cc3
zd6b1569fa1535270e25b16ba56fec02f7d9f037db55ee03a2817f2e4d9882bb1531ef344091451
z54f231fca4383d7067129affe993b710b06348b8b7da5f39ee81155d8e56c71afaa801088e176c
z6aa190731aa31437212c9d9e642381f863b4c07cb562f0657c11a76e874d111f395676e2bde4f0
z57c63b1e0e8e4badd69566dc6433eabd0d1bbf942fb707fa8c2d90b83a204ad79ff2a31c4c8a64
z8526edf597c92f22ebcc2a8b3bce09a6881da0d3da3449ff3615b2b9ef0eec96c9090398e80cda
z1d21d078dd840ba4192fbf3d92f27b3698e20a02daba780b0cca489af1df3741cb667a9f0bbea1
zec74e5c2d98bc72391cf7ed9a966c02567e36f80d2025d7218bfa6f381d580df7e667bebba7828
z7794fa351a604d1aea46fcafe2be2849b41f61ebf17e42dccad6aa43fd1b4fbe3bcda67f1498b1
z4e943318d767e8ef3cd076cfff07c5eca5ca4a7205f0e8ae6b4fd28eebd18c84bf33427dd805ca
z5df029bd21ff2c0f416169a6f65b6c93ac5cbed407d8de3ec4a7056a15c9a6386bac532911495a
z04dc121d81e57dd7154c37a6314aff2f7d65515077a87015a26e48b0047cabfdadbaa6cb49d327
zb11892e1dc4af86d24d6f7930f7519956822d5d8ca077304dbdadad31b762d5ec18e6b6eef4ae6
z0375c44ea17e7d9739b2ac2349538b07bb8a3acd8a5b7ec4419c1bc9813534f11a8452134e1aea
zc314af6ad40780d2066ca6394b118670987292fcb329a3b3cecca435f16eab983dc4cb5dc57ba1
z4271ce1412776fabb844e12ae3b9f7ebeff2c504a50bab9a336a24f8ffafad5a0f424177c66413
z775341acd4e2bc3a93dae5d81600b2d68bf937929373757ffe6089d0b0837f05ac536879a3ff9c
z66d52adc0fd9d89113beb38647d59d77781e2c53e132ec4d4ffe6906c9916f4a348ebf78586756
zdcbc8e44f50a1837508130b8c9520da5aa2e96dbeec93dd9d0d12ee62a468a7be4f95a4ff67503
zb90f4f5323d0e72ac52a9d7c7f19dcbbc35238cda36fc72385752ed6515010997a213a5c254c67
z39b9bf38cfd95e1a5b685516203d2311dc8eae82d0c8e26d139d0111afaf5e6c0fd76834399311
z01dd38bacbbfd55c150eac54fc3b8bc75dcbfb7f4d9aa6f97e0339887d2afa4152dab1b09650cc
zd3d87f3f85a7de2909bb8967f81fe22c8075e21e997da402f951cba64c100c6b522f48b80d70cd
z3cf2eca55f8ced6287f1e710c6f74b69bce49e55b4d8bd805f0ff3c661e0a4cd042cd52bcfe4f6
z1f206ac1a66809430c287c4ca94945ae9331aaa51b1f141587352e64fac3de4b1b5d1c39cb1083
z6703a1005fa232e33020ffe8cde91ab9d963b08475fdbf61735b3efd5f40644e729271cf52e849
za0f28f0e038d3b07a6647fb18eb25a97634a445309669f7dc9897867826863671bac856edbdd42
z4e2aec14032ef03fb63875d67d9ab002d251dd62fc95daf6bbd645a5c6c5b8b0a54b158c6ccff0
zdf1956859e18697a98e75b88bc65df4a30e59b31d45a9f9869134a5c35905936edcb5f19c2be00
z9f7aba69271ed0905fa082e8dc771d976a5d88693659b86d3a95f3f4a38a471d47de9f806fdb5b
zbc809884cfe5e1f5eca22d0535bd552ef2b3adb3dc20623f44f842c5b65f2bba48c6bb41403999
zdef0b6e8cd68fbd0d53150b741a2b7ddf1aebe797af117e60d63eb7b3aab5ee0e8e00f04832a89
z9d6169858f1537dcd9e383b5faf1cd716f794617a989eef7d6ed604cd739cb6cdb4edf460fd43f
z94fa352b224b63cae6160fa094ad4fe778c4ab93cba57bae2ef3c46438ccdeb05c5005183596fd
z4b3ebe6bed490a9cc3b4ac1730cce973f87a0ee8d20ea05077cf6efeba280534e6728a98b61c4c
zd9e684956d78a8167a5c365f86774f5f68a31f2d5ad4e51048b098f1f29e39524050bb2a89e835
zbaa4454baea5bfa58fba5d2f751c9f54b2a2965bf6ef7a113f737ffc6301b000c95d4d580c14cc
z03e8b190da330c52f9c6352d806090826fb93c51b591b73064e2c6ae4903870754f912a13461f6
z15d5212bde7840752a88e3b825d63fe53a23e88d57f6fa7cb4d1426f1a80577e52f51cd3755695
zb6a4891c07bc97366ed005bdc01b125def2c464dc2462902e3efd554414fdff5b2f75b1c6e47bc
z3bc7d655b5698d97b937b5bd3ed08d9305e58429e9ed90b5bbc1bdb7bb912c83905bb16501a941
z8da66dfd7891ab452d6606ead2202ac65cec29207494504c7678bf79c35187ad9b3446f1432dfe
zc1e938403a3e898ce249cfdfcaa5a20201cb35982bb5fca562cdb0ab257f8f58eca2300849ab02
zfa4dfa72be83195da82302a82792ca2c0c5db0496316cd15dd38007ff362c6d4cb9bbe80522255
ze371ec9e8049e8eaafecab21199c3b493a38f48c7889d6d0ed78edd4ab7907507397625f41053c
zb50ee7b416905d5a4789835b5a9400ceeaaa7c5203cce02bc26d76abb0d367be45cf0134becf6f
z26b09dd05bd3d4ca4f6c2ecb31d27c3f64b9cff1a2bc38af1f37b09ec2a6ec2e536ff91e88d884
z075dcd3e50075cffe376fb5135e0cf609c1a1c9e090b37d8ce53343a4ce018c7494e918efc5775
z476e0e821aea1e8c79e836055d3af03d2e1733df839c7361f6537c131e957dd9fb4f010b414e43
zf37e6ed43360ce549ea2799b96398e4fe37cf73173f323fccc24dbbf1bd82b275f74df372e77f3
zcd45f865689c8f8d5debb09b628b8148255b4ed7ddc73013b9ce4a077dc0684a8f1997f1df6d56
z913eaf768bc492622c4ade6f0ae91d6daa54a39090a91c2b0c7d7b12736abe640ea0faaef28535
z52fb86a48f3f5f1fb81e0a25cf87ac8b8fb36b54eef454e8d7bddd6a8967bd798b68a733d2e88a
z38120fbb309608b58245442a4f02868852bfbd8460ff7fce6b7b0787cc92fb71f1fad77822f104
z49feda97dc0fbb9c426a5b16ff9f13add907e987a65d62a71f9700dc3393f29e80d7e1ce45af15
zda10d418324e67aea55c92c59d4e91e61753fe62823635081ce1550aa52169285b05af114292f0
z73627e52d594ca7d47731716ed94def02e417fd2368bd5466ad78cffcd8e3c8597171139b0ba39
z515a40b865ab51c3de7dbd9c9437d2ca8e1996a34dc58c13bdffc5d813686c304d362d4c4187c3
z9fb6bcd82098edac19f952ef7b88b55fb694a4a112e038c5dfac7758ecfb1dd897f4f9e3c167c0
z9d15b4b5ec250fc3f0859444f26383b805c0f303e154be7091e68c4d1961a07757fb4d105ad450
z8f14fbaa335bcae6a5f5bb4c497d6929b7093417130143c662a28c449890dd34e6d989036e15fe
z22ebeca18b46f2f5c25a9fbf7d3df282200de9e1f5f393ba0581fc60ab9069d6df3a55c60fea8a
z0ab24ba92553ba33b3f009dcc887ecc7e49bef03297762f26d8ada6cc2d24ef18f2e676affeb27
z80a5b067e790b3e48c9edd3ef8dbca225739e22642d7a1c5d819e607c6fb492e1c2152dbed38d6
ze018ab6c804bcaa5262bf8ee7440d1de1eda99749d4714e45a9c5d322c455b294cba08e7c7df0b
z20e0d0d050a01672abb8e1f410453f3890b2c4385eb864792335d1d5b146237182bc4074df7817
zbfd74d66a5448ebdfabb9be50252e44730e6152d93a4b1b251789c1b55454a4cce7f5494dddd01
z7e5baca0e0932c49f212ca6b5e37d2f78e1468a156557b32557242aa0f4c63093ec0ae6e632352
z09d8a476531736a51e165df63d20dbc708afa39b515f597701779578bf8711eb7f58be755cd51f
z1995aca239d3a8df73228aec540dd3658da3832c71d9687deb8d3c96848055d4eac08c9d224528
za232082849d2812411db78bb2a68a6662f8cdc755bc23a6bb5a26536a65ede743a0ad16ea52fa2
zf6db6dc8efee56d52c5fb5d2e00a61eb3fdb915139c28776e2d29ab4d08c7beb416b37c866a6cb
zaa3db15bca181be22c9bfc6a221d1e6cf1e68dd4b34f0092451b2b4db53d4c103999e6835faca8
zcb124b772400320b9f9f930e2c1cb54253df6c7fbaa99f44af1bf61daf9d8711cb1cde532395ca
za8797d0e278440230346d690b83abbc9de2bd7154eb4c4690aec67b7398b6769a48948512c23a0
z61ffb8bd72facf65ede041f7d1d6b88793481831049baaea9a86bf6c68a4684c1aeaa21765e476
z16c9943782860b6c643ebe6fa65ccc63eae0fc12f2fc395294aa9fd255b31a84543e7d9cb30e74
z8be851ce0635e48e862ca6b9b2e8d63d5230891671ad07db73080114c2c47757b2d3eb7b4199bd
z73921b812b704cab1e724cc19725dcdd037f684c058a321029824e360f141e45c8269f31557f6d
z7ba60b0a20d5a6f69361f3b8476dad78a703ec53b15bb55c980a6253d21433a7186345c4ef829e
z3dd35b127614dda1b4e5621dc448ffbfd5451b910a5e7fdb51f7713042b0cd75037003779578ca
z5a1f25ed889ce143292af35ff0e596272848f8d1215f1f64128cd7cc6deb0c6280a46b8d1c6008
z4d6560c5c1e6ab89eaba5e68aa3bd936ac362d7bec3f3bba802c2cdcb3ca260dfda1e98496fdb4
zf5813e93aa0f7d5f1b00c8c467cedffdb608fef4a0cfec4f88ac06d20e515a0bb2b27b6dc8f2df
z258a177e9a5d3493f0b4ec5d60967542693097138084153c59020c422d8922ca4bffbc41d4eb9c
zbbb7229a06621a822df3eb9b84da1fb3ae8968f78e38486baf1cba8ae73879bd244efd83c6c876
z79c75154d7df34fb789fe761a1db4f2e0206fa69a852b9b82a7b27a1ae356ccf34aaa5e74ea376
z2f13a6cd2945d1db380f310b2c5400383a504a63670ee735d3ce30d4f10c8f42c567e30b800940
zc69e5a57590122c7fda193662ff50dc6de6ceeffbf752adc85f610d67c76baaa3c6574d612400f
zbbe21cd9793cfdeeb8d244c548737b68c949cc5038e8fb8b2d0263d5d7310907df57ea98989a89
z378738c5a5715d6904d11e85560e010f9fd3eb18feb398d4f59cd323fe61eafe3a0893f03ba6b4
z08a9353459f67566b04027776f47351cce3dec30837167ec684f6ac130228ac14913e431a66cd9
z2bac303771eb9f5e43237f14530dd743598272397eceac2dc6663797db2fde3b107cac5b636f8d
za8aace09485f74208f1facec84db3fe5b026a8dea791f7454c0474c4056501691bd28cc8c1ef92
za04cac626cfb82d121281215819b74dca19610575303b80c3f10f22d89973bdbe7c08e62166ff7
z8939b990648f63314f738ad0852784e3e473efeec3244748c55d7c988bc5d53652de592b37c61c
zddae493ac04e0fa4ff1f1563e3f70012c356df0dbb8c7b605f7355a24f4c62fb9e9811bdccc61f
z9143cb63ead5d22b516a3239add31dd2675b39df0b053ebdb37c0a4b7281c3f9fc19d16ddfca6a
z4e1fc27136ecdb006a9dffb5daf6bdb82c574c28f3e0ed69b75903b1b57ac08919e9866c3787a0
z8bba7662042ab449ae3a5170df56153e231e53b82ae947ea7c9190485667dff129adaee038e4cb
z53562a094a402de9855caf2855effc2a15b63678dc4ab62a7fbfc97a02d52ac8fd631488b47f6b
z22ef4f6136b4b3bb5f5c2c9f6dee3c224658d5135d37064e5a5f410d4f5306f2a9dfc2ef05d6ae
zaa98485f5fc6292b088d79a1ad5892de4d7c4b17b9c5a910db7d1a638901adfb3038837b70bf20
z03645fc486b4909e52151748f61fcda1da0cdf3c564754703aa3a84c92c58d25809c98785ff0ba
z0c32f35a5c8a299baac477008ae4ffacfc440f8c406b7e01766d4def5fa32d639178a4a666e39b
ze4c8168e65b1c232f5be626bc7db5cce0163ef9fad25b0961836cf29e8d1f21347877a87cb6105
z912b8d70ba8290f7e3e0cd0a7fd53a92b22abb5bd2ab122a312888f4b9fb40baa93e7b5307badf
z5ae8f0fc16c5ad880d13239354d9801d1927c8c84f199d7ecde04edc9f82ca93e0b986f4f9f28a
z014378a3df12d8569d073781c2399b4d120910ef792770e2e564b152ce3bd3cadf2c005f4eb1a2
z2fab268cec8a42057c51953a8a4e27f02cb1e3c6a58446cf7359889e9c2da4b819f04c87f4ccb9
zb73c89fe5c3d01e65fca1a120524f2d2fe1bc37017f103f6bccc6c00e854821a5378292ed392d4
zaa48af2f057152b80b75beb8c8145105f418765f4eb8d105c4414f40ef725a710cd4492e8ef83f
z260a5c92a0d6af52d8916e82ce0cdc36042d036d6eb0a6bc00e7771aee30f8c00506f7381f8351
zc17435fb144404fbb054665d7f48b94b477c2938925332cbd84fe3864a07f90d7b2449349d555f
z05e5ff093f3aaf7b23dcf36d17cac960d914d4b223c7d2ff10c9edeab5251cbdda22fbeadd4905
z6ceb327567aaae1ddb8deb9e08a3e413f644fba06004f346cfe750ce853701541a1bc2b2ecb77a
zf742ed810e31a2df06b9b9cca65a354ce7c5bf2636094fadcd8bd7cb9dd23291cb61693be8c5e5
z859b4af5d2207f1ba6fa8cdac98f20368d626efd8211468390daff0356563f38d586b88c476429
z246067c0560e1995025761ad451f66e81c8bb9517ad973afb74f6d6c5db9f97ad1b4e66b088fce
z015ce9c46debe07cd529e0caa6d8cd82802b95679d787f926cca5a290016faeb5f6313bc4fb185
z197cae21ff6f5d9e7a11896f10dee743b19973a6761532deca975821c5bbbe1c8a8032646d9756
z71de0e3c17c62f5c91b447225a5dc981a0fee414db426b7fee056a76cb08f0e3023a8c35569509
z888034efb84207fabfd56e7e36ffe07dbd771be746ab79a3cc8f3e736d426f9b6dc816a721f7fa
zd0a0b266f7e21170dc3a9982fbfb709dd1deb59dbe2b994ebb924e5a6f3c6a5298a6ea34f27b5b
z2b21ebb8a46d91717700d72c8c1156ec98469b1d93e7e0d2c3959d94dff2098fbd62eb5059b839
z76b23b7e32bacf55069690b5c4d0bfebaea1c9b88c9b6e7ca816a18adb703f09fa654fb2551243
z45b5d2fb8b1e3fc290d071a1ffbc1ae0896ead0fde7770158dfd02b8ad731420c8b1d2436daaed
zf0a21a88533c2670ca3ce69ae8e5dc0844036aa147ea59a22a8bfd4a23bf6fc97b3517f5872a81
z14590bb07e4a720a8fd7588576247ac1a69e8b087fb0130d55d06f59a0ad785f65cf09d2513c69
zab02e2350dffecc52279e908d1d995a0ac13ab958a20130059c9520d100ed77ee2da37097a5a95
zc90c4872b024f5b431372822f722e89989a92341a1751bf5a932203cdd3c1f846727583ebe5681
z432fe0cd0f3ffd873415d3cfceeec014e3dccdf9f31d9ff8a72af0e89affd32165f07216a8967f
z7e42216245e4a29bb400cf0083275b9e324a86641504b3d014522ba11acdcb4e041bbd59d0894e
zffff50e7a2b604e47aa66dd76547606242dbc6b05dceaf371b41afa3a006015ee02fa90a8ed08f
z2d7d4ec1f64034f966359ef4aaab600d38f98fb6be448e72d93ac296bc71a39aaff737ae484071
z5760e56fb49397370ec6049efd8eea14a3301f9df4610f1c1d39786cd8f59bfa6b425a8a8f9cfc
zfbcdc56e62f1868c2b4148abebea8b7dda32f87dc77280ab9fc29c23d8fd3884b5b319191277f2
z0db4e3e1a253204ae9fbd463a5a7fb909922e7625f6c83adf2344dc99d2fe5531abf9bdfb03823
z7add1c278efb6e52d079f8f44e3eff5dc6726d4ffa16e143be8e3d8a471ea992f8e624b6a12a26
z174c1861505fd21587bc2177daaf6c523a7220aed82d2a9529ac6cef22e81cce6b00b20d298fc1
z687c3a1a841c8f9df46895747be50fc0b0d51d7f031a5fb563656ce208ff0bb398bd902c70656c
z2bb30f6d9de025063cc69ae90c4ed62996e3fc2a66193d091afdb6bd7f06d7180fd736d8e6335f
z41710902d9b52a54e780d414ec3dc58b3840de79bee6d5ad289be80bbdd929f9825ae056dccfd8
zda21a471082dd8b504c50d28194861df9b00125563e7b5b5cc8d105723a4ab41f4a0a31f3248b8
z87a1fde0c412d4139c4b3e90b3e0683273208cd0d8166bbf77900aaa7a943f59762609b566492c
ze7c79758356358587d0e22b325d041968a860df3b3f19afd04674e55ef12beee274eb049699c7f
zbeb020808d21e68dc1bda2c7d6be1966ab4259f8845a5b93cf76edfe8e9f4dc24c3e081f99edef
z2678931d1cc37044a7faa3c278a44ae795ca1cb355cf2e6ae8dae08ba06b69a1452de35b9e6ba2
z4e843bf9972446d8060947de9d8bd64d13384f81fab068cf9871b74deed5898528ae98bf16ca76
ze1ee268a909a5d9bdc47cd0a384ba81c3df7bc76870bd9fa6eda3a68e663925b7dd84a49417715
za005944a7b6bdaaa98e5d3a97cde932c5c41a9129a129c9fea53c861eb637d0c3af7c2dc96a7ef
z4dc7fb2bdcedf7ad8d68540e814d75279848fd3e1a3b82daf486a94117dbe4e0b029979399ecc7
z71cc7a2b7e845b9c03dcaafe559173e0b4d709d699ebe01259c5c4649f68bda8aaabfb94a6eb32
z276f88493e4d04976c0382a488e1a83932d01150df85dcfa1d201dd52c11cd3e465dc86429d542
z864cb574cee47b500189d3b1e06c0910d697a3dd95b414d02eef3c854af710fee332360028da29
zaa64277b9b02095698e7211bfb31373d53c8d7713f21cc77344ddeeb2bfa674216f82e5f63b15b
z3d0b101a3d0d0a2c220eddae54dbff5a972b23c4e486ccefbda7c6979ac0893d8818ac3b3be47a
zfa82dc3675f55439ef622f32ab09e39f0164206d8cfc4ff8d00cf9fba6aaea36ff9d7add1f99fd
z08457de16154104719697b45887df47854b8e8c2b27d07aab4de9790d593d2dfefc383e712caa3
zba8eec7bd7d18bc1b391754b596b61a3215de3bf4306e717ce7763d396aa74d0b63222c43c76f7
z4852ce0fe03dc57c18db8c0ef6d64470caacad68999e7672fcde22562cf41531a62b296c5b405b
z366776b981106e23924ff647e4d3ea0f118f6b25a0a4ffba97629367e951de4f1acff3e2f84366
z58da12245d123db1ac2a59476aa98e5750f929af092cd8ba8e8899ac912c65ddf6cb5ce954fc5a
z6bcabbcbcbec5ea7a5d7222a0b44726500807e5a17296ad3e3096f0ec808df6bd6f263c35c76f2
z2b73f08b9a3bd464133dd8b9d810d58266f9d8d5f9627f8772072b2af3a0cec5014fdb8e79446b
z085f0ef97399777d076debe4a5060ff2f8a83777d2cb58809858ccb3b6da315e457de992f872d2
zc0eb92dec9281043b9e04311e6d562217a4b33f7ddeffa9e27252759c14f7961d4cb9a193c2677
z324092b3b78d7f874f54d817c781f96a862f66a3f56fb0ae43b57640f359e5d443369b101740cd
z6118d52a779b07fdf6b6bdd19afea10f451726f02188820c1e877767e65ab6e345c3370cd41738
z5a0fbdf28bd031ccc4fbecef9466518739603405a083107178a5db67d39de0244be382d56f0e7f
z2ea1e1f772b4425aec7be0c50c7c36304ffc199ce548d8c7f5ea377165deb494b6a0a964db90c3
z962b71aeb6b8caaf3d362bd557dccfe0d186c5e7707a37ee0a4a1763942583c650e66ec38f810e
z96f04c31a53ad238f2319d345c9ed3bd3a2e4b4b69efc1893713b4c8c68cb357c299324ef1dba9
zd3216311e2784c577ac14b1a7805eb7bd5e9c1f3316a44be1c5be230bae1c6a1bd0d33bdcafb77
z9e45bae62c212721edd2aad8bc5cf4dd0c75bd8ea8acd1ef81b12aaf60c3586b7452986366dcde
zd878ffbd40c706b572dd01276f77575dacd2f26dc88ab75aad91224c9c927c24e32b312d19aa70
z5087732bccb0ca1501f78cece3fdf2baff6bbd35b467297be28730501d4053a9764730c3d0711a
z9e0ced6b53f30f3fe1d36bf882953336ed9d860aa4d2fe2d494e16ce53ff1f5b04498338564f76
z3f7ac17738916fa75fcc966681433f36c0c4ea9d8ffbfe582c1a5537a6d7617d60f6bda7a467e4
zcaa521091f2fa062473a885e1a44d5f59b03c92add12f62e303ac47a361a9a892460af7c72559e
z6f056948f164407eac1fbec1ff010b59c8e2cd90658bb410ca686670462ed867e5b1c9975555df
zfe09853e5bc59051e12c006b29dfad202660abb38e58395a1feeb1e890325c94595e2e32afe8c3
z5a0071de173cc970c0d1ad85b20d190ad327a42ed99c7edbfe06e5554b3cced0e753af6dc82873
zb8478f01f73684fca28994e06078e83b4477011513c6b17b47900cc197c76074711c3e54b8cd20
z7af3874c8b9c6a28d1730ccd08589484911dee0870117d12fa7cae9ffbee92ce9370909cb72e30
ze77ae0074229c9224a5b4add39100bbd01f9fcee7d1be3f1c30d7ade549b2872396af175721475
z2a80a59a8df0f5b1d77d4f86eb017498b97e0b270c01533bb92dfd6a7e26797c1f73d7002fc4af
z21c419d9620a9d5a619793753b309abc956676c0754393f032cd60a8f7afe100f174a165543097
z9e32e3a61683a97a5e0e619218fcf2280257c85ae348b832afef731c25a2901ce1199914970351
ze965434aecd89b8861cd41bcb5d5f097df1a7b0c625322e17ac4ef74faaf0020df403dd00f3604
z24794481f4a7d40d6f200e9c75575da671be0ec6c04826d1bb85a013fd01d0fa3f63e9d95512af
z5a9c51251ce48450e83117fa4b2774e9ba9d3db1f70d061307fa1ce56180ad5c3e6198c83d7f5c
z6a8e0cefd32e365e643b2e1a0637bfb46ee0830349b51429a99f423ed441fadf047a293f6d2797
z63d61d93e53bd43862dda8c63600a89643a1ca67fea8ecacfcb0fb921974e57cbfa5a031968f12
zec970b0c2580eac4def6d10cfae3abb1bfe9861e10b869294695da476a086a921664005d289a2a
z77ae079d5bf110a9e73e4041fbd75a194a288052024753eb1f9f41acd6fa3b2b04a596b13d4d8f
zc7567fa53fdccbc22d352d2bf7c143ec33c9b9310a0686e124b1eb8c7f470f6b6d320484375e0e
ze284c538457f7626de0829971820211ed7bd6fd9bb713de4f49df35e84f2b3da07469f03236414
zad5c3024d4e79c166179dd57e422ad90c223157b5fc8066129ca60c6b3aa874f74884f56b3493c
zf49f7787723a341ae17decfbf9c0e84c5746cf6246b892cf4c8a3adb4e48a805733fe0db77e983
zece39962348865e9d19610b1d3684c4698506b32ed53afe16f009c28e241823aa215bbcdea6680
z35fc75398410b08665869c6ae90691d85d75532dc88b78cd1ac9b3d99a38ea7f787c612be717b2
zd58d5f183e44fdbb67ef25a75325d66901c8eb638942a873079e73a898399c1529619f9405bfa8
z70d59d9af1365e82e6a07042c3528a1afa849277b72d167e290fe5d214b3cfe07363ae97f0df2b
z164ce39ff47ce32085d4a819d6617c91ad0f85de183eb8a1703640609c22d7690d7df783fbe4b6
z9b037dfa7685dcff7bf7d9b628545c3103ed14ceaf10a424cf603301e5dbd1e4b2efb7e04d8c07
zbe9ad4c8ed4ff13c7e926ccf2c99db9eba4a74590344542fd2dc250b3ad01e2c9384df352e8b55
zddd6d461dc3bdd196fc8347262b160949ae8409c6748a57046f5fa8bbef0fcbd1f8eedf4a15a43
zd2c671d33d257ab46e7e41e01afd559f395adf87888f0b164ff2d12c5ecc1b3dd93373428c8bcd
z2dc678130890fc3fa7954840a699efc4404874692e251c200a8df642926a3713ff95c46ed317ff
z837a1b8aea3657aee2a5369258da44ca1d3dca91ed6825a6c84fa7d0ebfd9dabc3e777362f85fd
zae618066bebf49c139e5e716c126731104aee04e51bffc64d3d417ded9d0ac8020071b6f35e34c
z29f886625c1c1d21f624ced64511fb2ad8f2d22eb457ded0111bf65b2402152456429240d70255
z9b148ba989933befb83c82e72eef0bd9407f82ad41ce72b16a80942c48bc97a11fc6f705780df6
z1883efcaf90ef7c95448b4879696feeec173cc99e66f362f674b20dcfeb927568da55dc9eb9d55
z737434a79063df491d8d5f08c0c18d6c8231276061f904938aeb80587d4ca59b8f43718110fa76
z9cc37b863cffe09c664c94171fe2fef8cd992d1d839941cb6531be0b511df9a0e920ee782e4a1e
z11e7cfe5c6704d5ce47d67623c0f371f43b1552cd861b73b1e913ad5187bd9eeeb1ff46d663457
z865dd5e9c5ddd4f46d9ae736ddc2d93eaf7197d944823a141673fde24a2140ab823e4e234ab596
z4a64dba160f39e637ae3f1ccf76e99c83209c3efea9dccc8f0e0939583a756fe78a7f2f9875fad
zd3295ee4efef3907a4e441ea9293babb70579bdc03cc60014b3b0c6baeeb4f4602251d3ba6bd0d
z8835fd6aa155805298f6e875fb984ff9f3b5a639a14c30f91ed89ff78490670d5423d42bb95c21
zc67318e26343805027165feb991b55818166a5e0fdfc3b6d8159019461c60c818f18ecacdbf48f
z2cdb7bb9819dc39ca242ca36e5185e5e160ed858a2426da7e411dd819d327e842987994e5ee967
z97ff7c23c031498b0af2a16596ba71c9ee70fa64cb3a3e37dbb472ff742494579ec06634cb2653
zb17025573a7f32114505ce46a6f39ddb931c089718f7fee7fe01e86208dc896aab43dac8229fbb
z75698db813f758445718fa76e693b0dcb4e18121a568cdb2507a61928d172f81c3dc122a7ccd19
z9fd85de6f2656bfd038e4b9e92618e333e15aaefb2045364df8487078e4f131b65f9dbd4419885
z0592ebb47bc315039a17e8c2c35dffc20a75290b1c3e754a3d78873496e432ff68596f05a0ded3
z6609842df3fff3baab5fbded254d4e0efb0ea2dab39eee0c893a3803e46c7b879b68cf1efe5405
z38a3b7b30c3d4c0b0d92322055b0e98f960328175178f6133b98b754d778e9c5cc3deffe7b5d26
z35156fb82ef5639dbea3c24dd8652ae6656a4cd2215be122b0484f549afd604a97a7b7ca3e06fe
z53cb7f583580397d1e5d1adbc14418686bedddef207fbd6e52e9733fdb3a73613f5906b5eaffbc
zefe3da442a8d4b2ad03f396b438bacf60e132112010f8f44a65d6f5e1bc7ff1d1689eb529e9d25
z9b10dd60bf496afe301500407c611a8f4f31509876dee1aeb7c5c558c832ead7d4f73c2899226c
z21cee6045066ef3ef14bf32ef7c87376a3d3d1da46dba7ce22c39ee6e14661d837a81ec367ad91
z8ab765bbf12217b671d763747d59aac2ac574d3866d0ea83f79bd114e87633da221901b87cb3a8
z27f7597622a890609af39f526b840eecea722d615b8232403cc53d93fdfcb6d8bd56a083c6561f
zb1cbe5389c26bacea2114119503b71ec5c24fe6425eddfd3e63e251007137c7215b557735fd7cf
z5fba0a65654a747f07bd6914bcb65e63038c146b05e928d4040822e309b0f7380faedf55dbda98
zd5379dd66e69037faa64bd7c5d1413df68285663a527a4884be4cb68d872359e4c35031224d1d2
z8804bb39d6210be058c8a3815869bf6915273f06c7342f21b609fc0dbdbac35e706e5c334bca60
z98b2b3353cd534f2b31acc7097ebffd724ce704e15f9fde2ad17c930d9082d8ceef624b313b782
z82c8031aad0cd5f8b862d88e979f1be1fbc052dd63bcba364ba665740690d41a8f1bc779acb321
z786ba3e467748ff719d105c4ac97a2ce54b1df25de2f5a97b764c127c72ff8d1939ac7f6f297bc
z3c6421baf133e6be725291b617e7d9bde0bdb6688f0cd7115f3aea7108c902766b3c6e7670db3d
zcbe21a5212cb5be90ad9fce9d1b49734fb10f3cc412a19efed1bf3e3ba75d46e192d300375559a
z36b0d3371f6f17ab1d55ff75b8ae07b59b043ff3fe844467f19f4dbe5deb5ed48732f205908d41
z5762d0d386badcda5a1803451d62c3ca1ced52660c418e547ecaba04a4adaeb829641305865a8f
z172f9937ec172f9e8ace214aec77ca64c4a92286f003657bf716532ca953ee1c4131976a50aa94
z2f75df2d4b95f49efedba336701a05e8587ff05dc8555db9ba9a8c20d6740c289107061f3a17c4
zedb7700f66772d37878d690cb529e1a52f13f06066e709d86fe6820204b071c7c0740a7eab60b2
z9cef543461e2089ddf44caba4511b7b3f01498e60f52220d8e330bc14c5553dbd2c4dd14d58030
zede57ddb95b27263064b6c019fd3ac731c99bf6e220920c3f6b0406aabf5f27ae6f1ec225eeb2d
z2105273544da6f0541fe52bf171ddb54fadb40b6a85c19ad7d6d9ef5c1c937f084914afc30baa4
z78ea07bb7a79a051a4ff31615bed1bf4e1beabb8820756c293b3ffbbe3d683025c836ac2d105b5
zb94d159def16df5c8204e94ccadc126977b50224d825763e6798b62d0c85512c2bbcf037968f28
zcc12a723e84250edcc2dd56a0b37a6e1eff25ac5bf1b3f2653068f03aea6f65a14715caae3ee73
z4ac9fedb238485722e576446749d007af410412fd942e065b8e3193bae4a632688a034819738df
z3eb7689e96fd85e5163cb15b7200ad8434d8d282791dcef3e9b166b86c869d7579e5873551c73b
z3738ffee4b0673dc09e1c78ac528c4b9122255be709851aae5ee040f9c156eff8c9834b88765d4
zccdd9ad3f4ebeda396f45d11d7da303e99283d61c6086c2625b5156b2e1e1faa28f6607ec38f62
z852a42b35ecad7ec6680b41a15ada13ca91f0e583a10473e44a91c8f2521ab2ac48871cf973651
z8f1ac331eaf07ef0527ccfe5c9baad545420914fae2d5ef4e8e64e66e3bf53e77e636f1fabddef
zc5968047d9bccbae4a43a5ceb79da709a96383e217b13db140febb44f852f03bc2d8ef17754212
z98ebdd85a716a20d88ec16922310fd16c5be85fbce167299aa5e9b608ed12b7c31f67d34283c6e
z2202f6261b8231554c4c35def67f2177841b58d792ab792663c1e4ddc7d36b038f3a108e4a85c3
z69d3a74495f3b15691c9aa4b6a77dc670b8a22c3ce3cc46581bd046e0803b29017d757f5b3a1b5
z9044220fb83288c1390a71c4b32ac25edcfcfe4cf7ea1bbf1d413bb7a7c1035320382c84569fb7
zc58cfc30a39e1229c8dbf3ac0121dbf0652a17f98cb8f76e5b71bdd2e64793dc0db62e640c6711
z0ef53da3d9dd8753db24584651f706ac2d2dca62633a5c91728a89d08e28852f708d3de777ced0
z230c2c4d4226fb2266ad840525b338a00a251d28cd6228633fb9a9c2572d56941ab1196c358983
z001ca6c62307421c1388ad560abfdb3880360023cec3ef19f762d273d7e553665331e95b6a5596
z7f93d7cef518365573c188517a8b3177d930151abbb38eb557842e37d8b2952a04fdf024332f92
zf26426300f0021598256d6187e251d0bdc87d0dfb4ee463d7d25e42bc8b935c2f77dda37b14718
zd056f56dc2e7bbd142624c37c82f55fc0ef55dbd520068139724b1813a3300ba0a6540138c8722
zcd43cd723f712f9ce1227c6c03bedec986d3b8b69c7a7234d7ef59f16111624998d04c55b6c1af
z7c31496a9bce383de696497768345e104c90d16f74b1438b9badbde20c71b36d3f56dc21cddfab
z2c1491079a85608102d4d557eea97d9865635dd7ead014e3445396881e6e6c5ef18f448ef0c2d0
z7ab5c94f0a5960a19fcda59fef4a9dfd0dcf77f3016c0b7f55de4510862a8bffccb9afe54266c3
z409eec7c227d48714fdfde33aad6bc2f2a4637b5bf3d30f694d88e6ca3e412ca56b6fe31fddf5d
z397119583a1fe8b1a3803a3291f2db1e7e5fa5336673c6781ff0dc47d61f534b0cb7fd0d5991a9
zd2e81f80dd6f2c8b7b1e6331626fcb592bde52ae109fe964dbc0fe7f0896313feda0e7757b78fe
z015af0a569b9dcb97ba73636f843cb4e23f2cda9bb41337c38b52190f1888b7a67da36420c35e8
zc32a36e596e592b0c14b84192e65a2e1795cf59d8dae88fdaf93d315a783b8ef1ced1f7f7bc9b1
zb7f4bd7337769e081fae77d6ab7f1cc678b8643f4b23aebe6ee90565fc2fc59f7a771deea53490
z9aab1f4e0d1438c62e18f1e5e045707f9e8178c8a6f9ecbd0a966d3f56bc8d23f1b141d3ebccec
z0ff04eae9c3f2a82419480f56d6cda684e104d9d9dede5403f979c31388d099c9c2a9c8d8fdded
z35c1dad6b7d56883a3962f23a5be78482261fa9dc46f1b275829c12eff3c4f6f81c0f9e3be3de6
z0ce62e7aa99b40927b0fb0047eb0776c8f1270159d8fe6314ce927eb69ff19e2d722c99a3178be
zaec753bb54424339893f10b82c6251bef231280111ef80f2117fc285c010008fc9b8f08297bbab
z5378494004cdb7ae9c1f07eaec6742b5689e4f44e359ed50b72286548f5edf8c4e84859d1f64c8
zd318c0b52e21fba3fdf9b4c8815643b3386c638946004ca40c7331ce9e7d4b079813bca6a067c6
z8d01bb9a19b32ece903cec821d020fa0f194bc0b6f1320f55379145d7533d8ae507910b4fe4163
z1757a3d9849f701364ba8ca9ac1a605e2b7617f58c0d366ee43a7bfb416db804bbd0eed793f144
z1e62eab493526c85c6d8136e857b2a98053e95ff9dd428af0b707c3fbd38a61312867d0b09d8de
zbdf2aa651bf5c4975bef0f76045bd63a037ee4518ab91bc2b1863869945b52ba68300833d58ef6
z2eea438367bac382f8a2ba66708da3b8f9f2d73e68ab4640be76edf2c03d003e8e6a207a705aca
z511951d0c840577313307bd5b6b09cdb5b420ce74c16364542ffc1286b7d7e392236d7a7ea5082
z75e1c4bda475490e1bdc8c9268a28cd4affb9eec6fb39ed2e2d411544956f147f869f94377bda2
zb34e1faea62e4f7f221a62907729ca1c1747eea6690c31903d59716ad0d689ddc1a7c45feb1f44
z0d482e45096c9586c0032e5a1fd7643629fee614adaa267f3d62c8f60ed6aec5dee2d84cd4019f
zeb5e3c37afb53b2033b59b6711d3287bf30b88e5e01ae08092423dfeb262e8af09c606d9a77871
z3d17c43fa5afb2b23765ffe6bbb07d3e9b0d67545ba70d412bfc5af446dfd2b4009e9529f20120
z4afea94152dfd58fed30052fd8d7a70dec58883b94f754f0885ab2a381934a2f4f328819003ae2
zcffa00880d5b2d689d6193b8f9caf0756a616bb7fdba03bfbe39085842c26dc806340b58ac7381
z1c2220976ef0459a6e579713c0da12596c106cd153b23d28ba8053459da16ff2e2ce60a05fe583
z7378124542f551dfa3d6b938df18ae12c119797a1fd1c71bab29363286443c7fa5f9b715014e30
z6fd6d646ced8ac118a3d35f3c6de7b3962fb779a65bfc6c0b066d6d35f7d1b890f1104302edc77
zbf6c19ff8db1fc56a1b9263609014efc6e2c90e5f98debf32da03c86bacba4e380767634a980a4
za84d7f6f9243ee5442d1679232f8db404acb18ec13e61128178c50ce5c92a2000ec36cebf72c90
zd4ad8df4e095e14d0587da2e88148009e3197b378f1d0225e2fa23a14454d9df8d3d6a729aa00d
zf90319c53e5ac05dd3e2ab034c3c9855a94ec8c9c755a6b73bf9b1ab052a7bd8675e561f9d6482
z67047cb3e4ee511b8fa9a2e4aa6805ac0d827de0a92c0a9de097e07a33bc97f9451aff066a3286
z1a3366ae068b6bb4c736ab8530cc3f3ea5a1de296cc47dcc4e013f6906c681cdd35fa55250cd8b
z50a53be78aa5080b907de44c9ed3ae97b401a51c3c363516fd4c5ad1d4dab5c3336b2a8f8e415e
z94580ccfef31de68e615f19ceb76f607f527920d5a7f80cfe3184a50a0f4bca387e00a60bc0e5f
z91cabe6799c9bf9e6dd13fbd8ec2f675b22c59b5c62e4de7602d038e175695ba817add71689574
z12277d23a2b3a36aedf9dbe44c47fc9a7d24f454fadc6da8354032b5260157c63f3690dff0ab9d
z8b48466e8c1e85a07d83a58ea63f19397ca212ee11ff1092333db01c5670531d641b52dab1042f
z55b77fe7327c15501b941676e0cad863d178e46d4d293d897a7b378dfa3a0da153a9d7350dfb57
za8587f2a70cdf63fb566a29c664c1c9a2714cca3bf411f8eb551d8741559790c1e08e1265a59ae
z7562271658374e9100aea897b969b7db4f74181c0ce3618273f0dd5fd1c4d4eb114a0d5e5ae5f9
zdfdb2eb9182c1c452c24b0c33f3456558bfab06742b3c2e40831459cdad57bdb7b50437b83496d
zc09660ff087e945dbc64ed9b88af29488b602813ac8aea24339e700809704a9702e08e35063427
z98dba1eabf06624a5e6041c3dd6c446caca8abbce369ca987a7984c9b9c19246da5e6050c2d266
zc2d4827698f4f6fb3f8cc59dcfaf2b031e3383b9e80d0f3d073edd877ee0afa3dd98a77b15fd09
z93e9c85f0c66ab674a78962befa7bbfe858fc28dd76d751a83f0d60cf30d7203a28f648bbdc801
z01fc0e4d929bfa458a0fed1b02f6fb904ca4a183d978a80346680f968a09d6a064a7d6cbea312a
zce2659ad436309d6ec9b651c1aade070e60572ec0f3b9d43fdfc2b5ad873aa84a3e28e37ab01db
zdbdace0df3f413738309464a60622a05b8ea119b5b6e5ad461ea5e6bdfc26c3c135235f9ed81fd
z7794997caaf09e1f959ec46bd895be781dec90ab18ee7374f97e7a99c6814578af96eaa19218e7
z1f1609b8bd13ddf0e741746aad6f2b3812778ae931a84a676b24cc11f0f2a1f62e693852c664a3
zf22b5f2c327d04eb4788b02126efe3071b6935bd647f6ed7e9b7ed74fd47bf0390fc4ce1db6b39
z7609522d3b046cefa41e744120f223236b22e743f9ba2ac3a6b90f83ab2539395987b64039a3c1
z2c5fb7e3a3adddef2e3c53e8f45db15968c5b554a20108f5bb535ccc2a653cd54a75f3a8dd838f
ze76af7e71010b1250a079ad952662ddf6aa013dd974af9bdd8d8f06a146db254604ddd2768c1dd
z89a0b90e9c05117b060e89352401a9f3c53aac663772b76555a0114d357047d4b6f376187bbc01
zab5487ed1bf1e815e9de1f147726bf03815f4dd6db8d059c7580584d8ed874c4fd2bf747a38688
zf654036964f9b7b8df32c3861a96b97169305aef653a602c2c7dc3df181716b4287f1414eeb03b
z86062ff2232f04f68a039990d3d1eab1dbd1708b7a038d1d468894ffebe66af6645969e6b58767
zfb85571908969493816487629d3118a4521213cc191c285ecc0fe7c54eb793af2b0ac4cecb902e
zd6cc9833d746536070ad926ccd625d73512c3a6b973a5a8bac106d0a62153dfb0202c87f057826
zc944df6c88f53f0d7d27c800e9ebf115ac9222f4d0931049827252a0dd66fdf21255afbe03682d
z9ff9f82353e96eb81f46095775d43e16b28d8e5ab475c7066f90d1524c763e3607b0fd91df2159
za6dce508c510b805613d43b665b305815ffc1071b3643a3e6e7e7475d13d03682f4d0a81f29d30
z202b18ee6ca09586b47b971f47d1bb957ae949042460b12c2d5e8179d4fe6bafc5b2ade54f4164
z17eb465df0774e53745f1f0bbb0eaede1ecd7cd8da3dbaa958cd2e838b9dffa5add2fe8d7321ea
z93062f0fcaf2556b987360738a8388a086ddb5d1dcb81cf834ad67205c6875a82d20a9a58d3d2e
zedabc5e91e4246be1b7ce75ff00f039900c883abf4481b7d6fabd9c97bcc7927cd3f897e0f0e5b
z9e03970096422ecc0b42bf7cc6b1de0015c3c1da0d956cbde371bd2153d92223d72d32392f5c42
z9ae655012f6dcb2f0e8cf50c42306daf3af76234b8b7081c54a7cfa4c024d46cffb29b05317960
z07bc5a04025c8bb5b6a1ba16db77fc3f26296c9d9b2f55bf38a0f2840592cb401218b003392c02
zc3076e39e44f41940bea3bc3436a5f347483e0e5b639ecb52cbe6cb5d3d8524991016f43127127
z2e8791f2adb0b03592c132aa10463be25f1f1b0d7b5c5ebe69bde6c0fa1b4886e75cf1a81c5154
zaa93b7f36839240f653110b8b1228cc9043d23bc9371f9c375366522e8f2803e9f8252c037a848
zadbd17c85167e5059d6feaa7e1a1e7588d8f015881b22c587dc9a75f92efded6a1913b2ae72335
z3525834378885569af24d323a7fc27c88b0dea6c0665d27db5710dee1e0246ba094c4ec72364bb
z01bc1e3ba0e7750df9f9c629e8ae6257ba57689bf552ca4cde76dbec462b06aa58d58a190b91f9
z6d9ed9b1d53750c61b79d95c1ccc11b6da6b838b3aea6251ddcd30a072c01dce126dd09eb30461
zac6a7b30e09d247deb3917e92a1d00df3c21ca1177958ad4ca41d43309df40a92423b0875b0384
zb9d0c9b189aa0ceeebdac85bf358f9c3a35051b25fde4b5871976f2a643a030cb1c73910fd4dfc
zbea89377db4c859aeb43e6461466814e4d76c61a932bd4e57d04eaba4f4b2aa722b0ac9a2c60fc
z88d0965334b48e417249e8251986821f76fba89b06087788461cd649a8c50d3aa59123659a66cb
z412f039000a1abb1e960855b1e9a0f15f0529563feeb5bf06d4e66a25d4c5d9ef0d392be270afa
z3661ac70d51f05d979cf1165a89e3838baa79f7c8f6dcd513bfe2ff6c926b409c581475f472520
zff178d61e9140e87f7514c61e9dd6a9a37fd827f644f3daff111d7680d9d7897ed0b3aea20bb1d
zf65ccac7c50503d2cd71bbc02274fca2a58e491849774507209fe93815a0722d56da25fa45be3b
z42255524f95e369430674d36864d118a9f7729cbaaf31008524cb7fd1e30dee2cdde8cd2458687
z5e5fda8593a98a63dbd1ce06e959bc3989b37b112c83fb0608b0ea8b263d570a8c6ab895e544e7
z129bb147e7775edc6d3d87c70a5775669b98c89eb85d4d1262ce8ededb8154c244bfc012ed46cc
z8ca8537cd1a33cd87b7c781622a349f1f7e9157849ceb82a6c36196b6f917005dd00358d7e86b5
z0651d23fa34a6524cabfca5674e18f61baf3bf9f8f89b8d6084fe084bca7e82b760a02b8601843
z68d265d91a7b23fb1346a30204ad1f141c908eb88d38ecacf4ad668fe11866958e94796e11b5ca
z3cbfae3620df9136a275df471a00d6632d00d463eaa0987c1745a8cc07001dd71de2e7ad55432f
z73ff362621a5993fe8d4b53dae654184d05ffdc827d18fe72c45de3dbfa755b2dcd5508c0710b0
zbb3171211dc12a6c2fa02b9e28b26b66eb55dea144d3f3c6fac3577cfa76682f21570ac6d60860
z051ba208997cec2110649f71f120d23ae749e3504d85c43a3b6abf1a1ef01d022410e23ca36c4e
z8462349669b1a1984977081964de3fab71fe1cfb4148246f66b5915a15629d1253e8e3361f16e8
z8151355a2f9fd0605ee369d7ab722cea6d200ca35ddf86fdad6cf24e85180345ddda3219e0f60c
zbb8f45ff889483ae9a2b2034bed0d482bc01a9bd72c8a6c3b8e2b551b212df077b09958d1bfdb0
zb031d80ebeeace8e72a413e267f3706260286512024f8d9d979a7ab8314386e74703e53c1f6d51
za80d23e6c2eaa68fbdf82ca5ac6c74552e299464487ee2460f09f0eab224b962ab9fd749302570
z51dcf0d8848fbf61a177c10494bddabadc68818e26a51aed196a1b47fdfe6df875c6e4e73153c7
z2b62584afb4b45e83835e1aad39fa20965903eeba53ed485e2e10da3106680e9779ae16bca6209
zf91d03bc678d4bb5a70e95f197adde7c18baaa545334bf53d17267b3752f04ace3a2cd1e6d6dde
ze14ef75b18e2dd61e3727b9f875eabc82e495b4564f0d1661ead62be05f752e16bcecfd5249129
zc9f84de9806e8752ef658c7fade27ca14b9b2c330731d9f88975b9bd9dc27ffc49d5b060c8f2bb
z70a08cae972943dbce06bf95c42a911e92238824c46c5713cc7d451b3319c9c24b79377c1378e8
z30e07c00f193c97dd8bbb8a28dfd72a56840eda8295fe8c09826591ba35f1493a4a287d6f42b7b
z572645356a35cca05d485f4277888f8c48353ea258093a209a7d5a9ba50abcfa81658f6f13de9d
z72d9ab608f7f2523003873985815e878068df131b52997acd489152cba54e9aa988726c1618b33
zc6b7fa79f7d772560fcae380be3e7feb27d265b66528459026a4c54b797c119ee70406c3632293
z1b7c60698d99c6dfe7299db4d4c9b5a104ff1dc0d56c5d590660dac4d6fb2a4780f54a48861aa9
z8b9d739835c1c3f837bdee53a0247bfb88259c998ccbd1b4147bf778679a27341ebb64b40c2e93
z4cb5f5a8b6b09726a71126cf6f9942a59361df18b083a7ca469282f4f2478f1251693467b6f6e9
z32df85d460cc2dfb8c1df5144c9487e6b833e832eee774bb39efcefc3604028c6f966b9534a59e
z5dd7f8133f77bd44203ca40c699d4d4f3d7115ecdf7224b512941ea525220a11eb9a553e0ec693
zffeb9632ce8807ce3caaacade14ad1529da9c14806cfd4f2f7c5f6c0aa3871404494d4536ff4dc
z545484077f54d05d9f0c18d3af52355ab28e8b4febf4e83b7bc033c19e5b399a3257e9305969ac
z727ad63b52090c44f3ed9955fe8d9dcaa90571b7245d036ba477af926ea1b2ac3683a86d0c726b
ze0b5453778b38fa8aff0a01a7d4d7daac00b4a5fb4706b4ddca9322c5b4658b43ada9896493438
z25d626ea72f59f68706efa6cc8a9740e3381bdbc762f16c29262fdcb246d8b11f9e82d6ca9fb40
z4db3d5ca4489369f4311b71183a414116c4fd2be3c41bb9f3341b9b4ca36cd3a5e38a94df8cad6
z7cc8b9798bd1ca989b8d2013b816eaf88e3494e8c0b8aaff96fd3319b891bf10b155edaec08465
za515e3d75548bdbc48b857374d90b78d200146273e7a1f312a1b67c44d66bb7532501e9f40520b
zf6d8cf95d055f3b66875019f926de8119ec549b1f8133fc9eca1dd8953ec306a8a5e1ebdff4c2a
zba9b57cd09d77e53dc1809c1acaeefe830e8cc27c31c6dcc2f770ab1fac5d96913548996ccfd80
z3a22eb9a9d4519ba6f026911700c1332544552b27de20a276fc127110ef1c9a6ba870d94f45602
zf6d1222d3f4e81122235d2a155a969f95526c4557d0d528f5c133f083c814db5dfaccd036086bb
z3f7e0c41cfd078e0b53cabac26e89d7cdd51f08b90c983f50fa242bc9b2bee6712b70d81d8234a
z5dc5920738666f5fe83369279e93fb0e2577ffbd6abc6e769fae4cd6922e827a525274f14c58a2
z68c072e92f591e872f5b3da7beb848f5fb168e15131ad00241f54742ecef1215ee5bd3b156ac80
z22b8df8e81bc2cefc06a0083bb2124c0bd7eafcc156037bd55fe1d326fbc60d6b6d0566e72ba9e
z8834474123806c44e361476ae89ccbce59bb8d288f715a45b4cb8c6a50be5a0f2f4bfe275ccc40
zdb9aff6c98bf9e0f27f151f03561cf7e03447fbde120d394dd791eb6926074e2a1fcccfee0d0f5
za377e8d8cf27c76efb49de2c7ea42126af6831bd047d5d505b2571ef828e44ea318ce8030b03e4
z2e9d3613b799287eedd8d2bad31b9428d313847129e8135d7c7a1b5044f7ae63f001c1ec16915c
zd927854e95eeb538a0eb9ce7d8e611bb0e208a202e4c1da81c116953e7b7f2b08ef67f9ed24641
zdefda62390b8b69ea0e9843cf80f2242c72d21ad82769f81d2102a54fb04b5b2eca928f548cbd7
z52e92a20eea2f2f4d918ffda7b264d38b64d9de37d5230dd6db5c7c8b5ce426bf604606632bf11
z3745f87ae5ce9924cd5bdbc33f6e974e2baed20b6efc6871b4ed0402dafc99bdd9f279a838c8a6
z2168b91cdd4da10fc7f1dd0fd4f1e7a18002bfc3bc2d3ce1848903160c0b1acf4497c5f6312bd3
ze382356ad6e3c84c92700d318f0e83f5ebf101d63004f71f298c80f90622cc35af76842f93148f
zde749c52d3721fc26b64dc0f7e2016324d40680850a96fc7745e068537e1e73b44e48231295756
z9c295bd6c188b0eff1bb0941992d0bc3c44aa948c05e78a8eb68943cb1d749cb982e2aae11a8d9
z0571acf59ec497cd7f4cef217394bafb3ed711789156ca50ac55585c76313803cc8fd52c3ed6ea
z8b2ba1876696c204fe1dfe00038c58a06cbbf3303b6b030cf157cb9907cfc77d5caf487b1fa233
z177fa0c7f0c4200e7cf013d0af256715f3b567e1d3beb64f922fdba6b6ce896e0e302c9f7679f2
ze6e856ad6d12ad42197c3bbe5d240f7ecb405290e1c07957be060e814d9b342e61a72125094d54
zf95ebc513702e4bfc889dfdc364dae53ecc1d2b785246f8dec07bbbe9c8cb997a41ed5a095ce88
zfc5261863811b79685b18252a59adad881134c8bcf5e1732f7f07b73df1f22a3c035093793de2c
z8497b872ac71bf3f977db4cb9fe67a03a7f21f5efa5f9e394bec0d19ac2adabb09a53cbe99d713
z9ce3d87da11f7216e8ff57037078b6161723277cae1d76f9f2c06ee44adc4ce2f7dc554f3c849e
zcbcb7bca48e9a21e2be3c02bc5cf9c21e8ba0e0f4f3cc19bb9c4a0478c6ce53a3be06aeac949ba
zbd529dc247f033ddd4efab3d0304dc40a24d3505faff151633074e917dd019d9bdeb97641b8682
zc515c10fdbd40245925a87129c5f2b451913677a694ed8a3e653dfad89a533dd6b685c5e1dea06
z02b716c330f03c97f1e020c3452d2071e8caaa4f6a94a202ec35c946d0e9a4b49b5bbabd9f30ab
z58204ead111fc069ab9a0b111d342cda9df8091b7becbc96626da0cc608c60a0acaefbf78197d7
z82bf3b3a93e742e045fc59403b922dd0d3c380102b356d3240f8ec9a1f807aefcd47a72bb60d9b
z6a60d5fa33025ddd73934a8c184d24c36058f2c236672bf681e34ff6e5d7c344ee7b3cae4176d5
z30e9c4e63701f49a08fdd37d7d91fd0ad17c8be835c0783b601fd083139635bd8c5cd2b6323e59
z23a85453e20def9efe3bd61f4551fa66c39403b0113e8ed546db67ff12a5ff28e55de8fdaf80d4
zfbd8b416d8d7ad6c8025c90b15e5940f0940cce736bf3b18a52e326845a06ed62385a26f7437e2
zcad887867aa5e75a3929f64989072bfe338095a97debfae54d5d2c540074fa8a7f5ec585b09058
zfcb584f5d71748aefb658cd3f5e0e1630b47998acc09ef337c53a261f74fcaa39409241d80ee9e
z83efeb135bfe22470a18d413f3dee4ec095d268300d1be0457acd9176e121d193d4619bab9ead2
z7d87a7fcbb36728d18dd172bb2c93f58df79551daa656670cdb911809cb4d4e000f954547f7491
z88d09cf4e053af463fe12524985f0cb5816582907b1dc482a4fed068dc4a6b64dacec9e02fe218
zce995b1bbf127e041a7f76b9870da4e3be23cd54bf9716ccd76a167c11c5aff8d9ccdb3f91f86c
zf5ef0498f8467263f7571b01f5a1cb3b97602cdc2fc28c178621a73db805b93920f374cabfa6cf
zaba78b96cdf9e4dabf3fe536ba6b0b2885d7e5a0728a76d6d0a12c57a5e59648b7ef95bb6cce97
z128656c5eb16fe84174a99fcc4a8cde6c9240e3c67e76fab1a3204ae86c94780ab3ed32b348138
z6ceab124b893d48fb77d2e3c0d4b43163e39df67968814815420aaf4d8b6b389e5ac7c52d1c368
z39576612b7659a3f4749626b0a233e955fc231f389e9f897017aa912ae81a49cb06d8375ea5e93
z7fe3f8be9460cef396e232e0a568039c8a5a67ee5055d7b2c55e08d0fc791f67c87b2f92ebe818
za09892698097fb1ed549f749b043ccb199934b0bdad088cebf69631d84ad3c73f62bfd17b1e543
ze6e93dbc298dc3f33632f7d31fd7539e299c69be9691080ad8c8e6c330d3d8ed4a817dcce82b02
zdb42af23cc8cc3dc3568f42d03c62128853dd95782e839d5722e01ba077e21b3d7c3b43bfe8868
z825681d1be48ffef9b1f88d60196b5e8a931a1379ac30fab74fc947c4a05f36e6fced58b947d64
z40a30562cea491e1e3374e92a0ebd500ccfb8e85df58bc5188b39cb081b154321e7ea9962d9a26
z088ccf467f8b064a34fda6cbceb30814dfa5908125a5ae6f7fc3a030693bed67a01cb6b3251ee8
z481d5fe447cb80019cc3ef27a6985f026e75034433947ec166b81ee1a2a7c6f8cb3954a131043a
z34559f6a115a7a82e3fc160c03bbb36b6d2e74d399c94235bb5a918637e265214f99d9de746032
z2216980351aab9ba75ed74c55bd3a25bef18eef7863bd0b0527219f0857d951ec7a4fc82ee2d1e
zd4c387e0a5ed33fd580507c47b64204be870a0139b1d45aeaa6c52fd714eba689b94be5bd29911
zaa0212dcc49f7a581f615b3b7143317df11755e0faa3755d2e27e73b5d846842656edbade50f4c
z0f8aedb71a38784f0b33dca21f93f84a0a275d693cb56575f2fe15fe68a38ee8d93401253d9aff
zb75ee693328a9265d50e2bff47814dbf79bc9a38f20b413ca02d0b989078f00e8606064762b12f
zbeff60d1a7413da31807e87c935a123d06fc421c68c8dc9e647b5b797b5bb8f2cf5b294837cfc4
z265feba100d3f25577877b9ce1f7ab64fea8074a7434c187902c502e55d7b5b7c066fc83ea2625
ze489446ccd135f16bcd7cc3919d90ae2fab9601cbfaff25295d264839d1a83f0abe7abbe096628
z3750e00cf6c2a51e0e6474a465642b6bd20dc5f35e33ebb95031fadb235df447b8069a4025b222
zbe8ae2f6dedeae3d3a734ae39696b480f63007d58201d4dabf567473444bb240e23ea5ed506dcc
z22fb1a2840e97d88074b396f0ede43227ea5f8bee3103a76d056307d9d050fd5758d74ddfbff0c
z087fc8c2f9a0af8beaa2bb6a6756f33168ebccf5e855d7c306ba2708fc841005da3b50909e55eb
ze1b585b6dd979f4a5bb42ce5014fc171b7d46202856f39699bc675f774ce09314841c058fc16be
z3599b653c4d550ab2686405a12ec518a55cca19648913dc37508ee7fd342985795544acba40c4c
zb685d144be32f360e9fff25a91a79e09296297ff78c84f5275b1a9264d7618ea3adbdb42aaba08
z0c0dd414a8984e4904792b70dc1c9bcfb8e02160964ffd673e1f6efddf3b437da5c20817e7f473
zecab17f66892dfd061675f5831ec72cde029567d754bad1eb0e512e8ffcc463c3069a91cc7c6c1
z5d0ecec50e2fcfcf5036cd892a62bd57bb16c8aa6777325ff210c30604efa7e60e67b37abefa2d
z2af667e0748602034663cc7ac33f83fe176040414f362bd7c5ced597c8abededab2204d68af0e5
za64b7bd288c9483876583e3c80ccc89123bdd850d29b44dbf25c2830fa74ef455cc5f371a0a6f5
zcabc56ac0609776820ba9a953297e8ec9fed4553a2cd82a7659e20e9251c71a63323cd8f02a766
z7256185951831428e04d430399f1f6038e15291ac5c87e9d16cda10ca24acc4fa8e32185eb7536
z200d0676ccdcc0dc39b94b3e20f5f52bfcc1b16068023b45552c6e68b9ea84494d7fd078e0f5e4
z14e2ab2c04ac7adf5191d92ec7022049fdf00621e2753b61f36d6e9f98011c1a39fa3b48b5dbc3
ze33652276b911093159c6c77ec9fb30f9418fa31f5ffa5af812a250a9a0b0ac19dd40422df1f5c
zd23c6356dcbbca8cb97636c1fc213213978375e81e232126a8ec05269d104f9d851b2cb3ef9706
zb593bf03306790e72c475a0385b45d3e8ec31fe1ecabd5450f0f92191c1e1fc50543c1d42cc51a
z4b88fafb1c6641f3c4476bdf44eca0da4ce658dca8bc5f6cbf756ba40f60810a59baab3446a383
z083f7ac55e4bdb45e4cdb230305e6679fde8a5a2e41e93c5251678edca562500ae56db449c9ace
z54fa0d07abd3a872f234dd41c5477a0b0ee894bbfc0493a463962f402fa232a1f38e48fee4cd47
z3d9a7bacdd12a9834a614d22aec095d0e5f51dd622d7e0ba09126cb0628f466a977d822aa648ff
z801353f5d6aef2e12b9b485cef8affc6514c7effb2407b5eb95587cd4eb12d9ce7f6b45444979d
z6c18febd422997cbd40f37c98a6075fed20ffb53665c51ba67cccb1440601cef28f2cb9d471d53
z0d89f91e9f3cbd69745362f184716e95b7fc340cd027d394d911a6f2cedf2b0270b7c5a83c5d90
za341e3759d87aba9d18721e99cd3c5eaf4c280cc729dcaeb1a9af9cb99e69bb4691e5b1b4066cf
za1806a5a19ec86900291349af1fecd186c4a32578eb04848bad139216135d90b9dfc6c0c73cd7f
z46b452061a46504ac602312b04f8dda5bf933763ff30b2089735641eae00173b23ff3aa4cb9266
zc8b6adaa05f2af243789aa5e0aa39e962ce9926a5b0bc189f699ee375b33e2f2b4d849ecb17bc3
ze6dc885d481961d6f4c4477a8b5435a6ac74559b2a11731a40301548e0f36b9ea96a2e2c9a45fc
zbdc8629ae38b78ba2fd0fc7744afeb02c1739b345258b14b201158ec1b4fc22bc6defafd8264e0
z72184f141b13a0d682e2203f3df7cd8de2f5205346c4b92f327282f44e1ab46de5df08b503f27f
z79dd12cef968c3d68b565e9ade71b9742b65e397c15f7f642b24f4a451cbc1c129e9a922768307
zec7bbdf63adbef31d95123635fc6ef998a93d1b6d00af6000f6e63c8d0a86a80d936ea94fe88aa
z3d91d5f7a1e3635792ac210501a1408cfb1e1ee6de1aac273847edbc1d96d8dfed2fd62d1608b7
z584f757176d240a160d26dee13353c46472417b78997a09f7655bd9cf04101bd9cb7247a11ef53
ze47f03f3345cac2c4bb3429fda00ab3f3fd28cdd2c2d441514b12e302136995a2195ae129d714a
zbaa53010b837ce7bf4bdc3cc0b280c6ef633218cf6c8df30ed999b642c1116b4d3acae742819f7
zded1737daebfc1465b443c81be723ac380d087afb4fd9634e3d927edbdeb04ec71ff7ff40d6815
z546114ebf69b634c8a88997ced651f55e2e1e83d2b33b36408c256d6880ab6227694db2fd5e4ae
ze7667811ef9c32dba47fd74083093f72e0bfee0ef261fa19e3e3ba823e1c6cf0665de074c7fb17
za7fff654134f2729982658f2c11eeae253db40e3efd1b37a108a1ce85cea26a0ff0676b176a7a5
zb97d4f32f36281fcebd49be71cc8b90e2dec1b15084693070d769a5a5747a019e3c9bc790a2cb7
za1f6a01d9a5e2f701e4c74ee8ae4e328f95ee8fa373cc1a0e9ad5ffc2d01cbf9b56784dc3664c4
zcfcbe30eccc52117d1aab9464653965ef96851a6d015b5b7d05d70cf80fd89007eefc93bc923f8
z04cf8cd597d79e841804dda9697be8073328fec1c9773eda34d1d59db8c4f178a8c942fc8cf87e
z23de4e9b6f9e332dca18a05838d15a9985d5f4405e5cbd0ce1d29d311d821030cd20259f1e1cb6
z4e16af6b1bf35ed7c46676bec0be10c5dd2c3ec9967d859784aa816acfd4ca5f33134df4e63bb4
z62c228a15e8cda8303c13d5576dabc9d13a99243b11a334579a0cd58623e70256097f42f0f9cf6
z2f41b3b10bc8e5ba60e6156b495648a98324adc86b97d94d7bd16938a985f77e1339d2b998b01d
z0c353af6918722f7f292c2246c48ae946e8ab9f0c5950066d7548c4c82b65037dd01df4cccf0a6
z86c58c31b1752babbb0ae2eb46b77820d3292fcb57400be79bf352c39d50995ef527e3b4e4ec1f
z0432b422cef173200ec6cd6b2b389b195e381afea8d4a6459c4c9898a6bbe142131791efc60d6b
z46097ed83f8f7cbf52d46f589d3ffd9f43701fbd85daa5d8547004fe8e0aa37f8949636b6eda2f
z21cda593ef39a65a070208c655e553401d29f2748b0793f82bb96782d0a2fc0dfa5e52339df348
z974c15bdf9e81185a66c9538b40c1f59c4f8883187e9a22aa87a882410976f9989faa634bdc3a0
z63c98a9099bb4e03425013c57b42ef8415c04d3d2977bea050943f27b34f90bb456d6790a31b4d
z56cb7914ecb185e8913fab6c6e9e5628f79a3351d87b6f334e97c3da086e9f30bad015efb4fac9
z82d97a4975aea99ed2ee462f91e3d34bada891e75ae4f4d549fd3812fc4f1fc920b88bb7177113
z1e1ee0655aa45c79f08f4b46b2e8eaa2df781f78a212ef2580c0334aaff4201182aaedd7ea60b2
z278241ed9cba436de1b6d6040ab1e0562d58b5255a16e165986e4fb853fa6bd702bd2b253f92ed
zb5c6b334a2c0e9c425306648f3a370be590f2d1271c8d5796c9820042ee0b0a80586c0c2fb9e3c
z6bbbf5993967a51e916fde984da42ed12a1ae38eaa8680c08dca013f9f24c6fe76ace2dc493c2e
z4846f5ee507fc2b7da1d1ba460cd567ab43aefe40423b57b88e414dad7e92506c78757666b0adb
z45e940e2e978c9f26e2bba37ac2fd37b631d702e71bd8ef8c2b00d343ebedc352cb3a5148c11e0
zb6808d87ce38189d6733e6b53e03c0c77358b40e169dd9de35f7e403ef4ea772954f8d7516cd4f
zd112390bc7432695912f6d3042dce233ec96a107887d6dd61cee223e7fceb171e1d09ab2502a16
z6d7ad202e7b55b136e5cbf5a0c61e4bd50d6ead9851ad5b23004d2fb165114729ecb98786a3828
zdcdb1545d92d1381f654eae16a5f4a9324e1b8e7f21682622e57c771bde62b41102c91d1c611ab
z29cec2164f6cdf6946a33e99ee1614e1da9daa330f8c618ef3a9957df8df031303a91a990f754d
z51d4d0d3b5ad56f9a999854629f3086974f3b8ab8e78e7f35028012a2438cc1e32ddad96d65a90
z25eb7a71c13c4834ce0eb3260601ef075530ff62ca11f8652b9db5d58de319a398a4c43540353f
za3956adf0c3d8c7a4ac433cc79e4aea9b349aa22639eab63a6db69bbb5a01370f4f923644c6c30
z7c3dd43a5da29f7fe82562536a1b590684f5dd5418614d267dc08e086adf86080c7a8ca49279d2
zd5fb0f0f898a6c052dc6640b4ff280eca4be279085936249a0f756805c75cf0d06b2914ac41a04
z4ed884a219f03f73a6f899592b454d621057ad538f91585db8883382a96bb1e65d59b0b33366b5
z3f724b206fe5d2a9405584af9264a287ea4dc9c47efbb2fd93f084b71e08475b9cee0a405969f7
z341794c00a26570b4ce7a905931ce6d6d8d11c45beeabe7576c961c05199c94941354f36a73c98
z872f45fd2cc6236a72f466603c2da19d1aaf94b749393db3f30b90bde25c06fba7a9bd8adb10b5
z9ad1cf25da80ee9426a6d9f7581615a938c619a605c8e41fd0836133365a5cd3b669cef1315566
z92fce178593ee8159de074a42904729ea1ad2215705fc74d8b1b697bc25f08e183cc7497bf69f4
z10964c3aeba0016d910d50797cb85740bffcaf7dfbd3e481528c455438dcb6a451bf6075e3cd7b
z502c253dc8e5ad4ad63017ee1cae93146831d55046a7c552fc5f6d4f24de558afb9f8550770317
zc18641bff66651b6940ec8df4280cfa13540c7b1e08471e6f6c7e2726904660362028b83043238
z23b50cf3922e617c9cda06a64508800f07c4e03056b01e8d29973a2159f6e8f460117ed3da9726
z0be84f670cb32bc9cbf251af79553dd49adae4e5163ce79ce587a37bafd64cc0c5f496881a621a
zcb0fc18df0886d00d473c4f6c901b22499ca9e739ff44f0127bca0b66673b96ea058ee3cbaddcc
z192f4849feecd8fe3e4a0dda7d5166c1bbb6fcef7c0ca23786cc142c582c9c2746c9584c1ed7bb
z58175c11f127744a5dc3c2aa86b29cdd90b48eb1055e216f76fef43c97eedc33a4b47eb9460e08
zb882394d5ea912d951ece1aa261f95896bdb12e14fb9ff1db80221f3872ad86e07b77334f161da
z0d2aaea326d6dfa5bb646512f865fb95092bea5e7f0e511cc90f74176012e21799ee8b714867ed
z911d900cb55474d9270df30d00bdbc08940d095b7e5eb0c5ad8b3017467bed60ba11bdafd73b4a
zd7de48eb9df01d50e6faf94f27c2c7f7772cb3b45b0ad4e603b3e22c2e831729065e7617c56a94
z5b895453f9402f58801510bda9d7e843c202e705300cbf66d44f8610679d1a1f8da3036136ad39
z1a3bd4b50106c68553ea732dc4c35de53bb2bcdb5c9b92be22ee03c59328e2a667b4bfbbdfa12f
zda6d02d6e16d82c1a51470541d4defb7a06e6fa36bfc3c19f6ab1e15ff09bc5ee1b9bbd804b486
z0ab9c78e9a0fc43fe9e8904da0aa802d123e4ccfd9ba318e0dc8ce79f6cf3bb6b75c7c4726e265
z0f690847f73b942ccdd64d5b925e0018586479fd10a45f960fdffe2c107bbc9d20070de766319e
z893177a95d755b8f108186fe0b7ee50b8d4361ec6b588d0e572689f87951a652f773ca3d314dd4
zf5983e066b581976dca17a1ac8c30da1ce1a67a6786990634784b7b0c748ae007270bbe53c8d71
z8cbac712ef904f4e207e8e7b227fd288e1dca1c28460f7d49e94f877507fd2f77dfc9e0709d96d
z7e0c1ec7b5ba0bb67021130c92fa455eaf1f5bed9eb479a31b0ca5d21a22f4227e5d7abb309a1f
zb8152370938905573dfcdfe29faac234ef53f3cf32bab28e26e14e5351f19b2013c97b96349015
zb5d0ee6854347f2c710488caa20e0ec24983c72e29fcfc29cdc6a61143d9b4c5d7fb297abf34a0
z08586573bfec649f42415b2589d9f7499138f4d18a87fb3d1a5b1cb7653cfd9c56e1cee39b5581
z2ca66bfa9e3e04be7b5645ed1a4240a1d2e6a80f8699ab544699bff53d63db7d2f7656bed63e2b
ze0b18c480bdbae1422ff5e98464462ed24e534d6e9a02f9be2019386b13c03fd842501f50dbf58
zadd96992fba847896e203581e74c1443dd0b03c58bda766c5fa1b0bc5ab1d75c290bbc49d0fb70
z641173546e5efad18cf53dc8c399b919174ea63137bf5daf55c6fdef3c2ef0848e8aa8062f5da9
zd68f9e2b3aedbe217f83725e13150c94ecb8c8dd4d182fc7e6c8785b3b7e80fcd84164fbbc3216
z04bb51df26a7a25843c5db61ac49a7d08b42c5c4d81cf0e95b75f18c0bb8782084b9d38c55aa15
z3c2a3bc104f369193d325754bfd4f4a6f7328d331920971379c90c67a6b068ae20fc99525ce93d
z7405db59eb3314656f4607c7960c13c159c558259f8726166d74b5dae2d120736b9fb9ef1f5c8d
z2e8e31a1a8561aeea7b96a6ef8e4d8359c262fa3e8099685a99cfc08a12eec14873aca236249a0
z69c2f7740500cf7ad2dec9fc0432917fee1369a5ff66a2560dbb2b3f3782177d52416ccf93c3cc
z2358429a4304554a95380518341e785509977fd0bbd88c0867cf2cf2397bf77edd46b85d17d211
z396017cf0067503299f00a7e5fe9d7c8252528820f6ce797bcac181f9e6e864572bb0ecd01fac8
z05f5a3b2ab75291e1d50e676db7e20aeb8eb960de30e1359f61502aae63881d8d5339cee800c4c
z58a52827dcf9569f10f59eed7a3a4d5be221c50a9a9d6075678c781671ff6144592e61ce715326
ze618b3b6abf1359097fba996382148455288bd9292340fe23a018e826ff194347a2ca8ab4f73d0
zc8f1c9c58c0cdd477632c71305b4e0bfa25d0879bd685e664aef06960597c5ef821563e2f26ad3
za1bfa1effc7834a51507bbe0b734bb3865960eb909003aacba231561faa6f903b8d35b5239f29e
zae0cccf4ee9e0c0f16087709f5747b269b0e58dbc1fa87933c59aa7d1ef31f44c9cc85edbca27b
zce47a764703c006c924fcc0126228a182765f67cc83da31d6e0124bb2fb9797d1027296d146d77
z25575d617bf618325d04eeff519239afa17e5df9c8d1f7c7f46a573041e21e011ea22ec8165295
z5bb9d3b30501b16e46334462b03adc9f3f4bd7625a9cdecdfbd8fe813b56638f8c748464d65b85
z24b3a702d7141ca140d2acc4e92a68ecf54602b34755cb462efb0138993201fb0bc9b36fdfbe3a
zfd05270e61cbcb4fc9593c7f119997edd15ed98d57953a0886fb99c224a8ad5d71414b35865b3e
z0e6ca478437a891438adaf6a9113a85b582c2acec2351ec34310de7c9078b6023f7003fccecf72
zabe3c560d63ae51449d8b98689524570fb75ff575de04d78fbeb8558284db0da2d87ad6aa2b39d
z95dea85cccceb5686f8f1086a57814cec710ca3bdf1fd153f73274c4c7ef9a28e6964364e37f22
z5459d1bfbb7d76d44d35de35f14d81faae31386c67807361e5a827d705998d094afd47c1f9dc28
z7b839a94aebc6b33a5264d750eaf834d2f24779a78d0fc87977785170625ca69b514e10b3cddf7
zd15bc5f9c930c1991332603387d4126c8f37658766063d211551bd8a5d3929dc45ec458a24a1c7
zd8f556e4ca2a56fe20f4204267d0ab113b2ddb3a15aa102aaa105b70eaa1a6eb584d894f37ca17
z46153daec105581a48c54286bb701b0b72ff5bb9b397b6f62e08d53a18b1add8ab2b759076b303
za4bcb351d76449454a802b895e466fb15fa07b03b97c0d1c62e6352d9e7927b5a11570466473ee
zede799b0f24e4751e93757e77d9d82ac3ba445d0c7d26f725440b99130ae8fc5a172cc8ecd5380
zff74d8ba10a4e9365a612b6a6d6bb05d1a7d929b102076695f1870aed0739e2942a43bb7fa8b10
z038589a70c3138054b2cb8f8691305cc52e65b4be69cfde6c496e165e694d0d65f688992c48f56
zcc4c8b97ae7c4d8bdf59cc4700aafd6dac3bb755984aa0f1ef55f8debf06bde0868ef31bdd1f29
z99ad9f8669077c44feb9e76440c1ab92c679a6793a82bf241a5dd898cbefe951a6107aa2523b72
z9f2ddf51e2c355a84015d5efa079cb7a59221bf49077132ae1d3aa531f75d4f2eea61e48c2c85a
z27eee1152d956c32bf919b71e1684ae3041f59988038fb2ce391f5c8dfd97f8e75b05411938e55
z710417ac249fe8fda933467a9a3e0c9abe7709170227f49a146a51a5ff2a31f50ceaa1df8e7dee
z03518fecd996aa27255bc19de01eed4c995ddc0060bd161bdcd8fd2e083c7d913decf49815a2aa
z1f5a4c4740968e81d6d407c65954a1a607502b7f1db1b2140eb2c6242c6516f75d4ff33f859fe0
zaa704914a4365899c2740279e047ab028ef63faad24351ebd29ab49501c886e7755b8127ee4b03
z3a7013b1b1a31e5f638214035b8b082c3761716630095da73555245ce354017589091a62c6d36f
zb892186e91545f5dbd297e1881bb8b00e01c6eac1d1e175fde1e571389bfae9f616489c3cd6328
za5766627bd805fdb4dd86b86a5f2d7a8e6276532e54415133206fe5a0b79896e72a155f29fd775
z4fb4f647578b6d59c776304543251ead736caf7c852286b2b25e564e7b51d433ba44e3518e6614
z951c09e08459360927562b18be3674c439754ca4a3b297d50863426d7d1a5159fa6d718914d400
z4fddaa0fe78def03a684abaa3803ab0540dc4da1debc80eb0cfddaf2814695a916b35754b1e50b
z51cf475f965c23a2d513d0fd6a5922db7fea8cba98c60f08d1a9c6b0b1265fc26e674e629a4f63
zaa881ab2921e291e6df6130e7c4fb9264d56b4fe37ecf5240cf7fb3597cc3aa761ed47e6addc54
z9dfe9b51406f0e836ea25cac35b88f56be2f4f8a715f4a9dc9e27002ea97e2f1b4d67a6193dba4
z6fda768de7c25356c9599794f6021c5e29bd4ec38af02922340ec48883071d8592437a7e274743
z7e075d9d72e23e7581ae5273c13bc21a43a02c8b1614ddd3bad6bd88aae497cf74f657f5dd20b1
z4f0593efe2b45e0401d7783f63eb39a02d87839c14c2232bf65c2513f77206f9eccb5212e3c1ec
z5f2a04e6d6ed509e129ace61d85c9a772385c8e2b5a0eb9c20e5a60a71d02459dadb9340e159c3
z11d269fced119864f145f63849ea6aa1a20ba6d82f7eafa6965a0038578fdcde31677368631370
z4c1834f99e824de26654c24daff9076e6111144f87567174db12b83f180e5356ed9e2dcf26d48c
z94a66a56d98af00a1e408cb053410ccc834d94cf5f7f74c0ee8764fcc1dd244266c16d0f4ac049
z78a68cf0dec30d4f6eee7905ba1ecfb7d6090059cce6d4fb614b78555fcb46cfcdd546e409da96
zab3124276714c3a4dc3c8e6dc77fdf2aeb7678c31991ee676c7b7578a752925f12238e42593b8c
z49fd2ddadd952e31a6ff1e78d31be1c86111e27d21051532f9bb35dc3bf8a628b42f130412fdd2
z28742995871e19a62b0100ebe2cad8d28e7285410bcb525e6b3c5f7f1baee4b8a936e729b39ba0
zc1593eddb4e3743fecaf2f9174f0fe999b69a4c68deba1430be5ddb0446a693711fbe9ffc1c243
z01e0995d201d015afe22f961b4a2334661a27932574791938651934905d9dbb442e140da14ab88
zcc6bd1e3571ccae2b99dddb8ced41b2c2e8dd74087db0def4101d1b2ad01dc78c8e281b6b5a910
z28d134f4aa92b20fe98d31b3b499fbc169b627279dff03cbac89346da015978a91d242c7a5bd7c
z08a4e90cf3e740e381a8939a3d95418a9bd4b1a5f4ccddbd0d21367b40062fce7eb61457ab96a9
ze83b5498955003ec4f1ee5703399720c2136a4fd11bd069655b246d92666c03ee84be9c05eb792
z7c4f272f8528d6121929cae1cdf505fc711612554195f7395509609b5c760b584d8c26c2c74e75
z5d5f58f4ed8059e89558cb369e059b4d1ca55ceea060d265cba9d6d2cd87a76b85e0952ea1f0e8
zc6c04a5322f3810b250633f1bcf1af044eb4c6df8712039e789a89625a8852e903a4f9248003a7
z2a91f63fc9c002aad15360f863e5476083e626b40b5c84eb75331e2141b2f28971e31c7104de7c
zae403e2840a22a455ee999f7bc5e63a4e67aab1aa1fac52dfb3fadd12b7cd8935ed6ae0cc0e667
zeb3c2bb74920a86db4815d5df00bd08f3feeaf60eb5978358344a45cac7a5ecd7a88d15f005f19
zacce8000f7912cdb6d44613089f134d32fc310aec40950e5cd19432237fc4f1355d8581ba048b6
z752bafee7455a7e19d9e972273dac22f50130fd414896675c4c4fe253d193c94d6ea16c00d47a3
zd4c54ea0e01b7d3b02c5c2fb9d4f58e9d70daf5313a7ca5323f75e6102adf451c5bec7d4593e06
zb6f2dbf6b7ba0314d75119d89abfd767089004323e86d2958b71c86a2a2799c73b599f8ee637b1
z2ee0143ea81b6952a1254bf3df0cca166930dabede3fd6df26bdc75541b3a1532d5c6276552af9
zee6a166b9584f4f918e0973e7e9e70c9769d11ba4101ce247ff9cd92869bf6c032a9c959ea5800
zc960aa1cc1ecc3a08f26a22d54a4f252afa3cb3d17eb67b0f4c336b383b158eda16ca70b75dcdd
zab77cd98740ef67ce3c0261d6a8cddf3feb9c3ba9fb27b0cadc85c6b96dfacb0207909fd97dbf0
z14403e4a4b7a16b6225951f5e29b401d12088f45abf110a3fd4de49b98432c6b68d12ec75ad89e
zad04469e9f28f5dbb476575dd53e29d0c51139955d7a016175f2cd5af05739cd9d6ae1199c3cea
z7a137ec9490e1fab01f568a0b3b07ef9c769b76ed4d7c3c50cc821e9e781942d722e6fa1b9c032
z76ab33acf6b5572e047f9bdaf8e16f591ced9cada09924f6e07db4f0cd41970e853f3f207e9b65
zbcf8c6f96e73939ca7d2629a5b5b80dad33c79899ebf59f832e16033c8b6235cbbcec914c4e81f
zff2258799f556fcaba3d373c9b9f949fcd7969159971ab6c73f0d99e61c0458a1ba6dbef078c1e
zae82ac2b94dcbd9ba4a42282cffb5cb37402ba0a72645b28e265442822042f522a66aed8959e85
zf3c438e42d5f570d686458881b9981454e0ac396a92a742d73ec146642b11d4f2894acee43146a
z7554619a04bca116f0a553a03ffb7e5ab79018718296aefe2e05837d14efbfa911d7db09be8be4
z334f4a89207c8aa5db5c6640b52fee6d640c53418779e7a2decb9903e3cadbaa90bea39d439cda
zf6c571610b162a7d600d75ab4997ecab122e5cb21ad6af6ca25584846f9d648e524a0136dca86d
ze87011af105fdf2564d48642c3f5ad2f4d78ca99da5b094a9c9773991d0da086de9d9b7424cc29
z585952578e37df9ddc552ce941f42c7a087f5ce47b7a204920fe17dc755891941007960a54dd06
z8cd80b08603c4c92d52e87dfddebbfc071f1823bdd18d84b01d346d8e6d5764d91479a10c53892
z5d93f3b74f8ce339c29c52e0fe5a85ac346dc881ed96463c4d8b8d45a20ce6eaab2c6e1c989e12
z6406a3ded988d74ba03aac3190611a9d2475147ac35cf7eea05880756788186797fc31bdd78446
z0ff9474b55935fc56ce2a25fc08ed2a36d522b51a42f707e0d93b399b241791d6122f2b09fde8c
z54a5090d62ab5d23d3e45d849effed325f73afaa332d33fee5c59c0e1bcd582de7575cf6b14583
zc7056c35461462557069e2cd29f082c60f58840057002a4cc308df4c6510752a61f01ae1da46cc
z045fbecb9f318ffd115517b0e41e4f9a32388a9ad0ae8dfe70e71d00aadc5ed48c28e9ccc46274
z319cc24a5cb07c8f1780138b15d68df666398c21946fb0a895dcd0b05db5109af3c8ca96d6af3c
z9b600b024b264b9ee1ed9ff7c5f2aeac7c57347f47ef4a2ae7a57a35dcf1b4ba8e0b977d2c527c
zf9b947391124bce53b56e1dddeb8d13a6788b971696834a27b63be1b5eee26d593f1639052ecbc
z7f086a5e0b4232617dea6b36a1e40388a1ceaeec8008fc2705e3fa93e76886371203fd153ff1e6
ze30057029636ef4bf12b308f74d06919f96e5df530013cba9e220a75561ca65e7fb41a7ad8a581
z4b5d340f12c7524d15a60339ec682212341fe7edd434a02970dbacb6a0321782547faebbe180e4
z4d6f24980e51c1f5ac01f379e775bbfdaa5af696aea7485dd05948ff46fde8f3c06d4e4c513707
z029a9aa059b5f8f36e6903880b595e53f4aa2954d29595acd2a7c69fc0370474d5a62bf392e131
z20678142d5d81e9b4c03d0380fe3ff0134652e86942621ada4ac301fcdc66ad433a333e0fc1550
z0ad258c4209332a100d7dcbcd0271b9d076b3a891a6b46fa55b5b39956b0a15ecb35749e3fc6d7
zea2ec4eac46166b003765ce9c42858fc1808e07e3289e2b9f79394f4ea887fff8e112018511bb0
zc781db175ca24d4722b2f6f58af551c0d7e9ccbc0272e8b3ef557a0e2f3ad293ca308c83edad3b
z36433aa823a84e00f10ee81d7b9466fe2a853e71ba3ad80dc8cbc1bb3f76d9be63e8601bddfb76
z943b697b2046441ec38974e963a6add8704c168c6a80c6f649cbd99410fa1d5997dcb1b948d567
zd3a5d05559a3e2c31f329b7303dcc71550795596598d3e0064fbf7d54a77478b51d7a765964259
zc4d6877521033a677c926899486870173c7a368fc81329c50835b90404be82c0abd9f2a249367f
z3f4b5b72589545419460e9fa5d5a00689dc3296606a405f0173c9f1b19a2332758c7b5a56bb5f5
zed13a2b8b1f336f0cd20dfaa86da3cf61e98e3af61b10239ef5a77e7dcefbc535fa7918bc41d84
zb66571847587bfeeca239a2e9ac4e5656d41c47ae02d1bc77cef98b99738939a76a2bbcb4ee470
ze023959bbe284918679cce2686994f506323c8ad69af9134c6af045463ad81286c1cbe389ec57c
zce639862061cfd210881988665d514dbd5506dc0eb9e629c31794ac641becd690a16e85ac5aeef
z9e145eb71d49326ecbdd0797fa4e97f21ca8c06061535a4cb2bf2ff5bedb61aed5ef3014383e9c
z0451248c17a0e3263149cfca482649da788596cd4f0c3c3f07379350de7d3af54eddc20d229207
z66b6216cb2147ea219e122b458de6b6e730eeccf7aa1ab93c7e8d3e08de86e1382c8537c659023
zb6e5f3666fb4ad7f6db19888e172f4c0ce455433e1834d9be22ca059d7290c694b7b394026dc1a
z431bb47e94146da1b34db024534f813c0c06430309ad4879c31bd11afa97854db431575b18ad17
z753b9bd405b13b2f556acf19d60ec9ec49df0784517bad9aba9fd7753627a75b01f034c931d365
z28f6049d6a06ceb585cfb551bc0e2b9208fa71252757c4a962e491d0c5d15a4e6a39ee2bd92e02
z340d857624f775afefc332ff733c7de61532e85413e97cffa67bc6a2b71363e67ac599037e5c62
zafcbb7258e6fd9ab9ca9f516dd133a44babf2e9634e1c592a10ee1a31f7ab4a91d2233942df761
z83b0355d78630d8cdd5b533c628c11f73eea57756299c0b1d8a89aa7d588928db87b060f25d1c6
z0510b7ee6aa54ac8a2b9900d2b34bc84a26de5ea25688386c66c3ed2b13c5916ca7eb20456365c
z8874ac79977fd9fd35d312021c8c6f31f6bc61e5df45a3a29246a0c91f9e40f92427322d6e53b8
z3bdd64b29f2bf4a4ae7cdea9ef9901fa033f5a822df9f0ddea319b9444f0b5334ea6da79139749
z31785471d34995712a645082c14e64eddf9d2f81bc351f9db55b63ddda3d25cc4b68f9dc8f5449
zdab931ce3df1cf2c146b17dded52542f2c8cc523047107641a5be74bba4d2529a955d645820560
zce07ced7d4ff4f03c1c0db6cc335908f8617f9ede94131250e7af5c30735cd8544d38d6c72a18b
zbbd6886700f019da66f61e0956c31c17ea53c8eb9348a1631d017f126ac5032f0da57a73aab5b5
zef778455e3311e1bf8ccb8b3684a38ef7654bb97dbbdc2e753fe5b6b78eb2017ae39f887c42d3a
zbb29dde3a32d315e2d5574600b73b8eef335091350ce1e12bbc1f1bc2c3fed809bded8ff07398f
zc3db131f9fd79be583df665d283c1b729f739a530df7932ace474b4f08591989f316724ce2d500
z0de9783d70fb51fd653b6928cbe513d313801a4e2322e45bd4e797562accc9d9d79edc46fc94b2
zb0fa6dda47061a79b10fb9516d98a5ef6333c19205e3b1fa44a179efc30f7a399faa14431e78bf
z146b6c02116b3db3436a418e93342b81d06e372a446d2c479b11509746dc3d3b07d1e0df183780
z766ce54e8e4989526bae0a7ee2c5e34b72b0c98899f3802b3445263b224a640c5dd2eb98940586
z3e7b760196bd3299980693f3058c8b137c3198d8f10eafd16877511e7d37927b11c253333fc795
zc604e26ad9dc379b0d404298b3a15a4be7b26279aee1a8f91c5e6c73273977b3c2b9e4dac29f48
zbc93c6efb2a948303af00dd8ecabdfaa6d65c1e955c5c721a31110a1eeb0526a0980ff19f81741
zcdf23ed18f9cfba84f7b9a84a3afeb065775afe36a76df0b6103a2a800d2570f73b8ab9d4d8a2d
z7a69b090eaeb9c559486f3dd9e1362d4e419e8d198986f528fd320f96c880c09b115695cbb3ea0
z0d98fd6f538542086aff4577bbfbfa292938bf35977dd4905fb04d1f0ae79bfcbab336ddb8b795
z92b0a04addc2cfa218af188882ee8f6a88a0e46e466f6026f965b83c0346f229bcc84d3ec59fa4
zfa4703e61bea9ecca390a8bc5714a7c5db9ad520934ba547301cd5ced16e075eb3c14e8751495f
z37e65a5db412a3603a5007b83eb63dece79e57bc08a42a8860ca40a9a4321198a82f97bc03eecc
zf8217bda2ad60f51ed9da0d675a4a7164a7774e1dd19ec10a3302a898cd179f25fa9f329267929
z219800ee8ffe81d1e98703d6de01ab5a6673451556c0a9d9f88060e427559d6508383f72bde8ea
z58c997bd693c6e043cc61d39ed737dc9dc346fc6fa3339f651ff514a0b3a5efc65ad1d9b0d8da6
z8956c70cf8120d7ce7d92409c9523b3826269fc47d2277400a80f4eb32366042a4958dc65a49d6
z9be04b3c89008e3ba9599f153cdbf79fc20ba4d499679a85ee7b7d5c0bf70c40d525b186f9161f
z6ba1bf68e146a1900929cb39b844f107826e33114f8386a9c2668a66e1161fc91bb114ccdebcbc
z5f0ce6e1bf83198a850c3213edb2cce41885341dae252625b0d01a9d804a3baf5165e631377d7d
z77f90d53c24aaaf54b95cde75be2c21702b28867a6d2e80044a9022c6732bc5a5dc0bde807583a
z9ae635bfc5f3a3cb19a4f761d33668c96f8dc99d2a879e0075c089b2268ce4f4b1631070dafcf6
za58d1c2bf83dff282de67ff71a3e767e8a35bbaa71f5869809d825dbdf82436a480e399ad88f00
z11d03093652a9279d08be1bc01334a04d0d774053dcf16df8dc1df214c5ee948c1826a31caa1d6
z9e189773afd4c1cb22fc28a7b6c156cd53bf327ce5b957b5e5f315fcc96ecb31b9ceb9b86ec0ae
z36f205b73b651944fa5e01e30b7085e267618182ad3f407230f0f127e0425ebd59ed3d050c9ddd
z27b9710ea9e9d86a2042334217fced624cfc75492c5357db52e74e4c12f25ff62067cd2faf2371
z16ba5bf6436fd48169bd0397f41f333c8c1ef705f911a3fa712a0ac805c141b489bc953bb7f642
z7237238cab608a0d664dbbcef6b041293f3dc42054970af6af1faad1da4180fc4b6e233da2b40a
zae623d29e8769672da2506e57f1448893569f8e0cb88b4d521861168cdb7de370b8eb30bad4f1f
z0c3e25fddb7e8cd95e4bd502fa544960ea49b790da59f27aa2d59433a8c9fb1ed3cd1f511187e9
z32b8d8ff5edcbbaeb316a7641353b0239207daca80004e2004d168c3fc6ac558aa72efeceb918d
z7d3cec8a4ec3f1f6e3b809c1c016d726344ba817385b2855817a785ae8c45cd91b3d3fa37318d7
zfe539db2724f781fd19709d6739c815c980e6d5c514acf13179172fda0e79ef620e5be1291861f
z5cb552e29f5da9a345085838d157af8ef7e490ffa069bb48041066a03fdcf48bd54f9a1680e943
z89601b47230f495f81b0209e3488c02318bcebe9ef0e4d91c4fb09fc482c62f7c4fea3c74d6054
z32247dc674748d7437b075c5fd92e4458949532d202db339d7fb64520a47522c147a864dc9c93c
z66d06a5db782181655b852ff68c9be7da98eb1b7463e7c406055c67b07513bfc3c6b8c87789922
z724614468aa83d02f27907cae0fdeb2d2fc816dc3eacce80dafdf48c05a8da11097ae8a529fe0f
z6830398a98d997917010508c44818db7decba989966853436325eab9641ba02079605292e61217
z4788f92b522998debbcc3e66db55009393df901861cab0f0d47f47c7f7a5b6a21d05ef747c903f
zdac318c6b6b1ce03665bec9ea9c4f4e6af5ac54c04b6f84c46a5883341343062c6ad9b94808e1c
z2bf0197b86b2eac26ece55ee6fdfd87c2af3131a8d91e4f175f90585675bc01d7601297ebe7357
z1bff1326fd7f13ff3983667371fcfabf3625102299102a370d500b88abbb0430a84c56a99b44e5
z9bc4c47305cf3998c05dd7ca9fcdd96acf78ed0d6b2b94fd26216697a083fcbeb73fe206d30ef6
zad1c22bb94fc18bc9cd4631f72c39e41efd9d08bb6930c3669ac8af7a8a9d2455a940bc38adb4e
z8bcacac53610b400ed6375722f7ef649903f0e8406eb121416227645d75dcc5b86e50349b775ed
z633f0e17ece2fcbf67850cc3b31529c6a97f246eadaa293d34bec53c7906538dfac6301c7e2451
z457dfc3844981001ec74971eb6e7b0d39e56d845918b625a9a3da6ff60a0e9a6c3b02aa2c157c7
zee49033a42300ac339bf2d18d38731584998de1d05e061ba2899bc33f89b4ef62f8c9b83f67945
z1abe79e4fa1af1f631e790d394f7de56cb467327f617b2147a67f0047f7e6f304059fcf501d93f
z821fa8c3f829c661d79a6e29b99c6bd35f6d5315ee51d3ea554695ff00e3c5e24df96f9842ab89
z93a172814b54eae9296d71d9ce8696cbcf2ec6d71d43e587f240f883965f51916499d69bcb34bb
za1737cd1cbbbadc7c4878faf6ea151b47c59f79abb3ac43ff2edc6471da908486984e7d60e2ed6
za55571b6771a975248b50b5fd2b384ff070d8731d8dcb82794141baa52ec3519bd9bfb76eb3d13
z02f9187401bb04ff3d4dccb01250ffb9969850ab3b35a43ac01762cffc9b3efcd2903f635cdcc4
z412c325e558d16086da5411f4cf10495f57cea23f5dcfd09a5f4c7dc5b9547ddf5693637501e83
z8d0d52a379e02c03f1a753d4106a089c4b55a682d53996730d6919c9b179063f5b8833dd5a2a12
zda9d97f2963f3d3fe4a6ad5f94861234d888b80a60cf2c1722511f28e3d5da77a649b44a384442
z0a084ea34b33017d5f8fc92400e9bace527d13ccf9e8d611b9a12ed92b9e2888d1880d2f09161d
zeea7036191bccde0eab79e02e1db90f5167e0dbd627b5d2aa09d64f5ecf7359392f250b14513bb
z162eb6cf64c025568dfc86043e209a35babad1c1a01dfd024207c8ddc711631caa69f00377c6c9
z8f3e6b5991c4e30e04b616dfef2fae0a3f42e0b1d503cba3e2716c74f2b8409119af26768a16c6
zee3ab5342c9dd7a335e2687f6812e7eabe5a57dd853e93a562b95410b07007a830651b063af3a2
zd84495519f3505e669dae6c74870f0e3ab863c71f07d8d6c7512ea102607d98100062a31063e65
z9a4f35dcc7c04a8c9c0ebaa5f4f3655b121826053dc3f114d35c6b4152469d6b2a05c5d981b82c
z9dba3724758515e78706703c515f17ad0e376ba2154fcd0ab42a933a956d5d1e02e34f7c2c129f
zb0a9010a648e4ff799dfd66aebd0a198ecf004bc56bdd85f50d56e91106721a11ecfe5e8fde72d
z0c582276b833b6065449f32f181190cfc0e0f351211c50c8ac60bb19b474c0956e7755b296a70a
z5423006cbe236ffade80a0af065a9a75b0a152b572250f6b15ce2d6b6c7224f27536c67cdcae4c
zcbebb9193349baaebbe474581fa5c49b8b31d8241c14e6ca4697285bd40d8d03b88c7be51e9490
zb574757429a5997fac9ba776e03fb430e3b6093b7cce5cf1a8e19544a6e2e7da65f0dcfdcba292
zfc1628309cd0e603409f9e743f25c8f4db9f2186ffecde04d4899f1dab2213db57d99eae98a398
zab7b6056fd67adf0ef6df0bce8a1deb4534ff2375dd9b1a3f67388050e452d66ad6befc0282478
z37b4a4418e92f76121959a0a0947c923ac27b8c7551aeda7af2c98e717e40df0ffd0181f7cb8c6
z9b9f40f291621e89075dc568458e8d42a09a8b9417554dd7b3c23701a7098c7dd20efb1c630460
z1012e70ec3891128418cfe1ffd502ed25631d5a629122b96ca24f5010e7fec072fb16fe0551969
z6b1317120ebd2e9cf17f073b79cd1984eef0f2681babcd2d19853e82d56a1f1a0323f4351c31a7
zd4c190e2909cb3c11529c4ded042bbf9f54dc75da2fe3dfe1944a2cfa554d97110cf4f22de0360
zde1bb1bdb6014218dbe06f46e8ee8e45e6fdd0bc7c3c9981beaa9f11f9acea8e294b7f8189ece1
zcdc0cb7a82744cd15cd64b40754be4aaeb528b801f076a7f4e2817b55f0dba357ad4ab4d36b056
z76932b01b7f468df04c014304b5bebc4dd47f6fe976b0b57dba2db0070fdae34d1c1285d899b33
zd10c66c625fc3529b70a8711d49306370f4db04be25d1e8d9ff33ce470e50ba266334ce31e8f5d
z0b59d4a56e965063c8c0921535c0cd7dd415e780996e8c2489ccd52bbd168834bdac1f2c4b2a84
z0872220f47b29160fa1829f4ef2444c0b293e78bf51ee441c0b7925cf05d18f868d97ac3cfe52f
z0fbf7ebc93d397a75901435523cdca91225da9ea8181612412bb661c7b69a051f10a4d711480e9
z07210688340b4c090db89352d6105331963fbe4fdc5407b89c051868c3a3af235b9e39db638d15
z187d1645fc23f2bc2a0f356a23a57b2caba94c6c3f54a0cf043dcdb47a8b676aa24c47c87e7398
zadc78d5f204cae1bdfd44450f73e80da477cbc79efb6f32531afa093c45ff91febb82965778702
z132520aa9658e70991dace6534f3864daeb4034616e866f93d5537eeb4da38388075dfec5d0c69
z367d53e673421ed9f0d83746ba272cf7658cbfe92f830ac80098214d60b201587f4527518c7caa
zf1f615374dd46d88e27880633c58a4b5029508f5566c353820efe397344a6471b4bc3a610507fe
zb51698efd1d53adf204a12ccd426b51d8646a8eaf972cb088f3505c4e8847b98eee3d5584da0d8
z3f84da565732aae4f686e9595ad926eaf69b422669004bc995aadc337031f09d858ff4f9bc4893
ze08a8236a56ad30c6d7ca8408bbc3f28326d59e2dec312dbde2b5c6ca32a66cf091631d30f15dc
z32d786cd13b15e4f2b748e3bc4b8dcd156c4b6c422b0899bfb553416a9ac2245fef3eb00118996
zf6857767c0585b7f43bec77373e0cb5bfeb897900d4b3f867e608807475ecef2a5d02744d52751
z8d87f01b39402fd4532d4af0e293e43940a5cb461acd45a1c4fc16db62b91911e3c2b9b815ce67
zbf2d8603c36dc56440c48919f7402ce10949d0fd44bf182e4bf77d0a21ebb474a4f4b26f0b6ec6
za7c6096e37b2e7748f791eb059f7c766fcd17abcddb80521e902c7de3012b39e7b81c0884eae1d
zc0c4ca0f3a938f3a12d8dbffea804b52741d9a4614131d8d8dcbd05accbf2728c23c6433cab6cf
z295376cfc5528b95dcf55c9169aa637d5821c326b498f25ed7d64b4e3f1f055bef5539821ab9c6
ze484b26dbf16960b93762af6bcc229717567fcbbe9145edf416f59d8112c86d4c9087b4a4eb4ee
z9d30c78b1e4379495aa029cd4ff17730e1f660413b4d9c791717a41fa19c3b3f7ff4dcdf31f81b
zcf6df8922ea6327991edac852434461d854399b7d5d60b44ef77b330ed7291e4dba5bac6a18cec
z1659ab4a840bc9dae0924caca99861965ee96e518f2cc0e645a33b5490cdbf8fda35052cd0bc58
z944bc47fb33934c8662fdc7ae11054864adbdeb7e471f4f53667d815b1c8ff231828c9aa7863eb
zc14e29029e6165260f1678aa12e8731aae96c7cc235d34bd63df25de7afc4809d14eda5ff0dd03
zfc0f8eaa4db169ba7e56cfe0b4d37e55b084ddf5428b727b1fa3ab59ed9866aa40c68dcb00f1f3
z6fe55aaf3e4308942ad06f1b759371715e054cee15d5850d36c54e50b4991a027247cdd705dff1
z860c3c04a922204b4aa6bbece8bbc8348ef2716ee017298def483a2d80d6f860ee67405a8ac7b6
z9bd037c92025c27644c031774f95c4c6ea1c9e6ce5a297e4f6e3c4f536cf08d89fc05e9082beb5
z5cc558ea1625106ee65119cfb9b6e77c78b8adb7cf6e80d98d498a05d6dae6082f4ead2a4b310e
z3ffce40245b034b4a8f6c500ed46e2d560beaabfb39396d7fe51bead5324c0af6521316145a893
z817fa05048ec910a8ddb3391b5642c251b82e9e960969e07fe0dc62800a06dc0d0fd033ce96116
zbdf42a2d0e0169c63ff24776a90e4e97ea5381ff83d4e7dc7ce658e0be9aebde4de8c92a40cce2
z5c10ddd651b2b2445cdb225145d0728e5662ac723df22b36b27ab223ed7f148730c60b7af7087c
z948b2c7b7a3bc5c14f579d49db4791b74ede169049afdf9b4f76a1831f0025cf93eaafe59e9548
z2ba12a278ee15dae7963faf89f35ad98cefcc8a5287f774427b954a6a3fc0a54328d0857e5a00c
z0a723aee4ee95420282c365b3dbe59ab38ba35809309c50cb4099909752f557683d95b7be837e1
za2e8c7b1777771f21ba93e640137ec48d6c49b5daba1201fb2b3c1e70393afde9e6a676a6fd9af
z82539f1ca47486943d8e9b38f6d24f8e28b1b52dade7dd49587aaa0f51cf8d7e77efcce7550555
za4e6202317f8f2a8eafcfa7e5af282377fa4dc15c1ec06869ced91ba0370e698f025015c323aa4
ze3f15a77bf446470371f427271b145bf3ee4e226d1830a92e353cb1f1c5bb57a46140b4f2a3993
z00a5dbba6dd5ea0f230f9ea4b917cc6abd93758f08b293bc29a9951afcd7138248fba6a3366bd5
zeb74cc4e95d3035001d70c10bf023fa4bea149f0bef9cc4f087a1ffe49838a7241eb7cf737c9b2
z43134db259383de344abfc901c6f2a7db7abb75f69bd78ccc1b707a85239e4c75a44aee790b9a4
ze64510aeaf828b2175bf2f9ca7fa4a4049c2857a07ae29429c2f1bbd4d31e0b7fea9d56c1160b2
z18a88f154c31f3b6077671890401750f9bd6fa0e89fb8afd77b48200dd67ecf0a9fcf9f4fcc539
z15837f35b0bb4d98d969d52f2390b1134f0a8b92ed3d734630278b0f0f81d0e6055bbd8ce40df3
za80548bf4f19decab86e1003a8800b6c6db743f11a8782df9e57719365183154a70b3548c9774e
z2f5af8aa4bdeb7eb0d3fc5cf8990e9d851638a3f385a43e76cf32597421b2e095a37f157ba4422
z403fabd6307a80dce1c6af5f97345c989300430e929b9224cf9820154d494ad5e0eabef55cb0a2
z8ec823f4c496fbbd5e27a6d4f54854cc9d61ae6d54f07e9844d3ed2f89c1f186120b5020b906a0
z213cabdba5924b94a86a96f5feadf6afbb2ad1f9a9d92c7dcb3ff7f6deb487a4162c4bb6ad11a2
z41c8a817753fc5ba7da2153d38a344c32bea59adb158e5567871b203ead945ff90b545daaa8c4d
za263e984751542b4614b2c314e7a42e06e7e7ba8945a3f7a390af64dc748b1f074b643874c00c0
zd2199925775f6ee78b10759c2fbd6f1690ce1604b251aa629849c33e5b369520d6e9932bdaec26
z7df3fbbf14a4b7c987aed19a766d6c4c34cc3a417a6dfebc73071f8ffe595b8a59dbf67d1caf40
z7ddc3c4bc63872f54c0869d85b30a139b8e4796166b661f91ee0419ffb7a8cb509db4997a8ead8
z856bde6e916c0bb67987aa4859daacf375bb36ed5c67db0966639d6adadf8d97c165b9a2a6ddaf
z1bae67936411e80fd057d4ab87249a8035e5a488690143cd27b178db1a32c6acbdab78c433fd06
zb6a4ce325d18e80c3506903da8b79a28d7c0f96471bbb318750a8b3fac82a7900bf042e7f9c0eb
zf1fc43aa684f9b21784c64580e74791a0036bcf646ad66a35ed9cacc4d0031ac26738e3e86c57a
z063c26139cc4752f1811cb1da9ac1e27d4ed89abff1a13015647e3afe022d8a547816a54bf6200
z8ba6f65271671bb626dcc91f7e3d71c5bac014c19569c98e6edf0e56faf0dfebc0f22677067672
ze55b7324b515a50a9aeb346d364aac9a4ff0d16b06bf9808804ce85d86ea82188e269486e3227f
z820f8248388eca1afa81d368056ee0bc20a0a79a79151a1e544a3ddd954179918718d2631cf44f
zbae7d64ecb011953832948f4b9d0fb6a00945c9e0e79c8f1a869639eba80e8110381d41e20c4da
z76009457dbf436d1f760af37e0e5304a858992ee5b25c5b34b055f0c1c45da3133f24fce8a8af2
z997e57928ecbab59fdee463c91de797df8354f3dc8f2ebc4de759ffd0ccbee5f2bf5ded2722b7a
ze303a652913783c37e0195a5e7f4139ae2a271e58251637f0dd5f3752139ec1a6fbe0eb78b9845
zfd25f5af97a484afd3add9c317c9f5d8f4edd353dfc20c142bb0807e40ebceb851e96660bd4b2e
z214c5e9667d5a50e488ccf48bd8d7b5566f3df4675ff39d164947b6ed8753cb60c43155d62e9c6
z140a7fd9445878f41c1a345da535e26cea9edd6b39f3a33642174ed5c89ff39cdb809c971516a1
z72358c27f848efe02f5351195b1a6d9747723aed61381b637e8aa6b927823c26a8d31edc78eec3
z1d440b0e4d5d87352556c5bfaca84e5f7ff5eb8429e443ea01ab4977b5cc201a1cc7a48935d1b6
z5cfe3db5006ba268b47b036e11b9c74de15719f9a32c766731201f3b9d4fd6ac1e8432d437da1d
z2c5ef7e4e3f22024228d9ba867fd71e5164e2ae9d420ec0b9b9ea17f3100b167d8ef881c3bbd9d
z93fa2f4db1c8cca38e394fd32b0a25f2c45e56229bf01222480f9ac370dfb306d0de5217f5526d
ze30cca115bcff082ed11672333d4a6910adbc8f05a38dfae21b183aaef24cb5be45d1648c5f0f9
zde157231d1d848cd06d0ad6361899be49bec75af886e176f55e3ab06d14671116abef4d13e49f0
z01aa1cd79d3e149d012a155e03eee8e0340e5d5aa441f6fc2ec556ba17da3e11d695a6f0f5ffd8
z9ccf90e3bca1f956e78bce070f325cbebfc921eddd5c80780c919ac92f3000633d3f9035efd7db
zb884b5e70f9f3c73af75172a91e8760be823e3a14b8264a019aabdeba60b344b8656c9776de6b6
z63e0d8f1dc4b0cccbbe06ada6a4bbdbbd45d809833db7be6f6e231862b8a07dba435e04bb1c4d3
zefa75863e90a86566b2fef3b6b991bcf7de7c9769dccb1456e378d8a0bba1e3e309ac61aa54cbe
z38114319d3d22cdaaba2a058d557b134034407b264d0d6cab000cd28b4ce700df6ef65259cc017
z311f6fbbfa8d9f04aa8ad273640350c2ace62e71fe4bf7ae0ceb455dc6b5dd0906b6c1612fc46d
z5c55752c0b795b385d61ab700bc6cf686e05dbfd1f57f2b5787b533294c9233c1792bad0e7c2aa
z0c722d3df8ba95d4283303f1b4311782cb809cb5e7ca9e8aa74fd39fc86ba4950c3c0b1ed29bf1
ze9e9543c7adf2215ab5ccb78a7154ffebdeccf8b70b9c0abcff663eb1c4f3635f29e0700b03e43
z1dfe338cdef9e61709d53b18e154bf6d2c1e650addca6a3021bde8de398eff5512decbb787c057
zc1b121c45e668d4a15c725e2d19429c835421f0402f526ec3da38b1a7850b5cd0dd3f23908faa4
z5b45a4e8ee7ce8a8e4e5d94fa29e6cf1fc5e22621e9c485482abb6f4a6caa3449933db05ba5438
zfdafeb219b1ba70d88115ef5c818619f9caeea7e6ef385ac0c189e496552a94d69475bd4016ac6
z41660fc9b3974ad1c425295a280d6cb8d8d660b974588fadf91e0d218b91f911a7f65acbddb2aa
z78edbd95ec2f7e1ec92dc4d0d607f6b708d30cbaef8463138e92e24439c0d97e9580cd1d1ee882
zdf9e97f8a415f74f08e2ae31c4ba29ffd80322fe7092669b8d3a7c951643b04c7f61a947963591
z4365a2446c748bfda22c9b459a8caf836d46bd1631df29a69fed36a65ab6d773a6001f448ad9d3
z3bff3d86348a6485657ac3477da45ed6d6772600827067598083fb7ee8f83b23d4b2646ae6fb3b
z3832ce80d37f5d417cb2ea326179fcfad4eea3d913e4611dc03c1a5dbb25373c1666937c54a540
z6a791a5fd0e58c8f89a00a3e13009a25cdf1203fb1ef16e62e54519e576bf5120a12d2e5f07aa7
z0856721ff25f49360490ceb501121e4923f95032e8be88d92de033cb6d85fef5dcda8bdab23c93
z05756c88ecd36bd42640651ce454fa5a303fe67215c83743af41829a44ba26af1918194067d8d1
zc1f1062e767a4ead8349416826b2ceb7173653f70ee680931ca51708114790d63ef2a3d2c4ca25
z32b7401dfca84d5ba7a4714ff3df5c98375dd33f9a14359476950c1e4cd26f7bf095923ae4b71c
z5733f937bfeec3f63c181883d2061bdf0d80fc75b7468c5d3939a64085609780a89dcc1275b234
z8f4ab3debccf8f4e1bd63619fd83ce9515ff7c016c589da39ecec09cafc51ae81ac4c74eff3388
z19ee9c100cefb6d61682ab182bd29e36063d744839372669784ea28664fa1c3a5aa5e05043479f
zcba21c365b2c232544da1a8fce7c9d0e00883ff9c5511b46ca37cd876dbd375913a6554d510722
zc4f26d4b79090794b9d781285d8025c675196cf99dd6995d6743867a13ffa4b6bd14af628a1a95
zed05f6a2e15a47709647939b0d261136d82eec0c6183fb29bc85bfd64e4e3e9722d94bca5a1c0f
z3c1a984becaf3ed2c0b79b7905acd1085d0dc36b9b5051e5cd232e2edbabf58dd044c638d0b862
za9018f773b0bcab2c5837f88724341392ebcdbdd05080457c36d8c9cd6be8221a0d72768d3989d
z6cbe3fb35ed86f861f79d810dad74a73388e6d869538209fb4a69ad7c496702149166aec12a323
z4acde78c4635b6c9b05d989ba9aa03d6d664cc85332c8b98a4f8a36c3b968b7b1abe714250b81f
z37fe308743692baf33afbf168894fb92360309d336b3ad95f34f0ff3252263dc19a424fdf9b472
z06b8f892320777db265cd14e5c702e5143bb1d9d8ad21bc6a8a87574348e6816010cc0de33cd7b
z77339796fcdbfa973580d5ea5965b93dbe3f565c538a26287c9a1a4c44c01461a25fc74983d066
z32e66ef41e9156dd0d1eef68d3cba1edcaf4365cf2446c33947a4be0754fbde660b6b5641cfed8
z5f4ed3fab61065f078f2f83c2ccf60f12e4de7d0979597de83a20534dae3c53eb75ed8a8b760c0
zeb4204566b54b8dfeca261fea284cc650a04c1d64cb11f9cd0c9291a90ffd8d8dd08a5fcabc847
z593221be932ce54c9547160b8a0a12e187f60ce58761efb753d5acdc04921d6398775c8136aa38
z92c2514ce2c7734f3c78ddcececa3cd3d307186948cc1c394a25bca2f31ee9d4c71ac15a138f29
za74ca664677e9681ab00396f160eb0c8e986f30d25b8317fa7c14e61c0e514d70899705ad7009c
zb26c15e047534a8df1dc1139f6a50d8b6d46a6ddfa2f6a8067a12c94a0c3127983ddafc08d00fa
z31afe7a1e716df9eeae843be8cf3301b6cbc286ff9702ae969423417228f7cf3c275cabf05f31b
zb350ae7b969c79e3da42dbc67173aba3962fe916ccee526564987dcd9245776731c00d93166ac0
z5f3bf3f7af130b5bbf0975cf2aa39a30f745a2dc359fb0634d03eeb1555d74b36a729cb899f5e5
z36fb12f42c9e424d809a227ce6424151b0a00897ac57037feae04591d3f081af7d78c28932a68e
z5e1d151ab6d7b787539b3e4b7672bdb6265cd860e79bb31f6487c225a78a52cab22298c1c7e908
ze912cb01cd1b484114ac02bac4d9f72c99f9662edac9ad01551e5d67704a37bca6ccac65bfd090
zdbf02085ca82c1bbff62bf896c06dd72f7bca474a7ec74a50328ed9cf9f12dd54c52a0bb0d814d
z698acc2b25aeae80fccbe53e92730a846f615b7a0e69733675a5726b868e478d9caa2585038c0b
zbc45e2eb84014bfe0584b7eaed587070d274d9f3ef2b227c9845f7b41c3bdf1eb0db81a76d6038
ze94392849e5622d00d7ff2cced31774627de255212919bed1018cb4c61660f69a9ff7859bfc2be
ze1a04f176330f6b188ec11f312334bb0bf7792bf18a6ee45c04a15b99bac24e8c4c2a2b6218320
zec5552bff5b469620bc9a757a6b2fb28fd8064ce0a09363a45d814f20c83d811bbc78b5ee0070e
zadd344bf16142ac9a9b66efd00da55e2c2967b1b2036a4e22a7bfc995384123394b0dc64d61293
z0b97a8f510d0cdefa75e41ac7168adb3ed6989d4e0bbd965e0db13a6781d2dc60083a6f534ec73
z0697acc557d6ffba394b5d298790258484b6ebce37685c16638acbead3c3a1e4abef1fa05b86f8
z4a3bb81f76253dcfca00590f3197d172a7367d7bdb3ee497453b49839b68262ee687efb4917e55
zf7cb8d3f430e374cc68f5e37135ae7e9e169d6385d6a818e3ec0ef35334234efe278ec464431ee
zd78640a136ac78f0527901b7127183126a5ecb00ade5ae75d826c4c222542e41c7271bcf46f6f3
zbc02a48c6cbbf3662379152e876d410922a5284c3b653ddb19b718362a23261afadda400e75edc
zf7812159951d68324c5d0d698c25d8e0dbacd240c1c99cea24260f2648a77538ae39fd71990824
zb7017ad67f01246c067a22f3d41e6e80bbbe503bf97738da01f618ed02186796badf026cf4ade3
z470a67363453dd86bfc37a8bede1ceeed55ddf02fd011e355f88bd7a6a025858973568c88c1204
z931f76df137188a6230eddeacac47b4aabae4b2ba0211f58317a07fddf77f3f69d34b7249b8f4e
z33970006c67eeb24831c1cf29fc6382e1b0d3fbaafa2c8d879064dfa5cde2c317d6bc3779aa4ed
ze160a8bffaccd924c9e011d796d569449a00a6e6b8dcf2bd83534e56737039d8d471c14994fe98
z0789a09baf8a75c8c0078b395ac0816c3f81214483c0ca694def1928c74308d759df9566f59b0d
ze4a3c5426ade01d5b412ed1ddd1ce90dabda59d0e063211cf2954ba19bc7d96ba25a30ed73718b
z4d42c2625c541e0f30ff5697765a3839a1c844ca86f5194d71ed54feb913ae204ed4ce6c61ce8e
zfab6026d3bb077df0f573a6bdf234c363f05715db81468cef37deee745dab111fc3b638b28f593
zce325a479c46ece7dff502f0f1390c4bd94e7ecb6b0eac60eb7e1d8a8bc62c543f16a0224fda1c
ze957013ce2a662bcd5e816325068577176c056c409e66fbd70bec8bfdc6d3d454f6e3a4f1a9fd1
zb1437d52e37c0168a5a30fd1efd6c5b3d45c7148f5de2651bed7e9a90b137ce76ee4077ae18b97
z9476ef31dd0aafa18132097b65808e915fc33c0132f1e92eac682fcf4f25281570de5dc98113b0
z8cb44e19d4fa930d6833bccdbb93a86ffe619e570487aab46955fb157afbc9dc1858bafa1f90ec
z7d539c10152c150e73d19b694e2146d5e2f6ed0aee4db1704103a89d797fa010affc13dbee9271
z93b9c8a4dc84e96ba97ce863121d6e56bddade16ac612cfe60319e33b2aaffef1c58a8ba57cf89
zac800b7ef75f7509418916a22075d932a4953521b0e22359234d9819d21fa45c8ff00eb1a84f6e
z05b8c65c31b546f0bf166ec11615c7ea2eff14aab652c190a96d1a771137e7a44530ccfe8fa4e4
z59c14f0ade71bad85692ec9742a2426ebba1d3191ddb28a2e60cee40baccabde5e16bfce5f66ad
zf0cdc71e6201a2450d923755d9f52d639cb73878b50125bca3f33a2b57bd3e8a634fa9c38975e2
z241f4fefd4f7fdd9b731fec28dcffc71b2d18f61e572cbda6b8f7c5f1ebf7296e66d6f186b4bf3
z229635789c9ac81e1c6d804253539a973f4c7fc19e130fa831139816da4f76818fd75230f25bb0
z3e75fb0c862e5cf8e756aefdc59e68863383fb2607b37a12f3b47c36557b80079774296f3ed874
z56426263eaf625a410ea2334cdbd44086fcd675fe9504cdfb83d3b85694b169cfe2c6f265aa2a7
zb10391c5b9de4e0601c4d9b24f8747f56435ac361baec42e76b32851e5a1e952e73bde7a29c803
z36897d35d5e50b5de68fbfae44bf3b4026da38360db2dc7cc21fddd52b2ec4129f1dca039250c7
z1aeeda3bebfe3df90bac0ebe3ea21ec7a0669b15e62ce80acd0fa89aa2bf18030b562cc44361c9
z82136fd2af1fa6d343a765c4d60bf0c77bab42e342f3081b1e74a5d38f968aa46d65e2641618fc
zb9cfad5538761cbcab497850cb59aa0c0b63b1b89fb12497d08f447b6be4c0a2bc3b437b15417f
zd3f22bc9be6b6413868abd494b0c38baed953880d2d1fb770ce601150098e1a3612dded7bc5922
z6626054f69570e1a2c002494a709636ff33c9510a5aedd1c21fda682602ee71b718cf7e2ca2d58
zc5d9ed51b650aebabf60c2238492d124fba24dc92e6f69c67fd75f2bcc79e0cb4337d28de16d72
z8105afee6488318430902ef26a5bb1cbca88b24e356c29318eb04475e3ecfdf543aeecb834d3e3
z04f624b985e349d0020f57ce60f6d858b8b3fd34121c4157be0769c1d1243af1a9a9b6c65584d0
za9a4151fb270aea7074dd4f55c459eb95b0ae54e7c8971ee162bfef632e0649db579e6f7474630
za01076656c88ab62f34a04dc630e1ef65a53a44ab400a1957d2d17979ebc2b4808413baa48fa2a
z34badf40b7e568854bef1e70a98d3499e39f40b1fa010eb6633cf64d43010cb4d252a46ffb503d
z45bc49339dbba0f3fe53dc84fb34a824f6d7bcd43e7199eaa7db73708af82a95fff22cb8868d42
zc4e0560174854555e2da369e7587db55ef15e352b84d623f151046ce8be40c962c4dd9db6c1dc9
zdc854761b8ca47d7d1eac6556387e19b856f4df619fd5a9a09a9b4a2744a98ffc053d259a1e335
z290f9aea067de42fdd70ec3ee07e747b78d124b3cf54882f82b60e180bd3ce9621235d0ea0ff4e
z1c7cd4db2dda5c08fa89c214821f16adac07e54decacb4878107f49e314b4e321b22d07e81d162
z4e63756df1ce35f69ac8c7a5b0131243d08f951e773c4d316925be0c76807a328e11e25aef849b
zca7f6cfa05e0272f7c7bc8fc20ef9d55beb6d0c74d55dec12e30780160f108ac156c7827613001
z2d2fd5c7e7228d295d951c740d7ee9a31c0ac74463a4904c7757916b74e28a01215c5289dd2f0b
z4d7ce31f06b4dc7ccd3babccd9338454fe2235eea01b434f1b8ba7d64743dfc29ff4ef336b9bbc
z37737980b0316cbadda29c7fa57eb47911dcd1cf9ef2e0ccabf1c145b3015d88edca09b1c2f84e
zd48f6ca0ec59b90a39786cdaacce8fdf221b2c2a27e38d8adb94dd70fa360f45eb2507ad84b7a2
zd40a8acb644e80d7a064b4499e6019dfbdff9918627c67cea2cf1bc9f95a38c6b8074ddc2e9679
z6889e8ec034953a2950b58041e15f6cc140907eea27d93a34341d6130f82e9da91705c8b299c27
z82ecb5d85d11985b95a660eaae363d4dab32cab8c68cfcedc3734d81a570a1638fd083202bfdfb
z72574ae188fd0d997c601795ae1865cbb3c232d15bb41da8b1d059dcd18c59bc23c5f3b4b080bd
z832e24805b55e9c856d0b249b6fb34492d806723bf63b61c9f4a1e64977a130e895dc783bad913
z0ba6bdaca43700b5990289df7e42e798bab4ee17f3859dfaccd2b658412f6d62b2533d97433eac
z1bbe4ba8e4b957a023966f163b947ec0f5e8578a023f9cdce8e03c6217a21be06c1a80836d6ccc
z9eabb87ea3f3b603e5d210aa53431f18d7efff80198701146472ed2827ddf5d73633b44cb4967c
z5b8023a8c51511ac70b3ded9e71086fedc6855ef77e69b9cad378241c8862e8e06f753e30195f4
z207f5646c87016bf031ad2d916063eb9ea233c2a7138acfd34c2ea01e836db999dccf8db5c4d19
zaa1379e78995f6d7acbe6df4d879644896a69f04de6b9e00885485c229b013d5b46ca572434aab
z47b8b4582d0f24be9e39ba0a26fdae3ae580230f895a6f95bb3e559e43ad9ce2ad0c31d1355a2c
za823b297f7781e0a1e8163ca2910ecd35ff2608227937da11e9d17d909f703a6d08b9a06f0026e
z27f2f43e2133f01dc10b65899b35961165eae440a9ef463af060a75400ec2f13d7c0c6a4f5a3fa
zed9fe36952afbebf0a6f8a75bf7ddae12d30bdc316b6c00be4e805e8ef7b8ef7836f9c9ad7310b
z8ae7024bf57b29062a40083d3f17bde4be16f873bf2f4527299997ca4391b0c730a55c69b0426b
z585535bbe6f2ec89962368e89937efa96e3c1e7b35dbe5617e8aab5df76dd88922f43515a341df
z0a8bbad2057c3359ee5bf50de482f46132eade041d22ff3ece698483b4ad0ba01cc02266af6621
zf6fd6ff12a3ee9bc580d51882a271c46cf06c3224e13a5d2dc09f33ac597436a7f452610ddf04d
zaa4c2832b895d40ee8c5713ee2a64a3ba34800486723d89c6ff26f02ee21408a748eb7d4dc1faa
z6b25e24a5606c50299798e9a89c6dc2e6e19932abbb653cac36d24931efe030ace32408e6e31b9
zf6119999fce6d1261a290ae3e6fb26f9e4b7fb41c895b3e1e7cedb2e82f1ca5b80e8ea7103bcba
z1bae53915b62303538995f6159c4988ebc764fd591c6025dd569ce77c7f052a01b101801989a3e
zafb691a344d0dcfcacdd3dbbf305517675d1d7f8ce1529ba8f91fa84236d426d0919c1f85efc8c
z90787a0ef5b2dff194d479dd1e94ec42f346354a6e1505a7f997dc9fc57cba441c8e153d6093dd
zcb5390154639800df4ba6342e5260c3797fa768cbb762353356f9e2d7f2b7ed4ffba596ec40250
z60ac6b3a9e58217379217cde89c58e7ed8a56f699ff02fe87b252a98eb1c00adea067689448359
zf03383f7efd92ae1db32417bebc1acb4dac6275705c4062bc45fd374cd7276232933b825f30f30
z8e94614e3967e1d5b3469faa89909a645fc45b4e1b27c3fdd6ee0ab59ec3b8b35de9b0558e1425
zd606ce3118e80f6db65499c2f500fbda2d37ebe72de3ab35fb73a9b8b722acfe6f28bf46a599ce
zc7d0fa1bdd0b7438bbd294492b20eed5cf757f089f83afcdbf99f1d5fa78334edd0ebdfbe97d83
z0add8302c775b533e8dfb3c3b3cae8c09cc67a98a3ad1c9faf23e434f5efb3d3e104648baa3871
z51ed53353cf346482c071152fc4b7770e95cafea6f81a8424ebd8dd77db8140dc9bd793ff7d4f4
z21f5a317a59b2858d2012cdadb41b03cbf75ee3b4a51777659a8ae8ebaf7b8b5edbd25f473e6c0
z543f2ba811d343070f69bca3458df7d1f56aecc1831098db9f8b426fe8fcc9d367c9e7fd7bf1c5
zc870dfaf9237504f6844640f161a9c249db866370a6b60fc648bdebe2efbca8b97fe50de2a62d8
zcedf863129d3edad73796e06a0c40061ec2e4c5137b946e82bb58a60568746b0cb43220c9df2b1
zf2e15fddf4b6f007ba971d26d9b0525f6dcab501e51a595e087f21a8f423048dcc66acde96e83d
z342471b02728ecb1c57094868d0039f8600a8b9cbf2460abf29b3aa4cc4541c1c3dc9694a68ade
z6c26aeb1c23cfd2e98ef4c3e5ac95c9724628cce88b32549b1b750b1953bd083cc44775f8d6c3c
z1b0c4df598235200f010d72fc76e0d07a13755931203f17727a144487dcbbc0289aaf6a11d61d6
zf64a4ee13314792963c801863a2b477e8f0f5ea615bec0d3b7aab42b222419613b753a0df1d381
z89b390ecb150443af1dfd9ec9038c667b984d33558275be2401178ab25ee73e2ec5337ee3ab0ab
z5dd6656c8ae1cf7054d318f5a2bfcc8194709e0f4af10c7c127104b45f247c495450aedb05e60b
z1f32126903bcb174649d97fdd2a3c6c0295349cb3949bd3eb0903d8dd952b3e101e48dfc5e6fd0
zd7ac028b5662aa886e3102166dc0a0902f1642b4c5385133c061389314621ca0539da0375ebe1d
z9bdf59930ac5dc9e8568fe23f310a6917a219191c2d707732b3a3f4955b2210ac4c987371f082c
z4356db0e3d6a5ec0d9d5dbafd6584f717e801c2a3eff2a8aae013237fa1b6718565f8ca66d1b44
zc5ca3e47b09d2c2146f0bf211fff793a4e282f8611c647dbca4334e3c20f48d942555a418aa7a3
zc3364d4cb2a0b3e4ed9da1e1dbe669f740c462c7b7742424204480cc9c155310c5ba68812d5441
z7ccb849a3709a5cfcf2f0ec2589ebea19ecb5cc1706ec5ea93ba9b98715f7e9b932fcd79f780ef
zac016a597d6f17fc8d67e8217533c079241a85b53275768432de77f86efda9e63e6ac7f89ffbeb
zd15a6583e1a8066efe6a6ee808758855290d24a58e47e1b86f78794419989a8a2baee1045ea5cb
zc6af97622337a99440ab72ba1a2de05b9c5348f3331467d2d51a8b341a2d223889f57a506f43b6
ze32a90d7bd52685ffed67e133086b95e537a9ed8b9b13d9efe0c64accf691b17130930cfa1a720
z4e6465ca07ab0c5335d05824917f78b7dae69814b4e51ebee7229dcd864485c24666f0aaf61945
za0fb82f51c459563981c6bdf64960278da81eedf3b8b908e091a53a1a29422ccb537fe5cd0121c
z8ec8478c3c72afd40ac2301bebba1c691d96d2ce10cc4ebda866298a4d58420419a84455d7c082
za40936fa3ada5b70ea79c6860db077dd59447b33816f2b37ed855ebac9ddb79a267ce9daacddf8
za495597013cd156fc59907e20a2c8c4a1fb37701787dfde3c1521305ee4b52b3c618da5c7f458e
zef51755635daec21f4770eb66e84a87090a0100459b6ccb8e15f1a32dde4f45241b47d5bfd22e8
z9771e761bf0358a44d65ae54b88ab8b4edcf037277d421b253dc121f9e78fe10d51173e092d00c
ze68ed7184b6355e2262880a778bed1c27bf7c1570a69ad16bddcaead120f8fd18139cef99512e3
zd5870ff7aad56bbd2683435bdee72227e5b765372561df8612c1baaca5d1efb2d04574059b5ddc
zceaefb94fc690e94890f4305f08a6d1077e03b0b063a859b2ac553c455b89b5b3d3da6f90d47ad
zdb2b7c8aa169cc7d41d39c8ef714b934ce02eaa3aa37ecf621879ee71fc667867597ee736ffbb1
z4938b7a608e17f26d9d95dcd216d08a2a2baabb9446c573441454b4647a11525e72ae2168e93ed
z5305fb3db9dee6036d3bfe55915f8ad0d2e5e60c8485dd2211f35274000cd8b43946e9fc9c758f
z192c2d2b2645f4048593993c4e7b4200954dfe021e00a2ac9f1be88023024d8e41d8ec1aeda428
z2004596c271289ad52d3a327f5e105ec40fae67996242fc8cde47af50ac34ea193f2e9c8780f5a
ze32e8d9e70c78b1b3bd157f7a0df3649074cbfee4bdb2389176b1c623348fdc0190eaf32fcdb80
zc2febbfabd89398de561cd775934368f0f343150c7a4522d52b671d6770a9266b8033f1e774eec
z023687fa8789e9e4f27f1438d69a8c38e097a8f8037eeb6ab3902aa86093bc1f8e70701f8337d8
ze0101547c4bd4e59b2873eff2b7203c3402583375b82020e6cdedaa4b3c5138919b2d0917296a7
zdd93f90814a634c82fe15867add00487bd66883898aea24c2656194270df34896317ff1fe580e4
z0f6cb9f9c6d24040c84b886cdd8893ceefd79c2fedada9924b6c0cc76718ed256c1ec89f01a198
zc8190c137b53be7c808889cd92ec634a35d272ac15601c643bcef30645ed4d2d2139bb32334355
zbd2133bb4b22b3fb147a85a73b3f1986362544ba418495c8de85082844a3b0a878e4a3816e7f0d
ze017567df4955277fab2484d52007917bfcecd066d0034165d01baabcdcddf0dd4a87da2e4b0b6
z3ade96a23e0f2c2a34253a6e57b5341f31bee4cb045731b667595dc294461e79479e402c5f538e
z22cdca86f08b71d797cc99429a7eaa3888485997a715820f76bdc391973d6f002e45066186d4c1
z5225bb31ca715d87ad692831296ae94ccdd63162f1eec126f73b1d5e9ce37d4f7b425f1c578ae5
zbf01265654b0ca671cb500f7b3821d6ae19771b9cd6ae864640102f5a125205edf1862c8fab4cf
z9b6290555499e2072fc0240b149cd10fd79b38575581ad0308ac97c792cb4e10a039b350669e11
z7904613c738c3238e36f
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_sata_link_layer.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
