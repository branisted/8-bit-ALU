`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d5983e9214a24203e048672cc6c97760cbec45b6d4
zca47aa20da997aa2fc510bd0403e34db5ab29280056f7174b73e079769bdfb4703e1517a392c6f
z37cef5a5aba52634616bea88511d2eb9e1f3ca88a47744037d9cc31d135fb8a791de554efa3606
z361ec6faf19239fc85b7b51b23d905d30876b8217fda24769506b70b8c6b6f558cf002b1502a4a
z6b1475dd5cf6aa467af93ce968946efa7df20d33a5df626bf58d0afb61947eda0d5da080370406
z26fea9c5cac353ac32a0739c36c84265e7a0782f846a63f23d2e9ca93ca90de6aa00fe9688d1c0
zd421ad115f06d9e97e70a57c1bfa2b1da3a63347b6795ab7ccfc54fb152602af429adb042deee2
z118b874ccb288e19412e1ea31b0f7fcacbab13ad15ebdea985ae181da1e8864045daaaf55e47c2
z1895a113b0f47c13797ba57af5dbb183c7d4984b3b465d186921b953170edfe189a3d41a9fc988
z066b3a8008e31291ec44a1a143390c28d4912433f25cf7d4139cdfae1cd1fa18cfe1af1e6e9c58
z04807400c693407653c792c4e20921074139ecc0aaab935eb626b809e4d38829964e44bcea04c3
z23905b70d710661bcdb46de44b26ff9cf6a433ecfb0912086a4cf2030b1ad6142ca1cfc7347b9f
z84dc4c25b8498dba6f13e82e515d64d8b491fbc6d95024869bc873c67c3385bd56f43059df2b0f
zb8b459acb7ff495e310447f9734fe22293f203b379783d883e144eeeb032417f8630d78926679b
zf6fb16f6963a27b31216770c5139fc0a0181f313a7bf3f055ff95c55eec6255cf34cb5956417b5
zdebbdef2e9a3585698a3465424a856f0292d8ef385f2a61b2f2ef78ab619cc816e4147db81f478
z2413d8b99e339fe0f471d4b3022aa5baca2d859a28e95446b8c1dd9c50c2d623787106d931e8dc
zada5f7ce75b6e1b122d35f9799958c9c52cd54e5a90ecf5e644724caaefef0eb2669384a0ab523
z57517400f695c2c69b00f92336beff1c4ae5a35995aae35fbbfe171b222f91a009cb4568a5189f
z846157f0a3f27f2c610957550e7fc3b103f9343e6860014d1a886eae7cb88cdea7113ed6f4c00e
z757037ee351d1f747c5fea17d394f5ed32382e4ad38c27061416bb03b4555cd52e7b44bf925733
z368acbeae8fe339692981d80da59a65e756f892bebb8198cf6e860d5cfddbdf47a763563f19d2f
z860d1378a699c181a7d48e03a06b84be58297e1f64163cbb9009e4c31d5716dc45e978eca729a2
zb16c31ea6aff89841751fc239dd711e33d2fed34d2e39dfed43ba8a2cfbec63c0ed86d473dabe1
z0f3b7c7553fed66332c05556fa116c13876e2b9da58e69eb071626dc6dca9ede2b382cf1739c92
zb7db2eba7da4884e6432b4c87da298745e3addbdb968619a6e7a5c6ab3608410472eada7ba8960
zab937711d184fe7d7d0e75f1cafbc8298b58b8993ab23dbf13a5fc7d2b096f28000992899b620c
z2ec6fc3a12ef4eb090a4eea7f906678f2ddea27433652fdd066a6190bd70acf3e04f4ab6ac893f
zdb763b041eb52abd22aec6cfa71f7b59ac9137675e3338472140aae94a7bb9b60349df5559c91a
z4d4977d4d91f69e32f01f131da5729db2b23677122927b5b3f878ef8ca047a0010d30b6db7c7d8
z4632618b9e89fe72609c09cd8e57679e9a5e433b35016e33ab754f941db07069e8dc9ccb0fdd09
z173902554a46eaf9aacc369123eac68954949a5a198779bd9bad6bb5dfb7f2c086a11fc5bb9af2
z54653b220b392fe29cdbf7c3eb5622cba75a579f900a6b391290722febf2edef8870cfd7582c9e
z3be064d1aceca48b957cfa8928c2b0d452371e3ee0a13a12a8ce5b2f310f029347b87be5d25d5f
z2129ade91143012b1fef37ad4e344a8c1e0b978dd57642e59a4831dc6b2451bba18e61bb015e00
z7339d6c2ed062863e64d1ec910baca743b474c2cd661267faa7c94a3e1f29c27c9a916ed57880b
za0832803b512ec3215fbc796e0a155cc271f3554c4c53756cd4f127220ffed109b23abf254fd5a
z45d4f1c029c042b0aea91e2bcf4c4f615394d5b7e1d278d87fa2d7e1ed98c11460ec8f259a8bc3
zd6dff50f6a60441123e7e43b77940496077ccd7e0cbedee57498b513d2bc5a50fbf31d81013929
zf8277bb84e1f2671b424e748df13644e6aa87033b9fd6d8d20c04cee5cb401c8c967f6bb77e0be
z854cd50e2187d15febb3f4c66967ec888a140ed8ffb2244735f7c349c0bbf7304cf8edcc88a64c
z693efe2dc7f6fa953a87124a0407daac3f6a7388ed72a964f895f75b101a7fe6543a72847ee114
zc8a54dcc1286887c01cb48fb4faf7e6b5a104f25ffbd1ad6702e1ddd01a57883ab8a7ca8f58df6
z1cd641a4bd64ef32138dbb15e733c88142dba4fd9962ded4037102f868f10ee190e52970c5ae21
z2ce76f00485bf303845252a83909b39d9346e35189c51b41c721215fc8a7cb06e1e4b2e9cc751f
z35e2139a56201a8cbbc8796e14a3307536d85e382492ab0322221b234e8555c1ee0cb003cdf9aa
zd6364e30c8503b6233f3aab7798c87936d9155d1e7f5c4d59f9c2325fe5d1ecd951a46c4548630
za0c5906140b8304487a341191cfcaad8a9ba31c7a91efbd3328c3685d3ee4f47e27240f7f39d55
z3d20e2353944120dd54298f9bead25c7de3bb30b11d44cb26620341353c2706981f91574b50250
z72f7a1dbeda1ededb880a6444364425fe313892694bd1f9677d585848536ca042fff521d4799e4
za8427006cd8c4491a6dc73133c55d0b3ebb42383a1465f841b939bdd10f98f86e3adf73ef3da29
zafa9fb4e4b47837f4bdfcb2bbf5ae162c99aa1ffdf16cf123ecca6f363859efa9b1bd5a7e68f3c
z2d042d7778ed2cc82c4abddb51cb5540df2514d4d9a9a6ed757b71f1a3008ef72d944613eb69e2
z7113bb52fad67dd754b348dcbfb0672111f95d4a7b79210c64b6db55937dac73e777fa9adb0919
z82c87e9f7dafd2bd369ce3cd66a949ddc7bec5c92ee5155688727c55396d2c0d98e768f178ca45
zd94c47668e37114837f145c9f18892d8fca52d318bf3a96258b4eabb0763feeacc87220c88c8c6
zf1e57547f53ad711f7c417e86c0c990ae1da741657a0c18d1b9606cc57995b33e614ce7f37ae09
z4f81f89a7b38c714b93ffc97a1a0f347c803bcac89bb6a624c9780c54256629cff8f2326bea157
zac866eac53cfdec9e9b8f57fcf34b503ded59e92682a12a36c1c327002b10e1d3618d81dfb70cd
zf3d5ef33e4a10d94baeee11fc28fbbf1c3b078c5fbb28d2306c0b948da9f7b55fd77318b4f1cc8
z9f2222ed6573fc96a6d2f513f1408519f4a9748faee3f332be17f848cbba52023505421d6e7ccf
z9cad7938a875a35fb72999c6058e055197de800e9c987d263b54c23af09ba30f7ac4219e76f89c
zc2734517bea2c8dd220eee9c1b8148b1b6edb5afbd5b34bf6207b395081dc6e097a0c6bd42c39f
z2aa7a04b2e47bc116c8a72bea4fc16a93090fb6a0fd2020667275177718f6ddf317ac4b15d9628
zde5475c9439c72518e289009a2d2b73840b11fa153c12196b813965ee66d10fa74ed96241594e3
za6e276d0c7a9e35b27f9614424754928a72507d8cb183cef85de7d3a2919a63552ffcba8402e61
z8687365e3369e62efe39f0c019cecb0ac74be3054a473d7505cfbb1f903f4501b47ec6d5e355f7
zd71762c4023caea686532b56af40b52a2975bae447ccd30317a5fe6f5c9322790fca751685d080
z0e0f740ab1a5a7bb918131ea82c71b25a3e4f53d2fc9c1cbe180483bd85db62168841e8c6e7100
zb228afd6a32289ce541f4e70544e2cf3a616c6e5876703d5968e84a506b3da05ecffca3b0b82f4
ze091d0d4adcb1563e348d2a7278e1a8fdd657a4b2b1c8a3c291f770fef7eea7173ab24f5a0fe8f
zd05dc06521f7a7762facc6180e22df0f94c7d93f561ba077631f15fb469795b5f5da8dbcb31ff7
zdb31d509b3b8f1a203a528db2a46524b37a56cdd7311522cadc9233025ffa1c385c140b1ef0fe9
z76daa926ee1c6c1ebc055b93a4261fc4fede048e3080439ebe2d53a7abbc8e38fc83caa1e1513a
zb4524001c8148a25f70daef84cfc9c2de9edcd6eb7ff3c0a7a18ec4e2f2df4659e432610ecaf0a
z02bb965c4bf9112a0a458c58bcaa2e527152206fe784bf7f1783f35c236b9fc1deb2822fca57c0
z832da68a43aad8c268eae57b2658db1609c8e8fe338ab1025e3cda95385fbfe82534c524f93569
z4850c44b66ee120dedfe4573e204f5cf2f27d8619031eff8ca397c31c6f298915b0492e85bbd89
z4e8d432e2eca08c42760d1b7131afd91186e39d3594517798079a44fab9e7d69eb45c12a454c6f
z091a6e927aa9999142f91b41935ae626b11ab2f06d870a72f80d574c43fd3718b2a1f4659b81ad
z4a418dd9d0d04d3e368ddb97145a08cf30a7cd683c43c0f80c6ed7dea58df6e720fff8b6d074ab
zaa065f7642ee2a17f38069f83be030a0a7ce51e85d516c5cee0bb6891267c60bca256277cdb515
z1b9b20b9f6e50e361fb1ba79b8d96aacf0b77917b5a20cffc0416da8e992d3ee839334b099cb61
z77e7bd0d7be6d1949877d0f7cf82a8dfa6fa73f6ad484a07ab2502a68973f697a5d460b11e2e9d
z3aed8e8b13b548428bc0fc1e8a8fe0baf35b0f34d869baa7b82317489255e3d794220d57e16deb
z9d8e0998cca7baaaa5d3b52c989a3bcf84d6dae327ea54afe5f9f2b8b8aa3668eef9184be92eb4
z1897e4ee39a81c87eed23c8eb2fe44ede11457d98502a02a6e3c1ad3ee7e52633a0238e1d3ed46
z3a60c3137c1459eec07feafb6491add0de24fe2613fce75add559ce8bac59fbb6131cd3b8da171
zc238f028168b5fc24042bd96a8ff1140ca1d84075b1172cc08c797781b98bc7b77a523783e1f4d
z2b397e1f109e18a4782cfa803fea34572ab228e81ba08d96106f8a48487f7f502d769a57e752f1
z6c06ea95660accd2cf26fcf2b870c5962060dd131076135ae8d181229c8b9ffde02ffced7fb2a5
z1e8e0c150fcdf7ffeb9c88b7743299d15d98451ef005939edc500ee6a5916779aac905daf64cff
zec06de92ee508aa4d888929d6b0eaa2e0d4a3c917a4cb505480751d2daaa9e0f57812d9e28d997
zeb067ca818e330c123495492b193a455def8dc7b78afa046bc67f12076e157472fa521d54d0874
z809f8dba6a7128af4e5da2e50f84dd3a0b09bab480f050c7750feeee577e199d15d8990128b8a3
z85c02a9973cc6f33fc3b6a46d04660983aa40b996be704bfcaf2f46322e971e522791e9da815b3
za009c688874681614e4e49d1f29485c14e99359710915067ef32a819d65e3256c229f59c9a6e73
za9e26ddaf8a26a1c85e425bc2c1a875b7a62e423cccd8f611c624b63917c6a114c3033f7d47993
z6f907b3faa08c4783c1669f6248f9204654e3542d333fa87bb0530e8ea8c9f099b976e7a655212
zb11c43b9814f18537c05109c8b8fde7df3f5c9cfe710b0ea39059c6a59fd40d6191bac862bbdb0
z9c2e59cb5018f54a0f8438a2888606236d2c7828cd6f89824fb9c0081551d5fecfc06481cfc192
zb9dfac39bb04f89be3b3cc7070631097addbcc00890e765d9f96290094f3c348ca0b8fffb2473e
z79052c91451ac3bfa5ef3154d870d9ee7fa3614e89bb5893991626aaefe254f00e3e356c53004b
z2f47aaff855d9bcf5fb03b7b02de6b5e3efa0c251ba68e4a528474c01ba9aa60964369f1975c2a
zbec8bb929847fe6fd2ccada5a3f59ca132d3a0b906091c822f0e4b96bed5a9b10d07def23bf694
zcd3e9b2053781bef90f0d8296dd214d2e386db0a25d7b372251b77004027e32e56e480df6f3c59
z849c22fcc7794484785a035d03c49dedc3e6cf50ed6d4c3dcf64ccc0aeaeff9dbf6b546cdbf823
zfe2d0a13840ef4c7037cd9644af9d5f488b64ae109d42140205dae9060aefbcb68c98bcc76624d
ze9a8c309af4d64ea223ad960091253ff0336b43eb1eae48351f3517337391026ff9eb081249336
z79641d9fb7c0b83a0c32d65798e5ca78d5adb67d037c2b282205a07c7ba2c0ed588d40a9a09783
zb88160257a4ee8da6aa091d97ad1c9dd8065f80a3c3b46ffd9cb8c567ff4a02ecabfb99a694f62
z1e7870989d21cba0a065254184d00f59a8ba097613f923b4b6f39d84601d91d27ce3611e86d724
z0f2c6737796d9da78e00a0f2dc4904e16e8830976e956492d83974e2ed17b02692e5eb171bcf3b
z7bff49abd12e48e9f69b505a599edd7d48813f9c53c32798a0bc918d58a5ff9281db4259d32579
z9163011d0d81e3a8a6c35625f5241ccb0cc1ad84dc7d2fc407cc467e37bc46dd10d287f15a42d3
zc37f8e54101a8799225fbdaf9027d7075783e41ac6a04250256e6981b95399fd9e95e40894f49a
z8e06a98b970374c09baec9080adecac2408f0e5ada2d5e195f036dc177babe032e8307891bc855
z020a33a299ba70378e15d627b3a77e547fb5951cb101441c49d3ea4c9225a66e9751c2c6d8412c
z588025167d94b48b58a5cb75171003ff76b87bad6139aabd01a6a5a0968bda10a6d8011f1044eb
z8135ed9ce626607b1eaa57a50ff4e17af8a7ca71bd275a6adb404fbdfeb91b649d0cacad33944c
zecc16429dc3312592af5dd7150f7067fdcd50010e15561bff289516fa5c8f2440c13dbb61be820
z58fcd150f72b3131864817ab13e3963e4c7fd0c184180aef9ccdaeb536c9b7f56296a4b05c5ea6
z8931cd9847b2fb56272b4cab8bf87f9a3e217f1d4cc9341653c25b279a9e4badbc4f0dd83e99db
zb496ef57f2f95278cceb036492a07d8eb6900606eea3333412ee7eb0c28f7c304e6434eb1c467e
z3f37c87a25ab044c93996c70fe82eba9528cb31bfc0858e7391e9c672473061f45a786e0f9ae30
zc5492617e298c96951c58967ba8c31cd1058eeedfa96f2715dd6c66e8600ca69cee19ba4fa8f9c
z2a9dd89c877ae6b11309b288ec7cd33bf5b33aba991a91a27af75517d40fae4763890b9c2f1c06
zf9dc996a12200373c2ab79a999f1845be31e19f3fdc833fa9c58b5de1c5aa6a98e902f66d0ee19
z87bdaafc4f14db1ea35b0eeefb78d8a22adb5868a62ffae0df1baf5320b6d98d50de5f70ac57b9
z3311324c9e11a16fb624634d75ded9fabd7da423c86aaa534ccfb5bb548d88eded9d00394b1be5
zf2339589cdb5c507161eb3682664b9bbae2f42acd7fea7edfbb058d0aba2ce86f8db8533502697
z9a6b3176d10a8b7904c9236cf5e4afd089a935578f0bc19da2d3d3277f33edff7934c06295de16
zbe27ee0020ad5a311dbb97c46a9f32ff301c61d28b2f159ba8dc0f5945ea5007e3cba82325bb5a
z6956624d6a3fe79d5aee860daf7fe9f7a064d98550ba6d6437c033a5270aabf6ab9f76e1dbc9a1
z8901adf32350df1cd2996ba6915d531eb28357b9db04724428ebb6f3e04189bcb15faefe4da7a4
z205bcb839104f768cdde264dccda1b47ca639a7014e22af81e18b45651732a3bf2534468fa504e
z84625d87b5eb6a2c99b7f0b61bff0dd33213997b31bd8fe180df068e02ad2b60f7ce2f7211524f
z2b839ed26cb6774253f4bf7fe85188527122baa18eb2b04406180ccbbb2bc61cba9c9ed9b7f751
z61be97faab6a64f80acf01da6ce9c66fbf431c75d8141b1ff43ccd0d6008c511a679cc5b9ec410
zec6cae9d0af576cc3bd4e15311a29a2fc83093d19e3ee98733111d57298a76cb452d18b97b5a9e
z114ccdea9a1558cee0d725ee9e8626043ec6ec395232b29445c2b96bd75c8064ca46d6d8a19160
zadbf2205872cf063f030c8445db800a9d559d14682e97fec6b63c8ec2982ce1cbedf2a7e2310eb
zc9df40e4e3ec3193162c42136ccd9882dafdcb39e7affc439c9f980e9e3557e761358f0293fe13
zaf8ace1d189b3531e641959208ae0cc5d4d432c18f8a4f96f7aaed297f84dbb996577791109d2a
z7d00607c76aa91797b21b05199a6648e599f725986b19a244c82255acc1a68840a46357418c2ce
z88084daf2c3f551f8b2c8019de973adc6f12b346d84901f7ef1bdb9f91710a9d272ae9ae09d233
zef5b24c910f89f49b5553245f7e08af91d4ba23cb6dbc1eab4ed8b878f512b2e8a92c83f742194
zb4daa9ba5d58fbd2fabbacbb62a7cdf8e73b741d1f9b175c0801918330f84ada07551e2418c06f
zd0eef986e2408052e060185c7554676d5111771011e5d34d73791c5e32ccec858307b8dc1d3cc7
z1b0be3f80d064298b4be1893abc5b96fb39a02906d3ddbea243f038da220b5f333d607db7c0aa7
z0565ea367e7af98868af9d2f095994cd915267fce860460745b11df0f7905b836043311f567e08
z12dd7eb966b0219d4937d8a44847b9c634640304acb752da0de3bb55d8118be657fa4fac148d0f
zc25543cecf86caae5832b669e1a44f49a47b9a7bd4143c88cf9e0c70a203b2dc18b0a438aa562e
z5912bd813e632c36a985803175e962c54dd860ea204bdb840a8e84af9eff1ae0be3978ba747b34
z6e90181ee26d0795ca90de9312dd2465da94129c420f790a6a6432a51d0cc4b4611ef5557470b1
zbbd31904fce9b7ef6f38b5443cbf3570a9f6834d46bcaab265edf65b5594c2ad458474656a4e31
zf87217088f81d37f9796f536d1d06ba9fba118d308a70d7c5559c2f5f3a364070469cfb0557615
z056dc8f5674a7e685aa8ddf52d2441ff80f25dd3042502f1d33511972a6dcf1da4eb6a31165248
ze9e5922be940357c47a656fc5352cd95b3666495a80c5875de67919329c0e2d75544c125555995
z691d1791b6fdfdca07da4e3540dc65ae3673b77ef58a66ec6fc4e6bab9c7b30ffbab9dc631b775
z0cc90dd7c99f016dc37b83b5f1e41f030e4ff9c4f51e0e9e025c1a363ad8f305b521f2d10a489d
z2a1750e431727fee8cfffe86bb3f0c429ace90ede64eba1c7fdc2904a93f1d043fda754e493fcb
za051b75442c36ff0e6ab56c06745ec2ff8a9b6c4918b0ac5179616678de1f45ddd1e1795579059
z35e61735db04abea259e1288e3facd189e640d0225af583b693d61733d9112f6797ded55980ffe
z2dcb2d778f57efd50681fc38349d14c4222d45b6e73925d53b529a46525476e666a938414e67b6
z52d2a90714056c9be61fe22a5b08862a7ecc645aa62e2da9114f6c38e7b1568751a14b454d0cf2
zda4c77faf3d7f56d90032430b5d1187dc0932d2600900caf7bd6ab67a437689a8d1e38f35648e2
z58f150b5135cbeb99658797754855b1286b4d4e44f8beadd7519a8f4856ea221eafbeb710784f3
z3dcfafc35e90475602293a3a89e22b65769f94a115bb17dc17ccc056c0ff7763b6650519880f65
z7fc870164fd0e44d2c6a128ccd781141e6465e43f73d16c5d586b73ad82708041e9e6d566d510c
z2b254bd3d17bd005317769ad524d4704df30d5673a2820907537b47666360ac38e022b3ee5db14
z8acbb7bab6ae6a4505af6a58652296d351be01d6ecfdb86fe5483df9c86bc87372468e368c9dd6
z5a5378f94fb87d30ff6606cdb76bebc6e233aee15e6a5b2b65a78f4562896adcd22a39594b74e1
z3d4c314607dfdee1796a5db4960a6bd40972d4032c1ace4b34bc688a41283b469b90d371babb1f
zb85c4b6d9148be6dac474586027ca081c53c8c9b975943b53fa08d9064d5f770a6
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_known_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
