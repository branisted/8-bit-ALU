`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff98478405fcd4d89273452c559f93e5926bfbc31a6dc7d3
z54b24d4be133c2e8791d1a3493ef5eec5ddc7946adae891a373c8b420742b6a218758e6fdae1c9
zfcc0f88130ea479e101a2f6789b158b79ffa3cab79e0623a00ea43af63c2b68b90c14ebed7aec1
zc141effff67906c15a760ce479019bfe64b8cb937169d03ec80a9e71b99d78d574a4424e625843
z9de21978ba8ff3694ca7b3319c0472f99a45bf243b066efd00a192c37c2a6fe73fab2d14bef08c
zb5888c12731aee1846c1ccdc7971c30821b279ab3db9b8e5525e4d229fdd4a0442d7623fc79030
z19de04418662bbdf8d3e9ea66256ba565830d4424b73bcf9e509e7dc8ccc8bdb53635a6daed91f
zfb1dc689601209eba7e652b3bb9e4af4d46b3153f6c116e96f73e2a246ac17d9cb8ac3374f25ce
zf7726d539f16f0343cae77f6392f8a8d58f03aabe29d2b7cc96abbf9e990ac57177c41ba322a6c
z1598ac93372b89f370f6aff053adbf4d8d389b0cd70c737cb8d9163a161d876a217b6f97cadbcd
z739b1ba86448c6a72f06d0bdfe802ce80c023d004bc82db4d5f9fe1255c77c82e12e184688ab4e
z4f2242bb8c84842495e71ecf4c5614dccefd225012524465efc51407d548d6feba83208e5e830b
za1b937711984f9a7fe5ebb25f16d5569cf826bafa4be86f52fa042f1d09b781e110399c24b0064
z96b2c0bbaab6af780776b3e082d02f405ffd420d664f09fa75c453b66fe2a353203c15b7843303
z5ac4aa6cadb092047116c35bb9c17ed14a1027f12393bdf64637f08f476acfa9e2ba8c170d4017
za10ecfbc407f6b5cbd88b43149ff1ab4e2c1e29ef320eacc4b17bf996b2ea4d3d643e7905493f1
z218586eb01a540cfbe68546b763965b4c5493e108b5ac6ebcc583e4592a4fef4764b683844f30e
z314aad46b3eeecf1b9e17733694acb4b7690829483fc70b994aa63d8d21cb422f38abf209b9754
z6817d9dd92f452cd74876e24ed781319a870104add302e8d3b5a8f8b1aac08e0eb308b43f7594f
zd3db330204cb10250ca5529a7fbeffea7b6c6b017f918ce4e4d0610c254380469d681cf7cf9139
ze75123af473a4ad61b27c8c854d74eef8ddf7e46694b92c33863f92d08dec87eb6a10d0edaba8f
z91279c1a302c3d1e65971f9ca127aff6125f30b9ed91e6e600ced1972beae1b95e2712057ca0e5
zd1d1ece124e549ea46a2321f0e0928a3e046f2fa4752e5002b9c87755acb4453e4f5a87da32edc
z537ccfa23572b92e42e7a3877c8533e6c6b6ccd4016c885d985881dd8f0d5e596ab5153195c72e
z4785b7a898832b55e322beef3994aa48c775dab22a5b348f8110aad8ada5ab8e72283b2d4ba0c3
zf1e3be104e958361da0ac27f3717f69660cd87a734a4d0aab4a95bfa93461b75ecd3431ba195d5
zd6ee95612c903772b0040f718e2006eaeab2724e66cd088c2ef4d9502db524980592fcf15e723c
z1dd1a3b38e8e1ad0c529d944688f0aeb3814c4a2394cacdccb2f12b83f4ee56771e0dcf523964e
zd88e16bea1982de33a59faa3501fa3463628c57f5daf454486c53812292250e30393c7c7b37f12
z4422e479a9979161c4fd70f99283e5790a875914da6cc08b8fb5e5283d7c878e82b87a767020c1
z186d5c23d772dc7980510e7b1d68444b2d7067d74f978396326465d79802cf84849b4663d78efc
ze18224088df76517483af888752955f7f0f8faff073623608ca6ecfdca7578f02286c953abb061
z260e067d234286c2f9430f56af10dd996ea6ca6dca8eabefe104e569a4164fdffe400a9258d820
z0de56e9a7982780938a6aa30fc84eac3f10c411144800d1490a08ff9ba22eeff41bf27d0dc6e3d
z471e020fbcb72672208ddc2292d33be1ce524315de5ef3ce792a8bf3854963648c3970af0f0d33
z7931a341975ea9ec160777dedb0e8d76591b1d32391bffe871594c1f7343a5d9b51ea69c173459
zc5d3f3eb61634177091965d16c284ec24677a63495ab9591d4009288e124bd925c22c0cc107539
z02affc08d2c55c4c60dabf05ded268edaf763bd68cd8e35f99b2db50f56bed025fb30716fa731f
ze94ea1a4ffc55292312fbeaa4fd0a0c24e5931920c337f707a2411dd4704fa55135179ed0f848e
zc3b13b1d2c5a34a8ea1495d5f9f224758533a782a4d86f1951e3f69e07075deaf666de1ac1b581
zd00b67277e2a8edb0a2b25bf0ef4d22e4fbdcd94128516141ed552e26281907126b9f20aea50d6
z7d019f9c9ff1cdc6ad29c712121eba583ee6cba215c66fcc0ef9660d0400ba802dc8a3022e21b8
zbb409627fd7c6c7bc959417d219fba1827d1afb1a3a85f8fe859178f698a77ee23f8d11dcef537
z85fa671e3dda98d2a385e5a40f4c72a00e3d3a5a82101f16170f03b8ac8e9d1b03370889d91294
z0b5f8467aee5d697a8cf620e9ed82341db6d77108fdf140f717515f420962d3a629ed27103440e
zfde7b03acee0a6d7d22b91fde8bdf4ee14cd79889956ecd42d20cba2fb62cbf2fe225c374d7b46
z6bb3e906846321e9ed9285194f34bafc701b46f295fd0d138fc690148bbaa9d8e36d47d82b90e7
z95f90b4b883e616f271c46a2cb70a10e53ac36fdd110491d6bf20374fc5d2d9ee6b1b8a19dd62a
zb8aa311604b3a8615d603c6c21ec5033dea733e1c8347f5a109bf7a94070cd1be8586628b39f95
za79165df30412d0034b88b69760d7c5d675161703929df788fc917dcdb4905d411439612ba9d5e
z2513557d322a5181e10f245bb568f735c0ab7e5599f8618e73a303220f7dac9473e59d51e69bed
z365744cca36b273a2ca40f478feb28f742a6ea2da91d0689893e3e6ea0b8bee8ca3277af76ba7f
za6f0ff06bccc2bda25561b756e2a6647512e84aa05338661aaaf2dd4bd231208506277be35e9e0
zb358a72b1052c6ff1b028d7a24acf897202f837ad869c61fb67360d7f15b566786fa879ddb903d
zcbcf999047ef99eddfe7144ab67655529f751e698903c5fa9d68bbb6270bd4506a6ee9518eafc4
z5c8880f67c7406d8f6bc1458bbe41f914588556412fd89919262b7d2eb0f605eb49fd30a260592
z30db3d2af99f153f302c9a9ca78da58802ed883ef5838b50d6de90d55c73099140f07d85b675a8
z097545c0bee0428e3486be2194a0bdb0ff7158bee1ec5e7837d6c8df725c844dd797e2ae26db67
z2a93374474e11c2917a9b1d1da135844bbee2ec96fb48f8ea2b46610112c65447cbde0a7af6af9
z6fbec7ddfbbfb0d63867d3a6359b37c18b33eeb62135e606c6894be72fc25b7abb8c34d9385744
z4604cb53f235c9e6d3f207042121ca6c74e82cbaea0b047e77898fe3e413c4811cd4e6a8950b91
ze33a987b8ebf944a2adfb27961d9153132266bef2a5872f35ca5e4c49cad8ac6b4ded76edc59a3
z58273fa3dbc0898f9abb60857a3d412b1676a31a9dd911f129862808a6a6df6cdc18d2b3f3c5b4
z6d5085b9bfc40ea2e6be9e51be952c9776ba3ec4a2cbc60834f3d8d1d6f81eff803ccfc0ca5f34
z650014c9c457f77c56b02e09c31793fb92bd5b024821cf2361edf85c5019ef1d97ec54e8c5e226
zc29cb296af2f058c5cabde999c5c55239683cb9a24081bc902bdb197d4c7ca00e0be0d96c519aa
zc8c6e08085415cffaa99972fb0297143572b8da6a9178c8cecc251b5c59a66e1e00f9e60f5718f
z27f5d347c1fbe2a906b1281384ac09c64753db21333915dbefc40232085a941f0e5cae5d1635fe
z3aa8a6baecfd72869b5257daabd13b433bf4c69a16c5e31edda44bcb9218dcec53f398fffd0636
z89a3228a40b269267364d580214f437d7b94260e5c05550e5e76a0a1e1261bfb497db2c18ecd95
ze026cdb5a0c3967e2e82f7252974f671b4e00750c05d84dbd5f90ee899d6121ae12f843558f0f8
z5f93857cca9a4af7af9ef4e3815de430e2233afd631346b32782fd561942f6a3034577acdcc2cd
zf1ad2366b62a6c8c4abcf0982c65fb3226b9eb0e012b690bf05afff8f61c756cf77510bbc1dd19
z759960730d73253f7ab9ef9d0804277145998a44aac302832eae57feae430502b541de734fc9f4
z46043a6debaefd9ca09737968065262c6d3c9ef2b561cd6afc1becabd163353b104535d2249566
z52126e4ebe83bc33fcedfd89b67aa7d5edfd2a70c4d7e3f1f6b0f3af2aff01a0dc8fb032fe8d3b
z797a8ef5b6932c52bd75c1238c1b7fedd5ba1f1b05f473dab73e8b179c5ab1b8d9cb9bf6867032
zd3b39f820adb45da286e80afac956d469c19b65960e0f7b6748e639a80afb17d79e45de3702176
zf0d72e126ddac5301fa12179ed456d5a4406e69af51180fe69265dae0ac6d70d0ef8f264c4be46
z34820dfd60daf91e1dac31421c4af7b50cae0d5b41a5eadfb12812ef9124708aa262505e370940
z1f6918c44f20787b57ed01dfbb8171b01886fbe6784b0812b9cd7195f06f36b5c9ca9681b45bdb
zbc518b93ffacdde6353e4bf672d16c3b6bbdfee8f1cd9e46ade14b9ff87df4eb80066d24fb7559
z82a2ce6032bbadfcdaa76b94088dd46cdfe558937ad7d1ba8ea3d453b8587a162fd7c9361912ef
zb7b65425b2bf4b0d2b29c791f8a292cecb5de0085168eb832a1084bad9686cca4e0768124388d3
zcad85bfed651ddc551ae336a06c37803f4f316c2c421dcaf4d079be323d060af274588e66cf2a8
z72a02df01459221eee3d80e9ab73a5858adeb32598007a390026f8e9096619773742d7d54c6e6d
zacdee31b7bb40f3dfc45377607b0aefd0d2f29051b1d33a43d38a08c705f7f34a1f58bac47c73a
z50cd568fd94cfa8d8ec718f4718b7bd7939c1ee37f75110e2ef8d653336585038d67ec5a8fe3a1
zc3a5d0aee1ca2c66f46fe3cd85720c5b4cc93ff7b6dcc29eb39ab209183f0d95536901675d98e9
z684c8ba8f9a031ceb7ad6b01ed5c053fb119c0466e34075b9b61fc2f268cd2c6ae1b3e2bbbb5fd
z72325b85a78090b070ead2c20331b12eff220885cff463e7d6671775e2b15bc66e0f03f990bf97
z13932ba0a7344f505c52b29a8d1abc2b5473edc2be4347df47cfe7a4f46a7caa7da434eccb4b3c
z900d9f7ea4bb7013b6fcd77ea717f448612efa318f97cc805a9ea264b80eec5d2976264d9c79b2
z2e837dac9b9e199adf653bfb8109652ea92fb2830a2b0e17a510a41b98484f608fbd1e577bfb7f
z2da7bb6c60e5b41f0f369d0b025aac402db9b95a219a4f8e6a9d5eb4d6775a5b3e68bfff0216de
z9633d073bf3303d36bc5fdac9a7eda3e1d24f7c2b6360f86c097b2ee505f1bc435e5e903b12a70
z7d529cd1507a45edc0d4e4facbf1e5df09ab0a8a214a4d6b3397d6c6e021251d0789a82fede76f
z1cb66e3d9a90cd13913c4c2ba421d6d87b8948ffda8dd2a5af3e2a66125d39e71eaa2712c5781b
z52cea6ae93213cc656cf36c45d00993247982cfbbcedd2409cd3fbada26a9ec0ff13bde6f2cf45
zd0b66528f787e4f15c9fe83d1924897594e3ce4b908ebf27b8fc6c400c0c5d95ab71ab7b2250a4
z14f215840768adf3d1480ee99f47346d3cbcf7f89f095af3527e62a9a4e0885ed05313de2a347a
z47d958b866ee62315c1d2ce1e78578b9f04376e48b452ebb453d5ec1112d6592a2bc177cd0978b
za3121ca89c94d9d8cde5f513171bbc18ab059e2ff292118e7f1775f3b009cd9146b7186f90c962
za7e4b65a27af43f0affd2f239af85a40e2920ae4511f6e751d42fa296f01e65638c517ba5e864a
z3531f135406bdee46970879dd48aa5c78fe64f0dcaa56b07c7ca1ad83ba66725b56633243b4c34
z1e67c05e472451b27cbddd0de8159b7d723d7ac12d0692491a52cfd7ed751b067ff6a1e87cebce
z3a33d733b7bda654d4d42a8c8f18002f8816487993d3dbe45c4a918a5edb6417ada5e48f1ab903
z8224a96712c7c6abb1d64d56ac5a1716610f62cc4c1de78ed0a9f00f4721148e4e778031f55c6e
z9e96110f4052f67c1bfbd256cde46e27708145f8fd7070b10160799572de44b27431b34a37a9fb
zd6969432165c91678198d0051bc6d456779e30121bfc88f4feea1abf13f84513bf0fec4cee3fc0
ze5c31ac3cc02533536a041ee43ace16b01e67484b4118dbdfef5549907a1a33fdb693a34f5a03a
zbca774cae6d6ca19343552eae76225c8ca334303639a67b6df0e651a3444e7b82db7db2e9a3f71
z4cf1e2dda4dedd129f8e0e86c29d5435f1b7674048ca63afd83e8df88768fc00fb4b8221c4dac7
z23769f8f63d72418bd29853bb487fc4ef5d03743a7c799e822eb0300223ae23a181f2efdbadaf6
z028cbf48b228c0cb2d2e80c4e1c226bf23e8543e0fb3058bb24579ec37768faf1899135018ad5d
z88c4ada55625dbd80aa8decfed80c9a93e5591a067f9a74f162c930b273dd26d8abb2b21bf835e
za3b0870124afa3e025f1f60131d07c59a7ef81f477e5723bcb3c0c8f1a9467162008e822f68f2d
z1287a929aca373836ae4f7597693c0244a3354356cb6a5e468ed2db4325aa442c9dd5ef08a8e41
z8503949633c47c66efc2a40a5c3e9e0fed16823c777ba6bdc3be10b92fb7f00e3c4fb9ae5b36d5
z2dc780231ee5fc2e1655fee38d4f45b0b81a29031aa1f643c5327bb35844566d73b4d814571079
zc33e69ef9f24b508e6416da9a764a8b5f515228819e83011fe1c5d79741bbf1312683125a6ab8a
zecaad536926f04996d12504ee323dd4756e1f277f3edafcd6f2ec9852ed4a275551bbb4e754e83
zf4d7cedb389511d1425b38a9bd984b402cae934630f94be4fa3583866a6650fccb9ff14dcc8091
z3fad00b210be0021e8c93a6a59d7d79f2091e87ff8796519bc02e26bdbb9b2bf8503afa7bb9375
zbeed2c9254be1a77076722a9226b72bd5e601fc77f32231453131c8ce0d873447111b500a372f5
z861511472efef27dc2ce7eee5a574463797e9a6151ef387c351f1b22e7dc76e9645eae7fe54ade
z58b5504012aa008f81dab85e16837fd4d6a2fcf78a9555fb61b2d3a5cae2e87e7ca390b4d2b20d
zedf2d0d3ade37a52d1c97a8f84cbc688248a6331ac005e8c840c7ecf3d4e3daa6925c287076f74
z7b949836bb4409262fddbd612d804ccdf1325c5f639e08ef46776f3ef72a81969d91539ae741d0
z891f48651a0c758418e48a7f6f9ebba67b19d2d56f5401929c8c527da092bc02f5cb67999dfe75
zb015ca51e20df4ece60bb2923b537d4e3ecf1833eab488a8e8077c2afd7a9a8440e5eddd396365
zd31c82ab250e2c12f263a782377b3944405efad47876d0bcd9b80b4241611f6d572964b87668d8
zd71da33e1bef53690fee822982fa0c7ca6687b3b9d625d8cb917e4b443091db0f82a1d642354ff
z749491fcae5c3b0d04edd52167080978aa034868827bb867a65a0f29cc48adf3c2dff226d4f06e
zc6dd8f1ff05e65a6d5b159256a55aeafe7f8160998295f1eefc62f450462595416a71f7a9fa8fd
za30ff2f7c8f6e71939f8666ac181301f4ec320604fc007f796dac02a4a3ebe6385070df8743e30
zc84f3b2d2d937baa821431c656c3d763cafadfe53db93899c7fac948d22a6cac14e0adaa07fdc6
zb93e2dd9340fc1abbd4a11e84cbe7f01066b10e28f08a7803359b1a22bda2563643bb235fa49f2
z64fa8e618eeb5a1e31fa638c182978fa12991b638f55745c31eed9393752c49d7a25a5a2415eb4
za88b23b04d9d37e18da4345be4d7ab1c3821ef11d89385d236c3c60f02e3c4447e31348c5684f3
z59dacb26ced3738a7feb047123295cb00bbc7aa8db1c0f54ae0c89e4b61c70409078b0bd4f40c1
z8fcf9acd16917dd67453afe79635af43862e8a9b1a4255f75a226b346405983996d95e024e3113
z44c6b751c4c9f64597e0dd73b6e88c5ef384e9fe7bc7f0fcefd52bc50584d668f12aec400e4472
zc20b2e6e590cab80e76acc9475c65b3c4b1a49ba149aca1385c17c0bfc192737cde674aa86a91a
zcc4c5918fef3469d44917325498228e018b0c660a0abca994111ef8b6576be86f408af280ef818
ze20e2ad79772aba3cd7b612fd92188541bdfd36e59ca60a174018cbcc77feeb5170f7466970065
zf9043d63b13302d176da98ad031cdc4f71a11d9e56078b92ce79b553564362e3e0fde67d08cec2
za0c6e5ca95a389dac75854973c97f536459988f287a28a70c1fc7c0a419c6f0c64a58c99c55900
zc4ea66ae1342603841b38d4cbf7caff6c166b9329dae6b46ed6aaf7994a61bd531db7cc11a5a0a
z8c21c8c079dfb5c9d1c95092fce915000ddfe89b6cf520fd5eca9fc307d4e7f9d7c43d580960b2
z01f003867c4eabf1be36bb809f936387f2362759539abaaf5200848b0ca67960cc661f5addce60
ze317684f0d0ac55035805737a791a0b1461494e4369027504cd3ffaa3c25ac67d67cf31dfb72f8
z9cc48dadafe6c05f08e76ff213ef4b15a129bdfd03305b2137481332d49008425c568ef66b82cb
z82e71e97f8a2e76169b916e005f1450a1d25890adab609e64a53d8392c727114b639e5bf025675
z6d430f6d6511421a87a378d2eb504be53a06cf67b8b34b17710c8477b0fe550a59fe5688e0a679
za2e6c6b68b753835b725c3e1ddb239f816ef813f6538647edd269a7ab691297f28b21bcd709406
z581c8a870f99b7cffbcb758c524eceaca5ec7dc1e962f8fa92c62df72da4691f21a5ff127c2b0a
z417c8e5b92ea3ccfe2520204d1d1a4ff958c86291f91de37881760d8d76685c7c20c4d2d39193b
z5d9b84c8ac057f3ce709f098263a980cb97b3cf47ed347de35d2ec081f4571426fe05b29ec1111
z8ec159d7a2411bec68bc12a7343766416249b9053cc8cd8a91b0d09bcb04725e68f44401e6eed1
z8509e27252c08b114de76d5394f5d2d285576035d2d395c5a85416178607382eb9fe724d918ec3
zf0e19f66597f2034c52804e394add69caab93989abf6fe6617e379e21f9deaa252a0b18551d4b2
za0b20dfdf366dfca179c89dc7587bbccc56935d7a1ac415a3b93369f26d0e36fd6b67d4b1e2d67
z63f9bf79ff0d923b37c8fb9086308f0d839922221a4753da7d8452f9b18d7ac43d6d030b541e50
z7afe7503928cdef4d369d9ae8c2e3d2fd68397ecae207b766e059fbbb83ade43ce9bb41a732341
z66c7a2c8a0b18e5f96443b993b15da512a95b2911cd321cab8dfad30f4dcc6529f3758f3e9914d
za498f13b83fb977ff282446dbdcd23002c233e6bfa8b6033c5eb5f317aa610ba5ef2dea3745151
zbeb36c7237cebce8b97e1a6b7f0aa9969510f698254ae24cb1b5376d140aaae2673a4fa9ab880a
zdd0ea568d0780058e40676950b4a215a988093d50ebf59cf4cd813479c1aca70b7a65bf00cecc7
z4ef000162802ff0b4c49f9b5a3d5c627d559d5d2d352ae5da7229a6f3332b109ea3ead3c67fcf7
zccc641b638124ed3fc6c87afb814ad6d7bb74779bdfe39c540dc9b35b3a8e5a1f0955cf391209a
zf0815415e9d4d5012b908f36fc90e8057f18b58212f51115492240e982619bb33e03dbff32b343
z31413a4a3fddfa3c5868e18d0c23508b7099f73976a54bc565c52aefc674e7379533cc517d6023
zb36f480585f05fa54cc7dbfa5e3cc9689e59b263aa9eaa5f649e02bd0ff39dd45422d334263e2d
z9bec18d890caf1be65d44ee8ccccbad1a1e46486dbdfbe43fa6c3a7e32449298d5ef16bdca5c2e
z5c7482c845db32f696f7ec078fb9bcb101ecb8d2cb04152140794a20b6934207614806af982b95
z3f31617e235281520ab46eedcbfaabb6080fbd3f19f7af6d652abea3690355763d4099b3502d17
z32388848039934788a9e5d1db07870c704efe13b4f663b39229386cc9093ab2cdd8e6e3e1db5d5
zc23216d756b27ba52af6c30e75806a5a0327a31f6d4915c1c2a3df8bbbfe251abf55557f50b72a
z58324b1a0a147f1f7e3f4abf3081be4b340bbba85a30b438d56f5776c928490dc78e04685d51df
zde03707493a851c8dc4e6d0fac418f0bbac9bf4a7e5a44c7dd39abe7125ee82feb6d548d134269
zd27f47c35df2054f30d13015e1272a4f6a7d1c415d9de8dd23c542cf182a9f8d825a71f5ec94b2
ze3ce77a04bf3fd0abf8f112b9385afafbf2c15da6db5191f835e7610619228837d1c6eec23a0f0
z26b399e9864a304fc35f5b3f699a433eb5ae011f9191f3b53d8da46ed81e50fc7fc413b937aebe
z387a18856ae2afc0c2ac426677a553729f4e0ca6899b0ceee0e6c9f4b0e387194512f6525111f8
z9a8403946e4943224deeb1d8542573815023d3eb637888d75ceb68e5840f2d2d018f2da066f62a
z136380ff2cff69a233712b8a8fb5924457edb2d7b7bf601535f5c35d8265b5acc9f09a35e44b18
zab66c8451625c968ed1785cae22b98a37d9e59653093e313200ba7b3a2f44634f39fbfe4d9e8af
z34e6ea64004eb4bfcf00e70761eb34cd154cd71c1ab782b2dc54781c9e0f90dfa2770ad2dc79b9
z1abf61e49ef81263f0cb8e2b50484f63fdf3d1fcd221218ff2374aa02fc858c2df1449648fff94
z9c8ae05a5efc02dc200d97f2ba00aa74bc4c1ff152c1c4d323a9c25cf4e682dd7508373726e6c1
z4cc26abfe3cc8369dfb1416f037fc32086350cb2e3d86b491b320573d34202c24e6658b08a0b0b
ze49d9418c454c515d468b91fd818fa2fdcb7415ba6323605762e4a774f6723a87b86c26beec3a4
zbf1291afbc85a3ad96c5afda87326a45c23fb18a65c81d15d833c1cd99b0f76b9792c421e078d9
zc529a63ffeaa361b8b8749850ec203731d39c2b7492b805e7fd6b51d63a5f36ac86276840d42f2
zc545f2b0f6cdd3d16813c1144847fdf4388d054c2a0de38c650ba65f70790849350d03267d7584
z40fd45ab87899c5bb6cc68f35c75a59e3ee128ff7e34d3dc43596b3860fb369ee909dee294b2a2
z31a25d186a2c30bccfaeaa91d1c83c5f4a5e6c4e1a5303e65a45b0f4a0c42cd4d19d07850d43a8
z67a492d680d3056ad847652efb0abec9174915a1d44f99b19bb70a04b75b2b3f189e2ee6940858
z9ef0da70a4f9c39d144551733d9279622283e14190a913a8be3e127bea221280062d24423ca4b2
z665d4e0789b5ca845b2a1bdb40342a6a1159882ea6b8286be5efecde3242231451c96a4936c3ad
zda6d49a28ffaf4cc1918dbba0c04fd60c40788805f3c16d8cd8a45927beb5005d8a9b1aa1b5656
zd9b6af87a28b48a95865e41980ecb372d3ce510eb045ba975c5a95080b9b5db0723108648b6e37
zce68c738ac3eeec959a170c030679a526da7b004f9fce0c653dda098c3c6f8314da8e5a8e11246
z06a12fd6e7398594fb64781c99c3b7418231522f4b5787927b771b9fb07462bfcc843f52b4feb0
zbc112f76f9b2674b78131ff49b0479f47a9ba199c59d53f1ba1160d0fb33ac63d7501671d1ea8c
z7317a271e41b7bc7f72ee9f22240b841e01d91146c452888ec98b321a52779540cecec42bb1919
z19d596687de4f22b0c9014d9c0f72f2b5b6a2d4db082b294d5b6154d5415bca82f3815b23af216
z6d679033d3034a1188399570ebf2c542e8357cae28c6cbc11eda326c67fe71d979416c66602b0d
zb24003a3cc76226f474e3b0a35d4a32ffe106fc6d3d837c8ae751e44f7b6dab9cfb1b161be2c00
z8b7b29ad2e68ed4477d4efea978d0a6b6fa0a5e769243556b9f260bebf9c1fcb8f725d45b1e182
z31e2e7ffee319ad724253e65e29c1051d5cf7d8d4fd7019a7bad0e94ab0ff9636c9e31690b5cc6
z63baada013a936b3e1f26da52705d3da2a64a7f2348e651a5c0d22efa2dbe715753c2b6e07a6f3
zb8096d113340cd3476fab3bd21997c3b90046c63fb6319e6fe8a88b5d78a15062695ba7853757d
zab2edda19a74bd87ea0b534e37257ee70e5e52346965614cd33ca37c6b13ad2e5a803361eabaee
z291b5f3dbfdad489922ad285740bdbb075eabd7909f5c63d8c69e53b1121a8067d9fc75f1029be
zeacf22943f69257ae7b8c8a3ac5a0342c90083cf0b90e7266f5ada93ebb0d453e8569359f57d15
z80ea7c793c971bf42a17559bb2d79b5d405813b6c7c4e0094511ebde7b1818625b7aeeba287348
z45a9b14b4f2da74499ba6b648cc080a5e7cc1cd4ab521d4f7db3e10acc29e90be9ad10a64621a9
zb3cdb2b5437be00e68041154a3cec757a44e1fafa37bdaaf226b1d0a8c4f54c76472b3c31e5f1d
ze1536e86ad08a51cbb0a7e9dbbd386e1e019ef8356b04ee1f726cef4e86caac2ff10278d464916
zaa1f1db6a16844ca74ed9b4b141c5a1bff44790ed2f68f18ccf99b03983be262cfdc127230ad4a
z36973c7f1c3f5cf74f9625fdcbac6d6b1c7f45e33ee3d35c9b1c1c2ee342b03b4eaf8779cd08cd
z39100048ca0148eedb9a68adfb99047ac5b49cc1f5a84b1ab0557cb64a82df55e314a4b49ff506
zb38fb544bbc8c1329569aec60b3bdd55fd0c5c72b99663d64f8bdbf16b72e5a7be2a003565e61f
z81c618dddb5e88c568d116d1323839eea3cc572d15f199fb6bb2633e4ab528c7dbe75b6fe70b7e
ze91caeee52167e64b14a6ef88ea07c57c79269a4d264d9e25e7debc63fc2bb77f25b11fbcd3bfb
z21d28a60dc68cc405ce537c3c6c2146a9798a3b476642dda90584c662fdf73e57cc1590bb9760c
zbb938cbbea8fa5d025b5df3d0b6f4d254a17f640bf09929d752b667f7ddea10b7aed10ba07451d
zf432aa5fc5787bd9eaabe72eb4daad270e62c8ada0985909d5177fc851286d87b19126917f6ba4
z1baedf434f269ee18796ae36f44acadc70d76f4a0157068a0473729fa1a3db17841a3e95f24166
zddc37d7936b7d8029e2b90412a01b3b3d9d89e3ef97df1ce941e5de2413704f8963368cc9dc6db
zb617254c0e5d186ed5ea64a90303924e3c26a7ca87c0d9bf0de64cc3135afbdb5ed4e6683b44d7
z891dfe0c3d01a28996781715e39efccbc63f4f4e07692ef95a088679e9e95f7f82e02cf167a461
zb960f6b3e27349833fecf236555430c192125f6c4aa5762778bc6170c6ca9d801c77fd76f6df43
z994882a534d27395e723989f1f81b6aad3a7cdb18f5fb63d4247eb0e58fb224b0707676ae43718
z74653759074fc575f9909515124f374a84ea9ff31b32b54a43ccb2900f477037debabe89c6d51c
z974496c6407d3de65708b24b2875ae4fa556633b52a187c26fcbb4bf15afbd03b7534d1d662b5b
zb39a068ee305d6b5580948b85fd8c71fe8ae597cf519b08774dcc069cbc3cf99fa7d0101cd0970
z1b7be536813893dcac7048dfe3de25cd2fd4296c6ca3ba0b25b55b5f8825f4e4faab64248090d5
zce515fad2b32b0e2e040d75deb2a36a1a2c0b13cb53eb445a0e1a8aabe719e85e9c2ba5c2138fe
z733b48c3e805f7c4726ee3b48a64b1d3e5c2f064000876f9425d87e8da4c7d1165c2cd2fcb3000
z3d9fa3e0bd1d74dfbf49cf4437afb48e92e41cf54e1f1e850aa5927d589d8789c1a8dafd03ec89
z295b89ccea81bcf74e254a83bf03d69a0f17763bd3b75036ee5acb343e09dc1a59597f141504f5
z1b6fe1b6991a6e30a0b71977ad0cc4f084501a638579dcb5a955dbf413d6161383aa8e0a1ad4fd
za142d5745e1e01714b36a207838045cbe271d0048891f39676b121a264816b1b680f754b787de7
zbed657d41fa52847f672017b18905c95dd3207c6f40e5958c019cb14f8ba3128a0346aeeabd2fe
z7fda8d3a745f9c76417aa68563e4550e331eadb7bb8c6f792fd6724a1b74bdfe6877aa6694505f
z10877386681efe3a07ac02a5e581262f44ab6330beb95f1b210c241a2ee9b7ef044f31fa325d3b
z8424e6a61377e744eb67f0f357ab21f302cc5e3f435c8fdba5965b82a3c051277e91471fd7a809
zc3d391ea2b140ed69de4799a54fe65e0c8017d2fd870b9b02ebaa547c6d73a2c7d77542b5d1c9d
zfe113b269509ec3a0a8d8d81d3f180fcbdb17bad98db9e0e9c230125a66d95a9e44ed295993661
z6c6b100b73a1c7728bf02e63d83e3307f8ad5d1116a84a80456eab9d7d8e9c28cae22e8c1ce78c
z05ecfbfc66be5290d099494b9d248ce5548ee6b01fad1f9ff998eb3669546725a6c654c200bf8f
z3852cf894e9ebd1e080df2370ffcfb9e9bb3f45f441047327c5a47cd9f3d1b5549bb93b35e17bd
zaa08e6e97b6dd4c15839d4fe1d1266f806ebc0b1d87ec5458c646fe626f03cd0e7cf5ae851788f
z6d3a772a4faab20979a47883a67b602ca9b2a071c6e829ee289fab84e182adcaaa0356c3aa3516
z39f2bc9f83e18aec49a788705370d334ff01aa276fd940b5cab85c72a4197b0ec150c36345e532
z906f564b7dd4560c499b1f68c57c1721cf162b76ca98d248931f17e68ce587f4b37c8f56da844a
z536df7db60da5c1fb3af0b2ec5db5440c6b414f458f7abafd831d2f719f86259142ab70ffa344d
z0cff2a0bd4725c5732e4a3e61b9e11eb7b088057a18580bd687cce238fb0d61bac377f2e1aef0c
zf4a44ec33986f97c78723c80ea8188a1e230ff57b6fb171bec330b0453b90702436537a17edbe1
ze0ec0eea6a3e935f24ae0c8afe5a5e68ceac3a3d1fb18c52d05727193e16c075d635c4c8218cea
zce3fc0d5669c05abdd219e519c94d74c54896f5aaa5e8e78e8aa35015144db6529a9550bf55825
zbd41fd8964e4f04f84d1ea8aaac17d05ef5ff701c37920dceb7451ed7cc9853bb2a31aa8801e80
ze96caed2bfa1c02f5e92f3d2f1fefe18436fb650919528bb93ebd90707cc11714a86be8ceda74c
z96e75d74c555590f94814b08a3099b2c9dcd6a8db0cc4573850261ae705db388bfcc917e33d91a
z46f4649609c2aa22f9b5c0791e3566dd327d5b99fa8de39bffff95d80d9dc4fd8127ba55d35837
z2d1e74bb818eadbd5369414feb69be7c638fe5d9f205ecb2a092b37e5b51eb5c4427ee7599ddd5
zfea2717b578a0a2a42bad5f8f77b60f328e31b07e43e726d74e1463b2ca00b7f7a2be3a63a552b
z3ba1ddc6039308957723ab8cba879f351d05c1566168444095479f29f42e9ca4906a974d5a6bc8
ze17cc7f5c8483dcea18ce7f6bf49a032f5f153f5abafc8fdbae783a1791c00dbacb6f650ccace5
z192ae3d0d7e1829f06b7b546861103ec9da4a17d62593813db7bb8406942993f21ed959dfd122a
zdd74a1622e731c2ac447f90243982fc3b0909ff9aacc9522e1fb44254ea679a64d574641ec3d79
z12ea09896683cdd34b5c38e894361308170a33ea0f114ba083d33199b46847726a528a7bf6365a
z9e5cb9429aef7a5ad932cebcb2af9f10ca4cfb9ee3768190bd3340acd5e46eced5fb3f5fbbdc98
z414c590ee528bd88500d38a1fbc37602c1c6e7237993abfa4bc15deae944d9ce58af5e0d372c27
z72045df8f880acb65cc48e84de1c425638ed5f3ab46079516040af2aacf5ba32663034b3a1b09e
zc31b75c2e89b3340da9507b06fc680c27ef75f42bd803677bd0fac50de48622226ca9f512b32ca
z122656c6c5de2683f08a4c2cbc5d1526ffe46f267e7425fcbdf24ab51de657ee32d992dff536d2
z402244873ec384654b5d5f89fc7816eb25cf3b8fb8f61aa55a58e24a1fa24b55470125914ffb0b
z3083550d26813c871d93185fe9aaaaaefb0b99201b72e5602318f1cab7b07c21dea767ce78d934
zb385bc3b4322294a53e63b7fb23a1e2ec9cb0d9fcaae40c78d06afa7193b1052e628fa1bc8dfb8
zdd1831697b474d6afcc97fdd326eae7607a779604bd60fd60587a78672404b1d4588cea0ebb4ad
z195d514badc8f5a522095bd2a7560f581d7cf9f49a3437fee39ba26994911f226c7428867c28d7
zcc4b72e332f8d0cb13685edfb0ce491e6a7054b560413f6e30c897da59ce47dd0f577e52a4a3bf
zcafb8417010faa800ce2b2db8e24cd1636c7a7213301c94b545868bdd4e88259888ca768dc4712
z495fd5e162617b72328f252b602e221d234126e1a68b3ab67f9da688ae21f93d3df231ea6db0ad
z53026dd59d5c114489c775931d3452efe86344802337059ccf558448ac467e02fbc1227ded1ad7
z8e8e42a6bd1a7cdafb4b627cfd6f4946fc46a57ddb32adf56779a06e77002dd28aaefaf134e213
z10c108a2a2fc6402ecef2a09f2bfd293b26a7012e8ef1c7927989eb455777ab12fecc72bef6b00
zd2874e7568fa8cb7364f9ce4446fd088b00c9f9768ea601ee116f7d47215f2a7273f6d9958352b
zfae55224ec4108f36ace05fd364b5683d6ec38565e4abba096f736638e522c3a0aff46edecc68d
z1aeb20794774a6fef275de857c244a671ec1421ccce8ca79d3ab9cf4609d924cf41c5709c97be3
z04cfa96d87afffb88b4a064e8211e4d16ce186688a2a87f5939302f8b5bb592ed6833c7da1428f
z97d93cd89f473de162036b142dedd6a0a7f0985a34fdd8f04f2e3a46ab4b6a1716822b89735072
z880915b318b36298936d82688ce45f724810f86508fdf70754cc0fe1a1f4d01a794b16828ec2fa
zcb9f64bcce844c0cd693afa510981ca7e18c668097c878aaa6e3c14bea361ffa46dea665d15997
z24e46308f05b49b7a1efb75e07768eba0a38d9ff9ff62f507e3272ac76563a78f62a1ca0821171
z5f9f28b9ff88dbd964f0023d4d64d0022689935f63a6d97f5736eab1a1926cabeb315595a1b664
z71a6eea01fb6f1e6beacbb50f67c800d7d38f5dc749457a216201c02b745d8410d712813fa3410
z2fa9d50342d2dd284e2be981b307291827bce19fbb35c23181f9b03ca61b852af6f10883624d4f
zff6def7a128b01c03a99ce02c11c3b2b6e922411a87477ba2a49b567303505e05323d9aabf545c
z6799d1f1046c28c6e3a07ed7a119df4aaf830ee50fd6d909f5a1a9fc3fb6abe85ac99491c897dc
zcf99bf7b895e9035cdbe185c59d74af118bc43158cf2c81b84c3aaa686b2965588a87db7a94048
zb13fa18ea10322fbbb36833e4adf0345ff5c17e5ea1cd5c9dcb607de5c807a9827dd71c92fcbe4
z9b48aa2b29ec59f8d77fc1cd1c0255dcfce04a11d55420edf99c2e4e44f5f4880ccf0c284db7bf
z00aa60ad8f68fdac86fede375b7438710a7f519b2e79a7a56f566827c229dc8c5667b4b7d6e615
z50ec0a6a8b5e8699bb71001b63c37ada9fb2b2cd3c38a3013de4107fdc2991918bca1ef5bc4591
z1eddd2076c69d0e4407795b62ed20ca38f655a1c73da6095ce3d3662ecc07633e9fbf2bf047c18
z774ea45fc74aa8db83b4147c6d71f88ef807d716546ae94627c885f5864eb8cb4eeeeaf27a51ca
z5c43f436c4bdcc7a7d729dff0bd3200e4006948dbd8d0e0d592fb69a052db1d48b62a31bca5e70
zeabb35d7dae83519fb6278046ba643772f517d78cb4c091faf00b4225c1858575c49888b844bef
z31bc3c0c188ce2d5b533e404cd31a94f7296dccd609ca027744abbdbe1fb342527971c309faed3
zba97b22c78d3c895858dd22ae7b9314c3faf0d263f2bda923c74d220572c9c1c83425560acfdd6
z8d72f310b5623418055e013513f85cbd19be058fd31693516cd3fd9babc8810851b15dff68d6ed
z7cebef53aed9697abcf0749abb7de98ccdbc8dfa8389742948c92894b212e569ebcffcc9d9dce4
zd786c16bce1810ec864062ab09f5c9d235a287afcc06fed2b887dc78f5e033b29617a7d13ca36a
z9c6a58bb7604d3e6c9364aea20b2414c8cbbe238a103df3afa2005a0fe08771872b65cb1776ee0
zce79e52a955e8b2c32f789276029a1f3a9a70b91a2830f29b19d9eac36bcc53fbd4251c1b75cd3
zafc1ae8141640657fee5b87638dc5198259c48e2fc485a5d415cf514d88d547e52f27fe31b7825
za3f836feb578311b93e9a10cdf9a59472722ebe835a8ddf13c98cbb2e3337b3c88316127b58d0a
z7b20ffc8c5243a31b9fb35cc0db3aadd731e7439d2664f13ad4e3df59bebdc0a9491b7f7a21121
z6da921959e2699859eaca95a64223495c972dfd692d03e203479df411bf187db5eb4335a8e9571
z460a56c3b0763c2d76dc268a19724a8c7bdd09b0c9abca6597a9b49b91f3fd906b08e130d1a87f
z05370743994143f87435f63ca91a0bffd423bcfa46271ffae4a75a96949c19ce0f586bd7a2712c
z9b1af063c016756dffbee14f68e917b49cb7573ea456884a02acc85e8982df542971e213e23608
z7aaf4e5d448441dd6e964133df7c9d494f661111ae51ee327b76df10b4e2eb8af3dfc2cefc82f1
zbc0562ef8f8b8ff3db3427c5454b419abc583e750b7a1e082bff10a755e8dabd2258329310012e
z898ebedf01892991624547ed871d86a52969467332271b555d70d5e4ca51f016e5d1723ad663d0
z0b04fb9455dfdb5f0f82e35dce5bf01ade14d00dbe43f7b7583fc695b5bb7647acc72bc5dc1f18
z441711453d5fb3fe9e3839b5d1be1a9d4096abf906ec18aefdc0eebe1c787c3f95bd6703a0db15
z027df5890c15c48ab431e4c2e20f99b9d960ecbe1fb27294187eb97da29b6a4a7ded9a53168bb7
z9796cf52e902f9f4245e69806296263f976a7ee60ad7c4f94b644251839d05d0faff3b80a3788e
zaeed529c9ecd2b42c605fb6e34a650a2138a3507b1bdf3fa7f2553710c33832e0bf9bed9dc5eea
z7718b20d64452becc9bfcfc5939786ba81a7b59f0a7a8225df0657ca2c1bc3c233bb9b5d941511
zf35690c3cdf334e2c1342562b462a314810b63387e6c9bf9f99297ea9b6953b9ab7d58a1a7a42d
zdedc8b61c635050f16830b7bbe1fb4bd92b8b140c0fe38a7fb158b09943746a6c3b40113729617
za3bf4df4c9fd5b5e86a6bf2ba910cd3a3ea841b51baa6708319edb76d3e6e3db83914011f203e1
z952515356ced973460c57f81da6352787896f1a84a0680ad6780c35a43a65a1327e5e6c081f101
zf4eb4cc9655cf45532b4b2118b582c7b1005fe6b8d58829e7d8af8d28d9fc1549d3681c6bbef23
z6f35e0d87a55dba500c1d916ac193fa7ae2e2aab03cc2dcdcf89cad8acdfc8fb1d68a0ff81b0a5
zb6c059ff44a0be728958ea29829768251aa46c50d1146d3f939f923649131046d9b84f15c73da1
z5a2350885c60cca571e2c124f69aad90bd281f938b215e7dbc7f479c4c9e8bca08305710c93b72
z35337289cb230b6c200dddcb7c8336564cfeefbc872fa1b6c9e641b0874280f93ff080a1c76324
zc562fcbac800e1994ce14dde7cf5d4f834fd5cb7126e9a07ecbc36468516aa488dd9ba439df14c
zc0088bc3d2937ea69a49b0d1a3752183bd7169d33b7f45384a03a7ff10c3c1f8738b7c8ae908dd
ze7602f0b2011633d6a45595b6bbfc4c698e8b1b4a93c8255559020d1ed57a630f2a091f4350d28
zc4bb1f1e2ffe0cfa671ff9f82ad448eb2ccedcf3ce80efc01cb855e501441c172093119990dd09
zf9d041cdcf99edfc6033c61357813023fd48d3825ab9f669bcbb109630eb54cc8503179515df67
z3d2fcd39c8b18619fcb586779e406e04f55515fae837b46f7188cc38f8a1209b75fd88d20fedb5
z6e1c16baccd324aa4672735fa915b403657cff64f54b11558078a2ee982923749a86f973696c14
z09c7e4a9681f9497d7e89d3d604c4081866a5027f50b9ccbcb5795c813faad2474e3ec770a1c91
ze2c1e47948cd535e5cedaaa3a92081f458f41f90950d5587cc839f826430501e664cf1410807b9
z2dfe643830b8bfdb478fb3eb787c6cd65640b1848086f149505670d4ab10b756c663556149fb0d
zb4ea6faa09837784131e30ad4afc3d3e2de776a10d8802aaa751bbd9d5c4e565868182dffab2eb
z3655fed2da2c429b2d46019519340eecd81ee136cd92c6e352c2f75052ab34af10162094abb308
z25d3fe87a69b9cae62d673ea25856684cfdaaaebfef93158a0a4fc5f63fbcc52b06bab7a5dc744
zc3373031fbf9c339e3987a1eda52e004c97b5032051b0c69dda0fb6d54e6c54945e108c0d2c846
z7ee1b71b5a2a7f7d25ffefc2c01f3511595929dbcee6a9fc100795127f2b68c633a46f745705f5
z2724abfa61a6d67579dda8d0d4567e57b65a563ae1d4fe6b37e0d1c9b34c4783be64e7e9337057
z67c4dbf317fd2bea39fd4ada6087e8a35787e024e10b7c8877800eec54a449ff0cf1b16aa10bb9
z07647e891ae6191fffaa89efe3a8ddd085948c97043f140bf111026a7125f02033aeff2845c19a
z21861d9b277d5ef04d213a32e61fb94ba97ae75d9e676122be0367ede30c447365a4a79a9431c7
z8f7d2bceccac533e4f891e81949720b39e398ce8816347a33cb15eea72e0192707b3139c499f88
ze605cd41bb959932b3538ff68193fe0412281ac7ba07684833f95388feb6e51ea37b85ff5b696e
z04f70d5f2279fe4d75a65f06d482b734cb6dd5a939f1be0c1175cb4f3901b5569e306b6b3d38b4
za5dd0ddad95a704175b48a474f9d2485583436c957a72f2da7d85e3ca33587a2da3c37da4615ec
zb0640f7a74884b117269eeee9c06ab726b03f58a9d1d688c98272738764038729c6048ca5f601c
z29960df60f11f4a8642b3d6e92feb3d1934b2c356180bc65ac817b7ee5644385566900eb7dc7de
z7aa34b2b06aa94741135f4c0b2f52839ba16a10108f8c4038979a155585223c67f34a8947cfdbf
z3aa470df5abbc872fdf11d708d5da52b2c4ec665c108f1cad00df66fd26f89d9401b4e85e79553
z7addc04905adf804e583ceae8d106dacbb5fc82ac75ba671161766ec9dfd502e4b90f88d69c66c
z57befabbed6f315946d3f0d8e61c79d0204f3ed97e6297544f2e371ad150783ddd19098ecd51dd
z4d3ecaaddc020f6fc45030e02a200d8d86d30b9211b073266b64060a7afc0e3644e5141521e769
zbf45957f3eb4f9ce7e999f8a490bd6f2c4de4e50827fa194a20bcfb72d6124ea95adbb6c2e4833
ze096cef989657f757aead9661541157d732cbb2ce2cfc91e8fa9e7acfcee7bc3bba329ee67b944
zeb8e57e359621551503b999276f6d11e7d816c07d2abd50153fc865ac24c05a926fb6073f99d42
zae9dba9a138c5098600a47397229c18f9bc655886a34e46d3b1ad0b80ea6994096a9f434fd32ff
zf12b0a30b4aaeb83623b27e7b19dab7fdf0772456b79ecf0547aa032225790419a9d59efe847eb
z2c80ea1ae51d717845627ba6924db7bf1b533f3074bc14368381229ff01ceb5908f459f42a01e2
z4524891e2eb9d3196d5fa3fa855919cfb9ef8981268401606f3fb69ee61c9cbe0c3358f0d7432b
ze944be407e604baf966d0012003a069795948b7daef93c708ca3cb2ec1a966b1993818099caf70
zb45d11b26ea466d0495d45748539859af049b82c680618094f97e41471cf05a25fdc62cbb7d1ac
z4d781799accc303180921e6034ab03f5cbb97bcd0b9d773d1e63dda304e54b751e5ed699c9826f
z06691007225864f0bd2b2b046fd3ee2cdbab09ecdad520de91a8a4e9bc5e9dc7189a24998504b1
z39652b126aefdcce40e5827cd90233b7d6f124904986620af1434b266fb58ec7a99f1c07a5a17c
z4ddeedd5e2cfc7a5c2a33886d6ff5c7def7addaf4a76dcbdf88c1c63b655d4616e8a327b5d76cb
z0f0f894be8d103d16fcd47eea37c6527dcdeddf741ca573787d235fa8e63805fc14d3abdf34f07
zb79ac074b8ee66c9a4e81e36e49292b505270e6d15de85a4705cb95d1b3d0c049e4e5f2cd86f68
zc66f1b6712baa81919464c64b0ae899573f6308bb2ec5419953e4fec7f539d249ec409dff9db82
za9cb8927574b878f3f7f59c3b670e92911edf2661c754c186849b756f536a07fb871d23754d54a
zb980f9dd90e9424e1fa0d1c0efab03b3170941db12c4ca7410ba46cf2c7ee37bf9fb6c700b6212
z13c83884bcf918062a4b230d7836695fce63de8600d1d1445715bddf6ae1bf22cf1a92d5d976c3
za6157235d6e2fb014075882440f643ce3f66b425cb4711fa5f6b677fa2e2ea67edde1f8a86d4a1
z69ca5b90a3917e6754880f330f4ccf4437c02435222d2bf251ee7e4b307dd072a90f85167de68c
zc0dc39608763da062409f35b2b0cff0c3f325f60ab8e013a464796ec641bef0fab1caed4537da5
z3d287b3eb826548f7a66edb9afc9c8f8aad5d23985f58e538e0377735a9559c2eade5ceb604bea
z4ea8a3ae4f80bb40ecd4224bc1b1e44b047e499e4211ad073179a0910f893694a4f0f60202cbe0
z86a9323eb472508184efe69143647d5e224359b09ebaa737c6165ae9e4cd6a0adee2970e0a3134
za560e6555656a1aa9e3ad94926966921a9cc83d94c637fd0fe81ededb2b3553a5586e6afb7cbc0
zdf556d726c73ba4aee01d6c7494a75e5ee364ba08322fd09386644f264c05ff2e7bb45e79bf0bd
z5ef07d6dfb19a553537b96a56b656177ba04f67676a1de093a8fcf26fcdd8afca084482cec0a5f
z2783776647c47b9bc27f9c4387750237c31b58cf798f583a35b0181265b0ed4b4d5b541865aee6
z0f8809452dd1f209967028b4ef8e8431f0cb486bdd2aa30f32475a57ee07d56da567f841732fef
z29074c459a6f42e42cef3c5208d2a450e227528094f4ac7d38124783142741d64cc22e5b51e4ad
za446599cd0ce45c6cdbe5a1ea38183d265db6385c54c9975aa394f2cc986989f9cb2d08c980233
z1b26c972f7ff42795f2faaa9ca909dc78db2777c947a3e7a4c8b32ba1eb2aaad91bf693b06ca57
z23cc562e8728b2e35469d314db9943aeade560af4a3ca47d302b6ce66f88a23ef361bf23ee1caf
z16c589cc77564aae4a26c0bf0881e1a33bda6a63fa8247b03ea6bd49c85f4dd46b3fc52c321b2b
z745389086278a8bfa8e0520c97f7502cc2520e97f37cfb17bab9404fb028f0cb151548896b4feb
z38fcebb1dfdea5f381dca2a86399bc6d93a7c0839507a453cc834870e3fe1c294f1367faafbff5
z3f429bdef0e954afb2dfbb4cc22a2ca64d694221be870cd8d4c9d63441875de26ab9dc535578fd
z4c6e7101962c674d8c34ab05e8d3847f03cfe7d15a27722ae47e8a6141ab8aaaa4eecd12c4bba4
zf54318ea7e15c3e02d445e8f7d90474ce44a685a7c80e53e664e65cab0acad31721d9a1c20672b
zb6e53359e716d759c2a50045bbe389cb3aa15e272dcc00983171b42ffc055ff421a56b741134d5
z5804b6bf101276225fe8d318369a6987389f5dd0d1841187e3c5b339c5ecfebb6d4b5530f815b4
zfd3b4208d898e4ee1a6e49bd0456cdbc9961451ffa733cf609134367b492fb98a363ba0c4299a1
zeaaaba3b9e900c42e83892ff440fb3bf61eb1d8902f776ffcc7d7227f8f6109ec335ed358e1658
z21c124c6ec7dfd82b3a6ea6f35c818016debb54129cde27683d561703164c3755e21defe1bbd53
z12a1cdd73001c9e26cfdeda53f324eb1950125cbbb845bcd7813193eb96cd4437fb9fc2e4c1964
z8a2b0d5cd57f431221d77f0e00d6b9de47cee7da94bba3853fe4185abfe339d572ef57e85cdb93
zb531cbbde98264f339b224512743676063bdc897f0c28fcea671a8677c5e608c3258a841dfe45f
zaccd2f235063e53d11e0e3dd6c09ac7efa8039828797b0744ea42e5eb6eaedd64ba29da9835d7d
z8c08cb5a9876031aeff4e520563ecf26af0760666e3cdab89d4622460bac08ca86dfdde78f5650
z0c09f527bbbc0d3b9fb81f3dee3b84711d60a8375364d5c0402fc4d949aa5ac75a3dd63f717318
z7eac5be5b26691bd07b7c4cbd20f59105af4920984f94cac148be945fd22b1711d66b0c41500e2
z83f5a356f7da457529e3b77fb1b9cc0e03fbd0dc281e664ac86663a2151fd1cf1ac59d5cf5f391
zab35f713a0bf800672eddc876990e0e465f1d6aff7390a919e5644ad56fb0890d6fa7b1daf9344
z8b975da208c28442df29d394d737d4fba7530c8410529e0895ff955d68ed76d6a46eacf9515eba
z7c25a9bfabb50d1bea8bf8d934efee8499919aa00d2b9f59cc07d39d4e3533904006a1dc6bbcf0
zd7783f8b4c3b22b5db56f36a112c3d12664c707b14b461bb5c85ce35b05d1da8d25edcd2447c03
z0c24fcb25f9aaac1bb3d5b547b12baa0c09dddbf4d8f6426c7181adcf2126c4494f82d128819a0
z6c24f77da69d4cad32a243df0f677042a40d057b71ac9e9e5bda6676b5a16916610d35d5357710
z58d6f74736b46a106c6185991588b74d076b6cc70f9b860f8dc6b32d59f9822ee269d120a6daa4
zcd6b96775350a581018c7b4cba39c735745be3779cf9ee9fbe74a046bba9e725e02881e387cfac
z4492669a3c6531075b4d72470073d3645553874b320bfd49ac52a9172aaa9cd0727709dd49bcdc
za34ca0839519be47d15aab9f9e40105d348c7fbd38117cdc52f2c1708be87fe109690a11583476
z68248b28f27aba920f3ca5b9966ca36505c1e1b194a1c1d1a0fc1d6c9c2b8b426c676c3c7eafaf
zf766caf723d7138cffcecb6726d7bca468d256735d8c194b53669a0ed79adbea107d779c6c010d
z3b53b1b4f05597d68a883633e9c06e141fda8e2207f9baea4f3f3f88220fd144627a721afe0e0c
z259a9102ece73659fcf3f116e78836999e7cb2cb8b52612e21b9c579e905a94c2812068102c582
z7729e071e1cd5ee6fc92cbb8a54d84112b08430178b74d6f65b4458bf598a19e840b15da689448
z120f9799e5102818d477193d30883e5c9a236c20659273809857c68d361c7065b9611309368317
zecddd1a7fc8e6b73410883927a766847b1ed56e010d0dbcc49dc1062812987ea6303d84c272011
z8060013c895e098ca10440b34a9e5180e7c2c74934e89f3c391738b05bd5089cf516d023a26921
z557190ebb42d1d48b16e41c2ed5db7bc9c9aca7826f95886c8777ce872b4e759258f697e864866
z226ee0d3d2fb30b4a8f541894677e89867c3c7f16dfe3b8baf3e826bdf375161ad1734ca4f96af
z3fd3441fb90fc50198c59ac46ce2184dd1c7473460cabd5a89348d1e76cb66afd9aec3e46b54d4
zfc5eb8df6d654a6e0042c4574e259c0f7e62455c42516efb755ca23ed73218ee778f21c4986b48
zd2651dce3ea7cde64416fd2f7ff0fb53e070b1520d8efed47f1c6e8136d584030bda5d093b7ba1
z6b2bb7c6d4944ecccf1a6c1847f615b45c5aafcdd42dac9e1ad8d8813003bce42c2c6e6881fe90
z4592be9b22a64fd18c554efe0f842db5e5d29e400c70fd1edd1f541acbe7f5b6ab1f95de8205db
z871440f48e7e1dab40f74f2442819b6d3d26eac5acbca038f9f7fceb353d5b32378077ffd13455
z27059fe6f877648b194b166f4c33d7febb779d95d1a9fa73e94c125f69b20372002b23dcbc2b1b
zbd42306dba8763226a1f19e35c52078992ce2f26bd03119548e5e2382624ead49215275690b0cb
zc30ab7568f5f72301f7c186d94e8a4cd7e8b4e1ace875cd8f5bf5f341a3dc3b758b8f585e111a5
z48f3f3e030262bbd71f09fd713f0c59ac6c6a61203dc99acfac514cdd27b988658b9b1d43af10f
zda172352922df5105586a9c2609df8516994f1c84e143ba9f4e2b4dc84cf3f3f8b27cf7e563745
ze7ce404cd16a0069a98ac363c00851e034a25e9716b264387c36930ca31f2ef38796b7b01d08b2
zc725cc15d0f974935efbd16caae1395b4384f86f8377a065f34502189749e9d2c4bbd2420f52e9
z4052204eb3122fec7685074c47f81732d8226cdf4b77ccd4ddfd0392f3a6ac162b124d694cae60
zf20eb788393b5356d0fcb89b66466e9d03a9ace9473372c9aa2bc874949550a491e340b41cef1b
z82234bea4e19d253e7fccbabafd90f30d21557688539cd95711f8fbec2a8843f348400b5b8a248
z530d7025651f950419ca2e50e3c11966cba4c0f13b16d6dcc1cceaf1326c11b09ca5ae4b926df0
z9a0e1557d7ae871b2f95f2b6c858f3aa6ef7162668e35b3c21edba5d59a1cc6e52b7e37b36f6dc
zaaf13957c7751c4ae53905c67cf2e8bfb31d65e8083792a7eb13d4bd07a295a8f363651bcd71cb
za2ccba0e31af5b9194c34be83323fd2737f64f0e2491d092a43dec1a572c80fdd5e4055f103e9d
z3992e573467481335f98de5ad079a44c63680cfd0ffddeba904905581b3faa55ec19a30a6a34ec
zaa19c5ffa29683fb8168a59561cfcd58f2aa3e75b87cdc64ca8d3ef9305676e45720b64f35f2b4
z871a1c3098dde074267cd69b2635fbc370e7ca11e7c262324e7e666949285dfdcac7b8718eaab9
z756517b1aa6d767f3e36c7b54adfa49bfc93b017b77c1891ea70e89ee808e94d4b184196e8bd5d
z21c726d4c20c20e829eac0587e8393810fe4554b6760d8de7b306d79ab1d396f166698ced38160
z6625af57f8bff0611e44cb1c5e395ad11e5437f0041939fd25797cf02b141cc3043f7d0b03de89
z825a8c80198b363da70dee842a38755a1d6073801179d65716e2190449bc5c33c797f01fe2f768
zfae47cf4ed980e44203d42226e3cc8cf4fc66087b765b6ee9567b69c1431a37a0f94dffd2067b8
z31a76cd3fb8746827673dd5ec2f0e36b8797d4f7784e835dd5dabccf1d564e33d9590c728337c5
z5d88cfdbf5c2303c04bed4361c213a9b0133367114764edcd756ba737d8e56cc2a9e33df3a3a12
zd84504bc9ecf7700ca8785041d195305966dde0578d8f6e42d737b48f0686bccac90b24fecf178
zb81629819d65ebddb0a63587ea8a84a77f43b739dfec1f5d4be16e1ac5248ca79d39f2c1f6494a
z11bcd91462b434792db76adf0d9e0c074a8b1bd99b296eedbfcc7d7dcf55799728fd550dfe288f
z0c3cea0b6b70f7e3350d67abef620f8db38b442b94b718e13243997138cf4bcfe252776a4f2f7a
z0e5e7190a210e7284d664e403d1fadd8b049f35a610d1d56c26eae32093b649166606df4717cb2
z0b5619688c05ed8aca5c5f328a3b458053801f0e92fd352635f62e9d8f7a9614a81f2152269c56
zf40a82ebefadd2cfa4424098a41fc2aedd909815d4e4d5e45619fd88a009ce641929b1e0fe8841
z5dd125edc992d068afa0e6a2060afe00c6b4eef738c0c613bc71a4a82d18075e8c46be178c878c
zaf928d28702c601b02fd449df60588127ef4069cc2430665088b842632ad840e3b7bfee3047f23
z27aefbc303f689658f8130299f3f44007145aff5b7628581d4fa4bea336b3392df1b85d4ca7916
z5f49dfb74b93b6835ab79306e38fb775a774fe7ec00b92c2c119fda1969702897a8fbd0666505c
z2449f049c37dd23ce0c88c884355d0c79fbba202bbed6c833784615f2a59e01a03708500016891
z269b14840189445f545c5ad5489140b500c2f4f20eb238df3b3b5d29639ea2476daaf20be77e12
z6cd4c14ac6f6b9b731b3d270d8879ce5f0a466107ddf410445548e7fd0bd9f930ab8d38aa49318
z4004c6749d5a7c074017afdc055d1bf4f9ad860623b5aba68c998a66ff31d93c10e8bd0db9d106
z7e3810e7bc867eed6bc151823b19f3d4f5a7c23f48affe639f0bc733225d615af8d13498c3ea34
z15d4810240ebc69cf2d26f86a9bba271a67ad6e80ee927552fd940b4cbedb8f438d0715456fa1b
z4d85b271a640a9fa02db025bfe552f8bd60d40677e625bd1ae99078cdd6d6566229db50dde7a32
z8e9a2c8ebfe39589ba3513707e4ce4b05df814e1dce1bcb0058e93ff5c1704f711bd7931e8b066
zc807e32b5a027cb7e60f6cf6b478961ffeda3d995ae34c36ab1a8695f597fb10a6d877e8fb3959
z41746bd4daabddd67628a8548fe52c8c9eec3d416a9398e8a02e00e2cf1f98eea2a45937277f9f
zdc5cb4110cdef5aad0631f1c3640426c9fc04d8175b39e4ff4531378abee8f8ce64add8e9bf099
z7f2b0c9983a6a36a355b0acb38c9e0d69ce0d978e26fa7a61faa99ab5fe537a6dd6687876b3279
z95e51b66977f12c8c0295f6951bfdbe8be3ba547d646c557a139e0a6ded78aae9f481afa57a541
zf5c9b31aab57601e2d4957a108f566bf62ed084584c652de32906341d12b3d6f94e4f905f5cfc8
z9990ecd1277f9a1034b3a2147617c0d0054b42aabf32f7333463913d6b0aaeb6d104b65d9ac470
zdb599492d32ab8609309a3eafd58ca7a39e03f91277ba99017dfa1489609085856376c24a9dd57
z4e095088cb2ba6c027c640d70b898a487b95bc18eb7b076a542e2aa51eee6a282cfabe2def872c
z6e72dde27cbcca0e29844bf60adb8aa6d7eeea50a32367d015429090b576c5f2491e6443972b16
z5f2cc248bf6da09c85cab7dc26834a647acd0dc48fa0f248a9266fa2fbaa840cca7546aaeb98fe
z12ebef310091c42d6367915dbd65fbd4f41b3b5c9862e1001a522508d2874dd3e42b5ad07827ef
z4a3ebfc85a780d5d842b9e1fb0a8421cf2d5779bbca04426b12257ed9664e4f07f68b01fb810ab
z1b9ef8d38640d48de0790be0562083995413c7bfe82e79265b6c6d2335e13ca7a52391378985de
z630c550c06139856bba006c2a5b56157312e3317ad29e2c208b19a90f27088e030583daec0e0a2
z0a3db626bd77b3da3bf4416cb46a0c8221247b0d5a186184a38ae323b0884886d9501916e05965
z6ef4a32aecb8dd069c26b6656affe86f01390da9addbeecf39cbf7c3bde2f0a34dc7062d82fe9e
zf65fe6d9c1b633b3241d75aa999376faf019bf189f808fe3e5444639413f53ccf648155895a137
za3650a50df47bbffebec979e56e1991b612cc761749087c0fb1cdeca581b3611d004a86c4cb9c2
zc635582ab821038f0c34e06543f1129e0fd031d28125f432c084856cc6f2e8e7fbbfbd9dcdd832
z804291436a6cfc70af00d71cb805dc9de98df9affc2438981d181b06d03cab66a6fdc13a0ea75e
z5a88f528690f7097b8bdc40b47db247e54493f34898fa5b7357ebf696a7d2248ce783cecc92165
z344b3f4fd74b13481404b6e13d7df63bcc29134eec0c51730187dc1c7474bce0ae417840e5b80c
z86a0c861ce3de38d930d3c848741243d624007d4711fe544a2c4a8fe87e7c56d112b6915b0a170
zd3b25611b21d53744b3f7c1dd34dc3ed6e06eb8ffa1bc0f239f315143d424b91a651e55c30ee36
zd7bdd11f23c21ab796c8a519afb4dcb55cf9da425a84228b0874950b12dd7697c8d8439429d3d2
z69e56866fd892eec1e01876d713d69b95606cd8a401fd5d2d16bf60505fecec4727597de398cbe
z8362efc2697339311d230d239638b2e9088c0c32ac56b281a7a4c54c72ba837dc5acc76782f9d5
z2341e48ff66318456bde44e70e4d37ab13a0e5711e5436d5adc382da6c29b2e4acf95ddc1e507e
z8deb09701b8f009067965d7427585625ae3c105b3d7ce27a924af8a1a14a8a25458ffdf52fb006
zaa5594e728635587f59c199032fe2edaa1f441c1b2aced5625754007c6e91f868b588296c46dbb
z697234cde50cb04110676ddd19fac16ff7b9d356228e49c6237e6f6e192403e9b8640b2504ea96
z3e39807feb8a2db287d0c5bc7ec9bdb4cd9e5115b8dfe6c458b0fe36e5203867eda8f148ed82c3
z049143ad9675619fcf1368a9a10c2e07dfd960593d023830d2262750c1634fb975d235015b35a2
zd00865464c5b6722621a9447e94cd0627562d8d3d06e03a7f485ffca2c0e9f372f298ba7680e0e
z1b911221cc1ab3772411f87609bf918abdeae5b8c711fb14e515f6c26c91fde91f56524a69a43b
z8c6f68bc2d80fc48c46705a698b2214aa767259788d217728f0065f1671bdd90e0ba2b907629bb
zcca0bd775a8f7dfd47b5bc216df69b9bfbf4be230f73f7aa27be9b85f14ea3fdfb9b3d9862a3cb
za8ec926211cfc056148a4b52d3f1d454fba6921b4e1b61a58683d08528584f5101b65f0f60ca02
zdf7e9e2efb38d29ba16268986e02104abee4e0105d436acd43631442197dac6c66f75aac2057d8
zd3bfd881e3ea15bbc8c2924942689591d63fe973e911c604cf6baa229cf41eed4a5e832198c191
z0b89768029efadcc3d3ea5a62675650729227e9ab4ab4d685be07da8c07d644db3a62e3f513d0d
zc07ce217d72f5518afa95a0fb44ba2fdb4fb267aa6c612c4c0f4062b2b52773f4929ee854491e8
z18a61c34a3b50a8d2fa6a911e28d7c56c01333903266b382ca2bc27f3236b0cdf014800c230ebc
zc9c8a463da4d97a450c9e0d4aca77b30bcdaeb861c2998326d56467b396d48b492326865dfa0f7
zdbaf0b8e60dbd68376a077f5504c52ac8c9a6e4b1177fc23faf51c3e6cedb2e89475d4a7bb03f6
zb7770fe7dbba945633a897995a1810c58da97c2102d68fdf9643b2455f9d498e2317826ff8f833
z59f92f220ad861d675c54e4fc8813e81038b16cf420a0a2b0a7903249ca33209e262bcc374415b
ze61bc2f99decf06a3ae0eb555215aed6e2d685c0f6133b17cc46d54fc018db9f321f47bd0d9f82
z24e982ca4259cc8fee8549fedbd3f372c147c07fb896cf672ea80a6b89a00f686af7114d8ab5e8
z9f44e9983c384eef2b8938d33734ab2383c86944c3168a89fac74707f8682a12b35a65d4c247c8
z219c3d4c6c07383ed9bf44bb104af2844aeda5611dae57e44cec63157fc01d3cfae5ec01bddd98
z01bef6b31787caba960a5597b49cd6174359e3e55aaae5a014cfc4f47198909cd4436792729f41
z9744b494483cc29f5ce89177df0f31a2508b849c9fe80d5fcc534667fa9950b18b2ac2fa6778e9
z1e16f21706f08ddd03822776903f6045d432266dc36eb9d3a1e6a3674f6f076f1b3137f4cbb26a
z95158fc2645ad9df96e5f3077101b061b33aff858cb086fae017912d977896030e52234eb505a8
zbad7381501eb22a8c299ca450226be6182b0978819df35228da4b76437625369e6b951931a43ea
z2022e9a1072ce3d7607a4f87ece39e1045159f6ccedbb4a90511150d77faf6d5608d1b497fd93b
zf18b96878e67920c41078eaf97745766beb5ef26a5a3cc074030b73fa3eabce3f0968d93fdad65
z2ebd3096059e6f951ad4afe84e6f92a76d38d6b76bb71075d314e5ec89b265dbc7b86638696310
zee853bef47c1c22741a0196a6e3bb773170e130bfb280ea20d03f16c82152231886d884a487200
z1bccde79c9ddc00aa102820f0a3d78d6c5e293676adf39a4f291d2ccbe3c80845022d3de479110
z8cf738bb8b9ccf7765e7075107d4e56d7522da48fcd819ea762e69b719d24a5c0a27abde5764ae
z9b2e709dfc0653cbd3ab3def3902e71b56f4c0197057d557eb4fe86734009f714885f46f8d14d3
z1bcb2d034ee88e4f9128ba88b6b15cab1e2a6182a2a42861353a276bb13ac2d6fb764774ffaccc
zad93571c606d32c731c81b9a6d84107756759eea06ec9b280e2b79ffbe4e8ae5e39600a7b62f56
z46f8aeec42a7303b3f854f1c3ba88d085568f78ce5355744f222e12958bfc9878b2fbfcf17a72d
zd2bdf1ae0c17cafecdd732593ac505c5a6031f05a661de7e7392d8f13e668bb1e3fe9d9b298026
z38c7754a76920e3c58ab5fa7c594dd040dbeef3b6c40dade032849c43681397062ac3c267eba5c
zc19848196501b97277c41dd86ab9ce0fbbfefba784bb87149325b6663d2aa4715892b78fd0291f
z2006ff24101290075e2703d1f37d37341e5dc691cf26dd6a01821fb7e5697bb0dec8ef6daac686
z573cae1cd0c3b7c9f19c65645573df19bf300eccead6cfd67622dc1a2f89e703b9d3cbf2d59eeb
z07591f3a6e2f5633208d8f303aad9cb640e8513f56fbab0f68b956da234f2cb8e7808e0dbd2baa
z3df8343fb97a4d211bba7fe64376a0c5582adb094b6746a21983cdbbffd5370a7e8d97d25c5253
z1d8b015b375215c8b7538f211002b9d3619b75443533efeddce5e9d332cb4bd4a447dc166f1330
za7fb96cf48f4db8f0a545e9d3d2588ef8570d7bce1f1364fbea6d483e8a3acacb6dc71ce1d8f43
zaae08d46199a0b3af9b04c1b83d0d63480941ed35de84a089eb66243ac4fce75b95051089165b9
zc8a39f3789f4ba7412365d462cec13b461b4aa8d3857daa555aae0af5b86c173766c5ea038a6da
zd8dfea35aa8dd1b9aec2f501a429d7e36fa96031c2ea93fe265fede6db005b126c134b93dbe452
za6f1580e76455a8661ff10f499879af3d19b543ab8a8a10a702cc0b3c6574c3f1e6405d90c0db0
zc530e43356e323b9490626a14b682cadb00f8abd3a66ec77cc9cf2f2339d3582b98a88b5c9e979
z1d3375a4a328bd6256e96b19df2d5dd774ef56205a3ed99cdd29991111f7b2b04f86fe5fb828bb
zb58b209055f64933b4471141cf5b4e9fd7b0f63334537d6ee5745d388a4bc0bf2f6c0440e29ba8
zd57d091967b70c8d427a1568482aba3233c7560d755a4554835623cafcceaf725e6d2af294af1d
z3502e092f30a11ba79c527cbb86d7c64c560fe3b006788f163bfe123756444fcda04c18a8b0b11
zf2b45ad6695f9007e170daf429cca0b678f5c272a684780e5bdbdcbbfe3b77d42ac1a44bada6ea
z983049804487351883b35640494825e444b02e126f57143d6c6b4914acd25b0c0175d523b45f06
z018e9c3aff6dd65af282c164589699a6c6e2400a4c29c32d3b9181028597892d22ec38a6f6e39a
z7a472914edfd2233ae4bdbbebbd66493ec98896afbcc1cf9c1fb740a560f4d947123b305835c8d
z1e34066f10b14d3a0ef0968fd6e088586880c922270fbbd21c412888ba30f75782b35d398800e5
z401810a8bc516460dffec11055711ddcbe27dda376ca0f6fa8a05bf1c24b700a807bb548e827a3
za7249eb4c49d6ad89bc67a7dc00723fe7c6806c353bc0b1df216ff428d6f4f64a0ad35d5685483
z80ce35163ca35ebfda5c4e605d4cd042dbf0283cabc14ade5ea8abd2b1b3944ba09339beaa1d07
zf891dfee0b4ccd169319475221729a8a9c7758a909d4a329f571e4f0568ac74e35a74bba11f876
z9fad5dfc431e2a86103f9f601b9a3cb9ec4180213923bd640cd127b6d541427f8d9f07bfca5063
z79bbfd48cecba785275cecaffed14014d861fc38dcf8acfdf527bd0dad82b690295e3f4ae718f9
z102fccacede4e79a274a9bfcdf714f0daf4a11f77d600ac63bf1646b61bf8146d3dbb7d87df479
z2ce10dd0846957a8eab1d3307b51389503cf2e9a36f1bad2af010f2c244b70c2809aa120ddc443
ze78d9ef9ea302fd6aa8f102339280a93cab3b123a8bfd338c2771f4f4daaa177d7ab5687952387
za61a90514e022d6bd05f9f4e56270f618d2ce5ae79b8147558910a81f7f262024480cbaf4b3777
z0e5ee869667102d21426141fea452e8e91ed9e0bfd1bb9ff6c24c8f204e0d84b7a848a60dfcf48
z3fb6881e0fe205733554b03226ba62758b2fa06556ce0bcd98625f85f63c7bc65b2ec1dbbcbe19
z9cbd5421d6611398397b58d87268ccebf56181e8219581b828ae7141709971520e18af89bc84a4
z2d9e7721abf346e28dab5d326db1871bd87e2756311ee5cd1583598a5decbbc8583c6d21ebc44d
z4ddba76a146a08f022ee138ef73186d509f6777822c4b475d12992c771abd868a8942bee6c3365
zd59123a25d8d987f4155c0d306bb58f7940a375abb319e8f4ca16a44ba7838cea97324bec788c7
z818a53086a73acc4fe1ed22fdd9c44ed7ea393b44b0fd5189506f2ba7a88abaa5000e21df32ed0
z7562e87fa407534741e20e9161d25b31291fb2d88c593ba6c29f991e3aa7c8c2ae3820fb3932b0
za77e9d92ef587b2d58196dc7fee0c1e88ce7be215e72dcbc659667e240bb0af315959d8e4a9840
ze2a551aee9ad3e68d65bd54e0c6ef1fc57d19333590633252ea897f264baddfc305b81e79e2f49
za664e97189686c184e6952c9df8c90699655ad932eff6b2b593a0b0b4c52dfcdabbfd7214e1d5a
zbea66ac57247a97080a08101c125ac595c745e7f5e0878b4543d63b6e5b2404f8bce65d8eb0d8a
z271f555f0e2796ae6fcfd0d914b5d245d75e3f1a2287169d898737f11a5aca7fc40b775900d04a
zef5862ea781d3dba57fae6d743a827d9e692d0e3ab8b656a499a60736d3c87914fc1fe78390ab4
zb8814d40c970ac93d3385f4350a9f9d3bdb1595619efa27673e234ef2e1b1fa40d184cb1feb13f
zc03857977d28e825c4e4af0a4a2cb9dbfac86c3d3f44943929f23c9965232992118a8c1508b70a
z233211dc95c523b5b6b449e1832c5119dcf29a745db4adbb809fd80f2193c9c23186be03a23435
z58392e7ffb4cef91d968f325560e17cc9cf1dad831952db654381a37879c030d986f7a7ed86e79
z2d0254ddc2a1b26971c3468eb735980a3788300be95a5d4b59ec445c9efcc995480656719d4099
z361d1e78a3362db4495d6d44d636552be0f514af4791f69c6e9d37ee5957d797129dcad6ed6712
z67cb0bcd51183ba7cf838bb08a6f7cd24be69bed972c3b1abd1177e1e54e5a1bea554a72fb1930
zb53fcfb757ac29358a22b3e55497ca442c29cfd6b4e1bf1896c26a858cb863a3d7ea7c1017b0b4
z94f5a4cf11cbd97807a8cc95145f6c9497dd98a154f5dbeaf0131c5b0427a167272597c0bdf4b2
zc1d97a2364eb7e0165bafa49879591e2c6e8aa07263ea7a263de8c86a6b11fee9f9379b1217861
z1fa4dc8db39347ae59bc58b0412d8db253a2c422d78c9668bca33c211827916607dfa44e10b529
zcda59ad357051e5561a2086fb755fa7ffb492a4ae2502f253161f21cb101f6dc92d6f8d9d57196
z07c4a91b95cb8fc676608c3636ee518188c035bd599a99628c3d71d7f2ae4a072ac4eac1a8ab12
z81d31fc2141464cc79637002aedb3339baeba4bab15984e65b2fa46ee58969f2d1558e1c101111
zf35a6e386448c8449ae5bc7f777ea7c19b6e50bb86ca8bdd18aaddad4f77b6a0a35934cbdf7d4e
z2bdd2d7b22e818722c87d7c0cf5e4c9ab2c5a7a1726fcc6d7d9e1bd0cbadabdc863403dbb09b79
z76eaf6957ab27f543383d7017c54700e83df78597c7c2ba773bdd56bb23f196f816da658f2241f
z413f190756ba0de6ff5cea359b62fc2d4039e6d82cad509ea9d1c50060730d509fbe9ee6320724
zea353188ff1a13d3b3a9d2e1b1c74d5b716f6544544cdcb8a38b7071a993385718265f40b6c5a7
z6f79886abba47fc396d147bba3f44ac2ef5e8d122bb5e9e99c14f6d7381860f8be0f2c99871a92
zfb2cad800997a522f194502a372f44accbe696a0fecef9c02b58f327c18b985ac612647911ae35
z4274b1b62deea23da7958107aeb1e3349057c0e7deb441b90757d279b2b5ec580f41c0c05294e3
zc0ae07c671db35db333cf21655a042ebe7e37da58a5a21302081ea384ec554c5b1d733fb91e883
z292c8f52fe266171ad8d11c4f9c26ecac1ced51c8de532206183aa37223755e9f1d9c308810cba
z4614c3eaf90b30ae78123228e49fdbadcbce496ba0daffa01482720b051bd21c604f283c11e603
z25549700b788eab81e7243a946d63f95defe9c60b06b0322fb15c9edaf1b87bc3362e5ba113dfb
zd605500c8f7f3797d19afda7791e5f3a5a8b1d0d0aceebe16f6c404413b974a56472a4abcc7ebe
zd0aa4660a5f967105d98889962b072da3a431d1b9c5009cc1d57facb4cef6f8950764c154c7f1a
z2b09ba20baa3e7887cb533996a3e9dc3980b114bc20af4062beb876271cfe5a184882d87d57631
zf05d0a26b5b06da1eff8ed7db5dde2a296d48e2dae43364e1f27a1c6341286dbce62e9a535992e
z3c5ab2b6b7792aec8bc2f479501180046f6031b197ae42a386dfad306639aad1677be4920ed906
z2506a873d2b9fe8a86c3d8afdc306bd8dbf5c661622fbaf72596f7886b68d72d68893256b528ba
z415b25e4acb035dc29b441466e9510cd7f79f3e5cefe9732856aeca4f032543473b57672781b16
za88b4d383da387a8deda46d2541cb1ed94b86c6fc580e43256d510afdc3412a83b0ef42fe2c5f1
ze702500681f3cab3a89d11a627a7c1d397bb7e2d4a5bcf80f665e95afaf72cc8c931a65239653f
z2be04c41a9f8d703702a2032a20c5308e70a84201675af26e85294b933ead7806b004302fbc4ed
z88f55e17f0e38537912c95dc2435531609380cfdd306e87f5d595ae8d3be961f6ffd943a5b1e76
zb7e6d3f378b6978a8cd390263ea4b92a1fb55e46cac3f1565a5721861e6d799a3563ca3b581caa
zf7a9295c67ef8d1b4727691d4d352c9ce774e87cdfbd6e5d0cd0f15ecb323d2e87c4366e544e4a
za12f768f201301a8614ae90428925206b9492ffe073309a6a46f238a6329ab380c67ad388eed0a
z58fa9b233aba334bc1f2a15803e54799ff7b4b8fef980acb5efe72fefdb0db87dac60f775097d4
z8fb716bd74c1c553c4acf3e1ed256140a6d3e0d931df397137ca3775a456cb7d847df20528b177
z51f4787cfe5f60d51aff2e0cbbea8b72d545d9ac6d2a1e14ca2b2408a971f0f3e2e48efc1e63ce
zbc6a074b2aee94f5a68b42ef1560622187247c151f6f51c0f190cb5166a2e099a1f64043c0e3cf
zc7889a0c7f58e46919f3060e4e41526275026d4960baff46c0f0134529b20cf97fac227fa208e4
z5cc71d5ead34d16f096399e67102ec7ff8a3933fa5c045fc423dcf85527118109c85148929474a
zae6d7bfa5a8778256c8eeabf2df6b92d3673fbb067d727392ecde7131eb0daa4c855af49e55368
z8ee814970628383bf3170725374263d290bc74b554e3c8806c1ec0a437df2696bc5cc75db063f7
z58655d9b1b3e8f56c3c51f1a0c052a9f02a4a3340c4e371811f84ccf5b60d859ae7904c6c70fb7
z90079f21f3d1dc4974a9a4343e9e5f55873695d07cdbbf85638737febbaddf087f96328602daae
z5405b50c5779b187a4c26211885a1527735888405550706842b2fde296eb80ea7a41df33e7868d
z0ce2a23f31ba9347d5f5756203d86b4ff3bf48e0aab553e79a4d4cbd725acda56fc5e9f8c21762
z9333ba48d967c0ff81b49719cfa1289aa6e84aab898cc14f8a168be949ce8324ab38232d95d2cf
z011c1c521ae93a6bacf9518a4b61ef4fa636f00139ae3c19aba15aaff6f0f6c8a84da88891d4fd
z9f30230db16a54e08988493aa0007408bd9a92af452aa8d3b2b787e503d39075090b987d672d60
ze3185122a5ca67b7e438d38cc1d8082c1298807c48c6925a6301620373a5387f5a2a8867601dc8
z02c9da497558c22e13c90601c230c09c05d78200265d63742f8b0f84760ea4a4c3f3f6bf99208b
zcd25729692f47af294d7f97ff94946b4bda6f06ff360804b7b39e43f86a4d93b00ab70affd1f3e
z644bf1d91e6c2dca381e01a45efc4c0fd48f9c170e434be5bde3bae781f1524f1d616ce0b92247
zf725ff670129f80147e2f94129090a83440dead9b903f27636e53ceb3596655724d46a7b13cc76
z964ce7cd99fbb0f28ee9ad1f22c9764d1933932923382c99c6ca1821b91dff73a0134c2857db25
z043edf967ffc97a1736dbdd28b4f4541ce04ad0d08ab8ddcf9d0b7895c0d4e7404c16235f7c6e8
z8b7b139b484e41d9c62c8d96526a56a549f56bd98b2deb73e2913f43e3728d81b5595200413eb8
z696133d04a937c0d1b912a2a03bd55a458ceda5d2bfb4a131242b38e90069df746201a7437505a
zcab6e3b1bc241356191243ee2ee7926a40f3270f16f00064269ae8dc54357ea04df66d96771690
z1ac660c943057db52f4eba1861b3053db5a91f274ebdea5f09e5b8d0308fb37fb4cf6e31739e5b
zb136bb01303400d462afce61c0933b35b71179c30ebc3a2cc93902620012a50e36b6637952a085
z9e5dc5e53e542314e9c45070c6ae2d9c1a868e700c96e78430807f19c08f08195e98859f1f45e2
zd089d3588c4d2b516a4d1eb676f4a739faa192cd5c57fe1e5db75131381bde8df15eb2fa5020c7
z695d2166efeec9b9c5225cf3bc9d77499d3af33c8e2d21336ede2ec3e78d9ace047d6b702fe032
zdff21251da0c0f0a87478a43888bf86951954ac687021ea5789f03b16aa3bdfa4d1c63cd48cb86
zfc6f9e0b056332bd9ea74b187add2a19022a45fd52bf2c17f3d72fd1d98825e9ee49edaf36f6bb
z78ce2eab6972400c4ca1ae05c9ca60ebd45e827ab291c72abc7a982e64e1437395970ffd230e9f
zcd6f6371f8beb5d708de83d16011cdcd15cbf937ea776d68beb23c234236e489ff807ba54e8cf0
ze287ab57c8dac2e0095f16bc1909a5f9770abcfd884ff58284159bfc24060d148a8e9218644f73
z6c34d72f80f670779277a8ca1e654b66ddfb5df9aa9d45519d25e502098b02bcd53d831029d023
z54d9efde8829b11ce7fb6b19822a81c69e1474f613c3a601e54c993ab4e891085ea9df7c2a65da
z6a8a6d8dc9f7cf5b6ebe5ff52af699908c04ce71c4db6b7d340c841ef717ca83448779afdafbf3
z1eaa892b63b6a7e9bae77c40348de2660d34e5ea9307537eb3ec9287c7d46905be534a2d516942
z30c6c9232902d0a634e06273991d9fd6348e9499af6916f3403f98d07c8b3fa47df097b9d79035
zd986a4e67c2d53c81708778f56d44740828889ca93c0f4821d2f30ee4feacf72ecd63f527be49e
za339699db6b53975e4d4ab250c19c5c5273fed5ba4c93fc60de17a1b6dd79f2fc7b1e018cb11af
z1e8cc6d9d0be432f13644cf418f11c3225868ee114efb48daa2870f238faab15faf4c4e9023e9c
ze6527e2df91360c2feaa6552e83963335128460bf28d32d87cf64d28bda850ad2ef8408f201e1f
z937b8e2d02723567d963b5ea6c6870874c484bf4118da2710c7602bf9aeabb47156efcd0926130
zdce335652ffcd135a3b90b3f4124228471cac3d975f24696e4334ba72e4e056d78167c671671c6
zb0dbd4982ec3ecdbb144bff8a2de8de94a1b17fb30187c6e8d8a66f087086d669fae710bf0d8bb
zd15240f5bb871cc6cc456d324373e0e5e18a9e81cf72752f8f892c5b82ef4a7b84892177c8a55e
z5f1748e0cea62909ed0449e49aa46d455bbdc475ea98413cca2d7c34c5ceb2cc1c5cd278e95467
zf6deea0b10802fdca7c89b1cb22741ad205fd1ed69d79a0b6e68dd50e7b0de71996ce87dfd1433
z3dea046c03f8a62888c7d7ee0dd74d6e9a622bd71a6bc9a15a12b526661d5131f6d1eb941dae19
z6c91983d3655fd423cb039c78b887784c9e6e2329c3711da2cad059ed2194685c1e3b779e700c5
z2142eaab2a2245e32ba12323c1132d1ecf48c52714f2e549716147429a1b55fe29922e1cbf41b6
z7350c97fade7b38396739e656bc6ccb50b2ba64de7484a4e20cb7d673dd3b5b6a0f7e6facf6ec0
z9dadb66c37012b2e33fdf18028d6d7beb49fce7405eaef1dc6ad71e9b78fcfd2c641171b27133b
z45c8d449bd023b319a6ccdf19afdcc4b5108890dbeb1836500dfc7592517f0efd3eb4ac8573d7e
z4765b8422a72f4e323620dac01a176e26f9094704190de9d84ba33b3d19cad5c74eb2d0556d4e2
z677ea498a75094d7f3c790a6088aa01dfa83c46972cf93707b2eeab81b4da58eff3998d9b24ef5
z6ab8de142bed2218ad4e822b5a45fa62af8dcc7349f900edacc5d576efabf82f5369a89334a236
zef1cf7147309ade811f7d9ac64f345bbef9238af11f12ba62e8f171564ae1e058803ea923c0d0c
z79e644d909d6d9b74b2c6c541c487fdbac966bbd051274d1e0ec2e3bc0e17939e17252135abe17
z64b68c2bb10964a8c665b7891df49c4b6949b3ed09cdfd1c2de4f446f957faa3326c987d1cfa19
z0822c6f0dbd50173b4dc2c5453b542981d76744b48b7dbed1357f7e63b542aa7e3b6b8770b0153
zadfeb8c37fe058802dbe1453e788f2aeea0e0520975650e403359181a2b9d912c6c422e67f1021
z6447c0dd14c494bf61c4bf763e3b7e08d7349a4cc42315eaa6235789bd0fff57ca90ec966cfc00
z2ef4b105ae6e5b400303817130f32f8f39461ad9b32dd7c3acfb2637d1710854d5dbb4e0517284
zf440deef46d29c4a20db82e90896f24b08bef94736c2e50eb56a0526b198ec77782854f38c4f93
z0899b27c8793cd4b162ae881f69441045db8932381a26596e413390384ece50ce1e58f59521440
z6d62085212aa0784448292a5df38b4bdee38743556096118d9ae3afb5b98c335cd7e145f353c82
zd4fd6d335db6b9b1afa484c21d7ebccef5a36a6117e4b8c26604bedf60e33b5ee5c5345447f1df
z61ee3c5fa44b510cda483cba77603d74cf5c9f9f75056d27e16606d41fa3d3499fd4363a2155a8
z2a48841abafcb7c41a2d7f10878ffe5c544da216ed409d29a9bd97e184385ce47a02abbaf1acbe
za7684959e350278cf0253d4f94f2ba608b6198d12c30d01bf1aee2d7ca8d364a2bea41774b2ac3
za52c131c4f31e7cb71e11217c618095d00295b845c0353391ba826563c0bbb638a9d5f4a6646de
zdabccd9eb65d327e75c8e0046d5c40379205a645b04eed1e8d0dcacfba8c968ae64fdd7238bba5
ze7fad1c715164216418746ac2361ad9ce22bf7ffacaefa6deb062df4ba7534614204ad0900e5c8
z9861f7bb8b3b921d181d4ed9b15c7267e857b0679051c72a8ad0df2a5efd77ffd013af437cc029
z969e15eaa6094e631aa945bc87a8d98a9731d312e430399cb969aa93acfd26dce237cbca29e407
z7f8b2a45babbf65c8854f11f9336f603ccbab7dca433228dfbe3278153fe992a69f1fa505b7033
zea2027b73dbb1aa9ee8f979790685dd99a2dc1ed9b7271ec6f5792ec7000f26c629e4bec00fa97
ze59070d10547831b3d2e6f65e24160a5912e797a00c61cfac30a4546236e30eaccd226ec4dc428
z43d8b01b008ef0ab1ffc3da8c8238e20bc1039501d158876033544fa5358b4a10eec77896a0b7d
z15ce2cf1582f569e92c72ac3100c3cfacd3ad04318c77120f2e25e54508379f13af00abdad0f6e
ze2bbe6f27e9c815b5b597d8f451e2057892792d3e5de6f94752a9bd5c9c2fef5540dc7df8f84e9
zb03671671510fe0f39adeeec2250c51e2e8833c0f7b4e6b0e0072223753bc7e18bb68bc72bd7aa
zc134e972166d1e5f68bddf52af93244ef1c828b31e671bea598ed8c89a0eb7eadb5965fdd55a2c
zff7bbbf47888768aea4e09f7d4b82a0fe2a8d550abc0ec93fda6d5714fbb29e55cde541f9418a1
z2c90e4a72beefd0c1cd9935ae75e082a0db53fb051c2abf2b9421d17b768eafc5f92137abca333
zce3a2cd43da9c9c618bf253d5ea3510df2860270530412b7a3cdb9388501db6e9bbdb38747e149
z9e2c67c178d64b24062d977c589e8a19aa2b721fb207f013af71f633a3b9de8a54bdbdabf9a508
z46618ce3fb598b5eddb558139bcbaf138f900158f25b7f9f33b65a92d550c20e71c974fc81a5a5
zbf74510f398c25adb1031912851ca1e24652a7eec44ffacb0943553a2659697c04835d8cb4620d
za1379d1c8f2b4e5fcd23cd1f28e0499c907e23fea6cb69abc5c446563ab5a767070175c7041d40
zee5b935b7397b79d40a95c53ae43ab76381f5e9b94c6b35f184075908256f1182b33998d407435
z5281a45bde9be5444ef21ab8b821acb4d52d0608430c546f121157b3fce977678b9be5f1bc10e7
z19d615d15b2baf92efb53803abc9c1430ed0c29597eb9bcb98a4adad18551502b4a8b71aa6daac
z8853226deb56a46f0d461c14965af290ac52c33dd129efaf2a9f71991b1d568c8137a32bb1d389
z55a5db64606bf5c5239666d072dfbb650065a98b0d15177fb8fd89c1f7e10104054fc2d72807f8
z9cb6796379cba39dd4ea650ef8bca8fa5565f120a3b7ab2c8339aab9c8d9f492651df8572d69db
z31eaeebdf5af0bcd89c6b91fa0fd0777e65551bf610e7d6b44501ecabbe1d641ca79b780127d4e
z8d939b2013e1a7999f8921026d799af9dcc713f59d3857ed39b2004f5addc8e0c35b9ed55d8bde
zc05df89cc74b3f2be65a105a43b541c93de49b34c242bd304c9cab25ccbfe8d07b8384f4a10864
z7bef11ccea973ad4470aec9f977c48db81439bc90205c7fc63c323c27fc0fca500711299e79c3d
zb436d36ebc491c5ef2ffa168a052fd5c560c0d05ed94518e72df9ba3157714d772e3a95dcc0a12
z51d5676e0640aca58e44842440f0c8973d3c5b7c662a244a1a034a608d6723a82fecc46acec9d6
z8b6ee7e7a2c788e53f56141c2f9a2f37f6794cede4ed142d3d413ef33b55a05219a45227cb719f
z021a5ff8c775f9ccb7f2872d1e1d333ec29d5658cda3bd8899693c33a8d3b422116fea528b6ebe
z0f488d85f26517d2e07863ce1e990781bc489dff55eda94a0789e15bd7c33a7e029417ffb064bf
za636562621b0b86bb003fa785d2e73318057a7c1653c14976fc521711dfb6089218b947d0f2a7e
z06410e3561d3a111d7ec867e0a247aa5b648f7e4d2edfa0e625155bb40d835bef211df0c79ee38
z0ea43e1d592f4e4a3aab5567ab5d222cf6456752b352ede30bf50edf92d04cfc72ce0a5107ddfa
z8bbb852607a31b0b83474eb9418a1bca7a3c637797984c7892a7669e7acbbddc2d0e7e2c29a799
zb5b7a2cf9c1b5fc5c853b98ecb3a3b3d375d2a8808b92d58a469792a321c7974d6eeba7edcead8
z82a203702098ac9b05540a0a7b99952454b895d647ba59c88445b5b7127fb05fdb84b89095f57d
z721a482658ba3105b2021a32f0dded59aa6281db7001f591cb739e16ae73a774b4ece5fd6ea82f
zb8ae79440d003987aaa575ed4f9e86b9bc6decfea0cf975c073e5f4c0cbcf974f8083eb61005d3
z3b66e0636dadd53234e5e629c66b5720d2a445a9fe154cdbc416e2b17d2f6214c0cf9e4a8d0108
zb55473c1d323a2b665be63b732cdb305e191f9e5c1d76fac369080a55def949ebfbdca32fc619a
zdd12c8291b498b5fc687fa56f27edac77a2c8f1de5b6ed35fcb6664caf2318cccebeaddd2feba2
z46ade7c17ed52afcc4b24fcadfdfc2680febd68bbf4c7e5a31177055f53278bc8005fb841f38e5
z5f9a1bfbbf19b8077059ceedb425649e7e1ff85b79e5849cce1e666373609e16a5e9d2a10011c9
z6334df9a06af270ee33553de6830d0d37e46a7219a555ca0fc5194d28701eab30eddc400862684
z6171f8264960a0f794f1f79306071b87fe7059ceb28736f6904bb5c72a428b96710c6ccc20cc79
z747276149df6b7dc547fd249929f700605d60883e4b71fb59e7e4e0fa0e3cc30c0e148f3e64bb1
z412f28b5949a24bda21a2ef1edac73c8ca40dda0fd730c3e822640ae9595e47186ab3ecdd6bba2
z5a31db84880585a44cd6e78a3b9bdeedb06edd6e35e4703bc8c3186c1d17f161f3d884afb2124b
z69adf8822ad9920549f291f72e9d41a726649a770c1f48d0a939001d62adb74d1e11bd62328e90
z5c4713bafae54cd9be97e398a0aca94b2a68a638cab7d0103fa5dd62b43a7d79bf51a2197d1e57
z9d292c42cf976afb7535e214f671d39386d94e20f54fce0b59f6a66a72ad4d991a1777329530ac
zbb7d0d40fb6f7b01c13c6324bb5b0881d053a91582ee999d198fcba5e8c466606e50d457594d51
z41de9d3919f90ff7706641888605db9abbd00409863c212dac5942410dde73b4537f8e2bcc5b9b
z343797ff62ccabf79e783748aca1c030c3fc1b8c1ecd1e711b36ed07b666971c1712c68e8447c4
zd6d63a2f77cc9efdecd6ecda1241ee2c937f73f7f1eeb1ab7b2da808ddc9e3dd1eaac27f92e5a8
zaf540b33d327821f00451e5021e1edd43ac903a6eccbd45515bcede6f5cf3e1a4c50f40d2190ca
zd85534e664572ebb16fef76ba64ddd2ae4eac5183d1b593a16680996a776ec5959bc42178bb47a
z3334174c4c26730de71e88711e00d664898d9c8a17a1c7e999e00864795f82f760f8bc4497e36d
z299fec65ff935343ab039b1fe5b61da4ad8b24c8f7a6030d2ec9b161ea43c18e3d67fe5670d3f6
zfed097337466d6f8c111142ccf738f40571576b5a2945eeb9d3861090b91646f98d98136ffe08b
z351c83ba3242d96ca5de84a139a91020235bb0559c7ae7d094f1d8428d994f75bf2551fdab9dc3
zbf81e734074402cfb03ea965ae1f360712def9c49678eace1e882e3c4cb67ff307a289aa2719b0
zefdea00537114f49982c819b6779b21468761e7748148ed5b86624cf81c27465f1bfeb34c333db
z0c6c4da6aa3e7e0a0af00941cbd35dcd4c93f1901804ca5af1d4de2a5075f6931155291b129289
z6eda8b82816cc73ccf088c42202c0a5ecf333855dd3c341295dc333e0761f4984ac5a6a02d85ea
z0cf5a7d1acfbe660fb3ab4ee339656773bae7f3f982811b32dd87e7b2df4f7e390f83cbe5c8564
z7b33ce3c66006883df29d63b95c175856f4c6bd6f0f62459403c9d06287b2a757ad54af2b3370d
z302a981408cd97b41069cdeb2718eb57d542687619ceed5c883dca2992ad56ee2d664fedcbc90d
zee1c6cd1fea9413f7355a24f7af155b001f6f9d6929e86b721935f94ccdf2945d172a52e8270fd
z5d06960e9738848b1f2c2a611ad7025d75949aa29cfca233d2b6d2d977697f4ab2dc8245eadb4c
z17a3cea943702cbe5879e883e967dff77cef858702a37862b9811eb64d59a801773066e6f65010
z937261f780a62d5cfba13ecf0a3c5ff8febf4f26752d4fab38ec0ef03b4ad93fad9e13f3a3692e
z4c7d4c45da38be603cbef7fa4ed8e6cbf467b71d0f928b92153360a34398f197543584c31483c5
z26610c2bd829a6d433fa0cca76c431ce52c9718d8ed5a1d0dba3756107bb7dbbf4dc0e2108ced6
z1b7353405af11419cf57180e4aca83886bdc5f024f449af56d9c82e093a724cfa2cae116b176ae
zb3cff53526e6c396fc6ec720a62a4e6e014c49cd0165e2ec44e7e646d830bc570dd9ab232b8d68
zbaaa284209b3645d6147826081b24d9196f41e6f877a42a5bf62911f53fae18b63825d3ad88e0b
z0efdea0e7167ed05e30cb2f8de66a8ae4ccca868595c2d52e61120e36f10bb747992df2c396bde
z84c24f1baceb8de631d40fc119dcb4a76c6c54391de5db035beee3faabcdf79cfd6ae09ece5040
z00f01d72e7aebcbb487b1628b5759892d1750ae81d9d4f8e897408f78f242ba7021e5001d14fc6
z9a3e2b7e565503d03883ce36f7a6e1fc7ce7661a9756d87be88c34b43e24e1d7d1a597e79d553b
zbeb833100ba9d4a89af3fc83db68ed5d4ce73ca1e76db76abc30d04fb5c1c338ba8c816e9f86f0
zde6d7b4ba8057f7707a7eedf0b12fe9ab458049950e40ae3833266dc8161b412a14da28ef09b5b
z72572f1a5dc232b2f1fe1de4e11e447ff357215eb4ec9272adec976ddcb2cc243c64db19bd834c
z84301b8b342538bd120fd0a604edae0f4880c067de6f94bacebe1f675fd512b90d61ffc342c9a3
z8966f349bc8cc345f0d4f823896573d1884b249a6184ad9c11867ab4a14734c24757a289cbbf80
z6a823b2b3fe802ff347237adf964cc1d4d61ca2947c5c45fba72d0c0c1349a22ca5a473b76e942
zd7b663d6b5834de3bf0676c81581956261782f85a24ac56f33ccb664580a04ea9fcdf77f8d91f6
z6371d3c80c191cca20ba5ad44402f7efca8fcec36d242136d38db4eaf4151b842f77b8ace94a88
z30eb238de4f85a41a5227c4605d0ef14ba5bd7407063786353b5ecd3a9ec8121e9a94d8db6120b
zaf35d0737f33c5c7b7087841d02945e4009c30a7d3d9d61318ed68d0f75f64cfe11e97ce4a6b0f
z971be361b512434c71c54fa12a87c1dfac9f7cba3aa1ab5042de12f5319918bde48bce63207b52
z3da579651103a2a58fb48c3613862e1e7fbebb9a374f60ed903487d719aa1f1a495bc91df1e354
zfec6babc20215a01f312a63a846553d541d083ffa977eafa79f43eb01c26aa8194516d7fc74d8b
z0fe7764b2c19701f40021d66afcbc20d70bb8b5ec4ffd42a7ce370e7fd9d29fcdb502e3b2367bb
z5b8520b2c37894f9d35861ea62d857ae33cd41f6ff781daf6e2293a99d1262043307f0e467c76e
z7608d343a814e4f9b18a79577e80d60ca603ba95b2086fd4a8e1291622e5f83c7d8fc2ff10db5f
z4b21849bca47da9a0603efc8d70d9d8ae518ed6f3f4b1fb8a59c9e761e5c2d02ae059b1dcd1ffd
z008976f206450a4c4145593834a5e81a371731b8878ae59b4e5f75b55391560a09f0e1dbdf84b7
z1517b9f2ae56735e155e777a5ddc279fa73c97ef2ef00076cfa85fc9c4dca0914ea9e25788d98a
z0303a2a1e39049d9c48a5ec6d5c83a635fd17b2e2410cac68deaf31901d7ba5bec01f00e2bbb5b
z9cda909a5b38954e15d15542e5412ca4ca49fd1b73af8b758f3386794ecca5c1ffc4b49a19ad55
z3a859bd6e258e0916679c0e5a1bdf58bf36fcf547b0e2d7feb33ae2cdb5e5582193f7de6a77506
zcbd503da85819296a7f4f57cd828ede785756b5beba1753fff6333a91980538ed3e2af44604433
ze76f33e3e2641a5046ed563a0c9bf38031aa4964fbc75fbf2c22785b5b83cddc5fa619faf38192
z56c756e22a5c6e5bfa85e1dd2f554304a9c5f4c77ea520b1756fe83cd5c20537853aaddfc80419
zea2ade3965ac8e4ebf7e6e42995e5877accdd046b7a42b561fbb5f8576067947950914de3ccd76
z67e2be7e01440e3f9584441d900314e1f36ad22dad48c85fa9f276cdc2078376fd08e4de933bc1
zd18df5343a93eae7823fc21c3e197fbdde0bf3557a87434dbdc6c2045a2514e79622dcffa52239
z3a0093ebca79ebb99d21546a4e03bbf680800de6cd2c2a3574fb98af3cc608ed0747d8e794dd22
z2361d720aa818e990945e0fb33a29e22e0e20b06e6689eaa6fac294053141fe907dfdc2e7852da
z362237d5c3dc359afa7c1e766edb370e0a04a20b1be3e2ec1a8f6cac52be61da7133ef7f0106ac
z7adc7957f5381ccf846ad4fff4f01da208435235a274b510ceb84acbc640a3a26a6bebefe7849f
z24cecce8a37d74cc374d2dfe9e1a595dc6c70c73c6bc1ca96d768d2ebde2f7d61d283936a235aa
z1738cf04b4a14572f6bfebe08554651236922291de995b88d98e7024240b69272e1226f99782b5
z05465654c05397583e193c4cae4daf5470673a88be315f85debed474fbd84bdd8a6049f6f58952
z693aeea9fea73eb3b68de4cec1a36bdf2e8f727f7cd92ea783740438e986803227ed000afe1e5d
z06b9fa0c808865b172d83387bfc3391151cd995ae7897c5af472e01005c20bc57bc3e6ac3af0d8
zd17136fcbbcba2a39310180acbe3f731ead46809d56315612e076058caa570987786b8d13b75ec
ze9fb9054aa92778ecf164420ee94aef5c327feff1278b74a8407068c0d404acbdca4d820e6ba5b
z34bdd29a159cb4e8d80d11b69fe5c69f993b78cd65765295af19faa2e33be2097d7c0c600744af
zb2f5a0a4cfc112211381f3c81c7f310e0bf524cc81108e901ea7babe6c859401e1ecaca2a03a4a
ze338713264400bed04ae1184b1801c54a06818d6f4a52040786155e3d446770acea05f6dbcb144
z2d4df996a4f4ce1bbb17eb180069d2af06f114c44beb05a8a38d56dcae78a7bcd0cefa630d045a
za530faf90e631ec7ab01413c2c130b3feda048c08cdc9a7e79d3a38331221059f6392b9e183d49
z445cd415137a26e4491fd95657f40428515d08936e43cb1897533de65a544097c1b69388d6dc9a
zb854f16ec63327a49a889b90d603fecbcbcf4b9bdbbf5c22482e373e58e4e63b5bf87e52c812ac
z152685d131c8b0deb9fddd80f6e85a7aeefc71ea82588137eb1ca405477e6f44f3ec694970b694
z25dfccbf3ab321d9359461b025d6815a609863de4bb10e9d0a0c503b8d1c32d7fc59fefcac5195
z9309e592ea5c1ff54f4b37d33e72464d0225ef3779d3c8a75335f08e4e93d5e199f68f9de32c35
z53e4668ff1857a6eeeb71bdf572695b71b84d61a8bf6f071d31a24bdc1650027572fd87f77ad55
z655c347a94b5e0fdd85a5f3048c317d7af37186ca9b3db76b94c1ff383ecf09e99e7da2f83573f
z3fe97fc090796c1641d8a11c4cb289683779e5413a7511a56e9e4d7fbfe00c01baec126373d532
zd388bbdf6b903481c5ac16fa741d2ef91dea462b2cf299794e1ff8002268793a90835a5ce41393
z9170d5affb313480f7f2eebb1fabecea531b8f8e6e02a54a358eb320977ab0caa710a5598aac4a
z4b50652bcef984a14d8ef71c570c58050cc26fb38d7fac40d2813ed3b065fa9b7044c36177830d
zbaa617eab53074bd62c1c1ccd56912e2e13ec3aadfaebb8694d35577e8a4180cee72a2ff43539b
z295d2387e253e9498e7960cdf0e094f150ef189c9b69f9b08373b704803d868b24b3657b006e72
z5d47b3ebe8f9bf375bd334f78a3d4977274529f4e09245edfb9ae633597ead886f109907e17140
zcb179cbbffecbb2ea1c482fd5466bcf2193ba43f8031e23e0bbb90e7f257c32c12f91e56b25b94
zfca30fb438ba82ef4481ee09cb1a68491facf818bfb8c3f83d8c2dd7fae934a361bb62046a3fe2
z46cdc218ffecc7e3591c9f4d87d6ecd8f2fbfb03268c084e5dfa8f833309b66601a99f4b3f845e
z98caca98be51ee03db3b8fd92d7350f3330b94f66849d990f69e54955d9949a8849faac26092cd
z66a0a0ff75d6915202b50647b6af4a58e58e9e35f348c6e37a20168bf22d4137d5547a42466f4d
z253e6262b79de017c33fb2833efb0170412a483a3afa7fdcfcf443b5d26f41acae511a10f91ff9
z05ae9b420c71890a5da650978ce4f1705d0f458bbbbde4275239d6cff276c7ad94d85281560511
z239fa031cdcef2fa2d23289a66110c151d47cfd0a861294461f441949999c7f7481c03cb9d51e1
z1b0e9e7cabbbe656783ec932d4f496c95494c261b4a61b64b45d40562758bc915753a14adfd2c7
z21ece6907e263387a504d53bb81518383e907c27d42c57a7b46a5c27c6d5024e66702378285cb8
zb26c7d73d0190a5d5123a0073dee820673ba89a76654c7e8720de9e1eeeb2ca48982579da85267
z7ad4f64e0b814b37c3c892d95c260d25f296b676ad487696128a3698679a8aec69d0fd4329649e
z6af3ba2e01fde78fcdf5b0ed50c0ad31fc3c8ad5a838112532eb11f55c09d1765b02ca1a990787
z6355d0951bd6a7981e14bb6e10542428710cea5fef23e1ccf4d7957faf0dfe836140bc2132a5f6
zd95755986d40cff84d776c8d1b570fa5fcac0c984b3d5bf18726da1bb0fb71aa4eccd2fdfb1212
ze1488a8e8a0f46605f055fcdc90227d0adb0037245fa23c4f76eaa19c876d07896e8d569c672a9
zc328b3bbe3cd059fd168f9b6eebefaa3bf60607e80fc3c598d2f1704c21773a54d17438f5a15c1
z7916cfb74f9c6e08efc3c6359e8762d8ffb40fbd1d5f5507d979f416634b7126ea19cac7251d1b
z49be74563c614a2c0d05933b2dcb28dd910701b9a8535e56ccb7dafa7075b70adeb1af05c14ca9
zd0f762a10ed0e1b4c56e2f472ea9dd0afa82221f0fd25e99b050f2c3d0451b95e8b1b5d7eda106
za09743d307f96da5788d34cb9dc07924c9afb466a45f92ff9b7d33cb19b6e932a2bce99369eb89
zbfbfad9144df5eec7a458a8a711492d548f2eff2b1ad68b6606e8e18daa62d6ccac87c1dab7cab
zf88d779d91adcec245afd0dd09fb697d56e0d3f3b05c3604659fb28d4ecaafc34096af050c1e15
zde47ecbc7ecb6bd670077520215ea64ee340c867d7e5c6537d392597bcb718d09d4af46dc7a6f0
z1ac9573f190b83404ad76d33ab6509369a46ba29cb3691ce8753c13dc60a057a849150ee54f4a9
zd9f2dea75b76cc61524474ae380719dbe72ddaaf2f6539e092afeb792ef8e43769a74c5a4999db
z5f27e5514a7b4abf3cbc75d45141c0ff23385b32047a60bedd018002a5d2e1a90e3711be9509cc
z509243e12bdd74bddaa82bf5af054d475dbb236eb14d576257546e0f3bfc2346fda469f65c7136
z42d368c5d1d0f6176bdaf5dd3bb26b9190b7b1ea4146aa98152002a84118d3879b693352ff1649
z32978be8a5daa541c5eac4d6bd0068215dfaa831e647862324ba233cde9e5906f2542355a2b834
z840d93a27f30bc8a38f23cf60210595ba85dde9f257e4d1cbe5c1282a3933a6eec901b79f4962f
z62c1171ca3cd9bded912b7bdccd1060517d5e250b3a86c2ddf418c20351216c5fa368e8b50783d
zf0cc5de0ba83ee452ceb80437887aa2c24ecab4d8b62e8e5184948c6c956881fa4d7846fe4149a
z9c7fbfd62315700860aefcfea53acb07261863c240e9e963faa5a0dd3046f4af86f35372d8ec3e
z1fa49490396cfe63292654f383f27d95d1964b3dd2afcb506f2362e83201981fc1fa6c5b39c664
z0e43184cc87dd19df835ae6f53b85994d3518a25a04a11f41e3cc86348579a1bc3ea4830050f09
zee66af46e3f95a26b2cd649878800204925a40e03ca260ec367e0d9788f4c1da9687667c76a21a
zbec599855422f11f9f1cde044acdc4ecdb2fc15b79d7a6b6af6305238c030b001b4eaeae4769ad
zbe3ac84306791971cc94231e21bcf7c91e4dd5bed501229a8cd966a5538d9c17a79a2ae4178c1b
z4fbe3078db9bce9d86c0d1b67a376b3b50e48a2476f957801c6b4584df87654dac34185ab52553
z5d6b5da8544f3d310c7283b3e7988a2e27035b7b176061158590e0c2f3f328fd4971944f95a7c9
zf805235f535a8efb62a5ee2fee2ffd40e9c1d0e4214146e0a4dee4523dfa5e13ce75611056fdc0
z81a0e62abe57bc48a41b58ef5658c69d5aeac1aecd03914d5fbf72da5b6d68685d0c261e235d05
ze0dffe8b1eec46cb3c286776b8dba8726d10a7bf5f12590b12cd292b78f52e46473bf5fc0f71dc
z067fe5946152a0092e4c0e51c2ebb33f4cc43b53ebd5f612ff1f64274b3fcd5cf3b548164af352
zb2f5ce2fa88299535033d25da1b76247af6bc634d6b99ada4762c8346743fc0724390ea22b3f48
z15d6daaa4c3aa66bbe9fb510bfc7bd8b87a5248d984a7437903e5bb661f9840970767ef10087db
z2b7c103ea63868307543b0c8f7ad1f400b2e8a1ae3779abfc4dd305d9dd001e93ced7290b66c52
zf5590ef44dcb6b602dcb31d4cb51af4cf86111566d2e4119b1bfe788e980bf62ab208d5621ef3f
z80b8a7cdd5efc5dc00a3b97f22ef75f253d1e65344129477a1bc26c4d2746ef9c027c94a8cf38d
za3db858d996e08f52131d657efa02ba934530b103013fed1d05903218598636eaa396e0d1cb40d
z574de29042718b92c277db2bbc007e61b60638cb12558fe28fbcb2a64a8a157cd877f13882969a
z6177aa8526cf79d58af74f39bc5f5854438ee62c6973f3cdf5ba04f2a649fae9c2a6d848d69699
z7b3be44143eacd6248235f1f78657722a01cf962259b8ecca24e129fe35a936d1f4be3d8e433d8
zc4dbfde0cf6d7a8bac884a14e79500fbe3b1fb50dec6172040c12c4cc6fda23c8fc80bca74cbbb
z39f7f217c07b8f37dbbfebcd845ac6fa5c837b3556705d862ffe562479e8f58af8e11fbdbae183
z779a652356348f5258ec9d72108c33662b8f5c1bf4cb84c0eeb604f7c78f1c0be34db89d9cff68
z8799ae72389d0081b05476ab4b93c7783677163c5e5fde2fbdfcb80b80200d6c8903e8016e6734
z41932856e937c47aa4fd0c4c8fac85726134393e7a1341a47a0a04db84573667dc482a4b4f9562
za4dc92a129a1522dfce5265f0b17929726c07762c3ff3e255a4cffa2333ea9f948d691cc2b7132
z04f9b4f7677f9776bd8d2c2dc3d34cb68ae7f89cbbadbff60fb451c92bb857d2427022768d1bdd
z7f56e589775f54d45b4724a83521233c3e9460031a309fafec7b706270252303d01e03010c1f3c
z36cf1f1c8852d10074324d8640fd4b017d809d0eec9833060cb9a1dca1a66f1b659958eeded098
z741dd8cd89aa0f0466e6790c2109fd90fb571df91448cfb2e2ebab0c030857b06e7e9232e190ce
zabad6cc1ed61eda81bab2f90e7be00a10267d99d3f6c8cbcd205b779c1d09d69d447507250ff21
zcd11bf1e3fa51fb721778f29725f25fba50e3b21629302a411a9f56e242271156d20223e6cc394
zdd81b5e67c06b4dc6c0421dcc6ddabc8fc63327a166c23bfd4c323637590fbf9368ffcacf538f6
za920b31f03e067a29b1c82e95c040e1c9e2e6cc4ce60f4226719efb7e213782cf8ad91819e3087
z65f4a2adc2a4f01f19b5b81da3f93e2b7bea465df8ff9c3364128417eb616e8fae4f836bee2362
z64b430f9f8130f7ce92c35c933e9b92bc31af65aeec1b5034dc2bdb531356b81818dbc365bcabd
z333c880bfa122aba6844c637f91858facc24733c628f5b8ef9c1986e63a0dea5a11527032a079f
z770392bb13cf220e04a95e37189fc4bff75d9d0eb30ad95ffa0f641d5107ae6842156b2f52b1e6
ze048d06e90c71cd7ed4107e48822b1db0ce14ab711d31e112ffaa17190ad7c7b072137215adf4b
z2eca59ce742a4408a104c4e31d1d2dbb7a83883e01cd6dbc9a8918fc1c216a06ac67401dbcc936
z8e20255d78d851a013409b998c3211247dd8e68d587038ba6e2d6ac691056ae563766fc6100b94
z248feb1722b706241c47361b2e372fdd2b3d8f3dc9230783c15981d03bc57325e23942457632a8
zc5a8d7af6e667cd42016320c6aa40ec90e9e709b2f00810b54d207032f738c0d96a1f608d9ac84
zc1986a44da18c122bb8d81c99cce60992e1629898bb940bba41f7b0bdc34df986589e3de40f993
z191cda5dc1f01eda4b3cd97fba4c162750c5f5f678ab243d9c446191a9594a7fbe409013a6b4fb
z3bda483afc173f8f41144d580bdaeea59bad8d2f5183e8941310b3ae330ba8665a0132d4347d65
z460c6397a1d6b899fc403a399076c4e6404612c82053301d34a50233e0f0fdd09efab2282c50b3
zf9e762d7c1fad23855ab71c3034fe7076fa5d56f7ad430f9a246e92713944e9daff70586175291
z85df2b5e4ee01882581aaf21ae1db8e3474dd3ff932c37844177df2bfc9783fa5895f40bb39182
z7acc35217700db50ef812020c7693bb865bacd0c5e19ea0fc48dc9843afdb76323722bae3e135d
z4f1a6965e235c2627f4bfba6dac27c1b51df3165a26d83f0dbe4f081db334492477a424c5f62d2
z88d68164bf1a69a3d55d94b6f7abf8620ac7be3d4c80fb93d40e0e1ce447ee9673e4db493a8f9d
z7bb0e3046a97f2bc328fb9c8e8da88e7a29ef2e999dc27d08872d088153a231f03ccfc6aff98a4
z7dd1d7b68264a6cec403ec694ccfbff76fb93f6988e74101162247c5a4dae85015e5b97451627e
z0bec7b476a7a84dacf13f017d508538b0c58e99656b5a8c51a5ff0178b77fb6c4a473ab6af6f43
z0b003124bac2839f6d940a6f72bd347bef6649561a9dfb8d9cfbd540f727d486ddc854949174e6
zb05de672ae4a089c1f7eeae6c356949d0af9a16edcc52558d0e26faab91c2eb8b6244558571f27
ze656fb0ea4bf67519916a81a3fdd62d4453ea88369e571b7cbb6cb67ad0552426e844e55745fe4
z5215913c7722eaa2dfc5b08f94159cb3eb0e03e5452c6f88499baaf15d1968b7cb71fe4dfbf831
zf0852b5a33ce6ac4a7447eb9ed28e6a413779f12ca982019c422519ac2efffe75462ed14c11f67
z5cb9d563ddce665b6d67451e5d1f07580560ca15a02b7e3437b5f2d09e3646f7aaec12d4990d9d
z234eb92e539390f5c82142dae475c16ed8ebd1bd761bdabb5ea3e6493bbb6e7922dacef024e2c2
zfd15d2d30b150d772f51cfc3cc81aaf25243298079ad26f0fa2018afeb6ef23b2fc47881dd665c
z71246efce3477603febf13679d4c6dd231f6f9a3fd61dd4a422183b4bfee8d085f84211f0b2532
z0f482eba9a93ecf95d4001f4d2a42dd945a18cfe51c6d8c55f0cdf8790664fcbd471c25a076cc9
zaa759b213593f80f0015e627e1a2b24d6ff39507090f8d0b9f79ca9315f28962fd276a88b7fb4f
zb61e89ed09543ebd116f3a68b7da598907654038dadf3e5415d20ddefe525d28e19bae5b5ee046
z15d631bca600d9f0299d1e1dcb09ee95e3dd641838fb6f334cd49c682eab1efedd94578e044c91
zd23d24762ade7731acad6a2652b1071b24fd7e0ef3483d3539048474aa42d04a7f859b5f771ca6
z934cf4c4852a4197e1cc887b854f62c4a7d6cbb3b6c97498574a83d4df9e1712444f0b5b8c95d5
z2392abe59dde5c283866ba7a7502e19b2f85124ded8ce4e24cb595ddc90b50ffb4bc1a11d8ceee
z635f91df1bec8c391b27adcf6c68d230b2d784e0417d35b1aa950dfc1eb1689ad109564c9915bd
z728ff7ff749384c5024033396b05652899b3ef6db0180ec7f171df729bfd014bec2f8b995e7dd0
z83b6597433f429a6c4c8bcdaa3df05330ac3ebd0a74a40f0f45960edf09878f25ae41ee9f3cf22
z44c032d98601fdd1aeb162c91188359106dc6b6aa9d2f4d646ebb38debc6b8307f77cf2a044f1e
z32a6821b26423aa334afe678fd012bf64da2d42d99f64ce95ae52a4ee612b6fc5f1ce75020b7fc
z25f1341586c2ae7507d5cc9a9886b9b4681d80e2af0dcedef5d9aa15d376a6437ea9f0125d963d
zea87a87119f18ce1727b1b16eca9918e6e675e941a1bf507b6a0a4ffa9fbffdb7a77cbe54615ff
ze2f7a709664d16f560209200c0e6c175dcb4123165633d3197f0eac0a688c4214f836b41ce5f24
z1f17193a22fbd9ea2a2a8d644af5f8259da767f55fea3b4130b30a380c3be0e82d1de5221d4a92
zb0179c87ce1afca34e04e4297346145df0d85e9aa59ac1e1a4cf8b1c073bb15a84d62e726684cc
zd20f6efa007efd965289b450243bc7ef9f24a062bac1aa20c161620bd8fff4a0d16ea1fefc5ecd
z35cb0702ad61383f733c81b3190f70795bc5872cada190832dd6721445a5a5d1dc11739e78c092
zf6ce5cbf6d952d8c5e8e2108108b3ac63ab6ad9e16a203d1ddccd5a400a5c492979b5374dfd65d
z89aa10760234d4f3a77389379730c725a7783eefa84e58451f2cfb904379d67135f1664f459ca5
zcde2a7842ff97240b22daf5c42337d6abecda440454477e9a92b3b799b16bb7ad35e9c7030b662
z8aa23421e0f50ae92ce913a0bd2b28e9cec9dcc9a949bda5190d5faa2a99de39c3cf052e887b68
zee63e6f9d837a6f167afc6a3644af84bc13ff227ab9f6cc6942323e2e870f45863bb2335884839
zb59555e541305d7c85f0616551d005ffc3333d60b9a1eb130c4a3531a6e1f1e3c8ad93000764ba
z13491b111da3197be3ed9cc406b24e03040eef06ac38f97d7950f0efb2d3e3ffbab77df5b56370
z1514526c58c34e567378fd53fa9c61f5b30092cf600af8ded2aa94dc75f49eaa689a497445b0f0
zbf76bdda429b5933acf2b9a41d14e22e61e1601af11da5db8cd84a72e4d99408bedc435f700114
zd691160989afecedffab59df09794416c64191439ae705d2d4b4cee40019af64ac1f9fccb52981
z68001c533afba824492ef494dce3d680059c97e84bc06ba47ae433ad32ef945c5bb933e316de21
z3119c4eacc21a5ae95ed4b84ee88f6cdd0f60e9de5e09add95f5433a7c3e0903534fa1b5c7dbda
z9b638f9d28f9c2fdf03ce0d314e4c9174682404bec5d03c1190816e0329262ac90f5d541cf70c1
z49a7f1f64192c5598cf23421d0b8d1325c5f6dcd542015c038303afb248634d4923a757b11bc20
z774640cb95f8f39a8c09e9b0633858049f029172d615e79d71c0827ea4974fdcaf7a03727331e1
z2c8853788a2282c229e5157c3077a1766b1aec536322865081711fe0b2d2f0cbaa0097c7ccc727
zd59c58a30f3a4eea3c22a058eb28e1dde5c2aa1e0637835e9dd833a717a29f06a03ebe90816628
z360bf0a6b2e0506a2ea497407867c6fb1f3397cfd13510f0da91186a8df648742d2394c598a1ee
zaa9e436319cf89250224e403a383270a9b0c68e908ac2c226cc171bea014088defcbe9fd90783e
z534793c9a274d409ab02f60c938ed614973ba6c197d5ff3af4e70f10553dff927260c63b072035
z9d7e0b95350130564729d97f06cf07f44b370d7299c503481817811761fb18e02286197dc64aaf
z80f8aae9815035a8abd45a9777cb7e24f05abe17dd54f1edb321c22592890a4fb40af5b2446b1e
z0b92b7b6e0b6aa2c60977d996e1ec82971f55fe441b076d135064e782a0093f070c004bbe4a255
z5afb789929c0fb9111eaba1393e3b9e80836d10dd75f28e67fe2d53db967111594e5f7203bb5c4
z06e877b6544d6f157e36dcea5d10cabf84b778963dea67da0d6d8560bb3215883e852ed6587a8a
ze323447880c8762c553565c398e468772c33fc332a1cfdfdcd43993174e984e0461158d9bc4c0c
z29a1cdf78c0c86856283085f3670e9cfdbf210198dea566c485d51f0e4349f5e61a8e4ecb2d69c
z1c127049da65f3383dcce2a164bfba6b86a6b333be48475d29c69c967ccdad4927678b02d588b1
z5b12990effd57e707a9f9a897d6e86f18744b9bdf022da8f356de7581748ce2c9c341db2611de3
z5a530d41b970b879a0b52296ed7ad1f13476e43bb268be57d1be60f0d0172119c27467f2ccf3c2
zfc17727adb743b297e2337c51f6c6188c990c1ae7fc0f5dc9848e91bd6fb26276880b66dda48e1
za403cce2ac779a2003f17ec7ee4733ca50e85746d7aed0f4f38988cb60d9dd2df57ecaabed78ac
z57e5d7a69c7e426c84eedeee14396e468d7408b1c585197aa7c2f883d4a80f4b82790651b2ff8e
ze7d5956f8278f13262deb947e348ab877097844be8a3ddfb136186650204f8fbcf3487a880ec80
z3435185e3842cbef3758db2bc767daa65996ea041db0eaa3f90f6f9944a74255c36b49871d65ab
zc206704d174fb1194afa130beaa645d94d8fa73fbd9bc3d3017f51b93d1ee76b7b58530bf66520
zba215c48609fd230da7651966f1122fee73b6476ec93489b210c631815f824d94c506cd196cd2f
z83300988dc359c995d1cb0345a451b8733856b57e71180158f488eed997ba9fea1f51b7e7bb28b
ze5eda65f5f5fc8d0c7a4cc9c7f08d18c243cffdcfa3410feb52e1d84ba9260f0e0b0b847fab0de
zb5991124e97f7c72b61791adb36ef5d6c44b30f1fef2081b4b712c5eade548b4a08114e39883f7
z36565df1045158aab2fd0594b5e4efe76ca5e690aaf12a809da1efcc3056f9379ab5940f375b53
zab12be52811e1ad96b67d7d72085bcbf3f490058ab809b90932d19fc2ef8796488d76d45644dda
zcbcbf2e0b570f0bf38ec5116941113692183f80252179c9aea007b23baf4cdb59f4c68a417c57d
zdff3b7dc3b2bf4be6c3487dcfd834991671f4526e80111f214b8243b041cc39af296f90e24a1a8
zc202d79e8f9aa9d2792f177659154931cfc619bf09a2d0e5f3f3fe8f3b96436e1bea854e67b832
ze2c9b31ea049f6e1d6adf75c7d34df1fa00d34155d24ce3f45245490c14072ff627e6bcd64dfba
z3e10e09d26cba113c9806fadea47f1b495f2da46f76b6b7a97d8152344aa2330e6712e60ebb5cd
z50bea13b4d9206f758ffa2a1bdbf3aeaf4b8fbf1378cc7efd57528dcafc15e092b190cb6e4610f
zb527a97035b9ee8738bd54d44e606ed81fadd36160d6e6a3f9bf7d56804d0ad9fcdbbf8c3512fb
z4ed1415c541dd020719ac03adfd11623da23ac52d25c9b38a2309352bf1e579a3660030a679b36
z2739b529385ef4d993d84720fd23e0750cbd67a0acd214906a18cc2a3771b2f4e3468c39576391
z0044f0047514f8fafa4c5bc22bf9915378d88ea13ce85323e770c004107da238d4be742e78e734
z8dd2dbf8fd686c178aa46ce8482e889f1d7bb5cbaf793b36dff43242f4a92db94442165549dfd5
z68934de35c22ec18a64d4989d4125bcaae074a7f8ddf2b6509056ec685478bbea3a4541ac4c2cf
zf4e7504977c62f004917514401bbe9e1a6fa2bfb04f074a6112c5a891ab885d7464b8edaae3125
zd23087682b5628bc777a32d33cdf33b352015b5284ff582a1e44e2c0738c24dcb71951eae77cd1
ze8a3a3cdb1c5fd225e9caf14e2ce377d155a2ba6545d1459e32845a347ffe05cc6741db35f15e1
zba5cc1d632730e068c5650ca91a87196329129478753e5ae5290f20cf69c06ad6c2bafcddf3ba2
zce41c9eeb48d08bf86db1466087727c5168d7badf4ce5b3b22b012a886259af7e6d7e96a4f104d
z3394880b5a24105cb9c5fc3a899067d4abb63cbb62a18645d8ce8b782c45f2b90c52b764fad201
zeaaa20f3548c9566612cc9ebd0764abce3df0626932fe3ff062630a735b791603d7ea4991acb76
z7bdab528715c5c3eeb480086dcba79547ee6808fd8767f93d399704e55e336f743eb229ade598a
za2bc9de646f2f504fc57bbab1dc3259f5ef4ab2e11fe84902acfb15f5966b40506927198d9f8fd
z1e0f5e7c1b5fb95bd717844276a6566ba38edc4ebb066aa02852c95b96faa804701344c90ad67b
z4e4fa72e4b0a8ac20f124c5f9f67c537baba1cd54f06fddf75342b6460b05d549d045718075c61
zfa6f48d55705c5fff6bd47124e3a02511a1cdc3761b6059ade2fa097470f7ed6af7097fb3f2b88
z13c4d46fcff8d725f1fc80918cdd4668f20ea472d51115aebd9baa0dce8a281510e7243e25e352
z9daf292a9f1ecbe11684e71c97c6a14d12dfbecf433bb3cc80ed1aedd23f84cb7d99845e829b89
z7891980878fef2845fca5cfdb063aa5a43b2b87e7758da2199478b1f3ad2bf92e3d97e92f19266
z7499bb201e12bba7d748aaff43e239d7f0da77f8e410be57d4ec3d7f60e49d5ab2d61d7e73c22f
zf93c46f9a4541c1901a7fb9000623fbf26e9d40ee6bee3806e1c994631d435a83241fbb7f3125d
zbda68007830f94567fa9b99d41decfcf174091bbd3ba2075d7fe58652cff714050423a492c4694
zaec61d3f89fd8e42d21fc906ba755d7801dab87c18ff8b5966b379f0092e957df21ba6efdddf6f
ze66805d623b21935ed96cc8f5e0843b7d63b46f6b754ac98a0a5ecfcba3daa60587a8c06c436f1
zb464b46fb329bcaa689ce32d607caf9794f339f8e59f061e1daf520f400404d3eaf1ad013d1229
z516e7c537252dd2fd6aefa9a89b124de3cfeacadb7e98fbeb04af0ae7d13a776ac90d386bbe983
z9b261018484dbe43ebe6a941ecded532db9320158c72353268d3a0ecc426acb9076269e0f661be
z44fb23bc747471df01544d3ec32dcbe2d3020437d6f37c67ce437458e1e046fa8efb3a1591f7bd
z04fb4bfe6b58e0f5c3ad3054e2c165cdf1d6e746a02f05fd6ed88e433732446d1afe4e03c788c3
z0377fd4321cfa15d8d61136578079f9b00fcc4720e0a75f70eee7be996f1af62fcb1dc599fb8c5
z7a569c54791274708728fffee0d8ceaa9128cef1b3409d53d6bdc8156ce126eff01bd136427e60
z939713fb1f7d15f7e19aa41bbc92953c32e0c39595135759f2dd4dbfa6e6567f30c713d561d055
z471864dc3862741f69731532ca041bdff67f6d9852eef60d4266fae56736cef44d64fd176af6d2
z9e768169e6f93e9bbb7a228ca6a20fcac7908f8b0c31c0b067f9c7deb356e38370e1740ea31f53
z4da8ccdf66fe9d68ad126ead6338d2228b33d14c782682c8b098edb41d6e97120234cba578379e
zc7350e046e7820b9f6627a2af3808976cb765d2905aba60252da3831e67483397b09d637f165af
z9a04ac03c74938834fe6861218c355ae84f95e7aa0af54d74c0635b5340ee342dd1b32aa76577d
z25c71d60d69ad88e73d634f59de877a7bba28f793b585d327c6c39b084e91d7eb30e00f6d9ffde
z5d44bcb4fa610e0fedca4f48ee40beaa08f45121cb8f5a0fe4df8b2f221e2d6c6bdb59ff8321ac
zd0a7582178d82feba00b90a68ebeff3af0565df148f2e21651af3a4daf9274ba72d23fa2d762d1
z9f32ac5b5d07140e8dfef667ab667218eb91b98f1d01fcb23bb653e86e88518fa8f3b7455a2c89
z19c68a620a18396a7f1aea6efca2141b4b85e8719532b40fe864c6809c561ec3f5cfc0d2f9f6b2
z5f2c9f7db82b509508809c4b5d174465f3c63453641d094982230d40bb4e446762051bccb1b6c5
z8ee3418e361c7e24178bd5a5d272bd9edff2a1f49685ec5ed5a17e9e098b72ddd37d11185fd44a
zb0bba7ee120e92daf79effb0119059cf5ea4aab5e019ca6860a511dcd30b9229183fe7d67e2cf9
zbc83b0b5c634b6584b9b94abc334907eba92bee7f6aa1ec7c4e3026f30867f1209a6fd7171f1f8
z583d7db7703a52294aa826c1f69357898273c0e24dd0dfd195c2d0ea0190832bf5f82a2f84229a
z59f263429ab1f3e583668f60573794cc2565ce6ff36b99370fb237c351b589afae11f20027a45e
z0c44397c0706de4c6eae084abd0582ebcb26751f085b1dd6fcb16c869fa37813936f73eb9d8e09
ze536e87334dd1b4bc495291d3763bdaa7b009911d51a718a5ab04f58c643124aa419cadc93652c
z854594ff9223456681982f5e8ecb377684c3e4f7a81aed75ee1cfab5b5ba640b91e00a2c232b76
z31bd9b5df4bad7b618ae9786ef73851db7c6e1223cc0436ae746f38dc8506d037a0e6e96398f5d
ze84262eac5f7f0ca596c769dad3519cf9f0c0f8c78c12849fc98a5d705ecd30b4c504a4928286d
z8f0d0c645c020a0fd71bc26e2a0fa6bb2f283da3877280c58ff7d5aa88b37568a206fefd74caff
z06ae31a10281bcefd2f7dd86eaf98689f29e1ea07cf53fc7bc1d93b4ab7e0a7432db9b4e14245d
z3b9c136ec7c3d68afcb5cdfeb9f92020dbc0682f207360346ded502b7a419b4f7a34bdb2bc99d9
z03003e84e1b51f32add40938489d9fe7b26e63eac691058ff0cb599fb4d7e05ca96bf6401d5439
z9c238e2596fd4fd67614df21829256a8027f1a2cfe5280064343111858ab511395a959026ca8ff
z2c4b0a00ded436b3d4f243cc00a2eeea6bdf456faedf73632dc55190786b05c9722abb024c0a28
z5ebfc802071ad57782013d6b5a54b101c6c7637364186e7d0d4fdecb336c5d0d62699f360da2be
z15ddb064e32d8a0d10835a8f8cf6b2fa5bb30482b170633973ee16a72fc3fc1e4e2805d10d0bcf
z9f13bfd60a474071f3b184af1268edd053666999d2e390c5c291f73ebc8ae96639dbd5f68ae406
zf37d9ea6dbb5f754243cba6f56045abedbf56a3eda3669d904d9237c1fb38e923d496b41425cc8
za33519dfe6fa1ae0c3b7219940eb7a6c7ffcf4b0fb286d633f8b368d1caca8f7565dbeecc3492b
z3449648c2eb569868681139c105eb92bc6768441cf7392d2cfb3b3407f30540aeaac593471aceb
z0958005342699d21d842638abc9f479700fcdd25e755f188af040dc1ce11a5bbaa9da359deea9a
z59f6d672bae1d47fae5897adba2aa4560723d8365f90953767bafcbf3df2172bf0f20ec06a51f2
z13cda87b7762c219af30196ff0d096dbd0f84241f83e5fec230a4f1c520a453fe668d53c020f40
zed00ccc8987798cd2d61b7439f1a370ef4f138f4211aebad3212f5b63e1b1463db333340c46056
z5478bc62fd1e343918924fd8be545e823f80b3897aeea10b61286036a823d5c9d13da2df7d2321
zf099c557c36759627f9a8bd2c33ce9dbc411e22566a366d74f5acb3c5bd4b8ea618010199c8e2b
z59e133608af7e2bc0e3134b4da0e88ff3851e58db17cdd25f97cc9ac9fbd9e7edb98b4003602e2
z9c7b6d891c4ec5defd857a8b49ba37fe6cb198601ba837df0fa48b7afbae73f144a9e341f47bf9
z02ddcb3ef8c0069d8dea13d7f417c77c0c69ae513d9102fbb4e9490d2c7d9b3404c6bfe0c4c333
z2508428ea60be404b27e7cf805f8c5643767613a3d321626d9514334d6b25b45b5e3e2a5149552
z4d7ee343a216b2b0a73b773b866723260e2bd1f5466305a27b05c6adda75b095aa05be75f5b56e
zccc4b5dc8408f8d85092e8d1f5418b079784681806fd251c24802d6b1e4bcdc1c3296be33b8c75
z7656fe0e4e348378372f44561adbdbab2bc3c63694bdf75590e5c6d8bd95d1988f9723c194f4ab
z2401c793bd32437d431a3dff9f6368cfbd6706e4240386a9e31ec817870772cba9cdeca93e2e05
z948b393848c88e1af1bdbd98014212d63cb1027fe9673113ef16db01f5978b089d0ede34269fb0
z6a2d6f1ff9f03297af179cd66a458120b48e056a9769739435bd3a3daa547e4748c75760e86b98
z5fddf8229168cd1d8c07542cbc0f97ed73b9ed428883398e644346373aed3f65f5565269e8fbfe
zcb9193d99b45ad802c8ca80f2cc67afab0fc2c60b3a4b1c0af751dc89d452b8dfb48f2fc76311b
z31967ec77672e2cc92d33431803376e9b6aaaad98ee4562f2d2171c1e98ecc012fe28670c37ee1
ze664b1b89a3f496824a86ad00019490b6d114c7b851a7c8d8d9e060da20f28e93864e38d976ffb
z6f14e666b61f1a9b3778f8757e4fd9b55b75ab86c7cb988151af52d07488da03e7c2d4b8cc6ebf
zb19bea5082733b1d2be722d263dceb0fe04fea3456c4a86d0967d5b57ca307bd0e1c4cc5ec0379
zbaea2bd93160ad1f5191403de691783b505298dad092d11714d34a4303d6d7ce5bef3a1f38f39d
z750ce7a911cc6469127d7549dc77316cd5b80ca8b3f511444064004f6cdd2d7f70f2b74f93c12b
zccc7fa36cc6898c0ace8100f3b3924b009622b92359c000f94986a0ed9f4fda81843c063649614
z1e00988ff3d259abf1c66d88790cf5144f2cd8a48a993a58ca5d31276bedd2fce3950f867153c6
zdc8f4521d47402fabf3b7375b6645f754936307af16806b7136a3546c000ea2f8954d08099198c
zc0ce35106637b0d75b0b1fe85728e952f49f3e3fba63c72dd22d913cccd15738a8a5a87e1e8cba
ze5049ece96bb520d1abfcce44d27eddf71f321a60a16b7777a52098fd71ab5aee4218697a4b4e6
z5cd27bf228ffec49191af0ea99a1a2e7fddc00af8ca9a51da6df2ed39a2fe3a220ec17ccc3142d
zaf48fd460d113a6a9a2c9b57ea3e552fbea7db931d3e5ab4a43e7131c1b0e72bc88ab70d1055b2
zcd5dfbfcf90644b2f17ad07b174de5237b7aa7a4c90ee5b2ab5db0ae8c3f2924e4ce1a0444a544
z6c547b59d4973282f0238f2496bdea152ef5a7346cf422ca5490e4672bc8cdbe9e0fa63d60477b
z583c0bc4d640764bae245cf3bd715da64d36c9ac1d6e0a97259562028728302905b31da425baf3
z35fce612722c984246aef845639f7925b657fc2eb637d7fceef254b55c46727d006f623be3abf8
zd210fd3c0ba6c6d4ced8f3b9d43eae03b0bf0218caffa044fe9e3d49a6ac8bf77faf985a189094
z1c0cc1f44c9f44bf476c0e78685b0fe281932217f499e4f1797df96257a3ad9c3b4abbc3ce7037
z8c8e62d00bbaaf622fd8a4c3f8fecf808c7e61633f4d96b1e117cfa0527c24d792016c18336abf
z9dd45324014e10f9892c7ad6873300827d55cdf0700c6f08142cbdc1bae072b93072cfe1d61333
zee5f854419d3f98efd8987e65a32a9c40d2b131c932ad943074ae468fb23569807741312d14da2
z599c6f502c06ed0b19af6e2cc4c8b17af98eb4e487131f24c97580d778ad737091101c73eb4413
z44ebaef4ba14724740047efd8ad8fb7903948563bef531bfcd4d94b4ea0025a83d265b05a2fed9
z31a08044d524c164033afc79b17a85388d81a8c381c123f3f35e3521d5095847d22379cf2425a7
z6f6994331620753b93d8c550bb6f36ab6b5b566d24f5f3cbfa14bc2fa14c791006982fccb44957
z092a2dbb35f24ecdf7c593788ed271d0c429f20375846272e03228c15dde9475f7d66d32ebb65b
z1a9680dbfbb7f73bd57d80e4464d13b6222f13ae942e43158427de2770d43eb45810f4649352ae
ze399f0e247656857a4e8cbb985622f5b501e41793b60ca7459902280771f70612a0fb96b670406
z0c4d4f23577d458b118dfd9a42e16c1b6e8c6f6216348d5c715b7d6e3b8eda74473c86e9df9ab8
z6c65f28412388a6932b688177e61e781a726053c0a6e74e5e12580ef49ffa8ed06f4808bc21178
za4565ad15486514f397e55a9db9f7f0958bcfbd39f439672b74cd7fb08c6feaea307353bb025e0
z8b568a93dbcd469ed18a3859787e89ccc37157ce2226346759a12ff300ceff1f417835e54bbe75
z94d504b1b811168210367026c9c005311c0c6badef32fa2df788f40bf8715c93205d77f9778ff1
z58733171dadec023e66e37f4809fb6a59964eb21056c5f14b22f506efe8a3a486044f1ebe42af0
z45ae7e01f57782949123a9d7c63a3d1b2bb633dd4d32e2cfa436ee7e01518db5f5819d55de6297
zaf72d54b81ff87f527a05d22f0244719a0cefa9a9512aba95057461334fb9c790383db9c652a84
z76bce7bf5e09c50d151740528cc756193188221dd570b62285f31f96a52a7874571a855196d5b5
z45579de2fc70a334df434982d71566fa103a0aa936f5ae8b5b0923e09b78e5363475be0470cdbd
zeefdff19a516bdd81b15ba043fbd36075fdd721108c120c3deb3eb66371fd4e592157b49190653
zb891747c22307735aa7bd86c1824202ea843a537c3df9d35d2f1ab4fa970b6546d3eff87538e99
z74ba432191e615d1148d23f3507d3c61109a1377b96150ad183777977dac794e647bfc147444b7
z68e8c6d6904dea92ec26b9703e926097d1e128d642eb1b774dd4937696bf1ee159514c5c1be0d5
ze63d4a803a96c9717a0a5ee4d868a0eb1d875de4ba0669cfdf5a3a596859e8a0c6bca9ac5ecb9a
z28470251709282e711f8cd479398b291741910be43af495ebcec98aba85515f93cb69d9e224c0c
zd341c1ba8e0b76a4a17a3d2413db867e3c2d625c9b208ab79aef7156e8c3f1924c1d94760f1bc7
zea583c3f03df2e6e33b70c2fa1c5ce44826cfce72561447c86b5d2a799d7db24e5fe23fc274a1e
zd19d080bea3eaf030c6ff27dd150aa5c7158c5148ecbd5fe650a1eeb28848c613c4f738ab63db1
z3aa1217a2146046200c63f0cb9b0be66276f715e4b95720a730910563a5b4ad03905c9c3422915
z52b6a7329f9fc960cf565db539c6436819a7a5d2e844fe1e91667d3281f47b977868b29df1b09a
z3924b6d3aef5791ffd59271176d9ba095783f80522a4b69d94120440becdb02bfb07674db1be16
z44446497a34971c81815dfd22718c8c67b8c593c185959c22fe6e6d3bbdd65e29531bbd6fc1c70
z584c83a7f0e0f4cd0f8a7cbccd5ee0fb3fb3903cf4bd1332e9ff5c4009261b261de31498088f2e
zbb34659601c00521f6d4a8dc32c7ad990984e836f8ddcecda8fadb4c43bb15019ae411f4b5d5c4
z4bea311a1486125c97a4e79afdfa9fe25542fa39b27b8f712dbf46bf9d6ef6ff9287e324dcac54
z548a3c8ab3e5e874a3efc96c7c114b52a12116ecbb31c29927e772bc2a97ace6b6ada8a8718c92
za32f488383eab176471b8f9d66a7a45e0065387e1e2bea86592da44bd78fb1312114a44277fcd3
z380edcbbd6253d0e8656e5223ef5fdd8135db2ac168592b74e15a19504af5a01bf756874418f8d
z6106570cbf440aa9b9f0ad1c1a1355fc14d07da2298a729d66f769092cf92d50480a5ff4bc9b63
z15618daa7174e0d43e8bc1ded489ee91646d2e3411dab3c060560b909ea2e4e54d1e8e6aa10b64
zd7f0cfcc348224adc1b3ba2689eddb1421f2c75c63ff52f5458f2ca83615388ec9f0f2d65743fd
zd68ac733dca6f7430770cbf7cb9df1dbea515f73cfaef9809626156f8437a418255687f35b076f
zfa39679e2b8d446b56ab579e03942b763f06abf744bd1e6e8d155f70ba8a761257ce16959aea03
za49ba86b52aab21aa23ebaa2ef9f9c59af7618220594b22579d8bcecc6684f9357a9dd4c833a6d
z814ecc1f130f5a0b3a234bebe35665b4504df6214b40f7b575986f281ee2991bd1b2a2860f841c
z95ed1c980473efb5120d7f2a385b468ab723b08b72aecb07869d4368bfdc5152d321e071e6fdfe
z94636bc964a744b98beb7d5575a571e22253be439db896caf0df91d52af00e64aa2bc91063aed8
z2d57e0de401056baabba3cf32acce7584acc7fd5bbf1173f9e732aed1230414c82c3cc00e289e5
zd707e58f035e228cdd59f2b6ef78da30c8149f703596b653ef0e7d12397e1150b007744fd0c40b
zed98f68ed89d737dd0c5d0ecc2ad94bf3e28db5c7330daf521d5da156b6a77d499c5be66a121cc
z85a7befc9f4b770b37fa05bd85e16fa5545eeb216a37b37f288228949bd61749bc32e612c06b19
z8319528e80d8998c35f3c7e69d77871c7b2cda1bddd43beeec74bb423a26dbfe8ee0bd8902c88b
z41ef7f836028bd8c9b438ca7171d955f9f18a754480c006fbc318bdef57bc772b076364dca09fb
z914bba2c79b87fe79639b4b4d4b27b07555a2f7af8afe961af00aba45670183bb0078f1ee43972
z93e6c25a9186e54774d3030e7eedf08d2e3734fab824a61b1453a2b1b20854d2f057fc53e4c093
zfcbf485316ee584efbd895ef49bf1a45f4ad4867f8d3338a7f9f6b20cebba1fdc9b2d1386e2117
z86d46d6260245cd7a024c790d3c49b3c22cc72a7360e06330cd61474244de2723aed1970097055
zde570449cc0b6a92ee53981a66355777986e297b6d45252c0c17fd941152251246b365785a7e2a
z46af44307c74a0b470bb86a23c4ec458ee1d32999947d93cceb4f95c9d0026bda95c52597dae97
za273731f4adb07d46e74869d75dbc6d6460d47823fd7724e339a288f9b2083bf93868797e12d15
ze9db166795c00ed17d87ff28e261ebe3f31202309e488a71ae7aa9c1e3902375d0b16d42fe79ea
zbe1e60e696ddd533dc8f9be7ba3e93512e6fc52d4afdf9e402bc5ef318ba19babe1d4afdbdb011
z7186d4d59711e20296e77ad330bbf3d99cafc367d0abbda83a601f26e94587d7693648632b3516
za248787b46d8751fba3dc19d1ef1e67465e00c8aee4b01763657d1292a22e209da25f2c9e88174
z41280faeb0cf3f7095d38303e95edb584e8fe547de2bcbd8a5f47aeaf998c0cb49109688a09dbc
z1eb4b97e0c420de9513197b4cb586a02b6668289423dbeef6922697ee9c18fa68c94ac4b08ecd1
za6dc8a9eef061f96eceaaff808f52dda144ef19d7eb0f1f6d6690b4921b2235b37e80397b1a7ca
z780a5a84c71264fa92245c92631fe1084ae4c2c6c6bfad90fccd47ddf2c449009f7e9d25257733
zc918f9e9fde2c9b0aa85aec0e2c7529fdd3dfce0629b35a7b388b6be718721f46ab83cdfbe4b6d
z76fd6f97ab417ae453d2510dec5e4b9efe28bcc32d7097a07f964e5bf122b9088f133f711be235
z83d536ab9d6ee07a8cbae681f8f4502d09e410c427c13a9e20b10cfca55423f28b3c9579c47ae3
zd69883dadc2d94c4449ccf31b155095d83aad78561218bcf0d23d68cb00534c471df1b7cda3dd6
z57b4ffb3a0960ec18bf12501ca3f8bce691b0b44cf4e863782165bd2cb1b7c6d68577af752ef75
zb68236b7bdb78563202412b2b45b6b6e883f6da1ebfe1561081733f5d60f88a3da2e354ef35f27
z04f3cf497967d91442266f21add254e6923fc6a43d30378f18bd3969c50558c4b50ecba3360c78
zcd3fe3cdb34c5345234e8690f8971682630ed6b68e024233a77b1996860dfa7caacb2dd5321226
z2ab36009fecc220a908a3c731b04b501790884fa5be824c8159411108860bceb6f285593f814c2
zc1bd937d6a88259e38b5b995bd2486342c45a26d5590def4cc12a8ed27e260adb725519fc17e2f
z349f90d499d259aa5451e6531de865d363147b0d93c14fd7f6ffdc88a716cf4061a6608125f38f
z2340bd17b191f95aad44f335165252281cc8fdd1d63f638ba74794d1ffdf1566531051cf8ef18a
za206a429b6000a77b87a4c0bbe51c201055f69867c083b7f6baef3be54ccba665dfda20651502e
z9352ebd6c99afd9f72b9e2b69d470ba3ca71e8b743e423676644f6bee70b94c87de1a844787ee5
zb82238de06ff90c69f79ce63b8377823a5d663671f731ca6503b22e58dc895916d9eaa0d14936c
z19fecd75d6a4dda6f0dd1767718560288ba93cccf15f6c74f3c9b2fed89c6ab2f951fcfc509b5d
z34e26a7c306de011ef84b53719ad7c2020900e93a57a4e6ed4e63b7cff70659b326cae638b2dc2
z381b737e2a19d4a441389d54eba9204dd9bf9d7d58bde2597f2d137550076ad8eb7614fe6e3dcc
z7ea95d789b84578bcc5fbfbf419070e93876c8bfb0daf3ce94539da534a0a2645dfa85d8b233ff
z042ff6e76763b8886a484d4583de7d3ee4683a1b5c5da16eebbdba75c33d3dceb32c51fd253c60
zfe7764d5394a5f208a9f16831d04a177102214fdcdcf8ea5ff7219db879542e7c4475477ad3c02
z0df71e0baa41506780f0dea92d0423abdaae8f84bc8891d1683162a06ab6c6c8ce922fc15878f1
zf4b81fd0f65521359b6634ebd50f69793c5e7e9f1af489a3129f5a510dc2f64e0d2d0f0d149fd1
z0081ae4d78f6f07464d67b66389614574c803648bcd35c4ab26e4b87e5153e07ae689a5ccaddd7
z24330c442ea602a3f058db368957c15897725ca241771fe600137f2fce61a021c69887376d77b8
z1f9a374142abf6891f52d2fc3cec5e8292758c24f63ded2efd734bd48f8b45a008795ced5bffc3
zdd0846cf0581e4718dce665b143b4c0f457ed8ed19216c2ab1f5c1bb2bdaed5aee54774fd5acc1
zded2f430ab90bb07616c4e1396fe0d9c2bdc3fd380b287dbecbebdc0bdcb05324dd2103923bec6
zd58744eed7295f70ee77d14ab78c5f306e7ae4b89b7cea2d131e8b24e1a8e6467b2ee31b7e20f4
zd3db35eff6c8bf8c6165dd3cb3f212d9fd8e00108cc82c78d0a24208682d1c117981d35862c503
zc520756e7d63a33423bd085f4f15bf67a1b8e7e3c1470b7a19495eb3c6821163ecb24aa46b11bd
z359b1ec3cd1afbadda4cd401d4ed61d734406635d223f50b6cbff5fb2765e7c92c5eb8a9d9c3f3
z94518cf3acd13301e4564c2e4a5ac6910ee8ed3bdb72f507c8f5e9362975a1f6526dd2d96911a7
z4ebd676c59e13d24c0f3693792601ae43dbc297eb68496a3b9300a2c358bcd8cee7cf2b4375366
z561a57db2652fa98bffa72c090691250a8c0225a51a1605a82dcfd51dfa039911d79a1b614bf14
zbc8a309342686a3b629a00b1a4773f44f2f108c149d3f115b7ea0e617f6fea3861bc8c5d500e2d
z0a88c6b5f9b2ebd8c5e15b83fdaa8bbef70d347396c1ce559c063488a6d5bb143ef866399a4043
z97a321d5038d8a666b7f40aa5466a11eb5b0b34e0f48d6e8ecbd5954292ecec55e7aadd4d23259
z13d8733b474ac06b13e69f26f2a6a41c67a5f2f7085f817846e4d337e3ff26c360145fb6fb2c32
z6857c53589b2f7c5a79b85ccd9a3447435afad71fb722c800f444c4bb107077407e5b9fa7cbe00
z307505b3c7dec9342bb6e3a5c5fd17992311e3e76bd51d39bc1033f1626c0667371ebfe3907d31
z0c0ad373861e52d6e96b3f1690c6d5d04399d66097fb9d7ffc7eca4e979e19b2cf6ba664965c7b
zcfbea44bc2c09aef0fc9f79d88c29219dd09f4195238b50477e7fc60fb202eed237c1b70880383
z9b13f79d3430199eab7b8e1e0f5a5d64c91ef46c22c020bd5a4b1cca7568375ca42d7a7402f82a
za3845d9b24d57a13e8387e767cd79dde1887d48660d25ce4fa0383682117501a91da11283cfaea
zc154085ff21a4138e65fce1b30e064f48bc5a685503ccc3abf2b97715c56e956c65ebc96b30e34
z2e9f331268a0cce0b1d05ef6d0f59a83514484c413ca055337330de70b35cc92591385c7ff9d32
zb834ee6fbdb7d692f4a8f0109e34a0956562ec8fa625deefaa7c1c92c25a86ec0f4f42e86990eb
z685ab5821e980f5e299ecf28ffd358a82421436046c53f8630e0dc3a7dc8edfb47f49883179ba8
z6819ca6b27d8a3030030fb5a37cd49fe507b5b822095d220aa6252f8af32b4d857bafcff692a51
zcca98a913ffb8d39c3f3e511782e6b196790e455b3750f8d6754626acebc54028bae8864b08e0d
zff9aaee379dfa445997aa44b3b56bc0d8e29afc1fdd9a49d2466574893f38fff95704790ff4ebf
zb47ae10ee709441838aa1c282b5344bb2dbc463aa9db101bca3c3974a7cb7dc18867987bcf7209
z57d3bf98427a88cee9ff65446551e371cc2a05f51522937eb0b0c22d533bba395e0860200b3d83
z68034466da766fbe4ec943aa2ae20b77f5c28241e471578f62625dd39378c2d6abe336147fda9a
z4d867591f793eff705741272d415c06db85224852df489b1c514fbd369b97389341d16e9784ab4
z5512532c59d9d277971ae62473f3e7eeb4cad4d36b8c63b21401ba48b1586987946e7603c89c53
zfc75e02b1633b8227d21da8b66ee7d99d899bbe957784e9099cf048316fa78958d9846118c58f7
z3f4bba22d4eab298aea9fedbf441977d8dc9263051a8e27f6cabe98da3c58c658f5b0d454b92af
za94b5058984f210a849a4afeb5e81a537c9d4449c2cf285a1a3ace13e591aa178e90ae9677c307
z0b432d8e93fe638adad19da1bdfa97ae79bc36dd5207aa2eca74d742e42dc37b58672c0103da38
zb6709731694343146159759a69f4c2e88f499a3788e04b809f749fc94cfe9e507fa013c397a0c4
z177c650c1a82154e9fc6bfe3f2595887ae9584a86caced1b25bf6099eeb45960e5269c9c8b1e71
zfbcb511988f4d7ac19bf48a173cf7d8fa7c5001d725d795688ebecb847d25b1c7f887901a43993
z402b1ec6cbc8926c634826ed57be43e8dd10a9c21247d8f78ffd0d4a5791fb5dfb08ee8424304b
z31f630a5d6d33e3a782cefe45c7bf6b02eaa62efb935300a844766481b0f84b22d78531e6aad3f
z879ca0492d0b8cf7a01b2442fd7266fd01cbfd6e4df5de6e0bf048ed8c79c5b4aa87fec904878f
z408e00319123a22fbfa0f8de1a6cf5ed1f91d08107315cfe1b6236f004c6e63b5ff663b903fd1d
zd5d79a85501bb2c6eb54c1e027aaec14ee3806edfed7b086b0e76fcc8467eae4000c993fc62999
z3fddd436bf923ec923152a21a5b6f3bb2b1ddbf198f07fbbe139c5411bdbf53fd6873b42698502
z06e16cbf6d553ce75313aebaca7a325fb1d60db85187b7a20c39b96ab6bc13680da392765d45f0
z6cb60694959ac422a38743ebea49f67af3d955bff0f0540535d30dd4c4db88e7d8b6fc4f7e2b8b
z74e8a58c0b11864b9e17833a7ed78e4361d2342d91ab791444b3df224428a70f6b0f49782dcedb
zf7acfe63660e8f472ee38c31438c1601ae72590c6f2e8b2bdb1b5465c6d8be357242126b60d94a
za0a5b47784ef8692e99c3a0784576c94fbabb2ab8029da90e6296da1af845a7d0f7c3e50014097
z07fe5d3b8a12916f9e220fc82c5719cd085714e13b7a6dc16eacbf21b1339d3150f22d4a2df3e6
z7581c6a15f9669ae55a9259237e9892d240efbe85fa11b83a16f5666b23c52e4ae55668d496a48
zc186664114d812e653bd759a7815152910abb038ad3a171628c3bede0761eaf0f9eddddb6cd76c
z5b9a1148a18dc12415198f5fd1b648b7ac78a208aa5cecd62a1f921c59e4f8e8dbd1d0edc9ed09
zaa50b975a773491c0cb6d9eb6f13dfc0ae8bb200400c9042364effd71637a2969b3f64b59be9f8
za5d5dd47bede3681fbaa9745f26fcecda6fc4e46fec49bcee932bc58b1241b7282baa57df83f1e
z14199b2c04f53c44e358ef8c416686a1a85bb975db90712ec46f3cec73a9c0079f96bc5740d08d
z9078e033121ae89c59df26b6962a93c6b71c169bb295b6cbcdb840fd4775c1782e509c91f6bcce
z67628563ff3992776930df7487935a68110da648dda3d4140c1067f4f11a250d608fb2c967bcac
z1fdfbc8cd28825e2f29c34ff9cab1ac44fa99463a3a2b182950a9fe65473a5e0d51e61eb52ea3c
za5886a61bfd9e01a96248f0aab0056eedc924a949072b2f2b2650eb32ae4774a797e47db75c616
z51ab02e1cd39c10761bbdd0b858d5d38373c1d5a7e75e64b92d660a980cb81b97253ec3cdbeec4
z9aee8d97189d3b0c353171098389292067be471647008f63fa492c7dc0b2eb17e87bd8826ebc9f
ze5dc1d4b98fcf40932a155b0f88c7c74a0614af2bbe0484c3fce848b9227f28ab5f8f610fd0bdf
z49b3ae9b15202a890eefe50e6fc74fab19e0fdbd60a420a27fa58c16b038151d78b62a5aaca77c
z1174286391d0b04b9e3d62bce30e4840d4c094f6fbac95cca9fa1be33e1ced6a4f7d5519376d43
zd7be89da0ee629cc26cca62e2fe6c9632ecc979d7eb2fe3828b9bae0d9ed2bad2e2d870305b177
ze68d504fc2c23cd56218b9430fcf84c25f63e6cc66f690b5885119f24245cc19a618ecc4848fd2
zf0d1059af789fed9bde9a9d4ebaf54fa508c0149f0883356f924036d1e93b8c7da8352936d14b9
za8c463030fe62aab7a70bd503e75584c29fa2d25b1f26768c977c637085efbc7a7d9d847903149
zda70d08c34ecd0d8773cc5ffdfd88274df5e40cce247218e54f616a3a311b252f2cbe66db7a58c
z980f1792498e9c8ae1b7f79641acd0213ba311f590218d9f609671476fff385757d69a39a14b4b
z1bdaa578cddd037cbb6bd20830422d1238daf80cc5276c08b761eadc8315760eb8779e6628f44a
zd137638f1dc78cbfafafebe98f5c321f4ad1c6ebecb2ebaeda9f0b1f9b8a5cbecb3957d9662ba0
zc9a16449b5e5f6f126fed2c4559c156578e3e3d7edd40f076200c10c2287444f98ec9747e43266
z601d0b9d5cdeb1a218950250199a4510d9ba1067299ea22580c0e5416563b509f004b7c7390f23
zbda32406515c043099798752dd41d5fc029006ba79f425e59e2aea65a4df6b973e4e9d7a4c5250
z40b6dd9b3cd692a45113177f965fa63980509835b442721cf1ba17565e0087c2741633b8587c75
z62037d4376968dc9a11482808dc1abd39121511bf1953efd93e86d3ea13ae502b8e23fb26b0a7d
z23c69d7118c45d7e3ed7af091236ec91fee8ce26c41561bde68536793c954200323c4b15a9d3b2
zf0ca4aaf14a03e1a8026519a1560d12b110ad611f99a7b495cda22cfa1976bb27dcdee7ed4bebd
z3eb920b6106dde2e84749147dc2a25ca35e01fed767008b40b093dca44493e7f52f66a2c007573
z6128ea56d6622ae2e3c558e16654bebfb6a30244e0149afe0efd661336165706fa2409cec3cb2f
z1289e6431613fa0f31edb1f642a9bd882b4371c3a00917a2444f1814f9078a8db6b92927cbf403
z2b243158975ecc3f7d42747c96698d506f440e4b90b1eb43dfba9a68ea65be6b856321da914b3c
z8c4dafc4380ff6e93b1ce237904d4b67f11f8060b67bdcd6c9496cc5989fd3f25e1c9f79f55b58
z4351d1dee4fa3a52835d03dca992af23b06117a2c160642d433169f999d3f3e766c9481eacd830
z53178df20c69cac12f0c2f697db93fdf4e7d1ec0391f47b913c351d3db55bfaab2ac092816b210
z1378dac663dda00a2f5a3cacd9f8d3e186f834cab8cb76950d7784d3665b087a26f07b806c3e4b
z5c6df6faadae7f9125f315b8f5bf7cc8fe719d226f54bc21afc21761b399bc3d794f7f8a2cc7bd
zf332df75b1a27442075f74852b8ba519d647f84cb77954f476315134a50ec0dc8ff5c3788e0111
z1cc3600012638dbd23006b306612f7635c264e49e6ac7ad4ba7bf2ac60e37fb6e99697e3f4570e
z1c4a94344ff3fb8cfaae9efaf3c1d91925759330aaef2ea951ab2596b3210a95827a28bf79bec9
zcc0aff1cc3c98fb34d0c17bacffb6300e30b0400e12f2b5dcf70f77a6666379e731cff4116965f
z77eb2216413fcd620334bd9c8dc20e921a75997e695facfd7d301664004bbcfca792ce26aa4cea
zec199bfb6c1ce459626611a595eb06de8ac0feb99365043741813de3f0026b78b8b3c5d25276c9
z4b554fb863723166794b0b63fca42f745d1dde9f072672b07fa3b9c8d4766219650615a3aaf5b9
zdbf6602bc9cee4a79fb953c6afe978848e0a5e20b78fcf3c0be6696f8eda8dcf9da3662b788603
z19b9415e74480d258254cec4898eb9c177a7b7ead1e1c06c92d435e274401c62497bcad7110b00
z1a9198207f4b952ce9d6fbf4224ee9f13072f786dcc9b23bac61726125387240fb446eacd4b085
za67fb1b7ad22fd396b70add1784a67b338d5efdcdf1b05d64d7bf03f5a4c1d21ffd241639262c0
zed7fb05f3b53777df1ad1685a1f50026274bbf591ed4fa18aa5137fb1c01f2599d06bbdbca4858
zfb49d9326b577ef847ca66cb016de2aca4ad9076b81c44324301f16faf737a96d95189fceaa8cd
zdbb986b528b0a2575efb08ef833c3682b0dd4e2b5ccdf68ea386951ad1de7ef6e8dfe664079004
zd9f44b04736159a648fafb801122417996403f537652f61ebd50927ef57576db4d39a103d8a0b4
z962b8b5d305b64a506647a6798d4963cc2f7bd247345118735d48a7e2bd64bbd6173dfa10ed1b7
z6805d1a8f2e36aa338bdd7d4f984f8fac8a311a45ac679094e26854cdc293ac7d43d92f97a1425
z8abddb60faf39aeb77e656f2a04b00ffaf3a68f685870f296d8e3c66fa3e29fcb0408402037ae2
z68e32e69b2200846e1daa68216d0129c9706efd9978aef07d0fd667fc98e57c673befd974392c8
z1c7ef1066f18163e3fcc94bdaaab1b092dc6ec4a2e900637bfb3152f7ab19095321ec8314d909d
z6f421dbed54ab06a3fed21a60716211ac6a46758ec9c92f18b1c6d1228fad0b3db0668d7e4ddd4
z9445152ab061a94c0368dff66c976931820fa9ad64936e04903712eb9de3277c842c884bda2350
ze8bee39d48ff915cec33a133bebb5624ff42bfcab04ad571ad1cb009a750f6b117dfd38f9929ff
zf9b2b12d11a6ac80397e2acca573fcb639205cc2c8f96874faff9c82a0c03e2d002b635157a149
z369b8ea3c9d50592bc3a7b154c9b59df2de58b67bc573f75d3533f92ec9f922518e0726731c7f4
z3fe1fd48dad8e25bdae7f44b09b99218854ecb8aa32e2012fb5b7bc6123ab9ee980967e932b986
z7494e7a9c549a5938e48c846b8b8caa81ec2376a2229ba3c2253350b52399bb690af84d78b7b33
zc3c380e8eae2d9cbd73c7c8516b5607a6b67dfd24ebf1a23b675e24b5d0fffa7870f920615d55f
z5adc4fde9a79c88f3f4d8ef7023674f7d26c170f69e0ba3d83808621464332ddf1d2650a28c220
z03bce04d5117901bd4fdda2143de22f6e88855e2553e2e54da854f134a9d2062cd2ff18ad6afa3
zbf073e6c5bfc2076223ea7864b7acda93d9113195d3539838ef13c00c12a3ac03500f92e90e874
z86da81f44234dc9f9571fe5533fac446e51edfa16ba57689e30a24af02aaaae9a794162f480e05
zb8db14759b6b197785c094a89323d1b5e8a90db88de4db33ad80fb460e94042cf530bc55947ddd
zd9cde3db836eab2691f5c29e5fbc8d9e27245e2606afdad8c452cb04e8c19e4727c158bcb47aaf
z684a8dce5ffd65cae4cfd7241d6b8c6d76d197dd502e2780ad86b8680fae2c9667128ff853ac8c
z26600df0c23fb1867df3345474ab5f17cc4266a3e37fdaafe22550dfb1e83c7cf2f4bef03434a2
z9a854b6a17aaea518537d4df31764e58ec3fb2cebfc6ce8c799a8f5e8bdeb7e02407207c3464df
za4045a651c3e63b8e7959ca510b2b62ff04c733693015e238a566b251ed5fed29b3245d2e9cabc
z13bbf144a48b29fffc27f68e3b0b9de2cd92ab861ef4ef0634b74f1975f398585cb592936d47a6
z29ddbcd7159d2a0253c386ef75e4d8dd56a3497513e54d6a44228586298d8aa64e8c67c23e6507
zcacf264b8028ea391465bcb6e2200d80e27f6cecd3e378df77ecb60bc7b06a346e43370b1d10f1
z7e3df3c4094cadbac7455f2b08922b7de49a94dbeafca9f5830fd767948a46c8138862363a1112
zba873b9a24dd05e5c61a4d927ed292974d1aae983cb8f409d1c7c3d6a575375de1bb709f161dbd
zbb7b07807dd4f6532b03df9fdfbfe0aeaa3e41b810b126c2cfcdcdcf23ca1a505259082b1f3d36
z3c4485168deb44c398196b81e740a01a4f0e08b5c30b67ad5a9a9829e2a6bb8d6c5327688c2234
zdc3cd2070ffbf0287b5c0ccf33dd4858d13268be5fff22ba364a02efc05bde7f658400dfada127
zb4723c696d4592d46f675a83c8c0427b65ab02c4c755515261bb09c2c2e279beb715675d1493db
zf8cc5145222c6575e8e252c3130242aa95b5b92ae3927c5915939ed3d3df7f1d4c9fcf05af1b83
z890246e6fd4a826431ce0fe805545c1012913ef41eb76d4ccabcb14a00f282ea52fdb673822a16
z67011ea62beefa99f0334c23ce641dfa2a40313c5cd8bb6e315871f12f2002b4c9007adc0b61e1
z39578348e948a845af3d0916eb0cd03ec73958465c11bd7f42e94f4f6ba9134e148cd3e47bc829
zfc00b59ad0100f95cf63033f1cc1e6851536dfdd97ae2db0fa76e2c45d3eda3115c873d3f6554a
z58d476089ba6568177328f2fd033933ee81e1263a4b28f915b2069ccba08ca2800229b30df0764
z747cdc46fb0faa531af95ab2bd781021980ac8499b8c8772c5bd322311005f55ec8f6110018012
z76dfee1f99ca178d76f4a36c27eff9ae6dff4f2c035e9786fe88161a8f6c2833ca9292d3aeefb0
zb2491fc5a2130cbd2edefb0857bddcd0e7d7da6b70b11cde6f38dd52765a3726edcbe7e8e6ac59
z200c2d6ad21a50afe833dc7b21ec7da8915ee4a738887105088b8820479f21d4f24c526e61a465
z60141ae5b798158ba53cc6e0f3196cf8c175b7b955b8cd3cf4495ce446b73d148c371d78586a91
z94d21f9178aa937e4baca679b79af68f160b5590dabda12ab3b139aecc3d15fcabd39e336bfe51
z4b0c18a06c1f0d7e6367fdbf4614378ed4f870495ad8105372ced552de519ce8d37307172dbcdc
za085cb64a3fbbd528c6a0e92df031b7b3eaef9340876d0e0ca7954eb889e2e335c462b94756d3d
zbd69ee42e80bfc5db03e3d103ceeabaa34b57415a579d567386a12c3873589607b8425f2f99999
zf85951bc98fc8a383f51e3d6942705964c7e05a368eed048f34e48a053540aa4af9d54ae7312ae
ze1b37cbfc040a6c44d88f4e825036b4ba46ebe323e8bbf096ba761c2a5c39c6eec39a5a4cdcc23
zdf8002b2e206af399a0b8f7f9b92d6d0f7d6971f1e1a7fbbfd5de4f666567d2af9f23ae4baa755
z7519e8087c01f956c60f17c71703cd037c78c101def32372acce01b63e539414b4b43a39eda16e
z4c6978b1da9fb22ffba1025536ac8e67a999ac7eaf28a55cd40c070d1ff3620307ac8616f1304b
z60acd9808697c13be164a3b6a32c60681526e32cbc556d25652d81980f1e597b2f7cca08241d2d
z210890822e88a299e3f49af3397d01e2bd5941956bd61770d8f4d68bc53471ccfd98ac0fbe218b
z725ba94345d4c91dc2b50e1a47a5b726f23522685f3163736c0fcca72ba7486596b7c605b81b09
zebe5d12eb3a29f8361f607ab4ff5ed0cad0fc15d368febf2437d703bccc4b9b17ff9d2c3ee1b02
z3625e446fd969aa61819de5089eb3317f0b3cf923c6443ea79f827a965a11c3bfba23d8c5038da
ze4c612c2db1a795701b360fe61adbc5e4a68c1ff9b199d99425909a663cfbf33f0c7f94255bafc
zb56a6955fe258c8ef6281f91877fd05eb44bddc38fcd9b2440b04c38abd829d2462568e88161ca
zb47b4d08e1b24c77f7cf0b7c6043762756f4418f342efe6c7d5a78494dc1b71a698e904bfdc497
z04dc1b2f3a65a09d368d35bb1596717554b550f17aa844c38beee3dd6494b227a16160604c1b33
z6d6e734784799f4ea5db6de485e17db32771787cfb7fe9e86f4155471f628e5e487c3b985b8258
zb10a7c1e4939e88c7c75ef183772c316db461d8a60cb7b078ba5d29ede91ae3660186dab6e98d0
za13e7b7830efbd04709a88a8b44f3a4fa552f2fd78bfb9cd17a613aa0c8447e37b6e3dbde815c2
z160baa9542626d866c289c16142424e807e7600f6088b2b808de4120fa7b5d0d4b05db374a4741
za762ff53f5aafb55075d5d7d1d15cdc19dde3d8d9894004f83642ebf1534df982c751b1131b087
z6149d27060972f8799dc4890d1533cfa8cf5e846ef404485c8236286ab00ba541e0eccee595aa4
z8e0f3bafdcc3d3d75da32f2a45bc80509450b8a3975294e6b00096aa0f26e8bb006d7705205498
zd27b3dec5b4c546e74406f1aaaaa54b53295d086272523be25c8de1f05c8bfc579abd9b98f25b8
z0da5419f9f43517626a24815d3578f8fdf15ee55a9841db98aebe4e0631b23c393d7afe120ac90
z4daec65e70035d3d4ee6f931da653d0bcbc07f833973c36427a3f22790c00790f9718fc26344dc
z0a384920cb3da2be291cb31f8f524aaf1805bf3a327f3932da65745461ff546b3355358b9f240b
zd8971166d12484187aa63c77497563269385ebd7af6ddbac505528c838bc06c9bc46caffb914d8
zd8183bc62c525b9711bc7b75452523200dea1ae462417554414240ef1f0504548739163391b166
z0c0b55e66d409300067b45b14588e7dde55d3ac19044ad169d773b3fd6d16d205e31158380a6ee
z66caa2ad4875afcf7e8b7f844347c88ee64c28fc04bfbdd4a50bf4e046f15b07e4886ac8df89bc
z038d74df7ea147a9d53b2865cfe3efe69d738e6f5ad6c1b5e829a3510a9409d5ae927a169a6095
za5aa81acbe5ca6e5523abf07a439dfbf614b1d213759b2abd5f12c2f7b0da3715a22f84ad3a540
z51034588958371c6dd7035dc52bb5b6ad9065c86e2d14da27b2ac7968692f8a45a0814c58f650d
z767d2fb94b18013f16a77dbc80ae122af59d1f629bc08d25fc83f5b684f3b5c51d2773525ad7cb
z21972f11fe32dadf6d69ee1fe7bc62e30b015f0bce9402f0f9cc6efee891cf09e78a3d2ded175e
z1f3e0c9a59885dfb5927e52f6e88686ba18128e1ba6fe77d979f8841d566b2ec0037eb9af528b0
zea3a843249221a6b4d0109b708d2eeb293a88296ef11df9f3e355ba90eec865a7f8c87f03ab0f8
zeae570f4d029d3498addc1da0df7e69eef3e011a2256fe19c04bfe20a6249cd39870d70ef678a0
z03ed66259cba21d59add73b71218e9d5f47f807c68960b3bc599959bbfa2694738e0de7a8a2003
z378bb5fcc2cf0d9a706f0ae59040519e3293a66b496a617ebc15278221feb2ab93032fd5a874ee
zc84e85a7de47b7563277e93ebc9dc13d709e8592fbb146f54e1597156556969a8c49e01479f1a9
zfaed32fa796c7e363bf4385872e02591d9cba29a8d942be014f66cb80c91d832c0918538bd3155
zb1de400932908f032a006e00ef20c445a5dd855d70e41a3349f562368fb59bc4a9ed83e08bb946
zac1d0e955c07d9d36aba6018cab4b5d7858596ef65599b6323620b9da82368a129507296a1e151
z079c26bc3c51970ab975cbad0f582bc21033878cc22fe6f222c886a594f4e217e609f734cbe250
z4706a2352f7dabc39f024872a12b90efc3ca906069bec4b974e52eaca53ba2e49791ef2653fc70
z3104bc30877d26fe88f508e91b54ae0a301d5f2951bff6afe138ad7fb27d1b5fca2fbaa1b76483
z030b20e42883e45ca6223d1df7b087b2f2188d157317e3e2cc88ad74eafc648b771db826f86b00
zb8dc1752f7b0738b54ff6ef70c5389079db67be1420e320f00e9dba09346ff3bccdf921de209a6
z0a25a5c09c774ad317920f0cf3b9d367c7bc444d5d8e61a6bb96a4b68ecf010aa15336b2822e3c
z09eac7b9a6bd4e99a29518fc9ae0b44df78d5b7b86396fe771f6f0697e3326167d7f862126062b
z26d2f80bd654c47af0541d039974e538f9c7c72c9d7557f7a8c55613702aec8c9ebc8d59faef17
ze491c17f46ca39ba3aa179b3862bbf51e40e84e753ca6bd7f67d10ec0bc29cb4d3ebe5a0727661
z24e480590cf0419e31fab09706477f9ed5f47700dad986e69625e5cdae0799d153e2da1ff85f22
z8077384ac5d579c2df97f76e587743929e8c92d1010b145144fbdc4b7afbf361e4d6192367ddbb
zad4cc96a0be6585df269ffa97fd8fe06ded695adbc792a53b20e8ff10bd747872d97ecdcb47e56
z1f058aa8ddfc650a0c78a2c65e0f7242d5e39f9b2ec4a2c1b43272f5b054a086a5a06f61cadeb0
zd02398dab6c2c1f12d55780f11d4a84eac3572ff35b288d8c8a9a6343d92b2c63a0be19e4e387a
za49ed48fa05bf326385a4cbb1af3dc4dbcb155feae8bda071b3902f82cd5582505794357059ee5
z376415204b06acad4a067864f2ff33d8ab1b29c815470a807e5dc7b27b9ad4199b88404cdf3ef0
z5feb4d7545038cee655289f750caadaa6368087843e3be5b6310cf54ad1552e978cdf97285af31
z3727e7f33fc864691aea601ad5d7a0c2a04b1f085592ec6b0bf1649e56e1481423f473efc2a599
zf981dc6d60d8a2aaec52860c0a9d19044f5d434421a33815ea1ccbbcf9222a0a99b6ba8fa1ef71
zf217078fcf0db8fa86e87b2cc88b929b9250e5500d3927739bff7245574ab8be0765b8775e2fa4
za21fbd7ade84b147567ef28bf174fe6c247b34b8be2651ded7b6631caec04285a8e987c665e300
ze4a8585f2e515cbe34b01e786a0c0d54e34abf20e36b82af15d135c88ea0574de87b952f833bad
zff0a41b630b0854748500d27278d9198ee7d4e6ec79eb3e244eaf2249872b5fa60cbd8917b7b63
z4728fc6374cc415945676e5b6a1d681dc4b09fdbb1e3ba9f1abe80a7c985c6d03b028eb5bf1dfd
z0816dfb4cb92154d4587c390385bd61b91140b660b5e91bceca5c9119509b8fe772c3c7559dcb4
z93fda3f1d2f1aaaae4f43b335532dae2cde094d21552d1351c3f6579b4058f3d5691dae5844fef
z90756ffc7ae3a5d083f7d8d84bb8e38b511a4d5c376677fadef9ca977971ccd889638d63ff8031
zf8c9963bce3677fa576ef455cd6290ff1d1e418b4a525df1690b075dd9d54ed9eb97792d4e579e
z1f4f3e3c66daf7c4fd38dadba42c2af8c5159f884ad48f8782b3e368f8c334b85a690851735f03
zf1d15d8141681607714a544115025f484b86c1024d3ca325ab1cdeab8771075540e5d5621aceb6
z452b6be70af52563e5c94b74dc7d7b3565c81eb85c753fb570132e109baafc5f825bf2d7a76e1c
z413f1430ca2bf1ab6316cbbe6ea3852b451b3bef2b3099d9afc5aa148b23347ebb85eebf0e30f1
zea18837f4e5e244eebf4500e2a80fde68b4a103a7f6698c1122c2f6c02d8fbed586c13a2bae79c
z776e06d92d92924c6c07fb1254419b3633efee14d8c9c7e16feb498fae2dfeeed30084e75feaf3
z476a7e3297654c57a4920be797412ecbcb3844f76c0a33ee69e05658102a5186134138ac7323df
zf34ea61af03e0206286d819e4ccb1d6bedfe17e9b251e58fcdc648e62d2055a459e0c96624be95
z65d5ffb3f4fb777cac83a049746e82fe2f87c527fb0634edfaa1726c5889e1c330e59162eddbc1
z272d13532e22cf03e26dd6013b4004ae0d5a326170cbf17347c34e68e942b7577c1fb7ad8f461f
z0da41d199d7b0daea4b72831a7b5aeb7fa39bbecd7e3480aef720fd7cc759df2753cdd259ed75c
z026d9a76219a4cbabca466b591d8fbde7a648adc26ff459823bfdf13dd48b72810bd1616b0a251
zc3c0dc1afe2d0e813e342f7ef274cdba11e7993367a205387a34bdff99a6c1df4c0290e12e399a
za961ed16e186af652a6cda6a80c8b67d3cf461a4900d5355e4fb2fd100daef0b9b77a08e408c5a
z7ac8a6328b2e656452d811a9e6dd823cf5aa0a19b12792b51853c5017247134cc4ceb3fe16b04b
ze8685fcc0c580bd12b7d0311758ba13171ee86d174a8e02eb1071c45a7480d9381740044128d4d
z53d378ed2c0cbdf520b692b95a9de529faad41cdfaa41dbdb85549b57d0ac2831b3565335c4852
z487456a9e0e61bbecc8627fe66f82c262b4f8df7d91e7f4663a54bb6b8b2e063b1156ff553d4bf
z9bb0b082129c907071af76f14f831cb17f616f8c6079bb7ec24b83bbd7203d36ada547c0472e9c
z7c8216fb1532fbfa1635856e7209ec7911579db0c1da7861ca8f75132d43e0ab687d819386b889
z92a7db76c95830f3b8097d61feea1368e06755793f999de9a95e2b35693b643c96df64d9cc4418
zf6b4aea1d70622a9facf2169d1ea2438421a76817926682a29efae0d7c2d1472d85dce34422037
z5343c5ac65a315088d35eef0f93ef184868d7a8cc7768dbe53e2b0e7cf04c6291dd9df49b89de3
z9eb43edd49b24b63a9990947e82e0f88716571a7f76fb213ecc7837c07a866b345343caf3b03ae
z06c0a2ca61c2c2390dc06f722c27aee58d6c33ef290f43db3bf3eb6693d895ae964cf2b31e93d1
zac208c8fb36a4300504d5489b301773cf8eeca1b4038ea5c04e5ec61826de880591feaf883dd45
z22048dce90fca790eeeee25fb1ef3d13270d996c6a8ea2d278ecf57f0b85f2d60802aa50a70377
zfb5531f1231f4262ae46fb1363d31c33e41ff48b7166f38d9d3de952b554fc839aa220cd30b2b9
z5838138c3b3ec9cc6df7315a2388fa333bd207a2557a7c4871fedcb99a49de85f51353e09ee190
zb803e09f44498cff8c238fa92ba5d9fc9723d87db5c5822ea4a20d49cb05417d1dd89f80d9b62d
zad465a1aec58b4364032ea64eb2f0fd6827fc9fffd32e0ff2fcdb50d2f0495663faefb056c9a34
z8100ea800d86b2aef09e18b2f2007e552f6d4f7947a568e7ae980c4930e69e38037dcf57a9f38b
z1db74814f9ec7317d4edc4fe547f55990700dcd0aa20618ffc117f4f0a901d4af7ba17b417ed45
zaf26746be2ee6f4722c34f22e0a022d1807d373b05ca50dc7c332f4f04916b1e9d00f81b4804f5
zc950805c5c30d2dbaf642111e94e958469476e9deeeeca90b081778146f6da51a29e10c9a7fedf
z51809b49b36c542af2837065814d1814ec7b4e5a517ea0460b6d22f4fd67cb0a8d91ed41795935
zaf189de8c2bcceb7099e8a554cd092ebfbd1f0016a7a486039d7bc1735aa3c928de6df181a5d64
z381edfff309a54bd08585f0307decdbca06a673b1a5d963b3cb16bfe96c7fef5496c2809536015
za4dda0e76fe2b85e3cf4fa82ded8694658454f3cf172c16d0dc16e1d4be106a0b0e3472e71e15e
z2a8c98c3d0f0f3fa3aae952646575f1cd18e49f31bf44dd3af1d03467c867302a1368f64408ae1
za1f7fe37c9d2b47a5ada7e07ea318501318a12e3b7bc9ccc6fe2db721e0cc6ea6bcee9cc7b0e08
z2339bae29c0df25c0ae8afa1a8eedc5422f8094b3d9d79099467ebfa21633bb693822642cdcc9d
zc55cbd95837184291e0e4198e0cb981a58037920c1676b4d455c357a2d2b11fbd163d2c63df8c6
zab9f805516398d7d7034aa5bda15e208f7ff4eddd53917c4aa002208cff0bf12392c5e120e3f85
zfea4180a4a28ff784f9769e35a900e0cbc121b8b5c4e076e0032480f4a1c6e356a0750d7bb4823
zb2a56eb8836baeb42b360feba286625ef18ffb925d47395c6b873c51de78348269cc1551f109f1
z9cae386a5b19302cf82fda32d75315b1fa06fd663bcd219e1fb91d5b8fb68a8d0d415add400fbe
zb0ed4197fa86402ae92ca208a55b387b6bc50d3831de5e870bac81dad6c58086ed37baeb9f8684
z33682949df24593dd404f2d734531a5296341617b6926cd1011e0ed8c87e7f3f43b3dd5fec169f
z1bbeb12043e599e496592a38c1926464ec93ec8fc10ee668958d04ae4e1d4c5acca85f38a62b37
zc88d7777b1c0a4d375159b168194c2bc023a4887037755e7823e91c9584890e97a6446fdbb5be8
zc5f7d0b8085149e5a738f091fff764bd48a28a78cde737bc6be8ede7fed9714f8d22ea5d249bd1
zfb1a3e76c4b38a88f96dbfb9349e0f57b223201ee4fc9ca518600b3bfb81b8aaac1a45d61655d7
z8c6a30306da94206204d42ac28746224a2e9fcda538ad9bedd34c86493a782b799b1db7d8eff2c
z1955bbdd939f4fad70d3d1b131756f53206f293be26ebc3c1becf3be88dba61bca4ad30d9db78e
z0d031d8c1966b66b9294b9499e42cc5e269706645665df67744ae6c1fda7d8044c5c28356fcaff
z7cc6486825c94372ff102e6ea74694e751348429a1cd5e999357b3b6c85e0cdc948b7251ea8421
zd5df6c3fad20fad33c7dcd5544b315e90ea0321b0cc0d3097478fb7209b0482f949135c6e5cd55
z06e7a4ae701faa60af390fd8bcfaea59ec0417185bab86a1dbcd3cdcec4d5cfcf6df418669ca7d
z93e56ae02e7ae407f6d228a5482b88ad7b115a8f498c1b49c647e1b6a579a57c1fbaa01bcad7a5
z080ed5f56a37da2dd842867dba921d60eef7df0a4224c68f076f2027ad5d9e1cfe4c9f08e9a3eb
zac1b568f3fa2e0060f1663d64028ea65d8ea29a17f45704d6fb2eca2ede78daaadcd2746e198a2
z30496fdaf093b998d6b7967f78f9bc7ef01fdc63a9d1637d810a31f3a056599005c45832afea8c
zd0310e337fa2bc177dee2f6336275b63ba5e0aa451c292b246a07832e8e8d0d99dbca9936847ba
za28735417ba6fab8c67828ed2eb1ac83d5a78122bb86b5631b085a75088ccbdddcc683d0ac6e17
zdaeb03112e6570e6d463f4239d5115a6a30eb718c37a463d9dbbf1b849577787f70aa35834c183
z8c21ece566d31350aecdf9b04ad774fbb5b37f9cb0b16447fe426770b450dd6f98d9cefabfc781
zc791c501bb50205a51df54e346c6144c669649781b3d2d568831bfdf88af02397806ede0193031
z60d1f08901e0b1aad5ebb4967407026fd1b6f037fe8e860883f185694dd7bfe8aef4c64a9c48c1
z2a58f078a831daa6918b048c0040b82738b237a9a04ed7a3baf34c7fd63217195edc0a63652153
zb76c53651cc6a23d996a7620e8d6e756d0a02bad01d8114ee68ed9942f381e3fb523f578d9f1cb
z4f59a83f5f670e5051bde6b2dc3281776473585462021aa5a555f7cb8854daef9faf49865c16da
z1b76c56fe89f5d3dbd85584b30e5a14b989d475a5d182c596b5b4d81c7a55154d17e4d9a0d4918
z79f202ccbe5e1319da04796c73d4da193bfe39c709486dab08f104bbdef3fe18c834bb554ca190
z2c81ee33c09d914daf84a121c22ff0f2a5824bd1ade9dbe6c3e6afdcb0e4cbcdd7b8910477f530
z9932d91995c1ff6c579007f59c667900b12da57d1c32fcad15c64e20773f9982402ce7af51be51
z183556e303f7a614a86c41b2c20d1f0b961d02baf00ccfaae64f0270244e89950cb084581e3395
z99c6ef19c14eb720e71060928841ad748be9272e75f99a658cd4ee9489a43b536d5a6bc6fb244c
z099e0e4ce626c973ef49cfcad7225aa4535e40c1cde54edb645220e337de1bf69c544600d47d18
z70201bb1ac42e57cb065f6ec9d29662ce5a67da2d9d353f865ae122b5ce99069441a71779403f3
z8d247c9683dce138305dd1c4a86f48f1c31576efa34b1df12b62a7a7aae4dc06493ee569e3f6f1
zb2151e4116aed1bf8d262e49e7a0355ed6c0d5f0a409b6f5b0edcebd23adcc22fb56175dcd8d6b
zd24acd3feb3de7603b1a9c437613adb85aafdb0ab77ae316a381bf82e120633e215504c70d4341
z090bce99f998223981ce6af3af9229f011f105bdca4dee7701204c9721f2d34eaa893f2cee410d
z484f66de5fca56a07867df24877d0ac745240ec51402066b78143608c5beefa6aa6c2c2ad5ce5f
z131ab6c24c37d947bb654fa90007663228a0645d4b6f59050afa13e91602f5eddaf81eff6b8844
z4ca1c4f9645c17a4cf8f9ecd6768a9af374bc60660550fa2b05d1002042cc10850c5e7f9926e8f
z7ceef1d98e5deddf4f56f70d1ccd528a03a8fc9d1fe8bb2831598719e37a54c810df9ede2d5c28
za2b13639cd5205b8c591d54646fb2b001cbdf9a0b41dbc09b65044ce0dd8a86b467a3f13567e8e
z252841085f5b277f763a1d24930e47a4439b21be8c1876788f1bc5ba5b01e344367a0be2004d32
zbb1253e8a86613400b5f3c61b9baa5369c274be8fb10b7c7d0f06011e6ba85357b3c5b7a6f799b
za87356624f62cfdc5d606475fad389c44d93059594d97b7231f5a2e0424e2db5618d71bdf60d3b
z5025d5c5744e25644f1087e60b5f71b8fc4529f6546e88426a29fb758ca4d6378a0ff6e928356b
z9a59d3a0b98809ca74136ff98560cc18cb70b63ff82cd3d9e44e5bd1b7e77a1441e84c75727708
za1de11a9f6b9793b9d1f6b3791752f10c0dcfe6ac43e9662dff2d22bddc24fb3cbafb15cb6ff35
z557e55de21210479fec223f287dfeff9ef98f2fb289160f1792e67d6208d8f141060a34119a3a2
z0cb4b8464d0b4944346871ff1dbc0e18ef5218102c4230ef8bb40a0a4014629056ea0df51c5433
z7b814bcaa443c483e61b45a14b386e32e41215d3e0c83965fdb9b30bc8bd4d0208711bb9e75f79
zf528246b01baac50385cb87dbce926d386273cb9c1124c7b575611917a439d4274a7c24b0b79db
zaa54f7b52f979df2574d9ed21b94d6924aadaa4cfa478d12cdaa53d2de8ccd1c0bd0ada0bf762e
z4b62f6dbe12f4dd40c63548399010d4d64d26b251ce1c95f86d2eef78ddbc4eb0367fc23bc8676
zdd77fc81c38002d2c90e1914e3f637cdd2038f187f4809d2a3aa7611de1c8a422bd8fbe5074477
zd313dbd2bd98cdf260741973d9eec170baccef8a3ae1ddf96ffe469df34522080dbf7237b76e3d
z55aa3499321e95084ead281202b12a11584d216c6e648a990a70b1b3e243ac49b694c4dde521eb
z7916f4c6591b4df4653a3c4e72f6d171f0a70123d95fb2b498a1dec60eb64bce9d82afbb88c4ac
z0c1727482b96ea940eccf11b608343ea065a6546e53a915bb00b44d0b5adc7cbc31241e8484483
z0b0b165ccbb2c512f6c2771a957003937a3f3219daca9ee0b942deddb3d257ff825e8059264f8d
zbf2aead4719e5066a692129fdc40f5be2c01242501ff789ff74c75d8ad0391a727ba1243f9904c
z1a482910f38b3df4257bda43aade0f57e6f990cfd00847376320f8ee26e13eaeee1c0446136288
z728ae516607e54730f070bf5b9ef9fd71a5039fddfe1eb0a7278cfb3b920ae47d5fd1e532f59ba
z873151af4149b8f3a4aff166c0979f9e27ee9d5eb00aa6c59060f5583c9a72d5633d37dc77aee2
z8b4a47de554b963d8c04d45ff1629c494116b2e975e8297f1c01164c4c78f3f2a5e50ea282c85f
z8940ef75bbe6b2d2b19dd2c2934ba143e6a65988a0116ac3e17e5c21709028f19cd5d4ab760d96
zfe67c8ee4a189a3c1721ae8ddfb18a57c49aed8d05175ec57779d76bf98a40cd6c475d669de12a
z979f9ae17489e4df93579c96ca913e6710e1ccfc9cd2f87891b4e41e9d09e9d3bb1ae81aa45cc8
z7d10cb58dd291c37eed03c7827d316aea49f38f3f95f4ccd92532cbf86fb5d5afd64b29b9ee7cf
z592aefe935152b2d97ea69f82afdad05fc2a9668896fef29ab8f350eb1a8c06c741b107e222569
z0553e44bb9ebe7f101c7f54c94d18e04f4218000ccd58e4d8109bd6ffde08bf8866c0bb493058c
zc75a3e8a83ff1fe27afbf600a9dd85870a74cacc2adace1c9a6a019594e08eed28ae29031530ac
zd891547dcae59855e261e7231c1a31e9d24c29e9a6938da3e88dcd4627783f83a9dabbae38bdd5
zc7d02c99621422f4dff2f3e9244f8344532b6715b52a16c36c39e3773b2942da657a6c0d9f1ca9
zbefdae4f2100e98b109d840c2b28193f9ed1cd2e178b35158d3b6f168da29eff9895056fc240b4
za4412fcb3337be3133522a8464cd619ecf90da78a485130d1cb7ff772d997280b94e26d28e0f6c
zb3e31edd50934a5dc84741d21f167373e2cacc028b86f643e9ddedb7c4c65e8faccbdd07ea73fb
z8a92445a71147eca8633923751f4215197560eb2e6cb5ccb0ab1a878c34422deb382c57a4ae974
zfcbbbb8fa5e739a907e47cd1d1e82f6b3d9859895f3483a5f032930a1b3558e906fa1e954d9460
zcfd1269b5e58e68ce4be8ca43ad5fb5dbe79b3050db3757b50898cfdacb4ed594fcc0fd64ecabe
zdca6be9c50921e72d7fa39ec76c5606c1fd5dfb773d8a147ce72ecd131d72576796e4d6fefe6ff
ze54e43ff52cc7047a46e0c2518d5d51dd23fa0f7b45c4f6102d870a5adf608878a0882a84d19bf
z2298b0d971b61234cd6c64c7d6fabeff631adf3516397f4fba3096166e16e88abc0899aa5f3521
z4aadae8e210eb35c3dd10440d5131e743794db67d25b09879ef5e73bf254cbf27cd92a080f8a4e
z17181ca8e8343688e5543eaed1a65dc0039631d933f2ad519643fde10d8107b51478198d8e045c
zec104bc48e67a839a629becd3b34419fa42d4c9c770ff71663aa0c1c10c579277e1efc0be4ce09
zb5b033f2b10203aba83a2786f045a02a37dfa4fda14f54d83e95bf47f44ca225b175ec643b13e8
z33b552b58b5bd334a8162cf3cab74af291f555858e96eaac50b0f661705d9b19b71453f168213b
z51d0b389e47ade120db551b2f50feac42d373f785d5aa558e5a9f90ff127f100f82051a4821367
zadb4b6bf15c2338b036eaf554f52a28ff69a93c09095b0925ace58c7bbececd00210e4e7dd8d6c
z66e33e7a2fc2d4bb193e3f644e7c4a14f30ca8cdb960be260bdcc0c238416bcfb807f289c01072
z5ffb297f0e6e6e31523aa86375cd14c00dfc6854d04e9ab5b4e59ce84f1876a5cf9df4e93803d8
zca88308100ea4d1e45cceab246a85eb06b2ca7086963133ff6a08bc78e385914ae9562a32f8fdb
za2c9e97739c1767f2700f09289151d5a9cfb24eff8c42f3b2864094c2874956bfb4a6ad9f1856b
z240e2e226e87cf7056c007c7215933de4649402f549b5015593f79d5c0bba285db4ba9bbd5b2a7
z8f8930f019a20f119611a619bf8fce12a373052dda0f5ad44ed6edb2db74db0ff00f8d98b6bd58
z9ee67a90549c5dda12f60ccc7000a52498b4dcba8271241531dc6814a19ba3728f1ac2d5a2a263
z9561df50e551e893a5be304b715e9b1943e351339d566259e48323da10946130629e0d00fb2e3b
zeda1cdcd80ebc9f966fe95bb610808b479c730b3f53294595866c288821a27a201b4144811d61e
z95d0e106a63e706acdc8f04545d5cab7e73ff74e4089ca5ff732348cd7d1fe18bd7e064354067c
z4ae94c4029c51a90b9e8c09cb23eb8ef772d7d78cc23d35185464363c12cd9ab738a94b82f95c7
zafc245db9f6ddfcec1a39d4e3bf9bb096b4332ab4eb1f7cbcf7a24de9c627ad2c92a4c7e8d2b29
z36004d36327b91e12393b3447ef61df68f75ae1ccb159356da4903d9ed63ea1af8ca2b2cc5f2b1
z13912fa940701d786b1cb9ecf12c0fa4959bb2b3ed6f749c263ef721a499304d809bcfff4f1519
z70ce764bc7cddb465b486604a346a5ab36c6329cc63f7aec5d34d3a877f36ca09042ec04828965
za7923bacc09cfbac058dbb6def25b812471adf398fedb9129656fc810b86f7e9a9d78759618eb6
z5e7fa93d8275714cd7587334ffe0c1596b23dbe6badd2e3145fbdb5282e0624b1d2a080af28d7a
z006c8bc02c543db4fbbf1da5b5106e07ada8824dbf605109eb45c9b524c002bacbc326a7ce0f89
ze6badfa5fd1885496d941f642501145d7b50af23b6b35f9bc20660f2093ad8d069afad1af7d71c
z86d5afe4c8fb5170284cdcf960f33cdbebf988302ae156087789c5bf8d04850948d9e17b858c61
ze026e1ed764cffc59a69eb4423fc63650f0e88bda4c167d27e62a2892a1cc74dc0054be7d3511a
z09898dff6de44aaa03a4f13c828d1de88a83e65ff1c4628373bcc332ca7525f9cc14b0ed4fe96c
z1bba30061a0bf151fa765963c19b6e889f8928dc1cfad74b5a642955d7593afb1b7fb660500446
z4727b67fefd4755420c5817afecc31153fee3cc5135ddb54b97abdfcda6fd84e680b24930eca01
zb42b24e6ee66173e6bfb9c7c22357ede8478a5ed62faffa742a30bed0ddcdece16b90bbde204c2
ze4e6195463d8ca2562cc6b237375aa0abd3d1fd77de86b69941ed200e345da4e768b0fc338bd11
zd5c7f088092d4295451e38a36421b53a8d04b552d99611fba5256f302a52345bc9ea12d0b2fce1
z0e16e1465fd03ffc8dcf615654dbfcf1d2b94a3085cb785d650b462a9a54043e0fa7378246252d
z573aee61034305e5885bef40f5a3505edd8e0efb46aeeb9f49ae7401853ecf2a507987dda02572
z3078f4836505ad472ad60db9fdcf3d92f5836768bbe26649a3378274a0451da2c08932cd67c9f2
z68546a825e95480493836b9b97fa53c1f79257705f1e6fe160d4694e0dbe3f5e25d408cf01ca1f
z4ef905be0b860f0004f27a92025f2c39e076bafac3a9fe0823f45c26920a8e80ae71e08bf98161
za5a19d93906bace571a902dbbf8e22bf4bdb000d7b0fa62239bc43ad571ca6bac41d5a5ddf7d75
zd009335881c58a80c862d63b0360809af020e4ed8f6e732c2823b0fe9fbd48e704f2575e72e902
zcc3e4bea83610deedaa7ddfdae19532d83222a0745e5d810d5ff10451ee6f20213e30f5e2139db
z2da982f63dd481147c0b0718af236d10da4bcd69010ed0371a9cf03c48d9e17b9771436a6c1d5c
z4e85a7c0568f6298c45cf94a5e28490a09e7abb2bcd7d0ae527a0f987c8fbcd0b92dc004310163
zbbc5823631b3fdc9f0598303c8abf150a89e3600ac2ae4d78c50aaa48d7615526ca2aed8d2f6e8
z44a42fc98765842a3394e6462d550de662d5740335bd072050448fb8c53fc531596c0696d26190
zeb2af1d5b4e686d03a7c82c526545d30e4818dc11e4aa126c7baa720dcf26030432fd106d244bd
z17fe20a3243e126d91fc1b2d7d31defffc859dc53c16ff1a570149daa7031781dda19dd1cec833
z8f99947d9d33f95ef5efb41a60dc2113a2031e40b24677ed2c8679b1093bd8f08dd8f0df20ec23
z5d200eff076fc1445b8107720eb00074474c8379e3fe050dfee119f6b8b1e5964adef2bbffffc4
zcf645a2f07f8d9031ee6210597434bac387204b21bb4303104a19670837b0ba37b08fd12d0543e
z3559417e082ea3dae809443a7347ce886affe23191a5e937d6142552e9835902cc4271b4ac5f3a
z64ac3c3c0484fda42ae3c82008b15dc8137c4af2ffe4bf9a83df17322c7c6d41d224e43d00c61f
z79ce17332f59da5507bfef0d77c3263fd4387e16bdaee8555654e790e0deb0e538f5d812c38aab
zff5105bdaef4dfd978308528ac82129350e962865e5a784ea9f3f32ab3aca5c75a52c42c19e567
z776a8830146f8860a5ff7ac543280351f55535927bbb070224c13081bc012141f7e23df10866be
zad0a88be0994c0e7b6b5a40397e93798417479d1eee6b356edce2a8575b30e74f040338b050b31
zed4a23ddf5f367f880c59de3bc3f52f8d995802f630652dd27763c77188ed8ce189a2496435ce2
zfe0b845108ee34b8020f7792bdf91c448a898083071050471d776a6c48213fd09b30807f7bf2cc
zbc83a344ec28dc59bb6a335f23e06fb687588ecde5e8d3f6a5e4cae5646db68d7e023c86728d8f
z70662b0c2d3d9ad3eb6a641605b175613792817e6d9848dccba2a2e44e4332a33c8a2eae0686e9
z737f949d40ff9496c051a8f961ff446cb0ec1e69989a9d60d2113b3f9a8890e4809cc78e61f144
z77984882b29394b3c6d69a3c4a6b3cc99382d67e65ec3a8d71613f014722a0e83b44d800596ca5
z2b39a07155280bc85bdc1222fc4d670e5763ad6e56b3cea28207b6d7b8383268757bce6def58b5
z5844cff93ec47b9f7a4ea4e69b31b047bf72dabf19ffc57e3febc8144766d606981d429f43d698
z139b7f9544768c82fe54afb7dac54e3b56e5c7207cb51b1c4a4f2f5ffed817f687a2c1aa34902f
z3029c24c29d873e2cff0f25e76d561d514f193b81e459942fbf5d99bbdf869256a8fe1860f80ae
z8b4e5b4fb727ddee1316a6135fd77cd2a638df5686ecedc521c88793e9fc4a2fdb308fe2f8a4cb
z6b4fb5db50a3435d7ba54892929680cfdc77e43f86ec84ea6f83f27e2593665f41e22211aeb29a
zc2f3945545a294d386c548b4383a2bdf43d7dfac94841f9ef1faf63974f3e268db0fe772a87d8f
z962b5ec084948e9743f703cb592d201da947a3afd810f870a9a62ca218c219d999360b503175f8
z0621912b49c4f8b49ff0cb05e7f3b9e530c422f3f9d9a7b64bb371eeb05be927b263f9ab8ae8d3
z4ac215d419caf8b3e7e46ea63d1e6c0efe45694d41e9690d2a79fea11bc8760a2c555abf2ab08f
zb20ed9a22822a4c7c2568df79d95d73fd1da4526b73afcfc8c90b3717157bffb3d07b59b913013
z958dd0179e30ed3a872304692874f1fc77fc446de6f0382be435a3bc4630f62c29a0cb4e7cd31a
z9ea7fc68b7e9036b7f186134b42fa1a48b9c23b060162153c176ac2f7826e8decb07471013fbee
z61f2f2f5868628bcbad9951787be5d354316131252ca2df29c44239e84ef020df32be940ac111d
z6627da23a8bfb1c961a87f71423bd7fd880179b56a0315335a80533220d8f4a4af3da1b0ae73bb
z505247576b41bdb1f37b65a8c00f21751b3990a9599afdb0987d136755730d6758dea71964a6fd
z95234d6f22462bd12741d9a9aadf70146d48abd66c0f194c25ac9eec44e3a3dd24f42d55c1d36e
z8ecd701fc406c776cf2de174a7b4b6b3a07c32802e9ad29b96af0343c472bc161e93e11f1adc2e
z62499c171273041b9ca64dde806e9a7a889be68801fe974c17a94e1cb146ccbc65a2cc93bbc9cd
zbe36694d5e8bfb45dacef47411de871ab1b44310f364da0639356ee361a2c28d9c0f44ac813bc1
za7147db5d3971ca0140e3e56ed97a19947f1ab827b99c9f16374a7bff70ee5ba96b3c960f6a76d
za067b105de4616ebd557f4ebab568201a8f90fe17b539808b53a9ab9f76758ca88b1cc6fcf3dc3
zc6249be09337a567503aa5959c6d408b4ebdc32e9996b837a65130203d33f4cc2e17617548c114
z569f6a10555d0169e398a8171d81eb6ee1adb49a61938a7e79596dd73b245a797673db8bcf4b49
zc16294559402658fae8c21b795d7555e524ed9d1556a06386ed671af9fe0f09ec0921f31efd522
z94b3812e84a8f0ce3a442a7ef214167282f5cc389036a3c2178b2d757c296d46dcfcd45aade5c0
zd889a8fecb7eaecfa986fa2fa932e581f814ce9dc774eaebd1bbd8f00d08a1ecf8d9c2e9fe89f9
zbe0b63fba828454cb3ac4b6ad7d7053eeb8ec9fa0a47c22abd3148a493029bff3acf07192f49b1
z63dae2d1a474177fef2b834f85c0f776d43873eab70c274be466bc88a34dfb832c39c16169d6ff
z0b03f28b4371dbaca53b4e31fb5389bebfc5b683231c37c8e692213558491c98fc0be62e37f0cd
z655fc620df8fc6174ce578b606c49c3421e94187fc4b5019e23d4682ea7a8bbd2471870c3c5716
zc219a2375f93079fd05c0136f1989bbdba20c2414c7c1e3c67243da284f43bce6702788d1b7e08
z967be16ba69a9db6e59e6b556e4bb44ad910244037c9eb6a34ea271257e3a7b8719a48106022f4
z05c271604bb757977e51dea5c3fb17b6531cb16564b20e4e0bacdda4ebaa791e40aa99ca972554
ze1000237ba9b1b5c40b578f7fa99f497391e0e8f8781326fe267dfa545f93ec030262aac8da444
z78a640d7bd5f48943e7302a596e61eb6e6082d1e44c55c28f758caa19f676133075059f021d011
z7d19c436539825d290799a7bbf960f2474a7aa308545d8d89d056e2d276630fc337f9ffc9c5dc3
zb1fc347efa6dfbceb9c7cef73991b1e978ad5dbe5439860f7cddf7cfbc3a33a1c372dccd054940
zba5d249320786af1b5bc41d4ea77085e0a437707b035b0f473dfd92e5750b3d3a1a1ed49788f56
z1ec683a0fcfbb908299a0e4eedd7b18ba224bfc35e3ef5c80e30c8bfbe6cbb21fd076cf66c568f
z36c612a3cd3f6c42bea9fed1df83eb7c11b8564548686b189b6ce0c149eb5cd2c03a9afae05508
zeb7b108109578bf19a2ea2a9281821bfb0648914aa3f6b3a7d3dd35f94168ecaf76ee082c0c170
zc767f1d3224b2c04a9e942db1771a88af7801b33202b129868da9614dc6c62de7fba3b64c902b9
zd62bd14b3fba1ad8f95fc326ccf9177689f73e98a8c612967d6316ebaa93615a306840c4ab181b
zfffa5f5f1d0fc39b0311d3e8fc0624982e185ce4c525093f63edf91af91387eb1c7310f843950d
z0e45aff9b3c1d61f2d34521f9ea7f300d69f0bb84c576e28ec5dbc7a88ac0e1921471dc4a5b38f
za01c69b4e2c5ed8603cd61f44f566deb305afd715b8fdab03b622232a358fac7656f9492d1930b
z44169722b5cf31e18b435262516f5751f16364ab6eb10fe1b80aa28b8e7f56355e7a8ef11abde2
z53c35764209cc69e0a2ff6ee913f3d74b7bece0df06c373911972b6d270ea51786541d3331c938
ze6e0d8725f85a3e4ca93a01fdf0fb97d568cb16ed6ea0892f9e4e134d7b692bd784a2b5723baf4
zb0f2b0e21f6b5524ef8d177201398f28a6919ce79bd799a07e527b5dea81d9f168f5d5bc23298e
z55c6a6aed36094a2583869e1eb0d4498cf6a9ddfacc5a43aeec78fa88a78a953f84868691d0835
z07ed2679903528595948f151f480c5e1b58cd8dcbbd9a0f1e0e6365eec2ad0bdbf6f91a678e148
z7e0e57603e8a1a39081b86807719374ad5c57d713d237b35844c1417ce98d50a5b2c3a4df0cc09
z07c9ded2d5775638a417bbe065397332f363d02842e6c13616166e113a46fce044348134330555
zabacfe344e89b50f0176c566ebe0ade99ad9977c38e016cb6871b609a55915708d299bfeeed91f
z8843df40508dbbce20e1f80b91b48fbf01eb7cdde82632cff3b1795518155d887ec48885feee48
z04542ef379303bfc74b3048e8870c94ed984e3002378a4ba29e3d72418bae62989cfb7a3fa05ae
za5e862f7098b9b512d0cc9b52e89c0cb979a941335d29567afbb5e96bd132993b8154fb273ccb9
z07392065cc3e1838ea68f96fa015c783424dce7b7c37b783bf71ffccd9d95e9a9e15ff14e36a9a
z7954ebb591825f329706665b7a63ad776458d26dbc10bad4467180b14d99d3a980ab8a6b9ebe37
z5939ca5c67ae41b802051228cb20c35ff71150f34d6e5299504ef8f41cfcf508376a689658b3dd
zf88bf8833c888e0df791b7d225a6c67bc563d51ecc991e02a48ca7ba7173b578712c92e1c6bf80
z3462322fa18c682ed24a4be1a201b86e03d0e639699bfc9f35060abc4ba9b0eb16607f3f5fbae4
z88eeca7d5fa76f9f1bb3e8dd355c78505e552645203f5fddf925ccc9b9a44cd87969697c1c1726
zf1bd8aa6ebbb608ce5a2ab8b20db34a1f3b364882abbe72c16f6aa404e4864b4965762725b9dd7
z8745d32f0548b01d5371b061cba9e706fd50089106df172d65f2cf4363c727afb981afe1f8964f
z230e55b1c3d740d29f44288ba61e5c0c02f0fb78ef7b36de321fe8b51f6305493ae140d16e921f
z6a9791cace56f37de9c48c00dc44ad0cdd29b0eb2d1f2a005b6c58d6f06a56969c85e846ec920d
z5b6bda3ee5dfe9e09fc4426923a3c58247370e709e9f7989823fe496b1cc4e6d03b59077aa0a33
z050b8cc18083c531fd0c9174bdb2f819d712381e1bfeb74251f5ad072c6b51a7b3c9796bdc3fff
z20bbcb82a086b1e99c8c945c147caff010970e98f54157a4c727f527bce17b06b23a6b8ad8d3b4
z34ea3f2d4f72576d50ed77fc00bcf62568d81ebbbca23c3d2429958e3953a3cc0196e16db3b6af
z0aad5603fa8dac5e7998bc3c6d04fe08a3410ff7907c2ff0f7ff205c219ff59363e70574668a90
z06345e640ca3e0db0b7c921087699b1fd0af1bbfb781126fa00689e0bcbe1c4518aafd0ecd9df3
zf9b00534a4a667a80fd1fe4264848acb604a1f474b4d7d55109f80a4ff9d39d49d8d0856c6dc09
z76e2fe572c97da259dcba18ae036efaaf54c17b4fc4e990e3df28c0abb05245e3a10f5f67fce55
zdbc879697eae98c52b036cd2b4bb1f6135ede9dcc18ec6929f9c9d539796baa8f3b6784ab16df0
za309f3f3b354f7eb309a21204773144affd2750deec5c011dc8d02e21b12c14c3378c0ccb6344a
zf85c753a1519e6347bcd2d9c8aa2aa6a7b9bd51ba81b01ff8eb81cb0eb4dde3b19e5bc58c68723
z211c5fc32386af83f92729d6397f5e02507fef8d84cd962c53e1492b85bcf4eb3527ebffcec962
z3c66c792c60b76714effebc8fbd65ecd033d52e006a201fb11acadb6fdd9b3b182ffccd66bbba9
ze55786f64a2fb7b7fd012e8fb08a39fb155c85c61898bdbf7689c3459aa130c437f239121c68bb
z779cf75a266159f3010259f4669d1cc008624448a8779473091e0c35d846c3c3acde8d89ebdff3
zbd7590b4b7f7589276971e590668c66d93d69dd0d71faaa7cf61ccd7d3cbb3b7919b0c6d0c9062
z74a2d687a144a3d69be7bdc1643b4a47fd2479c97eab93a2290afaed0e31b7b87a5fa396c7dd5b
zc737dfc05b32a1ffc65ceb2b7087da3b53c472ca5b495ecb9d3506dc80ff18f6b65574f0073462
z2e13e183f8043c2d6a35a2b098ea5c3dbcc02ce396f3f13cbb96b82b6ae5eae670692e6c56535a
z373688188de3a8de714eb0b0ca0de2b0c03081eda2945918b33b580afdd4a1a537314e9c658b89
zffcdc8a55f71c8a3ca2c5a82461e3e4224218e08f86abc01d9d175381c1dcec61116d4eaa9d53b
zea82dd3c1764220990e65f6b3f380c177ef83e042a1eb13ddb4568ae35f9f2ad516c5b43401d2f
z0ee6fbf5b9233c3a09d1bcbd3a700a8fb35e6067d3bf3184c915ac5e70ed7241b60fdde577e5c7
z970295ec0d357405f6bef19861c273f720b265ae755dfc237ce7fa6f2ff458b8442dc8d40768c2
z49120fc8abc455c8f62a50958cfd95383134e715cebed5d28126946e4f1c2e4045503f00814dbc
zee11bf3173e276016d565534adfca2fa7d516c9e5f116616deae6c36f2545e78f65342fd295dba
zf7fbff587fd36f88ef72f149b660e9c42d48b015163e5998ecb49439268c9accd78298881eee0c
z4fc6a15c69d5c535212940e979746ae353e2f830eb9cd639fafd2651bf8012819909de9c5ff8a6
z11d64e4afb1be9c8476c657138b3bd3a91b44aa29bed6d6465e056a206707523adfaa864d6c224
z2ccbe1842b01124160d8e2ec1af43eaec0dd93aefb1cdfb91c82d1dd99520f4584d74e5332329c
z6c7a546b308a1b55189d7d63ad7b8e6adeed18c5f18b0750ba829f1f45e71754d0c7765592c94c
z45b7681802c4c131675427c6acb55ebf7f80f8cc49e0f305ee281a2d2cb188993af7a036576de6
z515599bb1c6d9f44a1d31469a60632decbd5d2be05c4a8a2e174e03e5ebfb574c58d0a92646a37
z98e9325d27a05ffeaa775114bfbfba9352539f0340f033c4fb2227b591b54034f033d831428bfd
z4706c88b0d437a3a84cbb85333ac3d862c97ac110c18dd714130996c6b6fb00a39863079f4eea1
z8fcce2b9aef163da47a03785a18a3b7d961a67430bd753d4ed208855a75d6726ade8c4337d8a38
z6085ae3fcff71a4b7dfad17254cee7c77629d9b6680090066b4ed1dd9079ad1bee745307c9a432
zb3511d41fd78b780dc533ec8fa743bbec022ad2af69eed3a203224f0667cf5040bb169f4c61057
zd74ef9d94984a46d617db57d3caa2d1ec730110b32ca8082e5fd548167c5980337f224927790bb
z78ef5e51a1ef095b5aa90283ff018ee0cfa72e0e8a3d1fb47af5f19f8e9a68bcd71dc2f90ee3aa
ze83285e77a61da2882632cec5c0cf058c9473938a32dd4a0dfa564ecc20928c447428eff71afb0
z0ea1814db3c9566762d7c8f7e27a2e1d357c70ccdb8a6a4c2b4b135e47dcca03d3cc042f55a8f6
z159b6dcdc3f623f08c72d92319d9d34f200498dbd62c340f94d3ffc017073d79bcd257e8b3592a
z9c56f71f61479ed33f64b7afd068dea10a4531b77b7ac25adc1c7458cb19db1e05e01d85ffa845
zf339f6f24811fc918a58bb1bee5c8eda6717e9edcdd44100a55be5412dbc39b8b287211f0e219e
z9191e77c351945af59caeb3ead0b65babd99ea8a1a9fced2ebd79578f065cec0b8e95bd1e2ccc6
z9e9632c0963573e84a8b34cf967ce8d68f1bb31beedb33c3d31bc2c561e81b46da3502568fe131
z861dee04043040afcd81f413440542de25a41e5ab5b54a44cbc369e982743f5820a8c0534a2a16
z81fdb724d3e68129c239f26f80552a7992028dc719242f7fa89e3aa8d4f9f9324276621aec3ed2
zfd629b955377204d4759bf9a65f3d9beedfdbb453c8b9eb5356216d7adc35373889ad2a0b123f4
zc296ee2bda79de67185ecda583c6cd28dba3521f84e4e8f8a4cef97712175994c38b1af5395f89
z4a07697204e7934677ee20ad7b633506d75e9c27110164a22a93782e5133e54d7b51334bfd1a81
zd3a8c2120516a105b38c2e833ffec396238806a5334a70a6d7955f8ac56c48ecd3d2cc8a587958
z52d4e36eda71718bf2689e27e35caa700e5ade3ae9db4d6110170f232856e9f05c386501a7653f
zafa5280535e64a0c5a9361d8e63741a491960b5187f247c4cf4d5f2893d87161de7ac2c4f59c2d
z8f218375bbc513d03cd90020d355e055e167eec3de5a13ba7ff0545cda41bb422ea736d800e591
z9854ce70feb3e77c8ca226d10c209e17a146e3b7980ccc54f6aa58271eaefcdd4e5f7692337698
z31f7a188a8b60e21d90f7fc58d25dfbce83496ba0ef07b0f6f59c0a9ab2e6cbde5d7a2091cd27d
zb223a1128bbf454d1b5771f42a0ecba97f790f3423fa8dc56eeb52a541295e35625cbb59db09dc
zd21985fffe8c523cc068c702b4a374ffc8a999edf31edcba5525d4f6e6f89f6cf9fead65301367
z68f053535f31352bbf7759b7cbfd86919d18c53080231d236b3f59305bd7db8127821dced5f32e
zf80c75222880caae42b6f18c48ee9fd8821798ec5546a4e80cc5dd24af1da0cdcddb343c47a1fc
z543f873cef37ab38ab894874ca3ed0e102471329d2928f1c4f03f032210eb733d711542f228852
z3a6aa53c261115997485013059ce555f386a3e13254970e9901d30e3e5a8644a6a5ca75db0515d
z29fbf6d7ec7ab183fcb74cac4d827165908c3cbefd604757cbf50949390087c181fe7b97ce10d5
z673a57670f83f97cf0b09e355d98362d1c019af5ed549d1917b6b5ba2d3bdb3d8eebc031557955
z5b12044a3ea7dc465eab73661c22d38d337e6db2c8512c1b3d6361101cd33c4426e797de418327
z1119c5742bcb554e660c3bb137358bf5730de616338acdcee705757801a06696d9240633d76322
z46a4c6df4f47251b714f58b80b3f2b2b3f0593a01f1451befff6592ad053e338b78b581cb6428d
z94ffd1ea1e5957f7dad16238807945e8c4b90f187dd0659679711a292f63ddc227fae56a349b36
z639ddc27769424c18ed1c58d293de082094048103163a25a70d85292f69f45229fffe88a7e93a2
z63cd2791c8d4ed52442f3968b6c411a0dde46beb8431115e45a751dcef41b153ae5c0716dcb454
z375d283c49e5589de477438e54ee3865bd855e7bedc6b5ff421fd14c285ad8b28b5e265c601b90
z9a71b8b2e17c803ba5ce846a09bc1c8a9c10424f8310632b695c09d3ff23b0b96edb3e61bb2e41
z8bf755aba844db486c92f99ac8e9bf5ae6ec8931352822b1cb52a17b7b662c8e5ede0a8d501922
z4e71ee847100057986a50799fa82665daf3b2fa5b8c29b51f4b11dfbeb70f50e0f32b9f86439a2
z744c054acbb1e9a327211833c74d6286f76085ddb96ddbf2b595bfbdaf510b4920a846361b4a7f
z170dc1f538ff698ae582c5c699cbb3a204f96d103138a0b6e59427d1485f33d0a278436d024897
z61c13e5f30d59db80d6e796689a7247585b68ff3ef99b8f68fbdcba8c6268bb82c15e9be462806
z54ad2ed0198e0c0f1d0df1fffd420d0295b952be4795a51fe5606c56618d63faee5c4795ec89e7
z669aab31f903e9583b3a482111afecbbf3f8802fd344931f299a0cf1a2dc87470e074c8b411de2
z5f97b51c6099b314b2a3d3d006a597980fe105e2a16e2cc9bce05bc534d8e57d4f4e0f7702f1df
zda94753e968e94e2e16e82d02e2e4e0f1e5dab9c83009a0c098cc2146d0145352487095860d911
z18c220831d6ba0759edfaf8428a95a1eca6ff5193232b193874047d5f2d37e9679c8200e27ef7f
z6c30a9163bc93ffc1d0691898643a0deaf89f07c297a7d3922e394069881a3f5a715ccbbde8030
zc84a70fc7fe5ae4b508e061916cd0f7c2a8757cf9158fb641622a2c1dfc4cf2cba1019df81729f
zf15a52dfa524cc4ec78c61bf95a8cdf80fbb4b11bcb504fe46a69340afdd456424a5778fdbbe3a
z46002e325ebb879f27424c3ad95c599b31b491787f66e8c4894ea37365285ff50e037535d67436
z8189aa6a5972cd82a898646396817a4f97f5596803ee05997c62012c603b4ecbfba91605e2fe6f
z9e5f022159a6fc8bbb15a141c02ecc5d5136f50afed8c86207d1e6a9666ceb9d819ad9e876ca45
zcd3dcaa4cfc7909e9e24857817ce8ee8782731211d23c4ca60a8f7b6880a7c570f4775aece1d07
z2fcdfd75caa7011eaeed6316b421b6690278e3fe883a35208dd04c1f89349a05f043ed4c01fdb8
zc009bb001e516b20f06e501a4dd960b2440a826caa1224d393fe98a5cd00398b4ca6cac613d405
z1ef63420beed00de7fe6bb7c4a5b0ecde0e223f509a3a69f1a120e08fa101ab6f6c88c9322c91b
z957514572163b68edb164eac80dc385fb7fecc0cf2fafac5dd25a3bb9e0bf6b7f0991b4c762112
z07719044110a5e095a5a1096963c3397862b06bc97ef09ffe0b1b44f7a91cdd84aca8fff57f6d8
z26a8f252da04fc08beee3219f5151159e741baec72a8e2f4d64a6a89ccf34d2563e46342a39f14
z680e2e95fcdb0f960f56c438002cef6e8bf6a4bcba64c7462ca7b5d183adfc48c8433f5c373f90
z4383102d346b2c97fa7909dae2d6e1a005c8d7f6307b0d3db9d91905ecead85c5ede4ff2ed37b0
zbc21d1d5b2151711789f4d984551f4126bd857a25b390b186d241a2f5ca8fedcc4462da6eda7ba
z0c8264ba7f64f3c94867add1637d62c2a0e143ba1ca94dfc01122cc19c98636db53d956baf0e60
z64d54c7c9bf641a02582d9bc2d67ffe26b3d0ddd0aacf19049b65376d623361b9142a94a2ab159
z0932930db7faedab0cdd0cbdf30b920fa2d5ab52a79fbf18332f29b047a9b9a923d553f30185ad
z4723894a3b1fd966da440c413efb149e4481d92287cd4aa6e711e213a0aa1e3ed2f1f06330919f
zb5c7684f72382d4b0787b60e9190d76cebeadea4d269c52d46885feb2e84f69de4ba978b31d2dd
z13d2adeca4dbdd849d8ffb450934a922ea489939e0c6b33c7ffddf24b8f1aa131d5382de4bf1a5
zcec1397fa348630d51ba2e5874b1b1fc466f13be7ff9b7d808c03e52fdfe401b394ee7e798a061
z9175a521c0b58bbe6f893f071b81a26703651ce16608f8505a62bf73422f58709a035a11e4a83c
z6e288773599bb1289d6c7e10e4299e33c4e15dc725408269cdb2dee31147ab45b81f4b71de7f9d
z8ced347041c0d97275e1461d83c9b893aca7994207a3d25dd9fd162557b4ae051ad5252a8f2c4c
z8feef1feeda54d0bd52d2a36018ddb7c1e970adcd14a8165014fb966fed3b1f37d2a979f49e9cd
ze5ada76b36958bbbdfe7c950ffbcc4ea32234ff8e619e2029b1b5c942045e3272b934a127b0772
ze58ab14b1e3f618b1e97963bc3401723c87172819b81a2b247f88597ec04dac3c796d7eee41e7b
zcf49fa257e5de94ed06fb229efaf1708b10a633ea340ddd775fa4838ee97d7b452a0c9405e6b95
z9b46a60d652845cbd2ca28456e8beac9f94dc45129ea8e869b7152d4d2864ce805a0b530252901
z2642aeb42bccb0a93d610cbb47366f66b0d5e5c0c1fdc22be2cb375b112f6a8327504d8b0d1c15
zcdd356b52f6df0cef2bbdd0dadec5d42f8c87ad58485a8bb7d9e31388101c51581559087c5b406
z7532e9869c588e899cf1279bf6fa89857660be166f337726c9cd6dc6e9ba511bbf16056e0cdb62
z432251da40d3973488a143ea9564bfcb327adf44812b346a1ba2b73a8fb0158af6399add177604
ze25e202eed040c69b9de1f71f2a3f7a0ed3ed1e565dcee07455f09a9a52a9650e800e6bcc79c4d
zc16c9fe0e3a0215ea220199b34e4c650d0a1466ef9a3edecc0ebd008f5e8dfd08cb549c6827c8a
z0e212c51a88534ae3a35ce94a33a8ef7b67643eb103acd4c37099551b028443c56d144834379e8
z125036622eaf39046c60c76110f44b39de9413449a1ccf74b64c2b3a4ab375e4bea064005d7e48
z684ebb56d9c7a54373e3c27871ad5d8df99f8642985cba985d951d225cceac4c8ebda834388e3d
zb545d5eb7a7a023799018aaa6f4b867f85b6b9ec698fdd1ec76291c75c260c94a5727fc7d44610
zd2504a8db3273150316bd00c12ae3425f158b278ae954f697e5ae829228fd8056c2b1110874bf0
z3646f320d13cf7bc67407bca186247fedda58b53ce2d81dfba13f1c2df0da75ca7db1dae5a25cc
z16b0a753a25eb6e95ea87830a8384f8e057178bfd3b24b17a4862fb571624bfae228383adddb45
z7711902855388a432818f2844275671c4916884e403983d056a42ca49a7c1e85ab50f9f02deaeb
z8e6729bca2b6b0c98e241f73c82c5adb540a458fbdc674d81a6aca3011776ebd4c02eecd5e5c3a
z2f077966b6a70ab995b53bfcc0371c6ac32b04fbfc3702a710bd4255fe123e41347e79ba844072
z65d42560295e41ff6fb35ecb76c4f71bf011568e623ec9236d68702a750852dca7c789cdc6978f
z358f5771068b33693df43faec955e244305ad34abe55793d134bca5d3bc0a430c36d61b95d5f43
z8d1a5f6ebf8491468d9ffe3d864d26256dce63f6ffb4ccd293a784eab4dbed29b906bb78c369a6
z6400dbe347d570e83ec52af1853f4ddf02e6f66915c5cf65380174a3e596a8407dc6c6a733ec7b
z4ff5a824042faf3d93ebd770586b9b5f830ad5778c2ac836177bb6a4cc3c2221594e69239d086d
z6bb63f28c910689f691fdf62be07c0bd18cf7d1877443f0b596aaaa1ea74f182bc5ea596a0e39b
za999a7dc38b744b06a3f29fd8a1b42d13694dc8a1f1d130e3b4a8be0a25e39426f1e288b42ca0c
z8a83c2c64481a06fd5b9a6c4006132786c354446a57d3cd785ca571dd1ffa42b33b1ecfd1b0a19
zdf89ce4bc913f7030fbc032ff614ef4d672b819987111c2a34b492145dd531d775b0f46bec2c3a
zcbaf484628c3c597fb8904d1fa0edd35e5eb635dc756648cc58d9cd870b6b3cef893c28499ff00
z232544f45a05694e5484521c488ac01307f14e7e81daa82bbddbf914d624bf45dac043c84d599e
z7f2fa7afd50cf9a29818b3876649e67a7ea6b3b897602c6add758cbf6f7a4d4324992fac9421ad
ze95d34b6d6c46854684ee4d8d65c86464a7b0993c32ed9a1122af32bf93e73708bd7a35c9a895f
z96fa46d341c836616807dd4c21a63895341f5d055943c3363acc796ba3d2e303cb40eb590c4e2f
z3e70b37e3f0b4209d7657c627a944c8e075fe5b4dd6baed1aa8a9da3c6a19c1110a56d01a61567
z8fab88981c9a7326a9c4483d467d1adbff4932cb08be9eace438f0bbc54f2806db26f578673378
zc046fbe4b38e6db64da2eb7263c709fa5bf7e9be008b78f2b84e4d0950f02ed2e0d02cd9265cdd
z8fc34994a109c985df63d702830f551cf36b6d9c86077b82e972ade45754cc39c88d6bb25aa572
zf7530ba8fc47e863e9e9f7e8621bf38465a06e81163c9d9e074baba58680b0ff16aee4e86509f7
zaab6cc3eae8715221ff76e5704025eec1b092f0054e7599e7435ddf529d229d4dc070035a6154b
za6645da52938de120cfd1f0bbe355fc13e42da8c427eb3d201257f013551e9be0dd016872be466
zd31d5db7ffe084ede443f8ec5ec1a84befe53d870d3799e876a3dc35fb5785a343299f8b88c445
z07a3dd035d909adfabafee264d62cf123cd634f8f8b6371fc106839fbee96d6a0e23b79c6d9a6c
z93e97213a80db02afcdb617444b10eeb887d903f5792aad2afd63d92ff73e03f4e971c2bb7e858
z3636a887a2eedcee05cab2d58f09d87ed5f4ebead857284f37087ebbd82ba29f58d217feb5ac40
z8ac677fee089ce4f00d39d10b94ae13818ac3b4b694ffb0f91aaf5ec7d54fb874dff491378d776
z8037ced261e7b7fc0b66c27d880edb083b154f4624f0e08ed6b5ccbdebdb80c0c0ead71e67df98
zd440e4ff6ba1fa985b6c06fe55e587a0a7c32a65440118a38e8fd7afc4b5f3ca4807a7825b6d63
zb41d180a2c803ce03d2a4fdf0fc809bf9aea14b7cb967a8e09113cc2bb95a55b68dd2767e36ff0
zb958936139fcffd42d5e7b610350a4b618687275bced7416f0033c929ace1b9f7ab1f2ea19291a
z6079e9b23422af628b52686349ad0e6125824d85b507d6b38b3a116cfbfca1880928711e04a6be
za38ae9eaec2849df3e8d97d5d1077eb9d5524c1b04a4ee31c26100361c50cff7626b9c772f9f1d
z8d5ec30d0f11046271d3372c68bc285720867ae259bb81665ef950606df86e5a5ec6c00afa2986
za646cea38774b5187bc5f7870904bdf1ff1fab2e4f47c388cd510954b37735f350cab1d5448775
zc557b94c30061037d6861d80069793d87132f97724ba9df02d09cb9f7c43bac54dca11a4d99bd6
z273ee3464def122902aec991a59907f3dbbe1cdef690a6da76d84c0120e357176342f77345d10b
zf871011d95154098de56c818d6fcd5b81af3ee46316cb48823fd6d240dbcd2e96f3695218a12fa
z937da2a36864852fc1f62db85c9a32b30211311d8774dcd45fcf7530a5a7315aa6f6cc67356946
zbc8dbbc61ab8514540b920ee2d3e86b4c9cfd42f8b75f42cfab065009f7f9c9d43153a1bb7453a
z550c7b5335867e0e03f59c9ece3d5890443ea3eacdc186a8c4a9c4e008d8113084f5e7bb60af24
z0c85d69471c8b10df69dcdc817586f6f1d74099c4b3ae8bec9d1be5bf9fc3c68f6e3fcaad2de56
zb534b51e9bd84b2111bc58c0f9d3ac00148ded76fd525237a01f57bb24ce24736fcbf8e04f82e8
z41d3ab9d99f4080afbdc0f9db4c25f1083dff31c519432fc728ee3f678ba84ad7ac8281e728ea7
z5ced415e753cecf9bbf1d0f0f0d2140cfb6dedd5d29fff0d442305a865951c479039f7564a53ee
z68d960aa76baca151bc40cbceb6f1f0bcc50a8e579c147aa9997a280aa7f65662db73ff4aced05
z2896586380939190cbe6a50fa1735cfc15f284689d0316e21f0f8411a8b18c2028c6e1ff439e48
z1a9f7ccd19b242eaa5e60b1d4a920510cb0e28aa0994e64c8af0abe706e610ac43e02ce1dadf99
z1e5f855487b674d51ad8829cfbb3ba99734d56b30b72fc14acb7e16819cc035cad1c825f970d56
z212037576c6a9227c476f94958bf0aaca93ce33656731e4a7e51adb579c464be28ec3387e3c9de
z78bdd63d20b092b736765f91d4021e3e90c1f53c33d08951cc217b2b43ebe14a62cd20076e0727
z2ed3bee06fa6c4510c6a0c8f781e47a285ecca6c294fa8669a7b77d93cf5bb6e401750374bd125
z7324c99f208b3a712d87de2c6a660b5e0f9a4f55eb7b65d5488b2064aa58a5a9981e96769ead2b
zce9b653d62156b3e27ab39cc1b77d8ab21602c836151ab78e21c098688c8b29a1da10ab3fcd140
z0c6288548959762b493e11c4993a72955f86b3f6a6ec3bbc57a2d5e8f16f2ec1af55e63409aab1
z3c6ec8aab110fec7d72482e77c9a6529cbba29f661ab4012a72c98bf0a6a1871f425dcef4f4342
z3e5d71ad20150668e32e05ea7d02cb61b5be3551935a13c5bf658105084c9d143eaef43ce08804
z224c58dd68be691655b94320f7cd52921a734694eefb693d848db34983c641a8ad1a041d4380e4
z318031db02f1deb4c219da2c87bbe15b5e68e9f4da2d9e8bdbcefc9c1037a99b5b52eaeefd5f35
z5e52f96d78e97990ba627666b85c1f76253110bcff1663738e5eeff5e136b4d4e9dba38aff7df8
z06c83303943f1a86f10a2e0ebd2ea3cb83bb5d1bc18708f6acb6901cc91765197186b84d968c89
zdf4532288318915790ae4d75a39cb402b5705eb55f0905c3444e471b3c7c22fb73e72b00acc1ed
z0a89c48bdd6e1d9614b016b2943732180114596918a5322ee2cf65c7dab3a5a540ee59a16003dd
z6104dfd5e960006833b5f154b727ca85a481540c58c8396d5d7cc3e11f0684cc46e6fce6b0c5be
z6ef68b4585cb8b923cbdeb3b62fe60c09cef1bc6d23bc2bb181e497c2b060575732e1306c140e1
z596451fa6dd3ce7fbcc21992f8a7f578c289524f296c40b8d26972b1e5490cebc10173b8dbf314
zc7c630a9a0885850b4509cd443f40ea3f66910f17affe7c8680df12f18bd2fedf1c7a1ad20d02b
z0db721550db6882e59af66e5eea47ce8f1d86c652307bf2dab676c44f97f2baab519a5c71afc88
z67686d6caa0ad6387375addb5f17a5af051aef2420287c90fbdf72f6b082f4c274301c43b6f799
ze60ec122a0b28cf9c52daf515d3bb223420389457449017c863b4d9a6ac6e9828eeb78714c2560
z277442f488c5288e956c2ec1959eb5142225d926281650ad35870b9395d6c0959ef67b1c68eb87
z16f0499b068bcd2a190d28ed1f7bfc9ad246dba431a0b45323f722f07afab8566b69201444b55b
zed8cf47fb502c4404a62709353f5bdc82fbef7e5b8f1c2ed4cb391b764c2f9e712ce0ad9179c3d
zbb62581019588029bc9aee8c1be1d6cfe9d6364f0da847378524df808b2b144ae2d22982335590
zbd8af66d5b65ad37ffe2231bac3ca2a6d4cb05de66af17586f43f3673f663df3794c3bc77ee5a1
zb97faa83f6e057f9ab33822e5e1be03fcc2e0aa7ecf1181d5b7b0a8a1281886ce9384dc759fd8f
zb98266b1f0825be0ec7c500ca2818ab0337c3a4ea434d839f4dabda50ba2f426a96e4ad01b8ae4
z25e5f68951e6249b0c19ce5ed2e768290841a451d2d0b77ef857023ef5d1add7e3d8671d216667
za3dc525f2059a25cecd5bf3a2541ff383c217b25b03a3f48cd32a5f146a9e8d652ba15b7f76729
z5752c9ee478c74078ffda741c8f7cf25fb820db8b423f07c2fca9af22ac36793c4507fe29cf611
zca98d93dd66ba75a771d4cf7ea5939c86d8ba392ab90b1226704faecde50f7f0187c8cd276afa7
zcdd697254d4d95b2a67e94e4c342c727673f2062286470d39b69f1123956e67e5e2230546af445
z54ce27b6ce0bc1c3df2b477e88a23d21bb57fee79e4145aff34009fe9ca4751addc8f8f40769f7
z9a3d1215f0e9245b249e6f0ca1b5d98441288b7f6a2f15209e3ca404200f5f1199ecfd1732e4ca
z9203d21e410a7a23dd0f4f0c55dbe13e782dc97c447d0cb5243d8a4249fadf32e6d4d9253b68a1
z085f0c10c0708a7a0b3a33117e0ff251feecfe16faf42d0d69e39c96ad891ccab34e48265c11fa
ze155f692f866890345b5ad74a45b02597eacd00faffd7c7e1d35e70f5d62fcc61ad7ecfa06798e
z7fa926f2e09b08585ac494973381adb59819006bc9091a6a063c4f8d7d4915b177ceb28f2656cc
z4e625946c8a3689a96400c65742d5540e4d171815b936f76faa65309fdd6d3e1a7ce5e0ad8b3de
zc17815af64193bc898f0818aa8706bdb2e7017b8801cda37ba638fac625a1301c2fdc878a475b4
z6ccc07b4e77c99dc992b1bc41b74c73eef811171a5ac6ff3ea1c47ff828e70d411f9b6d13b7bb5
z52fd7db02cf8145dbefd3d36ad761169f9b19ed1578a2d6d7dca33b888608afdce11a89f82fcaa
zf03b73696d2a9b60d26752cf5fbc24cc3415061b1c63a66856d096aa3356a5b33e46ab48f0dc40
zc7335cd772a470a3da2ca3356eefbebf8b1da0e184be8cd710db4a4a748346edca69a2d6f8d850
zab0d5dbc173b66140c2a5c9884438f3fd7047b3b622a105eb817f97566e50f4c7d6f4c7c9332f4
z2414a5f83c581f552b7f048d1df1febfb26729c8d9e3a3fd1cc169ff550c53d9fa3e5a8159fb9d
z8e646cd8b92006c3051ac29771d01092264880940add67356a05437e1406915b95eb5150f9c192
z2ed923de45f578e276fcdb7e1b668c6de089066cf8a23c0443e18a14086819b50c7b736d023eb2
zd6d2e63ac5403d135a5c986ae81bc8603088a003cb7ad83d1ef519a43cd45123dce9c5eb0c05a4
zf8b7e8286d2e856d14a38b8fa4ae00dcecb5c2a1760a282d39c0b774854a83bff4c8b5ebc80a00
zfad2bd30d21c61996ab0ae8c26f7ada64f87fa9b579974133dc8ce844c3219a780366808b5ec77
z9dd35c5cd7cbba3e9989c2a185e269d743e08220e2d95d504f85228ea111a50b801352e595f9e9
z9dfb115bb096c569b8c76aca335c05ce7d1ec135da80f88c91141c4050ed22a77184f55946a73e
zbbbae55910b04e1cb601563d9e3ce80cd30090165b937478531500ed1c32f994b95da6b0643862
zda87e9d80951585f534e2058b75ecd05de2f91134dac3b7d5a162fc9f95311453d0578e7741522
z7c3a05286080adc6bda4ec23aa1f48b6860546929c0d607bdfa28af98af4e0cd88f834fd93a38a
z5a68b9060e0b1f4c678b239703c83eff1306cd0d7c9f1d9d3927a4a3b0ab42f7223927c7c96166
z6f4baf92bf1bb6ef9975584ee91fce438ba1399b53c2c733e4ff53ddfc289842829529288834da
z6fb98d62b18ede44a12c5cb27f18a6d9f25578dc34a5a635a340abfd7ac1b024dc7fd7f6cba143
z50c121ad7c0beefab50da0aa879b983fee9afd619447110c7c37b99896395e3c87c1e8e04a922e
z2a1e10e9e3f87de9d02484fa5c5e3b29bd0572f790afd8be94d0680765dc06d1f8a895f707d044
z361489285f9d3dc5a4372ce9a0e627444c04c1dabd80024e536c15614657c045abfb6c1b160e1e
z5bd180c9e3f2155d1433489e8a9723bf0a6db104605082ea7863a055efe93edfdf637cf7f9bcba
zf4d4e27151975477bb98ef70986b4c874494dda2be79a79d92337d46bd0de50b6843669662b4ca
zf89f3265f8ab330fc8061cbe7b19a55c05de979eb3014f9ad138859c6f83d0a7ea5db454520c5b
ze7011d2b5b85d3e29ef8910dac23a49e420a78f8e2e24a96c16fd39fd1ce1fdf8f605487697cc1
z6130a2d2d0b4afc12d2f346e46c47a7bf67d91575e267b44d25301675b731101ec8bd086afdbd3
z6efdcfc4ccddf8e8e706acf8adbe5153b4bba042077d439123390aee18f24e0097fc5ef87b2462
z86eeeadb2d02acf55b4150a652e7b5964ff1a919c382e5148b3b8f47e750b7f444700ebac5eee3
z40621e654db018b644062a55fe53b8c179515d81e0a436dfa38a90a156a83ad7ac1f8cc8348548
zf638ab522cd42d0c8f7c509eeef01400c7783c375dc98a1eabe0cd033262b0290143b9c2bb892d
z9809c878729e7336c3c1acfb63482a7b6de707d3b1bb75fc80bcff54f146267e8480e53850c3fd
z239ac89dff303a3f3302b38d6fdbe6422fa2c7c1fcb2be8376c8854e5b5b3b5b65047d3a8e06a8
z7cb0da0067ec93331f33814f0e6ee3abb84af1c3df97551ef1dc22e2af5806c3dd059dc7beb501
z8c220d8e447bba7ac46e757f82c541026c4acee8f5017ce647bcdb2fd61f2870900eed9844170a
z2db956b1bfe10f4c4b78bb0092261f2349fa52559050d1ffead150cb67d9ad6d523ad725c24f29
z8586d9f93c6dace8f315a064df66a807e752dc454e41f645684ed9aff7606d58b50de5365ce485
zded135e9783d5bc9e2c17f501ce0d7225682c54200ec6049799d7d7727d09e5f6acc55e7bdccdb
zd88dff1d045674299c7b603d94e3f07049c81fb5ed533535e5e20be528bccda0f114bef2c72cd6
z126eb521479af23969ab77bc71c5968121c4c516b0397519830b517fc487d75d36c289cda5a98c
zf6f127828c8412c0ed97427421e6e849b3ac596a4f0d2fa933413a3ab87aa48043bde9dc2c1955
z555ed060dedf0ac2a862adc05eb60b0a23507b48617bf471f45c9d2d4ea5504884630cfb4898d2
z896936b5b222395fe4ed4ed1c3cfd6b8e66f07f8d9b7fba76a86a8066c23df02dc21e2e888c577
zdf3535a420d5c4c39a558c651b494590acf0a2c995f8dee52fd34e1fb7299bfa870e802a5da587
ze01c079c82bc21b60b0eb12a5c86c923d7af3d54c64829605a096ea58fd50eed4db7509bb47aab
z70323bc1626289778843120f5ccad940e02525eb5a787665a8e9f014a489fa140004087e58d3b8
ze6adb9ebcc2d7ebb1608ff67b4ea99c632232e2453df31ff47812a02c392836e560b1a062f0419
z6fa8bd21fe10cbdf7d8d81afc10b0af919bd86cee64ccd2c71e8b03f1115601eae625b725473dc
zac3467445dde840b8f70a270f3af9646d1f80b92782210a79f24b4d97fdc342002ecab83baafa8
z0c958c9b204cdfd1abd3bae0c1a9db9da8f5e843a8d8330e5d576e39ef86d4d7f12a19daf9fbff
z4d2afeb9040ada13b11cdf94cfff3ff4875341e3ee0483e3b1109f139af34e755bed9b6432b526
zfbd12b2410855faf77304d82963cef029f8da08d1e9cef08866df0af7e921a43a4bacf77964788
z89b9f5b8a408d9b3a04040ba8bd0c7f04fb3a29dc3d2a203a91a2486caec001809aeb394aa7fdf
zf09e1d1270537b84df266e6b862a6c1f875746eca38b7a30925eccb8f862d9f3bf05e1eee3743b
zbf073a2d80c47de75fe2e2308bf48f4e1efc399af6864641038e863e2a805891e7be8f075019ee
zc4cc52f9ea700f21f213fc3ee90c15cdd559201e34cc5e572c845f29659e65cab877e07fced702
z2161e528cbe0cc21673ce1b4afdeea45a1221da5fad6017153455d6e0986d58f5c5e9f14b3f9b2
z333aa05d46a39a0368d5383d54db493106f50c04405244f4ea181f29a99a26aebf488759aaa9a1
z62ed74a7dde3e94a7965ae78df27c089d63bf6b1074da16aed46a25e12128bf2ae056fb71dfcbc
z597d2fa34a2b13d9e9cde8f7cfedcfeac17f73b18afe601e4daf5903514e30a090483d620790d3
z20af12555e6410d531f7af61f70b8f8a1be117cce2cd0e8bc9580c91d184897f6d9e4429d876be
zc754756dac5bb65cd33fcd40192341864209d7664ec40b9c327486105cf6416d535df1d82c14b1
zbc1d4abb445cf1afcdb0170e4937a8a8e401b9e06010eedd3ac923db1b19480d7b441d9e1367fb
zf5198f14f73b620d705dc83f64d4d90107172a09a039b400c55cf8be6181952f1a9cc2cc5c4214
z84a2f870231a2afcabc4550b18a9d6a52de8d4f446c1595c595625c48ba5c401abacaf95228744
z1bb02f200d20059f2d0bbd97f1a39109b8ee54f165a2117494268e15a4ee6c57c360f100469a0e
z1be271bfee1f0b89c9c0a4f5df7d87b6bb10a75b35fec45c4f65fa9277d72803c73ba5fca59126
z7f331209e494790b87d1ca13ee327604472c43fe02f60fa39723433699656573bf53d91eb07153
z7d7140537a71bbfd344cb7f3769d829935951a896e425b3f869e1918d05b339bdfe78345a27bf8
ze81b992bca4df889b5211faffaf5ad9eb1e4ea60d512d91dde40f21ab6764d2e2830f14451f78a
zcf802335993ab8532805e9856f2f3f42a32eb581e772fd423d74a88de10be47070ff2d5dabda23
zf7162bfcf8f544f8933411679769028e8d8df6483f65aabfe8feb66f466366e650cca16ba556a1
zdbe09a01798487d3a2c2966f7a139a9bf0ba31f00869a32ba7945f52b03f7733b886b2c7da87f1
z8543d318c71ead3dfabf7298f253e44d3d9cd091022e6e51ba86d114895961bbfb98f528efa804
zb1e70c4bbdf261627a2971f393bfa610a1f0280717f1744997bf76ac643f7291aa5d7b07c66075
zaec2899c9863ed6ac59bed6c96552b9583b82234d609b015932031b332571a137ba74c2c30342b
zf416c388da55cf9234625cbed8ed8c4f22b45636aee42c762139cf5e2c4f5ab4cc0964e373ac71
z5af2c78a6967e83b15c968d7d9c64fa98d4ce75d9577a21ab7040564d324a3ceaba8af77d44fde
z1cdb38259661a6350322773de6c58df89945a2a9c63bb9c09279ab8d544dd37087878789633f57
zbbf4b2f868de6836b3a40f4cf4ba4c856f5ed16fa8ad80bd27fdc5c11402902847f2ab5cd0527a
z7744383e9e12ddbef0d7cb57bc4efd44da8810d8df71614534b2899f4f199248ed07b04b54ae53
zed077e46a2503fe804521c2be31431c951713af325fe11519608377c0ff6e482e2a69be4d60c20
z91d529c9742b78f1a46889aeedcc0e34ed2b728ce1f90668382c5c50222809c405af66cc03ab6e
z81bacddd51a865d3eb2881f65f013aabb7a11c94013a7adf837ace43599f20928bbb53eda5e96f
z4e41d2272703d78f4821387b54b96add083c4e2860a5faa0d46442a586556856a8e4e10d65594b
zb48f87fe9440ed24d641c8f3f69c6ac01c083860f01811419dc99ffa6544e60400d7604cf43b83
zff23bb159bb4955183d0b5537a8e2d4323bd2d7d03fe37dbe1432edeb56d665e43d090d4ddcba5
z1d2f78f97a56de20c77a35230c3687371490f4f746f8cce36ad2297c9746667030568deeb4e620
z4729f730c427a8c94f60635d22c05d9ed040533847ee0e18cd27079ba88fc15090d7dd628e1363
z689996529e27f8835707fedc09e367b1deaad6cf4c48447f5c123cc41be13bf894edd6e5266caf
z62e3a9e6b2c64ae1cd1650ae190b3cc561500bb86e39ef662a7b726c99b0e989b24f822a0126d0
z306ad28472c809bc43321a1e32f497d465a1e86f58eaf081b49b2e8d3e65ce75ba41e23dda16ea
z43bdb2d01082d074a9df70199ada3200acc414fd881dc4a9d36e62922a7f9391733ecf5801e57a
za54b70b07cb6370468074d600b5d34f1cc7e44bdb5c15860aa18ba8c145ea2a9dc3cbfcb3e7d7b
z5df9ce269c94abe9618dfc90d225b53b0a3e099126d3ed66135856c750c7675683357a08efd77b
z85fddf168c4f18ea745da860a01e2603109c550959781172811631d3458a161a40542790d9b965
z9ec079f9ee57695d9b41f59b5cbecef47c651d28e2544f3bf66d2975203748638fd1a3a563c668
zc2aa9fc2af0a01bf9704b87307dacf0615185d0546542530630c94513800b20f498c2969cb7599
z8d561f079e5ae1f228883a5939d32615e750198fecd60ae4ad195b5efe9a4c49444bde41ba4432
z5047ad984d0262ae5a5d7ed8eb4acca59a848170f79c254cced419f173dee772153c720e36e7f7
zca1e8f42d6725d001685b265287e7fc56ecf8010956df5457a5faa2d6d26faf6cb5ddbac209cae
zb29f961409c6fddebc64b9cfbdaf0e3619952e6ff5760ec8ca2a435a109bb8feb2a32f009ae156
ze071650f393b84d6cc13cf945a7599f973d6393404180e1e9677017fb02307135f76cdd68ebe81
z28cca3d0e2366c4af2a675cfff419358ebed28038dd8f83dec88852ba7601d0a7af4ba735d37de
z8e4183c3090d384f203fbf9900eef75fd73bfaca5de3c10169d9f2971faa832206c5bd412be813
z4b9929be0c6466cd7841077bfb2da6e969d75e77f7928efe9e546bb173f2752a6004bde18fed1b
z0c03bf1ae90f09432f9b90849e9e05e9897227cf4562fbad551817263038423b976fa483260d1b
z87f47350e522343d757eccd1658571113eb2c4f56256d9974fc88c5687be4c805a928c4b7e92fe
zf6ad31deb2872c253503ad8d8a445c1b037a0f0a9e8c378beb49c5133e2b4c164e9509dd2f2854
z7caea37f68a048001aa4d9aa78dc8117fc8fa44641313669790c378345ca62eafad17b299a585c
zc53d7850fe1911f6b84a24fa55cbe4b7984dbd98a7261ec4e9c91689676682ea4004caeb983450
z8e38c76dd754d24b5a96f8ea0977f5dd9e636e9126ab60f769199986574dd5ca86e39fc88df84d
z5853e4a65e7a0219a12014c98a485dadae5547778c54e0095fc02b61ee2e7a473d764c84b0f197
zd75802d0cf44fc6924482888fff7c5b54bdc3304b90b608aa14fb4aed819b275b15b9a148e1a11
z7b3ba8251c7fa1d66ac92b87413971b407dfb59dab8ff6044e51d0d054e2540609dbbcc2063fb3
zb0b33ab1b08012c65a56bee63e518469fb991605c45061972a3ab8e43cb4180dc28d45a8e63cbe
z1612740bc92e91325055df10eb548b0693fa6d1b1f30098c40662bd938e4e3546fc6a4942a7227
z8a18301006c8f65c9a9b0a17bc8ab686174d1cc9e6f5d9e4caab15c5b21eeb1be31a2d2c996af2
za9fcf42d6e1ffbd6d182c9950ef57da2148b6dd5f5a3137c87d326c6ee09608d2293d2c95528e7
z5ed3d9a46fbd3daa47114ca999e8701f9cbc82968ced1194bb348777542892e008015af3eaa056
z5a4e7e1ab754e874d25cc8551d5d95a8ee99876489831f2c7cf4bfe8da5a2e7e02718bc60024ae
zab2df4c45f25f365863fcbc4aaba1c56e3d2a96f3f5b23025b613ccb7723d4ee34a6faf9a8d0c0
z9f552a1cfca1463f54828af7d809b7ffbd441c91ebe0b64fc7ebdcc8c5b9670288787b4957afe3
z53d00baefd595fd79f3d1b0e68114bfec9fdf905f01cc04501485f1560f06950ef12a0db5b6892
zff0e06d3d01a8d874edee8751028a7c5545a855dc175b55a234069dade4cd314149a4d6fdcfa9b
z30f206f951945d8e67f4efed1956a2caffb459b2fab09e7b601afcf78e2df2f324f336caf42f6a
zf6ca0cf09a49acb29367d6df140d478dd4d177d470cef2da515326ca81f927b69704513ccae96d
zc1286fcd77fdc6d5dab1541a5d89328346725cde6d6113effdc7bb7efa0a61b22158988a1f2e91
za0e98febf44d2100d1c94486d799d466cf4b9037e2bebf38cfd341e703d32084b365838c6140fd
z693f8c02d0590babb1a57219de6cd78df8a9b626addba508ab460f93009768a0008679d917d926
z66a72b253dc39a109a4276ecc59047a63665cd9298422be210ac03dbd1cc8644cc19c503ac0925
zaa9c2ad3d4d74a90786c449f13d675e0c775238c125ea8bc2cb7499ba4c6e41836560fce21ce48
z293b18ae7f5ffd9b001e61b67efab0d424e797fc8fa0e8ebca25d5453df7bc0d61d45cf66c280f
zbb7f73a029d275f85e1a65db45d57d496ba66cd3699fb4a7fcd927e639dbab355d7383a4323384
z81f52f0e16b745fda11aa0c03ac31a8e9b7ee538884c4be6e20622e393c6c15f721f71e57d85e5
z8a7f5c85c417e2b07c012bdf9efd94f94f7f9b30f55fd3b62319a9abd345bf4a2bc6cb8febd162
z81f148a12acf779c058aa11126c667081cdf9dfcca7da60407a59942ed579992a7a06199c18b8e
z5184f547b2ffe3ca89b211a0c3bcf068bfb50859cce9ce818a3c7dbb386e1fcc355dae712a861b
z04ec3fab6d449f33326c0889d4932b6d7fa1cf5e73ebb8767330395362a72e9abbe1e8f4364214
z7b381f0c6c19b4ef8d3d447432c81e50f9254d281b72d303c96d751d9549e59c3e441c04751912
z73fcdfdfd519f1fc4857a73ef0f3ae4cf1fe88b1f29b48e0f804408f6833812787a1b222320f59
z1cdb587cec937e519bafb61afcf6ad3761bb3893fc6bb0950945ea435945fb00588aba56c1b390
zc2cd48a6cf38853d73fa6ddcb78ba8ffd2cdf56e32ad52930206cab5bbb8b07788320476abfbbd
z6ed57099db606349cf1aa77b12db80b3b727645ebfdfa33e310b11d48255586b16742c34ac0697
ze94ce435e11dbc9999614f5c3527d1d0c42ddb1d41b36ecfea1cb9ea7d4db2e4f0888c1fb47fe4
z107f5baee3c8e1d955900cdae72773b08ecc4225b668a3b25375e742faea3f2177a3b01f58626f
ze49d7d02a2a971143795b1622b69e5485e63c80e8a0549f3754aade14a45b6514cbca0e054afb8
zc9aabeb8208f0f14c421d29ad951d5e913b682999b3dc96ee2818a8bac2bf7c1cc59b3f8bdc4bf
z93556a3fcffb602567ea091cada2ba915a6bf8c6467774932b764b383b98a8e6f0400b5bf6758c
z851fd23e04f54d15f3d652b1839c54c213e749e95547579e4ebeec2dbd3f5d3e7738204b22cf7b
z42be45f11e207238c7561dba23072946528ccd77e7f44a08bb02d3bd26eee12a815f2766e7e1a9
zf4ef97364cb172ee5d6b9f918d4b9e5dd8f5262ebb4a78d301a6223a1aae6373ea6e51af866099
zaa1d611321c14664b122d6cf1663f36182c3d1b220c906c5b571be10bb3c98c549d08683b1a5b2
z93085355d62d90b3c72a3993176c101caf67e310a189fa941f9958ad75b1dc7f50fd087b0f49b9
z60d3547993a4a72cd251cc944b9dd776aa07d691866198cd4c079fae27b2f0cd9971ebb89d27c8
zb016ce6e379d8d47087e29edad71e8b9089df77b4cccd4d710d94599a479000117b40450f8d748
zee95a322ace226ee2e871a910a1a6a44734a37f16493f9cc1a09c9d69d0a5684003ddbf3abc8db
z37dc7194dec1ab90630272738758e5a28c99fb7d660e5e2ac91e69b9b4099ca5e34be7ad260f3f
zf8080af7b77bdab32054c63272d8ec2894697663fe96604ed3f1b11a58f6b76f9e1aae41d5f162
zfed127df136fc195b0119e60bded4f31d764849b3a26692114aa76b04e483b47f9573821dcdddb
z7c74657b6010d088c230018554b6d188d7d1d389b46d3a7049865e9076f7fc80443b355f982397
zc48840506e82884c670f11cde56af12cff6298ee14bcbe6a2ac5a622b9443b175dce007c0ecf9e
zd24401c907769edcd3cb64213af5f75ea59cb83cfcbc7b3fead133a36fad5162615a238364d6e6
ze50fac3cc7bc66b08a9ff5b877bde7f8625eab0a7d75c224076925624e90b40c96fe237e6e36e0
zc43a154bfa6e0c233f44bfa26fa7df8eae13cd4a3e91e81dd95baffb6ba2d0007e23e42820c5cf
z34b4e5bbfbdb5a51956b636335d94e5f186d094a9105d359deacfa5a8647f3f0410cf534b2a1b6
z0950123e576016cdef7bd2c5be5acaed30a32c6347a524b140e2632796a28a6c7c9c9d28e062d6
zdd405b5cc40f8c7526401f7cf0f21fc0c918d981604c31d8b48476561f3abc8f6f6e4240c0aa9d
z54221d06541b09e17f276cb2fe3b1ff1c70dc0e99a15e014ff860bb76c9840ed6d82c9713a36cf
zfce256553a644c466dbadbb62ab57b89bf5e2ad497d042f0ce5fc5fc2f0ba16cc39b559d97a42d
zc7f5e4408156f9761253f5446fbb908437b0fbe39b97c558eacc2ace8d24a29f1299e3924bb42c
ze2069fcca6ae319d48328cbab4078bcdc4e469730e04277d5b8582692eac15c8b4332306195549
z6d2b6d85bc11651a3b6ce2860179ae6ea4b54a0752cdd7d302d0c3f4854de67f0a170bb4cae3b1
z7963be2c1800f8f1deaa93ce2277670e68587f4198f60c1883eb2f36373088b529d0d72d8478c7
z7d8297a286d94e3a44f8edb5de543f9b3ff5fcad641dcad4f22c6bdfbe4f0e12c440d2dfced6c5
z0197c9f94b75fbfe989df8c0fde8530fa24f639c19ac444256731d8fd9f3464581cf09e43121c9
za884a8bb014c484f879dafc863a622d052485555908ccfe9d9cfb6a2854248b5e1b044b309d744
z7be6499add5c1bc94a899a9918d4e2b0a07d665b9646ae17e10c0892911a76f1141c543922d8ce
za02248b710d4acc5ba3789a87366d99a8b9ac8a9ff831d623ac0ea5c71740ab96a7c97b21053bc
z1d69d5389e990b0cd539a53359ceb1cb45c7799252a901f4a43138820386fc9300c0bc3cfb225f
z901159321afb29d6f12023e2a0391be95c43126bd91e32baed0777ff17af5d4a15f8c793edfe57
z182365e6446bb932825f7502cea60b05537c17c1545c18437bf6263fe3c5f40f49b12875c58ddd
z32ca22f9df4a0074e73791d393494fb17f53370cc56e329ff5ff87b097b8f32341a44c2590841d
z7f566e6d9bc0d7cec1f52eec3a71783e949693abc3eece13109873e78760ae12a22fbcc70834ae
zfa1aa0bf7c40f05b301705eb9e05a2b00ac371d368b9aedd65633b24dbdcabfe618c0f73a46d1d
zcc6f6d846c0bd241a585eaca40ee3b2cb19ef4dda5f7d131aded9dd3a6c2fc6f89939b8357e7d7
ze60ac5e00f5c534fdce7a0cb2c92998a9349b337e0353ad8540f58bd4270eb9df4ef91bcbd2b47
z2b125a6230d5aa6aea84ac6684c64ebd0f39e8b42cd152a712e31ac5894780763c071971e2d94f
z6d413b95974e4c9c059a4e7881b48c47ab7517911b4fcdf7b52bbdd7fd46d858ee8b022702fada
z87998091be585a0dcc17f1747df808204b817175e1789caf3f80aa358d12a85debbc59f5eaab91
z2fdf4cf477421562d0039b743a2f128048c8ee1dc5471352483fc59bd5919a6af6426b172ec9ff
z4270db616aa3826d6cc98502a6b1163423ed168b32b9b363cc3676ea71cdfb4927242ff39b6fc9
z2dfd6c763571515bdb83ff31c5a293fa97a5082ddcbc024e4cd267f6fd7db0b829325ebd4670a5
z45ff121a6735cda0ccdc1798ca5a4e74507715e1b827c0e48cc5fbab19042852e5fe9e14adff06
z11f2e183341d71623ba1b5d582bb2d4a1ede8879423a2520d5d25c4903f0e5b47f1f7e796d3ea2
z2a533ef6d2aa5e311e18a92d9d931851267bac62b9bb6621fb4191c72c9204524466e4b6240d57
zc130ed7191ffbce558ac2d0ed16ac822c9e457af8a6f75e8e0e73fe9ef9256ec89f07447e2363e
zdd00f2163ddc40b174ea437bde55f29b46bc69ecca8d4a31b867c4567d28cdfdbdc8b4e5810311
z7509ced88fc2b6b106eceb1177385fdb603aedbdf4e3c1a681457df9008afe9aabf23e4b951cb0
z80e544ef76adb394c1dd7f79a890e908369262313da57abbddea2a25754bc440295ea7029ab288
z9136bd53040f7c086bc4c478bf3a760f6f24626e7c2693de4628061a59e4f48cb9c5466704310e
z9d50fdc8d1c6146fddf6c8be707ecb24f257bdbad8bce34d75260ffbbddcab91b7a4928a91779e
z39c5ba2c99aae695cc54e0b222976591582ec118b14d152332b594299780957c373288f784f49c
z7bee5c46dc6404b2386c4ea36ec6294c263aec1f984f65e0afd1408ae74a14ad3f7769e15c4bdd
zf6b3d9d855c61639174f5b6810e694eac8f88ec7dd028a02b554e4635058ddd89e7ff69642e110
zb182166413e39cf0a95181b82c82400194b749e429d9d95ef2bcfd05e9b00dee2a8985c90b32df
z5bf60039a7b522153fc8ad507e9202a48f0cf8e8268b6f8249f84e6d33b59790aa4aba3e5cdd1e
z57d2f88887341f0dcfaa6e4ce733fd7d19b099c43dd06d18e9e4e2a2b05f26b9b6d01e608017a6
z1ef48792a5bfa63b17e5fc3a319633c5696e7f3b88cc0263a2dd292cd3b7ed1c79b681efc23c37
z3f45eb76218ea254839ff0eaa77fe60a85023d53aae2ccaf9721b985283362ed79cd2d8e9cd569
z9f3a381c592368e69f6026fd4d1193678e1cbdd5c4f6a982536f8292ce58f3f572a7bbc4b7d90e
zc6c4a3f16af0394cdc960c9a1a0803df91f23bd1f4f94bdd459653e8f1d71d0fe01f2ab6f7a938
z9eab49062ffe7c36bd317b90d52955235bc33907e88a8371d27d200e884991ac4c0d4b25482178
z84323febbc2f8950b62b21ebe840411ce43be7e2a048bff6b1378693caa91ce00099a0f71c95b2
z2735c5a4cc4333724942fc0b3f838d657a0444ec83f4384250d16a6888c82681f2b13e8f8deece
zaab4dacb1f678266c04eff902ddd1f1e26f2632f8bacf2c618a17bf8b8ebe5e24b292482d5ee40
z3a23d07fc7996388152dc62c933796b16f8c36fa1b6b043de65268f7c5ac5cae3b6b8edd734b39
z2cf27b2c44032ed218f234fe2fbb6cd3549fc7e52390363de8f185beb5321893705dc62841456b
zc17736331b8a0148bbe8f398c350a2d7095fc37a14a6c720be957cb7c0f2a01e729e527c5e0845
z14d6cadf295746375732f4aef82e3caffed2e026334579047ba2dc8017ebda58982f9c6034002b
z00572a184da6c72f553e06edb208d98fc6a64419c9f372f5498e463116eb8511da8da72e496a00
z92b7b33ba522fe6c5128efeb333105546e5276ec78111c7fac2e5a8ae852864c092971f9e6f5e1
ze375dc4061098681986ae44434c4486f42b7a7d16f3062ddc9e09e5cb5d8c1b0a18012b5cdf9ed
z1a5bc559c065eab1850fcac03c7f982414419bd73d3a3d6afef20277746dfd27c61fa9876c8c03
zc64f7440aa40236b621098cb0bc0c5e1397b75cd55a695d83440c9d3682e4c71e7cc615ef0e0da
z6a08df5dad3f025c92b017312e9cfb9c0bdbc714892982ea4e359677852abd84d370f148a5782b
z5e8b1d195ea3d1e0ba6fd879a84822248c7cf9cb8bb1dba0da9defa3e3f6485b62496b2e48df28
zf64e142c184d8374b5734476e8989a2c83918a8144084bd52dcb6ec435dbce6b6f0a3352841c4c
z4ad3841795eb2e5cbfa894458f4080e7dabf0e2f1816cf13eb96cbae63e3e82d56fd0ef8abc98c
zadd72b5e09ad3cf3a69b983faec6b1e4fbfae226b986db33b18219e79e206abf0ffd1d999c17ba
zeff312e428a22d199fdcc4de8b61e5422a897e68c20bef10add1c06bad8940e5b9ca9064256e11
z7475fb49d24b75ee7ae9230307847c36416d6cf6cded585e847c264c0689b92d9f485ec7b463a9
ze004fa043b4fef9fe9875afc1166a1f106c86f923bf1ee7ac0a2a7b5786ce80f601eb5905c0058
z4d0ab4b9bd64f8e992ca78378a9552904000848f2fdfffb5a907501943e6219be8a9149ce5ddff
z006d31e439107266a9d82ac7dbeeb546ce5de1e406063bbadc3ff69ff0b765d26ff8606c8c7b25
z4ff1f735b12b483ed27e9c72f3fcbf1f685489fe33bb4feaa1f2b9ca36ea3dbb1b40b617cf3d31
zbb339b09de496f27d8133dd80c779751f8b5a7a07bd335b435e3e5d0f2d7ec1b9ab08c48837d09
za5ece2a334e5701ec114630ca9e6891b9f31906fb36ad30ed9d3bae0c36b364f1b2040263ba314
z2f2e9822f1a7d29eec6eb5c0bb23ee0eac936979556fce766beb9f49d4d5eb1cc6944d9e21e2ba
z5f365f82f2d98381e85cc1ff1e121d1b0273fd22e594cc480fe3ab41d724b70b9df023cbbf7b0c
zb98c77ca1ecea7d18932deaf59839718c8c2db1f4c2fe65bfa0b7f51624bb260c6259eab9667ad
zafeaaf8ce6a7a8aa68180b30f72c95c9e98446c19495ad172f2f7e0d276bb10e69128bd38cfcb4
zde1bd398228301303631a5a2b604839c51e40069ed9ad36479cb7f350041919fd20adff0132f54
z05ad153fe3e7e95aaec5c13e0adf6319b327b35c8b2171bee548385186fbeb07e9acb34f104a82
zaa6f6e1eded3063959c5b64151a06beb044f33deb0aad3cdbd2f2344a6081f9f39210088d29539
zbb91eea52da60f77041c57266a0aa9989ad6ae87fe354324b57a335085e2463c174228273de112
z3f24ef62964b1a0d30c0776f8ef9e892a265a1ce480a7bfa740d44ce5cd4968ca55cd633dea5dd
z4c7ef0e6f8481b119e435d5824c859a017d7aa54ab9be8c5004d535b8f43d35fbb81c51f2c5b69
zf687973f8f5a8db8fa72702be6cd8da1762c904dd5d7fef3b7297150a2f84bb539ccb2ed6acbe1
zbbd4d60efbfb099ab4c6f124f0b57b0d911c84fd77012cc50957c1e8c25673cb6ecf3a7f7f8f0e
za1890f56b22e3fbbe8b972c1c29ba5b13534f12ad962973a3d953cb2830fe2bb5724a11f02fdc1
z2420e737b6aa272c809bb52549b115f976a2f085b4a48c671a2a52e39f7993b7f17c7fefcbb53f
zfbcfba65bb0aa210cfb176bf950d9b2adc368022a72f4aff50b89e1103ba08fcfcb43189d5facb
zacfecd5bd43daa9cc662e7ee94c8aed77045c4c5175fd31ada99fb2b63b20190e2ee2bd3d30d76
ze790a39f43f8460a61426132c04199b0949f8d680d4d08b87d0d22414381ef787779b25a120b05
z04bf57dedd23bce33f96d310bf6a62e31f26d7a9ccee99364392a9236164b379339926b22bdd63
z9ac2959dbd66a7d1648f3429aa0494de29b37b20afb2b14268b829059a2fe858126273766279ff
z3e93ee90ebf971704082c526622ca92566256c395cad532b2ef2cafea3b6054b68d0d6b72609a9
z29a124e6e9dbc79fad79383bb1ff128f138936ce8406612c5b8c2437da497a8fe14b348f2c55ca
z5d02628aa795f56f555d137c1836d9bd519b08a6e4330755c13d385c3befb31e5c7d0cf69d8a60
za4f1363affd407d89ac4d55b2a14d7123d9ab63f1b994a03c882d38d652b2651c0dcd9e56ef742
zd18b2fef098fe4852835cd7f6126c9b690dd14952a0aebd28d532f4a8ed856f33b9ff189d06558
zac6eb77b6c07bc9a17e424b069a33527c56dfb1523a753e7981649d26cd8027fce84b0287a8eb7
z9467fe7cbf55f6e036ee3a37024ed014a33b12c3d58feea6fd20aeb338ca6c0c0d85f1d91359cd
zdad815f9441d7d02273f24593c85ba28f25c6e779a4369ef78ed8a3f8ff6a79eaf6398de5fc41d
zfddfec0bf043ecb7451ae55626c4ee075b5ec182a1f7d822c4fd732bc6b69f556f494ab40796cf
z90879c5fcfc82e68f278105d9cacb4ee1650beeea3e8f1adf9b9f8e19e373959bf923853ab4ec5
zc5728a5d2602b95b2f2c404e9d50061434eac4b03891a19d39cf6e7dec55462bce6cf81a021dee
zacf569280aa7c396de8f4f1fc080fa9b7b590a573ada482396c8e6b01dca592023a27b2d6a4464
z70b43a8fbe46609a8eec24d1db51e75a3f1e7d6b6513aa8be2ca2c71c9193f301730d76a4069d9
z421e1761899e7b0169d29ba91c1a1cd51a39bcdc3875a03010383167a7df44653c305b173cc934
z4047df712921ca12559b1b98c52248eb4be09a8da943ab801eaf50b165bc382d3beecd5728a946
zf8bf3e041d9929fbd5942f5af03fb329e71db9cbbf3559089e7cb8d586213d58ee694f8cd7c8aa
z44e033ff2a42106a7fb6f72197b1422439e1c0abc40413e5de255cb5166af139bc517988c31077
z62492d6c5d559fde00502b4706daff9690c33087d1cc2f551f520a77aafced05f7d523c6783263
z12b23a3238d284c567b56ed93b84b091d700a8f21374e5ff20e99c791516f2c19caf8566f2d86a
zc29b28e50a4a0072d09130f87fe713c900f10b384e222c1b70aca2f3220bdce72f84ceda421e3b
ze6bb00ea9389445678b62c42b2f378a3a1ec728475e3e398ecca6fdc2b016690f68f732a0575b9
zd0f846149ba42a1f31770fe63d824e62b6b74711583edb1a807990f827b7337d5a10bc8239dced
z37eec8478537194cc6d8300b2332959d7bf4c4a532849ac7c88ac156b69a05743717fa323d044e
z3a7fa431c534e8bfcbd8608ecd8569f0006213b153ecae1e377c85cf53f81f53bf23be451952fe
zede6c3510e06d0096ae40878f6dd74c5ac8b45256d182646f7fde62f480d69ccb4d88acd23c819
ze33a5981998d24b4d1715eb6df7e5c4aa30ec56aa4bb3570b46f4abd98686c2948763c306d91f5
z3fc146cf2d03f90e81139ea8fa21399ef630a167520f4e35b6d91f20d7e72669c06d0391edb0e8
ze80b5ed0b65e083dfab5c0a0b8d3318b0865698aee9df13db95f3c696e1c9c9279d24b0b45ce62
z01f10a0334997acca9d9c0b08c13bbe5d85c492ba510a9aecb53c3ac6908d09895471678c42168
z67a6b06ac9bcea7f9d3043bfdb7fe0ff65bf9f3893f61b77d0ba008902f6bd2f95bbb11b2caf41
z748b39621eebf130960179fa6ff95442189da7db539690d1c341579e67de5e685a93be59bac80e
zb0c9f0f60637a4bbf63519f4d0385042386e2764d49dc330b275da2502bb445dc27f27ea319c42
zbfa2ef6aea58db074ac951cc52d4845633b0a3f72463bf0201d50866b1b05cc8b688340a3b8e6e
zddb8b118227f41e5784020def405e9af0215ea11eb63546f5ca461d43a39d1e668f13d0b2bc35d
zaf793ce13cfe6705586b19a9b842a984508be5084146826fb18180c68f109ae96b9f30c59f9457
zf44958d647cbf459a744e737fc0ffdff4cc6d2b8adb62d69b2a6ca2a72541fdefcc1a21ae17943
zd43137e896afe14b5a869b2d4e37dec54530ebc27259de4fa9535e466c57dae3d9b572463063d0
z157fce35f77cc3b53dc31f789508113fe2871622dd270ebd841bc29c20e220c1b66e88cbdf8dbb
zd58f668628b7dc95ebf87c3333446f72c200090c20a63909b051122de433ab7dcb4afd9d99e9a9
z42eff0a32bbb417028aeca07dd92ded6864be775c981b4b1d0e0a93c8ef0713bad3297be377260
z770fce582884a73a81a4ceae8d46c6c843bbf16b527a6ef7d872d5d1b08b8253b76236f10801c2
ze132c605e5b051ac054511679d876da17097fea13794b4406dd76647b05a23466c7fb7420f77df
zca510857c89925158f9692f3115309b100d9eb05f610c9c49fddff408474d91797782b9b950678
zd05c9bb4b612f27a5ac020db8d8a9e5c09ffbbf2f89137d5b92e16795a83d69f32f2849868186a
za13acef0bd5c08dc4221710c4186c920d04bcda339122ade86726db72995ef80fe2d35f90f754d
z48cf406f456c6789b0ebaf4101ef0ef1f9a169a80c55f263ec88f9f3817e7cf8ff96e929cc20de
z4c3e8b5e5344d5cdc9ce6b1489bcbc962e8da114987d10566307e95f0b2a878103ddee0e51cd42
z9dc1b8037986bf595159920c67ff1dfba82946cdb30b75de416ec9b93ba2459bd1577c3c38b08e
zfbbd22da7f31ca504e67484537036d3a67f39afff033e0d2a7a5ed1b40777b943cba04cb948d12
zbb513bf1e4a347941740529c26d3dd860ae1b565d4b922cf12f3ccbb7a5797385e6c537aad23da
zb12916a2d7e99ba35f7bb85aea4b6442eb1c6198ac5bb7ccfea0e10862a630e611d877498a0ea8
z8da78fc98e2a2f10679c216fa89faafb21ff0f15b62ec77d77fe49e5693619bdd56b775f7b7901
z72e57d6c182b2aa8426f852c97c2ee3603c842de00673d7bdfbeca20f456110ec4be3363ec078e
z2611bdd86be80bedae4e89352c9d33ab633ef630ead1c0b9a3800d1e27e3efe82fd0aeb360025c
zcaac2befcf767cc210ec9c1405605f68b219bd4d7804c9da440adae1531177ca1e1ce3c76bb7af
zdb25a3b258814f100a0b2e1f26efc32a02168feeb61b03460790c1b79a8ceeadcae16a812d18b9
z60deb847dfcccd532209b768c9694f688b137ca8b4d6b2ced776832e69535fecfa8ff16d075aa3
zee936dab2914dc91bfae50fca77b4ae1aacca57b490ff572fb5cd2a03287a8e077ef2a70458bcf
z5abbefbb79ec7ef13fc5ce2b5f88453419524f2e53703b89385465c7170b026e4a0aad2f69cafa
z82eebad7f671a25498c807fc3ad08a85644dea342d75ceb2589a64d21239f704960bb10664aecd
zc73f675e1384aad4262b8a33eb7b9adec9cbe96fd14e6dda0b25faa88522d6bc63305e7e18d80f
zb105c3ed80e04e1cf5b7c643f4427739ab62e49086842338b0ff39b0ce01f82153cc5d1a013e54
zb054c78262536ada83dd5c56cfa8b8f65c20e6250027695dbfbd18ce92ee29597910768d0b93ce
zcfd6708953c21d49d951ca4aeb279d18a6d6e7c141bc5fb480de7d45b06fcb79e0451230425d02
zbfe7cc966601a5b009fe11dd1ae95ea18acaf81791f5d29a787da0ff8d03aac0a86ff945aae593
zc37642c155fad16abe14b76dcb39bdad21f6df2aabf05d862d9da7ae55472e2533ee1d8df07055
ze8fadf33c21577804bd6d308c0f167132b6cea848bdca4d13ee618f7a9d974652edee54deaea5a
ze411b2b98d0e9f31dd6e35705563cc417348e4971e0be00835b9ef2eb7e26f301f7ed710dda68f
z9a5290a5bd01a5b544339a1faf7345ae9de3019e504c6641f7bddd908bb839437d8c8e0cd1ae53
zb93ea27a48eb47c12396a9e238b60e9f682bd683242c517feecf16ef9bb842c2def276549e83a8
z3042a6f1bb06cae75fe0eb47265f27395a10e4101a475c858088b92cd7b71809d1f651bf3cbdcb
z2f89d89be31f369f468303b6d79f2495499c98e65d37dd9e33143c84801d678bfd010dd039c0cf
z7f6d4e3642930ed1f4fa6dc98d9e52b2b37b40ae56805a066d21928c1d7e9406ccf040b7f0ff68
z51097a0c05fff994d5e7084e7776333bc3413efc92a11785cf0da02296da84e6e27f5e3bd21128
z9a7c763b75964ed41501d12620ce4cd7999d732d1fbd7f00e8fd2fa9a8eb19885c760f8a3af5c8
zaee767a709bbdc177d7b58d2d0da9ba473673d96e465ca616bbf56f995795dd9990324f37c1c76
z9ecae827c7cd4eb88f59a74e98456c92ecb063540b44cbee986723fd1e1a062e478f049365d99a
z1592854bfe814b605e781945a0de2623ae0233f422d83d218bbd72344f530f5485efca1821bf00
z26805fddd991ea67b674a73c8e81ebd56adcb7c9945261c64f1531fdc61c50eeab564c3788869b
z9473115dc2e0d4ad62d00b3abf4bd1e490b5013b2a2f364809a20e70dd183978c93a777ae8686d
z0f366cc22aff6b467d3a2f450076da8b93f568f01ec720e02ade7beec9d6c83a5d92949d81ee85
zd0927557f99c244a9114d9fb5e7e2267b272fdfb6a0525ae8d3eedf36c2daa472c1f76784f9c70
zab29916d7548dd6e5d547fa7153fbb3fee1ed23d8d1bab5a99cd0326248b668075e82290a5aea5
zca24d759dd00299a7fe1f60ec8db831f95fead6f978e4b589c329a84b6bf9a423d5aeaf638693c
z40228e44d7d9720f4e52da2cfddebc55a75f6dd52d3fbbed8585aa3529d352a201cb24364e34e6
z570c3218d45e4d09916139be1bf867cf9ed7aa8e56dcc3c76d0986e2eb2ef9d9fd1f5a51464e97
z6a0ab806275b67ee8a7b2295472fb745f2c6270b8161dd2415b65bcd70b288e8ae4c89b1bacc6d
z48757eb112d788e43673d7a9415c73fed7d447fd017a41ab7981129033e6257364238b1b2f3200
zd6a22e0fb04d7677dc5cf5df310d2c2dac4c93df5166d33f0e3fdda0cef66b68f9f20daaf7fcfa
za723e7d673475523f08bf4a108ed771a4e6bdea5a2b4b65758b3042561b098eb377ed1ca2da8db
z5ec44be1a10396b0e3f5db425182412e0e4509185eb9146a50635b6cab21b03640d50a48a13331
z6e8a11ade5f3f45f3e6f72e7d4aaaeee181a701284fec9462ef3b12b4bb91f6e75564153a6ebd1
zf9d677f1c1fcaf647d2ff75f0304731e6df22ddcab3237a1e6071038ef5a808c71475aec6fcbbf
z87956faca0690d49ec58574431f62bacdd400810de97b4a3ba9f925bcc2ab1e676ba5fa83e077c
zbe389b7fbe6dd0849c6544d8ae49f39b778071c8ebcc80f44a5dfc012e1dac3f1a06754d092c5f
z2a4f6e1fdd3e6e2b37a34bbbff529ccc15d4a2f39a0a800ae4fddf74172781b66d4eb80f0076b5
z7778e4d0d22f4de817f937619408bab41a7c642c794acf30b5e14f8a07a119928429ebe7562e61
zd157265fd75f8b2b17a3d37cddfb601cbae0f1788a66dd3b994d557b56e3742b693f290e7fc6a7
z77cc6062add6bea916e00dc14f6f6a96c85c6523b03f576036e868dcae218a9750a96a9857ca8f
zfe05aed6e42afe0beb53cfb2d743b846aea75ada8d1ce0e69e033dd94400d99b36d3207ac386bd
zc7b0f93780cd2bc15bc6d362002db2a319e7f09a0bab4a4f5a5515b0bb0dcd46973d99b14b9d2f
z4930d2aa3fcc8aa7b3fc14f27d3fd007f7809e4ebd3e521413d146c28a818c13a35069214b5a62
z39a5b18334fadd31fd72e7b96c4b3d36a8ff81576a3de1478984b79bcbcf3728a46711986e3568
zf49caebcf16211fea98f8b24613c1ae82d2d84bd132a036beee28846861df7362b816de2e9126f
zd4cef651f1f150a5fafce95b8fe9deac8719e31a924aab3533ecf7afa28ee2ed43992f0b40181d
zc7237fc018b5c1e17bdb3b89ede6d1d87c12b34e43072747d2d10781c4867f30d13dd7ac78c839
ze935eddaa24c3e87fae73e6b8695beb4c067cbff0f1eef5877451fa963d129486b80c0e98ba2bb
ze9b9e95ad883f1df6ad9d3182e29464337b33f60f3d3a62e9acb613f953683738d11fa5427822c
zec95cfc79acc9c52abc88e0756017178fc85d5b9b66c51693a6ea633b3eb6482ea846a32984ece
zfe5af4c79503bb0187564b2fa3e3a38d7535abda9395fb5cf5d4c63b1932f01e36fa1f7b5f8387
zda89cd1a161f0b6e56dc6177578bb69a8b7c476522348e1734025f613028e2262b3b624ceec248
ze0fefba39bb9141a6c336635ddd8fb154311d13a2f60acc8b01640a12016bd232ced4c48f1c5f7
zd2128dcd5e6436ca0230ee3203a74678ef1a5f2467577190973374eb4ba8b1ca8fc83bd3583aaa
zd72b68fc6864688758837eac966e54263aa92bdc942834a093840127ef2bffd90d0a9b789f71c8
z136713e916fc73bac0a9c481f0c20de3754b9c2e2e4cfcd6f0427c56b166c57153a3f6033d5e1d
z26d436b74c92d3cc995f81c280880889dffe004ac4f2455bc2ad676cffcbc9b893b2353c611ed0
zec24db40c36a66245d565cae73d24c61d8c94c09c7cd2e18e69fb6e580d0d7aed6ac9c1c1b4892
zea3bd7f544bf2ebdd99c8c74fd4e3f6f2ad169c511dd23c5492b0b9f1771e5c5ef928cd6c962ee
z2d328edb59094b8f5fa7d5fa4c7b7de0150e15c4ff9f8379bba724cf200ad2aaaf26aa9fc7eee0
za032a141c0575cbf7942e8874691125797fe19f2372e3dddf7ca4664e6158defff5ba49c2e9426
zbc44a6f9ac6e69ee4b7f940f7e6fced72bef9799877f0dca3e5610edbbba809809046bf38dbd2c
z6c4ffe7646f8aa3fadc2b406d3df7758c3776cb08c2a8c443ae52cf4f81c11a12a2f9db1eb2b64
z01afeef4441a7e115491d90a736af080e9df28269c8ad6753754102233b9469e96ed4771013cbf
z5da570581cc2ccd374437ca60199e70e1f2fc4fabdca09900981084dcbe82d98e27f2fea13d9b9
z26b53a48fe81ed7f35e3b4f9761957fbd29ae8616ed8028fec9a6be5fd5048f6429f27f001ba18
za6d456b950f4fba656b3bbf02c52a1cc7819286005746b2cff883e64a0911f4887cc268e90a783
z18f87d74d862586203b8ac20cdf9913bc41e534ef893e7f13f9b727ecd7c1f7188f23c231e24f5
zc734ac97f2be11670e9067edb44bdf42a128b6f065a6228872c12a443d2557708e9c141e84b24f
z2e36bc3ac94a677e17262e74971bb2e9a1a251b76adae1bdebde2f05aa353a9237695add3df1d4
za6f8673f6906e16475eba41eb447b502c5a19e1f49bef3dd0f505d7232803fa0f022f7d2c14209
z0482600ea75a44da306c8558858aee441fccc95011063b995c8684cc8fe70d048a3fad5ccfddf0
z046018d61fdbe31a720e44511d18a925c141e49b04da48101d9d5ce3c4947e7260d7e82f5ddd29
zf8b12f85f243e410b0f925f41d18177a4756a85f6defb74cb4f6d5e94afa8dcc26f1248481f407
ze72928ae33dff6833ead6279e4a4affd7c09ea9730ee5868571c10dacc0b14e5b3e6d0cd13bbfd
z42bea0f118f63ded149f8e03e47a9675eaaf531ad88765bdb4aa6224d4b93e1f341f63375785b7
zc1ded76dfe010de5414c7182d59e2fb1c4bce987881309f33bae052601238b099f1f15124ed145
z6e3f710b2d0c54af1d17a4207059a62a6c2c99d33a1b788ff0a65192f5906bc447955ce031bd5a
z17cd6eb2a5ad8788bc57830f1b8d0484134a6ff23779caa3d1e9ceb78e6a963a135e002a74e831
z012c9373ff05d927680c60d4af15eb541e23b2d3a71bc424db1c0ee235b4357013ba7b7228bad1
z1ad32ff0abfc162bc98b5c59e15489273924b44e8e519affd7607efdc8a7a46b72d6e7ccf747f8
z69bce3761d3c7c00929f6f80a5288b2cf49ff6e0f148c7f52d9c694ead3a1f53677d37e88cfd0c
zf443b63a986f96accc3d65ad1584c2a90c04774b4ad94360310dc91f681880056676e456ebf543
z422efd92a4a95cd492d5fb628998059c5e4bb6c594f1f66e8d1f6d487a3b1b181393962d5aa27d
za9ae592a45e53988be570b1694d65ab21b81c8ec54b911965b25c6bd7de9beb39d8df30534108d
z403b6841153098a198e06de779e1ed459286147d6660ab53f3adeb6cd7c2a2a616f77df7b483c3
z0c9cdc4379526d50f2770d159078de0798eed246a42aeecd282f3d74b5aef82c4b7dfc7f006d09
z95087250292311e90c0ca74d2a3cb8d3a3db5893cd1027348ab84c40cd11f2e63ab2a6f1c5acd9
z7415f6c39ee90418492f8490819468f33af60d25083aeed5fcfd1a7d593484b6179d47bce7e224
ze039f1b102544f96c717da341eb71e469e5c384dd99f8933244111d78cfaff01b5e22aa7c9c74f
z6f79a6da2641d4c8d944d5dbecf35ea924a984792fe125b911a68caf1da115dbeb7547fbe7ff43
zb0b8e73b479bfa7996e61e672ab3687f77fb97ea1c876d7bce158ee998fb83d660298817a7c8a1
z6a9ec725bd16f613bb76d97ca9c36cb03255a8b6b9b878fd59d6e3d050595a5ebfcb0d258a057f
z79534894f76bef40369b21a32fda1e5719d8ead2861958aba245beebfa05b7d0d2ddc0370f500b
z074ca146ddba79dbab57bd7ac01f2acd85e08a511906444d953ef411bc15025ea404e1530e4b48
zcbbd1b937cdac3fa7ec2b88786808dfcc1fd2864e91703cd70b0c5c2ea2e5bd12aacde2dbdeab3
z1c38f0d269bf7baa88d110146ffd3c2ee3975ad0102ed5e1cf8c74111fc2e8e482e619cbcd7735
zdf797b7ed1ecbd3f6bfa2ca097b39782606a31489537d357f8d30d7df2d5f189f6fc813fd35b6e
z7a7fec95ef9bca50c2f1997aa54f3c74b3d93320a7bcbc9b669c35a8166de7fcb324d2a86a7002
z5c9184e305856ca50ef17ad65b5e8da9a031b8e57ef7d4698cacbac2ff0cb54bc675e5832bed06
z8068dfd7484359cd7c6d741f52e7bbb5ffc7952292f99583ef8dfe8233579230cf631b73eb6f95
zc0be410d1b1054be334519ea26ce6c11a3803a9335aa6bc29792f5be998d964f278a0bcd79606f
zc986ca9a07472442d64032497d3d4f5e96a336ad5f055cf22a2eadec75bb51a12f96bf9386d0e0
z44f91c2deadfdb9244c934bb82156259449d5f2b9f83fcf6450fefdf6d8b0e9c87f275521ede7f
z477ef2c04dc1d129b8920f9a911a5eccd7d8d3474a229fb37ba456534bf5f5ee37bc88ede487cd
ze97e5be2a5a0e615c177fe2ddfbe3a521ccf45d74d4a88bda83d70da4da92cfa8174f974cf963e
z4c722cae31b4a023ea52ad4f080ce4af08d4e5e926d94c8c3c3d3fcd2f79d31b60f48937695601
z5106e5e5d3c5d1e1a4da9bf80a84ee72c1b46db3915ab34fb2dfb42f82d271e568c856271127ee
z9a19ca2c33f969f3412ddfa4cb80841ccaf5cdb799620802d9af113aa43b970f5e1c8f5d0b48eb
zc78419c4445ffc34427e381a80fec9a6715d2c8f6c4b140dde17290426bca5c41331605aba914b
z945903b18ac350099a34f79d4ffde09689b4355bad0ff68be96f8501f2b04520824815fe057e85
za29c915fc95c78425fd2a13562783aa422ad7fda13893b28b28c05c3a1bbc4db204a2651953081
z7cb8c3dd058b6a4eb912a9ab224a9d043cf39b315793a68e765e5bdb7ea30d5c9a25bcd7f0b9a1
z31cbe2b27ebaf8e998785349338beccc0d7aa835868c35e66ae5fa36a943b4da8e8b9098b4ae1c
z4c390e0549a1209b2e5ec68215cc6a3a7cb38e892f5ff71f09e890ded083afdab35a0608abee5e
zb5108b8168ac2a3fe09e3b76d1eeffa9e7eb855cd20b67f9d71ab1618a6914f0defc172ad4962a
z65ccb6a8b1b8c4d56688535a4d58b5cca3ef1977d636db84a92c23f749a1448dfcefbb3591f889
zd9f8cc2c12c25e6904ab9cde1c86f501131093b217c3927993e8f151c9569c55d2c9227664bdf8
z9e6c6d01c0cd1f29a40a35fe37c12890194e85c93006221744973ea55a921f751457b2e56e64a1
ze794a87b749ac9ddf7f1b666980f5b73bf8b068372ba2034fe5f08f520ab6fb446778f0d7b5e68
z0033470cc0ae7b7cf6f19d9407c06bb3dbc7554fa2820fe10ce007f4b9fefa5bd77e07dedbd90f
zf48df5e19e22af10712acd7487542d31189eeb795e62bc392a1ab9fe1d930f821e16276b4091ce
z390d974be931a994e0559849ef5cf054b1be6d4390c1b6eeed2c6e876575bb63509f63380ec584
z22ebb3b7c2049eff049d5f13db2e53aa5ededc3fcf09a7ff8c7960ed9ce7678682acea55e26ef9
zfdcefde814a49220d9cd9f9b4236bfd6251facc93cb74b3192c77d6cc39586a74c4103407f1964
z1e5bb732f0fee7b6d6e117589acaebe203b8bd055fb9ffa328773e6d620adf3ca83560743c30d4
z348c28765c4f5d943c58d932e46f100f96f838855150f12d527613eebb80d4d61f3428159751c5
z6a1cbf3c7e4d97a6bf7f685acc2bff058e3978b2334cfc2dee66467560f035f5a43fabcaf72796
z2aa625c86b30f26003292d3e911248734a3c10945f34f86734a9efc05b13ef65034c53310fb36e
z2913381b9582a4e16bf4d154e7723f64ea0ba468e5b2e09c228c902d393cc6ed116ed728e1fa8a
za724b9b7923b30ff70b8cc041e04b9114ad7ace446e75c7e396164f0702fd1c7a7611338b2567f
ze62d70f7ae0aa44968b33e6db3c49b0c265e6430b3908682f9ff7699403501caa22146578393a3
z3b8a361410017e63a1b6c51fb3e245984cc3f1740b903e794147caca46a21b72dd313e5f2b23d6
zd415460a5b1e3315a3d797e8909e31a9c25a24f3b6c884915c3b2e0c7aafbe8b77509b3528bebd
z0034ba2da51c738e35346e59fb73e2d8c2b2a6084227bd639fd0941fead3212d38c5c5f42bc8a0
zb14a5583695ccde851a6f44afd15c1571257cff1291e3ba989c29bea260572d41174ba63e7a8dd
zeee6978813ca7b58b45c8569a1124fd5dca5ff3fe9901e9f86bfff5f4a87fa0bf3eb94a5d675ab
z0fe9e5483c6830660e3d76975a09da61e62ca78446bea0f0e49a49c608d3ee5de9b9c98ef527ea
z92d0e334cbb1acd23c8a4719c19a423ba71bbed6776abcb592b5f9083ab16e8fb6fb8a178c930b
zb956c7150325a31f0e4a560eb796dd1135df4a503d813f2f36863d0bf5d12c91324ebc07efec6a
zbf2b6b82ab7142f5b5b26f8ea0dd140d4c3e4ca59be7ae07db0ed00936beedf1f098c2cd0f5203
z856359fc6b3d1a9a434d47d2f883e364e75020f58fd6559cd8eb6b53e47aaa3da2cfd00ca84398
z544d224fb35357a3696e087a4c0752e704e603183907a8cf1a270cc3dce31bd96f98987831f631
z1f9ede825ae599eb1ed84fc9d5272ed2e29e2ea49f23ecc4f0e06e5fae7e4b2d412f14f774732d
za57070cadbfe52adfdfb89728609d0df0c3a961337f65b87dee2701c415dee31ae81239f667063
z51e738fe2c16b154d2faf6f76c7ea2a690ef7c391a827ffe1905213b2b2c01266dffcd37783928
z20e2505767ece73da03c6de11be8e7a2f470c6c96ef92bd84636faa68b433e54b61b192345172b
z861344d15b81bfd9c14782aa97f0b3a51ac6ee07864b2ea2e68cbfe2e528ea689a4002a56fe531
z66e06a4ebe40f17245bda1b8c58791e19787f6f13fe4518dec5cfcfa410b7a7c994b3491d8eb43
z625ed26e43a66b5a52830df9a1a799fd6148f2adb523cc06b4740aa567b8bd2036c417d3d70269
z4043b25ce32bd36cdfa4a7791bf16bd11d463413637164a15121b7322da40ebd7c0ec7af34ceeb
zc44e4d52aee7985c44d5aa77254bfafa3ae7e18397e01bc509c2aecfe3c597c51c8108951a6641
z9a18c8c486519379771969bdcfd23858448981bd330c28cf9a84f710555f3cdceac8d7a0b4e737
zeb2a6ac470ef11542d18396f9611a72c97771801e04c06ca83b0cb2a3da4a378bc45b6c6950731
z731adf43fdf5acd82a4aeed01432174b47e0370992771b5666272f4a8a28908cfe13e56b0132c7
z661441361ac9f8c3d9e18a48777ba391930cab6449c0e8d9472011eddb6593e0b16924f7db549f
z7ed31b547e1fb7542a824fb1ff80fbe9b6cc75960a6c4362719d7e3ac9b330003728c0f529d0d6
zc681223443927ecc0b94bd154a8cd31efa4172daf6316e0f3c5f85eeef2817ecf376d533fc48c1
za0953a144bc5fbb3835ab823241041cdec94fde539e05fdafe8ab33f961bc63ba963cdb66a2e81
z50b81718d7e49549ef48f4fe75f74852c941d3606730447760dfbc916c2773e3917f8ae60243fa
z3635b0cf87981f097714b21924885bacd79ea09aa854182b3e98e84648b4d8d33d417c7ee47724
z3296346c0a28f0a2a9e1d57da1a792bd7bbd52c6bdf5cde63d192ce6115020ed992736a5bafec5
z85af9173089014cce6ad6b0825ba1663759a30096a8a36455290eda434654632f9a4762820478e
z46a2f04e1f5122d9dc5a8733f42584e30954d24af858750884546cf514c8bc3bbd78d0d448af87
zac4d8dbeacb23f864fabe629ccf304c1cb6cd1d618ce4deb97d3edf4afbfaf051b114b478f7bbb
z52578885de5b5e9e022ec0ab162a474e3222005819fcd6db75c1938a0914e23731d279482e6d05
zda4ab75901bd0cfdcf5a71d6f295838a977c9b3c7254ac02526c41ff886fa93bf371856b2c8748
z83c32876608df133572c1d60d60d00b5aeb27be3ccb327993a0bc6b0d522e2e90789ffea028917
zf9cf1fe18e0a997b169de229957dd1767df172e370f0203ac9126218a4dee5df0ea1046a045fcf
z72e8a059d40119be988441d06a9cebfd3b1bab795af468cfafd2f67c22c6277b96f3b63503781b
zf0579c79d18f4530e96d03bf631827de6fccc6ec3eda4b813c17df5f991485adaf1f5b10f19151
z4818e918d596de8b4786fb72d1872afcdbaa79938e090b8fb0c999a46e9d55845473620bb97e81
z0627fa72badc1ecf07c428a1a37e19ee4ee7e21c5d272d7716f71f931f25b3a4b8003b118a8a83
z8aa9df59bc6f17b13e62dc7c3f54a2246d54985abd1bd587d5871ab50abc7ebdf434e784e3edbb
z42b495a30d71b88e5a45c330f5813d3096a5146b5f06148506c8d26a4b204cae6b16d4f9369201
z419c40d29d30be4129c49ac7dbb05fdde524cafda955b6f1610be0f0c61d50c01e9dc427db5947
z4b4884daf6be358934ef678ab516f84a0e256a5cf3fcee502edcb32daad244baf7efdd59891a92
ze7ad9fa7cb0be5f08f3fbccaf6ad0a3e4fd4766440327c8d678a9a18bd38139f2f8c55681398ce
z4012ec4525c46bf6b52b4b2449dacaa9527a80a379a9af47c11147b52a8b5487d4414ee5490dc3
zdcdeb8654b57487418d078db2c37e42b94d26e561b92d0bb6f1c3e9b8da0f2cc5050265368bed0
zcdc17f674990690c82acfdfc0cdaacab27a09ad38f0e13122cb1d0f7143a547f96e5c55510e40e
zd7b07220cc5aab317a952ad506f29d8e4745d79c675a57a5b99fa688bfad83766bfef5ca05460d
z75f8045988d7940f56d0562e8f8aef80095f4579d99bdb31e419c39c64b098e4a69912f65ca618
z8061780833949b72b08431318784ebc201932a71e7ea38b0837fede3c4727f5d1a50fc6254fff3
z31ba0896b769ce5929fd975cb87dde05db9cffd32933e613012a3cff7a87f4d78884950a537725
ze96443a5fc9bec3323078823598b545e314fe5ce08819e9e25d713077050ce4285546274a6dbd4
zab7494ad2aa4c83f703be714a4a7663307f47e33f72de315fc33f1bf24c28bc427e9e19e9f5189
z600aaa963a97b291f02eca4a6fb8cd65c9b56606ee6112d6e0afc7aafb541c0334384c6b593c66
zbb41bf99f1ee2f11c4c7f7d3dfe5d9be42664d2a2d4d73ecbebab94de7cecb8a987d2d391f9303
ze7bdd281fb30e524435d81fc55d986967e5c919e55c06fbf966a9e84f4853c535eb9b0cc402537
z4b45aa71c403aec894f4e36caa766b34920618e9217f5a8c41d16325ca2d37e27e304518a1bcc9
z1ec1116c4695b2a7692a1dddda62b1ceb1278f860c0365c888fd0d26a67ef367935a9f48a28cd3
zdaf8b20d63c0d51770cb0b75f3c0f7a98976c15d65f112e4a71f17242988c9a0e89baf5494dddc
zccea5e9a044703974ccddce4724467472d29a61e094e4635c170fa0525f27b995c7d8ba32bf2dd
zcaa9b566abaaf66eb814ceee4731e055de3194912bfb8f26b93d64f0e0687f65235c2c28b06806
z323394062c2f187a3fa89eaeee222e848ad253ae41c9c6828042a438f6fe70b47a83b7fa0e9344
z61f59b9dd5c1390e8169233e45bed4c295a6059feb7e72fe851f26e23716280ba8266cd1962b48
z92d892b60c0aa4160528a0313b687cba32847917f9cb6695cc5fde4a22940bad2b3bcfe2b8911d
zd0c772a3d0b9ac7640424feb1715b5fcd4b34652fe1914bc57628cbdaf6037af701db16c06d37d
zc7cb7771aaca40ceab504284e2d4594a522793fb0fb5706b9cce84e6e8ba15f07b4dd431341274
z70235e9f049645ea54d4def63b4343969897c4d7c4f8eb445356318b71e3fcb149fb6f3f84dc97
z3496943edcebb42902a7ec9e567b341bde24b87612858066381da652f58786d967d85c40663305
zf2edbf095b71db4174b7af7508202056accc94e0aab4e085d68a91b6916f05e85df7e396af4d85
z9e1b6297e47be8091770c427c466268f21ee286a96f96e10c8514dc36e6f45560dfb10e7737880
z520c15ef6d75daf55c9fae99c47ab16b5ce9aa74615420203429904c8c6615f863f272fce3d2e2
zb993070c18c6006efd7fa617e3031241c6a1c184208e47eaa0921f4da6fe3659865864129f412a
z869f35853c76d30dd48ec9291a8404bcb33821b714ddf6e0846193d5e3a28c95eea293fe851669
ze4429cbf1b01543a462965dc8969e578843d7c37375ea8dee40dc6720c2335bfedab46c8d7470f
zd1e337150dc4bb45a7dc904aa992655f79e3ea8a8b980540646b3f3fda6025966ec53bd82893a5
z0f49db94ab1cc0731d5d741b4eca4d32ee452a070e0ea743117dd124b667d9aacb11218a8584e4
zbd6785d85adbf8d63c061d720778481ac1a0453584889207d71e558196b340402e1db8d5743953
ze2350f82b84dfcfd268d68ce82a24b639fc8783913b9ca6d2aefcc0dab76de8bf42972c3f6720b
zd49c282d11e0e9384cb15f23dc2ad16a3f26d82aa19f441fbcd2008e4841b9eea175a67ea88bed
za329abd82baa2b553f1bc69d366581bda83280cf42bc89e4045a5f1d8ba4f9e2806dc33e86fa80
z099164067902d3762e239018b648b3253b4d497daa3cc48b863a2ccffc04c85fd67cf7fce86538
z03d09f4d2049c15517ef9bd6e5f5628c5ec433a9d8d5536b6654093f536b882c6011d750b5f6b7
ze4b61d0369c2f52961e650738e7dd00c2e4a32daa439ee12f8f961396875975f8bf1b7b3db3add
z3192e6c5eabe3c3f95a03cd01d0ae695c391cd01ee501acd4216305bab5a9e7d98ab1150b42927
z698ac1c7bc46a2a43f6f81bed70f326d0812dcb6c26a74f88d8d7566f401c6213e9c76a3416c02
zde3537b93f2d9e8d1680c83f4df82db78265507e32333b092ad6e350240b34f99dfe6805b0e010
zb32082c808e7b3e413b1ba8ffde3c4ba1479fae2200e435fa5f4448edda23bc40a046d150eceb8
z5718b36fe81a3c7a2108958f6723ac04fdb9ee20b76d0efd7056251b46ac19016e9a48cc975ce5
z3e5e8abc4670b2674f8a412b1a941e49b79bd720233ad59d8116b404767833193b87e61f1285e3
z095b94f0d9c3d536fed886d437255b211d8e0d8cdd555384deaa88134c49e7994c73da80024b17
zd9ce76fa4da435fca845af44c71a24dffed4f979ca49ddf5fba873cfe58971c7aabafb7071d4e0
z68868ee06bd061786d528ae1619ce4b26ac38c0b2cee5fd3db73b017211a3cc9482678fa3e4cc5
za9fb75d6a2526880b2289e2e8ee78c1dfbe3111832b0cd055e878c7141966969b64e876cf236e4
z15cc79a1549806f3a45397d7428d84d212ab5d86a94969ae0f6dec46fcc991faa15d241ec7a822
z3c0d64d1ad890b2bf34919522e1bcbf4dd70b37eba86d83c51321128aa0ac69b7bf5db73a8d9b0
ze2a1d3d19b1a7a01729abb3c5349f17d9086327c8fb8f3cb4f5574334c416c230b7acc089e0451
zb6ed8f548a182e191f21bdf86eca2a21d30a0264a78eff1e464336a604bf69011d37640b778ee9
z5b076375bdbd92b1661e52916779070976add5947e7e1564555ff1dd21204cb9284d7c77814272
zf22c914cd86d501d0ec9ba4dcf2e9051560326aba8f4d1e39e4b6c2c5cff8463f4dc5bfc154458
zb46c5ff14d43cea25840d76d81122e0a2810de37d78501f09039fdadf295821ac58935c4e3be1a
za4f75ea87c15ebb3c8b24739cffe3e06124a7672edefb49a4a0eba0fee037193f04c7e99524f02
z1983332c030b1f06b44269347b1e089803c40b91ced4cb36f67313422dfeeea3bd38ac82b641bb
zb70caa51d582aa3d2b7789d3b38e4646ee3616235ff286de382adc258f5fa6b09c39052ab8f79a
z2a3a3a81370fa4f1ece19cd64404ea3dc3d2d0633e095e3d15ae8af97b927e753b8604d75ead52
z925a8beb238ffbafb3c994591b6a4239dfdf44410f67475cc224edc6cf2f41e1452fa29cf02ec1
zb53f33428afbb6bc5cc3092b6b0c0e962585d12c8b05e94a7d545a7c76f3de3179dfe16c1c0ecf
z9c0f18267976e86f14eaaf61afb3f3f42fddad1a9c41f09ca9e692965f71b71beeccaf6da3e60f
z230503761fa62c3e1e319da4d573c70dab47e3d441082a9041b9ef84a496f37b7d5bc183606afb
z13f7fa079d9aa2e5de1490b173edb4fbd8422997e62c7d682a489b8d1784f3d9afcab8160e4993
zb2e74d51f863acb8c2faf9ab3b6b518048735e120ef9e2adfd173e7efb7120546300b43061d89c
zb38034dfb9edad4be9cb54fe3349225d58984e416f908c0dd5d3220e4d54de903a8fa70f0c1573
zc5ab601e46d663af8766c403e17fbe744913b576c5d878e2e8d969bd573280bc472e0eba1f38bd
zfbddb8b2860df7e102817d99823217907f63eb6981d032bf7f6ac97f6a2a40d4cad2271dc15a02
z4a31b4ff304f1553c8f97718dff3795cfbeed5afde151b81441331ad22016bbe1edf862d33c419
zfc5f8b6f5a9cb703d6f61fd9cfdeeb40b2dacf5fd796b9ee4d8416135c8575836721e058b381fb
zc2cbe0cab5c6cfde09772f2856046b7c0b92029cf071f862089bb438678fcf088c0c05f9962726
zc65677c07185278f2c044822944d751a9101023760fc89857df0bb5dff034de0a79fc5d3148a30
zef4c446e494c325f57bd2bd8b95278cd890c837e63ca94260ba9a7fc9c891eb6223e33a5dc96b7
zef31651acc803d2b79e5e52c88032ee22fb5b7481c59ccd07f2b0f5c93c6c9b209d552c20e30e0
z32dd9de8df9a65b50a957cf707d64296a82efb445c2053c1b1da450d1df670f649e1f60721c2d9
za33b1ff971e233c9da626579f872ab81adb9fe389a4ae569343662fdb1d553d4d6b412a4598784
z10b3e8b1110bf2273aa31ec20d07daf29f9f32b608ac3d0b5cefc8132af0c7aa73da86f7a5e2b8
z57c04b37da4ad8c7b304e9e92eb7ec09fbe1fc1067110237d364c0deb05de6a269b52b865f0225
z7437367900e2d1e5e8ce34e7e34487473b2e6a16d47318721a84b320888dfb45ded6764b762508
zf4fcd2b15889b26d02b45e2d6d457bc7e1c2e5d1bfa3da68e1a8b4aac80eb701673d479eecc208
z6aac989c8aebeb66c3d6ac2627f1258d3281fb94e6a56eda41126c696cba7a5a9c16ddb270da73
z62bd850e732fd917d7bd7943b3ef57d2ed445ff1ffc0d2fdfcb97af699778c68cb67c422431ac2
z6539cd9d87d309fa967f29c9f06fb63b281e7c5fc89dd4e90be9e7b8819f02a8a2af641b2d775e
zcdc8c84c40c81d0c9231d1487efd9600cdc6d56fab1078558cf13d2679e263fb17579079dbfe20
zfb6cc502029f0fbca77315a9e2238f25cf3449506ddb7769ab308514d1da11291594d658879d83
z86a42c7cab3a05f7407662d0e26e1eef8e6716b871567fdc514ffabe85fbf91246d34e7f349bdb
z13cab30a6f1f04cd7104b430233ac7324e9fcca3b6bd68dbdafeda4fcb2e98441fb63bf96b4c57
z089612036a845e1d87d91215052e8f76fca7217a334aed18919e3fb620abd60b7ff965563286c5
zb1d39b308ef5cb69f2c99a06c645445497de53f9a48f09126c068525b321e9c4f809d8451afb9c
z74fbef595ce853b7db15e20d5db05109cf41491dbf5f0065855722cdfa4e0cd3350ef61ce8bb52
z2fbb5e8af9c59f18adad25bc2fddff4551cd4e42955e3e18bf6ddc141739e6c2453f210f4162bc
z0ad09416eb6584aa8cb3756c53dd955cbeed802b4cf1a564a2a942a3ae93beee6c7ccb6b420435
zbe59afa12a87dd5a9ebfff9aacb9dd846438df5dd4b0be655c5f429551844e1dd00fb1a79b187d
z41065261bec75125f24acb0ba221a43f252a01adc983353fa4a4ab57b7093571cf629896827251
z821767d974039c6d1761d701afbe60961692d2de199c45e76469c58eef2918fceedcad9de97ec1
z8c4c98b35e1211b6ed6ff8e0e3d80eafa9516641c109c6ddde6c1375f7a4f51632ebf61fbb5c53
z74842442fb25fcbe28f8f42e9721a1977b3fad27c88cc5e0674a7905ab10024278e3c07ca9c33f
z4ca2a7b71dcee01f62811fcb2e3aed746aad604c311535d80a3f84a0a1ad9b6f2992cb23fa9fe0
z9edf166a1c1f159c54f8d3841511ebdc7a656b0efd324b1477bf8727ce8f3dab04c4b366ec9a18
zdf55ad2c0a6d2861d2ea69190ddd071b60f5002489ac3714b5159381fc037d066f54cdc54d6aba
z93e41d5f7237cd9c6383975e0356557083727e795bc8b28b06be23c3507f24264a13eb780a542b
z6540661b2f706df0704f83eca26e1b1096b9b96ff0b68300cb81581389e7d09434219cd4589ea5
z802f036ccc721a9c9d80c9b08ebbfa5f84fbe7fe12fa2be07784e88a3fc495b602fc16e6d047f8
z26101fa1dc49ff9154a9903eb056729b36b58d73b2f5a656cbd8b622e9964a73e2156ec399919d
zfde7b7ef52d8006f96c2dc68a890d62f8294a0f37d0f47ec06a716646e4bc23fff224bfef803bc
z8914ee531c03348c0b0b7fb849d390b206dbaa79fd7198f0dfd61980c11a20e6a51e8bb24478a2
z686781f165892576960b5f21c12489e3e7bc591424af9d6e497f6eded26f9de7870006a8592d1c
z978b3bb33331a936d576db3603d21da78dd6e7457a97542ae6267512a869c91fef9601912e57da
z521dd28026c00048c92b4ad89ff88b35f194d7f0cbb428fa0df69106ffefc7d2a117d2ccf671ca
z1634763101ef35badeca2a4ebfb5c01e44cc69e0171ac643b5eadf157b7766a5747003249369bb
z69a3ef2ad2b1e17ac10661abeb650770fec3927305299a34b6a524905c6a9785f5afe0a96ee981
z41e584a4d1898c5f02383026f1f78c11c36f1f79e867049a0c23ba7242df6f4fa304a738c66b40
zb5302c464e987ba96c3201cc3b23f36f327e1371bbbc1cb6e5ede9925074f3111106e6caf58716
z3124cbb41ee1ea6bbcb7b1c3b5aaaa4191e5901f13a1fb3fb49c9f79991789c97f783a606f9886
z8e969a6fe3d52cca0f4378c305f7d52d2e172831ccb283443943a37212006fbd3e824cd82727e3
zd8e216e9ddc5c2d42a5fbdc021b409a96e42a0c3d2a03fa62be24119c20563a3483dc5067e4ec2
z7b852a495859096259b024655d8cd271f3c80ca136f0ee4e85edab6473487ea17d80f77b5c6539
za3b9ae446da6cefe5597fa5f4f91a4ef1133add60afdedf3a0c7e6ffacae76f4f463f877c66c9e
zb48e4987d3bcf5bfa7e0f1f68f59ed08cb0f7df83873041c4b1574a4802cb30ba767268a2ddcb8
z0e29c853fa30779eb96dc663616fa80ce96655713484bfcb999c4f7cc66936631db708c8575ccb
zcc58dad1d1b7c92871cb66d1b22d7b4b3dab8167b6b8375645f47d4b146e2e92513086fe957d79
z80d2fa2fb7cbce138177cc32f39218e867fc30d3531f9badbcf78f88c8372344398e5f83b1697a
z3ae8d08ab69659529de059fd9efae4a115c951a12ea29dbadd3a99034c6450d497d46a99d0bc84
zb324378c84fe659e45fe63bc7c932321e416ff4a9096b0004c94694d182374dec2d20bb755374e
z0f9dafae5f99722a4fab1dfe2562af7a4134f4705fbaea0225b4704153d8cb49afa206d7f01584
z8e56eea8d79164ea5e38485e1cc77202b980e6f8c7a688614552fb853461ec25351c55f44023aa
ze2971c8ad76f52282a580ea8aa87ae8247fa98e6f4fc678ce112432a532d0086b4e99a9a287d16
z83e0464dd5e22a1c17de3bdad0669685957448e7670f847ddb3755a12c5452321727e6610b4dfd
z974d01fca44e6748f6b32eecc438a6f0775cc2a62178929cb735dc4d511212229535db46c06ed8
zd260ff572b44b414fa9a8c0022825490145217087ad3ed5add97690b256bb23d0a10cfe06d1ca7
z70599d13db13ccd487193b7dde2b5d3f17208a5147a0ca86daa4059c05e04423f1776939b95c2c
zcdc11b7c6e669cb5b977400f35776299f2836a4ddf378774adae10d96f168c80163ea8124fab6e
zf388230bf69e7c23eb2733df52848a02db7b1140b06eb67529fa83680a84e36c10e03709be2bf0
zda5235dc22af830c27f6520bff2af9e6d93934546de700c66e841e7e65daf87dce03031339df2c
z41e86534c446ce52ef5471f9f88872dc2ffda5b64b3aac115b1f3d264ea03da7356744b80bc226
zd75a27483e86d43e7e03ddd887d30ea5cd72de1cb147abe0bd64d2797b3d59f0933bc66ff4c9ed
z56732ed68d2c89b34873ab9348e664d673b8f986c3f82e6504f5d110dbb32cf43a3443e8f168df
zeafbe116ef10464062b3898fcdb715398c5a3de7785f9d73febc514cdd13290555628816211a04
z5ba3affb5601ccfa7b9d38eb43e4bec73ee4d5b7c30ae0d3f548281749b4be36e20402dbb7a456
zdcd3898ab455b076b0dceb4688ba332fb79f36c82d1748284e95122c4cfc89665f641183dd3772
zc1650a807f52fc9c5700cefee4bf9114ce4e826365a31d874e61b6ce05ecbc7abdfac72a8a7baa
z3fa0ec1ab26a9395342bef9c1e300a7a2f221fca3a702558305c427f81b718eb2eb3e5365340c7
z3708c49d06fba77951cace36ca7d18a0b782f944a5ff6c1d40a4ca8b8b6b860edf36be18dead84
zaf94bdfeb6eec5b59be9a93a643c9e9c42093886d4e603f3c0ad3d5ea0911e2fba9742f9e071cc
z29e59aa39d74f13581f0cf09864a183cae30c393c28103be246cea57c3cec730410688af6faf89
zc79e91e8ac4c9f029cee0c2059b935233406e00fc6fb5b7afed9958697ef4827ab17e0f0bf2cde
zd8591883e0cb30936e4a1871f1b791c3f969a8b6fe1a72d3358541c0cd68586714f0cffb8bcd95
z69be57bad0cdf9bfbaf79c6dbd2fc2be99609907a41864708b575a00051ea2325057aa279b744b
z7868d797601d09bbe2f3fea398fc13d5125e9c708fe85364903ff26889b50787abcad2e052e12f
zd837789746e6d2d3f310f507d627721a0ac46deb1c9ed5773443e52f0b12ba3c8b8358630e2393
zb4ea8cd21d95bb94b6a9df3dbb6a4d8651dd1b784995f915f0fcefcc8cf109757de27ed16bcc89
z31476e6f66dfe45224283aa9050e126fb279689f2e0e851daa5c2e7d7d96a60c48b01f66cc6a3a
zf1a9a092baccc51378a4d11b93389597f8e76b6278a746c8d31bcb9297e41cf5f0382af6080bc6
z6e7b2e0757b6374020ffcf5dcb1d20d81ee38e8f118b32f20d5c46bdb4dcc59ed61a6a9460504b
ze217ceef40e4140847f884b28e04ff31499969f97a1f77145d267565f232012cdd779eb31ebe2f
zaf3aa07c8a69e373824dfdb3cac43a5c23c7257c10840fd9c51be9117e9451f65648023d246e92
z0b84d9568625bf6b15b0708c58d65b88198bcaef0ae773faf451952e6a818775811674fa134c69
zc603435fd92c8a0ba31386564d28d5b425e5aec8778bcf8370dc3639abbc045ca6aace030b57bd
z957940cf1cf1ce3eaf86593bc67a30005ce6d788fa04b2c625c8ed8545805697248b5aee0e4e9f
z57685791dfae3c266baedbb0bbf825e4d4280ce09ab55d84c8a7fdb43c6912e928e0bf870e654f
z36b0d0403d565bdc2c7d85e23137da4ad5a3639aaaeb302eb1a1181e6fcd4135b0dd3b05872af7
zd0d3280e46f92c5024bfdf497ea9d6ec6e3a755785cec57e42d0785a753b54fa83746818b95b0d
z781bbbcd6cb247a15768865415bd3a6d4f39a6f8e690ca3e6733259a9d5bf177be25274f044ecf
z36238c48cc5e34cb85e03838556e7087b7e518aacb8fa3418c5de7c0ec26274a9f881dce72a03c
z1fb18776eda1e87350300ab47fb722040acd0344c903872419c1a7a7c3701a7222db8176a14d92
z719fcff31fa10b25f6243041c1e5a4b69aa5ff97456291abb50e8b30ca81bde79990823b10670d
z90e1c6e44dbe2cda3a4670dfc1fe9e0706ae6747c89dc7a530d5817ec089b72131e334680d38ae
zd85cbaecbe00f44545fd3426c9a899d464f4dd9ac4e74b3122ba1cecd9dafcce5fcdaac7b6203e
zc54c03a33944c0ff8db448b23c60f27efe05e89f56a02b8ff7ca5e5451e8716d8f65ed99d7f79c
zbc318d80fa6f7d58a7abcd02e75ff352cff5781c689afa2d881d32649a40b489f168c307ea81c8
zc531d067f529a993ffa3ab71f804e47cf9b9937966b8ef6d904bf3359cd15e9a6c0af5d632eea5
zf7a424e57cab4a7cef52276ca084dd4bad3546b9b26afcb6d137f26755d9d5efbc2cabf70d7210
z8aabaa991bde896accffc3c24584429979db84dfbd39376406b1c831eb803c22d7f96baf65f98b
zba38b2a81cd91b47930da7bbb11c8caa5a606a7b0a2467ac3d05b03605f6d722766462d65311e7
zf1a98330cf897daeca294d275f753306ad725a8879f4dd6109ad1b0f2d0a425f6b06395fc2da5c
zadb3b3055d9014097fa17c2a104b68da119b50f554a32b4d6d51f2fb43fe55f83bf969681db771
zbfebf9bf7437313c1c8db87641fec601db6a3f644fbe52c8e00ab620a763b5bfb7fd1557311e5e
z8c53b252d5302835950b7d4d059de6c32461b742217f6c24e83754da703bc35ae8d2a7f94bac9e
za1ef535aaa8e06923f4d5d9a5439a727ab5b62b8fdbd1353d67ed5c0f245bdf36b474282084a05
zb7c0a934b9304f8d11d61c25eb078b36882bb24aed79b6e710d75b3a27c89085c9619c772c1fd2
zb378171e993a4c9f4ca72dd03cf97b853e36cd2ab111597551830001076917544ad2d9f021f2bc
z30bd28eda89d4b1893cc027e74ab58521d215cf0da52234721a46ec1f442252f062a7f2ad3cdb1
z05b96562a47a849935d2f9e6937de24d85eda1b3dce4ebc6fd0834576b0d11f5145403b36386db
z1d56f4ee335277ed93d153524316d197b383ca7609f4cb02b5650ea1722649c2d955565552d8c5
z50c434ec78ff0c1333a2c18b6f303736924b6fa0d3cb4a11abfa43a58c823b5a33a28762ba72b3
ze704401f4e7efce0145cc38d929addc866ab3648fad5b3b32eba152fbb57e06c0d4dd3c47ae22b
za642843bd5e79cc97c53fccf339b894265ef3dde33cf6e2de0837d8206d676c19f5d9c64921d16
z6935b5628b411c2be27e82d9bd0b1ba392580a6160fb5d5cc19432ce239c14a8338608ab309011
z6d3693f3e2d1ae0a89a349802202f745cfdf0196d71a8a455601caa98133cf41e9a203363585b5
z91a3894578b7c6f0716bbdc37ee8e362beb60a2b55350cb260212112891f0159ef29785bc5cefc
z07770d0f8e2d9709f9634d34e22cb65856a6d6e6c56f96405f5bbbcc030c202bc55a227bb7971e
z8223f46e6adad5903146df528fe91f6086fc1090a93ada3d7054ac16577e4a99b3858faa2d1066
z4bc689c3ffa2cc12ec0d0a8151b288699a91daa6a63a5f2969165a35368f3b43ef0d8f302130b4
z9f2a2371bfbd6b46687dc81f59b5ac1f3e75cd11446bb602dee2648f6253fe44de3aa0ef355af9
z7d11cd2174df2a7103fe6d823cbda7dc923fcaeb13e7b7f928073d71cef1d4759b8d92b1b0d9a3
z21f10ca5e3ca781e131d711600535da5f3d10a3c6b913a4bb9f0b5536c20b9705d24b5092a2f71
z231c3dc26d7ee2bfd38d9b869585a3d3b2753abe965af2031a805a582884216dc0b2587f922d86
z3ba6e77d322d32ccf4ab3658f8a9207c5ac3fb5e037e24699f9a52e2b5821ccac6ef33b4189c16
z4f9b3fef1c86fa68c83cd634cff75a4b8f794edb71a10638bcdb2e8bd37ab09df6fe9da470de79
z67a5d7d56a720e1f3e0e25014230b4ca5ba7b7e9e133078f6553e553d8f06d8868aeb3530da758
zdf6375f37e3117a517e6cc0d4460174333c94ed3dc26572f8667fee78bc496d8fd18684867c3c0
zba8418be2150a864fd1b8149c1a2e0469d6aac437ffd0f05d9bbcb4cb93311cf4e73f7bda9b6d6
zbda4736e71dd8a4f2f67472dc2069c28f70f7ad360dc08fa68ad271124e3146757c2fb147b24e8
z1b2bf38cb2aadd739b826016bfdd2473a89c6555d1ed72530ee5bbcc5e0e5c58eee481852a9d3c
z8b3647d9a2a0b2759ec2e9f7580432a6643d1a98ad15d31d0dcbc1d4fc3b2c7ab550fb2f1d22a9
z9c8d33af2347684d773b80b304fcdaa83e71b7eba98ff1062c733c5a041c6b08aafbdee028084d
z4ee7d3645f5c96b595917b55072f8c3c5857da0bede0849c4e3787a896d0a1b6e6a2471012f9ee
z1472c584c6eb2f888a2ec2953d0a7bc636484c2255113ec27f369ff63b87c73526ed9059ca3ffb
zf7bbebe9e1f771d9949c26099227fd9f4795ccf5785239efe7aa6f6961f7301021858fde35bfd3
z60cd1451af5270b029893f86f46e42d6a930a23f0f01b99b8d2b8083796b5c82894472e86e1a0e
zb5ebe627978da7f3bf3caeca2063ee7ab80c975291506c1ac097e6f45b81604193d2fb23e5e7d1
z7e03cb7c76b82583b60b231f503fe912d7b698a0808b58077caae64c4d52ae6a5338dbae961f65
z584b7143a4591c0e5d9b5839ab2fa24cf88ba1bdcb301f7d2a99aaa52c2af2fb38e6b55f74889a
zeade3278d19bec2bbb56a30f0bc4b48bd31cd62ce84a18c25d9380dcca62da93ee3b53cf16ea3e
zc6b978642b85def8cedbd9890d51c7973a477e8c17b719caf958e691c69232250b45fac0aec435
z0b24402bafe3a2998f52b1e0e89d21ca0f12143b44d41e62f12679b7d0a6db0420083695bec747
z1833a3dabb86c5939d251c97330372c307c3683ca3c2d15c36e09b6aaa2dab200893d84e2edee1
zd87f27d648e54867dab1a97757f45688563d85a3a2bb0cee4aceeca17682aba64f83ea602018ea
zcfd168811213b88595070bb10a16feaac755516c470ef6803a6966ef59f764234c14842378ef59
z2fce55466fb4abf60792eb870d0b1820e13be7c4b4cceb7e2aaa64dcd7def349f73780a12ab23e
za4434a969971033355b1db4eca7c2130eb76c205cfdd1d0cc4dc200c83f0bb98fa4307d7135d5d
z691f1c7f876286810b7fe8b9900779519375ecd924fe57c27accd8e7ff3860a29e9e6a8ae12d73
zc84077bfdcfc42a03562f70533c63202b5e3bf9c7f741dda16c49ed0a0f40a0513bac1a86650be
z8ce743ec3a9b56a43349f131df7df2d6e6fbc0841ca6ac8d0dc295fce614892cab92f5be33e19f
z3a6152f8a3220241f301b007703ae3015c4b466d275b094cd5507b89bc5028576ea56d511e51c3
z14e5ffae4febb6dac2253568455dc965059abe73d246e5a253c61d3081f268f5d9594921da1ab5
zc9eb9f8fd1db7d0aab36dcc56d9378a41f80e124bf697ce7ca237df82216be4d7b604ab31f454d
z08840f02c7ce966608648ee5497bca19d16449b432feafde7457c8e56afa15bccb3ebc284f9bd4
z8a762a15bead47d7083c328014f060fead1376a52546c6a9b7ac00ec635d2238476d841fa32df5
zbb7f86b5919524ac7eed69a63d5712821ed0d4c708809ef1707fb29f51f070ec1249174b9a6676
z038d17b04599ec33e2409d3069b87d08f146b021c2fcc0185234937d1794931e04c2ce1ec27bac
z8e08231a083285db0a1b85794070e576f0793da85100c4fe9bebc4572b36ef3be8effa8152e748
ze7c0205e78fb82d9ba91a5217580a8256fa2f69293bde24c43262b6d34eea6703bdc75f8fff39f
z32fa75ba0e1a331e577c8c75b3c078c1e5dca344398c57651fdbff94c73a664e5885df34a0564c
z7950b0dde5010272bfe8ed61de817697d8cba40d73b874a8b99829a3264106cafce07ebc6c15f1
zd60224450fafd6c8312ec692109d0e8fe42806bf3e196a3078960bbc95d8293bc70b1fc76796c5
z24b3ae27901456204ce0bd5cf615ebd0599f75f9fab593b3c587ad1c0432b67932b5b5725801a9
z4c09106d5aa17ab7c073b9df777e38c8581a91e31916e51a9fd1c765f4bafcdda64e585ac3175c
ze652588551b6f9c394e90cd140ed151911df5799c0c6af412387356f471fd537bcd5e309d45525
z730760db057a05b6f6ec0244b635f21bb82c93007040effa628a5e8eed3754469f590db7f9ecf9
z282dc76b3aad732299b6098e2693cd15221639d61fb7b74e0e98a650303e94808af6a92e37b1e0
zc2bf78abc6f905854da6e8d4e4198708a36bbf6776ecc523a48dd8ba40c3c8204eac78c2d51200
zaddf72ac00d9912b61ada634f394580bf9cd8ab7207122614868f65932a0fc0f96f0773203e50c
z29af95a96e5f840a66ea51cfe46f2e2a50f285093033154260a9dc20061db6122a90f9fe5f521e
z4047f5d5a00485e91434cc38d159b98a338f8aaef7c9e1f6fe843578920eed85434d4c6b4d2fdf
z1c7893a983850a69a66413de35ee46e9c68a8ecf0f85b146a68acac17f82febfb04aa9587502d1
zd3ef39b572f769de31df22c3c4164f6d81801e2c5e9c1e9c7cc68830c28a044a5d87a8128851dc
z6cb1729aaf2cc3de69bc0833466316c2a5c80a1e66ab2f00946fdb6f236b4c7d79196c3e564d7a
z28964130e35c64a17a93cc746e44f9996857ee037913d55a99d74991c702328e3d2acbe946b9e0
z11150de5aa82a0158b14a942d90e4618fea7689a2e1c0465cca73957a0a5085dc52258cdddb293
z95f11532ecf625dedd5e4b16210373c781ba7745f732141683fe5882bf07859d7d5a01b755c2ec
z6c709900be44c26469d838cd8fd7efef719929a4f75216bf1d664db94098c9d8d99e22fd93a0e9
z0c797638d4c346cb5c7338e92d392b13098fb0c3eb64b00a4bf7bedb5eed59acc9f8199021a120
z00129437ed14b651a25256abb438f6f74f2ee407b16d581913df366ce220031c27b22e36f0599e
z33a03bee6b76d8f3e6de78c9f8ce8ef60dd290ead1769e163ec495b781d0c0f511c0d63e099ea2
z8d3035dd2ebcfaf0acc5a247595327ba279e552d29d4d75a4550942681c99d3516540dff0f8159
z6e4410ee7d6b2db0ca6f3343b2967acd4ab0d5a88a77f67f96f7a2acfc8ed0bb5682d7ac4af64a
zf5a3088fcdd1c9ebd6ef622bec10b1881e4adfa6fb3fb263b7b0beb02d809a74cc04496e3454a6
z00de46cd434a59f9994e357fd3029ac7057215cb16d27b5e055724cb166021ad619626d19dca6b
z609ee43aed17dc947213aa3c144d158b18e763181828c48eb495d0f264031a8be5c7ab39c138be
zb08b9380af8e6aad728b30f233eaaf2dca4737b48ed8a3538f2e946fa95fc848e262bcf1d27cdf
z1ecd4056b15bfef68e49317fc82ac4fe89c153a220d275827f5b6b2a6e52646f6c38ef2dd54fa5
z01e64d98979a3d6f1b96214601eaf8a0d7bf08503e71dd226218d6c5c1303f45e38fdfeaee0026
z3ad8e62b1579ad14366ed4f03d1521ed13dc11f767edee791fcf2001b0f3081f1e7821c8e18b97
zadcf6400a3bf0935d9b4827f241f6364357b0053ecc27bdf9614e65e76f8f8e312ffe1221e4b15
zbfdfc7dc60edcee14aa1b968b1f617f980fd97c21bea31ed03c77f369e0b656bdf935f2bd4d9db
z7a55ad04e517a93c799912af49a3f8cee34603e71ca012fcdec77c2cd6b9f3a50ae12aa1fd5815
za842fad194f7f99e0eafe45484d74dc8f5d36e73b434880110b97041ca43fcf1204db7552a4a4e
z941041c2332f2c69a68bee7dcc5becf6020c0dc2e45a9cc9f9ff4f02588f876c9f0e99cd0abe6b
z67bb5cdb26fa2a2e86379bed2cdfc5774fad3b7f132d12083954b54edfcbf0a85fa00d573405a3
z7da0c6d30a4352ccbd4592d7082748e9423819509645cecd18e2df55bb120c6f2b47f9bc5d214f
z643d73bac33b6b972a818f8ee36e145089a8d9993e5ee32fc8691cfeb2cfdd4424c4f094157f89
z10d6dbeabc27d03640352b1d6c372fecb24aa390ea9a4026fbd7aac5c9bc4b50d077f17e9c0b23
z6299aa079726a6e4a9ddaa50acd5b2dc2bc5c533c6c3dba5a5e64c992c20f18f9539a8009dd125
z332197ad892a14232165e26b7d74a89ed5dca0761cc58a3a694519cf14e263801bf12ac1345738
zd48359abfbe351fc93ec33cf3b033e449cb7f5a6ec1db8889e3dc0aab9fc1323ad0bc5ea4571de
zccb915c8875631478dc88c938357212159edc20e999496325d570ebaa762bf6b188c86c31881b1
z98130591697e9f74d08bf8ea5a279bfcfe251ff0a707d75c4da2335d3e2ef5dfd59afa8f342068
z75cec8c315f60bbaefe8f01155d8351ce32772a264538967db4acaaee8540fe568ec5c5a678419
z4cc0f3c0a88156d0f97cc68bf9608dd507645853bc8618ca8a56e3d559d8082e1976aa3dfdc533
z0d7d8fed260c8c4ac34c6c4714f9c3b1d5ab7ce99ae26b1c78dc37559b69635af2d16bc6ca39f8
zd561c572aaf45f7bfbc3bae8679dd5e24d6d3d2413a047e107d50222189ff2a3f67479b068ba96
z7bda9a03a39f2738ca10adad48ac3a08ab86cc8eccd3e5aec1a718c7fab45a32a6494bd024b2ba
zc3ccd3d74fc54613d78ece724d1daf6e9d60ead7924a43c136dbdd5862e668d77d483582d8c741
z56d9629a2f65172baa7e6282a0bf53ced3069351f5e23d5da9c57731edf048afa5d0acdfa1e901
zffbcba77c3c1b2589dec4aedde25e1c27a0df103ca6a3a52cd8671af1f8cf7510ed2bdea7baca7
zab6d4aa20f008a3749d831a6fe4f0339edd6638d0278441b913372b1cb8bd8965cc9fa7a705fcc
z0825ecdde1291960e9e8b19a1c28dfe5c2a1846b17cf38492104d2722caa0250f4cedfc135f0f8
z59b252a747061fd5716ed02d88d99152b2070a48b91e954dfb1fe70f0608cc21eb491044ec584d
z3482b0cb5c9e04b4ee396b42b5f6b4bb91c67391a5839f32f491d92f735cedbc0ade35cd132a79
z185b636f02583d679fca1e9b27627a237e0b60b2e573eb046844a78c77981ece8368a23ba6db22
z21d26b8b45d327ed4369e46d8cb4fcafb1f10dba488f3bf1daf75576f630e399099e47c1390b26
z72e76c0eba523cfc0b22a578035b490024099f6e5de6960c4024aec8143ae529fedaab2b94b640
zfb268cfe05b70f8fa8a09ac7b6e8a6b370b0cfe2797c4de0dc206b95a7f7629fa9f0e472de0ff4
zb5ad53b5821db31ddbed163c9ef120cfb0487f123002c5275027dfcacb117cb7944e86cb5481e6
z9ea2be6bb47ebdf5f0ded343806fbe5568535cb2e1e97531f97040fa6ee781221fc5469917db4d
zc651a8d85312015df57e5819c037ffa657d4f1d99057f2af96114cd25af7fc7c2be70b21ce57b3
zde4b3b9d82935ad85e92bbd58522146e6898f73b09c2d75b7ed6f12b045d785457195498a90ad8
zc61f3c593a39f456e6a466b3b098e1162a64160d13614fbaf0c7def7527657ce74341381c0e5e8
z27cf52fc27f8693fe58230c0b18e6a2b158fd600346a38ddc1e8556e58dfb05eb7b7fe73e005a4
z04cf0e1d79bbe5ce8805bce541c55499b9a1f99cadbba8f2e4d2914bdb61ac82e45ae089a28ea7
z9fc51754b7f19795bd00635d1ea339d14bf6c7e839f82c671cadbda4928045c9128b8e3ecc615a
z85ebeb5bf6e135dca86821acfea1ebd53491602fbf6c87a124373193bfa634b914d5cfdfec306b
z0c205a2d7920a48f30403c544f60c04c3965a7bc15e3227f628425b9a94782414beb089ab929a9
z58ac97e43cf6b4d5cdc2f4d12a1e5a881891108e519351ec4836468819a551be24fc55f5caf799
z079c125cb69df2589d89d1f2d170e943db9dd66344aa81cac2c944fb643410e33ad9a5a12938a6
zcf098f27600460b8a13b7bcf09d58cc18f10cfd5ca231a88f7566bd9da1c45cb2e5c5fad610225
z4cc87087f7092b639937be7c49402b138cee7b40339bbe7a97385e3fb7f134209406282a592877
za96672ca0588407be71be860fd508e1588336ff079a51804e0c0c7d3ebce7f0a27bda553ace168
z02a64cf63ca57f509423570e6bc23233afa6b3e9fd54016b8abc3f94bb2adf9c572c00f84b8298
z19d6c8915c30b11e0f6e27b6403051054def6b62bd36ccf44ccc5dd42a5b1ab271e426eeb3422d
z27cb5cfe88315c22acbc7dfe2f13813a2aea1ee695eb2a812857320f4f47c3f9be9b4bb51105c8
z9cd6c78e0266c3bc347c080d1842ecd7819618887de9e111bd5a53ec6db374a2ba96d464f93282
z8796a8747bd781ff57e8bbe54e0be131509d3213467977b1a1ae56a322b5e998d857636a63aa7c
zd505f5e7c5ab8504977dcaf2aaa1176af9bd82c90605fff8d2fba8f482f8870908dd8ec62dfb00
z347b95b9588990df4176592396c81b774795904c350070c0c9184e8bf46f074055c29627c0393b
zcd3c745d3603f7292bc4bee74d71ddac54aead7e8239db89eef5f2f518a53d0f4e8d2c0fb27892
z9955d8dbb8d09c0af9d6f0ceed03738202c90975077f1f9252da1ca76dcf29c66edd90d6e2c513
z6b8ed4d0b08233cfda96140b6ee5a107477f2488620a62b0d791e2e5eae7b4ad9f1276a8140ddc
za24c58168bac6fc0714a0a93645726ac64140a866e25d71c996b0704c5ebf869e9300420df985b
zf730f2e656bb8b8d400d118eff93216d5bd8967d10c3b1cd0e602f72c101ea97117c4532c05ace
z19ef5b454ae69dbed67db68e0ff1a43a949385dbd52cbc581a9d403a3cbf538fb6a749a99c5695
z2558c3430a72021c554bdf330733a54c41b4aaa394d052bde4381b28185347f8a8fe7f2e48f845
z77ccddbbe34d083b919ac190094a2d755571aac3396506c865b1a3f2bcad55b9a036a4faade3f0
zf78669ea3c3a124664180ca706b98f8437496ff504d6cea8c13f67c5ef8a2d8947f9c273b06e8e
z251b1842d7afabb89b6d688adf2e0500ed101539ce999792baa469c87fea3eefd548469c71df6c
z7ef1d95d6aa68a76f1ebf7159ceee0d7cf9570c1cc8706de40d91861de6d98491bb3cd94ba6745
zfef248346a057f2f72423561d54496ebe5878c01abcc34c29ecd0ae50a011268fec9b5c8886e10
ze3440e4ecf3a5ac5e8b6020bf2d61b913f6745c5f28e3be3ce4d084c45678c64a1912ff2f88a37
z08afc7218629904bed7a9f6198c2a8d1fa275a4861c949d71dc9fd612bdd6f82638e22833599a8
zd5eb50a1f3df0ce4f2374d907a24ab310feddb69474c758cdfa97b4db1fe619afaa80fd74a7541
z9cad08fd20ac74c4134079466192b75036a39c64e58d5f46e3ee48e3e700aafd7508ab705c9447
ze8f60e978a9ea47a81fbe9f0a5e378049052e70ef777cfe9eccbf4d68b6a3d997ff7cc7a5ed3c0
z59752ab914093f04c2fb778ac720733e82e142c9d243ba7ad2c2531fb4b920b418643e2bdd388a
z11b87797680824e2cd5b70eae1bece797015ecd1177e5f4e5b1ce69b9696cb22ac9511f3fc6039
z9a7f94bdabd6b9f004fce159c352851f5c54a06f7d6f5833a1b393304e1b18002ec46e98e4f5ee
z4497a4744a9900ce27cec8b7f4178f2e01104777b45ef67b6496ebcbc1f2c8c2ad4275d5b50483
z3b83ddc4134e242f1dec97a125e88a615349cab5bf9836528408ea153b2f4284da0abae7ba9545
z23396160e9fe1bfa53f6050468ca2480509934ae90317d114944e951b9ea375f8cd334f0c81e61
z20dce949450cff7f45c78bcc7f8fcb3e55f34a52ad7c86b57564aaa32a4d96de539dffd59e59ad
zf99250034e076b152bfc4fced8b2181cf79ca279e0274b4d1bb526a99fcb7bc115b48f37c36164
z624d42f3797ec1749e49edc38831c45caca8f87e79ef94316e5aaf013260de35348aa4d509adcc
za14ed145e68bfd91b7b0aac9f959ea0160e1477e0e01e1170d60161df159962c5f95b4bf4c4d02
zdb269e7195d6848fc443fa6a11a231807e844ae848d40fab870b8658988b0a4920972ea4e3b046
zf12c94285bc97407749bc155447d440f7d22f5d0e272d4224af53cdb970a3c0183b10af16c6482
za106d1440538948bb5511b54f6caff5eda052da309ae4628c490f6d6e46fb69a934973577ca735
z8041a4ac6d33bca4b91d678075753ba96b949deb07dddd60f757be5685efa7aaf1164ebac08611
zc9e50c32cdbabfe1229c1c77463d63d06aad75e5b918496438a8c23b25e40b4e03f35d466c03be
z3b4b7d5ef182b0910909251d3271d39ad05de79923a28780c67ab92ed12ce96360d3489e120a51
z155642d7ef27ddb432dcdc29ce5b3e1e53011c9bb0b6c2cff0e8b2c69632ebc929bae10ab345a7
z76a418859710ca1809661b071559979c10321c40619c1a00491e9dec7fcc1e3b350559ec40002c
z1cd836cf1510606714625833c7c1b7604c1d6ccf96bef5550f0c06f5c5ad3e6a6ec2797d14ec32
z1d8f3603d072921d6d6d0caa37c456db45dfc2c10608c43784dd6da58f16aacb1d6c3e16aedc36
z90865f79f272e1bb807eaf72ff154e12b416d116a1d29caa3b4ebcf2150b751cc673d0cf400f4e
z7844abe947a1bdf4af786d3e5bf62e073b69fbf20b576e8a40ddf5bff931d9b15e8a73c9a33fb7
zee3cfdc4a861dd128d42fc286debbcc9b560b9acd11366800a5291a3d85c57eb84da53b9fe7e90
z6e8fc28ff528da1ae3a6c847b705acc2a37b04547f483adc25c5f56cdca171a0d2c45db9696b62
z6b633fafc6295b33ea9023cf8a0ba4fe6d6798117b63bd86bf263a788535c959a0cf2f758ef1b1
zd1e26349bc2f00b31ad1571065389796ce0a14f14e6a38b0eae4d9ffbc884f96d945c31f980090
zddce386dcf9feb64cc5f09d5c7e945001721a4bc83fd441877c935cd9a8ba0987ae306232c9745
z0246ff4a9307de372d3c5cc316d2ee6d286225944356aeb9f0ef9126c8e1521c3325690d230007
z7871554e300fbecc28b86526aeb0b3a20abf2dab1ceb5ba83d9d03bfe8c04b565463549a68b503
z4e8fdd68e7bc723e41bb0e1f4de8021ea7c6bc6b98c08b5df072b3c05cf784e6d7716366f83db1
z626cfb0e5ffc108260bfabfd19faca53e4d91b8cbbab3e70ed02433f5e8643cc9b8123bad210d0
z2a24114ee751fd8fa5d877d175a8d019853c624dfad6c4f5ddd75ba87225420ce7a388912a0ded
z41bafb6ddd04598777a590cb8d36e29d6d21d70a62de34669fd9f43e767f91db63c866c251711e
za1515881291cafe7851a4697bcf6f108b2c5217623d8154e5e6a356e3554f0a36630a736f537c7
z6e9d68dd72e60d53a4a5d82bb82b00f371b4710c8f6d947e61bce23bf65e9047b66768d8f56362
z3b1007b325b8533f39c972c9062be51bd078b8293abf2c84d0d54bb552e4c6015bbb1ea1ef2dcc
zdf1ba329d8d30bd9dd118995b59b63d4631b1928ce55d185e7d9ed6a5208cc8d0409244f43926a
z49e91ddab58cd6949d0325e2a8fb5794064661970b34e1188087e0d35c275e0fbd38a3d7f7d6f6
z53536e26ec19a574a287dfbd8b16a94ff328ba6443984ce2b086b16e14f816b3db7053fbe13bf6
z041d166888728d78a8868a70358153ccfd078a90be74f948c7a3d68fc060d5568df2a598370047
zd912ba0d4c53702147c43c183ee940c94115d5c62aaf611f27ec0832d5960ef019267576cf257f
ze76f07a364204a5ab2b60c937dc936dceb509d5d6e0f8643cea83cb97769198708e99e4e41fd15
zf1cda14798a8024719cdbfb9acad7e1167dd8f4a7ac3beda2529478b6f616dd87773f1e4a8848a
zd4ba13214856a6393bd48bbb776f73d7362102efebbf73141d4b8c9cb7d9de2d4413c52b158cdf
zdc3d31f08584fb1b801fdab66e9e29e37c485c25a69d531926aeec7b04415a6754aea26d0c2e24
za59b09afc2b6461e3e914306c76e7af421582e9e42105fc576955370630be80e594380296dfcf8
zb87bd7be0176d9529fd9b85581938a47713cbb2672c55b635bbc0d0189b57a297854b9748b4ca3
zd9013785030781fad0a1490bc55a874affdae62c69483f62b869d640e29bb1173fb89de8fee884
z87e654e694492a0b8858be7432c10f98e96491ee94d15fa421bf91d91977ffe4eadf06130deb26
zae1712c6efcbff845c6ea6958d2de5cf1b4fa345e7f3cb2fec68062c182091add572f7ffb1efe2
z44f1bd27f493d7975d173fdd171f44e27aa1e214532d8dd99955c22f75248e920f6da6093b893e
z1680df4b7a83e34e2b4238f85af726c9b5d114424c0a6be8272f0526b74a6f889f0c0b639d55fb
zb15780efb4fd8710d3d437b18e60bd1842c93f60932452927492f7525282493ba7a636b8dfa29a
z74bef4263d6158e6b1f2719b6778c09c225a5fc38379dc45a541126dc93095492e70aaebe32a1b
z92b47eec557e410860c288f756f82e22e7110991a94c9acbf449cd37c136bbdf1db786a24c5e5a
z41344f7f4dd2f4550963dadc09a74935a08aee2e9bcc4f3bf4bca3b53b033421670d512b37f861
za99d70b8f0a89542e570f915023bee5631ee89acd3d1e2bc2f948904eea76d4fc4f23f14a314ef
z00d8e45af33c7bdd0a2f0c8a9051ec643c4521fa7317227c2f2db457e9c248416a916a1848e359
zd553080d21ad611b682ea982f81f989292e3c2d63d5c9a8317680eaaed897b5572d0ba1e435dd9
z8643e308e1d71530bf8154a474b834c72614f562429a08c03344b6fed7af0508c2730a2250384c
z89322b705bc29c4392a359461eec4c7586b8e40446b0d0c281294a1eac37e1da398ce4394cfcba
za0ef8df28f60489b8e9cd03f329d78c526782612b273ff25bbc378e4af9d0073beb960cec11884
z6513094c22b89dd868a9446a67b40a7cc022925b3e684dfab2fbc62b1d023f60a62851f6278820
z6aecea85336acfd738f8797207bab3482f4d56289f4705cd79a859c67dac46dc7c9278d89217a2
zc8990a91729ddb5972457c66417ea18ea2cb3753d587ac17c173d36db48a8b41f1d3aa5dc04e42
ze85e727ab385baabcdd2450568d50ea43ec58a4063142251bec35536833d121f7efbfad812cdaa
zf6f32f963c1f9ec73fca3d82e8f285db58e9bc1bf92dc2e87642493cd3df892e02db11abe460cf
z267be4e544e92dcdd666cf3727c789240cca4be23da3413b43f4ffcaf1b55457cb795b8bae9bff
z14a53ae9f626df24b1dcf11fd1d350dfa431022731e70760df419fff15babcac6287442612f8ef
za5f7677560e33fdbf97107bbcf2ed3dfc239e52ae249f5d8281ceb619839227e0ecc0d4d2e32a3
zb9fd1f4def3a017cb1a7381a5d6d4472a16fea8ec2beb0a5c179315144decb4fc5579c2f461740
z9da4cd08ea9d9870a869b33bc5bfde54ff2eaad4b4e757c5977b3c1360f0f816cd7af46cf39426
z560852097cdbd144b94d2d418d35e8b5c656456dff11b57424d6c818e5004b560bb74a7030a88f
z23ea30ac0a0726770191067237356436ccaf12ff5d7c33ebf5a30d9fba78890d975cea14d483bd
zafdf3d6259a0aa866aa3de545c53a70a708584d2fafa193e7fe4a904c2dce184b7bf1f8af3a6bc
z8e489f5ff199899940285f699a397f7635f8f0dca506a1e7d5b9bb8771ee3a7531eb00c4a1b204
z258348f0468d2f467fccd7cefbe8c417a5120d95bcdd31ac085f6dcc8e9879d55c2c635d4ba50c
z42c81e9c55ead9c9d404db95b082f80f1c044e0a635236e7a4a21cbb45614b82ce0744ad1a6c74
z19197041af8dcebf646a4e2442a727773045e9b4df75ef35ccc31b88b00a0bf70fefe7372637dd
zc8e41ff7fb4b01b3a43626b883754ee4217501d9170064d0f03ec00ad838464a856a830de5883c
z40ef035cd0051a026f95c869e8bac6533209f63e82c5e5ee18e721a940816c065bbed5920b6bcf
zecc3afb09b2f0638eba3cc40cb34a94c58b3949707bf0dfa55df786d60bfa6ce3a703c7aa18521
z0eb5f21c5750f03939278ec08503796ecfdc97b351159ada8dcd337c05376ad464d32f0736b2cb
z9b023a24473ccd93ac7fb4eabc2c3a4a2d397bcee2a0a66729be6bb0471655a00eab4a1033c2e3
z0d420c5e80f67a9883541c0f9a2fbb160c78221689c5374695abc3807afe0600073235b03554d1
z8a26bb1c153baf6cf77f1e00108f115796f18f43f9e61c68dd0fe4998ef7a1d75d41940d64a961
z6f9855553b5ce7bb95539ba2c510329cad0b8ca948989013c79345b25f3233ed64295ef6eb3dfb
zb73a54e2a469c6f24b91bc32bf7d3197b14a8798cea4b1904c141940ebce5e30bb506ac6156861
zd97e1f6469e5ea940b6ebb602363afedcd633aa8ad3cfb034f404af08a799849ab8172b42dbe0f
z5cd013d56e8329d3a0de39e6a51c77dd46a6b34b47b0a4d2bf65953a25163d1950cd4efc2da3ef
z2365ea71e34e1cbe6953e71df52ccc407e320392bd71fda6be55d6065b007e5a865eaac075f88f
z5b5abcb8a550ed7eee97547ebdeffd65b4089a2060542d6ae33370516293948242776e17a91efe
z675f36f47bd7f4c331ee202461f32a66ab084c92b50a04d9cff46e4997f57c6ac86bca984c2199
zfe468a186f6d82dea95b358cf4aff516408cdd8449f4a2cee95a4645ac2452053b5554521bac11
z219b2a56cccf10326d33f8265f0593f1e8febc491874ceb7708ae963697c8366abfb26ecb3638b
zd429b03d2b85151e15a3a3bd760cba219c1f1e036811b6b95742dd048f2b0a2255e59d854c4853
z0889148124802de95cbc65fb525bf10685c604c676e965619e1ac31bf2a0b73dc3e0ebaaf979a9
z57e033fad413edc5cd1c8e83360fd9650620288ebaa6b9a1a84cbe7976c22b85c9681f3092007e
zc340c79faa5bcc165e41704441c6ce6efeb3b38ee806049e84c864fc2b34f50b92d503f1a47664
z4f4c4266f0caccb0f914de777468b1aca85981de9e58bc0dab87982ae6fc37900a9db9663ef5ef
z9f67abda2e0be0ac666926c18a659fe19b295bf9310d06b01fe2c321019f4d1247affad61e73da
zdd4534001ae5bd05608b07863aa37cf7c4bb564da9aedb4141d667b06ff0784f53d9d4eec16831
zb0e55abcbdc0dddbfbc58fb33871bdc259cf3d92d241bb3092d195c63e920944642d9711943437
z5e4e946faaf42dd1ec23b3e64dba8a246564fb6826b8ad24050a24e90bb493fb43b1225d119487
z23f8be0edc66bf96fae983a327af6eccb381343a8dafbcf432c7be7716b6825b6a5a618b84cc58
z1a13232805d536a050d21717c6562d910eec94aed352cdf7bcaa5af4a5f26bf9baede7f86bd3aa
zbb4046719e7a72fb75300240022f6e630b6cdd311d6568697492f4f8d232748deea0037ab3e07e
zdffaf84956692c89fc0ccfc52a38c27e0ce74c51727ba87e807abc567c920f945076c6a41027fe
z106302e5d8322ab5a0a7a8def74025debadbf82cadc8bd99ef008ed86e4b769c843523e3cd8e41
z059330f489434117117c07a15db28734ca83e6ebe1815ef1281b03f6a869d7f43cf4c558bd1d1b
z33b5534439824cfaf7fcb6fd475250f809a23b553b57c2b87d315fee2605808459eac70f70cf30
z8966b0fc98616e04503ce044f38649c42ea22a6b75ac09b929f5d714ae8e31a0344f42dd7bd599
z2f409180fa081bfe6ea45c6a61770fd600cfef169e89ca5ca9c1bf4d2325757f92a5a383a44450
zf0cd775478bcf921c45e307d839a0fcf2b15f43215aa62104137b2cec37cf219e809a4f577523b
za987207835a9d1c11c2c5741babfd595b001c714bd502228efcad0afa413d7d45899d1fb551e6f
z76a354416753fa9bab04c1520cee0518153a7f2de1ad7398781957e9c225399b1e26f6ece3f01f
za18829fe969d0147f6d400960bf485e048dcfe8c36a43394537b22f0aa38ee5ed2aed54bb37e89
z6d7f452a87e8937518484c6ab32f30ac923dd27887443a4740e4115e67fc17d59060d0480a8253
z01a10943b58dc894d8e39038d0948c4866a2c799a00b6c3ccb8f78745bf4660cd92dfca69e7fdc
zc4b30eeafabe81c8fc8011c4fe90de82d7484b09356143fc9b584311cd71129edc070881d8f494
zf2cb6eff945e6513252dc19a2fa448b68b7c95eaa832df3b85e70b75b146a6123e52d439785a4e
z26b3d548a1e6e7fc9b5450b1b1a6a8132bd7038630edb82c8fe08617b28c04b367b2b49e7714d9
z03f244303e1709265ff83aa2d0194afad55ce9eaae39dc9edd1aebc56943962bbffefff2b5502e
z1d5738e2eafeaeb2e3d351cb1a6d57201e1764395f0452c6f6b6370f721801f03bc5224374cb0c
z764ba521f45127139df41f5819c8ee2143051ea297b4cf2b72cedc2f2a62bfa0b192a73cd3ae9e
zc8cfc0b065a4d057442fea9f07c4d6594367fbfadca5be79e3bee59c0d8b84922d193a7339dff2
z636d0f25e31eee819e5db98bb76f37509073a833b9ee9bdfedd4164a361dba69a0dbe56d8a671a
zaafc85b32e5926c82d5e0503efae79eec8f33669ed5f5746d8c7e719fe37d3a12cbaf3bb3e2a34
z74cedf0460557c45499678972cf609d95515f2967c8b607fc798533221f6b7b815c49bbd1e460f
za8224f395cc69bf6d8aec2f59a98e0730b2104a6142d1a4a5ad16ec380e95cfdc0a0cc40bb0f82
z6fe9dfb7180454dddf245175b751d76aeb172e0d9e90d55f66414c677a420c06dd4f1bb23fa1e7
z917879c6bae83f702b26bd33849d43aed13d9ee6aff8cf85a1e26c4362a0de4d3aae8b566890a3
z0f30729d48a113c3426b3554ae0b840f7c23ab78f759c578a9708704fbf5c21d8b1311b0252bbc
z40dddc693bfed79c404ae8783e32f8a0a5c9196645deb47b17268a627f780e027e117236e05263
zcdb0a5607d021c9ae14757c4d5bb0abfcd588d777bfb95c55e023863c0ff22111a1710a2c2e1b2
zf6a7a59774ab5275b9ab7093cc9650bc9d47d6888baf0fb75bbeab70184b98e4cce6c3d29118ef
z4066faac4e7c45d166e406d6945284f966abdc90468f78fa08f2d6617901cd6a09cb4b62b9e222
zbfbe6e77fd49476725b3363b48baca51efbd69fb5a7e4508780c3b81c4b094fe324e53777576a0
zcc3d8424b2dff5a4cc2b15de5170630f5ef3838a049c06ed03c5ca6333326174f588219b2a8e0e
ze194b32c4aaa239ba440e3bec158d403d96f791b3c1e5cee72b7d5bc8e08335e3ac086ed5955ab
zbd6a99f66ead6f2bff62effdedd817ffeff4904cb53a45a361a068196a68a612f86d62a4cb5b62
z0a531e63dc89244de745aedecdb03e8ea1b6352f56cf3aff8b62abcfd38240b06e554a20dcc907
zf3f47ca581ec8e78710420ef10bef3730e4ae54255e672a8eaf5bbfd48b428f881a17c07a108c2
z73b65c81d74e7d9792303333c9b233af072595007d083689817f8126431671e83f95ad7fc93f57
z5c92e548a360719c803880db13cf5ba5f4bc8263b141f3ddbd64aa08c9ecbb45f633896b8f3a47
z6b20205dcc5054872cd66c55965d4eff35d18963bf4b675b407ac0385b03c392c2368560fad478
z75077d98e1041319dc1079d8181fef8e75e0aee822423404c02919c1a400a8eeea2dead41daba7
zb9e48962cc9e81e3cbf395bb4cd6311cf3c0dc3b72336c6c675c389c1d35b1b8c133afca9f2244
ze1e3d11b923a238408ccba5456df91c87373032f1d8377cedace504e22dda3de9f4a6701b59ac2
zca339e41f1c7288b6b6ed170657d3bc8a30c904cd407f72a312990ade7a457009cd32f41ce512d
za1def8ee9db4296b6986d6784f5418ebe105a0e04df741b00d83eb1b97a92daede9b8b0db7a0e5
z0358797bf7a2519c238f4501c1ccf94cae3cf7c8ab3fb57ea9ee46d22816a26b86862d62309c35
z42714aea96dccf9bf9ae48c0db50e86d68321fbf001d6464bb73bdbaba975d031c3027d7e0515b
z1ad73efa140db79411dfea0f29ec040a7199ffa7fb4ae93a13a2d4f5c5d8acca4d54f98ceb52e2
z757f207029f3026720e5766ec0e76f3ac103702d31cc2fffb4a0bf90f76c7041bd1744980c9ad7
zf655575243261604132a975989754b44dbb000fd074c160ea9cf3ec7db5c1d1e50bec1843b1f54
z177d61551866d8717f0fb19906389961dfbee4aa8ebe231732f7a6cf266eb9602c2dcc0f78979c
ze1662a551199997098f860720e47b050d39865a159dc394f4167885ba8b4e0a93d4ab93a9e1811
z32045cb02d26b3046617168879ef9b39f264853f4c452e4eec16f1ecf9ec10c019b47f6c4787e7
zb128e9a9c68de5e4ca0bef36e9c7839ab4821cb04a004886eb2020e48efdd5bc5312702ef660d8
ze4ce0052faabdc909eb24ea25d6a9d661796aac1cd1a067966c7aad26362047651b6849b68b291
z5d2dd13c13bfbc74305f0456db81f8022da7ce353d6e927913ab1a4363b8947fa2ca7b1d76cf8a
z18ee2b429c76e0a7edaa1126a545cf0551759ed01cb157c2461d806c5df71107765b7a72d5d5aa
zd718551741ab7d98a70701e33dfa87743df4087e2b18315984d94d83b920f321f5f38677a9e121
z2d6e20a04bae923a56a78ee450568946b1ba63754c2d4a18fe6d91b1f60f394f80026db3df0f76
zabaa5d0a69b8f819fcd5472143e4b521af919613a4fcb084af7d62c681d257c1f6a0f0286ad408
z6de7a29686edf0950cd8d09e69ee35391917a98c6449faaf73822aa4e6acc7c1bdf4f5880a0f4c
z1146edde18437407baafa853a42ac472cca5372ab3e84607549ac28a3dcf7b9468d69a8c914d61
z328314f123c4d8d788dd12a243352f27f2daf1f7b368407236c69fb2564afc96af5c63fadd4c25
z2b4cacc277a05e11c685be83f0ff1d920d3cb63da15d9c6d10cfcb573788ae19d459683ca0a7b1
z8cad3155a4993c2ff86fa05137f1e72563baf74a2f9a0d078a4bda657e1aeb3d54efd31b16033b
z5867236f1eec1231f54cc591ca175158ff4ca6d597a2703b95a556e3508d43f71ff37bc38181b9
z7670b7a9e16eb9a37b6f906bcda698670400f34325aaec9d41b5ddf3410a4de5d6fd7c48ec364a
z627634b951608b91fcfc525cb870287b724a4529980ad3c78267f565b96e138d1e70cb4d7c767b
z7819defa762d67236ee36fd139fcd2f3833d503f662b8458a44751d7087627e0664165140ede78
z17549f5642eb6c93cb9fdc71f49943d366a63cc3f0e062546c4f6fed0453fade3eea75dad8fefb
zb9a73ab16b3b04a591106d78c0122a8eb49b93a7940530b31ea9608e924483dbd58b3cdc043dc8
z6b0e49947857a03ff6ca9121405b610cc83ec9c050fd84bcd3a5a41f49637086751feee020be8a
z8be6d4d1678984beb1f8ba1107be9f30f386dc1e9586bcf006708fe8233c0f9de9aac3f76b16c3
z480710b8b9fca3cd29d3440e7473e18069589c1ab675ef5298fa94b487489278556cb45d8dac0d
z3d13b7dd7fc89660647067aaee0d9b94de6459de9a67ca04b209c31bd46d1da578de44cf518858
z6150e6cd8d7855434065e3916493062a934b1164733ffc73388fafc10e7a7bae243dfee86f69d6
zbae793b6af88695e592c3d7919eb4af8d4141579fd5eb6f93619ffbacb8a0365f7cd05416414b4
zb0a9e4a0d2534bc122797e663a5abae605fcc0cc3a3aa1f46930b6e2c89a2a0292761f0279671a
zb1b271f64b9ab38c99bcb9849ac7d9d5630263f07289b9f26feac0f506dd743ba8ff327b75cbb2
z1883e1da3166f32137f73d0dc4f52cb18ca68228f0cb6f8905119ddecb00f13922947d6c1e6e67
z0800787fdf7de579a88b96d7a566c754f27fcf1283ea549201e615538be82a8f9b3ddbadd7c067
z3bd84cd90f9bb39620511c3790a173c26413cf36263e5a5515013e914f311e9f6cdabecf3a1520
z5a6fc8756d877a7f38bc45a4ad125a06ac66e33885624ca6f827eeeee311f40cb5cbc1033719d2
z97d8f220b99d896e7a1d6c9b8513e915ba751beb1c6f03e67505546e6fe9810f3c12850a18ba8b
zc281567ed5aa22b25ec9dd48798261735b0b246addc4ae7138bc8f36e04653db75fcfbbcc217d0
zd1eca529aa6102979e6e5f1780a1a7b7684d64f0d51166ba49cd358e9c995e5328a067cd202d61
z2342df7c2ad8c12e6e5bc615795221222c84345b68ad58bb07733ac9bb13b1ce4fe30ce0f43b3c
z8a3531d9626c602846d1b63ab17a7ce5214b87a7f2923a23095633e7a12c670da74ca469f1c140
zf11a0bb8dbfe3917397cb97df222597471289772bc703d4d4e0676bf4722b0d20b73968c855996
z85b3c9c9067af38068bee5b328394bb5ab4b9b8b1db91c889db368ad325a53a839d4d7beff93fb
z811afda9b5326f557bfcb2b929ad421783e5a1291943db7d889f2ea776447df14f77eb5dc412c9
zf53846c78521a7f0e3e495472072039e18235290ceb13a1dff9d16038a6c14f0fda96ca55eb50e
z30d7e8139ef0e76b13b096641d4905974e564cf2670f2d101affe0ac590a9644ee64c52c2ea1cb
zf7394d9652c2b6463079c29ba994e896c24fc34e98209973b95027bc5eb14da1a35dd30f627313
zd1fb7e91679bba6927d08cff2cc58b74c77db7fa9766b3afff248d445591978a1282bd12853769
zd86dad6dab3843d90025f4ed5911486753aa2b9379fd57deab05ae2de49d1e43201374f9966c40
z9ecde31a6eebf0d8337aeabbd57c0a9a3363a658c52791bffcb7073054276963e742ff6cf3208c
zd8af977b0636e778faa569a30caab56b566cc2939a06810456c3d3691c6f51a10470e8f57fc9ed
z7a4123ed92ba9dcf60fb43deed18d198245317288492830c3f7984d498627c2cf228f49bc1733a
z12d86fcc8e3494eb89e11a516f8203ba4c13f0f61c0cf78f74c522e5ecd76e0f59ed225b1115b6
ze9b6c8170a577d13fb744da00e28f4d79462aa79b30f446f6676dba426de783db12d08f88b124a
z1baeb8b66213faee36f108231ef7b3c6865a5e05627ad9fe1bc34ebed2eb57dcb5a753e0dd1f9a
zf8265c5ac98b84fc4aede48788586f348ff9553eb5be3b5f340c2e4b72f62d59d959c9b7b320b1
z3b3fbc1c67d62298e993beee4f2091f6154ba08db4ffddf99eca25527a1f6139245a4622c8076a
z8b65d2d2a71f995ddd1aaf28fcf55b5fe436ac43b99814928a7d1aa9353483f3f20b83725bac04
z1dda0012678a93cd607aa471e0f68251f0c37a4409e9e9108435f184b5e498626ce09246743b2e
z388b7c6f9955f601a3a973f13eb828e9c624182ef836263acaceef09da598b1e4f9fcc55152450
z76ad5fd03925b25aabaf1c27f31809c7f3afd0284906c6c618f154530b1018d79a99e748662ff0
z5921f8791858e52196ddb452be9cc6443e1c051c7f81a5b596db2818cccdef7fae2921cba361c4
z6b5e3e41680cd6067d2c2a8b406ad85a2c2322b70a5c5f23c736f95c1991f15b1d752fd359ac81
ze445d91f55e9cab9ccde3be762feb4f0add1f275c6ee178d844a06d1090fd547284c322bf6a2b1
z0305a337298d646692632babbe15e976c38f10b4c9fda749a256b4c4dc8bdca1c142abbc2a5ff4
z895dc1e0d544b8fe4b1e900e666e04f29bff25a5edab68855577219d149a3737f0a71bada1a46c
z063b2322345b4c7b23522bb81318ea6dd9d37b1a77b0c085c60f6ce5a360b1e00cd53113028687
z65e0a9e3b950205a24b17ee7420c41556cfa1a46abf9f22961e74bf5422e120f7900e68e4a295c
ze20d0475754e3722c30085fdd38213455d5355ec98c1e7a50ddca93fc41ba8ac85f073fb364cd6
z4703bb90ee5ffd4c0522767235afdd09bc6709e6205599b79d5dbda7f433cb7a30746e1f39a11d
zb9ce34a05a1b7a82e033374d1320a1e681d497d1f9e754d0bfd2956798ec1e8e8874ed173df14f
z8c996894e1a48401864c8673dc54a0d9015ed49184d5a7004a4879943f44e8518c53fbea039b3c
z5c4c6d58076051f91d0f1107a9fa637c24a24a141232429411f372a3bcf62b4c3a669644bd0c86
z88f0969bccbeebb6b31496954805ee00c2a0cb6912f85b165911699de74fa09dc5a6c163456e80
z667ac90fefb263a4841b2bcf5cc7031b1e91df206a90bb90ff6d9342143790c57f2350a6eb3ee4
z5d7e200955e5faf1b77c77f6bd23d27c61264e2c71199c3e70b785357d9ce8563a7c5d2b499266
zbbc3790027883840b76a1be502e0944391e0c513f893e5fa10767ea451df81918a27170ac5e0c4
zff35597347b8287576bd87f9744869ffe262d261f2af588b40efc7dfa6b818b8894507d365dca7
z1ccd55761df637c1ff1efa7d244fb8c4f9fe21aae9173c39b218eacb7a368ba934737ba67f5511
z455e1f2ca79d4388c348a4105913541ae82dbf9e57378ede799138fa799ded2ac7ce7d3aa44102
z493b85447b2717d7a3a57912d92c76a05e8fe7d112f4921d6dc3936cccbe7cdd6b51f887252aed
z6d4592ecd029f74a83a0a0de314cf9467ed7216b6be401e427df30fea58409c20d3f5c69c1c387
z37397a3174a895a4aaaee0d6d168f6ffbf82aa2468fe026c93867f17efdca2342435b6a5ba2ed6
z38fb162c1044231507f8f400e0a7d6748207d5ef844a47a465bf71b3c88520dd43c82836df248a
z7a6ed0318b5e25a7ab2875f1e7d73fc4d99924be8e2564bf19c588bb28b1022db71bd91dce611c
z1c8829f0e73aa19de02f07b406fab9da518b7fe696b272a9fc71a5ad6c09402ff21d1052a984bf
zfe740c740b25c80cea34a89d2f07fc5e60142722910f41531b1dde82cb9fcd5d43206b586f071f
z7774de86118dda62886bf2a7750de8cb9b96318da4db8b362b95488d446d914448558eacc5a527
z423b61df090e10e72a43990dfeb8f7210b1a1254d860aebcc4399dfb9384ea06f8ad99ecee0e89
z0dac2ce02fb2cbb5b14d3b741c793084d5e13ab1f51df5f864d40723b2969fa09866bcf0e6a1e7
z0f534c71c9a59eb9e00a6b7cdf59ad13ee120d158e12aa14636d718f5e9c30b9de4ce886a14818
zb1c72cfdc1a28cbaa0407f0275f5cbc9d66c2b8d95dbeee6304b2293dd72bc9e09913081a8b67e
z809f3a9beac39a857c4bbeca23b789792bf91ff0d249a56ada0269bbb25b78e0c053095321a8f3
zbff470c92335acc03504a5517483ba11657d0fb00817e0e67a1f36f4cadbca1da47a9415c2e1f0
ze542b21ae5d5ace543e8dc02adc763b0f3271cb9886b6f7ada89a97ece765e8bf67f08b2bbdbca
z1e6298c5dd98a624fe68e07c99847fb101aaea66c2b0c545d9b76ac473a641500ace5871871ede
z96b953a16d166fc7f301208c7a0a689e4a57a18330cfee4d6bb872a1468b902666122431f175f2
zd01bf2e60db5484028672a45e68fc546c6cadc3a3f02d5bcaff426cff4cc15a67c9b422768d389
zd4773cae235e07ee1f46c8f4850e489509202e21311bf1876e0291f6d9a7fcc8deec7e3c618090
z486a2d823bee29ff38acc767b97b041be1249a34c981a68baab955c4bf840c17614282e648ca11
z378a8c69128fac6e6946a0a285e9462b623f05784725bf8f1dab9de7abfdc725e98e3cccd2db4b
zc6d270de2d5697f954102d2f980870daf23fd0bf6e30185f4c47dcb07c689b82bde37d7b920c5d
z0ae628d96373d61bffc9c3b60c39a9184b8a778fbf2f8296691bda31aaad5453188a47e62a0a0c
zeed3b95b47d27c40bdcb79f168b780f5978de345986b50eaa8b649d4091ec28321e70176a03e72
z8c51c16e01bd1f1245933285086de19dd3f25c7ac6173bdbc6bda24bdbceda4703c2237110a710
za0132fc4fea72be1bb27d18556135085a63e5e3432b65c7deb1727841f2707b0a9f05197219ef6
z0e7f5a91b10ae48566e1b870f8aa3f6a08badd702c678c0a6f0bed5926b74d301e99178e004d7b
z505d752f481f59015f1c0895f884b51c1bb591506e1e1e17aca12c536744041c21c7f466e70ea6
z2c7ac999993783f83be8b57c83d069860b2ea8e238546bc17094a80cf726f916e96cac48e76002
z59bae54f1a8b33e1cc8dff94e5dab493214520b709a099f89292b406931e9985ca3e8b2804ed51
z6a80df9eadb304f1f20d5cf2db5b2d27c8ec0e62a166c846db475cf3675f601933fbbf625e5597
zb21e50d57b1385a3e5704b011b9635ad7e08663b52ac081ae95aa6c8838ea51478d9ec1bb02da8
z44f69fcf6f32c181da127f8d813b07ecb949c514bd0cbff06828ab777f4b373ae3d1a4e8cb380a
zdf8d8c26bff3798d2e9e059921e4531681ad138dbef0a18b0fde6bbc8dadd4cf7465d5bba6dae5
z62674a53f309622604c696392451dc60bcfdf88e59d780967a2bc5cdf8a2c4beca3e24f969076f
zf65f508de31ccb81849808e8785a33a1f6300c4bc82fbf1a5c7cec2d8c4af502082bb8bb18515a
z6533c8566b417c5966362b379306db8a8ebb572887c32a9919592af9c73f8bee25ede0d089b37c
z6f85246f1d88efaa6ef32610f85a9c9fa8dfe63ff1ba0b366de33d002ad114bf2f6464f8e80c7e
z7d51075ebd80bd0406655d7de485bbdb254bfde9d520da0b1c720f4e43d95635e67fab9c43d9a3
z1a6b8ee106ec55655d7d348560e38f3fb187eca7d6b0e965be4e0720629024710af41cfd869611
z400c2ac728a9ab38d2835173a1c687bc7fa20bb426e583cdff1c39d5a4afed91f16db54a596ab2
za64c4bf997925a2aaf773de23177b3f3ab02e165b936ef679ed706adbc475d9ce7d7af2c2fd57e
z601479b63c136d943f9dc8616c079d8eff14f3bceaa7fc0d649257213778c2cdbe6da2d47a5df3
zc7d637480f82a598904fd4826f31197d94a611efd95f14e2d8eab1c1b443b7d8099469da63da4d
z7a0c377b9a0f2f3ed4f4c5b07fccd59fccbd18303b7a5c4e626854eaf73085cca1e75d123f30c8
ze4fa31ace1d9c66f2510900c47d052fa32abf61a027451bd637e94fc5b7aae8bb84de05477b908
z3bb582c814ea1b37d1a2b1006747ac2f4ff3fd2677570e2e5f6673ce614edfa42bd0f48622f542
zcf9e041ecc08b8b7d2faa0db2c4617e9f5f53ef75906d269a3d177bb689c1df0ea78794d95798d
z6ab495b4ae1299239ff3b407bbb849fe42f39c739f510d8b6a20bac4d7b4150ccc45b0a9fe6a96
zaf486b3da5c59d12cfa0702e531464f0ac8b4bf268667a1b8abb39bca144f713338e8ad30ab722
z04b3b27b964758677817739e5785d096d2dae209590d2f5c809a6c6dcfa3d21b394799288d2a6b
zcbde0ef179b1162a152d33d5d4e0a8c948586c6d2eb5ff45690c398195ae78a0ab6d60dacf0dd4
zcd7a4bca3228b9a23637058bb244f64d0efd3e259145fa5824564e6d1f19ade88b0db50aaeded7
z72422a86f4791aedaba2d8234ebdd9e604006045e5affd4ca7d4ffb09e28edd49e0d996158cb63
z009cf43f41dbfa416110b353ee9cf428c91c641ed431e1c852898d2cbd4b2245f2927db2e9d620
zbcd631543335d99e3c1589efc65e6186ff0e584f2e95616650a533079a32c630e768592a2f2d9d
z76a3ff7dcc83b80aaf4bf94bb2df99adcd3892358b0f6255e3968266f7ea5b92da672bed65255b
zf72002e0d24718a9849af238d0c40e7d03ad7419f2f589607474fb8d11e4975459f8a8c7d464ed
z8dc2e64ce1f068f73636d8213210a2f3b1cba2e54a93999371dfd602bc2ea31c75af8ecb8b8f13
z8a0d451092344c4a0c90fe5aa7e7f748f95f92132ebb5a393519f149dc384593c5bd3611a2be64
z84aa9fb8713bdf15097304ec89b085ab2f9e11ee85fc2c296a7d98811eac76cbf259c768a1e140
z5089ca30ea3431e2510df9ef64b980cc3d4e7398ba0d60bafe303de6c2dd28b2702715e418fe76
zc88fc07b61d5a7a0e56582cd4bdb32bdd5e0032150215f0274b59c55d6105551a1c55a7d923e6c
zeafc7c84b90eb203b192bb41795b084d868daa86a79f7e6dc78d7be73a2b59da7a863f3d7c6616
zb75ce287b800a6ab7f185addfd8568ac7c24590631c37a09fa2f4da81695c462edb80d4b97028b
z7c601c088cd5f7c4a4fb22888357c916262b29439177df68df52e1fb4b5f8a6c8a653c5cd89735
z776390372788aaf748c36e7308d7975ced769344579c6e524927ba3f23bd88986a00018a39ac65
zfe5a4f056feb1a916e4f21f1361d3dafa32157c37e94788a94a7ca2ae08cfbb7edc83410ef9108
z19c1486961393d98b25f85b5bb75d9004c1d600c11f26859ccff903684bafa3458ec26ce566df7
z0e31b298a6c0fccf87407ec37e4f22aa8f97ce9453a3b3d616d250d8d444dff1daecb532f385a6
z6a52c4bac9030af3cc75f25dd8ddf88b88a6b833b2c67f107a28698ca94d52de7377d165d2a7a0
z0a8ff4085a8359150eeb3181d44862dc14608715fd0a50a3af9bcbc691ec195da948b6293a20a1
z785816e72c2f6c6d5b71c40c8ce554f237958c505f1da9e5a8525aa920ab8d505dd53db4fc2e5e
z8372f9dd9e781d1480aa99192414e763b07e33d5b62ba1c38e4ab62c05c57de15dc4678083120e
zc73f4a674674183608773831a8f463eb0d6b5d2c713b377160cf32001bede7b89b9ce9f8ac8ef2
zc6499670bd6e81395a9625f35a2a4a3e3bd9f39ec3b6498923610e6c72ac1432f24204861f8358
z9006081d516230fd21fad013e05721148ee6f01354adccbf81794ddd146f4b770e383866f37f70
z10028cff2bf7cc1fc8e9b22d9fc892fefbb39f350920b1543b1b2fcf7423a0410bc021bc34ec3b
zeeb3aba83b76c20d6097356970aa5cd065e80b7263a7b2a5d5f6de396ad1087b8b0f0540e2334a
z3ac89e41f58001330a884d0ff703ae64dd33d239bbcd74a869cd16e543a3d870464d86479a7d1c
ze985c7cbfc6fee1d09f70bdac77fe568cc903f0b60f415383c4ec67d7bbed539f802ff3c9f64ea
zc963cf5f1b60167678d47eae5bf05acf415cd6e388a707cbbbb7a45fcc466ec1d773fca93495ea
z8b149589698afc52d97a68d2359d126f7d45598472a7bd127c0fbaf0a4f04991bd5eef69e081ed
zca232b3a927675e0e0e49dd232e36c6410c41056462b851b8dbfea7606199832fd99bc44dd799b
z9ad47d13fa13abae11110d57547e39d1a277c67fd122f141793ea87929398ee4cc5ecf99a18697
z6bd2089408789cbd5192a882e218d446ce36b49cb2c0590fac551855ed84e4052d1053b84b1717
zb3d0b12f328793b404262ba9df7d6b8737ff46f7bff73425688912251b2c91d404e4560a8a32b0
z8301550ee1a0d7eddefcf1fab60a05c41f8f5e301560138939db6e649045f28f07849bdb8016a7
z12273ba8c82607fe2c92302b732ddbf02d46c88af266291c437a4cfcf630847704ee216ae66f4a
zcd4c5600058fd518bf54519d5b3cc2b0181ec573b291bb09a465f55d4d8d05b659d13ef499eaa5
z7f4af11d1cc39d23e1f4ecb00bf44713d04307749c4f91b7a423eb5401988fd3b9eacb38726053
z6b32830874ae876c16c2e1100d68fbbc5ad7f39ffbfcd50866297d21751c042553c4c164d21c61
z640d3f053ed37b11443e31501ebf8327554201862745f41fa09ab9240042d62ae0a11eba5e740d
zf41a129937cadb67b25cd00e30cb873e7051f11bdf79e91443aca0169374d84a3fdde10e9ca219
z2cc18d402c81c8c9003d2148dab828288d046dc4ee8892f0aa661dbede4bf98559df522b64a331
z5802747e2454795124388b62424554abe3c41f24ecdbd36553b19a1e5e8223ed43c4fa30edf088
z221392fbbcae358a16114ec515f605453a79393fb91aa3bb5051c30510123c43c7a703d423fbc9
z67b473b8cdd4478666aa9e2d594b7558bc4b28e76f0421c0f8d4e7cacbd68de766d4af789216fc
zf2407f3ae211fdd71267de2f6ae0cccf57e4eb479d4f667ec19afd0fe0408c7cfdc807de1b9ebf
za1d9f587b55d2871c4e7f88412b32b4918e38466356cb98a1d021c012a938dff0c05dd0329e7ae
z56f8f03384ecbd45d96c4b84961d522a1b376aacc8f169e5f2db0effb378b9113d43343afa671c
zff1ce49df1b5654f8e4a896434365f904c753a9385b150accb018e72d12ad47d4d7899cdd89ad7
za094be4e91e8271c7f59d8b6f0139c5cf71a379e186f8021790376a87da884e25a1c60d5805102
z18d62454bd66ede6f743c8ba1c6a5fa16d830416b7106bc61d3a850864c0d0cd3d42dee386536d
zccf0b995c1142d67ee427770e89e6dce6b17fdfd8c285f554adf5ea6c4e3cba3ac92e38f761157
z488e8cd9ec8139b38efbcb7001658a62978b2bf081d5246b633aa3cda17a15da9233e01f3ae5ec
ze1acb0bbae21362957729781cf3eea8045955f3d23aefaa4af6d17731035da8256a6a32b25556a
z34a8f34e9db526cba7c11e4cb5a9e2d00963ccc5f8bc06d2790a2cba507915612a3bdffeca0f1d
zbd1e02fe97315606013c6448eac1b518b9f4dcb761961e73ff06f2022cf5e34c86021546d405e7
z2cde631de44fcedfa82f04cbd0f3635865732beb42a8049fb28537e51bdc3d095d93a4ae818d3c
z2a319ed8867a63cedcfdbcf674e21f0e0a641ad4ea097a08701cb1632db2f9b244d0c0e85da72e
zd54772331fa2aa8169d1411a930cc136e757b604a4926911d80618fd27ef5ae9272eb681a106eb
z20a32f34e1c5b9eac78e992b6d767ab75bd44448aa061744cb06e140a9288540c0e89e3e7977ba
z924f208b711a9f9796d15962d47a6cb5a13849f0a9113520422ac7feea1fa9902a1c72a84f88c1
zd60e10d9f28ef42346960c0be4c2d7f558fd6feda00eb3cf016e200637acd7606f190cfa9fb028
z1c3c50d7058fc1fbbf3af59a65fd98e0cf5d542d74abcd2132b8a64daaca2018399578d1fbb2c0
z9b00b7ded7324ae34e153dc7332c0d64f642ef788c0c5e1072745744ef7967244005ec443cf1e8
z178db056c45f3d0ced1fe8393ad3a62aeeea06d6201bec61d524b4bae1e44d7465c30b03c28ba4
z43adf8d5af07dcc05662b3e72d0b2db5ebe73c62b2abf1a9b7257d18025579a551565013f0ca91
z7126775122696d7ca971f620124536d2f0f525a956edce7a6e06935edb7277cafb4aa2cea9ae9d
zba8c0a9076e3faf3d80935c9848e79e91749814e2ac4f56614bbc3ddb3fc216a226a20222a5a35
z7174e6c419e929621050d3b3b97b50899a557a8f1140786683e0278e25fc6e47fbadb31748e451
z1ac7431ea213ef253a9db8005d968d3b6cd658268ad40c6348cf4a624cc478cb607fb67edd884b
zaae7fe77127e9537b8fc0d7b97ffa8cbe255d401197b9bbd3eb8095e947574c54ac5163f8a5add
zc4912008bd10db9e887093154c391bf6467442f779721f554069487f4f71bbf61c2e011a6601db
z75d3a5d9d1cf4e857d739eff28cbcf7941b78c60c39577318d79ff82e96ca126ff7337cbd80ccb
z7d52320be0a55ab030b3a0cd4d425f060a6847417c5e16276192ea97e4554c2cfd553b070d1147
zfa4872d5781f07eb857784d0a9e8930cc94d03b217236c655e2bb3b79397a0c9aaf4609f3eae30
z28385e34d7355a64ccde4a287a39067051911a27c11929d35819ea9caf7421fbfd42baeb00e682
zf47368e20990e0364fff7fa0d83617901a21297329342377392cc852843c7b47dff2413b853358
z36ee1054be781b8567a14735b9bb16c884c9f0205f0941f347f893de9204d19732ff1b966c7ff2
z2522fd847a84ffc67e3483ac1f36939ee51aa316ff4342d848959df490193264aa38a515907cfd
z519364c77a923b01f95db6a6702d36a0d2183073435d54fe587babd5a727dd4d1f268dd3c74209
z2756000d22840f683082842357c6a046f8eebfb94534668401aea6ed046f1a22d04101799d1141
zb0c648ac229e612adf70f56eb4e2c1251ebb28f2b8a3154a4b4fe764df82e3edadc08bd691855f
z06b10cc7bd5a63c553edffc296095cdb756b6a0316b8bf72b14720502f5d1c5c38ea44beb2149c
z747f68ec1f60022e7a1ca137a6c62a8c97be1c677eeac8050d8c563c2f09fa9c48a72f98709e71
z0954a9c09829160cf4f20db688d5aeadd6eedcc72dc874c9422f868e6265949041e27bc4a48aaf
zb90e882cc994ef3b66b3c3057a0cd4c643f2c04d03fe9c6d224ea772093802a98650b84f3ba544
z895d2ec660b6514f331783b8da650e740feb8f10ad3a1e47039be56f46162ec86efb29695dbf61
z947aecb4e57658479a436c7a2bd5a96ddce3cab19b02d0cf8eb83d012f5aca70e8b498be80bde3
za385bbb1e2c9c037415884832a3f7bde0f8bbd977525c66439e8e6afdc39c33f443a8562a5eb85
za603cc3f6ef1671240509dbb41cb497fc7eb441c8118dec2d5da98e12c5b34a67597ef2873e4c9
z9bb44b63b440195c0a3db4b191b7fa10503a70b377dd16f7c048f7d9ae68c6299b75c75bb39b7a
zf176f2e46022d274e45ae936f898332682abc4d17a39769bee65c21b222e765d55de03dee5f075
z9ebef2bce51bb5ffc7efee094d9ad780b0d3f1ac90d3d1e436770cb5eba292befdb640fd220e54
z0e8cf7889ab36d4da2cc0f818b9941eef347d769235c577957c02ce9070e74c695c676d8bfc2ed
z571a88fec91473e1a459cb6db29b17ade66ae96be100efb216d7c61cb5afb686f176f33c7a1e98
z0340bcd0fd3ea0c464b9758e0dc31a64141edb3cc89fd814984b7492bca4f616b410e1910544e9
z5c72afdfec43584316a05757cb29ab233ed6bb12dfa76907f75ab11a8f6f75616761d382d0b91a
z44bbcb5592073d08df048f46a68f5ca0fdc789b57091f9912e787f387a4b23835d67a0d69049cb
ze607f4d56d3eacca7e54e980b64c2b4615ba969e2bb6c93fdba79dd84ff96d70f6abddc89de9c4
z2edafce05d493272fbfb8d078a6f003a10f7fcc932c046c33ad36e7b0a9eab8f08be1c40dd036d
z9e2298cfd774f200a39e00d3cce9a122e573c05fb0e38727ccab9269e377f989227373c34d8bd4
zaa0adbe6caa8713e261662f871deae31b897c4faac6c9769df562d730cd2ad9837763206cd5e07
zb26b460eae1e99c50471e4bbe2ec6154e5da9bdb5e6fccdb11c30e0c8d4877c1015b18205f8ecd
z0adac7004ee8ae1bdb428b09e9b07e9c7e53da3e53f19d3a21e44476fff8bda329ff166e79d44f
ze26d84f7dd392c9bb03c62b0848a69ffc4104e76a0312cd557d6ff7d5a47c39cd4a21ae991803f
z0e08bc7cb4ee49c5f4515d3c6ce5072a593007b36e4f914993b65d55f9225af0bdef034978327b
z4d67c441c8f38eef29ebd2eecc90bb7c61839c63249727401185b571b9bcc2c5190655259ebcdb
zc80b56bb01ac8fbad03d84d3ef6514aecd7817089f4aad4053125460611107ba4201a2289c3294
z793b439c1f72081033f2131fce925f833421be8e9f0de25df0d884dfda51c30fae83c33e72946e
zdd1ead6510ef94b3e83e3b03042f9d6e2359fb4947c0bf87e2db32c5644b271d9ca7f17cc514cb
z5b1fddfd77c575e7bc03f977656bc45da798b0dc81b5ee336210eb093cfc6c44545d071a6116b0
zc2018812260adfc6f49218b2093dc3b0300bec6e74e6355d2c289048f54da5ea4884087b53def8
z651c69e2dca1bc16e1a60298adce6a2cf7212623583da6f250d04521b740e39b2c8f00710f8e69
z241302e0475cb5e2acb583ece1352ca5e580877e428d31a540f5cb43dd7b609a9e0824f4288875
zed79b8f7f36c7e3338a60df05a37308823c5a70a00e7254498754b0fcfcde6f25cab6845892ca2
z9010d3922521514907aa3b3a2c5e0203fe88a76004daee49cdf9d2eb9300a06193355868474366
ze6312e09bbe5baa7ccf6c031709074cbc795765f0e8043a16f336b47f60ae466d4298c24ce2983
z477b8aa2b240e34617fc4fc26e8ba93a224370a20f82cc969c6746404644e33ce8a0f294b03ae2
z710e2f0d6c2dbcd262edb0d526202706a07f41b0999d932c04d7a6ad23dd99c7457120c066025c
zdd87732f57b7ab536157a22303442fc4d2e62b7edab4ba479f09afc0b4c7b1a5a800830238b411
za1d449a458ecd9f14e658bc919f3db57c9d4f9a635b818d1f8cec5de408d361b338b659706920b
z5dfb712499f7ad147736ad027ea7b6f51eb5d8a915b8ddf29e292a8d39e1a2df7aba15aae0f926
ze075a312ed9c8b90339c91e75611f458138b33019394ec24528e3898d7d90543842cdb6b62ba83
z7a58c1dff1166334238eaee9976a0520340eb201ac44cd0e6096b36fd54bebc02de70c82ad1dc9
z8cb1f6ab7371e7eb5c57534b3ed92b00898908151f98adf6946cdd98d0bd683b93a5d4716d3279
za5ea559aebf0874b42965686e83b5dc44f968cd7bab750bbba84343542f161c4cdc8e48a77e2fd
z5c64bb742a8e7560f7d6f4c11441cf60b5dceb739d6b624d8c59245b21825a00c67811fbd2d47f
z38b4e7fa9985eb2efb78317a1cdd875b19c4021673eead91f45e0cec00ccd82a4fd32bce7abedc
zdc3decd483d4dc9b152fe36fe10f2a1c14f70e1095c5f58b533bb03689544ad106362990605fd5
zfb30021a07c0633824958d161f3028ac90d0009f269503e49a873502b8c71b8892d3da9946894a
z8bc0cfaeadb60a949d0d705e1e4b33ecd5c81e26da8f08ca8de930605d1f28709871983c64eb36
zbdb0edfd8f3b41fd34fd9cb892762cfbbec821d7ff70fe192a0003bbc90b8cefad3eff82684f14
z1c806baa91455f96f9486db9eef878a67e8cc2176e538d510606e051876cdc212b82f9792a0207
z0b0a619ed6066d623e26216bb1ca22f89ef480d46ab705f580b1a020015e5183088b50135e0f79
z840ebc6f88481ffc709bcd54723b2854eba4cd13ee922439cfd925c01016e6864d921bd70773e6
z0e7d9f68265bac10107bf7b7c7b2356d9fdf3de771b7450473e31b607d4dc36f7aa68ea64b7190
z9faac277b9ae7d7da00e79f986745848cc527af6dba2192ad42a40e5d12c7cab1747bb7cdad4a9
z8c08e9212eda1e3c3532082a2cd72e6cd6112fa9e539eeca18e48414987998951be1c7ec27c6da
z031f8dcebf998a3fc63690bf184d3017670cb72251e72e60f858e42ae5f29f3fd2d18f1fe96870
z92e6f84260ad71abee0cc414426e7e21f21dee68a4508db2ead7a55cde517391323cb9e25deb71
zaa97f2b825bb07c516b6814b278ef75497b3dd97eed52f8d6778b01d2bfedf1366501f3e78dc55
zf133860961b3d18c3c0340a8ce5cb9882790c4974e3fa4d025756f237d2a7e28422afcd567cb41
z03174ea5b7b591f6a1852a3247b6fca974376075975fd598f2bf68201d1b2eecaf32d328d663d8
z9f8a5096db851bf009ccf51c4cd88b3097067a14de6883535776b4d89fe65634436aff8bb8ee8d
za33c11e5edcb491871e3f9c348275dd5ef84470b7b23c9323edd53455539b600b403d6d94ea0ad
zf9ab23e037399e212071b70543e7a2b11090ce2b1e0567d7048f22833c7bba202b8b87aeabce9c
z1f9716de96044acd9ed55031b6c0c4ecc2a82844ac8756ffe12ed1605d3724e9ccc541cb281678
zd85ffc67c0006950bb3f070dd538abbd3806167db5fa575c0dc86c838415a477b21fca4745166a
zfee4971b278e645b3b3dfe37e208ab64771905bb99a6abaf418ce9472b5781083c6c7dc8b7bb39
ze40e527d897c28b2e8f280cbeee840821668753a9646b0304dd36c92a0206d076c825c75be8779
z426a0f71c76dc584f4ca5dd6e53763f87f0c79e704c639b6b4b14c381cc93103d0a6740657c19c
z511cca33bcf548fbd9448b0fb57464a8ea15d890fc0bb9b61459164cef524337dc9f1bd8ccef6b
z1d0f8e7805979e2b62325c1d30fc6d400b9acbe04beaff1a48bc44214ed7fe91cea545e2bdc5ab
z53aa4c63e4ca4b3d55c375e9f5fec4c5232fba23db6d2d378adc0e61f470d022f801c8784c9970
z1cbd5887ae24527032351bea85f90b1b52bbbaba236520250790f5b6f695e054c0cbce8c27667e
z1cc2774719799f002a6b42dddd1bb2f7a0964505a56abefddf6c005a4624018b77fe2275021ca5
z5a94bbd339c819ee32abb0a3dd5648876fe9b60e47361c126c3ba83755c5dd1864454bd8519285
zdeb37bf6a8092ea2528a6169cc528fcf523d28463a1ee39244f10ef62a6b159d08f9808f5781c5
zd0ed7e7f3920f6fad7d773a726e8f952ad7c781fb7681e77c2978cddd4d4fd034f68120639f74b
zb104a812f9cb459fcc2a1543c564d4312de9940b414b722f12a23f0692f8583514de45d041dc94
z73e3fbdaf347ffb5ab2d8515535fb0637bc39262c3fa4811eda6bdee580dfe255b45e22e82efe5
z2837962be9b16b540184df2bdb2d544de506baa146857abccf1f9afa866c93b276308f372e34d5
z7a9bb807ec006740bc1a45b365dde22b5fb9e53ec1a58209d4cdd8bd5cdf7b0e0993b88959ec6b
z3fcf34499239bdd0839d6dc33bd74177b82ca5078465aa1a0515c4845af7710964b87f6b304148
za9b7ee2a196cbedf2ef8a80518ed1d6b163c52bdd3c5b208ff1a95f8a35e6485e315df1e0bf7c9
zbcb556905be9397fdb63ee9205c2f2866f520517af25f1c0f98bdfaeee40f37b9fe2bfd3975aae
z358d32cefd57e3fcc2371cebf652f9e7be8c6a021a558530d0c21ff20916ddb01c89d0c5613350
z5a7130a8b5cbae45bfcd869a362b11fda9f10fbddce8eed1074fad8b0f47c5feffa9f63189f2bb
z63bbb26d886bfa09d3eb29d0f96ff78d8699187eb18b06c6ffe5180ca825304f05c9681260e078
z413e074800c550c9e5af625de2d83b6c346596d5c5eb5a70a4d31084b4c1d3ecdb287c44909071
z36b28989231f80f3309e4d0eb64f271db92a3fa962b1cfe9a098d8ede8d8f0a8c33a0eecbbb254
zc5298f44a829602d5e8cb66c1a806d5468d433d8904342fe89ce9ee4d2884d2b60e680eb457ae9
zbaa6f5d0de61801e7392072fd3fccd1296f87fc7317101db33071f45a569b74c3845f4d7abc566
zbe8bb979ea5005077522e04856194aa69107860b94f1603c46ed41cc71cc84196f29869975573d
z1df08964395a34fec9b4f06c3f29419c4c0ed5b0513309c7d573cb5f57d8d96deaf830fb72cc15
z19516241c85b6279b8383f1bf36cc5768cec7d48c893d22362fca39d0f93a04760d0cc46842a68
z722fd327c396f794474974718650f8fc60c595e5164fff35b7bbf6d432187763c7413a6eafb281
z87700ab30c25dfcc4974bd486f113b0d045713a2036acf80accf036b15018abe48f40be0b51b7f
z9fa8caeff08db313c6577af89e4e91743787cdd1ad28456ebe5ecccc2b9006a58c34f345dfeaef
zf6a113f321cbf7d2ccc0e9d7532a8cd344cbae3bf0d309e16b64b749a162d1b616d029bc0d348e
z6407202f6cac645b35455d5ed70da356b7dbc6d91c35792243c2df94d19fb2b03d7f56900cab52
z180a0dd9fed14edbd069fb65f2749f84fdefa2c7e6ff4d1e37369abd3b1201a677305c2a4ba4ec
z93c8bd33d2c2b1dd47b9c871a4a1e494e7db0cd82bac2444b69a07b61ce22a40e90abf3a4d033b
zd8882a27ee5280e561d4387cf89556f82aec1695ffed0563ed9e6b5397568d2c741a2f555bbefa
zcf705ef3241d431a6c9ef6db8068daa814c3c742984297faa6cf6f3f953a68f7c684bcd4e556c8
z901519d6ede4bede715afbc0df0d5fda9b6286b6ed6b4d5b5ae85bad47fbe8a053fbf22b5c6f45
z0c277c2f0e77f81681fdbf676ebd4248e5f2b0ae546f0f1d8d2ca815dc382b728b893b813e5389
z967bff13c76aed9457b4012be34425510f1b6b322bd46ee7ae321ddc557f75e483cb403b0e2805
zdad36020d19db5b36a6c48dca72541410238b3f00077b0b311ad7ac2e05acbb9d9e66efd1a7412
z2dc624f36b904088a85a3c7f830b7845b2807972ab9b1f4f22d66ec0c4841f4eae3b80f4d4dd5b
z18f1e4433b75a87c174ee5b2fe927c48638928f38a07b93e94e0756dedf081fa40a13033069b7b
zb4a7a8380fad16fcfc439e8e4da5cb8f6c77c4a548e82e148ee55e09b77f4561dd270814018cdd
z97ea5278490562d686bcdba38a9c88ebc82bbb4fd3b498c21dc7dafd281ea1de779ea1743b5704
zb44dd4fc2e841ab9d2b6385c61355be0e541af7bb8fdffce656e5ca01794f41b3c08e082e4920d
z17f8f783d8c82b37d79c8c27d4bc494df7a199e529c7915ea3f04f0b8f38304d685c355c3a998c
ze298eba16d46c043430a9e3db42b886e68d6d60d812c86d3727f3823f22c510d6ed088b60311db
zeb8ce5aaf8d09d3846ede775009c016284a01bbab4454c8d7f6c356d7958f14422b3180c9bcf83
z700d49f444e4ea13900fdb0bf58c12af13f95a09d5772b149b746f93b79573b7b006fb0786b914
z70b208f7069dc3689f8682721d5767244df0f45bc1038af811edb7323c88327bd8c5620c6f7868
zae1a0fe66107b1f2e01115213cc74fc5b1148dc210c7eea0fce44b3acb216ff58da6114157249d
z6426e4874d93c243f7994399bdd3392a4135e8c756efaf8d13eb2990be5c7de7127fdf243be2ee
z9ab6c751a26ee5123e6723314051588a5572f96b9c482f3ded31c59c07ff0af7734475bb06d55d
z99461054042bdcb6bcf342edd741328a3275fc5e7d4feeb8b5a1f27962a3269ee324bd89857cf5
z6e96091e8c3234120d116b4fdab0413c34834b16f65fa84fc119f63937b1a9d44c9c8fdff431b8
z0f43e4f491a833a7ecdc965fc01cb0eb073ba1a0b9e1de58f2c4bb12632d40e95cb597125464de
z8c71d077261ba74a34bfb8d68191360c2b98ada7b11be9257bf960360161bec32da8c6ca3acba1
ze38b694eccefd102375b1aeea9af80e92d5307b277d29b0bf7d9e6e39c7118f3a85e3527b8e6e8
z9029f52c7bd85c943a9a42eef743530f3da1176fb45bd953c36932d0007485f19fb0836585f162
zf34e0f909dbf7ca810e8f230275e268ccb86f7033148558878f24f06bfb88b4ef7f817f465e7c0
z12ece4630e4070f403eaeba6778036f871b05b50760e83324cd9bafb43562d6b5795f4689f86b2
z9c1b75284cb54c01a00dd4f5fe3a6447d9c234e370e2b078465a95a17398066c1cb89a507be33a
z4969c36e2ac912b071ec54c7524fe0ff13ee4678891840f9d522a5d36b7471f8f84b4a3aebdae7
z09cfb38fd27bc7a1adf6289c9773c10e68a211ed4af282b797ec952042f34144b33f0923576fad
z5cb08b1c81121f9282d0746883685f50b29817889529a097b78c4d162462c2d0aa2550ab5aca8d
z684c355450ced66bcb209e0cc2cd1b11ad9e009967fedb077f57f90f9783a9cb74cd9d4668a22c
z39b639c18dcbd08e70acf82fc3df6f2fc54f857296924aafc5b49340dae293025f461b65c8c196
z7784813f9d81f692285554f582b5d4f0e165acc6d1b86e60db8fc818b24e91b8b86ef644402b37
z44a2aa66f5456004df93eed191efbc31ebd7d9ff6eccdeba2b32ad8a18d18393285ccf8998e1fe
zfd2e28400681361ade8c2b915beda70b17900c2b989eac11a874ec09fb8fd2e1dc167e77b88376
z5eecee8470b2db35f89aa9255f130548c99d878e703a675a066d8ac3501262552e79132d5691f9
z0b90df2f3db7664e52835bb011e71dd1d0ee493e07639fa58021eb5bde33bcd736a17312588709
z503224bd751c06e73fed4286fa0929b2c8c68dd3b22c096b0ab893e848918b3c3c1fa8a32f9610
z4309e904ec9be476c9e0b9fad1dbb1786cc25bd418374edf48191993eb8189a08aa7859402a489
z9d6835cda6cfc857b8b3031be8c11a2c7cf5b0fa591765638e52e776622d51935176821586e1b2
zcd2e6a749fd39f1db851219a2b4256073dc5d9a1f3e076d4558f34f79234eee33c50699b9472b1
zf6492200b944afa96983d74901eaeee15de254730ae55eb42826944a0a5c8cb69bfe4ad9b742d6
zc6a4a484a63803c6f44813f45f29f507478f1442473504a218967cd5653ee6b89d3ac7ed773851
z17a00214f5920476601be9a15edc22bdee8be8008c9f335786f6bc09bfdcbaf53410c244e1509d
z06aa0c54fe735e01d49b477cde1c46fc595e33a17bd39018b1c1dabcebede99f5fc0e11e354f51
za045e758b708f5dc6b160eff94db7368f129e9143d9c2119d12fa264097edf32ff95afea4cab37
z8b48f250cbf3c2868a6cc07e52d11572017d118104b6b8e2a23cca9003a3030b36b686089556fa
ze36c9e0ab0a997b39a0388c1c6931a5bbc0079b45c13fa1d89d0b1b507dcd86690fa7bd3a038eb
zece726a50e049edce05091646c5f619278077d7cca41ddddc092fc04818da2dd7eeda35f0a1d48
z5c3c2986e9b0b2f248a64bb595f9399c57cea3e7ab1b33f66c3c6dd105cb04e4314ee2f32fbd49
z0d9c89f9e5316b1ea01363250c9c537ab6e3bb78305a95819c00538f552215206b035e72e2b7e3
zf30e654a90cc882f900ecea0305f9902e1165e859d3a704f72a6d9ffc60a5413cde5bee7ed8c3e
zbc88448aaca608a46465c5659b8d39af602fe201246bb45af14db3fe1f6413b787a00c93f9d879
zbdc4431489cc622b7b09d25356f61f3581f13cbefe776d043896345c77636ea6f7804aebaa42f3
z85fcaab032d9e12460c5a208b41fc35f39932ff1d1c184444733095246bcdb568831727987fbb2
zb61b0d43300e9ab64cbaf5cc4172666b65101a569504a69ae21d68344df21c2076aa65f67e7e0f
z4bcc8705fbc561a57f570eb39c4560b18697576d7c876930392f2478dea3d0876602d1636d2efd
zeb1be3c13db0a430ff4686649c0b6710895c835752a8d0f51d3f3fd4950d25db54b67e27212d81
z984d1fb0f46d4cb46a378d1bd22b1d80e6b732ab2a9bd0f4130ec28bced61bd16248d549d1faf9
zcf1fdcde75d0a95f95fdb7a6d354a01359295b97cd9672d11ddb2ad90fec3b0df4254361a085f4
za231bc0e75877fa2f6058ba0f2f75e3254692ee322299fa9565a9a3d1cee0c9082890ff7f5aa1a
z992546a11c8944a695eb2264b6ed91bb8830f49e18db5f623164ba59e7b5bdaa12428580605093
zfdec05c1e1a88411771037d1b72da26eb20f1ed0b0ca0310c7ff9f1c439256d082b1d6091a796b
z64815d88fb2872b30d7a6cfcbd7f3b7174f5661e7fdac84a514cdb9d58a768a678a3ef882f0160
z0c13c60521808864023666e6e98b858ee51a41394312bcbfe107ad817dc0e8ec98aecce7b7aea7
za9ac2a9820d0bd18480c1fc4a76d1e738e1cde918a35b1457a4b4f7be6770f5863fd0d7a377939
z4c23b132f4281442cf8022b994e111172d8a6294d809e487d6b2186e89623a6d048c0404c249cd
z367b2534ec3ed5cd59c96874d3cd47dd9b8b728212d6dc2b119c20b1cd50a005608fd31faadce4
zafef8df232e519f83f8a33c5bf8368326c3e9c72dc914312b5d4544020725938ce79c5c053293c
zad0625755960b21c67cd14df1842397ede1109e7c61b197683cab9d712c8393991c080067e4864
z64634ac64b023411f27f272d9d7dd7a6ba94148f2c2e7c4921178f3caf919ce5ebfeb1a1216f26
zff59735e5543949e1d0513ec640feae213a271c9d11145ff0f5f782ce4d5087a213db8c11d3c5f
z345d4599cf245ea4779f26b8d019908868ad903a576ae51bf48e73a11e24b1368fe423754a22a8
zb725b37c38a58d28ae885831af396c3ea3250335c4ef16fe2699a59a694657b7a551dddafa14e9
z6ed2d062352dd7e58fec4195a4fbf980532718940c7071baee0b3634d9202f886997869ce4e04a
z34e89d07d56381c0fec4d2648502ac9a4ab99dae028ab0e4ee894380ed23137c0fdbaf895041f0
z970532c6b453b90eb0b53294440ace26f01c15743d99a3299ac6a9509b3b3f124c9fb22d8e6e74
z70a7f19f0de1585b3407c29ec92a41c14fc4b0f12ccf6b0cabe15bf5a4999e914fbed4ce70bf73
zf7699d65ad41638e22c2356d532e308390fb94af1ebeca839c9375c5a65f9d90911152ee6d4f18
za2fcfce003484679ca8e04be9f83c50d6293574a29b4e15db63d7a7d093aae24d1910906b1dd7f
z7cdf4cf1c18f0c5b7815569355cf66ee0ad79d8a3005684a5220baa6d8742dc88c2bc86cdcd93c
z25f5f26581b54aae327f7601e6e138b0f262f8dcdab40d6d243bdd9335b3e5b5635a7d985c9335
za988cfe5384e65e854cd049d79fa7bde581a3d0b7739c2f9b87dd230337d586d30ae15fdc108b9
zeefc799dbb23852b009558cde0654b84e86e308c2a18c791c5bf9a133ea87d32196a40bab13ca3
z073325738a6a964629a09e8e9a395c25b4c65352733e3ad156c0400e6f398c25507cfa4f7cd577
z40eb660b789e1f90d99d127f683f1cf241eafe222f699e80e45a88be6e3bd77fa2dc931cde9dcd
z43b274693f2545c1f30cefd5059f704de79d2e85cd36f8e62535a8ec2f643cb51818c8a7e1fbaa
z51663afd6c884f132319a84b13dda9ffab2563ca749a075e2ef1fd8dba8cc3ce042d6d91652525
zace122ee61791be56288f06923da0bcf56a48548f24db0125b698a25616035f70d3c7ac86c2bd3
z84ad56c84677255fe59d39ea08900720ffde33bbaf060b21a7ff086bd8d779bf50b19d39f56127
z80d16e1ba62136251182ba5852600d37c76eb824e1a415d79bb33c35cd431faba81ed573d46817
z82e127750a87c4890248fbd6a742f1ab5d5e2ef13932bef35bfd1221d6fd23b4728666eab2ba0f
z5c1ccc99806bbecb44b71563bcb5a5fd89c4fecedb930624500f6b609e5e344aeb78fd4054f9c0
z344267338e887dd8350fefeb829868acab2678d10b03945c466468186f526ef6c50832f58f0384
z796babee82b9a000dbf60cb9c2b05abbeeec13775e36de527fc3b26d376f8df4ade4a00c0fed15
zd33cf21011f428cc54ac656812756f2af96e53d2ba617c444ee0f4a330b0f3ce6133af1985e401
z4e7c1321e4b425db7ff51c019a721e77574a16b8743b0fdc4085dda635c33c28f1cf47cf02a1e4
ze8db1bf0b16ba05f09d240f9bb50c4c70dd0aa5476b24c5561ce4ebdc287392a913e5b7c683dd8
zebb2549843ca03f1b19e5cef266a67cafe05b72d518397e429e50dd0adc4f3331cdfc50fb7fca2
z73e198a2507d8c1c01fd76111244ad524750a1421188b8ef9a30ca17484302c3117341890a96c3
z160aaf89daa2b425bf6a91b8a19dd0275b5efb4c39c497b53b1b58147aa7524f05dec920e565a5
z03ce65208a0325c94bbc9ead00429380c801b7da77ce7192f7829127375f831e79eae79b07f556
z086bd921fe74adb2051831c1f2357fbb7f24b261460e61b5b42d3ab7a6f7a696d3c8233d526212
z84f43ffc234c0c3eb8e9cd9c62c254ad3d86e8227bdd30979086ff009e46f2c9b14fa141c83893
z8fddab672a54854e7aca0304d8aec53d2510c5140a5d942104fbb4a30b647e09ac0ee72669baac
zd61584e222250d88a9d9a485c3eb9392e67c071187e65ff84b0602af7f353ab7413da144aee155
zc4ae60d4a82ee6519248a8ac0e83a8a078789513a6b35c6260a327e8f95ab5dd206e686bb0c69c
z429f41b96d6b0309a0ad114d0a2e22509c676c08ca0bb9837f9ebab6640e604fa3d5ceb38103c1
zab7266b7f038bb706ca70a871708fa5d1e266ca4fef7877a9549e9b8911e1e46c3d58117392627
z3dad1ffc7613a4558b18587d7004c649b6085043ce881297f7909a1aea313767a5d36c73343e04
z8ac50cb163c769a2e195e5a774c339f2d3116d63904e084a7b45b8b7bc897d18151ba2274db40b
zf439e0f601fd7a07ab080568bf1de13eff31e22c909fbf4af33b88d62eca4b4a89cd345729645e
zb088ef9f13866c2dba859e672238af5c261031dbe453e96f31c49f922c394ca96f5c100f89c36d
ze2a962b24febe784e6293cd3c2e28ae13f6b0112ad03bf77932b7ab3b64a113f83d8425d7eb3e6
zc21633f32ef34b2d2ad23625566814fd4a1464b0e0fcea68aeaaa03df282faf0abcc20f9e993a4
zac45e15c60841bf581f448de74c8fcbb99fe4902113bb62dc41db59aa9f427ec0535f00ec31f97
z14f23586603d1b542a785c317eff542ae1ae7bfda420941fe1034b55e3d08f63ebe083eba0f228
zf5dc36762f4d2ca0548431d77c12b75287b4f4f9fcccf4b3d3b1b15904b3b3c255327d2a1b8c4c
z7863eae99708f48227d51b31aa699ea99de6395df02fde9a2841f99c2c833d78d7a9b3310c7f8e
zb60868842dc6d64f3603d796f6ffad4631164e219120b6006a67bf086d09b4992b914307b9d7c2
z00fd90b69befce33d94b7343db735fe78af4b62be338bb186c88d71e48d068956e5aa4548d5b85
za009a93c460a9bf28bfb6640f767bb5cc58609d89a3a0f5342d512ba4dbede2bc252daeb589232
ze799d544bfb55fdb548de7a745f2a12142525f076b5fa89f1acf74c375d337e5a4cd9cd92dbcd7
ze8e87f194c1995f6c83ffb496796bd47b91a3a27dcdec519508493b8ce135436423c6c6944a6ef
z16cf681498bcc575ef3daa84c49568d117b5183cb374df2c8c1e84fb1ca8f80bebaafe8f06d64f
zcd60c60a1e79d6e5a88a3625be0906c46dc49c9bc7ce58fa0c632fd55afec613537022c654d9c7
z383de7a61794bf23d16df591eb3bdb9d67cb0a1ba56c78d4d8e0c44ba24c59e5726129c1964a09
z2dea6257f028ee5c87c17e7e691c3d59d08770049aabd1d7dc160e3e80957151f606821420c3e0
zd5bba3a56aaa9d4ba5c2aceb0c3ef213c7be86a2d62650250f1fa773e78b854b1f407c17ea2b56
z1cecec9e93326aee0b9883d268c5cc9eadb4e54a5836998b06a7d843f8c659b948cd6a380a8978
ze739c1dd0cc81be59833e7531ab65733acc1910fb61fbc15f9ff47d0077fcacfdc71787fe36755
z64ef5b023e93132a06deba9dfd1883e08b6c2f9fcc0bbf525c2d580719149bf17fa57e71448777
z187a3128a5a09206d7b4e289d2323dd4db56c4468144775bae6961369c2819c166d85d0a327479
z7e1856bfd810d3b66a9b712e3eddd4b7d6a79d44a9dbe7c7d50b78e65b2e4119a2d5975a8c8f6b
zc8ad7ef3cf2e224cffcfd935835a2fe53a0f9889cfc52bb5c3ba3fe6c5547471ae62aa1dbf9bb3
zc1615ec0211a523c8502a5ffe51a8102e411a5e8d089a987ff14d10f501f704aa875cc91f303e6
z7b840bcbdfd77ef8a47fabe0a5bf6ba2cff05746f6b995b7bdb0fadec44047a33f805bdbce07d5
zc7880de6b0d3ca4123287c236548ce12a018c14eb02ace6a04c62c07b9425af0c5f4086190efb2
zec019f5f1a598e6e782b646c98e882fc6374eb56036afbf6a0ab8df98810bd470253d12161cc1c
ze36f13fcb943911709f27a5296136ea973251e14276379af79238df81a40d74429259e8df94d2e
z3aec5d55309a1a34c6f1ea144df29c623c793153c1834ed73618df0694f99203d0e1365ce0fb31
z50876155670f39b3480a467c0913498e1197c95e9c89e5af45b01a945f1e3b100a8d9daaee167a
ze9033f95baca26e94320425cf2c0399a5ee798dac58da893913e259834e03f36c7ab5f80a86725
z26f8ab04c95f60c14a9c8894c344ecc09b8d32fa4a63e8a4afcf549b206aa23d98cbe69d2ff7ad
z258dc320e671cb1170a1ac6dee194d12a1b3a1fbe430d48289a68c95410dfb2b1ff03d4170b040
z1bf2210567438f85ae178e219a2ceaf0a2afda93c31d9f5d908a500687de913447dfccac316b95
zac5cf64abdbc5fd102bf0369f7f1800dc8bdac9d2306ec67d4e5315718030362b09e99d150738b
z77e2999595303543016416c0f99eb7fe582d4b6670ec6da26151413539827f489f3e6eb9bc483c
z593fcdb6ba3073f4b47b540fdfd675ef87fa5953d039b61577c2b3c0d9f55ec5cb30f465fff6f2
z1582bbf178286aaf1607fea2ea300681e1b3170cfae9698dc4ac753c213c9cbb2785d4e332b8f3
z12c40af6f42b64f0ff09ca15f950a8f55163f7fc38c004ce08b8c82941243463bd4366063dafac
zd2593e869d2b1c44fa4c567361303fad075f98829df8fe535123e6fbb37e60ed5e317875f57cc8
z6423d27bdf0991e1baae7bf955707e4a78f650427efe66850706901511cbd7ebc2ad344f056b7c
zc6ea0064fedd6b8370e79bf906a05cc7a5627149f2b1a97cd85fb86b2652f4cf090661f76dbb39
zc3561fa78663834d07a9af8300a0d4ee4b4eb8560da794216e17e9492fd0ffd2f22e981275711a
z144c3b1604a46c1654c8b1fb11ff62a576997109eeb45fe89037295bae547a49753e7f4099c57b
z1ff888cb203bedd32106f4611c23e67917b25cec5619387f331fb38292f73e17c416456b3a1002
z191d1207d9d8967a1a79d7a7370bdfd7135b3510c1f90fbea2d820faeccb704a18f821783530b4
zd7423689faaf5f62184250594d094af99969e9515d904a381c8c08f9d2f91bbd678c5a1c9d39bb
z3952ec00e195136b8d9a9c2346a188b88a64a163d97671e1072511c64853967542ddcb1b556aef
z812fb1c336f85f02ed0e040ee51f7447618148ae6d2cdc4f58ce184f13c0d7ae8f7657ad68218d
z7325b044f0cabf19bfc8b1e019adeb0e7fd648ee32fb3c1d21159ababc9e3c81202bc028ff463b
z6690eb043c6c1f521e2d152d54431113d9c32409d8a55d3e5ad2f829e358063b7fc12b21a03a19
z4e55b5055fde9d9c7c1e434a4def4418a944285c5be7de8e510a1a0c9963ebf7b7b57937f5c73a
z8f37d83825e4189cf4e8ca493a492702578cd3a51c26004a07509d88b182c95b0b273c69e584c3
zbb214ae01faaccaa33c483886c5274527d1fa77843efa120486d66eb628b2b48df315beb99deb2
zc5bbb53c675e3e7eaf45a74c2b6cd47b47081a79d8d11e78b064748837cdbe654babecc255d0a5
z22a93f1b8811c8de97551ed1ec4a499740abd1bd4692955dd7a84b89b017f569524226779dd401
z40373742acc93fa2feca0b3002f7aa14eaca4e493cf1486eee9f355e768b14bf4d0b7885efd475
z610e758e24cfc8be95a5e9c3c28e157672fb64c42d7f1920ad702e02c2937110249eb0530426b8
ze9cb3e810de6202e91f50468c3a61185826ca18a6e7f46fd43e86e156b5724d99d3cc8ad165f18
z758d7ed6aebab83b2755622c25182598aff21e09a6f27856a38877cc9cfc404bb4ce6d823f2b65
z75fe5a25dce9b7c3a0b914156d5f574386fffcac9ed7ff66a1b419fd73f392c2fe17672a7e4440
z201481ade145f0beac2b7023c9ee40cff32182c5fe05e7568a26e39efe1863cab9164f1898a166
ze6ed6321a42d04a44bbb68d9942fdab6b4ddeeabab1767641fcad74a53aa330f0e03a4e8471b14
z84d73572b695a6281afc08ad105b94a4fe5763810c383d1da14a9bc51035e87a627106d9d17cf0
z26ebe056edaafdf56638b83988d0b79972eb67c0bda037272d9abba42a6fed54db6608c902e8e5
z8acbfd28838f2ecb6da636421bccd57e9044fceb10e59ed47340d237b5c5dd935cab5511828e5c
za819cbdf437f73acadd56ac1962cb49c6598c07010549450fe093d55dc4a9e06b3abce5cc3c08f
z634c325a6127d38bf84dc1cd0989f9d29195a1b533bc45155edf526b3e5ee69c0c8f097d4f7899
zdf3451a8743c583186390f629a6a50f5d03d5aa4baa89251ddb9bd6bd2a4f6c7700b9a91825e87
ze7860ba8444a22ac21d13391b3949dc9f953419a315e808e5e2a72e3ff81bb21470fca46c6bb6d
z800bb42fab4aa40a4df9b4df0791ecb883e1e8f9591b4a8dff02143ab06416781292dacd93c837
z68eb5788586e886c5462dffb1a84d2097a1781690000c07b5e01d616398755407d54abeac53fd4
z2a5c510a40a7066ec6a8585a45ff9b77d4f086a883ba0444a37a644c834914d582929052b31210
z1d8d83d8b37d1e216e7c0663fa48ab9530c42f571c8f1cc2a8fe689296d8dcc9872cebd8fbd623
z77b7d2274a3cc1101ca96e73f4f00982caa28ed0addd80bd040de813c99d44e798416050553324
z3676117c7d8a9aecbce2b6ef6ce74b620df4cc43102d765f5eb037800fa6ced0a6fa9b95eff93c
zf6f793ddcb4ee1c7f739b7edd04dc68c786890be13692365f33728b3c60766864d77083a2df277
zb0bb7234a861a47f6f00a8e6f91f266ef43fc7b6aec3406f9467724642720e30c6260bd2280003
za629624c81fcb4d212b57ad7381172ec99c3f80c4308f591493198bb4437206a7b2e64ca142d39
z1383109512edf23b5d7442dc0d735a1b080467cb2068e5f501b6b9ea2f52c52f139dbc31cedcd9
z5670ccf7f4dbd9566848ed87a9000e83e117be8645e1ba0f71848dd160800304d477f652c9bada
zafce9cab3ab83a6ea97bf22c0f57360d1c708cbdc6fd45145ac2376f5201e20ddcd9cde202aa49
z990ba69c72d22576a387805785bd1b4213c520a46db1cb1cfdf1700ea34c842aecf255a2c3247d
z85b6c5ee555832b58aefa35151ead69427007bdfc6a484d5f3e641795a5f4806afd8b1587cffbe
z5dbe7bd09baf6dd4e7a0ba49acdc8d6d30a8030a33a01ad642f0c64da9add5f340b195d3b0d131
z9dd3cfea0ec95f3db1daea8fb98f1e917deddaee4458bfbec1fbdae0dddacb03a7731c554bd3ae
z2fa40c0d265a0520f7e901561d7e0ec456ba3656d11fd2fa3fc2c2d61ef4dd6a51f5b39235b69c
zf83ea2dbb4fc8d32072ac8f59c867ac861f085fa8bbd54a86a1461ead4fe50035ae3f638143743
za5c9e688c274a518b410c30693fd6273328b32ab24f7eaa8bb52ad55f20e810f2e861b711d1545
z436247f4305cbeb8d2604c93ca59e0d84d7de9f000e64ca0739986fbd1beef955eed94825cd0ba
zf22d0a7aa84a77d3cd60622b684d936faeb56912dee3d74565c6aca4f7b444b5660ca658043fd9
zee17783f7792a9914f83d0113be294dedccf3979e32398bb6aacf8cc99ee775f0d85cfc84d1b15
z2670dc6908383c866875e3848318dc182621b8a403333995bf35cffb8d3d091bbb07643bf880b7
zb1dad1115d992f82668af52a88bf423461f0dd3e66edc1d81b6b5e6058b18d20623764445c385b
z71e753ded3322c388223932a13b736a7ebbc735b227ae34221999978557c3d446a6f3243b014f9
z8ff695a5f56afcfb4dfb689ada8cfea88fec1c49fcfb528bc91ee2386435d1efe8dbfc8782cddd
z1aff269c780a4e38b9d0644ce54750068bc6d5d7d6c071b30177116f22629e5693608753021a58
zb63066ea8c7bca64f8566946ddc8e8b4db8a71447cda89890ac2c8e667de8b0e82bc6235957a79
za9e7087826fc80b2b7c499b51c8e05abf7aa1f6f7b522b1336e9657d5c12fa27409470a3223f3e
zed17e227547b166ee57a102f4c6af2bdf50495c64920299adc5fa4594fab089fb7e5696ba236f4
z9af3c6cae4b1df3a0b057a5eeb0e8421716db92aaafb7cfff63971164a7611598ccafcbba322c7
z5ba121e29d67334bd6131e75a3880798c4e68d938a9b80eadfaf7e94b14f86b8d8dd7f8c31f422
zb0e0e1298fab04020b038737dcd3f49824aaf016943a7b6d46604004541e34d02ec1161ee355fe
zc3a9b848290ee607a1c1fc33f1a5463877269c0aba826163fc981547e6a667b5af864a8ac46457
z61a68bee70d4d824dd2033d845ad44a6a670817d0513993de3c03ccaf8f255d805facd94cc113b
z36f136e2b818056de740800c74311d4107a8a282b712aaa450785685ba93ab88f9b40387f08c17
z88057ce29e28e02f64f87ba8077b7a604e9ff948a094ff68d43155c0e32e29457dbdf030f0bd11
z25becbd8fad2434ab8fbe11640352604ae70858372b3febff83a3d0a06394fc5d8ae8d6293c301
ze2c2f5b582c8c762029f8f30c9c63f2db87ad0c53b1f2ededdff909212bab4656b3c201575fadd
z5f50cd63d59cad246287334fab053414ed33375f06166287ec38bc1397e657ed9ccbd66382d1f6
zc297f0dfd10a210fc1ea7d26134cab8ec4b9c917008e501148e90da4c154fe236180749d36339e
z0fab43afdc191897ce92ce4c4df98ebf20d187346fb66d24ee9d02cb83e631751727e0d33caad7
z03259e60ac16b3b8f5be6bc602277c85d48d5e7b0679145044f72f3b68245b9d11fa6eca3c8177
zf6ccc56b73f24e2b9d0bfec9cebd4f18737b4d9a8d793e8d4abd7e661f6e1daf671f1262697333
z7fe14ed4daa78916a4fa9572437f854ed6d3c617a607995503740a8d7a10f3a8856367e7cfd313
zc5d9f3be02cef891ca37ca8d7138a1a48295fdb5e6b88c13a5132e7b5d94f9779ac8a065983743
z6d33ea59d25924316ceda8bc94e705c01e4ccb1faab393b9002fdcaa535aff9ef252a6036ae231
zf27f0e076068ded96976c1c166d20350699804a07e453ff4225405ea150e400305d3a54143b756
z3f49c349f55da81aeda716bdbefe9e0174e75b6f6d440a992561a1e896796d4505bce2b9ba82ad
z41a538adf6582af0d2e02ae99dd9a346f61e1c8c5f85e0dc2da4391c4b389d3fe8e729942568b9
z72855477616ced49eeabbf4253ee573900e51fe4baa6663e9c74164c86cad80d3b96c9e5b9f1ce
z3c5c71350d8ba3644221ba12cd17c01d71832bc56d26e4e29a523c58c95262a11b3daea269ce18
za7fe9fc64fa2fca3abf551f4d5b955126dc0fe0563f585923fc33214af9fc371adfaea6e9d1c33
z8ad64ed71c5236292f72a42f9c40a614b510285f5aa230f6290ef2ae68cecd924040c0c2e1ea7a
z5208cdaf55e3b78c3a0ff599a350c6fef9beb9e29154d39ce48f4524ffda6415bdcb9f7086a8c2
zbf2feed073ad2747fb28e4149314d551a42831387cd67e88be4be9006ee6f55e70ad89dc2b36b3
z7d41e69571d03bc63599f3f72c0f0aa6f8e038ab14fc90e08219c8df8ba43d949bd2b5c225ca89
z86cc25c62927c28806019ae464189895012bd9ecd31284490a0805d7c59cfb11481692649d5416
z73c54c23543729fb14897d888cc1e0272d7337eced65e0664bb633778f6ac5977a7a9e02e2abcc
z433e983ef05da368877ab96ce994d7bc6f2bc50a241afd2b3399f3a28d143db2f2cb75aa581420
z0a9482cd986b4ac40649278579f72da5d09eac5c2d1b0c38b8bfc0a45bf22bc72018905751349e
zace711dbe91ce57f8784617e4e5a65897cd37d78e94c9b43f48d2673b4f5c3957acf488d8b687d
zb311ef749196e771753ae3eeb1d324daf452361b7f0e40f5a79aaf3de2ceb03cc15135c030ef86
z0ac39794969eb62a8dd821addd4a9c100a1eb60db9bb350216ed1d394e71d712efd265fdfcd807
z4aba0c769ab41b6bce8373cad5c4a1e91a8d479214ca83827ccbe230723990c40b74f4e678c8c8
z57872702778ec3f25218837d3210f78f118d0936083e6818d6747ce2c0e8a7e6f6dbffd1138ce3
z0a4410db784cd0ac91344d38839858b951f86b24e7bc8b5ac6955b1b852ce8c6bfe004e21d6912
zd18e2b8a4da972f6e41679a9f6a57bb51c5a0a851535aa8c8e2836dfe14caafc59afbc8787a653
zb5d420f8c3e631ecfa79ff7b10da3c7206a8e44df79193d402d3f6223863296fa230f49885e3d3
z40d1a2470cb25441fb0a823c76573b17d00b1cb4a1ccda89736d3cb04850e5cc0f2d653eb194be
z30167942ccb2644071e808f138e1489f50a967e794a7e3ead72e8d83b33c96ef60a3c54256d89b
z4705bdc8c94c5e2ffdcfb49b5b45b17e48a8eb34049fe4e9a6fe1037bb60e04c2947994d0d41b0
zec391629b0a6493674dce352c812851cd881001f4366131764ee24b2ed72cf1a80f98e79a82128
z51f35b351ea936e18312bf9d01863d5c887df224a1e4803d86285e43ffa3746030ed6a026881df
z260b7abaec0eb810f47c207d18f164ad85d338bcea2e270e940da5fbd9025b965a707ae7b6f789
z62814268674660d5d4f4367b395380a2d3c538dcb6396f2de641e7d141e0e3fe46d648c88366da
zf2cc256cca3d07514a644dd1e3089066de544b8ee11dbedb050a82fd4f8001a00d13a68d3a8f4c
zd3168fca8d942727c864d4abb26f7fb3f57b9e804c4374f24b48239a0579e536c940c626d5e212
zd4bcb2066eed26155d29655651c9a17535bb58da2ffafd61dd349bee58484aed97955c1aa98242
za0795621dfd26e7ba0505562eae20de1914d93334b7b966fdf335346fc0fb6586ddd16412bbb9a
z5c8307e1c6de2012ee3a9384a332f13e8840acc54f47fb45136a0b672dfa579ff7874c34ec7b1c
z8c596bea6792e57155fef96aa503dd08adeb7ceae049ed40d66b3a7a035729b9f25ba9cac1e134
zd779141dea2fdcf0931890f42109533e1121be065dc7c86d1ed184affedb0dc61916ee9115ac7b
zae3e054c622bb0f0358e1b9117d9a25444b024b8e830a2da50d2dc8d1d18369d39cfd850f95455
z82a2966470cf2338dbbddc74e8229e5b2aa006641ee7a5fd44a8eba433fe3ce8a00aa4a1e816ec
z05778cbd7a546c84c044f8032ad845c38c3b25ac8fe26432d856437966693116d212ca3c540ae9
z80d17170395ef3389fc55f9a3fc7d688b500308f421b2f073917ccea730a6eff9f31d9c757bf2d
zcc954399363287ff9a55b2bfc9306dd3a4ef902089d2b2f47e9defe5dd1b39171c450a36c80101
z027432669a86ddae007e55d3e476857256e4834a48116e71e36eaa10215f460e2032a7de4cb4a3
z28044fe63a0afebcae433bbfc11740a49746af91183e8ad182e8115b9a858259a52e8640f76832
zf28d87e7f39710e39f54e6ed45ae6ab329835ab8e7c22a9ecd96a83c60773be1d2e4c57b8ef350
z3a3dfad178ed65ce60074e454e28b6d68d2417cffa84c179505410c2580b6ab28a332c5035bc74
z85084f6888fac5858995e1b7925de842a23cfe6e4fb3f09b3136fa591eb00452e7672e66252ef9
zfa84cef451f708c7ce2f6ea07a320305babdcc15f5f511510d175ce5b0160cc27077a1f35236e5
z77b683bf696e52f5fb0fca3b4cb17dd1777eb21f3d201803d9145bcedf3b49fd8c51eeffd8b115
z5512c66ecdb2e6f505978b3394c2d1a22a7e9556d3fde0b88bc5cfc6b44c5c2501dd648091358c
zeb11ecd2c0256fb554eaaed363eb9507db120bf10726f286c72f5198c8eea04114f5808c9f8927
zbbbd4e17866784aece02f11d3bf79f0bc4943dbf6f52d92225c4e5923f5a3068fb7b0f5eae9670
z132c0d5f2fbe18909e0c3aefa38e701b4b1c465db9026b25540ea467fc54c3954466ce914a1c4c
z627f9f87ade078bd223480962c3d58d100d31b977337f84f069f8cb53b62016e9a62e467b3a210
z84604ce039a42e51a13f64533a09c288492e11ae3ff9748d7da731ac9cd5b0bf6c2c4f7dbf7ad9
z853d37b8b7a942db5aa3b4a0a895267004753d4685576c620a82ed5639144d5cb6c808b78c6c6a
zd36cb41b22dc3db26b51ab7685244223a4480251e68838d432474a4d652826bde5f2a76815c0e5
ze9ab717351252e58d323792f50857ba9f5ca88686a23d737fbd62ca6d4720517ffc3cf9ed6bb7e
z0be42a74865459bbe21ff90ae773298de58e3c71d11e5b7fc9c3abbcf52d75b49c7a0f6ec34b92
zf74b2b155ad9cf841f7f65b2098658a7f81379ed7238944f3ea0f7ca6cc5cc50ae85853f3b1a8b
zb1e47c59ea046b7ea93105360a6ae8f3a02648414b716552f45882eeef0f36f69909947c40b9e0
z350bc339ab8cafae2c837e9f8406cc3d9795c91ac6351acbac567872b80dbaff0b5d7a84e68403
z54ea1617b123d60a45832f995d0dfe42a95064dab7bb90668e852f88c90d4bea3f1c462271aa03
z9655fe4dd306ab0a99d819b27cfb4e718f7db106a3552392e6b4c22672d7a8e980e8f47408535f
zce0d0f4f64a5d0c1897e3dddddb55f525c8a6586827ceac636bbcc5bc2ff370c773d0be1cad203
zc851ba3134ce920fc77e4e508e44a16eebc40acec6587fecbafc7f836a9c001d54463f9cf0ecec
z2edf76a4a479d1eb869cb2d96c39be3ef310e417345a23caa82301c5741effec22abf5ce50dad0
z83e40ed5d0dbe383a9b426670e0ffc912af8a4718b5148d8cc0a305d06bbc68de56d6b0bc634d7
zfffc1b8b148e0248b1b8501cd6120e24a07697cf07e5a8c7123c9bb86361f4e1c6769e5a3684b4
z23d2ff9e253291ab61455c6a70ce8b7d028c2eb4f428932c4a6b318d2f4114fef650e69e3be753
zeb1c07d1368eb313538468c192da502435346448e780859a3940f07bc3a97a67ddaf99a07eb731
z2027a05bc567ad8c79bb5d3c8be1984e7392e43725bf9808e7b41636cb58dd1abd80bfc0c0b883
ze16e5232c4b880b48b68e89407892e3d28a040503e25160a5791190398fc596c7425b11048e27a
z0a58043e7bc7a3f8fa765ca85c1b02fb7cb0f4f4c6d56a99fc6cd41122ba1f0257983bafab1678
z8949f470da801cdbfdd788a253f01e96d6272071cbf38b21f672eeed45480d6939ec8ca24ae972
zba06e2b55941d11409e65802d50ad86828f46bfd43cf02f112ef6fb2a1e9c21bcf112d9e488dd2
z0ad44e72a7b76c3db6479d0104549232f7254b15bfb9e348d3b2b70ef20b9b96e6236a1f901b3f
z850e7b6a45ef1a5bb3149612fde080ccfacf53a6a05f6ed6bc280732174353a68430bcffdf61dc
ze3fcd2b993b471afeee7aab65b9fd0754a26dbe7331fe2352912a6ffa52feb1b4ef16630901dbc
z75c4c395e40618764fe03923d936aabbf48df8a37d8daccce8eadaaee2d6f7e5b35bc9ed2dac36
z91c7d5d2f6c0b104f2f6b071f97d6f9d7525125b81ad2debb0da129c156d958600812756932fdf
zbb67eb01543259f94ac7b263ec6b95340ddf7219748daf90353154bc557cab53e70fb73086b08e
z6717e14d899e138fd154f586890460b86317e405d44aa232c07e35bf3313a6baaa02a05cb5a48d
z78c92daac5320f1bddaaa88b2c1b81c5019a921c0a581ae2c3fd58ad31ffc436fd1a4b8a9ac06f
z49419303fbe2e10c8b76fcc1275c741cd2be8170a0efb57d02c4fc76b96ac856db7e74b0578b16
zf8b8718a260a6ccc3ffba15ab8c86c5dce44d6f4cc1314e1704a8f4ecdcd1eca90d8d2b0454a51
zeceab38741c8e32e2526d6e09044225ec28f14dd57cf75c2e2f95f8f79be7136478206367413e0
zddb80f4ff26cc3ac96d1097afe77e1231b9160bc3c95593d3fec561923b5e099d1922b76139057
z006d6c6eae7a2d4f3968ccce3ff291d3edb857856da33f471910de5737a80fb7d1eee81efcd63f
ze0f3acf246cab7d29c5711a2f2e25df817d955b42a108e8ce35334e4a70d7a3b6d846024bf083a
z76ad2a1ec2dcabc396373e9bd861495bf154becf7aba0c0b3864991a12e2ab25c829e1c135c02f
z611bf075b1e8d8549b95991144acca7fd2e73784729d3dd49e11471ab11fb00f9207b421d1d97f
zc03f1d1dfe750d6af31e351a94cbbde87ced0cf1ffc29f637f52f600095e14f7ade4096f25ddca
zb8df9f472122977039ad6bae8c03402b1da755f7e40de4825c7bbcdd2740e9ad1970addc789e2c
z7cdd3d319dfe32bbf6dbf1bc5086796fa190d016bc317dd508cd59ccd651d73520c5bee468f499
z1de9c5bd8e35ffdfd5c5e5c8d75fb949a41dae98521d5d0bdf1bcb9cfbb256cbeae8da93594f7e
zbcf0fecb92db3138d2428b585561de7febecc5fae0b3a759ca1d38c0f8368c62bc853152dc3f4e
zc5c396fe34b9dcdef13894bc4f8cd49948ed87e6ff93bccb515d90d4247e039260f250ef76d1cd
z3b4c359c340115f33f72c7b5d0cc177ef9b521d6761e3b65c397e9410bb98a4e1193e928e5e981
zf2bc96cc8b9961ff98b6312d5e3cf81109c806bafec8c061ab19836e701f171bef23677f4aa6cb
z93d72a80932f56b5b4e142b09b47a0417141d32507b62629c31e6e052906335db9e158b84f4d8e
z096faaf30a977e9185f1f109c9c2c2c854ea7c2dbeab43522cda630ae49fe0aa244a2ed9e68e6e
zfde4dd2a1cf1485b3201f98809ee0e5296158cb2062d469c2a368177e7ee2a4acc94bfdf602c57
z46477be81dcc1698fa953624e95431d2ac2a13585caf8d396de1163902bed523ec6e20d67f62ca
z597c67f75261a1cf988076f2ccc3ddfb9c7fc435ee575bc06b4bd3769831ebc0fa653c2cab0398
zc4f9f4e3844e552e6b4349746fc49f7023b1960d9dea6310b80ae33b920eab6c1a8ca794e73542
zd4242a9d965baaa2656d76849bf1473b1af7c2acc1e9177129d8e8db009cf76cb29fc435ce652e
z905d6cc6b691fd0742a33aa2dfb4bc0fba0b8fa505f528c33e1336044a8bc0ce8982408def6e43
zb8b497e21aface808350151bcc603197c8e844b4245c6ad9b2215f2534f0ec1a8e747f22e74803
z93bfe1babd74d5539e9cbe616b430b3bbdba2ed6caaebb291d91341477348f93abedb5f3e9bc7d
z0a3eb4f61286fe35e341cc664043a9078e70892623128b83a11940bdc0ce326811c2801a2b4ff3
z20b810872c7f632abaeae5cb8c165a09b755c7cb0960705d58507f264aa97baafa9d466bf98e35
z217a32c52d9c31983251ef74f28b7431ccaff77a523d7dafcb6488185143d291bedf28b529d8d8
z35a2668f13fae9cc59183b796719fe2597b6168e2c43d9b14776c559bfc2400dcf222ed0a31c8d
z8365eadbcd6a945e29c463ef68665bb50ad0614affce56acfc2f873c3c070a295f75a1de701ae2
z2d05cf14251560e509b49d5f3245b9ef6f3aa06a76d23c14efb980b937e98cf8bbe465107ad1b4
z54ad8059663657034b8ad1d4408fe98ba6eac41f0f2af873ac1bd585f97baa01d4013940ea60fd
z17592c74ca20941debda66e79dfad61999350a897c003738f612a1bf201bb16bbcb6dc4fd51874
z8c6d12097e2e62d7610eda40876b7faa4c9c4fc18d5f35b2f63e99fdec48db460b89a5823c2485
z24bc9704a7fa57c999087154cdde4301d6c2d41866fd367cb351719d4e8ab997b31688aa941ff6
zb85dc7b56f3b60d11d8ea9c9ac956f1bf90cfacdf1fb9950c222d9234852d0bcf52ea55b88169a
z80ea74237c1c26918e2527d0bdc354c544f99b9366c50558995bc0ac9ba06c69fd7fdb271f0ba9
zbed153f5189dabbb98ff341184736055cdb904413a9d2a4350293c3cc5d7074b86ddd3f4cf8091
zcfc472546cecdbfd790beff0d73093450b437c6752b726b913f27bbed85d4d8bb0db884c228325
z571eee0198ad83ba1b22220279fb78158b70e8d6e2407f44e68dc7b582f5e3fdff46a5f49585ca
zacf930257b71d2a9628b98caf05544e822ba97b9c28c2ed05838224bfb2f55fd378fc84dd74590
z011ccbe2a15973a71924cb100d3b24bc298aaea540a151339d538c3d4322ea7d87ed3d1eef4e99
za042813c87113ce6fd3a8a2d64a92f5becd2da00a9c4345a158bf848745342294ff0125c839409
z391a05793a17e9715e52a6080ad192a6ad715ee02bf3efcd951c79599d71662fbcc9d7a8f4eea0
z95ad59a7ca34a9640b54c9cf10cc3b29795de3853be731c377e4e256fe64a5f435b53b82575d0b
z12bbdb3b59b68be40ed2193c4bcb6c5f6faadc97d5cc381580ac5fc76b997e7e9474190d7210f7
zd2132a88f4ca6a82d5d4d57ad6382f9ac63171f7bac55080f6bd383fe99de879a42d4c20914d73
z816d64c540aa2cfdf319a64f3e29060e097c5e6a2aa05f9820af862bc844bf3bbb3ec3bcaf109a
za1de294537bd2b02cab33adc898ba4ee1f1e530b9fde768763454865319819f013a3dc32755ceb
zcedd57641f67e89d727c225d3779ae0e146eaebb7f5f8979f76ec1db038181fab37bdab9bbd0e8
z8f1b0d5354e505c7df1a40bda0b3a25565c2b1e022c7025cda2a0ce923d01f7420c39fec615a4f
z3b52a7ffd360841134615e29dca54fd3dd16d4359afc2474abbe3eeab18ca770496883f97c7df1
z3804fdb7a419217ea63233bbe259bb239fc3a3ab83e6a76d229582bf74fe71d5f4499ec60fcd1d
z004fb1b529ec44ab4a303a7c58a65b82e8117c45ff280b7d6369eb70a2edd9a5dbd906f4c40bae
z8ac3c13d2094d63fcc7faef5c6b8cc6887220d81570764ca1be19f63e385499cf6454b2323fb7f
zf6bbe3dc09d05c9d2b930ac3c0aa91ea300de81c6012fa2cdd00798dff2a5b5ea8c53a87f203a0
z9162604a5f742eca5127106cf99d720f8722006d84f95f6c2aa750b81d50588c36d36a6baa678f
zd3249139b9ea4cdf370e7c32504b20ce9f07e297d202a833492aba9f825443a6bc56568bc29194
zc56d9260cc9350dc4d5ced4d72cc1b788a0bd2e7c836fb53da45ecb0612c00c9d4c4ba44b72db5
z3829c2cf425777d317fb48326ebd7daee2538607c004118538b8cdea7d435f05b2367aae07cc11
zbf080536bde17d42f68aeb0b2af94d542c545e05af84d25deaeaf8f129c9819213920953e9ad0d
z2089cbd5643e68870254ed43553c72e43b87857383faada1e1e9ad215ee8c017f5a38549f99dd4
z69406f6d9e6ab67e9049b229a2a111aee50c9288b1eaf15520b9db40369685c7b9a47baf49f18b
z28d2bf594a473c9425ca184c7ff30d14072ac1187a6890ad63b0da0ef13c436010de78f686598d
z32d8ed08c4c15d03b8556dc2640cdcfec0b038b9dd5799d76414988efc9e31f68386071236a818
zc10c28be33e53bd8d52b50cb2e47a71147cd43f6b154e0784437d2aab42d05b971a0141e65e911
z585ddcdc3fce9a894b0c580e480d1ef4aceb23b211a9f778f55d07f26729cc6bb340b7cc6a21b9
z3c51fd8aa1141be9d2716176dc6fdcbd8361d8900ad1715b7fe6b40c2fe37f08210b3b140e89c4
zdf1a05540d0c4d2e8c8e63a00adff30cbbeea507f5ec0897a4f32d2d69cb8bf7ecda2932e29526
zb6829eeff8216153df21b2a66f37b3dd9220169dfe4cb9bc84ad0e12727cacbe5ddcbb022b665d
z611ea6e8f4afb047360ab641332f590d85993e2a9078c89c7485ca5cf5d6f543fedf8ffa484699
z69a3442acee478c09c91702d32653f350494e28f91c2d67a3b6dbab93952ee9df84e3c7d17a4eb
zfc1d308e95f62a057fefbb40e5ce90a6af87ab54ee9803e86bf76ca8f54c046d71b2d7a2141a1c
zc987ec5192943aaac04a7be8de40f2c307e045210f5ce733f23a219e49bde92aaf2b397cdf8c65
z9db0f8f92c094baa58ac46e0de86b700e4a4311d9b221bf1940a748f39143c360a71c0131a2578
z13e886c89c41382c86d24eba8f15d93c07b65e7427b1228325830648b4e776d5929724ba791bfe
zf39aea38e7d3dc47c46b8189166f1e6693e632957e5bd58c596f75238066ae6bea27f78c74e273
z82effc4e2750bf5f937e855d03b43a9cc4ced946e7cd13916a3c0551f050cf32d8be45fd22ed51
z612394960a641913aa01cadf85ec6ff33979295aa4c7549a0f5f10c801996b5cdcf191a1210116
zf4dd3393cba6d161399b7ed3f13fcaea745d5eb66f80e3245fc971ff414a543af8442b61d20ad2
z7ac25a521066f5d841901f1c01aeaa7c026b3e80c1022a7b60ed3087b92d4211763791e456cdf6
z43a77836f2c63c6f969faef3a5be4d3794d9eb8cefbccf45b88b6e91181b5b24c5af6a23aace83
z3d73649943d6d15cb561fd994ec2dc8fad54fac939963635051ffa8407b85901af869e896a0a35
zbab94509dd0cce1a5e9044b5cb99f945c76c15eeec5c2e27dc4ca5c54d5a0a859725c2bdde6bdc
zb1d701e0d6b8d09c0c5c81ad4c663cb1fb2edca555677e44fc288a5c95d050283afc604f101a8c
z4b85af013467b9a760845e7ae723605eddddcc9f2d49ad7e00a92d6785ee4c80568b77ac84cdbf
zf3e6151c16fdc91164199353822d053ee3050579ae365ebfcdda975134962d0f9c30808a7a2b69
z12cd5759fae7824cc5b9eca72f8070f368cfd4253b1498f381bd177e3da4a1853731ceecf79078
zc01c4e16fbae73961b00dc3ba5fe44fc433a675b9840d43951d823a1fd0c442636db4d0f738f93
zebd90360b348fb45faf548fa94753509637996269b2df747513ae0264ffcc1964274c91a383801
zac972df0bc524f83acdfd7a3d6c2b8e9a5c0a46e6cfb245031f17594dadd808bdcd0eff0dcded0
z59bb9809eb00bcfab85a730ddf68e9c76dc407e1dc00b4788743c8fb3e230f89924e64ecbaea35
z42b000a937bb2201540b06e8c2cd61dc684aa288fc817ec60ac12956c2ecfc97db5158d2b01f6e
z80d189e7c946330c8844e40ba0096f49fe26026581edd5f2d1a77f5c417f984cf5d2cb0a8e6112
ze6fac3d853c83bf09892eb53727e63922857ca522d3f49e624fd669b247f8b9ba545083de40d3f
z83671f6fc3939a181d861da1733e3e31735a28be0cbf22b07d4816f490dc3c147dd747b0326cf6
z93db23cfd83da7f950a46b3ff7b4183dd01a59477320d7ddcf2ce8dd711f4756077ff904510495
z751a4ef927f5c8cc622a047286feb646704b8ec0c5f3ffaa6ab838cbd1a1a08ce4bfc89ce12dde
zdd610812c3f5d1100f6215c809dac6819dbf8445358698c2a01289c975822d1bc8f4b6c8abf31e
z8bcc32a21b383090449af96ec37c77115bfa7d1544ba475d3256af9a462f290ff3ac8f36f01852
z54c017bf9a9c5e17d53f95f63b6861c220d5d0620c848c892e4010c9892fcbd96f6fe846feb959
z54d1cb37fa1462ee34c2646315b83600a2d0906a878a8238de20f031d3bd9a37e81c24d3a6cd3c
z4c8043c100e38910a0fdecf307d1ca937e0c6adb957b2bca2ee597772caeacf284d5ee14c06c5f
zd05b63fc15be0fc817366c5ae5a04cd95734f248564e0277fde0237611fcc01d34f694a1ab3cea
z7555fd5feed529bf74ca75dd7ce914489dcc7ef5b73208a3b7aed5f237fd90fb262d43032ec689
zd37ab7167f1eca57e370ead785907d0e9adb44e5331cb6241f69ddb8b7db28522e8bfea42e0a56
z190865b22657c937ec432fda2b1f75463523915bd2dfe312f2cc457b724a7c4b38a5ce71291a10
z27962fee183c0a042f608f0a9b6fb0e6cbbf963dc8bb72dbd7d8b4be2006036dd976b3b3711c62
z2c4eb0db6865a57832173769a7b61621fc359ac8474fe49fab52cd18c33b0cc739ab954533953b
z419099d4c76bc3d688e8ddc5904bbe7aad2086924a4bdae0506fa3797862bba72064125491ad59
z2baa0a29a769b996757a7869dccdbc69cdb9268061e63a26d1ba9c35841edbc458015668b29a13
zf96fb06fc336b94b645e1be8bb1a72247884b4f2e34d8111ee61363035ace27b65c4acaaf4d450
z2de97c349582363371cb72e66281278462ba9343e0b6528814cdbe8435a60781a4df093a0ffcde
z902359fc7e4a9405f7e151bc78d3b598c094baab219fa9ad95d1f67b95af1f56b7c6d1c13e06c1
z702f386dfe7d4a2a26abbe11c2978cbd77743a796c9a8ac9787fd221eb171af4cf797c940815c7
zc9f5ac4835a5579f65f7be0de1100ebad1c980f1d12ec84210af6644c34ae3dad11c04a5b4bc8a
z06d9589c6e10c3bef4652a9b11ff4d9b3556592e736dd23669b4270696434cd0da068fc82e29fb
z6cf1eb4de0f1834652809d5cbbf45c8fcb2c40ba654531832b4db3e089862fe56e68d7ac2ee590
z640cb03e314a10dcf63b629877f87033942856ed7b71a1a467bd46adf0f0b5860ee20df6540742
zfcf42674af438b2b3842c086bd76a613606bee9d39449dcb0d2efa4f1201fd232e748ff0773ac0
z0b6c90ddb93e58b1a1fe278e1c477d2df26bb69c06c06025559accb8ca76b3470787d374c36fea
z04a47ab1f3c8ff09c037a2f96e9473a1c5ce3ffefd9bcb5730387d2db573bad4ca6410a273af6e
z82bc2395d6392770950d73cdf943b48bcdd64e7a6d3c7b2bbe620387499f1ba478d9959da5c92b
z84ff03d3dad0f4aca1a6a70b49e5d9a0f6cb3f4620cc2a119291795f8429bb57e4126508e18027
zecca4b6f380e4baf438ba382c299964d88617dd16b158c240fe496d9016ff9174f61f0f5230955
zfb722b4b4e8514d6038f6f4c3e7e6a40415937711631ec197b6822464a878d9dd0307363968663
z202089671218977f082227fc40179704334b3326dc0f01d19e323138bda05517408807104a85f4
ze1c9106223928a4d4a2386129a2cb591e42b7e40155c3040f40d4d5fab1699fb5a4b8cf46510a9
z5b8652d3f5b9961e81133e4a3fd0621a4d1270e8f6a12499b72ad91a2f5d66e4f4028c95260533
z48e50123f14091b79aa3a7ca4e44ff2c6ade7b05a36e7d2b0a7db7a6c447baf7043c86dd056774
z978f4803308f5c8916a8ae2077be3c886e67b11c206b8ce28e59d11cd6ff06866761402089efcf
zbb4e59743d41be2ea5e53919ddce2398498b1d815b05af592fb6dff052e9f5109366f7d0cdcc87
z26cba7fa3d87e3b4798981d84280d716ad38d978cfba8ab547c6fc8819dc7413ebe4d47f93fc8b
za2cc5220b6805f4bde31b7e4ed900e25fda34358129a49e33eea3c1c9bdacb748e7ab26316d943
zc352faea0770d185a4837eacbe0e504ec60d2a66cdaff4dcd58635f2fcf47b7d5da749cf98c896
zbcd7709acf2e41c7af80c9a26b7026569aada5512c0ba7d6c67c2d20c766c7b177b54961ee8303
z7a21368bef28aefb431d8afade31b4dcc41288a667b60331b97581d4f7eb63a62ef9c07fc66875
zef79682eb9a709605a84d840b552aca97b47e784e062ac4bce3e43d3f39067bb257e083d2b3a42
z6464b26fb499785d2e0c95bb15ce309b57e09da9c83e1482ff5222bb29e19c1fc13e4495d609dd
zb2ac2b87949290d8c42514e724f3c578103e802c71a95b702d778207501fd914942a3dc5b3a68f
zfeabdd5843e200f0f3be2b9eae6e5fec9bc384491fff64fb44da6b2c5a1b485f8baa80722e1c9d
z80a3b424c95c7ec41f9e96be5bf4177748a4b8f1c6fbf77543929d73e2946a13f1fb31efc90f18
z3ba894a1133b5cb70836bd7193f38a5b4c9471e95bcceff2e5ff97e7b3ec80829d5e6618ae9ba6
z0466b54c63e2ae984a1e24f8f96d02ff506ca9e3f09f350d6c95ad10a299aabdc4eb31abdfd755
zc5eaa620251517a52d4e0cc167aa01a31e42286687394ee3e75b7dbcb57136f1ce0b61a576690a
z761517c3d938183ff06eeedf28f390fe382336e7d43cd1e517e9b535498666a616cdbec6cb71cd
z7a62aca856cc3ab1e5d785f2b3a94c60019ea47895ea5e942a3455b59607c1c4c3da71f3f6aed7
ze2ce71ba7c7ed04784bd0cfc237edd6f3647cefc33ad5affaaf2ab6709cc55b099a8bbc00879b8
z04fa56f3017245a6f92fcc985eb98751ed876c8ad0f372a0ed9505a47245c5f5f8edbb124b01ab
ze84681a2ca974e3337845d9bce3ff982406b619dcb90bb9a501dca42d57293d8ee0955dd595698
zb58554187c50ef571ad0fc180045452dfa8f4634592c4cff0274c097962531df294c033e8bae66
z1aab00c73dcd8c47a1c748a29b6a5b17c671329ae6d0bc8bcfa79051bbc362efa1908db785548d
zbff14a73f5ccd3c01e26f111ba386a84eab95bee7523b60c2239c14742c20780034c34a5407e82
z67a31b2431e248974ed49bd1ecaf2b3244a6b30cdda6d796217cbbe3ba9dd3a0e6c98bb06a57dc
z85fddacb494f6d5cdd259f7a34608bce6f9fcc7440e66465408e6f7b0902bdc9813ea1baff2c1b
zb4f323a50f4852753ed5755a70bf53ab404a8a101bc362835827e26530f1f0f5a7383bf78418b9
za4179aa324d675929db5b2f990f1429baf752de43152c62fc8cb783ab0b334def60a2a2c809588
z2753d4150d4d729c0d5ec39374b33ac1a7cf52a6bf5ae1d18419144ed5534a468e555c61734b8c
zbca719bfda09e1ca54d0f7e550d3c34b63bc63f38a095aafceadaeffb431b09a7cd20f80ca0f96
z41f26884c6a518a8b0d78d87f7d77bb3cedd79a47f70bee9565ed12a135bce0f592c3a92abb52f
z490c7b76d5c588707a724f106843d06dbcceb4cd6c501e2d007398b341deb99a6d41b01bb5e1fa
z218474ac3318d16a5b08d2a4116d6cde96fb344f3e10c01ff7dd2329a9397825dd1492689529e6
z06ea13b61a1e22e6ba4d63a266449c245038b1b3d7d3d062ee2fd99e72a743bfae4a9cde869717
z6416766f7a44c3845cea73af1a20e1f97cfba4a9431d371c9006663e860f21c14bb810905b55c4
z50345b021843dc37e6a267d323c0366a29f94b1cdfd0482285c38bd78df2d00b75e0b0947369d0
z343b09209b2ab3d8ffbcbb4ce2e5201f1ec4a450eaea96a9c5389889ea7cffd067ec1bc9e57988
ze01319f22aed862dffa473b92fc5585063d5fa393725b194b9668c6229f99e0b95dc81f3626e0b
z8bb86fc468704f3dde9bb9e00b7ba239178a9b8acb3f277aeb5a115da286b5e306efe891495864
z8593bdd9dcae9551c4500e70cebdc666ce823a4d04ebac82665da829154e005c5ca6c379f4befa
zf7e2a0afb7027bd9760491c446c962f663ae678506c5834a89f2afd0cfdc8b7ebbb9549ae923ea
z15a0ff8411a1e49d20db7a179cad8e51a0906a1030340cb2eeb1e6df36f9040ac96a6dbdf4d024
z80dba3def3765707978760f38346466b55c74dfd77d35a1c9899dfdd97d11c5f7e3f327544df9d
z4ef37955000616bd93223a84e726a4853317d2979f308c8f17f2244bd0ef75aa2123bb16e70afb
zdbd9f67acb9a29800ffa9b83056998bc217c9667f4ca07f553dd2c17bbfa05fc7750b47260b183
z8fa43d5a8ba3b194f3046cba4c45a64f8c3df6d4a6bdb205514b4a7823a3ad0bb2dacfe833f8c9
z16288a6b4f620abc733d06f29d8d2873e0920b26c3a01e5f8e0758f82d894c8139043e08e467d8
zba8c6fa01ed8d99596a94311a0123a4b0f2b1764961841924ee57099faf4dc85904cbe419d347c
z6ee8e87c29ec342481a3bc2f2b79d11b40b2a0c229da5c007096b3138cabaf7875a5cf77ac64f9
zb9d8990affcd8aafba6d80537b8736aea7888611cdf06e67891b950823a2c132647cf194fe3fdf
zfde2e8113251dbc0a9c8bc6b85c1df8e97e5c3adc9c6cffadbea04345674427fc3f10640ba188b
z4c9c23c02464742ecfc62c7c3425554e1fea8d230d310b89522c4172be4eb2c3580fd933fac7aa
ze850a19d7dfaec94eeda73fae531715120e2a1865f5f375e7b84a60c5f24d066809a51af04db0b
z96d594bed3ab046cb9e487b44f4f3e88657284cc6ca1b3355099d571ea1cbf1959ec937f6d21ef
zdcab91e1f8a956bbb02ce20d489de820c2ad7781179a032a45140d4eead30ad131c4cf5990f1d9
z60eba060a11c1412cde8af4d1ff022c96c8a63718a0236600f6956a445517aa31f363070c42f7e
z3ed40b2a1994a4f2c40654949d3db869d6dd61c48d674e9cd2a423371e336e448dc8dd60d2d761
zf03ce9d056ead75194180f0f555b0387a8afe0499ef7c77352fd76da1e50bb0a27417c335e3c77
za4f675b96494175f204b88900e5109e82b0040a93c42a8372ff0c43dd1d3e3e57024360268832a
zccef52eca85d81b7d5673402a62457c515bcab407af7c42557546b48daaf4dc5482c545b3cfb94
z7c2466e1420d6937a33cf78008fe73e6765722eb0ee2b7f2455c29f06c269440ac9cec3c236179
z728ed23b76f9804518fd6d3f7acfbf563535a30f5509254c264c2ce987e15c217066e5c684caea
z9575469e3cdb5c9802009f30d0206f3f583b8fa62f2c8f37136fc4bf9a8dd532ba36ef834a0bd3
z56752e6ef6cf640404896c9480434a5f4b0387f0eb588aaced4f14f00d3ceaed2375464cdd7e77
z6c993874135f19dd293d73fbce901b602f98d8064df733cec76f951982fbcfbf3f513fc3f4f1f0
zcbd0c7e1da392474e6c86f6e33e9b116624e9536ea531734966da4b9ed913c7cc9db4e37185f69
z5f444ffce8821b1b54695c75035360a45fdd07ed46647b9ad0e4e79875b592f5a4721aee4ee218
z543f3c973fd56eca3dc512f12baf7e3f53b056e06d58f6ec3c7aec8af7386307244efa5c8342a6
z3c50f668f4ab2bfee33689fa1a7c360bcdd72b1ec4b51caa1251d6c916bada011aa7fed65cff7d
zc8deae228c5bdd538c61ddb3cdea95fe7eb12b2d55c8bae1ba546c5cca1d656b1c432cb5b35b56
z5b5a8b4dcc3ee404b01af8409be03df75974f101cee983f7c9e6223af29e83030bb9bba203b9c1
zbf6bb200ee0ec23057f7db3f25c3a8ee69aa056ddfa4616cfd8456d1fdd02b4a08b39d13aca66f
zb6b2df4ea3ff00198fbaf85db7e1c411e08635b610495adccec5ed72489bfdbe658eca7adb1437
zaf28fae0f615ba69bee67e1c7049d1292e32beb96a8a4bfa636ecf6ea1c10056df9f77b85ae771
zf404d0576d6cfa661c7b6a782e4d4c9b5409177f2354ed0d3aa6b8c18d08767624b53d194036be
z011045d3178792b1e2e74d94a4612dbc30582f64b9cb21f696477edab19b5dbdf1eecb75d0e812
z62e210a22406837520775df154ac12d428fcf8697db79a00f928eed7b6e37fdfe455d7d4d546f9
ze6d584c4f14121392974c5d2a0a2c8b88c189c04a87fcd87cf71382be6b378b9dd994e72ef9433
z429b88b84f99bba809931af1b693089089ca2000f7fd1426d22bc9ddce2eaeaa6e578a82b5e45b
zca5bdacb8c5f7e5e5fae28ce1118f106c49f8fb5fa05b6e44e628930cd474cf32bc9942d2a1b2c
z3881306150146928157677f574891db93556bd54dcfebc3fa49782290a30fd8cee0dfa8c00d988
za3743af2c8c786be4954fb91fa52f6130e393624c3b9a11c7c285a3caac53946b4c8f34b153fc0
zbdaffb147f7f7b6ee4178fa35f68c6cd6dd2b095b8493e2cdf435f209af81bf4dd3d33e5b97d26
z1a62294620e77a3b004b0657917d48e8b86cbcee9644bdc4d812e41c1061e1cc463835097f9d1e
z095b91456c00cd1f81853b92d95f3ecd172ea5521d86147078d28d65a5af689783663f65213eaf
z5dde753fa0631b07267539a031b4ddf9759bdd61c1de6a98d4b967fee461834abf3588480cd83e
ze993234049bd0b8cd6bd3c90018f0d6720d145af510f0af5e59b71e018b41f54c1491e9b9e67a3
zf762775bf4b0fd7ca0ece9495b7bb14df050c8b0ee27d2cadba40fe7226a078a594e17ff1b6366
ze088c4b822160bb1abec1c31f1855b3d9797b346c2303790956171fc7658734d75be9e21c291fb
zab9873ee88cc4acd59e19ca795cf5e1ff063bb449e9e9c9d462a3c4036914e888cfbb3c7783290
zb9ee2a20c7789aacfb054bc7346d18ea14f8809a49c1225bd7ab82c89a2a252dd01286db1e7f24
zdb0e881eadaf38185b9bcfc6191deb0457975200b420a82b7d808679c8ec95c56d6dcf3c73c74e
zf1edbaceb8b10508b70089a65fcfae9f45b1f0af672ce5449a74ce74a36952e859eac1b8e9e2a0
z97276bd5f906173f44e2c7fff4729986718be23c9832512ddea3c54580db1d48295e4ba10aeec4
z15d07cf189600b24c1c8a42e08ece75b8652e4aec1cc0ebe9e1b77029a0edaf8cc5057a02ea9a7
z6a4f97c5a9590335b8968f8925e01bea9d1fd75876b7ef8f756c9f5a24b4a47ee6bae2bbc32db2
z2ca08aa1cb3517e23d377c4f84275077ac7c0ba0266410d45cbb94506c06c2ebdf040b498130ae
zf1ea2ef5a1c665d1efa47ff36741b8835d0f4ab037f1d8477dceee7f670ca8c85e39b03e266004
z4dfb3055bd2eee6c723883701b411f9619ec4aa2ae8380d3715b4b037c9f1fe60288deaeef12bc
z59e832abf66c5cc67d2c95dd7561018d994d679f3adea2ed14472378c7c00525c35ed9556382c0
zac3160a48907d098104ec9e02420e420275cba73a13a32260b5935ef8b2277554173c36508ca07
zb63ef0d6adb52d89b2e81ced139aca75a641af81c6a81420db58032c30d6c97dd90271794fb16c
z304e3ee68bddb098666ff3c88c9209ac78c30e0111876603f502f265d450a1c85269bdf5c68129
z6d24a4ea9336ffc1cbf385a89aad3b708f6384c07af7fe093599a17b481b770e4e26352c40944b
z8a0cec734a0f1211dc46d77344e86f8a7e4b713cdf0001aa791b721f791bc5d81e707d5361f617
z062acc760955ebe300cd91104d17fbd78181837bf8de9ab0dacb9de7ac13c33d890184448a1d8b
z69229f9474ea1056ea6e199f0218e40d1becde624aaa2d9b6890b16cf1f6e1d243559fe95eefc1
zcbc134bef7e1f977a348600a812692d3d6923e55ae86bde8dc11232f47a075ce39d4d257347781
z4ce68e12b997329b2674f67f12fe798f352ba61ad8c561106b8c68a53b34ee981c85fa3d25f90e
za20dd8526401174a2af889347d1970818c8cbd9a1af3906995aaf615cabbd59081f389279dfbb8
z7909cd10168130d7aa77a8bc87a16159c1abb48366e033e9aa836d5b642508ff6f31c07ce1bb89
z48471695e7216a8b57e163ff008ddf4d62d454ceb9b9b30dcb6397acfc7beba70dc315d8f41a7c
z490c5d85999fdd5043728373019ae30c90b985bfcda5838afb6516e453ee0affa822f0af147d18
zaa8471407d5e7358db1b8e01fe9b488277aa450245c014340349c6050ef7e78ecb68fc26811b1e
z0e10d1bffdc864cebd4696b771055f25230aed715477a8c58903aa8f6877a2ec84e95259817ab7
z53db8fcd89641bec05564b869b0c7b60d6647fed2c0596466e8fe5af0d5eab36b35ceba57928f8
zde85e2ede95ca00dc0359c99c1fc640e5eee3bcb83117135903282c7781b69185ad38f56ff4b80
z6b387de7d753ca2f994ab1381d2f4d71ef01c287c7f8b6676daddf6b375071390e34fc4443618f
z57e4603babb520e661ea5a471230338b694d25fdeb980f60d580a6ae319f08f62d5f2e1d6ae869
zdc6d0c1f7ce05961b447197536e50498d52920ebc748210a4206e5f05c30ba24e8a4ab12dd234d
z4aed54bac2bd77429850806faa03c1ded31b0e820e1256da1154d7566987ddb87a1412e1654b4d
z0c3b0e99b593d8ff24a9faf47fa255ac4a9369d6422a932a0ec7df034f056444feaf2aae819294
zd35caa2dde6e7b648f76dffc115bf5c3de51b41f19bf7becb4f06142dfc134bc7e44d3f97deef4
z614cd4121feaf81ec4f96a83a6e0c52e044412942ee95fa01f52117229951e7c8ea71e08763cac
zf393d61b75da8fbf28fe2b9c2afa735077c55159496469057b6b0faad16d48123eefa50bb4a71e
z7d4bf02be8475c970fdeca826b0eed28c627a810603f5e588410d9eeafec272a288636a070b154
z064eeb7670ff563a6e3374fc35a902f88a6ea2ffde9611fbedb47e47df22a1bfe3a28b653184e3
z3b7456deb620434faeadc729d8abecbb8654dd64de7aa7cf9cf50a414ebb80c0d5e18ad8d40f9b
zde51a24536f47bb15723fec4129e1660868f9d147f092bd2122dfec5858fb14681907507201f00
z8ffa053fecebcc3f8308677922ec77f14c4436b7732dcb7c2b09e08e238fe8872c25197a64d22e
z5670c8ad0578b0f698819b204ad2e9309b49677168dbf76f122544220c7f6f3ce8ccb935fcf674
zcf589b2843fe2f0e7e576b1f8be34f5efbac47b0887acdfc17119e59247101209d80b54de2180a
z5c90aabefc885b53a90de2d92a502fbad6abc93b576dba26ac94587b1ca3ec0e90b6df882d9461
zb3c11270fc50bdd059560de3022c025e2049bd6f3ac6cbd5fc953d3ecfe3c77c17c5ee86d7807d
z9f9ad95c6275384c19a53d69dbd6a5be92fb5503f935702adfc09c5a29336a6bc4b7d5ebdd6a43
z6314547462223376f6067894d5bf285a33be461d6f8c86157ca929e71951eff147069b2e70d2a4
z796ed7edb0f9f01e01a7ccccdca297f0deab0d438c1c638f0951540d64bfa2deb9ee0b2f7f35b9
zba53e1e4510f9d1c211b99cafe739b33bec49a27621fb7b5b0b4a4ec4169756ff7b087422e896e
za4b722d888488db18e7b9014bf0fe3c83d2b11899382356342c8de64b486dc231647c6c79eea16
z87fcb4b38c4d8df2616476fa77ce80f1e4a666e5fc973a3571ca4dcdfa7a091b353805b2f2b240
z8ac8b5d74956d5656a22e576244f04bca0198d8ce0ba47a923e823a896b81ab679d57019980e0f
z09503812188d215118292ddbd40491de0dce81f78f212a3264adc511a366b8bffdbba3ba67aab2
z3556059881ba0d5eddf8a2b53266d1dfe55385af64f3843a49a155ec28a3d151b8c790956992d9
z21cddcfbdf3c43cfca41d81ab83180b08991c6d0688d6ec6ff97cceced87a06cf47a48cd878d33
z4595ceb3831c571a98d5af5d3176ab998cd8fbc98933b35209398f34aa33df6b5b3e551d1d35a7
za13685b57cbe1807a4f8ce8e1422a652110a796ebc2a40b61d7cc9b6cfe457b5c8f89d1b00a833
z8109f83f789d9b355519baad572f2775b6f9d3f265fd2951457456991da63e704de741b94dccde
z95e464c65e2a3635ac27bf07bd6ad94a2155015da990f4a37cbf0ee6c2dfd378208ee10b2bf460
ze0b3eb31fe82b2766e247243e73537fcab995fd5518f7cca81a24dc375d1ed9a01817c88941070
z6562d7632ced861442410745523281d0d194318507faa49b45885664c7bdd8f268294cc7fe4141
z78dfcca09e478ebd1e720d08321fd14e95ccbe0d7df86b26377e27acf691b5dcb7d38f5a180cff
z4a5d833e2dc1f8d34ac393923cd05240adec4c8adcfc94071cf0a32a633c5cbeda934b4780b55a
z9d223c6a6fdecddc5d3de8a034926d906db27f990906f540286d22b069cadcb423e683bfd1a73a
z874aece2a021c6d1543d187ebd5e44b51570769d25c64a983429fcd7bf6665ef5d4c43c95d86ce
za906ae6f9898b28ace01dcef50ffac61fdd276d56864125d61ed62585a886c4ac5d264c61fc0d8
z2a85bf5a2b6a24b6a14f8c765f5ccff74f13f0fa1d396bf364f9b90aef7d91b0ac7a85f8d93500
zefa701213f968c2d23316d7d830cb2b6e9b0b5d3155a4cb335507387aa73f8b5fd93e3675aeb84
z2c8eb804a5ffc376b662549d50f9a5d3c3692a0c53c32a78bf9208c9af2ade6fb617a52106de32
zbd201e94ea3c184f40747aee46804615be3220f23748b4e5b784fe4d1833a76e375beed9e69693
z25bd187b886572180f5b738aaed908076f0112741703809ed5bbe25c42a3ffb66655e1c2fc2a07
z30be796b415c5155ea02222bd40211ed0439888ba3baaf4c30935bfc35fcc2f5f25d179047fd0a
z8f924c84a6a7e4f07fcc41399c44bd07270b1ece87be5fe14573670a8cff4e11107e14cbeebbc3
z7d6034824e07716abad6519dec408545c92f02f91c2390d1a408209e15d31bbaa4d9d14528919d
z385edd6d6727d20f457c4b239be919278df0eab3490403eeb694bcbb8a51c4811334a1d433b43c
zbcdeee0fda718fc9ab439001e004c19f9d614c68650b47530ccb399863509f626900d030c1e991
z033de1027b18ecc37e3475d57d89ce3a3763c3a0582fa868ffd48d82c03c1ea86095e2af149cdb
z74c2dbb0ddfd578d0dc5dc45dd3cb32b62e0333d708d9dcd15aa72cd66873dcb3d8c8727d7e52d
zf385b2e7c1e23e5058b0fd032136a761f49f20f0dad3500aa30d1a6849960199f162a538f82276
z6484b5bd19bb5fae9a35bbefc83f995a6ec70da1b86591cf79e0d5945866b73c8134939cd3fca3
zfffb0dc879e109e6959286634d8d4158fe0abe438e0f619bfed9e1972097b74ca59a366374cd52
z4f7592d2aeeab1d05cd1f51948a43209c67d1af2ea5afba14ae7b206057ce8ffaafdd98e212320
z7aa50e86044637f1c68c9907163c396b2010e43bd313b3222a03960f16b7674456dca874137a21
z5691d097d4dd5d0aec40c3828c484365d3005c60ecbcf7f36873ed0712a471f4dfb6ef6666f229
z51b055253efe2c0f17b21b0085ce023bb7f493836140ce7d52773c293ba427df74f236e5b64dcc
za459b3cc998a34fb9899028ae9108941847f14f726ffafa8f98c269b489e77c3648cb16f959fa3
z4a075ef3a1e5bf306fac413707f6755a4e68892180c2082af6e65967e03e509b64494f57f304d7
zfbcf0d9fb61069b263675dfe91f2fec496345f3739c63ae7cfc14f387e672f628ee3378a66d32d
z626d62ddcb41f4725155fded8b41e394154e8ad3d7c01d8f8afbe38fb2fdb0cf3c5e277f72587e
z313f9c95cabedd812678fe50f497b3c79c0e8c3c7183a0895799aa367b57417b9fb53f730babf3
z50f6aebdfa622121fb5a2c29bc627441b69d45797aff3183b814e56c9f1d6fd044be9ff7a93c86
z4d5fce843abdb9af0c4b4e1885bbb49f4d4e7a97663b3e04b8b5068ca624152bd0443b6152ba87
z9fafad50ad62f8ca29cef03aeaf877263b128f7fa6197d32bb2fe13969f8388c72466faad1f0ac
za33bee8ad6a072b4f4db098069ef4f4ce713e8c8a179cd193b87f2ffefd595cfe1f0a7952b315f
z5f120d8d221e7bbc1a0582746b658548d7b19fd47c1bbadb4ac3e360ad2c6bcae9fdce0283e233
z05b821cf2f66638fe29ac3942047f5461923af5977701d4c7f580adb41428a415f113b1bc47522
z288fe916c13638c443e09a8aff6561be978ae283f7bd163afc167d676bdcc0b6115dc34cf62536
z5b6996e4fb6224c198f85cb1a668605819d3772a66f4a7dc54c23dd9b9027c6f879492184927de
z6a8b2d9786349f3354ac63d0f0619e7e98cd240a438070470508ef3fe234dcd10ffd34faf1071e
z3a1fa0b43784212c434c7086dc52648db7e5310b7c87b5a608264a9ea51babf049d8d08b771430
z55d25b8ae8872a7665239ef4a643bf016cfbdc382fcc6ce55f478c61a60bf9738e29becf9bd173
z4bbdf67cd73034d4a0c90bed9a8999e3695941c4520780b2e8be1208d17045015bdf6ed097ac0e
zedbd1d8e6f917d3a95bd3a3d66631fce5ee1752474a33003c17fb0b8023259a8a922b40df0e92a
z69bc11b0ec118bfd2f80b80136f4585cacab84c656e8823ee72fb66648852fd14de00e008474e9
z9c79e6d03ae8d654f91c5f9568e089ab8849f48785427eaa10b76cb35d5cb48a30a424b7b4a957
z15ecbf0be67ebadb96f386bb81cb95b0ed62fe5f8819b98434e8fcc0e5e5d3f3920b961f7cbc34
zbef72fb99155e0b805c1df5c05a7fa0bc5728738be79cceeb0b1d70f3798b5dc3b683b128878bd
z7fc0ac0696efb7480a6adc841a4d248aa9a194ca0c353f90f20b01a284673707d7c0ed7ff026f3
zc60829c0393efb0199a733b08389cc6b3c5cf51fa58443b37023882c369ba8ca4dddc04d089ef7
z93a3a065a7af7ce472155a8455770e0da27116972632b425b671a91c7210af69f7fb7d5b634b98
zde7b723608273c186ed40bfa345b75e8fa676dfa66abebe55cca7b85216d625355821f45afa997
z4b52a213286aed9bde4a293f2173040ecc11649f9bab98c550b34f5e5f42db21e9c07b5db7c4e9
zf01b62ae16c2fe857e85f672c2782d67826c679fd72c9677fae38778ff4a4c43e1c3bd6b682bfa
z9a810bac465a0246b44fe940065ce12312c2d0abf9060fbed1f46a38e5bbd947c235a1e4c833c0
zb43886a7cee3e31956dd689e9ff85743c6f476743abcf25c57377ef2319a3f602bbed526c14bc1
zb76d127a77cb9f5206a1b8cf019b60620e90a08b2e0427c5f1bf57d18cb1c04c314c3513a7100d
ze333ed607bc4a3845730147431f698299d6c11eaf1f10faf6e03e5de326be88f05343783691ead
z7e9eb7a142e39bb471f63b46a294a921425bd742b5102e7c1f9fe889470f755a4d3eb9abdb4a78
z8b08231b8571a49be4a47244635c9560e95c2fa1d416ead2cc7660f8e682ccc554638a49b6e982
zd709954112736b74ce02f58898949ef8974f183f29c3ea2bc02d8ed5a4d70de05a3d11fffdeda6
z96721c9547cd462f9566defeaefa3425da197606577f0639f860a50e046d92c89e243acf9dcf40
z489937a9efaec6824a008cd472d1ddd7c0e69fb11a1d797f4af6a0fce4f669b9ad18c161c5ea2c
z3f838523648ab8a420b981d7dfa9bdbea2be8962e3f3613b742f94dd23ab013062c5dac2831631
zbd14391dda4d9006a33b7f98536ba195f363c82f8f7e15a7edc4a9070130f4fe303a7674c611cc
z6d2db9c16e9b86a2f6dcb3a3102024e7b121c0582746fffe53e2dfce74ac2f57bc5211723c537e
zfb97aef45fce8c506eb58f70da942cd0b7a8643cfc57607cdf0d619f0022bf5c2960519ae34f06
zc52e7f7111722c9d7294ce8717029b4471444e71f78566d3d8240c01e9bb1b99585caa1c390285
z70d4bd9be51a6d12d3799f4769ac6825ed7327669d4365c9d37236bcbc6a05647f1a1d0f3a4463
zf6d664bf8c31e0751fba0110b41dd419d37ff323b6d672d4de75b16eb1d1b69474b84af6392507
z542192c9a97452b5f784b2821c08643133e1d7aae24c56d9171390b13e61e1654945dd8823e195
z63b503c602a61e9ae5a1a28b8a6b1a592f1e0e0a419b447444ce396df6bd44bd09ac726e21ba8e
z36bd54c9f38a4bfa6f269aadd7a4f6252fa1571c40177020b8f8601c2bdf66df7d3dfbc9cd8667
z1d625042250e94fd70e51bacb1acbd05c2996c21c2cebc4a6bbc663161202ca91db70f506de3df
zb752144cc76145c25cb30570e3e2eed99a47d76e9549537e276d54f50f61040b0e6ec6ec914b97
z704a288ccb3eb5fac97c2755686635041cef0265cf3af3af803c59dbe6876e2a3db927f122f20b
z5cbf82c49335a9c8af64ff159eb9334747f7a21517a1f98bba2227c2de5912117789ce8003f2be
zdff08ebc1e717aaadf40baa993d877b76849c0c8c202233393b7766c418816c18570b3074ba498
z5b3b14bf5bde7a114d600df6db0eebcf94f7cc74f95b958e55c58f91f6410426e1a592fd7aacf4
zc0547784c436cd0c8818dc7f0846e8f2fd6731ff6a01a971dc8a6523d662aa33fac6a197174db4
z440be01fb13f18f1fe912e3a7bc300cc365806618d2cc2218c7a1b6c8948e046e7710034b3df2a
zdad714b171bfde133c1432293ba690a1915e3ef03b8198de918a6e0733c44221cc999e0d36c6e4
zcfc333fe38e3ab1479ca42d28cc4da6a23bb2c3d0b2aa54eb8677d69cf9bddece5583d705b2b9e
z17fe1e94483b7f09f43d8957a094ee035d038511a3ef88b2992f7f98592fd6c7f7f3c2a85bbbd9
zbb48bf99ec72c0188445506c5c7cc866c4828fcc33d405ec18865c75c1a3c96a7c1719c6587a5d
z8363f94979917cd8ea1a28809164c1bf6a8ba8453f65a7607f373415047fa52b5cdbcdfbd3a441
ze7fdf206f5405d4a76350c0e9352d0736a0053d0d1d99e5df31bf37d3a990aae1e041c119dad13
z1851e41d0bc6b1761397dd8812a0bffce136acabc06d737acd08c051cd56f10c6f86b21669c3d4
zd7b96b0f7d3d81b8d0a50189ddbf27cdce300cc4244684aa9b1ab7481f53de785e54bb87676169
z197c65da995828412de4c527fadd43c9ad45ce57d1e743ddb9af5d39d35884ade6a6418b0186b8
z95d6960468bdbd9c6c541b661611a81db523313acd9646df3cf372fa08ccf671858ac42036c63c
z105ed6af3e6df8586ebf70f0c500e96af5a93c96d87ce108682715f20fad64fa867f5fcecefd51
zc6a079c917e6adba9ca2660c973f6501b3cb970096189d82d57b63280ad392bb41d73899a31490
zac1612576fee05bcbce65326a6e38a86f1bd2d8d1b32f90b883dde29f5368c021c13a376f1952b
zb01f9d919f3f977df2af628427302d674bef8d08941625a4b3375b8c9ac95b9ac59649ddb489d2
z621cd37d49e4ae37c4716d35b4bc1555335697f13eeb38370524dc4dd747bbc7910f7db5ba916e
z4e26eadd0ac8f8c39fb19293fbe94f7b6f5e0493f84c206a2ca731fcc948a598a1da3c6052e48e
z83c1cfb8289a6146c3955c795b1b4710f727297c2155b49e4bcc28b14316812d7ae351caefc62c
z97d067a2696a776cd478477ce4d9cfcc1bc1efbf4ffbde798fb5861a69554ad9967dffb7bce718
zde3c001057428653a7471a3fcbcf257b824ba0593846e3cf26030f9e20a5b1e58357865deaf256
z156483ca5583ca3b5ee84987577c002b6dd4e3701fca27edf9053a648d4e625b55d0b919c73ae7
z24e6393e97787921bbaac5c85e0bccf1a7b9feeceedb0f160207d529e4d980d20aef145359b2b3
zba0d78f68ee7736858f9109cd951343854cbd702fd498d1bce50057d7b39a9679041e299f84096
z106a28fd895a0b1f5c584583c613121a2e14de1c063af34263e02970ddccbb2b2645ed34a1b74b
z8a5ec7b504f0ee749d932e33be5ef2e3b3abe7229294ebe90f3b8dd0e3251f4ab63166b7b44de7
zd8d19707c89a7000c1551b3ffde32d4017e4a75339ea74c307366a3827a711369ab5327a9f7cc3
z9b1dbf709a990f4c99a794f03b871b9103045613c128fbee6db9a58b28cd17b3075c73476e81db
zeb1ab91a70168a30de94118dd958b987cd95def3f456fc0608901f9c70903e940c24617b2ebc72
zd816225315eb855bffcbf62185b45bbc0b6949bda3a3b12549444222af082bc1bfcb34c6b47b69
z33e79235641808b68287d0a155d2b9c18c299b8ddef040ba6c0bfa9963125a10452b1be88a2c65
z9555c1aa9f02f2423edf4cf0c2394d81eece31c60c1fc7c667400c75a668b06d8376c94855be04
z5d869c53985ab70392db3614e49e903e5f0458e396324799043930ae23443f91d797a006a686f8
zee54edfc61a20cfaa2e265f81aa8909823c7bcdaa1c71919c2c33e4d4fb1e95887d123ddd3c373
zfd775120a5bd5152a69a3bc4ff1454cd97722cf8c1127326ded7dc7ba0cf13b09e1af5d9f5681e
z7b893af64826a71abee28e7519038d15eaa948a77767c3342926ea2d3072e96f69a9d3ef074876
z77cdb300f81b3cd0b682f6b1082ae8434831f81d20058c2fca56b92c5a8305a88983f8c0f4c006
z826cfaa338a7b5070b6f6bde7c4845415829a9840c89fa26d872ad69724f3ed0ecb7d60a1946de
ze9887872d4fa8cf386028a1120f872e5d1f07fc5d00b99e5cb3ebd257b13a739b74a21e5d83d0b
z560b0f63be156e7db68f7d0ab745accae0bfe67e8ada0b4fae5b22bdd7dccdb12bd1b9a81cae57
zd80462cea7b8235e81aff67f678a4f762fc092e4878ffc9ba0f7948e5db2d5d5b8c0363c1ce15f
z4b4c7f3239d364ba571ce4d9ad88eefb2fdc32055ecc1edf78fc81751deb2b431ddca32757245e
z6f81ee0ea51cfe97773c3e021ad0dcb8bff4564ad029deec0cf099e6c829c310f1ceadd19edcd4
zc4d0bce42affcef3ea193eb1726ef1afb4de62692c2b8bbe3ef974692227614d87e976db9fc90f
z66e418a8ab0ec18600640ccc6288211684f3e772391009b474b075df28894c7d9c6939daa64e17
z7c7252716febfb2cb782098eb75c58ce60c46613a512c6a3c2ebf59865ff295564ed478e1423f2
ze542e01b3a8ce7ea48f62131dbd7489b540f9850122930888f81d1205575bb757032e7e20c2663
z7492b751f53f5b02e8c756dbf09b180ba174153c78148feb7d5c2a74b8a66ccdd567a02097e5c9
z8fe06e4bd289e3079a2fbdb035c86d52e7011e35fec7b91468d07254046bbc6eec4719b9a1b052
ze9da94302600a5c2d77c3fe3b1fe73b831fa22576762ea30c539968c56126deaec0bdcbc85d393
z551f884efb5bab51b75a617807ab84ab8df2686d09e3e1a9a838c49f696aba35b6391274384407
z9d1ade9997355177cbde6f7f858e26cb3be28385a9b38ae13f912f86f5ef28248e88c4aa373826
ze84183f634d805874293d6161db9614d67fad340eec53058effc3cbfb67e59803bb7af34809051
z1ada92c8ffdfa61ec6cd0c21f51f8978432b027b1bf1e6009cbfafa33f223f0d7761168d7e74cd
z2308fd9dfba4c0fd033cd5d7e878e416901db09cedc01dd2f0e09e4f1bccaed466c34e02341b4a
z1793ef61fd0b97376c5c520cfb0d9c3484a7d8a20bac2596fc8c6bc468933832ef3584c5090da8
z1efd712bade611a73a9b1068c3847e040fbd8d91832c654e733d48cebea345723bc9b26a8d1798
z2dc708c9243d1f7265d5eb383b70df92804c7a766fa08c2745ecb0944dcc5cf9ba3aa46bee8fc7
z233d001620b0538064f286b9aa2272fb013952cf344151a380b34afadca9e4a020ff4b0772dc8c
zf27ab269291ba180369d24dc365c735c30f8e932e5dccfca994f95e2d5fad30b0dbb28fbb9b1a5
za67b15b18bb84a5ffe09a450a8167f9a97c910c53e180a859b3066809d5a195a4fd7751c56cc4e
za095b149d893ea45ec9d2edb6f2afa266e17c5f96757dfffcfdab2395a7c1b17b250a7ed77e375
z82d96d2aaf48334b3b6c44bf737d98e08cb0f1f188e243d6c3aeb3aa251c460c7900efca4eef4f
z44c0c7804a3ecfda63291bf3111344509080139651ac9a0b4809975414523dc1eee20d15835bf1
z5bf4de70d775431157b3230277da86c4717233efc5d97a8308ef378fc7d10db7f09dbccdaa2d55
zba29a59d042f3ba0ec128fdbe2b08d2cffcc6d56e2a2748119725bb8f88a491a6c3969570f0bed
z570c4af0c6eb14c89d6f4b2e58f9bee2bc8738ba94f69aad663dfe62b48fe7cba339e0753f478f
z5acd0ae59c16f141f3fe03ada7657ed2d443738cd355c2f614f2531d593e8211fdcc0ad9e4fa52
za66ee2d29e08281f5e311122cc4507a705f9395c0a97f784772e4b7ee47b685573d7e8eb13eb0e
zd1018580558eaaa6b81def4de9bbd3e65e7a3730b6e707b74221e60b7c8edfd799cf25be5e7e27
zae52aad5f374185f9178a642629f69c09eb26b2777b9ba848d4fcf61aa6aaf4a046c25a03b01f1
z73aa213ce834c10babdcee099867f31b370d6870d787d40fc23293e2ce640a43da0968c4575c8a
zbeb76c2655108bc15b0b4054367a44dc4aa2791e6817692d3eecce4aef2c734b1cfebf8b2cd90a
zecbee5aea2fbadc6ade6918329c3f6e75142dbc8971b996534c1eee23cfd0767c84108fa872e1f
z0677bfbe6ee91ece3445ef10ba431519f71f2ad6b8dfda1427496bd2811a1bafb08657122eb3aa
z16bcb2129cff06a56cb5fcf4c794b572a5d8ffe99b0ec4beb46d45df1f8da1e354109fa45b7dc7
z6f2970f104a79462e255392befd1461b91a394891ca47d73b7e9f626596ebd42a1bd557f382852
zcec8d6ae2bd08ba75ac8a23661e60fbdfcc61cd322a2baa6974f859e94da3bdd0ed38a4c7a924f
z88bda1e7d5b73bdba1e1b9c32f1b23b8d23539ed461fef5cf51eb45c1fb770949d2f13da3f8971
z56a1f53b1840a0d2e93e6ace43926d68b6afca8d48d9ac02c7214492071d9156b2fb002f9540fb
z272b035b16970d14e1af36285836ca0c809ef0311700352fd23cf2d2dc0bf6383e1d1b78daced6
zf1b02da93c7b148bc9c95c414cf32992525135c6163b0c45bd252069a049bded89576c65863727
z90ee2e904949b338439a2fb89ad1f749bca7190991b345aadcb05d998a3893d3b40489e18cd8d3
z600e82f5978df73e8e4a3cc6a81c2a330c425c3967dc9582a2c7c1eda478ef22a379ecd696a3e8
z1d2d19374180f59a875f12b614a6eccdc4ecbad1a78228ea68741377b9cbbb60d894ed2157fb8a
z86d944fbfe12832300f5571cfb962de6e91d396f3b7dc8cf0bf19eb03b9607539b4feacf47eb2f
z6276dedba3ec6d5d8582827fdb68d8d1cb9024e905b889f6ef1786fa3c148b451eb9dd63a49b8f
zc881be1bee512dea79276deae6fb68a07ce7feb363262ae170efaba73125b235b9eee67fdd7d16
zacd5bc898a339f3eae57ad1b289113bbc49e571af619bcc155cd9dfae74e486a065a51cd42bec4
z7cfefe6dc4a0f442580019ec66e73aa61c114985dec74ddcfafebbc38485ae96e8b70590ff551b
z9d1d3a3e2788133bb8440fe87f30d39bcc2908e72a8ca3525c9a0374e25b5a61db206ba1fef200
z40ece978381401af15d14df7d360cba221ffa86da2f79fc2c3cea262de5c2fc2e637add804ac2b
z6456cb5bb637ad3e6f80a6bbcefb23bb66844aac4b552f2624daa532fba45c8b7bf6f827366604
zfc7286babec8b50a343338b430f78eb4a7b8f6b1ae48a862eb36a03498fa1c2d6ca97f8b3b1742
z49620af351d0d01204906b28cc78e3974809f44d7467a0a16a8d58c2bd70e612c4a1674f70d08d
z8fa82863172befbf4dad64330b6263822adf294555a44c5e66ada8cc60dd711e9a7558c3e08fa2
zc2583b302431ff5ba6a842033a06839f05f450283f5349a9be135c01e168a60515f982209794a5
z0c95a1c839046755c193e9dcfa7615914fed67d9cab802282cdb86ef5d2a480fa4f3f9355c8de1
z7feca75cefcf19d69cd1a244bc00d7f13e5a7e5e4b229e8db4d965b52c396a2502e780456f9a2f
z3559f10eb5287c0c4a94fff49ffb8018cbd71e589c95455dc41bd45b63603488316eae33a29476
zaca5a1cfb91114dbdbe8de1ef6f21f138836d3907651c17104d7261291240ad162168b55daf251
zcf63bfb446cd82c90579cba5b51fa60f462e86c6ce08a5a4bf2957a7e7e3df484020d2bee0230d
ze97c2bba82584a0fd95d3c797ddd1db06c83050dbb095889391459264c2a264dd8b1d17585fba1
ze000bf571faab681e934429c843f25f9a7ed163639b70d0fed9787c7358bb8bcaded403d6a7506
zc625d6bd2f7c40836e61f0f906170312a0691e3c5b849d83ab57c9695cc5865b369818dcd1cdde
z7eaa6787cab588cab00934546c1316a08f9c04920a7ab8e6b62d41dcf199048b2f97d3833bc5cc
z9de03ee414cafb851636912cf14482f22ac8a637b41f524fb9459c7c908b1fa4a6ce75cd1d20f2
z549b74da59c52e457e34b2b9ec9974e49ea2cd28925644068c4399dd743437ffcc919860238b94
zaa0dbcecde8996af3fdb1c1828e3357070e9415d48dbe0761d3d28f677b655d10859aefe8d4404
ze0e290ec58fcb110e03a0d37980a15798e9d82ad1826f6f273b9b9b670a3883b36c6b83e1d1331
ze6599b2efb835dcf6d4a2b6fdb24bd5276d70719f2e3490f2fa57e0aaee81485d85c6e23e0374c
z3193a0feb9d08ba4002ee3874cbc63b5bc7e2c909b0e076dc971a2ae9500891a3be5b9caca475c
z7517164b4584de6605fae93322b6c5d893ffceb1641bf234013f5ff3fd76db9fb29e1d3c23ac8b
za636b25d009740f6213f85358924aeb28b02201c3297daf63ca9165eaf027c78d4a73c4f1217ae
z02912febb03359bd25bbbadc479c5f24ccd5306ad2d3ad94a41921f3d29ce872f4c62452fa7d16
zbe0f5ab403e106253fbbe901b35da92ca9cfa7dc3b31bb667b5d579730a49598f6d7da4d05950d
z4fa070eca194567ddf368748cebca3e0de220acce2f864c8299d4ae0c8ea4f0d71839f8e0e006a
z615f712b314ef084d082a9d541082a2505f79530d42657c5de0a0e0f9881c2f6f7fda330e1756a
zb835e612b91afd5a86c2624c0976acb896b48a3e352473d8cd11ebbf6b92ef8ed84e0e22e889c6
zb6c62938b7e92d6ee42c03b7e12c16d668bc5bc7c6c70add78fc24c79e701a23906ea1b78c6179
zfce425a560d642df03cb931c7cef9b073fa33fc0c05717733a24cb85c790fe3f8161db4a5a0307
z226d7c4ec8ffa8c1dbb2493ffa30bc1b5b938baa66d2d9dad8ee27156163768c49db297e571497
z16776a787f600b8496accfb73819bedeb190a5ebbfc9e3ffdc3295dfa809c481dc72214f84453c
z742241ab9a019b627d3d8808186c6b56990cc0d995022634be5ed09b279d6e1a1f484f340b4e0d
zb513c24e89bf6efb73bd075982249d61a015b5d0afeed030ddc962ae26d357a1a8bb520cd17c1b
z762bcb269853f9e6af086bfde06af0b3f09f2b8170ed60b34bb7c98f98a77b815a512952d47783
zd7f948a93299e7b0ff5b6cd1ecdccaffbadb7a5b71074cc0671bebec654d7c7e6f9236f7a9b36d
z17586113643aef4537914c35d6d511a4f41c566c941a4e3e2ae449dcf00888b19f4bda31577100
z41712ee0de8f85591194c23a22191728962ced3a7a930d976111f9a716164335011f5e96b1b10e
z3cffe02a5bd29ca5a64c14c1c7d23485f3ee59d9c3431069c2ca096335bb14a45983e7e6e14f28
z6c8b620cd3321311bb0cb8ea94e54338425a8bf9058d2d066ff496b86f088428114db3b4bee485
z8e3161a57c828933697c4672820fa1c6e2aa81f67ab7f173afe923bf92612478e31ff4ec8ea1b1
z421f367a272f98b36a804c07e978eb632d3b3d46489e0dd0dc5341e53688283cdf73b9a9f23fa0
z9ab573a2411357655ec0cecfaf6ebae577d96df94072a3926e7f5ed8b203099215e54a5dd2c580
zd19be2c4ac41a74f953711b6a5e71bbfbf1a91a286a552a42623009585ce9ab59c897536d6e934
ze855e5e1beda870cf7c07f0ec8f3af326963550a4e54c214eb42ce040aa605311b5e25d8cacd4f
z7942be9b475eca4cbdbbe7dc2333f7e2de7afa6fe0559fdcfbc49798fb44b302294a4dd76de3df
z1bd982e4095e444aca5ff4579bf81e06d38a264b3409b034aebcdcf6a99b1d75066ec5b294036d
z7fbce3b3321f10bbbcb0df2ca0acebf722ad7a3dad5bd9c45887173396868a4f8d4c524e8d8e5e
z1d8a355939fe2626438dde3ebde1bdf5216edc3465cb4e91c25263d57203b83b59b5f2ba51c5de
z586a855d19adc14c68d1f1fa75e10e877925d7104de558dc3fcfcf1479d9505448d20b0193732f
z9de42561393ba35177cff2de53e0454432e643f4f468dafe284340552ff9423d2ba69394ab7c55
ze43c013601f1eb6ff9147b240a3aee05020f2b5880243e50286b52e404e7fc0b4b8aa2efcf76ea
z9625333aaa1d2201128042e928b3b88d33d59baccc2c4602a05c57625a9889fd12eeaf942c685f
z4f00935154ace94d02ac3579ae52f8ebca0ab6653875361337e9732998505bbf89d06815a8856e
z603f58042bb0518b0506519ded8f795c13bd4c38202217b63111256b5d51607944d3bd83a46c25
z0d91830b77980e9dd7426d9f727b47e907f3490deba82fc9f54302041b1e423efbccdf92d8be63
z1f1e007e3533b745f61918c76c5fe1972391cf4d480c6b40ae9a8ad46d4b5cadd71d7a074c715d
ze997720a2a79fb0a9831dce328cb81318e190989c5d3c96e0fa87de66e58871bcb227e953f7b2d
z236f0d1ab30e7645dd1c34ffff5401499e5d777ec3d5b06b3c5ab5c73a18f0c32bd439f46e7fbb
z0d353d12794fcea9a0085b234c102cfaa4394ba0687c28f070ec9807a4bb0ad8e12a6dbb5d22ba
z16f86770cefa337fb3e8f65e7a14d2a78ef1286d46a678c34d3475807f9ce8f9744c3a5ab1913e
z9eed97a0edad52d0fe8ed01889fd24c9d559f676577eb9955506010ba8e2261a43e4229eda6e0e
z6d7db8c1cdba106c2e032cb7ce898e7bda86f6549b22d4ddfdb5493acd463647954fbacebc3e83
z3f32a43451c3a469ce100791c3cc213cef585799e1ab97c017813cf2273ea732c8b6dd8aded2dd
z896271db933e1233d2fc3ed36e0a4a8ce3a1a249aab778a4ddd28cb426d005dea29e7f521039ea
ze03c280efc54e2df7734bf56202d132ee401e8049ce8aa33a4bf7873ba6d2d4ec8accc1c52ab67
zaf1d8333da9f98c2d1c71b3a599fa41a5002364d1c37d7fc49e72e1c1b0297dd6fe1b86739946c
z8ca33131f959f809ac29e31791a347f88dbbed261d839b136f88cf7fd83bd0e5a33a71f47604ed
za95cb5cbcc22eb7faee386af0ff6f69f788b5de75dd58bc5c57c288f5d48a1e69f833b55fae5ee
z040a2ba5f3b9ec30241a59d11b97155ec635ec6c791eb37247857e91874edfcd6df40e43c89e51
z782ce802ded5a2bd2c144ff242a0b251a21fafe101738ab6e918460535b2d5f3c81df4f1ab585a
z9b0bf26fde008f208649520df3971f3efd9b541c06cc256570b69e89ef77a7393c5642a1d09e30
zad0fb92a778c705cf2c981bc732055fde7b6282dfa04c780fa5b6ae0fd4c2392be34a2ef46b130
z4988d5384bb49e4513702211ac0afc5b5aa405fc6093e5a7d7dc9d660be8b02eecb28ca9e90b0b
z38131d11b8c8c5f42a0d229feb93820d97c470a565f0fdb710bba9a04d14eba2d6ae6a297201e3
zd8451cca0dccaca211bf64bcfa998a06b17ab576d700cc049bac11e7ac091ae78ee3c95fb8357d
z1512060644853b65cd06c86265da29061117c06d4db3f6baccda1944247545e275170093933bac
z09ad7a8178771618ca6677c0155fd5853f6b31d6c6ed920363641273f4852855c08942e284065f
z91291fdd67e41e0db97e65e45c2fb19c84c607e3d7adb4cb0fd97ae5b3bf1b2193fdb921555d87
z090e0c0a2618c05b704d3392da5294291983bfcee348a8e2c236df0ffa5d12f958903c9970764b
z14c225bda4dc08b35039fe260e32ca19d56738f2b9ea6d8a9d4b5c986615bd935d8985375fe5b6
z642a717ad4ce53320790aa0f1fb71cebbaac387c0de55918d1aadcebac9e8b57a826d8a870db71
z6f82c855aaad834a411e9e963f70be9c063b73cde1ae5e0b260d43c6dc699aefb4391f252d47fa
z850396158780be1fab7f12316a1f27d90c373e5c5083504a4624fef673fb3ebc09455674e0aa68
zeb16a5bbada56d8c6439ac7a0bdb3898df89f1188cc5bba14b9806ef06078dabbbf34a3ef84962
z34c21b191824973ed61334de014c3c814e80cf179ee4d41621cacb88c9f275ef8403ad4db3946d
zf6892ee02ce1dcfba219b27090edd56ed05121b72218ad6f67c12fc2db31888332b671b9adf769
zbf2b6b841ab2fa1954eeb19d6696cabe29e56e4c8d6946961fe170d9940e7ba87ca780fa64930f
z8505534eeaba0e4e8cfdd5b579bf794c2bde58d008d1a7cc3b226ff216db67c5053dc2274a0cdd
z2965598baa4056486146acc8f2d437cdb01950700d120ecabab2ab85741740f8962da4fc35fe82
z05f2790504767f0cde65bf97f7d80e2d7a3a35ffffdd6e0e0f252e5eac82f1cac5475c23490031
z095f42839c46530586f884193ca620de31cf44bfb0c7621e13bc7ab006473574cb64818cb402ea
zd238ca09e319554cededf1a0c13b694742e9865c85a2b277023584247cd3b92572c3cc44dd8782
zaed5b3e00c3410ba32273308263b79e0c3b586f9680a6e72c8cc540d3ce9450881ae301f28eb2d
z97113e7b53142463d4438e1ce0abf85d37649d143bac7c25f115830c04b498661c8c6aff9b216f
z345a09fd8196f54e3340f5dfe3f477980e32850788cc2b091705d52e24add316109fda695c7d56
zb2abe90c7b31860192fd7b9e197bfd06190a21d80e25d8018c1e91227481363f3354a09139221f
ze7cbf5e8b80681e2170fba7d96f8e10498c6765eb2f82f835175cc4938a03ff3633bcccbe819fa
z68b7e71cdfb3b7fd34e2db35eaad42f180e5ef1824b9395aeffb5684e3d277946944c409de154d
zf90d3b3e795da99cc987589b31e07b826a21782c5244d0bba36361422538997eda9538a1aa5f78
z9fcea97f87587015f90ac893545f941df7328e18ed1db369ea9836c9c751f8f693774a4238a392
z3690191dd39b114838828cd592d5fc9ccda491350430855b2f90e79bc03163be81efcdf1eef775
ze2d2794882062d31574f5cfb52c07065c38797cc42c8605bad6ab1e4409e035b38bba3e484c10a
za991844f3d5f4c10d9e6bb441b496259331249f057e8c8b18ecba8d4c2a9a9ea60d37e6fcd2d0d
z629c81aeabaadab39fb630277196613f1ca067446ab2a27805e1215d5956c38870c15c877ce3aa
ze8cde1c899f712225d3bcc62b678fc41cc3350396871d1ff51e4da10ec47d14607f6a63e329844
za06bdfb3282a3675e77ec78d4444559190cd6105560fa3140431c83391a3d5be65e1d0f3780512
z682bbedfb8061f07e75b10a6fb72edfa86cd309fa199a464065a7850e289dd7a7d9175d218dceb
za9ff05a6ae885c31858760b60c3cc220994195c7f5b8e049517648eea331440116b5421fb28765
zc8e7da5d0e24d3c9c0c3fbb8d8b1f8be0996d6f3ed22afa8f38d3b323ca11601a8c3426df37a28
z5aa2a24b032295c78424e0f6a18e34dae9e9406fa0e9b201ec0b96da7dafc89fb659dd8f30cf0f
zeeedced3fcec7360346167e3522014d442e6ccbe9e7b4f4a38c504bef15869466ba077be27b41c
z7fca496978d6256395d71b851f911fe47c3ede59905eb61906b8462d2f7a7804ffddb542742567
za7a8bbc1422dbf511c82f7686e213c3e3c2640647745a9c1a3009154aa55c88fdec12734e109a1
z5379c479ade5d19fb823f8c8c17a40e1159106be0a83c3b465a1d110183b9e7ffcdfcf7cb0d09b
z773b6edcba15a2eb21401dd3de83eb3fcded9dcd1ffdce4e276832018e90e6ef726cc45198b876
z2d7e50c03a7925d6eb58198aa7ece7ecd5b5667f80bdcbcb87bbea138f657e729ecae0bec0d9a9
z361f3a80aa209a350e2fc87980c9aec00787bd87e3f368e89b79925551be949b5de7c5595d28a2
z10b759426d1769033f73ef37062d502b16f6b6cacc2bfbf9d4c343dcf7e83e151eae53c491fd96
zed716282752dea65fa73a07dc037667b40d9e689667850df6c08d68d96e32f8f11659a1f31b3f7
z555edd20bdecdfbe41b98be191272ca9725f964a95d618c991f36168c689e28a8e46e55350508c
za1e81c21c408c68238784415afa39194fbe08da2ce54db58828d8f8e8926c21ec8bb80f6d18d87
z31cb886a47bc060d7704d7e864e832724f8ec444aa7b00d6d061878623c8a3a784f44abc504149
z750c513669b5c78ea01f350a7fb410e6cc9e1178c89507b41e6a872759f8e0a7726674431754ef
z0b0d5c3b1bdb1e93c636d9d7a166b1db425c787c27eca42a9c981ac40ca84eda2e409e7b0dbfa2
z79d2785100fbd0c8c12b8a58764ba2719961fce8bd7db7743217575d8312aba1923dbe8e3552e9
z312aa754887cb6cb0922b0a3ce6d8f605c85c168f86d154ca3951cc19309effc0c592bd3c695e6
zc0d8b9efc8dc80869718e19ba66298b594a2cb244a0345979c0cf076620bcfc6432f1481e15020
z5870569d060272932e49e929fcacc421964e4365fb5badf3595085526622561a181b1111738ff8
z8113b27e4719e45bc1fb8d61627f14ba2b0dac147cbb40f4cc710628db3c903bd64dd4be09df59
zab4379cffeb7b7ca3a1699a63d4f9384c0c813734dd4ab6edbfa72efccdc5e864569cb4104a728
ze875f061849e618aa05f280473977cb7159e6af4b82b710dca9337d3fb27a3a060e18989dd98a5
z70aaf247d1d1ac6226c9972942e183823187d8658e3e9e761e0eb8da8970698fa69bbd2db515dc
zad18f50af293774f5af5fcb86ef0093a1dfc61810dc1767cec2f92a465b3250cbc30e8f448c17f
zc9e843b837fc0d4acefd09e3c11bffbcef7bfb16520573b855a18d7529113d45f954af3ee86fcf
z7d614bf55e180d0f01becee452576e0514b690e504b9a377716d9f8b84d76389730c6e5844e7ce
z830fbcdb580052d623b86fedf40fd9e2e70b97f8d1a48d120ffaf9d930612c7c4d4a5a66f827f3
z69e688263993561132c30e8d049b10f5acdc983e354d8e1973225820e5aedcc8568267008de145
z9734edb6982ed1b25bc1abf0e727757094f11c29521b02841a51a9835da545f62c7d9a82d05214
z7a729b396f4efd3888a51b3b86c314bd4831b1781e9f3079e4f2774435bac3941f3fc172d5ef92
zd27c47f09f0a2b28554235ed355d0d7a7f983a460fc9aa5d6ca2f51b9894e1c22ab040827e8c45
zc4d40839ab17d4b5fe05994ec9edef6ecc83b744a80eb0262f022f2d17ea6688f852d933617360
ze146b60c0c6dc028a71d00a8169ce32fe72c56b157a88cf323e8625aa3fa9fb6ca8fb0cbb301db
z6bb5b2be8bdcf0583df8967b225d9e4817f98fa58519d23b181afed038fe8bfa841ee48c9a2e78
z77f93b3619293412a075d047d4409f2ef15af394fcd7fb0b87b888705a1dc63b3e42af1e2ef2d7
ze0f71b4743e946e6e52546206cb35add5994a5349877d8635fa73f65da48edc8921f07a14babf1
z116c819649c9680d772c6001782f607c1662c3be1b3d59a554df767d401e146bf8c7b5f913397a
zb5a4fa1e0d443f1a73779c86421269762aef213ba3c3c557960b514993255363a6bdb5f44566be
zf922e8d771a415160809a7c03315c9ca60183b9057ce890cf39032ae99b7235d5f27aef2f404f3
z55f61bc1e92688167efccf3229d5ee4b3f3ac83de354d09fda0262645b71bc52e41e8f708bf671
z37f42beca1f7e7aa790fff403dba438f5b05ed9dca82591b4efc0dfa68bc449e0ca5d02239e740
zda54cdb50c1d1e8b062e3ea4540f43841d3139db467fe6f19b70463987ba4bb1ce9bc6d6df4e46
z84060dd602cd2611e7c9e27aac8505c9bc4c135cb3245de91b13d95e650a1ad6c37a364b87a788
zc36bb57e23c4058b7618b6a7cbb340bf6da4dc7577a96eb97b2bc9e560990e2054f5bcf036bf44
z6c11c7de60c8c63cf9e8f1ccdc6e8fef8bbaa2c5015a646d4336b8734a44af5ea6461357b9e4ec
z0faff575440e03e5d45ae208b4f759702d99f2c654542f5762a1339f2753b0b9d717d0f0642355
ze5c1b13719ebb03ed60d25268c611f9a8150cc3b58b4791ba4bbaa3420db40a3bc413ff1d1cd0c
ze776dc57119f15a372992616dfd84ecb003150461497f1c54e6d5ccf8bfc195c547b735e9a04e8
z2aad7f4b62dba422f00896938af67a61747ce95cea7c41c8dd569ee2aa25726dde36bb27b70954
zefd1435c4a38e46901fd4c0247b3f9d5f6f4c1bf41c116f73a4315bed939d92b94c1888e4806ca
z1ad7112ad9391d2c0cfb0135fa10389535171e19716ff791636ea3510dde869d15259a422565f7
z2dc5a515c6d27c03a4a19bcb8cdc079762256920a6d6a1993e9ba3e58e67fa8d44e4f1b88599a4
z55b0d07af81ac0e3906ac181b9f2e369636f37245b04667a7fe9ee2ba48f2defda1b23f9bc3230
zdc86dfe79453880b2c8a22d1f688fad309b9a8a2f641325bf7b2754b5f45d91740eed4fe0d9575
z38611102a78a8515882109acba776403c72808e34b8db9012b14b2f914bdadb82beefd26fde897
z24e1e7559df6fc3ccc3f0b8a59e37fb805b31ae3e8d3f216f88e6687a14c6eb6aa1d639196e834
z49a1dc3141b2ca9794e3e6cb264b5d54a76fa32319c98e2cad3fe5b7eef2701fe7ac8b60e9820e
z3f5488b7bf7f548d6631cdeee4c355d0676ef92fc08ec9e20f1ba8dc4468c2d63cb89ffa178f1a
zecfcd52142db37399834115e7cf1385335223bfdb87f4233e6c35e3076cebc6a664ced789147a9
zc27736aa60d5dce62c1bc9bb2e2515ce98546cff2e92e318332dcf93c44428d7724e2b02103fb2
z4d9fd266cfd4718e18808143e928feff8403016a769bcd6c26f9de0283ce569a5198ed7209e8a2
z3f1376e375115f919093f88de6723fd7a1aa14e414cf8ddc96485ac584ac86f5bc8d83129e2336
z8bf59153beeda374f754bbe3d744f570467cbee4b5b595e6e0013810b6c65a5d53167e0a94647c
z1a646db4b0604333a1cca90deceec1de8c96920b12f9de4182f8dfcf7232ad5e65f4accfa18acd
z4fe0ba662ea5159d5e234017f5ef9605572c8d5602ee338c4a52b6985d63be5775849f8d8a851c
z924904c077936828747a50a2a943b0fc35cf3acdff63e26ac62d61e7ce68b423afff9e590edd1f
z7b2293928ef44af6ad8916d75b57c609ff2d16f6a84d0f1da401c3032de67da52d1ea1e0795d71
z53a458fcac89dc64f4d38faf0c536aa2764cb64de78c922bc9045afcbb29764c7bf357a565387a
z888c106c841cda7bbef842987231c6cbb42c37b2de5ddc910b9b5da2a27edc4a0c625f115eed23
z1e578c64f242e0c48c7db43efbbec17c81960749d3ab744bc1aaf83c3bc5369f55bb3ad4c794d8
zb28eb172bb5b4efcd5c7221a8f3fe3ece83d431b7201e9fe62a8cca6ef6f7a08d4680df2b7face
z999d788079c5e072718440735845cf844f320d4099b128e5adc81853a40d2f9fa4fc06e632bf81
z260f087cab8563fd08fd0e931b9b6b9a89d810620e29e9cbae37a6fee171411c4ce392898c0fc4
zf21f83e9d6dcbddf3019957cafe560a71aa54e16cf4669a60cd64364e8c5ed429f06d6600a4a9c
za486cce5ae3d73555dd076604bf8abcdb9b95ef20be5496c9fb50e3d09bd626c69a6cfc2c6348d
zafde4e5446fa09d3e665eabefe5da2511b242e3bc4746565b8dc96a8247d0c3c83aa0f4952adde
z5a6d4225d6629cc9fb24f4efe83fd5511454f812ce0f54ac1d709c1aa449a037b3a9ec934e7074
z07fcbbe73d1ae24dcdc320b6e31f8b371bfc9e2cf33c6d919908d63b33b9961fae077981731d6d
zaca2f1c1b25b3cb8f5ca4b8a6b1b1575ea54f658bfbab53b73771e2933afda07a1f3673179d1b2
z1e38cd50e19a2a0a42c3fd37dd7e983df2db539eea7c93ed271798aa9b3921cf9689a82096d029
zf83427710f90605b73f30b3903194a7d2e9a4e6f126f70cf02c91aa84421d698b1a2a01989ff3d
zaca42267a28773bc87c24c30be9b5cd2a28a39add163d088ec4f2df8b866c097532e192d7181f3
zd188debcb5532064236d358b9018d03f95a51bede8ebb99117da6ace059b69729f9d6cef3a91eb
z331eac52860e93695041f911a4a2663ecad908586f610ea3669a0fba0bf5b068a02c3ac13ef514
z46be04b9eeafe28e9832faebcc76e400c6694386e372b8bd5345b97a52fc8924460afde1ef0f7a
z95b1482619fe40a59fe1b541a4cf9ef5957546e238015711f8488d111497f593aafb8496035d25
z0427bcba44bd1c790543acff4c59d4ffdfa2c4d42f7c1da8f08c8b94880735707d7740268cd100
zf6f6581252f527f2bbca13ec570c0b1767ddf32bacab4ceada8e63c6946e423b26c7191e753ffd
z3842f0230587328d73b3e643131cb740f17dc19808474a03f015ac6db315b697f698ff2ecafc34
z211c9b3e2bde2f26da2e04b583a9826b62a3eeb3985c2ccf22179f2039c6a3be8f147e01b77ac7
zd96f2c39d1a561448f5cf53423a444cc312ca03e82c3f00596c8c185cbaa6faee45581071ecc17
z5475be150970ac2641f40a434848d9c3b8832c2f4dad934fb8a23fd8765fe5d61e11efaffb915f
z8280c86b8929bc96fd968d140f1370996afb4f4501385d3acbbf92b1ca6d62822b17c0b814c5b8
zb8bfd4a65004b950a301a7ec1431ff42a97b6bae490932668d5e04ef1608ef73007493baca8c3a
z963e625e6354adeaea766e104082439972ab1765bfdc8eed56b3e0bc48874039202e645e165730
z069548c7df07b7d08ce03e4593b10a811aa59950f7f01e4359ce302c894061cb207b3e15fb4c31
zd18c3b5587c727406a938ff5dade9db8a987d01ffb05fe64d0ffadc24fa9bd1f77629377b26b50
z6435068df4f367c004df4cbab528245cacf114ef0e7a8de3d6413de453226a743c7dca6845e8b3
z235fa0f20effa2d313ace24526c29571b5540bbaf104d87bf9c12a4d752cfd860b7c19b3e5e337
z77d2bd5cbe8e27f4df276607e31fbf78832d536d41bbb672d55589aaf353b65c5d8e7a010e80e7
zb32c298afa8331f95702d20e0d02dc6529f68ba64cccf33186370ba8e9ad7f3a7c320763937161
z1a298f2067856b1cff95e39bf0a2a3eeaa0b079fa4a5349fd61bc9ff473ba50341c93c47ca76a5
z1993091c96426acce4281ddb81ee65386b08226ff6204eb3930cc87b78c0f9a6c346b4229713ec
z0b008a0bd40a71b5c93c4b844ff2adba6d3c63f7fbf5925b1acfd8767670d89af10195e3258b43
z179d6147456010fd73c50fcc40a6e6f66ac9943e9fedfa980df45431b83f4331f3c84d2abf310c
z14dbb3dc3c40d0a4551ac25120c648d655019e1da2cd2cdf3a093d17567147b504e62af95f6ce3
z20e281b66a6e902530125ee96a5001e58883232b21f2939a1a63583fe5044b306871a7f5300212
z0c2f7e51c760e7d9eb2cdf829f7d74081bc7975307c8b193ca655a471724e37fb8666515144b65
z76702683b230ebacd09611a745897fb0aad23ea71c296ba1b875f2ea9ad9c4eb050e4cc81eba38
zfaa8dc04cd90dabe6eceec760e92ae90833648493fdac88a2569a96b11e024e570f459123978ea
z8fe980226da64b055376fc7d41a40f03edffda3ee7d93ac6adf061d971a179be026341041ccbc2
zb26e1e4350d954c7aa2b49985f3454bdb96881565a85746683343195c3fa5ac2f6413eb945eb91
z89c149e7fa8ff2db54687106a32828d55f27ff1040238a72f325ede15e643742ae8137a428b0c4
z8606492fff409b0aa4e95b99be9227e388ff6f9ee6da78056842f683712f725b06e89147f3e9e4
zaae6bda08c9060711774c0ef36edd971b43e85a63fb45b19e7e292b897b72cefbece93489a8811
za473a291197adb0430cdda66107b09d0aedcaf48910e06924814bac4045062f132359df5eca48c
z0624143e30fb2aba931e1c2c87fbf5776ed22620a85ac4c73bf0a517e8bfd19e1b87a67578e72c
z43e52ecd701c359ed5404e6f2eb4a2cfee85a0349d68e73fad5d68c05f163d40d3fdcbbb87b2e9
zef84772a8a0b16692fe11029fccedeefe180140cb0f7f8e82f6ef53a5e938f139f9d470cc06466
zfb7a03ff05596f5527055488af31b80e6e0bb3ca4a8d4d2d383fb0d92a9d7d3c2679f7252547a4
z1fd5c218c1127bcee642de4f3eb3a28557ac1967a4c18c930fac1131594ecc1550b1bc39f3cd16
z4309750e873ae9d80c411d2df725649fb47260fcd54c0505f27c9a2d5bd8a56edb236fc742c24a
zf26b51982b311b443fdbd408a90fd8cb28994963772659e74d0e2ed3e6ab4bc275055ed8251c13
z51db16094eb1f9a29fda3aaf2603580cad69f8b736ceac3a44fa20f90de33b713d809044293167
zc21a5b9a0b2b6bdfa2857bfa5c12d66ff9427815765169159f74c13f9f6d1922266c67a062deb8
z00b8a35d717230567718fdb108385a484699c767142e6c4d51d93b901999d5697f6cbf8a1e685a
z8eb9c19b36d1a868e748acb6f3b2a304817898295ae50226f2a820e7e091f35becac4388972f68
z1d6f27dec4766f91a3752bd5b5f14c9b06c46e555e08f189c164c8989bb9756bda781125cce6f8
zfe3daa83b86dde9c42d7f7c11114be2026abf4bfcca86c53f7775dbaa7b3dd444c4f23a6f013f6
z5270e85b211ea223a11272ed18f5bab03a46d437ca2fe263b17d8b739ee90c911a0d9f897886cb
zca4438400759f3bc0ac30941c99854017656697938747c3099d7785994b01d8bad59a1bff853d4
zccf647d548f69affba5f1436790290dc766dcbb5c7e001fafcfd50efb5aef6afdbccf456ed3a07
za92ec369664157cc8bbdc4391ed7d2ea43ecc426ac1fe4126a0df9bb11b7386b0feba44d6b34a0
zc4cf05ae9d252dd271eb46d7d5e47502312982d6f48ae7398309115bc1e33ed0bb7a613f7ad645
zdd7047108cb74b37547d0007d01d33b683c034e6eabfd073af5e680a8ea2dadb6a52d1bf96f608
zaa9be61b0ce43a9d4b7d2b1f8b6980c18a0f7d66044f0476fd77c3a3158d06a8dba4ee93d531b1
z6f627f4eb48c807faa2dddf432ec2d93040846dcc5d04d9930e3ef1f7fd38b399901146b2ad2e0
z5405eaab63217737567cdafc33797fc456d644530dbff3dcf4e0ee3aadcfc5108cf0abf88b4bb0
z7296ea91f3d20b429cfce3bbe20cdd18d0e3b371488fb39a2d9dd848f7c8caccb233b53662026e
zd524ec50a15487786da14805150da188d90871843a215b7fa18de477af96225d608d4580c1e2b2
z9800670a91268a8895203542488238e6ed78c1bf5d2d733066cdc9529a1c3eafd1b3a9ecdf426b
zbc1791c824103fb2403e9fd11a8f36cb67fd6cb548f18e5d091f8c98da11b1ee6caaca03f03dc9
z3178ae08b0ee04db1cb3641ec0efbd42012e0516d56870305498ce312c22263c5212a12333e09e
z24e90fb5da8f583821e4743f818d471f82dd162fc2298e018c0f9df1995d7ab54ea168eaae8303
z811f8074a5329d3718bdaafe2f85fcc064e04b515b70c47bd493a7b338435abbb113bace676ffe
za646e06b9c81adcdef186b620c13f0da1656482221a4892c4e822d6aff777963d4b8f3f5f376fb
ze569800f8f7b4275b0fe464bd2a1aea49f861f73c1d4790754fa9a9814732e9d4b7dd4a3cb701f
z75ff5e1a89f3acb3d21240c63ca2e9e2aaa5c41119f91e0cd5203370fd294c5205931eb60ffb1c
z9e228267501ccc6372a1bb279038e42f537bfbafb00c3ecfcc103eeefad90009295593ee2fe53e
zbcb069fd7586d2098d4ed1188a42b0634fc09700730c476d9eb037680f2e0d29095b3390798271
z6e5ee408b62248cee8d5dd2913f66d34420f07e99446aee9dab6d9d68ce079db41ffecca2a7641
z34fa4054e46340046ee93e304513f67090a8d19496e8a7c1a039bce54f691b190d2c79395ca991
zfae38239b8ede64289ec6cb719f0b918683b6fd062628aa60c541d902dd2fde817190d20c718a5
z9fcb309f6cf38832f0dd42edcfb96787eebd68b05a0dac470d0f3e5dc568107f364fa7d2febafd
zc442544d0c488be5bcd6f17015ae0b32e0f1705aebb3fc0b1bf72634bd22c74f6f3e0103753574
zb6d92c70f9cec693fc7673efa71c39cba5518f82646610f2dca5debba7b040534f9bef8d3e5091
zd631ce592b9bb2ac2d6aadd55e781e2a10025a8c950f41885b2bad06acea15bf5ce83a74462ad7
z44dd0e261c9fca82304c827238554887bfb18beb18aedab3083ead51a65d05a3546a8d3f3c1823
z856656da0592edbdee694b76dda91b30506585781ffa426d5bb9ceffc94f7d56af6e14def701a3
z2a31ae2ecb1b8c684903d8810b65840e395480738496b9d96d3c68655008c48bfb2f0523564601
zbcd62a4fe4bbbcc32600e509d40ce9e9ea7b26c92a0a0b637605d6af3cd04341cc4ba4ab9a507d
z243b5d346a8f17bf3b0264318e84ef20fe98a7f1dcdb95e15d246bc694e6f59db00232151a2a07
z6a58ca92f402af3b806444cf959a95daa2b869f1d55aa4cd5f49bc04ca50f0c29f35c47f05698d
zfc4a1a877c14b8afbdd6dc89ba90d9c2c178d085b4e1bbfcb39d6d91a28e65108f66738a9ffc60
z6f9463fa29d896f933f2515bc070a180390bc114f77a22a0f604fde4482b78f135fa610f72fb01
z556af5432b2a3e9502ffe0c64d46f77761f2c571f6e12170748f0e71644acb95a75140b393a478
zf2102a23544ba595849f3109675df8359cc785db703fc6f67bd01ef2045626cdfb9ab5ae663d27
z87fdff35b06d4bf850a5eb8d873f9d03e425fb1cc36f90ab792c5fb7b6ae577b3855f6dbe1a867
zf7d76e0e26cd4c4c377b3370feee3b98b7b71d50967354dc8371c98c3297b4d51f56841a97286d
ze7fd31b3c7479a141f4567a66a0660639f5cce8fb0229fa03a376777cb7032b5f8b95517f52afa
z38ae50f03689abb7a9f623370e8328b075084e7c90b6d4bc872efb5deb231a99dec30edf9c4946
z0204f6e5a50966dbc582fe5704172537399612089464930087cca9c3ad06e5dd6dc6385477e480
z425353f636ddbd4c84b50b3ba2a9824d3829ed799d35423da6b80866db7f8881bd5b477d98cbac
zd993d42356adfd0327460e8c3fe962447b85e17bbf97f6a5ffa3f94f7f9dbca9fcf8fa938fd545
z23d569980bc88293b87a04f895b01e518a06713f7163255237e170e62e2e3c3b85aed8872c4409
zdccb9d08cffea845680b76367a0e7b2f3d057e2b02341698bd9f9118ec2c904b4054c739f02eef
z222a5a0ba5ac11102657790509a1f6a4c0e3a5b24eeeb7ace16e29d91f898a7bc2432c8d7c1e97
zab0dd2713da64781ceee1280edcc7fefe8640bcd932050989bd8bbe096d18747d945948b3848a3
z12c5b374bbffa06d69510f908102d015f92587a0ab280e50c40e36e1b4de31d263e8556c33524b
zb59b51f1f73548d0710fae52d0452434201fecdeba2e0eb73e1349f0b6b7e588fe652ee149449d
z6c0c8597fac57b52166c350d479c6e7cccd17c850c08faac5e2144133b1365624840ada79a1796
z246e5365831cb733fa41d6fe4ed81965f60fa83d88470aabd7e16ca9cf8833d4ae6efd137dbd5f
z8aae928c38ab473a5a6d548476114072dea876fc798d603ec8fa60e257c6d75b8d4e0fa3378c5e
zefbdc67aed1833250ea60428b97b3350945cd35e343cb51eaae2e2e29c4a16f0f49478231bee63
zf2c0fd6d079841fae1ead900c925b82df0e2221cda2e2fbc296b7a85a0b32bf4c6f13a76651608
zff311b91000f0d71298da17b9d407c721a7c8d120644a9534a1974fae7ee1bba5fd56176bf1fb3
zf4c3a2b0747fd351b49e3547beb66e937eef72dcc0788d0ff815236e21359e7d0442fa3b3ebab6
zebf5925daf063d2548506027d8345d7f9f5b215ecb98e72439617b6dac2c80c75e31ad50841f9b
zb82fa5805e72a7408095435a1baad33c0ebf10dced164d7b15d7a0520804b22f3b98cd9d23959c
z067a6219e2990874a661d1c86b290eb1643281f63580d8a91aaf0b32b7c1fba14d852fe583c7e9
z060cec00c2a22a83adaec1814601948c5cde3a06986b6574f607b3457d308208f4329958933bfb
z36404e66c0338f008f0f5ca2cb4f95978c1795a5001520afb7331e25e7539569be1475d5bb0945
zb243b9458ef6e651c0fb44cfe075098388ce01a6681957558a0700f01b6b1a5ebf69f1ec5e0fda
z0e37021e56d87407c01688e006e2e43479b3f5b7bb048fbfa1be95fd4822a7feea193a19da69b7
zb4122e7b809359e7a43ba9b453df80ce58e1545f204c3467334e71761458451dc24c350f13780f
zcaba5a1417ee1b5861efa2c4266cffd78676aec25291266caa2971c715d0f88adbbc17aedea2dd
z34da32eb67933ee5df7ddd41161642a234f3231e784178f472c34b231dfd972538de4df753e66b
z71836dbe58e25f19a10d3aa988ea80cc3cf38a72611f5ca8ca2d74f79f296a10d7183c6fb605db
zf4b2f4d551941f707fd9cb5bf2fba79afdfe07c47fb8f1d63ef88a0863ba13b6c9a43806fcfb9e
z574e574db26d98b11c22f9855a276321fd9b333294842227bd15ca5395dc61b264d0e6c24342b1
zde7669dbcdabc28f9cc634140074782c3b44f0984e5130c1a67919acf9fc49ea0920531126b5fb
z52874ff75abe9cc88b1b92f04adbb3234d06cbd122a3c1ed936443f5739e0b40cea20e15d8fb18
z077f4fcb7a7ec79e456da9299725de63e84de5989eee99a0d681c5c033d41a4d7e47ccfade823b
zc51650fe3112e80689ebc5f6fb42a5e22ccc4f464a8b89ca244c45eaac8b568dcb773c84d08087
ze17a7fb8c4953edef3fa7fb1ca76896269147f3f400ea19e148e41efbb3582e170025a4115900e
z997684f2116ff9aae06520e1467b59694f6b243c59154307951188c817a178b9e5b24eeaa18e15
z5c94b2e81c227e18a46c17887e55f9ea7b5a823bb815110bc1993219b404d1eda7781ff7b4206a
z378d6324f28802a1f5f186818e6c7d7816d1d9b4d14dc1929149db83677f00a188bb7eb9e8f0eb
zaa7078f5b175f37dda2c4f2d3b3c69fdf7a24fdc5d01a583f01dfc7cb214241f673a4b22b45a8a
ze2f3e8351cd48ce75239add7559628d2e6d17cf915572518fedbd5eab8cb1f5be3d06c5eea48ef
z11b0935c824affe6c04463dca2847b447c9feacdf436ad32fd512aee0ae0ecb5b31beb81857eec
z91d4d86e4dfd53995e2988ded4acc30e9ac5271e85dbc1ea30ad1cf727ccf2f87a06434e89107a
z712b6303fd047a9fe00c21409eecdeba5a875c1805af079cdc83868788e4a7528f76b2f97bf15a
z1bc14ed446d9a37d9397512627e43da1e3ad33f1912332d01b899fc3847c98cca307026720aa70
z1c4e1d5142247dac28ba5c00df573f84d9070a11204ff7ffac448f280b346a12d57b79ac0d9321
z787d318cfc85ab628de9505a26569c58cd802e88f9b58421eba82ac98b6ba30680dee9e0c7d71e
zdb0238a7e8b9da5bc035d77b3fa7f69b540607836e49e6d5b7784cd18dc1977dc1a174f1bddcc8
z07bcd31c3a6c4311df72a97c727bff4ac1ced964ae8cab4b78d8ced0c09c33dc10ea47f818c3d0
z4335a6d0eed0c00572be37c2be6c39a3861e852b8b568c6c25d579702900b3d12f534e15d893f6
z357908c3fc48b7223d2f3143fb437ccceb20cfa193ce1787fdfea8456e9b9c39271ca2e93332f8
zacb0d92eed3e16bda572019fa3335f11ce99ba5e72c9d191f929dd03a582fafcfa7b1070658645
zea5db4ecabf4a6cb329e12a7480c0f1e0d62411b1a3670e371690f8c44d560ef11b7800dfd9bda
z7e0e7bccbc0d7ee0355b69826b0deb9d057992812e559916181dc5477052a0273202dcb3165438
zd3b6435bb6495d2a2953b95c16d5f1e950b9b7326a77d38bbe8abca17146993045b45cd2b79e98
z1ae43cf5d23342f8902ecfbeddee68f6ff43b37f257048b4fa48af2d5f7f49604805711d4bd4c4
z929f9a173ec91babb88f92497e2fbea93655487cf7a6c3af98303ba9bf5ac6b453070cbe149262
zbcd535f607c5d76e06d2444b12f82bfa6f47068e9783bda2c54590a4ee11cb216fba4a47edb253
z17561e91fc83d7921dded74da9381252cb706107fe6b78eda72e615cd807baba6f33de864ea5ed
z58dbd4c3b99a00a2f8a721312ff9db0c985d61386ce13712bb280538b31fca0e7f3d13dfa639b2
zcf7a3a672745c82aa40f685575504d27808425486f016a35f42096b60ccc1a999130fb5912b328
ze86819a87d863675be6b3771efdc555917ac5523faa8325b3994d5d605052040add873815424ff
zd76c6cb1f4453cafa538f9f04a12b1b3bde097ede2a4bc1eb94ecf462bd5be951a40d537837b94
z1d5da5e7518d4dc55645c14bfdbdf6d51827000f3bd5a6420b99dd1b7f9967c808eca6959cbdd3
z34abdbb85d96957f6ef5122f9c11d3a9abad6a4726692589aa83028394687d05d48c41b2fd4c1e
z04ffff52f2d5aea18799ef78f13567b53fc3ed4804fe748d96d87df9007d07ef7bdb8b2283ee8f
z99d81575ec80a4a7372cb03a525ed95f076b25d3785daa75eb2c4bdc5b5333b5aabba4f40f7b12
zf50b427458a3996d8a889a4bd1932708258419a04c8687893fb3f975363b6ea1063098a5409274
zeaf4affb42b3985f93e4fcaeacaf41426cf48a01282212843ccd3477f5bbdcd0017eb8d22a832a
z2e5794270fa7f71979f556ee2e8fa32823ece5a67170c9a2ac43c8846ee399527e9e8c2d55ec0e
zfd5fba4c34eb883bf83e13a452d024f85dfc5bf04fc64d7eca96b0b0381b4b9aa53c038cbc6426
z726b44d6e6b658cfb26f53b33531834917e562c228533974aac13ac7766abfbc77b74f6e85f524
z604abc1eff53adb529673dc48d7408610ce07b62e0e06341cebb094e9012d5849a56dd5c4efbb0
zfa3c129a5f589b02e8a2aae5ae4e5d0fb0f308a0bef03d6aaaa6542e76b909bad1b17653149274
z367ed8930f5494cac0967bd08c66da932e392be59542943fdf193d67602cbf68d13affde1a22b1
z06a7df300e75f54d928146928be14f0b5c32444f948e2995d50ad4cc0588d6ccb9b521c8636b7e
zd38bcc7839e0f0ae393ecde0bee7192b4c941bd9e3e2d917364e88532ad3b6bb4055910c2a56ec
z6b862f35de8fc7e0d8052acec87f8adc2eea30c5e8cacf3abd6b1f52c221a0b99773e0fdf49145
z8b9abd788f16e1abd972aeec14d8b6a95bb0cafb99ec70d4b2adbfcd43920600aba697654341ee
za6ad871806e45e0372e47369a18d24eddef533922729746efb980b8dc89d2cf3e3859848fd387c
zdd17597ffcffc9dfd1d2d38678ef5d06ad82f3b80e6804dc530c3fd5ac14462f829ba8e225507b
z8fc682d7e9d55eba8f62f121818c36638ec7202ba2f9c92d629366796a87d2717ac50d46016a70
z40e5319c3976d997be1ccaad9689fc4026aa2364e6778845cf12378e1a23147b31c57bd936f850
zbb5d6c841ffb7007e22758af11ab26b6026f9d4f2f42bff073666ac50127a966a6cd8d9dccebf9
z5ec7360c4b8635660b69fe257f8fe5224a62e3670a1801f579dd4bb18df9237ee062d851bebacd
z05ce63857b3f3a761301c4376fbfc3655408c23000fd6a54f6d818211f3417ede59131afeeef69
z8b815076d0c6960bed4dd004d8981dcd919cf5d9f8198f6bf74b9bc7158be61ecd8e0823e678bd
z67a5c5fbadfec56a6e3d66366b8d3dfdf6598b457b700b41507c15ddedba9095267da41a8d6806
z609b2b332a35f5c584403ee17c9682f821d21c4c2e2b23abed80f0584900f2d57f2249a8d34140
z9104dec93e92f677dc9802c2412854c884ce1bbc32de5befdaff2bd13773728982a02726788598
za80605966c9e815cd174662da51c6c90f74aec8cf67a92b03a4df3af553296b8afbe4c8310be23
ze209be01d49fc1de4bd586f6dd17c85b7aebf3e1b9f647e7825acac6eb42d4861a3bb2bab08c19
z03ed96f2f46df1ad2830570e4ef10d43b770ba24b9166886ee9e12cc18d90cdcf6be047c5001a3
z8e05f5d9abfd5940879c48e4b3863282973e54bae94aee4b6f9a51ebf81c21f6d43279bc5c1086
zc94013ddeb7c385204dc8c7dcc85e01ea96abc024d0adad396dc11afeacaf18f8c1d2bcebd1eea
z84279ec9867bf486e4c5b1f5158b35633449c00dc079e3910fc252788fa2cbfe24ea40148bb1a0
z79f4c303f2b3119128f938f363281f7ea57f5566c5d07b864e6e46a048aadfae9fb39c59cbe14d
z77020440560b1985dbf8ca7c3e3ef6d658e760756741c9020a950f2d4a6cbb15c1fb0bf2cca25d
z2f87b2ef3b4960b6266bad875cdf57e32f31dfd0c0521c3ec579d29ff640cef7525e3585ed2131
zdb7221af8fb81134b0b02d8289d3cf93a1a2e3317aa9217386c2f0cc81ced8f54c16d6cd540932
zd40fb6e73ebdccf92590da442fd1f745d60d9da4073a0d39b2908a6c11abeb2abb2477d9753afe
z6d44ded48f249cbec9e6e0527c182f90895b2c551805a5c00417778e3e3dafbbd4580633a1c7d3
z657ed3c017c4250c77411ecbc1bb2917993ccf86d559f88f27695887d81a6ca3db8e641d3f153e
zd7b3772b5f35de9fe587b0238d21bd8ff846abd3779ae92deb106c8c882b555aa0645b54d096ea
zc02e66efdc594e86679d5fb502fa63394364fbe58b6076936e06c650ed63bf0b730a430f89a08c
z936c9b7a6eb75218d853d8be3586f37d6d07d3a70c9d64f30cdd1c2960df5f0ca0c2423c7e5bce
z29d4eb68a35a78bdbe521b4432e528718fd6ad4f1aa521edf332a40759096303766ee90a9eec90
z56396fa542098e8ebcf0981c5a87f9a7cbfa26397a7bb9c57f00d948474353b14bbe2f643251b7
za39fd3439d551630fad5863263ee46d0970c33f25616a9d906cb09115e538e8263d50c3172bcb4
zf61b141454fde59d7fbdb4359bb1ec67bd383e63a6d97f95a04046cfff880637cab913f6ac0a84
z1a5c8d3b85244b59bbc64c24b0ad197035977e2193ebe099afed3ab997587cfbef0464403c88e7
z66328bcb4d582ecdb1304fb394d3299d031fe2deed6b8f05065bcbb6db787230ad2535a84ea3d7
z39b4adfb287b313ea6ef941ab618e5a0e28ec884cdc3f5d99fb2a69189d16d10a10ba4eae16f4f
z6150095f20871ce4cbf58efe3ffe424eaa5d2aa4c93d9a871768eec737c6bfe50b04b2fcf12c44
zfb2ef011c20792446056ce653e82d9e03754edf064a8bf15bd88ed2b4505444e9df1d481d3ed8f
za733b763cdc2f00246ec0a9683d430e78898bc586b0c3feb3c547fcbdd6833b0d82d3d71c8f981
ze4567e81b7d9e5d09ae443f7d1ddf3fca4b83df89f40b603e4b6d26008e6a7f74a6e8eb4e6a229
zf55bc7172e79a4f7b188cd9ca8d53a88eefcf05bcd74522bae525d74dcb534d52f73283bfb2023
za2b09a3cd9e49d26caaff0aa5ce4d2d7746111b04a85eafc77cd3a8ffc94d21faa0a1b0f3c59cd
z301559360631f8e221bd96c309cdfe60a4b986981fa708d5cee5f509fa30083a88c83aca84829e
zd08c9b1e332683afe207e2493609b7553215dca0a43d061276cd2bf63b5de512b4a3040bcb1ab4
z5fddae587980411937c143eeacfe71f01e2c9895d8207f7b72b50f43554067d5692c2e83ae5154
ze1988bd831de84ded272f4ff937a3da9c7a7dd043d22aa97f5509aa254165e5b073ab4122b6e5f
z73789fb173b8cd4fe428953225203e0764af85a48b90249e4e40bbd1ac9f5c9872d64d1da9f567
z36229e375c7c6e5ad21cedcd5fe0d3c831d76710dfb173cdf81870fb8e803c7aa6d7694e5de005
ze3abfa8f118182b58e7a832fed1da8c74f724707b2ef1efa0347951c1096f327645fe1c94dd7a8
zb908b956f404434b3b7fdca0b6105e4932716d905938a2eeeadeebe63fc82e265ce2a128ebd498
zea87e854a3d6fbede792e9044936e7ca3d0886ae76c3192d11d3f8b0b53a2ce5eefa404ca327c5
zc4b05bd865b5dcf69c2c1402eaf9cf70fe8bbddd5664c9c695fff32a1f4d1ebf78ebca9ccd5a31
ze4b3cdfcf02be939c2ddd589381d9c7e01428aa5b25e10ccb7f2835c9aba1a7bf19a0ea92bfbe6
z901339e72ba08e9045f6964096876a494e134986ea9cef39ec4e68b19d74d58f3850664988e7aa
z6e52e98416d8206ff6e52c3d652b7207bba5711da0d80685fa1cd872dcae7754e34f21bc98c69e
z28f04e71ad29cdd46adc15f17142d70ddf20d2dbdff03720a7511864046cfd0b9b74ed34f5dc79
ze2083055f79b12ff3a69085d8df13be881e222dce47d98ae559ba632c0864440d0bff89f3fce0a
z148acc1a0f3390a0b5310ec70264fc57ab6db031862b335e7e6d38cf663affaf3d607fab96470e
z6cd46f126d117c378c545621f3b1566bc00b3ae8fa2fe499b24dce9957af20a6a9347c9057cb37
zd318cbcffd2836cb7a40c3b195c601fcc73d904437949ec1408a887982e628d9419c5d87b70de2
z3cdd2ed69691dbcbfdd3d22fb051a43912379619b760474cf14ff07f926e20c832bee790b26161
z034c3e604cf274baa066afdf13127fd636a486630d2072c8885d0e95395dfa07918b4f8f4f4a72
zded05fa8439cd21703acbaf177d94faf87ac6038d3d897c219cc493c143109de966fa5371ce061
z5c70238f1bd77d5145990835b77b563bc30c84545bdb4450a1ce54f03c0d486637cde28763b746
zf641dc5b9bf3ab6267437aacda2a4287f09b06ccd1210f33418b4e99e030a3955d630a761cffbb
zd5bbc9c87b40c61a759c88eeee7d4bac4955c1a62af647258829a445509fc2d4d62cad77703808
z71b453b3d410ae17cbb5b88f5ee26d993544f483c2f5dd710e9d346b5055af161c98d6193137c1
z108d2b87f50000d53cd62bdd0fc00ba04f9566a15bb10df92186255e8ca035fe744bf5921de56a
z5aa79bdf5c4f0356a8c7654fd030f8fc1d3d658bf84604abdbfce836f201a72cdc8e8cbdcfb5ba
z47220b0f1e95c7bdf5bab441c3a34de3618fc7af8bc7f92542db338d5593f9756c64e189fc3833
zcd09348430d0ea789051410572fef88e5f0e25c8f2e719fa96e7beb688a4d31e7ffa1809235c8e
z047d6d6e1ca91251b5dd32c928494811d2ac52cfb6198266eba56f14933e5865910375d764afbf
zb2ab8cebf232b35068480e1380df35d4f5a4f92c78738bf2e8ec648afdd9411113b00b6af43394
z651849a04e9c7178d540c4f882ee941a1625d5e9e64e069579cf46b34bbeb81c0337dc1fa8dc4c
za7a055cbfaefb2c3ffb5d956da8ad13a7e082a966ac0ccb46f4f26852039fa311f9b7231c91102
z3b32ae16b28b2692db21295287e48eb4ef2a7b3610904376838e2daef684129822c60457155fc1
ze9a7510ba4055d295be6eeb050afd1ee41680b193a6a21cdf9f1df9e69628733e7833054e9d433
za7643c2db4db14570d7961b492cc1ad3f22c6653bfe71c55567dfe04e8fd1fc2d5b77b15ba9303
z97f1e46dac8106bc2fa8c22f5c6bf7b49af2ff9ffd3f26be6d545b90151554222466cefa814f56
zef0d4973e9dd4103739de206a4f1ebb3db0ed977489e1dfec1818df3ba2d0c28327e1887ddedbc
z97742fb713b4b75ed999bc76b1557f69b8615222133bab6006daaa93fc72f20b69e68de55f4547
ze0dc49ea3d84fa1f4f83c369e03b87f132cc8f6637cccbdfe8db793c18fb18379d8e7a3da18931
zb72cd2f67bb98b99348c0846cd14da964177ecb161bdfcfe9757860f26babd13a78ae6b0090124
z3752ba81cabe74f6d20c6dbb6a37a4b8520cc2573c22cd6bf76875426df37690016b6ffc03fb73
z496138fd354c11d3dc5fd3ebc65e53de70564efdb660ccb3c68fbdc2bdfaeb7c89b2b8c1a39a49
zd36b481993dc0724b5f7f458f5326efc1aadcc0879c47365ac5ac1faf533c709916a940a3cba25
z841069c0707dd3c50f9c8b57e2ff5884cbd00e86d12246a43254eae670713f25d6491b5fa2e072
z9f008e9e8715531bb381b2b146dcca9b5e12b452eea2c28af54630b2eb4b1ab5b55c578ca731c7
z315d10e99e7e7c6317cc8155847dc4af43338d23fea417cec33e278e26177c9bcf37c400a7d633
z1857c786f606ac37f3c3b86748fb44001bd13a906d31ed1f716fcedc9a031f4c1e76c1b898976b
z56bfca409485067257db96705c8708d1eb14035aba2ffcef07702ea0ca54fc4e796d605ef89b2b
z4498c7f19d5ce81a4ffee744129ee00dfcf6225c6ebfc93a1c49532096f3a91df6ff7c898396e8
z9966c8a3ff90156557966efaf327f3d4d0818e43212fe36df6728370de677136484195a2b30dc8
zc3f63fe479de7ee0b5a45e3216204cccdc4afabf5e6650725ba2170e2c03e5adbe1c4b65e59242
z44c7d9178699c796267973d4f784be403d4f60ed442642777a055baf7fdf08ebd085cc0ae69792
z4c8e56684c7fbd0580c569f6ea0ec42d19ec0f9a34722ad51beb7087314744e3c8d1c5861f529c
zc072e1763da5fa8ccf82df8dbd17042262e08f893c35fe17c313770cfd00d4f225af4cf98b6c4d
z23278631bb5d5962551a0ddbf644b33e4d7e120ad1da7260add6d0d22bf67d8dee39e44aa4dbfb
z7ca2865d0d171606dbfa49e42f0e581da7ce7945bc4d42f0cf762e5e81341118857223f4896e16
z44e496c5fa3d0e74a879c06f90030092d7f79acb602408fb527224075464634651fbe8d86119b8
zf76a6792d7ef288a478357b494edd74c7d2941fa26547485e1ebf5ac62bb22a0b238f7abcab86c
z3fcfd5cf2950d36d9ce7e6740ba97aa5cba3fc183d3cb437d679290a7df32d287fde88d13f0575
z87aad62a3bd568f9d3f3f8babfcc8849f56fa062f01a7d61321a3088f54c3a64a59bdef213b035
z6b945d0b10fea9a1c679c547531355725cc3c65ae0ed09e701fea07a7afec625d8fda2bb0910c3
z066be3566be2a21ed295507bfb30b40d6276cfad08ea592aec7e71a029823c2900785223feb439
z1def2c30aceaef3f3671dac3da10cd02bce50a81410f200f7ac8475370a4582f35ec6d70f8ad6f
zda14b3a16822b4940b3bece7e0afc3c6ee523882edf966bd77071f9b212215afb8d0ca9f2ea32a
zba6f074eec3c866220c316f95a17e1e533f31217b82a7adce01ebf95ba683ec1832e13fcfe82d4
z0f58bd6a6a1094bd8ceb634c512a9fb1b07d888bb0e0d2a55aa2ecbed3d04743f56ff1f791b8e2
z271be0ec954ea0d97680ae17eab1be0b691f031299aa89605cc81fb3234004b72b3497b3a7580e
z690da0e050aaf3a13478b9b2bb95d947f9b38f51f320f86d1f4afeb77ae250dcaf273d6603ea17
z4d83caa68672b2ce6b0421a7a6f6ccabaf8f707d40fb62295d9811f09b973b3f54faef5b3178f9
z7287748f27a46e1f13a0606bf9a7c4e0e8c7fbe5b81980a348cbfd02ee755cd39803808b8991e4
zfb030a2ae2f0502353229ab07ae41aa3dfb6e8a2cca21e989e121b67af9ae7baf2072ce13312b5
z980c551ecd8851ab1afe47b3d3e7de2e02ee904d141b48312bd8e2106f6cdc87948297c437c6f0
z0951e2f2343dd67fd8f6852268158c5844972f378719a98c62480657da1d1dfccb65077bfda109
z6c1d2d5b61b5777878da5a9d53a6a83260b1e6cec9795b29adbe822131abd5567956710253e058
zfcc338770b61d1711cef302f16f009294e7b430ba52f38e8fe20521a2b4ac6d95c28b43303cc13
z183c927f1135b1708b80c17a50eaa3b33ce5b9b26a6283e1cbc5e665116623f06797e57979f075
zf467a97f4b22272ace8be389fab6442a960c568ffa61a4a99812dc91df468de679dc4cc9f048b1
ze107c04b2915f108138ae5336408584c5f07f490b05f43eeaebc231e92751d6b1308328018e23d
z00f2d67aa9a8eae67008bc08d9f078d12f2c727b0f9a0aace99b16df5ba7fe85732534aa75bbd6
z6cc325a34a7ff7de91fa9aff4abad97ca3593c66a8fc247e8fe17db5621fee5f3d9de172f663b4
z7073cb534c868583266099e5cfa47f16c0e6afe63bacc87a3eb039b135388499dc665d24466742
z5e1695cad543427b6166185743395055a04a21e9d8251333e4160d3b6cd0552fc73c5420fb1e99
z7f3f57f9541123c5c7fb4d1ed7a3d7d769f7053ec5c7dde00786b7e985a0208083689ea7b6b728
z34a57950906bcec828ee0be33ad7e9a4053472aec6ceed9aab305d861787a62c90017dbb547258
ze6cc6c217b1bded1411f5673535f46c653d160a9a615febaaa0c80ef980460498915c41f2a1d0f
z5c0674ee195feaf582c94091f12eb2ba47afd540ed0e4104fd751e75818dafab72708e3de8976d
z87f02cb3c81a880a257754f10096a8c14390d84de0d084270173ad5d06a6418a22254b179e9942
z424e1c94cd5e38979bf6736878b625314446d8094cf56986fbb29561e0e2ebe3a144393a6a9e6a
z829ab73810fc3cfc9bbeb5395200b5c6ab30dfacc10dfb4dc021280df5a021df247b6b9b6ecba3
z05c3629961ef068bed15e63985cf1097b445d6814423273cba36938936cf5c4ed753fc6f39ba9e
z9085ebee170c1f59ddd4dcd96149c23627fe4bb9efee96239e8a0210c7e7febdfb6602e475f5cc
zce2c568d0a37d8e426d9bf673172624c7af0c3b7ff733f872b84999f88afdac5731e08f6de6216
zdcbc2ec9a2d132420721489877e5ba92bf6f7f24f123a6d9f54555dbfc3c4cb82e6c53cca85d9c
zc88102c1744a1dc9b81e4caa0f0e2e964d5fb5626838c445eaab6333edc34e65f18c65d89e932a
z03d4dca40e2bc4e5370c54bf9e74646fa21adab1d9ea5850c06b3c515d120d4ab8c20a6ace0c16
z3bf5dfedb264747415d5d203750bd6b2116c4c11089a64d03b53cdb425bff9c1a9bf849b389068
zdefc0d0e899f0c12ea18b30312cb66440e70ac19063410b012ecccbe82abed1271887b9cfb6e5c
ze05ce158f88d4eed5ac2ffb7e396e2e93f62e12204618a57dc755c89fab7cca267ac72f62a432b
zf0dee8cb74ba94f2468383eabbc36d1505c9154225a36bcb87a7f2eb45768adda7814f1da8b529
z661c5a25536392ce8598191b997addb7b825af55f37b3b6f33a664d21efa90553d99f13caee7de
z5fddea071612cd97a11df49d08d49699cf5f6525a6a288b32619e0a7c176942985098e651b93bf
z592dd2549cffdd9c37450e59076df5436bbe7b5eabec06823ae649bc73cb81fa33d059b0506953
zebbfba0b1c6bc0ea17c8ce48f0bb78bebf36e22e2a2299fb86e860fc44635f403ef0e933e741ca
z7a4e33b6e28642303be62ad1534ce4c3fa8c4e56a998b0eb86bfde258a9ff1468e0eee4a9073be
z5d0efc37d7d6c00cb4e19f54953ca4146e7d634455467550e9cef109d2ac036c400112c9553916
z274853a17ccf0adfa23f81c989c3b316c93805d04457186c3265e26383a5c39c83b6b56a738dde
z05c6306672b9271119e6f67d7a7f9a822bb95bb4d2fe66be1d8df82a12d5d03910be82b64aee65
z5f9002a6268586975a21c99d61de6197e6d008504ebb0c0e397e573ffb6383e9a86a43c14346f7
z1b6558eba7570e137c96712a29249ce075d3caa686e92e937d4aec59b3cb873a414eff34beab23
zb371f7d146c2fa2b571de2120eb71d85ee5b9e89fb98c827d580259c3ac57a1a595bbb03cca82a
z8167811a6a5f0574ba96a00803688c58efe460428eadcd68313e24368a6e9f2c839fa4e582427f
z967ea5de6f7efaa152cafb28c28198af3a1614fbc73544e3690602c5c04d6baf00c323bbf6d059
z60d4a79f0fb3594e2a51f496c347593aaa786e6f17684c5252c89a0eaf0325c03a8b7754d8790b
z14efeb23c68224f4f07dbb42a13e8555264e310b78162f6d1a588417d454c7a526e324182c0a23
zc063f87015eed2280bda6883eccb1de839f8946be34de7e6a2e3f768f99db96050a264e2b45bad
z197c14646ea6d42de7bafeba7922d4526a07a440d0505b13b98a7d3bff001296b2f2434b13bed7
z0e1f72604b0967c32dbe94fd770b0aaaf1e20c8ce5d8532e47f221ff833e4fe84dd64a547afbd8
zcb797d88afd62394b60e455fc76e9da1ed399a432d76f816e82bbcb1a7baa1997fa1213aa1c385
z8308254b8717a615471844b78bb17ab98e223e09d696f5221d5701c8fce4d8a192d671959cb532
z897cfc0c2ce365aaa7bd221a31c4ca21f1a7a354a38f62f8134dae6597210435375ba3e8c3b7e5
z7778f065110d8de0cf213799127ee88cd4357a3c1845cf93c16ec44b98a459a24dee544b2d1943
z659901e0f4634c7e00e6b5286bf451bad40e06b4456a15f6691878330503e8b6ff2f6490f93d6e
z5821f615693cb9d2492aeb7874c6aa5b6566a0175ad29faa148cd43c84c8c33082bc4e7b6ae3fe
zc5bcad9462c6c4ba03ae2a65c858ec5b55e6029e777b3d41a195e81ccd92df4c160fb57b8b088e
z93d8d950d3db369579d34bb1fac9620a8b7bb656371449857750a71a3f1911924d1d15e48b9228
z4cd12e792ded8c7180be37b9f476d083b4fb4435beb428282341dbc4f585944a14636cdaa79808
z0d1635dedfe1455fd72a41123adf63ed67c7ac6a2a261ed029a65706a2aa80b8af03dc79b3c945
zabf784d7c6e5722781f342022624711ce31bb84a3be08db8b77bc8510fc7eddc753f50c0dbd71b
z0c43d02b3b5ce914184b66f6abb9ee0b0f628ef07e162c7f8213f647f15e482dd7b65ba87af824
z5122af359869eceb54a8ad1b9773f4b604153e6addfc1c07625edb2b7cf5d5b4273c0d5298d705
z39becca9b95b322f9c7a6255dc7c99f0bee468cad661f881fb8665ad6ef9e132e7ab6c8ca12cd0
zffd20fc1e96ad4028f8e809b38b45400c9b1d713b77e1297b41e0175dcdc4377fc74f190da5636
z79851a49673e3740388a3adb82e5f55f1c601ad2faedc4e6ea9ce7013b500563cabe4605f492f4
za17a764553e55a14c37b522e258ae48868b92ff991be16aea75dd6ae74044997bd49c02c108fca
za953f4b9f0ab1f51820e5c26014fa9441a6ba3b60db2af759cb8543679efff39ec1cd366a31d69
z0818f73637c9524b51a097e5996cc7cac941b5567025efeccd6ca6059d544e4dd28baaea7e64dc
z64f5ec35caf39275e9fe7934a53ab90543e9b70849f9a661919114956ec84c89c122b7ae737437
zef476786fb5f3f774fea9189d190f198b56f3c1d41c7f627af3ac3916ddfdcb44ea2f0f57ba88c
z9cac7f6a2893ec4143b887c81b9a20aaa3026a7202bf41452285fcc6807d315dd64628d3ad0ceb
z726e7b65abe7cb4cfa87a128fe82ef1b5700c54d920f84e9e2eeb9dadddd50cbde181732c8d41b
z0d06879aebc68236cd949c6f436fc6adaa6a26299536b58876caffd857115f2463ae51eafe18c9
z5cedf51c00159fadcda071ebdb62287ea35eb4bdf1d80104c90aef8d5bc5c8fc9ac07c7f212936
zc5ac57a3186c5dedbc7d5e49ae0b5cf78ab264d0c4a5a03e8f1c7516de4b29ca4b443ad977013d
z58d2b02dce8932c1baf5f49f02f1aab9f15047d74efdc0d9b16808e759ff3e9e2bb5a8fbff09e3
z0495a76d80affb2ed484792f1def864acc06fd3d7e1bb0b5b5a7cd5574c37758aa6a33f4b5da21
z7db773e08d1e41a4a5eba7c46e7716457fcf14472f7319a46741499abebd31183a3386377330f4
z37db45dfa6b72c6f85ef0bf01e352ba63859d92b85ad8bd63aee8e1a228df7e3be07de911b5187
z32d51842198c50e932eafbcef13110c82538b9b26da16d7ad33ebe8315e31b38d94e03ea79ccc3
zb3df5706677c1ab9fde1e4f83be95d9e94ce563bc11e2b4bd169b9d111986c14c0f4576167e901
zb0cc26dfd6e36eee49c0ad2233b08f4480e519a27d4e5e3c1a9c4be421669f25875381afe19924
z6ff4a45f520745bf6f72673443732c4c5488df27b12218106ef0c0b5080e75d94234185d798cd4
zf2759df3b7e95aa5b7286de59117354482889b270ee92691e88f5b1d25301d0297c2c60e0b917b
z4df472072f78aab06199ecef9160162a4e0c20e387f742d4214b876486c8bb475802819648c609
z2bd0c9d319ccff445e474ab8d9858e6c5fb76c8a3e40e5dc073bf43a7bc2699213a90bad0764eb
z897f863789909ac527203c841707ad520296dbef6e9033f53f1069cd88c324bcd4842b0e6886b3
zaf827004c9d20af0415e563a7182f4ba26fe8879280453f800e9d5db708fae85a2aa344c44406c
z6229d1438aa75c07e18559145f1f72c6c240fbff122a7d0ae2bb280fb3e546093e1a1f3de89e55
z094cc46ba7a1f281f1c20f8fe6e72da8c9444e2951c5fee04f56599f8ca81edbff62aa428655c4
z5cff91af80d59d1912ea2604ac624b439c4bd6a789d55b2eae0349bc00bdb7df064c06632a1968
z0636b7d171f44c5a8c3f4ab271ed0aa91b1e71334aad919a7a124fdfa36a5ed5db9321a9d1d738
zac90cd13bb9fe8474f81a51f304a802a3cde56a25721ba8f9cc9f2152b6205e0e800673b78fc05
ze4bf5a4f8e44948c3d2fcc5f3adf91d776694013c8a0bf717da1b49a83086a4738e2228aee2c35
z13898e7a4b474e47e71740c6507aa14561828b5de6fe55e42664c2914a14dc86509787323b7816
zc82ed293f9180ab188fd385f8cde79879166f854d05c558e7200cd68a829337bb7f1597daf789e
z8714c8e5935b6b7eba2c31f651134da25f4207ecb46289d4933c49ca23ba75910eb52e8be5b39f
z80bdd5c3370ecb795becd18d80177ff8cbb4330d39987813ee6a69051818e274c8da02e3ff416d
zf8ca1e3d10d007d77b8b58879636bdb021d183e0e582d0972e53f90d0b878059df002bbc71a639
zd0d56927f2142509c90aa7f2be88985b072a802404f21b559d06c298b99ac06f4edfe7f338e1f4
z8783732da7a55693c3a5654d47a15614bec501b156f8fd687a8a10b48374f0d4b02d89ee615f7b
z5fc2544607e83bf67cbd92497bfe8e117ea4a03a3924b3429881ca7956f6c5c7f57e7f8eba9ace
z468dfa2206e0e2709ed21b6848aa71888208b41a1778b93959bba4733ca5346c2fae27b0aaecae
z593c569fe23a49c2728835084c23dacb6767062a0894be4aebc62501b878be6837d093f9c7e24a
z1e19331e0cc34383be67a0a4a52aa2084f572ab824e6c212eac88c36135011014f50c2b6bcf387
zeb37b03415440b2da64d1a0766cc3cb8d0a1d61bdad90a0853b1f23b1ca854999d35ceb9b908ca
z7956b4133878c7d633c5b0a2d2a71ce493533d654c6b658d32e1faa911823c04eef2d2a6f33c80
z19636d0f4bfc40cf1959fd020b01d1d58c960a3fee8397a129c1c5007f3ca06f356a0ca540dca5
z945637bb1519aa1c9ea3952c5a4e16cd204267b00b80ab2eb7d694539e57c1c04522b820824398
z04b5e940ff908f862d28a25089896c928004b97958f713b8d2b9f2940f9d3c8cc959e91dcbe837
z046aebcbfd4bf2f6b0fcf7226d451e7421f5866cd96a28e0513480a97235b764bb4b415c08b25f
z39142e10eff7e9382ba7890621e0fc0a34b9228062e5d67c3c75f64f6b6d80542319eb062cfa53
z02c33a1c0cfb053f8ae89bceecc61c98e8f85634a1a4b6ca561914a678c641ba6ee7393691dfaa
z276b6c933eba1899f95a879a73129e6f80fa5ed95ef2a0f5e90ba92ccea05499762249e3414053
ze7cd9870f7050c1552d2ffd9f892743a3a8d0026f6dddea8e2b6a7a29407b81e07c0eef37b45ec
z07f855920ef23ed1ecf225203f45002019c7e0cfca35c656d3f3c37489fb7c22652f7693a4f3a2
z35e1bfde9a128636f76d413924bcfb3a8751268371797bcc042594f568dfda29ec3d395a50a1ce
z89bb7d368b1212a064c131fe44c2159f751e1b8da56888f3af39564bc0217c0c8391e87844c5fb
z289b046f8a60c39e91f42489799b2f8a825e3279c2f586dac42149e215b58a4a1975ab050052ad
z4c24c07e4969b582ec02eb1adf111f6ad0eb7fb1ff381731f16e0bc1853d973cb554cbc550ea53
zc13e8a3c341dcda218587ab93e9365760e79a7590be55335d59fee3f69a533a4fc2649cc986a76
z74d0265a8b6f336cab8b3a0d1e1374aeec4f1ea783d89174372247b8c187e7f0362b15abb9efa9
z4428531ff7ce8d4c7d188e4b31326e15d021aa710ed0d2c34a1b517c58cc77fab5bc37d5d0dfcd
z776aef2300a410e7c057a60bf10b87a6b6deacfa91b27cf85e48bfb166dbce7ccb6c78da43cf43
z6ec3cfee6c9d7ae97fa6ea282890b934f1081a86d7aacf1b52c504690a8f9111117a54011bbb29
zc18cf1801d2c547b98f5bdcd4db97d002514fc6ac3bb2586fdfedecdce794989068cf758666765
zacbf60ad6e7f93642bd7395d8257e04478517eb9b885af31df67adea1b60ed7134980e4cba664b
zc8463fa59d9f80646b39b32c94335ae3e473191e1c29c815d76bf8f9899407ae22b3cc298f9adc
z879e27dd12cb928b0167ef843ba4556bef212ea072cf5f078344b038163b34e75b6cb1968ab5d3
zd2387515ba623f28b4aa8b497f8d06c40c8bba42c9d1762ee744f94cfb7c0dde8346626e4423c1
z3626062864b0b04e4a00e670f841c70e3c73b6af864a2aa12c0d89a89b5cea212d2fa0e254d5c3
z7d41e39bf69bad2d530270661676a79e1425c9e897b14d5f4a038c039226943e61e13d16ab7cd0
z1c2d0673917367297cad5093fec3a2dccecd10cb69af23d83c04fc85bea703aad31d563560303b
z71a2da1cd275c6f1df122eff17263f80563004f8d579b8cb8cc15bb8ffba6072b3da0c7e7ceeaf
z8385d1c7f0740b401d8070689f7e85cbf347698afad1ec145c990db5e96dd46106e2874d0fa306
z93b7a50637cbab32e1578fbd6669416a6aa04982b297d3b3a5b81417202ffc88d758001a126f2d
z8b3a796c04da6849a7e087f78d142f82cd2b1d988dee2a45eb3fadd56e35c5d3b81c583dae7101
zb8b174fa3245420e0520e4d16d2ac23475a81fa937eced53c0266b17b0ab196212962ee60bfedb
z35a18548476fa73d8d6d9b01be87dce89c2a6e3c68176b65e404a4e87daf8bc3f51511b25d1543
z56ab0bd37f19e559ea117b294d0c5060b505dbf5747278e330bf28a6ffca5a54901372845215f7
z19ccc9fdd36240c2eebb25e18ac8ea557c666be346c28ab1e87d2796d2373b8a6faccb1eb1ef6d
z78582b2961fd748a2f4e59cf2163f357a721c2272f06b75c5f5d3b7c1176af86e771e6bcfc656b
zdb670fefab7fca8031006e30d401a25830d60d7737b1366b8db82320d90f2fcb744cfe1bc7caf9
z8bfcc624851385368ef7a5813b47b5916abc33ff05f4c4f614f278a8fef5f247b5515dd40e6d77
zd96880bfd57c948420822b22c7d53372f487745aafbefaef18e8297ab910c2fe2598fbb074c303
z694a38067cfc2995f956e8127eb05d181793b4e02038c2f5ebb653581c2caf2bf4fc74b69fe848
z0904c4d3b8c9264b3ced3a3aec3b93a2c522fc50c09a1e278ca2387e4d760929058b0eee5bbb7f
z165bd284a50c9832df0cc2b3b1a382b5cf837fe116959d428a4c2553dbcd81324074ab8df18984
z5abd7da89f5f352b5d5febb34fb38b38d896424260c10e2848ed58cfa746bf01a32e99a1724a23
z29bd03f228112313a6b157656c5624c3da3e078ba4868914f9228518b64a202329b0622a229c93
z5515ebacd856f0a0f1a01a355733ec4d5700c671d082e2d58508cbc24c844b77d05b0d44f85978
z5b6f8454b0639734e89150702a15e89389bd3e03be3958a31eedecd425a378207783d99927c2db
z810e1ba62a1d910ed07f10bde77192e48cfff0a1769a98a6cf6c09e1cbe0552e746524fe825f55
za185737485b0388e0910de18e9c782607d656923768ed3d05211c37d362855611574e3ba37cf87
z76e4253d2b6aa21de2103858659f5be6d8f9c95d355ebafb4264dff5af7009856a99276f85b463
z7b358b02c5a43498a578fe1676354e09fffb321d5df1c557d38f2c01cbb72307aa9799f7998fe9
z2e4bc9bef045b3c4276cd90287195bfb64e3735167c8f4e514f55aada3acdd528c8915962e9207
z4ec504cf019fcd0fe4ff500d54aec8e89f6616f80cfaf2189d5e769079999d826fad1f21da9e48
z903683b4063e32b3b9e6b149c083767bce7a675fbcc6b2e336c804aa39d7149da6750b8e211826
z0eb599275ca6b999d4dc3779393dac30abd732964d6036f113871cd59789d25f33d35433a9459c
z40be0cd5de0f7050b6354c461f00b7c5c88af2acfd12a7a8065da7ad4866816e8f7a3ac94dcada
zb9f56162259225e8de1d1f84eeb2e349ca0f17de926cae653fb4ab08ade4806e5cf8b7719fc940
z4ec93dc9b816115b0bd7f822d7df9e79dad04aef5689a1bc488cca932517b4da3a4bdec9fca91f
ze98eaf3cc775f2104f984b252ddadeb8aaae5098f0a83fe1deb3442508d1089cdc51f6b9bf9a9c
z3bdda4ce4fe7d9bf30181db80435a1af392b7099a8a2876c06c9df288414bd3c01a2cfc12163a0
z56732bed15d5072a5361a90ba0131582590d0e21154c45b390aca05f6662c26662213b5a7cfc3f
z3397fc86c887b14c685a7eb4eebe261c2d5dae423e9cb173532405deddc198949455cd494a4810
zd3ec6b00524e50288702c4f73ed44636765b0b210d68045415f273fdfb91f15dd870aeb7608b7e
zf2d5195f9492e18f25817448ac29d4ac831fa4e5cf770a7879a859d67abdb5fae62852732df82f
zc1a997feed22e3af102c2627d57b590f3756f23afc44f7af6d5af28b72dbeb8a7d2b6da5c91e10
z4fc56ae4939d7bcd771bf5f0e5d78a7e8562f00a368ec5bff5b3c3677e6dc60f078ec5c0088df3
ze2de581db81b66ce60591140efe072ea551f4fb68b786dc1166af5d2ff2f49311832b2ec101f79
z538eaee936d5ec671774c9d0da2b954671f687abe0758bd97f5c6b72d493efcc35867e619626c9
z2bff36bc8e05b9e66230dfc212ec07ee4648eb50ddefaea343a38b27f12ffe7a8ff5780fdd21c2
ze25538b8180ffd79b4a22689ab7d0d3bc736710c8a87291bcd6948e95d696e9cbee0b3673f2e49
za0d6c3edf138bbd6d1c2a24844c9eb8f16b4ecdbb75bf007d1849fbac6cf4b2c38236740a75ee6
z28d438b5d261a24bf4a244598283fab9338a5be28a5f2d4e6fa39df28f8b75c1102f0293344494
zecde5557d2fd03a9f1023b14bb687ec4700dd99eabb61a54255302f1b575a7ac3e9b51c0d100ac
z15f38471a49345c4690259a72fb2d51b01909a0ffb923027022c68a491377d54540ce4e54a4bda
zfecbf678714078610895b3f42654120cb493c5b7d56ce647c738510bddba012950e4323c0c680f
z1be1af3f127fb18c119b87a273e788c6bb4b133b2fbc61eb9aacbb2f38183a432aa3781e5e0238
z6ba93aa6ae9ec1488b0dba20b5cdf21c8c4330f821df50adf7b9a99d385f826b5b18ec9b628122
z89a85be930abf74006903e7ec9a2f1f2f22115a43acdb22e5927e49b3765788964dbd4030b0bd8
z38f08860fe2e585f4b520f1c4818209ecb2f133f2a1cd35538077912fbd632bfd6abf89b271bb2
zbdb80726683dde7ccfa2e4ad4638b754ffba042b5d1db4132b8da19492b08c9ab49778a34f8cfc
zd8b77b16dc7fa57e97fe89045a98f34ceb82f39c9b494ec5ffb2e8992ce210eedac453dd023493
z5e8fc9bdd19f1b88863655e7d766a7aa364d310853b5b4cfd63d1e9f65db714df9bd1da2646932
z146ad435bb068854eb5e21e2d0cbc81b15fc746c98b103ce76cc1ee3f523c1bd774e3ca97492fe
z8f0a44cf9bdb21a57579cc170cc585d32aab456d12079ca56784d6e1b9a4007c08b327f62b48af
z33746077d7c8ef2dd7ffee114d52e3d31fb1010526afd22ff2ecab8af456dc9dbd814d77f7604a
zda638805141cc6c41ee27b15b6ace4b4c1b95257ab6a690411966a20776c554c2e30cd379e3384
z22a25074b324fe7bf429e5a64845039beb46315352feddf4884f0d066a518ba93ecc24a9be63e5
z38dd7f0c3f1365f6d489d9ed0c8c49ba2fab564c399f85598e232ea8ef75f0ebc6f10de078499e
zdf818bffbd0b069500bdcf6ef8c066045aee8b5bbf25b62339a2a4ffd18bcaf83b82c5ee63038a
zc67b0a54d9508c870a7bcb5ac6f626892141f4b6cc62371d3c32ed5ae95cf26fdfefa9fcd60b00
zc8f01999f6ec7bc15ab3270ca9308056bc5abc1a4afd581efe2116cb71fd173dcfd3f50b078eee
z5fa8817514f3148430edcbfc6aa8c4433ee965bc7768409f50437443c8146b58d1088adcfaa866
z4f01b677e1e8ff58478718527eddf6e589904815db9777eca450ffdc1db11b734242a33523eabb
z9591a19062ce9c91ca25a90df55f8761b2d6f220b068349444f7490d8733fcce6f394d5f53fbdb
z217f700a27c49da88a2ada7097fad4f21b6fbd7f66cf44f60409d202b503e0b60939d094c3e1e4
z20174178912d6104e6998cc80dee5f5521a7269bac152cb98b0e08ef03b08877ed2489a644eb59
z0a9860f5555452026e2dcc9c45f9f65af0a38281c833febcc754ee08eea9014af9739a9a95f31e
z7766ea3a33b51e70b6e2852dba8d8052212d9cc070dd966d302defc6d123abb5c799d42200da0f
za77d338174c451956cf3c9f25f52c40e02da1a63a5565cb33fe385eb0fd4114cb812ba3ecf15b9
za3439dc57760fa7ba0be92152375bd9a4de8af63b0a1e68b78e0150ea2b39c43ad4d84aa015cf1
z3cfdadfe20b072d376210a4a4a309d41e628391bd97f21107cecdc342c5e13ab2c87aabe9c4001
za978c58c5b05a9cba7fb21f8ecff6670d5d1c1ba6d88597c8bc8653b2fa74563a68d6d62f31adf
z0c1e8c1cbe6355801b3050df386a6c4c36e9244c8132b94e020dd08b3e371892d7f950b7382aa6
zb4200f3f05cff176ff587c29d0ac3b9d05622c1ae704912aeefdbbffac17daa19e4805ed846bad
zef00ef0522993e9aaa2061f35c8cf868cefaf9b0f49f33938ed0686470901d950c7838a1c4c125
zf46480b7931db8f49f29f4b361cef22443063fbcd039605b2d2a11729c74ffb00327634aeed264
z63e20637e77e41b7ba65c67e60b3202c7bcbf3ceafe0ddb73621c2f172d0ea8fffd16dd321764d
z2671dd8b0cd1250d78c34814ab18b0e3c92eab24e776d3e4ecbf9865bb4e1857a9759408cf677f
z91a847490dbbdac6e9a8e9f488679805f70e55994ebe2ad821c5fe39251785546f2b3e53a5d89d
zaedf52cdb824a71a7ec5fdc96e0a39a8819681d9e727facc935eaf61012d45aa61c7e98b3d0899
z86866313941f79c76af3d44241f16724543e0ce588f01c11d2a4ae2d35270af9a5793a28267cde
z5fab93aeedc62fd9387322a7a1a62464924f26157215270dffdf735ba6ddae02e67e743ad383af
z0791d397248077093e0f77d52ee8846281f0500ff909056f579ab1d218537e729614f9f286f605
zd8b73f8f5c1df12d99e615259eb74d2265f4e7ffc7a958e108422cc62e6c4d0997a7e3a343d657
z63c7aea5e0d0416825d5b4a983c02ca2ee7436437a63e1f5614b25ade6db1bf14530feeeca1357
z26f3152ed00d6906af01e31cf6539e9d0a3da9cf6bb212f65627901b1f6a88fd9e5ee370550e80
z4b6a25a8ca852a0ac3b328ba9861239e009a5562bd4af1b5fb8b9fea562a5b5e8db66f8054bb6f
zc16729f3f82de9954983d5f1f74474baef8cb2b6c4f6f563b8e3a24b00bd7f50521241c680c947
z5996704f044b25d40d88dada211f35d6a49a5929234864e86c09ab6e62e92b573561de72b1ad6b
ze46373fafa7fc0e7ae7ff8ec44d01851bbd6e46e65f5f3685b74f7e938ce4367a3aed822798e49
z1463aa7070a007dc1ddf0c9e2a44b1e395e8d5f357ef01c7741e4ba3ed9b2064a81c0a1f952084
zc4b1909fe8f857dc8dc9c4dddbd4bae56e12f6cad9746e3c852718ca8446481d2611e78f5916a3
z941c35f641a88b20a0ffed69ee778137d0210b1b3c3614b8bee0688cd87a55ba239790f3548c8d
z01d9653995bcc9b0560ffc9db0faa43f804c3127ab8a328dc639037b658fb08bc2bfe353173ba9
z0f246b9c9b80ba7216009dcb9aab0e434801f636cd2c3e54789d51887a34e0bc4e588ef40c7cce
zacb7a60c48df2ab91f2f9de8031f2b0fedecc8832f67f67554056951d1d50abe10454cdeff6abc
z3175976101cdccddee2f66fc01ed27d1f5c004ad5dacb3b642685fd4f4f5133e06f36d910e1d48
zdc33487c8634d20708b6ffc46858093d87fcb6483f9d84dfc225aa216a70404ccdc7f1d436f7dd
zd44f60e3169561917d49e5986ab583aeec30644fb168a1940c66c07fdc7f6b5d7bea9ae0da9c44
zd79d1a1a4af9334c3242a26732836ceb9cda856ad72e29afb40d9a461cb7adf0aff729918408d5
z1641f845a7f4a67593afe0c9e89ceb2e8255c0fa85599274da39e835b8c734057e3710a95591bf
za1ef7f0f8d497cfc34a27d30944f8a5d03996b29a91cdcbdbe5c1e7a861e7d7507c51ca3747bfc
z73d7db62b505df71a7bf83a37f2c6c903a867f304edbe33ace240ddf3c75d5929ee4cd1ec4cd8c
zac5e2971f20adaa45ce4b93eca1c1b92302097f5d0d45a4cd6ac65c21a504c3995e4fedf2f38b8
zccf8193fc5cbcc40fe29b4764dc34981971515d78cd513d9a6942320d1dc32874e0fc308e105fd
za20f878c491e4c20c46f7f7492069b30ed85bc74cafa91afe278e5e4f36fedabbb57fcf7544367
ze5585647cdcaaaf2ceac1ebe08707c344ca1c8459e7dee959f05f3957bfe3201fe8916a88440f5
z5597e841c08fe8c0bfe268f351d2076b5a10b04d97873d347b69f60056c9dd56969c63b4d2f97b
ze90e6f8f9601113971d8d6ecff613c48d3f2806dd8af8df1d284d8cea80436359a37b4f7a6c56a
z011c2d282e4fd3b589d31000865b7ba8963b214acecee1012991a12096ff4a3b6be3274ccb4e05
z8fac37ba43b1b83ac585b69ccbc58c37dac7c8af1190d130bca8a98733f316633df4c1765c48b9
zb57020f727221f9b779629218728c41bfcf572ba8d1d381fa07ea041dd1ac19a674e827da576f5
z2708ffd12bbbfb02fec376ec645d11e6a6480e1ccd11651baba0b6824733377f36457f924ed308
zb7cad6bc7742e8cccfb87c2c097a8287f464b830680055eebab214c3787ecc91ec22b58adc70f5
zc4c23f6bf9d175aa096887645fe36c1d12a9b2d074b30b2d95755449a7dae90c60a0dfce6e3a57
z24c51653ecdd3a14b1fa61c5806067468746de2d69d876fc9aba9845a5c2204e13edbbe62b5809
za077a7804dc305cdd597bef3693cc41221bc3075d65c82cf53a7ad913899a7306ee033796f0069
z17980b515c97e4436336f9bb6594031f0d46770a4a95dea72afd3ca6350c38a59836c0ec585eec
zab802496a86769681420476b6361d8ca9598f2720b0c540b8f581aeb9066bffb99cca6534d55fe
zad284c1af9dff2a292560e9870fd2c2703f1ac36632a96f7a2baa5a4636877be930211de8eedf8
zacec1b440b8f77ac3f4f7e95d981ec96dee3fb30fc989d6ebbff6ddbdd0497377d3e73a8a96f10
z47db5eff916431fff88c77034c1fc3079832167ae88475289147d87201b39d994d1b13b51b842d
z6cc98d940132a2a16be023361e50178ed0f77d92ea26fab56fc92e0da1865bf5978aa50c11a3b3
z2d5bbc17df8c900ec6c4b3ed62c14be779d8380e8ec0fb7643cdbdd1f3acbe6154e98fc9c0628f
z467f5beeb00ac3ee98bb33cac58b98bd061a76b5993f8530023774224b21a5a8e110135baa6876
zf337ccf0a55c2434ad90cf27eb8b2014a18b9c7c086709a44070e1ff2385d9ff403fb523a4947f
zdc01aca3ce7500ea3abfa5db066c9afbb6b14077537b197c2c4f012826e3b104dbd589889a184d
z12462206bcfa97e942cb107a73ab946cc6c6f3993e638638e0b2c9bc5f6a53f144ce7949928cc7
zfb5a5f73d44751f2cfc1218681e09bd87777caba3c428ceb6ac000f52c29e548155dfd6ebd17f1
z64e6af9eae40947a0cee216a090ba8fa65d9573f61049baba0f2e3b3beef1fd5fd8403f40d2174
z24ea39f73660c7779e80fd559ac3d56b7b7f046aba209b675f67055a5b94d0cf15f4a73986e73f
z4cec62f256a9fc841f7e6a54a6044a16c1afc65f4bbce47fe732309347c8982706e559a1e9849f
ze001f4232dd34262ea1485fa60f60bd875d3b0f5d82ab9ac20eec37631a60e2ab02c5d5ae639cf
zccd7478e88da4673d9ef5fa037d28e022c73f20113620148e212019b1c8fa6d0c07ffeaf84628c
zd69e3f12fc5e3878463e954082b7cad553951c448d8f0d61aef0f2afc0ab43e02f3da0cae72667
zcf9f9591af5441c3ae88478f71772c66629691843d4b6eebaec60ea0efcab25af4c8a24edc8af7
z60cfe379cc5cb754ba58a05fd0f51a4c3a5fc33c2cc1fc8d404c371ba02904717ed997aa2284f0
z94ca531c3a238007deb62c3c0e94b692ca4b86c9cb875a845b2eccaf0b427781d9ef236154b7f4
z15b80d3bff3d515e1724d5a994ce0a0cc7d56447a5d219cf3588ffce3d27dd084b32c347d3fa36
z9ad90a955c98ce593e0b0294645fc045cc77f8e8924d586ca5099e2c8bcd4eaf01858ec9443fbf
z199881a26f7e88281d2ad71c3d3ea8b1dc5da12cc27d1ca7d11e69960b750ecc9ed716439ec1be
z943685e970c2d906952e2e20adf5286b714a8dbebd9820b657ffc1f20b553ef1b238d48d598856
zc92671dfc6af757e08f05d254303557addde5e80994bc869b202c09184fe720ec23eca15ed0068
z709c1acbc456f94d8e00b7fc7ef25a3b8e49abf5de8069fe793040b0c028fde4ca1f9cb9626a4c
z958b7d2fc381e04610af12bfde7103591b20549800e84f6ba685ca409c688856b52e854e5a8edb
z84efb56b9bab6ee0b54c50249af89dd26b8929f6c77fa000baf93e871a50bdf0896550b093ad02
z46b8f0c0660ebc130ad4ddcf377bea21d8bffeeb14a565ce97fa094672fc21b959b54d6f7dfbba
z98c745b48ae9b802e8e51579bf1b7a24ac8e6a52c9f993863160660bd5e29af9b6f3e8b77e920e
z81ddfd637359f30369894b53024635d3e018aeba59e6a19d1114cd4ee2647a7934bbfe2227f11d
z6eb701a880550309d285b38f8af91216403484d1ca4fd14b48c057fc0104510707d1bba401af8d
zf28e2a0862c80b2c49a272b1687171242a2d5e66fc80a4c99cb5450cf9824021e236cb89b03d9e
zf3a27dfc83d9fd8517f9269fed2bf3ed368ea42122f8aa27b4a95dbae5bd4928edf3931aa3aa7c
z25845ec3b2a9882b91fbe1e6edf9ef08b37a0f6fbd77b53745aaeb3b0bfbdacc45f33f18be28a0
z935ae612bbf93621e787f8397fce7872f12f0f8ee6d3ad57c0196a528786e24ee1c9dd69114827
zb5626f9b23c4b3195c66146544ba746ad82f5585d47cebb757c19083d270bfde6de225ea6763a9
zb9991cb23c30fecbe15aed849f73bc3488f71b646fae7180b1d801a9a12add8b759ceb67e8065d
z90334ba28ff05e7c7a7617c74ca4351622ecba4c83f5f853ffe297adf1b02e41e4dbebbf5ce57f
z323877f105502ad9d1ccd9ac42bef30da7351173e31c5d1ae908de3b54ca5ec79d63af176a08e0
z614a00a6e97e9a58fe611b4eaa04ec69f0a48c72cad809645dc893d3d448a13d86c3558e5b3149
za5b59e43e4b879e73e001cb68cbf5a396bc1ce8c16f96a08030ef4b8c68af6a4ff64a0526193a6
z428c82a5bbbb91c906b67b49e105fd113c3d76b205d7df2dd1eeaa1830237b23344ca536b135f4
z8d9e2d3aac3f003dd2511a8d48f8aa9df18ee6f43ef460f755399e3b645147bb20a913b39894ad
zef7c22d39f13fdb5b2e56af766695d4db8cf40e8af81a7af48e4d07f5560bd079388d9d3b1132e
z542ecf2223ceec68a16d6c6c86c1aeb2b19da8200f80597aa127033c5de3222c5bf3450e6a0d9d
z193ff6439e2dacfda537adfd0cc02c4a9eee0bd9965d1a98bc5224495565a1ead6151ea9cf5cc3
z667151dd0668c171f913b53ada2bfc2de79435f6a1986836028aea559092f12100fd2017bfa4eb
z4a141574a884effb96bdca6b3fd7a7c86815644c5d4812efe503d3ba5fbbb54068fbfea2146b01
z5f7454a413ca16936fb38ecdf7d11417a2d1f2b89e94aeb9a57caec65e92ef67598e4c0c67525d
z3f1a0ff6e4a045ad58353252a6988bf3736ea5ddffad1c81bea79ed5bfe43e81c2c8bbe9829767
z93c5fd0278147bc4da51948b7d0ace1cd620b6feabbe330235040d53e23e4f29168ade07ac7741
zb673b9ac139aec615e5a2b9b76d9a0e4935441d5984f7b91202506fa571a2fb102fad280929b31
z86c41120a36d2eeda60ec06fa49a54156dbb00d4ac769179839a0ed2ac46a3baeef24b5a17771a
ze476521b3018f0dad50ce8172baae15a965d1960c0ff9686ea815e8aa7a3848fd97f552d904446
zd490f00fda4f94635d29e887479572e90e68f332c143d79e7604d8d3af16060383e68230140548
zaa0a89e391bd394666b382a25b33f6b80b69881597509ad6895d0dc42f0d5469de8b6287b3f80c
zb7867f54469732d7af8afeb1207b9aa2a1a437da1f2bc109b43082e9f6c9df79a0eb6ca7db03e6
ze983bc3eedca985b94ae0ce721ca7bec918e6280a1ca6bf5a1ebaec2251d3348840dc06ec59325
z087d766fa84116321fbf21b546125d16ea821377c6b97a0607f77e03b19b1b3624f277c6c97070
zfae2e40f7b5fd4e97d34f5e0b43e6eebd883b4e16d36a22f558fa2e86d16d7fa28716e6c7c2531
z9a168e2d74d7e418543edd42ed6004d516bb1bb1f91945bf58696c6986f284078c1e1d68f77b6a
zbafb40f30c437662f1d1a1b40a40d2ca1f78022118794ab9d32287cb048b482bc6e7b217debe7d
z240eb9732ea520a1c985b474d647bfb18a87f69f6a7931ee0c4ce2a71cc9f4a821cd6f02353c42
z6d4cadd84317d4c70e604b8f862940448bf73e446c83f59ea86d2391ff62a813aef08696bbb75e
za28e08df8a86fdbcb8f75218cd0f0d40c7d1df08bafa72b1c99588da4e701eb310e42a804f5284
z29ca6a95374931e9ab05624a98f1a81da75b0933c69c6918f0397c8ec6b4136bd8db7f5e7ccad0
z6e294760f4aa067111c8b82c3c4647be8903673b8bd92c0e1cdd4aa68f3964bc8936b86799414d
z4eb5aec8b438a3ec23262c082eeec283b73056b308d47aac197639c3e4b18978f61e6bc748f727
z140dd9a81b806b1ae6e8f759b2e496a87c7881f952aa48ad8499fd942e8ba9d1f9d8478694b787
ze4e982c8855111651c0069be1952a08a80fc7f5a82bc5d8cdc7c019a85918b4fa335bf25b14e0d
z1353c2e6b8911057105c52c7bb7a41ca697df4661325b8d2498bde38fb568cb4332d0b2f07209b
z685fbf812c86a16fb63e84742c488cc77d06a633f5488b4e5c83e4ae18e2d1c74deafd2ed62944
ze5f1fc26eb02b9616c0b4752257ea8bcefeae025b82ba8c6f28cb18bc56f5eb02291a6bf96d9ab
z0813db2ff36a1628e50e91fbfb0f2e862aeb5acad56b4ae2af500ee5014ce882526ee38e8fa26a
z0af4771b552e753ad124ac43cb0c746895db6d0fa07da2594835d409eee014c51ce53b00b90d84
zdec24f88782c72593f425327adeae6ba09623ba4136243f8e9edaaeca87c174224db977a35ef06
za6b580df2c3245ce471bb29c9b1dd3fbc8a7f82738f02f6be66d51964e6c42e1b096079b73d553
z368a6c769ef5376053688702b7baf3af168198951d60305c71dea3ddf2e38e6ed01af47f5c3e64
z3f93d956aa779ae27f593f8ae2c74958c54208a4aa2592fad0652cb65461d007ff3c3cd9495a16
ze177537c60e9d01bced76104035507876abc21aa0c6d4c034b2d32f233625fe3fc0a404f052af0
z024e724b92d33ef6601c517d8151bf239dc7076d125d5e3b46d0e88a6ee9793e33567753851ed9
zc6ea77f4c860164d9a592ac13840191a958db33d24ac006af849f1f077e7e2573a14fb89439fc5
zabfcedf3378ad6ac5aecce9bebb51c4e332d6ba95134b53a325b38307c377c1649e7ffd52f99cb
zd10da341a076e5890f880d6ae28bf0e0b519b38bc008d3a70a1d706971fb5c2a90573c520d51a7
z8380a777d875e84b500de1fd66cc728d6340be8fc74f688697fe47e6a76df4d6eed10e17961224
zeb68f5006a853867a845dd8dc690b32a2bd5a6231d00662790b1656872a07617f423666726b1b4
zfa1e6223bafd9a182d72e64b03f3188cf60d42cf759fe924f5d86b25e2c0176c1c33363e4edec7
z1a97fdbe0459e868ee4e4797a89c3e730ad53c72264f5d51724b362be833f2a988527d548003b8
z1bb609b2b4771c024f2eea835679cbafff2a5c9b86f7dc802c0ac7f7ef27b5e79ecd3b82fb4c4b
z5d01776ccb410c23e1824ba11c4a9d861140a5e738ee74a8ede930a34db2a86c9a272d733538db
z287d7269676d9aa0b6d848c3df3469b7d08a6e7f96d7c5b437f7247384821363d5744c94ba0540
zb939a28b347209feb269d3f9ea66ed9482f08672ab3ff0ef99cf4eb50bf438e79cab3c5da3056d
z0aa56e15636c2e939a29b8237f159af62341829bf8e273ab618867b3aefbc9facbd38aa136b7d7
za37991ddb89ca4cf2baef03a74577d6f1f76465924b873a5954fe5ca219d9b484f79d31ce49a50
z68468e86203532778fbdd7818ebec21be0d332d33cf71cc9d123320dc56121095c2aa30b59caa7
z1005a5a8aad3877faf4cd4933404026da2dbcaa8187a878b2cf0778c95eb4a67d3b34267778cf8
z68920ef9e7dab4cc5ea37e846b42fb39581590fc54954ac7d687f367577cefc80749822932f370
z185a0f5abdae87416f0d4d6b9482fe4a1ddfade35708dfa0e399049732348fa1a7c0e382c7d585
z6d93822c56121049e8bd088a83f67c3fdac69b532d0e4b6f532ef781c3ca1468506fbc49f5b75e
z8f4a42226ba34cd3454784176c91824230c191811b0726268a6d1ace45599bf9987277ed153860
z03078bf9ce07fe560d6d6c1b21a3614529bac67b8a92e736b9d6105e3b7464b8256e0bb290c4f0
z00d85bbf5b3e5938dde6def57d0c4d57d20de55653ae2795c65b7a99d000832652544d83da5035
z19d85cdccd40dd23bdd77e96ae54c7b8566732087534f1e3108ceba08176c51d3de77be508b287
z39b2a8ee3a4778ce6062112c8131c5afe5250abf9b74c61f5b10421771a8851dffc33e5e67893f
z6da39a5761e63b57805725675e93b7af384c6e28dbdf2811f4fcd9feedc41978365719c6bf2425
z71a676d58f0e61ad5c5988df66548a48d6a05cb8fb492af0d9e5dfb9f2253b99e2f34c04342dd3
zc302719b13a0e4dd075066b97085c17d3546aaa2df1324d39623a4c0caf1dac652f7dbdd58052c
zdc2a4b77d31883dea1520b171af167da4b20126eb6362eb549793a133bf773b6dad3c7e5a10693
zc5fa41cbf88dcf2a04e6e5978fa863544c482a1ec6d7c415c8dfef38309b740040320214b4d635
zf30194c5d1c7ddb4ebfa91985acbf2c270a81cfee3dcbfba598ecff8a72ffde98224f03f2749d0
z0a99b44334615e0326f205bb258341b7dcbd31df63fc663aa80c62acda195ad1686ba78f3b43e4
z5dcc10d89a231681f87ab739c43d23b7dfbc68df2b667721769fb590ef71031aa31a80018ed0c4
z3313d44dd0c36e7ff914ac0493384cf3f548a3095d186afddbc2100ea7460ee48605822d5e9020
zfbc0a64ccb36877228b0093fbf9747b4c9a28cc2db15d51bfe56ce87e4f7373032c021ac1a0e30
zb573b8dfb2ec5b08e768345892d63f39772204be54b269c842122115a707da5e5ca11fc3718a12
z3a9349e384df027972408d44fa63aa64a2d066e2d5f89fb5e41216e62f6c778f55f10dd73f1bd8
zcedd65a54768849cf12d2228411de8237588120f386b545cd970a78f6f77fcf57e56b971c739e0
z2163573344a5cb861ce24186dcc724df3545efa39cfffc2d7922cbf15f95a3131e32175dba7b3c
zf2f0f59f18be727ead2a02218cafb13bb089d1d7cf8ef700f235b28d2dae786806f660d75d5836
z8ad7150e5035e18db656cbab5afd8e1802b71eb41e1741267f319a9e4bada76f23f5fa36894bed
z079d83e77e1ec02089841a8b94cbb97d9224a15e71be4307bfb6219b9aac3369dd0c4cb7e48105
zaf6e10f56320dc6bd0d2bc5d9c3fa5885d1c763d3837d51b812f82587b815ae1e493b9572c5984
z70dbe611742b809b742717ab781f9352b9ea78cebce79f6c2967cae7322fd085d0455bb97228c1
z03a8899d52964fc9f95e01774077117baa1c5652250f517f767fbf21861a9236236053f61e842e
zd23a5262bfce60d5f27547d4d6499c6cb1786e8fd2c1518ca36a3367ea2833b82706b04d10fccb
z4f11346db44ab74b02d4e7c80f7d448c244a9466506a048df624cde2948f8dc95d2af8b064ff07
z78c34546f2a181e148e93c4d1c5ef377933a0aef5bf303a15e068c21927a138499abbe866cefec
z4d1ee4f769916046ae4487cd776c307eb3ccbde425e14c30164541a983950550a69f85e4fd9856
z3fba26ac211d95426149b8df4050f6cdd78765892efe1c7c46312379bb7e57c65bfab4fc54de6b
zf0e020410c08bb488f786841a1f8480c56d3900100bf8a338b37ce0a0eb75f06d761048ebf6c30
z44b9bb3b8cd08f42be92cf8cfe55d002f2a2be554498cb076878842ebe3947a3fe02bea0af130e
z224cd3a76e16191c6ae9597a189fb35335884c4571387bd9702f2e61fc19970a30e3eb3fbdc755
zb9e88355c36e48d4109af15e057c725ccb4a5a5772ceb626cb5eaa67cca58f0059046be7228806
z599e4be1652e8e8ddb3c24b1452b5541985939ca85e95cd4f565c6bee16739701202d46e328d05
z7f2c708cee85304c302d177f6311b9808a77c991eaf25bd3adf281d1f2b7344f86fef64935a4b0
zcf49d5b776350cc7ae80be8907ad9bd622026b447ee8b3c4b531d6caffa444c81195dfa05dcb8c
z5b3bbf1f8ff46dbf4f3e1305c7c9dca61da0368b1bc9f08baf4144693112d189288fd4409a0e46
zf13a8ded6703c8664b775f0bd4860b08c1686b96c1b85f4b268128d11dae0007187a91a459419c
z0c6b7aefaff09d3d2d9804dacfdeb10afcf94d293375ea79bfcbea544c097a957fe24e16371c70
z21e06c5d1a8dff023db636ef67712f9443289973962dc0e499f9c3cf4db11c6d153b35da6b8eb7
z72dd67625d9aca892a0ec309e1e93b36bb52182cd8af05663a5badc8994c1b8007750cfa620105
zea786eec3926bb86fbd742328bff6aa3cb41da68c476b2c05ca0f4653558263eb5df62ff359cd5
z845b938f517e3dcea84b3484d4416f17130f49dce813b830578f5dadceb9afaa07327998c29970
z38155acd98bbc46730205cc5e22bae12e86411e79fffc188aa7b3d1b3e8c9bd729a7840c71d9ca
z8275d5f26e74fe2cab7ba92bf5319020cdea0b02238c449b6b57211bbc0d8664a58308a73a2aab
z53880b0274eb7e9a7d63f785c53cc2425b69da7c37fc57bbacf9f959909ad5bebd35c576225118
zf1f2318dad097f2cc00cfd9daba7ae4e6ab533a043429138c3f958d3c59ffd8ec2b2a589e304e4
z7176efdb68b1ff2f40c1df51c96510ca88665ae7ddd4bc9fa05be16b9f1789694f2de2d40c1af0
z5b731bb47ae3c6eef0336c0a22b982933ccd2928ffa36d0ce499fb5833b45a21b20a1bc9d6085d
zf100f6e7ac767b16c3bf10d9e54c040ba76dc7d899fde19b32aeb1eafe2ef20d71b698242d6540
z2c55ba63edfeed5d695c11e4f78c3174a2f6e6ed1472b4ea24b51a9308f82d4e871245a17d1426
z6f39adf6770ac8c356a243b79b026b19ce4e1c6fde46fbb27d763a21e6630b95bce8c979a2f048
zaeea409ffbd1682028475211ff922471a1c75cdedf94ddbd32a819172b3b7fec6334d9bef01ccd
z50ac6285a7f16df7c98d8f6726dc591c399a110179e241449002267602587da32c1734a278e4b3
zfaa60caa1b83f86443c72bb98e0c17bcf55e30d95e4f2660cd5fd3821bd3219d0ceaae437961f4
z61845057417e536c697aab7bb6097cf18831468581ed18dd7dd394a184af536a6acb4710a45a16
z8dd50bf4f6b735716f2cbbce3a0af9d8da9e8edf8a0addaead28edd45afabe9769f669cfba0fb2
z513f27721637a627b3fad4500467b011831f869865f05c817f8a7a38a0c45a69a37365e6d64d66
zbcb846adecd965dbe5145645cdde1400784f9f6b0692648fcebda1b5d2143c90b14c5ad01051c4
z8d85e87d1d968cd3f3c576c1e5325a36ec034c8eab7190246f70df4b94b570a3355e593da2ba6e
ze937af09db82f3724a00f8259c909adb6c839d6e99fa561051af5dd3deb284eb5d138d45d62028
z17e7cba115ed00d907000823802746b6be3e8cb554c587755bc95ee1e0e232393044ed51766082
z238c7ba1b7ecbd46dfddec068011b0f2ec3b08d2cdd5488d23cadd8b8e0bd3929ac9ddc806e955
zef6a475939a830f5614c1a63bc71490a385d1a24397aefdd3fddc3c4a0e0367b0e56667f5ef7bc
z50997e6066b73142bf9258aced7c0ce2fe6fe48c6147bc33ba725f5e917a06d14bf3967581fe0b
z6ccf437c556f19bf5e8ef4051fede4cf69d64c0c80171f6a43379c8700703126fa60c705d6abba
zbc8fc0c4b4d93aa1ad1e21f3b4f6837b20cb9f408845b4e6a4ea6abca6188477a62273209548ed
z8f1be5d01869c827060a14445c8d5b8afb8c7f40c706d98e9ae79d38c2340432d5da2f354d3fbd
z4985bc2b23d00574bf28db2fbadc47ab799b33bc508ed8b68f4b87b943ca776e4f24f18474113f
zc1f55cf29a9abb9b710c18b801bd73990ba0f7429515dbc5504c70bcd0e6934d9f0aafccbe8b40
zc2ad266720d47e66aca6f8e554832aa4a74cb11f22dd8309b757d3489925c0e22ca1f14a446c9f
zd052b9868d6e793babd3773b2d0bb24e120e4058f53f07344236c2665149c91e9aa4420be3835e
zf675050549f9258189993bc6cf0a8672218d7e898d6fed37042316a30b7b9d26bba5dd82aecf5c
z445ecb0c7c3885d985879e91cb4cfa7e1759114ee93cb6d8b4acf4260450f7cd1562ffa6b08896
z114fe668817027868f5124669333a48e9107a668ef747f0507ac3318cdd5ec12f935ef1312c6b2
z344be7aaa27d15938219e854d8472f482587e73148b1c652a0fe76c4a06d90eb433a5acef86de8
z05c0baae06e51f5064f94a3d25ece7461fada1196ccf45d17b3052771f94c012cc7bfaf2b1611a
z0d45573d89adaf759eb24aa6d7a6b76bd97f8cfeb552fdbe32580058ed105ce593e37d1ebc93b5
z6445024de04e374bae7494f7fce85c8152e256de15858fa231c651837f8ae3bae17571f8303e15
zabb2641cf97e7dca967e6d698d6ed13aa39c53ff0afef81f1c6b9c7a8ff23861cac79b09d07a41
z01a90c3adceee8f1cb683efac424e523f55b70db5db0332cd12b250c47f8ddf0c9b25a992f5c50
z15a8169b43118df357d3a4cdb25a4a6d0e9286466884ee4532b1051a334390d146830f558c8ef6
z3cd535932a3078a9f22d05099ecf2d24c868b56eb2e790cdd3203de2d35c2fb7cc0c8ffdc2a51e
z59eee0d67d4a2aa86b1286a865ea9dc8df21b46729c2508c1f80f9aaeac29e21794a3a9b470e5f
z5c4cfe06282eb449adb05ce0d813e9492fc8883f241ee31aaf17fa2f9d083e6bd4cff5293e70f0
z59ecd611d04b5a355065f59d6f35e21aa5fad713ea379399e0ee78fd94c90b4a3a15ddde734345
z2e70880b26fccececaae5f9384fdec3cb2dfa13ba18cbb5b7090b92e5619d397c57522033105fe
z76fcf5c06ebcf96de8b089c0ec932fa6b914790a12db270f747e35682d52d89d4c0ed74a687f5e
zc87ad6dcb80d97c6549ad56fe04f64e03b2abbf9e55818d792b2998892c188803d928aa43f9f67
zb7038e89620b3f97cdf8f26698cda962eede6d0930d12fb89e7e99e6828a60a45e43927cea5f15
z184bc792dc275c0664c75d23861e5bc2be73f6a02358be8bcea452f7b7a1bc11a8c10ed6deac42
z0d168da0371f381c34c974333d5efd77e0ff842b426f7706a080bea407317380eca1874fd89fa3
zb7cb0e7ddb5fd904a88a40357589496fcf63810f91d7b3d268b1a91e148caf5a9ad2f48ce8b3c9
z35d44a414084cc7e167c1a6f2b28cf6461eb3df06984276427ec84a6384784655388958565742a
zc3b258fccbb60c17ea4db547fd5f3f98d7a7cc8a6275ad8620a4884dd946c1d90d6ab9f89a4d28
z776205456e31180ac77ff84fcb230b4098d51d0e098f52d82fe3854031a39b53ac98c835e50145
z7e29c8aa96ea28cdf273177d44d653bd28ce94257ce24f9a334ba87273b56062b6bffca82f067c
za3302b296f6e187600554721854fe85002a853aff7cc1577f14a655c241537500453293a13fd11
z7e24dc741d00d064599056b5cccae96520864f0a6f2c84b51db3bc610c4c6ebcecae0ab552b219
zeaead9a59a744b22aae6c078fd075cc695d2b4d61bd5830a6273fe381445a66c1aab2d4df190f9
z6c74d65ba4513605ffa3c3541b1383acc97856b0e22e5d76c585152fb68ec5f4e257af87e3ee1f
z8c72edafa87d1238cb1de5b15a0175aace307fdb73b87bb201217737e001249581d2fc7db7439f
zd318b2daabd12cc52463c51602906ed6129591a9a5ae27d7dfd2093b62671350e958259a6e6bc9
z8dd14962d85b63de6ab0d38c67bc0044934c5ae61a7c7852dbe025ff817b43a965f866cd287ddc
zea36c0375d8f21896aa60f1a3894c4da5996dff09bf7b49e81e07024beedbd73a41a23c4d76268
z98d4a353c35b8a1829f1f5949bf36d0d6d99e9ef6dc80e674cff50c02fbf07757c96a4b00fe1f8
zd3254194fdf40184468b1b7770342cf1485005722a9959c80b7b66e47117ce0382b45d90629f9b
za2fd2b670a43bd90cdd38511397a5da0043f1ed6e54a3955ae69bbfbb5917b75fbcbf4eec153b5
zac0cc436727028e338d89696f1e49daadb96ec21a5ffab95e2ad1192f5ec6e50d8665a7373806e
zf6acd645ca8fabe09a38ff253600aced3569279a040abb2ec3cf1a8c98b97e4ee431af990ce7b1
z62c2ca1e57017a23b761d86299b4cc939c4cf227e8236953eea306a2d561e4c5f74a3702acb97c
za816548ba2dc34c9219afa86a4bc315e5bfcb14184fd7f304b280865aa69f4b6fffe6562890369
zf5501f760e5501802c4254c71dedc2771c50c7d7b521554bb5b8651b83c6646d5c669001f3707d
zc7c3db155d57c7bc2295670bf7599242466bd18b3951c5e4ec2d205e9a3980e03afffd8cb73791
z1f6ab75c000fdbe8a7d805a982045409c0797052bb8ad651922e9c89327d77a20e1b5dd6ddad7c
za2c59c150bad34f87ec4d0f172c20854c6c7f6aacca3c00ec03d15a6fc43651377c65011f7a822
z486cfb44e2942fb9358e09deaa47ce3e8fda3a3fe326acb141223bf4d481732ef338a0b52ac5d5
zb1ee991c40b37e3b3d007b11eec248b53402dc485f56e464b036cef14926769b36fd0213cc7af6
ze29e9d3fbfd62ea55e9a56196bfc404659f4305ea4e14c1deda45038944e6f039dbec6d6d71e0b
z4adfb803dec290d8ceed613a37b58e943fa22b3e7ddfdfd68b1f9a483b4f8bba9e8cd54f4b5586
z7c1356d6d4bd745dabcceab42b8291da0f4cfba1f8fb29ee78e53227a32a297b40dab4bc39875d
za38789e01a9ba06951c31b7019e1e217cbaaca1b0e2d0d34215d15a7b8b4f117b5931c574b9b02
zd11b14ab67e34896230cabed593f0c65d4aa2c8b968924bd85c156cf24191797d9775b625ff66b
z863e79aedb5a220223a191cb7874ec543c0a7a01cde59246ac1f5f086422a2a35b2a4621fba136
ze9112a6f3bb779e9c97175446e5ebf3fe50e3ca127f07245099d49d2b0ac583682d5cd1a469308
zcf42d991d42a010a52867117805a068182ee15d05ca58a9daa470f5b87b6a968e4066394488eba
z6623e69f70cea38fa50c40835673d9be997d75754336b2b592706c0015c82482dd242a97d7d1ae
zc39aff81b4f946697df61e38672d3f71f53992a21acefefe6208208d83f0231611e0126c64c91e
zb5b04d6ff71193d64574d7a4adea4e8a3f26445b789e48372cfe4db887fefc89e5558f6bc01de3
zdcc7a7af53db259583330362f08bfb6977c4c9ac22444f82de615220ce8a5161c94c631fb6ba0c
zae6dbb7570c4f06051260a7083a765fc3dba1ced0773b0f9031fa9502d809a1d8632148886bb29
zd37961ff9ec675ea8bf0e8ff3fb3475a896b99acb546362cf2b1b22253a09ee8fce4ce1a0b381a
z45d59c01442d31101d9d2c650c1c27b2e0d9fff4cffc010abbb79831d478b87060e5bf54b97ada
z933451134a9764da12a8845d28743227c7c843c22a781e1c103227be87abb7fb4a662f7c56569a
z2b03687e7efdcd81c769d9125853407e44edf9a95a198f643db9e45e0dece3ae2b5a5c9f75afb2
z9919fd07e2ed96d906cc57555e3c45bd1f46e153f0ecf3faccd3d0bf312e049b6692b7fed88b6f
z3abb59831e6446025e7b2bf9f2ad6008c9794bccd299c7a1182cce72f5c8cd6994b9e8a3ca0409
z858f4eef3b8a954b788ddbbe7133a5dac353e898c77f441f8abd0e31a1183810608f55d2f7e74b
zf24086158cf5d7a195c0008b7c3da639103375d3d06fcbf1039abcf078d93d82b1c83668057237
zc5a22f57c99c1a3d692a359b5eaa6d37748791792a8de82138a86b03e792ec4cfbe876d7730fa8
zc44d34ef8caf8a34b2a1e620f930cfb05aea1c42ea538393a00c631d75e13533ba52ff433e6279
z59275b0465659aca2a80b0470ef7b351cea9abdaf68f94d08d49d77490fa061dddb077bc0c281d
z9c2e5efbf2d165a3b2b5e22abdbdcaf4631568c47db6950cb4f9cd18885e8a9de0dc4c8a1a2b8f
z4112736866e6dd9d467fa0c2d1b1cccf3f740eacfec81ca0331873d7c2829a24e09a30d4bf35b3
zb046d886f1209376d36b22e60483f8b37663a9d89f1607291c4555b37b28056de4e250771be4a5
z95e469529e69aa779b5f984a6433c323215276d33031727f64ffcc841dd9060ad2003f445b720e
z2bfd5f54762cd58c1576b5b98533051caa6771c0c40b79a3eaece584da071245e70336f7eec80a
z6a7fedd646cb8e38b6dde9984dc94b554bf6d50060a9891164356104cd6170425d6f8f923264b9
zb7599dfa06690277e4852dd68658b37ea13542fa7b6061c4a56fde2ce2bbc64ad63afabefe795c
z436870c9548582d05f8e8b7f2dee99bdb528b95c7bf1fb39429393e8c8929e6ff5050d670eb574
z2d4d486e0637b1c88fdc7492a7ab9578f62b7f7559fcc9aaa35608e1a1320129475b34a302a691
z17d10eb0884c4e2c8fed84f8a4142557f51f31917dfff66ea19355a4b196f113a1ffec204220e1
zf4629e456378b16fd5b61c6b7f5c857757afab6d57b714e991554ba64fbecb8a8b444626f77db8
z5e2945899e176ffa08555b4b1ea3763c694ceaee2958475837795cc1ede843be7cdc4bf0d551ef
z2a90bdbd96512c4298f1c356e9e35d5292730124df22c5a1942f822b5ff1bbe9f5029bcb4ba3d2
z28be62058733035aa8f84465fd502de4dac7e3540dbe18fd5ca23c266ff133ae84475b599ee368
z14bab15d7ba9c61f4325b8e1fea88a083d0f5dcc7e501f41baf2186ce0c03c82473f339f892c48
z1182a3bc8c110bc58bc23f57f17eeddc914a4df79da8d9b7937ffacc7aa1f8b059d05ba543cfd8
zb421c325da2179b20c5bc2c9b611e04870a9ff9eac578c0a16805eda544d810fec91a59104a08a
zf8d3e98875e7380fa08e05104ba76d0afd304129cbb2b9c9d19c3ecfc0c779d8572091a47da16a
zdb1ee5ef4be2f1f2a6065d9b1a1987cc005efd7fe2eeb46c37b44c66f8c99cf03a833ef3fc2dac
zc870e960b4f8d6e458350754c4f1623bcdccf70d70ee68b866323c5493460d52886458b8e833e0
zb1eb02ffbaac22d546cba33d693184b0814dfa8f34172cfa4f299515b6163628072bfcf31ccb2f
z2c638a636f397b21a3ac40dd3cb68e39d1633c53df45ebb36dbe3314778c1135c862abc56a286e
z6a8dee2e661cdfbe04525d508ee8bcdf9df73ece44293f73157ec8ca443fe1991e14252d0c2c72
zc7d624be0529ea1b508368d728559bce016f6aa26e2ad0921a163501512b90b26adefac751e66f
z32d4c79b76f8904994013ad20b3ca6d2431a4283c3cb49cc5f88c5b9d4db3fbadd4fece506edd4
z51304dd65d11e4c729c09a1e1848156dd6973cee8a548399f941e9a04463304d3f05aa493565f9
z003898f4bcc0dd9013ff2fd4ab651360439f5f92adb00736efdb1c6314996d91057eb49520f070
zafc50f6cd87ba92d29d3006c9147dabe5f858660949fb01866d5f2d9470957e8295df3ac7a9e53
z7fedcf258f19d8b31b9a967a0733ded175b612bf30a9d00b6a240940d83aa5b72d0ae593f0584c
zb81d0b11f26c6505864e48c3a81433d7e637d41a75f66602d4c29b3d00f7b64897944daeb79da1
zfeec563e5d1bc5595d93bc888fa8997bb4ff55c169385370e4e3a426213ea6d8a242d963628706
zf4f63cee4bf5fae4c3516766928ae245dd64280a61b73c7d111e5a9d16d65b9813a7cdf9d4221d
z5b83d5dcb58f6552201a036b9a8e41dab85effbea90d3e3e62d04bff7a56d75a81551c17b5f800
z2e2637e9f41fc400a4ae0e04d6e8e536ac0a1adad99982f2d6d3ad66a1938b97a0913d6c86e19d
zd39ed214b525f0e82347952a40bdd0d546ad155db16364476b9605bf372e22e474636a6b641f4e
zc7cf70045ef23cc7ac48afa556a0c80f45a5698638738519f9f6b629cf53ac89f4ed5a70cabc9a
z1df0a57897d62481c2814070be5a27a279b0b5cc8059a65961d0d72945d1632eaacb9b8638d9e7
z3edc430f72a1cb01ecf652009de18211d888c862bc055ffcb4b91f445604e73a320a4e773f4179
zf84c38dac45abeca530ddb8257af8c75b18dc5015eb778919b608b5286d6e28e11739fb24da964
zec8f8a70f5b9c05d2ab0026aaa791a23845977889ec0f5875653df96f33e14ddd99dffa6f1a250
z748d0f2e88040866c9a698ea6d6b5a2e2b8711da066734737de659e3a65eb20ff0964914fd1b4a
z9f2439650dd5e9d5ba2a35e62582a8841e5a9f426b97ef33960601df53b8392473d2cc3ef0a81a
zbe2ae82d0eb3ad72c8400405fe245e509fcac1b2a4f31c2a7f76ca87ba2b472446f68cfbd9fc46
z9ef3d639ad07f5cf560a43838bff69c56bda069d2f3fd724008eef5bf0481a1aa3b7d819bdb39a
ze089bffa919d9b4a01ec55319784a832f540a9253f9cc8d8effc0344ee6a571a575a7078b6cc35
z9dc2aa038d101a72bb9cbe99302c1b96bbcbb1c99cd752813c3a9e356bfe0da8b152657a597e5b
z29ea20f159df47c507cf46abbe5639dfbd9d02a557113981ca6055e226212bc4be0506966e1133
z8764561541ef1aa97f145a432c8ec5de9b02865c882411a2c9992d62bc46ba3971116dfc0ec89b
zbf2ab7f0e765982dc294a52bb63d373c0493fe1dc4b641395df994c6bd734c6403ab6afc699f4c
z41a69bb11f85c56da3733413b60ec347e7596ee3132705a3a5f5bc56eee4b44726e27dba5ad428
z68fb96466688631984f8d912eb1be5b6169aab1cfdd98189512e71632d4f3f60ffb6bf265cfd4f
zb064dad19c5d5d994e25f68758631c911b28835789f3ccc450e35d2ce0309b6aae8503b48b814c
z3902ee7ddb99c2ae2ac1560a7be2e03aefa36d6125e73cc954691b725ba8199bba1d81d5671ca2
z10be79cb2b21e6c87a75384d29d41f2b71ef388abd22a90193e1e2ae29969b5031ad01303319fd
z280b493d05caca029ab2ef4b2a2f3aa02d977b71c944fefffa5d46cf3a65e05ab5d2818c7ce05a
z2f4877948a2edf6032c21b17c0595f271e3449d1a13bad5ce6d9f2e363a0570c22d17f62ab3508
zd59f0e3b1019924b95af4a4e5bffcca5de92df225390c81a51634523b9fdfc6d6a420805b0057f
zad8c4bdd6d477af21794e47cffebe81c57fa51acae0450a3aea1375acb39ac74d632583922a70f
zf8a51026ec8b667f487d55677f0fce0e09f6b5fd10ef3cb921c17b45ff967ebbd52ff9d2f05c9d
z030e7187bc4bbe4ebd5f71a50b5c80bb6db96e6fad117112db2a80a8fd7e7c160830a0640b853e
z2bcb04033658b5577a733934fb338ea4fc8be73cd6555d3e0ad32aa949d1d6a02fc44a3667d1cf
z226906015c5c5c498569237fa9f9d09c06cfcedcddc70382fff4fc32f66ecfe556cdb30bf65849
z6ed33e1cd22a6353c5250450f4dcd9f370b15441590726a3acb77239d3a74ec8ddddb57fc49906
z5c7f5cfc875586f122f2a9088536a452dbf009e8122edc1ccc14744248217781330619801734e6
za668d273c7c371a4b6f6568e4ad3f62bb42a67190ba99f573a30f0362d54fc527c94f844b66a9b
z00564f3c0fda23ef5abf9249a7bc93c89553f536ba89474b059039d2a57851fbad51112e335bbd
za4d4470b4af085f9e1e047c21454b9b44e5290da7ce0a47eb1a10e40d002a0930bf2bc6e028633
zc551d8c823a8f35f1891da628e95160b2467a61de3d83c1ec25e21fe3674e68a89eb8ca84d5a1f
z2f1ced60002cd9ac34482eb279d3dd273eefaa95746ebdf2159e7d561b9f7a3c8d6370983844ec
z2c42b2472d9b559dc50ba54b6329e420c4b8ca2050548ea2ea643e17b0221e820f6c4c39ae18f5
z10eb093bb4e4054755e87108c7c04d6ed5504272ac6f17de7bb6f0a8c94bf4c6a7bd247a27d7bc
z4997c8fe446ba9c54b88fd710168479c3f23c96884c1f7d68363eba0a732dc67486ced9e5dd131
z47fa9e6b8107ac21ac2d42bffe6e8d7d365167dc48a609a3fa0726024fec8407c4a859b340217b
z917edc7fdf498da31d0519ed923f83f6bd66127ca17bcfa9d568036095fcb5a0fa742465e32c4a
za07b84f7f71683da15674097f9d8f1e16bdd3450944d3e9db4359037fbd6f86c45621b6810d5c7
z9a4de6c525b2281ef59ca22484bfc870015873720409d8c467e8dca89120949f0bfcf4ae0f9a38
zf23b3e319fe6cb6cc13f9945da7e74dcc9999d4e5cbd3dc4f9ca505d0a551bbec180566b4409ad
zfdc43257419c3181df502a50c0f60f5b7d2bde11553f1ef6bba8a83639be2e72c66d422c241598
z7951499c08d8af88cf7ae658c4d615201514641c0be13cacc90f15ca08d540ed2f95908d8490ab
zab69a391696d4a4a87bc51de3dfcaf0909e98398c1c7e64abb562b4c800124ff2a353a4c46293e
z27d0fca2ab0977726c2b722a589d7188c47513520e4d4b292628121a696ace1d585d59e6821231
z833212d2fbc15b3c2911a8141fe5828bbd3001edeb289ddffb278670050209c3981641acbf96f2
zcbeb4e7bc8ed1cb003cd5393ee3de7192d2260ea82881c9f1a888fffa813348889558902e8165c
zf27bcca919ac603d2f0b09d1cce123bf824030bf50055f9f50be9fb50f2c325bf9d98daaec0c63
ze50516d79265fcd5a7b4904cd7455a7775efc98cc67a294bf4ed4e242996e9ab72466852fa67b1
za57e843c07483ee347aa85992c8dec9605445b9ee270fe29c62535c243e3de93cee1f51c3a4b07
zae1aa1e83d00200e815246fc91c5c052d5b7bd111d60ba3d40ff76f739b8dd4a4efe29ca442ad8
zcc9e5645288f60801f919d34573dda9ee618b83832986a530e1d83453957be34f7971e0022ba6d
zeefb7fa78210afde8b591de09310168b9058429ce9849c5e3e8dac35083a2d83c9923cdd1a6138
z49a2d9fb06680d9838f3666fdf84021cc5110d217e9f5f86ae706b45b31c443b79e7839974d1db
zfcafefde10a8fdbafc04a7c48cef4499ea7b07461137e19ea9db5efb692be744aa350fa97383a9
z926198e043cff1ae9e9a5b532fc0ca2dd39581ee7e5be976fdc1e5b23ff49b57ab04de9c669bb8
zc92652e9582c9e92ec624478ee06accd668d6953ed00c38816e6f838d38e0aedbe67808f5c233f
z53e60b7f6a88633990e815fb43e8cb337b0fbd7f3de3a26fb8af4610befbbbb9e093f4ed1d85ea
z9c302996fe7fba0fff2eca646f8341771028510f383c7cc0480f7bb09cc6e1af29b5e0736444f4
za0ee94cc732efa8239918190e59c797bb729882016dce8ace5018a1bf57eef496050cb98c4cdb4
zf7686c165960ba5421c5f16997d3226d753ffc157f9bdaeee99b5e9934d0fcc43dd5403fd41fc7
z32aed570bb2242eaba07a61270d2c6e46f46b57cca61e6223115227d48fdec6edf2bc9eee84db9
z06e5975edeea19eef160e29fcdae344f7b4a5e6ba7a43d0b90b8e32fcc3df3155138ab20fd17a8
zea6141e368f86dd6f5ab71ff7b2f8302bf66268d089f796db2ccc2e9a65ffdc622d398926c5bec
zf184f8409c7fd6c2d699f2590a4db9734e53275552363baad27a0bc84442c19a74a9c012456485
z9186b5637836d95e8d6ec76cdb3b555c85fbba491550b063c73778e9a14f8237fb20f460174dac
z55067d77ec3c17ff6ad63dd960678a31090f87179432d7d0acbd8a2bbbb6e5edc88351bf6ebf67
za1a0d1807842b01f5401215510fd2ff532648321efd962b65ff04ba58e84d761c6522708fa00ec
z2fbab99fdf378a76ec4b73dd34e302800043a9acd9229f0b0319ae8bfe631773e9a091f206d010
z9e6e94a2101bd5ce221266f32e9cdc3b3f58a7ffde775f76039d5629a9911233631c7417a9caf7
zd7a95d5394de43530bb37a73d46b1d4d34bee71f60d6557da56674b6a4664566dbae30c20d9257
zbe694f1bfffa74b9e63ed3534578b0c2d552fbce3bbbe939a6f4b9c73db2032b76e6b142904b33
z48e4f470e74a0bc23554229bff50bef2765cfb5fbd75d7dbad4a3d2d9f367294887c53eec36070
ze2b610855fd99e76c6574a9466a8c5d456323bfc547a71a78ccdea0e0ae8c31fca50dd1bdda1d6
z00552595ed297b63c0b734c577e1a8a1cb04445d65dd234d397befee0d61f39c6f19fa31d1bde0
zfa2d5df71bc51783659abed37adf468d5cfaa2297d1e20c1fa015f0f00ce4a762b86b003b1b40a
zcc91d827917ea52db7189cec7cad00093f144455e92c1493005c94c54e0226746b85da2efc40db
z286029b465a9a5f8697acc78f8e95625522925712b12788c7b1427612077c0edb834dfdc445279
z96f62899f5b6929013908baff7f3f2e77f55f44c5b8e37ac844bd6252cd1a099c88c90ea82df10
z636c4c69afd67e081bad4715dae93c95e10eee119171b860aafd062743760fca301330512689eb
z14b635a74ae735b5fd6a6187799afc586a5bd2a4bcbf448069649698d6f4b11ba1f9c138c0ed2d
z3f2e59d520de6d5d58ce1931894e6daca71e461119fe9b826bc38e772b171b574fba47b7de1fb4
ze2364098135c5417bec7ab75d39f7b7ac85b5704dacf39e8c14f77f13327309e2824c7ff36e64e
z395872d47495c32b850fb1e9ad9b1c824e461c009ae4b0b4e34ce2d87147d76d963eb303455a6c
z96a13d3df58fbdb434aaca19a19f47de22744017281ffdf996de9a6526400a2d68f335224f2f86
z5d2e8bf2b6f0911a6ea6cfb78b9dbbbd6d456c59e2b529cddfc2f19d32c8256fd844ddbafd5c21
ze54ad1047c63182bd31c13ab5cdcc5abb19c377a2a83bb86e892a1fea9aafb86dd2944a5eaa88f
zaf35b11c1dc77ab7903e9351ac271d9d9b872c61ae647246dce6607c4318d985cc6646a483786e
zaf3c59c311fd16639ce8e65848e14d2f11e2066cab9d1e19520c625c6bd860661a7cc1b81b1216
zec270d69715f6adc9bad0fec527e01d38cdd02f10ccc52bca28f3932bd07400e76a3148cb0eded
zc2658bb6943f59f83a7cf64dc11fed44a0456be4c6f87bc126c0e68ea8386cf60dde86c0680ed0
zaa768838006ad765ea7602e57aa66a2cb42882d72bf64bfb4b8450f868b2d07ebaf4d7d567fd7d
z138f5d065a890e3f2eec1ee394d9172628919acc4f8a793d9aa0a66428aeeefd2ee8df76919464
zca0c207e8f8bf440b9a165ee60e689d56c424d38f225ecf182e7da442125bfcf29ec1537b4f1d0
z8ed54ca80924739515a94aeadad27cdb0185cc3051e1a14ddc94b4b82711db256a6550ef51e013
z0941681e50ed8d50ea98e43657795f2d7d0a0cb6b70afc24a0ae5d4a092a48186231f923193281
z60cb38314fd07b820d222d81f68c34ed7a5a0acd649183aaae31258b509361912f3bea9b91c8ec
z1c91e97c9647527f92adc26bcf6a539529d4038fcf4a014a9cfdfbbb016e58f5e3de0720b968d6
zcaf824132520641f8b1b8a1715495383a1e638dd1a7f39eb019bcdeb4e146db056167eb454220f
z98275516f521e9540efa5657ad0ec87ca4c1cce8f22742e015e21d72a3d8176a21b95703faa70f
zdd728e61c8ba5a9ad25fec29f5bf225bd29930140a0fbadcc3d0345e0376697c1060fc9ec12e87
z7077b7a7979477ed78da5424ab58eed914ec51b92ff1de42d83c8ebbe7e5e091db81a557703834
z4ca5306143d90341cc3b5e294f8d10c8597ffdfd42911ce735393fa6831f9985d4057e8cba6229
z451408acdaa5ad8329825906f563e411bd1f77c08ff9bc7fd9b93ba76bbaf1034537ba5d2f1024
zcf2d0a04e2623c022981ec72da9c40f5a09898ba11d30bf0d85b1c4ea53a3b5fcea6a6b43f7445
z8e9b44b0374500b0c8caf6394cd15fa23abaf48616f789ec8ad54bb5a481377f048ee784467b19
z75eafcae0e9aece3f5d1b2b586fdb1a3d57a767865c30dcdc1376fb1dc56e02df008684d128d6d
zbf3aacd1f4e0b8df23d194c8bae3eeaccc7658a2fd469d0fd0738ba956f18cc934960187514366
z59e71bb1b9cd053708f5c86d90dd16f02ba9570523040c68862dec932253100f04f1cd115a4911
z0eb66539090c3728da5656f12bbbfaae62f1c8b48a296f90cd933dd26c70076258773197e24f5c
z356d59c0d705e64dcd1c4755fe89076896d61c003fc52f2288cc76e2a1627ea4e64fc1a4832c8d
zc2dc7d3f1ea9a1853b274fb905ff844994d2be7d081dc625910a9446290b3649ee43980eaf454b
zcb944b80e1f6306596ec220352cdbc1d16f8926f45f7c88e842a8422e75ae43734453e3cf50d60
zd835f92d8c10744b47261e05c376e6b420ece917824a4e7556243342635cf022ef121ec3e3e209
z1be4d3d0f4b2706b44a8b645181715f01662a8da1e72e5dff3e37406634f067abace0cf3ab73dc
z2dabe215c05946082d4b1a7ede92fee2c3c9c58d4e4951375568ee9630c035a4e848b03b0f6343
z1d386af966f3ae273bf8e7a720e0f085e7f26fbffb37fb1dfdf2656c266e60111b0f6a1fe7cb9b
z6aecb372770dea70f57452a20bc9022a30583efa5fdc6cc73ada0c1e1bb0861117254e5521bf52
z10192d492c5a65e773ac1495c29f4e9f970594b432932a890dd9435095367c491e25d2c26fd06d
ze51527cd13cb7bf8886252edde3b0d1e2f85db34e221d1fd3e04973d4c9e842b8e71d918281dee
z82b5f67019caa4354c23d685628467030ef15956fe5307110c676a594c94e26069438d60b664d0
z5beae996c900088ae1b7ee0ce22abfca0dc5649bf325c6f29a97744e3fca3bff45998d37411d03
z37ec613573a26d050f979df74aa708eacd8e7e26c056d2ce43dc1d9332868a46d1e7d11d96d72c
z1bb51f1b7ac2ff26fe44079068b4f286fb3bbc58fc21a90c94914ae8b689357c0de7ba480a6d4e
z9f680cbcbeefa167b31e6594816c7420b3a4aa9efc4bdfa69a61bc0261eed75e06f4bee326cd94
z44a9123f02b713bdfa95632db0cf7c8f78c213a2e342b5f19f5abe424e59cd775488e212e11b94
zbcc0002a220353de0566a3e8f2fd6da44ab123aff377110e01eadc46184d7d309c6fb68481103b
z7de430fcf9d322ef24a7863af3bec07b464597f4d94927a805a77524d7f40930d28782300f6c6c
z639c30bb367a1139b38e8b4cacfeed240b6f66cfb9b24978806ac1e90e087d0218d0b46345b37a
z1a40e51c0b3b9ac8b032731d95e6aa1d22ff1976b41f7ce60bc315c2b8d429162dd97c27ffba9f
z0784752a16637cc427fbfcf1e2ea46c033e28b1f73893d3b7ef363a1c4c1863019b2dab17b941b
zad918f9e1e04191d91428f0c0ae6020d61c0850ca8313d61c0f0fed6907263bd85e01cf2c4bf24
zb1c74d6e8f6efcf52fa95f51c98f9e99f8b67a9c0214ff5fe8653273968bd15395e1a46da3606e
ze9849aa3c3ecef3bcde44563c132172eea3c26d81f8e3901de058416d3086260a3a8f4fb493bdf
z451e37a835a9d7b99e9424154ab46ff73cb0819ae95d4104ca0d24a80be545bdaa5d927f0bf458
zd7efa61c11cece29fc6bd3cc2588e44041f996bdf676c97d9f058fd5ed758ec87eb98d4503311f
z2690a686d35d61cdcfc9f3919f794a005c66fad8e534b8584d81de00f81141aab142a66b445b44
zcb86e04d27dfce0ffcf42012d84bbac4b94542fe65700aa37d133906fadef44544eba1de1956f8
z315de38e5756a84c80038ea874b16e26fdf237c117cab585e765c2e044f9b2bfa96f1607b7e0c4
zd5d9e39d55f23542c79f5ecb4e4fd31aafa3c9f4ded5a8f6539454f19d22675ae4acbda4d46344
zdf9c4d9bc324f612cfdae0775789492ae026fd5a19e73f14c60623aa83fef6dba52698b0fea7c5
z03fc79033dcd36a144851d96e3b65b0ff1446cbcea163d062ab9c910a65e9aa91ab3ded1c48798
z94f73f17ac80b5ed52bbe84ef614e4cb8499820494e4a518b7118567fa39779c2d4bc36bf1bb13
z1d64a880f03e73afc4e75c601736241c1ed05035f059cc9e28a63f63b6701f0af9bbf1002d503c
zdda3c072ee021d739455dad6924e12021e08b301d8be4e5abae4d4ea4e74c9018873802f955ebc
z8c0b15a3bcf93c13570ce15964f2c22032829cb8f6c30e744952170336a08dc7d4577b8518441c
z5971a21740711d395b6d335145584e56cf772e9baae4cf27170953b8fec06137f8da22fff1d42d
z14510bec0b53b993cb8b3eb9d885acc697cc783fe75b91d5833d2c72b686872e051bc952ac265f
z82288392c7c765867c824fe41310b1d6bc18b3bbc2c59e107e55fb19a9026f00efc655e65d5a29
z74401549ec7f509843bf1b7598ccd0fa27d996f1143dc4b109075f7e984c6a372f6f5296ecf6d9
zbdd8912c6b2fa665f5254bf7c85db2446bb2aceb94c1a2f7b96889c0a5b3e022244c9ce490f84d
z0f3a534e445d5af158fdc3840bba492f1501a29b4e35805b7ff4917c56b1e226725520ce068fba
z33c3973ae699cae03d9c049ad7cf01abbee0032227b13c72accf4a25fdec453bfeb799ab77ca71
ze1590ccd25c97cf8491b370ce843d67ad7a8acfc5aed4e895d1dd24eb652014adf6b5b072be6c3
z6644661496f2bab34eeb57d714a78903625ac96c6ed8aa57b3f3f3a4e6e348ae9fb7e4ee023695
z300a97b487d766ab4f0274276a6718cd09e1e5b4d2626dac6d4d26225007dc0e3531e82b2ab8a2
ze0aa55f861ce1601ac6a32d51e2728f06d34fcdd9344130b027c3d8d13ce6ce55ab1763e2fd34c
za7412ba21fb9b3ff3b788c2d9bbad267d959303613a2c40f9a8afcf7b52195d6c9f5155af99743
z2272d60673c5bc4ae08564555b7d26863fbf5d986733ed1b6f745bd58684f230077055ccf6fc3c
zefa8be46703c6bc952c4cb30039666f229156b1a51ddc2f6bc4420c6f56a8e5ee6111c63dd6637
za5c69a5596db91e9a3833288b714ac843d03fa35d47fa6c20c14a75111e0dc697f6687e7871120
z2273c057225bb50bce05e01cb6609c746e2ec04c350f9a0bef6b45120cdc769b407b304a8923d6
z4e1f494f542b567fdb817c6ad77de6b80b0bcad8e4c4c24899eeed39dae966d2c1d16516ed53b6
zf96e7b80208867817c2dc77d010a0682222673308641e4fc3bdb2f20cb3d1964371b58362eec60
zb3112c7cb9e256e7cc7e60f2cf09b86cdcf90ba61bc026215a5f6b297857f82a646e56063b33ef
zb2aa1309c50a020e7155960b0125abf72e6855724d61af9dc5fe08cbf0a62cf059443c4c828173
zd067daf3b5a48678b89efa6ae649b168547993d674c4f323bbd9ad5dca42366cfc7a8ba951f416
z6c37bdd93e317818fda02331ce0bcbf5517e04c83a0204aa363f95e9f68b476f861889ba37c5e7
z721f2842d6c620a013409c1674abd4f9e7aa924f7742e56dcb7804fe2eaaed3e4bd1d8dca9bd22
z1ba107e170149d5c45748f0d42766eb84ae9082f796538fbcfc06550bb9bd30cd4d6420d494da0
z247e01ac4bd212f4d3f66f9455c6eb6ce772da4612b38cf75993ff0dd1d1681106d024d9f2d42c
z547e2868dcd0cae3513e5e1e437102a472927861897f2c30ca6649a070294fd430aad9319abe0d
z906a2c6783fc9860d029bbfabce20715612ec55303156957af6ba2bd25d1c099b6f74861a735a7
z3898b76728dd9c9df8b3998d1b102e024762e690a7c7f35494c10e1de6b330516f689cdc4ae439
z8fd5af175ba1e4af8b50a530ce92077badbd1784db24d7042d720f05fd4de0d886f178039906ac
zb34d695a6b4a8d824931f147b7d3a810a878a40b2b68215bc78632e449a73b4627149f6a1d16de
z108ca7b58e856d2ed772c178f88e8f853bcead69d8c564e5bcfd21ae748e5d4190918eb096ee3f
zc0d5dd757f5548c100cf1ce504efbf943934e0eb573784bd36ef47f5e10cadeacc0b40c9da180d
zbdacc8e9407c36d787a464d70da4833ce689ab810f5ace0586471fb793ba161f42299d694201ed
z93ccc921ceaee199a79e2f6b44260afadf6c9b403fbb5289d96f7ff2bd97cae2263e100a05133e
z978097d0467995f1f8091b979d3ae5323a7e9914fed2078a7c6dc30270027bb008eec8c4b6f5c4
z055959047a391392e0ea3b8a4fb4fbc14e5b2ad41a5f62f9ea634c0d878c1ab2d07ba6948478d1
zdef69dbb654a5080167d955ff2b6db11a52ecf0d37a4dcae545ba275394d63a0aff255f60d9fe3
z44fb12f469c3084f669162a9e5740535c6f4e4620aa8808b71a1c550a391daf5656a1cd025c4cb
zd4acf1d718093cbfb39c360ae542a623e7951173c7c9e4bfe1e56bb013bdf5f2e3314d430abcc6
z16262a6f433f7790e4e46255cff1e62fb922847dccc84ac8b581cdb2176f0fd8531c92d49fc4a9
zde9f7c84b9df996e818e833a1a0120befab9ac6380c5b81b27ec42e975e5c4fa7d2a3885d70d7d
z60ce790db26e24d02520e21fcd8ac41ad90badc8410d58dc01cb44afec12d6668b939e5665682b
zb724cd6d39688080ea4141a8b9fc908ea3d5db1e28b79ad7b4bb24c5f2327c346b5d10c3484fe9
z00005eb716465f8db7dfaa706b19a93e910fc7dd890f13bd1d75919ffababa6d39f8a762b57bec
zd42f50876382098383feeb8652ff383950279490925ce13c07e78db5442f143fca5af0cf8bfa07
zbf680749a5f7e3df052c03447691927786c2a21a76f00c54bdbc2a950afb1bba13ce68667b93d8
zecaaf86610c5562e8292440697bd9ba8021abbb4d5298b960b3824a5d9431edc24faa3ae1b7f5c
ze28b74e338721183ee20a948a529770783e756634e12d355e4cecaf5894941f6aaba4408244aaa
zaa7f56c41a9e08e8d3db83c1574e01e62cf13bc0a4e6f33e74edb3144ad44f899edecebfe2ca5e
z50d1ca4f19e0a6e888a4f77395310bac88ec681f8c62f0a70e19beb933634e67b3d95a65d2cdae
za1e34b2229a1ef13005a49e06799c49c0693bf0cb7074db65cc59af1cc8e3b0145d97d31dd21ce
zdcdec98573c282467985474cb2da877a259aab535591fce6eb4498decd8ae044c5038dfd8336bc
zf5147ad13eb0e33ebec83f102152f83b431a4b3b38cfd6231e070ec7cddade10e06a252b72e307
z4f92878b1bf37a5a222c223c7826e48cdce881fc188c3f4f91b564e3b45d7a3489302250d13707
zcf4b8ca94d1a7644b53be27447cb4129e1c366c2badcc19a92917c5e3a27bf142af35e9f4cd117
z44b762cae5dfa56a41cc3195a7d6056a21b7b661dc9e7d64d9552adda99eac8d621b9c43e94e62
z5b53dcd92edd3df398dc0b1e39b7790c64a6e404612c99426509606e3c6dfdd98505c93632e3f2
ze6bfac5230e6dfa928719dcb620b12a34a9d2079537a49c00455fb30121e6dc582bdea3d9d1295
z85f695322f8f0565199bb860dadbbbe1af67b18b10dad49ce4c5fb9c33c833daf9cbf6be3370ba
z9d021bf58dd5361d46bcabf4c9cc27e714062c6a095f4e562b4ee9a680ea420bff21c4c71c7780
zc2f0bae9aae60a959132ab6dd77ad02b50e2483294e641b4e15f82c46cda2650c9dfacc14add0c
z415b20872a764b4176010eca0084963c32dd270abe3a0e6c3501c08fa456e34b9db1a60ef16a5d
zbd7875d78adb94abb9bea7d8005f333201cfe8073d8db36493edc2022eaccdcbc23116a1837792
zbba0a22a5afe1f8a9a42ba0c77a76f145edbd41bcace333ed59e783f3e19160f6f771390d8cfed
z117fbd153780e584a5aa4d39d6fa90236a574ffdcd62e19fe61d9417fc2e8ce47bd95b7fafc8a9
zec961505db12636f0a0d88fe4689c4d1bff9bea2d8e9ef073b9ae0856759eabc879713d2791a02
z11aa4cc87be9ea4606fac784fd44ebf272e5b057740eff6b6b928e9bb79b4ef0245961418d1091
zb18db6f4e6d47dd2d24319c69818e69c74a481df2b0433a2b5d5499ccc85d9f77905af9a9eff8a
zd2f561caf988f07797e47c2aeaa54dfa3681c29a4d9e14f0ab7592829b420bf3adc558e6632e21
ze3a1dcf04ed28d17a49a3ccc755f9a6ea941b066dc1047d103fc1174d0582d143216316c7a630d
zcee70b8349f8fe87e13cc1c16df80dad65643ff9a382956ea0fb5286e93062283886531c1e9307
zb6d01ed05cdf021d0bc534ed0e1e4404494558bb8b2807a8771d8b3d56be50ade0834a335430c1
z88c5868a34a8eb51026d359dacbdd49df34a86f09fe7809309ea8b949539c7b618182c15edcb1d
z8d8ee643b8aa2edbbcabc8b6e20ef9c40ad51c61fa1374224a50ebbe6b3ebcc8976093e4b2768d
zc4188f3c3a3c6a822b013672856ee47e625b90588f75bc54f25e86275eaa26e003b7456aebbf48
zcdb5c98e24508e5e06a25cc9ecdaabad634e6ce378272ef587ce6cd30448b9049d14c8b540d254
zf249aaa0092fb7bd8a1992d86fa1f55a41181f60fc2d7c6c1eb9225452430736759c6abe6651ae
zfe7cc553b7486d3d9b423b37db0ae6592fb9c74bf2f61de77eb5b6eeda6fb125ce05980d90e38a
zc5608a378dc00867537656e450ac06c1e300872840b3f8fd5eefdc70448982f8c395a2a15cf222
zdb3733fd460c4d19bc782493e1651f1ad9d85cea1543b2ce708545eaa550fee0c17be97e35ed75
z5b52963d71f356a98d3999607f61106c03346394184d846d77e23d768fe5aa905cba1347568e44
zfd812258c629d802a6abacdd0dac4ab7489c63001e0326a09c2442ebb49617eef14d2d9100ebfe
z12ad9c3ee0cf69fb490c252fab73879fc0880c9467c57797634c6a8403bb6a16d4b50a61c66fac
zef07b472fabff4676c303cd6452a5fdd615aafd256423f9eb7092ed5f0b6912e1ee061f40ef534
z546ff7a1d64d2ace7fe5451d424b4c7b621b1af4c0803f3919690f86f50498e4cba7a0c0a05400
z6534b8c5e15b5426944f479e9bc0d3b356444027f756eb1a9498abc176cd8a49c755a8b63c83a7
z7d5feb54a6f4be4a5d4ebcc28359d5cc90c1fc6f8d64fd55b71b4d22d6060dafe7fb84bf01211d
z541c86b810b0da46222fc2e621023a862e243917fe7a79176cdef01200cfa932445e32bc258401
z97cd096d29b07949c1a107942c3bc5a1094f9de120ac8e5628b4a9a720588f89613ef37302eeb7
z97c8fb2c2e6d94b45380f683a0ebcb5263bb04d4fc248e0015faa8ed220e9c1fdba09475c7c633
z00f0cfdd801c3ba0d7e7796f285c659309bf75d398f8bad4570c329a46962017db9d3562035809
z352b7233e23803a7611fa42c1ff91fb50cd5fb3452b9b04443d4001f5861d4b8a5424915e70bbe
z5f42e234c7f4518afd380b92673b68d18906e4e25c26e4cbeac564830e55faca20057252a5df82
z9e05ba2cdf845ceaebb3ccf6ff3d7896d664ed3c8e066cabbc2c9560bf92748dd175ada2f56826
z6b910329aed231bcee80ecae461f093a2d29bf8192b0608104288632f86ac5d74e29109f8c6787
zaa7132c4f874c97eb494c5b1c5bf1875d31264cdfa32b8a3a339bafe6fa9c7e2b05452b9ea656f
z957cc87d83694f125e9fa40de51ec0f3cfe16bf1eb82e3779479784f5426bcda271c585f384c86
z296354a43926c45261455912adba79cf25f055dbc9fd07ae2eb294804004ff53881458b81b268e
z856d9d289d6a56758a1bb69b027313894ce7a4bb3737c4e59bd36ff17ba77c0ac4445ba640f6a2
z900a5522620b5101ccdb3db8471d2a9e8eaec804d9067a46f4afd6450522ef9810d2e1b0945094
zec1c78a606950d63560496d0a5357a124802c88482f113e02c2a0a9d0fd79d55b61d0137ec1601
z87e23e270d15ea9578d96a602e5927d74dd2c71596465ba45519bb19440afb12d2523695583d81
zd23ccfe3fec285106829575b8dd697400916a8dd59ee6de001c44f0683566b4082b6992f1c879e
zfb492cf3b77a4e19d2b03c9ca9efa2efb13360fa267e11d0608cd26b024f75fd41ad269ede66ad
z9a565ac4fc6f53c5071aca1babcb71511a2eac8f10aa7ee692713734a71caa842126feaccf4c4d
zf09d85f5bd6f8623bee4ff3296a068ceae86fd750521d59e4453bbf6ee1cd36e8754f326251e86
z25a69674a370d4c372ca90fdcec46f859428ec5f8f4364032cfae870c4afe207b57ba413fac58a
zabc2cc492f31ba7ed183af3e925d052237363ef222a92847ddedf26013564966fe52ac0170a8b1
z8616a6749e67545daebae8d095b0f646d3dd006a6042d601543010c568255a58ed29feb6200ddc
zfd15b60872f020ffcdab4b3f09ba4a3a0b05fed1f1c26509bc1e436275bd3ac82088c3f2efe68b
ze32fc91ea53674e01a91c2457e54461c99936d2de34f59aa717cbad999b8f024a5cde4f775e7a1
zca51c24a7959444ffc26748266e86457ff15f4bcd3d9d22cddabaf1a5491eb9cfdb4db5eefedc5
z00c4ab3192329902d4d62e74fc0172862bce1f22628cf46adc0148cdfe896a5026d91117f10492
z21cb3b1b5e263de9ec411b64c0ce88454eaa1e03226a300620525ebb2ce8723b52a3e453df63e5
z735f7d0f9a816530e2eb85671c9bd910698c2e102e24274cac0c4eb5d1aaccd934aec267776d15
z456b1924eacee6914497e6c12e23cfe98155554283308c353a936cdb5629f744702a2bac53ad74
z0701571fcd8add3202ba16d045dc8ca88e4fe39cf06939cfd60c7859ee4f3e5caca36a2c79bbb2
z56098a8f6520773c175c1b755140598432fb11577b49b53fff162face89b8143d2f4f14ac2937a
z1a7a8c630b25c05297540798a75cee5eb8dcc24cccb6651841a45d938b0f039c095242b934e9fc
z08d73fc41c10aac2e1c54208cfbaa1eaa30ff9e67f2cfddafb50c460228544792d16fb8fea9630
z1d6be7c55574aec65b96db7e4b4270e0c5f0e60a2ad4b27b6d86eceb0312a7f5285cc6b9a74739
zfbca6d90a075314b8946df0c2bd45ae0ec4207fe44b44edd8b378a93b1a542cfb85b7fa8f8a342
z0f3e3e37862e3ff2f40bd38b06158d7c71f6d66920b34e9439386debf3927c78f3e140cefe3420
z83c611ae13629473903945b7644455135ac81c4c1bbdd69403082204df30ff3b4cf068697eef8a
z60f3e5d1227c3934c4cc40a9a6f5a859c2a51e0cb262e14f32d4efe1f2b2c6852f19eb12cef8c2
za7d1cfbe2bc44833e2edb62a5616a68f5241b7dfc2a935c932a081e00e7029a460bd3d09313e0c
z65ed82cfd0a20a07348ae88f05f0a8bd32c73866d7fbec35d8a6445134f0116ca808b93396b0f8
z013a1dee745ad8c2b48e5df7142caaadb54b3b48883cf67182e34f953f09eda14b7506be23a9a4
z10df1ac65f2899c6735a34168532a58276dbe5f52be8a2658cddb3b75b6536a96eccaa8d98ff80
z4d7b44e10415b61e281ddfdeb586fcf546e7deab7404b9303a0afe8e37f894f8d4b162af62ade7
z71cf8e1a3cdf79253eef9e61ec8912e85ab90ace1bcac419ce5e3ec7e6b79ed6e2b50dde52684f
z0e6b7ff5e878a1909522f0ca729224aa2fabf180dbc513b9df07c2d15cbd5da768c4e113a35032
ze939d5367b6580ebb93662bf0f9cef71e4198400fad2095956b909e61eb23d6727130bfaa0bb1e
z5722ac850b4d088fd8562b9bbd82cc29f629f33977feb334349fcaca03ed7af9a4219c9a842e35
za18a955d684eb79270af965811612ca0b92249dde5659bee98bde3757a3d74d80743fe3f59e8b0
z79c9192045d5a56dd0a1ff67592178798060403287db87ce112f5fb7a4e42090471a019f359f75
z7158856c6022f477de9b5669e8534ce7dc8958c99c5419414be722dd04133be096198882c16663
zd0b5f62767bf0ac72372d7a6d113534fbb5619c41052e5ed40e92f77ac23a61dab8a25c0260624
z25111ecb964b3a20148e787e9f17e76f2cce7829aa299050b14f4d3d703c9a5aee5a1da8d5d476
z2e20852d0e813faf2e6fd344b1b0e127c831a437f6155f8b1bae9b2c26cf71771d0e63716ea234
z3fa6b2b9a7324b8d7842f4bc3caa37a362f1d106064cd7bd5d799f8cfae46afcdd176bcff6c810
z6e442678ce8e6ea73a1c42204df25e4ead8032a74450b8214cf321481c9577e228f8ad69bff04a
z14829e39ae476315657ae69bd1a557bad5b5516291377ad481df2a83f1cda3a906480ed004e9a1
z1695938dd7b5201f4bc40958e64a3216ef2e1041b2648d3a3ace25b6d21a858abb2bf43a569840
z971b36a3de821c87c307f873faef3da21ecdd17fe418cb635cefbb4c678a4294595f58c4572c54
zc17d33b4ee7e7674d108fc37ddba8ea994402e0f29ea9b8c6bf8e95055b17de2f9a73633173023
zd0e00c424a1fa5ab4d99776fef79b1d0dd90d6a13b1fedb2f2761d97c0f32fa9e65161251ecbbe
zb820b8876ecaeebfe9375ef2ada7ae05ce9b4e8d7aa9a988a6d0147d3ed1e9fb0c7468d1f4ace5
zd7b9f12bfac7388f1426d42be2cdfb0c02afaa0384125392ae907c90b3bf637916252bce1aa5c9
z0dda75aeab885ecb8ebacf6cfdcae65b5707de9dcf162306ab437be3e40e63139e5deda3095bae
z06f428b3d4a90c4ef90bec33e742c7627ad48552276d098dbc3904d5dc1e057dddbcc1b2e3e6c9
z58452e8a884fb9d6b73622d87a1ebb1747afcf01fd067c96822126bb5623fb08a64bf8af37bc73
zde79532e4daf81780e2182d28f9bb1d0d347f830ab1de2449d53c7855abae58c4e8ae38e8fdb88
z374823ff76eee7b7ae1ee7d92876c65e9d8fa8cad9f709168afbd663cf763d7b23e6605547f012
zd8318ee95f5a2ae6fd2b12ed9c58de5adb4cad576578093b6653d3e1b24a594d3321524af40691
zc4ebbe079d00903e1015bcdfa429e751d2e785235b9c35c288c744c74adfc9141365c82a0af0ce
z9fe41a072a1619c4ea552f6efc9a6c391ef57407158d48b5d9d609f678eed4afc3f48cacdf60ab
z60e7ff7ace0c03507c013c5919266c797e2f4e22372541d0482ed099f7b6215a189606d9c35212
z9e74b743c28244113d9f783bb87715fa1d9e5b543c3b0a0d545a5f6ed063f4978848eb5a37cd9a
zd8588cba8019c7d1924cb441d9ed4522ae61f204eb9b689738f87fcd5274321cc9ffb2b17a44dc
zbccc30960a411edbb355b0013a0b10f5eed2c9fe0af9a7ba8e941999dbabbcb134b733bd9a686b
z6754c5f56c7569c58e56b81bdc579be31a1932309a6d59c7c8e4d45bd2df77850cd8b158deef14
z39c7210a73752d95a132bec268c842311eaa880b7a7b8658b5a7efbafafd2e44175f058560fe78
z300fc84dfec30dd6bf991d563d4f517d071b38008922ab179372c52080015f7dfb6c2b9bb1200e
z0dbfa927c1f7607936bdd7931a381694a5d9137aa79979109416379da9095263d527ff964cb6c4
z4ae241f288cebf33342bd2cfbd6ad60ca33bb220c58df498343e575ab8afc741b451c524934798
zebfd0b3eb355f6fd62bdc377d68e6d3cbc088475ed1f5e541ab8e3f76200811003609202b5bd89
z76c8ffa3faba861fabbdb70695d279872021772b4940a2951d38cc125b2fb79f462f612804f671
z14577b3fb05916590e5ef28ab860e9a71725252633cbb356c9e9fd8b091450b4d57dd5849a55eb
z8563821e5cd2d03b4673617fc7fefb2eee2abd64d9ee26d43ca6a9eda5779f51b3cc4c789b45f6
zf9d56f075a31a0ed47d2738fdf4beb88e650b8b794ea77c870b766ccaf0d027a4c5cd70f0fc7d4
z5caf4aa34fddada73fb134b981ebf3352fb3803049f1e0a5d906295ad343d87b0a65b35d88c73e
zb96664a7d52ceefb8640033c821a42c277645198204fbd4b6dc433bc1d97529209f246aa83d168
z4419b90940f9831de681bf22bcdf6092dc2408233aa6b0b7412ed897a89c1015de6d3a330d7cf2
z1a013ec8554ebd057cc0c50bc703134f0d81d51b3cad3fcd2d601b0039fd46c82100e632d68ebe
ze8b5bdfb776fece56c18671acd0a628d3aba8a1d07e8a397be09fa99127b3c41f83f46fe7c2816
z8a6d37e8ead206de2dc3c1da090d0164f50acc90ea3b50497252003401ed881308e704255ea7f7
z2b60fff125edb656eaca97d6c5b67ef5b0ac63c7966da482315858658c4e1f21a0f37aa864685f
zc6ddf49fbc274d27aa9142cba029042c52b41c4d02561e5dedc00f7a12bb310e7b3402f9f3c6ed
z5fef5e4a725b71df32716c10617a403fc5e6a4549159dc587608f8cacf31538f1bcdcdd782ec63
ze428456c6c6dcb5ccfe6a73b7f79bf0b0522decd4195d43347d56940058c800a4ab6fe3df7c49b
z5feb19399eb41527b7acedeb078b6a37bb987c8b0e5e01986eea301a032ab7478502ec08926c72
zbcb367697c13145b355191d3ae8dea0d97764fa5ab0f793cc4134e090e377c99ca2a2d73f04556
zaa37533a64583bb8ad795d57e96b89aaf1fc84f461dda5377595ba1174d7438131841d1a735cea
z21d9221d3edaba0d6e6d9c3f04e984cabd98893809177fa04a93d6f2a693fce7af861e1cd5011d
za3d2528434e353855b759466b8f2bb481264d98a0aa465aa8a957bf214230af2fb056360ad03a9
z1489ed4fb5441e19ab12b76bf77aa8d64d3b17c2153929e8a23219b2537671c77d9ee33141fa97
zbdbfc9ace0f17fc5555873f183a3e8e8d81062ab4c989c8042b5df4fbb2377a1490501172227d0
za58e9592b77292208bb9351c9d98153ae437cf3ed34007280ad5170a9a6ceb2fa9d957ac78a2f3
zb1abc215159ce1888d7f72a2e827d027101a9b4351fe08585dbd0ab60bfe4357da33fa8600af74
zb004b853a59bc133d716a24bb41d9d234705aca62c66d6e3abdd7a83a5a46b77f9ff4d478df79a
zbd43429e5fd6371ad662dd1464998db08d3f316845a6ceac9a9b107325eceab4ee066434468eaf
z2c477e8029d94aba5e9647bfb6450ba07cdc2dac53630ea9237883ddc2c7d2b60183cfafa8c9ed
z7ab6e46dacd12b64f2b7e128ab3763cee76c4f5da9cc9d6c18ac3ee0fb7eb13da59c2310035089
zdac14c5fa3d65669806124b139abb320f1d30ffab65897941414a60071acabb366d80116235979
zd9471fd7e98c8a893e5ec9e1958f63d031e3922fde284f94621e48dae9da7842429fc7ec00626c
za1a908dd33bc5f23d4d89649cffd52bc9038ca7cca21a348d8d035ed490d70a1ac1e08f674ba93
z60561a0d6e36677abc380b0740b964fbd5513f462ab7a9df17f7f7c2f3f6c64a898813451ca9ed
z6f5a56ca189eca968dcda72fec36eb1fc0635f71faa77a1dd26b03269ac5abdf399c20b8f398c7
z2a8fd7c174a252f889898f56f4cb2667fc17869a1657722368caecac56c8554902be5bf2e9ac79
z8c0a660cb60577f57b3bd29bc87326b2464ccfeeec1194098b0669b287089274fddbd781a1a7ca
z483d620879f8a8bebe27e862c28946be15c960679b381c0eed88111036e8449d5875ce90504418
zea624b83e8b054b3799902fb3cd4d042ead9f7bd45c29a245c3cb85450df7626380b1e2d44f12b
zc0f02af1536146e18e3feb5cb55b295ade6b067b0e7e9679e4dc1f50d62cc9277a51f5ba73a704
zda09a09f3d3f33bcdbebc06a4f6a5c3a02b7f29472e80d392fff123626b394332dd51d879c37e3
z46bed7b356fb05b823233fd2ddf06a39f715a3768dac6a8d58785225602f480a1ac00dc6632eb9
zd7cc447cb113ef79ee9a8b0451976b39420cd98528f06a1bf28b18ce2f86e9d8d7c3aebd2b47c0
z19027b69fb8aa75fbeffa4bab770e1402eadbe474b508b7f27b727e849220e650c043326dcbc6c
z9a1a76802569c0cc4ee2fe828c5a81862eb4592aaef2eba672487a59f42dcf6e1c9a1c4fb0ea3c
z7aa436aa8c9efb2a13a226463ed632c006974f85421a8415d6d2832bd39e5799b98dfdf2e36d2c
z882c5ddeaccd04c45a395447cc76d317ce0c972a244ec84bb2fcced67593124edf998bf78c8537
z21732f9770d6ff8db16e739eea9d1faf360cc9df72182ea4e8996da0500d8d2d790b911265bd3e
z4790d09fa2796bfac3e51928b49db78f6351dffd06c668d4cd7ba1466c188f23fc0889a75c3683
zabe22c7a8cf4c4ea1f0cf47977248cfe4d690cd2e5505b17b19b2bc18c279fb036b8713655c80c
z9281e7f9f053e2356c20aaa0eff2231d7a60248710ffdccc49e079df4836e430420d2fe91c6386
z190bfd2f5d64ab3797601ce5198e18b8281b23fb8a64dad782ffc4789b2a4781be4e2cc5e24b3b
zddccc566d00d603d73385ca5fbd466d7bf8b7bb6716c7f2fb129746c2641628fdd93f84aa338e4
z1d99e95a5713bcf24926cf109659888e9c8edfa2b8736aea86e2a9430a1c2603ff0e7f145707b0
zf8a3d93403a137a065e542a809fa929d262bd9eaafdd9b323f5255f3b4beaccbf556f18de249ea
zed259ac86e2d4d7157855621a93e1aa3272a8c57852f5ba26ad7b53f2e7e3637fcc9f9cb1cf97f
z70ac56c0ea3b08df136bddf44be803c89d4c5b2eeb28b9fb218fc4da30e18a8e69b6e49788af37
z895ba797a6eb7bff82328f0412874cd5076f69429e69cf8939277ee59a53b505763c59a110f172
zb109c26a8f2644ba9081e092acaf42d7f79e7c4a747be76625b7a61f445e7954c87391eee8f19b
zd8ebcd32ce11af66913a266b76fa72a3da484982df089afce4337684691a7aee84d813c0e9046f
zd3fff5e14a8a4e4f68dc7ef0f4ad6cd714a6c19edcd571a1fc44755b2f210a512787bab3c47841
zccb2cbc6636b6f50390dc14b6f8b628b3e61e44bd09588c2932262224ab920814905e4fafbab10
z361c784e28d659e4535072ec4bbf6cfc6c40a935545b3a9a0b439404192d890403187b7aa00252
z623d05e8643d3412732f10409a3561b02ae7d7ab652daccab7edf1118f2b079b3794ab99bb728a
z3333d4a086ae654abba701974bc37fe716593dacbcfb2b33da13249c0b29ae9076773b7bba13f0
z36962a430c7ded8899269d1e1f931f4417651bdcc59880bcff2ae77eee5e43c25eea48dc9a06d1
z8c645fa47229ba6fb5e795f17d6168035d7b70c65355c22a9463c09b10d7a9b4aff524dbf706b4
zb6150e5f1c53625afe1f8e9a1ece27bffe4e2da768b434a806357a34ff3af4056dc50d633add28
z63e724f7ae99655f45d5899d99f29192143e282ef3536cd82ed1394ca4f2dcd7cad4c318d54b48
z8097f254a15b87ea0dcc338b62f657927d884dd4bb9011f6ea44f39e5fd04d64151f79ff10b514
zf5b9579c258a745349c66089fdf01189ca0d4e0067adb7f0c1bbb09d2e8d1d59c0617773c93776
z8a0e2014d32ab9a312355d1c620648ae655636a069dcd8ae32c9e9c461a54220211d051167968a
za3476e9acb1afd2dd1db9807f39e89b5360692f609498c0d5fd3e79206a31cddb667a16485c86c
z5ca5eeb13b96748f9ff803f71b30d0d4ae8fd9429daf01c90518d6da4def801fb934976fb9ceca
z6d5da383768514a3e68aaa5e55aaaf5b7aa8c0bf533362f5f86ad6518d3980cc6c548c796c46e9
zff4594c8127e29fd3c435c4af1fb64cfa1c4d6ef908b08d3b6b526e28aa1d3ad4924c8b698ee3c
zd56b60495b0ecb47870ad60cb697ffcb5e84188498e53fd2ef89f57dd744fa26f34e8c291b4422
z017a5854749faa5398021722db6d8a677b78274f232b6d660a4148227fb43c56f762d06473b6f3
z7444b577a9e8a4ee67ea5d63ccb1a73eb6574b26e220f43e14ec7acffc4368cdacf36466da8f27
z4e551ba3974f858fccf05d62e4a1d2670e0962dee8226683b517637caa15538457cfd830dce643
z40eeb6c8cbb9256b6d7d4e22c6c4c96ddc2d35f5baf3b8d30a9ec6c07d21c08a2195b554083de0
z4c02dd2dc920bb9e79e23887ba769987c3a7c56a165709a6c8180faffeb594b30ec411cbd0ecd7
z9c5592e4a6c3512d225b9be7023d3c6248669afbf05e6267e0c7a12ba3708aef3e0e7a95a9dcf4
z56a1bd8c2fabd578bb7c402c1d68284b652266130d8e2620d07c132ee4d8bec8ff367545edb89b
z6b370a7642fb18e749eba4a8ed014e3d28ed3877d283c0481eaba5a6e12e20e5f877941ea9e2aa
z8eac2295677bcf50a2d976997e747cfac441df94d20e3e42eae557f1386cd551dc7d87e1f44549
z01764475c37915a80af6b2d4dad7561328333177d045fc205be0dba3f327581ce33366bfa79ed6
z74910b3b557e062e10e8202c11f2e4c927894eae212cb7530bf1c023120c38ef38a6cbdcc09be2
zefebeb91aaef3e5f15fcf0a08d742a5494a6976d102506eb55d963243d0f26abf78d62e8d62032
zdc0935f4636205a63b0d13dda8b7d182f4d842f04195ad3804218769c1d4a60e8b3f12caa13ae2
z888635b73808b9a18d7974aa16e5a90a7c33f047f3a4767a0ab0321bf5d0f873310ab960de66eb
z622542bbe42eb90cf8028d9314a1060053a1f6da6edf532921029a1bf8702495260f030e6d683d
z91829fb4cba3cca87eca2dded3d8ab16bf0a67ca12125ef2abfb4155c2c9eb73dd1d8ff0436194
zf7054e9f31a42682af767bb9408a066a13cbe4c3cf2da4053772ea8c39c9072bdb44fbaaa3ad57
z8897a93db1e9674b74f6e2d5e32f8f76aaaccea63a88abb8205a8ca8b9b2cc3e20ac8d9f0b0781
z6ccd8c514fd899b2798b885d0d9334ad9215b31aaa870f15b20d5b62bdf48b69b1bf9b74be06eb
z7ce5643292cda0a4dc83abae20ce6130dac9cbd0ee210ab6f2a647d869f7431f6aa27ef0edacfc
za5eede24abba55751ceca6d1d59a1d4e49196322939c367544617d14621c503651c3adc31d9ae5
z5682beddfd6a53c4175ab2573a2820a8f69ef33b0c28bcecdc72c6af73324cebddf928a622ad50
z6823270e308bad1279853fc33f6160e540b5045cbafa7b80ca816689c443f5bc5405ffd5b97d56
z48340dffd24be4e3420b262f71897f588a59c5fe8717a479e694c8554e183f00c3f2be2f626598
z26995dcf5a93f1af6761411dbfb39128ef9511f7d94e60e11ec6134c3a3ce2d5a1dedb2e464d89
zc33d51120231bd215dc23297be9111a7659e73f89d733ec838ca3ae8247cab160311fd4a201785
zcbe02657a1227fb2955d07d0eee1399aa15c69f9aa35b6784cddc12c87fcb5583ed69e1e181c87
z0e839d7d40fa0cf269d321baa849a28556d935c0c6511556be44df18b60a0ee599530a55a0b045
ze168c8bb32c14e42adce3d359be1da868686da79445f3b43336fd407cb0478d995a0e1f1f9ce18
zd7e5fcd87d2bae08c48dfad771a0acda5957e47fc04eb03e28f93cdb801c91d77f4202bc04410c
z606fab2d86d408261ed25ef3a5872ea8e17ff1254581ec995a287ea503f93f0cc6a1c691a55c78
zc912bb8c9a59938aa6385ad0ef2720cd4097dee5919a0ca2bd40fbb481b9a1ee22320af6155405
zc1d57b9226fe3ccf35d23ee752de6df08f22d855c00aa7c81d8d321c3e78c1cb358f0494b2d59a
zc5067dbdc140b6508a7085f7f1fd8f13d855ced323c615f8fa709bed829e4334372835bdaa2b8c
zdc8ddd2bb55147fcb3b4296f9699e4332584445a5a19f1d97ca1f55e5ae6bbc961ac46236b66cd
zc30558273f0074e37e59d7d948f69ccdb0da7cc17f36f6fb79644964eb12b7f6cfbcc1d249faa2
zb1750101d619e6e7c58b6f2f76f153cedc67883a75b528213f3e48c4f3ff17c80930d213ade2b7
zfe6d63d15b49c4d61ff79a9ce1c1309eef8a06b6812277e997656dcd8cf1bca578dceac09e675a
z1123d73d1ce92fa8785197d8f75863b25dcc22261328759ef1357fe8e91e290afd4098accd1f26
z65ae54f8a0f6ecb54d53f191267842892fa7b4c7a65b0f2afc722c4f92efe1f361e9b9bb5cce8c
zc54b385c39e81f423fc6f1b4ce96add26d8a55e86e85db6e28d6823bb2a686fa2dc39b38bc5f50
z164fd41378172e1766b412b5b0d457d2fa2eab6293ce4f7fa4412718a5109f1e0fbcd600959b8d
z72c62bdc8cfdb4275923de6cb3214d7a82a62a001e156cfe54d7f6636c1a0423ce6b582738c374
za30d4a8e5c35f5ef9b353580d2b8fb9ed8fe8871c995e6a482822148815197650dfc3ac1a2a8f4
zb1d86171ef45dc4647e7857c1b8f9ba79728fa5d418c9ef7ed26dd56529ce0705f066af52ce262
ze2de323ec84a028d9ce2a07a8061a08184e17edcd4ef673e73d56d26a3ef7c48df0734ed25198d
ze633650a3251cc29b7043bc73c2c61e9c307d3afef0c937a384873f3b10db63f63c21ba29152d0
z46c4c91ac6d805a224c32d9bac9fbc812b051ff60d861a987be167540f62d5f870e20ef5bc034a
z22309c9d4c8a5ecc443ef10cb5a8d051cfbc1128189d101e7a40b3e36816746085af37e835c1fc
z7b8f56458d309dd14d3a35e32f03d575cfe04ae92054d14c516eb364bcbc49536b2479793d8db5
z0cda7a7a1d6b381e2589437e972497aea46680f2ca13422ab8d7cb1df30722673ec59a65e9a997
z14aa0119688dea8a94bc2319018d77ffb41a8d6dc33a0af5ff8c8aa418b08f758592ac77d9b3ee
zeea6c974843c28af7df154af2196dbd73861c74f803794d2348fdc6fa040dec20a4b2b9d05c382
z0bc56aad33e57e23c3a25fe118cf416991ffe60cec0c39ad12ea9cbfadb43a3e2dae887a3f2108
z8c5a9a30f559776acca6b415dff9e7e3becc193419e0cc0ad1922601e52ccdd8e513913d764aa0
z7cfa091964f6796feb27d25f742d4da20dc3caa014e46440b310cbc05175106a6390cf48fdba3f
z2cd515b5e21eccbba198ddb794e6a97b714acf891ab4e0fa825af57f071a25f03f830a0868022c
z987c378ae2f96ca90d5b45f44f537687c187d1084b88bc9d9ef8d00a58ae68e87a4f33a913f4cf
z17c292d8ee48421496b3a721eb72811586c100270e907616dd00441be603ed20900bbe65648736
zf06182b9a0fa6d0d37ce13c2bb67a3f6e70fa6fe708c17ae9d81db91280593b91cec9538643382
z445850828edacfe15a98df7b70ab1ba51e31bc000ce5499856bb3156bd295f23e2247f4adf5cd9
z08413ca5ab6202a4c06ea7018ba4961e1049dcea603fbdddd79acf5866ee5619491f3c4df0f761
z18c70f4f35228b393fa59765d11695e78474829b561deb915dda186507c45bbc03b0097a4494e4
za3b0992f7330998e8b323c8cb240390b41711c8342e2e33b6d596dc97b94246c06ae30ef0d0fde
z7dc4abf20c4af823914e9f8cd2aee63ee22a338152df792aa8b7f85f2bf3ccd4b4bb96766d9004
zab933026eaf04922055c1fd756946c25b416ab4ed49535afecbe239387b577139452f721f5d71e
za028ed26a3fe67fa9e2b7d8bbe5fb4cb40f744732c08769bfb6652f1fa55a0f0b7e31416263bc3
z01e301634e8679be737e01bf1b4d8cf3411b01d0e1cb76cbd7d2090aae73810adbbbdb6cfaba46
z9ebeee18009f7adf147110507792c7c91d863e8d2392e269cf34429a3d424b030014230b9c0d08
z1f7afe3c4121d7897c24a20be97d196c820265684136cf9cdb4a9e2ddf27823018a11ea895140f
za1ab24b033822ceb1ea0379519b6b1aa5d9a1d6f5a89e304b7184e8372fff19e72ee8817d9211d
zca2745b6a5a4a415d000b4f1557c956d4e025097f2b227c421e05a1abf680c2c10d53c6a6088a4
z20ca84334cd5d8c35bb91afbcca014c0aa0be3e9dc41550976b99841f38b3636ca879bb8762889
zd1cb70776ebcbec6c702b5ccc044759a1e457da71be5be767f6ff908bcac7d7f6cb9ba909041f8
zaf5d1c33ff951539ddc6389c931db734cb7040e6b0207a014af7c40434c69d1d33d87d7c46c158
zedd25ef83c6da8ecf647afb23136117a994de2411213eac40b168f70dd13b0dd57fd76c18f8faf
z2c1c440c59aae988b52fd5e7f2f4bed28e36a2de9c8c3a5dab13856314004dcf549e3524fbc139
zaed2f8f67b894c374f77cc576cae0162895dc9ad6e2c7340bdac9ef1211915e0fe22864f30e715
zee221c6732391d7bcc16122e9987ae8842181620d3378d068fdab134f6fc277d69e5c6f3e7cc3e
zac1bd62d0e4988bc8167b5a974162974ccb78dc4895cc9a7230607cd1a949a18d8e3ee9ff39c46
z4ee0913b19abe8872c6204455816bc5d79c9f1c0bc16db8e234908e49629130c003109eda34011
z7e679b515263994eea7f91b35a9dc5efec86028b524651c556ffe7f98773339949e71b1bf318f5
z83fd5cbe20a2c6c41e1698219856b7624eb669166caa6c0dee8d30198ba51525316ef259112e39
z95da23b2d2aefef4ed3f76b55989848feb5e971afa73d8209e856d12655d591af90c1854c83411
z897cbcbde21dafd57d4673b91028ff6a51f9d4f88d9d2dadb85417a5ddab06743558633d21ce72
z222727911deca16722745f4512970936dc580965ef487eb8c8410b87c64a99afb799c8d58003d4
zcd824bbfe82372b2e21b82c119e8e1451389c762230aaf251bdfbe59bc245adc49a2e039cfe50d
zdc0350fc61ca3a529734227f02576a555dc50cbb3909b4db641846c0bc625809eee2d238dfc29c
z78bd6d349d3aa73519fe97289ca244813a8c54f3795ffdb99798261e2dd0da55a9c4baf9299ce4
z1027ecc743b6d9bc61d8b992fd38f86667ae8951549e93262955bf7d13d5579582d5907f06667f
z096a040a24917c9c63ba6399beb0405c496fd9b88ffb8e7f19881381846e1b3371f0f447b68fd5
z61495504406d0691c767581839abcb48557b27ba2f624d2bebde433f0c78848e96733e456e1247
z8fa615df6d5b7a601cbf63652da910522a567afd44fc5e7a3724e8e44475764365d680f31a78c6
z5de8994f2b75c94ed961745b3c74f34ae85a24b7a2ed1e38affd2a8a4900a7618a20793777f52b
z50845955c8653fe6bc031b8f8df2dd22e63a9d642e56505d6d6630fb706a35e6682bfc92b3e56a
zee46bb50a16cbe8c5c0754f91203f069f4cc93d4cc40389b200c03dc3cfb7a7edc69096ac762f6
z56041a998d1fac326dbc5010952ba0bb1f7678e56549f66819508c9ac19e7c183b051fd50eef49
z250b4e161889170a81ccd079ae414f2a013d1e0a9ea8edbfc67cf3fd922aef6bfaaafcb9689e5e
z1af3e9dc06072dd1825c130eea7c3ff3e5944963b4d664ed0130b16a6fb303feb1e13089d67064
zd208d507f3b199812516600dfbf780ea7eb19ddc4c62ecd087f2cdee4b9e1fe8173259de501f39
z7a4879870e052aea4adccd4d1723297fb43b6fc42cc7dcde7173c4137cacfd4d999f21bd133bde
z6110c799f72ac3884959920e8c4ca7dbf476c6f6121a192313ee385a4bbb78a136f05309b95ce4
zf4f7c4bf39448ba1029bf529cee9fb9e0177293545eff105be6b8c54a02ed0ff05f4021073a9bb
z1b77b64752a534d955ae8d3a80c1343422b0e1e482e18f4b28bd876be15911077a69e7ee8dfe98
z38657999a38aef12be8a8d24da236809d21e0734790ea8fd43460d3a525a4c07b3a944e9fdf088
z264d604e544f8558b87d6dfabbc02669cc159d238acc6a798bb916d29adcfe4f9c7b503dd2bf72
z23a13334245e90238b4ef6ef76b6d24b3bdd80f964f859de66f8650aa1c1601dcdfa590fce24d6
zce4aac18087fd8b5cd02a63429670c59bc49a845c391db31832d1ea4df2634aee3d74e9a90901c
z3775bef098b61cff2c030f04552601a7e31c7e8eab546b0cbcf6037103164de79ac6fda5a51e22
ze64a0c748315fbbc166f531b9deae0c3ec37b038f5de0fcd2e09318f3f7eced83eb8d8fd206f95
zefe265ed71e5df2a5004cf2954de1233ef89734a046e10e638cf906b420eeb2fcea28510ec138c
za23095cfe8829e6f341f830cef65507d5d4dad61a74a1d75e6e31097b0b3f4f2c852b206c66c87
zac2f894f6875026496942bd4fda99c1cf87670c39913c346279326fcc52b695450a7fb9c5b659d
z4b2cde736cb14054c0d27327ddf22303e75215b5dfacc2876b8405d31c7a44055128fc90f46df4
z86f0baddff84898fbc47b7d7e398b38c4e4001ff5e909a2cb232229f6339c2ed3c08348883f7bd
zd1890bcd705d59907de7721d1983eb4012408cbc4557a3877c7cbc4841cd771c39a3a7c794552b
zac31f1be731c91b3106b3cd3da8e2c21d046b137d09789c9a5c8663466a879caba0b6b48e93b84
zb5b5e3c4cf31b388d0950e062d799de3da390e46df738d7e9879829deb86df940f1db33897d908
z8bcd53c7c589da128024c05e8467c34c2c837a434c2e550211fbfa59178c875ef2c4e197f51168
zea319d8b31d87cc6b95f6c8fc572101553903a7de45a52d87c29b4d353ee52bc991af218d10594
z3ad0a249174f8ba74f479dce15a48eff92cb649559e4340f5fa549c81ac3abdc13bf0884afe376
z30eb1098ac3af707f6044f4b7952646769a2e37d00ed1dc9bed575a21e3b8d8fdad3ef50bca406
z96c2cb931e93f15106f38ea4182025a240b14aed35f28fec7fc806d2e0060258b03e4e174268b4
z07970a1779a619bf6c436b3ec89274fcf4a6403d03ec20f0082949dd3c43df898d69b1e83c896d
zccf1c09f04d3d5cfccdfb9b8e4df40b130fe80c02ffb799abb1b5aee2b873d4077be19131b3ff7
z27a13c7404969d9fbfbdbbd44e79f28f62086aef68cc035915c89964df8ab2f02bbead0eccf406
z42e152917cb8cdc9f6bc1464e6572ba1b137f1393cd345f10f55619f8beab2a48caff0536c3d42
z5c754108ac8b59798b765c5419ecda5154254fceb9ad517aa70bb9830eab7e55e5ea453dd6aacd
z0356d7dbdcb5a356d831527a5aec3c990f3fa5d5d3cdfee3cc1f2b10a60a8671aa1696c241e38f
zcc4007786183eca0cd062381e5bdee9bd4a45b1cb51f260b076850ab413905b8e7bff4704cecc0
z641e599f7050779110dee71abebb13e2b3786c24d55870d203a648dfc49320639a24bf6fc84e14
z322ddf6d74f9d78370bc7299977abe02be11d7dd9c6fb486ecb73a1da06fcfd71ff2fa05a46ae6
z9bf615290028cea65b68dcb77fe7ad2f7bb1742f6d9afea1a256048914bfa3848937732a97635e
zccf0d3d92f482e0dff00317b7f7e912f0945d5a34178a863139c19908a228a1a1d7559f8fccdca
z825bbf1e1314530c1a20530c6c91cafb7d554ba70800fd9096e73dda577be935168b0822b8c9d9
zc62c6a66a59a2a237e2598be5a5c758b3488ff6376fec32b513a93f0a608baba28ae812f095a1f
zdc0d1f69c3d61f94a891ae1b88f946e6974057b83f9c27a7cd08074f9d1bde98afed73c00e79e1
zaa78ad7b7a2441b5c4b575c1a8872320b9fda6db948bd626c27f0ee0895f107aaa3d5735f5b7b4
z4c882a420e8bb1c4cdde23939958cee403537b4ace2eb4a9a2c2c84ac1c26137d89a1dc34fe194
z41e15253af0116496430a6252a5776bc52d1daed875bfabd407c6fe8a5f8ee046c5c307a5603eb
zcfaa832c38343bc634d834c6cbba4d081b2ed428c5ca8abcedd8883e3782e834789b6645a1c541
z024e19190c0833ac6cefba7a2925c64536962772c8673609d9d4d93fbd4c44296e3ea7426f567c
z1030557c2b04caee1f6e270dbffb6a640a4030d836a96c4d7961104f5869a17941e1873d5ca5a7
ze6928d7b14fb091d986fa192676b8452aac65e5d2720ef7cdc53029fd5c42bc9626b0ba9b54eff
z5a964c1e9584e698a5e4b04addbf1fec98cb5b641ff48128cddb7fb37506230a5476c53355af4d
z0bbf7d35acf8b4186a2d9982b8984812f75c4212edb2725fb6debeb0be2d48f5e53acf07e2e218
z98303faa1021fca8cf2fcfcff0e781fb61251fd772186200bbdb818365a4d36745a83821a266d0
zbb2b6be1197903876f20c4b1fa308dc5f340c0d92845b525afac945ae64d340a290aa0d8f3142a
z7a98c3839cb13e66dc37a86e14af01827b7f5e1c09bfe57a5d65217dbc113d74f60f9e461ad9cf
z20490311445b68e272ef71a7380ec60fe1580bac99a331cc3ba7a754d31ccf8d03f03f08b758ec
za2f0b9c691f542404f0750318ce6d32e9745a89eb1956bdfdd2e3cbc8be97a7418d738a648e1e3
za7e3e0ba52575866c0ce8c9184366c1f633928d6d3ce321c16de60116b8d1358e9864697557155
z273544844146de58f4c362516344ca6e5e9c2553982415a1906c4bac57afbb600bfa8499cd2bf4
z312b0aacdc05ebc187b24eaeab1a18ee3cd3d79eac949a0aeb29edd60a9b05156b7c762f3236ba
zdd65e133b13623ffa1c802b2e5fbf1399ceb973fa39856a0049c8cc4da1c73682b68523838d95f
zb5f0a2b65aa99aa03a7616cdb6b72afe40b62beef3811c0ae1d9536034d66210dca71dbd3d0d9a
zbca9cbb9dbe83650949407e2f11f28c8aba435addd6ea786395f6f3609673c46da9b3849040d4b
zf65a9b935f903bd7864de10031184ae39c340f9615394a90769e94590e7f68b65ef1d4019623c9
zf59520bf7815feb8e06bc0bd7b7e2a28f431fc7e46c9a2f202d4f81c632d9d0353807c102ea9dc
z48a539dbf65b12170d16c01e9d37d7ef686b09837ab1387c2eef8cc88e1374e6697eba2a2c4273
z1755e5660ee1cb4b7446029c72e2f94193ac66cc90b9e2139e355f2d1546abf3c6605d660141e7
zc2c5db0bcfa9ab2e994ca61547c8daa999d2d7ade8c874e2eda6d6428dde26635b31c0438a5aed
ze0d636c0289977c020306de712ea72fc37e7da4fdf63138d294a7c236086ad8427499ba6e0fd18
zd705b16b2888e72d4ff0d4e6bb72687c1aeadf98cf30b066742a11e0d7f4395cae0df6130401d1
zfeaf5fdfbe74f56f353c29bd3d3b56884d3e69539469dbdb88c76451dc457d8359cd8bedd97590
z3948bb0d2133a55f6733187d5f3b91194fcbefa56a242b9cd4f44d1f5da453f3ddd5f8675646e8
z2e287c49293ed51fb1f58b43944342abe44020c38e624c181352b5e9695e97a5356fa082b46ee9
z29b65797e979f5f9c111583e9970397c39ad652bf08fc91185ed1a29c4a7bda4e63a6d8dda5eec
z7136279cd42ff769fd09aa28d645cf9189af0d8c614015451b4308167c4940761bb53b5c56cd7a
zfbdcebf22ea17ef31d76efbbd5806dda7f4f2f04b36664ac2378bfe7cfd3f9a19433a6a8a08cc5
z8e3b2c03315908014acb53f357c68358f0c590a2710f4eed40decc2622b646c1d3eb8839960441
z3cc35a84996badd3e160f6dd88d891fdfd3f161cec79ca1fe22bc229cbf65e2473937cca3ce692
z9883877e902901f44c28a70213ebe9e6546c805e33c839d6391264a7a5e808880b948d1fe6e59f
zbb5b10a74f2f58a2c2768eb8c105b6d52593dad2c4ee579fe215d9d5042f11ea022d03d48be527
zc051b656dedb2dcb16020dba3d2080e74b36d91a77273aa8716745f617efba5579b9d9d545d502
zf495f1eaa33b6017a1c5935b14bfd313d09225e203893a3dcc19ae3008029afe6a8f9d9a2faaed
z9a454b57d47cd4c096ce649a10b8cb098b6acdb0bf77bb1780d7ce7c9d961c5c061e835c59b99b
z04d1e930c9a017606c35b0692cf51e833c309326601cd47f8a586704a6fbca0586556177d90246
ze6f2c21956596f7919137739b80dd699a3bac2edc15a10b770cef51700eb4427b2a2e1f22376ad
ze5511e17af99bf9b46219f6eb1e0ba22c14f9bbb9dde6d65c0b831c544959c1b2a16d525b27da5
z5681429a0f9e66c54fc41d333e9e6fda2d25eb0842c641778fac1c853612272b63167e3cdb826c
z541e31cdac3884885b5c854431f3a0e770a141d0e787999cd8b53bc86c3653aa057e2d859e720c
z7285e706656c362a463b777ee5280a3f87ea8afdd2312f42c0de4b633d2f5bd0ea6fcf6c051fb6
z5b2e846f7a983fba01df28774bd9a96447aff935749c87f4e784d05ee7fa899dfb67f9eaeeb947
zf8a2d3e9e108e287d837ff5efb05afbc8170a27eac6ce64c84f1e4853717995cf082a77b6bcb9b
za3f693c0e7095309bebf169f583b4041834de3f78a9bf394838ab49961e11f36f2b303853302a6
zf497a012bcea0224ab2f59a79d1ee5d73ae0dd134944ab7f4e02083f59d7f95310507d080423f1
zb0d969e21641e92daba781a11ebe41af6acd7639769a3af1efa236344ba46594bf8c2ceae4046d
z98a13e9890f4cdcf0c11314c15081ffc422ff2f065407891744ce631b8e9941c9fe663520187f5
z1d94d91ece0f4447f7ecad0a7147a2786caf334da79d6e893200defabebbbefb6cf766f197b8a4
za71264dedab6fee0098c91d78b1c5f45b4f3d412192b17e12737af765a5342a2167ffe52fda685
zcf8aa3c4160a63dffd7eda0ac3c8275ddb42eee18115b424cfb44c7b200b284911dd394199abee
z99278f1579166e2bda8e9a724b8e08820079b9d814d98af79fe57708d32e2c70c2dca2d6c6fc5e
zf72d9e854e7635ab8386b4fdf7eb865487235e6a258080646e639db562f69205b351af2b180f79
zfc390410b4a50ef2eb64e420ffb014db0b20663c54a236acce66b7ce946f3daf24772ea50605f2
zbb06ef3f3463ff36f2fc2124a6d3c7115ec87c56931c3823b84d997eb2ec25403d760dcf800faa
z2d146a2ea994f53f246ccef13b6a1ed566a780b0171129b7cd43e7908244abf79f2202d007ef9b
z92aaea4f8678c911183fe35abfc51e0f646b6c0f70ec4299d491e7d16bdbdbed53e07692555447
zadbb0e14d79af2ca3db080002f31cf14e72ad629a5df2f2d45f62aa2d8c6b8548363a8f2d8da42
z8adf1d4cf8e800e0fe5ebf399087aff083f1dbb1053f32e4f29ace2881b90ac916733a2230740f
z93079f3f76deeaf2defe256027985f5c8d0a2b9d344c9c222c56534612c61756d5424fff9f857c
z0f963179103a47331aa3d900b59f57dc56078b8ad9fa847ef2ce190746a1e8f965ea6a66eadf5d
z0dc2e607b536cd5ebf3b8df8efb6cdebd584f563d064d2247a59e63452ef71d5adfe6ffbfdcf8c
zbdb7f750454217b5dbd3620e343e253d3f50ae7e57ccb877cbeb8dbb9bdddfad614372c42cb90a
zd70c01bf9f51786aa5f20e45f8741613c8d3082e60b585bc4e06c07686b5b29a30877f7070f5e9
z25df21d8c457649c0b4553faa9e6cd272db33ab229a90976ded263f12498c5fcee4e1158615d7c
z44e006f30dcd0d498d9e02023155b5e900b44212f744ff5c913f595687472224a1c492e911836d
zc0fb06693a474ee527511ad3331b52bf41feb0e3e45bdbe5c53ad74e3e84c9f25431d8c0cf991c
zad3fe4b6a819cc799ab389d16d8538ebed67e33e28d6851a859773473945ca6742ed57279b54f4
za7f5520ecd753472caa518e54a628f6542bd730d3267542d1511a8bd861774f79e9a778dba90e0
z4a2a210913023f95e7bd2f374774ada6c066ff2e8a553d31f0a3da6ec8cfa602bbcb93dfac37bd
z56578ce08d5dbf3daddb4451e290f99b70eb76699fb0b4628c3c55423e7afa41f93b61e2d97bb9
z403abd2f08bdd333594aa97d7a19f588e1f76bc0353c30f48ffe562e8d6890c324e8bc421382db
z00366f17d532ed3d0912676784e27f939e0bf95b8ef8b49fe0c49b439d72460c4745326b8502aa
za926ee884dc359700979ebbeabcfaa0dd143ab815b4d559a09808f795d1e4ed30d082d1aed8e61
z19b0e0c3482c669e68baad5f2cd42072eae4d5fbce65f42fb1c15d2aaa5f169c2ec2d4d9826bb1
ze76c51afb0af98ae92a6244afb7170b173887f1d03f45a18743cf0f2fda7abfdf54e745ad1516b
z8f87ebcbdb97fee3797d294b05e4c911db13ac1f1c75f5f51db4a75632557136357c04638d9e2c
z044641f2e350ce833f85cfb513705610c5ced7f8f2fe4a54bd58db49b791fb9cebb6c6084a67ec
z526fd92fcd9e973f315455da34e3de93787120c209b4c08ae0b6d4374c258e4ee1d20899c894f1
z41f7eea9baa2d388bf99f1cd73ef86f1b9ea3ccbb746beb9244480c7a97532276da1af2c5e8e51
zeabe10af1ec9680d5146c50c90a2efb7ce809c40e7a7509d8c325b79235e7dd8c747d849d65cc7
z6b66137acf761a29fbcd86d0ab297298880a8ab366615582ff22a566f077a5fdf93fa2f713a097
z851f467adef0932127b667f71ea14a9070e0020ca11a9b9f87733460d2b04816b8188bb567c266
z5b3b456afa8d26ac894c1ba5b7667049506fc087fe236165169c9dbb3da9d5e9898afa960c98c2
z08b186ab67243a12d75154bcff7c4d5b489a04f3a2fe675db194a0f73435c73e341c08edc95706
zba0d1b1383a3c17fc18ea04572b0c349bf76a43efebf0ff251aac239a6b9637d622cac38e2bfe8
z3195ac93dddb12d0f302044ad1969ceff07e4d328a6905f94b89756ec78c33e420565aa575b779
zd02191da32177f53988cfbcfade94c27ba5f8d61e4e39869a8b65226584e731559178d430a4410
zb9148ca5e9b6ef53e9409a95ef29fdf4039ad3b39f62a76d55239d3e277102673c100e659197a5
z02cb691542e36eb23f4ac0f3937470d2ff44420dc12d04cf85dedd9346b4619b55dea34b73076d
zceebbf374805c761e8f0af7d89acadc8b82f27b5c94da671d469b2dde9c9bd51c0bafedbd26841
zb785355fba7e6655483248d823e1d980253bd5ca3f1ee9000f08d241f55f47544ac606ee5133d3
zc5e3ec1b29d73e836303bdbdba8ff967826224c85a253a7c4accfd64c618177558e0787564fdb9
zcfaae0b657e3488daec8c6dfaf187065c3e4927ba3a766c8ce2a18a2f7cf7c5e982ec8d7c05504
z8b926efa4598494599d57e2f2844e2f10acd455811fa1d0f1ad3a03c4febf2e02ad56c5767fae4
z1fdd78a2aea67ea0a9c238bdcaf1b12530fc1e3e981c3177a55a70bdd75b4fd54c03e429fe34cb
z2dbc4e05c77ba3376823a2a93432f4d783111dfd429e548e147a8092dc4e9d554431a4c1134488
z820f6b1a0ff0b25333721b0b4e5480735b70f1559d084083fa4f5323a2afbaf632130bad634b3f
z4d1e7dde0dc7cf47daccdf0111227ab15ea483248491e97f615cadaf51bd60359eb2a3ffb3bb0f
z17722062bf6d08be6250c3dde0e2bfbf4eae724fa64b57d3b2310a2278e0f08e54dfd03e2c00a6
z54b0f28299bcf091d14dd424acda544f3a66b82a2eb0ad07e26e55c2a0332c3e49f3309a7497cf
ze5567550bbb6c809054b4f5c71017a9657d1986bc4a9230c4225189874f6ac0c41c77cc1bbf365
zfbca3384232ba1bbec73d018326462936eee8a31d02b1efea8f7bd03677258bace0247421e9da5
z14e21d46e68583aea4d506c660ba1d321932f9085d92a03b1b2159523e76bcbe1c6fcb129b8e5f
z8a56deb4caf6fe01349d74fe0c5a811899739fa2f3d9fb40e758cf1be8bc9143c8335052c8798b
zdd0cde0e7830e4720a3ba1ffc8f53205e4b320c771e2b20dc64df00f2f207aa87d46dd4b115878
z81fce45ac0d6211eea08b014a757846633af3f215a68d25731ea8ced0738d89c2276f56e7d1958
z0d59d3c7b4da2f234d283dccd0df0aff408d66cc8bb597a5e74d9ca9cca4b74831760c5e23e300
z04233cc491f90a893e33015356a773b764c41d152e2cc4773ab50ed774ccd2ebcd0c844b990be0
z9d54755357616bf8e742a090fe6643db551f9b84bec3855ade9ca848ffc73ddaef2e958d6ebff4
z4e8d623afdc4a4826d6d0137b610212df5bd9f0fb20c28d3e29356a5bd45fbd0aa349ce5a8f9bd
z9b3a50c971135c33d34588935c1df58a22445559fc412723be4d3d686d300e5fa7747ca1a0e2dc
ze4f56395af4d188ac058dcb6166017134960e66ff37cee7cdb85cdd2f6ef9770082e1c037a8532
zecadc8f8e9a5d3e62e25705baa731a7674f51774d95c89fb3f53ed12b41d07337ea9c902d01449
zf7f79637089cf86421eed1d7096d9d28d9ae72081caa30b6c22cd108a7b1838bc6ed9beb7e3e41
z8781b624fcbcb572134cb0a2a7dd71c961f154b1b9aecfbf62ef9b003dbc72cf0eafc3b20c3cf7
z3a4144149fa984f6236c919af620c37e269464840876b238050f58e9824f4302d73a1de0fa45a0
z0e33ce0797e37be7f9b8e3a5059f58a209d778cc2eaf858d774d0d66fd27452cd47318f1801c3b
zdf0ed5a5d60c423cb8248b42d1683c3fbb4eeb0558a53f67e8856d813728ab241f7319e8aabdfa
z5fd8fde8d31e3305e90bef8b025e1068c0f0017e34c2728d2df2aca537c6160ff4f919e84854fb
zda370484e4ed0035e7bfa4bb76c54a6900236a5995beafa8ed801612ea674db4f008f01cbeb5d2
z9a29929523ea98704cd55e88b1ad845a799273df0ee1a231511a0d11edcf18727d5d0a2a9c701c
z4414dd05f220867c3e6d4c18d611d38647aa117a4d69b300869a5eb31709ac77b57f36dfb3d6c6
zf4023552057262f156d8b628a6b200eaca9ac7b02bd1f5f24870dec27b7254a111f7877d448a87
z3ef6d2b009d043392d1951f8b96928d75bddf8f90c39b96cfa95f44519c3807a3444616d7b9121
z447c1b913437a268ee72ef7c26ffab4874e1722b31decf54778899071d3fb1939aa8d7d62efab5
z5048469bc484c823c027f51b7b5e82a6dcf8faab7c3a854f86030fd512b1f5a0782ee0fe8e2deb
zfe5ee7827424dd93490cf7d22254df18bbe1a409e5af0d87a705679ffa57f805e1dfd0bce70e04
zbcad75523353890939cde0b25a38ed05ce159845f8325bf98a42259150db599c09423fbe619ccd
zd6d1d6f85a4406777a939bad70b49d5a1afbea9ef3aeb9f6bd3202d09d990dbdcc67b3ab6ff475
z611580d45468f6b72775da933db5e84f05fb5e4b0e35cc61d5ae178358b2e608db1c891126aac6
z69d02948b64027d015578f613702b1959521fc071485f1f5ef8878a499d8b3ad4b48309b08461b
z501ab43afbc209e54cc4d82d1425b0673b0ce3811211a3b23335aa654e094a6c0c0f36062639d8
z9c03f671f6101d3003ca1016987028fd0c321c5e396776c915dd25fbdfdf7aa82e4cb053cc5e0e
z1cd99e1fadfbe12c2fd956083f1d33254ec27c0e3df865a4bd1238692b16097ef67eef4453fd89
ze67782e7ce689ed44f7066ceafe8188c4c94ab8a00613b85d6dbab23d28ece7f71b14399cdcf86
z4f23d3e77057686f4294f7ceb00c121db8b5ee07b928925f63389771ed5ed5b90e502cbda3e925
z8f6f69c0fd7bc87fb8bb224fd339eea12d7363cb83e7b08dc0d536b7f9c416093a53996e4912f1
z0009ee7c434fe5140c1f1147c187705aad98428d9f17547d5655ec585862fbe677d9583b699977
za86b9abc703931d3d96582c1973143ec958be205bc626d256c3242079115e80f05fee18d27fbc1
zc0835b3fd712577167df8aa1f88706966ea62959fa9a898a0477179a0b57bb272ace0fc4edba2c
z8bbad9c8296bb0800c254d053989f83aa43128c12300d35d75fe602beb3186c985bbe92bdcd92d
z7fbc1ed5f4e42a1586635350b39da59b83e2f9040a06a9d129868c39434a1656eae08056933280
z42782350a537fb43882a352665ddea833344db49dd051546b19720e2870d6fc3a8c4429e3f705a
ze566a83ab9f093db8159f079506dc5bd3b7042cd3cd740a3441c44cccbc8c602cf3809f4e13929
zf0499f55b8697907fb6f12f2697ca14f5504fada4f097b92fa38b27a64d29fcfec005aadbb395f
z6fa7a1d669fbb0babe32beb3dea52f921727d24a803bbb7b2a16e7b727ded28eb2fee34f02b95a
z2c4359fde29de935b62de8aaaca7a781203f1f0b3c1da5b5d572bff7a071b919fb2f9972bb3892
z906c693a6fab8dcf3ee580b25d249e609167711173dfacc7b4286c311a77c28f78e6eb2952cdbc
zaa3ac2179129f4f8839da9d83e0eec76ac34baf6107798e67d9456fca5a68870a21843c22dc3d6
z442be8fd9984771260d29d73478720380b32ed13064724fbb07fd4d3c0206ec53bf5954ccaff63
za8e0f197e4cf6fd6246c7c8127f8b1334ecbd7b67f480743b2252b3309759e8cd88923db3bad33
ze625a358f47270ba1364a7fe3efaa7dda94c44429080aaa4ea727433c024eba450462e35897db6
zc9ebf3425f9da199589823f3ba7548a9f3f557fa0e9d3d0d5008b5af9f8e0a5a77dfc09e072dcd
z95efb13518b878a38f2e502d33efad2c38efca661cf887a5e9d3a9ea34bb157ec4989249e2055f
z0112c373c7700a7193f4ad5c6a2197d7296534beeac4645d836a9b558ae198080528fcc5d5dec8
z7183fc22654dbeb7f6e408c9878cfcdeeb28a35ae9539db905740acf8cde725df9ba3beaf76bd9
z2aecd4cd196ed249c4f3237cf9b271a1e76b723606ab3a4cd7d686278eb64e51b4d64f94272e78
z71034e88bb7de7a6bb702fbb3f8379130ec9e2d5a01ae665cf5176ba963aacebdf9a2fef2c4c99
z2b107fea60cf3c97b8a93797a684cc68f268edb8f1a6ebcd0c4048b9316cb2076175a0d9f68c0f
zec48b37e06842495eb42fd100b5ca4bd24db95e42c2881cba39ea88fc2f7e0c2e9fdae5144459c
za656734f9109d181d0954e3ac9ba7be7dfc2068db871fde58381ad6046a4893421b15a87d79f9c
z74f2b47e8e8467e9c395f6553df903eb88482b311e09f56ee8617fcef285a7e7266daf1e8ca355
zadc4687ddeaf4efe24d2d402f85cc0d27d1c978cd7eed4af88fe310d10888f0c40b3a5143493b6
ze32ceacba92caaa24fcd9cce2c888a4d0fdb40923600dff23f776882ca4b153d0bd61dfda8dbad
ze71f0d04adfb56c6da57be9e1210839c2beb500ca527ef05ad3243ea945ad9aa49b8ecc8b1f1d0
zd7b8513e71f281d3e0128446f8d3181b9f929f450e375849ca5d1e6ba3768b0ee42edf0ebd25ac
z46e7de40ccc322c4c51ffd2864a69ed1d164cf8699bf02adad05b8106b44cd69ad563d5a715862
za5b76ebf1691a01e5cd3fbf6c3768bad63d590bc4c1683b2a7e600fc973451b4e0d4ddb4dce1f3
zda0edc77d79ad0274677e31e1d090cb6ebe4c649b42bb56cd69f8a150178f51762a210d49a2fb8
za4a005e659df8fac26469c343ab911799b65ca77e9e7f5eb2c1b35dd9a64509927ab0b87a5ef07
zfd1c4c2f29f0f826ad5cef710811086d210b15c24a49523811092276277642e2dc2f8f6d613e3c
z1e2423f4684d4338e1e4c018cb01ee3fc2998b439ca563ce716426959edb5fbdc77140816dfb85
zb8ed2674e65f510a3e9f0499c17d1ca0b0f0641fe3e2dd73f763ff39732c470875f6509688ebf5
ze83c88f68f49b2a46147f2cb69bd87db0b3f791ca93fb09998a287d002b86f86071a3ce579c65f
z27b32967e07b849d93c1fb869a06202fb331619dbe397bec68371a408a9cd27ebbb721641b1a8e
z6551a00cc0a3a3941a25691bd83aa0d5c393918753e4cfc34ab1568d79dd249a430ad136ef472f
zae6747cee031f71c2c0f1d5d620222183beb61826e2493b9f98adcb352f6a3830f881b344ea346
z1cc98a928a6bd46ef7261c2bc96750d1fee8804be44b92be8fc80bd6252e01e84442c5b2d6de3a
z977b828b0ef875d837a654c79642f9d9e18986370a7b0151dd6e83337e6b447950546ea720a626
z06cf10927a3fd5cd063173c4eedd97aa1e510b21ad9396880ba7de08e79cfd118667fc5a7b8e50
zb0e040d458d7c7d0b5df0362077ec6aa7e83f73e4bbb96121c6e4491e7dc5e4864a2d34ca66100
z40281701c2d70db1201ce7832c948bb8bc088f4d1af6fa85e3d664b74f74eb43fd0831eeddde13
zde2e463f8e8900ccb309aca7ce756e1c97c9e50f7defa0f6f5a740baaa1c249079da132e39da89
z9d80e788d0ded127752d0d9110797d498db5ca7a6312f73da55f0f07a192844feb2745cfc1d793
z95b15b525d7aae7c223de50a8c91e2763dccbe90f5678df4da4cc75ed56d9888d612b3c74fd709
ze817dbbd5c9be8a738cfb9a0b4c783ddc65eead814086a834a0fe5983f0a7145cc8582b10a6be7
z02965d179888692e23d64c080c555bcd20af15599698d4b03a89c1eb6a5bafc963084d35478ebb
ze39312b2ccc1feda2423eb1ca160b4fee8efcb59ded6615ce5989992092f61510aa002904a2571
z90b22089b4ddc32143a32bb60f879f11eab1b818d71da5db6e3eaff78ae906c8a080f2d921f991
zfb0e55ae3573f9ed7a473364d92919b2cbee9eb69828d4e2b8995a5e487a2c6d35de835eef6c23
z67a3c09b3e41bfd84736e91397da5a15dfcd17ebe6b2749873f7df1efd99c26af83241d5f1cc80
zebec736950f502999cfc57848012447df9ba09f73b37ddcd425857e5c5ddaab36095e82ce46f3b
za282c6640fbde4cb170ce9a69bbbb854d0fa13b89c4c5d1430e24c5fb0114a417639da3a82eb92
z314b00326b2d7609d273f710dff92eb553749a14fa76cbbb8d95670ab1818db66fd1f9ebb0a634
z03c9d95e8040435037e35d68fca0a385050bfd49c1d7d85aec4efa48cb2bb10aa9de2a6fa64fd2
z1d6dee230515b53cd46071d2ef0f3dd17eada0c17f257bfb25891df251e22b6ed338564730cc3e
z7a2ca89ed2dc330f2d58e31865cd174b3eb67e2c0c0bf5916730faa2f03325470bf16401963654
z5703536af9df2ae03cb63a3a8cb321796232b14ea7d0b5e67a4a87c993a0d9c5ba86c7d090b4f5
zaca80959f8b6d6f1e52d74505a822af5781a0b749df9a9f165c5e483c0b0a05cc47d6c1ed26fd2
zf357810de4857b7509192b2952fdbff7f2590de4000949d6257c2e28c7f24d80c2338c06fec4ab
zaed0ea169a6a95a4d3d497860dc4c112f221a0e1e1ea6de3de0f783d11da97c486685ccdc4f1d7
zeef1ad7aebbf1c1e798e0d5cdcda9a3372cd38939bf2872860be035862423a593ac872c9798e8b
z06459e6a741409a40a843bb0ce6b01c1ced8cfb37c3569055fd6c91bea0902438c8d3002d516d1
z1bb4cf6ba36b29ef767058763f5a142f68b7d1ed083a747d0158a5440ca5f029e891453e422db2
z1065430a167693b72ae62b47f08218f4dd5637825481d392af0f7b44654238f882b951e111d88b
z3a41555660854b166db3411d724b43a54db6df00fb002111fe25571e9c5ef1029c1b482faa477b
zfb2fe1d1983961ef59e7d8fe1da32e956b31aa3c3d9c12c669bf8c7a8d905b98002688af132a13
z36a86a51828fc9db2fa4a98f95773382b6606c3cd461472d3d4325fe44923514d244b55ee3c58b
z92f5ef84b3f43289fb2f59a590dc8d6a020e9f5c6bc739e1bda8466327da85e3ac995739b722da
z7986ea71bbb18450048cdb39b72d0a6775637f47ba40741df93a07ed57fd9bda41286197e91f66
z2a7eca7d662f6182196911879441962664d1bc795ece9a131cc8b167def5277bd634bfa6f3e0f7
z91e392c84ce42317802e05617789072e8f4cb88b7aa5facf2f49274dd9a22326e81440f10d381e
zcc643f9bcde7651e6e6fde948f0d8fc1c99250fa1dc11f969c94bcbbef4b49901db603d2cd4419
z2637ce88ff88d970cd071a5918a0805d0c65756741232ac38a09067880e58df95e5261fe8bdeed
z1c905531f1ccc0a38b6af0c9832b6eb4ebe1144df2421f407719b80e5538175c41b5d3c7858824
zdeb7b080f6e9474be5225590505aad218705143f51592f71b65ddddceac6499d531b2164094165
z29a3603e75fefe235d068312348b1c728b7f3b30d2249c1d9dd150acbce0a626515f2f9964b883
z30ed82d04d24229553e7e93e47b5dcb5b2e130031f42859aa520ebb41f03f8fdccc12ed3c9424a
zb4fdb83cd403525a82793fc1902cf247a422c99d657ed6aa66baf652faf16728fb7a2a8f4b5c2b
z3f301671f0df71154c5dc95b72b61b8095571527f9c44df105cfca62da779f6af9b2cbaeb33b6c
z0b967e10b2c51b1197ca2e477cc2de70ec361a305281feba7a045c40b3cdd363b441970759d909
z1f355c0453995e710bdeb561b340f70474e8d7571975cf4824bf5850a2c1a24845a6d2179878c2
zb85515f145d46c7a22ba5d561c52fa08057d2326fb86fb5ac3b1a389a0167348f707e75e8fbadc
z6d0a871b7060bc39da25c6786ccc628728cd1a7e440a4e0f8fb7b03d1b7ea502d60a2415cbf22f
zf52860842c92b43da0fd00465c6e594ef092507bdb762de88d57c1ff7385b69e4d0c2def204d1e
z872cfd449174d15e2bd8441d0f88008372ef45b3c430e1ef6d00a4b2a063c20f4a68c17d542489
z456bb71854a1dbb5a8d4e58ee9704c417c3181e9df3ab98ccd5e2c9059c0f1f62fd5fdad5fe951
zf5e1a2ce15bb23b1f9ba4262338944eb5a0c29f48e367c690adc495ca51eadf8ef133789971bdd
zedf428139cc9981b120ab9133746af6de09fea139aab7a9ee7634550f392d7bdb681660d7cce28
z6903a687f30338ef923f746238318402b87d1caaa000dc24151476697ecb00c650b4103b7e1e61
z2379a5b0fe72961933e27e676ba05dca176bee225fa52e4b31eff20743732d1e61a585fd72a375
zb19ea2870ad8759a41ccff2debbc215e79e624cbcb917cc46fb8d747ab1638c01a90c7933afa8f
z7325fb393ff55e023d84d8798b4b0b13bc1cb57c0dde86816209d08a409d0a85e8aeca844843fe
z010d962c19d39f3d062e1ecd3588dff033357b3d4eb9d9e77967b190cd998f96b05ab3ca959a40
z9019f4da315419da60cd38b8a78f5a7671227f9b40b71e30858c1325db20d6149b10df12e20783
z993597e871b4e6c5275cce589635cbde12c98d22ba5a0da1b51119d59001c57b10394efa504a8d
zc72baa8501f15a581b1591659dc437dd3ebb40e09a71a03010998fb79cf9036309f1e7f610066e
z5b0904fc914d5dca952c1e3c85e2f5801777b9545d24221d3344e5473380cb2413d9c403eed87d
z6269b5ab3fc7729c661e16aa04784024f401377d287e767af2a3a7e7c226b3aef6885427ea5d90
z554ed280025421f2ec5839c088e9d243ecee0ab02771e1906a59fa636e0b783a4877f498a60b7f
zf7e3dafcebf77344fa144883ff9152a2a16d76a39e089c15a9cd0ee5167f670edba85bd0b58f65
z50038b3a25c82db2f323ca9a1cb8fb785851e5d99ced10adee2c3ef60cc15d4190d20e970ec981
z215fe397e42666c796a408bd70705909ad1a5f9076b1ffdc541ecba14495afefd1e839b50302a7
zf936cd164331e93438f2ebe49ac15aff8c4004867802af130879fe04d81a4be29924d79be80209
zce3148a7a4bd1d22e92c4342e7437f40d91381af66b2b0ffc23f0159ec5c814cba40dfb622bd9a
z63caa768758bd0b8e752149b52837eb43856979900e14ad495c78866b6f900b14aabd2ba4505cf
zb725d16ef73c655ed7af4936ddf807460fbb1b28db9abfc1c1139ab3973b13f39ff9aee1dfd6e6
z9344721680451a531b07e44cd5ed6e05efc3bb6fcf830035dc878adc56cfe897ebc0372ab643ef
z3baa1d695a5d622b73f355557d3c73bb5d61d5affefe3382c9092b26557616b1228b4b044b35a4
z5ee1828eab30968ed654bee5294f280ac666d4c61886dfdea6d14966b58f44d5fd2ff34a9b0e74
z2be7453c8b843dec539bc33355bbe1a2a8d19110f7eb9ddf4c2373c7653fc2dbf8acf6abaef8f8
z06aaef870f91e5dafa97be5a49a31f69f81be3abd2091704dd16185785f2718db1439c5118de65
z0b4c51e0fc63c75d67dcfc4db17e4d1d45764e711429282a52b40fc1ba9155828c2acca4649f5f
zb1389c8171ffe9f9b59499ce67f3fdbad4e4c76350aff1ba0abe01b69fec5c8b1900ab3a871486
z0f3ea979db585f77539b4025dc95fbad5bd0239b38ad1c29f4ab5135241f9ed21696befad31946
z2959014e6585a82d7bf952ec5733c089c9028bc55474eab012c240329c8ded0d773e14a16f2780
za397e7aa15113f55d1f8b5aef95257a629f23f6fde271069b772761cde2ceaaf6092301d1d1ecf
z7ea85c0eafab0f10f7d339912bdda85229a25ddacd204c2cb8c5231ff2ebfa61001f3794aeb149
z4b37ed3b7b50d0e16a3806593deadeb14bee4ee94663dd6ea9de518378624bf971061c16fec3c6
z553d01b905ed14dd67e4d417df29ca08acdc3636ed81391acf1bf37c8d41c7d11b133f4514d362
zcb95050e4cbdd92efe090bb941a706720890e67646a9154ea28c3bd7faee4efc06b6021f38c487
z7442a998c52370684b3a19da70637603dde506275bb51166a7c8a20da809a9222facf2dca89f77
zf4f8bb987b6884832501279f042db831cbe6fbb0dd413fbf0654004ae86521ad97537d174ce448
z152133170c4d091b34de8308f85933ccdd059199daed4933888d499741c8a738047ad0b5c2d234
zaca9ed9065392d25b857303b2203bfea926b8a7fe5585bf197f8d8da7b5c3286e485a86a8c9c3c
z88b7ca7e0a9edd1d40312e07180be188b8a7babeff073a7cab168ce40e7174ee941b78872ca9d1
z956df52d6999dfd27da7230fa605616ead1f531733d9037c7d13d7f1594bcc98a5b157c7bbd587
zc4e0ece2f0ea7846c0bc6285b1708696c23cd5fd3583c8039cb1de2e3aa866bc5d88bf01fec095
z459f95f3102333bb8299c4314ea8e7b943a074cd59ea69250a98de5096b1a654af386341f26b47
z004e281a4a0b42189191ba65f43a9718bbc301a01dd80346c557d18d4d3470eaab0ae1c533ff21
za9bbebf0fa16e02711794f35bc00751946ee911c350f4812eeeb2835caf806730b45eb26ba6fb2
z510c5e373e60a386c2ab9815dafd876bf8ce3ba8ce453c53b99f58c12dfaed74e01d5dd042d34a
zab7fd4c1f5cf251ab67c06fdbe0f270d56004dad7bdb7e134981e2d9a615e0858b4bb428ff9d1f
z333ab082d2d9e4fe6d24266f002f056f11d1db1fe74e98d92d88f5f66c861ec41fe012a212e2a5
zab23c16e6a56a80904fa73281b87839706c26deb480ef180cd439df768d19ed528ae36c8441d88
zddb5411841ad5b6621e69ed693b91e70191f8d9a04eec9bf3468469018e15d3b11c70e7624631a
zecc29f4c17b9fe9893039eb8aa93790957cb1c0048af3e32224bd9a90f73271f47ee97dd4c5d5f
z85c118928cb0e6c0d86f616ac4943f0d1cc284327e218a70032c62e128e58fbdd69bd2190ca9e5
z6d777c86b9db299bfdb17611d323cbd3e26df2bfbb60d871effd17fd3cff87595ee11bfaa66493
z14af62ce99dd5d200eed1bd87a196b6c433fa75220b65c9b6cdc47fdfdd3cecaf979881b920aa5
za9256cb2c648024b3532b502fb7ecf060a2397ed805f032e97293d87b16fd5970e0b2fbfc18987
z8306a4c34e8f51998bfc5390194195429874000ba4d11fb36d0187908cf1c230ad1ac6b0222fb6
z4d6990af37513c525b986295bb773cba1f0b18bd75e615f4283e467132f59a819b10d8bd23544e
zeb120f2d6f89ed8b64ff6ffefe44d4fe2057b57747be2ac9217feedf45e7a771542e80cbe987a7
za86d50001dcabf5be2fe3a51f10ed524338cd4951ef02f076a4277434d0378ddcc8192faaf2257
zc70d0c11ee7ca57736e2deb45350fa082105e3a93b684d86d49dd9c2e235ff7c14d8cfceb8f772
z245a3074f57a8f65a9c4a7afbae72b9de20abecf0d76bba5d6d53247cce112e35373197ebff463
z171bbb423b3ef0a3c6a69062282f668bdff33191cba6cb3dbe8c263babf6440faee815fc9beec9
z07f82b9e70797b730a25d40f04631938b9694a72dbd636b6e5466900c6b19b6a84a095d58d3181
zef83c7343b313eba16854e3e71fe50b958b4c6c8432d2c1e6dffe1a9bb32bf7fe30b0f228984f8
zffa06c3f5a5cb3a97de5ef523fbcd9e6e1aa5d6251856b065fc41891a15cc172194c22e8905dd7
zf5a7bdbc9672214fa61abd08bf3cf8b17f9819047f532b45f42154448fbda641fd9c254eca7bde
zcfb78a80ff5f9c938759a070a19a91d55aa0785d91049d016e90ad766242ff00c5d39065a59bf9
z2ff04e6bee08f8922e7761aa342eb4dae021e4a72c216b0ec16e833b418f2644dcb3bb4b5ea293
z0c2abe2f8c241aa22c5bad1cc7a0a5f15764827b20139149d722f4af18e7a75e80c0306439003c
z4247224b0107ff407e66f04cd8982c1c931c4e6e0f43be92ec6101e7d7fc98d4a604963d4e38cb
z6d131ee3214aa64a0ec898154e24c2aa537c287d4cdfad2ae108bec364cc513427ee510014ad87
z188dd87e3f04360c844106a87ddf5e9855eea5423db7a9f68fc2b7fdaa05b9e21f0b6f9e9d4d71
zf65eadfb1130af7774df2a49d517b9d81a7a1271ddd912a910cd3ad05edd5a5621491d3c8ed77a
z5e02ebdd90d5e26bc270792fe25a3d1eadcb304ffb3119eb63609aa96821c08c213a7e86019f7b
z434acb4e1f891060077f3589007d2401efe3891ceeed573c7cdceb195dac6fa72e94d882a1fcb3
z17bea30fdad396144f965bf1e274299f82e90a681e3f195fc35e3f2aecc77dc324b2d34b6a51a1
z3c7fec091f3259dfd51461e43ad25dd46240d19b0e2bc99ae748a289929a13963db8a2002d8896
zca004687606404ccb3ea873d398557dd84c891808821b08250a3392335708e5734e3411823d34f
z1cc2b3738200e2af78a65512ef0301344250b97e486d07c38815a2a142ddd73aa260f2c0365ca4
z60960e5afc503191855e4ff21d40bc65e6b5701da57a4077bfbbd32955d565a3ee9d583040be24
z72f0899f4f4e3f7d55e52e636c7c529681521ff078bac994ac4512d4be7a6fce3d853994856a1c
z3ce0f3b13f2cc917234184a50a020c191a54b9cc1932f320e997f9e0e21a2226d0073a2293a32d
z770975b1070de5c4ade6ca7298f27b17499492f3acc6d87c9ee37f94a38e101fe2ce3878d93a82
z02fe425bb1712d16a961548fa0f9d17050df1d736e0c04e7dcb0a48311805fea366f6bf5add9c0
z36be24b0a624283de10bd9e4c98daaf38e7b142a5539d9ad971fc828333b7c6e2b4908b736c87e
z1e0dbd800d0cd2a97eaa88eb2634cbc72176413be4c28d344afd15d5cc3d680e5798b5468637fe
z7c81fb5dad3a7bf6fae419301c56aeaf5e50422e704d2af2a08e59bd4fdf14f66408a6a2db7600
ze5424caea60a1147347f7aacd06d0d373d1ed1551c3e3ebb84ec2fd8e4ecd389f270d38abdebcd
z928e01bfd5225eed940a1e7fff407b3574c9bae95d3822ea7f28fe1762366e4c440dac0f3f1157
z1a542a8ed7e2c110be2958948ca7d163f6a163a70a525cdf60c32ebb155923f7a88bc90dcb8ffe
z2a6df039638230d49c58c8e1ea5d27d156a4fc82b4e2a83722f90917cd2d3ae5133d32cdb8aee7
z516d36b1782378fdbdf7a15e3ff1d7e5719070ae92851fe8b608252e4b05f49d2ad3363c545f84
ze86452d0310797b150eb063b78b4d5810dda14091f85068b1a2e255c1fd4b744f17c29e03124ca
zcb5ef16e50e11766347df11098128b648d7200f162757a1ac34c1a5b8a50fbcdc7e28a75f39d80
z19d870a233b3f60ab0ab68f106e58a03ee948d855026be28dd891f20637b7fd604ac46396f7764
zf1b3ea159774dbeb281432822a41b1737d01d41a1dc301d27d7d7b02d6934190018d0f029e2345
z7b146788d5b1385863bbe734e84b6f4d269a160e1d78394be9195a1bf95bfd8bd99d1516c9bc62
z8ba12cbacb99240bd7cdf3fb3987a02e61e3a7eea0b279988c2db7416f320824929cc072236142
z38ed3d087283d7e00262fe1bf2318efc32b01b7aa82cca7675b737037cefc2661609b2b25fbbc4
z65717039c5cb6639bc36987ca236abcbd97dad8c00cbb0aa105cd67291f2645dff06552b84d2cf
z87f73eb545770d2a6762fa488185f486e625dfe1633698efe1a8e9ea59f09ecaec4ca43951ab5a
zf6730ed53ee1224291c5ac28a952fee77635c8a3afc313194a9702abe0379602397e3d4592c2f1
zeae50d87e8dfae5f6b09edec744e9d0337d84ebfc526460875ab5b5905eede59a15a056738dce6
z692c1782ab0b63ebac7751dba7d844cf7200ccf40d8bbce43ca01852ba8e43e1e80c6f4ff6d2ac
z8e1e013d322d6baf8ddb90e0f2d698480ca817cbb51dd29de4f599444f7044681692ff211fae3d
z099deb90fc2eefe8fd52605b26eea2f94276fc8faf1c54c2e220318996cc8404f82efafbf69581
zf93480db92a6027d1710200e42f3b86eef50bf20ae4c01583b85cbf38edfd15dd1ea949bfd746b
z3c298169749365ccb1983178cc0e1f2d6b720aaddb8fbb268181861c9354ca0da3a1eae95131b4
z92d64dfe12df70f3675eab09c9b34648793bf5c76d2f87595b92b344fa9326572069c2fec95881
z61e5121caf64927f2c3f68848783ba1364e53602558d26aff9f8e0d29e9cd5b9ea3fe19da7b162
z36a032916a5b7ebdb38b0dc3235cdf13dff9e5b3aa96e584ebf2c2dbeb58bf8036c8de39a01036
zfc303ae0340bfd936cb084e34ca73085ea9c68db02d66618a62f13f8067b712eee641a18bef99f
zb0e5a0f90a8a1220c00ea061654b1e4f086f6ae2a64d42ebef6925c6281f0520bdcac4331fc390
z6035e343457793460ebf285ca6bcf9cbcf7b14e17a73c48c35e4423ae4d6bf72b4d2746a465622
z043f07aa9328ab97f9b521c410903e24ee84a321df7e6c69ad20c235a2e3ad7b56c90cd1e40564
zb5d30c3096e66f6459c06dc367e2a20f878066790afab401d49c42e5f9be1bf022a83e713de728
zf270190a2992be856fb5e5012c9bbd27809e14938c74534e747b9d4ad093463fccefd338107253
za5edf3baccb95c2e9aa1bb38a0084717b9c0c4e7d059b6eeccca7bc54d080ab99e99a6c4944300
z3d10edf295c7f14c2d804f486b3f94c50054998d43bcfc992f7ffe63820c34e8ee98e9d2067845
zd97895049a5bffd0f1dbd6ba881074a62abf77dc9cbbc3adaec7fc0464ee86aba1703d0a63d938
z74a1e5ba096166c14ce1c39ed95fc907cada5434e06133454860e98e1686d1a279949a1ad4560f
z6ce0d44ef7d96263eb37b143763f14fded3ee40b43ae8bc6999be68e6714f2694d56c903e949a8
zf2bca50f0923c8e1eedab4f76ed2ada07c70023f9b8be5708cc0ab9ac773d8138a6e821da4b164
ze04ff5269c30cac5536b6eb0f3170f804a7c1f6fb1ebcdbe895447355d8af73f50eeaa5d4e9cdb
z5b15c629c6763aa09e7a43cd622baefc078343a571ecad96e58ff09dc2884024d70165887d27fa
zfdda6a07758282fe52e9524399e98510c5f9b7fcccb3d0d397058be2c99cf4c8cb5c1c6e1f20b1
z0fd236253e830e4db16b38c7b78acc92fcaa473a726b5a92c8974227b87ac3dc7fc072fea2b9bd
z5261f3acf288d80ac205c4fc707e3f623c58ad1d39e2eef4bf4422206ef67588a81a1659779570
z6e744eae02356ea2b4731d81542bea91f2effe0869c05705af28a38089aac5442b0973163d96e0
z8641f2ff146ebf493446536a93a344a3103d801ef16ce1f9aad0c5aad4e9e8ace2ff65c9582d9d
z8cf301e613fce9de577480ad3fd27ae5c9ca4dee006dc30fffcf55e629387061d99543e8d2ba3b
zb2d80c471dddba06b59de0efcb6b6455e97f7d0bdf7b13e42134c64522e474f2522250aa2a6ef4
z57dd7befe0dc475e6871255b93186013c3e35fa7f030e8e06c27a00c0b113cb38205e4727850e9
z26bdb62e24862c93c130e9c94600377eb9c27da5f027b20d149c95f710b268ff0c62b91231e8d1
z48070af3f16a35129268fd2587d89b317ba9e96bd4bef3972f8a95327b8ebd25b1142a309e8ba0
zf77deba101eb74a8303b4c4580235bfffe73430c04e3fceb5d82993fffac3b4768c71caf148ec8
z843acf03f9cce025b94cded970b3c030aa115835221a4308d12fe1e404e12db7c03356bd2c408a
z7f0288b3bee3973aab7f78d9f074be9df65f4787fdf70ad5784911eeb9667edf9181fac592cc96
zda24a0d82de32138a93b8df065e8728d584356fc7ac5d623d91095bfb6a4cce1b41aedd20d4d84
za1d1f6ffaf8d3edc5079fbf8dc4ce637ea779e934589c6c9ffe187d610bd0b6be9529b1b1b8e8f
z42de3c348861546826d54a7d70bc523def638b78c64f1865a152a719da872539b02f4cfcde6085
z3c7a1a52935618eb6c7b52107a5a71bdbc4db8f841e4040d4e8d664272984860b12033b63a80c2
z6a884dd655e8b93663755bd495f6ae7f7ca45d63de8e7df72da5d175e0163f1fa110099786c282
zc1eb831f308ffd9e356e49981b0eac523da4bd2fabe3648f49348685c4a4ea1f3ac3e42494200f
z93d8044c034bc6f6d5c00ef7959f68390920e11a87c8d286c17face43662a9e2a69eae461da571
z6b572af9f5d1810671c39df02292d806ff1bdcd73c464ffbd226177de5f578557e866cecae3dc0
z898e157598550de5f873b3b6f9a38c0bd6f935683d66bdcb41871d96dfee5fb02a89a7400bd37a
z65e2be6303d87e44cec07413bcc3a83511e5dc1ee4f7cea6018696d6ae64d865a3c44206949de6
zd95ce6feda9b84416cea6ee61f5441d9686f78daa4a18d25522397ea5c24e3ecd470c8e1c47006
zbad936def2969a5febf71ca78b53c9a25f9f2188a9176a212ceab10b4af7389acd9bcf98eda1c5
z736d036dd219c8ea9497d7a0e5033e7ca79ad9094e4af67c8a47c50bcb63ed032667ec6f5a6136
z3363bb410cc60c66a5198e8cca3f131c68d429fb74bb7822ac2d0b77117d3eddd13852ab80e04f
z19f9b5837f1ba8da1eb8d801cefa707c6e17ea3263fc02f9613220c1a8323fe47a634e46e9f51b
z5f2fcef92059d172547970314e94e99b5bfa62681d0c0bbb9a6332dd66f85486e85cdfee486170
zfa0b7867ab1cc4429a1c68261f2598f7f74f7d46950f1a487cba367cda5ab2716b0f8296699bf7
z2c90d9bb8b9636044db895e3d3f5c2ce5cf1ba728811937a32dc7172f6e618f363dabaa61d8e50
z15481c0783a21b66cd2488dd0e77615bcee4b833f74aa163c1275713dafcc282a3b49891676a15
z90ede6960c5a30d00ee3378bc63b5ada3a97cd1bcaa07ceb5944c81ad03ad9a1ac9451d45135d0
z2c8263c368c8fe92548e57a284409878f258a1c2532d18c83158b1380b78d7d2e3b0889657ac6b
z28916723122603a859a00db9e557b246efe2d487811e3d612fb7aa1a9131a2098cf5dadfd9d50d
z0d662fa454682de2aceabc64ad902bafcad2076a8d6beabdea81de9bbc21ddf0e6b13077ed89be
z6bac48b956959be62e8e6d4a95dcce416544f70788e5adb556532e55549d4a4559585ab410e883
zd900292274d1698039644de0f28114da6eb8c8b201ca0b3488c1548f7bb169572cb709fd78205c
z30ce506c655dbbe7e209d511c276fa39c1102cbe92aa99fa8ce3704b7c137db4a66a798ea09b48
zefa83af2fe5d9a5bde7c78e50918d43fcff23e02781a77e895c4b3d75ab5b4b8b88a11c8e98186
zc5b94a4de675112b003e3cb2b2047324dd3b3ed262f1e030d0d2d6b7d470429d251a66217a706a
z876d8284feac5cc8c141f2b5c8a005e0d327660af42f8bf309a8630006da5243c7be8db73afe67
z23abb4d62a671048a3a80f3187a6ae4d3e28b2461da876a9f40ca96dcbdaa344402954b0e06888
z7872c0b5471cff1bb7b273ecc41305b67da1fb780963c014df757a34361dfcf0c8138a0f026961
z63adc7a61e2c2bca54f8e557830962abb5cc499ecb5a992b7ac1f7aea9c41fa1ccc32d56c74891
z6a77276c404e201443709c77d099a5cd4955b296a2f25228625f4ca2c57e4629d22e0b5470ebcf
za51523406288e0c8b2a3412e997b38c9fb435f8e81f58c8cdae6a282e209a1e39a6dd69fdd89f6
z9f5223583d9eca4d9693610642024e104b7ca9baa6ae88831fd108fd86007d0bdb4285fc546fc0
z1f2177752af4bc2efa4560f24992f7d90f6807b83cfe82dd1f8973978b054fb462fcc54cf908ab
zfcc7c7018c58ec818596369fbc83412d2333f27806c869a279c74c9179f87b2665058829074a76
zbc52505f14f9bd210a721c28fb28dac87a13e5c160a82fd533e054045f902766bb2b54ea231567
z9dc4b27ea482d13973158769ef369a7093c836d4515e16c8fbf04616d42f66a47ffdcc620449df
zdd1d2779aa9b347690bd263f706bfdfdfc93868d9e21a03d3feb1628f6d4b8a78a6a5535e515fa
za0cce51e9fe7cd9c5819a4c532584e625a217672fb2849a9c8d63b10603019b86ba38136fe7ceb
ze889dba2b030b0b008c33d88d1e3f1e8c61354cf597a88cfc4e93ef9eb562a0193b3e42f78032c
z38559f47a75af24f29fff61d650ab937fcd69361d1ed1e6636fcf31c61dc0b94c72ccfb67302ce
zebd06db6c118ebb56253f344f9c9b10e9a0797959d707f3dc226c8c8ca608adfaabf6008ac4146
z25e781917e24793a5c4f746127dad559d26edb28058e7c4ee7ac7b8aebe82a39740986710f25aa
zfd8f1e49054cfd9f3f57253d8c57df13dcfe410cb287f4d5d94dc18006892284d05ffca2c94fd3
zb3a4bfe23d36a99f49ab75b06cc7e2ccc6dbd025bd5f6f62febaefbc41b01db90b83a8795512fb
z12be32183b7531f6bb1ff2dcd5a88b1ad31c4ba963b678cb8dbaa67ef443a9901e698a14904c4f
z539286ab312a61b3f8f5acab4df24031556596c93d769e96a62bc7a47917222af8a00c54577a69
zc501b96d340ac88e9fbc0fcec5f2a6a87194ee713582400845d1e5a9da377f4d63ed1767cfb952
zfafee710acd13631325324a9fb04e34fe88981ee2a95b583e5ebc24de267ecec9307eb878f06f0
z268126cf95922aa5bc36ed1cd84074bb4c2498dcfecaddd480eff05059f48cc246da00f2a4f4a7
z72d048fdb0de415a325d05071f6766018afbdd35874a930c2623999e3dc88ba904e97c9474ec99
z8d69142d6ae31a6b1635af974937a87e4b414540d9ef2eeba45a25301956873afbab1eb5168d50
ze7d63415109aa1ab35122a2531e63fb21d4c69fefd688d08c1b942499fa35b60415cfae3969970
z07cbbc62e3fb12f0d7a8e616e675d2810c07b0d3cb28e6d073dc686ab0c75a016921b1498ccefa
z0fde9a87fd4743dc79adc2f97a99c224e6f9e8902f978fa0961d664bba91cac041e463ed29d3ca
z2e37cedb2d4ff4a0095683a234d27244bd719b8c80bc4b1fef4987551efd92495061948b72c4e9
z3eb8b5cdbe1a26f1ba37652cf11aae0e099d365b39a80486bf14318714d37816da9c9af8a61644
z982d749b370751ef38c380260f876c36b3ab7212b08225a522b8431f083ae07ab4659378a6b140
z91917e087738adb18d72813b2bc15f1294ff1dc9c22ed3c0f4f3bc56120f07dddd6eef9a392dd0
zc12c79c8c7c9e1ef823e2f02e866705a2dcde36796d87f2ad3ad471fd5c396239cf8208d686a1e
z2b2d14f3cd42d22cf19e51ab953d5ed4c0019bb7f6e14186f31da3013c36aca282b1cdd16378de
z99999c7554a3e9cb11e026002306cc117ae4f8ec72be850e12fc9e9631ed7acb9a084fb5284bad
z58705089303794d002c3f9df4e1a02a96c76da957d56be343f0dde22ba652d70d8450931dec1bd
z8d6067d86bf945c05be836611ddb056904d2fb2ac79669779c8d22accb21d4804d5f0471906c84
z993e5c9c18e05f6f18cedb4e3605fde056716b3a1ff208dc649b088b2849cab4f207af25051ca0
ze36d3a2ff064b022ef60935f8c966704461d6d3252fd0d979c83f82c88e6283dd9c09e904c
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_amba_axi_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
