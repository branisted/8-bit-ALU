library verilog;
use verilog.vl_types.all;
entity mti_cstring is
end mti_cstring;
