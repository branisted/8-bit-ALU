`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262e96b75598c81b19220790e3a0d
zac0e9cec59fa3a7263133e4e4c54ed27d6f010cd2be3fb7767eeb444f708ca477cf85d225b3317
z483338cc9eeae82f9dfb824e1f141e648770668538b2138cd99227531ed113e33d2dcef1bcb10b
zf455eb9866ddc8709b87c30e446e39255957dc030b8b7993a4b340a3c9add5dde303f8c4126b48
z037ece6695fd4de69ebb5786a0e8ea19034124ec30f21bb31e20cc9dbd07490ddcd5e0e8708a1f
z7eb436832f866195b21071581ae532bdb5be5b63ab5c1b94a872c6ed8949f7672f7b9016e8f30c
zb3304c03bcb8acd193f90cfd52a9c1341c21b0269f1f21692c29ff56e82ac85c79c9fb49e5660d
zf127a66f269a2fa1d228670e299c178dd605bedb4a4e9cbe114a4f9b1626e2f96939112d96ee56
z00897141aba1e6833da28a3f526bfc33ed2296967d2a58dfeafb1bf8d1bc422b091c8e672c953a
z96c67bd4f53248d0e9f685aa362f9ac9cf0fbfcb021895e6c80d3d332925aa10736e73cc065ba4
z6ad4c3345978f11659ececa52ac516a08cce9e93c30c2e3597446aede49a5b2493944e743ef856
zd02113d182e4e5126c20081e0e0ed18b363855e92e7f87022ab4d69a27ecdcb37cad48d6cf746e
z6d810ad135fad6d87854dfe4a3f604b26778aba4b5d4af90154614d8c202d4ef8fa79a74d0dd1e
zee59c6d188411da107caf5d6a0a4526123f018a1f427d853fc669e0e0066e45180f07ac4db9f23
z3ece57d81556ec4f96f6a957809b154e9422bee2d7ed835a2a10ea002d17274b94612a82a6a90f
z1ee9f7f3b6cf6a1c8f78f813c6e519c6730a3f87eeb59cb82545e050a3aeebadbed0f9395833fe
z442d803e5c908ea84076996ae6ab24a781653f480d3a285c73cc01df63d671bb28d1d705be0012
z42004d29a8f5f124ea13f77ac4475a812ca486aff69f0d20b27707bf2b168bfea1636408f46c0f
z68f5b8e44081f5ad31c5494ab94f74ff0f8307a62f61bf4cf8005241a14a827138132b8bef6326
z44f91e283c506c722e9481bf4ae8835bdbf1a189b496b3acbfbdb83478e2ff7e90b4767d3fb9f1
z9ecff137c711300b8a0bd51eb078900119f2ac81eee19f7284a4d267ff7512cdaed5850908a3d2
zbdfa322ef8cc3756e5a607783b2cb95ac2ecd8b9ca92a5202f502629836b3d53d1831079fab739
z694bafaca865cf5ea1e7ac932af810ec4cc7e6e28fa59191146144372c26d618e1f022e9625a46
z3c51e96452d28b97a306b4fa340ac7326b0a841762d8ca0cad74d7b919bea01da2ee1dc6ea02c3
z96fb8fc6c05e0774f00a59eef5800daa4eeec51b026d8d514d3b5eb8090c76698600f92fb5db22
z4186bb12a15d166c33525c80d7442694c2e594e6cdd9009f38b573bd4b6903b39e57dc42122bb8
z42aafb2ffbb51a4543a02d863a8edcc2a9425b896d251d112e635697eed68ecb8b21fec96dcb31
zda493ce291fc4575856a92045f66d5d12baf3fc5a1a59720cf23858688d51406b44dc798aca90f
z9d58f898b9951fcc730d88594bfe216bc398e388834ef85dc27f8e56ba7c5af464d86ef273d5c3
z89fd230911d444950311c075c3e5a4e2748f0115f74f686e941b393d174d5c538a9962e25814ed
zffc61c312e47cdbe906300e8104081396f3a30bda9edde3b4b8bf14b027d81b88bcd4a2f5f538f
z5242618a97325187354cab0c4eeeea0a53f477c368e1c775e04b88e5149904d2dfd09845969786
z5f8f6a258eb120ff5bdf189448cf335b87015843fadc7fc7cfba2c1f6b11b1166c13991f9b1a2a
zc48926c0bf1e5d3fb55614525d8014896712fd2d33f5980ed15e16286ad8d0761c5009a99e6a68
za93a1ae2cef58182391efa3d50b16852c38331ba591a397e631aeb89101eb2817f374404abe243
zc54ddbcbf1d11abef4f57820b459d2ef83b5309e8a7e3671f567a57ab81fdba6cb05659f1a6ea8
zed3c203a9d169eb42d5e8deff81fa6ccb605dc9f280c9dab1917120d8fb1fdf20cb0468519bd3e
z1f582351cfb90974a3e0519c309b898cea7760df5f7934b6a5deda3b67953d0b6b2522a286c069
z8b83fe4c405c826a9faec56c928903dbcb3fd02e7a9b7bf6fd08a64611a31509f8162d9783e342
z13775fca4745769ab5666759f92bea180deb521be662678fc004e7740b318235bbc921ed719db0
z1f7660a85a5585fa3568fb4c46bb23c39a00153f15dfb20baeaad4c0f483275c1007f1ad399b58
z125e659b881d80406b66df4de051e9aec1c9341221b8eed83e72a29a339efd17c5a354c428957e
z1116d833e3b2058f6cc7f680f90cf2026de87de40d64d7d0d8ac1a000815a4098c2e74fd9e2bca
z42a67bd6dabe291bccc8a5deedd968a7b550da485aad799b611e601b8a54da82bbc287c1e935d0
z9eec09a7d4025cd3d89a4ed636d5c3f3066c4eefa6a86c1f116e2961da6be497042264ef0012e4
z024b30509df326096d9fa7fd8f723a826bf2112941de543cdd86c16866ad798be0082a6fdebfce
z526d6d32f3ba675a6f8488ae8ef9f2b7f5f523827d4190c6ea5bbd13f34a2c7c570d21e541f882
z38b912ba31a7eb568c5a271d6429a3a1aa044000cf6d9ecea7a9628bfacf70b94ec0f18ae1f2bd
zc130f3df07f746934e758657ca97e6f5204a507a17358581b0b27c7cc6bee9efd4de5037bd4b30
zcb617a4675afa0bd00263a51a540e6b93ff6708d5e3f9e96ac5c64ffead00e9044058a1dd484fe
z3ea83a038f6c04d4d7c866d47f8d24a78abd9ff9325943f579a2fbbbad1c61cd0a4caec8b2c29a
z44f68c9fc144e7cd240245b5794b2dcec8aed1f008d802a5e90575c2502dd07f98e73bda37fa33
zf0f8be82c9e1acef44a006c76738759282a4e4777715e44146df6d3634246c44c62c5b418334fb
z6876cc950c21130af44c683108ca050f4740120ac3cde1b548273a5fbaf4cf04be5a855c242f65
zd8a1408768d9d8fd3ef722b2507e4694b9b3b3060ad0d6f5b84ce8ccd26a01ce15a05dc60ebd75
z3136a95d7767e5cd2d44340773a2b0e0ec8ff7108d769288d54b572589faf8699d73c8a5112035
zd0437f19df6327eccf6bca0e9d2ad9a74252a47390c09876bea75ba5fc07a472e2a34bbd47554c
z3d85aa4f79dc98b101e978070cc7aeb210d56749658f3e0f192e5e303cac2b1985c6e51ee1ed08
zc0977720f0f165d35430224f0ffa2f4e4f0ebc5520be4c8d6e6c70363dfd6320e4bdefdfb932b4
z56e022c385b917864eeeb1e3d23108ce42db4ee194eb8dcb9e22dc88edcdd53945209bc39dcb5c
z386d81402b2f5869dabe0e36cee2873b443541c92bf3b2dd0e5079e5746f217c9b562c840a9718
z311133bf2c39999fbbf4705f5658296a7f927a3534fd7aed097cabe26a2e0c4e945250ea46c4d3
z00f14231b534c0307c10165284cd689b9cca94e223a790d093c9be88e39a87d197f892f70aa976
z3ee8c47946514e8c3d9d6a17383a1745485b32cbe14ee25b69419ed677e75f86f1efae70e00e92
z162565b35d149f7d1e91dff1e7ede6449a0bca2fad462d6951767b0c60984923a7f6f0b715f3f7
z248c4ef88ceb06422c46243d54b43d1c520891201c036df65cf17043997a7ee837112532808a82
z36d6c57881f07e08038e4a8d4c746975a9dbb40ad684dee7bfa5cd7348bc375afe6cc26de563d6
z4e7974d6e35b276c42228059ecc9b5ab69805802f63a836f05a58ddeb8f3b213faf8f062dfea98
zf29335a248bb15327d1ec3cd9b6fcef0dcffe8b1435f46e035551c035896da1a7733d4338f15be
zad305cd5d2f3b0ff92dafea0bd6a6b28939f173696242b63989bdd6446d4c9dd2e5ccc56406374
z7b0dcfd072e0f3b1651647a83f9249f813488b58c829b000badeb61c04012cce70e7cc4f041fe2
zd81d03ba9c5cf99113f47d34ea6968d2e23b6730b7127f5608bafdc3acd940c55fdd7484fe5566
z1818d3606bb91271e17476accc48a98c13306ffe0d0dfcad457cb12055def86dd94d97171257a2
zd76f8c33b1c80a9bdfcee74d2fe06aa1a5c42775cf60ec01a5532127fed501537caa7309b59aae
z9aa3debe52338c4e0f7cba11732f9eb7cd3db5e4e76e4fea176f9f9c8a82b0a876a6c3be383b79
z972781782cc470932d583dd37f10c2e9c38de5d631fffbe1378b4c37ebfa5302075b1beed5fa39
zc65d9fc6025dce01bf3b4cd80e636a659d0edfd389c21d0050b09dd278cfee7c52a0aaba6d2c69
zb5238c75529643d1252531fa6559cd71a74f707ce227492b208c3a3f14b5d2dc961117007e63b9
z5a1ceed438914470bd2a6bb0a35a65424dc573fb174566a5903b4502b77d2bd088dcc20c60082a
z12b263db60a8be473a4a689e5754f545401ebce2a3be6261ce45eebb78fa1534c0143617c24a69
zd2a8013adfe11206b5f3a32aba356123691503351d661353c3304ce701eeb13b83e9839d93214d
z326e939345b69d3f8e90b84c77bae46eae6a602f2b3a3edabe6af8ed3e58be764a751f547a22ac
za43543a370596683288a1fbeb5ab3463b67cefaf4380cf111c65205e605b24ce4e0db0b8425da4
zc1ccc887799788374cdf733c924ff6fc359b442a952f6b7905c08fe1fa239698b7f3037ae101aa
zd8a2aaff200b68de3dda0e8da903f4e3b6b5c6fd93316db38735f1e1236c51775d93862342873e
zd71e97c45d3fcd1b280f200bb27405af486f6bc2df51462e68fbe10cd301fdd52639cbddad52d9
zf161c246448ae46bc9a60e7a766ed70cdd8325cbb7fbd4504732fce5749e2a6c3a90781da7b319
z9fff4fc844ab23173c956d13993e4e1c384a0aee684e796b16c1f438077fb0563000130094a5a2
z6227ab4330aa49d4029cd6e8a5e9ba0a6f4c470740ab2ec1cfa4fee41c4bece9f2c65ed13568d5
z719ba4512f22da9c6213ebdb4f5ad3d05ebc4f796808472c7d84d98d92a53e0129a4a9d8d28768
za6469def3777977afe4db36f1130c5259cf2ea12632861acbb1872e6811ae873997a191135557b
z1b2ffc06ae0d086b17b9364947d4c5efee773d166140cf6da2644ea33802014e390c7e94216fe9
zdf7282cacab455693c646fc346c775ec3a0dae47e919ecdf39dc5f2b7477cc2c7e9cd76e765c07
z8ea4a7971dbcf74ae9d43b8d97df28dbfafaaac2e1985e5b1a4f3c108efc35de307db88a213614
ze3e817754b0fa7c0a8385d871740017209477f59c7263491d8c2dede0627b69388738ee7f5c462
z75c6275946d655c9021ef0b634ff904ef2c807591c5a9c1773464d4fb2a323a47bddd8b1bccf79
z237bc57378c1d875256d6ae847703cdb49e1bf9b30ddfe520a41e89b15a1e6a2cffa8a80a73580
zb7d4eef6eaea5fbeb593ca7dfeb4c1aa3d605d1106612f70edcb2e6a180f25f2928b6f63fcafa8
zea7902e590aa841090081d405c3e536d9d86eb2fadb44451a4397e0cca65371ec39481423bb7e6
z6d5cb8706ac59457b4f88222835090952c30528606a16a86fe520ce2af96cfc26c32ed4d23334b
z4ee02453aced2084092890f61bdcc2a56e33fd8222b559a1faea11d1a6bb57c269c288b4b23928
z4930140a57cdd98fdd2839ea4e425506cedae97f72221b52662af7f5594478bbe88bd118ab27b9
za5349c59caa5979064594da7b4673a3cbd67b185b5ea9c4cb6f69780fef3bac34764d15c0a685d
zd914317ad0833d026bbf94327393a3acf59089067c4c9752e495c2da405326f677098cc1be51a6
zbe4642db8fdda2ef49358e5b0c6a1664175413985b00acedbdeb07b55b902cb56d91dc5450040e
z8631ee80d1459f2e112f8a86b6bd2aef7a455977ce9c6360242b9597d6427e097d12b4c7d7b0da
z158e80ec27d6e9af50000acb821f224d5d940c959faffdcab8ac5d09547ac77bfddbd0ac964779
z005603c3b2a0ceebd22968615b19e537d6b78a2259760fc0bcfc1c467c53cf7c8dbba15bc38de1
z9f5cab1eda4201614220b64b5b0c061c37c656f79c278084a0e89fe2b0f7461f2268b5a6608234
zd87c72fe8e86d12160830f380ae89bf29b5ca2c77ea5f0dd4c1a02cc2ff6bc6b94544dde9823ba
z6fb992ba2ff93489cd26189abf7618c6caf352120e37a9832b9d63c74d1896f363c3d9183262b7
zca019c1b554048d77242bfa8516f97335cd0c19a48d60b6dcaa4a4d0e817d199eefe72f422c06d
zc70981e111ac770a6931da34aa72e55325d5ff61c6ccbbb372c7b0aeb256c03d95a9203e8f3942
z232e8209665d08f4f665d1698e39545539a1623a72242d7c16f133a7bc3e43e5e81001dca6ff98
zf62b25d09cae058779cc8e1989ac969a821c343286e32ed4be385e097b34f5f237b459ef21d802
zcf41a1f4f5f1fe41dfabe2b6f8b6e8133fe9af1563813a519eb33fe6d2bbe680be851221ea641d
zb4aa41e64b7febd22b7f3c1ae51ac3b81cf801a6ed7d79f3e607b608a4c1dfbefe16e1e80c24d5
z7c8f739a35046e32b647d1aa1e00a9ad894f49ea1fc308edd234870323610f0669eec01838f754
z1681a4aa5588b3793908ab2bcbf0eab1007d7c72c849da641e56638bed84e53e878d65cb6c0270
zc0090224bd8458d658c7d3c0161ec3b806565fdad62331f77e15a0eaf0e2ce798492d636c1c89a
z87cbd77f5c743f8c957419641ccece17530c2814b3bb97ea35a15cec090ca2de0acf4ba89cea7c
zfa3199180c2ce9f91b0342ffd0354a0a8812f8597d8979ffdd49a16dde58619de28b7ce4fab581
zd3ef66a7f79241ff6964c8adb14ebb83138d61a6693706701ad776de5c349b6dff2df687cf7477
z5faba1d0e69fed7d3d4fa14f0efd12fb36b73cb58fb3d5523a88135af9622736732f0c12a97179
z437394856d1860524619b1879e26d2719bcfb1ca21192c48223690eec4a5631b3b4edf8bfc4997
zb4c7926c809abdbb0951d14a41ee15e36a2136acc7b192376f585baea6bb52e6b6f4a52b27ca0e
zf39eba3181f6cb12789b1153ede59aef2691097209256c3d80796430422f9af7477b001460a36f
z82e8463cd72881d1e4dd2c72241d45fa4be603a4e2cbcb7ba4355cba536efda040264aab961fc7
z15832cc67bbfdbf601b68a547f6103eb691aef93bcc59833e699dd3acd7962ecc6182b477fd8c5
z7a1f1d1a728f3bbc669d5841c56f7ca20f1e22caafea1c7db2733665390225915d61a2a2afa3ce
zc99f4a4543d7714db17c43debd1ebdedb13de39960c27eb26332677124620b419fb7eb5c8ac50b
zc9079317155859d9a624c77aee0eb33e09d59499aa62d53f5a6c6ff4b0593b41500f069bda1cbd
z102372f9c4ed39adffcbc3cf83b5c0653ababcf85fa07a0fb6cdec4a91fcf232aa1aacf4cf6f35
z7d73021a08ce5ca0e6860760fec747314f682165a4c9cceaf8f61008f86fa8af83a54abf4b4000
zd6d75a45bd5a8db1063eee5d1b5eeb5799bd6a667a500168480a27288dd7f96fc4de3ca3ed0cd2
zf0e91e517a477c6aabb3739abf19a288b656182803c76ba14241b5c9633efc40813568fa80a473
z4f460b9277b0c91476ca3134d742eb751732bfc4530d8d2c67913a4da6898e3fd763335b0f5605
z4ea180015e9e469b36042a3317149cb21977fb3d6664cee21e6c8c3eebee6b8d5e6ab2460facf3
za93eac17f5981fd63c01c51777da9fcdb937fc51f98197954f0dfa72f40d6da67fad8adc0a0be1
zcad538da23c52b2f470801e9b35ba76ae18aef17b742a458bcfe263e973469fc7334b6794f7086
z01f2992f04679555d2605e86010cae0cff2716125a6aacfe07067964750a12799348407bf162c8
z380b29c67e0f34e8959ce5ae75c509ca816ec451aa44401de7e28b20dde7d250ca4e5c8a2075de
z9c499dd4bc50513d9d2c8b4905ca9f7857ca6ea331e144e6d623c4c066c617d3ac6a4295bb1e38
z8d3a518938bd7031a8e54381e0999954af8df3a509c669ab83232b11075cbb65140267b629d94d
za89600a581f722feaa4fd7b753cbb5ed22be8294e50ea6e8d136a5c1b49f879f371c3bc577fb32
z20a1c15ffdeb3d431e9cd5b956f650b14a6be1797f697ea0e2071f91be7df7df3db4808331f9c3
zd4e540058ccf1d0705bcc673375eb06b3daf0d7e2a22dbc41ca279298fd016595e751c69bd9749
z567ec04f813b36a04c2a9ad5168d164fce4e5adae48aa5402e73f0654d759cd3f6f77e10984160
z1f5b839eb2fc176988388099671dd62710aa7f0c67c81feb44af687492613b1b5e8a93a9f5bb25
zcc98c5578af2bb622cf5fbabff8a49e4994009b80f2ef286e487bb3c40063477a455894622527a
z5268c66cae6f0547236a057c22d06696a293523937781b7d5276338c7404b2b401a2b011ab3f6e
zf1a04e469f32c3b74d16f975a923425c20aa03ffe3e9dfa1a229c1d65812cc9fd027133119cfe0
zae123d5d5f08234cbf53815ce197663837ecf8a7198b415fb233992861c5511d080200e419ebf0
z65857e97907ea2ef0e80be54ee5acc83e3c78fd654b66a640751eb8001f1ea61a1c5d6f93e3c16
z748f97a29843fdb90fdbe47fead72a3007058140ee6f997f5255284cb91f81420a6d6fc5135048
zcb7222560372d0f276225f9a0cf37d8461bb5971f36be84df92d3d59e51f1d5ea93a52c2cfa886
ze0aa69199efbef667dda73e24ec620f32cf7cf6c016bdc2b0a992c734a5016755d203e743610d0
z3b5948f7176c78595d5086f5a1df11cae5b91e948ecd590d11ee1e9c19445576e1c81286c4ff12
z75c7b7c5edbc6c1f5ac020b1ba14d6312ad50fea4dc3b146add6ec9602be01467e390484b6a03e
z65223091beeb4c8308b3aad1e0af7ca8f57cd16ee7a91e9dd30d764f2066d582e7747f2c1d9475
z9f091a1ed56b7db712ee9673406c28d45e9613aee8ca7c1d9616015fdb640d843790d1d173d2bb
z9f3807d1460e5de839c2ec95bd9d55879aa5442de3feabf3eab5d643649b7a664e79727b09034e
z3daab4e11ad9e8cd104aeac4dfe59a27bb0970fb42e5c8d9d87bdf4eadaaa1031c52f656c6ee86
z21178d58678db53f9206fa0be25432d2aabf23fb4a0c1c2f0ff966ecc61619f9f2e67507fdecda
zbe14a1e26d945bf6ee240b7e7f0fe3dc56a2290a8d9db779bdf0999b98edb6979496fc8316ba74
z5b54f13bfaf9dcd80d831c9e8226ecf3e558d387a583a5720c5e9093f9fb83e76c0ffec50327ec
zdcea289e8a42a51990f13aac08a2605953aa05b61863472da87591e046ab0273ee0f10bdb8640e
zd53e259b816db519747bec9d16a1ccb6108595b1d407177de430b1984d9766f1f7da7360cbebb2
z079278a4f70d8b0b698cc438e5dcb05ca3da57e0cd63bf269eea67c5e399af77bb1f3fc40d8f99
z08081a1b14672a999de60ca19f1e0169db545756f089a405e5897a12cd43b88926fc9cc5906562
z6406a50138fd7d3ccd012642f9aec50fc2e99f155ad1050c24aa56bf9ecdbfa672ae4c4bb202e7
z99d94028d657440de408bb580d3d9c087fb392d26aa84db3333371207bfd563b880ce893957bb5
zb8434e58a7a2f6a8ff46bafe39cd571bda12f3379d25dc81cacdcc4cf773f5b538db517de33eb5
zdbe47bf2c8345e0feb7094e97085e375a0ab2923fc30fdda291dd435c87b7fa31516e8d9a6ef8d
z597f309cbfd3528acdc9dd78c121fbd55cf1a7fc7e8fcd85c6cb21ebbdced784af1d3069179c79
z752b04de93347ba1838c23033742edb989844aa5a679b73cc2b9cc6e058e68f5be2e7ce6da196f
zaa2c47612ded7e5f1bdfde2b76e08c6de243c2f669f78a3005e2fe9ba4d2d126f7eb438e5f87de
z8bb0423b7ee780ab1e212b72150b75d124f2e83897dd34d99da1c8c04c8b16c20adf615e8597d2
z05eb52d46b579cf0f22499b4ed91f73a655019e4153cefafdded04f95fd63d6e924b02a57bceb7
zd622aa51ef0f70c35476816cf76ce2a4159e76ce1a0f752a79ba0c0a11d098af012d4aeea0cb64
za98ff79aa35ba0ea48cd9e701f555f96ec18dfa70869a7d19472320051455f823907c9dc26542d
z1225b209bde104c279984cdd3c4be20c4c5ef4467d984965a09f786c000d4e0bedfe70a30dd580
zf7979a699f114140b2091836fca8043b2f16b839272f2d4bc0e3eddee3c7c02839830fd53cce2b
z44fc18d981f4764f64b66b60295873539a0914821fa67bb7b1f55e98e54b1813acf7c63c77968c
z86ad9a4ce81c89c7fe98be525a3d5d32f396dea0b5e022e22d5dccd85a37003e3e8782fc1c4f0a
ze6ce0d5211c69bf49943d785be45c60b7da2d2c949e8b3fd91c8f051cc1832fd605964198f58b0
z4ba39bb0eb43153002c9093443482c806e802725681259a6878869716f604fee287f5d4a0f6fed
z58ab837caba457d1cd3eed430a4af3c94c0c6cd71a7eefdb0d8fccd5d3e1b3ff399813fe9f48f8
z753d093ab4f725598ca06d116fe9ecee122ea5136f6fc5ab21a46f67ac5e54633288fc44e6a484
zaf6ca24a1208dce8584a4e12e5aa55e3a290a7fad99a5be75b1fe75ceb12af5022ead5751844c9
z7dc4c604cf41a4f6f3b1f4ea241f12a3b752149456c4bd57308a172d6ce1aa090ee348eaefbc7a
z19f98f53ea244ca6f1edfe79e3a4440289e724618dfa4cd82cea9b8ef9c197b0de9e53b5879580
z8a26fb22adaae3a460e49450ae7f961a2ed115e80356da320969f3c4f4a0ff6d64dc6dbd33f48c
z7ce7d113cf4834331ab30626eb0d1a53474872419875a2516b8107e35d68980cd084b464e99e9c
z97ee5a4bcc41eec4c72bf521b18d7150db81b54685c78742b5a97fd3058157fb996180d60b8026
z8bf93e6c403bf81cb4743f9d51825ec82cf2159c9b08b2042197864494c28d7469196d0fc24381
za6d1e3a0c1d8a738a9b53ed7de924b581b585952911ac9adb7b6072f85d307a8f61aa9cdab2b1d
zc1af212c9ee072028db0a9da64502c589ef7b66e75c717ca8628371c24bc2722ee3f47ec24d70e
zf52097a87c0469544bda9f949434247662d48f526ab3f6752b226635b154c8013fa124b8f673d9
z6ca6e0bcd410dd9cd709349bbcd36a405813a48eaf644fb3ae0514057db6065e4a5f56ceab332e
z755542c2c4e4754acbae8860fe5c776626f736aa2c3fa2ddc9de4d55e49958733ace9996a95d8a
zd23c14d109858d7ee0698016c87cd567efab309dc7d889249432132b2d43f683ef26ea713dfbb0
zc236086ec0f37b0481aae4825c16d0654edc33634e0b9b1aad0eff4e13bc9e81841aa707f69b9b
zbe1ee31e6a85000d24d274aa02b2aa7a4ffb02d36e47fcf8a18efc522847ad9491780cd11cc5a7
z7a2ea1c95333c0261fe68688efa25ea7f7b53ebdcde9609693e277b2f2c0f3dfb35cae8166efdb
z513a604c68557e5b5c97439b9f67cc0452f8e2d31c402c5e1887e64ca6ea81b19e038b29905c66
zf1ac86736988b8eaff11e95ffe5d646bf2e3a4fa6fec96af0ce7bad36999d2c4a7d3b49c41023f
z06aea41fd4bc6266ddf980c7b4a68bef7a56365d8f3fd10b90de98bb3d1ca191b3dc786ad77dec
zf5bb247ad62063235d2d04491b1f0f8a59f30a51f977369c03596107520186b8a6c79da51db6c9
z16ba19efe61a8162428741f9794db529adad5b4f4e277ac6ac449dc231943cc533e7ff9843a8c2
z63b8ce9f51c9fa2c6a514a64006d45f0f237ffefb4ad71d65174a50bef1a63bea981f56b635d43
zc0082bc949fe340766c9a7336b4c02cad49a8949575d994d943cf73da1e6d2281b59b8fc1f7039
z0d3b27bc43cbd163bcf21bb1e7474cc0175c133d93c4b90883ba50d3066ee528604198fc5fc48b
z8c13a5eb44dcdf1422c98bc49fb3c44536a24dcf297a1365d5157c35c0926ca6d4bef3d8c60a84
z7f475ac12a42482851a68dca164f061a59df9e1e9feb88bd285bcbbefa2e54375fe505a0907942
z1d670909ecd86bc0f69b15af7b105fb300e26cd2261fc046b89e32521a5f80f18af2325d57ce6b
za9c10d41c33620fda19b21af80d6c8c9bd40ff936631963cae89fa1554d476aa1d230eef459273
zcd3b38f8d80b21c5897bf1af3eaa1d604756b6fcf8059af12f18972d60d95827101460de2160a4
z3154a2a38a0fc99030f3d60f0a9a1a06b632d4d8b54cdc9bf9626e4b90a14932ce642a8ef2e4e3
zfe561d701fe410b02e0505a3d2a5997015658d65a34c561b305e9ad809d1e1ff42efc259b19b2d
z0958e5f45699dc549ff1ec6caf5b1ce24d0fa32dc63fe31d629fd22dbbe72f5dd401ad14895157
z9b846f723a4cffb862330cabd8b1e9994c7237b6f0e00316a0dc138a7f1ec98e9acddb72ff0c4d
z1062b8975cf166338bfa7cfeacbf62e6af882716b658e85bb95a2f99db63827e3fe5a54ea4e10a
zf299dc5f886ca8c4daee5d138fa3a0e813b09ae5219bd73f966e13d02352dfc46a92e1e8b8d830
z5be2a2c87e3b146881eb8087c6377a1b6544d9fcb4074556c558a932974f839d95180495503835
za9527ab44e07cf7276b53b2998ba6caff465bf434f258da92a6280893b0d1616b495880227b417
zac8cd50aaf6873177bf70833b500e0830bb58e8fceb941aef382603107e81165f406102e
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_xproduct_value_coverage_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
