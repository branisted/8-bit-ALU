`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d5983e9214a24203e048672cc6c97760cbdd6befff
z0c3188747b2287b574e4000415a25480b650cbf0cea357f97937ceddf19bcacddcd1bbf128c8ea
z738e62a93410d596b8c70ffb9ac4afda12045af64e4d311fa389f508ca6f54a8a062cd975123e6
z13d4ae6db2843d659598bde04b6754142103b0f4f04706d4df18341ba54524d593a313e7b58280
z7f77e51b674fe8947b5076fe6ffa9de1fac226148c24e120ab4a53e5c036c95752c01bb0a168c3
zdc6e5ebe9626aba68fb555d959b862589e1d9f76d5de9aae3128875401f06f70b4f32aaec4fe71
ze36a1674620113fef2deea020d5906c341da308ad7c71e4b49434e350dc5515cc84905f023feb7
ze47da43885b89d19576f53200fb7b3baaf55cb82da729dc5cd328d0a68e1d902df9f8d3b68fb1d
zea87461957cb1b0ff2b2f84621695737c81870dc778def3a18d869cd2301dde48c559e06f9874f
zad7d851309d8703696fb65005dcc38e13dcc7739ee14d855353c8201893e136d21a4d73a22efa9
z655f16e39528aebdb806be74818ed19f459d07c3a4ca5efaf8a0a5efb81825bea4ba4620345ac1
z46a614c4f0f85ae5e50c65949da581d95ebc3e3a843aef0907b69f830faf036e0bc542fa7c1ede
zf3362c1013037d3a00b064768fdd54a76ff53f9b1cf06801598349c2ee451503506daa9690ca42
z2b318b5bc7d98032f2832b101b45f154fcf4f091db5f390450b4c7e29b9c712abb03b794ee1b2f
zf4a6f476f4abf79f254357f8fbdff9cfa6e679f80cfbc9d902e07256f8e14e8edb46930e202e2e
za356fac0615a6a5692153741561e6e2c09934c7490a76eb09c2172f6029583b97b6526fbf47d04
zd6f32323f05d9d580a9c309a87c2a6f6bf43b82dfcfd9a88d12ead2313512fb7a06e3147284d43
zdde4236add2ae16d243f68dfe7e3f31948a7893532cc9be93960ba034cadfd7a8b988db1894c2e
za75a7b2c090baf33b086645fed92d78490710f2bfe200c4dc3e969b4f35fe52d37d6cbeb9bbd03
z2037dec869d936247ef3e0ee7c8e310495d84971ad0e909fae7de4b56a60e76e1fd3e9dd0974e1
z022e9761dd0f030e609009d30399fd948cf84a822710376d42112f893974cec9c2ca1c6e8779d3
z9bb9884f31bf94ad0bfcce215a65f0703446c521ae8069f084ed59d3e675a54d68d11fff7c3722
za0dc5452ac1a7608a10594d651f4c2d43dc607ca74f38bb0f854e734cdb7cea01d0a43f6be3bae
ze477ef23349e7e651b2dee9a4058e5581fa7800b4a1498a99c2c142d656d26916b88f4f7cc6ce6
zf4552d7f666a5b3baf52c0fb30a82f8ff74f11290888cc526dcef61797fd9fdd218a790ce10439
z233b0dcfd76c8a9b96b14523c0a85bcae0f25d03d9be363b60b8eb1c2659622cbd9c0871d81576
z85077741f3142f55e1e477be63680ea6ad3d7dc4f383e210e373a0484ab3f0e2a0efdb31c1d2fa
z423ad0409c1d7b2a1ae53ed91b46894ee0e4346a2c3b11bd2022fc0f3022078bf7c9e425ffc92d
z68fec6c6d34c33236ec3d88876d04384fd209b169856e4135c9e67ac90e63d6b4075fcd82562b3
zf9b00ee2f57ebadf3c85d0b26ccb27d5f27eb177bc8bb1f60b44409bc8680ad11f96c615ff51e0
zd11de4b077c343043161e1eb37bfdf6d590a8ea26f4585a5824f2d978b13273fa34c26a1f8c335
zac2027cf08d8277dc200c7a63507d9926894705c7402549df9d527a0f4a22aed49497b3b5a5c95
z0abee2d2f47c1b9e55dc56cde207ed19e3cc9fa90d67c1ebcd43cda01f5e77370ef290fd2a899a
zea23af851a8d895b9bc78b2349448810b52e738d96bb22b8f74a4b3ac9052d25bbc82dd7cd7bbf
zac617c55fb836f92eaa67970bda8a459704daf763d170543b47e726b8ca8f2a794dc7bad97b475
z2ae9fcd4f432fdce16864d1bc9e455c175dd0e22044459f846df305132a2c3a9cd767677325a4d
zb66c7f52d3238839a2c3af4a29570ba81974ecdfbc867221d4c5a0d91b090d280909faa7a103f1
z70d58560560277087023828a9ebf43b82fa75b3608ce05a735a9b6969c26f0bde79feb9a2a406c
z3bc230a783a7b009f8ff58b389df8100a23005e0d0e30da567e26958498c50c921c4769b291e56
zf47f4984ffd9c47ccb72a5313f997678f30e48516f3455e371c2f34a8bdf4b4aca9bf5b13da6b4
z21314efd639d1c7b2cf8289a47f661be5a5cb46a912edbc7497ad423ddc7dabda95d914d39109c
z275d46b08f8ecc6c9e2ea187f44a1d9357a993031c0b641cbe604b7f8667766c34955d62534d52
ze1e5021d9b77d04526cdce65268ef5084873283927e8fe5f1ae522d3c8b97e33d2183d2019e94c
z65242ed89d6eb0bbc74af6e6c1b23abdea0b086b39e69bd2d1aaea96627c3064174305b8aab59d
z0feadaeb5918747c283b7f1cba298002b8a6ad082fed037c77682db56b8722d74d03c660862af7
zf26f9fed131c0b54b746bf17dffcf35e2e7ec1738eae2aeed68d47cbe2a04d7808a95009f5a2e2
z2fcfbd3c3146a95afc93a5b37df2fc07f87b1d5d0ab41222aa2cbdaf3c5311fa2d3fcffe492b5b
za2159b97547c135d414afdd561d14233a9026c55d159cf3f771bdaf18d0defde332ab732f2ec67
z032b563c636049325eeb435c26e7664ea6889a59e7388a54f37e0a5d18f9792a6ae294e89f3218
z31b0d5aa5a7153910f7f3dbba9e076bfce9ded30001340d83b04b714d298771ae3a24316d25bc4
z1806ed51d9cd3f3bdc137006946b896602eea442ca415276952c5adb055eb286e972b784034eec
z29a89296e08cff9351261bdcffda303f72c20940976d9d014057e04f313174f1dabeb010859191
z37af22e24c6f834bdb8e7c6695000d2bc3a679b3685d19c0bc77d946c1720789918df8fb83378a
zc64feb39adbf54773251a9f7a07b757bb123ea42d71e5aa92190ecaec870d441e21656d0d9cd9b
z0f91b308d3ac80356dcf9b3498681c2723b3f15bf3b58f61b041bd13a066146527d49b8d9bea36
z550ae197c7b6dba4278cb1e6255a7cad24669aa440885fa97fe0a4d93b3759658039a08435f16e
z74340ee15ed0bcef7a69fb085e0bd353067af33432a91042d2458d2e20789f08fac4e985f44628
z490245095b46758c81ae63756a0f04a2e877d43bfe057973f37a5e0445ca950190a85c89f599a2
z2a9942b8ca432f26cf2d1ae99bf85f67bf61235fdcaf9329f5aebf36b5c5582546c6a126bdf90b
z0f892399feb2b642c079aaf852ac86f8c8fe20530413bba5e53ef9ea9488ea4d7730a5472580c6
z9239586c115f489cb2d3174a18e5a2d10a761f341f66d27dd577c0970c70291e0c9b979bf52535
zde704c692bf307d97c245a8b5422fbd8363301c968325e47601407904f1dc454e686b024087050
z109fcb1e8bdb27430989ca35b368c49d33558e4641665dc21a4e88409f03e1b5b7d8659a548916
z4d42989c6be23949d8b1d275557762f83d3f464f733dddb785f62d1a4284a4b7b6afbb662cc554
zee98cd5506b2007af18e07acdcfdec3f3ce5a23997081c89f501b7dbb5a030d2e328e1b12ce631
za4f2384e032bee0bd913c2e3c77428ecc5bd283c26066d17852dfc23b80a4b6857a58c194689c4
zada5daeb335ed3f29d20bf0a13df7200290a2e663ee7c7c8948be2a82c15e0b834ef28ecf1cd32
z14e02ef9c440a1b59c8c0fc7f96f953df3ca50301199b62b90de80c8186fa6845e6fb9a13cb381
zb56b2ae127c10c810d59fb903bbd2638b063eed324048e6a0fb7ccdf53f1127c9970918863e443
z961c68c681b997cfbb76b5431a397295a0aca79f048f8548cfbd840762db3124ef922502be7f8c
za89d59b090743d0bd8820b9a21baf69a6fe6471690631815094d4bc92bc0e5152b8a976fe34850
z57c8919b4f620792c7458fc7787fa7b41a5126474411e874b446840042ed159c4eecde72c850a4
zabd442ea5c94a62219bc7669742400b0e7d5e507b8e693ef24424d17ced423ae660e7a632f0251
zd9be3216c717ffcddb30408bb3fe19ca971f21f8c9fed444fd3a05d94dfc1f9b1658b5455ac6c4
za063d7c82d437a84f5b1ca857bd7b969e434faca45540f4177c4334d827b1632f3ec0eada60beb
zcdbecc8899975c602f1722a55f34fc76b26882e529e82bba14c44de1e80d17e0b27d02c4b6a51d
z030786aaff5b95c52183b2a2cb6b0735578e278f46dfbd9aa3744d0a5bef7fe339fd18685d2153
z3d8bbde826c5c4eed9500a2fe192240d22e01533de18e4040a123470315aa866a53b7bb9d881e0
zc440e91706105497b5839603223c3a8704f8d7fc476ee5a07ed4ccd7e7ef025432f9b1dd2e1702
zdf78264b3302df088c4707475dc38ec45d4b5d833604bd3777451eacf45a0eaf673701c65b1f8d
zd281ac2ea0834a8c0d355bd0053397d0ab904342ccbbfbe71486eb8949dc8cbdb7a81ffa30fbbe
zc2dfd87e61cb1a58f9cf583bb8dc2d42981db57091a8e75a52196ead61046da74116025a874139
za9b3bd91be5d947675a5ce8c4f43ec0dcab25b802292f30cb02854150fd3e8aa86031bb433c2c5
ze3ea2e8cb90366742642d136990a425100571fc1fb5ca14e357f50a6fc48e46fb49bba16f105b5
z8294e30a997779b46895357423a66fdadc5b3fd19200633c0addb39c453f9e00622a150b4589f6
z8d3f556a9e84a5bbd946028c631d399fe150c2f7bf1fcbcd083faa4b3a03576a33147f2241fbde
zc5e7a7f57dbf3f88fc8a2b816b1575fc0cca66e05815e573293f5b28034c8cfd18a51dfc1c02d8
ze67424b4a9994e126a5c0a3fd77628fc386d8bdeb2b3150ef092d76910e740ba3e0c2bfefee63f
z5053cd3fcecc7dc1274b66dbbcbc3a84409c46dac5c1f22a2244a2de404720439b1c22b459cf99
z82aa00203c92ad0de10bd5dfa48ca311f037606d37369885a55c214b7af5e51224542e3694b956
z40cfdadb5710bf32454512ea4700a63bf5e5e9dabacb219250110a2cac7b4f5ba92a0704acd8d2
zdc90ba1c367cf6e3dad02c666a6d6e94aa326f9171f728739255a2ab6a9f6658e869f772557089
z36c77f922f3aeeae6be6fe4fccc0c83f700c8aae03d6682741c8076fb347abed4f17e7e3ecc908
zf72d54f7882cfdcf0badd9d246fbe2b2f6cb5c07e7a02af1e0e07a2b6b12f24be821cdd5d15fdc
z57db230a28e4fcb2ee3aa945ff0ee65c96735c9de7e78763136c484d555e2e8ea17ffd4105a65c
z1c300871d0cd72e8c9d16d8b39321cfbe5865394711c675f359221a6912790a64b36cc640fa9e7
z300bfb3067457f471670e2121fac9901c9e190f60dbc1557bbf93ec1167a324eaa856c525c9601
z5bfd1d95e83da66b091f598782f2272b03f0ba47c3e7f7643e31fdfe6281d7125f4dae747b140c
z4d7b739cd8374e9617fca211e131937944394516e75ee881af8b4ae1d912d18cf8def2ceee80e0
z27b0888777f666a13523cdd70ae006ca6d6de580f3d18f97315572ce299ceafd6f15ea598579b7
zcdbbb5fa86232fa405548de6b223e0b94963ceee30b147b25f15ab94ac4244820a8096cb966ea9
z3c543984bb4c9fd4efbfdc1ff88e0102acf9a5447fa3a3eb46a8d160c75019100590119d8e6d32
z568b8b547a10461674082710d4622ec0e377f4bfd72422cb188c03016bb0f657e03f1c2c47d0b4
zcfab8ee88bda65b8540fb74ad1dfe7bedf85e80cfe9aeed1b5a3b678e8c7ab3aad79aa81d0e53c
z1a997ddf2cc96fc23296d354a8239b0c73b5470d3842337226dba5c2f3338d9986e4a0e0e2dc96
z6ee4858ed93ab556ce8a67821747230e4ed862c70c9aae3424023cba78740385b8f86a18720973
zd60f811ab986fd7e355d128e859f54fcb0c90b96e2b0fadc600d3633d60e02a5a9dbd12fd8af89
z51e232609b5be2f8576bde9c886779c20b89f37d3a6b2c9452ef77b02f9c44b2dd2dbab6c5367d
z3597c69f6363850e4f4b7230d957d295b2af203028b1e928d033a1ddde37c688fc9434fd006d42
zb243e6003967ab5f11fa2f78fe45a8c627c6e638870469dba5fee0d83128e7f76dc957455a09c0
zff693b8411b8444fa0fa031c7cbf50a14e17a11e1d2dd13c801480108455f7261b2f4a2cd9d770
z623d8bd870866fe23e9ba799a0460ee644424b5094ca20320792060243cd3abe4ee9374dc3fccd
ze421cdf14e47b0deb761d538e72c98975bd50aa5d392745a90134908d0a106d9aa1bfd4c4b6522
z84f2fc76c114235711bb1264990c00e61802f9b83d230b2d41720855716596023b5cfce2983689
z72d4961d0b2254d5bbc39bd64d8106b5a3019182cdbb4e12325c2773ef6a4e474b6467e2d2141a
z4b461e56c0c66c3b29997b6de0b05ef8cbc06dacc9e43548c844f4948888a020908f1dbc9e912b
z7460dc6fd0a453fe200b23510400e897042e9f32a0543a0af1177ce9af2c4535a1a48368751ff7
zababa7ddef458a34be493d7d43573f94ba3062324e9d7d88d2d1655833ecf39189c8dc79d55ac6
z408c9bf50d8197aac1ec007d60b4fd8a6092b95016d3e03ebda3285ce2fe8e0ce569e30b1c7a3c
zf7e84c66d8aad5dcd1d6c63dd4d5f1785fc435d50c7fa18aeef5ce3bbc40204d639deed60b6363
z38997c24513ded6b2831e708aee7786407a14425327aa9515b55420c809c151b5a7dd7fdbfa24a
z31a8ada4e13858c8082f3cecf5e2d34b4eaaa3df69016ba25cd0bbdf6d05520a5a7e1c372053be
zc2fe557eaa7be327a96c16ab675604c441c947fe2218212d71222a9601e698f483195ec4157b8d
z4b6428ae1dc2da04fd719ed73305be33bcf78d19c58991330a64ab6b968d440a82b4f24f5f891b
zc40945c97fb3b55d36f1a94bd0d6d1f9f5128eb40a0a73d930b2126f22585025b980a3c393989a
zd3b26b8cc1c23e634e653a212d8b0218e279b27247cdfcdfed96da6c098748aaf8ca9b4c99d56f
zff611c1c2fd9e78c2a060212dc3ae53276e27833ecfeeaa859b3998784f4fa8af202624bc4438b
zefedb5d375edf916dadeb3c500abc186f1f4c29e590e731bea5546814d65d7ac990f86228d5379
ze2d6858d2f2028c5f063fe083ec7d71c7844a5c4d84ee4871b660ec7081c0820357b2337f6d1ed
zc4249e55f9a057a815af274ba01ee85ca7b80f8b1edd1f610897034381254d180798a5375e9c62
z7bbb5b85844e309967ac4228eac1378d74b410e3cb2abfabf1f650c216859a58e2ff376cb78be9
z8f3ac631633177efbd551abd3d8271b820e764eb6cc73db6be568fc709c7c63ea0805c43a701a9
zc78425f2fea5edafd6f8492d248c50d1567f8856a3f600101feee5de7de7ea12354d255c1aa79c
z0fa3c2f909126165ad2f0d1916d28cceae6853a2df9349c3b6e9f35e4cbbf284e58cde6d91cc41
zece7769e6588357668b85bb2671952210a90a927c4e1b4a8a46c9bee9f5c5dd596b49a9ac0682c
z18f17a761d8f9b8788c54dc2ddc86cc89efc555d32214b74d9b3a569f2466bc5c32c3f3ce8ec44
zd820067583fe3d11beb3b54886dd8f2f6cc7680ec81d9a3b501a70dda438145329cbd24b07dfba
z1b2a7f1210c02e300330b4a203e82abe8c45ef1c902885f6efe4fd46696086eb5e8714f0a6525d
z38e617b967c62b7a0b4c7b2fd1d09b9d8735cda92f80d32ea6b4fb459806a2f7a83d6fe489523b
z34330cd7727976a5b8cacdd0e188d149bd7b57b51d83537a5b8f314b04f757f317672e4c91d996
z0a01039962a072c5ca531f621c66ca499b0331ed8a364e2000548962d4f4af842ccb367694bb61
zdca059b20e19142e03c6cf9eae803c07d7181981e8f5e3f4ad71199c6ce1326e17f94247f4397e
zebce8728169db70c5d634a5a81453157a9d443beb219a1d52aeed2b9b833bef7c6a3929fddb6dd
z578df94af0cc4d988f4e0b4c29b64e351a85ef173fe96a12881b0dddad24ef1a176e626b6672a9
z3db2809f6fb2b55ace82173aef163f9472556b226114ddf61775aee0e1dd5e31114bfd577fcf12
z29ab44b3b627fcfdc38eba6fda5b68ee75022bfdeac4c476ab5114bb70ad769434d2d217db7d2c
z12477d2904ae7ccbd3db7b1e075336c04289c5a7ad9305c61480ba0320205a8e801eca8553b63e
z696416d37de379d12d6481822675ed3e11b261e1e341095779d211674f01484942bb978f9072ea
z255ab52b1bdb6aef4350bb2b818912c5501c4ecbc0ae3eadf15319fe6af226b33b475619932cf0
zff701200c59c00c6aebcc7c2ac0953b33b0fe3143202c1fba7a6b3a6d202e1ef4fa8557985388d
z955f384ed1995ed430d63c9e2e0c6a1f58b1d53aa0d4f37a475e1ac1d6d6b635ee519684a74d5a
z06a77cc505e1833d218131d0b4e5214158c59b7cb0013c5a14924e1e6f780739fbc0d3ff4075b8
z63cca7eff6cc26f95920576be180f3919ccd401009f5fa8fb597014d0df7950984115c1460af2d
z11764f0ec178a599cc0c263e621451a0a84d2ca7e8d02d4924452a97a44d68e766f47956ba8c55
z68c77574c216b43e29622e500f38f788b962f3ce79e4aa34bb036b1fb31788e598434a779289d1
zd906190a52f890f4ba6c159115d8095b6ace1ecbeee883c6c624b4f7c3216a570b38f90f57d6e8
zb69b19d4b85511e2241ed7133b4b25b8ed9c5d6987eace3f80b807aa09a6565f108a88f10eb4ea
zec2242fb0614f6944e24efaf66c4a1235cda7b998069b94ed59fe490b1634119d472587a1e6321
zd3f458aff20432333a2b01f48673ce1da4eaa8595f0db43fbf9f85361dc92ffee016f0ea484722
z0a29a1632695e0b9a23958599213b81f4babe9601a1bd98670b7bb64989a9b37c3dc31ed7afbf7
z3282685506d220f7821de9c65e0f703536d8e07253cb45d3895b9eb649707630b22e21fd18e238
zf5bfdc0912730cc81b43b50e07950624b82278fd849c5efb9b8b41e88248e5620419414aa22590
zb0f0f1e5e78704f16bcc3dd0885ce87145b9cced83ffb25465527cba1c4520a304cf42432f3c23
z98e74b504f1ed9cb104f67d8fb536a40fc11ffd92e73d51e6907f21ea5741d30c35af494d6a0bb
zf67d3a1e88d22e545eac6f9680bdebfc7a467b300f137e7ef6c71e5bb7e40799a354f19f44e78d
z3fefdb51e1c39550771fb3cc78e9f9d9e4f6e9273dce38481fdf1a39873b9cd75ca31ae7678510
z1bd26766ac16b7bc94704a356f7f6520830273d5fdc372fb357b80dba8a7e5fc6f734e55f98424
zae5d341d2f77ac777a762006cec46335097658184349be18038b9a662019f41827103ffc011306
za0ee6423f01833af937f7fce8fd90614ec0c7bc127bfeb9c3513308ed7f9590ced74beefd650ff
ze7549c50a0df242f7fd508004df41bf6413cb096d770fa823b49c30166b121c4573fbdb33460f5
zc036a55096a5931506cbfa527d0bac6d195dfa9d1c0d9ab113a94e1b452812bcfa2486b93941c3
z1a51fdb354f824af51347f738b70994234e0776bd0de5177c4ddddf5762021c6e15e2997a100a4
ze3eeab6a912fcc63f03fbd394e65c0f98ea4bac0de1da2c6eb818261cdcb017b23d32a685d20c7
zaff757276ca09bc1c917322a4ce7fb21544b4299c2fc6d3150b4e3adb1a1b4749675f96916f595
zf3136de08ba87dd0f56ddf5cc2e188de9b1e62bcbc1b1b6808a6a3a30a29b4830825b60e5ff637
z74fac278da48269f373d1fbfa11bdcb85fbb87aee03c5104e8d0240855f5eeaa346e0de6e9a36f
zeb4e1199f2b23f9815868f27f623a5ebfbe137150add74853b14deed46821a012310637aa4365e
z1fb22fc2f0de5ff45ab141d1d13ca581c67de51adf2f9e09f8a5c9e55e64b077c1bee8968eb891
ze8ecce82f8f5153d53c43a759e4b527c4c413a947b746ff90042811869bc4ce0dd352a7713e8cd
zb2e4750c4dfac76e7ebd2c54069bbaa3bee841c4e71407483ad288216cf10e4661da4f337dc5e7
z909efb4cfefec7b1ffd8de842dbfc20d203f60889b708daaf786ff4605eead3a1e917df5db5ae9
z5134a117ccf9fa9107a2c26d9b45af815c01841447644054d97ce8463047c56ba8e0ef93af67f1
z136c0459df869e724ff8ff5826fa483c5490722b987abd9650605f9cc247299ee99bfd3828b305
z13660158c6e5cd58f85df02d827a21f020ab33fb16ebbe6dbb4431290da87a78c88d
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_driven_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
