`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff98478405fcd4d89273452c559f93e5926bfbc31a6dc7d3
z54b24d4be133c2e8791d1a3493ef5eec5ddc7946adae891a373c8b420742b6a218758e6fdae1c9
zfcc0f88130ea479e101a2f6789b158b79ffa3cab79e0623a00ea43af63c2b68b90c14ebed7aec1
zc141effff67906c15a760ce479019bfe64b8cb937169d03ec80a9e71b99d78d574a4424e625843
z9de21978ba8ff3694ca7b3319c0472f99a45bf243b066efd00a192c37c2a6fe73fab2d14bef08c
zb5888c12731aee1846c1ccdc7971c30821b279ab3db9b8e5525e4d229fdd4a0442d7623fc79030
z19de04418662bbdf8d3e9ea66256ba565830d4424b73bcf9e509e7dc8ccc8bdb53635a6daed91f
zfb1dc689601209eba7e652b3bb9e4af4d46b3153f6c116e96f73e2a246ac17d9cb8ac3374f25ce
zf7726d539f16f0343cae77f6392f8a8d58f03aabe29d2b7cc96abbf9e990ac57177c41ba322a6c
z1598ac93372b89f370f6aff053adbf4d8d389b0cd70c737cb8d9163a161d876a217b6f97cadbcd
z739b1ba86448c6a72f06d0bdfe802ce80c023d004bc82db4d5f9fe1255c77c82e12e184688ab4e
z4f2242bb8c84842495e71ecf4c5614dccefd225012524465efc51407d548d6feba83208e5e830b
za1b937711984f9a7fe5ebb25f16d5569cf826bafa4be86f52fa042f1d09b781e110399c24b0064
z96b2c0bbaab6af780776b3e082d02f405ffd420d664f09fa75c453b66fe2a353203c15b7843303
z5ac4aa6cadb092047116c35bb9c17ed14a1027f12393bdf64637f08f476acfa9e2ba8c170d4017
za10ecfbc407f6b5cbd88b43149ff1ab4e2c1e29ef320eacc4b17bf996b2ea4d3d643e7905493f1
z218586eb01a540cfbe68546b763965b4c5493e108b5ac6ebcc583e4592a4fef4764b683844f30e
z314aad46b3eeecf1b9e17733694acb4b7690829483fc70b994aa63d8d21cb422f38abf209b9754
z6817d9dd92f452cd74876e24ed781319a870104add302e8d3b5a8f8b1aac08e0eb308b43f7594f
zd3db330204cb10250ca5529a7fbeffea7b6c6b017f918ce4e4d0610c254380469d681cf7cf9139
ze75123af473a4ad61b27c8c854d74eef8ddf7e46694b92c33863f92d08dec87eb6a10d0edaba8f
z91279c1a302c3d1e65971f9ca127aff6125f30b9ed91e6e600ced1972beae1b95e2712057ca0e5
zd1d1ece124e549ea46a2321f0e0928a3e046f2fa4752e5002b9c87755acb4453e4f5a87da32edc
z537ccfa23572b92e42e7a3877c8533e6c6b6ccd4016c885d985881dd8f0d5e596ab5153195c72e
z4785b7a898832b55e322beef3994aa48c775dab22a5b348f8110aad8ada5ab8e72283b2d4ba0c3
zf1e3be104e958361da0ac27f3717f69660cd87a734a4d0aab4a95bfa93461b75ecd3431ba195d5
zd6ee95612c903772b0040f718e2006eaeab2724e66cd088c2ef4d9502db524980592fcf15e723c
z1dd1a3b38e8e1ad0c529d944688f0aeb3814c4a2394cacdccb2f12b83f4ee56771e0dcf523964e
zd88e16bea1982de33a59faa3501fa3463628c57f5daf454486c53812292250e30393c7c7b37f12
z4422e479a9979161c4fd70f99283e5790a875914da6cc08b8fb5e5283d7c878e82b87a767020c1
z186d5c23d772dc7980510e7b1d68444b2d7067d74f978396326465d79802cf84849b4663d78efc
ze18224088df76517483af888752955f7f0f8faff073623608ca6ecfdca7578f02286c953abb061
z260e067d234286c2f9430f56af10dd996ea6ca6dca8eabefe104e569a4164fdffe400a9258d820
z0de56e9a7982780938a6aa30fc84eac3f10c411144800d1490a08ff9ba22eeff41bf27d0dc6e3d
z471e020fbcb72672208ddc2292d33be1ce524315de5ef3ce792a8bf3854963648c3970af0f0d33
z7931a341975ea9ec160777dedb0e8d76591b1d32391bffe871594c1f7343a5d9b51ea69c173459
zc5d3f3eb61634177091965d16c284ec24677a63495ab9591d4009288e124bd925c22c0cc107539
z02affc08d2c55c4c60dabf05ded268edaf763bd68cd8e35f99b2db50f56bed025fb30716fa731f
ze94ea1a4ffc55292312fbeaa4fd0a0c24e5931920c337f707a2411dd4704fa55135179ed0f848e
zc3b13b1d2c5a34a8ea1495d5f9f224758533a782a4d86f1951e3f69e07075deaf666de1ac1b581
zd00b67277e2a8edb0a2b25bf0ef4d22e4fbdcd94128516141ed552e26281907126b9f20aea50d6
z7d019f9c9ff1cdc6ad29c712121eba583ee6cba215c66fcc0ef9660d0400ba802dc8a3022e21b8
zbb409627fd7c6c7bc959417d219fba1827d1afb1a3a85f8fe859178f698a77ee23f8d11dcef537
z85fa671e3dda98d2a385e5a40f4c72a00e3d3a5a82101f16170f03b8ac8e9d1b03370889d91294
z0b5f8467aee5d697a8cf620e9ed82341db6d77108fdf140f717515f420962d3a629ed27103440e
zfde7b03acee0a6d7d22b91fde8bdf4ee14cd79889956ecd42d20cba2fb62cbf2fe225c374d7b46
z6bb3e906846321e9ed9285194f34bafc701b46f295fd0d138fc690148bbaa9d8e36d47d82b90e7
z95f90b4b883e616f271c46a2cb70a10e53ac36fdd110491d6bf20374fc5d2d9ee6b1b8a19dd62a
zb8aa311604b3a8615d603c6c21ec5033dea733e1c8347f5a109bf7a94070cd1be8586628b39f95
za79165df30412d0034b88b69760d7c5d675161703929df788fc917dcdb4905d411439612ba9d5e
z2513557d322a5181e10f245bb568f735c0ab7e5599f8618e73a303220f7dac9473e59d51e69bed
z365744cca36b273a2ca40f478feb28f742a6ea2da91d0689893e3e6ea0b8bee8ca3277af76ba7f
za6f0ff06bccc2bda25561b756e2a6647512e84aa05338661aaaf2dd4bd231208506277be35e9e0
zb358a72b1052c6ff1b028d7a24acf897202f837ad869c61fb67360d7f15b566786fa879ddb903d
zcbcf999047ef99eddfe7144ab67655529f751e698903c5fa9d68bbb6270bd4506a6ee9518eafc4
z5c8880f67c7406d8f6bc1458bbe41f914588556412fd89919262b7d2eb0f605eb49fd30a260592
z30db3d2af99f153f302c9a9ca78da58802ed883ef5838b50d6de90d55c73099140f07d85b675a8
z097545c0bee0428e3486be2194a0bdb0ff7158bee1ec5e7837d6c8df725c844dd797e2ae26db67
z2a93374474e11c2917a9b1d1da135844bbee2ec96fb48f8ea2b46610112c65447cbde0a7af6af9
z6fbec7ddfbbfb0d63867d3a6359b37c18b33eeb62135e606c6894be72fc25b7abb8c34d9385744
z4604cb53f235c9e6d3f207042121ca6c74e82cbaea0b047e77898fe3e413c4811cd4e6a8950b91
ze33a987b8ebf944a2adfb27961d9153132266bef2a5872f35ca5e4c49cad8ac6b4ded76edc59a3
z58273fa3dbc0898f9abb60857a3d412b1676a31a9dd911f129862808a6a6df6cdc18d2b3f3c5b4
z6d5085b9bfc40ea2e6be9e51be952c9776ba3ec4a2cbc60834f3d8d1d6f81eff803ccfc0ca5f34
z650014c9c457f77c56b02e09c31793fb92bd5b024821cf2361edf85c5019ef1d97ec54e8c5e226
zc29cb296af2f058c5cabde999c5c55239683cb9a24081bc902bdb197d4c7ca00e0be0d96c519aa
zc8c6e08085415cffaa99972fb0297143572b8da6a9178c8cecc251b5c59a66e1e00f9e60f5718f
z27f5d347c1fbe2a906b1281384ac09c64753db21333915dbefc40232085a941f0e5cae5d1635fe
z3aa8a6baecfd72869b5257daabd13b433bf4c69a16c5e31edda44bcb9218dcec53f398fffd0636
z89a3228a40b269267364d580214f437d7b94260e5c05550e5e76a0a1e1261bfb497db2c18ecd95
ze026cdb5a0c3967e2e82f7252974f671b4e00750c05d84dbd5f90ee899d6121ae12f843558f0f8
z5f93857cca9a4af7af9ef4e3815de430e2233afd631346b32782fd561942f6a3034577acdcc2cd
zf1ad2366b62a6c8c4abcf0982c65fb3226b9eb0e012b690bf05afff8f61c756cf77510bbc1dd19
z759960730d73253f7ab9ef9d0804277145998a44aac302832eae57feae430502b541de734fc9f4
z46043a6debaefd9ca09737968065262c6d3c9ef2b561cd6afc1becabd163353b104535d2249566
z52126e4ebe83bc33fcedfd89b67aa7d5edfd2a70c4d7e3f1f6b0f3af2aff01a0dc8fb032fe8d3b
z797a8ef5b6932c52bd75c1238c1b7fedd5ba1f1b05f473dab73e8b179c5ab1b8d9cb9bf6867032
zd3b39f820adb45da286e80afac956d469c19b65960e0f7b6748e639a80afb17d79e45de3702176
zf0d72e126ddac5301fa12179ed456d5a4406e69af51180fe69265dae0ac6d70d0ef8f264c4be46
z34820dfd60daf91e1dac31421c4af7b50cae0d5b41a5eadfb12812ef9124708aa262505e370940
z1f6918c44f20787b57ed01dfbb8171b01886fbe6784b0812b9cd7195f06f36b5c9ca9681b45bdb
zbc518b93ffacdde6353e4bf672d16c3b6bbdfee8f1cd9e46ade14b9ff87df4eb80066d24fb7559
z82a2ce6032bbadfcdaa76b94088dd46cdfe558937ad7d1ba8ea3d453b8587a162fd7c9361912ef
zb7b65425b2bf4b0d2b29c791f8a292cecb5de0085168eb832a1084bad9686cca4e0768124388d3
zcad85bfed651ddc551ae336a06c37803f4f316c2c421dcaf4d079be323d060af274588e66cf2a8
z72a02df01459221eee3d80e9ab73a5858adeb32598007a390026f8e9096619773742d7d54c6e6d
zacdee31b7bb40f3dfc45377607b0aefd0d2f29051b1d33a43d38a08c705f7f34a1f58bac47c73a
z50cd568fd94cfa8d8ec718f4718b7bd7939c1ee37f75110e2ef8d653336585038d67ec5a8fe3a1
zc3a5d0aee1ca2c66f46fe3cd85720c5b4cc93ff7b6dcc29eb39ab209183f0d95536901675d98e9
z684c8ba8f9a031ceb7ad6b01ed5c053fb119c0466e34075b9b61fc2f268cd2c6ae1b3e2bbbb5fd
z72325b85a78090b070ead2c20331b12eff220885cff463e7d6671775e2b15bc66e0f03f990bf97
z13932ba0a7344f505c52b29a8d1abc2b5473edc2be4347df47cfe7a4f46a7caa7da434eccb4b3c
z900d9f7ea4bb7013b6fcd77ea717f448612efa318f97cc805a9ea264b80eec5d2976264d9c79b2
z2e837dac9b9e199adf653bfb8109652ea92fb2830a2b0e17a510a41b98484f608fbd1e577bfb7f
z2da7bb6c60e5b41f0f369d0b025aac402db9b95a219a4f8e6a9d5eb4d6775a5b3e68bfff0216de
z9633d073bf3303d36bc5fdac9a7eda3e1d24f7c2b6360f86c097b2ee505f1bc435e5e903b12a70
z7d529cd1507a45edc0d4e4facbf1e5df09ab0a8a214a4d6b3397d6c6e021251d0789a82fede76f
z1cb66e3d9a90cd13913c4c2ba421d6d87b8948ffda8dd2a5af3e2a66125d39e71eaa2712c5781b
z52cea6ae93213cc656cf36c45d00993247982cfbbcedd2409cd3fbada26a9ec0ff13bde6f2cf45
zd0b66528f787e4f15c9fe83d1924897594e3ce4b908ebf27b8fc6c400c0c5d95ab71ab7b2250a4
z14f215840768adf3d1480ee99f47346d3cbcf7f89f095af3527e62a9a4e0885ed05313de2a347a
z47d958b866ee62315c1d2ce1e78578b9f04376e48b452ebb453d5ec1112d6592a2bc177cd0978b
za3121ca89c94d9d8cde5f513171bbc18ab059e2ff292118e7f1775f3b009cd9146b7186f90c962
za7e4b65a27af43f0affd2f239af85a40e2920ae4511f6e751d42fa296f01e65638c517ba5e864a
z3531f135406bdee46970879dd48aa5c78fe64f0dcaa56b07c7ca1ad83ba66725b56633243b4c34
z1e67c05e472451b27cbddd0de8159b7d723d7ac12d0692491a52cfd7ed751b067ff6a1e87cebce
z3a33d733b7bda654d4d42a8c8f18002f8816487993d3dbe45c4a918a5edb6417ada5e48f1ab903
z8224a96712c7c6abb1d64d56ac5a1716610f62cc4c1de78ed0a9f00f4721148e4e778031f55c6e
z9e96110f4052f67c1bfbd256cde46e27708145f8fd7070b10160799572de44b27431b34a37a9fb
zd6969432165c91678198d0051bc6d456779e30121bfc88f4feea1abf13f84513bf0fec4cee3fc0
ze5c31ac3cc02533536a041ee43ace16b01e67484b4118dbdfef5549907a1a33fdb693a34f5a03a
zbca774cae6d6ca19343552eae76225c8ca334303639a67b6df0e651a3444e7b82db7db2e9a3f71
z4cf1e2dda4dedd129f8e0e86c29d5435f1b7674048ca63afd83e8df88768fc00fb4b8221c4dac7
z23769f8f63d72418bd29853bb41b053ba385c106365262d006b53dd3d18379a09eac3530dad615
zf4492da6a47f9e10a512a15cfcfe52c1541ed69f928b1481e49857a2cde13c4d0b2b20305a59f6
z4557d9aad887b0f2076c30551e30c745aa0f03305330c8c0de0e9e63fcd7bf1ddc20949dbe2113
z8cd587841856bbf666dc6e420dcabbc599effc120742f2da26b023b834c825e6a56e5910e0d67a
z93537eeb07c03e7f733848ce31cf5797221c9fc23b330f00a3e1f5414b8856170a4392023ef972
z7353e0ebbf88c2c958d756f049efd4c525f364b8bdc9efb0d274f52b2898a988187144fbded629
zc2e857c8290d38424e2bcb050a1422e72d0214afbc89d0f8260232b9a86c1508f641e9adc663c0
zc05db93db1685ad105f62a331bcb2b2b3d4ab7c58da8218669d718bcc0251035fcee6809fa2de2
z13730aa66d1d3afae0600f4f596a2da0edc8e4d5a00cfca8e5b343e27f8548c9ed69d0e00e5ea2
zd5877240053399fec8dd54b6e1af920b145c01de5d314a66eeebb635a2408dde3bb97cb36e685a
z2905a610d15a9f895c3ac994675f93297db0f5e60faa69714541883c1498304cc4830b3c8010f4
z5b8042a5263c72292ab114c3b8ee25d50971da72509044a72a2342831db788ceff4109dd4e567c
z2a55c99e1585f1ca0427c20c2c4c3ca06f4dfac4c4e7e3b2f4427207b8b3f53fc2d9833b2fb9bb
z2beb56401cce3ddf5d8ed7d13ca7ef648c9074dbed901e4af5b0091fd4255855c83cab222750fc
zce94ec9f262d2dda230629b71d883c94d6248f18d5d7796a4a6c0d7dbc9e7504c351f59d5962d1
z9a2bca21f509a623cdf8f4db5c5d25179a2526016a415b7d2c295e19590edc82969799efe40db4
z2e1c0ea0daf7e5aaacd09e076153f9fb87a67b0598097416f34a9260bbceff805a70c0b242eb9b
z21fec8d6aea511fdd0ef1b8f87e7aec4bd858ec07e36b6f33fc580bcc71aa30a74357e84042e1f
zf166ecd9576ffa0460e8811ed34f9d3f85fb710f941949cbb6a2e65ac4c40b9cd076ca3d9cab32
zd5612c62f84790927278901cc9b2c59acf8342eb9a9a995a160bcdb43892df1c339b7d5054e4dd
zf5c335f2cc277fb2906dea16be3c1aa3397c6ebe3dea1cb7c4f1ff64f940fc8b66eff870c61db5
zb5c540e3b44e6001ebf9090ef6c65ecbfddc7f53bf9d09e8d60acd644764a530c746804234f50c
z4e49ea4dfd7add744dc3d38cccb4b53b53341148f311b21f4bdafe7abafe67f51d065af35faeac
zc39c09e0fd50f56fd855ad50d83786e623aaf69b40801363d6c50fa6dc4833c99350c83def4ae9
za9dc0458af8fae63746c409ac881cc159c510a5ea612b9d82775686dde48a5cd812f4e60b045d4
zade087b4ad4a214cc9fe565aabc4b784db3a2c649edabde8c3d6a93f0a8f7e3340ba4791b8161e
zb705103816c6cd930eb0606b0b15f2da9137e65a73c316d23ab45f66c8e57c2a4be67f4df21c8f
z3174ff498518caaf5b809d5008e62859b5165625c03ddba50bbb02f661391e39f9f4c6072123ba
zb9bce3f51576d4e8ab82370370fe09dee5bd804bfbc229a6aca21e0c38e5fa1b31be5ae8839e12
zd7d6e27591193daf31ac374338048dc40b42b03da7843bc9b23953c30419d1b89a23825e40a735
zac5d62a35717870740b50887889bf8c7819ebb6a923f9b4a1728be04e3504bef8dc44e413b7174
z0a72c23a0f9bfd04b92e9ae9d186d19185806fbf6866fca123cab039254fec88b5832af675f8f8
za233e8116b0396839b87a4306668288a5a2a4ea5d4625769998f997c12934164a47c2af923572a
z946b4c1c84d365aa841d308ad7affda8772272edf51a00278997b0b587b48285d0aa03f00c764b
z70763d0d583bdfe499c27583229b9a970c72fcc6b02f39e215ef93ee219dadc63ea99fb59ce55d
z8e4dcaeb08bf5d9418d540ce761ab356ed9698833b28e4b30dc910b820676f4ba62890500d1cdc
z23d1156948a6f348c41b5028baeae1f338a704790b73fafb6956447590e40c35a78928c4ec1450
z151b226289c2f2593d8ad88a5e83543970c746f9c0514acf8eb7ea59f772729986ed17b5389728
zb3e50edaf5786134bb6b1c5d4b7971c1f468f4fe96c1776008f8134781081f9c4636d9e6ca2485
z7cdf217099679c92f1fbe4608a2d6b29db2091c09ecb3f56b934efa1db0d2ff248c581d1bed5f0
zc02990001a62951acfb1b19576eb4bb134d582d33232d37fba919049aa84be59f77b7eb9a5bde7
z34d629bd3cc71b4e99760b64f4547d1cfeb6536959cbddeabfe9e25347b6b76d6a21c9fa223fe1
z7695b9e49e93d92ac457990ecb3a91bb37648388d73c21f267197410ecb995821bdd752612c74d
z77587b4f9291764122285008f9de58a388edb36fae64c61df5dc1acb5e039f6d5b4e4d6dc11a21
ze584af74352cbcca68ebf11336ccf252fd811ff275a5b26ed80f74e46f9bacd91117bac04146fc
z394e44c289f1f8ecb635c2c1a2ece7fccd4a8108bc6dcb5017a2db0a3fef7401508cf5fc196410
z2187bfdd9895989ebbad4bff8cafa7df50ca3db69be5e80582b2feb4a5ca666398806bc9b15421
zb55b76fa78c06eeffcf0aeb232de0ecbd000005127435f80dec20b9eab9430c81be164eb6265a6
za8aee243fa1bc4b378195e6c3e32ede2d13d493369b8c78bd7147f5137dea8f3e9fd0caee61b0f
z35f44ef2187389362d1fc0337f07e28cc85a5af924b57d56ca9a967e2e026a6e90ba0f44ca32bb
z21538e5c9121736edd11602477b0662cbd37e708e4225ad8de8f7f35a50b8094add389507b1af7
za858fa9fac6154d68b0be9438125f498ce32a115b856d49f5ee2aae8e0c028aa32591177632d51
z827f6912cf7f0f11f3e1b327fac560fef4a8fc59bd522e0047783de53b784159f27fd221127d5d
zdcfc19c746f3bf483c3b5f5ca4f5b9d4c1a7a6280d016cc884cb5236eed7b77d5c3215568dc859
z89617d0a796898a4cd464c95ed5277acaebcd02849410e5fcb380d70f59f3bdd89c36128dcac5c
za85a41dd568df93a236724a2d4663b99aa44865817511ef04d664fbd75c62d51041b8389197c28
z7f98218533d72361a691e2ac37fd4bff172904137cd42cd5680fde53befd28ddf7c4b9551cfa32
z7adb75568f629cbb3ef0f3da871d3f238f3bb8b6ee1e4496d2eabb9973e6d81f43f5cbf1bda5db
z1a5880fcc57712a9e6cd96c5c65c2c38fdf7322539c4d306f63f45ab48c6ceac5d47a0af2e90d1
z447bad15dceb0622ed01ccf11979cf2038b013194a325f60529ccea530fbf9488bd80f3da25f73
z63ca7ea68eb468c7f67dfdbf6d89e47d9ad5a854f897e9b70ead79bd26db755fb52872b63b7ca8
z49d3e120a8bd871bcdc5171db8af028f6fe00b27fc1b9c278c1a9615e0258e6aae45d0b8a69387
z81189ef96177b6cd425a2d600689932fa1b3d741d6a7cea7b512e5fabfbb25de6f459feffa2753
z6a82f7087ddbaf0a0abb6f33119ed64d22a04744b1a990cdffaa4412de18eafcf29cc8471c7dee
z263ff49f534bd88a44403f4a2ece197095b0a765d2c5f2feb00dd9968d717de29928fa34ceb93b
z0e84c41a2e1753cdc2747fc3d1720103c138813b00480ddad2ca988e7167b34fbadb3b839d1cb5
z265695849450334188da4b9480b654fdd587282ec710de21c78641384e2f5440b14a5c58be497e
z25afa22caa5ae1b96f9ba781bb8122434f2246019dd73a7bae154ad1fa30df62bf588a20e032e7
z6b1633872dd75df501ac93bed146068ab2c3274a7834ac3676672e431f0698d90c6a599906c725
zcc9fc43b4a2d729bc8c9178c2758b0e1e5f51205583dfe489271e0f5a8712cc35d91c20b1b4546
z492369556d3a0db2ea15647f0f8b2d5b1261ed0b689a237d730577e93cf147d4da23e24c44dc06
zd3e9b551f9165f1c4188ea0deb9b3386d1e0ed2fa55f9adca9b2b39dc28a9b7aa01d3943c3fb5a
z940716d6d56fb5622bba8b4d11ee3e54a4af73765aeed2451f84d30c6f6efdb3f1803536ab29b5
zfbb6478cdb4cf1b30671dcc82bcba994831382648a1228df402d889525b68211880a3afec85e94
zc487f852b765a94ba1e5a40b3550e0e8beb1c214997233a9c157f7d4907e7bb24e084ddd898260
z5e8229979f23d3c33729dfb030cad0efde40e38af7eccc2aa10218c5538e7d202b5ba18b3508bb
z012c74a4b09ae7a9de300dea098183decd969b822b28dc77716875096b0f57a1b088dbd2311f48
z4bc4efe33648006c7c52732ca6d8e3bb027f93c598b7afbdce82923ba3e3594d9edbc66f930037
z5185ee91f672e38203779d407458739808406501bad70af6d2b76338024d87ac4b01754a3a8c84
z33897637a6a6825677941e5653c6b1a542bad1f7112ee8767e671aa5c9ccf73a0ba2834e3bfaf2
z4baf4396a7b85d7d5788ff9e9b8ea27f6244a52851e97a7f7dab49d8c944689a0fcf6b0fc04048
z0407c408ecee85704631118e3369c96765ec0d2e787e81fcf9c877ec49d3889fecd8dd830059a1
zc6b32f955de6391759a6337efbf8eb8ef1b030194ce2cda25bac1d68ecc1de267d883c0fa82ee8
z0766fbd100bdaccc10f2d0354841fcc7d5c7213e20c378a538212121c227e2a4bae05c2f26623f
za02cd616bd60c4c90bcea7d3db7f704cf05d126dba35e9df43d491a1265870e3ee93d8ac36b347
zaad86de0979d5f3260fb505da90093054951b1eb6e3576159739788cbdf92cf2fa404d28dd99e7
zc292ecffd1b17008da5c039e49622239ee62406fc3a319b9d86d17cc2f2aed23e5b661b772576b
zaa081ea88543c37dda9569e3d83b728fab1199374a29997f9f41286d7306026369dfe40dd6d89f
z302f8ab27e6e930ff2263062668cbe5d5d978bfbc7cfc119d23d26715adab6eacee8eea86732b5
z0788afc665a28e1e1f5b80fea962452ea1b4a4d738499e7ca8efd889a227233f7688a5709b9cc6
z2c0c0d9939867d0970e8e9a5a57307e2f94b53a99e97d2bce3e3d0402f1e525c81b1d99e8e580f
zab270bb5e828921cfa60b6ae20460dac8850045a8df6320f476b4a43dbf5c186413b2a1bd29a94
zacd8ba06b8b29777efc07c5b7ef8c8ae22383f93555af5aa095926551fd3659db789746a15b089
z479af9a5b21d59613bea6d45d2f494e305dae772f374b72183fe08034ecab206fd09097248c0ba
z854144b45d26785039a221b35025292461bf816bbcc31d28bc2a97af9e099d5f3e040bac4e4438
zed393161f971d350a9e65069ce4944e111530c7368a032903b8e07bf5d4ec9cd90352713a1154e
z8e55c020890d282c1e67266bb37888a7c582473218b9a86acf08dca278f8cfb34512cbe30c2fd3
z269df4bfae10fe3277dec8c738f6faf49c758f250b66091e730d1a4928b94bbe69694580059ce3
z42d1ccba8f055cf0d99dc640c4dd586e70322ffcf67f822f38c777c0aa722e2e25125584d4385a
z722ff6547bdefe76a822a03e3f85bd21e4e0fb7aaec0eb3551f8a6b4029d803ab81999fdf1562c
zb71e215db5539934aa8bbf33e4eb05c4f14e8683c7df416ae5eedeb544a53a6ae7c92f5e463563
z6cb8799e3f43ac03d03ff1cf33ddd7fe8b689c9f5a9a6562e0db26085fbf66c476a9b76c3e141d
z9ad45a02082c99f607b3d89333ed4d1bd1932d1807d7a3515e69c68ce151d390499988e6cb6147
z213679e9fccdf0eac6d75fcab8bbe7130f5680e6202a2edaac345fd2219801da9ffa4055c5ac6b
z0cab7224a23560e4feb992682cebcd24d51d61d610de8d1ea7ccce596fed4f6a0d93209b575fb9
zb88ae29646a09c08f03d8b7cd2f9933da914ead47d76d6b89ec18dbdf522d6aab950db8bae1fc0
z21ce1f61cc2021b329a17715c9ac2e78852dc100561d8eceb4cc2392837b22b8f2a4da89951100
z09024a32c2ca9e7e9af167d3f6733f3b2d8ad52c07ab4681be78ff51db1b8aee871f3efe24ef2d
z0e101b47c066ddc783b4b65dcca56b3d9181b5d447d044550441c040f46eb37d26465b2a3e2958
zce3c12b9cd6add1c1e3cb3df698f52516cffdbbbcc0154920630b1e54d4172cccc2ba8c6cf02d0
z40d503c0888e2da293467e804a5f01c21302e7170e9f45f8b637902819b6c952b91da31211c392
z02ac6561f60984ef38b2549e207f6f49e48a8310681f890b8fb951d39f9fb02d7795008a1b14a5
zb76c0cdbb82a1ee0e0d910b3547192a334d2b6b28e422fba8ae82ad3c2eb3936cf1a5ee3fe14f1
z13e259605bad37ccd0924f0ddb94d75671124335fad1accfb30af798187a33e31a45f867fc4e20
zbb60015b5c7eac3a8d42afac09dbf9159b4e78dcc92f294b1acedac8d37a6a72e7916d2026d007
z5a0ba813913801fa0c7acde56fb73a37292e7f2ec9f4b6d3904a3d8a505d4d37bfa0122b4861ba
z67c0c5fe06500f2f3130562e7e226f41bb2e1fd76ec12658788a99bc03d6bef1522ba2bd5c8262
z53ad67d0fc9c457b68d5aa67be5f6779deb59c4b9f6e52f6e128f7d5f3b43bf0279d60a7f84134
z64ce1e8c44e4a03c923cb1379f1675404c09e545b9484f5b864b94096c9cadb502cc5a2b693570
z064697f7420e703f8509a3c01a4d0df30e762b56fec0ef00477e4da6bf8074e0abc374340d2430
z2271eaf17b4cd31bcfdbc87120e94fc9c1793d326acbd979d463165ff8d9e07dda173c1708aa5f
zb3a74eb34e344cd12bbeb6bf86dff9032d27b46602e65af5f3e67acbcb0e820a892f46c33847e4
z2da325dd763b412c25e01a9a49137e11583f1730886027b2809a037e715c662d6ba0d58ae21f4a
zbbff46325fa5c6d75267c674327179e383023520d8c6bed243f9376e5d9132dbde8c813eeb7182
z8744e98e9a6feb04ab646cb26aa6bc85ecd14afca9b330c62cccfd35ff7bb979c46075fbd3f005
z21882dc12c8a87415561529b9e2d4b64ea1e88e664f87bf396eb5d59c1530ec9afde92fa1cf6b8
z417bdb58614d1553fd3b97ccfbc9ec1e33572878f01aa00010620080eb188ba85020d4e2594019
zcf3df46abf74b4a421d5189cc562212f60d0775dd0aee24de17ec52f0b188be6f02dda2752060e
z5967ecbd3f9e59abbf1bbae9b7a7507b3a25b79ae848db687178c4960ae3ed4e2d63fa829e71d9
zeb4e56c74547dee9a88c0ea6ca2dcecd0d33818dd35778c0b583c2d1b4151f1a0ebc0f8cc81fe5
z15eeb9095cb551f367890a25ee5b170d1546acded080c729b64e2902d946ce4ad86f51a704ef72
z1f77ddec86c03ad02c3a829c345aca4b15d99aaa69ca5ee54974efef9e561d107d508e3f7c792a
z9f9b909d31c6fdf1b9035901759300544adde26ee4ab59df75f9030e1e4c4fa0ff789bef4ac0fd
z6fa4c11acfcf966824f518d3b88c817d126677da4c3325b61b7c3f9df3afe2b6581e0ddc76ff04
z4af4abda5a80dc576f2f8c779036285481bade858b01fe9ec203c658d44d615e2e58a0bcf78fc2
z00d2c533e800fd6ad9c244885cd2f241b1802443e7e22f4452572c978332fcab49f6fba6c7d74b
zdb8457e975eb53a14c96142349d1d2de69c1e731f175c3259c1f262c6e46328ac36f4fc90d53ec
z38f7b0134aeb151883533ebbe88996de51ba22c4cc7a653f714e392dbe7246bbad6f3ee9e00be7
zff62e588316a39cf4959973115d7777e0568f0de91755d737c48ccca1fe9b2e4e91bb5090a553a
z211a05430539743b556db4353bee29fe4379e47d9c25e3da11927100e26c1c7f987bc6c4bbb64f
z4ff268cfcca6e0bb95117bd2f5be8e2dcfae357e5d4fbed75172a015fa883f69c92876035471f8
z548dfce309691e5bd020c51adb2a2c27ca2a7f938738859159bf040dbe4f4ddf4b637a9a0adba1
zd2211245503599dcf70881a105c67ec4afd8f8d3305bfbeb67cb876415bf003b9a79fa8d0de032
z1eefec415b668484a252238fa8a457cff7c195680e7747ce7ecddb523b909e3797caa71cec7c58
zd2d87cb80446bce81eff01ec987673c00f2d5664ca57fff9e04cb29751d5b42508d07c9daf6efa
zb92aad8be5c5fa89abe672a95f826a9504e84f3ba4abf7b8df151b1472e89880e5662d7c2abe9f
z6a269df65a6d280ec3b10ae08047209e3a8fe7c036edd953ecc9773e7a75a18a5404e002e77183
z04b756d064f3fb330efd817d0d2f887b15aea8fd606f50073a89d8245a3fe6acaccc53786b19fa
z066c28403dde78fb1311adc11bdfb1923eb2e5a9f6c87bd700d4cc6d931264b214163327d4b937
z39961b0a02d3d08ce2fa6616ced5b8817cd1d7d7d97d83cd427cd773674b3c28069cd8c3ee35ec
zc1f9f383e83c9500ad5e9a9a2c39eaeb7b34162b536c92d6d1770a82d1b5999a6be832adb3a532
zece5163b9fd67121fe4961e426fb4dc32ef863e910e4e427254e366de5b4a105baa579601f093e
zcaef5e3e3dfb7824d8e9ebc42b41506589635c703fe8286ef82f4554a922e30461a504515db81a
z83c9d093d0cf3bffbcd792f2e5b719004b1c1d9f149511b035712a1cb9ef437eb5e98b8f06a84b
z09bcf61feacb78342d3674a9b9b1120768c819f4e0ddc4391ef635a0268bac30ec1cea7165d489
zc8ed6502bc1844fe9a328332176fe13697d09258e386b35a5188a5ba9015f3b1aacddbe987811a
z13a818c8e7c39d5fccd3ca5bcb9a09319d987d1badc85975781ccf77383d94dd5dcec6ce99dfa0
z89a2c7f186cf0900a11b0d067fd3796a92162c4326f55a433cfb65bf56ec3938b1d251cf954d72
z297acf1edc948cb3aa975bdc0781cc493b38281b494dee11d6a2a22c340ba54ba2441a64cc6610
z6e8ba911a081591b51a46c75578857fdc2f68896673696e86e3b86330c0de2c9203a21bea16093
zb4305f36f6821c7d73716b15e0f821bd13f472a5dcf9fce54153a999f6ac8b0e30b713eddb13fd
z799378426e4a1c4a929b163ae3e8e485a58666c5b87a650f5beff43dcc18543e2019724494d713
z3ce2dcd467eeb61e77127c8e38494ddc2bc91d23ec2f52ef593ec0f3cb17839f26877fbc225585
z71ab645c787d36c1c74e6448d08b54cc059cb54b70c4c093b488b3be34cb577a587a215b326f8d
z1dab1be9a1ab2fb3e5324a7eab801e4efc8733a9dfa43c08b4d4ccab0c401eea87f51745145a4f
z46fb509e9fb41c7fe7daf1c952130095c6e0bb9fff9338776a41380b8e5ee606c812b1207c7c37
z8891bef4e46c3d502efd7010c9e146b5d744ad7dd615c82a6d6d8056405c5efaccc967db4a7cc3
zde77b00d239bc97a9a9668e4c756ff1434a41213f78043224c114f2aab7a89c1cdaf3450ae6064
z6e6cf29904bb7d2610eea1ec26f221e095d57d7e35e50d7239cbc71b3e8d35be214c733aefd5b0
z7aaccf22a9f5e9d666dec44cbf366873aed55c2032875a633e21fd5a0c87400dcf5902111d11b1
zd97601125b089ff46ff54773112448e593f584c2fb99a5c48c36585bc1ef32b7ce6952cf1eea50
z0cbcbf2c4166da0c7a02c4ffc9d2c35eb2c2a6f240fa8dfd5a82cdb22d18be701ec14af863534d
z00369ee47c92bdd294422bd6008bb50ccda1b2a0696cb553c6406946764a44210e6b9585dd75f0
z4845660490dc8cea168e6f86fcad46f7ace61879bb664a46b421c9986f76544c01a6402b82e636
z92595fe3cab0a303146d2cb4975a7f556fd5438a252d726da31a7aa17c0c200645195340709014
zcb63e33a79a2d148d2a0aa87ea40ecf21ef8bc669bcdb0e6cdde23a79a67dfadaf0717c8c2c983
zbc0ed4bc0fcc06bde6e3a279d643fbc01b499d8c60d5b54f64aa2cdbf406a0f988429d71918395
z953f0171b0d36701f2aceab6161e578d0c5337d67d60cca91325be16879589bbbc9f947af5b3e5
zf247ab9f03bee1c88a3937daed388efab3aebe9c0fd60264b8ca478b9faf8e188b7bc0a49f1fb3
ze83f595eecac3aaf05ca7711868c26b40eea4b7e1592247f702d0883961406fb1e41270cb5f3b0
z3a6dd3fa53a83643325f2c4d86ae6226c62cf84afbc757209b0c69be62d0d6a733c0f0103aeb50
z946174ad0d2762cf385cdf5a3686238c54e499404f45d7d531be2bd31a598a09641898b3767d10
z2531be68b82ffebdd2b494b44ce3af95e23ad4cb0da4515d84ebb1d5950e8be417e4a24f332aab
ze7ca0618aa93eb1695c1cf85add0d6937b47234a0d072ab3938c23185f1e1e0fb1875eeb3ef797
z0acb1f46ccc384be53dd725a028cb83b73179cceb0464e9680e14b6fe5fba3541927a358764567
z21efa2e0861841df942eef402f27d1eb98ed2591132ab6e9043edf1dfe2e0855eac9807dd927ac
z2592f3001982c3bf12c0a3a2531d6efe04944cf6151c1a9b170522f8a171a431d316c9f3be8073
z173dcd5d8882eb5c4de2b3f95d4813ffe49999305f005b1fca879443018dd2e5e411bbfb4c959a
zc9dea14bbc38ece8c96dea57c33b967c701f5a0a84342ecd57df4cd2de1d46688b30305ca486ea
za192faf1aa90ce9fabf7c2b6d0f87540ca38c02d72d0e9c3df8b9338d8f11968a5e817a7f28938
z8d334e821fede0e2f108f8c78c1e69eaa288010e8878db47e691965a11ecd8490b9799f8bbf1fd
zb1522d14da8a64f841ed7c19f660dd6d0be8ad5f2a1c6943892cdf96ce072dc5a8e9107a22b092
zc7729b4bacd9d801d9c7aff40c61b02afbd133445d8fe56ae2a6c5ed10c36378e9e158dc1dfd75
z72c7e2dc30466384104fe623283cda685720a8c12e979ce8a19ef58fc1f063ed9a34ca500a5c72
z2f50889a8cee08c0ac7133d165895e3232428444fb5af50aa3bcfb6ab6498f287827ec8dfa81f5
za2663930d4ae494b6d5ebbd3fd98186a67156cf5ae05354b69219345ffd92bc0d194b74aef1b84
z920ab51fffe665910a142002b078c187221ca582a5f8ef79d923576495a465dbe9d3d4ae47b6bd
ze0747fbacb25f1d8c29bedf3979066c169137f38a57d18f1c49159b0a3b3347f0b7725cb86a0e9
zaa947bb2421829f4eb3e00a81eaf228946f013e873e6ed9383b03fd9afb95f873647f7164d4221
zc1826bfe1688c2a55c5385398523e42afb60d8427c002e98447ca613782e31eb38ae7dc6b08a45
z9a6f08d4baf8a06c56be43a74f74570b4468bb42a55bd0bd2b444027da76bce81e492eff15ab38
z19b0dd14c3059ebb1c1a47c6d34f648bb446593b6a57efc3b0fa6ef38ac0b82926a322653817a0
zea6b9838cfe9fbab247b008dcc20586345b1c25272db1675cdd3b6668139c5600f63cb47775674
z1cdf25269b7c05397b1b9c78c8657c39f37bd2560fd2b775242eca9c01d369c04f1bc216fdd917
z295fb27c341cb1b236208f6855f72b6030105398fbcceffe7df06e155981b09b9baf4a7c45f351
z97343bdce9a20a5e08c89c7c09321a6a08f056972d52b48f21f98523e0a2033de6fb0564b42740
z04db0b41fe23cd51d4f057de276808a858704c3daa0533591d1f2a826f21baf62bc8fe74cc7dc4
z859f9ada1702215717d8a22d5e147ad4fcf1c951145b8d0ed5c1c959df0489e4bdf696929da510
zafe72ae61e2b52ff9f45af6b7142184057a6b810ae060334127964d24106f0ac516f35e42f421c
za46eb0223f0eeabe4ac537aa6f4b07fe5415298163bd6d6bcd8b131401ff6c7dfa1fb207290dfc
z4a9f692d00dce0c17f7e44ecb0ad77807aed397c6fc630df52dae3124fd08f9230c44b624882f5
z87557db64c36c3b3d466e9958bb5137383da2ec3e93db586a98b2092ef5860484339b974ecda94
za07e893dcbdb2d5420b7fd095bc2068df86a01cf104082d9b2bbb9d1fe129c6f02743821c67821
z6826bf76b8d86c31c7fc6b0a30daef1f2929fa37c0ca343e4650939bd2c1db641b7b273d592f66
z6a176fc0c73e17c77a04a04235b1eb2ff40d608ebaacfe00b496e49e9365fc4f5e83bc0918c616
zdcf4e21af2bd09b3b9e0a5d2d1bb62175d1365570b57b8902091920f650d8655a6ba7625b2d215
z5e22216979c2e95a8c2d081e3dbf399354b59feecc3264074d0609cb8d49a1a80c6395bad8f6fa
z1c63a6c1eb95830b4ab48582677bb9c748adcdeffec1a59f73643e7d50a42a117d245ee4a11842
zb1708cd0f877e4a30c82df7b4ddeb709b0925229902f95f403f618908681dfb71e42afa4a9e823
z3c765fbca3fbc29bbca42fc9a40145dc00c479b39fef821f9437cb364ed3d3c89706ea13411469
z3c66b0ff4fc46b4e525aa3cf3567aa34e3c39be21398e7b7a2a5a982d01fff19331a72bcc63c61
za5811bcc6c28b005bc309cf9abf0875df29962316845bdf5afe0165ac37a95b7aef8cf657abdab
z1cbf982e720ac5f8fe507dcc4f41fcbb6d9262a4f1b199f4ed64a6e6a38ff9e4821a105b92667e
z2a477e3b0c3f9a240c866440627f11be5748c896b4e11397435e47cf64d0671461f602ebbdb086
z2e0594abe0c0f2842f43a14a9cc19728b910633d9661c8857440f7a02663304821129c6469da15
z83d08ad63b7ca94e991538f80ca73b42e954d82f8a488b3a0ba1a9e4fd46d5830d777fa66dbebd
z900dcbae04870dc341a18c9b8a26e49176413ac90a254e6f6ecb398b0bd22b86fbb3efdbb24777
zf4c132978bd06aef5045cd499ef98f72d89d3c6cb11ae83bd259c09240443ad5f517fed8b59747
zdd8318d2fc5bbdd3b1016b30879c4b56d05e816080c7f2d8b8baf927c68eee0749f92f31c0c932
zcb771c10451e2c04be6e077d0e8dd4773fb244962c0d13c26777f03de9e9a2195ef2dc7316a47f
z9c165648990474473550f89832838433b91dd0b5ad16e2fa93d546dd0d3b938c5091190e5edec5
zf18867df51b7458535a69f07643f4fba7ca0f73bd97727d0415cf79985adc799272da2ee144c50
zf5148e4875af57de117ec6af5163accd2dced6fb93f0527292d5371f443f88f25b698f335280a1
z7ca310df26eb26eee7efe655ebeaf13a7474f8c6a57f7740985805089581d4ef57bea6a4fe21e0
zd2613b170737a653bca9242d04885afcb3429e71dbf8b2b9f0d026c3d909240276d1aa37dda750
z40319a8b569de61e87ecc3be623eb667e1a36482f52b8eacc3ac9214e8c9f3eddc000950d3f1bd
ze7b882dd85765f7e11941504541851739680e8292bcd16753484a4c7239ce859be2028b79f9063
zf5cee152e504e55901773c771a95edce01cdb19a36a4a447631ae76ad4794b253dbf87b7f8e2fc
z5cca3e5580d0cdf3100ab4fa114d9e9a413306ad24662dd477b2bc3ff06d2468f8f5fbfe9703a2
z5385ab509b268a1327a8bf0df5204844583d505edb25e2ccd45cdfebaf78568981c4b876f1e192
zf0eee008e3efb5b7c0e80e85551f37e9c5cf001eaed43703d7f38c4ae1bed209cfcdf6cf743200
z3d3e750ee631f28e4a47a2c1c9f1330d04933293c721a01e955128173da9aa9ab2035655fc4dd5
zdc6e669e75adf3c362d1b2070230f7ea095a283787943ccc52443aff7cdea8bc6846ca327a8faa
zfa23165451f5bd87a5cedd9665d8e0f10d2f246d0860369e7c24a4e8e527a125eee51bbba7e53a
z87c5c61795223af264bd45d88c5e4b28d2917c3e60d9bcc4bc09e7a6eec8195d08acacac186a44
z2614184a93216d1cd994ff3bd3e1122f00f2ec1bd105003375aa15b1fd66cc1388bed1c59a3f44
z9ec5104eb63ace5bac9faf91f6318207327277df8435fa409cf6a8a77a0f7b609da3588cfdcf1b
zad612276742e6e14e7a930854b85983ac0f06294d7cd880c75ad55132cee17e96191e60b3d448f
z051da9f2773fe7fde53d393e03368d0a8945dfb2f47c869467a00970e4493eed1c398b22f9b6a6
z4a434375d4a218f3f225df6ea00d222dc2310d9eaa3c4d8b8afc98f244856cabb40ac8ec6bff94
z61001895ae06988d90117c28add08e2abab969787e3daafa13fcb3ffdb77ed3c0fb053d0099e5c
za03231b761380a1b1693d23ca33779a1d686658cfbaf94ccba3e50f379451cd7a03dab10871c70
z22dc8402c15f9f1199768ac3b25cb873cafb104dfc1da19cf61367817a1614e36793129272f8e2
z42ee89961499c0651bcc77d073037d4ff368fc37755dfe2eaded31ef557195ffb83b8d7d70f813
zf82ffdf275adedbdfd070cb34fd42a7ab7e273a09c56d7ea41c246730d9793e0df1549ce366c90
zeefe6ce4ee3a5e75e2537217815d7cf494ae8f187d84e27d8f6803ef120ddfdce7750e6ef85854
zff12f0a6d8b9cef1885f2177e5cd611d3f74f078ca3114b66284cf869ead03e629b20891b92378
z5852a8e7f6f1fd8ca6c4080ad9445abfb4efb06b3928d5a732c14de7f64b69d09ccc459132a1a7
zd27fe21e7e8fb1bb15fb5d802ac333b0ad36fb9a11820f5c810f4ac19160b6b54d7b79769b2389
z0baa9ab500c37a5bf022eff69dfdc306a02f03f96c07b33864eabead59c452ecf1cdcfb4c67552
z70ca6678a763cb43f310fe210c4ea9fec5e0c351e9f08b06eaddbcac5b2ebed71a0b0e29b302d0
z71685222502430b0289368d15a838fda439d4a40f39cf1d77d391a2412b87891ff30789b7e9ab4
z888850af79de139b7f2f25468d0b2fb508c70810d662b4c7c70a68a25a73ea575216607c52a9af
z72b0ca9b79a169a64b06476b7e818c243ef7ed7013bcc12c07e543bf310b04097147ef4e8def6d
z8d380dde57e766ce3f44ae0175c178fc78d1a620b217d4bfd44e4bc0a37b4391115fe366c39bb9
z5e4a337b3452d7f4d45defc437c27b14f97bc2afb00c55ed37c97011b2b84abc99fe6b39b18e75
za6a49a44a36c6b0ca54458d60da24c4e7c0e31c0babe4c2135f88fbd2773ffcdaec69c5846671a
z531a261f9209896b9bfdbe9929e705536c115b2d24dcbe4ef5ce74c196cd4a62eca0e58e023add
z4d441dffb8c98a1e252eca72c1056602b1b244f66f70f1362880ba555b5f1f1b6e627fda308008
z27cd30e09e4b868ef1d5bb86e694e28788da87d5dd030e0d443ba540d56dc276db89d7541fea74
ze84c860404b808910e6761bf9c7fbace53a5988ba1cd670a2639cda8973dfd3027c81186a78858
z9b30690ee2544848b35bcaee6d024c6fa160d631ddcc7b70b34473757afd9cf64f8c40defe576f
z69c364a84a1492b4e23d9b9ef3f126c7fa25c1847a71e986fd8b022de4014da8684adb3dbf41db
zb2de53dc1c7e91d127ad90967ab44372413616aa668b4c2cfb6e96eb8c2bf7a585c94bbc1deeb4
zec0574bc68bab13b696e5caea0927b165580a4c24025766ae34c99cb328c3901fdb96a5da55361
zddae479aca61fd76e7f722d09dabc95411527280d2833d435abb151a878b3c059dba688936a344
ze2ac1e824f8cb61f5d27af299d02fb90507d8094ab7106c7e5703b2f04a0e44bdf82c951d35bab
z3b343b34270eb9c207404201852219239532cfdd9889fca5ff61f2add6c89685b3596f2d827d50
z0c5e88cffc95eb8ceb5143a20321d7d629060d440aedf64745590c89f5d24813c979cce67a43ee
z93e27ddc9cc62e9640e2f1e164103e255bc0550a06f7de48c3d6cc6b6f273bf3cce0354e910d0a
z020e00a60be27cef6fe6e61e82d70431880a0fedfd0d22afd68b674f7dc25975d0ae5b4e61cbcd
zd932dc9d59ad69b2ed20a8099cfb1d5f0cba9f39df6d2b8a5dc8373b898124827a9521abc1bd56
z3afa66dbbd418e470a97523dd13a0faede1159619f6d7504fe79fb3f66307da06777be5e165b38
zd4fcee2b1fa2279285c79ed1ec57879776d5cb872d70decb5984b7050bb4e50b21031f1c12a11b
z82502dd45519c1ce2465d809937e7803957dd29a232b3787085f8dd3402db171aabd308cd6e2b7
zb6ab3d2653f15c37b445b88068b63a10a4ffbd0c6d9ca786eb40fb87e9efe4f132014d4f198d24
zaff57e47c7a4c2a538280fd8ce9e807911236bee1f07323c0feff7295b5f9c5b4c9455afcd432f
z74df5e4d6159b2f429491bc9d7c4f28539c24db5283c3c268348a1935479bcec9645dfe655b11a
za972234b52b4fc6ef6261de4b79691009d7edaf41c29c228d77246bc000072a9af2a8f8bdada10
z69e3dfe5865a6dae41fc44564f5e570c6745aca1d25adb3733fa8f346864ee5031c65d06a8a7de
z96cd4b24f1e7ec3b0b42e27c7a2b9210276e2a064534d274869d53da074ae129244efc3a404525
z95eae868fea8b10c36e2dd0c7acd3d78e90d8166958a86791be08bd3d492df7fc6283d852edd7e
zed1bbb9ab88fb71adf74f812597dda79996d54ea665b88fcdf5b740f7f4398efeae38e34ba8e4e
zb6f13c2604befbd8c68e0edd8942228d13df8643017e2a62a306afe16cccb47494074cdb5b23d8
z66fb924d8e8d8b047171c753e9a01f90827d682d4089473297b294461d8e7eeb1a8af7279a9d70
zc5300cefe0dc786174dce9a976098a5d3bb74177e4713faff1c456b36e310e87b5281fbcf6dacb
z73d7a001a16964283883981c14e32d7fa0637b0190f64fa60ff85133b56503f552b8af0df6cbde
z90aa7ff63609c18ce9aa0b15a0d761010ff9b97c58d152a5b502e41cd92db339a5720b0e1a596b
z3cf8d263210876727239e4520adccba561bb80a517d379980fd259bda5667976e7f5b749b595f8
zf39627870207a633af6c3f78845445e65e8fce67a84f205676bfbca66dbfba80849f02a80f118d
zb81afa4aa9b4d2e03cf81ebc992b88149c6c307b49242d1696f050fa4d943d21c33b39c6cc78d6
ze2c9de96ba25da34429f61e33b6c1f0024506ac6241a6126bf7d418a2b8aa3272c10b4536cea2b
zfac540ce8f74bfc52fb5fecc6ae488a3ceecd62aff51440d367d356f186e56ce8323f613078a2b
z7d88c028e46fe1199d5b55c547775e5fe97078e849e7ec48f5427e6ce02d0501587d543cb6e4a8
z905bc81617d8f0650a74f05486494624ebec73e58d77705a79bc85508602a4653ea7396382087b
za41ea71b42ed89789fd8b6864698e72508847a83c9912e122ff5b08d67b286a174788c2e71137b
zd952340d9495e0249b512ffffab73ff0a0fc460fb318af8a340c12fd2ad41568c20658c97b7c5a
z6761eb1b1979496824f12734c4cbb03bfeff5fffb8f69b43d36ff943c79337e390de1c20cd9318
z90cf7417182961af6fd5e9ebac07f2b1bc0d46722142b64cb4a5d54bb5f66e9c78d4ec5c8153c4
z381c57ba374ae0ad4bb1c5b40cc160c143e93d33b5ac0de6f2582bdf3e2a5b99c849b1aaef78b0
z8e9051046c630b4995134ccc153c7b564b5eb1a32c366ad7bbf1ba738ceb2f642f3c95f70199c1
z353d15719137801ed0bb2a4d946d96d72247343df43857f24816483ede1f3225eb8a5c15874641
z852a34adb81b92c8c33c8a4b54da802f88a1148eadd71ec2964e68b54ad7edad8e47d3537502fb
z0e9261c9b579501e0265daa0e35154a90c2926aaef453ce74421cfef6fa30655704200a5642898
z2b6fe60b6e12e9dceac32fbe8e5fe8f2f1492f22d5fe260897308f278f45d8455fc52e8b918beb
zf267695e5eb7ebc09f8c1ff81b89e3ac719c6e3b68b15ca1c7394fa0c664e5f6325f1b0641a72d
zd53350da9cbb052fe181cb30b6972bd826c1f1209fac925ab14c14e3949ac6c332aef83c7d7783
z4d1828d97e3cc04d8c5409d708e7576fbd995010cd894b3f6890a709ef392572d7d6d2639f93da
zd9ae9f58c2ddda1d5ec31bc62c7fbfcc60231779d53ea5003d942b89c9ae72c14c9805e36fcd79
z6cf9ce27ec44b91e2cf062485c1669a3219f27037ad5725e9fa6a5eea890132b471abd19d0cf20
zff678597db74e8eef278eb46bcf16176e6f6003ad03f00d5170d8f2913930f25fce292b18bdd2c
z5763550848b4755182b7067906cf5de3a8ed156cff5abecce6c889a2e9fcd1c614e904bfac85bd
z8858f81193be32a88f4cc36ad699fd69861ea1d839e3c910db2fc991178d5edc2f8623ca50aa4b
z306b6004db32cc24f1ede68148c770f8ba1444d219aea61d40baafa01ed0419ce7c29fbf8edb4a
z6a009e03efbc837afaaf19fe0ddda15d7d15cf68e321179c7f09b5bbf0167a3a46027d979e3fa8
z90443d09c3b6459c869adb4829ee51e286f5f8a9888dcbdf8dc843c5af04cd037fb170d7f8be82
zd42cec055621caf6dcd427973529492a536b6e5873df4b6e96749272a8827996ea59541a114497
za4da0532af558018dc87be7a13277853b9bb954c311dc876e637e94630015cca489cd585769990
z1f3aea2f74bda26cd3ecaad5c90c03615bf950b82d707fb1a6ef3f149fbfb745d545c9c5095804
z234aa7e82d8623e69429ea4d0c659e1385e79046e94a437d3067256a84c414556b0e9877d0b89e
z2888bd9f858d5a23f33db8a783a57081e9b2f71d9cdf14573feaf9328588ff56b7140cfef0cf7d
zd186e06cf8f251e13ef21d786282caa1f12607fb2d1dd51c4dd06c418f5c314d047f64327e49af
zd1cef8a4493426cd1aefd813b84030128e67b165f34aea697ac653ff71d9b8f6bad747adcfe8a2
z90f26194000804a755fb287ea03df5a3494f234e1b9080c47275085654ca9b4fccb6337de855ac
z3b58d1a03cf1330690d41eabdb1d3ecb1521bb0ca9df28877ebabf6bf5b761d8a96d8566ab7357
z4c80b6c2c84e36266b81e5ecb35a78df254f77d7125afe28b54cd3ecab03b848fab9f256ab0830
zc391b97729a5dd60344ee737da36688228cd20b39953797513f5314b2de8d4a16804c848bf92fe
zc98c70e0527a66bb30deec8fcec7b7e92ff430eb8b56039551635b852f9eda1f464dc781e019dd
z060ffe375b71f04bd2729ef10217b8f3ecab49dffbd3d07ac9b68c2341120c19992a14ddb944c4
z400e51443998b3c9efbf7b1e3fbd67c950f001eef1f08ede29ecde846229180dda2772f49134bb
z065fce4dcb33585f539923e8e14fcc8249e955e9e5f860057fb5df0ca4d8c416739e3e22644e3e
zcbd76c2da9daec1e2a724271e5d64f47cdc79f53e25240c818a8d0b37e62a3d34cbaf177bccf8a
z8ce0ed7b203898a3e45d06d75acb783d15decafb73c7f28716344073ea4d419fba7f2f08833fe8
z46dc861f78a63a7f8e8588936ac645e09baa31b09903ec3d05b617d69d32d25c51965f91a622a0
z77846c35dc7b725bc64e39df813895e008c410fe844016b59c34ad62d9cd0807bc00903b3fb404
z6ee25f1d4a136f231d0a3f3e1253104cf262895c31112361adac0e4b1f69147e1f5e95274e7bed
z52436c663fc4135f5f30b1c2b63190b6ce355d04b2f82f910a91c9d26700fd7f5d50402a1ed1d4
zc1cb71279a0820440845442c33d52d30d95b0c9664a3113e8b1f8592110ef56823ad8da53989bc
zb64cc58831880d16538541626e48a845a7196fe95d3b6c125ac688c4b874da3ca4123d58a2b9cd
z3299fe4dc3a8db0683f63807b2f60c8428d895f9d70b1c4cbb8ce3b7be9eba1b7bc797710dedcc
zca3d9c438b68ce38d8812480f7a7cb214881d8835133f2428b0cface5c52c9d8b22b1433e165b3
za3a548c67267950a342edaf4efa16f833ab1e8d1091aae4bcf2dbe2677c629925f18404f454366
z5cc5d3a5fb5884bf89cb0e4486e70d8bea632c49124bace2a688cd563d360c4ed5f17ee00bb5b1
zb5501b4f1dfe2657a84c6240949df34f317a81f9f45e1f2a70b81e5aec6ab8d08d4db513f10ee9
z549da36e9615dacf61abb116058a19efea2d95a8af1cbbd11229fe953fa7e59d8d03f3f6772ad5
z683bd830438802ef87af398381371d4c3e0159ba7e64a72140990bc2dc1acad6cbb873aceb504b
z416c921ff9ac02b21881e4fd65d05a9dc4a8a973946d275e30753781353de678c79b40b291c300
z3d7af4ba98136b4f204f33d24d1e5cbda394d33fe70860af7729bae9394a5ebbe0383fd06be6af
z539af2c9751733c1f66513cf9e92fe1d3166e4da41af271d7972c3fed6d33e4801242f917a0dc5
z1962e08e95118db19a7481b736fbdb4c9fd3078467f7bbe1c2df8fb2f8b80fb153235a02e7cbf5
z32b3ac2d08d9da3df2773c7d874ec86773424e4474097bfb4598d51c292885eb0d1078e753b6fc
z6cbb71f36107ad659e9c05c74919331ee05701a05f6133a5d7c97a5b1d069c29843102bd00a910
z7ee7016796b429e2fc0bace67a83f3a97489dd7940dfb7bbff78e8aaef3617e7b28e2248b6c070
z4ff19c5b45f387c662fb5fbbd47c3bcffa7a07289f3335bd0ff3c1da55776952ec3b170490e923
zfe94a4e47d20b9d7120f2847d7a4e924f4bf719866c10dbd044dd0c44874cc14c35e5ca4a766ca
zf6a5e289ee0b3fb3103e57f59e3ada38744823ed02791d2a5732052b90c37a37959b660ef47508
ze9b516e717135711cd2be543f56b59bdff1e0ff9323632d325a0d3444759bf0913560a68871502
z9ec2cffb3280cc873042c963e56fb385ac5d3778929d07bcb6c82e05717310ffffcf41db97fe7a
z924901c05a7415244339c5c720fd4b491dcfd3202313ae820966cf675470ebba355285c0807a6d
zb72eb2ba5f32c5e2a401516e9b58d73883572d751951e815180452ad24220af53c96af28b2d41a
zfe610e315b4ca60c87b576d0989bfa09b025858f925d10e1afe345c38ecae5fe2dcbbc42575fe4
z5c799403dee8e7c14feb98d6e9ac476ef14f1061ae0a0976e0220d836b9a056d964e8fbc76d6d3
z433090d4778a7cf40a62c915fe36e67194629e816e530a9ea2f5baeaf1fa133ee35fe8b713c998
z6e53ade1171151537e1319d5727514ed1799fb58d7bc3a7437c4d541f59072d43d8dec7a13a6e9
zb229c913c9a8d47c5b64224b4adbb40385ea42407e473332249195abe3d9b9ad9ca260a6aea1fe
z13c9e8182a43091633142e4b120900f82feb371923b6160323ca520fe657066b03ced81416f696
z4e2926e1ede866b077694760ac71ed0a7b909274c4e8f7af93530c81aacc6a5085ec29cc16676e
z0c06e02adf310d8ff698bcbd24882c7c596a8fc468184ed43a6447694e3063e563c9c31dbff202
za22a4e72865fbe22f48a309296d931478d4cc7ffae8b91a51fc032395f97121bee97c15483717f
z6031d2399e1d21394a7916385789a99c149ead24efda95e16640e0bbcec12a300e435847709860
z2463439febbbdda1aa72c952bc332a7766428ece052547b85a00ddb25743240083d230bac49e87
zaeffe975505755dad4030fab61ddea871414c1f1fd57bfad5fab5b7d2d4d7d6432f7eebfe829a4
zfa086c7952b87cf798149ef1f229e5f0a9e4032ff6d1197e17bf1c4f5982b1379aef9a1fd0421d
z304e03eac5b5e000b1d24495c95ca47cf0529294aa0b24c9b921ae8181ee303e09bca65ea92dc3
zed9f00c47fb55139926e9110b071eef0fe88131948473616deed147612efe178f1d4604d09a62d
zb51e854a96604d249be50c20d411875601898dd5b9def0e90401d09dbaa544f5564328124e8b72
z31b877536bbf86aebc48da22f17d67f9d573d982db79c5819a5060f99bfcf628b7413b40852af8
zd92ee927b450c5b83814d5dcaabd5cc2bf4d079220581dce11644fc315eac511334631a71dc3d8
z09a5220368641581deaa32d6e65c24d0db649e8a1ca3d3befade200d120b2c72fbb9ab20a02b12
z350feeb9a591289bacab0ed356ec7dff6daae58726bcce36ada203dff840bb8c89f92052fbb432
z95adf0460a34e6b2eea15b9399c6f89e940dcf30e5db137939e76dff1b57eae96d4ba6b32273b2
zd7a600668df02117baef1dbc0f5db90f50b11ffbf91b6d75f36374fa9ddadc54fef7a01eaad165
zf1f5042aa9aff3e5c2f400457d9e77e2616f55ab90c0e31f228b135463355fefe3a2c108b521b8
z3795a8b3cf3a8bd24943d65e35f5b4c47f333ca5e9b774ee76ae9eedbaab479d23e03795b5a438
z11e7f7bd23ee2bdd900904231f44b58b594c95ff2172e26ac0b4edf1feebcf5b28c10e96bcf3cf
z8132d660f187746f350fb16bc7e1db9ede08dc2c3395d59895b55be8b17c782013035f6b98b2f8
zc63e28c756a30ebcc44ddef5e3f66c37ea74a15a2185f38a78acb59d2e40c5aff5b3e7a0df537c
z8057daa5470a5580a86a4d3a0babe78cd8a72707a8d516b371aebdac9b05cea6375f8892f1c91c
z55dcea31049fa888cb424ca17342ccfb987d25b1be78f006bb489cd38e7af98441a3cda10b0272
zfbcc79fbc12a2de4ce45931c84648ea109b40afa6ad4574a94b3b8404d3e8650f2e562999ca9f9
zd7041a9e1fcc9c625664d665a632ce15c92fad0f00548c4c161345644ea98c915f754c36451fdd
zf0ad91e4acfad178b519b3b56a51939f94e73b00373184c1d5a79fd94f4adc1e8d53c7d50268cb
z15754ed27ef8ae005a0e98e1dd1f41e2002a1cf4805a2276c91ccd0fc88fdd9590d7da531b0fb0
z1d6c7bf2cd367a5b607984907b7af43ec1ba5c73758e33c9286105387bbb2cbf37bf138ef391b2
z2b56422f92dbc71cdf579899079845a6f95b50e9eb0cb98559a575e4763f143ee56b54b6383bdf
z2381b5f40c50364a4e8d1022fcd96339a591b3eb4e1802b659d10a8cde9e561912d9d521b4ead9
z548e6b15d20dfbce37af99b8ec443c3172b6b85b8d32e0d9b688570eefdb292d12ff0c8b5fc4ac
ze63f84bb2c0dc413a0f62dbe85158ea1e5675720906d980da1843e2332dfe29c21b0d25ffb2098
z39040caa6025e8255bd29f4973d875a7055bd9d980e39ab9a9f60e9441a3c44217a2007122b5a5
za5ba81b575f350a736e4bf2724a1c701315ba0bd6cf40866a3cc8fb7a45bb136e199c6b0961f0c
zd19694d87076cbf8414a711568e3bf4557a07e4328168c8d26baa53d709eff833f549177b3a54e
z9681db9c845e4c5436e982fb063d33f9153c7e3fbf00380e25b30f66cb795be937314759f1a863
zabc5cfd270dd88c83cee3d1f716ba4fe6025b0f5fee9bb74748146c5e4b910221d45e95b359cbb
zf84837c4c320f43931743ba67e81d95ead816ab132c8b2492610814663dc5e7abe3cb5df454a4a
z58a5d2d1e8d0fda68867090c0be86cacf0edee1c7c5cd68c9d23ddd013a040251ea6f775ff861e
zfb86ff1ec67ca3af99babc909b3be6581a8f6b8268caffbebbae2099b0a46b1c384fb91ef66c90
z423dfbf4f00909f7391c96eee92349b133209bd760acde11bc0c39a0e081bd5aa225b94dadf341
za78e7e861edb66e20f704012f35d6e642ce1a97971f3cb1af5f5cff938a8e552d973d709046449
z1555d680231bf5d29e98242918aa213a2c11006fb3625a75cff873ee749a426c32dbdf1e76bffc
za81a1ecab694ad7d780bcff6cd0e28e7bc06960d1a247fea8f76c9a6c1299d599139aa75664150
z86e86740632adae037a15537c6ead91afab0301f0c0b3f2243f866c227f574d324191de7d1fdfc
z59b59bc86eae965007bbe7006ac875d64330ce594d9d130a159992ccc55e8a1324f36a4f1531f1
zcf5890a76bf3eccd9f76be00b64895d6ce4da25f81ce6787ca6260bd644977ee5903c707571230
z14c013d801321695970f25ddeb1dd6cb487a4444f2fd84bd6c0b749c92e97f5bb15fbe52e345b3
z1bd052fcc801310c0439db4ae4cdd80376c953cd1c62f1c14824b69daaf42aaac3e6b53d288d90
zb4b72eb97880efeeb364f84d9ef280efd2b7becbaa704b6bae03ab07f60088cfb42316c4feef5c
z07be007e5a652b4bae62e1a4e04c8cbc35de721017927c1826626fdc1ebf22122af4025361a586
z056908846af33f293279a37852e659412a5e15e16807a0cec01304733b8029922d299c3cd5f9c3
ze806db03d3ff5a6a7a65a05cbf7f2cc80fd8a6df60f061035ed515d4b8cb66da0dc11c1b1e70c0
zbde5da9e1d6bf61e29a70886f055bd43c2a40c5f70b541592b03498b78249d6d5acb9231495ca6
z71b8b9609d16c7c02e802eefde13b34daf9c4299845eb245e94257222e8eea1edfe42b96695179
z1b48466466443a680423aeee1fd3e1ca321101f6a34c3266aa9428e3c26ee4631f567a02d88779
z1a8320214b0853b9127a4890b202dae3950b6730956b04dddb58e69896395a8313b5bdaa655da1
z9a501a1b5345ad7097295deeb1475d92a07c7f411ed948a8aba17587743afe0ebb3308c64d6bb1
z8d57be889a63058914af4388a71cbddaa243695d88f0c6f95ba6c847ce875f97b226743f6553a0
zd9b66a5a217ba364ab9b2360b88c45a10870c449276f2e5e766556d363c988bfff3ae0efa52371
zab0e2999bfb5f6a04f3dc06f85e9f80e82b8d4b109438d54ab38cf87493da8ac518660508d4a4a
z25882af5f150174f5e4610746a7031a3d5c9a0c80b8d372b3a1881dbfe7bd01b7e30b28ff49be8
zf556202e6f5ba06b8abb9f1f28adc14f36a1b0db5e54252bec2f3f5b2cf93a0ccc94bad272a939
z948b6c7054d8bfac5cfc55dd5dd8212852ad915b40ce9face093fc66dd16cae54193634490e424
z1607c639c0f645d20a544630a511b95f485382c9dc9c0c01693eea37446443a1c8043dd8bdfc3f
z6ab066e1201f2530400c36f5530ca29d04f4555282f5a2ff616d0d4a8f079a0aef74c4309a8e89
z6e69bcee66ebc931870f84f441fb0743251befff12c783318b6513836a4363069f29074e48562f
zeb4af4b0e2d76366cc4115e271abcae98d4f2666f6ef2fd0ddf8bc5dc54b1fcfef0ae8c1e33cbc
z57b0ce252e3e1eeb1759b8940dc1875fed676b127b09d01807138f60c73acf8faeca932636c3e6
z09e974b32f33c9ade4e125568b257582750b0574ec9f83e9f57a4001270de940d19c3ca39030ae
z48c8fe898af3ec4759b65cfa83bba4e4a32ec477526285dbaf787523b27cbc74f74b17fc06c6ed
z0ddcbe64d80b67610fe0c16b2e42013cc79c2f55740b285d8f0374582d340bfb191aa8620b849f
z99585bda0e4e1ea4abe5d0d1d8ad76f13135f7cb4c433dcedbb8d88f826738d202edb681620c1f
zbc710b633c59db838582dc888de1aceb7d8eb2e209da2ad7c8791e2eb9f89d9c1dec9847ed0719
z674416cb60b898bc488bf3a94df588fbe8de6c379162d07446dce2547cb2522dcb8b7e4538d9ba
zfa77f968f6e05f00c564ca9b56310b593b29a2b890957f15ae45d521aaddfd17ce4c57b59b809d
z61e384054af669b34513f90799b6e1287ee772e8eec973057df403334d3b6918e1702aa7c736fd
ze305faf3d192c3209cd0a2077d05b4d79872a64566d0dc5d45ccf7cd8228d30aba02a3d80bbc74
z07845b164cfed084f085b9c5d10ab0565cf422745b96ff699f93ac492c227315dd6e63f7819553
z6aae8905d4810278fcaca32cce7eb6403031e150950c0faa025b90c00b3ee73326a4b4783a2afd
z8997a209a6795ce2f50731228ca965702a40a9c269a6c20e05144843e7efe006f9288974075183
zc9f7667a28dd071c7bed87dc9fc34a32315b1b9581789a4ab0cd26250dc975018935cd7d62398b
zc41b38adef1e5d9f7d16bb2a0b93e71eb0e69c89f9c5d54e76933ad25ee9eaddd3200911524468
z0c7076187441e0e5bbda9ef7b0059f2b775adfa16f563dda84dbf206d1e934e36c15c7068b2f98
z0ab17db5288384fdfbaed37ae8d7a97e3cc56441078f63baa0036de00588e891cbf08df39024d0
z76e1117b35120cf5613f619dc270cb1f4d93f7ed2f1a21c31d6a814f95120cf391c224a7251754
z61c4245d9fa1e17e3413febf914e5115d1c816b767c230139c7f980b2c0461080e97173158a58b
zcdf5c60c44fe20258e5e82a77018c004ab0131c4eae4af8c6cbdb88606e5ef9cb40b017f1f59a6
zbd1419b53160bd2347c7367351b6608f041bffb62f35b21ad6cdd8228cbc7f40d31ff5afaae10a
z44ee9a97caaa80c9b42539e0f3b9de820c7a1adf96ce17624b0362b62da58d12147b6be3ca7d99
zac07729f5c15ece6f326d107f7ffd976b034d1271c745adf5dc2b446640c893ffe9793c9438790
zd82a00f58ff617c7e27db5996b9f7abbc1235eb7a70db3a3460daada86eec9825f40b907c85de7
z65db7e5ea82639a7e8bdd8a15c06a94106baf7b2f8a1770a6c4db471512a771ec801689ece574e
z52ee5042e4c941b91979c2f0a44c2202af0ac36403ee1c2369f95aa55709e6a7734b3f6856f117
z888859ed510026c5dfef134bda43872a6a8bd60b415c10effb7c87f61ec47fa6e726756d57c528
za3c1fa822ab9efc5903e0ed4bb6aae2ef020291c4f40700233ef1bb751be1f5d95b6f54eb74abb
z1848c9899ca052287c94b04ae017183dfa24563715ead7b03e01a61d3afcb5fbe1c32daba3158d
z5546106edc1458b1062bed424a06c7b1f923aa54515a3dbea1cafbc4df42556788dc868a69e8e2
za648fc567750b36ae3b9275905f3fa432e98f994412b441a0eba59f5ec7e7b3847008cef7a15f1
z643d12a9e0b71c9f45845c25182425e82ab4315bcd48254f2891bff17043246d4874891a317d42
zdd7fef5ec7990b691a548cac0da3febd6a15adda345b3f50f63b1965182e46fac8e334e956edc1
z3b84880e702ca35fc27b32cad926819d271269c50986625b92e5537e5a4101b933d99a0741c339
z1a92d7f6d2d6279ff524dd8a691520247e5d1757794c0e22f95c4037273b23708bb8e47f1721ab
zb29858f9bb13bfae88bf75034b3d60d987abc800d6435a7664c58a623dd6e9e85b5e58a8c8c8be
z5335a6c310d6d212f9550fb201215b101471bb496a2ed5868fd2483364750cba17b4be7aa64937
z57092c128960b76ffd7fc9a97a6227314ea028a9f9904c1ea71b0b8f25737524c2174d70b12ceb
zc1fb662b65d25b7af2714fbfa862bdf29739159f0781aecb433bcc3fcfd162d86d0c1e276e9b51
zddca2cbba0793d449b7a7b45dd78f5b3668ae093fc3b9e645d0f22b01e0816af21a432ce19108b
z9eaa4b3847553059f0d181ba320d9eda85571b72a943e5ffa1bd466af4e0f0ef194c0e7f5f8b23
zaf0c0ed65a773644ece95dd903080606d676e2071cf48b834f780b097b27697c2d65c602987fe2
zd3d051427fa0ae6535f10a4534c664520e7e26fde7cfe205801893e68267936e7acbe6febb448f
z7d90661848f193a9cd7ba302b885ccfa7ad03058ee537c91be304a88f1387d51c3baf0165b92ef
z9b8b0cd10505721b682e73d657cf50dcf95416ba9516a8101367e1de918302124128e3c1d75855
z42a99b4553062227b193b4cef58e44d5b2a8d457683f9067fcff9425c912d950f0589048f71fcb
zb18970ef12f7189c64ac68dd26bf56e959bc1aacdfa11e0f11627a643aaea67952ac623f080f26
z2c87df81248a56d2f1462119052cbb603cc7584e49bd15dfa8cf9252dfdcc548e37bcc97a919ed
z9f810efa6276af5b58cd7258c62114de07467efaf66b89b182186ba54691421fbb4e1bb43c8a40
z080f203de79cb199e129d551e9b58fdd101d151c1c4fb721955857794d2838d59baabcf5b88789
z2f8906c6041b0246b061b7f0bdef831616a35fe7789687aac858fdbf01fece942c70fc9fa50127
zfe9a32186ccbae0bf32197c24bb5d8d6825a06aac26ab13989ff5d1b778b30617d78e369f68952
zf011da7020e7af983937423a213630a56ad08902e53d95ec212c6587098ede4fa0ec568b5e46b4
z5a50f8db083a50d2fa127e35808f90bbd4fc5084d585549313377c328c0245471902cf463d499b
z35fdeac7574db31edf2f18600a9ad0ebf39e3e8592426e6ce11f2c425340a1e68dca5106ec4931
zd33b9024144010149ace67c5eed80890a66b9184cbb46725fa97b547430b9995384300544b0f0e
z280f6dd8618aa500e1c6f06b7487b99eac4bc3482cd0c5637cba5b82b523ea1763e0455059179b
z3d6e453aa0ecad3d90a2894b1a91f3f22474014cfe17fe08552b501f28193d8e252c431f45d181
z60b6a75b353de12ba7e020380b19a1a5240cd7b542824ddc256410506e8a9d2968a68fe7608659
z4aa957a50443d9dc980d1eb91d76065ce2d4c1bc59c8e9be94ef4ba0e896f5c5e24f76a3f9fcde
z38d173c35bf842e6a23b662ad9b1d688669af7d659cc88bb9047d6098e4463f4672036edaa189b
z0e326fc0c87e367fbbdce69dedaadc233db0cad0a7158e7eb6a3b63456ce58cbe7ecda99a2f068
zdaaa33fdab91cb321d0dce633ddb98bb7a0bde00f100884b3fb178f96eccbc3f0de988d598ea17
ze024c689916128ee948921470f09a59cdbfd55818166797b64610dd90a46b66a94450281e19125
zfeefeba6b9c04e0128f13a57a61a8b5e84f2e17989c822ac3b69b82cfa3950f0c67ed2d1614664
z18ff8f29ea9b83a6040ec7dc4aa93633a35a61950eee6f951a136cce2d895c837187299faa0aa0
z15eb103a0a225308b5e61ad3a9eed8b0c20316143522eacee34abae027c178f05e9056af6eb7c4
zbfa85d9c16262c82756aa399fe5ffdc6e2f953fc430c0f5d20905b2a6ced4106cd0e3f41e1aa04
z95c224f355a466ad1d8913fd2f9977d60478ed7d788228222d87d9f0328868ed8c3bdbf99e630a
z9b45e30d69c250d12f63f038b4ddbea3b6a995a96e665339d521e8112c7abd789d9707298ffbd0
zf7d793be030689f1eb3e6057f0d59169a74b7f7ce108b95e357831aa2f01e4b823acab8608b5e5
zf9b564df01cf59a567d9046616d7eef00183d5823974cc820b9aec501120b0de4a79b97b9f2008
zf24245ce73d1235d84bb17c480c7d90872ea7f4d184e126a9cd88884830aac54d70331f1200b60
z12de03114683be2d756fbbcf9245ae4b6a57363584aba5a98e390e4698bd3c9d01432089528077
za15056b0007e5b479771fbccaab30075e36b548b776f7226a87efb128c50b02f9bc9a935b89aa1
z30b5d3246463bfb1f94638598f97630667f28899cd4c22c59d34f6908335c3c5fb64f15a627b19
zce926b67effb8791d6857c07cda313f055de107deaada4d6ee4f37d1774122c460a5a2ee74cf7d
z0935905dfc587dabafd4aa468718b09ee066deab74376779db8c92ff06e31de232055ada3f0b08
za4e5cbe121c2a8cdeaeeb956f9c275a33884e2399c6f4f34a7b903ae41dce86229770a3cbe23ac
zd5263ccc879c9aeb6b6528e2c896c8b03d19c9ccc9c2f139b3fe55bcf6e457c0ee5bdefd1d0788
z20b7b66a1940a7035c4d20ea3f6bd14f3d10efbddb830ca1cbed5a90f5a9fa504b7a6345f5ec99
z1e0f2e6e7d282661541e5c88839ebd28738774d6688b275faeb39fdb70ad9d308a5ad687dad699
z2a7854895af35b6a11863d04d152d76b3737ebbb80bafaa32b3c8c0fdf0f152d42d94489c6ce86
z8f994406525ef0f4fe5296c12d41a27788a31ee031113f43602290ab50cbbee5718cba15fdc749
z830048c887b908cdf429d020e3023a70cf007b83f241c800c07fb8039174c21f0548b32463033f
z7c33e34918e92b7d422e9e885384ad819c3c49207c5104b0f158208c7d7d56e796fd070a9f8008
z9e46cb059ec857906ed0fae7d625775ff33f0a0d7c0fd6bbc982c61321b14b6ddb47acabd09dce
zf0794e426d94b646feeb6fe84870d111cfb83ed687d00d2a4140695751c0f36f4c496329c9bba1
ze139610a3c68357367b5f6d4d911909b35f524c6919fc0e991155d0e32aa65f88837cfd71bf2e9
z9cad467451a71de7ab4c8f0e8d4639840dc56a9660ad55a76e315ba751d37bd4ada638f569b4f0
z1ea83aba41fa34bdccb95f8eeeb4f590aca1122f4e6577993252ec07f6eaf22ed1a775233248c3
zf209e50fa2ecab8b93b59c2200a25154341768424cfc06186258fb0a266c60ffa006903c3c7995
zeffe427517adcffccda998d6db99cf1bc4cb9e8028d3b57dfde0850e89cda518bb362b90a86703
z76827c8a70d271b4e487c0b3e9c00d5d5c408beb89e9be217b6eb3587799fa074166f5229d3484
z760713cc2f89e2cef5bdfadbaa5282990cf1ebd3e7dfb5ee5361bda8137016fa1e8a65aa7d83fc
z7ba0bf31c3fed826402d4c2524bbb44101fab97e284a412e4a927cc20b7e6fb1dd155c48c347f0
z98655d3b66719a7e9dd6127001702f76ed348a53a851d4f6dd6b2902a056b7fee5f88dc1fe9197
z6bd21025d1fff303e9908c8de18f1fb68358677d84eba8770db19c0ee3baf7585c99fe15f56f8d
za3d3b9c64309f4014ea089e889cde81db5c3cef3649e8ccbab1bfd1c4160904cd43687f82e0dc3
z016ede544caa12fae807665362b130d85de94bd7c63765cb1d54ca259d23c213b1216c65a1775c
z940ac403ef6c7a6a3ff9366bc5fdbe0f694172c44d3f35ba156a95f4a6bcb92097dc426fc5c842
z3faa4b6f1a03e0633e195ba26101e601ddbb197b677759e5f5f901d0afc583916710141cdd135a
zf3d2a6566a86bcb8a45bfcad2f1fd659cadc7ae2f161ebe1ea9b72233399eaa5f8df5fab8b3d2f
zdf923685ec28020fbd357a8db4960d41352c08f0e620d4fba76720e4d93a54ba68f1a32f77577c
zdf0041aaec7ab539be8ef09c6d5a7acaea9ed76798fcb1194eca1bb47495c9bb79321ccb2fa365
z7bca1633c804864d57c75f86ae01076bf5742274510ee11a7f4f9ae963e32a2cc703e2dab6207b
zdbaae49e36671cfa253f4df194b921c9abb32e2f5baeafe969121ee48321f3c1cafdb372fa12ff
z210e122aa7ea40d7abaaf34e36d612a86abeb79c9ecd5c98c0fa4606edc60efda087d4f95d9e97
z642b574f7285520552284c53deb677262e5b74f9bf63779002a651d4c2a8c958a8d5f3dd39c86d
z9c5c864395fd5f300973a121654adde57faf837f5d3a6d9dea6d61b4c7de631b698ee4ac720869
z7ce522dcf66ddafbfe5fffe6d456e2397097b66d8106bcb9521da4f03950bf0314b43e36288453
ze95feb3f83dc07738490768e551b6f6478daa2aa09c1d507627d2c1d11136382b991b5330b001e
z7934facbf6f41b5105b7d85ff44556f42d4cc14bc1f763ce622dac6188d46803946ce76a94ab12
ze8f14cc44559875ddb9b2591825bdd8b727eb0d2269bab227bb6ea0d54265054963e28ff119374
z58e2f7ae42fef1529791afe3c52757bea5f3678e06494326f0c4612b6fbf1d2d9ffc574bc66486
zdd57c075aa06d77dace0ff304c25d01290071d6bb0273347d2e63467ad099ebcdae03f79dce06b
zb0c389a38a9f7edc2d7ee2d05a4395fc2474a31c93f201f793b765edcecee96963464bc0a7caa9
z66c052d3e95d3a78012e2f31a20a55ecadb048cd037635ecaf05339a42cdd5c4a543d8750dcd36
zd85ea0391f061d595febefe41f03747ae20cea212256873a8bf8339df1183dae0718555bb99618
zd783bb0296e721494daa224f46c1bf2c4bf2fc40f8460f07f5242e9c1e4e0fd28ee9b9fbed9e1e
z7cd04512006b296edd3ba64f152cefa7591ea6f1accb9500dd33a033cf1b401bfc7e1723329cfc
z656d8a702dfd947c0d0cdbac1c8178fbd2aa7b7416c558631db4b2811ebce0af2337befef16010
zc0eecc5938499a4379227f53e2809129f75c9ff6e05ab212cc28bb48a0d62d0a8d815a3b5657f0
z8f124680acfcfd0e795fdd8f7cf9f30720fa2fc625a8e52e0786aab2d206f35417e4d1a6ca6822
z886493b453052773254c50acbe123068c13c776fd5747c99ec15ca621d8fa1e8c391ce1e2c453e
z1c230e48151aa6a7e2f28630e453d10c0bc2f46c672858f44f6345c0636a8aaa870bfe970ee457
z74d293645c18c9fc8a56e695e5bae4033fd174dffa758eaea016a072e223122ec8cdbdb80309b4
z079506f3f78247db1fe205b3a1efaa2bf2bc361ff38de56b00458dd3052b7d5825444ffd613be7
ze50a331714866ec78630470ae8cdcf3b8b701d9ab587feb9dffa16783be7df5f1c8a6c683327ec
z94de95e0a38132abc8fa4215be3a0e23beac13b8922ebefb66e5d65ccbe1c2d22e20aca1fd66e9
z9181858206e0aedf34f1e1dd04911f386d6cf02194671d4d199bfb8860dbd6d5e6bd6e941748b4
z127cafa28329ecf5d090a02b9db8eb2032e0ee5d4f16418372b218667e748d25eebd040bde8231
z42d4d00cde89d1a1c5dd4000eaa64d32761f97f8a765df45bce7369ac884bffbb3df1b00f2b622
z284e11453e6e8d18e4ff36d00c3539d81b54447bc81cb219a9b6fddc92b82ef8e5c4063df5e2a2
z4fcca3cc1e7341f6c008846d05413e65a264057c14aa9ea505d292f474859c86d207f389a97aa7
zc7d6f262c9ff7556c20a8431b9c277d27a14bd42aa447970d276aa8b301f6c534f3da611e174f6
z280b518ae4f0caa99fe490540a424137f1b12b1e31ece3afb72f75644051510fdf61548b22ca45
zbf441815cdb8e6b04147d15ceac0434b5a663cf4c4294baf8bcc3231a08f06e2cada8ec8ad6c64
z20a6e124292114c3626ed2c73ebdd95d4b13a06889d98805e37df52fa86fe077274108
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_amba_axi_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
