`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff98478405cb2c034d92a13b05dd6952355a8276837fe1ec
z31ed579935d1f03c8aed1f61cb6f74edabb0b099810d7bc07560d8599c00d4ed4049381a6e2b8d
z86a7f6abb625239b7bba7d5cbfc5666e6b305ffb196abdc98f050cd1496e9e7a9b8bd29150791e
z328fa776ec981c1023a4a6b0b906d92b5cac1c55b6298044a221652eeef177a4db4a9be3aef948
z0d5197faa7d81d340a91df6af7cc47464ac47ad744afe8d7955f53a20d7dc2c70b870de3c49109
zbd37bdf88bd89d4c520013049826a5ae443afc225d5378dd93426f04e28efa6e0f8de08f960ee6
z349b2eefc11b1e051caccfb9523ea03bbf7871b77b6315eea8043e758ac80a6cceda9f70ce31c9
z29c16f1142785f52bff8cf2223c113ba95c30633fb1158cfd0b2731d8349c93151aaa2659c6d4b
z36f2176f6ea50ecb06e3553100ece565e4459df0eccf14c18413cc057195c25bd29da5459c3f4e
zd2c990e5c5add741e799a788b33f495df88d1b2f3d1ba83bb4f22721e4b9f7597f027652c1005a
zb1603f1c5d02c094c412f98caa1ad2ddad9baa87dce839c7267d16510e2d9563daabc3967e0f43
zd6da55840f2ab40409dc4c26f894843e3ee4fd3025033db5da70eedea0d16611aaf71e0a08793b
z670176909010c72591fffecde8a5b87174bc9317dad63d4b9520bb01fa36672965213c580e9ca0
z5716517ccaf0f44984e97ca40155267a39135c0b7406d0e79918ca5a3a8c45010b24a0dca4d54e
z8dbe866ca1295456fb61c8d152e50e2418d8461191c361c236af2f04155a4fc3dbbfbc722eb814
z91606681e1990432e610873d88de53a4600c08de9f20f6343c8c2bf154fcd9b8f7a8b409c78c97
za3e6da6a6beb0f551d4daa4183c12c868dc24d987da0a3051b596d75c6a463f2afd18e244f160f
zf86810a2279c4f6ac80e62ba627f4437cebb5978d1a898fb79a942113e4683dfd7a4b194897e77
z3aa434fd4ce56057929883adc256e532e06aefaebacbe2f2768eb6c69fbc1e6bb74f8e77bfd415
z4e2c4f1d12e497ca04e0e5f03e56f5cb4a9479f0e7cc01abe46238da61be0c3d40ba8d7e573795
zc6460e23658ff3e77c2a082d2f479bc512d12ef6ee32a2eaa5c825d1316e64edc6b225510bd9ae
zc57777be48cecac370d2d38d33511fc545df4ba376ce064589d42f81927f99ced4b6f2d2645e81
z951be29ba2c245f6ca059a224ea1feb94074f44351b79c7962b342a95bd101196d7a1fe3eb3ac3
z47e0ccff0d86a450e6191bc683d639dec8d476390c079102559d89a91cde20d9f9da17fdff44b0
z0aac538cd236b0fa52683b23ed1659326fa738d09ea248443f35b9ecd6ef475dd11968904c7947
z20e296c123915b962ef72fac74af6a75d5cbd21a4f75a535681ad2538a80a7fb70846962fc5c1b
zcf0d4912aab44e04cbac31f3a8065e7d9e30c0a128305a062f827d080c9853e6dc7b559dd04518
za134f2e47899b6e1295b859119ca93af08e93102df8252dfda482b50cd848c2370d1686c9b9165
z9787003354e779610a2ba208d8c9a4cfd937183a740e30fd7139c73fa66d585db7e61e062e9852
z6101bba552b8c66dacc3a845627b37ea91d63f732e61997918b8954bfcdf0e6b68287db9231a8c
zdc824dfe7cd196aafbfc307d393537a990c2c8e1d01741feb86bbc74243c6fbce7dc4dfff844d4
z232608e13fc5c160b027a8ffeb194608436c5416a6da33a28d7afe201f5596c5e35935b4db3b26
z176f0269559f23c51a63299c545cc00723f31b4560220719e4d979c43c40d4884189428a4e6922
z63643a01005283f14d31b6b0f712401fa3e522fb8decb30c97f5005c03b4cc9a658741b5f1f1dc
z33e9ddd082758a0e600a682d9467bdeb5576e255eac982f9bd92fe300641f09347c7f562098189
z3e06364f1e2b890ca85c6ff25e7772a473763598f4d5022f33bc5e940efb82dfb60fb2c4435dd1
zacf1ae8c0b1d3f87552cf4d486c04f5b58fad9b518c6e01ffa6bacbf3b321f830c54009fbfcf90
z3bc79c17161d8c3b67b626dbc33a9a5de5399118760de6c6caf63c2f853180a4214404f807ff62
z14e7a89a2a4c51b21ceb6038e6b6c30d1cd01cd2cc41cc8adcbf1a242d528c8e5d207a67cbee35
ze33abbb60633c3982536cc6d7c9e77133a0dadfbd8c504eb5c77a1036d8c6728ba1e8688352ddb
z76c5aecd84b9fa0cbe4aadb5edb8cc84de066191205ccf5624126fe8c04937ab83a8ac8be061fd
ze4435aec3154b88b4aacb40965488454d4ca7a1a4efab5f1967c6b5bf74bc3af93c274343030ae
zc9f505f3055e8273696915a531204eab556bb61644d9a420f8607b2a5667eaec1a299cea49d6c8
z4c777c94ff3198e799e199fafbb7c2bbd2e26c2f9e6d1b3dfe91a3cf821433337f0e89912bbd93
zbb6a8d492ea956c988dbc0124b944a24d5582be0cd6971ba2a6aacfc15d9afbeaeae5177db2aa7
zf72b3b3341b4f594799993e5dcc1fc92d842bc31a6529e0ee2383fa7a0eeedb186c2ea5ee1aa4a
z05077fec5b22afc490d3d23de3ae335e05967fabd92c71239c57f8e90f6e06ae4f3e9088f724ab
z2dee1d7ded3c4cc2a91d3bfd79d6ba02a6c727364e7db4ffa9e506b0b1db1b0e8fe52b269b340b
zbb91cc15dcb6a9650a48492ef08fbe860277669443f833eb9399b13b881a764c8e80e5af773911
zccceb6a065b2661b1ddd4f7133aee81c52fb0cfc330135d941e42e8a4240dc3b3e1a08f34f2d3f
z629203121aefa3d565a63f731a2bc174a5903d0dd9719c8a9a183419ae9ba0e1cb4ba9bf2cc2d0
zba1547cf960c7939ee64b248feacaf6690156335450b58ab6fd17d141b07ae58f8c1a9da7ce614
z7c3b7df86b87fff422b7ebd4b9e8b2f89ed9bc83d913ff23a3f2134205dac7461f6f6aa1801247
z5eae1345726e1c650ca8fdf24c42313c294caadc64a129802f74bae75ca42cb1b97922070efd6c
z216b1c5ab724a6f9ba1ab1097d726d2886fd9c992c77be2d8573736e274f9936ebb3dedcfc7416
z9936d286130c4ffa788823913d8df1cafefdd503d94b7ec14d9a7c86059782678895e7ed92b3c1
z3df69cfc124102099aa67589efc841b3874a83a32200c240872ebbc6a58329cc4177d8b810a0a2
z1168bb7bf0c7bed7e2516be6e7922ee6b7d715d66be8d127336fea76d5f334005f9cd141a38add
z0eb7e3248b555b576daccaf8b4c6bf21e2f5057808e4665921cf45a2854b587e8e8640e58e4525
z55c5bb12a52b71912e50bb1c5feddc898e5bac9922df7200314432829ecdff379cd98eb584bacf
z4410ed93f98b3618e0c7906cdf5714a46cf9db16a14efc735d999112e92aded2365792d147f5ee
z05ed04b671347d77467f57e7cf08285d30406ee06c72628e06fc22747466cdd5a9503e4d9b93c8
z5ae8e1cd3b6bd05e4f77901a98a860e7979012d3f3df2fec49d9de778d9e698496355fc5989fed
zadeba3efc01e0b71ed0ca41fa48e0079ce8a8c1ee6473d0af1c5fca01466be2d95948beb511393
zc81eda47bb12d295046772d87fc0ec78cc65a34f018f6fadbc02ec9c53a9f54ce0e0d84d2694e1
zae5e3dc1619359801b4f99e8d8fb750e244ed62252dbf7906c98fe82b44b03a3c6a5403d25ca77
zff3b4b902a56766b8cdea9be6d60b5a05e4052c980147b710517b4b5517bd2685f4cec4b64265a
zc9b88b4c248ce7c46b6883eacb507c0a924cb3fbdfcc768d6c4f7feddf8d5fbaabfa23c2150307
z8d0f2e5bbe6d0d9f00fb16232e9e50fa963ee2ac9584b296e206e919325603f4400a95410a2632
zb64da1ec16e7c98bde94d85df2ed82c03ff444f2042238f5bf3ddc90c919678b39a764623b45e9
ze890051488a9f7cfb4126d4a832b038eb0e35cced25ff55e1e527277d622c836ec53bcb8c256b4
z8a9d2faa1ad28e0ae4b48d02a9186119795e83c12178e4b2ed9ef7a83128d73bd5332bb318ba35
zfb80ae72f18ac46264649cddfca29d8aae14872b1fbd8f0df6b042aeb168b7a23fbe19c8db659e
z9283698ae63746bd8dffd033db188b5e19c8ebbb197b4b62544cbb9f598e3e31afd678dd8055eb
z17b866c3e67725f9142973799f591237109e4171ac6bea7426741c8031cd359224c48c9f5c3cc6
zd59d18b40921e824ae27ee8d370870df92e24307f8101c7774788fed2d0f016792614d0a84f18a
z062c6a5ba93292694a7fc7deedafd3284fb55b6af6df46be6483dbf2bab9060e968f8a4d923f4c
z77ef117d37c1c74cd485a4efb47a1b79f11fb2a1fbb2b34ae59c82e5f76d7a1f6d8eb159aec216
z61766908a52ff248fa3ea8b0188a79e81a335a126df7f664503718a3eac33607f58995a96e9a17
z30e48e55d41dc1490301ca1a02f2243dcf2bcd77e00a08220c9e84a47ced113de4ce76945cf868
zeaf1ae48e67a41ac7214cb38ad65538b612de8eccd6cd695e493524d81b04ee6a8e6fcd55f2450
zd7beff95d6c5d23aa589f32d274fd7c8ce48cab050d3856abe0fb135961fd3495c7f95b1849eab
zf2a97db0b594077ec38cc783fd62a82699c9252c85365d79de6cdaba98a18fd39568d013e423b9
zec68d9cbb85351e1f10a0d834c4ecce4eb5fba7ea05ca3362a6a479e268d703107344feb71807d
z411a3913fa07416580e6c5926ff3c0e8132b52859537d9c0761471f80ccb1be5a0253455086d52
ze383582e80aae3b1129a14aebbc76af1ee0e5ba7e9979e26b9c7521e14fb81f2067bcd5a921d22
z67bcc1878fbd9977b1aa01d310beb4a51a8ed327598c55a4fda6924a7e49c18bf6de59cbfb0493
zc83370e820d46bbe3715687eca861733d7a3b24ff65f36b3edbbbc1cbbc8361985b446e74f956d
z20b5dc200aaaab04defbb1cc18755782c68c45292b199255f0bb56f27a8ae727dd0513d5b58a18
zf90e2c0b4bd6b9e30e867bd45a45e71b471030b3fbc70867ad935ca54a601a34e3c2eaee5d80bf
zb916adefb5544c5624efda26e3b2b1764bd5c71ff8d761af637342aec2814e4356936a659e0b1a
za2e2448baec64c3cf1b93bd20e16677ec569ac53adb12379a627f71f74a991e90e3933cd80f207
zd3702c310afc058faeb7992a3498b6b2722828518cbb48addf73c2d9fd7162b20e0ab2bbcb5902
z74d1e246b651fc2c1ee0d6f1a4b00afda48fc31135c59b2fb5ca15b1ddb8bf2cda12f2fdc74a23
z60e0351260e252cdfbbc41a61d7b9f09684d434813fbc385dc65123cba9ef89ae9eacaf8863d06
z38f9fe8717c0aef2a666a368c3ab5b7eb36fb9b95ff5189f6aa420e7ba954c3d8dd3a21a342c3a
zfb89e6b31b97f404e52db51314bc915249cca74a886f39d25d1e93d48999e0889700e4d9553ba1
z8dd3f23879fb2277eda43f0f2287d539e7968aaedb122ce7a7246c0bd3c9a4334ea3fd3524c1f9
z6ccd3c474d6ce1377b88cd5790ef44a83b37a4ca4eb308afd276f91b2c1970301d3cb34d85ddcd
zc45dd54208a3e6fd5f536c46832b5c0d8d06e282b53c6ab9320cf54ff9b723c219f13df9d51fd9
z255b7a7a87b5aed80922c60aae3c2426794bc8ecc47c638cdce1e98348f8b4bf5627e727e109ff
za9674bcc792aef91ea57997a4f73ab24e0a740a5e06d09ba55221f0da51b6143fa97dc60681225
z00dfb4adfe836db3cb7aec6de50c8ac4dee6ddff19dda82ddd6a967cf657aa1206dc0d21e49121
z72415848c3ecd344d965de8985f1d4fb95b688477ac840aaaf4b0afdd955d9248af4e3ca7531ca
z7873c24fb3550fbdd9bd533007fed90774ff62fb73c261123180a4ebe9ae5888e5728d3e70440c
z1c011136cfbf919a52aa19fadcbdcfd49808087c93d4f4504c80cbdddca99bc8726ce8915b8df4
z9f2639e7cab103729a410365eeb6d8ad4ed1769fbf067dbdaee07911c990dd74e4fdfb6e58379c
zb35eac3eddaae63fd6c309e72b5f1eec16a61a2afd19910ac6d219ee5fa503eb642c0494bf9e4d
z6d33dd1afaf19c5155099f6d3a1bd33d51a58a6ce008bdf08b8cf50b691da05d265e368681e411
za6a0f344d619359ae47d1a8de09ab60104aa81dd46910017d52ed0c4bb3aa135cbf3689e508140
za1c97e5988f21793ae54c5aa866c867c1c12dbf5b9490ffb8c0b71e046931420c3efc87813ac04
zbe5d98b97d948cc57340d43d7664a7c744ac07395e05996b4e4b2ea1d8d9eb5613a523189c5efa
z9876319c596899f4d303496a6c6f3ae7f5fe5367c11faeedb963efa2827bfa59c5283b84d2447d
z72afe558d61b9a54284295d22aae38f62d6007b0c5bc749cf29b17f03a50e73533ff61863ca96c
z6fb4d682b7b4c278442c1e8aed4a4e78f97eb3b23ce36ead918b7428ba93539d636f12c57fcd5b
z0651b3ba3acad4589be224672c661fe272b84fd07eab9106bcd0a58019510aafd20d1800554248
zb63de89d0067bb3b2ceef84f781c985527b101c288bd5737b104626e3fe90d787c4b3b4e6116a6
z1bbfb3d94216b003ea7aca724ec8e76f1bc3f22baa76b0a554107bd766731c0b59eaa9412ff5c9
z76c73c9f9d3f4762d83dddd2ccf17fc807be6d7d11b34aaa82483c6eea7a19462e937d1067803d
zaed2c4ef4939b9496328cb60e7e8e5eaea2fdd86fde80ac137d97e4a439b79605d179a9c5d88fd
z33a3dc06ff280a2b440119679432bc05ccfe205d646343ccf76cc99b558b6c439da754dc1861b2
zb986ba16aacf0b87b09449af90c518635267ce5741991a3530e458a5aedb33691843fe9bfd3177
z46f2a61ade4b61ac53fe3893d3409085bdca1962c82d3d157d1649cf58eb8781c9f2f7a5493e13
zad04df3664e4d93be029e30e898eac48cf6691a996e983d0c516f15e796283dc4aa57dba80a9f3
z8b799d7429038058a606833ffdcb83a72a14c5c045c19e7a33edf6274e04b9ce7b1e573b574827
ze0127fcba3165ec388e0d565a6e6c0c184872746338229e28cc1a551e6dc66ce7e9a58171a2a10
zc8eb6a52cc4f9ef80f4694f004afa8aa497447646442bc65dd11454f6fdb31eea0a6b2e62ee295
za1a9a4efd6c314348dcf65d21e669d5ae75a4ee14cfba4a2ca9cfdf4523a75cd032115044ae29f
zcaf4e61f9e8efcb81b90ae81df9ff75998fe99476a4685d9b50855d4fcf06aeb82c6d52a6cabca
z409a1ba9553b96454e119f0c85d38a88abe52d575de825f72c99dfdb88363bb32a2181b6975474
z386ae26a10a09f83a886f46b54866b8118939822d6c8130dadf9183059a4995588996fc5bd8160
z909df9a5a314625c5e67640f1260e122bdc0d9d264ee4f2edd0c219347661c475215c66c8984ae
z38dd869cf3cf70a3bd25cb97952eefdd8896cdd7f380037b7a98b11d8327c492e73799c707b354
ze1e6c4d442c95c3c1c6225b129d2fca1705165a3ac4102b9ef893a6a8f02c6a3c16b1420e73956
z1b6337e2210d8704ab7da7c0a6d685fbac4b3b8b5657316b799a6acf7d95c55db85e04164e3fd3
z5b36516edb6ca820aa8889c78380edf6e6b2e8d52638f077f1805f2b6caf27e81a8644dce30edb
ze0d04974af7e4be68af892b95bf22085898d1bce2535d2272601982e81127bb21e6d82f2795905
z220510f866255034dfdb0257d6f091dda0259d6dcfe4b63b04d795f1ac17c27245f67c127fdce1
zc6a8c0d5fab750af2d83dbf45a17a5f879eaf39c77970e104fb43d698595158a4155d322736fdf
z07cd5ff5012f990bdf64f7d7be95739b331ef3acce89a88c40182b32827a80f23ac7e41836facb
z5bdac36f07f22f97a72cee6ee61a5745d9e83cc9ebeb386c9e9c565c68b5e420d4e2ae2ad58bd7
z9c9df9a6d90cc350a969be5b6c00c659e41609696f5ce1dda3a4a22ec485fb04922f1fa82b367f
zb1fe2e8394c932449d440f87f74b90e91710f4c99795eabee7ac8ae69ee7441cf346c264058182
z4a9a8d7ab711cbd0a3e6e28f56a0442df4dd9995c7313d6a638f24ca35d2f9abfadd5f850514d6
zc14a616f3165ca2d4289ebc3979c75ace9584500d8b6ebc3c56925af13198a3da6be8e05504a74
z663a9d1097750c1708692d2a9dcd49b7371764ffcafb9337473ed2417b4ba7f345f7e7db07a7dd
z406c8080a60a58d02b83b8cdcb057e2cab649873830f602a5a7ff8416d35a6624a2d63cf2dd994
z7e7c57faf6ed629d32927cc1ccbba592007746610e0f8f1489c440cfc1b4fd2cf271870a2d180d
zd9465534b43f7f0ecdf74cd2881b5c3d42e99843a8b9e48693bf21ab46ec8c2675c1daa7fef3dd
z9bd4b5fdac90c4a92f101f8a1acd875e26523c272fdb0421a3a04f713211ca7c707281ba6b51ad
ze181c4db94a3fef8c86b2a6b640c0e2bf0d6767a8d0b05b550c9cbe3c08e9dfea6cebf4477e4d8
z32a1e188d6a7c7c69e7aeaf9d12ae1cd1cac7daa7c0a8f27f69c18e95c652b238c3ca6c83bf63a
z30a9aaa5fd0d5642179ba10ffb88f608f2317b86a6672ca0f630b9bd73134947b0be8daa826c17
zb8e84f717a19d37e4c78afd08bc38efa719459d7b31fb45bb2434dbf19adafec87f8bd11a29e2b
z0d04a597dd7f7f1cfbafc48c1967f4d3294206cc3cdc6395e7c8568f62f89410771de19cf1e270
z9c596b1c051733ff1f2d2b0840171fa14956080cb3b5f6ea3f156a4be851ca057f8c0407dd3a44
za83542a3b52345884b0665ff3f186a82b394f04489435d4146faa439a6e4aa3abbd269f4584f89
zb43a6378548e8160c2d59e7517a47b5e82a48859f1c1c638ae85e019f77ada2c20929609113780
z18bec2701c7b9d4fb7bbca0c8a37d6a08fc4c64fdb1acb08b66dcb55e4e224b8269d7df42f90ae
zb70e009b9dcc7e6d7a84e03b77bd89f70f5a9273507c0355356926cd680251ed11d64f62fb450f
z82240dade8851b9dcb1d4882df0951e81e1d89316d5743226516b991cf42673f62362176631132
z2abea6826a87a87634db20d0522364dfe8cb172a373a9008129252be15941b68801e04fefb3894
za2b464464b8f8f2031e06471d6b7e4b22a936cee804d6c13ad459a01ba70abc10d833bf32701a0
zdb40ba0d911880642303397c5682873e1ac37705428d7c5366896f9e6c465fd9b511d79fbf9cee
z430b5bfeed8af955a6341ccdb80447bf5bd067c85b7088537ee809a8e5cdde8121093a1e1b2096
z6d52e4812dbc56308cc9ad4aeda2d3c0d79604d95cb131216c4359ddfa9f5c26815fc5210c5339
z3f73b6a82da27556923349f53210d33257ad693e670e8dfb2a154fa6b0463cc823173d4036b9dd
za53a61e445c60f25c5837353d2350b1b203157a84abd4b59f1adefd8264a29201dcfcfb30ee390
zaff55bd8cd102c8c86669302316edae695d8f17489df905a00a048a5391c3224a8dd670b69ee5c
zf8951258833805fb6cebededafc598bd2b40368da080dedfa42b67ac0e7f454cca7f2ad30be45b
z13283fea465b3f39c568871a8e8ea723a8baa18a5006c00f7208e38e917477049dfa3ffa57b6cd
z7f5b2ba1d994a60b34a039ee9979a4bc1da2239a9ed8cde457e567df8d7e4367484aacd5fb4389
zb608e02a52d3b6cc6bdf61bc92ab21b41084be9652cdcfab0407ff054f729186be2a4135b99225
z2a1429c360a003c8652b7af821a0d0b6df7751b2e04adf41b44f3914ce4f01ecca1f0f8648044f
zac36268a60d0c641e1d172da943a44b350c0cec7331d7378250d87610e18d1f87b4c1453d3b9f4
z7023c8cd8a903a9724020e521e32c4380132054d0dc9fade84209d1d3a556e9d5fd230bde6ae74
zfe3b98e4d01938fb476b2153422fbcc6b98169a67543dabbee86910b1852e796682205f67d7b61
zd7732c18d1312568c2fef2ab49de1860e93f65708d8724e8dbd5c0907d42f5e14581b4ab7bdc0f
z4ce883a0b535e819c8bda3258f6cc00dd981ca34260b9454586f62968209e0f47c6ac6a595f48f
z168d88466c2650086d734cb42ce186b47f455c6fcf97d8599bb6b5b6cace61967a243e8902680f
zab96bbe5e8c41348babe5b07bb10cff6b9efe39fc185f7e05118cf7d3a39233133f68752aad75c
ze9c29110c73b7c638f18ce88e42f67d829d9b1ec08b2c37c0c1e8ddc8bf5336401f7819b64e825
z907a6a1f6183cfccda3d91322e2ea2a6eec276e71989359293a4282f43bbe7ba63cc0005ea3ca5
za53e928e683d1563808ec197ec1c54c1ac8d04636ef0a1205ce3996547c7c481698c64f59f049a
zfd399b1fff61871a2d880eec64f529e7ca30ceac1487f9eb147bde71ca87c37ac0d998cac846b8
z3681636d6a6998649bd985a080f7ba2fcd38b47ceaf3ca2e59c69e8151d766955a1bbaefc73996
z07d49e5c6d7a6a77b5e85d511ea0ae3cff7fe2b9314309e01f60716842dbc7ba152fa6d2914915
z53d3116ead005d853d5117f90e254a80da21d9ed14d5d63f3f79ea3d2e06d90424d396bc01622e
z43cf813298b38eb4f6d020b1e68baf395c45e426e0d188bee2bdbd6639ba94a87f5733230af51a
z505fea4cc0fe7a7396d7e98a0781f49bcabd7638ee0fd5c0d75c6a1d9b225a4b106737caa73254
z2a78d010f77808c10ccba1194fdf6e6370acef5d440753c8dde9e31022eb02110207acc148de3b
z95b5ddfed3f1cb32eab7ded4eb7d19eef671dcb44ff67b7352f0341bcbd05ac2518b4ed12026e0
z905b824918ac0726473250c3fc8f82ed5688d841f05205f27281544552b17edab6e7dc00edb2b1
z9a9a67bb23bd8b2803ac0df0510ef64200084fe85731d5599608453eb34b73417888eeb9c0d05c
za17ca4304102172e89c1cc75ecc911ea2460e50175e85f63262ec980c81e19f46ba73629daa3c8
z346fd6bdfbca67764b51eae62c37df5077140cd71019e3cc87a342ac1231b54b73ce7be94376a9
z1bc499bc16de1f4ac4f9c2eef7b8e072c2aedc1e696314ecdbfb358047507da8dea3cba2227b1e
z9558d7d78c18c09bcb1056e9b6cf9ad01861add54ef3f79d87198002d1918bcea4a6a0252873dd
z8fdcbe70082fd82c54fd398eb54a3c4820fbee535637bad3b4ee073af48d0b2150ebf3a26d7dad
zbb7caba781e405f136061cc3b1b75916691bc22d2f8b89c04c32935872870e69ce85c3f5d95cb6
z1bb0f38fc0bed50ea44a7e86ac6d1a3f3cab05b8a35a37114f6cdecdfb50d105c15b1f98ba0a53
z5b68d40490b62a54c5898c5ddae5b0676c5759a452f4526d03ad21b366966715ceec3537ae7b4a
z2670d9b943569766e1b954cfcc5896c8b7775181513d675f23221cc4f912dedabb7d6d10a2940d
z2dcab2a7bedafda1cd7a01f0d14bf92e7e9eb7d2c700d8bd9f6b712cf1a3c57632276b94b38e3d
z581142d89e7237e93a74d4ce5cc7aad3f25103ab700ae76e3ea75759c9573ed75501fc2f2f033f
z110ecaba5a413aaa8ac320e1a4a7f14a51cac527b4f53a544c09fe0d64244340fd95c682e2baf8
z99c4fe2d8be73a3e58657ce7184ddcc1405a11d7ee74351c29d9c4d0c0e20845f57e7df61e7dcc
z0369e23e85be423b29098b2c6ab3062a987d527ac5e08157720aacaa21c5064ed8547e92345afb
z13bd2adffe534116e3143ae9b20d59abbb18108a2828331bdbef35c5045b7df9e9075a4886fa58
z0d01f18e85685e59360bdaeca245c69f8846bfe91e5ada57221907ce2c07f4f05f3a96ce76f0c2
z81a7e427d379e4323dc808dc407952f9851d8bd2c2940046e44e19c52a61a8db177411a6805d9d
z3a7c064cb1f8a18dfbb83a38229ebb39cfffee269343b1c15f7415f2dc71f3f9624569edda25de
z4ea80b06af6c83f0e2b02c932b2e47753fbb408694fe973f06b433ee3b299a85567a8852a3b278
zc644600eebf434d7e1126faa724690a153845cd8d427f47f59e92e23d372edcdd15c5865cab261
z5b57fa8d5e555eacaba3bfd89c009c0b233a6a628e3c80a4049170a85c77ae088e8ad0eec20138
zee74c3b0067c9da9fb6eb88aa44662fc5772877990c6f1d6367b24eb9036794f530444e99c0619
z43c3ae0ad76aec8ffc6336738d58b72bb007ce6858c2e2a0697065b1a199f9bb1a4732ad3d9b12
z94df3e539bf8f12b365eafb7ad16770220563717b4f82676ce5855db7f21891e415f9ce90c39a0
ze4b0534e8c3acf2b06709815006ddceb2ed255165933d0aca34fbbb334abd8d29797fc2f05e3b2
zc5ae2b8c18702e754a1d9407281f323cca2c5e05f2b1201a01db7f4233874eaa072a5e098cd9b1
z7bddbda62ebec17c7c2ec6d2ca3daf194d4eb518765b789d969c0b5d97f6f6a93630aabc11def5
z2b426be6f938b9f7e7b09ff0bb2dcab65c5fe5f141eedd9727ecde8c3759bdcfff404864d65bde
zda2c79829c917eb475e3e90260f32206452dbc8ead6620c0893f52e63e4d4e23902bbdbb7ed632
ze8f7b04652933be4dc068b40ec61376089c9cee2d9d9dd0ea2226addd8393b4bb98d3b5167cdb3
zd1814eaeddc12978c784f357ae8a87abd84b6665b1e215a649f49e4dd560668ee1bc9081692920
zc627f9f38bfc484ca479fdc704351737fb618b6c29e342e919770c7c0f2e5cd994efd2f736c3dd
z2823a7d4959b5bf4b60cd570e7fb966d64db65ce6e2dc0460b1b5803eaf679303fdaf4442e43e8
z4b537da8fe751ccce0429bd976b1424b720baa5ac83163cc624c14a12e9edaa51aa3ded0f4bf05
z1fde078c9d2ec563aa3ba4f309178ff1d2889216eafe88e7e721febb59498379eb269a74c0caa3
zed04d97b10abe8a164c7954ee03f328a035d454d884791f02ce14015338f268a44ae97b9517853
zcef31667968fa36e72ce13c601fe6e357e7857571825837f1d5261d4ead6e7d807f7b25dbb4c36
z46d4e2d6ceba3d8900a670e25b10370e8f070bedc30cc3d2e661394453c6edee7c3f89f17da678
z8a2f1196bfbe74842fb8f35a7806dfddb0858389e8a7ea718ded088e4bb2d60899683ae64e1286
zcf8d18f24396f5a2d98bd4fe742c3e30d47a98339c71c48f211a9f9ab29677db9fe3e461d9f8c5
z5b59323c9fa3c179a7434ffdce2143fdf4887af392410f1d4fb55f22d9bce308510c353feb76fa
zd889777ef6e8861e7494497e702441bef1e28869c0ca3e54dac72182ef84a85bc94ccfc95bc41b
z4d6ecbd132caa9045e61b14b8ac0f74e5fdc3f6d59a111e84feefe68d51282b01522f525c3174f
z63ddcb1b16d1aa6ace836965f9d7596be5d26440cd6cc2127c57f68a8d01230f75b28bd4a4b347
z7a87f9096e6a0228fd3276a68dce36238ac0c5bd8dfd52fe00c5af4b767e143dc17de85d26d1cd
z129388c1ba6463d66004bf6fe3c74a0a35fa2a9b4a9252077fc4c33af11f3cb9e1aa4c0b6734c3
zced4b184e59d5d45a2f3b9491c61071bfff7f4f85db3cf3005bfec50128e3bdebf85573f50a548
zb725d0b83627ed7e05b15576d186c5af47532353ef41b4087ed83436d4d31dff478b3aa4ab8ee8
z2c8460f7af1ae201ce5b3d91fd35f7b192443c5fc5a91eb5cbaa081b6576f2c521cea0ed4f8895
zd3d71be2d6acdb97aae1039c97f554e2391671a247715882a159ad0612acc08c448d94dc675b0f
zd05b6a1e53a3d3395ee1f4c910c7b1d55f0a74f941eaee99313f8c14b85103f8d09782074eaee2
z6662c577c9dfe9acc53ea7fc5ea8c53c5ecc4a85f2136739084096f2598da1b62715a162c39eb4
ze745e8e1eaef77a56d1beaa4100e62e5b959abc423f9e9df548e7608d1850a26f236bc46a22298
zfb66aba88f7eecb0cf0fe8675827d88528482e75047e605d8195c9733c9c1d7b40e2fa38b639f3
z23dd6a7733906bef6bf2420ab1fb58fd7d998157a16774ad8e183ed08a6ecccf443f530d79b2c0
z2b56c04dd1db2f1b7f503417be95fc9402afb97ef24ec425c2d631d7f3615221a5ace249497e5a
zc2e21d62f14786ddbfc9774121114358811ba687dedc432a0dc2ab22149d6b138b6aa545103932
zb70b5c038c88fba531069d6bc7dba1bf96bf98ca8e48e5dd6828b76d69dd571054c481936d58f8
z5dfa40590e0631a235f93574411d36e8fd7b398ab39ad64879ae4eb800aabadaa46a22dbf4c335
z431b4d59d89463443432f1d9e0e434871d00b80e5aa3acbeb2e42253705acdca8d69e297d68f82
z7e20d48ac27bfa8c63081bb4703b62c9f0ce81d10c5b98a775ea654cbf222327556a202d2d5d3c
z7d76a84fb09ea823820e539806d7bb1230bf50c28843623049c197ee60ec79108658d524059d39
zd97a40d2f4f96b1aba66c292e7801cb3479b350a0b36a38cd3f3f560eaa3da7afd8d43d7f14801
zb4ea9866d1116aeb4704665ce955222f3d82214e879532283ead5191fe27d43b0282e7dac2404e
zf18f77b04416e6d3f6d6ea2c515053093b3ef912c5a91fba039a28f1a2f8a5608dd57ef96c6a1c
z808709c4a901f883ce79c3a0fac918620261be306d8b63c370158f3bd7dca27adb64923c2b4706
z27d8c772fc70e867ae550b334b64195dcc3c75719eb6e620a12e906e925c37edcdb14f19431104
za69089610db441c604d06bd24d96e0bec114b10cb4eb94775a9c4d8020a57c0033ee616713de8f
zd2c879b4a85ba43f1a4dcf2c2153c055181b0ca69b9e0268556cbf07a5eb34e7bcbaf3d2ac03a3
zebe1520495189c8c5922d1d5adf8c48955cf4dc65fa73b5bf3e1dac2df60df6e0f372a87fca599
z431998bde1183f36545d9c821d5d7364f22593afba4c133e2690cc83af20dde3b91f4d4ddd7cae
z7ef8acb7148e9246e69be0b54bf39bf8bd635e0a3d0868ab2bf2bbaecd6c3f05c38ea5bb1d04e3
zada157ebc9fe97bc9ca8afe924765d38a2d124f608bf3668c3a7d637e3c22d2c2e66b3adca1676
z2a438d34e1fb299d0f6a09ed924ab4d20eb525e1dac744f2e4d107ebafac70673cbe1a90e73a18
z1f75247b903c886e4d455321f21834b7a5ec8ca676f8a33f63ca7b0332b4eec5cbdd6fb59cb6c1
ze2f0997be44ec7a161ef8c1a143b51005af5a8d6fd81a938cc28cbca1e4d0d69ad08ceb9f74e0b
z091fabcc919b81068beba1df4bf267f66e095a5fa623cc050e2c6280200559aee192ed43e308ab
z1d90ec3cbc75d006ff0ce87413280ebda59b323af6de5df8c809bd0ca5b07a68dcae67825ecabe
z829f5111cf32b9dbe731e96982f693d11c17d5356229a762783c7aa1bacd18b0107502a6c685fd
zd9118586457ecade55b5954be2a3fdec5899d329f7def5742408c8c421ace0c84f18d8223d2afd
z0903d34f4f4169e6df4b176d188f91dc14b0f4eafdf5954c611e980557fee04fc21af1bcb47921
z17671104ece153f7c076d74a48bd61c9603c57b4650670e15b58b0435bfdef215e365d5edacc83
z64ec9a4c208eb9a69f752b26513ce8f61dd5a73c8a56a4828d5701bb921c21ef07b01189c2e167
zedbecd8035682fd2ebd22c25725aab91629c5f128bda269924ed0c9052d1b7ef37afea9f2d772a
z37bf69c75fc76a1e9dc92b33732de82bfb74a6d679271944d75df75a8b98f03f69d55239a2086f
zdeb9345ae0b971e5e2db7a7b0514fdbf52dc6e3f955e287358dbe3b1d6c3fece49ac4a8f7d1cc9
z27f671325a1191d0b3ad034673b8cae688477598ebe2c169d828ce9c21f59a729240a641ef52cd
zd3be7e505e95535015dd93d19d26cf9e157da5609da9ac5180c1434c11cd730f4cc525176af535
zc889f4dac51250095ca17ca2432241c0b1d7066edcf6769974bc4a7ab09501a2140f268e3c619c
z560a51aca5a22df9c70b6444814c7428f2d3d2335affa00bf7f278fcd239c25663534ce15294eb
zd9a286fe300d88ab94025ec1cfd7714a246e4d643aba53e587b45d79556afb07e79c405effd913
za41e5d583815f7b84051eb76e30fd207ce3796d38f6501644dec388c95fded5bc24d46ca4707d8
zd8b89074c59e3090b4e3391c09c201be9f37b4e6e84527fd76734a1aa0caa3b0dfe8847b91f4c9
z83b1fdae10674e904f8802735b546fe178560bff03993dcc8e8e207426066e505e876dd6abca61
z576a4fd052592943a29544e2f3856ba921e95a96c8e5b1198f7e0652f94453b8ee262145a4b72c
zf20288e7cdc15e51e65631c4ecd55f8648cfd3df3b13959e71e1b2427522154e75ea4d6c8ffc5c
zbb87c2f571e4a82930063b269808ee5f3b26d67e5dc7623ff8831bab5f9b52f2b4ecc6a68ac934
z1ca619d6852a1f250d61a2ff49e39313747643b4fb1a852c97b5dae05bab8442d4905e2a52ca0c
zb8a6117088c44470d0f40b192748fd7206f447ba7cc97e431dd84172b324fc67e30ecc6aaa70b4
z6c917dbf90670e44425fbd855865fe37bebc98d84d02458609ef82498c3c6bde4fa05b6a4fd465
zbb1bc9a5edd4b54bfa166634ed9ef850fc5be987d26d7cd58954c139bd506051276fa3466362aa
z793f3a528068e4b8cb7d4577b9edda392a6e6ea9782b535ff2e9da951ba9f4a59025645ac4ec61
z8315f323cb49aa0056645a26d75eabfd0511cf9b6ad1e12003e497bea5099acff301fdd810d200
z84b5c597cb587f69e5d8c9d08c1458b4bd127da6cebe431b3dd44511182941099755a9224ae96f
z7013754f967feba8cf44662c221f21823a805d535808404b852485e03b34dba2cc952f1e286197
z20ed37e3b5772ffe614761a2c71bda59d4912045e8d5bd5ee4b3d3b9c723a6c0f510a55d2ee6bd
zf05e086eed5a4fc080e643f10c20957dd970ec92f3c3247c32b73b7b59f701c76c6cd66324e9bc
z66004ea03fe828542f223a97d75d6d12275c467263442fc82aee3ce144bb57af68c9964a7019eb
z9e274ccf38975a7d16dde4e324f92ce3781a99a2776b0652af8affc2c1251addb8e23fedacc44c
za564342edebf06790a3ca80a21afb26de452944457df765d458667a50c48c5e3c1ac47ccc44460
z5848ce651cafcd144f16ac9c885f9a7aca6ec231bd5725d046869f9f2fd8d1780373ec948145e3
z21b1651ba281d0ab6579c9619700dae7758ce5d42227aba1947b342740929e477a8f6e4bee99bb
z196ab0ece964de8111c7b49d8f85672d555e975de792e1dac67b8619a0b8691ad35024fc3be2d7
z5ec95f728c12e8664b6b3e8bf228dbdfe01df1f126d2e2182cf5ee9474e157333bdea56809e338
z58aace3c9bb6c6379ed843f601dac68cb99d2c054832f260cdd283ba8ee109193894000050f95d
z3c1ba6405466658d39152a5ffb1422723c7da724e43832074ee6bec71edfd014151ac07f2e9186
zefe8f64bbc4e5d466a6d8c2428bf9bbdefc2c48618709cd2d3bc11b90d402eb99566cc3d9cce45
z4902fb0a707fac66732fb130cfa3c30b7e323506f68ed71a8af41826b8fbfe9e6b93a7afed43c1
z94f829e673524d68e918e4604d09d340270c09f1b5351c8d4f01a9c467868a83134a29f2217b5d
zb3200de788100cb6f74c578debeb41d45749ddb92617d6d24f66788bc160f8dc89640f9380ca5e
zcfa68dc46b6e3517c055c4e6f411d8ad97ad8a026d1355d6d1a4f5de955a420228275407648326
z9f53e01e6851745245bf08476c31d18e25e35a3240e50270fb04bcfd2a650cd4e1ed5d6b31dfe3
za6bc7686ffd95e84314d9ff8c900db964aea294f6dabb1fd5ce1e6e5ef7c40d72b379acd77b1f8
z0492774ca1383e5408ac9dd3ac4b48321ba9acd8d81990fb738c2b46bb67b60d857feea1f703af
z5e28e8e025a512d9f64d3b8ab8e6ff00f1dc0dfe7ebaf74633714cbce126fc1b516b9ff0648fef
z37a1065145a0466491bf35d32edc61242e72a75873f2fa9d9e09a03705c6cb71cd577ae368002b
z726e7716273719cc1acb216314dafebd689f569e7eac98023010d5188aa61782c506805445dcc5
z2e380a9227274646c8aa7b7c47595200e38c3f9d8e51300f9a27ff40513b2f68e26095a7520575
z58ed66d599840c4ec7fa8e6374f3b4b9b3b037fa9497f62403b798f416806e7ba929feb290aa2e
z273bcca95d5e287910c0f3225d0b9f28ff8b7adabcf5c5d99223c4623731c7424e34dd6593acfb
z2221c6355ebf46c015adc69e741b3780038519edd9b60b41db72d9e94399be71d027bcdbb4ea30
zb53ec551a463bb0645319517ae375b36cf40496002f3433e6e22ccd756b8fda3b25a54c54cb8f8
z83f98c74d301970ecfb534fbec2a592ae3407848e5ecdbe786239eda4ddfd3fca2062fe8879c68
z5d694a244d7a34824920a80898b7355fa2c5a3ca213eb4ddbfa253c23017be4bd5cf96a6c5b623
za899bc0ee38e888715b02acf8892e578a262019d9c2ee67de435b1cda8bfccffb342f7ff73f1a7
zf491f49e262021dbb8e61db7f895fcb3132937e5483a519aa8dee0648f026aa1c72564d1f303a1
z3892bb08b3fb1dbba05d2e2dcd3bd35ca53bdeccfdffa0fc4da9ffc965a5e10a5e63fd730b4355
z9aeac30a588459624fa161ada6c125d3fe594199b1d94494dd25a4d95f5c64223e1e8ce8149910
z6c5a248bc24422942ef2a28a800ba072cc71beb7ad64e1f1c3f45b4c32926f90363a5aaf754fbf
zfece5aee2f2630aa192ad57fef4a1636125ca782eca693bfceacc66d2c40ddc8ee1d0443ac7ecc
z1f1b15d6e6d6c4536b4d77969c92cea852d506d3395474615e8eacf69ffdbdc2f355743c307c28
za600b2dace9df153c5ece7b3b82bb8113bda7e4c95ce534d713b111b2852ba1e53ce05bbf49a1f
z15893c72b141c1eda23cb70fb4081829fb53a8b56cd71268fb249c9876cec490242ecc8734814e
z5863f1f01f8773e84ef05ea8c166a6547a972ecdfcbaebed84397abbe660852928ca39318ed45e
z06c16a50ab215d96b841c0e9735a3b11197265160d393cb3736bf7cab7e9572cce5513fa0cb3ce
zce125eeb0c962a422ab29d92f0122cdbe856b39d1ae369fbb9a135fd2035044be8221bf219e185
z7460df47705e9595bcdc51608db3a94c38ff96ff47f4261094d4456c09a5783ba2ffd1e06fe4c2
za6d49ab694b70e3d589dea3de70cdd0c8f7f351ca2419445df08c7255b19de958b0bf5dd1938f1
za8ee6f79490ffd4bd4e96e16cc7fe524539c77438da6cdc0e3a97dc68f410851b58d923b6ce10f
z5e85e2e25bf828dd6ec3ab1bb8e7ae47b9aba945b603d4163b63f4a326dc5694b86b12c9f5a29f
z850ffa4f4f50cddb3a04cb2b6162ade90e74d2978292c7fbd1f19fae5f394106f7f0c7c2b127d2
zfcce98d6f0748aa266309f2cb03e29d6342f40be97e27449dae7f953b2d7dd104d4aedf19c8b55
za28d0d1c2e0fc091da0b70ec59254c2cc4368b5fa6d8c71e3b8602e4d95a78ed4417fa1f7de1e9
z7945e3c789ecb953097617171b9c98322cbc45a04862cedf24ea7e6144c95914fb0cd7528509ba
zf26ffd497c6acff28dff5aa01f5856f06d6b2a41f20c7640786fdf09d3e772fcd1275a1be3abef
z54f984bc22d5f507171ef0e153c097b25df09195bb7d367a2d35422201a93442aaff8df0237472
z382b06733e29aab58233c8415c1d78403efb6ffda3e94396f0082fd23fbfa72d576f72327172b2
z67fcd4434eae033003d3df9f7e41b1601b5e00ae677dbc3d8730b3b4b1f80739d80d2a76528030
z498366632df79257a65bcd188b551dcd4cb92c07ce57b35ee6e857ae4edf8872a00a5f9d278e17
ze9ea72c1f2045b83781ba85fd029e8d73b483552cb6f4f7b09b9a3a8c43bf5d230e58f37e984ca
z6d0014017fc02dcf745340bce524e70321ba973af351ba0d43ecaa63cefffb10e95728fd1cc52b
z3ecb7d468a6df615978abe8bc90b14e9972351f852550b8607d270872db7fff55e7339fb62f732
zc0502034602895bf629c98e12d8ca15e7c17300f16e82a061eebbebe4593bb40e005b6fa2ac46f
z81cb1245965d58fb96d096d406b72f020458fa1212fac793441be7c2cf0dd3481bd50c1d55b2e1
z3c1dfaaf615e71a7cb41f4d1bfd988d3d28ea9e2495e7ee44d9d810d095b43b3db269eee669d54
z13e65b7d5b09a4b72a5fb0efa51d3d2d416ce903049d49f9b0b51787ba0131226d024810fb724c
z670455fe940930c95ee20ac482e8e3dae6800cb09ca3e260859a053a9a13cdbe4cb0181feb5131
zd9135aedfd0cf52091bfc5c4e4777c5ba4c2f60fb5585d4c87f8c5c8654752532556f4422fba4c
z224fa365a14227f86dd637dcc7d324cb066ba134d8e4783e554b502ece4c82e3c2792c8b4e54ed
z5045b6cb5e8a2f8abfc6f470302cb9adb51c2d0b92f97d9a4a922b25f296e0f34f5752fe01d4d7
z4d42e5773e93e7691399df8b50f146370353bc77a8011eadd3f682243a9c8a49e2b04508dafbea
z552e94e632de79624433455f7eb713f004b59b11035b65e38fd8986867f1d64f463a8ad5b168c9
z90ba465024c097ae4fd578ec03c5f787ec5e23ea831362aef0be2c91fc5d565aac77fc372052bb
z094ccf24d01f915b4aac12779e97a52ea59f68f137b569fce0acb69172974a18d6f907bc9aa3df
z35aabc6bb1a08e9724058260cedfa8ffab1af77a0883366e072b72ca8833261d9644dc6a6cd9c5
z4c4c1ead47904787bfe2019ca4f537d5560a0f7acf56bb654f7aa7591998d2ca5dbff7bb8a852e
zb02df60e2e8a5f95f28808bd3be682db4a7d57e1f8f62be6f1132df963f8d9706f5dfbf50dd0a9
zee348744acabf9449bac1f02eb5ea5ece2bf310d5769f7731ff8879b2fac4891b1e0cbb1483552
z54480332b49028ea0b9d47f069f5769c08933bc2f51974837dbe8ef5a9d1a7ecdd4eebeefabae4
zf65657c29970d7dc946ffe737247f77b5e8d8eb76b51dea5eecf5401407d7ff3f33d37072bcc10
zd237ae9b767021b7a33f6f3d8f48259ce676cc9f027185e0a42e306ea092113b9c9b34e9f46fe3
za5e4fc90bfb7c549ea56c649b4931d04c2a481b622ceaaf2c99b4baedd63ce41ae4dff0dbfa05c
z9b5ebf036ec201ca873fb72b9904270dab1c53d7f9c3fac7e58a1b00818ec94118afa0d0093fbc
z542b2e18d9f6746823942f7ad2546d2d27e0bb4d5bd83d532240d844f5352e367bf3560724a29d
ze6f96bdbb125aa371e232d89a87b36898f0efbf6b0e4bb83f6100132838585b64bdb2aa8565c9b
z4fef536c170520d83967d5941c441b620e56e644099779a4128f30edf76a74280f47f3e451e303
z8ee08cae635c26734422cf8a0ec4fc1ee401a3d6721f79d874d68ec87b1dfe8acb98f58b1cdd85
z2cead302ee6dde0f9657e622eff6a7b5d1311d31cab24d7a1000b23b99a24a3944a036db090b6d
z5c8e0f7c71ef4f1af43fd600d36a7af5feec599949b28b3ff6609dc3bece62202170a23d07a803
zf8763ba694b26717b94b4a2a3e2ca26331f63dc7e9db44329b02f493a15cbc7e1872e75c1b151d
z5dd510fc825c392b6dd83e4805004340fa892829b07c809cd31c9fedc92b6031cf0b574551da1d
ze9032094eca73a8a02ade858014e43f84440e09d5cd63ccd17a00ebb376848217b66bc7474e725
zfcba6ecad4669f313ba9242b166b3ba390fecdd3f1451270c3f32eeb35967d825d8508dec459f2
z9366825e993584a6d2d379a07b2aa2d1af4eab6e656aa3accc9d7da74a8c72e7b182973356cdd9
z791503d145a21f3b4a6aeb947736faa4ad056d39f47b5151c74c14f549e9bf5bd595b99802831c
zb003289f0b16921abe35a1a3c4e64f423c522bee83bb6470a00600f31d5a94df4717a40b3ba403
zaf7a16a1ed54e7ef09debc6781ca35d60883700f5f888bed02ea5537d5b0b6c629869186658a7b
z636ff3ca86a4eb85e30965d7a457991db6f2311e910114964f8c22edb373b406e823d90e615a84
z40998103384233d49d9604f74f8ee657f9cc73b59228ff78aa855232861df185bfec96fefd8a2b
z8c60d755294aba679489697752bcd7abf74f3fe2fffee808493cee3a9eb0d381c773f9e24e1641
zf8c96c91a45e8cb662eb6aa3672c8448ff3f9ed95d0fa867c5e765e2d612740948be79a072ed0e
z322dbfc108cb98b1d7906651c872d005732b3da143bd7b84782cedd22258a62b34529382245f88
z1f883d5eb05b691adc36af5794583edeb854a2efd253102347e61f77b7d206dd98b55c7d2e9960
z2a2d50f82dbd80c9b68efedead75183ba2c7f0edc89538dfb7f455d417ad6d9983f31742bb19e5
z84805822265ff765bbd2e03fcabce660a002385d326d5ee3b56868f909e9885fcf61e8d2931e8a
z1d004aa03ae3057c51ad53d09209ab785f61deca80abce3e835b0b73f2435c02aae6c8f1642dbb
ze57f413b633f0f872c39271ac9a72676f651dd49b219df0f39fc05737444c231e73218dd75e12f
z9a3d727a2ba7ac8eb7fe8ffd7fa9a9843d61e467832a87418ee178e1c9619c4e2d4acad799a93e
za7678aca7a38d0447a08131cfaf15910e87a075f502868f7fe61b9460b67ece888c8313e442359
zea20ea9f92dd73f61d4e18b0be9961f2adca1b3ebe8f56adf1abeb1b68b53c586f992900a914a1
zc741a5ca78244b0b5570d0604ffcb46ea0ab8aa93e9d088b06093b111534556ac813e7cb3b55fa
z912cf44575237625657d050623c134a29271192ec15471d1ff325353b9fe3f06d93828d296e7fe
za4644da900da0106a3f3ec47606ebf6b3ecefbf6fb42dc7a7da0507513e059d153bfe1ccf03644
z66ce4092f14d124cd423858a7586f29705108fff79178a5f4549abfac3d0ead77799a6761663da
zc68255b1fdd2c13308c54ab2ee795f91576d182be9e98c10927af315b018ae9b2462897999a244
z9bd2059141099ff85f414b06a9c243638bf86a599a54e9023b8176943b14d05336d5d39dbd602a
z05fd47c43b10090d7171354b26c2f1a7465540b3b82b6a849965b2a77cd6b5612916038707c357
z844357e5f495a1bffdd3bc65edd8477fe78cc01d034a05ab3f88bc22943370482927a9b7c5b511
z316462e1eab80288595089ababcc88fa2d1b12444a22e6bc134dbeca6e7939b4321c0b40115bbe
ze39a7311256fb479611e57d1c81d8ca26b2c34d28cf0acaa520edf98b8dccf335884fac0f03e86
z86a62a44e46a4221d4956a4f03e4c41c57d6be6359345aafe531a5efd995a68d1282ae6ca1e159
z183740875b2c89b3b449ffaeb1a24327295c482f65efe7199d9729f688eb679c669f16fbd748ba
z781004bb277f47388b0eec2071e6c6b4802360f0355c4d5ab9569bfc933a90fc95a13eef943ccd
z18bd44911076480783ec4a912055c9f752795dd16686e77151610ecb37eba02798ca73f9122776
z40f10a33f8cbfc4fd951fb73d70dbac3c867ccb18b62f81fb9af92719778677dc217c2f8b8b8b5
z93e735442be59e10b4c52f28a377995b32e62f6ac1cb17a6df6f9f0ee3c4cc7e89b416d956a46c
z622ab2a012fd2c7c260219b84371de4b35fe4b60ffd8c8c364174b4e15220202319c8ffd514023
zb53f027f3267e60a9f751f077c3d98563c971c0644455e9db659667ee0c793f2141021f472d214
z38fe9226e89718471f69665105c3c11acc84860c2dc0ab5f4653ee057e591276b93059688052e8
z4755bf0d9d633ad7351c2de8b8bcd7ed0d2cb4db931c5792cd94bd3340c4261fb4838e1fdcc368
za69d34889a9bbb6c4c220ef92fbb92633d9cbc3fddcc02fbfa5491dbe9c1cc8259703c5a1fede5
zd47b120701ba7f2ad1215dea56b394087316c466ac26d348b7b094c1fb7dca461814cd35c1cf4b
z6c1cb05de52a17fb94a4c8e8d777072f4732686946c7d5f7d1d7b8eab13af22689580d01f6c06a
z44bc5aecf42c287b3686b0646236a1358945c9b7fa700a3df0a044088af1d2577da470ef0cb019
zac235a2d7004ccd69215db7c44ca70a91e4dd706acfc5a82e426e9534eb911ab6924a8656a8b82
z800b4f1ae7a057071e413ece07b905172e988773e6d40595b5e96f08fc851ba31d74d48a9eb77a
zd528e74d007e2f989d1b88e0e56da2897bd093376bdf2eb47d85a746ea738e259e5f14b90de69d
zcbabface9217cfecbf0a7d58af8db1e9af2c744104c312c62d5d79a04dd2bc2aeb5fecb71d2f72
ze6a0ac08d6b61dc9abde6954fc70b67a5cf0a2bb1fb709b21df36eac45cc02032f43fed969d605
z6623a0c1e645f756cc369d02566218dd85f1028d63c7ca67f8146eb1be1287cf97cf2398b9f40b
z9a8fd3343e757a2c89267fcfc9ac42a420817caa456aa9472105df5651a75c7d1d17288ca60794
z91c84486a7db2ea1e1885a12d5c383dc32b2e0ce8ba32e4d0d69af2560f8fa2bd9143bcf64b30f
z97a33bf01ec2c82d9b276750141657c8b7f4343a378cf081edc2f4f38f4b435c38eebb6b73b266
z5ade04fd6c9eaf7b156a192cefcbedbe6f50f6e6e0e17b315522cfe8a2ff8b20fad98279170fab
z667c4c5fcd2a26a90d4cffd6034d5a1e1e4cde76e80d228d978c65a5dd2c954f027824328f773d
z9db08ac8f47fcb7345f44793491706aff35806c38e50a8bc5ab0ec8368f005cc191af14ff942de
z82bd3339544ea0603037164644f2f0ba08cd386297c85cdc360f7bc915a17a7ae876bf598af21d
z593f4fd470cbec29253e16b8b30fe29d088c27d808b16270b218720c0fbf8a79764b0d579f9fcc
ze07447f5c36523e8823c55c5af667346fc0a945d61bac7f226e84584df174495573cf16217a1ea
zc3666e1bb8e3ba9e9d29dd2011c7d8a2a8cd2f61733c3d9113e7f307a8519d70646a68c8913975
zf8994583d322fb255ec1f7b6568e96d738ff752b6cb50a94828c2c2847c464e6c2a92bb06db810
ze91b015a9e1281dde3e948508bad90341b62c8b2fd19ed59ccb8e9b6da8390de11e6db8dcb4a09
z397f5afdf2158b931bfcdd861cf564c6897ae6b707376ddac799f745d09f45d4dd0c72437a8749
z2e23b01eee82b82a0253a8848865038d3a67d1591b08ffe7b377f55045fba9ef3ad7e48b218fd4
z5e488f305e8c1b9ec3685dae818774a156142fc41ded5e48466e5b46d83147fd3f07b1716bb8e7
z9826fc1ecf8a8e50afefea28444767bbe82fa392d049836e768b1edddb51cb1ce124c39daad83a
zfc95d570fbb1f0d88d2e72c7c443feafbda081a931e9582dd0b8d101db1789361ba71e408d8407
ze88692c2a4ea88200fec6c544b525f9101091a96c4fd017e5cbcec09b4d8513ac7f13c926454f1
z7989550bc147c2b132d2ca2124a0efce18dcd8e79b5b0952024c59abbfef096c67db65f1960abb
z39a4d2728d1b2abb0d533a232ca27aecd31587682469ca9bfbca37e04fea633670bf6de9370310
z1498cba0eb38850061b8ab904a9c554ac68877ccdf0cc5ecd6268c67edca740b654e56d62aaec8
zf6ba13a1eecac94f5ae074787199f1212484d6b54436d0973ab1f360c148e0d8743ebc6194221d
z2112545f029018030f6c72ff2c7b2b471b89bcb7bd31dc03b9480e33de0b5762d0f6edfaefd06f
z4109995e63b1be0e1b813de1955a1f2840bf09c332f4bdff86d743e905e6332c00a4b484fef6bc
z708a2aed289263e17e4c55df82f392c71d4a78d681bbd2f708d0663ef86b772a8ac5e033688591
za549f8f827aeb189bc243bddcfe2a2deb0e0df1b702c297f3775755ca642beb016d3f95674fff1
z81918954742acfb31b9ad46ea8c56c0029265da2e48a12aa98bc5c3479e1678401cdb2ba04c8b7
z584247cee0fa20513134b34a0a7da2239555d5524fcdc9fee931c753e41eb7d8fed917a4da375f
z06c3bf2490ac5c8aa269a01156bf81add0ab931970eda18d2b4bcb3101a4a3e985e2d2a892d572
zc588ae7f876507d384747c5aedfa899a345671c10f01b5373d19d76c8d8af48fc1287ee7f6d3b6
z11a6845f5a22d65f67155c4b45d880cb484860c14e699be9a5a804764c7aeeb5eab6cb22e5c28f
z5ac76fceffc499e80fb0468bb5f18fcbc3fdcfaefd2f152e4c70604aa482c82732f066a4315a36
z5d74ad2992803b3b91e2ea3cd529a25e10e527473f021bcd8c0ede063cde2319cfa51b8d335ecb
ze7dc2e73e8b36df02b43fce04c6e38df1cb7ca8c36c2d0e7b0370b09f277fe6195744114944ca1
z800e5c435cbc82cbe2dd7c62b00ba85c0ce77181d16b38ca8a83cde4f12d90cd2da446b8bd8e85
ze93b420d61100036c0cd1cf6d647355563332a836033dbdb7a4922b1f44571cd105c950b62be01
z57977fcdaf090396119f1839c19af1bcc8561ae0443d961feef399732f6f00a1283aad04369756
zae909fee80c76a5c030cb5661478ecc18414a34d637ddc8844c0f26fd2d2064ff9621b2a1f137b
z35f2a95ce734682fa6b8d1c3f31d55990a2f90444dfd0fcf3d55a2c91e64b8ce141840f1ccdb3a
z4755456548a3dc53664b0ac40162d7e36dec33ae6b179654cfc5af06728c36da9dba6a23cb2949
zf255d6fa5e2694cf03686695168fd8d9516499329da8e78b10e1b086ff56f285aa6cc826630379
z7fd712d5f6c15f6110de2fdb76b8a2c93d0e59ae68b082e9c9e3b3433ae97a4cc1d3057dc891bc
z00ba6b61d2db9711b864712767398c9fcbda45ec60034a4024597db067d7d9c3f7619f61918916
zfa71df48275d53d30ad8cd466b76e95c678de78f1432b25cda57dafe742ae97e5d15379091c0c9
zab05378735fabcd3032518d299aa00be3990ce74770cee1a4118acb6ea2fd9f876a32dec08fbbd
zf1375693daab969427c476f9a847cb1750cd45150d90ca99a86eb7665d1189056f0e8cd3908cb8
zb47b05adb5c2eb201c75304d23d1ee63a5975bb84b78114f429be89205a17239b59988ba838666
zae3e9d6e6013b2cd4fdd9f815ed7f0afb6cb48e890b5183716bbf5159b0c1018734fec04f7a915
z5c08c798d07c92200fc6080dfa8b6969ae9f6220d85f3a8174bb4409c2f188fa77208c0c07929b
z4baaa5fe4b23b42f87b4811ff140f2d89c4ee284db4edbc72c9b1d6e8c44e524d6dcb8c401009d
z63b47eca7faa1b929621a1d22e02c1c222f742f0ab40a5515af308f420197e50336c877355b2b4
za2bf6230ed09d2f4a375a9ae748cfe2ff4018288f1bfc70465157ffe40d906c0338b8b116f1321
z95ca2d6b1a72bcce8d6441e7e8e8fba471da1c1bf5fba415d0f81bb3903377bd89ccd35d9dbec8
z549830b1707806b672ac2db09eb24188bf0047b485892fec8959fc67b792e0a11dbc93a4f7abdf
z8573f2c251bf7d48ca0324a999006733c99ad25b790fa811574ff0900a7899931b324ba3c2bded
z6cd1fcfc937e30179f442cde86c51cc3bcbd4d2c047c5f185946b9a878b6b6b364f00928e10bdd
z844881f1fd9dffe6c12ae33a06cc4a3c4548de9b10180174a281c6e99f6a5bd63f655e95518026
z962af28dd20947acf0cbfb2908e30537ed4d16d7d01673f3471a2dba72b584b94a49e6d0f5eb27
z46a0cad5dc42eff76b8e11c7c117227e065a9c17f0b2d4e997f0ec5addd3752b38a581f284aab0
z221d20c4f9fe2868c91bab981dc15bab2bafa2988c8f3100b2c43fe4784554a5ab5337704791e5
z85e154a56bdf21681ad84dfcdb4a0b4d4b17522a823f74cb3e4ecce1d85c3366cda2ac196c213c
z5ea13b118886e6477eef9ccd31d20eded9d0e79454d33248c517f8b5f4c09f9d946138831459b2
z48fe2eac147678f892a9426bbabf64b8f3092f6b440260625e55e2dd263b25f1d475f8ba7e711e
z996d71498647a8359a0841c02d3f25157f638192178caae2c22e849dcd0a365130ebbdea65963c
z13c112ff8b07f29188e46da2605c016012b108b829c6752be38870d4f382157b7ef5e1a34c2185
z73cc6382fa5803c8a0e72e714fb221a1996afcb2b16b3c2364772c3b3b0d00c68cb83a0e71a4f9
zd17a80bb1ac4fd05474255ba838254574abc8308ef8800408b2b2a3e8397c4fe1d5d31bfe44eab
z56df56412672ee1db6d5d19a895212a4460a78729e68e7ab7c89fa6deb9ecb87399f37fef17e67
z3359bed0d6566285a7c962febb3c155bc3e9289bac842cb618087c9100802e53f91e10264ca6ad
zd7f81e7770d1bc17b7221c1849e00d1bcdd410918f12fd86cec73858b70542bc9a0ddc1661a3d7
z87494338272a38634e40ef97eb6c9b1d73091302fb6a9fe166863126b2749d441889a1fa6a369c
z707866793a0279f59dad696ed0abeb03a8025d3683e7fdd898310f9887cd84f81ea747bc485486
z487bee212d508c7545ac30fbfdb735e3892628c1ad6ca353b003cf031fd5fd97cd20200cda0a63
z5ef1148363f5790516400efd4452d411d68d7e6f24d0642916964d816bfd10e7c92c48dba63528
za7122f542cc59f902737ed2dc54aaa3e943afe96e1da04cf7b6163646e1214a6e00ae05e50f900
z900274f231b5d515e048caeaa1d9b0491f463d246feb3b551156dd11a9378fb414ab76eee86f37
ze75420b3efc2ede1fe20ec8bc7b28e470b2d1331336c7442ecc9e9cfff2c3abcb84879980ff563
z7aff3b1c7861f2b0de2c881f1579f166db256b4ef08fbbc0e906a334f763c1c5fad72e1f99e099
z1e447ba2a1756138821238b7a7b45624abb5d42bcb8bf36ed83c1864868ebfd4a840668e1e9ba4
z24cacd0442f55e7b27b4ca8c7f3d6060bcba7166d3dfec718ac33c57ef3d1ecb310a16e30390fd
z80e8c1da963331c8828362e9b97b66fdc5e6fcf8ee2198413c021cd944a8f24ab6b28e4f9af5a0
za8ba3d8f3d9b10e8c084700ec8723667db31c5c1ef14e06e573f79eea91a6a093b26955396e2ad
zc190186d34f626f51f34470d2ee6511dcbf0e3adb3c63a74e08b22db8b24cfde6150b1d3d4814f
zc681d44b8d3341ac4aa644dabd3df19d9f3de47bac1d715859031b8d63704313f8b3206519e916
z42f536ce9291124d8c7a46d036a14d3bb4be86e7ca9c49d4107ad12e87ac3cb18e78f708ca7f8e
z524cfc8cb466aba309b0d25469727aaab3b1dd9a5aafc71841a3f84dc5c20441e8a705aeda07c4
zecf551cc8f68f93468fa5d0da12c3114d1775be44ddb898cea4353eec8b51eb48d2cafe25ca579
z4ca39f5e526b8b2e3f70e4789508a359ae8f2677cba5aaacdfc1703c57df5c7687e34834ea0494
z6ac843f22ab4e8925395b0bf052bee7bda9bce4fa858efa34a40b7c98a50a1f37774d152bbf5ee
zb03b0466a5c49003c1d65e6ebec5b19f0978356b674f2e581522cccd58acc5ad270da771d6a3d4
z71fb259c8ac9a2ffa1864528bd0b28f5b66c652a2e8b1f6b3a61615416d6d7f2f0054babf6bd78
z3d885bc168871c574491ce067c3fb9ef83d46841de5af186e811fc2abd0fb0de6ca2d879b61e60
ze87052d9b9e65c1e23d002219bbb7925439049fca49ffcb1820bcbb74f55efb0f418006979723b
z3808c3b03ca4bcddbaf2498040946e5ddabc8831d96534305a0c09ea47ede339859c21e9d150e4
z7116912a987cc37c2c8dd66f6211247aa97eaac7402642b2d8b82471021a1d5c66d23d2686959a
zdb743a049511155b4d29176a920e5f48d8e9e5b84b325816c8ec55efece19c4a00ebb27951145d
z806c6604628d551580601cdf5d6a51383abf6ba7e2f6579107d340df47bcc504c0893e3a9d7661
z37e33b3e71e12563f10a1cb61987919a255a69c645b5cf845c45a22a382dac3bc871bdb85e2c5c
z199a84d2aff459f0e859a9e9fee5456ffd05d4b8db49fc4fe230a9b87d323793ce0d85ff415c70
z97a73fe60a2228ac053c3c1649a2c5c742c2ae44b67ea28d56b59f892e76d20f620829fd01abce
z96240b0ebd5be22789e06918164aa3268be2ceb2cff8099613d407ef752deb2ceb901d6b897491
zbdfb1eeedf21ebab7ea981057f8648022e06c25b8572c3a979accd11b3b39ad2a6ed64e1c1505d
z5581f754f8b483a7a96889fb1b471185ca138df0dce6c6b9ce38729c06a4de061e072eba274cc0
z236e4c46362873211300d0db5236e6513ce274b84c552c345deef064d975a705d29b1cfdc5c4e4
zcb48c4f3a153c195eda9689e043ebb7b16689df3db6eadd2218b20b751306a4a394fe0c9326294
z96d6d9d7ab40538094376a735987f9b122e6fd164ce5754fadf6de7526579e857c821c1b95ad41
za979da70989f1c8aa1e36046ffc16d28fb5d65e45ce25f9ddc57b2cc914df3ffda32635d1c0fc1
z9ddc041128356004a8cadc9570f43cab1f53f1bad20e7bd90bb8b57dbbf1fd4f0984c4ef1822ad
z9507dad379361fc7d02a08114d15ee2ebd75006a0aadfb9f13811e4800da53864fe9d24ad360f1
ze8257eaa744ad38a8f1494788a4200d1ff34597d08f3a665488ffc88c53b6075e0790228793d8b
z4ff3b597e5debe0f9e43dbc45492ba435805e11d1521ac6e93b1b031a340a570b526458e3638f7
za47da9039e3b9fd7d8fedc8d38d87278f224e44315584d6343faad25903848e0662be2b681fd56
z1196dde47325cea3c8e4f72943173fe58ddd4df8e7801d6c8153ea6e8828e16596887a93697e28
zd89c6889930377b260e3f048a04a9d2cc8a3bd8a0a0f0bb7966677cb7b1e4e921117c3a7ba353c
z4f32c049ebc47179ad50e8feeb564d2463da0e34f423cfaaea598e89364161bddd179feea8ca2e
z235f7d1534eb5df0582514b0f6765270de5818ae5ebf325491535c1a559a70da09783a8c350251
zed44dab6fe4e6da5052802a2a56e6c12f3a14554907a81550287374a29f4aab9c4540289c1eeb2
z1458faf9906c85a92b2a2f2332e7ee0dac11feb07a06eea4665e6c2af728bebe3ab3218ad468a9
z91106215994a4c4e024a730d86005168272d2c776c61ffdcf409d623f0a70fbbb2b8510b318fc7
z406795b3ad75a3520aa9a79dbf37eebbe137554aa1802485f58313f4c78e0cdf2dfaa198657f75
z12fd3d8f54b8396a8bb46e6d28037bd2133f424c6ba01abe4b890c5d1d9f0478ed195a01dc6ac6
zd2949433a7aa5c62bfd8d075fe53c956dac385fd8e09b43d881dee5fdab98bc985a656c59fd235
za41264275f894c9df65c54ddabe9e69025e2aee5938aab65177565e269be11acd95c142d421cb5
zdfcc44b70b74acc0ad06d7d73237ea55b954fe042236ec935a6e8934c344ef16a05bb96e92077d
ze300ca4ad914ba9b5c2f06be0fd3c733f68272239604475fa5dfb3ce4565e5722f571530340587
z57a151a2a37cd378d87334b6606cd8c884f04c0747cf4e073847a5cb4fca0af299d7248dea0d6d
za335007ff821523d7dc0701042a1d4db322163568b3d615d7b70cb58a9c0433468b7e44b37dc99
z0a99ee9707d05fcec2946baeff538c18f79916ab729e197f870496f34ac727a61aaa05b35b8095
za899175e02c5e4afc696684c076b47bf1bb26a4564c5c5f0eec41f2512d2e7f03d322022aec722
z208dd9e651e02e89958767434398f5efec0c35178ac8acabb123cddbe65bc2e150c211a678d4f6
z8c13f83a98affa4aa947efe126b85f309eee3e57aa1cee92d0a39deb07510533edcacd314e050b
z5ee49cedee6b7260e50196c74d09eac1adc37e2b4fc5067153bf90e84b366b38110bddea4d09d3
z96fc4179db43e343e53b0982f9fb94c559546cf98009e91516caf668fea63bb50819ead801d749
z6f3b1a11989b433b5a1588c40a836ca8044e7fe8111725274a8649264a8d852a11067fb4a492dd
z14f2a343923d13db4b4c956cfd257210f4a3e5fa98c4888394e1e95d75ba54dcfcf782600458a7
zd23116251c36d272cbd256027a1779f1b065aaec884dd5a98eaa77ae6c90db4e72b1822d045e14
zb88f5e9ceb0a81524862ab6b64a4cbe99aa4e25db0539bb5ee16f9a586ca20d3ee64fa3070a17e
z31984ea17e9997eb5a4a5fb2936caee826d9e3e28905fa01ca274925ce3fdc853623d848074252
za2a388d551b399ddc8149f1bcdc32a6d8c2fdd5aefb5bed0e2a92dd44d86b4cdc2fb6b77f48447
za891a9f986e4fb7a1d15acd28c66a44eccac49245d43d7eac4aeef348d85201baf846b9d797df8
zb6fecda9121455d12364e7759e1efa69ee362e27c7585829de756002bd2999e511b149f2a53c47
zed8cb43d57fe686a7a95face5fc9ea2e6058980d06c7f7faf3f00098c597ecca37271e1064ea76
z93fd0bebf6f4a3156cbfd3e9248427464da3ab3e8baf5f9531952013dbca68d06b6e88627d0be3
zb7e1da1a7291a5fa450e2cba5927e84fcb6334e7e4d4d5ea405dc51bbaa5e50ad173188a1a3d24
z3d2436cbfc4bf6082cd70eebee19f126b4964ae184943b2e9f793f86113d5936666807af50e821
z3cad3b90377c865772de85fd7e96c556b755df57c864ac6809a74715b58be0a0b404e5c10164cc
z1a90076c027932e4fdbb882fa6efa85e24765b9b5eba8b96c9646f663f9c3a4b20a21598bbd917
z2c6f372c4b6579b0310bb1a03a64c73275242aa62a4226e17627a1b1918fb2e9f1d923ccbdb753
z540a2e60415c9968645dac29c261d25b5308a3643cccc4acce752c664c7211b0fd0106a11d9814
zcefd4b56332c2a2d1c8f5309a9d33858f1800a2391a0ff2f897fa975dc95fc339c8b7a2ce4ece2
z0a4c0f2c699d6035c56d460b12bf9ebb5dd6f3be9482c69dfcaf70218a7633e4dc226afc3a1305
zc71833fb4f7129b4a1097c74318b0493668666e72ef9e73f5711147b6be2621705f78b859875d6
z8cc294517ce9b7d9aaacdc54be7a854cfc746277eb508c40fd6facfe1a0ba03472e26294964591
z49c6703651ffaddd690b983a4b34c42575c7712953d3c5d7a5df9390a57f5e568d279ae2d8921d
z61bca460754641050d5b3e920fb6e94b530d47bbff036b0e0bbda3f067728ab818d77133a2a76d
z46ed41ac225e989e9c8164c0772e4ac6bc65511a0a38ea067a52465af3266d11b3019adf91e821
z97657a243e07ddd69a4f2a5bacc7683bca2417717e3e680d61235c787334f28ef3f6718fd34818
z547d2e03157a8196535aa922b4c22345a28b58b662029a408f3eb127ee9aa0e6b8fe2a0013c4ad
z871618ab9742d124191676de380358e6964c5491ecceed30b4bf38a530d2170a31f44a0483bef2
zcc5f17633276289f186fe579ffe35cda8adfe5d6ea83528c26d5c23b4565c8435807a530572f0b
zd4faac471c4368b3a84e7c8277e9cbb373c3a331ee98f87b06efe1a6582b93e9ddd269ff22112f
za7817437441c9be450e9864f6a0565d7ace67299a75f9f3e99e87881b5611cb007c39a03fc440e
z01a6fdefc1070587c2c11416f90ed57bb38e3bf4169cdb25593a7b04b098cf12a7c0adccadc6cd
z8b7a4f73a53c2f75c8233c9a2943699cf7d1c8482ab65917fc30533819dfac286e16ef06d6ea13
z4873cc317891235b3dc345cff74e57b49b746f406c763e842d068b1c6a7e0dcf66679050a1aece
ze4da700c0404aa57520c5a9a678fdf9b94263be86f58df9c647afd1c2d497dd2058dbd51ac91c8
z7b82d266198755bc545035a0e1c471785442db5d85f2f5769ebfad9be27c2a234a4ac6c267e168
zb5fd71aab8e1570bdac5c4c27fca1f7b9fe7715930a67d54d40de743afb62297de58d1c7c26940
z54766fdcac4c4f8e34055e303381e3171946cfa668ce8ed850ad9d7a530174a67532bad2eb75e0
z511cb26b125a8f8f9640723dba2fb306c351b770ba4326274e8b5672b02235207c7b7adf755c08
z7d28a640c7034701be66b5a2e5ebeeb1855868da1df6d1eeb28e3063582b6b7b61b8a45bd9ab6f
z5cbd2d4f613200b203294932664b493fac6f3cfd7465ebaa6c51a8648abbaff573f57388f60507
zf72757886d1d6b4bf7fecaa420c194bd1b904a1aff0c3f4d8e533fc9fb18cd3d6fbc6172f47c96
zcb4ce7584da7d8199c0e43a32f58ea0c03228af29e8a553bb257dc31985c5c4964a903930576e0
z1b31b028e59d6013b3894d35bfb72c359f30b8efa7dbc80f2f7252cc68b353dee734997b5a9fba
zab74b9ed0a97f423a815580100c56a08af9fcd08eb76a6804951af49edf13f0853be386e80bdb5
z22f909668458eadb08778ac6b72874adb73301b1b71bd8b0f17826732c232f1c88158e566ec828
za095faa839d0cadebb2610b405e49c532e1d45107376c687fc2ca849b040c318cd162ec19b1af4
z5aedcbd9e000ddfaf0370364c78b7f822d4902358523aa45338036283d99c0782f72c6b95a69f0
z4d33314f9b4529be8c8bd6305c0ede0fc3d37200a2a3205ebda5942eb30ba15eb77e5fbc6c57a6
z7c068e82f6925f98639da23449cd05db2c7746f01c3e23ed877f85421ce7f31ec63bb27560505c
zaf4e8334ed596a948c525b5716b9a2b4e268e8e4fa9c7b39a498d6c639b72aa5d8417a803b8582
z4530a88509da1df2b78b86558b073d5bb9006621d83a27666620356711d35250bf2fa579313ccd
z7845ff10d119254e5206cee2d73e8d89edfac2f1fd21feb53949309988ba28c5a9cd78d04431df
zc1ebc79366c832717389d88e4e070335021a0f036f89ee1b7b704adb6fe54baabe8a19af843a82
z4a401baa6cd27a64df04ef056aad755256fd385641543746d42875cca9969680b5a9a34f40e53f
z79f886901ab78f38167fb4a584ba44e5308492759c3b01bd9aa6869bb19fa636f6ca1071028137
z4a337df4feadc9ad28d39bf2181edf2ca349df2cc6a781fae5bd25fe3b0dc704572b0d01ba0401
z419b935368a73292e76e89d62d7bb3bc2d756dea51b61f7c1329672ac26192ca87f0f31edbd5e6
z9a2af301d1ba9811eb85afd76d8e1dac630faa47da7c2c450d7dbab2021bbbc032e8e29c637c7e
z0796c174c2501b4f195ec61eaad713ad94d79bce4d93644594db0895b244209ca6357506fa7b08
z16e74f03640661592c86bfd8fd96eb12b91a9524f1f7d6bcbcd14a5bc2f2b7ef98b181a623e4de
zb020905187e66ce49304407e0265528318b2821d3c142c4813f56f27fd2a7725b90aa665725803
z6f59580333643d13e1376508641e2435a485ded204958ed015e38a206fcf96a1213cd552d2db7d
z436410edd14b9a3c2e7dc3160f1b336dcff60356d06e5d888fed9600d0088e7a82b98bdcdf6c26
z11cd09a3cc9f4af506f71d101c2ed0cbb2a94af6e538add2d66b8d59e6e88c0ace2c6fb80d3591
zf06497ec1a1dc98ffc4b1419b7ef30d0fe622535745d25ed09419416822d03a025e4fb66da121c
z9e989cb340a160c6bc3e069d8c6692c39b2c8aec765971427f2c4e6133e5c163e05a2f4a4c7dab
z3ad78bb14f4deb82365aee3c57c8d7ee8680beae3bdbcee14537a7bdd6e58bc0b87521c0816c3a
zbcc1f829822fa6547f3bea6ec080dd70595590d0cd0bd1c082fd98154cfeffd6beabe7d73a6ff7
ze38f7260a19ec0a79ca6b7486d89dee71b2d26b8c34b63f33de7982dbfef8cb94571fe015fb654
z8a88df06c9e70b121e7c5e35ff5fea54be7e6a28833be721d180e788bddfbd4c31809e93cefc9b
zc2bdfe41ac15fd8936105418b61dfed346313d42af93a33c6cc009d9ead5c52fa8096a29ef52c9
z443f92305b770fb34cccccfa71707f0aa16f9cb4742c7e7e468ade9a0b96e2af00ac78816942c9
z802302f8b900c6b153d75a4a1d6a95d81b5fb5154eb6b809a19c6453d36654beaacc3f6ecc34dd
zf4873a2cc5113415908c49cf9fd71d970a187d2564b5c16c8f6eadc98f4760531ffc8e8d5a921d
z9b066cff773a39c9c1ac07b644b0299865b8bf1e82e7488955c3bb87a9dfc281abc6600e45917b
z1d68a46e74d38eb69cfcbbe60a9645aa42b14b30a5f186b412f26a8fbf2c40c1c935e88ad4859e
z4ba5cb797b2f439e7ed57077a0a6d33e0cb533d51aa55df33e9f7408b9ed748a512734e206e9b1
z16d5bf97b95dd7a7a75cefbc83c486e448d340866ed8059fa3f9e8d0650640748c6fc6a14f28e0
z6c632ed742bb9ed4388445b610f4b862a7c7f721068baf72e5a7b50ed4ef5944452b24e965bf69
zdc231d5a61de6c9fba371290144702031076e2f86b863d7bd5a3524a2dd534f3261a78a5c1dfd1
z16ea6ebe73c4f02e113642a4ff3b46ffff00928d24d3fa558c6c1fff068db712349ff11c8d183e
z01711625c25b34ced00cc31346b24406f796cb13eb844717714fa5126c8a8ee4d5d2d69b4521ed
zaa531792972aa18cb9fb498d55aaffe9ec37c03758d549ccdb4a92b58562432784d996d32b67da
z68ac7686a48f805e8cb00a2a2837031566d9594eaf7e31b1ba71c10d6a23a2a84e874f0b8e0d29
zde1cb1cabbe6963eda7336b6b6c733f8a6ed711093bbc411008594decf27e04cdf1b322bc6ae2a
zc4bb867ff9fd3e53ada1a57a3fc0c77d15a23ce099141febf925889f5f4d192034f6eed7ad20e8
z192ad730de4952165414c073e49db56cd21a6aaccfcd8d62ade2a6493ae770a326327c52daf84f
z1eb55f7d037c509743dfc16b97295506237c1d735e7fdd823341999734ad124ffa9253a35da4ec
zb4fd3d0f1ceef580f9954377c2ee85304b28535ee696479da4396593bdc040b42d112907a90a7c
z88eec59175e46571d7e8d77410cf3251edd1fb1f16330c9286961d7e7b4a4002bce4c21e73162b
z1b5f7379fc7f21b5d5c5120ceb935c5894e977d0dc243fabd4d24151afa14a1b51e4aea3775706
z411e24a429b2b4fcff6bce226b40f44dc41b900da895c50cdc43303550c8bcbbfb21f34fcfc12d
z4750d155008fc8e7b7b188376c9ef73aa9c9cb01ae902dbf41636b34413e29a3b338b714694c15
zcdb4604b36dc7084894f49360bc23a6d44ca7da994ad3e0cc2b53467819d7168c9d8064f6dfa89
z424077617a1f703253c9e71ca880062e6af12ea500fae79a92cf5f3eeec7228a7f2e117c074932
z616da3bb5a4399efc56607b01f9b1e5b162bbaee52a06d98735e72b911071b55d936d0160d83da
z5bdb0eda49a55ef4b72dee980927d497d540d7b06b879a31681917ed9a50a8a4f8cdac1a834a77
z43f7833e7ac230d8f5a7d27f67ed06b91c491112ecc660d3604812455667610f508e6f88f23f5c
zb79d03f54a78642fe06eaecd3984f03ca9625fa8efe093c756831c806f679f7aab9c3e4e6b48af
zcfa050d01449425e1606c716a48359790ea62e4ac3b88faf29aa96056809a9a4f91e931e988e82
zd08bc0f3a5e1a31d2541dbf28d9f7c5c4bdb0e3c8c31ddcf65d8e9d253e70e3dbb182b2fc9d95e
z8c0b1c2248b5fd2d4b3f8d693143d341dec99afade686892592d7d6f5241ad9a4df4d8594f8d29
z364aebd6fc4f3794c1c2d14f8a86de1abb879c93a778332ff6c5807115cffd4c294bf9f5e9f28d
zc305dd1fd3cc88eccc77f55891077b1fc1a6ed514648ddcb74e2cc3ee0f8e0c7cb863367b793de
z04919eb3a612946e3c592b8ab934179c2f9f1e9b894144dd1732ea50c280432f13a9dc0f400db2
z276603844d6db4c9b332b1ff5eb2015acc1af8e4ce5846c92d454a9737b54dc7153b6be45b834b
z76a4f87d001394f1fea3778ad4018c7edae32edaa59b8c9febb0a4731cacf8e2f3e876197c42da
z499f451120f0009a5d0b78b7184dbecb23b540519b92519a5f9c013b720d98223f2be21dd7543e
zcf7ec38a93029c6dc31532fa9e5082f124daa92ed56be68ff404600fa5307ab8ca2aee9b7d086e
z570cba276ee1b9b1b9e3c3a022cb755b0b2a170534b74d3ded4fae46ec97e13ec7be742bc69699
za7866b6333936b5cef0385baf1ff28f8f895a0ea83717a89c5073d106410578269d75dacd9bbf7
zab8c679b0670f0004c41cf9d23fcbbf999e22b48695f8d183a0135fd9670e5da3ea24ec13841a3
z697c0d56f06f463f90a35a242edbaec2363acc78630a73089c27eb5bd7b1124b0443beb4cd6543
z6be6ec4aac589227977c2d40285194a52cea0c8c208057e974adfeb9a2349f9ba5271bff60d2dd
ze77071a565af3f3246632632eee8205023ee1d77cec739bdc849796fb9152c8d801d9a8ca0d75b
z0939d588ff00c65cd7cd63cf87bd9551d21e7653fb10b851c7086de502b2e90c70827ac78ebd2f
z48a537fa2b78bc597d42dc5f03a63394aa0580c820554941e1b6e42d6f5fe2ea2e17581790df4c
z34f1ae14b23ae8d12d742e2eb5e4f93f24218609bef60f3a4c8857a8ca677ec199725389adcff9
zf0da8485f3c02bac43c6c595eb27442936a7acfab607017ccf5004be6ac6550e9c713d350e5af2
z3b3744d0107ce515f0c10f4e6ba5c475c49a437b1fd43ee7950bbac8eaa166112355973cf78653
zb2bfa0236d43c02d7595995bcf0548026a76771436de1d828a6a0c43ffa09cb142a19d3028e07d
z48ca7028bca89060efc23491ad5596af12eb1f7f2a7203b864cdf5dea5a5276a73297e6216db72
z4a3b11ac641eb8ac499d01919eda5594ad738e93e66862b44fe0d979738cf4a9e33f7b33b7e277
z3dcc6fc9d597c6a3a7f383fb68ae2fd1a98c22d984b57491a5a83bce5364676c231bdadce49ecb
z35ca58aee7094d5dea7026d2c5951d326b8b7bd5bb6d11b7f5521ce00060290c82f54fa944b14f
z32e0ff523b7205220db7cd930bce42b1b4650449715deaa4d94955f9c43884ea0554fc2bd4a171
zc208ddeb9e212cba5c70616019757d79ba6bfda2603435a0f6dbf7cb5897590e6c842b5274b894
z5e31a0bd119aff63ffcb9a855ec551072b969070482dd4b706514e70d18d11bcc909f5d97b7e2b
z9ac7a6983a621398494830aab50e5cba032c1293683f75909815211d8c80f4ae37370a1e5928f6
zd9d99a63a238215ef984ce064171872787bb18f470e3aa346665716dc849db995d70571caa6dc9
zc002f83f678544d5cedf091232302f07b49d7f7910c09d42a98090c78373030c236293bd4da94a
z4c44f17620cdbca92912bedbaa73aacb3bbc802fb1063f43745906db0a50dd82fb9d2d11bc410b
zb88b509b6eeb9d1eb09defcc4ac09590ffe1b75db0f78f146fa145292c7fc9f19879bb3d898e2f
za9d2ec2e2e178a5cc1d6f8ac1e7e185ab1864ef2a75b953dffadc4931c4e1aedf5ef8c95fa61b5
z3113be8a71526685ea751642332017d787b30717e0f34824a560b2395ad0ba50fb35443ca73f59
zbe82c96c71cf3d737e8b634e8e0cbdf2c306047e48f8352a8c937e5d872e9a19fc3627508e810a
za001f259a8b34d1d7e16e9bf64d1eef90f5a8b11527fadc1ee444741cd9193f7da12d798097815
zf1163b6a76453fc79373f17aeb3867bada68f6cb91b0d7154f44214b132a866f0e0ae122801990
z3d36d8f31a51b35c31518749384a3846c9c4f1958f3e14e00f7d7351af8444cfb1a3b96a4c40fd
zdeaa3f1d858271a35094cecb2e3936ac9cb0b56548930f50e718b8fe45dde6fb24103752aa6530
z25cdb2388091ef3d1da094add4154d72ca8c0e8c9d32609da9934229c209f64ed38d6e32f24095
z6c984fab186d1d982fe945c670581553a2d68393408bdc5f8669caf4950aee6ec7a3b7813f9a50
zf88610459b868bb68eec850e278549dbace6cf93952427d827671c5e94ab8303907a2a3facc73f
zcd96ea21cb557239e2a1e2d81f8c54e6517e7019faad23e2c3a9046ef6f8c1c3e92ef152c0b2a5
z553bab3377a58b8a16fbf5dd47197f3943fba3b4fdbdeefebeadd637dade43d7fa410e3f494b87
ze4392e902d790c2ea9214f23df4c45643edce73736a43315eb6662018b338d795847eacd1599c0
za7550c12f5efd640a8296d7b04078af7af76899f49425b39e21995a3dd2dc04cd8876820b2383a
z2a7f41747e309d281df3ddb82b9c12356142bad1176de3e38ec9644e3926e8804e6e7dc68e2290
z744b36022258fe0d7d21077f30ee08fea54919473fb0b5295831dc358a0cdc9c40cb4fc6220d8a
z9450ad602d355d28ca5eda56f67de52c81c33e954ee0787757b4fc135639f3e62cec573d1d37be
z6b83d76de8a73689cf6217b294de7de927367a7b060a198882746b3226ee8c3592efc1441d68f8
zaf9d2e472e337347bcfb177e15f8dba3e66756f27a016389a8880d0556aca2bf9840f252e70b9a
z84aa25b8d11427e132432f5bab5b18ed26a5100816eeebfb4416b0d77634924db5ab05781e4842
zd63f712e311081efc909d928bb05d9593aa5ae2d1fc53a66a9b3aeebeac7f7058cc7263a7303c5
z71f7fe7cc9a16a0c2931b709cd09b0c4cb43237604cc41b669db44902dffb041b6129e6b4177d8
zafda3a86fdb7b2d67959fd0215e273320432d468b1e5aed6a9e32c51f4175ae064164cee8c7c6a
z416d07b58774dd861449644599f3b2002e8f4823e1aa1c97e193fced302c5e338c7f89322df1e2
z09080ed6c0caa526c9eb70d033c37c25a8c77752cfe24a93ed5c7761a19ef75648473b96ad5304
z9182381b4993b3a34986a6f40cc3b190bec4de7adc598b7dcfc03e5397221a9758cc9f983fbeb1
z4723b03372a5cb75bc1cc69a4a20fe4373489057cf3b387b4eecadf904bef918d2b509598e7724
zfc61299489e5081d69017b351e43461eb91f835630d3dab00e27c3082100378a19998a07206a68
z82065a4bd60456b5e0f4bc13db3e8939930f49eff267ac1f19183e8ae5ce1659c75905b6c2a70a
za7c879d27113b2825c99b208d418365b46a8089b757931eea2d24257871dc8c29c7f69e6d802fe
z240ab96e7d3d816aae816e6ed955481d7238dd424d3806a43bb66d12e74fad42e2ad3e38dec6e5
z209602cd85bb4a52faee6dabe2710c8ca0f38979967202d7f1fb05bf8a12de6f113bb06b3fa142
z5d01c518da219664ac807f07bc4d4dc42ff72e02932332063591cddf48dfa39692c87fb06fda27
z3991652431152b5cf4693449a923455c8a6fa6371d968622ca118aeae1861a51554ce1aaa233c6
zd1a4351a7eea9546241c83b03e8c3a0493d42af34375959a9eb4379e3f46ded2d9e1aedc663d82
z0864a126d4a37675a9ed68e7d05cbafda1f2eac2b74c1d57bd297359122cd0e3ea536520351adc
z6f1478542af446e7fb36372071df73631f225f3434a634db1bbbf7cf504a4747d477eb4a872181
z7ba69f6edf5d55aa8054a42e45e77ba88bdd82430711169a00203d3079fd342bf4799dc5617552
z424d198e8dcc0b5e198b4b550f6f15779c2530719bce6e5fef8131995fa6c3f8b138f694dc6817
zecc499e8da3972c150545cbda6cf851c0b149bc53190819e188fb6ef385eb8ef774aceaea0ab3a
z22b3c5db0d3f23935ab7e1474ed4b0b72850b008456f69be4b45b173cdcd6e2a3a8bfd43998db4
zb7206e15314f18958242092a0bf72d74343b991e06acfd5b7019444f93558575419e68d1274990
z14b50707983addad22463a76a1036e7128dda02edd36de6ec44e4df21bf5a17e33520062e2e4c8
ze6bff565220c62be8cacbfaa6db66d9b330565a5d4917309c62a58e5f850202cb4e62ec332768d
z98f38eabdfb3eefa0909fea35189c922ace5ae3d2d646ece3b6cfdd769633d16d2ad065423f402
zb91621ef932da891f984431a35b80c557a299750b14f755bc57e7c455cb62ba0ea9fd2fa6bf76b
z0cee3ed08e2f3bad47992d5d131a036dc3eb1fe61ef11ec80032aa581c9d16aff55b14a2c314be
zef6bebd2f9eb9f3bb3902f4a59fedf4930c4a9d6a1cfd58407f812df82997eec5eb772bdcd11d5
zf2a3be99084961c09b262880f04e45a4498c44d57214167684a1f47339116106f1b091c0492e71
zad7d1f69bf23be04ba264c94d7c5d3df5d4b74a9f8b12d672391039a9554f42575571ad8dc7fde
zc971661045023b25055cc738c78019475446b0ae2ca1c7a57bf15a6f0ff69e7e41b8dd47da6be4
z9ec8da5d190b66036302375ff07dd3b76046fa1a84f16e09d06c00a4eb4753dad18ed6077ff950
ze7fd6f815ad26dc06f6dadc22b39907034c13e7ec00f545b30e42984fe913b8749fcada1a4513b
z3d186cf309322b1d8e9e4435a332dd98da2ad95952a5461c1dceb06e2be20336573d3fe1087b58
z2e1ee0e669ea3b828ebc7654c2fbdcbab77c01b5810f07ce2c4920a344b0ccdcebe04d36271a10
z07d9ef46705d3ecd2df5b4bd3296528b99485cf566eeddd9db41d330bb1ae3e049a410684f775e
z57aa6dda6a2249fefcd41d70eb96a3bf4a17f1f3651c9b656df0a2e5ff6bef8dc6aee11dc509b3
z1ebe83182ecab0fb7bdf0b27a6a90e9b6a380d8e260e67febc2510207415ac8354f22f850b291f
z4ad31269d83cad9b9859baf3b2b69a4a47b878676cef52107944c9720181c3e9ec8f394ce962a7
zf853eae0bef456b13ebbb61b1c3ffd00f8a4e3c70943a51b3d99e21d66ab982cd5574f369b9ab9
z3e6d9163b0390df2cb7971eb5e722112ce10133dd77f0ce1eb3c709bc982226b6cf802d177dbf1
z259f1e96315d03dd2904b3087e7d743d82495311f8de5c3bb063ca7c6659d127cd853605e6ab96
z635af3aaaa5c9435b4e31174ca91b091cf27b2bcf23044a622e26aaf2029800539e88a6c55ad48
z61002066601738a3160d6ca323e06808539c168f148efbcdac300ad43b4912bcfbe8a9821835da
zdf5206f8dc938bde45705e5efcfd12e7d2ea000c6b3858468b54cd98f1e495fffdb037a5f126c2
za7ed57568c9e6b449106b0739c093f03936abca877f8120359134ec639ca9c11996b2b0e0028b6
zb92bf375a75a98259be35c5df85a3826d1808b75c19512879b3a85abc5b5952d3dbad03296bb2d
z9e8a3fbdaacd4956a856ef3a0301e796d382735fa2b86db29bef46cf0c7992a5613417b8ef213e
zca677391c84a3d5f96ae542cdf4a74805a590a1dd79559de0cc960819f96b9ea49e2c1f05258e4
zdd61fa8e82f423697af77a4b73c729a16e366e7bfe860f6117209d9dfaa0a458bb386f5ef4fc2a
z7f0954dc6fd5b2780917533778e2248eeb464111d3b340292e9f442dbb0ffb2c5c567692f90313
zadc944791035fc3ea67b6b94d2dc014b04b9c73481ce07f0a619901481d89b819bdbb4bc9477e8
z31ca1cf060cea00bac4d231143a0a27c7f73972772983b51e7e3b60613d63e5c983bb647fa2788
z40874d5cf5b8d3ccfee3e0d340866bea36fb427dd3f7ad4fc21b0de4e9c81b396f2b2c0305bb8f
z22c97a7875f6d8edebe99d6b73c6aa2c49e3fabcc81dec398540551ceb71de5c424f8211b8dbb7
za338302c62e3636252c6c00e472236c6b89943de09add3ab2e758c73be4a671ac6c7a93f2a1c67
z361722d6d87950fab437d604d295864a968890e16bb12fabaf7b48605f08dc6d86a4e214a07fdf
z96c7cc0c480d33719b882db01c24b2ec71ff6e817a051cda519bccab3a0cd564d8829fa76c928a
z06cd465e8849ed09ec9a2b828f433045ae7f0d8647193c9d24311a0ee85393238a4571f8624e8b
z27e0bb969c95390efa63c3fae157e97f0ad693ee526676ffda6197bcf867945846cd814977965c
z0967af86b49fab7856a8283b6416cf057f6faadc4a31678a61180f4e7ec4640ec587db9093bb08
zfbb6cfe9954895e924718b52607a5b00e29aa494494fa9f05abe062589474e4c00a45084aa291c
z05a9b1ccf85a8b75a2980bffe04ff0fc8268fddcd21b66709b63c86f677f1cc38060648163b808
za3fe1d4ca2de50abbc2f875a67871cc1b42c6049d76b4fcab1ef87c9e64a22b593ea8c04bd7b97
z57e69f7367a41ce0222a7237039c670535bbf4e7ee63a36a7e4880dacabe142908eff41e9c87d7
z9b411e800fa3d2ef60db569c2e826b585785e71748151e5af0c39a0386298f7780a8d8529efc50
z6e17e022ae2682046a21412fa1258d111ce2da74e709f011aae4f19cbd0857db4120edefd63fc9
ze9640ce782a1b316afbb614fea7609c07c0343332ac0abe4374ab86eeb6e2a21ab84ecaec72c5f
z8f5077d8d0780d3ab511f26c933c77fd665afa7d1b2766100a7a03d401e236403ea81f33d32646
z0cb93ced5b28b6c992a36d2f43ff5f784953d6a8b9dfc9428a9f8bc1fb6ec98ce1145c25b7e24d
z8c5725bf917fde22a5b1e3f25e6467822f28169d60eedeb5cd649df22355757773c4b4c4990355
z0056b9e89c3c5ba08efd973a91caec353e353d8da47519c9e7c2466dfcaa737d3d149a9a4ad4a3
za3a6c35da18a4c431777e8909c1ba4804eea895f0fa17758354c405c6b04442adb28348ec94876
zb063d58486b9f942cc7edff60be05906ceff6c58cb6dc1c426999a465a2991d003b9c07b13e64b
z69b80ccc68eeb9d3ad7a04be64020c1a08eccd3f3ebedb3962ff0826db723a0cde4a28f569bceb
zc0a9dbd321577f015651f078840849278da7a13ab6b6b0c2e8118ee6fb9ea670ab855c7ecc4915
ze1601077d16094fa048d07ec41b9092bf6f6d59e90fa23f391bea045236ac18f7467ac30058e23
z17ff1b3f91310efaf031ecf8ebad37b29e8d045b8754dcadbed464147650267eaba4e9fbf49349
zce0e9e90dfedd8b1652a6733907d5a2fb52b72b2e5190bb07dbe30a396a04213f62d7394c9d4eb
z0479b40eb62845f1fd1fde3c65e1b37ee1a506a7d3ab5887ef9f362c5d8240ffff90825721095c
zf6862e71218ea5367dfb5360536c2be1fceeb1d4b0e1f6459c287714e1905008479842b41e053b
zae907fdcd9c24ca62d8bea41c79521aae479b4f10fd1853f3f98a7441ef9064d7edadce4ad06fa
z8375fe3eb04f33cfb272f517cdac723e68492a590be5bcc69255177229bb69babef56c215edd31
z915af055938f96802447647cfb469272e3f96ddd123c3f1de7fddc0c3a653b52abaad13541ce2e
z13a167b6b0fddc4b29b0a9a85ac0cd01e129ef5cc1976b6411941ac75cb108b49135c7a9c05eb8
z983105d80bbabb947c1eacc5003d6089a68a9722d14fde772ae0a63b77170162dc49911c38711d
z1766441ef49ceda3fbc2127288c50506d58324c0591f757a0fdae7e827db67da581b073408b7fe
zc009fca451ce23608121060c27ecd57824de93cd0b2f0a2f990c7cf5b774adf15a52d3140b87ef
z65b68b4b74b0fe6f86f9031eaea8cd396d87a119708477a14511e829c1008016904f16e63c33d6
z8737ade12361cc11639e334d4e504117a51889f4b265fda1593bd9984cd083b1300c72f4183ef2
z964ceede77f674254d2227777d7ac6c21c366d8691f5383be1795237ba6363270fd36fed4e5aa9
z63d7175c64a6cd3fbf4fdc49bccb34c81f3f89b83af8944cf5a969493209933f1365483431ac82
ze5b08737bb725560b66fb7a1a9aecaedc54567a72d6f002966d19bf352b7642ef2976b65bc8380
z5aaa5b2407cd6ba5f4059681e9cbd0c9fb91233caef8d826778aa95a38866781d7cfd8250ec893
ze07c979de8146e6379b8110962d9e6e992d9ceefb09f9e4778f4a78a45d038c00fcb1294bc2397
z0ba5b389f92c4b374b287f61a6ccadc4f018361f4bdbe1f717a9015b3560f73cb290dd42b8c50c
z4681739e034737f37855772869427771bd922ea83b8042e7ba97d5f07f38f517800b4013fab0ee
z546550b4dd28621558272213c20eda18242576bf0f26b164753773cf784aecf4abaa97d164c1f2
z45e997b14ba622c6d33ac5a17fd2335cb38f13d843e98744e45774281dc19b1776088dc2cbe792
z61efd66848b5f3863236189b060a7552cb09381aa75f244dee99a1697734a45f4ac1a9b831ff63
z92a6215e13fa6d92bc3959d88acf83f05b87bdffc5ab1f0d978bca47f05877195d03002b91c5a8
z3091e8bf912a5f36bd3dedd3dea2d732b771414ee8c9d67c3b1e12205ad00725c8ec56a474ba1b
z65f46bf35a53438b04d276be7d1c4c2773a9f6daf709934301b03067f22b585a42f9464ca9386e
z0850da8bf4cbb3526f3ba5b8a65837a244f55bbc5398fece8a5ae59218d2a31bbabec317fd441b
z244464cc458c6e4dba85cd4345b20a98a2f41ac6719194ace2c78112976fd6df79b7cf7a00c631
z0e2018019ded73c33f19434bc67f4541a3c83b5df56e89d2985e0612bd57620d4630848870c633
z5e48064eaf4974be2dec3f67be9897edf9cf628a139fa848200b6980e003b41da741d2921a9840
z1e00c1b0bff4942af09ec5ef92f78981a4540f04656ab63b58e8ec8de54e06816edb0f89dfb028
zee745b3a22e641dbd571924e70e0b1953ec54565ce60fccce43569d1453c52a3c21f9152240641
z9cc1c407df162b1803621d53702c9f10cac1aff858e1189b28fcd05ccc1e21e01bd5d1b9b3e73c
z50ca65de1137c4cbe24f6097cfcb74700e9d991d46b9036cc4982bb023edb65b08d68e7bcd9122
zed8e739a47a2a7eb3c5977e3d794bb8613bd8f910f26500c1e9c322e764445337863d33947c881
za30aa2ed5e84642495c88acb36fe178a0818ff2da1f35ad08a23f37b7a0f754751061acebe4854
z7f367f8c42bd7c46bff85fa053c8030b982a07ba75f7b7a962d1838b958146ff911c03f1a13bd4
z16e9cb6a66f3539fafc5a65a71f83577849fcef1f9990d8ecd9cb0ba90b8aef6bd1f8fb452e288
z12293ae4bf96e1db5d431070dac5623d73f1ed763a759a2595e933fdc6bd917f5e5bd384cd337b
z29f6e33dd93e0c59e3990cc1bdfcbf1169cfcf47861ced77e151e0c2696daf064f8d620de79456
z2a2bac91c0bb07be10d8d81b662f4f5f6b66b8ef35fe18272383809bffae09c3e9e23b0b8401b3
zf81e5a50fd4b3f2412a35e87e834b0a8f4a60b13e32d86bf74a33e9aed7dfe22a10d17971612c7
za45c3beed699f9e8d96170cfe4731349d2a93733f0618d7b3717e3914a2df1bbc65090623ab882
zc97f2c0a3c6e4a77ccbc4b0779def1da473533c45ce40f42e93b43af6449a1625ee093c4d4df59
zd31fc7999f6de5e97f775ab8dfb25927420b4135e7604435d309860a0c0c49b50c70978d8d1ad0
ze6b6f3c6156432b227fc402c0d1d2092a427a54bfea58e984cb34773e63d14d1098c90f00deb8d
za608d5dbf288d254451cae816409b7f5cf31a767e1868280f24cdf124a5cec7b72b9c30d7457b2
z8893e0fdab720864c404d8689fa8a11a80d5c3251e34cd5466948db48e29f370d91a5f547e5dd7
zab6a841bf4ea6f47eb888cb405f07a2817379f0bf9d228ddef5911997f5e8aabb2509a65708d35
z3848edda222ef4a4232665a182d606f6531b5e9acafa9e1df7db0746aa90a7c2185e4a05583d7e
zfb529a1c2d415789cb0deb792a068f34251ed24f8c61f1e9417d66bc008308a82b58ff8a126c7b
z2131a777b43b5050e0df2bf2d7de8b1669cd6863be1ece6972112d33e4f986b528f1082153a694
zba8aead7c4e599b7e906dc56da5280286550e346ff9151b2728b701a30834cf1b9cc32beaf4108
zf7f1c6319fea9d1b659364f3ddbac072aa7fd4ad8a9646c04b897e6592c6d10a4423d9062f1e92
zc42916de88039f178638cd84637941061f24b3046a1c08cc719f8bbf5f0e87d318ca6ca426a32c
z9910cfacc192222559d5af88d8059fecb6bd22a70e6b1a425302aead7a53a3dcf7fbf69e8cb32f
z828940e153ea474979b3be8d426ecd093caa07d057f7823df7d45cdb5ddc3b031edf8a01c837d4
zc3ccc722dea4e9a16eb95ae97ff73409874a34a1089e84167f25134ffcf0341ebada2a9aa32448
zdb8d876579969727c896fe5ad708f1ac1ba81d4d5e0ced3c8f7bb0463a66788af0ca42e2a9b854
zd2cd896396a99f61c9e378bbf82ad9075881299efaad7365d499caae9d512eb3e9394f2e8d546c
zc42da738e2dffad9ee687aafdd609b728d1ea6df93da10adbc3cfedd6938c061d8bd73d9aea107
zb1c6ef4867d3c5045e5d9bf9a52a34cbc423f046996e4374c5492feb88972d7892281738a5dc70
zed633db573c064935aee8660dd509a6e87e8dc9a6cb4fdf0d1398abe206de862c4fdd1dfcb0d34
zc24eaa5d98ac0d0aa9d015d1eb83462b182730508b2c753cb441052592db5b46a946480c4c3ecd
ze6a83babeef071c985e3bacc18bc6568fbbb7f8eba8af8ee951c14ae08b47a5ae0dfe0934a7c25
z0fb66eda5499cc0c9da8b3f0b7dcc397fd0e5274b6b4db7ce02fb3bcaab68553a8024f15e27179
zcc42d815bb775ebe1dd787aa01e55cba5c52bc3612ef003906ca62df641d88cc45ff764c326ccd
z26f63f3db120b6f093d462e6743c0c6e7f2c7e305f1ca24f338e7040831a873eb575b83a22686c
zd56b469419e9e4a9dacabd38ad42d5c84a23f47730da5d9f33f91caad4dd27f22a638f9268bb09
z4ee170ec6f394763b07834c59fe0641660cf2987fd28e48bf1e178a689ea787d2909571ea2aee8
z6d2e07d1d7e338c35d418b471803d7badc3e4da1f26f71b98e6e73d8b45ffa5153268fcef0a8ff
za1225ccb937973da2ec9e8d705add102b95f7d31f14f4ea843ace8acfc6d17b1df156e0d97e51a
zdf4030c97a5e2fcb5d4c9c4d8ac022b5992de14e91d8673bc0addbe283f5939471596f0ec5fc5b
z69d0241931a1a7764376acd30a4714d1fb0a80e5b68542030b1a53a88196b76329c3674c8a7743
z71ecb485dc8fde26baafe22fa0396cde0d6c3db18d5c36fd64c55c5151eb561c8bd91a30260bea
z480d23357e717e2f5c4ac810ce6293d0a521c252ed104b9db360797780d36b88a34d72f7947b7b
za88388f7586d047acd5b97c98075aaf372f1f60cec6c7d36a4c0f7c608f4f854eefc39154a9910
z7a9fc6f32126dee7482281a0cabb3efa9ae53854bcf16ecb8764d8009effe66569445c20630a02
z7b424486a96f97c14a56c6125a4c07a0498a6aee3d75f5da8dfadf23f651475df394ebe3d2d503
z1741337360a620b309919d4a9fd1079ce415400d919587696914b0cf27b9802ec6cf210f911932
z16f5433525305158c8172ce4c8cb741462bc2e569e74b5bd30a726b15bc43b7590fabaea9840ff
z9cf019bbac576843fc796991381473bb03a16711832b1c736fc7810d3fe0771de7c66928c8ab0f
z03d52cfcec5b1269579b568376349cc7a3a46e56ea5ba794d9f650c1e356cbb4497f67074c183e
z3df72c8c35a3f5ed03a5bec89b0f80921413fce83899cf8f58a8cd63cebace6da2ece8077684dd
z434942f27a11b2d96430ca0a74a7e4dd2282a35ee29fc0761f54e20057cd0f62808ca66e361b6a
z45698d4c0f1bbc7f9025443b12bc4304db5cfa756191c306f063573a2f13ff5b8c5c962f319397
ze28c1090d83b8558124551237d42502ef39e9549da1dd67c38e4728b9fc8b5eaadead18df3b551
za469d03c21e6492768ad6c627cb35f35a642d90b61b9d4db1e555d358e6f1d37428db8e3ffb384
z4e145064e1b8b060c0c72ab48cff9214de629986178dedce2024290e20a091b0e53d4cb005d658
z3a55c1e282bbbb4caa3adf532d198fd88b984d22d46261a2e35fa9aacf32d92d724ba861dabba4
z210061f15ae21404551de1da5a250735c9c1553467c4ffa58906f4388008905b33120b8deb9026
z368950cf2c16cd4519b72646fa44b9ac9796932744b0efd55126863fde204ead912e2deb77f26e
z48310fcc7ac43732354b802b4db83fec632075013148746a16f46b9d1b1d6a491f1a8f2e6b2e56
z14a233e02308d485534fb439fa4a44ed807cd9a94aaad65484221212e806ba535ec81684708e38
z3ca3f5e60ff47aa853779b9d69620ee9c9efe76f20c7b9277f0991c73cc002528fadde7fd812a2
z111e57f929e317c872e24e15a822cd79800390ca397dc698357dcef5ca53407f310cfa62b0e684
zb454819166036f2253c1d46525266bd988c831553aefff5b431eb9cf523ac06cd57d77fca6616f
z8cb9321965f3eddec1d3e3c95dced9123ea921d68b1ff1fec23665b0a75093266bc7251f92e69f
za4158486e724a26bc1361c6971e2c032a361bafb863561e10160159bb03dcc633f2eca36b6d5f2
z77cbbc6b5e95b1d3eeb1c65d419fd085c9259cd349ef0ca3d7555b65b316b20931b3a4ea648497
za77485f2a7f837f55d0e12218b0bdfcc268c90bead962af19a7de0097da387b94b25437c42c7eb
z2a86f96ceb654be68c9fcbe9b683c4fa6f267176aa74559cb31037d843cc4e92b87f4d56171481
zb246c039dacea40daec5b101601aad79c7d03dd4346982d826e2bb123efe9c7a5cbe20803a58df
z705c1444305846845717b51fa0a84bb92e02b4ecb7a7fb02dbc5693811c640aec6003fa75d7f9f
z1b2a54510726d7d20323279390c59ea04d6e84af29543e14f5970426372f13e8263e0c627d0f5e
z794a24c7be6bcb406812b5c15d1e1282259b3cde7bc73c1d7bd1317c2352c445735457b8233b1e
z274593338d3ae2b181396a2b7bfbe5f6ebd5835d4f7e16cc2736fc26aa90afcc86ea69f9d277e3
z313bc5464a2ade911f29c0ff48baa6bcb017a78450a96efb5133837a18e183a23d7760b113b551
z657e2f489bd551c2b5a338eb72875d5a121a75af04bc3b867e8d8fc6455f718b4266f24f70b494
z3318cb09134bfbd9d98ba2ce7ce9a43cb94b1173f3cfeda6b492e69c12573c35fe2ee42d3cc41c
z6a56d88bab00aea0e3eed9be6e443a302b111db68d63b4977441bcae6346fc323676cdf7879704
z4b201b6d6c9607335681bcae90f72e802328326fe2441d930ffe96d852d0ddda6c32e2d13bba2c
za03cf4a29261957446d37e69f79caf90824c84e6b4bdbc683f0e5773a08e7745274574596cc15b
zbd547e6ee6ff26f4f1832a2571aa728375f8f58f4e472df6b52768233fc2a3e41683b6864f1a28
zcbb9105021967564ac8c9335ea5f27aa6eb30f7f9bca51ec5c127cc34afda0cfdc9732804270d4
z19f680bc112e8b74b1177cbe61a7e0426edbe85acaa96e8fca93f0f66d2748e78c12db1a2899f5
z35832a13fd48ad21410f4f36f847eaedc4d61b04b558c27d87a7abe56563bd6b077117b6d17415
z3bf3edf6b862784c4036eb8538a95cd242b3345877d660a0f0c5df45743df4a5a7559001308be1
za7ccfe002208d066f2e6539d5f9755d7294b3273da75b58643d73a3bde50c0d14f16366ea045e8
z48e72915cb12161de8ac4977d31e821ba7716a8acaacdd49baf92b77692eb5c0fa70804ff24b49
z079ec0996c4fdc47b3adacbf328e14841f56ba7bc3b8dd1932b5d8d12bcc77bf2ebd9ca525b827
z7cd505141dbb96ff8962ae10dc6b8ea9c4e47928e9a47947226774b4c75d2187217e514b9bf216
zdb8795b237bd04bebe840e1701f17bd79bed365ecca31b9491d940d93655344e8d2d7e52ba1657
z1f967fafab4d541a5e1b9a8c67c190b9e67aae6c76ac845e5f9610f43d860bae1abbfc474d2378
z3b94d29cb78a56429493ff105328f54218abede60295c7212f74c2e7f74d4dea994433fb08bcfd
z3fc4f5dba5d9889976deac0d97ac59e41f307181e1bba5f5a3ff05d0d9547ad1a3fc88ffc6523c
zfc5a84e4ee16e56dd5bda93dcaf3f6c8599b3546e6bae22fca2001bf5c944869a0d1786e020e68
z91122ccd5deace45870344a39c47bb4d6c8d1ad7b9db17601d8397e80a40fba57f1a39d72b7852
z4b1a3fd29cb97967039c515fdb1707516481c13844983d00f21ebb25f012f3cf8ea1f5b8fe1e26
z1c5fc7cc3e8e9da510150274cbbfb4a9b2266a419983eafb4101a31cc55ecd990aad734786c26f
z41edeb12dfe7c3629bb422264f59dc41ba60e4b58dd27c44882e4799572c9100840e043c35cfed
zb3b66175bca11548b73c44cd71cac6a6764aa4bfb41d21459105a512bac793f91fcef20cf7cae7
z72bd4947bd4045400297a674adc19ec837803916510f33e1c17a122e8eafafb0c2161d6b932460
z358f8979e564dcfc6dd5b40b670254fe5011ee51f0b65c597b4b0d78f4239320a077ab71d05838
z3678ebbfac12a997d7bf94f518976dc4802be5a7632565c7b84e65456ed3f277436b88b9ab7f5f
zdb71faed0dccb9e7f80ca4475217d7d331d751122c8b7a5d5405cef9e1d63de98f4c1ba79d180d
z953e5220676232644744ea988c5d7ec9c286065e0a5a369afa74dfe03da8762534a7416422ae56
z5f82c748859588bbf2280977a11e21fb09f9403bb0fc1fa531c3689da0f900b48647511965768b
z268df5f6bff51f9dce72301d94c8edd68ca326c5165d06affbe41eb286674ce62b1747a81228a8
z6494894724cd3a86a5df3ba00339e53ae435cc16b07c4eeac03dd611b76deb3bf9f96d9afc9d34
zfcaa797aaf05829d2fe210216f4edadc0fba0e30888f047edbda2f4edb76086b2e2daaae8bc31c
z8b51a74e163344b5f72d48a0a696a6328293cee8e4138ec30a9485a7a6d8ed10b71e4467ffe3c2
z39a863c44ed91edc95dae542be728c0b18cc184e64d7489c7017efce8af9bcb4ef5c20717c0a6d
z59a102b5ac4885118291315dcf6652928a29ea88e5014a7ceb94e1462d7d7848d8d17f8701dabf
z983b45f9106315fa5f6da629e4f0374041f8999e5627bf229f9a774f7f462713733289c6e4b48b
z967c3af6b0eec28eb62e592ae560d8742be24ff77718c85f3a36ba76fdf9c5737a4e4dfa8433df
z9a32f46f4b58a7d2183552f9e9fa07e8671e8661227204bb36aa4809a4289d1a3ed9bbbf458c6f
zd88ca2f2c5bdb7f28666a8aac5fa0c0732e959be182c2e28996a4806238b6d014d7c488956bf03
z0f8551cd2d06faacc70a443fd7c57f5a424e9a775102c8960efa3f6859b76747f3de833ad1531b
z3b95ee8bc51902160be5ed1730c94a596eb20e68fc031c53750ef65860e41a36846f99dbe58cbe
z878f7a06e11ff87f77b6e387f39a223948ffd9247959529d2a82187754fe4d0cd08b2253475b67
z60a6cfe7295c91a5d91d3215de1a2f0a60febeddba442a2a838a0bdc4497d74e02e9ed805a2934
z967184694dd5ff954c2d188ec56be5a75659787b3f9f27e23fb673e09f01c753f09a0f940cabc1
z6b9d46da2c7e5895bed55a947c8263d92c44e3900cad2f0481dd7952b8356b9d1b8042a9e9d518
zea30ede4951ff1597f6f3c26e3c7d0a4453b242a5b9060260b12a980d1090825a6332eb9d87f3e
zce649101a870b6533c6383fc64ec489c323fbf7d49cd5f4d373ecfaa29c7c5ca3718fa8545ec56
zabbdf32fa89f1d65d5755e91ca3adb2f3f9b299541b744ff8c633849f0b9b7a741e1266d9fd396
zc6734b4ebe0b3c0fa78d8df2494fa3ac8d586625cefa54e6c5625f8cbd2f54ff724c979b1033e1
z33b5c1221787905cdfcb8b2657df85be69abb5927f71dc1b29d3c2f17f969f703dd85b5b4c0e0a
z7969e1f41630d65f81a38247ed9a431de9b6c7fce079fc1109c851ef4030977193eb22f7355c88
z033fb33346948612b143e8d5eae09428dab7d38361ec8d3af618d7a67cc77449ec41721e4bb636
zf26bbfa09312034c2917266657797a5872f154b49795c3bbffa8fdeaa7d266854fb5a166d82d37
z0e48f810bf38e1c920e7c816c462a452103a3dabf76805b873072fa5615a4d90e7581b0a7fc15b
z0d4cdcccf8f4681f319b47268a208163fead020f9bb423288579dc97b18d2c162ecd995ed80549
zb4bc47351da503ba09f88a76516c3df3b0b3fe073fc1b94959f3c47e65c875e0db96bae2714126
ze4e0b1517bcf00341d53fb8010b562df9cb5bb0ca04ba20bcdd0f855dd8cefaf0f8b472595e190
zd7a095d92e44165a2d3c180924aadcfab977554d82e30a2b9be616df9a33f9fd6c54007a92638b
z718dcab5a5a81f64b02cd2bf38eb4a0a5da69cf2ffaab2013797e8fcce99abe0d096c6ee124dac
z22c6fbf24d45de4126a11022e4d8f492c8364df5868df06e016285c963f32eb79ce0420397d2b5
zb65b6eb8bf4223378b1ffa4a56ac3d09e132e7b983752884a6a08d7dd85fe2e60f040b59d7c625
zc81f681ecd71ccdf974e69aa8d32b9ac9abba48db61502ac7c0d12f55985cf2b5a1cda8fd5651c
z29094d443782f29fc4ffb4980929d1178b58f12ef33289369118dbd0414e80f1193d988bc466d7
zb4f228f8766dcc1811146353f21704ebe1f778a691614462829d178889ed9be0bb6db358b6b162
zecdac5b0bd4acfcaeef09427b5b3228ef104b91a4c11a93ac2f68f8acffd7bf10ffccdb5c6e13c
z3e4754da80657640f8a27e8e521bdb68cd77b3891b66949eb8dc9ec3b5ad2fed4d4457980fe5d0
z76a8b35bf44c19ef69f908dfd4d9164123c9aaff9e3c815769134998623a602a8a574e2c769924
z875f469b5b98f9e9a6631daff51c8f9c079ca975329e2954bd6b27b7e1edb161ff29214ae87bf3
z6835fb161c83f71dabe9fcd0417e2ae6fdcd121ef8ced92f62cb59ea1d35a03227e0e1f9d6e1ef
zad436d1454b40a300e14f225d6e5e9048b920af57b5aa55154aef6ca0d7db29709ea0796cdc1db
z4f7bdb640055b8d821814d6563bcdc6e9be857b70d2b3b0709eb28d65f80bcedf6ade7916fa5dd
z42b65e38d44201d2a392812543800c9cb860f4d784e0d87ff5c034fa6cba5e2230860968252b66
zcdf942819f774dfcac05fbccc0437479c2810a82fdf8b9b0b9234973f330aa975d5067a4e84542
za65c5eb63444548a1741e5bd5912ad2ab54ef6a517a43b4211fb2abc8603f66afb972b2d885e82
z5992fc65b6487aa1b705b10879e6de5c9600580ab9cf3870b7bc4e666f31fff5a945f0abe28f59
zd4b9eb0bc2b377944dafca2bb0588386a51a7dbe2a5e4e74e130b7ee9bf4636a5fc1a8f005522e
z3b5f7002d28f6491c53c7abc0b50661932b7d04fb34672b3c3b7edfbd0ed694df8bfd18740dcd7
z1c84600508a2b021bec54c177fddc6f2164ed91500f30513c68f6a71e5cbfea5de21ce0df51402
z1a60286d93422eec63ec924f0cfdeaf1d8d97dfb4a851055e8af18b0fb50c68ff17e7eb38a523c
z7b226b3a3028685d031900b0303abb06ff89a2428a6e169cee3b7f29d120150041133be8551302
zba707bbe1c09da9f1b85da28a7371a41bd47f300057907358cea86bfdb65ec542b52c97628835c
za9269f6a0d846cbe309586090d37ef161c6dd15b8b1345cdfeeb5515a748a0fe3bbca7b832dd42
z00b7684cb9564dcd8e96cfa9d28af1b6dcb8e66f8885990243a7e19afd68147306c2e472f93ee5
z0bc3b0dfb336bf8f08fda5bbe0b6731dcfe1864569bf6fd5089a1ff91c881f2439dee90a098448
z37bb67f7d93e1a9143f2d3d6cb3e6e9d7e532710f3ebe113eef936b3f1724fe71c05101eb9218e
zf7e6b698b95b2a3f5bc4d3f06252cdd1dcd1dea62e48b7b167fc9a2fa2483f3160ca3a2d687c75
z9c8b5ff8aa2bfe12d05ac394200e87fd83ca59ccbd9173e84e2150833343aa2f46ffb42bfbe56d
zc9a3f5647b11eab797b46c9399d1fe1fecd242326fe57e6604004598ebe423060edba147bbeb3b
zf7c5858cbac89e3ebced63d3dfcb75dc67cdd5f85a716fe0efe941e714e9b16e4ed0fb18e98ec9
z952abe893adee99b219f7751e1040c98a0061fa9d1640542021c256c3cae12e0fe32e474f26597
zee6d3b7505acbc25d874368d06ff31dd90be90db9ead58b398c21223652e0480c7f30661336914
z62a857c9939cb01b21a67649777543ce12d7c951aa26306b7bfdf7ab20ee18d1c9b7c82dae3853
zd109f61cf89baa1c4e1b18b160a120b3940ba8e68ef30a7d7ad5966371f9b332da87a729dd2e8c
z697bfa03d0cdb0918e75c1c407419d95c2615ce00216357403e2d77551bb8e42565efb5a9045e7
za93b1bff8d966ca27bf0cf559f2c9168bcf6c51e0c4880ff721b7bfa7c5a7c32fa2a722d36f3e0
z4da64b9e38a661727680c2b20991c56d0fe800e33e9fe4679b47b1b8a9c100ebedda8ac7ddd2f1
z73dfa0fd3fb79f022ba3b2e91487b88efac3d2831bdea8c5141ccee690059063d7290c84fe7cef
z5e7a2ef3f0e68306693f222dc1dda21c8ed6c91aa822d10bad3167e6769bb063035c4a4a6455a2
z6f8a9a4b416ae192e5a39f6d3ae08cc672d7a9058b1e531896479d8b1bc59727bed31d40e61385
z1908b4eb91a3e4699496d812408ce5b8612feee882472104198ce28216e0fbad2d88e994382763
z3cc67a0d1591055de69f703b315dccc94f776edd70e771c6324d752f63fca08795217d75878cc3
z3828e30dc7fd611ce9baac0da620f1dded24bf7575b2848470dc110f0c259cd750d7c9939b7798
z1b7ea7d9d0c8c5774a121c0efe215212fd44fc671d46809f4ff08f343af5502eb2641a162f7ec6
z14e9d54341a61e4fde233af4e770df280a5e6fd6eb7378fc7273430c13c9244a703a4004c7c89e
z916d7a743f084ee63348db3cd70c754d4a2c7d95bc19f2d34320ac9e535486f62244d1a57f7afb
z62aacabdc1a2dbfea4d981cb6f5f7a22aed74a6c8cdc0f2e9f4b8bb8c74f1e5f242fdbc340353c
zcd328cae7b058c2150a1b379491c9c2afdfd9f2c1ace7acd15d330d579ed60763cd0785eeccd7d
z7c9073ab8d8e1a3c4b176624e8b3079ba48d48cf3c12da870cf46877dfb5c6c1322bc23f695745
zee4b4e32f64c3ad5ccc13c0fe1a13eef67baa51c73d65da7d1f83422023f9d436be394211679bd
z3585158a6672846f046571e310a8d38f33a3ff966cbb2929d07270c9161342854dccf0874cd2a3
zbf369d500cf160d1c24532526021f0cca595fe05506320220353fd343dca839ac06eb73945496e
z2a2070457c4f0f7933d53fc20754f061eb5c18c3b9d68eb1ec84121b0a83b54e133ab6f1e84d8a
zd96a90984f005b412cc93fd85df01367cd07d328f147e1a2264d5004339ceb2110a5834a54c870
z94e6fa8cb7501f8c45f4c550e2a0e6b5192bd89d9c4a20d28b728a35deff4802f2414bda02ac2a
zb8c2026c86eae6a9a0d4a2ad762b8e0ccf66dacbb9a7a2af1f79ec60abbdd4fcdd22a83f8e66bf
z0b144369fa34960debac02bfb9bebe40916597a08a3a98fac92edf6d7ded91167a5a523c1a200b
z6d8201d4152cc694a000ec42f206ffd26eacb2d5114e5df105367bee0698615f64b61e6304f621
zc28182f774226f690b5828484e1b829d37dd245e19b643a1ff54d03f24720a8d3cccf9fb7ed34e
z08ab23028ae237a801d038006ffc61bc3d2d30cc372819b106d03b271c04d6a50c34e0bf19b36d
z07f4fd3043207f2d8aae3bcd6b70babca9c453ec953cbf606cf71f3e6d1ef962188ca5b615a6e6
z3085977ebd080b9242c753e0ae5bc3a9887d23b0e5fdaa66d8dde7dde85eecd6613eb8f2c741c8
z975e0455ef682dd1785a489ed546a85c918e1d379afa21563ae03cf05db301794d644e6b3774ef
z6a10712a607dd7df9f9237462386b6d4931291e18497d39467ce61d53b3fa2a356d7dc32abba0a
z207f5187da0a559a51c9a3b877395a47ce4f00b55d40ef9ef11a76c5e7b3d8635ffb4a821b8bea
z325e6024ed529d7b930038855ebf3e1e2d68002d2f02f3327e9d185d5bfe8e56d359c3f573ea69
zb7bc7415f295e4a839f8cfaeadf583e98a8b6dc272a63e5f5e3917984503a4e08b63d6f5e61539
zb2289fadeced968aa3d3c5e3b456f6b0a38935e7ab25969a7be88078dddd5b31e028baa4fdaae9
z7e6117b6a67e5f8428723ce74c1928cec2ff154f1f406c3a2831698c2bee4156976a075b10a910
z44c53c17a8fb2e924040868d2501e5cfb03646b4a24c96de138c02f93333bae6eea14008845f27
ze99be4dcd64b337c9f068136095b9b02bb0098bb5fd728486dbd07db9f640583bdc394b88ecaa1
z5eadce28845c301f5488b8f41c3c2fd3db8a098bf20bbfd1b39abe13f83da18bd3eb2dc5cde3e3
z779879c99f817bbabde9ae8b008b8b454d656d9733cb2e11887075830f51df857e0ab6f56180ce
zc3d877c2193d68e7cb0c1570b355b907543142f0d1d4fe1d6109866a7ea7436a9dcd857867b5a8
zc7e33dde251e319e28624d147160a21ca64c09bfb4db02ae9cefa154008b468ed61e008e9228d0
z804139d64a35b65bc4d5aa9e9f0339fcfe47f92314d0cfc3911474cf54a1afe142cf32a11cb5f6
z54a3eeaeae45a5cef5087bf604aac6e9d04498b21794ae64a9b8ac8a83813d60abfd416b6bba5c
z11d08507d54602b4578208e58e2e5ee1ec626d71ead06bc2b10043b05ceed409dc717807af43d7
z7189f200cfe5918b80a6f5648fab00b250cbfcfdf7da0cc5c993d7f60b323e3da961999bdda904
z0246aaefbb8c692dc5705ad833b2813354aa5af78e75d24c024083df1ccb6971066f816aef9a32
z45f87a0eabe31e4c7892f12322ade5a373b6355ee73363e0b324f6063a8aa27552c5473dfec3a6
z9bec95751429844da6b8c9a290bb2747af8698e59176bbe5bce00c89fbfb4e1b93666eb4c7e534
z46a63dc7638af7f4e267e4b6f810bf19ab72ce10150ab374ca60ec38b0ebf3e0cbe02585a73c71
z8dcd978f7ce51d14db1e6863edcaa8723bf00c92b22b8faa1a8d8572f4736022e3f3517e9c3c79
z7dcc6e8391595eae5ca318b5ea9bb99924852cdad34c95148091b2bf087ea23859467d1f210cd5
z03744ec17655822c68ed51e48cf21b9eb7ecb82e372cf52e0c6594d3ff93372490b1573c72bbc1
zbd9267c881f7526c066b68b7ac4cee1db5aa2c05deac52c50520084853131132358f7035964b04
z6899a44975e093a6202991cf7c26d3cc588c0abeae61028fbafe9f9b70db142899d8394409cc01
z2ce3205e2f5fb082cabee79cd4210249a2ae6380742bedc400ae3ab18e939775bed6a15e04764a
z70d4a3266ed282a3a2fd1cb028db199fd6611b91e63681fa0598476c360015c2567db652d1916d
ze508a3456157658f3d39d0df600e188480ea48972d8fe24a9fd31f9c9ee3b37e9e1f69196d30e5
zcc97b3bd23e08391cec92668b5cf362636aa25ba92ff3d483d53ea353c955d7964134da411f324
zccced409a910c79dbfd135ccc6f8297c11a9853493e649e3e87aacdbd01bcff413da89a6687250
z858d47a5eb7db5c2d63798d7fedadab625763c689396a9dd4b86688a0a7029fa764bd0f4312800
z22dd8b76d13be19117865d493a4e9cdc614a21ef53837f4ca6bf757eebaf92dcc5f1ee6333a5d0
zb8977e2c460d78661268db97fcc93b6f983f6ad2a6706907a6d1ecbbc85d32317ff6b4ff5e006a
z546a4be7b22a83b7c258bd1c4b804d873887bf5f7aeec87476e90583af965bfa1c8fbd2724be48
za7372542525f415236a212fd97cf9c5e64c4f7aa79907e89f9c679da8b85e34e5bee3d67bc83db
z49d113f584d2e00bf7f3483ae2c648b21a05e7d088bb9f62ef542649c26fbe3903b0b9f6a9f879
zb817ac88a8777ef93c35f560f338221dfe6cdfeee42efef217a71c13b3eb793798cee132c07083
z3f5c2cdb71a1125ea40497b1306487bbe5eb5b20e037c391ffeddd0cfcea0482d1e950fddba68b
z98b742ff08c99675f0e37186f3522f7bee0b04e5aff4145a76823be29c4353c735654bf354baf7
z1aef09d0e868de4c8b20201db45f2b8376f9d722c99f806dca06405dd020a287a8f23beacb2149
z696cee808c410cdfbdbdf888634f1ae123356230c4dda26205a6f3a4c9ea85370be6eb327bdd91
zaf847845c83b51423dcbea5e3afcbf7a4e842d7e37124c350ddf846c40d8d1198f4818b5a22be8
zba014702fc1147f8436cb4e3dac1248acd69706064905b0f04b17276520311d5425ca58b49cce6
z70ac9a297b29752c1dec33ca6a85e8ab8b0257257974417a7ec6c42ef06a8bf68a5428e2bfdd1d
z857273a6714e39dc7b7dffbf6a61a8043459674dc9ec40b0f59df0379ebf3a06ef9c08ab4f7b66
zb8bc034efc3f7c26d50d848b19dba1cdf31bb0f5dc8b05c1f6af68fa5a02835d049323f372920b
zfb0c8d3c1a17cbdda8817fbb89b23c61c5b32d98c5709f1c8740502caaad7b84584375b55eed6d
z4aa92aa6d6d4f7d4dd386f3016501b41e98ffcb58989623932320787737f7f9482271092be695b
z092a0a95931b421a60874855eab44e5f94a3eae50f1aac71ffae4abb3a3e0b783506fd5c080785
z02593e9e7ef006da60fc4ed2d63a191443ac37c18453c201dc5ed36177dce4f38efc8f3576ab36
zab7f08234be8715638a81bf1bdc0b0429a353f337f1472d1860d6e3ade92613b88cfed237c65db
z242dc16ac8ba38e8a69df40c3576e9c1b76a6e364491749c64abeed0846db42529f29cdeb9e636
z39fafc5b7cab2e164499542c0ddd4d5d3fbc6c419b7356d9c468671f1e359c1589ccf1399886ee
z68135653b96fb2406e3c3ed278bd777c0774dca52ffa3a3a5408409abf940a68cb38e8d48494d1
z0c3565c66d6d586cc9604c17f737ffe3f34fa540c9dfde5dd1961f5c975cbd9c154121c66747f9
zfd448dda5d500953d041fd3f51bc503f11411c9cdb88fa6a8ce6cdfc6096f61a76575956ed8b3f
z96233e4febbb8c1e270bc4776a5db0f05e74db08acdfcac4868e74f522cab78456303c522540e3
zdc99b5d95327c5cef29c1c473f43440e69c69ae2304bc114e5cc977ecca67711d25ab3e0b449c7
z15693379a0d49ccd4b4c35624255a76b58c731b3b0687a92bf8ad4192517225c2c50077a90d6b9
zf10f3d0830d9770ca1d33883e9ae1a22e9fc19ce84f8d88c9d81428d42cec3686d827b6c02220a
z3004de236589113e1cc0b17bf317fa5b00ecb2d4f3cbab9759a24523a45e628e94cec09c66442f
z78330a726ee5c43a79b929256ea93ed5dd71d86a7aff7605b2f8b5774c29018a5b9165906f7c0e
za20c7522fe3e5081b74051d29b478b27ec4f8a9c3b88eaecd5365b7f998374593f82fdf243787e
ze315bf871adba2a5608d4058e70842eb9dc1bb0ba0896f4c2bbc9235edbc3edfdbb02445aded86
za689953ac88e9cfadf6f82f6e5cf6c90d5122d7b072a5ad009c598955f7b04fc060e3f45899732
ze50290ef2206796e3eb5cf37426fa5cf6d58dab509caf72534d69278daa4e25df9f158a74fc58f
z616f8177adbbbe52279dee61c10566fc528b0ae48730d6717f6c8370f8aec7e7ba06ee2063be4b
zc319d8511071988a4ecfbeebdcce1196490d1f24535803af507a310474219b7154851362840a97
zf12b4d99c0d3365894e1e94d98431bcde14e8861a8416c8d74b2b4d1fbf1cfb1f326d9d83e69a6
z2fa3aa9f7fd958fbe29070e32211db0713cf17e37a53f3981f6adb9716d4ea2283bc7dd2f12438
z55e24b7df2324542bd790228254906bc1a6222758d7951809c2ec397d1a8e95f6d74b729ab24c5
z44ef52d2ebfeaba64baecbab6ec34fa9778ad0cb28a21ff303ec914bc35c43d8c8ccf9024e9258
zfe1dbac227d92b97c2fcad2fdd4fa197d91bdcbaf4efbb0b1ddf5012afd88e55ae5f48945395fc
z44d9de86e3a5f48c6c62b1ed51a656baaefe036898514823897a30632d287c849dde8b633e4764
ze247ed5f42fe13b064bad0bf09ff901b848987d13db8ddf5ac46259c844137b7fd5a588db3a417
zdd5686bfb45982ad9271e969bee94c3026d064df2fa6e1cba8376d892a26b7abe063ee952e1d08
z43599dcf1793387a2559fbc0323a28b62488c53a0f50cbe56fe5724b2268a3d3b73e153bd4d57c
z6a24070e9b866bd69d3169e81f9800dd90a82471996a52ed18c81719ec69afe5c0a27430638edf
zf80c821bb32a9847a47a439f56269ab4d7e1778828abe06227a66fab0948c6f9637d7c92e89a18
zb48e56b2068d1f60a49ea3887bc51c5056fad98484e08c27a83f00964dd8638ff07f16734a6cde
z1ad8bde0f341da1aa62e95aabc41eaa2d9ba63ef4d8893878aba814ed989aa51b1ca62ca8783b8
z4f65acd77901639e9236c20b71e49a77e3c1854e23fc90663c5ee212121ba7bca81a78988460b8
z7d8112647161b9a0591481f9d1068e934e299ec484ac25fcd428c3125cca1cc2e4344717be2c06
z2e11a8d48d8e70f4bd07b5004521f1ba9937ca1ee6da276b9b47381387048103bf3f2877c38ea1
zd3e074400683675514c7c7c9d5e5059281144ac3df60f984133c683bfffdccb5384db064c12c37
zb7ab193f6c6a5f8f03d4f06ee76560aeb7b4021607e8677c2578b0c7c77e806c45bf6ecb70cbc4
z7a18b9a05f733db03ed4683f93f2d01a6b2df300493660bc9c5b92a6457435c95e7f1c85d0764a
z1e487e1c81c6de1d4b60f653c78b96b05918120cb3e43dd772370519935677fca51d5f0cd7980c
za2357b1cc3ee6a6e1cb185866954bc05660b445e5a3d79d9576dfa9401d88be5ac933f6e34a5d7
z484bd343c81e2d608ad2bc87175169aa05096fc52a67658820d92bf8ac4841b8941a93cec7a419
z8710315aa5a2099e8e188f7d5aa02dfe1d81ef5609bc3490326d861dd44f03ebd8a2da38d59213
z74dd521b21c902d5fbbc44e6f1862a36c31863cd1f34897fd292587d52dcdd16d755c915b3ff7f
z33b9e02ca78e6c632d781174eda507e1a922261269bdc59ab1ded5a8edca006e4825db1c6db7ea
z6557b2b61108657463b873f034214f8ecf925952a80c591b896eba9797a2fd04407fbdb488d9b8
z6672f7217d0de36b5d5f4b7fa035b643cbec1780017b022f46d82289ae09189e1c11ea4f520324
z06342c072215380f31df07f8b96f96ce83c4b16fd52f411d774a903aaf7feccf0e9cf892b334dc
z514de041b4b25df78a5f0b968026ef9ea385ca0ddcffbe881bb547721afc48e7f9335e9cd5f070
z370abc191f1c07113445ca328ad4b50b927224ba9426a386a66c25a232179c366868ecd03ee429
z0a1dd0b58a5ecd75a11470388bd9b876ccd6f079fdc0e185a7b85f8ff23626fd8bf65c1a71b2dc
zae94b6e944fe6530c3545084d1fa477ba89a0344b0ce89f8086ab09f63956ca4a12824afdc84e6
zbe5cf6f293bf7229000def3bf15f95830c19d49e1766bb34d2e9927ee3cd2c9f8154b0fe860724
z68cb17d0c08971ddd81c940a8b832c9d50aed6249378976b0ac0abd63676eb33a3024c0b3a28e6
zfc84a765260d5228a96ec3b0a717ec57aa2b0a13d5c452769c867e357d7084df7cbe8df2e18770
z803fc91e9570e91653e7d4a88de6dfc29fd1e41630d3ab4e1f768c344a906d540fac9d6957fa60
zabb1a5292ee57b36be8f2e44e5eb7c0810efbd7a759bb3e9029691a19038620a28d7cfd62f3333
z7f4799ac7873b5d5371112fc02276ffc5b7939d1fc118291dfd13262e597db02bc4d72e87e31fc
z5cee53d9d753a0a55ab97aa9ac6c35f200988adc94e9b8bd1f0ce17252ffe529447c4b478bd37a
z6055f26386eacab266c92a69748209032f2488fe2f3d0e3e27d77bd0cf544daff5c921ef621fd1
zbee46bd81c28a3c5b85c952a8a0fadc7eef86728cb404769aa031b7eb261288c3436995afee3c4
zc135dfbed2ca47075ce0920c1aef299f0454bd7b92072b19eb7cc23cfe43b793659fd650d243d2
z84829085ba2eca4d415b32334e805a858bbf8b2bef4dae1951eab201ea4ebe986bf54370c0a986
z368140073393df176f13711d413fd5e04b62618b33e51d45295cdd5750e1b95a9dbb9e7bf3d311
z49bab3bc11cba1fa33c8529c1e40af7ee8476eacbf237984dbd4417807370f38494fcde55cec81
z59e6b4fcfae7c389cf73de6d5c98aefe0ce0092551c78d66c4ea81d1b8e82557bd762468175044
z59c7f3dd8e4c87b5ae7c27ee1079b3c119ed093763e954776900319ba13a9e438323d40f4180d8
z8c85a4f697791d61720a41f33bc9fa0e364861236ee4fc8d054b0deafaabd66aa49873da90ad09
z462e3da9986408034d92fa1ee3113611f4cd83dfc7f4ab9103affdaf83a1ec5a130f92fa1d9f86
zcfd81384263792652e48917df7aec0c9b7f5a3b476bc87a91aaf4eeab53a072452cfe0852dcf94
zdbda0387cc16eb25d54974af60414c3329b71a17931d587481a1725263dbd58b3d09f1ce2be379
zd52ddc355e837152de99cd6f38df8215ef065b9444fc3b5e6ec37cdda48ede51b8c8d0f956f623
zcab6dc251d42bc6b3edea97682d41e7e33fcf7878178c2238670ef8ba06985de6c4bd50be727cb
zc639088bf74f1c72611e7e0df5405e3beb2f721a9b7618673bb91abb9a589b9b7937b75c608990
zfcaf121804fbbbf70d79cb022b578cd0c78a64076af6306227d52ed3c9b711618b8f931392fedb
z831bc0d0813e08f134f8183c49e41806c27703ff1980870640bfce1339211f729daa4488f8f3d4
zed0495741277f65f8c6405be871f95adeeb04b866844c0dd08b3912dbc90ba0f4d2f6733fa25c6
z01ad714b150ae4653f533be64a533202d7dd662c422085a70d13ecb3f69afe40ca326461517d7e
zf750e5e8222b863a41fc65fc209d9e8d9224f571a1867f0e32f6599b08d8628873b6e4b3505553
zc94c354301525b1cfe78e5efe6eb33f9e35ce8f9a9dd1e7bc232a5edec5b81c8d6a010be2c67dc
z8ad980c8690e0e7a7f04162aa81a17760c76fd4f557613ec3752a6accfce18a817e7776cd2c5d8
zcd65faa6ad69dedd705a409a59fa7a0e53e85dd52ce48205cad85bb9b60928c5b361156469cf85
zb77c2b92bd2c2bcb259323430714bb2da469c893b5982c518d9ff926225a993ab2233fbd24e0e0
z02045b37345cf83ab82beb6c57db88f522cd071ed1b9eb62b0d377a30530d8316e2797c0d0656c
z6afbb79f4e94cdf13a3abba6229488a134978472d817bccf841b74771a3c93146daffb40395d4d
z2a951729bbfa8b63e12a73c55364cc7b96caefd63ff4e268f9fe0a15eecdcd3a2cf5a7978d9739
za8b3ea1fa0f12c63fc66e37ff0afcc6d16cfb4fca53384b35b42e502d0701ad905aa9c8d199ee9
za03fa505e8229a8a60edc56cccb4d9d138658f6e60e134e346415c650086f56315b18a15d946bd
z7f860f1d69a80ec067e77627f9bfb845cb8c41ea1af1b0bb0ea75a535cdd2d739ad022fd021141
z91014797facb1bbf2761ddefa8f9e04fd35ff6026ebfe3da7b059342db287b91a49c3bccb2176d
z4a86ca82cbb4a5a2d30229abda3d76c6ed9d8aa7c199b9c08f8e920b98996dc95b9815f2b66ba5
za610eb72ef8084c3855a6b982573522e8c2fdc1ecec72e5d8aea765929a85895746fc36c61dae6
z1b43f85c2a1bd3c130cc5d0e77396d23e8e12dd8080c00bd55dd4ad6ac4fdc5dd0a23629395248
z0abe0f88ca4bb2e488a2c7e32dfa59650a56a3df4abac3c8fa4e0559cb1ffb66a4a4bfe7f1d66b
za0488a76f72ea051e9954a976ab3a9f27874f4ff8cd6ecfcfef4230b99d5f55a1bb8bd69a30832
z9b5036f1c665d8af3579e2d8c0b95d96ace63454fcca9c273305c9773822953e9ebc23eaf628c7
z800e9bc0dac047972824e92af95deb24b65639d98fb8012101e9e3db347cb1de8e39c86bb777d7
z4f6713ccb0bb5bcee8453429703e7c201fd268aaf034c7626789cbe495e13fc91f40c6f8e57598
za963f35da2f6b2ac78e78fca9d81b14eb313e4d8c65f6ebc40d97026501630cffa02e22f42e7cd
z3b5e592ede2ddc0d8481afd3f7a24fdf69b7c1fe8e8b8a6b16837f534d85fa87b915a7e250cc99
z0de793827658113bd909d35494523c6634050ceaa5599601199fe6b82f1d58c5c2e9ccafa6b4c0
zc2e7e1febd97002e08acee3cc995c5bd6b4a2f6a468945250c362db818a8c71eb4a076c87e4344
z47930999b9f38719b0a0459f5a404f65e1e648f022425a44078b3b4f645a0f1e9bb2ad0870c6cc
zfbc4f7ed55ce18241ff02cb56fce41a9a67e2ae9582965eccef0d2ea6178f0bb2adf901910d6fe
z5d335dddf02d9942b01c87cfec9510dc0b93b4f18a9703af91115b18919effe9ab14602e2bb7d4
zf95e705fb60eaf2d53ca8593a2e32c5014b64f1f17d61f7ebb716e1a92e93b02600dc34b87827e
z99dc52acb67185af7196f3935f893eb5bf9092b86804863cb3396d9f148bbf958e2e0f7a5846d9
z8c6fa46f6026a5c2d9600460a41476ddc017a1ef38c766fe7a19ae1547ed1153f7ce029649d596
z963cd788375f653d4c277d210e84fd46fed24e669c187fff3cdb8759f1789c53876aa3749c9e8f
z3ee4277a743630a7be2620333c3f8d5b8b5b070d557bca2af8856418ef83d3fafce8f9821b10cd
z15b634da3fe21cac4b2ee8c47169bae09707901c131c2b637085e6fffe008b8567ec42a8974366
zc529abbd2c583432d8bddfa72b2a20acf6f88db7208171d30b671ab2df231ef96c55968dcd7bab
z688b4e4151d4bfa4efabbffb45e19dc29c53cbe4752f1b7892d2b9e728aa9dfa5926f9a55a1dca
z2fb12245eda2443594124566213127493bc5c9962c041d0d795b978814a0418f85d4791b95bc0a
z9772a8a1b55ceed161db3d685b26392af1f65e5677f878d5e7ef7a1b10745b7edc8e2668c3d880
z07b7a9e507dbc356c2a7d509fcb34c6f164d7d746411dbcdb2d678e313d18bb1197ec1dab95f44
zff95fd5daccec2a13bde851165121fde6d358651fb2610a8ad8cff4994655b17d8e72e656f8450
z8dd2f5b3d80f9a311387ca6ec26d38868bd758423311d830f1efcdd042a0941574027588ef4f51
z2c701d7cce82ba1afddcb34e49e2634636b79121230cf302829b940bea927b4150b273d1a7a6f4
z7056374643df7e8e4aff2e31c44900bb17adde52d4feffa8bb0962f43e812be32d7f11d39df279
za06e09f074aac0a260dee49de0189a1bf6ee4584e94eaf9ad1e27141caf0e7591277ab276e934f
z1a390399d60022509f18d74a78a732b2be0d7cf463d08473d5da85df076f06bd40778c1703f377
za4693773f9325589728cb25d6633cf7e72b4b6335bf7e4efefdeb49d58a6a87a158d3e19b59b73
z69662f9c0084d09192b87b91b4a0390e34a7db461015b12b5e42a44914b62d8f9c64aa2337fbec
z387992ca9214ab6ec94f090704fe212c3ee63dea578c7760b91176d647423ece39595323a469f5
z997eb91881ee8f6609c152c59fdb2a3a5b22ccb966132b0b7cd3105023d1d1877126e0312a29f8
z5c9e1ce403a84c4d43d50b4ea7291ecccb788f1bc6269bc180f77d6260c6a1c3fa543ec67754c2
z3da2695329fa7986f31b82c87c1592447cfaabb9bdb20f7878a45341c513537399bdd238e43d27
zb3287e2443969c701e59b8b0223026ed9f2d12288710d4012c07a47770e5c4e6f5434f791ce339
z4ce788ce6a40a81913895e2556bacf9f0560b45606fb20e0f302f9746663fd4dd9dac749df4e58
z77a7c55a2190b67205a1cb40a1080de9ef5431f33f761d8b937b2ffa8c2e05474368b9c912fce0
z75de5b2f2fa17a6c93a177c79d92f977093375600f60d812682a8b1773709566e14b92887f672f
z462ab2cdaf71745b1f85d05484f729b4419450df2e726e9b06a50153dcc9d253691c772cd031e1
zc24557b73041b12aea76399068d141bea6dbb01a7a81f58cd4d1d7213b3a2c860ba96398edf098
zf4357b76bc2443654f0b22a18522b04d21a314ba01e5bdef29a27d2c51913243c7f797c1802f84
z24c037be5268b0a93559d1c2330571e31753be1333aad4d1173b8b83a9b4c3090b990c352b26d9
z960110a30a2328dfed34a7ae56229d689ebad3a0a55778b23b7766ab264bf8cdf03a97d3414cc5
z9bf0b7be348f70ea12f94982a7b2b597404e3877356af2773808b71c149c880740be058adac1e2
z292094406631fc41ce39d9ea08f5fd8c91d8242b28c25ae0e0206994e771f50185af6e6bba4e1f
ze6b9f01495482f7c7433f8340e79d9b8d9ad4c5febb80beebba097f21ddbec5f23b233cc990cd0
zb055f3fd58aaeb7782fb58511f29dc5a4482c8afb81212f4f20fea195e8653d35805bc09985f82
za0c9bcbb6e41ff596a068bfb7834be7f44d3bd95d59075b5d9cd98b89673ab2916725e47e1a103
z7367dacf7d58d90205d651f0608fb84299b0c93d1ee5d71865a9d62c406a18a99124ef4acbf642
z4f0fae32df0ebcb99dadd452d5f7b5002b195d2e7e415b188600ef544c2e6649813a1e112b7875
zbb7b1311adb89b066edf365161cc60b2aed845917e5550bedb330b416c6b0112bb6443841d8bd1
z250f7c2cd32f8015db19c87aa8b5506e300ffbb395289c76ee22d58f5f334f69b63f68ac4f46db
z29ae5d61765ebeeb388f4adaf33c4435e0294534d4a74205fa46645c7bc2e51b8831a99a9c7f3b
z7c088590471eec48c4a6695af7f7400b79c98478fddf862cc9da4f838026fe7ebf76adb340e6bc
z9fc95133ca85b19c439ed97d3e2eaeef52fdeb9a86ef624a30a8b294896129f6a927383107e073
z90c00a38d13adbd0cad3c780f95242cd1f29ed2d41b2983974ec4c0611fbd436addcb80e5ac9ea
z7cf8ff2bc1ecd0a22b4c3e79687742846d54ee0fdf4cbe7409add555d2907a3999dc62122d4515
zd2f0cbcdfc67a36a8eb73c93b97be5a2ea785958f38aa570bbd2241c8454b2b316ebdc69600196
z61bb12df8b7cc4ebd018050c8ed1693d72962fffe831e8a13d720af04ac7f33e8832f8e51c400a
zdfe7d4c2c5aa986c3454689ac5b4da2d6c2089e69ca431665aa1669d8fff586f7a6b0d3d27c0f1
z678b698eca18e0686d6cbd1104665c6bb043561103dc3d19149db01007af6977773713ea6a3997
z7efca20ecd6faef8f1c1eda642dfead86fc4d493e694dd13416f91704e237d9603ae3fb97068d7
z6a33d5174455f04767dfc46dfcfc03bab43872cf2ed6801cd31f6ffb9309ad51ada1b6a014c3f3
z5ab4989c122cfadf7dffade67723bfc4d09271cf065dfae70709eb54cce7c5295ff94a3536daa9
zfa328b86396d26be84c57f1ee26db40940f95b932492bf0edd721a8fa703fc22d4587ef788e0de
z33ad268a715155905b7d0f89570e84fe6b2ba350a6a2d2e04f4e9ecb69967ebe260f4906cc58e9
zfb8ea9bd9917f3a3aab03df141fb2ed4bce5ef1e723052186e583f3d1ba387e3e4a6fbef5b9cbb
z9671cb60b7c40b5e9445bf0cd4739228e3c5c9af439b74e15aff35ce2b411735244c1db3f44c5a
z5207d2bb3ab405209d44a4a70087e56bef7392946c539b7795a988bd2e10e4a1f74faed27ab477
z21152d5c8e2ba40f1e87a00d2d59f6e256e822d326941e581a1714fb5657c52e4358190c24886f
z2b360af5a11eb6d349f959de3337eff6e93e0a8255ab303c7bdb46678dbdd2c3d99d04be7672fa
zca48eae2bacaea3ff49fed053e93c1fed3d3bcbc8b262fd52ab5af71d76e9fd695aad042db3097
z61066a3c9dea30a5f1f10442382a66c2f9845306fba056a2238e8c6fcafb008608baee44b5217b
zc392e05ff0761f730b8417e2a01a4cc872b930cce590b610c975d6ab9787e58d39837d242c3a24
z663ec74eb73037a2d3b513687dbc7ea7dd51acb15650a0d5a43c18d21e41f0eda06b762726f7d4
z0f1b4bead5811d841611c58c1d55826b24f9787c0c373c180dd23bf6409923bb74e099b2103f58
za94b85b50a2cb8951d5be4a2f1c7d8a53418ccfaf55811a838db83e7acf9e60951b35f9f63a506
z2ad8ae6d3c658861fc91d5776e3eab00e7b877bfc023f8dd9460a39b5ebcdc90dd71f947815b70
z920116bafe9f66d3e5d91d7267fdc67046f7acfc7f583d03603bdd4d0ab36cb25796697fa52773
z2d9f16fe900c7e57e31c1a9290a49d2936382ecba8d3feef2d08e69e20aaec772a9fd03bb0e661
ze97263e7a5eda2e312536521ef0d5de2b33c66e3ac01fa15780a865b36451c4370253123b0d937
zc170b760a2f5845a68d622a4eafd09138dc34ee91e4f9abf8bacbb3df8d03cd342230d2b42f63f
z61b8283a6c9d7c365b6bfae9e6ab2ce49b63dac3e8ca133a1640382cee39fd41f2a52931514a2c
z19a12d0a59c59c7a4d6687c3a097bd54e96e3d6fb7c3313a3312b40449b5f52ff363e5a9650515
zed2f98da99ad6e776a64dd36644f7ae171b893e464cccdee1c409cb5b9ac57b22e1a34ec834547
z003942168ab0350ac94fadd8d1a4fad249460d65474827450c920d68945b17688d114b5579f95d
z483ae570719848341527cfe503facf2f0bca044f038105f9965ba0823b4a2230ea3415f710ff00
zca74ef09e7799ffbd093f3444148ce81e735956de55e4e23e1915737134fd031475a7b9c45f762
z043df493b9c764e8fc898da8966ed984cb4b031fe1f2153c8feed5666e0af0405790c34dea3ade
z3f0fb0ebf3eb32fbb76f2826908ae0b7ca6a4a7d3799d83fe1e400f389ec2136c7cc89209cea77
zd025c128f4123399e46c624a154a49f13ba82aefde163b3d76fcb797e043584e58b3c2b20affc8
z303fa54f1a8be961593f6c37f8c54f48b55fedeab1c435c2c1c9f16627735002024e301778c2d1
zc64d2a5477544e3f8728c2fe260fce89f301b466ae865d1fb170eafbeaabd81c6c64be9c741a3c
z04720797729c6cf9e50a41639d72fb1e68c66c1dc6dbbc1f76ab13664dd9bef03a17bdb39eef40
za01b0c6384b83626ddca376284b266efce688209f5e0a721baded08dceb5a22c0b75e1d57c2679
z1f0f4559011cd4c79ba0e61eb83a28e63e2ea73927cee08cef9d4dc002d77dff15595c469853ea
zb59371e783ccd1822db726fb5623968eb43518e94bec504179e5bb08bcd9a1aa7c1eac7fb817d9
zb4441f0992f78c4069e17ae43bf8e44bdbc694e0ed30b2f1c09f5369752f769b19f32f3b13debe
z15183d9e8fa3a1bef0e51999274ce92975ac2611c2b0561bc69a3081d9fbab6b67638b121afd11
z0504df32de78492218c8a82571bad524ff470ca50b694087e2a066b5fd06ac23596e7f729b9f6e
ze695aeb5ce926b28239fd257b7627225e27d6bc6ac2c4a8828a52390a6ec6315c5f57757985105
zf520a086219c44382cc1016350ddb48e176e2719205d716bd3770fe5de9d9840052d70f1907e1f
z3b7d9aacd31ce77242bda227728ded312af163aab51456d99f7daee2cdb829a06a9b81a82fb1ca
z98cba5ee9dec5f53b6faf4e1fc96a159e060732266b9d71492ee6756d36b62300e5b67170d4fa4
z8f156b4cb22757725f5d725b8a0f22e644d5cf22aaa26997a3cbea8c11e79431cf8afec59f2374
z8f9cfc271fcbc219ce4b3acb2d2d38e7742732f2eaa469a96e43eee9b75e361f9da88fdb69f6df
ze2d0824dde3f7ea8d6a3d6cb4abb58e152f816aa8cacf80626ea3a49cd333cb784c91c4cbb85d2
z698cd9b9b38693b809425711727a72807dee6efff0f90643858d2c7605ba39e277331512fd3251
zebd8db22a9d6118b42891c70a59ae7742c54f2134d0dbac025a27a9fe7bbd2c1d0ea39c941a3ad
z09e675557bf5c1ae9c3300316c02d119234aeba21a102f06af1d25e94cef504ae2bfdeeb5289dc
z6299d3a9b922526f90dab0426c83c59951fc6b34d959ce4535f4dfbb238dd9aed4369d4e85b277
z322fff60148782b8bf00d38a97a26d4a2807bbe20df429570afbd7ed9a305a538bf02b412c23da
z7add06faae99b54ac00a7d6d59bf10409032c92d68a7d100505d7d70e5c750c1d6243037a74142
z5e853ca10db7da6501bed35a9e7fc78adffdefea01b33367af787ada2823bc686437a3498f3f17
za88329a40337ac3495d54b806e9328ee85d390a562e03bbeb2435a0a794427eab1fca94f909150
zf37567c4cc7a480a01d0497ffec553c20043a133835bbf85d8d4b8fedac2e64548e89c5364d722
z85db2eb17f37eca4087db669027d05a73def7c48fe16744e07271192d9385e04f3aa67084e8337
z3daa3261fafe98b2667c6290201140b9f56b41ce8dd0106efb9d66bcda05146b194a36bf250666
z00d3247bf39e38d650a40b2df2180d096aab6b6ab3b3a1c0153ae95f655a6918e42eb6e3d26f68
zf3f155c4e3533e53ccfcb2e43edd2f3e7cee7d9fe06112cfcfc5038c23c5591fcb9174712fb0ec
z70261cde0aa70bbe5774a46e7f017f92b0351dd527982cc439f35796a5207ca322e24595eb35be
zcb741c6d170cea2a1b1ed336d82fceb90b1727ac52bddea6d9dcdc443d4441e95fb7456c89b3a5
zdbf38469c66881975d0fe920847fd43231845fba9c2302e445b4459f58619c237f5d72ccca863d
zbaa93345e2af2886f3be60d1b2b79979e636160e5c1d4df3ef2a98800bae7e8bff7cd5f7d10fcf
z4130919a031181128177f8070da1b7c424f501988042e2f5f233a19794116722f25fb3c67bccb3
z26a466d7c0cf41d5ef0f0fdf9d4a2f3293cea7137e9d1b5e1470f99b50c37795f73e864def30a2
z7c85c2ed5fd52998429b3fd8915c2aa8554bd6caf755ccdb79d00107c3c662945d7b69e100a0b2
zf42c1b7575fc472a7084439dae63f36ae2c0b028e8cee196e2df00cbff0a33fd8db583e5d3619b
z8cd5e4d0b03a385d99110ec724e7a2167e0f47d2fc7ecfbf599b7840941da9f7b2ab1feb418485
z89cc8d9e38b7b8c4c0c3a8610595fea0f7089d66a8bd5e2c0403a3ae3b73ff1d28b9c5bc4a09d7
zb79f67f328f3ec38d338f9fdc8f38b5c821fb0999efaffdd7229ff2e9bb940986b9a499d153a48
zf148bd6c355774443282ad9c17f361f6b53a2a18693c9c32c2c98016900287319e524617281127
z32f6575bcba3021118fbbc7fdcfddb291c091051eef68a90f96c919a9e9c4a380e5db3890dd8bf
ze45982bc3836ebb79ac1afe05a362586842cc6f7659a05f56f5b642dd3a843ae2dd38cbeb218dd
z89e5b4e59dd1b6456eee6dd372cbcfb3d054f7382a4d58a69eb00a9da0a9b93bd11636cd1c4902
z66a2dcddd9ecf4e5b838e2e24d04dbec4ffffa061ae54a3a89c7f66b11f9706aaafbd6ef626afa
zc75d60733997bad19eee25d9d638232808314cbb7bf11aa6a415e829afbaab34ab9244e9c633ad
z6994a68be80dfbc9f0378887a14f6a71f02c67c238da174226cfde11e13efe36d27a9e2c63ac72
z6a43b940177a29e649868cebd3f93be0a92d003f1d91bbe6e522804010f2a2c9138282c6e5c38e
za0db81f127c6320f6aed4467b5ce3b8403cd10678cc66c2abcab4c6289d7001237271654372344
zc6ef3908d646d57f9151b51ab6e472ece2babc1f652b6d3224544bf7f9a387b413ef3b9a641cea
z5880ceb5e659bf33faa3466d09cd1da28ab53f00ce7756757359c025c37162a0c121f9c2551b48
ze0af4f9b5e3286daf252b9a112b814a27bff8ccbceb5019b150c1a7c143bceb14422f17cb9350b
zec406311658cc61480829d80c890f15e64d8a0a25bf44bb62766eb17de3a0bb5add6ca9c06085a
z9b5727b489cb00b538a68088879df4c5b2654acf9723d9a3fd2c6b5cb81c6c694ba988d9cf2557
z271d452e8fd326a85000c91c0cdba56c9f2f0a69765fb26338b5f296370b5de9e5e885ebc0701d
z54123c5fa4d73de7c1e626d339f17988a109359aa9665b61f2573160fdecfb36c45dd4832b4ba6
z0b15de2fbae493569524ccfac5d44a50a873986396933413f39f5bd6f2a0fd2f8b8c5101035855
zee13811fd7de3ed0af4fcafdd6367f3d73402a9a19d1d8bf3bfddba7c2c2ac1d342276532b37c2
zcac309784b51be8facb57d5f206bf4e45ffd8f1dd19a08b045a504e466101c8b662dd77b9eee8d
zcc4eb659c2582dd6bee90345362b448f5e7b0702a338d04636f69d5e7436a741a0ff2058d2b88a
z5041fb1996b6a27407f1a6f7546a8812b3c4877a21bc3ad16e4d402746b1def586204a2c5ce5d9
z6bc228b94460cd47b82156f4d4b3f976a04cea7fda81061e8eac04f326f03ee5e1c13cb9e8d30e
z3541565f5b904eae2eadf4b2bf4daebd891ecc359d1453fe48cd24d7549dbe2aa2a3693f3661cd
zf551c0864e5ac507f8771678cd73ac0093fc6bbee02fb69aca326e33ab76eb191adab6cd1eb2fa
z2abccf09c10fda4c38f5bd8153d14b09b0cccf0dd68468e2d7280d4f26df8cbeeaa7956dcea40a
zf9ec758d195ea4b609dd4418f678586dff3f6a5f328f4c3df37f429aeb9aee8bb8647b51822b0b
z4af3adb56759a4af5a768e9471ebc40e72672732ab277f6286743422262da4936b516bca364839
z35dd7faad3b0d30f56db8504d6a297e371d9428bb45bb9eb31be9e05883ed770ce7301d81b6703
z236b87989efe59ebed355726bd506b6a5c5d574f9ae405ddce8e68ff638de90a95873d233bc514
z644dfdd69a2bd9f488dc1a1159414106ac763d6772c0be79e17e9302cf87363096d9f858dd8ec6
z41a11d0475b11ccfd3311dc1289b8883c83f8016f8f025f91bfd18f3d826761b1e684805b7dbf1
z6932fd838f06b8bc2cbd1ba1ecffbb9f9585ce627d52bcfff11d5d6088619e28fc108d56ab557a
zcabaa2fd6bbecf6f786c62149b32555a33edf27713a6a3215b9eaaa346f0747a15aed1cf934a06
ze6b29abe998cae4175bd5ee034b8eaae6295d3dbb8f47c0cc8c044d921f06f6de21987f7ce2f03
z07476f658d471c1f39688cbbbc647f5d4cc0c353d6907f7caf7e21f9e3bf8e88c429cdd7e42ed7
zb8da107f85f0cdca81f7e4492de69b59493e6d0748ec2c7d5ec6e70c2b2285152ad4063f93885a
zdbba37c9c79eb310018f0d6df12582b1790da737d5dedbd0cce738e40018e38fc52ec779669006
z278cc936e18431ee594da21ec8c7ee12e6bacca0fb82108cca7b4f04aa10a7326e41ac17e8fc46
zde93732edd3501c321446af03c04841e0f472c04dc0a59160b4cd5e1f7d1611ffecf7178194715
z798147d56f89a8c53e022a955fbdeb00266d57cb814a150031145e851038d62fcc78da09590f8a
zdae38f39ca6d7dacb1ef1b5019e988196e8f6279d158318925a639b5a8fbd7003b26f028209191
z22adfadb4f26157ef7d433b3692b8381a9a84c2e2685518b6213f3518f81c3b79b017b78cb7aff
z83e749157b418fb522f6dd22f14431297b7c33cb529660e18ed8bc72b36849eaa01f2a26b71bc7
zd4073b7c2821557803253186cf2bf86bd505d1f6a640f10730f33dfee88b70e0d409fd6d372f74
z542935ade1c7b0551b06b455149d136e3b4c84e94390ba81593904ba01d92a04cb5f63b270488e
z06f669b4980cc482eacd222b980df6839802b6d3ff6017da2c1f611f1a296b5ca6a67fb722b1d6
z5361bc61696d1cd5fc60e0357500f93e296dc963202eada912723052e1ed99e6112a79e8cb1099
z833bbd78900cfc33dfd157aeacb9136d7fadd9bd9e288fff823816ca101165e6ecfa4a4b8d26ae
z49e2ceba564792d29cd9ef30aa6021f334801c95d12b67668c74ccc42d06be17ae049e4b68bb74
zeb8d1b550ccbf40f107caf741c34e16f1ba3e1d8667d18a388d4caf2d86f265f6a77f2923f7f1a
z5db3f353b4e7bee68870eba2f5ff6bc85a3a98d755b8ac1a45f3a06dc13117d5b674d0d8507fe7
z5ee757508218135142264d8dda59bf522509c409c2f528a940f33e7ff66898ad593ab908578aed
z97ab576cb85a783058809d172d08cb98e7ef600edc27f864e1ccb5f0fc82a2e9412983cac6d6de
za3b74331e058d3fdb81bb4c5bb7702d0b316cf63d465bd392602a5e4d20c1c60714b837e74009f
z89c07bd8643120df95134c9384494fc14064be5b6f82e347af8125a78572ba60ff5367c60fc52c
z73b7d890c7246136eb7f57d6117957b5af633a4d4fbf217330e73f0115c84562378aeb02b6ade4
zfe042e2eeb5f103ddc76d9ab2e3e1d2e1b13f7be5050c4b7ce588066a4152ab12ba949da2a8f3b
z8562687c20292ebc31c9341eb1f8ba576758582f6d4283ebd52decbe29d49b0341d09096ca5b3e
z7b029759630ff01233042ff4f84f57c602b89a45bda929fd1c3123c71a5f5e75ebd1f98e6b076a
z5ffa2b0fa62194040ee7b21f44298d335d9db0511db2b3664bbe2a64bd935d93803d8bf2f5b7dd
zfcea7fff47050d3bbb1f68b82facfbd65fcf6712239e12ab2bcc8a5816b52c91d4df60e8899eee
zb805e5eeb341a4734d8437b6871840f6ca0f6a7784677359e1653ad209b9385e219c67ca9dd04b
z06e2cf3f6c418fdfc14c3b7fae5bc4a7828744cd91a12e810308f71abce86f83fed1b73fbea62c
z89e110544b4d45641e30334ef539756756d6f4444c337338d37962480c27ab4b95e8f20684f4b3
zb5290942801b06a0b65ce5608019b99ee5e54f7d8cdf47352ae4b0013db1213d6cf053e598f8a9
zffdf1e02d00d52550b021f3e290e04c9ff26cb3cba7217169a0bd36d073f1c0cd2e4aafc44c20d
z3c937417cdc96db2a1b3aedf38c0d79f53e7f2e82977d284b64338d936a2737247dc7ce7b68460
zfb354408aaa15011a038eadcb42884972b4b5c53cb3c4e5d3387455cab1744a4df561042f89b88
z25d1acdf206d82199edb9703cafed1aa52e380d7e40035f5c4eb936360ecb678a1f9722cef6c6c
z007881e285fec4048f2a0a972ae451aedbc3d67f0b4c2635b3703c57b7df9fa0109ca21f2212d0
z053ea94b30455524850d45e81f9afccdb63a17e62ddc5767adf15933dc093b0e89f347055c47b7
z93772929f896300ca4604c0ecf143942687f578bf3e98e9842463b77713c4f1caf23610a17ee72
ze28e2a5d98ce64a8630c3ad7ca71edec64dd149f0a5f9a4c8ab8347b1a919b8421cd97b1d545ee
z76bb13c3b4c4e57309e11532ae35aef536104ed891d57b5d1bd5b43cfb057d64144fd0f5e1c6b8
z3691c642f9b4fb057194946fe51c512e46b850c71ccbe19ccfd74a7c6245bac52602780d485bf1
z920c1cd2ad0dc22aa298a7b39a272cc94f40e3d7787c4ea9e073186e5fb3a416c3eaf79efd5ab3
zf1621703ae95d5d94a321cecc538c7cffdd04a4efdbc723323eca3baa49ba1dfcbce937cb6a7f1
z7df19093627ebf7504fbdc09eca1b4f0908f04b6a4f77ec5ee1013fa66ae8ff71927d1cd47f353
z0b5362810c89a82704ec10478463a8eea8a901bf5a6dd90d893849488c5252d096bb243ca329cf
z8d6bc62c1e8cf0ed93898a7877623708625d1365d1ef7a4e7cb37b7744ebec5abad52a3f30e5b3
z6213e12bb65acf1eb01c8e5a4fb9354db32ee1fd0bc907e3433d813cf64fbbae383bc701864515
z32bf465b5b9bd0a57d66f829461fc24818306adfbdcaf683c80e7e45c1fb402bc93b90ff291758
z279993f787fb1622a2533d0b593ab52be300a0e765b88cf33fe3e57e575eeab6f5cb743e1cc77c
z107341a878c8b25fa9381363c7319f0fd661e2f921dc8f1fd162510ae706121f9929682793832a
z84134eefce6eb61568a692d92d19f71e3d1195cccfc37cbed3f502e3506cfcd84274fc3c2fe271
zeb6e37be733062e1fe08fbf6e574947fb154a701790e111e3575c2ccab1bbaa5aded98d2003807
zea88b0a3b6f0dc21e0854e205c507201ee65e4189bf9b2123ff0485129b753b967798861a96918
z533f55efd9364ffc62915061742d2430d2ab3fc7058cfc4bd06924707b766a398e91573de229ac
zf8be1b1a2e1eaee76e1c235517c80e35319c4b624ae8ba7091646962abc2c542afd94b1b18643d
z9eae270daacc02f82a9ffb31f2d47ab5c7b4250b7dba65a50cb68f1252a4e2fee06b180c60569f
zde2388cfd325a37ee75b0d4141e5315135262140109c030b90e8e79b4060f4fe5963fe4cf96a27
z650397d4055b908490f7f9aa3c079ec8caaaafaf46c358efda8c3225cc750a53e954ff4a561dad
z31849d2d045a793ef1cc9f2d380e2357d143d858ffdc31fba1fa3f51e2883bbff0d3bfb0330ca1
z1d100107f69bba5388248b1832e27473d92f415c13e29465a26d6d8f2c76b6776356734e13ceb9
zd586b25bcd76d23625263f9e8c62a4c6c408bd2c707527f24174af8ffeba81a28260c5e3c6df36
zf515dcc369001b9b85dd3e9feed3d3c85877ad942ac2485fd2656878fca64807c26a23cd2ee730
z619b9053748de3866b582d487b4f33dfa85f1617cf418a63c5f714785d199bbcdb605176a63c62
z8cd5579f7bf4a799b484d03f0e89504bd77df65a1c8c00898159d669d7bdf9303df7abdfa30771
zc1ac25c2e79eaf85d69aa2cfca4fffdfdecd6b454a75c7aefee59dcb481aa41bfc52ac2f1a66ba
z7550146763978d76e270ac6e6c35c58acb54a9029836535be38711c96b57a618a053a1ba159308
zb73ee5b949574042dcb341a95d8e0953dc64f480793c3f59831978ed61c7e074d645cf9892521d
zeff0fbd859a5349cf7500f146a3589da956d70dd7f17bd8dc1c47fd21460a672843497d004d0b3
z955e106e2bc3403017c8713e11bbad6aaaa3b6eca68b2ce359ad059dbc4864f24efb4ef9e40b1f
z2db1e5b7bd07f680994dd82b21ea61788abe98388e775f8bbe5e16659e7bca1edfc304270abfdc
zf1760e414db0ba7810cca58297bed3abd40617067da40f55090b1579db5afafb873b05e06f26e0
zd317d78139fcb4c90c1744fd4d32b50fff3f82ff879b69e30fe3509a9f9bf553745e34215951d4
z3ab35770d3177c1552d811ff5eec0c2016d0e674444623f41942e6158b1d9eaf46c578a767f45e
z51f06d1d3339804f0d2a68e1aa2bf997154e60b1c4ac4c70bb962b73f8de6342d98043f2169f5d
z646d6415232ced946ebb9221998848524550803cf03632d9233c563730c01919324c87d7490abc
z80944d64b39ff5a98be1a2b122303b940b6134d187a4f650752f603aadcf42a419b494ad4f2d6d
z4e94c8cc6e4a03263c2c1ab5206f555af73b878345316070c59d9ffa3801143117daa1a266f904
zc14375467fac802f048280b6b0c2c1d5a704da1e2fed34d9b5cb535ee9c3b88cf1d39709055e69
z1eeb76dd69658d7e4985fb37d559b917c5f4cb278bddcb33a589d2e66b5aee4af4216f02b20d49
z17da590059e341f6025d83e25f9b8fbfde3ff94c7d66766024ca8a294adb83d1b2aa6bee0f73fb
zc85172c3c35421617a3c25cac1f82763550d3227c8671daed39f8779a7c8ec6efbea0146018746
z815c3c6dff1e918629af522aa8f327e516717486f83152d3deed85998a50a7e2b2e6639d893902
zcfdce9a248c2202119bac1453f6530cf165b13d9dcadb7bc874eef5b820aa8c650143885408331
zbda706b2601f23097895e54123a6303b3e3b5eee92b7ab01bdb9c5e32abca8fcfe2fa4d16543e9
z46722fec801067926c758fe559e5b034ba8cff5ce4fe8fa66810d694150efd149e3b9bea8534c9
z76437f18607ca919596bc2d9682a24505d5c82cd23c375b3ac14ca22a04e4acab90e6d02a19c87
z213764983bff9ddb6514349814856e45c1fe47242d9296a4f58db93cdaa16f1a8aa698554566ac
za284410bbc313dfbd9017b07e3d082139cee70c750a389295b2e39a5d46778ea9bd9e3dbcfb4d7
z9b3ed30d0da5f732311e4e39ec9d07e287a208b6037fca6a3747a0fa7c7db8616e388e07b3f7cc
z9a2a539dea5909f2c772ac84099ba8bf35f8925d1c15015772fc8420dcc7c49c3567bf0b4ed828
z39862fd3fcf89dfb3123b1a2818ba68d4978e77bbfc7a373611676af7bcd8f8a78308c8f15d733
zfcfd2ea4e18d40d618c93b9d7c1cee3417a2ddba8ff33b7d357a431f801b9092e6c0133628d29c
z304f8614188059031ee110bb23bc0dbe2dc55272f567374dbf3c058e8187b1ae134740cb0d717a
z8572471afef6e2f844d08d6e251379868f4bf6ab76a7545d66b5b90286ee895299361b03dfb248
zf8663fc57ffd710088c0fa9d40d4cb25299a43c0c156dc69f806f2e8d5d72234d797821b307deb
zad1b81a4dd134b4732306b539cc0ba71675e31963350e94f9b4f1f67be81f74f7559da89d07ec7
zfae1f9fce9571f27c66963dd4aa9ff6bbdd6b7d5085b45355185bad3fc628b3770a6db949ce3f4
zbe3e668379bf7beefb1bff5a7983657986cd030d953207534eca2b3cd7f75b6e0892a41f11d2fa
z119bfaeeb1763b8be51e76a076b6d5da1f583441770005fa8b3fda951a92681b16e45ba90ea8d2
z3062f00188d72e42d4d42975001c8e0535109790c072038667aad08fc11d452ecad27251aab473
z6b69b3df5952e2325ea4b0357233622d9be6d53a91ed652bac152068fa97d34896e6a3ab7c4cdf
z18df8ecf013a3d2a59088468db7ba551f38222145f22ce010f0b1d8e7a95a70bd628dbac6885d8
z6e72bf3d9418b712775c9bb4bf48fa769e32f325710ac345d043e90a422e58b4e86794a84157d8
z76fd409b45c3a136a263f04784f250bfdb092c36c964812543dcd3675d76412a4947cb04500c59
z5f651b5621b39a85bc4b19a341788f68245e1f4b33e68db2312a47ef857413755ac34f9a186ac2
z07f7c1ab2ce6ac9bb63d69f6e6c9367e84ac78ef3fcd7475d473a98ac454f391f99352caa8390d
z189e5d1eb680040578df684c5f201789caac58becb1630950aed53126597e58f85efb307c1fa6b
z805c73e88159dc9d8e49fd704d5e787c05c66a68875510001e43236f86f11f393ab76771bee4ea
z29322f38d8bb2c98a800af560b36edc091d7e9794a48a3a1eb3416a18633fa6eaec01c6fec534c
z4e2593f301872fd7ab32ac8be4fcc5521210a88745bb1ce75b1e4b984c1ec8f0d946ff221ce02e
zb2e8514f4fd558598c3d4a29f43e6b28182c4fa0480ebaccce01b4ce379183ee8f7e150969882f
ze166efbd1f2847312c2cb2bd7d6965a71758b921b809a937c02fe17fe9d57b7e75bd2a5939e57e
z1f3e5b770cd135b8a00a5a82818ecc6c6cf024a25127094dbc6a19960fc46e3704d2e06b53e188
z93e7cd7ef6f3e6a29fbc27ccbb5b672edb19ca6e911726963e2f6eb03e3217acf13ed8edd479ec
z3595000a60edd7081703888932bd9b634d5864146d5859fdb8ef692fb3b0fa77a3c141629682c0
za338b29f753ea8638f8dcb2d3ff124265f78c754e54e522fbba74288c025bbdeb4f8032ea7d4f9
zc430e06db3e3d67e0119bf7e43d348f8eb63b8f8bded8e105f49cb45e4f9d3b565c19246e17857
z1f7943d8db8327a1e8035755936624e251ec0602cc1b11b4f65457a2b4c47fa1214af9494cd4fb
z9b59936e929d6d5161c1fff43b7a8c70556cdbaefdaa33a287769264fc8b934712755176a950e2
z05ee9d32b72eda88e862e148c32c8617007498e3390a6f2f6d39c68602d24deeecdffc4a9524a7
z6821e777942392e7b5d5ea3b829ab2a18eac4d3bd93d83c1817a3171db9ce3e50c0022bccc1ee0
z240ebadc6a13f15b0258bc985b81b2fb386534c7e38e8d76dfd15c80c4d77262ce0278178639dc
z0eae1266b69efb950721ebd356e0d234552f93422c0d3c669edff23231aee9d9ac278cdbd7d031
zf728c04067eec1337ed39cbed15cf05353f905c5559cae7606af68444dbb8959dd980db2557b86
z135476b9b5f9853c0f9d8cc8c60c05a9b6e9d27fb9737b307a4941711603e0e1348bd22809eca2
z79fcf7685fcd23cb5614f0b6b3ba8537a6e15bf8c35a17fba310b2f77ff0a9388b12b8b98eb8ec
z3fb820f0d8ebdce98247636bc68d9927cfb1db419966b4dc8b7d1da48348bdbc57bfbfe70bc6c6
zdd6862d53d9982e2f0314bcd6efbe0fc860e8756e4c1bd1bba3c49dcd7dd9332a4335138ec3254
z0cd9f5176560269999d19e10c2787f65f1931723926a9c030a7a4a0c3ed3d3a8b0889b247bc999
zd460197897f6a26f1c833d7a971e77b7f6edf9f3a59f0b61a11240f0e9993b1e6d49fbf509b0ab
z07a0e2e82a9b9bbddffb63f8265e30ee3fcca85400c92faf77fb4c837bcb87a05a22c6c894ea4b
z18b5e99ff6e6f315f812fc1b9ccd2b9a27ede3a74ebb2a99e3f8c92d25643a55cd506cff1bb9c4
z49bbac047228b861b2cab4f68cb1a577abce5c89532954f3e79aed652e40f88bfe3000d855b973
z90127c80ebc0e0f9c155375f9737b589836b7e01c9ea60a0fab9f260eeefb10fa3667d570a7925
zdf7786ea086cf9ff50dd34db04f6b3fde5a767eca3dae6b8827413f17914144468cf2be49cf8a0
zc373fc6cffcd9b0ce255ab025a2c4e7a2c25e1ce84e4f26b6f72cc873115673f15ddf40f848e19
z10bb7bb358ee312233854c670798d94ecb985e6860d605186591dda30b06dfeffa5c29d4442013
zc7c891f3a31b9641fdb1d0360db5fb3bf3af13a62e8e9a8f9e1adc659af4fa8fc648a5624b07f6
z8675c37689a22b301a94cd6d11ee75d1b4380824215d1e0d21789aea81b971294b395d2432a8a1
z299c593e0851549ccb81d4e106dc1594eb8961fe717bb156e9c24d81c8c8317311760e0d73ca91
z92df66b50e40125d9717ad1368d0186118d756220de129092b28a10f896a16dbb94962aa6d4ab5
zf5e108d7bff6dc6621c09b8cfa8008d1872edc306f3bb9394766d81a053fb2fea4a911175ac0ff
z27d553e217c5b0b5dd82dba64b9517c1ef0c914b0c8d25ae49dcff367c240a2926ade2f9c2930e
zd63fb6818bd55988c012770a691915f9faafac92ad3b597e851c5d7ec82a109dd112b694a9e8ad
z88b6a3131dedfe7a43466222d3d015e4e1d8f0b48e531f1d0e7305690be4e979ec0333d76075da
z4c351f8a5429fd8d8e7e4e5a3a71ddd976ca74683a70732ce604e5766b1af025901bef2bccc049
z1eed6937162a42a36c953caf3373ff5c166bd5916f107e899c27390e523da4021e4b8e4756d3a9
zb88315a5fc9a2474b5f67ec817cfbdba558427f9668d42c7914d1222053a0cc8e1e341dc246b3d
z89d5fd1fe5747eb5f48ceb5108887fbea3a103015e3de5d610e7ef8563e1f0d0cf703987fa16ac
z574eecaeede812efde25bd5e4f24213e9afa7bc63d6b6147b31110841b9fda5c0e1e71effdfe9d
z443ab5a12a4c0c2c50811d4aa05a9ee466ad7fb5aaec2923954e2813a98d2b55a28a94b791b3ff
z6fc1bb68ac950bb1b8eff02065544b0b86dbf566a74819a4d8d0a5e682c7d6bb9fd804e01e758e
z70dd6f6a9b70765e9bee50a6ab0423feaf7e335802aa2555a0273fdbd58e48726a2c8f04cc23bb
zcfcdb2ab5c1b7dea25171815162532d87fd8a4b1e636d11b4bca941ea0a9f125ec5db07df2aa17
z7170419be0ac39d17b85bf62d524774b12269f425458c15a5f4f7c0df8bd00add52f663a4b589b
z43b27c969689c4dca2c798f228f18d2b0ea1a0fdcf314abf5c2e57f80effa18b175068ecc4d7af
z9012a895d989b06b4c5a3a683958e891999adbbd56a1ac7d384bc762efef798aed0902df0bbb09
zd2a8bbc2ee8156c914bea3b0dc816a625059414cbca91e86e6eed3ba65f900f2eb90ca00fb2e38
zc65d167e0a31f1b2e0ba67a91c446c84864ddc6127ac2379eaa390a8ccd80726d61ad7deaa3285
z30722adaae4abee48f62ad9634ff1bed92e829247f714075fd5c6684bd2767af3159f0756586b7
za299d81c0b746ac7798f52f0e640315cebdf4ae6b617ac153523b29cd7ed66659d69cf9d11a43e
zb3a2e35ffea5fdaf144e8cf86dadff38696888db0d2bb68f86bb5a82ad389501642b772892bfeb
z0f98deb41fed53d346fec321ef477a4d8d48c18d469c46cf0bc8e0118c6054607261a2556ab6aa
z27d6d36ec6826bfc1daff8da9633a229b4ce171da0a0605d2f15dc4c6ca3e5da2d1e6f54953501
zb9dafa1c25633a529f5af8996c3f6634f03db125e56a4ad02582432385da5b7967b6456da357df
zee5bdde8a0b999388a98f60a96dfa9cb5293d318a02d625718ee07733d9f645613268202de86e7
z62885cacb39fcd46deb5880e6d7758767ea958b10658595883571c2760925e95cc88b287d5e274
za2bc7e3a9fad61a8eb52b3e3033158ce249f817d093d15223173c4c2b70e87bd2a94d7b285a3c4
ze86c817f85dd73fccc300f32c8a63ef1af5a9191b6adc4443710eaa85a63e871dd0fe8fe2784bd
z9c4f2f45e5ca0d120bb23f722044daf413e07ec5edd311960116d7e28901a9bdcb0271436f5eff
z3560be6007a5cbe0f882f8afc76d7180a97818a76248a151abc9c12b7817905f4dcbc4ffb75afd
z335f23b25f4bc7508b6b1abc375275b60a0993e0bf48561270640fd4d103866b33211c3d5f95b2
zd79ca3aa58fb330c8cfb25464f1b1f6e3d363018155c7181143b67ed3e72c00734d2546c0c7570
z433a0fea701203a19981833e5e52c82802cf004eb3dc8612da5d468f91170d9534e57f54578294
z31ecfceb967f90a3d9e3192ae9ddc683fdd1d55ec21dcb34813a52530f789c4e428af01d4d1d4f
z2e92161da4eb460c1b492683a67286e3e7eb6113bd6043f8998faa317651703fc81dd8dda94ad1
zbceb2dc1ccbb50acbfe064da50dcd69d61841e8fe0c3b983c26b7ffeb57f9c50c84908a12f1713
z372403007fbfd20f4349f1bf860365b29654f80aeb2c1e1a3957867bc7d8c627369637967a78f9
z9ff1afb49c9e788cb3d392c0f19fca6dbdd152eb843d73f4b4ed701e3de549a26cf80d231dc442
z8eff5eba80366d26d013f1bb74f1164eafcb36beedaf282016bff0d118ffa8b1c09e90b87d289c
z81ab492863dfecbab82ae753e3a11c7c1aaaec6b0bcc52c170f1b8d89e4031eb0817a2e9999680
zf511e236471c3c9c6e60e2679ab5908bd4d2055987d8aa11665ee3067d9219273cd23b19454169
z3805e0a447066e9e361bd2ca9e810b599e5b2307d33199543f86655081124c461f861bc8c4608b
z5fa93a9eec15143ba7964bcd1c906182308a781219e81e299b5f4a50b964fe93661829c599ea56
z2dbc3b095d3cfc91715b334ff2a0340f0f1a2ca5e5c05bb8850eb4a34e6eeb2acdc0885d0bb771
z702feade284172194925b2b75366406f567ff2750b4e361da4dff98a406ea136295d353d8c6667
z9d7cd4711eb118b77cfd44e84c9793ba0d1004226b40bbf2514ce847595adca9781ec61bbb3dae
z53f0bf63512be4084737ddab1ca3cfafd0df869227e347cba6b3514625b4a874935d13030f1495
zac0f4ea3b34702f7f04a5bdfb2620685c2271f9cbb15941b851316adc921984b1c601a07b0b919
z664b1f229990cad305d939c8aa129605ebe1bd859c089962a0cbc08416597f908b1166659f0c49
z8a5f5c5ceefb0194fed22c72186f18aec39dfefc9ee56eb4accd880d6433fb810e0aae59709e78
z5db3dcecbf730ca811c2348a7a977a0ae62bd32689c0c2275b1c94015278c3fb4ab439c1f2b740
z5b98e938d495f9d6de44bbdfbd296cfbb29aec1f64913847a7e824c6b1ada20ab07e3c7b08217e
z318012403d6c8a16ba7eb17752ddcc5af7c556641a9767d4a9db3ed71d0043f338a9308cbe8d3b
z3e4ff9deeb257a0bf7937037b78d729f894af2b0dec592a6b55d2047bab65449b832bf1446940c
zdfddebcd438d16213726b3e5e5b308d3fb799fa4563708013d6598729672fde450803a3aa5babb
z27e15d4c9ee970ca1fa7177be074528f193572ba95b6ddff41c203eabeea108dc84764aaf13e3b
zf81c32c6e84a08ff5964c5987affe1d20ab6be43450139522923d57c3561651e909526ad73ddf9
z3f572da2c2307aa8caa06e7ab590c19f90479498922c6aa710624ef7d27815a300df669f576120
z62bc1fa9ff25c4adfbdf4cd565b6d80d5d78d8d838d676966b3b73b96f1f5971a113979b012e77
zf611105e647adb79bae067f609e64a055016007ecb5a2babf7ee6a759c25c0cabeb84ba4e3b3d1
zc20c1065c37c48e34b49b60e805bfed29ef07b87b5bcb102178c1eb1953f9a5f04c1c61f514eb4
zd56eedad1874cee4525679d0dde95ec0422b19f4946476376beb7054264485223637477c2fb6c2
z4e8553d2214c9014a31f72aadfcf85286e6f3335adaccf7b4774922f48cd4532d9c2eb08653986
zec023e805e5ee806b2e3350b9727539bb9ca235ffec008dc4ad789810134cfead69188eacccf9b
zf94fd7f2bcf37bb55dad0730f7f97cba3d46548b8a87415d1fd036c923d91075424bae672398e5
z9385c7c6f5bda5fc2c0bc200735e47d92920816aed41cc80d830a5cfd15107ab66279280fc8bf1
z269f57d1ee709cbc0bf30067d532323198fb8b671e11d8c2da5fc1fb00adfa286d2d51307990cd
zf82522cb705253fab407dffa7a58b924d9f211711b07ab88b6530353c1ada6fc7deadf87a72c16
zf3333e551aeea71c0361dc6362f98c4554facce205292c61b60d3184f8960973a0a6b4fcfdc80d
z7f63355d45348bdaf298e15f121c98c1051492b3df2d9c6f27fd1d8b2bc9fcd8b1eac2f4e15bf7
zf8d07c661f2d1f96f9d72c131e9ef4c66b294a95715118a1c7ab2ff7611c13106a31d4db0edcd0
zbb97c9c8bd94c340819bb28b9c63396c843fef6eb8ea62fa646a532ad9696e5b2e10f873eebb74
zc4ed10964d5a10836eafe58645d4f0a59cd3001f9a0201f9bb7a04ef5d8617697bcae2ad5503d2
z75c3600679b6124087e1a957a6c3e7a4b711eeedd18a114fe1f322c07ed37b93b106d36cbc9301
z164eb2a433ccc521269b35224b9d740d7b29d34666190b83151d72f29c9ace0c709b52b331d3df
z33f5d70b3c0f6bde62cadeea510fd911cec563c13c67220c06e8dd6f9797e28a671cf824586ea9
zda3d6a4ed98b7498ecd4e113d0ed9ad6f150c3dac3655c302e812a16d33e817ffeed3f4082ae7e
z148f3b5f78257c76426ba41009c27aba2a03555920e39e7239a820a8e05306bd913372d7bafd5e
zb9049790707861fdbafe7961c749a8aec7a17b24d12a970458d0860526b27ce6f67c0f77d1e47a
z2fbe68c190be39d634735cbf54df7fdf9da2d4849fdae9cdcbc7b8ab870e95317a347696dd2c80
z68c907c5a54f9486dfe7406b92f843ddaf06cc517a3b9532a0835fa18e10ae589d2fad6e430215
z4851f14172ede40fcad448fca6fab6757b90b81c19aabe6211f29de66e83da7a6dc2a0d7c2d331
z483abea229e360fc2d13c0320c334f1a044fea5c0689e99a22e5ff7c6581496f7d2cb8e45c269d
z88401810ef9c1bc4e25f01f8f99859a059dadf075de8b2b22a9b6d4376148da5179e682c1bc610
z3643940098407e8f1b3d9291d3c5be086e9ffafe4307b477274b74f2b8700e84e4262632d67bc9
z12451fd98590259218038880f4dac3fabbe92b9041ee00733f5d12836b642aa457c657fad795ed
z48bf48389bd38327a6448e7191308aa2d80dc07795438ffee9b0e69327594341bf65824160b0cf
z4f2fc8381d1813c5db39ab38ca63125294969977bd3ba8561750f2a84829e3ecc292b4e0b3ff96
z8a2d866584a048d5dded9a29d47f6651bbe14791def813000e1a44c49061acf7148ecfd3387f17
z6993877486d712251c102defc29ce25d9575442dc78d8d02a7578bc1478b3392f2db6b3d978504
z5384bf4adb3416fd6779a22eab654bf8995e2da6f431924ae7734ec711ae4883b51c1ea3447c28
z54f530816203200aca28270316df85eb3e36d4dbdda1871cd1856571461a3343a40fcfd1396335
zc083a8578b57502107c0dc18080069c894e56f2dc57e27a408ca9acf368b13fdec7f6c3a8e0c7f
z89b8640b6ba51f0047811174039d5213ad42060c293da508aea4dde93e54ed2f30ebb435363643
zfcc8ce14dc88534157304616a498de73fba289344e10e370a3885bf9d97a9e0104305e10a1b8af
z4bdb301d1f79ec7a295617a63cb33f57e759d06aea327305f9259dd75712b7257dfe3e72c872df
z9be4a9da0ed0e36ac1175d68ae7fb563c05e3c073a5b44c9ebf01767254f942b082246bd782fc6
z4bb503f816a5b678fb8b67fe80aea586e98b06febcb0a1ffaeb0e601335e3beed092812ee6e1b7
z923816736001d615ad5afb3c001ec07379df90f13b66e21e3f93da6d45f4743256e5ee9c2c46c7
zcd752950146c262b6f0abae1e3e247c9edfc48dcc0f563dab85540c94bfa2aba7d2436c2680d76
z013302c6bd3fdf7e2bc564190fd805499895870e2408507bf6c4441bb4c7b143b08e53b0d479cc
z8e72f49bd522f8c5ed59a13c041643fb388367a166b36b2d751248eb16743bd3d0150821e39064
z1f15d2cf396446d559fa703a764a00db6a1f91e05eac7b7d5f9e2d725e43b6afd01b7e8cb7a18f
z1abd35d4e72564c572a4b2159f388a2094e88aabb850b65edfbf166d57d6f2fb05e4afb9c5317f
zd95dfbe397c513b70ae9e005fea3f2f41a7e4bf3843692ac9edeb88a719f02b6f681284dcea28b
z5c518057660aa0c54be79969469b1105f88fb650e037c3f0c1e2b338c94abc5065cccb2e0da4f1
za105158ada6a1e68dbc8489ac1b8dc29d220c410bde3ac4e77cbefb44175f4020b59a940aac276
z99ed1a4a0bb24797e12b08ce16cd3f2615f05b4687a3d72fb4f687d7a632752a50c58667b4b3ff
z71259293dfb93421c3b134cce437002e7c4d0e9805c498c48c9f67a83103c36918614112814d38
za6c86c766ede750db79c6d28658fe3864c2f6ac92e70f654c3616a5342c132fc2f0308b158b056
z0cf0963b0baac782f872194164d1ed251e776dc9ba94a2254798c1b123522839e5cfeaadf7b822
z917eb3791485fde1d4ad475f7995c2c344f185c5bf57dbf68df60ca02284c417c759ec2d1cfe21
zbd65d47f81cbe97ebf3421a310a756c56449740a53126298a1d81077c0cd662162a2189235cc91
z8603dd2a3c4fc629ca1ce516e20e631762b67ad215531836409fdbf3c5788a83dcaa8a9592ad11
z2b9e15c41f91a431d8bca7f5bb199dfe58b5fcd5cd0f685a9a085ac519eb35faab5a2168f1d479
z1636aa54fc3919779512520cfbc96301e2a7cf74309276721676e62f27308b6643ee15e0eea50e
zde40117da6c2f04cf1c5765cbdaad8d3ba0d1c3444bc2f28e80f1425cb92e34d936d0eb5a58a7f
zf18540b2fb08ac33eab50c6c8c4b140db052b9eee4f289e60331946f44f701a047b745b5d83420
z9367b0d6890b3c70717ad994e5149a2501605bf6a13d32d2f5c13fae137610259b406cbd491b64
z41d8df0f0f5b74b2ed7a9ba33a24dd86ce8cb75c82a6b2c745beb72c07b3db102a2cf54e938580
zc2b2c99ea081fe518cc201392439b656c0bb29a7b6d9d6989f8db75603c3487fc7ecdb68f496e7
za462a190196bf46973a8ea351b432a1aeb703c58bee5febedae053884ec8cb84a6cb0bb3018d69
z9585b56ae188746265063832b14552628a1bfab5938c44a4482da31b65c12db03c608ac98f7230
z8d554003d5ac88a71ff7136b10a0a72b6acc2dd1f0f9714179d0f5476113ce45fae1cb9c445be8
z68758f8fdb52a498a677008a4a28083f4c6233719cb993b03ea794d50af304e7017fad3c2a6ecd
z87fbf3ea28c320fe429cc21ee0792a0d81ca6c070487311373ffc70e77fc172e62fa3406f66f79
z912f46aa25a7c40ae90fda9fa0304cb2e9fe28d4b4bfd1934eb06e83b49a3cf85d0d580501c891
z7bfcf49086c0dcc492a31f13c934a31916cff668ffffc77147f08f8655ef10807af33656cb69f6
z3949500d3b396c703d0952ef846ed3945871f0e5ca29e2cdc0af9afeaf36c4f98c2877672070ad
z6eb4c336842d18d7b2be1d14e4260a52c12872c72abaa863bab06d7de8a322fa46fb117e5d94b5
zf9d30201daccc80e9a76ff7b5aba7ed0e3d1941fb5cec55e78bb3134babaffc1af38ad4c46f635
z8b5fe81e8cc573e859d5f85e00e812db9a92e9d24e7c416832149b1d8f40f736f12517c1bab286
z2bedae6d5b54405c91a7df91de8aa2ca13a62ba894a83fbca81e1f7493cefbc147ebe5bcfbc1d9
za015ddd4d56d764de844014c3b8f55e4333fece6c3d11ac9ceec749944d052ff46e8ec0c96df84
zc7ec7b269e25d678965619513da3f59119cffd9ee8ba9bd8d96ab9fbb39f9326e1253f28be17c1
zc945698d9eb066a1af98ad0d8d99baf977466b9b83d6d4a4cfba0fdf0002dba991c9ac2ef58c59
z5fd416e783ce2e5b6b4794348b954249c65fab3430aa3f32134d99845639f00850cf9606ff0896
za1a0be64b52db0bbaf0b00b7bffdcb35673428e44fa3338412b16aa0f705cf0bcc13e82e89be22
z3f2dd0ece8dadb5b50112275633b8125701d67c74a2aecd18ef18b8d4986e1d7883770f6947bc2
ze19691445dddeada4a26ce65459959704be990dd39d41e38b9e909c2dff2b463554368afd519c8
zaa9ae6ca7da6f70905e1525b167953a7a72e4551187afc241f0f8fa9809c1dd676ee78810b7f66
z03e7636a8ceb3c09c10ab8e8b24b4abcfc6dbfc6cf548aaf1645ba14792a42e953f743c4c1ecc3
zf35eb46309f7c76001732a86d3567a85a2ed6ba9db0d23196d33f0bb8caa4170922b5ef91ce2ab
zbc11c05c4c26ad32578bb7595ddb97d7a43983425e291af5d1fa7edc0a51c18effb44425732286
z7be8dec3d3238c88df0d2763c05a1a2bc3713f8858c979e728aafb7d54fb199b03920c03e812cb
z6aef4075967666fdc3a931cecc1090ffe3e02742f3d2aa5460af7676dd3cc3d585871d8b7a396a
za00e6e8f6254538ef0fee1502aa7915679959630b39bfee913ed9d4eef9964bb747c0b9e1f22a8
zf70d80ce4e211bc9e466c89995846966d2a396ef6778606fcca80bcb8137d7cfabd0fc24ef9300
z83382fc7b4471e04ab93912284201730d35b304597212ce83c76b718e60f328e8a441b4ca3d339
z9b8d91defe453ebd671d47de0c233b445d58269276a34c0ff3152c62b0da81d760ad64dbad9d98
z940effc3e44e78d3ecfd2fb7eeef6e801f467e426d4153ca10e4616e565406f42b612d99f61771
z2c156cda1ffb9dae84d9fbeaa5c73a0e6b3046b524f7f7e361832cb50ccd6c9e53cedaf6c8eb0c
z56080ee006abeff7b4b6ee8becf172fb4b99f5d9eaf5ea1d725fadf8a3c1441077d175364d81d4
z67b26a1fc7daebf3ef972b8ea4052cc312acfd16f2c7003642f958c5059aa7c20279b78a68e775
z66b2ed82fbfc4cef61ac4dc8a764ef7c92cbb93c788dcd1c840910004caed05accbed731d43977
z6e60e19d0396515d611928f165a5d7e19615428798c939b3238dc9da315ad84955620f7e29ed92
z28a16ac8cf95eae7feff91758794b4d95cfcce101d75bbf24670521e481f0dd304f058d8f9376e
z1850f49d57b26cfb74fac5f9a38aac364e3f3179d61de0ebe2631b79f454e72808ea279366a6f1
z73dc25695b7e4ddce37b0872512146e700bc21cfeeedf064591957f6e18211661f6b7080a41a79
ze50e5b1beab0ac5482f3621f4f1666ba12864de5a5b3baef758ebea91307842aeb3238ccc8da8f
z1034d3e730efe4be3c97659c46c3f13037fb1155e7a01e217f18d98b03db00be3af9a20dd11918
zbdeed6d93207ca9d8390c9367d1ce71ada9c8e9b4b544d4ad86e4c087a7d061d7ad814e96ca28c
z1ae3cf9ae1dabe56ed357115437dbb7a8f18172da89cc996e28370178e5bf51e449daa8abb2019
z398836e9f258de37a6469cda9c07a363196aa568ea462619fc55057d14f31e043a1f45fa1db28f
za1a78027d908f22793bcdf4be2d43117ff595ffa7a84a5fba588046e99f6e7ed23693084822ead
zbd5b1fadc86ed8232c84007a9a91d7066bfb4d7c0a2c521ae62590ee5a1e748e0ae9e950501e3e
zc3b4e29bea40dd3052ee802cc48a12361690b7427c6a10c4e34600b134245c31b48b7d0c8b12d6
zc570208968d9ea42b19c48b1854fb419b588007948c04ad2902af6a75e36ae69d757d6d4f8873e
z00a0db2adac65d78ee925a17cc928a460f452911add4910713cc37983b0304c3f7674a67516a54
z8fe499c9f7ac1c96b32ccd864a452a3d5b1ab82bf6df3260f91d66d364df37dd1bee48cca0478d
z61c5762e518d6ad7bfc2ee67cbe3a5eac80fb28d89b1717d6b38e44ba28f6e84d51631d75feb0e
z01b0a296ff8cebffdce20917c21e0dfd30961b62f1b22cd0b7c5f0566fa4a64fcadd7e3d87b048
z397c41f21eb0c180cfb39fa499a33caaaf904a69f4d212e1a5e5056e2652f4564f13cff5b378a5
z12845f570ec4a2235e2914564aaa46d5afc7f476db01a41b1620fc850c6d41b0fcb8e55dc7928d
zcaef2f48d30646c8322e2ffb9ff1e75d35513e9a8be3d6fa0a2ad42a58c2bc97c95a42f1c9fb38
zf8472d734c935a340e6af7d82db42fff1f7f4e02a16f1b4962718c0005401cec93a31a9fbe98cc
z1c3971a97a42a8139a542aaed10d74e1f419d061683771986a2fc0cd5e6ff4ce5db6d002661d7e
z607ea8ec2699f3ee654632b07806f04318eef9ec36881a0f620e6aefb2ff88e386dc0fd916d8d5
za77a5f7d9c97d65202923c6c3642ed1e4c0907e9f556dac70223e6e3a3f5a6141c9271c509e165
z754fa9eee2c41d49b4a2b93be3011764a32666db6473d950de6c44af36f1c6d44c829f5a0a6d27
z0e2a04316272bd01701079cbc42e721e9328d979bad02ee3d6fdb547c1bec7a32c7e7221222a50
z6fedcfe3567b8584739eaef0fadbccea9c7f1ab476cb53fc479e2c9c818cb95342cb24e48ff2bb
zfaeec4b2321dab43325feeb2230dc429c1b2b68fbf0fd15b161b39e3ae490b6cb635b0941f4b08
z328d1674e01e2a8b147e82ab58bbb2570be11c03411cbf087e0e9f9a476d227d7c278f0027347a
ze4e19ca833d47dbf706812f35462110175f7ce77744246050e47ec9a3aee92bf864acc04f2ba1a
z2d089fd5aad7587ebde4dfd3295afac528671b37beea6482525beb4101c83c128ef78a89a5e9d7
zd205103227209872846ea2972c3a2650683497789906f1fe683990c5ab6b483d3b0d8c9be14a4f
zb78a63ce6cc8b29c266379a343b9dbd386c530f2b3dc8919a1387ec50a9c2fa5be093aa50d1309
z2ac1f20cfea675319eadbeb2f1dbfae62ef04fdd359ad725ec78080055f18604ac44f272b68809
zf8c47b35dc127fcd14718d1404756ecb0ff6a3ceb57f6e7d130f579281c1b0710df479b32d5a4f
z4f2236d1c26b76d95fe65788406eba3df5ca113a3debe2caf79326b980f8d381c7214b21753cec
z24d45aae2647f4309bdffa76cb666ae719faad73bf80ef88ff8b0fdccf2fb998a4e75984e2dcd7
z6394a39cff4fbe3260f99367c2b600d9fe502e5c228eeb0b23a244d82d00ad3ae44e468d8460b5
z82341b0205c79072cf881a8fd9ce9c07b8e935083987f3d08e42f000c4311b9186d903fcee4489
z5c64fab772b79685fda584b617c2adb58d647e4fe8d80464032e6bc47c64a568934c00c56a54c3
zc891c51b12a5bdca0526439d4efccedd4bd53e25c9d466e575c2b5dfef2adf393342d8f1ac0916
z05ed4ca8a56da97da9365f8740420b6d3ff40755442e04b85d06912260f258957b94d24032c987
z6b4dd1511781da17cc6fcce78bdb001274b897e41556fb2251e1f587add3eb988840b82c369d4f
z2a39bf5f3fd3e4bd2abe2c9504d85c64bfe337655fd58aac210bd824dddb5718105b81ece58f8c
z0304182dedba34fa7c837f2cf1fe19544fcc2ec14339482c70fd57395dca087ff8d30975f2dc48
zcba1f356370e787f1a61b738c34d832ef5bb99e52916ef0eb46514c55991d2dc5807ffbc915290
z38a35d8ec2951a31eb885bc2ac078d6ff301cf8c87a07dbe297b66e4f3894a68cd03f4a5cd2c33
z1d2ec48d05bc1cd3dd4ba5c87d80f1d938f9f78ae386af82eb54a93da7e61b99b91419324bcbcf
zfd1e3be5eb243230e951c169b059857e44130536080a89bfa379605216ed4014426e208b3113a0
z028e8a0b05ba2f6098f30fe5ef89601beb0c8ec311d748b105e7a0c84dfb469c08a72bc6a8fd4a
z656d73236d2e1e7bd248a46a306d62114c38e9d62d71662e9e2fb8698160a5e04e076abf94e289
z44558f931d2663be44d6d66078e7bbbb820bb362efda0b502ea5b937b6161cafd2c3613bd75af2
z7dad1bd9bc74c3ab8c333277c1f0314a518afd2c7989f0a0950a3b1fb0655c6a31b000b5680ad5
z54708f02eb3dd48a22db224871b0e183c286679d9956217de3abd5d4fb9ca82265b5f0b61aad55
z7a012c43b77ff5952909e3602ea24711068fc2a6bb90af091df232201f5179a1dea6725229a8b8
z1f460a23abd2abc35e6d3fbc5e4fe0af16738c6938970b206182c679017708301d42a0ddae91db
z309d841cb74e35d2d636b863fa8e0775349b144c8edbb3e5f8bb24e2760d7ac07d9123946eca0e
z3d449118f4dc3b058913ea75d668d93355cd65a00b77e1e813d63b71406f259634198d6ef70740
z30a90a75b955a6d16c60bbafd9495e9f6a7b78f564465a091aa78431a77dee0e7adac5c1c3ccbf
z4a256b3d156e2cd66fcd902aa0e1a02ed45c589fe048dcb994942e1a9397e546a04a703eab3c33
z99540055820759e4fdf9be06752bf52046996db3ef0e5971af77d07c9eb729edda9bd5028f4d56
zb9e2da712faf758e20d5b946f9524c02048d5d50ccaa77d4d8d9ff296318d852c1e97ff90ab5cd
z323122d38ad7ec3f38a2f06dc6c55b5d24df49c2874899f4a0da92fe493804b457d9939b0fea66
z120cf132d8a26e7d17538ba82104351b9a4b588f9488c890c924ddefb858e9fbc36618c4bdfffb
z86ab84d4a527d3b22db3d90070d1f5a5abecffd9a4d5bd87a6d567c0795d8b7729b7af89a483f1
zeeb1a4564e6aec24e4af7ac9846061e5f5f375929d612c23609208628f0d424a39470213c75314
z26cdadbcf9ea53ecaca821ef0b9fbb04bab59b10cd31efe46a55f5da4a3a6c91f012cadaf34eaa
z716b3a9617c45d04571d27df37222704db0fa3f44fd4b18ae8781b397b6e67443174b3578272ca
z0cc10ca0cc97c6ec470436139cb8d69c6d7148997ddfe7d786fd1cc424c729af7d2c96b8c32cd9
zbe938cc94cfa287d33e8faa946babd6abcd8f1d043eb70f89c91c12ebe413f6920fbcce2f2f1f0
zd53886c0eac27391cb9abda3d35ce611df9ab5cbac2a472558543c524dcd318f47de6a0baf7590
z06456869d3efa164341bd4b6071027873f17dd7d03f22086adbae72ddd711ccdc70706a27fa644
zd81ed4b3869fef05b65a79896e826081ca4f75a397b7f1ea820af20c95e0e9da68442b83d15ab4
z13915e75e0847f81fdc0a26e2ee1e5154d1096176083eb51f75f6cf0bcbcacaa72194f5526b9d6
zb49d871bd7c115ab5111863f71b3d6039af67638711f5894013496b8a322c0aaa834b491240751
z5943c507be7a033281fd3a4d86e1aeced2624f7c16827e97cf53467a1ce8f784214b342fca0771
z8c905964b785bd863e89b6e30fd63cb5b64d82c6df7ca85618d9b731b70483b5fd63986517e4ef
za9eb5e498dff7c7b12fe3df0f18d3a0ae28c7638f3c3f61c347d28e29647f5b8eded2553ed77d6
z8a022111346f540b2fd5e45228c68a4b57469ef4dd5ccb42b39efc076a3551f32bbb7efca74f72
z473e76d9268c111b0f31f95debaf0d33d186e59aeea57bb48eb7450a01decc5ef1761b3b201699
z2e580260786f4671db10ad8884881cd486c9829bc79664d906e8943085ec69c83df975cf17c503
z2bd7931cb6176b4930e4070ae1a53b84f6ef13cab92b3910a8b55a8959a4cf4a709299ec1b3728
z65fab2b297c0949d45f49c6bbbcc14249a3e960faa6ddbf67dded71cf2de3d744a0b9cd9305017
z6e02769cee3bb87b9b0ba42ed714f90db3e4d04c0e690e5acb2da2544eef38d9ea7b77e453e066
z0d67c6536619b594f6799b7a493d3dce454b65665d2d1abf8b918a049ee95300bba760d882c55f
z279aded338e8d9b60eecea15185e8ca1bbde5f2ed1ca1c826f3aeba774c1fb2c90b18292e6c3b7
z8eadbd620bf84a811973c1604b5ce995650b00d115c395e5781afa18a46dfb153f581219462d5f
zb0f7a91083bbef17c9c0b6ffb0ddd882cb299fda8bbd68d75e8d4145a3df6df0a6e944c470e50d
z1e45b2c9ced7b9238f05dfc6b85036833ed3b4d4ba80ce1e8e02c92b5949a2d215cf01db3b33ee
zd39e732aa53d4b3e8b5c3f91bf416e5e4f57d0cc7809a35ad2bc337acc6293585daabf00d7e3d9
z2f64e8d924146d5a05dc9100a4d570c4bef572914c25485fcb3fbab88a664b4c01e42a3e2ce398
z2ed27d1db68788b590e4ae3934b7585d1b8e5442020f1fb1e55be4997e57d7e5f24cb8135df2d3
z64f4d4ba10f037b413155b0b28f7718a34275c965c06ea3444a752a2b67ace85a06c904140b810
zdf8c245c9269a37c3ba5810630d4cdcf31957f6f34deb7ac603d328f5c832787a6f9e96461f96d
z3ab15134d28ecc03b169d204f73e01ca164d34e2fac1aa8c07361ae2f15d0b172bc0ca46515cc5
zb576e23d13de27c2e477b0a0e9e72c3a57ad709b789dfee01b9ff8d4202f88a093b49f855c6638
zc94ebe0a3f384991e0675728ba80c3df7cecdad773c6242146efff739a387c460261abf264b6cc
ze16ef9f7925b7f0c9853cd9dd24bbd76ea5ced67ca1c2800a0b0c5f313f60a85702463538fe2d7
z416fdbb22c1c4fd99ea792188ffea12f8b4a2359fd37a93ffe7d34cc50918f14af404c711177a0
za11c3aac359ff9e9bd00e9b6cd59a3f6a5ccfddf3071ab7066ddce85e742659a9c178350633fd9
zb1794ddad02dd3b3782334abc63bcc46f96b836edb029e8d0c33ff622ea5a631e351beea06f429
z3c64007de6a3a2531763fe50869a9b1d059381b728fb60574e6e93e595a09933c4ac4fd05f7a42
ze59a347d3d6eddac7268d1952f4e7644bff110f6f94f3785bbbab690ab9830855afd854486a6e5
z5db17f34f6fce04cdb6b82a6ae8c1f9461db5d452a04c2647d0224ec7e8c0b815bf0ef900b6444
z560531abe3224eafcf023e7d927fe7f596c185b0963cb0ee023c8bc2291214fdfb200a80e059a0
z079306304b248963f15f2c2d10e996e8e21b252d2eb6510ea9ba9e587e2b2c654f2129a78a57fe
zcd5bb55e9e6386722f0b8a5b303e634b6016032c381463c2d94506cdb457687af7f2bddd174951
z23a8ed514f4a94c15389f20af5919a417a41b94cde2e91cb6d0facb204be8cab19cdbbe24f848a
ze89d4eff295f2fe7b252627d7bebca03c5104ddbc309bd1ac1fd3feafd8982ddf3237928fa86ad
za789f9bde1a35a8863ec7518e27d890128aaf13d28434a4210e3e8d78023eedb7e8af8da9d3438
zb35973fab115e3f65341d647623ff321ec30c6953a95421c344d9825c138e3b328dc0d78575184
z73046034da2e974641383aa8927025f9c4575e9bb8c2d9ab2c4008b02fe96db26e0885b90b6199
zb4772020a5ca548bea2f877bebeef7a9cce0c619bf88b32b9e74568bb980c9f977b3d68c01eba1
z3ae3b221e5eab76b190899f3cd917ae47e98fff68d58e1189767fd288e7fd0dba8174d20c269d5
zc198b1e3912f40b4e9528994c2aa2759efd758c1c6ab8f09b249e4e874df7a4b50a86f8a09b43d
ze1582a9740480bb051c3cfe517312dc83fcd352d3eca881c74e21f1c3e135da17dcd136a3c8e4f
z7d1ff14044edcc9f499d44964e83b510dd2b02fab0ef7b210bc33ad44fbb70a91d04623aced583
zd37ab2eaca41445cc63e7e277525a455c1694da1d48b214a3e7d711723674c17d15dca03781982
z9d13f12b2df575c44e63a0736e8cffe079cc84f6b067050f7c9368a45d0685e318c959aa651e42
z7dd2d3a668cdb89aaee4330fc75e49adb38c9512ed7a04fccc9a3b228a092fb0494703a5cd5730
z491888b749f629f56166e8fe6d569d37ad181de1d1f2ca99a5916771780d10d82c06a7e320e797
zd3a6a1935ba143696fc1924477230a5c4d76a069fb9f8d5947ff670acd5722ce59f0b1157f14d2
z4724092627a97b9e20d47baa54179e5c166c7e87494f8fbbb82024882918622df2f520d0dc0dba
zb61b08bdf6d81b407732048fb349ec501d3ed05cacfeb08a595314a7ff316d186937e8b1ffd9f0
zf17ac86becbf5b1abefabe58cfd9b179537558ed11956d0e13fe021d8cd828b3e8bebe0f954b2a
z28876a880e05ce729669658ea716b10e8ae260306cfc81125774615eb31ec9f815b06c62c788cc
z74d0b5a63fef62764be0b93591a0b3d203d41a43f6190c6f876d7aa0c6ceef92a97f38af61d0a0
ze48fab462045f5f5ec1677c3dec9e9359c658c9f6b713517b8cdb89486efa149bb95bf0b2b1485
zbf5e15bdc575248a6f63a105ea335a053c4951dc67504c205e2f0aadab476d691cf575b4e65cc7
z19c6faf81b791f038513725707a220c2dc10dc272c46c97507b295b0d0a5710cefc8788e974843
z2ba71836a8074979f3df616a32ee818b5bf94b77b592d2e6991e6c2585e11a5df407c3c3b6f481
zd32c827aabd85523e3cb71c53b5b4f14375544acc2de1394c28f53c9145c61e48b00828475bb5a
zee36a755a3979b870ffcfeb73f475dfd2b7c1568ba479b55f171fec4ceca5cf695c54e5913d3d1
z78ba4ce1fa7b69a0973c96c1ef492a1339ac1aafb7d09a56eb293e7ff2da9df96351e5bcb356ea
ze542a039f4b87b735bb9a5883251452547c95720097f44945195a368f1426c0f239fdc2a2df8c9
z45cb6b3b27df748aa1356f0cc4e93d463d15f9f8a4089bb94df8e083f48a50d9d22fc5c2dfbd7a
z1af1d7ac8f0a9ea39d5a340d4c28069ed5debe1c0fce917601f5c7139b594b3afa250360fba303
z8730a65bbc52e49d053406f64ef86a6622e95c911f7a651834c95318d101ed2486d3ed5782e65b
z83089841d326d66982e8f88d56d8bcd0024de24a1040ec9c57c039e04c5babc9129fac56410311
z150a6f4b4591cf9820b3aa4c20835ff964fbb34677e1bd4f6ff3e3b7801afab893f6c4e8651798
z723460cba5377837f59ff72e0acd584c2a32ba003cf417abed2b4418c83eb0ada89ea0e9fbf0a5
z9c1a2abca89c9439392e5ee0a394ccad65b0678dc2d0ef1cfe61d69ba175dcba37091ebad56fc2
z8205cb4a6cf88b169b034a3915de39729f1b7254cfb8e2bd3c2b5dc87674f76499a904d38f10fc
z468e960f50010c3d55cbcb36f0f1fc77a0a664c376ca250adb1ec1dabdeedf2ba5bc63334c72f9
z0d813e3ba213c96e98a6fbf13b9e715aa7411d893d9beab37a0d629facdb265014e09b8849fe0b
zb8f26c566fb40c5c9a835593fd4b1ec98554e41db452a7c38f9917e575861b48a7b707b27a26f7
zf4f1bcf268cc30b45ec1e5bf694cc89f85f44ead1163a9fa004ad145e1e47f628b25434a2406ac
zaf8665c3bcbadfcecd377fcf855f12c593909840dbe76fde5ac9993edb9b327cda6eb52272f49b
zdcf0f668d82cd31998f1ccbc5c6b7f7f59166bcf7888b7a1f11d3b580534600c70ac57449a4592
z96c9fd57cdb77ec7d2a3fc8bf4a21fd1ddba61435754c19d8bd7dfb98cd28d7ef7f1a95c5f6bdf
zd04f3acdff95ce856de252202a2898e956cc28d0d4f96371220e1d91fc583f5da59bc307be9ef3
z3c8ab734fe2b5dc21c35a0680539c5a044f66b30273401bc280d3db8a553102f51f93515079efa
z04ab8827122d7946c4aa8d027f921988c7d436adfa92afcf5158ceb5bec0638c1f54b5f4dc7cad
z2c8432f3e57cfeb8f8a315f17d9d21479e56268618d4abc95ce0815e9d2e4fcdd9a10ba78ec782
z04119d382d2e88b2bdda6bb6f465418f340d37154d24fa03dddce7a63a888a759b62bb3961551c
z1c08a51ec89abdc9d882976bbbf99bec7e1dc6315ac1c6d5a2a986ef08abee31414ba07c6c53f4
z31d4b19d7b5fd0479c0e2a949fcbae6eee079ed650f57dc83c46a3fc89ba5a3a123a89afbc5505
z879138246f36c04efe6b570dc91f4bd1dc6d73a5afa66d4c593b0d98feca812738b61d2efb1290
z902df1ec64b5e00262c7257922100c9bf3da22861ade7f7ff6ebffa0457397caf5b3120c08ab9c
z316dd2e14a7899205a99cba24242ad831dfb639bc017b156e75387fadbac7ed269ad5c0d45546b
za1c4ef3a1e1b5e0f468e5099d04888fd2d103cec9baeab97f9c7300f2199fdb37b19f8dee209d2
za740b89f0cb29c6e5cbb3037f63566401fc1bd92bbbca1b83f7cb532e1398ac6081c7702e301c8
z4a94a8bd1db65f57827cdd71201972ddc97dbdbf5cd5e652f0e00ad25f3ec9c7da59c8b94bf4ee
z1acd6f53fd1075ea490bc6ce4e1dddbafb3269e144daab56f669768d0d217108ea5daddf4b9904
zac61aca811c7127b8a49f766182cefa18de12ddf39fc7d0552e3415553ed822191cf5e367bcd56
z6d9112d276ae6c096aa630aa6e86a3df304d86ae5757ec188e4d737f9d8052984dd22279af8b57
z4bd887c534ed5edc83bb90146ec04e6d161e294913ae1b854097c6b0a4299274890c38284f8842
z4f29db447d909d36ff8c37a1dea179ef02d3623888fe0c5fa9ad05aebc9859dfd0554c0788c830
z146c64079653a6c2fca88210517965f6edbec1cde82a89e909be8a7ed85a4214bbd93b3ffc3323
zf8c06fbf81c2713175ad4be06ed9bd9b3cd8f15a051e3db6c71d3bf7e81a7304b431f308c33f7d
za96e660ce94c3d5048036e3fbc32b674cecc92681c510c0abc5ab68dfab704f3f111f0de61dbf6
z760902aa681489148462675604a486aeeae63e742a5ea9301a8a730038a31780ff3a8a4b222b51
z27c6893beeee0ab392c41499c09f182e984bbeb01013536e5cc2aedf1226cd129a939746caa500
zd6db277f10a95f7e20bce3b0609ba8a085d856739b4ff20947d68739e24373a5d608e39043e808
zc9831323617dbd239c25b0a759164a4952186a9e3ace2e4e546dc5e9bc6ac7bc3ebed4b094e1d5
z9fc25406109163d877c88efa4003a248e37aa77c65cd05fe74a6dc7459c40806f007c01afe5a3a
zd3a89b87dd147f92d679a68f4a29484b19dc3b00a725ff81a9ba3762ce5f50d25cca33f9051e42
z5094c4957e046215faf0378122ac568dd1001fdbabec385a5ff222f4a3eac1e3640fe31608602c
z2a8cf40a9ab6bec1b157cef6884235af446239ce0cd5790bbb1fbc5e436bb17d6c901af48ab112
zdadab2e795fde79621e2c41ebe896686ea6680f555bd42875803f63abc9e9173fadc84e3510869
zf2b876f1d29cf6a719fe4ddd2a28028744489943ff5560633f29748412fa9e5e023b8451f9a983
z9c05baa31e389239a9f37b8ee79b72662e9ff5f275ceea0e4916132ed5d525a6ec6409a15d6d71
zec4970e0b9f7d4a1c610be7dbeafcf08747b4bcdce97ffa9a257589e1d23aa9568ce9d48196207
z05931090ed2e3c8edd64e71fb0543d19ca7f4004323065b55d148dce3969b5ca3e65bb0fc1b0a1
zcd07a5e29ca1898799a9484cb928808598316043b8c677940855489d0020c9d46ad986f598033d
z25d50a0c893727e78bf81d0676c0cbd8c742cc01a4f21453a58e4e4946dae934cb1f16d88dbc43
z6da5afbbd55bbcd8cd14210ad789a13ea57df34ce24eae01af1d3f35fbf01325bf3a8ef8448a2f
z0447bae2d7b8ef6f0065cce47fbe897292020b90e2f2a5ba97d81aa908efd63a327eff673800e5
z83ae7ae08c243a39881e1ecc259b6b56c989b51ca390edce8ef5622e46ef709198e040752f6f7a
z7a0db44469d28d1958e398fde28b58c04190bf53e95eacf86e9b1e36a3dc1a8b5230a938fc21fc
z960f34f0c235c85d6c2d5d550b1121669da601ace5db45f3a2e52432ab735eafb33aaf569c8274
zf66845b9ce65aadd113726089b2f67788ab54e481d76e2aaff9dd36d432e135ac578cd6eedf803
zee4dab379562793f286741c8df1832528de38d1ee992578796ba58ece1862ab01aa74435171651
z76a7c66a59827f2eb3656131f96a762d1f616451700bb92dd989d97fd23b8864f17761b2258662
z9933f9696cadf3d20a3413908bec25a2c0c2f3b738a883bf4a04df9737e1138334570bd397a94e
zf92e1adfc890195b8e7aa88ab98e160659dd323d698c09606f8b7879c7b28ae863df7767adb9c2
zee87887545b43c987a912f25f76c90a4a4e9e088f045c3ffaa92687f94d9310f6be617f21f39aa
z5f1479e82f8649df356c6c741562e9a7f62a1c814ed08e3a9cccc8d11346d3acb9d7d5a1e50b96
z472893266485bf65299b10d0d09e5cdf845671d69e5cf0100af7138bf199e727e984aa1fac99ec
z97dbb7ce06e913bd45e38b049c1fb500e6730cea722adedfb92116c15bcfc261a60fff6498be63
zd9c120b1d54641f653705a12646fde6e9362818e8de08614858d5cd52caeed8f9b967dec92141a
z49c0b4fda58b8b2dd13a129a707a541b3a198546e08f379f99fb8bf79b5307e3cf544a38f9da70
z276093726b5ea27ee38b96e9ada5a2200293fee7194b086a210b592e7460fc98aa3ef127a1aa7e
z6164489046c827884b001a6ea51d0c3fcbd97c1b0c7a461e2de68eb400a79f84a975833bb0c09a
zbdab4280395c0e6ee88064aab43734948d927e9b2e2b242518fd28e57202cfdaccfde46e3047f9
zf3896062d9201d12fa3bf750ba4cb4111df173ab555741e156200a8905569ca29cd717566a846a
zd3df4d646fa58b1054657e1696e4f22e4ab559e8be32ac4aff943ce390d9f85d2bc9a57b8e4520
ze832470333912b0ecabf52cb3fd0d2941bda7cba8132ca240636a9a856e8a312b5143c6c7fd2fe
z73dddab821a1b4a8d28bb505d0bedfb8f401840a0491c54b3510591e3d25bdff0addfe4e13565c
z8a36c457b6962d09507fb8e902cb6e6729e2496578e3231acc8295ebd978505b1e11e458d7d477
zdab746acd79886a1959d6462f6184e18b96edd10596485909f3d502c204580cf9961c9f617c063
z0cacef075de4e88de8596c7bcbfb152677b074093d281dc9d21916c9e8158f252e7ea242f61b8a
ze04eda7fe14586caafc2cfd98bbf3729ac24b1c8354f258408c5eac9386456e23544bd2c939a0a
ze4d5d395669433a6f3c45da185edc93174edc01cf5bb66872d6097554bb4b5c7cbecb76b999d13
z2beea3c71c1c2dd00e871fe3fe796fbec404983e2c524c68e80c9fbc6e5047310813582c9d25b8
za362fec41595baa54df279630114bd4907654bbc114c7c785c5a0dc3e01faccb75d1ccb7ee2b93
z593e8bb36ba5fde9bf867d1a4d9688c1d444a4f36cde51b47d0403d30bbe34eb23995f0412cdaa
z200a5c9ecfe182ed492393ad0373352144a5ad44e62c206262407899f3b675bab964143fe89e48
zbcaec8cdb5738691c74356748fdc24cda7f48c9721509d20983b7aea759d30b8b3880b1b539125
z7689b7c7b7ab5d04f97b563608a753467f09663f8291fb6d03da7b47408a3b573523c54e1be5d4
z97dcfecde3335997f83d77152b8efae92d0c0627d580b823928f619c0a0e5fcf23f9d3ba292baa
z2bf61fb155e0a957a380d1f6f7cbcee8e1f31743d09a944225e78a881ce6a93f65eedd6d1a79e3
zf3bdc206b37d4cb69bdac9e0314188b413eb285d03866ebde0e298d2f2d0ddb65009925870ac67
zd68e9752da0a719d741c200aee5fd164dbfd153594b43d8b473291a2201994587fefe2e1e2108b
z9d45d27a9132f99bd5f63b3d9e128b035765a87cb8d9178702b53ce9fa9227ce441352f97ecba1
zab8ffde3992311d2b5341d4b0f80237c1af927d3eb99a041f2e75aa80b8a78cbbb487b0f1412d8
z791c3b3c920d2acdaaedde25bbdc78539a005973d13048f50ee65f1ac8da1412cf2857eae2f3db
z0fae5fa386aa14c7ade286272e1c06ef688e735ec11bf0741b5fe927ec8304411ff7eb598106b6
z290086e9c1d8d244120bbd759cc965f4584445926c0fdbc0cefe90bade5f0d8ab6174215196f8c
ze8ff28bde7b2799377d0ba8289fb1beb879a50515d604263c5a3792ca3605afedbe72d13ba26eb
z50e871bf25acb989b10a5c4831b065cae61ef7a6d048421e408d29e4dbcfa4f40e515109908ad9
zc55510b49c5f9dd139336ef3e4ed89bca4df44b63869495e8b40e038eda886c7fd74118a1dd970
ze24c9331d8c2b98091fcfb01d9f3f085ee48daa565c6ec9ae991b0866f0b3053fb43e37979e1fb
z5d8d705da1f1e83d4b3ea1473a72f57c57713d039f41590f242b9da442c4355629830f7319b553
z79a4c44d4a67c3176982c92d7e074f88ae76ad34fcf0ef47d60e5adce36559df5df7b20148544a
z4af7ee00e23b8b3fa0f4e7cf8339c3bc949d3e68278ffbdf4c4f2c0698d13c35d9f07f3a672067
z6124a3c5cc4ac6155d4ef08f2f58649bedb098f00dc3d5b2ffe1a0812bd02b5ab3eb6930b24a7a
z43d506e07fe02efd5b462a180f97d3b945c35afd1644994605f80b412b3604dadbe6b8817af545
z70ae3505dde75599f2677484be4e3e4e8f57544d645e4746a1599eb27b4fba36b9d4e6cf7fef85
z81607a7063785e74c35d9292f1e12cab1fd0a2929c2cd8c35084f261f586a46ac4d642a41da24f
z9f81c8d8f66d4dfc7fbdfd345b4926ec1f08579ad78ae14bf0ac7ac752bce34628253700210e53
zeff4ed67c6f29f62f97c05b13270beb243bbdd320f88dc3fdc3d267138242ce17c6804761648b9
zca71fdefa059134b84cebbac14a9e86e14a34782356af26641162d5afb018caa56055fe7678cc8
z68172d2c1addfa930256e95ad1c8252aa846ebb0732e2de3ef7a9a1dbd4194165711932c2472a8
z010d13158308ea2535e9d4200d983a465fb1595d21c4fb935ef2cdb2625287285dd802ece348ce
zca3c35f95d1fa363b65131086408205f2374772e1ebf484c6766879e525a3e8208a42eaa3177ac
zfa22372151b28415fab7c2db304959709a06f602da6e6a21436e3aecfd45a44b0b84dff63acf03
z06e56220f7f514ab9b307e67934aeb0536068541e008eaa534d9be76f6a6519abaaf541b2a764b
zefb2a8e45bac88aa71a32e8eb30c1a0e046fd6b3ec1f424689c7f3e6f7281da34ed5def0e0671e
z462fd24afc39638dda608b67021e8ea4b359739dff86954039c02cea2e4774377fbd107df4dc86
za7907b910be9932fbd8f875383fcc684538e9c20e3d13f41707a0e39f7ed9bb2f181b414f423c9
z766aeb205d301668db0a0f2fc99a8dab222677b84fa14738962a002a08a0419c7b03039591a368
z0d00f17895c6ea8916c2df1d40d5c30c8f3d0d77bc82488bb05109a0e0f33d99f5995ff98e4264
z86939f35c4a4b2d43024eda89a124e3a96e5b17b7d68bcb39d40fe0a9f4dd268fdb1731579078f
zfcdeaa40757fb9eeb6bd2e30b0494fa770f6574166f22000eaec8c41c27aa23cba1307e2f6ffe4
zbdce6a5ff2ae0683456513fe846ef5165406cac4b6b212601e481330d208373a9db733440c60f1
z0af28bfc96aed144a70735b7c2fef8b0afd3788ee58828d70a7e0da787b07add07d22ecd9ed2dd
zceba5fa29a9d1c10fa9feeaa1226e4bcd5407ba7598499c944c90e4d0be9ad0df63682a1d5bbc2
zb20461604e2a7b82b6465ed02a2683540c5385b260b4deeec678246db3152578a693866f7f4d06
z1b66d9691002cee4074159001efecef19bf0b64a78ce2aee462bacddeb1bf5cbb722329f6f5697
z4865b0129bb2ecbe3417a0e446e193c95d0789c4a06ca89e01c43e000b4446938231adfa2b6830
z73d3c576cc168143cd7865d8eab156ac5443d2a76663eb00fc8aa8d10b1f5ec8cfb551ea8bb8a6
z9b949ae5a1933f3ba20f9dabf320d79992ab6f58ef3584d0ac2ecd142d8cd0c96f36658fd8ffad
z44441586219673b7570a2496b4a643064cc47455825e15f19053e8be5468a448b1c75e19c1e3c7
zcd628f154560d6dc277e0aeca0093480f07a1d4bf091b53f66cd1249cfee42879b1e1f285e3d7c
zf78a7bab5220f0cf5f32bb4b7d406c27eebffa8dad987274d28ed218003fcfb684257c9a2e808f
zaa76fca5a10eb573503d744f8c966231ed771e59b460f2c787069d59d69013341b32fcb4c346de
z6b6aaba2197f2fae8539d317064f26eb6ba828b3578c93b62adbbf5c2eb4cb776d29c0bb7ed22f
zeff4503d039f3cc92db4018604d9cbca2cfdab94bdc45fce816a8227228d859dd54c30cf02e525
z096948c0c50fab4ef94144beec4c44c0cf5a990f8e0cd360fb2cfac75b3f7ef9da3f8e83388a80
z21d0e5e47565b9073553c0f602d7edc921cd7c8f70ecea4d95f04b6aa7cf332a77f45ef8b05bbb
z015dbce75855d84c392b906153b9da3369467083f8268da39cab6e743b56e81abe77793c7dbaa2
z41e4c30940cac0ec7e0f32f5e73a3f98902d5d75ee710547ba5f5fca4b9e6306a6c0c40800e15c
z8f801818afeb498985bfab722cbe36c52f1f4dc3472786e6a6dacdcface1a5e3b73c1cec3c2c31
z736ab18a68eb618de3967ada911bbde829f6f946d5ada99c2a823bf4acdbe1acd23ddd87bc0ab0
za69e958c0d5732eacc91b1c7a7ec95ebd7c8e35f62370bd10bef28781de6ff0ff7d247a2152944
zc4c483974ee41daf065414f420275fb990c0201dc251056937bb8c6ac57a2390c09c4946b62fca
zf6c0ed64e9c452d86d59b760fb4f486142930e216e902fc1265f2f08033840f84aeef45e3a6a1f
z9b25076c785619a4f276059d352f1112fc674ff1980dd85ec772da2a2eacd35003c7fbe623e313
ze3c1f4cb1f82b3b5b7fedeef51a08490bb4577af47b2e87893029d1c74fda6606c1a0b404a9f50
zdacbcb6ac61b73e3d7cde4026aa70eafe5b472a6054647d8ceaa322fd6b8a44f178770e0eb74aa
z773b0db8acc17e5655daa403bdeddd43c8ab91741cfc19f2f337def03056e603a97e9173ab70f8
zc8b9b87223858bd5347dd8c8f63fe0f57694942b59fdc548b0fbe4dcf47f6543a589166f7fa961
za3d84f2eff664c2de7272c465a04cf9bfe8c065e63b83038c76248cf8607985fb9bcb264d6ef12
z39605e091f9d7203fdf1302b90522b67877d306dec3e491ba64f8ef6fbf18b4eefb60542c73c8b
z58d1547175be81fe3acc0add7d4702b5ddceeb5baba10ecbe58ab422fbe892f616446fee401b1b
z2325f0d5de1219c27a67de8729e24568f237319405208602054df31659fb9b58aa3e22e68a3f94
z751d5ee18d5260a411a1dfb312a38d50f182bb0b1fb8b5654a1c4a6066dac8a3811a7e8871b778
z11c743d4a005b077f85fbdd9f45662c7490cd2e76932f841026ec604a0ccbc987ab5f708a8cc51
z847b88e98e78a3676f957a956d9c9cea0620ca9b32623a0f72db61964dd8be95d280a6354a8abe
z2e58c5b1710559988ac72fd6c127ca8a77f5e8db9e0361e5525462d595dad250e773a8f9fa845c
z48f2939e2097a6505101c981402100cc888fb779504db9bcb753a26e975b76b848e90062a29fe9
z6a248af92180cd40872a83edc9bc0042460a6e5cb62bfa387bf98a69accafd37c18a552e24b559
z9382c9a6c02c7e49fdd8b2b3947396f075753b7ca2beeb22b2dc1ee7b2fc88b021dc9a38d7e6a5
z108dcfde1aa4b44456c0dc1b8c392e297215b5077281542d59147a496ae2145b98a1134f82d07a
z0e8206a0426fe99e76c2fae65e752e68880dec8dda6970fde77274cfabb839d2ba21b2ef7e1826
z2a2c5f0852703c938a4dda7901d930bcc173b26a15f706a4205e403816766e8eebe3077e8f4888
za506a54e2afa3d79d45c08b12d46701f01b9bd9515b264a8b6c8f646b7b0ab83fa32e2941402f9
zfe9cf6d81b6f45de9ebe2546290a5a120fd1b445ebf8f70b79face843999ef411249168a2a51f6
z440971c81ac653dfeae247702be63603bfeb397b9f6b8c18979af4df1310fed4fb145269a22dfe
z5726544b8eb210ad92d6b96de530eeddbe6c14ca1d4fb1e326d00f307794c88d862ab8c2f9e08e
z414554fd4fea4090bb47fce6778043c913d534406d88ee4d11c94e01fe0fd6b6992daad6bab06e
zc2ceb66694eaef719f8013d9f998eca15d98da9c880f46a4d02aa64013e8b3bd3528ac7aebf460
za9fbce464777e25ada341e0440106394556e2b6bb4d1c99f2b6771ba04beebea47445df644062d
z7549990b1a1bb0a044de8a12d7a66f886bbc4d1c589e6a2b9cc989683e599e1f67a3bffc71842e
z6f09f6848b99a33da131d9a8a1b295629798d4fa958b6bc771616f8b5b0bcf7c78f77a8349a18e
z1ac07e5a0dc68e1560f7646a9c9d3c6d09295c87a20cbc55c9a55881c79d12f6d1d1caeb8647fb
z7d284e68878eb624d93d50a7dc562153e3d2a772ce89402a33caa8956ad124c75dbbb05ded1c69
zb6ccf19a47cc18165b9dd5f9132f2a487250c1031662de6fe1b40503a9f768e0e63e7a23846c6a
zf063283d131f7db4a44bcff8a8e79bd8892e87d48a58ece39941acc8ff915933acc8db9bb6d000
z0685a42ea8084725b7d492d65937735055ca7c2491de2442728e0e3c9ce4d507ec69c0d5d0c9a1
zca428f9cc0fa1a76247d0924865ed02bc7504c7839464a20571b1803e75ae96e7d8dfbbd31058e
zfc6a3ee8c4be5d54737ea5a009607355346e4f1763c070f605d7e18993607e241c4ccd9401e9c6
z66617d702f390fdf4345cb2b5917571e45822526c10c0293417bd1aef9025dc9441f08cf5a9089
zabf5e263374512ad6909ae5715ee93755dd9db516ffeb784ed53dc78e3e2b2cddb54fa07a8aaf3
z7b249c31f60ec8da02026b5cf86091d6b8ffeaf4599f9c010c70284308df1c71063a36dd9a8913
z74aee16b1cf89f8aaa9c846193726dfdbc0ceaac0f563190f7abdb93575ec96c6401e1eb04962d
z3b937058741196b4f9b23466aa0e44ce001758a80179d39b3f67466a999084a165d2f598183ec3
zfb5aedcc4bc1eb8d4d2f40bf2c434d909a23317450551716ed5076f544ad0b7cdc5a971b691caf
ze592a04d7498b04dc53d29bac166044c1b66f3b8de91f1b349ba3e884e435c0208ad4a151da749
z0e0102ae2f64c9b2607f4f413aa1475516ac46070d81c9cd35c478b3946944f61a38a7b82f7f38
z4fed123f95f6523ed322074e1fda545e98119831367842483d561ccc5ec321a29b01026663b7af
zb02fa91371f54ecb5714c3f6bf1a4e136c9f698a43743166225ad3702c553983062ecd51be645e
zc86061176dbe99d31789382b2a2096deabb878e4acf72216006b0201890a6dd9391092edbe714e
z522c91b93a6f6ca45db69310c2a0814ba36cbbe044717201e6056c9551604be0c31f16f77d5735
z73257637cce6b7d3b3e5cd67355335ea8e6d7851722a2ee6ee76c2cd0090b09f17fca82040ef2d
z099d5ef0a07996bc9979d637934d8532f626932fa95dd2abfd6de666abc62634614be65bcffe6e
z3bd74a91a076610eb7436dd8ad339e1e79e80ca42395cb2a8a134fda8d3b993fd2b80d18a8604e
zd9dccf41a67f0e9411dfd424c2b107bb1acf81fa68bb60fc62b3be2d0d6c0923e172249062a7d2
za71bcec5a9bbfa04231dc4103d657ffc3ab33154ce7fdfec08e11be2bd4fd634cbdf039c7f547b
z52f3e96c06e38ce725d13b8a9b4c152345b11497a5c6b7c02a1ca078c92b320455fc055e06d8ec
zb89aba583a76bacb1960a35922294c4391d71931426626d131f3988cd73db50454afe1e42a7a59
z204858f9731a37bf98cbaed93cb5eb13c97f25c34667494d1d89e3a7abe2eecf358b34e38ad6dd
zb5840734361f6f7337eb660bc208398490677c67ce46bccfb61fc5023d0c05d9a73e472b684903
zb38b1fc0f2b56e8de08dc76e68a54a936ea5461d60745493427fa28e1d8e22931439cb3b2645cf
za68e5be2857d859e450297f72477d79d30e7e2ae3023a15ddfd3d4039bea7a085f26fe0e1f00f5
z2f64417f673d48cccda1c132dbcdbc562c92c04c4cb1b70dd2a9e025c235ec8bef760359bd4610
z34fe7072ef9d5b3ce0725eb26f251d78b2dcfe812bb93a0e7da0f2ed5896eef4fe7ce198196c72
z8eda84ac97552fba82e5e845b80221377a627c854d09ae4fb46235656a49cc28c9b0a104851fe8
z78b461cb74343ff992cc13873fee75fdf05a0ba334918a524f1d8b2d650aac86e1f80d0ba63fcb
z8a62193de33edf6c8e2cb7a917a983d254e239a605c89b882469dd62820f1d1a512d201601e563
z1d14cf7d98083249793a266ec52640ff9fd68ddf49c5db4753ef43b57e590af83812a8967e262c
z0c58fe873ef37ee431dda0af97b187acc5c98896bd235b60e39903f9aab5ae4909c9317cb426dc
z0dfa6eb6a9628a838753c10d54a8192be94963b5fac1bca6795ef30fd03eeb357316374bd7170a
z7a4ad03567ab2b4b1e615d9778cae6342ea87f3615f251cc7958c5f9648b79cc7ff7639f3105fd
z3200c8e6b8260533efe1f925aeacb3be99a8c4b723400fda07ef055bcf9ca5c93f843a9d4290b1
za33dffb0e4545c1686f22c0a66eca431935e94f8c88a10eea76a53723d40a4c89ef7b0214d0cd3
zc27f0e31dcd8534148b6e0bb280d29919d3203a4c8014418e96874c1c5ace299dbdd5090ded2ce
zb5904702c46e1e72cd14e7dba6768484d4f206f1511ae0bf143602758a440fbc12cf6b7ea4bbcd
zcf5a4d47bbe399664886464365a68949a815e124214a493bcc9c42ea9a5b0e63f78908222ff9ef
z16e2fa67661c5fa57f881b2eb30369085fbed478d6eb9109069a44ec02cbbfd235955d491bb485
z9a8159a74107c650a631361b5d52760a2bc09389c67640cca9126ad22875e6f251a403582528c5
z655ae15b0b8f921eaa225f4b19b903fbd95c5e4ee69853ffbe71a6ba5790cf282f2ef38dd98ca8
z7bce7ea722979f8a73a18e5f0ca7cad527d4669696efbbc91f9a9138ca88fcf82be141e4d59ee7
zbe03e051e31c68d62aafaa919f453b2ec668f9920381ab4116322c348a1638f3e53d8608f231f4
ze8baf1f55c5d7f72e476e0252294eded34906b52772d7118c8f257021e16adc2eb31822f5dc9d5
zb19541d7577b28346715f078c1cec247808e490e83f5854ab4ff897b9df89416b9bdc60332163d
z762bf326d5c1873fe5328d2988d0625ad41b809487c1dd1c37294a61de1b25c5f0bd445c837c01
z50b6225851fdd752ad809e03a6e2f8a1c06b170e8d6e38e341fd582b5e2b239e4df1ed89003be4
ze06b8d658ce59835b768bab5b3edb56b900f1f623350065a04129419797c378521051787535c45
z8caba9458a499b48c1ccd3966ebdf85b050ed0006c9b63d1883a9be167d9ab1bc29c158102bced
z5d62766787c4fdc45d758734cb07c5f38362adf3b46db2684e7dae7204362fc343a5aa77b8d112
zaf40f650cb7598b6681842f6a32f28ba4d4caf598a8b51271fa660d1e7b9e10bc1ad9a3dedcb5c
zf5ed37e7501a27c41cae630b1e51a7115a7d0152e0b6108e8c6ecd41716ffd91506cd9993c1fe9
za8f073815645a1cc84d7d6d96d6ca5babe2460b399d10b48ac1f9564d6c75e4e9f740cd1a9b44a
za23507081bfe2be6c795eb9fe944b6b52fa542911405d0da5603b7746b614cae57de0355fafcd6
z927b15d129d2935651b029373d26fdad0a1f97d381d44b003542a5ce8c5fb58d2d9bac88dbbb04
ze3b96d0c316add9dd5dd0b5cf3cf230d5047dc97a02d7803e1adec6b5c0737a5c47d40056f0e4b
zf9c024c1e02fffff48b112496656c6cc1e07d15c8d825d6a16a8b1c941598ea9b47f906a0e38c5
zbf6406bcea2d17065cb266f8a62cca1775f3143e4f74d50efbc0a1b8cc0b4a94fbb5a663924417
z8ffbbb76a9213049b2fff1ccb546765a0ca1eaf9b06ddb73138ff02349d4af08e50acb1b97fc9a
z10ed546db83d00c5d82f7e85005fc6727fd76ece529c29995d3a14376409368dd2e5e1e98d76a5
z0ab745b5731ba0d92ed93b94ef92e143ecaeb00c8fdee16d23f94d4327d4eaee634373f5282663
zc9d3f6d56c6a9ba4aaef0005130f5f3c3baedeffb1eddd870b2b4572b3d7455b54f6b0753ecba1
z1c653ce1311029bf04d420da738e5b4b767815ecdbb733e0ffacaaeb6cdc6233121dff7620d88d
z055ae4df607ba86182dc6d7a59b557e34b4c76538569849bb45cc0948b244c34161a9e6b7de487
zbb15b4d5c6153e4916ceed249d4f096bccba837ba5f304c3bc8ffe830ffc26302600d3858e70c1
z4200cd043c7ca693a7164f4340d90655fa3a18c47b83c2624e0022b34c3753f71a6df05bcae464
z7d97aba83a93521ebfb08ec954ec53b7108548d835d2d18d4fa27a6bc2bd8a269fc489bb9af0a5
zbb953330c6b2f5dc7a452ef8ea653650300e2a77f0c06c189d6f0f2460e8496b8bd839db5294a4
z9970e048bfdd0f38f2cea9b76f823ecd7a61db2694325c67bdcf6eeb1a86051556e674cc1d31c1
z6329347eccfadbf81f4b5140a9e3ff5a77c9d28fa05cf952a0f301cc976955fc478c9ff5ca3888
z33d3712d98f040ea17fd1e7ce7c43490bee52e3355cb64b667184482efca71a15e6dabbf2c2b9f
ze8f944cd20df0ae8df9ab7b29652c7824efde3081eac424ae243ab9d03603c209c894f73fb8c93
ze2bd29d038857b8ff4663c5eb35277c2bb0675ba56081145843b83ab2316bb8e746d70c061b73d
zf6a3d1cd90189cf3864759a266ad9084b36adab867a17d3f108d522c81302b4ca8389407d3876e
z09e22850f7c43be081e91c7ae8899ed1712f8689708715fed7f553cf579884c339d33ae4581a13
ze888700c058380e71d82c6de4c15708fed25c8972d503bcc8ec19a253888d7fbea9f7edef09a10
z094cd3f60eb329056862d7ae0ad33ea838503a72646d38a3e97c4215e448dcaafb383c59342d0d
ze74c8d6b1f9dbfcc17d442b6081132ccf08c8729dc356f7d40d234a9d4b1b7c3718c4be32ff674
zcaef2886e1d5069938c61da460ced52d9dbde9774b8c2b120f17b7952f6163f7ca1a52c999a6dd
zadb74747a2ce20e0f5c02982426c0b5d7d59599b9cc818ad3799bb3f7193e8baf49cf2403f8362
z4e60dbcffa9251cf06f04c056678a4130e9ef1753699473977ac372059cb40e5f684d4f16780f5
z113c77a2bd7bbc937baf3814e70f909930523bf5ddb4c0c58ffa7eb73507cd915852e7b4b80414
zac894bffb39f41e0c52fa024a97a233dc93d6bbc0f67ab3b2d79bb05e0c42a01eef6f20c788166
z1bb288e8dbbe32b95aae69b4466be636afc64b6e99671adc8ab1817da34e82771fc4190b70617c
z255d6edbff088adbde2e1ff520e647554378ef1c3f4544a71fdda89ff894f771baab0e1aa4d000
z36735cab09567ffb9ecbd7512a41899637df8d276e67d15485c9e3dce42a7a315df5c45de9395d
z282896c2d94ad8d518dfafc59320ef733eb0ecea070245e20ff89defbca51c39306be421ac86c2
z5a2ecd61a2937cdbff2d2c5e65e70376e1f5e1804d67d26b3c6c78e81c8161f86499d2b80d7491
zd41d6be4f18ef3658bf26a2182500ee536cddd49c93644fb174a7805362a86b7464fd7cf66adaa
z007998b14ad35ec8bd4dcaab348569bdc06ed9618f371fab731c009bc5a724edc68102ac3c4411
zfe645b8828235bf29f57155f6aa25dde079685c1de015f55f539762ea05efc07f0cf39917735c5
z6473a8be89eae7f1489741d38033d9f65a92c42a38e071d1a0d7cfa813c8b36ec5acb5f746b746
zec198ab1784320241c314e87ed2d4ca3fa4a34677cf0cb0a1cb0ba50981907f3faa3cd3f3edf6b
z6a7ef1f429df9cf99def6ac0be0b02127fbe367cb641ca6917d97b953fd27b96c487512be4d1d0
zb66016b168eb44a990c2e27081f5255432ffdc7d25c020742c82a2548feca92d0ecce8c0b9fa79
za60ec5de1348a7191440df2851368de08d1ba38e2460530faf0f7bdaafa0907b274d5f899abcb1
zd46d39e8722712503795f16684f5e514a5dccd9d6765a8cbb24e866e918bf63c0c53f605bedfad
z677c4705db18e5e151a56411707dd47f23df095a0123370b1a38e7674e13e71b117e3074a9750e
z1081f3154cff3fdb15fede3f50b815fbb76b630e5b6bd33be0976b41d8642387a2dbb14173d9f3
zc195a0efd9e3a824a88726733b8a1f8c717df0cfc781182a1d4632db6bb982b2c8cca506c619b8
z10bc3ca43d2b26cb3227be296c83a286aa50a5b650c5d93d974599bcd7036e9a1dbb195cb79ef9
zc4d3fdc1ee30430da8c9f73cd72a94677cb8c61168fd17728c75a31bfa9beea0ffb832859f0e5b
z3fa4df9d218d47287327ae20b2ba629cf8d9cd0ec2f460140b0fbef38b8b24693573e23900c614
z702468ce3e3c39dc948e9bebb755b46b1b604d058e1cffe9307d8d09af6a3e0954b0b4ba7cd846
z3480a1edaadd2a33c3740e9609b838cf6cdd0edefff1984f5f0b34e4fe8436e09d8a2a2849d9e3
z6d7b020184612547fe8a7f5712323820672b69aa072e85029fa7f5909eb0606e203cddfce6dfa3
z540946fe24f4a8d5ac88446cb75677f09aa4795a18031e6831eaaf5a2600951b69c0c3e3a46531
z98f19b2ba927f8d90a0cf25a4ed9c055d5091902c816de02ed961f9f22f6184a156933bee251c5
z3da35a8903a33540784a9376c6a249857a2fb3c55f038596264d325153e43695eddbbf6f9f6d98
z9597874e7ed12812fe7ec4e3a9e04e2333d8ff2f15277846628577069b04682a3cd255f84c0dfa
z593f716d0bcffe28d862c2c742c53e6eedfb24bbc3622e7dbe9edb734a5546f3b970b1e3074e58
zb1209fbfa61becba3caa04ed0661f11b4c94e8930273e02138a32070de8fa651c139465f6fad80
ze183486730b72add5362a06ceaf22434dedcf4456caf41e593ebf7da64780a6b407be18b609c67
z709c1ee55c7ca389f279ab3acb3e4ee50ffe07835d9218ff8c1e7d5772d816da43709e043a65fb
z65d5d3e9f3dbac8b5f141ea540fbf94725f52e4c9cb0704c184ec8ea07824e1cd838d1dcde058f
zdda3ca85b02d95181f56992c824dcaf16ca836e34b93081c8b31f33ab90c1c455fc4ad758a3b66
z38fea8cee7bf20aaceb97d1434b6db474a05867076324e0ce1fa5280da8a9f0e9f633057128dc6
z3b497b44de917f646958b2d72457cb33c5ba0c72a633294f5fc1878a8ca397d0cbb0c273c90da8
ze578a0c76505257f2b3655ae1379794329248eaf86cc2b6ae8cbaae309c7be1ecb0b897b5f8378
z38a3652930c20b7a9cc9788f67d8ed40a67e025ec4fc4955a60892b06661de425df94aa7624355
z3350daeb260ec087e678e949f83e6ff383177050def8490607de8dd1a57566b9c82a299595ffd9
z4fbeb753e3f8dd0c1a9ab5f654809b7fe953bff1ec7f834b6a9afd175f10a0b455891ed2f91462
zd382f648addb294d95ce0326ece8e6239f95df6d30c1734697481a33235f9f072a0808e41d2fa0
zb104dc7dfdf19d5a54278ff01f9c0d936baed7e59a37702e50d37b4ff763c152714ef9b7b6d2e9
z79012db27a93c1f9a908ad2974bf7ca0e84672b14d5e84e30f32ada95bc9226d7359391df93d85
z828b5a245f3d8c771b2a3f1e1783683d42716c30bad9e579dcbf95b2a18f6e19504d53b82c1077
z7739876d8569e28c26bf130d00eb0c75808f736a11287be235c684bcacdfe5f41bfcae06df2d65
z001ff0d76883d08c846186c66a92b832f162b107c90f86c183170d651aeb14c82b35ad9f7b2590
z7661e02b84e3cbae4e2e8bf029321d3f5b1c46baa9ab17e5a55be714ba6c52304168086ac129f4
zbbc3156bc49ba0f46a360d31df7f0e7098c078f529d15f597829b495d0f132359c9e97d2e08a9d
z1bd8913f7b66e3daa7ee53a6b1af2058dfd524d7499f7a1469788e4e081a0596e910eb9b8858ca
zd648968c1bd97e0fd89e97ae4f49d2c5e60f01e44766aa6dc2835665ec584f03e5037087d9dff7
z7cd18c992dee07b88b13a3d61d8a10c50f374d1519c63db5822e048342de209ed9f1149039b38c
ze09dbcd56643500ee66f30bc9d7534a156352d3fbb011a9afd4a116c8f03a0760be5310acdd067
z1be23619bc14a9f8bda59f5cfca5147017b9c4aa7de56a2e47a20b4213c673d826084644cf5ccb
zaaf500de0bb879677d9eac7163efc2571f3860c053cb00f3d4d7930ff14bad54181c151e72e2db
z1ba15ebf91391478d899af042f8875cb8e5918d2994983a264e3a403d9e6a9d3671a2cc4fb27c7
z881f8a05fbf9d0e2c7aa2466c3bac82a012a3202e352a4c5c96f560f7fabe5f213b35830d41176
z49dd53270f79bff93106e9c7980bdf5d63a4a82d2b90656976d70e48c789bc08f8268ff54b5dc1
zef8ba88ce4e9db85ea468468c67f13ca30e6c4e0f6eeb4b9cb91ca5c7d4c370cbdb894d228d1d3
z2fb9d20dea9b46f1c27b8fcaf923779eaa9d2c612d98f80257a31cc447711b876620eac2d1bcf3
z1d76248ef268dd29a1fa915465806a9d7e5c60f26ebb4475fb16eb5942b6566c37a87175bd3c8c
zc8ddb35fa3ddbb9a7a216c2733dff284bf52ee780c101e632aa0ff2d331aa63ce6a4c6795a95cc
z05ca1c775f27233bbaa2944d5c7d8e1eca84c89dfe05dad3a2f5a522553d187f9876e9213f97d9
z8a493e3055020a8da765db3562cc6022fb251a1c658e949a67516d8e3a0ba14bc725ba4f805df1
z8d57650329003d06a4b387c538811f3bffddb72a282f4e6805740dbf3ea189ffbabf13e0ef4753
ze1fffd6718eaf87b9f1e1c0230909ad128e7906a1dd3015681d082e22e7af85c41bed68449158a
z96da6ab5ebf6c0b727907d39080768f7eb6a7807110c99c50c0aa573e041bffd0a97b5528e593e
za5b2267d218a0b1d4b392210a9e609cea4254a800ef4f769743ace6a719ed6c04b7c2e0d8bd3ab
zc6734a3b238fefb8ec4becb3055a64f2ab77bdb8d6010821c9a3dbe43d17c714337d0e7b22eaf1
z320acf48d310da5a4af75349fefd2d4e2ffa868896e325313c3aee1538278df7d7449702745a72
zc917cbb07d1e01cdb6409c47246d8c35a7a283ff33298c7c5e3c9961fa94b5174d19f694d60148
z19cbcbca840928f8c8ec50615374d55caab1b58106cc1489b6ebbeb6d03b490557a9c1fc19d353
zde2f9084fb5e61ef0f18d943b39383ff864b0f4fbeb3f20ed47db541aa4c240e03bea550b18533
zf4d1add78baa5eb27cce698bb7c8ea05c2b900d7095a939009902a09321b5825ac2e89460ab9e4
z017232dfa1ff192fe22203b80e4b1683fa5dd0f5404f6590a88e0df949418c0cea26432f0bdf40
zb47959dbcc8d117e8db371752c99b60ed10d1db9090ee508adb59deb0968816cd948d2d3a1309e
z2b52032d948d77ba69090a3322404db89ce65aab9e2e87769a43e2b549f1af845825bd6caa57e1
zfa035229f0fc309b12baeb8fb843fa53865e31c8f786596057fba3db194e8d9b3fab50b0f527d7
z5177f1aab62a0c97c2d9b2ef5715843ced661c250c5a1630136ce1c0a33a6f65d74d4e7fea92cd
z011ec886f3e55ad742f94656edf4f8edb5eca1eddacb97ba068becdd5fbaecf8a19c54a9bc6ee8
zf2febe3f761c94afe5cca7255f48a6bda33e841db4724ef6a09b63d42a12c29570656aea533947
z3df110c243b9314a5f7e982e3a2c2db941fcee68c511a5ca8ad3282a30740bda1e8143f87dec78
za5aecd69b2bb161e1f6be39af957024961c81e45b4fe5c3ead4f9a6caa869625dcdd9b72da011d
z4ea93819b446e5a3e7c3487ad4483a11f5b1ce7e3a7fb4b8f14831bdf7e5ac611c180b22986b49
z1a6d9e1d4bf4514c22a0b72acc57bfc8d11656e54c066a10cfb5b6dc8fb2e1e44dc47a365a00d8
z5c97c17aa3f71996c67ae8ad6abffc81b27dec689393152d3ee92813705d996563e7ac9edd6b31
z5e9795e231246192a1a95c9ae463105b6954988e5231d814bc53fbb7d901afdc7f5f3609316817
z3546bfd7e839807d69c6ec533f93ad8288c06f14aa75e41b3358e52bf78b7f9f441893463ab07d
z46d726e9b57ee0de5aeec5f9841dbf27463a8c3072dbda083afd46b4e6a153ef816d39b2f1f7e7
z3ff381d042274b6f2f12741c09fe3ec48f8f85617f44169ae52606dba680e5969ff24fdc4e4149
z747dafd092533b4f99e6f014974f4e2d95a30cd789acd6e1e7fcb226553bf818a424504bea4088
z61d323895a0d68be29a8b374769f9bc98f09b578786c1b0d9a0788b66825e30e8f1c56c4d36e23
z5f3490e326dc37bc52cb1603f10cbfacdf5bc8b91d7416c60d2dc6ed28aed4b69039fcde17d3d6
z69521fc285a06acbeb4cc4f0f0b729d64df49c2d525045ab51fd26c656a9c5b5cef78da3a21f06
ze51fd3a459189b6871270f70781a8a122f29b698e9d86598603ceb602fd95060053bf1b114b483
za5697ce420305d7c8de872ad0e9a0a37fd1baa2e37cd6369fa642e09398d503092157147f11325
ze025b5bc22a78a046c7dbec6210d9194e837ea20d9f47700509f3ef68381913155ab22b8a798be
z611e1b7feb617022a1259853ea36bad495fe3971ff6bdfaf5e3a8cec6f5c294786defa2e066455
zbc02c2fae4a80ca1943f1be38686d75fb52d472cb7d7674940ffee25ad62d4407d12e96d9f54f9
z034930d3f87c2c222bcd46bc70b55d2ff677b3114b9704e46843c64aa18ba73d5dd0f3446b3489
zb468d950a2cf9bd32f0f5525d79e046fd4482d42d3f8eea33f4ad2baf033dbf3e20b4002c029f2
za01de27446abe43307b9e743adac90422e83e6ef9f5e5c6ad6a40e91027351efb8147c90e2c2bb
z49208aaacc6f290cd2bff96366bf973a94111d432989ed455659537108653cc5ab3f2839b1e5c0
z9ae4fcbbdf195dd6c752d191b297afc8dbefd99e8df81f2e78a30e3a4c63a3c4ad16282bab56c7
ze1ea62474adfc884de9acd46ad9e1df0704d29912a3574d57fc80fb316525825af9d11d9c25a74
z5b54f9c404ca79ac87f49f0521752b54ed374b927946ccd5ee58dc65b907004316982104658c31
z8618f4008e21e49d57f5d982cf5d29d8e052f6974a9efa0f2d4659a3a212fa35894821f74eb799
z0341b8f01f4e4475deb486d734bab66b4940e6cfc7d77980d1ea3e37c18d1d29e9199a5dfbe6e4
zfb0176df643a7003bff2b06d8f338761f96d005a5c02cbdf46f2a724be39108b770354f16f29bc
zf808f9f21eec09b1ec9bd5288e0fbddc152c9f1824487b2e4c5b0cf98ead1b094b5525b55a08ba
z1c3abc3eaffa07dc021cdcaa570edbdeff64f1edf5a3d265a6d53196296873347fdb3c998f54c5
z5940dfa90eaf108b71635e2965d47c33376b9d04ed16d03a3984f21aa1d39177fd68327682a8f4
za603d4cac480cd97fed53ff184caeb04a319ffca5277dff7f06d388254f0c5665da03c35d11282
z33dc88cb4eb98672f052aaf4cd0d85c7aa2168f0808f831cea07052b487f09733f22e0052f13f7
zd593921e49bc9c3037fb31fc60a279ca132fe0a60187d19c92fcd06dfccb71de0ceed417695396
za72107c9b01baa90a624a0e349b175009bc5ba7e287617660ec0295616d1e60c78d948bdac347b
ze6d45a21cd4f2f043b495283070c203b8d161daf6ebc52e4c7ebd0f00056a15a1320763391a0b5
z6d715f2993d1956f3eac857cee2eddcaa3fd3b9c0190572a65957099fde7c0abb87d31ca103c1c
z857005a24ea87fcdd4172d1d92ac9cba506d12e097e9d82ec328e9956d9b6649b3487e13582fcc
z15d86bd13c78c5b1aba1712e95a66fdff276b244b3eacea2e409f269c91ff3204b735e42e8e73a
z928090575c8ebf1d987d06027cfde4c501f0509ed64e163f3f2b71dbe4863a01a4c5e3d639fd1e
z0fe11a1b1ef3f8073139aa6ecbb570babf2098a2fade7ad80bd1959046b8b71e75c92586f22b8d
z203209e444f9017e553acc289dbf780342f0b1a64fc0cd3ebf1e3913311bf1d83700888b2f14a3
z35da0c91a4126575c15853b516416ff2e6b86e9e4680bd35a63fe419ce539e0eb820a49c97ddde
z01912cf85162259a6887ebe949b0a742c74df350a44ed95c2502cc83b4edc26f9f77fb0fe90c50
z552fb436b638b90c0cd8ffdfaeda9aea54e8763eaf5a63ef33e08bcbf3b7df27cc87b4c8cc9617
z0fd779329706fc4451d02331e257376c505f49523f0df26afe5386d5e70cfb319c61ab65c617ec
z4e9b0f95c9c15a61af3eea979a8d7f5ff162819989bbd3156dbb11257f0c00a85d8ceb99904422
z0c0c67d6c9b4a082410c35f316543b69575dc6e068451f0f5d593a59d825c960a4f71aa06c7ea6
zda02f2afec444d4974e2b739d916976eab9efb77ba60c6b77db0482302d6a9b8271c7f216b5013
z9689fd54c6974c0d6a1d0553579bb40ecad46ca2d8e963f138d4dfb96f36e5679e2df570d912bd
ze6896f2f9be15f62a3280d00a58a7648a6409ca349a9f0c8a8b4e8a863f14847c02bda1a77ae51
z0ec9a9eac5e363d7dbf31949e05a51b49c05bcc5f8941003d48403de3eb6f81f13228adb7dd9b7
zc1dd836930dd2c7d0e64e0e5d2482f254e23472beba34e53ed4eff1ec53d4626ff3a83fb767eb6
z2734d9ea0d6db22fe52cf3c31ecf4910a3327195b931fdba3708ec95c91e44266d65d293e6e4f8
z4394934e1074ff3d0b61e87854ac33ac91e998ab794f24f6ed75c847bbdfb42a68c9442080c792
zc186259e7c234903b15f032b88145c3ab85c6b9c12af05e612af1c803e4f00005c79de7f0224e2
zbd702e28da566a6b249693305d1b8cbfb6c2959e2c11985777b52cf4068cb187f24a1cac3acfb1
z1f019b81fd37247ced69c26647c2b39778a155c046193b7fdb6a7c73c65d89eec2417a1003386b
z6ee641ea20428bc0d962f363c666076af29b55efb5848634cb28b4da3e6952e569c2a7ab83bf91
zff566a532555859b008a2cd2369b670ec1246852f36664189b24fd53040005afb0c235a189abb0
z40f1c77826f340d5239280c36e40f9daaad27fcfb8fa003b437047beffdaa212ffee8c644a612e
zdea3eca700112a4f4fea4bc44844a1a5752bbb2b6b7669b4b0db599645556797f91b56e3cf78bb
z16cb4a17708e2e5ca2b3e7524fe897a17892c611621214b33a85a0211a73f15a85478d74e1310c
z4c45a218f40e935452cd6728977d0538cd785638b8c8ab11e9410b6f6d94e6e26e9ba9af71c6d4
z20c2011cdcebc8331a3339267aaf07608fbe484d90a570b724c0d21442a5b02dfb0a0d2a131a34
zee86afb603ec75bd2c132cf686ae1b8de9378a2de14ec8205ec432e959362f799007a136af7b95
z8c7f360dc8b0e448bb4333ccd4e7b7487d32f3d8b7b17df0d6c8b119f53cab0d4bcb0d1671ac7d
za30eec158f6a75db33f87e5551c14e8929295644d90129495054be7ad0070c5675435c7956d35b
zf7408afab2c5e799041a279504b6abf9ada82a65247443c6e78c50c71a182e4220b559e87de7aa
z7699d73118ec7e9de477478ffbabce541b766ba28728345cb1c158aedf666f2e265aa58c21e83a
z66d075b093cad1fc9bfc9d2395fd88583f353a142e9d09e37882d39c934dbf0770a9d29b3764bb
z1064d9109d68d02ca7027eeb728ba45874ddcb0ae3c655d98805e7fce07a4ecbf2c0c51922ce55
z37a14026dc7969f6c7bf78ac2cbe95d8ee4f63938c110527b9858d1515d877c532ebf88009ff8a
z2273f4301077394eea79caa82c0170056f1a68aa315b59cb8874f8335ceca8b96d6702c636b561
zc63a127cbd36f59e5a428e7d290c597fec34f09b1b4b7a75c8ba7d9814127655c553ed78bbfdb5
zc53663de436d273c6124b8f53324c3f73ed2149bdf1f1dc2ac57ee38246f4a6b3fb8e66a3680a2
z54dc487e2a3249fb79532b513cb2741948834cf38f5c54dc45c78decce0cd76dcddd5c738ec34e
z2cf62e2d25b12357771ffedd2ac1190addb9bb314cf2d3958c3f2cebb3fae6cfae48c29ddc2ca6
zed07507011035d814fe8f0990a983bdb16fe0daca76882d0324dd71b16d84453c648c004b38c81
z694e397a04f07921f4f6fc32b6d6669d0c3f0b696c5e1c5f0091704a728c5ecba7b2f2b01090e6
zb3aa7fd608692e0a9b94bc2275b30295cbf53e54686cdc14148cf70c8f43a5ac51fe3e1e2e7e95
z520196c80f47064ee244a0469e1ee0c45f8899a85bcf8fc8e1c9447126ce49360bb518f31ea72f
zcb19b0dcb17648ba822e4705131d9fcb937f0c18f64d4a5b84c4f48952228954d4f3dfb70b51e5
zd9352d2248b993b7c5295cd8b9b16bb4f0bc2145a958867a8ae29fe95f7b8ed9697137981554e8
z1d88f7703152d6ef76701c7c8ddee11a13691e55b88d223fb1a35e7bfa28cc7398c5f685f3b59d
ze31aa9c18fcfa2424bd5fd2db84302c0c2c40f7ef51f310651c86b063678a41fef614fe777d711
z4aa81cec8ab8bab9f73bbe7e462f47ccc784832e3266b00291a51b381f45438f734561703e883b
zaaa152cd0c39425e3baf5fbcf00a333573e0d61cc3f1f2a21ac3b0041a35b8e561121dd5f84769
z7e6c408e855cfaad18e1a62f1ec50712d18f4378a6e1d606c8ff0e020f86bf95cd9f22945b7804
ze9e46bb2ba103f9592a601760c61769691cf63be2a781393ed9db49e35b310eaf730a1f086f771
z780cb25330d5001089f428e6ae5c6ec1e342cd886b3ebc4dcc0da7730dce520f190bf5e6aa5024
z22d2c19e751bd1c33389384c73ecd7876925f45691b0c49cb66cbc9e4430720dd659a675899974
z5f874990ecc96a96d1a133b488b057b29e2af8128a0787e685484ba4d1707f6d3dad18466a962d
zfc8e0fa30d7b027857cbca80f7532c2ec3476f7761f7fc61f92052420d15929a8e53c4a1639fa3
z7730bbac245a2b360926403e58c71f2def6516caf63d1da8f53a1f99ecdd74a05c047009a704d1
zd647e4356f81c0ef15c544e8aa7ed918158f2f196d5bbe0581517932118de65f8c4fc9221c2b34
zdf3026fb745306e8357918a1fd4aac865e2c73aea0a74f9751092472a2bf98eb2ee0cc2f6b09ea
ze8456e39f19eceac5f77113ea4fc0fae0511a80965a9e8c3a39b9843d5621acf99d5fb3ea3e56e
zca890cb10bc0987bd9c05a743831f1895a68fc29c397cc37fbd7c7bb33682d2f504cb03bc4f93a
zc6156827e98db978c1ab2592b8cb97dc457abb456d3c80efc467325f2ae0ebaa750b802dedecaf
zb73c47f02311e4a8242ae18dcc2e41ff6c7b7691ec2d4c17b50afe90210f48898c823efcdb0779
zdb55ea9789f6d5ff3f8f3844868b0a0bff2ea39907cc5bb152e3d46c53eaf8360b0b2a1f8f7a4c
z2dd2a63de1b8c16d2619036b678cadc6c5a71ffddbc47c2cdc51838efe60b1eca3b48cb916e49c
zb8d4731da1c8710af37795f9e9ec2c4088d8d0ece80d50468f017a20e8d2bb0e7568c2f9485d00
z7c0e1575bb1274c9bd2d61cc0999e7ca665bfa317709cf97c0909e6b669b8b9e7df0504fab3c46
z9ff4dd2493841111d32d53dd01c688f6e5efa72237e279c788f7522f7fa87de078008bd8e74681
z67a0783eb6ced0c49efda616f75b3aee7703ea3d848f64dacd58e62e3a54f12ebf476cec68e75f
z59a0eb14548f0b125cb1d922019e4f82866db8111ae74a8637deda4bb3cabdaf9e855ea22bb811
zc5bb816b01cd5e01ab48cf01c6071363950ad944b497cd4dea0729e3bb93141c9e84b6d1e63431
z9b3b16b3642c9f9bdd20f205eb8743c60e4953f1213b13dbf32d4ed67f681eec3ed8d5fdbaa12b
zb48f779d186432194de1399d44c417a44bd5d9ae44fc00d27c4ea736f82bccc362b3840129a2e1
zc3a38926bb9f599befc8e4c6d9ba36e4d2b29a1e635063c3b538838a0b6b7c7682a02c5e32ea8e
zce24ad5d3c30544f6e7a72b66a3702dbc513009f919c365d9dff0b2076d2faaa079312e3aaf51d
z95729ee9512675b2bef03f61f42affbdcf9817973f5eed5fc5decccc293b4af27b6738259d4e1f
z5b94bec8d1fb96ea7bba32be13fdf358bb75e7dfb3ed3f2c3594af9a5d52f1c53517913bbd5fa7
zcc268cab072ff08813d2d99691041642027c8c1a97da93a12bb6c7db3e3549ad759188129959c3
z5ff1b10f4840476a0999a3d9731b7cbda7b51f7ec183f1808202853241c737a034722b688617b0
z596b4a675920c9f00e13da4445c17ebe244118eae583ed13af455665ffc8abf6062c53d40194b2
z7e1022bbc77d075ef2197fb8e6c839301bd39f218ce24625db8918680a602ef8cb1771a0eed109
z566e11bdbd541da56716a0c719e806229e7421b95009b2d9d35d72bae81cfa6385e5bf69e2e4f7
zc71d76885b27ffb7386d85b680ff11a6f267cc8e7626d524a5e685dc5eaa379f059af0026a640a
z9dc80d3f87287f6b24daa0e2a5b0ed460b8a1f742b57d8ba4e3af92ebd73f893d8f0c06552fbfa
zf147d8d3f6630f563883dada876ad3a0923c2cf2451cb077577921becf937530dcf5da93000455
ze07a31cefb3e903f9fd5851dc45b9238a2b73e6ce2af8e19aad51a7fc32631cae550dc159b04b3
z903a1b55c2ae982e6b31a16da7901afe9d218a19cd8b1c13a3d453f09f72b8134326bdd5772799
za27348e3171d745a06bdd6f23b5c6e127e96f0e3ff72f9a9d862263e34ed15f4196dde769d9386
z1376a710a82e6cc05d71fb9e5ee0374a239ac486db2d8806be5ce685e9864460401a61f35234ab
z24a58df9c6b53259548a9d857832aeb2e1644864ec9e92213b3532437fec780f27bfa13969ee38
z8830b76d524c941db3cee159c93176d361986c3f10c87bc6363b9a52e8ea54a561c62aa17d6319
z7f6986a3015f4f323cc7829fcd3e109cd270aae167542b6d28e5d938d660b6db31fe747b06a16d
z4f7b111b7acbc749f3ca875760a8f18476cb8bc3b79e54e2f08fca70ac7f039487377a3ba46e22
z4ff0b849f9726dab4647c71e3f41bf9fdece2f57c13054b7752cf51ecd42c17b66a14facef6054
z8a4f7b4c9652e4d5eb489a5486f0809aab330807edc3493c4ef4545d967286919bb50fbf368fd4
zadd0946e9475f532b42d810c8211698713b9c908919da8bfb47d9e1d279b67159e0a4fa748eb76
z6728ea47cdbf30ff1f10bd689fc50566e54aea40e65f0dbc656554bdaeb2147b8d5cc82c42e948
z6d1326afe87fb56b880b4aa26cd05d652192d21071e3aedc7237858492c5aa860ca1f2418ebfa2
za811bf9babc6f66722efc42b3621bcf0a19c6707c4a7d485fe657c73a30c40090919325ac18826
za22a3feb0cfe81dc0f95a3cb3fb5870a34360e4ded818206de4fee82ab2dcbace2b0efd80b760b
z765461bdbfedddd53ac27faf7c9b1ce63d5e5ace622e219884847b45166771fba971808d4cbe45
z4fcfede5ae47abcb54fee1d1466ebc594f8d1a427ddde443e6aafce4920aab9dd7fd64703297e1
z8cce171f7f12d78a70f4f11a0aa3603c58a4ad35d3c8170595e0b56bb700fbca4d71ef8e026924
zc61488f3ce5f50b45d7ee6233a4b720f13681dc97c6d2e6ed0466a3c779f0ed7a20ed4863cfc9d
z276a7c97aa6a9964637bc436372208eebfb42d061da2df1cd8caa82d41d0fd05ac63d7dab3b9b7
z95fc6469ed398de4aff965ce99a27b6a4e5232e00840309ca1b1f80b7502930eb2890f8bc33787
zc4fd0c9b496a41a34e8d5464e502ad2f5056d2b14cb9b35867191dd3b707a5bfa82575678014f0
z32cc5c401cbaca45f68c097fe4023c98fae22303d0ece7b82fcef8042ff8ac789b7803fda44045
z3823c0f3c0667e9292564c8779cb9a4e523e726fb46651ea6e97a0700658f2c878098fb246f94d
zbd9445ae3a5764c72e217562e2cc499832520587b3dd245d1a16aa0c160a713f3fb7192d6214de
zc7d9df1749c058dfee557db2569b114d08098e4f8eb108ab5980e7960bd5985ac7429760f8981c
z6dc082c80703eb2536b2037a1130e17f3858e38f2ea287ec8b02807109ba66f17eda01115104f0
zcbb741f7213ffc06416fc65609b6a1de92f25814d06c85cc0486d499175de45d444e0f65e1c186
za847dad05aa9860f6b3b95ba12455ef16f59f1964f99ee9bfb30e3b46b8e8f5f33c7a63ef35555
z9f70c1882010e050d1bdb65256c319d22af3eb6b118be44685d617b4b8205f547590138bab01c3
zc97617a68f186ebc31e4e859de5e762bab454dd58a99e3c156b164267f13e09bb7c307fdddcb1e
zb1a842cfcd576ede22459700e0b23a3a9fba97189e70f76c74718463b4b2b8ee848c318384b6aa
z85de47c8ce8275f1a9ecc400fac37d7d8fbeea45a50352a798f9586b94daad0f5760060f480870
z2e9784f27bded79888d183853f964a022bb8c23968d411cb13661bd41686e7f4a871eb72812bdb
z0c86ad9436ae672f925b37ecf9a36d3f4013945fd2170dc0a046971937300897da35c7d3684322
z6f53dda96b48d984779f067cd19f5a2f7f78afff851831a9c16eb52e3571208e65b677b51b3138
zc3048c09629964f603fe4bdd7994c0448d06f4358576b5b9e8e238a385afc5edd4fdea1323cd30
zcf8081b25cbb3c6b43cc1741da809c99f3cf1b2cb2b2c6e569a6445e831444d28fee9a5d540bcd
zebb4d54c701cebd7b652c2415512a8032efe26e241571f397aa26d407ff5ef0a98a53c350539f2
zdd3d937a8e4935d11539a842751ff1a12e398ef9aa2325d3c6c48126983db8a2af4c2dd8eff280
z48c2083602f25d5b599ea6e54f107fd79442a632d4b1f6937f4021f48171bd3968b2212751ede5
z164303723c40be1535050ad9d623e21216aa4cb2e144076ff2effd99784d0bf8822ac74623af0a
zd3f8f74e5994d6a2a768ac294908b0a48a4b9f17123489ad2ab3e96aaf30e19a86e7413ba18ca2
z8da7a001e6439d557bdf8e59b6d04cd59d5430b4597b3d775f9e84978074841af4682f469b209a
zf2196ac7b43d2df8eb13a36c27464a9e18e925bd76484888b551e2b11783cfaee32ba93e729590
z2ceefc76afb3fbf29276e0b0cbbc3e33ec9459bc78efc81b76877da5db0a50259768b3d40a8b90
za46bc832e16e47e14aea4530395eb86f9d6b1ad034a946fabd6f472c4fb5ade4f624beb2f6289a
ze15f40b422f78ab237caaa30ba233ebdc3b7372c2c49694f0080ab19c99bb94dae47592e25b43a
ze82c3996fb375c2a08b4d93e6c4903c8103a6c5674be49f74c437778eb9c9a4586aa06e15d1247
z644ac3f803e7c2358d9331386fd9283c65ee8bc66f569a80a1733fa73fdef468168c40899d8133
z8b48d55723f429fec593e401df35a9835f55bc4411b2839e1e68bbea0e40225a985a27a51a31cf
zb791527c9a0d681a232c33903637feda94d9d9fccf010aef13d28d1305372683bd7ca512f46357
zeef2bccb14fdc6faff30bec483710bbc74955888a27b3389fbde301c26c3347c0ac353e133220e
z5d1ace48aa64268ccc7bc1257c3733693d3f289d5e59c63360ee1c73f463ff394b32a4934fb8a8
z9eaeb4bed614472c3943cb65af5472bc88bcb6fe0fc1642d9ecfea707d86cddaf38d0360751bd8
z2d236e8ab07a1697d354615e83bc54e2010f455855619734425293efe08ac13d3a18cde4b16947
z5949e6ad1ef253c8b2caeb6fca22c946e890ef84e6293b010188125197148df8665d5ec3502fd8
z32716f668c0ed1b9864d073e8c84c30f4093512dedcc521a383863e2aaeec70ffd1fd645f9aa3e
ze6c8ba9f2b634c79b47f684eddfa6b6843323ec48c5e1071e145a52669cd819e6a8b33d4592c12
zc8f5704ae40728e2506b02d73004f160ecd6c34b93c6195be5d4e73d492809bcc10ff9a8c69cbb
z232876371116cc3bc1c2e4abdfd858c45fb5dd52b3f749331b744babb41499c15ae1e2e8102b02
z5e0b60da1abd7936aec22e9e33fcbdd1f9ee398c587e3ae251dfd072c45c8b51d7aa1929c76c5d
z4706fd8016eb502e816b8cab6ca63bc62dba2e56843ada1e276707c73af8ed5e3f59add660a774
z9f92b3403b9870afed2b919f89c670ea164017cb50610494228afd8d019f5af25a928f3573a1b0
z5536f2a22203338d9b5c4e03618c09cd27785d905aebc4491abad62062e709256a0d643db4318b
z40f4b8aeb1b5c44262e3f6ed5f079e22e4eb195d2b2c2471125e8989cddef0e1901d94efef0738
za3f423c73cbf25870482d348027d55f7f9cf2b3949761253ffb8bb5a1c978bb3dea5f1d9a8b1df
zcbc7d1579346d951d594ac0d039d20944598b333421389f733eaa95697987b81c8a42c5aa960b3
z0796cfdb226eaea5dfb3b5fa10514cbdd996daa10c822c807464dff568c3d14bdc3a5b91c1e8f5
z02c210f66fabbf8ab0e6b316e7f9e95f6eb1e3792ef12be273b6efe8e4a9e221d13ec4cb5ce307
z7560486cefdd3e74e39ab4418ab2f2f7797e23792d6d63e83cabe4e4882064142ca19a07515d38
z750a353541585c58c244a82facf7c0d09a32a7f204bc6aba62c9421fee906b6d03092919cd7098
z3179e886c2651bc7b6017f18c7f1da2d5418600a6e10e4fa95a1a127c8baf79a6d24d857269133
z84400758d40925ed857e42f74d3e6c9c417e7d895753047895b904d8ed631c0cd4df7d4b57e2f7
zc5efbf97c863076f8adf135ac7ce6134d75e80aedfb5714fb8156a93493db0fc784c0d2bc01d40
zc51d9f9dffc30159243d73778c46b39acf975bbd2af5655f9feeffe8d2dedd5595215c5831cff6
ze72b0b30c68f4c9cca762c7b127791a81d6af15b9edb351d500eff3bc080c855548d9019d78b80
za3750d4b401a9883a50dfd586806ac15b5cda133b952f3808da5c0e7c7e635ded3ff30a5b3eda6
z00d737bc1e7cc2295d3f3b5f402e0772333924e59114c60b081c8963cdf90972bbbf2d4abe0dfc
z6d8c343a25e7024b4e046d7a71ac8e6f004a5febebe8b302b206e127ee4b699a8f082fef6fd7a7
z5508f62b1cec331bc03454afa89b2177ea5a0ec807190caa2de56ba6a9ea3751cef14661828533
z99e2d04eca31257eaece886277045e13a0b934c79c1201e353e324fd56f229580b30bf50147792
z2d467d1227666a938fb91735a830700e93cb0d3700bd0efb44550e9b39f303428a933f911815d8
zb6d5c92e68f3ce4d95f6ca1b4c9313d4acb02b05abf742691f7abf452a281fd682ba2716680253
zb95d6f30e98405290a72552e52ebdefd720345e77625c7897e7aaa1f885eada7660f558c048908
zf0ddfc2266b01db1e581ad4daa7cf9dad87a876b6e398a976feae26afa918fc94b066471fc512d
zd6ca06fb7910db7cde59cd1ea4ab8b8dd707fe078a0d9038a13de3b1ae6b799f6f35277357d923
z3afde4b3a92b61fd0bdd61b99b0d9e44eeca9daaa7d0cdffcda058294c46a9827b19e1dcca94ae
z167d818c9a91ca09b30592953ec69dc4e1c6b2b26e0ecf0766be790c8e5875120ede81e16638f3
z8497ed8f2b570b7b569ebee558be7397e5acea7b20efe1bb48708f71245519698da765a6b81c98
zf5aea135aa6752785018bde72312588200416d0c3d60a328ab10d6722175723939021dd7fa3d35
za00dd7df19c3c98b26438caa5823192187b31307070f401db12d83dfc3a596a493a11755785c08
zb3eeaf7745679c0e3a6d7ebcdf3c9c57f37f1874514e2d3d503b7e8867789608cc130bfe901f60
z93e8e2d266bc5945dcb27654ed5e0f842888aeed15d8c3f84cb98a74595aa47e65f7a115af9e59
za2fbba23871f1cff4c833ed52b14dee09fe9ed1633a9792410fa4b0feb7d91f901578e4d9781d4
z087c80003f48a2ceecd36baa3d4ac0eccc60f4a52dcf8c71770b36b9ab21b3e6077e426a5efdfa
z2cdfb0a593e31808da648219eae1c34ed82758887a331b767671686f4da54df7413f65516c36d1
z6ee64ebf6ead034e325b9649697abc4eb0660469de073a2a294f416bade38e503b6038c76df9ee
z1747c76f0a846c95615c767439d9cd77d0558c206a30763d362296fe97c0bcd3ab89868f9528e3
zb456e841164006a4e4248c1ce3c2a29b9086d9dc0842caa16a263d8065642598d990873599b178
zbf57c9625d38d1367e3cd513c334975bc070539a48d52fb54c5a2a23908665fff3591ab6959372
z87ff70fcc57835d1666170328c8ddb6ec6ec91a40ccdf6cf8a0dd634bb8da43f43558b4b94cccd
z1036cc3f4ab75ee0afcd2f890882528c783b9ddd97f626e54227939869dd6ce902cd6bf4770c7a
zd8923dca8cb930fe530ea2f339eeaebc60dafcc988c36c93aebb9e686373333e10ed779a6c957a
zb298cc793bebda0d3af98e8782d8058803d3827cf5c8846bd92638ab9d950f9ebf22573e275b8d
z3da3db92d3a795378c00ffd675dae7d329d9009c9630e01668e9c8221984f3d8826adef06ef87e
z9ff909593c5364e820b284ee8999fe177571ec48be906f9ea21a6de0ecc09400a026ed128505d1
zca01a8f7f33825167e22f0cc0301c4a23c51801e7bef22bcd9be77414e757ca1d5b495b9e87eb8
z41927ef532272c1372e2677deb34f99f0376a51b60cb57d8f8283bfdc0900f11fec454b65f2b47
zef68b0e36210f5c4d0f40762dbfa0dfc918965edfc449d5255d05fd95d2ec976f5452d9cf05157
z9edf68b5102d881ec46403d54baf38dac48de284aac7bc96ccfad0c11921626b18bad439810cd0
z4516f34cfcec095b89fce89c02dcdd92ec2b0fef3a7bfd00d35dca549b2f9c7ba293f7c54f104a
zad6f2f9ede10b17cc10e3126397da66eddf92c7e91a124aa1ce2e15bcb354529c9b3288d1af931
z27cdeef02f4233e6c512a2b29e4db23fdfe75b9c279f32e3c89e8284b7fe11b7e8938d9538bbe7
zfd5c051fa587ca1ea7d6482e80b4ad77189228f27a31422d3a5f0dc2b570657e90c20c9c3f5510
zaa7c0ec0d44e2b8d00893ff03f672ab6d7bf07deb493f2c038ff95f954b3e7b7b3a24628085e47
z12be12c5fcd173238b732d176cba74dd7359363dea261202975ee1220ed70d2e0aa87a930d7d98
z61a6a9b957bcb912a19cc97817c07d3a60cc75a5a6a978f142d4b1a4b13073eab0772038eddf0c
za7b517a73b410f67f6fec7029a55a934810d8bce4d4f4fd7f9285a080231c9e473285698be2d88
zd9e6efa56013cc8c1ef3db112f7db9daa5691e8c7f6bb82d4ac89c34da8e2267c3231b4f0919a5
z0622c8865701741e871580e17890a1f998b1db703f4c122a14e47bad7252eeace5da4d71940009
zf2c9dca0c89c6c6cc7af81cc4715f4b0897591d9ccd91fe24575a150f4b1b9aa55963396049764
zb32cad92eb5346112d88fcc7ffd328594d22309138803c06850b6da1dfcde9373ddea002a24a95
z216985127e982bfb3ec559d90335b5b7761c4a2dc020019f4e2ee4f46ba8627804f3d7c561e47b
z1c329270da890d5a22ffb030e8b36c08ea007a7167e3914973955f4e794e80dcbd22db3f035100
zc8a8efa0268911a42d564b62a9ec3012f4ea99968dba376749f06282061d7ab738b5fecf61ea19
z85701a6ecccc7f304eea9ffecd7cd38aeb31bff3eaa38f9a5b8660442099c61ede8913f854259b
z7cd2f5ca5a5835513ef4edf868c4b1e15e63a8b38429be310dcbe1068a2e1a98d925550062e6aa
z2369b43a1d0f8fc293e848f5e1f22ab8f3a19e9447a5f776e79d39b425383111d69ba907cc6fa3
z4caf60530d55738da11794213225d6bccafa48240067a4db53ac31c2e73f2267280822606d489e
z0fa7975270424dff73be500ae554b19f6358f424cbaf389b2f8c54b554b459ba1a4bc41db70177
z73ff92b1a71a07a61317e3067cdf6e634352afbe884cd888a5230a36722b210392d49178c0f7f7
z577157a00fde89b3e29b382629394fecab9adf414eaf8573ddafa50f379a0ad0576e952d5fc1c0
zd36549f6671031c2e02c0a10a5426cbca6de30fb7841328ba864ebbf044e99cb6098c99033a7cf
zf3b0cb3c3f6cd98d7e21cd98d0e31b96251d73cc8c19d8950fa36182e7ab3165d91e3751a3b9b4
z450b04b23027f3ed8e11c55324ab00d991b0b19b00584f6b1854ebfc0dee9d517c709fbe4ff313
z62b0c4845ea8d5fe59f83ab508eb8bf9d5050384ba46de16f3f4e51a9be507b76286c15786d989
zb4c03961f86c388148dd9954941014a6675aa5d9bcb0e5608290b839548e384f6dbd6caed83071
zfb862dbd916d497cd6711c8659e36adb0f4b8dfad690ff96fa64f6f88f86e7e5d78442f054a170
z1a3aab7599c1ddbb70a4dd8eb7819ab027a5fee50ef4df3637c80c93a1d01f6e19f74900b5c927
ze22fe1e9cd69590b263d5a4071119bd8f2908a59289796d3649ce136684c5eb2ca0ab4af3b974c
z1d40efc781ee9d528df39bffe63f892e9f088eb3e3fc8fbd7455dc7a3a5ffac47228113b917d2b
zeb898e6f74a885e10bf2cc9a5d952279f03e4abd22faab15e0546ef99f910e3f1df38fbdcb88db
z48555f4c3d9245aec14d3ac1939580f196f82d90bde365af6357e134b871fc9744540ed5e6a1da
za7f05fbfc68e64c8d1759bb8202ed90a068b205d2fc21db346e0912df819587d829e5524dd033a
z0fffc91abef526f689c7f7be596a45f021c14ee639153f90f6951d50495559235537ef80363ea0
z91f88fababdb6587518f03d8be251d1dfe1f664e0a8a785d045f4f36af2f325c7b89fedccd65ad
zb57e1be2eda5ad6909cc9521b249e7449654f06142753467d6f92a9ea619d9fe5ff8510e187749
z920baa383cb1cb645039d4d7135ba028301610bd06551d495f1a8f73be0bad6ce96da75a2aeae4
z2548977065a1c6d091cce6a9b3ebe78e4ac3bac64680e64a2e201c4663ad3f22382e51048931cc
zaa95c96fa62108c8d6d7f7c3d143af11d9854e32a8a602ab0b88e9e45cb8d0976b12516731716f
z676e8c469793888212005c7ecb2580e5fa81f954ff3976cf47b387992bd2dee350698bda20ccb6
zb9f4df0cf44f111d09706af73e19647e786c0abc6879707f7918ceac493536eb9f50785b9c293c
zee1dc3762a5eafdacd181ef47079375b07c5a40c194f4fd967415f55eaf80faf8a9cf4efc1a543
z2c7341093d8c3ac8903e3efd0ecbc0e4b230c111576c3de55c196986029ef24615554098f241d8
z73c17175aca725b0e30582f5066d1c8ed10ab26274588dc5f5e4510a2be5fc299b1aaa80c2209f
z8a40477d697b16ec72b41ebb39fdef2380990139c6711505a3554c7b775b7c7d1818ab5805c62f
z52fbcda450e9bd0103b71a1401643e516aac33af4b81034d3cd4685abff9f693c3055420f1015d
zb1ea542d808c0356c18fd324fc5f7e9f281b72c076c6ab4c9c15cc450e14a4b2b9e0cbe1b41113
z4702a8154225193a9187ed09d7d9f4c52d6b78335278a23c9c7848cd33a841e56f9eba62d6d80b
zd99470cd5dfcf903555acee46f1a18cd1180e8221a1f75dc46cb997ab72391021e20417335ea1c
z902145c1600556ea73af5a74d62397fe3c07f47e7fc3f0595d8d952c3885c6e1cc485d9f623e9d
z168d664699a54713ed4912ca1600351b32f9e2a7b6704f8eb9b7108f587d5efbe12d8ab025f1e6
zbfa8f995c9d1eca57e2051031fa7e7da428956ab98bbafbf3eca9df64ac6752c580c3bcae36b3c
z50e0301654c49ad45f69d352e4785786591041fe32caa42cbc4098af3d742eddd74bb581436a5c
za1a686473aab30d9c872e1eaa778b3053c1c05135a478699f8a71cd33b38436289b1ab1f44bdf5
z399c30a4b10e4c3006fc449ae318db163646426d61fd471f46c5bd09b5562272c93fc35e0497af
z22ccee4bf1ff6822f957f01ab5f6698474003132e99cdc0ba38ff8c0235e3251655fe93e070f8b
z564017421714a756b9e27387f135f6e801fafcf50415ac629aaa658005f86445aad6af5bf3f60f
zd6579197807a9eef6b3ef2654a992deb8776a5013bc50f0d918802244325053b11a2e5c4d3e703
zf17632f6e754d7f314369ac3bb07a5b1f326dbd2a3171e46d9e4e4a058db6843e6e4f4eff07fec
z546bdf1da06cef58ca3a204a1ea2e52da06c0e97eeb09bbde517c04ed8815d37703a462d7e2baa
zf09d4d1e2fc1a3ca1941a2baa42149e0bfe045903cea180ab5c57d14ec0bfbb252a831a97743ce
z422e5eec8f9c3cfe9f07108147a61a2893757b9873a8819aa80018d97ac6153d9132657f43a742
zf6828895c98ebef08914e9ce69e6a50512304cd7ddb1d40db41d7cace8c63630e6f827013a8b90
z4113e2de1fc79f46fb8268bd7e86ec28e1c5bd1a08bcad632f0d86baabc808fc22f6f00bc3c54d
z2bc55145b1930c59ef9077b22d402174265454ef67cdf89e95f0bb5e0a873214d4e54dcc08ba07
z7f257b872608bea8e88d1cf0ca15908afff215db90fa7671d3d91a6c0bdce32501c49930376877
zfc6f5047caf226495f3551029d109fee2fcea54eef7c055899a8669e0eec26cdf97de0302cfa31
z992ecf54e1d7d3d073c71e1ab3109e403ea1add3124740876f4538e70db58f70d00252aacf1ce4
z84f61472609a57fe67bacabe6870ebf382131d18f0d8edfc5c41d0e2abc090005df3e12ac12b7c
z1956906ff6f992a593ae2d7c8ea8f0604422f893584de0872a58ca093765db2499312a5a3e8cef
z5c561a19d0a813275c195dda93a857f03b7dcc7d2470d4765de0fa8a46e6477ade499ceb784b7c
zf38745c402a529c0063fdde5009a5208467d100ce8388557a3a3355ade6ee862be3be7624e0433
z02b76b02d5cb488d85f8aed60ba3c8d0d90884c0c8034dd8869a98ec457591268f022eb2258197
z881341a77132453a64bd0805a3dfe45989bb778f1f91e52e9c10c31f9bf714d6abb92d0374b703
za39e9bc31bb2140ea312a17f2f692c07ee0df4d376e358773d3a425a42f158f61dda51a99f7482
zc63bb3469889a95bf276b36756581da44ee42a01d804e2180f6940cbbcf433c8a0d3868d397fa6
zb9ef949515beb692a0df8f2b463259c4c9321c27aa792c89b6a2ecd1ff99371391051b28bc5d5a
zf60c0ef1cfa8bde5004c72a175220e550a483dd3f69195d70950d17dc751a872e30088fb7f7865
z3de2cba43d0bbf1513894cf58b5445f1c8dc332cf48c7850d2addb2c2b0c47a1edeed0a62d9d2c
z73d0c7e971fbd1ccb7c0cac92b72e8a9e6b247a1cc3a2d7f9bbf91cc1e1ce8a0408d68d6304dfb
zd972134df0293339c59de507b46f80766a9a1142584c24532dfc082d6439042972a582ba206893
za8ba9679996661702cc9c4ea216a40c1069b4de6aa4957f055b1d5a09c8e72bc90776e847917e3
z55bf93d7864d69092e57129683b314835203bd212b134eb004061fe8a7fe8a7ea8220e2ddff4cd
z1b89b34db1925123acd8d1adb82da83cd5fef39a954736979a49a737d3887dcdd227d0d0250cb4
z111fada61998df32f29c010d7c6b13d3896d0e30f6b54c1262e080cb2899801bc02b9e3ff74e7a
z60707d7e0d1608255d7dd6eb42fa1437eabcf6faa5c060a1beb7ee4aedaa1562cbfb8ea9a9cdbf
zc2e95b28a5d652936ef8db111cc8b18dfb21921d133d469a073569a7f53a2b926662ee8d052652
zf67d5f7d588bd6ea4eadaab338adb205c2ab83929996df4a7423b0082a5496e61c95540874405b
z8c71957503b62243047d9619c329bd133fd8b6bc60825c36255251e37b6cf248c665f82a5062fb
z9dbf1d221c500ff8ad6548268ab35ea4316b9d81d377794fa7cb56895558bae61f10800fdbc22a
zd4e8c339775750124d136024ee86930ee18ea8e99d593afb2ab1f8d8fa259adf8119bb5ec943de
z948d8ab56189a78e00ea2820c569c136bd001d6262fb6691942434e255c767858405459b0ca76f
z2ba6329c25e7cd5223d1f418c174a68a2f83c577d7adcd177274e98a4062fa514e7602555eab20
zf3aa680dba5d045e328e11e5dbe836a3c8ccc907affeaa67e2fd4bbc8d675962cffa70f98a9c66
z39b728b0199f5f261ca8972ab74089606bf2ce88d450a17dc7d04aada6252798b1692e1a680e0d
z57bc6807aa4d2dffd47a06fedeaeb94a799682d89c704b9f815ee3cea256d3048d28c8a4ce7416
ze3e8e02a76efc089929307003c816ee322f0c8cfd39a4024a89149dd3cf44cdcc5d1a89f90a2f6
zf516e0d1ebf38b0ae189ac779376785aa806e01aea994a4f61c355721ae0a187e4a1947fa60bac
z6501cad79c969c162f9b35d34f87d9d242fa5efd984abe090d696413a1514a6bd1d960021bb3de
z0ada2f17d96cf6d07619e564fda10a7dd07756efd9099d43bf5fc0133985183d9af945ea656fa6
z92c307614359f4d05841ff8d878a54e65bf34d025c590785290c70008b82ac87c8a45e0b4624bb
z4456d45e3811e199cc78aba1a3b33a63cab3cf81927578c01afcba37ddd3b667d632f6e761b12a
zcee52655cec94a464eb584557422df7b74c3122fc7e2d2fb23d921a574f6641922eee7ca850146
z32c7801ac2b69a36dab223d3c1a11c3fb6895cf69631c88ff28bf2eab3347f65edb54069bab375
z98f6ad264411a348633790d003c49b1093312374ab7225b7a2db7526b98c05797497f4d3446d36
z41fc4442338d9dd562f623177ddb41dd718002980f184a93031bca36da3abb7f43b34d0db42a51
z35562cb36a951ef9ffead19487ed98ac5c12920ebf87bd1a0b282b6ed5573ef09f4ebf23b5c592
z7d343dea8839213245b37d34555574a13a4ceef31d5d8b623fbe4ef93b95941a8e98ca6d961b70
z5d699345a9edc5492d5a2cecc86191a37fe28f8a6287fcc361d613a3f307e9db9ccb05f1bc8e0a
za1456c0a8d2b3a0905b0c72f290f800c4e8727b96d3024091088527eba2b8532313f52bf8adc7a
z96ee018cc97be49eefffe2935195a75ed9f8b67d08d64f93275dfb6dbba214d98419cc493f2c11
z69c89ad2561d8863a2d171bb6a88463bdb076c702afa065674770c79d984cc2cda70fb358456a7
z4989926a6889d1c2090ee2d0cefbaa7a1044e36d8bbb1320528601b1e05fbd75117f30b6401475
zc077cb49c20263661e2a8ace79e7399a65acc81979243bc18c42224016bdee6363fec7ad03aefb
z8856dcbbfd097fd1490f16f6c15e43d9bb91cdb9dabf33a7ca02f04aa430dcd4abe4a76bd3e4bf
z970c8edeaeb861f9b4861ef0f5d66919cc4ab89cce047851cc12098fd7c130e1f0c29d99c1fb18
zdbcb450b7f69bca28d564deacd4eac4b67d3914aa198cd1ae245f1e0dad895703613dd9601a27c
z1941506c479b491d57ca59b9b1aeb1c8ff81b6bcd64ac1b5972034463a2766d71b07e801828298
zbe0a1f606107eb6af5dceb5c029ea6c96b7d5ff0e43b179df3746324671cdc24560d4de707af00
z0b98552f0804881a0e156e1130e008c529a0456e45bb03eb1420c724111d472a2c63ab18cf659c
zcc40140e333785a54ff01d33cc47d0f8e7140d97d0a861e31955251d9c9a8f096ca6c411c845e3
zab32b119c5a55b57e3ac0739c6d634edff8b19307dc8f2f84fea05071664e10b1be8cfe27d566c
zf51e51b68c513b160ff2d5849052c539f54b11edbb266e1f252de07afd0c2329ee8bc74ad00c64
zf2a4717d11b815c55339347fd14971ca947ff5ee6991f822c66d4c6b2e5207dccec6608e016684
z4f3fc172cd4d3740e26e820aea73b05d2d1f37b299746d96a4536650562024b473564afcbb63ed
z60f46b988c202a43d2aa32ded752204794fd8e7befe2c38c6e9e4a446648cea637e05e07a55366
z21f112dad9784b483072e80527aecdf2b08f03aa5b4427075c8a1f2df44168037612cf2fad0ed4
z8a207954159269802ce9a50d14cb37f476a585e6ce806196378ef95dffa9d637d18dbaac85da37
z0a6c98c8a1965f8fb4fc63377acb297117a4f66ca0a9de8856e97fd713d2c8ed1ed2a92ff72d20
z48a433b602177987e995b0f54c97652f4dfda6f0b076244e2bc6b1fdfd96560ac867bc04c28106
zc952804c3914317383fcfa22befb7c3dfcdab56247ca24a4e57bfe8fa5e9251850c65a0be33fd1
z2dfc69cce1a0f74093faa986a7693fc9178435f3bde4859ddd3e3bd506aac921ac80b15a48c08b
z5c4113d328aa0f9780ac2bde2734c87d876613cf37cdb163367526ba785c11f2a6f2c22e224cc6
z317dcd6447417562e06aa5b76f575634c90db734669b3989d3ae337bc5506fbb0f979c26734f4b
za5482140dc1d1d601a172f7a7c2a287b0ed572c837b48061bc895f3a36f8a2334d180260805922
zf1ebdd260f5d83fee17f23c06a12b5212579e1f010d2a97f95de5348572366b1ad330dc8e1e2c6
z5af215b5a695b95385c9abbaca2b66b1d410c398294dbabeaaa6d0d4957aefe16493ce6527711f
zc28f76d1cf64b1334974d67eb0ff3477051f671ffa452b02b6f84ac6b489d1064c8ac41b9f7d96
zcfd14517fd6b4c1a74983da645e4ed191ace3874e982ea8d8b3d5611794af70eeb8e19577f962c
zee4fc22ab6f1bfb4d35337bd96f58615283fab60919a300bb220723ef674b233f799cc3dfccf1f
z6a6f3c5c94cea33fa956a2c5ce68624e1c15f188f1590ca19bb41b750e5f92e87ae07976f8e86c
z9875139490739f333b22da2d187fab4823098735c15ba5393b854f2c5c4c51df411ca3d198e944
z7e98c1cf3bb9fc5a1b4c5d73ff6e56fa80d1dd2bca8e699e91ca99fa7534588a82fd56399ed071
z5aa50cc0af6d2d03a3f0d6e8a61c4e17c8718c24b6247a7b5756897c638da5fae37e6df70c9276
zf5668316fe2b5a629a98ed5c391ac078fd0a6b9941dcad8c7d09583c9383c6d5449bd195d9566d
z9e7d54b17a78bc42d07fc4c44761603af128a1e64e2641044b2e805aee870cf934ac7eb399c0a5
z4636efb0555d5cce5f8c6da74e861f5f8fb95f44656da39771ccd7360eec1a585a2b89723eafc7
z992b229155ae88e0ca34d4753cb3dd1da4aaefcb06542fc4c13cc0e9057c4f910954af555d0733
zd0a36ac3b3f9c0749524ec6ea4d1b23b0ab76ff38809c424204a40df8b3a0e67d7767f5c85f6d4
z071e8b38ef0d9bf60525e6a5f65290e53cccef47472a41a26a7a24ff0f0e11d09e1b4a04a2eccc
zc464a0ebba1923620daed7efe46880bca6dd80039dca795141512d57df4fa1c27a28a6972e99c7
z0f095604693d685a185987ecb8d7d68b36320cdbb713ded6f89b3114f149d3e0080c2d32b58d81
z8855346dbe97ccf9a70f723451933c23c2d958838a8fb1a912b879b821d49c4b936a61297f2e4d
z5f2bf800791d0110a7eef098a92278e62e03582e6aef38413b908f352f7407ed67801b6893bf98
z408ef0294176be32f10c244d6293cb6f9b15777e2000566abeda71d7a370c81fd361a57734ebac
za8d0cb6a9e265d0f88f26e4df558ab681db08dda21ace5fc7a5a8cd4957640fefecca6c3f2dc0e
z8818ad7c8b9be2e04798dca6a2a5848a3f32bbb1eb969f62b6de0f5afffe845ba878a891317169
z4d44284530bdb5b4c16db53e073eb59bee08df3dc4a6a07b419fddb07d6557f9f07f57b3785125
za235598b7b733b5c092c0863f94716b96976ea0d7f203fe5c7868ecfbaebe4f16d140d2af0c167
zba433aa721013aa91b6e4f3b058219e65181c7ac8ae209bc60d3b96c56a3aa6e7f4cc812e1c87a
z9b01f1906a05447761cda3e3a85c8903bc1cda76b82df3ab8b8de5fae2bb46550c7791bfd0bcba
z7e33162170f8f565c3b3baac67683d69e69f9d880d74edf30c87a9f9f489ccf7d3cf82daa2f496
z892085acbe5ebc91f800d64a7ffb0ad5fbdba9cef6a1a4424f133b1bf5a7ca71ac17335c57e82b
zff1b653845d81b534fb72542e0c8e4d82b995c39d6a339027ad491b0178e3b384a37936e4c0572
zd0a6e92ae4e6aa5e6afc79cb29cc454c2200764bef97206c855e918fb0f92bdc0200c628a475e3
z959fef3aca9c0ba21fa31e1ed233e6c0b8f8c118365d5e41991ed230e372c1270b14ccea714e5a
za43164dcbb5b1b232626680fa2dae20ca22739f8135840350d2fad60b2a21313ed9d38edf01705
z58e9ada7e3b03ac83a1f493881539efc2a943037eac4a9e5edc9c2d4529f0abb26365e34284597
z549a422faa21152862440f48ccecb5cf72a829f7e002d5081889d44bf29f956d6f68610d79c0f4
z63072f704a0db6f12c956837e7d725cf70a34331626ced053290331fdb472808a89e42f3a19ffc
z77c595b8770950d8da740a1f81a9ce668d8bd701694f6ecfa6e27535887678b4201474ae1ce659
z4dadc8d476637dc13a11f55522da5cfb737eafb429864df5a9f07cc7e6b2a4a3c128fac5bae60d
z957c4196d74c874781d8c3397d98b746f3d8663bc5e719de246919f8dd2f53dc1433443afe1c97
z5ffbdcb6cf34ab5d601a0bdca2bfdfbedd084d7932d95b7ccdb4c6d121b1a8214ec76fc3e4bbb8
zbe2c4d3506b4e6f0c0024cc287316aa4ebe84df1598bc7553b0e3ccfe62b2a13a3728b99e7064e
z7522ba53620531fdaa16c26171777cd23f458a30f9b992bf9128a7f74b03da44750e9f21d1cce8
z10d4da6b322a8620ab430ae3210e422f1ad1d5e0671cc377ce02291ef586bdfb720db98af9bc02
z5c68c8774dcd332a5ba381ee826ee18758902d33b03860092946726e0d3a1c02c9242cf9e5607b
z9913dcf11158bcc29f9dc16d87403fcae9fac944ea0ac628e60d0dcaa55b85875ed3a8944530fb
zb860a65d78ed51e84929dd206f9139aa0fbca0ba2dde97c0524208d951ad7b4fd9d0be462da1a8
zbee52bad5f81a0e6f3e7b3d4562baf5f5bad3f0884b90034167f7e4debc29fe27faac893527640
zd1b42b0e559aea59956c12b5701f9edce34b261cb12ad1c6f5d4968b1b601cb2f079e34454af3f
zdb851b73ae337aa3463cfba0d32cb5455bc6877bcfd407995bc36a66e8f3d098e8e6a6168cc6da
z31e333fd7b3ee3d14dd4b58456dc8be6308f8c178345611ff548827572dd9a9186407e54439fba
z4f919e37fd0a390e12a62f18d7726d6f60d2ae05ae77ab4b6e2ad17a494f1ec350be123fb6c6bc
zf19fc687cd28fc4affffd2b4e0995f5bfac1898d9faa772c9acbdc6c0942698ed222d08b7871e8
z6380265404bfac9f83aa476a0bb1fc3369658da6dbcb8a8529c92182b5707524cd680433116015
z9d22991b4e736c2a439f3c1890b9ee87e1dd29e2c8c20a4f826537831d68c440d3ff57eb687a9f
z19c9fec86aaf00ad1574f0b4bc33f1d3cd2702e071ac871f1243492b8ddf347de9a94a816245a6
z9429f01eed50f80be98f91b83a21d3dfac192d3646594e6cda3c8353bc5ec23938d2900c20d2dc
z4a3e70cd0d226af934ac3a0fa380f86e5e790d732a1ec1fc7ff181ca7e3fcb1caf85c50c8d6ca0
zc16cd6e8297a5dac45ca99cf21593e2e5bbf71f71cd47f560e9d54e3d11fe064877fb62892f2aa
z894841f3ce7ede8ba2bc7e434ef170c01a3a3960eeae276d20ace18b4019ba28318693a2e5b0ff
z55a62bdbe1bb61e109a6480bca5d554fb97c5ea09e45d6ad22f7306acf4588dd72d6f84b0b1e2f
z200d88b3a05ef73cd9598dbeabc9592c3a7573aa4b7ebf40a00da6b549edac8e262ff87d22ae67
z656ade6d219ce15e6522f83bbece5803b823b67dc312f76cb9835ed7e5ba78d30737cc557fa507
z781dc4fcd5633e4d7533e8805b458858a931b4aafa6af502d84c3d6bafba1116f36d78e335eb7d
zd14f0a2186d49e2f8088773e0d3a7d43a3f57e95881ca3126863768db548a8d83d3b584e9ae505
z7837b569927b07beaa6ca6cb572d1398db3ebb33ac6cb73e38cbded193d17e22c4217aad5a3ab3
zd6f88a396ae6f418308e63cf5910e725da41f2bfcd4396c7136604b1cfc5c7de40a399c0fcfa68
za94209e6c90e7d892d1de6ccf1265d40fff2f0a2b97c03d6c6744ad5d899b8486c0f251eab7715
zbdcabaeff1e36968596ce92fba0d263b7a8a37f373604eb67dfd2fdf7f8644b8a46a2bf83ba7a9
zfa4f5aea5e53b98bff35956fc9f3590a0b9eff8bd1f93b8b20b12fdfda27c2fdc68f04603ffcf1
z39f00ceba54287a9d5ee9c54146d5ab16317c0f76db949a1e9e875df567838765a68b3b0b6cf6a
z6ea023365d3ce84e679cdb8b789b9e785b63d2c6f15ab4f480b31341346995fa88ce25a7104819
zffc94ca1e1ed9d2124c4fd066545c6d4bf3b071466b23a2db14dc187f86c4600b36b3b118a4dc6
z405d8fbe53336d71d2fec7a96c9f4eaf8a8717481e322944aabe886182b8ae6ef1e41cea6a7f3a
z99c56f7f600f060d760277ad16103306247d0e8d4ce5d3dfb82add7e0d9e9e381203391d9a9e21
z7deff5e311762c15eb3c4e312d018966f30697b927b1e1b8ec72a5da5a16ce4d95acf0918bc4ad
z03c500f3ee4a621bd403f4de361303991cb4497f83a3922c82f0523c81a1a6b3462b73307df2f5
z41d631516d62f71a90e868c729a9ad14a7bba06c9943dfec6decafd3a4dcb11f1c8e745c915cd3
z3e8349e35f3e45d4db662c9ac4404dc39c60868069752bb29ff352f6f434b4b97adae628c60ca5
z8ca0aa5f81fc21abc7446cc72c39a3b21096cb1fa9e0750172d3fddde4afe03ff518118f6f8407
z64ef246d2904cec44018639d5c7a30a14b80aa3b611b2c059cccc9423a14d067768099473f3d72
z7ccf2fe12c5a9db39f6715b49b982d56adcb6c206c9a63fb6c37ec882092ef80aab079dacc2540
zeb2c0497faf46174834d42ed980c683152bd7bac1d338fa054c7a1bf93ed3abd4f46d24cdc9321
z19aaa9b219d6943d0ca8614c53abb54130f6a45e6a72dc96745adb28193130ec358d8ac8ca6d93
z97439e17bcc983408047de5a34b01e09786a77bb669ed0d06c7cb65fc9ee728692f006ff51a967
z977c1cc4ddd3ddfff0e8b48c524bc267c7dbbd9eda646f356742b0c25b0882c164fc19009b398e
z44abfbfefe23fe21f71b0375c388a7afeba58e98b27aec2c1064b1aba542679cd909aca02fd7c5
z5f1a113e053cf16eff083426eeca916fd8dd11a75ccdb45151c801a115a5fab4ee8f030f497c32
z4c47b8ba5ba5b8eda0200fcf968f258eac778da0a0e8d43229deba504b9c65f4d669559663a0b5
zb59ed054e58db30f4776b2e43e73b9304d05f7f2912714cb80145f5f832e32ad468db0c7bd11f4
z8288b10adf8320dc435b90577c3c852acd06573d4cfe42a37af4ae210f59120c2ed828267530f0
z00f0820577f1fcd9b28c14c31e8516caf32e5bc7f41197b82fca9ce10d824b1e3c136fc21aaccb
zd24967c38e1671fad0910e817546c57aeff62ad84c08dc48c6472cb1ee527ab401a9b101319855
z7187de59c8e6888fabb9218ecd779bb52e3afb691b3f0f52e1dd3909c893a85b9874e5e4498a29
z1b46ca0636bc2337639bab4ab45dfc268e4711722e521909eabc74881e1fe60b649285dde68d5b
z1eb261ace5b464ec9a9fc986f1e04c3ace59d84324b4d896892197391103f3847e788fe26cd4a1
z44b061baa4a8b02c2e0d1586aa0c5e2bca4b4e579c41e4fd4c8abc343ca784b48e7bc1293ead3c
zab88c73d8b3383dc6cef6857c2d69025c447d2dd0e1dbec334847225d204df83600fc33f8e1b83
z8bf79a11792c1862ec3d46866f29020319effc79c413287ce15481f90ae595b4911840246aa920
z76aca89c156fe776bd8075e012c0c53241647bff44c372f813977ac960ed446bc3f4eb7f49866d
ze25201327ff247df70e5df2d0541ac8952b918f85b10937283efb2106f551d57bfe8a919ceb2af
z44b316ca473ca46946998fbe198def7917d9d0b6db84cd713206ec68b68fe48f55eb030830b836
zeb3e2a3195ae4010135e5286e917e994764422b3349186ebc4ddbfa4cab01548308286fc5abe4c
za073dfea542579668c48629eebdea2202ea7af0190b1872083b4160eb9b12a60dced24b75e365b
z5fb7c6825036fad3c22a8b42bfbee23b80f89f9c99f9084b13ecb0cdf30fe45dbee5114fb1e7e7
zd7a16aa2f4a9bf3a089fa929dbaf4ab1748d7bc5aaa012a9d1c20c9fb7bfe102c5fb41721e343d
z674350d1911a17129d166e5fb3e265e97d82768d54d889ebf280949d4c0128b68183d4c1426bce
z68ec9d1125b183045ffde3d90820f98e5624969f24b2a8983e6cdd690c6bc098963bfbe602d52c
z173b62fd1179d0b0f97124cd06e2073ce5118578aa042d223ebf25b312ebf1f44dac20e0a58a79
z3e4a98206835cfb6359b6895d40115dd2e06711e112fa1d81aaec899a89b49346994c2024d117f
z45934db222638439652f8497fb58456d2aceba80af628764969b761aff1beac948576d30d3e52d
z04107ca6af9c901337a9b2e59c67485cca4b430ea3595caf2f5e609184e4e28458edfc4d2f786c
z47a25be3974213a6c44cb75ac6eea6c3265cd1f7bf7c9d0dc94e86b7cdbf6a0b3179e52281e589
z5b368795d9e9f134a2f428c31007a67c0fbfc55df99e910b78e0996da30c3de1dfbd7949f06d87
ze361fe7836751d1e3ab3cb5d573f4c943af5ccedc10d8134691d9cf468e82c82cb880b52b21f1c
zf93168a6be6c5fbfbf632520e565ff7b38f68e435bf060831ff7682f9c85a14957670889a56563
zde0435f46f3d8df7db5cc47d705b0c5abab17614b16a370a71d9f6d61bd1360d6f518cada8a0ef
zf2e568cfe606d1e70b3b88cd3f877c71d303d4aa1a96d47fa03617ec4d0fb2f30737b9dfc80221
zcbc4eeae076bd3fd6cf1711cab9b549bc3d34c941f224ae18ce260e15116df34d12e81e05ef8f8
z04bde5612d476de2b35b5b3e59b8fe3d75089be470495ca56003dd0946d7812d951a99fe7d062d
za04d5665cb408d54561dc7a53831baad5148c98989d5c7fa9d5b80902bbd6108293906bb45970c
z14e8f5d6b46bcba2ccae1a4f3322debe96d13d6f8d7af6d9743ee7541259561265107396e8ea84
z1e818122915edc0c1eb22dfc65a5c9582e059c7ba6a61fa05200625c94a8e9c2db9d4fcff39df9
z611a3a2d1dbda5316598e333e2ff8861db1f3ed935537e029d4c32e1ccd5a4f4b8400fc7d5889d
z6dcecbe60918274748f3fd46fd05b70ca973bb9ab5b75eff92ea3f68e24c535bf3a3e7f4776a58
z58b14c9e7bce1aa46cd275a4fbc7544d6cbd9c6edceb0e45126f2a2e0fa7f0ed608e41c6826a91
z8dedfa7fcf3a46fea63d90c01b8288ca5a85a80e54bc412e7226af75f609b511cd53e2abc83014
zb96d936dd37a0a294df82736c317957dba5d26f5623eec461ab711b506cb2f79904a698e8a27ce
z31d509eb9dba21e36f58cd6fb303703e4abea0c04a0c6641f42350a07fc616e6c83d3180a5ddf5
z7109f095a81e82107eeba8723501a7658aece8218c87e4e2e930e09058ab3902c14e704c1cc8b0
z0c96a7d4855c5a20dace2a3deef41f4818d0f599339a828a46716488e497c095bfcdd23ca84f44
zd5350506073b27d683f3d0e2c97d1969d0f417f4719eb3efd8549b079dd1aa4a7a0e85436d5abd
zc04c7542356ef7b8b8fcaa40ed6d6b6669abb9cd76e80f33511d7b20060688c4f5c3126f4fbea8
z0d9993bd897964f3459010682b5860790ae68f7bac569ada9be0c8106a1121412105a5bab47eac
z041e1884020808d5aa61181bbb6d22e86d8aaa73a415ed93e9f4edead3caede28e29251d5ed062
z3b8f0930ebb438dcb47673172f8afe015d83a3a00c9ec3961ea2fe44d2bceaeee561dfbb34ad48
z0706fdfcf17c9152aa83f85c15c97060d11b739075f390960ba9d45335167b6d7986b28c0aa356
z407b5bb009f2d49acc2265e012b67af10c520b7bd64d144d945bb0246f27b1ed1af80cdcaa0d02
zadc1a9c328077393bb6b16f5bb56186771cb46663c6e857d5f356f9768a276e11abbd39cb397a4
z84c25246bab4a8c485972bf85d93fe0fc22101d0bd70c835ca92bf060af543f8b46afc3d5576e8
zd69242a1ecad270e87a07b2b3fc361eb18bbda63b2a7290565a2d96ca9a208812816122f2c6fb6
z7e149a64cb6d7d92446b4427aca0531ba5d0a252d50251da59e33e439163aa2caf373938ce332a
z908319d0736cee7ec2010499c02a1c9b733341588c0be1e1f0f51d57e92db5795a0504d6ca8f82
z8476fa4b22da585a13f77266691d512032406699ba61b4032343cc8ecc0af973b261565e4612d9
zc58dc80e827451237c84b66d7b349673a8c0ddc73331db06dd6e11e438ad229313920bfece6921
zb3885ba9aca26c8f5af5e1e38665ba4a096044bced8f1f826b21d19397cbac42f669de7f9d942c
z60c08c5ded22434c517dd75308f1a3f420b97a5fca55989ea3f2f6d826212639c096a057e7c416
z0fd8d412f7845625939c5f8e2d572efe9f0127ccfcbfc043a524ab86fe6fc967623e9e3eba1475
zb6c792759e5922a306ba9e55af31793ecad1d826e29fcde7c1e2ccbc28f6c3cb195a6c389574a0
zfe3c82d399f1745ae0ef6320c73f4389e21c7038f272c6d4938ce13f08f16b450c03c632e225f0
z8c0cca39985067512f10f81c33f931d1f7f29197f9f1f8f42a78a6bbe5358d18f57da390dce796
z001a0aac9d6e9e5d00b556f6005d19444be10e62373c42fda13a020f5a48f042a6f2278e4aa548
z770dfa87c9983a035bf32eed9220353a2f3225b79a1f6e392027c8afef940339ed47256fd97d4f
zdf683adbf069127b7e23ffccd7c288d31de067f89dffd65353041e0389d41462c7e08a09a0ac83
z828d78a40593e4b0b6c8428c7e71190e923bbfdcd5d167c0412b61387e2f75e4eb9f186b90b566
z90da0a0e0346eefb2fec626ab3886fa1691396b9b7ab829b7bc0dd603eba97b9073ad04dd07f50
zb8b096524d6ac0d5bd2d8f15b38d82e9614de19e7543e43f3ba273e4c9579c60e12cd15f214e19
z1a438def0fc96466a6151e5ed4e4d3557788b35cc23ad7bce207d173539011c392307a7a6839fa
z79b638a8b08e1acc1f3fb0998e22b23eec6002918476f2608ee6a41c4fae00f175e2ed52a2cc8d
zda86c9e83587e51f010012ffc9c5c15052f267cfed6e6f3fc28af009fca6be677d89aabed71729
z21674099d0ced06293ecc9d170711b5315da16c4195240ab5a1fcd84727ee03bbfb8655a80e95c
z3df7f820c7335a3549b4ca5369df0384ac3cfb8d6641b209b97678ee0a63aafb33a1ca366f3283
z8b6da92307c2b5247c8b73f2843516bf4b9068a266560bcbc74a0bd395df4661571ce16e27a315
zeef2899c89ecd8e7c2a75d30bf5799f290d375a3fcc0933e5f7180b001ca36a0e5d98c85eddf89
z9aa598375b86e0c412742afb56b014e19fceab0e27228958dc1aa94e2a14e4d7acd4540d33cddb
z3445ac642712059edabfd1ffe87d706ada7879fd299778154f2d57d232db5048982453280d5cbf
z45874db5037a7504189ecadefe12c6788c5b098f2810146aaf51a0adbeb33d38b87406d201a54f
z621345281c9078ef87f6f0bd1bcf1d333cf1cf32df42a785815da768695c4151c62ed3c3de6cd7
z142a598bbef239288123c169e6523497c95f54bc7215be5a33bd2b7d73df3789cd2449e9d5ef82
zbe96958540c472b10baf303f757ab27399572240baded4a31e6dad077b52c82024b75dfef4daba
zc1f86d4311ce168642bc3e79d6b161e2547fc41881e2f0ba087f0760b48b357d91399bee536a79
zd10cd2006754ec736f59fe19a8ddde21c7e16aeb5f23cb914e020209251a5555342a0d5fcba499
zf88b505006db5ec95eefc3a5f715c5ee650bb8d34278bdddc282ef270f9bd587ad2b42b6b15bb6
zd137e294f7e9cfa493c3b34964aaaa2a0703788a80061aa3f3a0b79fc2fc172ab8da38c9be379a
z27942d2548e5913415c1ad97f62a022d3a78d2b00c4db6f858505b718aeafd51fb61667b45d192
zd5fc330728d0527c4add7866c88298186aeec7aaf5e36723c585cf9cbfef579ce65c1763c31a21
z37a04c2125f2c83106d010876a9ffbf622294c709fcfeb60664642eea3dfc192204ebe1cd084af
zf70f0bf4916be6699236ada7e962f18cd1b1c895d0b29fadcaa76d11bd4b5ee39123ada1f97317
zee532f001bb7291d4c9c78c003417896cb50292c14b1029be3f9af49b3ace15553ee59d92e1dde
z1352213c87b0cc40261dae3e9f20ecc06fd77d0c8f3c2c842dda810c2db505a318f885861bda68
zf9b4827c163e196b800c25d70acb5ecb0c027232ce7434b9e0cbcda2f99969960fb9299550a2f7
z9f83dcc46e5337a77e2bb35c31d6b8179b5a4938bada38b73b22f7eb13ae1f12d2b6525eddb1a6
z38c1fa7937869e0442bb78aa8aff67c920d2e4db56ce5db56b71d7192e9f5643411a2aaf8eaaab
z6c98bb61bb215ebd6166d654cd6dd28b27e32feabcbcdd0d4948ec513b33d97337349b3d4b1eae
z8816ffe9f22bccb7899e543510f19c0ec834fcad9cb104b88c33338764a73ed733118ab59b9805
z7ba84b2093ecbd9922de60e0c3c15d724f8933a67c54b3c8afa61bdfa305105327110e8bb14882
zd05108a6fbfaa15277875f1405e65b29e2118cbcd0fc1248f37038c2fedbe63650a47e9182d00e
zc431ac05d568f4fef01b9fe0d9eae2bd386bf6269912a9f20688fcca0aa3cd38e9a55c65914b58
z4439e179f9449ee2c9d7636b13fb2736143598da14192b08e3d53cd0b9abc68c8c48778d88fd8b
z1c9db76565cd6cc3bff004b6ccdd75d23ecd1cfa7c2d8b7ffbb1f4765a3bf0e74564f15b75067d
z50ecc0953625de200c678407c3fc23396317f50419a15a2e6c4161c666ef3676aa7378f6baba47
z2c0aee3c62d5f2a98239525fd9a1ab2797dfd1f763d9a3f22ca213593c1654200cb4987d0a5820
z7eba57d1bcd92ac242716e9308909ab87e11d7353df5315bd202357e6433a0181a8f55e040bbd9
zaa49b6e4a2a8c70adc5ffe2a7c9ed3b183e08e91b6160439975ac681ef7af47189b5b529981239
z5fab8b7fae74e13cbeae9ac8acc4896b58b83eaded589fe4a9eb4dad7a70d36b89d8b3c1b9b4f3
zcaa203f8440ff1f24e835465abec3d6c27a1a65a840c568cc91d4ffce458c382122c39250c7816
zbbf8f749426e9285e596d50aa7f7d3d2738912c639feb016fd84f7cf7512691918bcba5f9e6255
zbed85531741d483db127a7b62bc715fee415474ac660c2e381b377b93eec3115af9e3db5a9bdcb
z6710a1dceb30901a38a91878d2f1dcf2b8f6a7acf90bd6ac7fb05fffeaf1453f7185bd23a58d47
z531548c9fadfe680103ff48de1bf9444ab7e5f40f632b0abc044ead40396dded40ef3423e4771a
ze695e88dfbc871b2223dad0a1e7551187eac92435f4155cf4ad4e74aa766fc0a7872cf8a093665
zca5caab2861279f1371d1dd9f718a544b4de0737273abeedfd307914f498ea15feedd951defea5
z5e9853856e52c8eafe5e08c6d08b10930fda125111b4789d01ea2dfb03e98d953d464bf3c4e48f
ze2647ca5a12ee9bbfe86e43327b3cc1ad53a43f0abd248a27b224c9610d5ca968526237ed0a3d5
z386a3042d2be8b872801778360b1e94ae53b5adbf851ab89da8f28f9a25258894c904474cedd7a
z5dbd46e96926d2fcddfb2b39d4605afcd3b5bc6a758fcac85d9436935f412473550e1226640c31
z42b21b539f25811e1228f8bae48df123db6c4132c0e68ec5f57536360acb50e552466b02cd8224
z1452c8324cc8095ffe346fd1e313e7c63e4147b5fa92b174370c0a8dc744df3695a729def34bed
zc6d3af33072ea0548cd9c5d519019e870595cdd2e9c24e7fb8d4c079e3a44cf1316e0881bcacd1
z95a9f36bf4701905cf217d2e204749c8f8b5be6c7f011b4165721bb69f30e8431e1b9378f56182
z601ed5d33d877966516c00efb45ac2e2f19f02b86b348878be4a7a9e5ac913e0a7db13b2ff7390
z0c664fb406f8ae64b8894afde4432ccd265c96b80589f983dbda3a156c0be07545a43216f84284
z850f041df4b78470b729e109af3b9e26434cdf8bb9105c3a317cae8ebd8af5d0d0fb6e791a7a49
z2570bded258f7e08fd37490d78eeac61291b7d7dc8774f7bc523207360bb874c44319af9dd3280
z1b4842c982ec0a280910489f099cb41a724ad9b8e3ec1ceaca1cbfab786bd90b45d64da19d4dbc
z26ae7cbf2792b851da34a9b47907892b77fe1cab2897919f99296246a0c0ebb5ff4dc16a55aa4b
z4f640821def828278f4edb7eced3eb0826400d60e48fcd92cc35fa3cc6af0b41c0b3772e1732ab
zd28323de657a9c8c27fadd94f58f9d63d1cb282c9234c97720644c7476f20f2271a9adf7f5e2a0
ze1bef91e011ecfe99a63f10b175856a731712684dafd81e94f64a256c7c17b034b6da4a438293e
z96ca7b540e077ab34a5ad513f1a260ae81e4e34d0ea4c880a43d0f6cfdf2f90119edf81b6f5f00
z8f7bb1a4ea8afc544eeff21a3c18d03ee172d6294b0b33e8940635620ae642afded9ab6798b21f
z7e4ac653f7df60487e2c8cb2d99a2002baf3f7bbf63f1bbd51a4e3b147f0b9dc9fd149453958d4
zb16e0d259f153fa8dedf701b841da5cc194f4cf72ead787af35e3276b16babdd43b3e43406ca5b
z2bcfaa7c8a3d1300b313121ec50ad72121edefcdb9c59fee86eb7665d6efa17e738706fa4d9a86
z2cf3db2f1eebe617aa9c4aa6b9564e696a0177e2d65068f1f51e50afdb888fa6721b1d60e82a09
z677e66a586677fab7db0ff0a52e6a667e17c2f1f8a7a82af35088102c1b9c57fbea6cda575e803
z7b189aedfe326aed09cb23df86288d3ebc874d0ebac0a6e40874fcb1f903c1854646905d3c054a
zf0e28c8833963ca4c939c16257574d3c302c487399d436884fbf33f8b54d54dc31755fe7b667bc
z48a70043ead6fe1cda333c484d741978efedc7165e4007630ec6797ea614f08e974617b6410021
za448a79f94762c31e7aa504f68cdb4cafa3adee77633526f7057d0cf878a94583ae6a6c09ed7de
zc02c8224d8f5438e1e101094fe502bba6cf8a8ce041bd08cb141347ed049274df4fe7456022779
zc5bcd078e96588dd95df2a0aeeefd2ef0e9dc4dddefee59a456a829f029a75ce80bc1817211d7e
z04157096cc94f9c47bb134876c830450f77ae6c4c285eeaa71f4f8b20f7242bb01f55da9dae349
zce52b53569614bcbaad100ba336e2a440a2ac14e9b571b995cf31b038944b2772f5808d618fe27
zf2d8691867ce1ed7708b00aa4620964c93989d61b784e121bd10d456ad1654c0ecf2cfe86566ae
zc863b637defde3b83b383d2945d40222de232ced36c72db8b08a1636ae4d0dc0c94876f035db91
zdc495d9bb703c1c46362ca663358f261887d6704258e22cea24e6ba85e245c9cdf1153905d2980
z8b06fb1f09bc4c94fca4f850bfcec036daa699f6d7277670f5bcaeddf263e39048a7463e4b35c4
zbc4e829654ef4b0eb3614ddcf6db1f2b41440a5237a83b52dc3dc9f6dfdf2ffd13558035cf4f53
z7d775d2e9a4969b2dcb268f1d4073073aaa68f659b369c0376fcbec53250a35c4cb33a26ac92bf
z0ae4afbebbe296a681ad064cd4af3fa049c009d7b684c5db7c4bcaec8b7520cb3de02d88fb2679
z5ad6e1551e3d9057f0e04c2bd021f5978bf858da25c2dc288747156b25097cf6ffb99f12b6ab39
ze44e6ec34c278fccb0acca6b2361fd89c53b5cd2a6a3c542c47473a7564b9f02488be3a5faa746
z0c993e76c7b807f7ba3f97bfe31892b298cdeb8aa6b4f0cbd583c19cce0692da8c855f6c9db191
z9a8119918bf082bcf83f927b11cee3bb6be54e5149f1cdc915ba69758852266685955181ecca13
z30c53aca9b5ae475354d5d6a024bc7807d0c999262ea3c98ff94d50c9450f169df339e60fe2128
z6957c8a6934c97024844c1d4c588c832501530bb1f7f1b77e4056daaf36660c758f90645b8423d
z37f69750a5848343357eea7b0a6715b83a895a5a0be7f8dba86bdbd2b856df04dce9928ee16276
z6c2f0d42cceba8f921a6b1df79bbb99dfe7688c2a349b877afad1fc9d1a13ea9ebab10e7f66a03
z5ade32eaf4496b776a1030394e5ad56f486d4129ff6f8180902839645a94a265b64b407620dbb6
zf5a51f50bde1141b69153061cfbf158479641418ea2e2183daf5f9d3ef062f416e1ae6c813e83b
z686c3c81ec9c772d76c6915e865bff9416b253b756125b7f5c9d5b315dca72223f25ba9109a4a9
z4c4e9c05c9728ee604078f3a0783e0edd198676d3e47768196b40592fb5986375043f2eb533ef2
z58f8918ef84a9acdadd6436d66b840c17c4525ca54358d4e782e25a226f92b9e3c31a6805fbdab
z324b23a30c70087b3c1486c8eb8ac59f8c081cfc4429d01131ca3611c25a270994c408af548bc9
zb49706d886eee0f6784b949c36b4e4b0498c82b8e1f3d2b45be645ea54e7c4c867dc4858747b6a
z0f5fd870ceb95e0e1b8e9174dde602638aa216d7c0391c2a8e55fe72972824613d32b8b197a798
zcbfa76bcfcdb0dae810b4e6573e82e6c2516c1ae569600e59eeba84ebfce7e648d5a5ebfe32677
zd8e4b2274d02e7acc42c6876082b6dc90159fc3bbdeb05393d7598bce1296931dcac09c7a9816c
z05e468a9dbb1e60fc6df5a8fdfe838c8e904ba6e73962d20537b166a75c6f4ba24ce072ede835e
z1c6aa315ce1606650e54a66eb5646c86ebbd8bb34226d635f30a591c050a235498ab0efe9c7c43
z27c70c7965e58c705740d297632e41a2d4adb82091624d6c6e1cce20df009e5080c522f0281cd2
z41ffc5011797e786d8030c6fb9ccd94b3bd2bb37826fbb2160e99eba23dff978e34739a3b6801d
za02ffe2f95354dca323650c8f380d0d7bec6000eb493beccb6f504feb0441d0dd93e93796c35c1
z09465bb7573b6061a8464a228ba0aa29f7c073f9d7adc37a18d32fee6b191e7a4d1004a843086f
z3cc8e2ecf7cc94e1a86401dce5654c35924172c516d21699c4ea9a5d5c56c378d73892c23b61e2
z4f37ce1c94e0c7063c757dcb0cc4d0b26d5e82d5dbd06f2e1968ebe7e16d42ddf3861005a6f8f0
z63001fa8304447de1ff57102bfc73f1ac6602758486fdb31b0b4d0a34c1e4b4f2ee93f732ae5d9
zc76c08cdeacbb3fd542ffbcd602e7d5508bbe164f8ef470b63e6bace583ab12d673226f222081c
z6f63490d099520ab4f102ea629d7adf84b832a4208eaaeee9d397aea35321a42b413de1f557061
z12ce288910ba85a2167e30c3232b1af9d1f1be6ea1705cd68e6d10422eb10646acb0785faf943b
z9678fd0f4fbe9c59df0f4fdd7d09b396ef7d1cb92a7bfbae0ceeb55964a13da4709eaed9c85953
zdb61b008f8bd79d36fcb3f6e4b01e3c83a502b4ec9d230f0b0ec7335740254bda8da1db189455f
z305a9ce2075ffa9d09477331bc25fd96dc636f0b7b12534afab9246df29402cf37e891a99b9e81
z8483db46b568270eb8d43509b757db332fe722176fc761ea75516b14bb772c9abad31253826084
z20bf03ab6ecf97170e6cd9aef6fcd0206359948bdfbf11b966aee6149ab6969a876d6566bdb91e
zac2da6ae3b1f7f421cc876e55e87e541544d8c26a92d7e32a33f2a16c0a38ebf0b14971352075c
ze517a6d312704aa537b164fa3de57ae186b8f4687be041b161916f0d1116a47273d619e2d6ff22
z8e6955aa348552711e00a740138efba3bea8c22af2f478624c6105c4f5bc0744ed08d8e5e951ea
z5fc1167fee707872d3063e11d9dfcad34056a28919f5a127a2e72fee68e45b1cae140771d8d985
z66c9c57d7825b2bd107287f1c0e8512bd6800d62ffbe7bfeb4eccbb95bbb622e4532cc83dcc164
ze8842bf31d361f98eb46ec8c406149d7bd3052ffab75121514fcf861f120a8aeffb57d6a37bcb5
z0ce0b1d30f2debcd70b5fce2a2aa806dae8dac076c9ccec994f433c60feb6719eb22707891d970
z7d666767de2614f8d3780f93d5358c88ea29827f6dbdcd3e1dc460d6bc114cfda6d65cf1b40535
z72379e741ef43bad460cef41041f2bfb37d9ff92d21be775b3b6fffbc5a751b44ed9b12d419217
z04c4f52106abc4eb5f6b87a157877cc53d9fbb96c76339853170605c7126a1edc083306566f216
z55ef980e0700d62ec916bb33bf4d3a422c6af455c26e343ab8d9898e54fe1983e8a72aa9ff9394
z550b6fa86dae120bfc92b0dea897d937bf42b009fe374952a27dbafe6bdad35089c783e4c09643
z1376066c746fd4c542b0b2b3de8e9d4796ef374eb8618b7eec4c8301b800f292321fec849fb8cc
z71bfe8991b08a969f9d3347ef9037a394e83811a31b8202075d465efc08768dc77f145320b8f8f
z262b9c21851796f6a94edcaf225d2cfcfc8bf7733aa694ddd100472baa2efedd24bc5c8ee5e5f5
zfcdac72afc948dfd195f9c302e907a4bb6e4b6c4eb486c69f97dab3546ead628a38901a7b209e3
z70a6a94f18af07ee9e95e3e0241448a21b561ef0be99292ae342969946645ad35d0cf6e08b93ed
z4f00176afaa493833d5e1d2e61efcf790a4e4e55ad4d6a566575f480653e573a878ea2e95fd699
z978b715b9af27caed7b6e911e1d51e6791869bb395640a0c6a713f69c3c9ce5c77020017828c90
zb7b0b42619a0ced92c66931bdbfb35164e33cb5b596f691616ebd02f0414ff524d73216e08c8db
z72f8086bbbd82d4e966590e0cfe9d445fcd7d6550aa732b8740df4e0854a41d35118ade69c9613
z7a1e67c2984a90925e0013aca27f8d601e4dd5e6fca7297a6fb7bd51aef2c69a0660ed3faf1fca
z180751203dfd5deb2d51578faf2a9a6b3de402333a42d79d0a60d23a3c0070f4c8f15f8483621f
zd2682df2c1f4dc14e68747ee0214169d08fa57b88ea86b3d7396eba7f4e6a082c0c2f5c34cfecd
z72afaa77ffb877c06e01245ea0de1b391b43ccfbc42e39fc720b2b7b3d4682dc02e516df7ebb71
z0d52268cae8a8acd87776d68de6f385f19be36e4992151c661945f86bff446305da6023fa3dbd5
z5a855cd7c8b69bf89df389b076e158b1b302f606a3f2306e06ed3ad421d7b2c4dea81368d0efab
z0cf8bb920eb2e32be3d813e420d30e9eed3c7bd1783bdab5c7cbd690907558b559ea1582aa6d77
z6d51df3fc6d79378115744d3c5445a25530763124db8c2d17924b132c222a10e08da0e484a5d97
z9de3c279620e2704ce255e72d7f6fa03d24a5fd6c2f0269d7de7ca0e84ffee792d22b7fbe7c387
z3354e27869b84ffb961a852929a33220f140f0f958eb95452ec8a3fbca5c4ef4abcabaf8ee72e8
ze6e3dec6cc48ab1a48257c87f9827b6f2145b09204ad36a354a5c9573398c4ba48d40870560316
z1b70b91d024360dc9071b9f1ece3c96dbff68e76c0991087be54af98536b11ff0f68b8178fa857
zc15d8df4bee064aa498e45e4366e239c669ecb4a483be80c7201562660c22056fde7afd214b8bd
zfe8dcce9cfe8d9b6feba851e62d031c0cccf8b5558f57ad1cad445d8f1f8fa13ce70e62905e560
z92377b4cf24ffcfae3fc9c73f67f6c0ff549609206c8b7add01a5c8b72e2090bbaa133b4636190
z647254406a8ec0d19d9351729f864cb0411f052f1defb14f3c6eabac92cd0a442e9a9f359b4d77
z5cec4e2e271c8b8a9643b81cae97660ec563c82860c12e24ea6f428713190474d7a01ecc0b8d97
za8c76253bb9fe50df934ff7b5a59af414645b0a1d8bc41b01ae5a49464ae982c8d8bf97a03b063
zc0cf52bf24a2b415b645ec4fe66fdfb5d7ea4afe439a9332083a9ed960cf10b7876fa7981c7fed
zf8710948c872505a8f6c7dc839a0eb0f6463c9b4e069022cab9dd2de127faa66ae0c9d46f4e071
z0c716b796a4dcdaf5db881c39fcab798b5e265d5fe8eb8b8e4c08e04cef4bc94fe44c99252528a
z9cbdb291bff47f8aaefee60388334dc6b91416a658f87238eebe5098d38f11bb62f81e9d4a7222
z78d9b07b2e8e27bb5f2aa6493a489ddb7b3830585aca9ccd34edad6765a444d60d18f3757cd40e
zda7231177ce5f734f900843af49794251dacf9a048fbe8e5ed88ded3f5ac010cc8a4e1521de31c
zedf5e9d65f1564179b0dcb6d9a91dd458fe32f74a9359741a09f3f21d8bb67f68fba7bc016d6ce
z3dab83651688adc0ac27f9d4a6ad3c1e19e95e8e665652c8fbfcab3ce4bb33c43f5d54544914f1
z906eb0131236d8c4d6b4e2106e74e6ad6af131849eac6567ed68324b4b8eb38efa24a958e53005
zde5f5c5a64b2ae8246ae3047bc8a7ccc57009ae608298f1b4301fe543f04c31664ff5dbc77c640
z48a9afbe7ebd935960786cfffdcb139c9b378daffcef5fb0cb25016c49acd457b8d98c6ee67886
zc89573c4eba3760a6079ed43261f81cbc282ec41f6fa544f0b2a4f0bfeffa1d68e9c0b7a2c0eba
z325bd9af04ba75b6de4286c99464852d3cc9d391bb705d0492fe658a99168a26f916d4d6372439
ze29c0134ab7c1b19214bace3f52139f73a5929ded11b8a7734898ddf7630679e3a779ca7daf740
z2c9d94cb198f5071189961f0d0d5e079ecfa0a096de66f264deb0416af139c045eaa845f0d3afa
z395d693cc9c9433e1cba0ee19ba839da97bc2cadea24b69a3c7dff953c08c1f19883946201eb2b
z3069b94623516a58a53a268d9ddbcf403f5b390e093a1a9cec340db1db0d7dfca5c0b1068157fa
z4f32caf14656a9563972c3a7ec64a566e5e8b37359f648c5a69cd86b90b8a218f1fc65dde85faa
z9e74c3cdc3dc80a98005be91fed14ee717e05f7bcafede5be5f366a4d5d02e1c1fd6da56d62ac0
z0d69dbca4e102e712e93d4adf3ecdf368fe7b10ad8017344dc2e2e5e6bea98ec8137de21bcae88
zd808daae55b0b015eb2163124b69ba45dd51ba883cb3711687c7199e340506ec979a15bd87bb42
z1d7c05745bd794e75a328d7d8f034da9f3d9c8756cda50c87e374dbf7a285f28cb2c70e11e65da
z8d64398293f7300bca228e373b22370c2a2e114ed25aed686f6d7db8669e9f847e48301f53447a
z846aec1127622557d059a309ee7a670e6c922d176d567d1f5fd32413cace74cf160f08888aa5ed
zdac81465df3f92275596838c84067e7cebe04ec3e064c3a0f572a112b703e57c866f39c4cc6856
zb06033021239aa7fb33363da1c9c34ab240d922188d2329ade26de020a21c382a2f3687e8361d8
zdd3c4b11c248f796146a3c7125a4babfc1a21ec695be0c3272486fe5bbf77ddecdde3cb4c0c9fd
ze37adb57db6cda761992c7f6409be9f0141614461a0fb944ad12be56054d3b485be7fdae3291f1
z668c5a5a25ece59d5219bdda65785e9b0bc4054672cac42888178dbf5a36aa3bde0076fdfd3130
z1db2e7c4a96b1e1294fd60c59dcd6f9e57ee9e26a74c110f2025e2781c7c0dd7e4eac798c352fc
z8471b8cbffbffd3ea07261e2d25e5f316959d75180422341dd7432d0ef74b4dda5665e69ed4317
z7a5efcae14235f14917e41d1bf95532ca7cd20d649de3865b4811806eb9fb0c5fc1e7054725ed1
ze65aa283a87d55d85e63ae2f380aaa91dcb9e38b8fd1477674388cee8cca870d02b40f22837d87
z91b361476191c5a5ea9beb1c79b79412036396c669ac7c161d8b488f7c1e32dc8e0a25951e3d26
za03e3841c59045300f224ae06cd147b05fc3b3fe5997e7380df1c24d57b3c91fec6d419264adcd
zb641dd2849cf377e2fa5291bbef57563bc8ce932763bd62363999c153e9a23032b9d418e1734a0
z4b3371227b8fd1981931c767d3f3be47b3ff7d705a2b46432b09da1781082fab47c8879d7b06ba
z4a7d778a54d8239986b79fc42aa24b2bffc6e1f5450cb549195972cb9d4e0dc06ccd2701d25dea
z2bd6c55530344f7ff80b77b3be23691e89704068c7403bd9b903d52f0fb4e9e92aa6817a6f2730
ze6aab6b167e091e171d8bdc9074eefac7fd548d45d002946a11e231edd44f38bd2f4a25a30013a
z0f13b8e75a344f33af7bf573f07a1b343f1ae497b99762dd461c457fbce040bd595d8b80bae972
ze223247a4e2ee016688911d7bcf960c12dd22bb9da23eabb4552b21ecc03c21c04b7b4f48c183e
zf1f9a16893db9c366d284e15c62ff62e4e2d7d43db3764cffaad386c19366878b3bc9c3ec28bb1
z9eb4db6f8d7b1a31a8c3173fd6fc30be28c56fda12b6fcdec2c0227957938b88e4afefff4cb37c
ze0c5786f8dc8274e678c302650955ffd782c0694f15bc899f9ddb30419355e9faff160890b2238
zf4e4bcb42d1499f56c45a57dcbd9635cf7b00797f0d3cb178f14523ef31ec93ec124deeba116ca
z5b42e6c1010dd4f779b65a0c79d71c298f4be570b6bd3ab49f9fd716470ec4fde8820c1ebbe609
z4e0ece0ebd7fcf68f93f635c98c8894abc7f361269f9541883f604d0f4ea12d9304fb2c1ae4b6f
z0f3da82b64ca883754554f5347986f77e8fe65bcb7ad7d7089bac38ce384284432cfe0711d1ea3
zb9005ac23b8be2a5cece5d9abd2918cdeb8a95b895f129b3938d0e9328867b5ab6c71151577ee1
zb42cf0351b296657aff14a21a51eda4ffcb8d46c03233387805cf59dc2db28a4a364fe79e659a9
z6dbcf8553dc4f44fc9fbddfd1d5fa0344fc3fec2a36f673a97ed18fab701a9a22b253f87039596
ze2a5fb75bfa754e3bccb909117ad3b28f3f9ce668a9230fe8180f11c4f3acc962b9e6689629909
z96e4d919efe069622166282cc4baa7c49aead3e510e42b2339f574384e92100e71b83bfa508c5c
zf34756a071284d8c31a3188d01822de5995282d46cd77a4de6ac4f516b8602e3ad557532f07e45
z8ea92a7dd3083c3328665ec5cb2f6d298c41bbbba34ac249baadd5d909bcae606621c4af88a74e
z462de95045f327c204685882342f12c0d20f2e9dc0e1521677c0e729f0aad60181cb5334254f1e
z97656d260f4375c37cc4393582da686490747e683bb4ab4d7ee74d70f08eae033035a36f8f9fa7
zf9e337a6ba964ee1aae96147a47bb8d793db5a298e27a9b3ba52b2aae564281a9bedbf8a9fbe22
zf9000152e9dc8fd53608ff1f2cb9576c602628bb85bfe26dcc5f5b42e03420b42bf236631613b9
zc72a2204fb33dc7033f2cd495eccdbe1ea02e7b1ac9820476d57c06e0bdc51b4244a8788ffadd0
z9982977746e128aec4e87ccf540239049bc723b098e6793796fad47314b6782c54ad2305956f40
z8f01d0b8e8b3b291007739e3512923ca1441c36acd5d8c3e56dd49689d8f0e1277d4e878173479
z594691b3153bf961e688e12047c25668e264cbac4c5345772478feee7e30d16a2f64ca16fa445e
z9925f4db443ee8d6d77895adb33ec96dd9f5d9b8407bf9b97614480bac4fac91f499da306af8cb
za3a5e2bc6c3328841450f309531b0023d36bbf28a5a4b042aec7ff5345ca36046c5a53fffead6c
z6582bfea587b0548d4b5946b5d24714cf0b16dd5ad0dfda6ab28203a158e3efba88bd2f256e2d9
z33681a6139be325666f33b127827362f2363e2b663e9326b57e584752bffdd3daea60e65036711
zd223abe880c548a7b0ea3a464072fa8083c7ad7f2c6b2da35307b3f2165e423320bac4a53bd7af
z9a54f4361f599198be661945e933d8d3cdb19ad8ae67a672fdf539d8eb502c7b811cd162f110b2
z7f778d34b51ae04f8337bea1c5537f6e4a085fcd83828265b1d07de254f0447d670f9689eb597a
zd1c2f4f04f38a8cde346a1f5fe5a2e2c43cd101d942abde2d3dbf9582b71bd0bbdd3515145f4f1
z0cbb1806f2d15fc3ce90b7fbeff3f7c3459b488d897532d01c07916422890e77ba06d245f72fd6
zffd62ea9553b4ab7ff6c28bb41251ba1129f695b2c1e9b7b02ba3cd614a2ba7b38e75d9ad4fc46
z6455cf42b46352244380aeb70aa0fc82146a23cada702498b828a20034a9d3bb2bc3f594daca12
z88a4dfc4de80f47c3ae737f2f4936cf22fa23e979300dc687b4863cf90f5e311a988a0e3787666
ze221a6e57f87cfccdb0eae1454245a2212b666650433d860b8224e1f27c5aa34df7b99b138541c
z977487594a6e2b5e91aaf92a91d29ef38559ff752e834db54689da8e5963168704b4c400226ca7
z85b280f19896d6eac151bf024ace6ece93e361ed9fece4adc9df36c20d9bcd93f45ea602b8a165
z5adc6513236e91f73be2e095f1bbd559a65d026c405512babfd8f75122e33041ff2ab71344d0d2
z234dc411ca524730677e8a1ec16f569155d57bf69101417b76e42ac79d13134c9dae03504658a2
zcb6fe2c5edf8b668cc8e1bb907fb1d9e125a61bb703a0ecb5d7bcdd4ab975c208df1430fa25cee
z103d81739f6c3c6711985312700ac37f47f343b292b3cd979a6fd260e5827568fe5bb9ed979359
z08951728c6786bd016af6fa46b0414f22a0cbfc6e814fc10630e4c1fd64c751ba4eb0c96bbb003
zb85a437118d0944c0e981bc4b4b183695c1e965c476844fd71ac487a11874cdfa336d9cd4253c7
zdd70d65f13185bc9cc88e8cd17fd41ccb81919ff9319fd3294d1511c0233f59b9c6716d204fc9d
zd445eb94bd5706d0debbc23d66e44d09b591dec7fbc9cd086809c002970245ed4f8c30e41977d7
z7b43e4267b167943682cb9186b145831be655ad619088d2fd6316b62789ffba926bf280442c9e7
z3b7cf7b6c845fd7af40f4bffa9cc6b368d89bbe2bdd040fd462a60e3811e70f370b237a83cd909
z87794a7d4f1aa242798ff2b295681c46ab53ee79c7cb20f8570b0256a5ea3e080a52a27ed94100
z8672b7c438370c159a6dae9c660ad101c2a1ad408cac8a7523057a167168c1a83994edcdac7212
z3ef4d2fc64c0216ba5853f76a914a6e1507831ffe556d19f84b35047690dbee2b64411f593938f
za5c705e68dab295a12e994c802d43de2d8be69da57a6daf182d427c275e4991d82ffb20bbe1ceb
zc951200311c2ec2bb4d1ec06cfb810cb3919cbf89530919efc345b7b0a7fd2a2a03389d4546616
z8565e1cffb7736da209639e09703052642b8db911d4d5f085872a879ed6998b85765501b5064a9
z3cfe48888a2215375d7b4e1d0be6c4df771bb5368c774d3ed551db0147c9dfc477d3c592c63b99
z67aba312e021039fa91ec36fd6711c158952bc7d453bf9bfb2d5dc910c320095b7236103aa259d
ze8af3fbe5f4f30690bf67e802b30b7f1b9d4a004560035ac225d8d4c4bf5fcf18d3761a29f4b7c
zfd978b550ee8101a398a21c6afbc492ceb639b6cd22ccf2655fd6776c169202414106236b0f474
z30531c80019deee77cdfe891503f956fcc3c51ff3418386c5058f376ae8ece0417ceaccb1c3ea6
z9fe1a725bf284df0d4cd48207fa1534a82fd698a299c484b01e3694601e52d481ab536300d0b95
za886d5e355a0f1c5ada5e05764200c83901d1b9b7912f1c60cf93b366ddb86491d935d8763f9e9
z5bd0495e6e4a539fec6f9dae3fdb865011c5c6e2cca325f73aa387796e8554c128d769cd517b77
z3fec74facf62ff52fcf2b05998e41356fa43851d498fa43a77c74589e58be3c2b2488cf245b982
zd64bb7c62773b35cb2806a9df19d279c67d0bd5ef5a14775526435d41c83e0659b0835c000f1c7
za67d7cacc0761a37cff565f8269bac794788f54c47314555cbdfa451b7450b2c18966be6e5f48c
z298de3289890e1b268399e5fc25ce8c1cf18bf758a63d683eee915570bedc46a611765abb1a6b2
zc3a28022cea3620e926b2286c9830ac7191f467748522345666f9b98b3c5aa03324f64f65be81e
z53aea086614352aa5b14a87d8c85cfd732000a78eafb6ed413a3c7239956f90011b2647fab6e22
z68c7a871ede434472b1a74463a61fc1f4e20e5df30010ab2bd7f8d5b7b64c1c0fd8c727824fbd0
z7c8c410aad47823d67ccb7f7eb9ebca3741ec9d401566718dcc0849eac959a3ea777683a53ab11
z64422d1b8fc6211c69ae3231e3fc7e917a14f713844ee4434f0c7261627a33127417ccb1597b56
zb0bb50be9ed0337eff2ab1046ab73b58638b4aa5df06fc620987f2994d9f4072b5dd273b6b0942
zd61cb93525fd11bc02594a8c29f5ec79d4c281317007230c939da7a621270a6d38ace3b4b8e4b1
z642617894ca5998cae8b4ff6b7d2904c4efc9c5d6eb6c0c7756bdac78ba62cb95a43e0000926f3
z1186f89c032b32eacd96597963849ee3463882c64835828cb75d06903e94f6ab3762e05d2e13d6
zcf3449f0d948f3815919ddf4a0d504c5bd07c62fb8413dbbfc0525a306908a56b96cb73ac002d5
z06b5d3cf93ee0e797816bd5265e539a540776a0fbc86d94a0513e38b01d8fbcceabd54fa3176e7
zdba36ac7435bcbfdd1742dbf34ac4b14790a3798e8346ab8f05ebff19de6118da55fd0de039110
z9aa2b06a90f66b6591d5b3c0ef6fec9f1d0a7018df002cb287ea88322d7729f8e159eb9393c76d
z1f7e246d868eed0101d332a216dc074a5de0465efda466a36439656311f989bd2d222db6d4be5c
zf5407e4769dfcd0a3e42326f93adacfb17e125a37b9006f93d2355a3c23235d55d8535bed4964b
z339e6fae0552b402d6c4b04e016f6a06907ed837938a243fac222e4125d6be124b17c10dce0471
z6b69e9a73715ba7e6785f7e07627dbae9dcea1dd77e899660d6998218067d887e5d2f8ec64cc73
z7ee1c80425d1bf67bd13899056ac9098b4be6f56a819b7984729ddce8c0b11d3874a1c8d5f0ec9
z30054ce064d016b653a587d8f0cc3d1042ddc0049dec8a03cd39a43f8ad4deb8b5c3e99e2d24fc
z017a9323d5295a1b99950f4a6d2aed4ed30430e8c50f6e70ae13dd78e29f9056b0a55ec9603009
z6e88d5d906521c516081c44d606a66d357fad594815e65cfd72c8b2d38f5fc5f24067abe2ab587
ze35c2a2291eba0954ad5c6dfa1f70a9cd0aa5feee52788d425596bf7d6648ba5eee38239bd8e43
z072b6beab44888c9e89b547015c640aaaf16f23faf3e0d82a29b94a3f4d5d1b600ae2fed72e113
ze977cec37ae82edfb3c93184b24b5d347fbe57e91f7e410ca1cd8ae742d49717c5eebe10cc92d4
z95e782672a509309a2e98b861b8deae1baea9df3eeee6fa9a48c5a1755807b2d193df6525354c8
zcfb71f119191a23dd123c6732af3d71bce02bed459ac736ecd40f77eb59eba67564ef97e02f55b
z71e8981dab2d24fa2e96c517ee4452c73bd8cccea2649858edd3ee1aac44a6434f4c845a61fbb5
zf9d5aeac80999ddcb7432d993b649f99bcefcd6a2a434ca0ca66c45fca6ab9ce42d35c2e513289
zdd74b05307803d520d3be729fed99d95e72ce804a22c2e80cc4c41efb8552f28967e85bccd739c
zbeb5c0064abc415a691430606ed8670963ea9580e8abb7f0a1741f9b7489298d7ba36cb9a07f4a
zebc035b40cf27cdd7b1b56b0ae454c2206033ceb40acc06c2e785badf87ab665e6e99a3aeedf6b
z0b9b0997f2c3ba63a9efc6681604c673651c8eff6ae3f9e0c6c99cd6660bce2c07d37548f06552
zc2efdd11a057fc8e1586bbf6d6b2edafc05ab03dc33b1485feb7010bdc71a03a2ec214083657f1
zec37776951c5e922accd935501b48d69eabea4cb7f0d3ed0114bb5dbf057baa3c57811cfbc2466
z9a972aa6e8e0962773bad4cbe2f48e34591463e5d32fd64a5bf19d361269696d2faf5504e2492e
zb5deb79ec6a9a231612c43b6ad468b3b5cbec400c8713798b1c32ad61d130bf16bb8945fea4adb
z58c1803f5925fe07c021953fb9490eb06bfcc1371cad5c7a4f826f34d877ab1b5e1b93e2638b6a
zef36b61056432c349326bcea9de60afc3d148c5af070ac69ad29371024c2cb6ff2ac6753f98c90
z2f6cbd12b677ef84ac209d47928940f1cf299dbb8059f7fcc39b368c4058243f1c6688e74d51a8
zad939f53e0eb58db7127da7802971af6a505fd4d40e247248f102dc63b5d374ea48f00dd9d45b6
zea50a6ecec390ff0c865b8c64e520a140b071047d8ca9ee998f5a596be99f6cb1329259e63ad59
zb1ad3026e75a0dcd9343e972187934f96690ffb2a89dcaad308d61ec245f9e3f989d32c4cb3afc
z6f24aa3ed8280184ad4fb8f3d1ab56e49303a10e22c0844da484f99503cad8521156ffc648d828
z3cfafeffef767f6667f337948c835ecb06d730339ed3b24762963da433b58dfe8cdb7be0f8bea3
zf4b0acefe56fa19cf65d59161bebb2f782d8678e7e43cc6b4d1e0a63451d032b3158acb6af8be5
z1287d52af747d6beed74c672efbb1b91b48e24b9a76e941b0e438810b2f67e980b42f11b8607cb
z86f188bfe3690210175e08f3a6032dd62a58fd828e3c871e2e4a3d9b5ab3ccd5285dee761e6dc9
zb21edaa7e9701c9547b6cbf5b70cd460e09de2338cd51a6e83aa0f394316c42554c4c950f9aa12
z1b94812e502b0f91833b96c9ffaff90c8085d84d0ed792dac3b0f5bc55dfeaa0efa26387dd2230
z1e746b1fc0ba26a423468d9dd419703d81a6c346f9df46786521c0d8ed4e77bcc56b93c314acc4
z1710a93c0a080de380673288247bbcbd294071a34cfed10a6593db0d4d4c2c0355846fe089ca6e
za80e8b712e898bde729db83d3e6460be8e68c5f9713a17d1d109f3866a5b0949df3ffcd05cde9c
z2fe4314e7eb34e120522fcf8b255686bc397921da1a44cc5673101bc0b65e1fa217675928a7667
z40b98586086d15f0a343aa078edbd4c0bcda5240e60080e9aa2a67aeab0a4bdd4adcd4ca1b9415
z11a1301a3c4d17f1f4ff54de88355eaed894fa9d62d51d35d09bb0b5e64668ae047f72067efdc0
z34c89d2cf430dab8ac9a597847686592503264665c22a9fdf9bc8f9609a4ab769244693cd520e6
z42f3cc873f67d4a3e27d18dac3584467933241d8d5f54ab7fa5a1f2ed606c38790fe944cb874f3
z1a30f9b438f20c7670f671c68a524ed1020795d84a12e96fac5f96ca60423fb6f88b7da5267ebd
zfff812fd3c5ddf86e883c2df9040055fd2f8e4298f12bdb8881ae907bd5de393a6545f213b3182
z73b2a35561d78f37065a10c573975717ca5ce6ba835259a49557d94386bf91d01ea3c5eaa6727b
zd369eeb05211dd280a4042a38ca802c7ef0e201bed2a9331091b91745f5e0955dfa0cd7732573e
z6c51159d291dcbcf722328019fc60e703474e963aab04fa7e0ba39ac9ca5689e241e992c617871
z949bfa25a2483b97d96bbb5a1fecdd23027531a39b713f54fab7da3febc561a3049b1a0fd52fdb
z8248afb37b589b014132a4ee718f531a5995840e443cd6aa52b378c6cee82d3fb249c4a4f3de5e
z5541451671165104049801b237cb7fbfbcbab9fd1a3b110efaa9d9d81a76f7be971e2d096d3609
z924a85459e121bde1214542066b4798ec81544bea46c6808d8560e1900a59e8e2b390985db4b00
z3e393ea5dbebd0389294874e126350cc8e83fec70696f06d51ebe2d770a993f1599afb017afda8
z5c23c6196e9f34ae4d4b41323ffef2fa5a695e867e803869615a98b88b0ca5e530513507d4f5a5
z2e578963d63fe5414580e9673dc614d9aa44ae754bbf513d7df31384ea6cc352af7aa7e3f7424b
z94d50697ff49885820783e287425e47c94640baeb52f09438a6be6b4b135cfd8a7bfda6832de62
zf0ce60ea181bafbf0af88b37b6b45f1f6d4e9aa5067ec794898dd275cf76dc88d27618f0ea27c3
zd2f0d6d23de23d017026ca8cddb0e128a896982dc16f873c37a37e4f00ac00361f993c33a775b1
z979b8367819415b82d07c141701dcab27b1c4444b727b6cbab420ba88562ad9d326af9854a19db
za5c47a743f0bc6e6f05d4a97d868a850668cc34a8d7d69973cd644a62b32e0fe93797cac57ef65
z0027365417c8f9e6ba8a3be86024401194c68d075aca33328421b2bd7be4f7cbac4ef1093b9c85
zb1592fdf04ff15bc2c5ba13d27922bf09ab5b72deee087ab2a3163311e35614262a257049a2142
z4488d187bebcf5ed9fa223a109b0c992a6f981786da4d1491832e35afc7dc3b6da67019c2a13dd
z1ffad79f7dfd9e75d3ea3f0a8040f3fb31ccb0ff1fb6b10759f5e7fb9195462d46e793dfd49375
z1f31d5de9ed26a2c5bc4afdd806aeddee25abf90b984aa66e382fc9084b80fe46117ec67a73aa3
z3701e189c6baebea09652906a0f848edd4722c48671dbfe789eac99ac9900adfcd12754e902955
zb01b87a3a6282f12f380de05273c8309423428aae792cdd3ebc5ce91fb97f7fe36541c774de85b
z887390977a2a78aa4f96a201fd65803116ee802ed6276f554802a19038a70c86fe57cb5f317085
z0876002438fdec15b341acce3aa9aa0713427568dbbf1349757f091a105adc2a2a1097781d0f2d
z23bb6bbb4d9fdab4eedea96982ec2e31efe9d4a93ea4d1d429c55b6b20af29e2514103f542c249
z9eee05d832129221144ab8ec01c183fd10c260a37d8bd8fbcf92ee2999107a98658f711550456b
z4629f3ea88fcb21468e697761e346bb987dea9a90b77b7939e4ab0ac4c0c5d0b409b6c6dc35d79
z4bacfd3e565dd8f61f0575e7e6c12f185a4658c43fab83dec171399451411e131e5d5da2614bce
zcfdd19c7d32e161174d2985d3947a31ec059d510e4c9f340fccc30e55ca5f3c45d4ad36c24f21d
z7b35a459fe59fb40d8e04e8ca6762b4ffd99e96b20c457fbd129389c5a4d8098769cc53c3badc4
z722810d99d77d5e1b80d48cce1e2ab72297da5009efe15f328d7acb3b04e3d53ec8deb1968e208
ze21533c0467731561db76c7436fe1b7dcb01efd448354da786793920460c99edac0032bbf320b4
zbbb52e7386c696839dfdfbf0ac3e28d849cc3727dd33ffaf84f812016350afd6d3121548646a6a
zd13eaaa17a3ccbe39f8326c12d940b317152425f3f20b092b371dd01f7d9700e0c09fa96b46db8
zae438320866634f775dbc9e34274a5cde5b61374f6694418cec5e02681313ac0a401bf04f8dbda
z7506fea7a3a66685d8d27c5162033f82c24e929f9bf5fe32c985b22d09c76e136d162d274850ff
z72fa0fa733f32d089c0a6f8e9815c6f82bb076a0e8f2f4a212b98d148d1a75611485df096d874c
z15ab41e358bc6765c7a84550f02feb144fce82d2aa8479fcf30bbbe66e72849ae10affe12e7278
z89c7581ec2b37d70a2200bcdace24fbfaca1e505af148640cc7fc17a44deff2f32f875f3b0b90f
z533baabeb944bfdba9451ae03891c299deed4f5ce3e7ab5b4e15b957bf269f109d4b05c0668402
zfa280ffb8cb8a8b62e252849b97713c4232147e68903044aaddc7245d51023c42fd8a4da225613
z6b85b97ceb1355786efb46af21039c55d7f96a4649f39f066544d295f2556df7f6347f33cee067
ze956dbff57d45c65ea7a25c8b4f5df167c1bf833137528fd55080e57131fb529a34076d2cc9a16
z35f18c35901ad31258f2e9fe0c16c589be4f16df351f77af7ae48a328e7a47ab1f9b433d5619f4
z1be7ad8bd11bf78f354c9d203641e07eed86f8b9abf3d289aeda37274267628a02f871d1f6efb3
z0e5377dba65c582ebcb8c12b3048c469cc9733a29fc8dda2db9a40b89bd0187b85c88e601d6689
z5fdfd31bde98a9c437098ea6b80dbcc7cdd1fbd447dfad9f6ee9a31ef2f9cbf8350d6aceff2f18
zfd3379e5b1edf72831398630dd625504dc6f0142d2a73ef428dc1c0c3a65a0800349ba91779b73
z3b26d0bece484fd7df542c98e0a02ec6da23649ab583f0ea0eae44efe3487e15ad514cab8a493e
zf3433e3cc953d7bd4f715d5b1a389b88f7d729c6fcb09ef2880897cced58fea5f8ea798471123e
zf0f2c83418e18d11f1f32431de2f838d79ed52a25d992f9905d020f016a3621c6cabcfc9760d18
z304dbcd37f551a4abf5855ca581f4e458d58df2c76af7d8b9fd088e35fba793201ad485f91ea8e
z7c3024dbdfb96105e60f019f7ec641b79051d06ccba413189bf2fb6437ba86d27698f35d5b55cd
z2a6625e7da9487f794ad88e022d6eb4c2256d2fb23733d6b59413645cea9af2bca9912a0d9d93a
zabeb5395b9263c7f3a42c68ca4390592a1a844a2f7b490fb09950999e524d4b691ede876ba1d51
zdd11b36ef1bdc4880171473a81464006cb56c32dfa434393281f832930ca2ce561cf3cb3dc551a
z4eb4822007128d6c0bd13cf0d171bfc6714aea74b11d3073ba75d2c83a028eed96d5dd4a3b57d8
z017370b225b9aa817c8f27f18ce1b5bdfb96a327fc5c82e5babb347a31dfa9932f2b80dc4b9c67
zfd6d996aadbf74ddffae86cfa61654ac4ce77ff462e99a8e3884a8a816e50aad1b757ee072e9ba
zcb1ba82489080e42c36b2d631e20ee1f68766453095e7d1743fa3ab07219cf12a57ac54fba3044
z0d984d73f957ed85ff716ccf0c80b2eb0ff820af7433552d4214cdbf73ac30f3027feb729ca260
zf9616485811a79a2a2e5d308f96ddf4add40a203b778fcb747af4ae28344c9c0d5185c693ba1ef
z4550a02012c00f34b3c3eec275ef1ea4d780b653b37802fa58eb3f6f9c151f828771938b73f8b3
z4464d53d7e03248fdeb139291d71b161c720161e2b328e78d51b44bc8a60e23b3e4688e15fa209
zccff3b3418782d39224e40c85aa8829361f48764a578f3fb9e9da75bbb3da5b0d2ec4a45bcdae8
z8f670468193fca5ff61889eb11d179513dd57efdf56375dbb29f5ba3b9033bcd20360f6e7238f6
z68eea88d6a739bcf15c9810cd2b368127249238bbe9168f56a16611e22d1dc99fbd230f5315547
zb1c5fe799af0f6cf6143ec8338f7e942c52001623d574506d1f26f6079d691bbbdc7f3323b57c2
ze7e23ae419c2bb1792030ab9593940f8b0e55da053986b5a651f43e783316f10f86a0eea4f380b
z742188da79329b377496c28121be2f44b7a1d951885718f9f75f8ef0bede9bb848d42927a2517e
zb1c729e76ae9623ede144d8e8202027f2747e6f40529ace586feab62b118ca20d0db17d9bd966c
za7d6628b660a6aec90a54d0f3f91534c0cbc2915cb9caf0dc3355757c2d477577859280aebe343
z9ef15dced5e748ba8dcf41c9ec9d94bb6d28c7aabf8122b50bb4e795f69d38766616e38e7b0b39
ze47ee5fac05bde7cae69a1b3ea42537b413fc7c34a81cab6c680965b9e515d5cb79da369ebc62f
z8f24648f32d1b9f94b6c621a9d6426fc253a528b847d606a8c2135db629394d5ec18f16faaf281
z40b09cba8bd53159208036303d700d66b7ad483b0ec84f42da603a58ef34bfc529de78c029155f
z006193a70827afaab7f8bd8acd6c163d3949cb2697db32e305726f79ea3788f25f74bc724c671b
z0a4a8492e299f2d0a62a98bffa3a9dc7a68eccb8ea1f39d5dafe04a0d2f8c62aa861db6acf50ca
z8514365e9443c53d49e29f1a5a391e154dbf7cabd2224fb7019d39db44b8b92328db0d358810af
ze51d382205da67f45a2f54c16b095969b217588baf8856864f1d21a664e510b8d7bb331e81d1c4
z91ff1f23f4bf7fd187572fbbb795ac99b9c9f67fdd4f422acbc6cb174223f9de8e777d220430d3
zead723fa6294c0a261898eb6e66f3eeb8177c996b037890da97aaff475475d96c13f5cdbc4bebd
zfb3cc1850a173c9ee65009ed5d0433011017af32fb87440b559f534e785f9b85c015eb4696145d
za2143ce99650ea325eb55c910dc858b1ebb6295611fedcb9018324ba29a9b983bff4d45e54a9f0
z72dc0cd155c600ba7406cd6b010af8ca09c61323fd97d38b21611b1ef2c512a6d35861c94c362e
z96b302f1a70be15bcb94eb1bf072f43d45bec9e83873a810e4dcc98b2d080231a8d122141b9928
zf73ad6eb7ef86de716c3a4a1f70b129fdb4e487fce7f0b4e4809a14e5a5f45dcd58bd47179c8f2
z9917d23e9a544e8b73ad32f76174b9fc55c60f920ecc70113978787f4f6f42f15d20ffa5d458e9
zb14bd6477b40eecc4df9366ecbc4355776dca6473e153163e64c03e44ac9326b43c0f8c08efb51
ze2f37be2584cd9902e295901f66642d14c6c251b4d0a8f4e837ad14fd697c05bb7190f1c4aa4f2
z448cd752471566793227c23fd764546092875e5c3013232ffba9fde9de43e4a431f619bd5a2571
zde3d75c4dec6589b071019fa3f469eed299f2ae7924d227a6ebc366855e23e444424c5d62cb8b3
z2a18fa85de7f1436309b1877295ddec6f6a433358268e36ba904c1ea400f5caf31fb40f0847a6f
zc42ce40089abc26365b838fc0377d1c7e4533df2d344980ba596f3fb06783d699846f1941346a4
z5d8ee93be2f5842cae0a8e6c4e779b340bc63a78c4236de0c168d4cbe848468e18484013912e7c
zb6c15c35f713576ff5250c5a80210ce35d155db62b92dd1f9e96311f455678eda4ed0df1efa942
z54c0c9fb4df356cb37f005d54bb02fc87cbaa1931e6255eb1103ad6c6a7a5bd9170f436c6e4365
z4063810db8eb6feed91c60cdabdf527afef253830a37d218245f954d38c798afb35fb3437dbe44
z975a74e93dfe281256f80a6daefbc85d54f2165104ce10425639783fd480fbae6a9f1e1517f410
z6e41d713e557036433e5b84960b688faa9eb9fd4936b9f57a38bfe09216016b49004b2fefdb300
z6bef0627a643021f94a4f3aa0bb77e822d8755770fcc12d8cea4657420ed53d91fbe9862e02b1b
z0da57ce942b368191679eacd8456f3864100117926bfd9a8be5605c166ce7e4b06194a6c437d7b
z4c95e3dfdfb453d364d6b6db6cc5c8b979279447cd9396c0e33e68ab4211e5d54d672fdf9adb7d
z384ac52cf2b14f776007a1fc01665edc27eaf6c128b04c3b5e12b00d2bcb44b6cd5aee37dcc751
z375a63cef07e9ee1d311626923078ba46d88a1d55387e798a1dd03057c19d2b939ec477e4b2694
z90e5f52ee10312ac23461f945292a35754972a0bb9b344b2b91c662b1a301c8e46bab49368e98f
zb2db2426ffd869cb851124b533375dca26a0d6997c8de75f57f72853043316dfb2c74561975bda
za0bad7280a73cf863a4987848297577ff1ab843f6835cda2d9aab51f7e7ed71e161539045f37c7
zf92bb70000266147d5a26aaad15d4930d7e6a4dd3d968502deda2c418b7d519c3f1d390806e214
zb47034597f6952e4614db50822090e38e1905e1bcc7d22c0e78427ff88993b7344c9d4df4a63e0
zc325b5f7409594a875f3a4e378967db90c4ef4bb24339f3af898a80abcadabcfb3726af233b03a
zc5ff60c8bd489b82a82e499506f104de68d4d45f2735c5e36c918a8994a9a9640bab305331e3a5
z3a37986dea6b9293e203043c3f9f7c4edf967b92387d67220e7c1cae4246508c1c936e6ecf8cd3
z4ebd5ae61cf51b0afe6a3b6934229b8b58e59bb529acce8f87e0ffa3606b222246253442c5ae79
z70f83516059814a8350b2b1a78bfda753c4f334f710c8342525b01823fd7a4e9ae7b20d2c40105
z9c1cef46cd1681773b08bc5ce08541c3236260b9b47dd5b5431b54ba08b72295d19cf2b505a08f
z9ad9480ac382143f54c4b2719898859a824f464c25e1e548f8a663520a15a58631e1e0c05ebd16
z246b4649c4d0d481bdfa209e5bb33486a0b6af4193d9523781e9062e55d2101fb3bdf0c0ddec84
z2216c0c58b7d46c150cc92874087d347c835fdf92e880576195ed158428c0c4a02fe1746a00bb0
z5989781f46c7834b8c1ea7a2fa9923be3fa14855dfe0cc4d882f027ce5ae9e9d96c8487f5f92c0
zc04119e8b3f8dcbe358714ad541e2ac2727f1e373df1778632cf01a4be67540ffe9678b80d734f
zb2773355ffe206f21ba305a45a1c922596f844844bf8d96bd7ece4230cdf029f4871cc6ccb8a6c
z1bcf81a75d376bda879b03641630cae3030c7898e319a3f0d8307190f1ef9c06eaf83e7ea244cd
z85918d364aacf2283e1e4b296d7923a2d6c82a0e0d028ff9ef1f17c1b1b044088fb84a84e2428a
z024c8e8e651541dcc72aee6451a8901644df2e475da68d3056b7278dbb20fdca287e2f4cc94617
zff2aeb0c8ef0862a58ecf2ffcf44f2e3a78c37d7b1e5549dc98a4fd0c4293176c1a56da0bdf3c0
z62867141e64f901e7f986fb5511c9a80630cedf33fe481de47bc9cf48a88087b6ec2698d42a95a
z32cbc6040b87d9c35bae7947a93f518f31d4d86f2dd0fc9e46468456a586a4bcccef58066595d8
zc081866a2a58afcdc345e6f612934a8cecc1639e5b6e1b018c4718e79dc605a9c85c8f9e091ab4
zb9a39bc28bbd01d022f8710aa79301cd9f6fac065a1302153c870c6d6e773df091c5dded729552
zf316a46810c6f0067f5bf356c6357abd71b06e3c819d0ff1b2e84eb51185e0a4dbd2efc46f3158
z4bd5ea964f00cb62f381b6a398733bf9c4f2082b0cbd349779837aa0cf8699513479a7b0aed2da
z2102516670d771f9004bc1790f90511848e4753a1d1181634ca16c7531ca797211d976ed58c9af
zc5f2e7b9ab19c0ba2234375702c71f92356362b788749705a05b51ac94a6a4a273a0d4a40bf674
z33b5bccb2f22655362b7a965db13286c91b8f1703924249f5294607842701eaf208c7dcd434a1d
z9d3b7666b543ae9515d5640d9a8471f62384e91c803e819ea901dedb2e485a13ce540708128173
zcc84fea6401fd4553800055354dc77b409bd4cc2cc75e61d0b1b75a2332293e527f645b64201ce
z76255744243062db892efb0c45b30912f7acd01aeb977fc8281952e6786216dd591f15bd8346d8
z9ac7f4fa815ddf58e2b242b7a18dd9186b355abd7620ee19f055bf6e6c4f6d06b68111bbc75e4a
za5bfb83e36965ac92f654c56253317e0cc59eb839f3ca4e1cd4f16f0f1a1bfafd1f8d1aa68c23d
zeba3001ad8c8db91b8ce8f99a69cba26fb8faef743cb5fe622cd50a71e5ce874e217b74f1b0dff
z59bd8990f09bd54def89cbfcc40e654f8b1cabe1d8d68ead89513007c40d3e531cd90f1df92146
z11fdd506cc2ed06b8c7ea38361bfd3a0ae6a9e1cb4a58c00485ea2e851b343ec32871774eb4b22
zc7d78b22d39434e8ff8c85f2a8762a8814e3fb0281cee52b8fe0036df9322895cbb7d5e672682a
z91c06dfab97d06f14d63a69e4de49e3cfc3660b6759213191e91947f6d5aa402d4808c1e511eec
zb5277bc3dc185bb3a8d0580912caa64031230509d10b5b19df6db78433d71146217754f9e0af97
zf3f4a650a376e73fe0e6033719d542effebe01d84c7f17e9098af3caf2a30f8c23ee68935f17d2
zd2570ca1fa81e7f2b927ed9bdfcfa9a843b7acfc33068d6313281008c6212825f6210c6e1a8fa7
ze64f8e6fdbb484618ffef480b77694bdb7e28e8a0560ae5a8747905cef162b470f22842aa99149
z00229c69c098c76803dfd7a67297bc60af8563061763675bd38e5b1da8e0db7490888a60070087
z16aaa231b03c54935f7cc23d75ebd8feb6e59085406091b3ea7ff82a857d3373d9e1d67b6fab80
z58170aa46c29df02c6a59e21762ce5a65f599c1c1c3ae64ba4b7f6414b76c70810a912cab07765
z0738b17a0a316e491bf0de8bb72f8d5a396fde24a24e41a293301ebc96d79de25e09028322856f
z0067d4c8ad653ca99a534a9a00d6545474a38d206db53481ed2d5ecb0166946039f5f08f3ab0fc
z3a53292b95fc8ca5dcfd7c8c1016e1d4e9341de7d0d007f155f735b696d175176fda6f9c53257d
z3a4b571518142b197d071aa9cddebe56247860a638fca6a659de268b897ca9e42af920338e1218
zae1d211ca801f36477f04617081868f052affb148d7a03106edb0565ab0ed7019951de84df60e4
zd1f51a23ad0a7741d1680cfdd104bd0052fc0531e779110477d3785699e0593567f652352f5a55
z403b46302dda9b4f5747a8bf74e0cf8b2a71c73abb01b43ccbb7d1bc05852cef9547d1c749ba5a
z92c26b446ac04f228b3e8407eeb1e3aa6c6c5bed7659b9a09e278aa11837ffc9c8fc1fb0910ed6
z1ea4bab3a5c6118f4bd0dec7477e5a57707d48efd2ea97a846ca933c9f6de9b1bb5a72dd53a5d0
zb63b0b15fb2f4c212b7328b4aa137fc4f3ac38611ea6be27f36fa58b978925e06871ffc2c36718
z01818f6bf282194db721f10b90503b681370338609b7bd47243dedd911f2d058e4070877644127
zde5d7e118bd3f96d5a2d7faf68ab5ba5f6910912cb373f46cd94d82b3efc3766fee5e5721d0fc1
zfa2afb0778a8d2dd94bdd62e144e6ed571544e0eee070a1c0ec85d296c2552f33907f71bafb074
za27686e5a79698c70db03e91ebdc60ed39ab0a8cd60915a732c443b3ab8eaa71acc3d60b28bb60
z182bd54e8a9a8f1a4e6ad6f7811318ad418ec8a03a2bf2e82aed6083bf2eead56cb57b55ce3e01
z31c88d360783e6a66561815956fc309cde666b275bcebc48e3ea7d09e8169d3a24558d36196abd
z76b68afd1e38808bc999d144b163486c96c615c3d0d329e2cf58ec074f4a5deab734f4c0752a3c
z9859c372b360fa17da00910193d48667b2766b2eb219fec0c9648cbd2eb2d896267d8b9ab5d0db
z338f2f72369414da6e005f7bcc7bed06ff1fcb595f0a02907f5379cf8c463c6d8baffbb06efdf5
za8ab007b11157ab771b492413227d5194ea8ada5660f88e9b14622c8089b371feeeafcca0477bc
zd465d46544fb6197b30a33da435091f6ae2498365a019bdd7a3edfc53bc804b2e709807bec351a
z3c5f4ed1ab77b4de6948b60e80372d9cd719bcbcd5b7243276ebd8041a9d44833911869d93e86c
zd383edb4c3af0ac00ec97a93f399f08241191379e29f56ca1903a642090bcb43cb4d91f10f2c5f
z6c72402b9f622f0736ab2f3894030ffc1f24940e2e7e600a48dd9352cf327ff819425044cd4adc
z00bfbc50cc11d757c600e0bead62a2ec14948bb2d825037a9e557df35c6b5923adb4ad4637e904
z9f3748d7803c5aa18518282c8e842b0247899f79aedd39fd0ef6b43be24f01c38d4d1f4dfe9fb1
z2d01f7314157b3b434d25394fc2725931d1d7095026b9ab2b8e0861f93e7aac3c0ee28a0f5954f
zc55e7d581c8ef405dc81b4e15b830b6636daaead27f1cd24a9f4f046dcb5b2cdf076f539b17bb0
zf68538a71a0e5fbb18a28f1795b66f0e27f211ef1148208ed78bc425b8e61b868f1dcb3ea6971a
zcfd203d5f256339db2cd752e3c7dad8f4d978f4434603bdfd2503bf8b6e3e7b42161e6faa26a2c
zc5b8595622dc279944de23a5f47181b79703c017b8d561f55b5042351230b02ba542599d13e050
z81e736e4ad1e4a26f9a88cf430c9e0d551e6f027ce548e6dbee3140df411697da1868188a2b658
z0ea5689c0cace22c09e954b761675ed3bd323a648c06f1a9330a52a63d388fdc7c805242daece9
z094f1aca882332e68332afd6b7ad6cea6f710e9f5f3c4b2e3b065c437e356029b530273410c6ec
z2fedd0865cd23201f36bcfb9139b488ed95fd656eb42764de1e3a325fa9057d70f260c64505117
z4a6b5eb7525562266f00519336c0d0f5c6d237d93a85524cc3aa611d824631b172e972026fedf9
zdf85056b67606153b7c6d2ccb1ef5b2dcacd6de440fd4408ab481913520ee10d6e5c583a101fe3
z6c649acd86de45a2801cd0fff4a8367f0824397328ad9c6cb50877ce4f6688cd442e41b084080b
z1956de31dbce15366643d1ee6fcafba7e0b4514f3a103ae4cbe6be10caa5c11a229d60d4459ce2
zd938a8227c75c2775ba569a7ee9a37529d0be5405cf2a0055dfa5b0cff0876bd19f297b4be0349
zc313103038b07cd0e96f74ffe43f6eeb3d648e0459c116efd93c2aa50e36cce46730cc8e2678e9
z8cef45aef8f55935cf890ad1adfaf730cf285161c005a942163f69f27fa3fdc75f9b50922e33d1
z3e6894808886342188b023cd839070ea2c6e75526bb7dd2abeacb7e1ad15b836c2128a4822dc16
z0bd7a21bad86222e5b1168b4913b946da0276df82e503d24356ea368335a5244d9867226e62ed9
z59f39d4d2a3867ec3ae4749235518c03714c1f5529eed1418f200bed121b902c567d05d601f1f4
z48f84961ec95cad03c48987856e187d5258b9a9a9f2b40efe0317383db2e23a4a9ff4fca29495f
z5b06941b0559176208a828492dfc6bcd94b94e27250ef3f098fbb73ee83300865065431f485f8c
zbb7f63030da712e89ef603cf051916bdf585dfc2f6a69c809e9962473c791fedc81f73bb89f9a3
z651c026009c765c6883dd35d0e16fa261463b3939bda78514a73769ecaba8a9a88fd9f0a3bbd25
z38ec20a8d90b0d7e8b78b2114d6d4bf1f7a44853e33b34d20043ec2b810366acd7178ef6946be8
z394dc224a5196576c817cba795b782da2488da2b3d0dc5d951105b8381eaafb45430630a49565c
z46e07945cec1e72ee7f2bb23a839195db4131977b360d83f2a51ced5c746bebed8690095cee7a9
z91c3a9e55ab928dc127911ae93594d0765ce0628d760c00eeee9ffe3f85f34f9a35a04a6bd751d
z38f873d6c0f6340881fd6688c13b364f20d7cee4dfee83ea1158449c10c12c76a8916376878554
z0048a525a07063f558de9c884e3719522ac2c86125efdad15d5db06d4465395f240bad517b093c
z835bbea53c8141eed529a9694c2a876bf6395a2ac593e9a673c75ad21f45c33350b3dc91bcaf18
z5165015bcf88ead6e6f573ca153194f6928714691ba209642235e5d7f58c9a0963db9ddba5ad90
z79cf78b5ed30879789387addde1ada1f55db8cb9ee628dfc45f99c3c1575b703c80b97178e96fa
z311e098f03c8508b9bfef52373d377b7fc34877f380ac3406a7d267e5c84bf24dd3d2ef7f9bf68
z6a3bf13179a37bfc15f09e1a387d0f94d93d09cea8a404baf90fba0af3e03814b248f7a7229cb7
z1b34d9d7be24b480e8b0ee1f23339128c650094de9d04871a219dda75b01f434c54d9ad3358429
z57c4c0521b61b6ff6522dd05ca343d3cb635e1a7dd65ee46b021d2590de46312656a2392a0d69a
zcd9d40e712c392455a8d98f4b40958a502b0f19c73a0237f81e7f8a056e98166ae017c04db7574
zd0d7c1fe492087a7a87cb8e018335f8032c660a9068a01b811bf2913cebbbeb8a390d18892bfda
z18c4b051c192391b33008f51b379e3b3d6fa5b8160a7aa3897d2caec25228a1dba52acdf4d1d95
z8e6083f4b1471d93d31a71f1524426e533d4d0db60cad11e6d15cb7b41eb71b74340f04667559f
z4bfdab8318efc5ace26a62db33431769f44b617add88f32b07395bbc7fdbcd716affcff0bb47ba
zba698250421a48aa3aca5788facd8e671e0a9085e60e0f09c0ec4f8ce17e2f013a1271f758151c
z5317b1ca3e7d62ffa4ed47d6184eb60712e64927792cc70ee8bbf480b29e23bbe3ba107c53af2e
z37f9263b0f0f0625adf7795d0ba7c8beaf51de2ba16a2658a5632dab80e67eb4197960b3520973
z64c3f5ad3ac0a64925f904f37206c0d76d4f38a80ee9f2cbc27172413746d90540e662a1d46937
z473db73a60d57c00cfa15761f14a23aca8a41f6ecdd28305b6cfc8c177d733b7390e06ad4dcd33
z94dea0f4a039e1df4d83310a800836fd6ba73cd71eacf2d1caf625a9e4622b5f2c82062aa8e262
z9bbeb93a18c21ce4b01af9bd17887ed5cd767614f42b60b2de07088fad3b724b84b2fdad575c3f
z1a8a4fa905b1b3e72035369d56ea6116e9922210516f30470bba187f585cec076e684159cefc0f
zcee7dc8f93c0e43ffecd6eed382ca474951dd120064f0d6deec5a3c96f88dc31f4e1a735a96305
za891604c32903d5ff602f425f5ab7778794c4b26703939735c5de3515003760a7669beb381005e
z7d0b775642d10d63df707579c9f339659fb243d97bcb8074af9b004dd67ac052c2a8f98c8541a4
z85d2c5d5ae0301272f53784ecafce820f26084d6a1b645083fe2f59adb9c17cd0b63422ce161d9
z46c292e7364a09d8ebaff86f1ae39c06cccc50aa528ac98fef13bb1e5c71f663a2e58b7f77c6cf
zb9a11641fdc3c47c0302fcd15e5bc667ade1537fc9a13586dd28b990cdc97afbae8929ddb67dd4
zf48a00d48d1c7d835ca2a7d435e9ed0093ead4f16bab2e55e1572ebb00e2bd9305e013465fe685
z1b08d7bbbf16e893f4f16851d08a1a29c509108f3a0714f994c9d883053fafba25455efc7dcfe3
z952f344c8962cefb056c884413e22d540cf341dc2c1b4d3625b0b81559528444d2e806a628c004
z53174cee5e81d5b5061a51ca9270920a7e04763e5d5de29cb4775e29855611d4b9947507694be5
za4a4a9131c819ccc687a3eaee632768f58061275d8ec32877dc2a90c1119ea3829456ac4010d42
z907cc9458e44642a0f7731b788eb94eecb37af82a5445925e7a8807f6f8968ce7d49de4ddae374
z35794f7bffad4d6d9273324171195c44a4f3e30eed81e5092fc353d4685a9d38af0d0d6877c9ef
z47e2ad8f1a7929670b8cb7fb471eb6af3d7c52e4b0e556aef67d692c4df642169ed0d2a2e4def1
z22c594bd56072158ac5c4c4c512995723e46c76986b4816787e691a1320916974cfd29344be96f
z5ce27ba5e33213f62ecdeda7486dbce3f3377cec9900ef0b9f9cb9395ffb03c19c3822f10f8e97
z1105a6e0aa9c0b160dc1f0cb8063c94cfb3be165c744628204abd5da9e9f8d1e38a6dd6ac741fd
z1536bb99e3dd138ba5bb77d5594ed4519453e0dbc6979e6e0290737ebf768b5879f04e3b160d8c
zeafe760603d1d4e253f74443dd8bf089fbee24b250f7ed10143dd2f7765680f0fae96e88ecc930
zc1c7b52cb42c4f31befcb16aaffccb1eb5388d65e678670a524d46bfae3735f9b0d0bef585e39b
z8de1f412235d70d829d92fbf88e649922bbd89c995b75554999bfe6869a839a5c632888077681d
z300fc488795fa5546e1db69ab18ab8b0cd1778604caaabc2b475c9d686ad10aa08611c61b5a0c0
z24e72e34e4aa42d33e39aaf4f5aea85112ab88f5afb7abe551be51967a440841ff3b8154b71362
ze7cc735aa82a13bfebdf517eb7d48d701205e3bda96da9c93456f8b716bb67382a82f7240c452f
zaa24648d26ee8cfe0bf148cbcadd07d7ac97eda2508b77caab0449ab842ee6b07e85a2e1bbf599
z943ab85b4e0391474a5967258dca9649222fa1fbcd22f327e32e3bae2fb73c252b242f37a277f8
z4b9c674145f956a3625f29403ec844a9605d1adc3f41cc67eadd2f0271e76f26f3314fa44bd509
z3932a6a82fa9fd06072f9a79d47bf0f0abb83fed1fdf1e6a84a87bf7cb03c457c951bf335e8c5f
z84808044b728ada55e570e000d7013877ab009f5f9717ac1f19eafae35eb07b940b4b7d5ac9a61
z8fe375740ab9fd7f00a28e65122354942be4e24bf973fd1b87ef2bc77ca4b222c7292067bb7554
zab79fbda31c6dec0492ca9d41cf72409d02aba20e62890c5b49f36bbba514d21c1ab0d911aa986
za3d64b92bd2bb23d0739bf43ac0befa151521e1fc44eada7189dd35e3363b667067ca2ed98d1dc
z55e8cad222044711dbd6973e34bfb78cf3a2898c189f146e23dad2c874650ba40c2c3f3087317b
z6261d254104c4eb0306e842d2fe5475292d4b3934a2731ceff89a38f7daf362c108a4b572be09b
zd7988f86d13e62af51323c2fabb12d13daa296599118d217abe9171c64ee09aff5681be8510d7b
z0c0cc83296e84b18cf99e07a736edf6279e1a65ab28844f0c9fc3dd0a82c99e6e3ce6dfad0ad14
z58172bbd59fa07abf4c20d55298b4dc09b1f42cfd949b07e693b8bb9ff80a872b6491b628f49c6
z0f20ca67b7b36831805ed416381caaa5a44c92c8361268a9d95e592b0c0c40d94a6a64dfaa5dd8
z6c4b1876f69156f99429edbbec977fe79f65c458b0aa2a3f6183e8c3ec0d9137f6f311cf45b579
z9a5454706316a377fa7d24c9820907fa6faaf8c9353d58395c4da3615fea985de5f5a640895eae
z6a1700f349968d56b767ef82a4954e0b68f0abe21b0f7f459e3333a20bfe26b8efa2135ff10125
z1591f026ac5409704d009bb0a59f69864e8a589fe915361f9c283950b144299323a10426c6f3e3
zb766c51f664718831c9c71745c89ddc4ce7dc82a9b086dcb0fa9cf5218ccc514cee15132694bad
z4c6c2c4fb1a0ce56d2cde54d91c430db9db90d4b4c1c92fb833f13ebe9cf49deb14410d0131a94
z6c52e62a8234eae46ae0c09f6f54841c4b730282a5dd7b25f34dec09a75c8f3a0bb7f01690c58b
z923f8faf35704010c8aa9f4a95b925568d35e169617e04106edb205447d6b009848823a5207627
z4b8ae5abb367d5fb66fbd08baab883081e0d8ef92a13c2e58941aeb0487991ca8d8b4fadbd8a19
ze097ac55f40a28c4a26660a574673f1a63dd4ec64b59a0be5a682f57252eaacd3ef34fd4215325
za32d7b63744aa594c6ea76788fe1a169dd40ddd81cc3ec482c37fe00d11cb76c0efacbe1b46569
zae9afa4e3ca7974c377aed477e234701215231c7184820b66b3a0ba2ec0487580e2c4957ac8feb
z57e5d743962778c79d0b2f94b9e93fbe03c751bd0bce1cb561c06c809c6c409d3f57eb7f8888eb
z63f645b5e5e5e48ef612ca419573f6c5b8c2bc78c0b707658ab4857602e3326bc231d772c716de
z3013a589a3d02ce6632c7c6f8fa12a2863257692db9f1748abaa7865eafbf5105f36e15110b958
z1435ac7f2cd7dc7998ea6a935e1bc85b729d87b7bfff3e40aa8d9a0f7d63aaea679d2f643004d7
ze69280edc6167c8485e6aa4fd2828bcd1db5783188ebee689bfef7d84f2f986b22354a352b1c47
zee819596d345eba34eb762d7c2747bd9d34380a5e9159dbfafb1804cfdf555cccdc0d26ade68fc
z33b2668fffdbf8a98fe15b7a3c5c61b7e92d2fd4123fc496f30d6070d237b2903c3140f0e62c09
zb415a19943c37bca19c0949badd39eb0d8592f7db01282657a6f0d6398744b7001a051736036f4
z8567a64fbeea3c8ed877a82e5b4de50c629cc4dd4fc41b5aac40093afb9a89bb47f6eb3ce1d62e
zaea36c5e45813a7cb62bfb3add2a5f279a670b43994b1d3a16217f735cd10a8eaca6cf86da92d1
zb6f8f0c4e0cb1f7162b063c6dc6a18499f2769f3ab9dc3735e10982103345e567b65f92e764446
z04519d9f4784aace8492ce31ce33294ac007025f5470093ba75a746b09ee53957ea69e56007243
zfad62dee32e79209af2b0749eb5930ca215789dc65f00f8305c4f373703e09e009e5b506ae9377
z2051c6289f00b4fc5274f342dcdc66874184cb3bc58c85e9e2dd1060e6a2a51dac77ac86b8a9cd
zd4f23dbb6ba34dbdd7bdd2fd1cb53a75e594c19841084deb86ea579220c7d67a70eeac97992b26
za4a4ee64b7cededc374e06e9082ff9665ce6f42f1028c03847715afcf39ab151b9bc6a2323cf59
z61c4571dfc4a72fa52e26d4f60198a5a2242c4c79a469144b7721855c23c8d77626658584aa614
za36166658a4ef5992b68d08b8b5c8321958f6e5774231be8c17a1b5c513da9d745a3d3d258f72d
z02b5740ddf06bf45b50720f7da40f3906883be5881237e7aa65a0119a9c6654784e79963dadcec
zb6d53ae396c0f522dcca3610149b157fe7cdd981ce5415c6241b1d88c7e63591b38292c80fad24
z5fe0698266652236555e4c202c27e017cf851bbdbde646cda725d48834e0b28654d34a97cc1234
z9922c2fcec002906e8f0ef6912f074efc27bae4b3eb699c6dfb3dc5fde9baa8a5fccbe58921954
zd58c15b8e0fead6bf2a68661e272b7f09e6b73c863b371a888ffac7feb57e32a90225afe96af64
z61dec20469e903553c48b971c13a14f910b87737cc01730a8367efb98aee60aeeadc6989404f79
z645cdba849909a6c8b2aed1751469d4f22905796a18ecee4c692406307c88df5a0c9182999be44
ze8128190b6a6821fa33f97f3cd5292eae8b516ec4af2dabc66063fb28d400f819d737c33861d67
z3b299a368d3db991a70c0b4bdebde2ee1306d9f10cf3d4902d43c417eb4c7ec348707b958bccba
z8f09269cf5707f3ca09e8e4477c19384e209479d78d248a459c9f985847aee81708f6ad5c501f3
z7851d0367b763345db42412b97ca472a93081af0a91d8037a9e1795c799b40886d092de85a6004
z3a1ee687a30de73269ba6d0d0a76b19133e9202b1a10d19e4c20749cc837f33f680978be3d2f31
z957cdf1099d49b793f8c101ccf0092cfa698c2d948cc33e83c2136fca1ae95fdb81a40a3b7f7d1
z2c00ef7960075246411ed32de2dc9bb0154bed7db53e27af40995e95a7ba270031817495175b62
z8701801093967aa9bc6a4d968e762b6081c40d2edaf9d9a4863f9e52f4458e71e2129e30417937
zd35ee6726bad13baae2f4db19ca158066fc4552b9364ce466c3817f8024f311bea7c5337d77481
zf70b70651affaad83e4115c86d014765aabe36627d2ed436cdfc6e98618eb0ca1c42579da0c24c
z60e405d9dde99165929e01d06f81366cf336a8c0adf664d885dee4a9677a0d4a46d8d9f77062d7
zc872c8d06346b2c9c0a79959b0897bfa81e717fd64380ee43587e97d84e83100ef35ba6c871d5d
z9f444c53da069791594a531b1d02949c90b9ee8bc9a48ab4fb1fffcc233ca51202095bddb8ef3d
z32a70b7eefa96002bd312ff44f7d478c460387b666a1ba28359d1e371ecb35446ef1512e4a7c41
z3fc7b23860d9ca33978c731126c350375d28e91fde04e23c1003be62629bbbfda993d9d869c0e8
z26f62bf72f941e68e5b8dfa298e2737c07ba2899886e2479ba18c81230de59b2687165e6166e18
z3af8760250678d729694d5663af3264e61a2fd8b6000e987e3ba29af38222ddd38f3bb3a9b5148
z75076328f73eb244af6e0918d1d66c35032912e7efcc66933ad70e7582aad9851e7d06e08874dc
z4df5672916cd092cf5207ea20983353d849d9853a064467261bca6be932d0ca4fc863e83c8717b
z48c260c661da75074ada00e885ae784242287e25fece97a95af7bc1591496638dec953996a9cc3
zaea521f356957c88b2f6280725f931231703eb65e9cca8a728cf850d193d3f6473bf7c24500f87
za72e3052c1e37106bf828a3d239c9110b8ad1df1750de6a3fc12180669811b7e6b44ed81817871
z42ef31aff1c69fc61fa0edfd67b7827a83857687dd684a51ff3c0117e358b11347f3f8c6a91559
z4ac2643725eaa13581a0409ea71e2deaab95862b1a21f37ec4f3511a5f99d674f0e2251575bb09
zcb9e6e22d9c31f1c31567226a6cb456641da2bd01371740b47c15ce2875eabcfb61af10316e201
z260aa8b512193ba621866702a05781dce4792cb3385d4703c37ee223c77e529e1adef653c84e29
z5492a0d8c5216a6d7bea28b2afbffff3608f4331eb040e55aa3769e41c8ab21de8d836bed8c05e
z3b898e848db9fdb3a5b44b2e0ef165ca274c9de4ef0c5add71c0c395b8daa44e6e83190d16bc30
z8cda9718ff9a74ed83890a64fd1688dc8fc44cc6e1afe0d2ae91704bde78aa0d4786c9526cf074
z7712e084a67305f203c72ebddfeb8439e423a405b59594d6ebc3e85816746020dbdaf9d801c1dc
zb6c27dae126cb6f9e7aceb1271a53da43510b5a96ec805c9e89d9d04092975ba4c2caa464c63a1
z1dcecf94a99a6d2a4389a9be9436e72079c79985612045ee171df467f2729a1a11a8715cff36f0
za8ee96265947726e230860b0bcf32e609099e04a0733651fc7dca5eb108a65d91273520e4a63d1
z1b8088e2908d8e8c3af5ffce92dd0d169cf9be4b467efabb8f1788457e8787c1998ccba85925c5
zf51b22f053bde8156da7bb61838e11ed5b1f2a47d674f1bcb5ae8b6ea97543b713f07635b6c523
z9446f6f724f04262dc964d3323ab1494808a8ad60dd18c56aa6aa7f63353e44af979155433af8a
zfbd728a6873f61af5b7e01f3ca0bf1d9e2af3138b7d40fa167aadfe43440f09ac3451f9db07a01
z96060914c8c8649e229951916c4ddb549d0f9d2e0c6ee2f3486d6a9c0f48b66b271a91cc1b83fa
zf4fd675f01d6f1b60074b91419b6c2239a0f98f671e32c1e185afffcdbfbc29e4a18c44f36ebb7
z3dd44f03c8eb0541ce507bad9612e2d50dbddbff4a26f3bb8d50a5bc5a1ece58a7441f95aa633a
z509bf313648e99c3f40973e061049cbff54feda29307bb2c4558e2b2037f5703faf855c1c6301e
z2dd59f429bc64ec5b46c38632591df5c3305d4a5b0ad3837bbb68f81143a8e86a4b0481cd54ec5
z4ab085e37e81f985cbcd9fc3f4890bad4ee4d10448cacdf25cd24b750989299e59603aed4d27b8
z0515738595f3a287fd1f6d7d197fc65d67e7599418066394fb71c1b04036f1b0b3c9fe9ca7f564
z30a1626a573fe1a585b1f2fa27a31423256332f0b8cd700e6a56538466f65cf3f1a6863a93fd50
z96676db849679d402407b855bab8783ee2d80e93cc77624e2c78d0cb7c29a0d777283b8d368851
z522b8993102727be71d4f8fa4d075416b0a78c4f5fa6e7d91d522202c039ec7b241906dcfa173e
zd0a553ab546a07ed1349374531cc2503dda7e669775904cf5eda1e73dca1a5848a3be2f0f53836
zdee2bf4f9ccfafbd155203998dfa6b88dca796936cf198cb71221debc0d8e6ccbe8e21ca758323
z0a893f42b7a0b18a782ce79bcaf6468ec21fbaca9882855634493297d09666c90919fc1c3060b3
z7739117cbcd218a0c6f667fe87975632ea59beca5ca562e1498189e41307bb82377398df25e984
z305e41c385d1f40e4e29318acc7aca79f975280ba5d3b89ef2dfa9b6cfd363365adc047bc61856
z362c3f087a130e21e816cb539f85fbf99d8efd0a3ca85df847c580db71c9af8d510bb2809c8d19
z4284a66a4807b428a7d6305dc16d6d62a4fc0966d1bc9457acb1d985c84fcdc2779467069df8dd
z143f9ecc5204e9b8d4753bb325fba63f2c7455d02d55ecfc94942abe3c92f5698e3daacfb7a6a4
z3843615bd009765fd865b4f00eaafd96a2432dd6f68ef96ed589e0ffdf1afaaf5f73daab3d5c3e
z9a3eb896c1ce1e14c487539202362b54aebdf5a266066a39a14daa53ca748fec5ed46938ac0aed
z8d5d61ed3900ee69cff80f33de732bce6b2cbf3638aa0aa842fc8206010d9748ab72578865fa5d
zcc21118822c09215e913b7dd52d6d6ad72d0cc619b6a48e3650028bb03316bc5bcadc53737b571
z30c146c0d4b99a7b167d29b25d83c69171aca218f3eb9af549a574b2a95f66fc736c857051b2ba
z033546e767ad88a2ea5b1b694e5a88d0ca0c87e6cfd10160be83e68305691e97ae68a43bb0898d
z71d866ddf5b52a8c94b609931ea6ec20f7bd066f41fb560984569ccf8e34d02f2e8d0ad21d2d98
z4992a65434ed31f0684eec1c65a01742b88360aa32522bf01c532cc501c26e8f6b187eb85bc703
z3c0f417672566b0817873b11afb13d7e30910351e28d449d433b09230111a2c79025de40c2cd37
z9be978ee3221d2339a78684ec797df87143a6e1cc8e078556170701e80da229fea33b81f31eb69
z0517653e4f480ddd401d833ff4e423caf7d789b5cfe0d64c413148ab5e67bb9b386f14f4f238b7
ze8143c8e820a0c04059da49800664fa9263f7ce0a40260d089b52df7abc7e7905447bb5d47655c
z125ef77b47de3b7967b9c284c0ad99618d767313dac7c93ecc72d51353c080f6b86b1b3cc706ab
z75c7f079847039debfe22b0d56ff99346fec9c3c658a5818a89d3e6015f15c89d7a38fd8e11c5c
z5326c1efb2cfcbf65adefe9ca83939a3cd81d9ed3bd996059847af2fad37560661edac46a476b3
z0f8d8ee05495e206789dd1b80d27d863643a4d8d4e1ee0ec7abd3abf179d3b1b8e43aa322b3dea
zd1577ff1f23c4365a213ef0af1a3af651e249dd84320f618912b423a9605e65d151dfc0ac02046
z35cdf42ac57a63f331cf2b8bb7ad412205d1f4037b7179c7a84672cb5b16fb47b1451c45a7c656
zb04ee08bf2f7126bd1b4d85d0f545906389369943fb5a186046e11f1370a00c677221883a523e3
z3b400fa19d27451c502fa700c306cd617da2501eda9d7fcbb465bb11f9effeb316eaac8fa8ad5e
za7a1112a0a14a0a823c8d6af92579e30731ba5696bcfa54122e12d37d17a382da013545d8d39fe
zcd9282e65114d235fedaf22b69b3663b2de6d41f67d8c1a945bc2c9f19ad86e10c4f66aff16aa9
zdbec36f37ce8acc4bac457a0fbfd3760f539c1a3f6e5fe5d6f77192bce348ae68d30146a10fe86
z863a380305d0f115c3b5986ec7b6dee3d307aa7fa2b7a46ce6c065a1d97d1f09c514379568e635
z9ce46c934caae105a230aa9d16b6d0ef499ab947ee8335a209f1a7ae7e86b7116425f3119764c8
zea2e7e83ec9797a15c491a09e6cb7caabffeb8b7dd24ff94cf83d12f65e7679d95ff23c841c68c
zebf98e1c1ff645208d288961202b8158da3001e31019f80cfd2097a2a7e183de3b0cc532f3dcde
z1d67627bf5805e4988a1b13cd69e3e2ad6f0786159775bcbd5ada9d290dc5caf888043e9d9ae76
zdffcb06c7360d461dc66c976d9f6dc362e199863853ea4d5a18248d616130f15a62b446268ebe5
zf1ef97fd75f38b3709b3253c576c89d544352da8c60b72c5f81247788da661bc25c17d54fb8d92
zfb7a4af1cee0683a184a86e1e48a9e3b16a0e180a841b067ff5512488b87efae83d1fa5ed3016d
z7e04f22f7064d01516a56668d216ddcbaf7a770d7f706d5c308a0d38f94f3576a44d99b40e9a1a
z39e9c4b0284ddf394660c3d540d481c62f5e6fed76df4d75c2ad494dcf63c468ce82da7ce6fc11
z722969d994a0b2764c7f462d5dd1078f012c2c1b0447d3842e4ec1222729626b1ffd5db6ee87c9
zf40f1757fc11b46f9eaad08b4164ebe9157add221b527f6b8bf317e100b58178fd74e45914d04f
z2c36be2078ff1d623cd84f05086b46772eaeaa73bcd81b1341c615a6285a4ccddb105207813d6d
z5037ff718722d61cc5e46f9273290b42ea4b1fee683c1dc090edd16f6b14b8e71f229cbe1be00e
zd3d4f005a97f26cc5834d89802c83f80506ec74d7d3f64217999fb24365538dc43912f2395840e
z12b292fa006dcdaa515f857699a7b9f90473b92feedaa2673d71259be3ab38b5c9cda61b4c9122
zcd6c7f53177d15284e37b56dccfa7180ac3f750ea902c66f87209cab6faccbe1c03eb0f46c5a7f
zf4890ff0591bfcadaf0a61ddf892192cb50923eb723833f5caab45b834a89973ac37c83ea41ec0
z3bfd4da5bf7898a299e38b931066de4e70490b043eec0688ff4e3df6054d4c98a07654ccc73609
z71c900f6c6f4f0c3c86a5a855044b6ad7f5d18e2daf325e187aaa83b92fd29af334ba265c206f4
z7f98371259d11a137b9cdb8e9d2156be15c27e33473f985efafe3795674e4aa134f99c8e3e22b0
z679de2550f963b179c572040ad93a4f1973cfd0da3d5c9c9a3235a6cf7b0512f72e8e8e0619181
zd651752c1424e675698f668c8e4ec9f403eaf4eda4936813ad759f0d8ee068a2da1622f56c05ba
z718121fbe6531bdfebf87ccba86bdfd68f35f5887efb71f0b383f7c5f88957250a7a1508ca1494
zee191152f92cec01a14b4378ae67c53e79811ef49c1e0e57b80d94f91d688a82f3248f469cad16
z358994b37234fb1ba844e1d347aca6692135d46d192277c043baa52b03c28e0ec278769b19846d
z7075b86b03a17eeeafb53f16d1c182891ebb3c3a37959b0f7f8b53f38b42806081468ac00e457f
za71967e2091cd87df3ab8b1cf4442f6f1047810b3c4aacc183cb078056ccc2a888fa2e743b81b6
z90bc14633d2e3dc1dcb89e3ac7f67a4b4907a21d254cf5471e4402cf26c79e78bec12d4bbc2f8f
zc6004764c3c2d43283c8e345df1c1cfe7eeea8bd1b593f07d828200bea5c29d24f1de80beee2c3
zaf9c972445e0f35bc106e8025479333056dd72999ba1ae29f9ee81b759fcdeaf6da30e22f5ac86
z115d637f24716ad612d8bafd8c6e725aab6c26d65107fd0855079a400c21fd3990f5dd9f9b7de6
z76f2176e9cbe42fa92a8dfad90b0d17da785c4a09136674cd9c9be67969691dd9ff823fa3e3ab8
z785bd68a42827c1c9d7a3fa2b5640cbcbf912fb35cd63353bbf45db36609b2cb8ef37e0e2113f2
z35e69f33c1846f05a3f4472a02c228cdaf2a8465f1a15320910d4229801d83939fe0886352ab3c
zda39d26a05ef551afdef38c39039a356103703f8808981fff238cf365d2e14844820ead9afc528
ze7de2d7bb5f85bb10d9a64584896c4ed23b1d7b1962804571113abc08bb33b00798cb298df35d6
z529533e1cb77edc850436ea3f1e0a176a365f9ee1328c61f4c08232f99b6297bac96d4c6895002
zd61f597a0c5b5b6bde6fe5776c34e652fb38018bdee4e0be5c5ad5b180ba366c8f7892883a00fb
zf81fca3f1b05aab0b2374574381d80607dc518d27b2081585fbb2f13d60000044dd88ed305a86a
zcc06d28e28742d38d0b41a5a4291558775c31d389dc4ba7e94477cbb2f478d72c4e87152f58da2
z76f02da401c13ca89aea510a8ec1419af8245d463770638c65f893701623d0de6a7dbb6969fb4d
z8ae0136fe75cf9dc7dacbb10d6d592ba23669f8b9d47d7cc0c7f4beddd2f17b3d124a920965821
zfeee3d3fa045fd351475cd625a5d8474dc6736f827a955dbcb9aee6a478a44f9a67078497ad91f
z929d00a89be49279424714190a9496ccf6f6cad76fa67e0c8c68f2094dba7d2149867aa1857eba
z9ded56bc0c1b23abe003510a1308a62d71cc0b8fc53c93a15675f3045a73deb729f774190e144c
z0e3609f2dd5084d19bfd6a90c959ee870629c22caa2df8d9fa86231c9f2f9cd6652084dda94c5c
ze0ad55a0b0d59ac7658d434a17a57766f3fe75b15b6c06a161814c0015eb727b8851a4120555da
z145cefa0eea02ab46eec32ad1e334f5bc8195cbf98182d9bf4e4241569c70dd475439e8fdac161
z35a8c8b2f90e3fa583da1e3736cfee24ced08954d786fb6791c55768de422b4e13d04635c9c581
z1f4e06c5264694799b594641991e6efe8771830cee59f8e528cb76f12d0656eb3d9e1ed4147f5f
z3793c010cd11c9137124bad367de06f533210514ef606df1c62bd9073e02bce1942948d0731216
zfc2f6f7ea200db272f32c89752e24d629a53bcf339accf58d71b9fd921fa18285f74f183988617
z2f5b17d4633e40608c61ac1e53f60966ac30da4fcfdf9e14c9be10b5c40aacd8bf1a1320114b5a
zc1e5d1fff267b01d20a24232c3f05f6efc89d5c11d046a345b0fdcc8a876669004cdf94e8fa6d6
zc106c681155b2ef2a510b0e5812001230e97d628fe1e997762ce6863a9c48d407c5ac35094c1a3
zdbec8a3877e8a370ef1745968aaadd0a0ec76cdaf9a5518a7ec40b753d8a6eaaa5b49f452a312c
z61fbb187c899c936f1d92667c2a789fc66ba43463809a73e43371cc83b314004d51f9d6059ec3b
z5de77039fa199582efd97ab1703e087e304e61eb146ccaf7a137ab3894620d22111f6b6c9451ae
z92a7a94f4d80b39f83478d4ddac7983a0fa9db75e0eb6b6f8dbec12133ec2f13999ed34172296c
z21c023455e5fbe427b142926de0ba0845399025ba2dfed045d17b451b0ad0810d29ba635614bbf
zbfcc330d601eef5f82440fd41d77e3d198cc19beeb0bd380cd0502805989874a93a9991fe38648
zcd5e1c29ea50cc59ae365e3934e05e7030dc85cd62a6fbd8e0a252fad72fe41afa9facdc07dd00
zdbc0cd07d147d4d1b6955c65762eb62c66855ecb02ff7a7455faa9314e3b98f5e44f4c0a772212
z0877e77aeede921791b3738ee2edeb2188d07c571b7390477ad1763290814c3a3e616fbbf1150c
z1277156a388524ce2b8ed2852d24f0d20bb888bb6d041be0e169713b6ebefb9bf8a04c71308104
z9f7e1e0b84270c7dbc150d6d426fe2095416752c32dbb5e23dcff5a6031d855c8d149ea0df5695
zb1ae5e6decba8b4ac3210d5a7c93f1a56590d9877f1ad87a70e9adb1a0dd7bcdf06707d1e06c31
z64dd1ee2d803ca176cb1312d23973b3926bf71b68a9d63d7dc1a2b52994b8920c8be59ff4cde7a
z167433aca28d6f83d3b1289cc3184255e876b1d344e34055dacad921aa39516e73f3be1f2589d1
zd1b4ebdd3d8da9f04d0fcfde3faa18c7e7f6d71a82de409a70dd9c60faa5c33d9a06b4552111b4
zd03f3226b9044a626499db0727aa877e80088a9328ecd6e3436400e88233bb141670c8c8f64dc3
zcb8ba6120a6c5be4cabaddb1af88f3eb57a5614548610790b3391b728f734895c20a39e4e7f72d
zdd7002dad026ae2915e1bbe650368971cd1e93f17bdd6ae0bad4a00ce0db7bc290aede4fb13d5b
zc36dd7cb6317be42fecbb271e478777d3836739452aa69a197bdc24d3942248f15448f70fb0c7a
z2234869d9bba18805dafd8a757ff6bbf8b09acee231e9c5e8df06cd79ee2e6fd8e7e815bec9742
z10812b9176a017164b96e5606fa2a795ba1e6c7b4ca44b18a8f1a782863264e29cff25c4cc2d4a
z9c86440cd0f63d3571e8c6de195cd5ff84a755d3b4feed5a8b9dfaa7de44349b90436749c58d16
za3bc2591006d10bfea709a863229ec7a04f97e7ce825d671ae6197497529fabf2627559c3d8972
z656926bd9ff24be618d37b1faf0ad2bb7d1ac1346efb84b56f5f567c28a923f98f031e14931fb5
za74726db14a6230b98adc17581421d8c4cc2083d2e3436c8172461193fe41ddc821c79475cbac6
z42254979d6c1e5d40f15035f81c7c697cca932204bec47facf388a8dbd3ac22ddcd4ba6c486ab2
z7b4547ac89a4b32d19424c00e59135567a642e24d93828ab52b968ed7b0a9c6854f0d5af7a7a73
z6fb244c4c87975d0f7aa29508e85a9c8d59cef7ea8d4838f2119b89849e377393c7de343b91413
z656e29d7fabfbff8494bbd5ce5730bd19f4d433e90d39e21aec666b672d0fdd27f6316e4fc3657
z2357f31ba2355f0816114d6ff39c1620b07bfaa3af6be668fdbf44d1b1db171a69eba7a9fbd89e
ze29546a1461513e125572f7bb3b72547eb5a3459978b2060d8d422c50ab4205b8b9123124d664a
zcac1ac317c33d4933ca841af0988fdb9adaad52031ba6145cb537ec155c97653120137a18f968e
z6cb24280828ac0421f395d5bdf01832a9199b5b96f76082c253c81f1b7293a790476066b0b37c2
z1a9742ab19bc3e4102c927eaeb767cc27f961eee1a0fd0f17ea0a3ec815c6b6d1daf4572ebf068
z10eeef912641ef8b9fe12d980b42c0e4dee2030ae41dfa9c985f0d73e211739057c779698f0289
ze281925dcbf76ccda52d8319f2fa3495fef36a403e8f4a6959cad86cfb723ede0956a35ace99fb
z995c7fd33742950b522f89b39254681be17b9a629124ec465a220fdb6e2c302ac14861e40a115b
z8ff9039ec24be94a2e36c92dc87ba904089b9458e1186f049b326e4c8f4050bd67c2041e180634
z1c369294637debcf6163540509b26c2a08171a9291d7eacfd68035c9f97642d89e7d555f375a04
z1687d5698568dd48a442ea9be2332d196bb5423270e5a570045a32be1d3f03675bec33ae7d2909
z009ae905254ab3e2fcae333eef1895b6db22f115116ad2db1e7b6f7c5eaa2681996b0d122c684a
z490d49c9f665c787f2e153f7268e1ab91af06a9d4ffc8abc73f6a66516fd0832921e7dc32ab759
z4067e952322076a0cd622ed6e88ca94ba2b29d3fcfece2bcc8b1da0d325530321e46b833d9a75a
z827f402e68d44133c01a82a05b5ef1b4e3329579db630764d23b79be4e6f2658b5d6cfdd636e30
z3241361175b0250f1bba4d1194b2f24918024cdad729da9da3b23686acbb5a242fab25fd16cedb
zc537cb36c79f0437b862699e092144ca981723b04ff39f3d2ff8a2e4c451159e28f750b52cff86
ze587dc6d74c3892d508cec63a74f521af2ddd402eb192c6074f5ba93f53395bdf460e5e27dcf8a
z342bf61dc1ea348a384ec5f4a8a128484c4b4cb63a58cbbe2513fb48ea9e191b45052c07c350b1
z6e336facb56f9f2a17a5315d909fc7c96e4697af26ceea5e050b464d15517d63a493713e9c03ef
zc9b1bcfee00e9d6e9c24fafc2268afda642ab4b412d715b43fa31e8b20e44d010f74b1f8702784
z713972878b46bcde7bb9db3747eb622f9eb3fa85dcd4ccdefa92224aef9ee247781ee1884d0a85
z49598be976ced8b0dc5ad31c8c07ab3167dadaa3f8f65023623560a822f77fcf69cdbaddd74419
z14dbffed3d1881507cdb934db9fe7bd16fed54ca38a6bc6fe577c229c340b2f8319939dfa42230
z2cb84272f9fe4e5f980b66c67d866f316921b28619dcd8cb805e1959f154a9130453d8b9a37f46
z9e50181641139cfb9818b20387a4007f5b73f23222638f394f0cb31628ac950613d262e28cc84d
zfc7dcfa1dae64106669158f9c976bc6fedf5abc2814760e878434073588266648387bca6770472
za9849fe3648b90f6080e44548d32db131f66f8ed7970f99a705ff76d343fd5dd778c5c3a0f66f5
zbcf91d5bc4d87ed26863ae3ac9ba3bcbad2fa915760767024ab087ba234edafc3862a17aeeacb9
z20aee05a17740b884f050057127b9168a7f356b580dbcf87be90838785d323983cd19ac50cdae2
z633b239c4b4188bbe1a8a1ad53344269218aaa597055bbf0b914f248287ef0eedcfc60d4131af4
z0dde32864f5506d4a21c4fe683ef8f34fd4b68cafa6183bca751e6d2de768c8bcc3978f967292b
zeca28147a47d0639839919c1327e11db7681e42e70e64e51ec2d25699f33fdaefeab2e107cc933
z637efca8ab1e2b0f83a987978290e88f5944a9d7791603f66ca1b32a52602e2352d86d2f5344f3
z95ed04a25f4300f5d3d91461cb2414ba48999ea4a3403272cd266d46b57b75685b685ec14dc025
zd777da063259c0eef2ce5560c16d175b9ecfd89a1e5bd1483bbe7eeb117b8fd39f5f47c9688bd5
zae99d41f5b357dc78994bf32aa2f960314dc467a80b5e90d62c6f185f86563224634db5f9bb7b9
z7596918f272da9d3141d4f682f9173075ee8d9c62f5810f658bc2b96f43873e1741b823e296f27
z19e43ed1396238ff78e1b431811f24684e1ced3b4615feae937e6e481acb13a85b2bb0ac3d8e2e
z6c4509aa34e417eac693cd00595ce4d8b2bb2f9c5125c91d358b2222cd3f9ca8cee5f154cc00b7
z3bf25aae8d7eb693e4c4642a557f5c797df8b1d604af661711ade0c6dd4f49a86a9a05fdd12e80
z83eae377308325174f84b45554e6d36b9fc0a512defbfec78907d4a28a35359b907a1dbdde243d
z227e677af138119d98a5755cfd632e46b450418e97b2a16f82d9442a19346b9cfb2358719bfed7
z0fc0cb9c76fbba5e47c073d31db0c22b08aad2c02e51d2be4b9de014af5f8addd718130d9764eb
z034f0597a97dd2bcb926e38b999b226af7a2956e303980e047ba74abcbbfac2ffde626ba90f3f1
za0e18da6e8fddc8c352c7fa072f255d7959ae7471e1a0dd68f1dbc8c16c33f427b0e6aeefe1d17
z3224af4564bbfd770791641573a85d028f580e236a96e9fdf1d3d144a2c70b12ca524efd5d1081
z1eea4d7fb3d2fc1069c67ed64790041fdb19aa0613f68c984b4c441d9eb7e451cd0d46310ef772
z8a00851d051f32dd41223ea706b8bd31f85fd9149c0fbcb9400a25978d5b86bc289a94ad012e86
z644ba835c48fa81f7de58c776ec691bf39a90a8afe1b4034c98309ed1cdad8f0f568a15394c468
zf047766ab7fcb6f1495cf953e197ec49c7ab5fb0d6a3c4f33be291095d92d0d039f125245c91cc
za091db1ebc0666cf5dd844bfba9f502ef030d71bdf6246d960f3e5f90a216717453d54467c1de6
z1d10a9bb00b6b31d19c88ce3a8043470e0b96b79d59c0643724d8f82b11474a75e60c2a1c89fb8
z49b3b0593d50b15edab8bd2b8d130b11172abcda87aa2693c98b1f95a1efefa21f4850ad29a450
zf8aca568296723f6f43bd193059fd3c04c123c53a870217cd0747cff56689264978d0bb2316144
zfb0944e4d81fa2235e4d851adc1d1f93d5ca09e9baa4d6f08e3a7697fb2a8b61432af320eb42b6
zcf1197b0e9d55fe53cd492a00f92b08e7352f503cc9bacacd37ee12a79959b696dfb8d8c798982
zcddca4a490051128125642d0ad428c949a7bfa001e13e8795d0a99b477f31d69c3194a90ece1db
zeb02f7be4e25bed60b7eb1bd5e4bf3a5bbd1074b3862c096425677a7c80c9979315be0d748f10e
z398ab21915038f7f1dd2923527c337cd5e31ce7ab27a3ee6cc7017e4faa5a6d22274bce2d72e93
zbeb4870c8001a51708038294f63236987ada0cf7fd2559a13f29c08bd4c8453a6c8bf5e1a6350d
z3c50059f409d457ade2c708927f7316ce683936838654d2e15eb3ae6881aec8c9fa81b0c5b2723
z7d1c2bab47be17ab77b5d2b06fd8c6b7e67922a0995aab941fd30855e300c8e3b4079d1af22765
z943ca9384af5c34f91e4fe51c2eaae658a4a1a362ad1c889c1a4c39861c658c0e935b58344dcdc
z4b0e1f16cc3ea91e1e853f55f8f5687332f90b30fca1fffad37eb5007f1f180a8a969c4d4663e5
zcc8b4b905a10860a2501abb5bc4a80905cff1ac8919f414c9257276012dc4d55163900fe6be2ef
z9dfc60cee4c8cb56d51e0509baa72456a135394f22d0cb78e83e49823481f516e33942aa4aa635
z24dac9fd1c473b1cf3ad36e0a762946d06dc73217a5f21f1cfa7693d8f7bba7fe61558bf485dbb
z71762de11a79e8c611a1037b2943342f5f39fed65403a346ae1d4622929d4104e509aaf4b750d7
z586e11e88c152380d8421d266fc91284f09ffb2cb968a6931b646de42adb1d1d9f017339bb001f
z82d04defb2959e0daf49a33f14f51a6be42c666a1c41fa876f4294b07503395e07cb6f4ac8f681
z52401f107cf843a6204cba3d9495aa985645a4f4ff47831b67da76866bb9e38c51660c677765e5
z9694e95eed2c3acd1c80e07db12a05f1529c123a7afbc5f201c2ff11bb09163c719ed0fd2960e8
zdd62370c14e2a1015265dd50daa6130822111902e1eb355557781d0597906e82e8b71edaea66c5
z2ae5d0d7671605a3b287a5b3664a872cf4d1d5dedf1713f2cfc979719cda51de2b925b8da05e78
z7160e33713e5798882c0fffe4a0f8722de8ddcd0d79b0a3ba29fd1c09ed13141e85b1bb3897eb6
z28aa1c1fa08604d2a539675c1230308b879ee8c4bb481577d12eae1f541b31583fdeace7f09565
z4deeb102e70cc0cf43f0995527f83552d3bc9d8234c8d1a709830f1968ab8c9ddce7855a6fabef
ze7ec564b1516692428be4a1ba429a9baf396d47f2b4f9be072099be38a92ae3e53e80dce60827c
z13ab00b054569b3de6f722e22a5fff66189bcbb8b292bf4fa144fb7b3d70e81b9160e367ab2493
z37f97dbdce638461f6c663ba3677b9ce7252e391e8b497ccf6caa7f61e15f2eb7acce6ebc93af3
z102b569a6696875eaa83b4ee0c6c4c1a82b21a361a56442b03f5968a9604b639100a2e2e138027
zc04d9dec0c3312c4c7930504bd1ae418b0833be51a81e9fba9c3542b61111747805dc827bca181
z7e27195b96901525b3c73f18ef84e4e7f772bc633f3010cd7af7254050a881275b995a72edea9e
zc210a416c4892240ddcee6f15e8bc3bd4ba6b896bc8078c4b039b02253a280c59a24a57011cc2d
zc16593456c82e5733cbbd6ca0fad22f1223fc6fdade497a1e1132f3174da9623471a8f20a11e23
zaec662cc36b4a730d0d255ede018f1491e1f8b310c8bc58cb775ebd12a0a56153821c251062d93
z1a65fea9199213af6f17ff3ea5bac949795207b95e267c91e5371123ff2a2c39c87f754bda946b
zecdab437b28955abc5bcbe8ce407fa08dc78a078d2dd9c6822ae4d0a1329b4d1fd4e83c3243a69
z2d278d1f6aa9a6eb9b175a05065a1925d3cff7853e630c50b7fd7e45fee6046d711a7728ee39ba
z98e78fd42b57469f3ddafdb2c12c553d12a384e5e58e358326c3cd6343acc0f1347c9d72bc4b55
ze704b08337647460c9282e7f2651c0595304b41c2d76ccc3f8b83b7afb903362579db32de6a052
zf0c85182766252a2e99860938b8a5ea3e5d8e89b5b996f566b55f143382003f11f42ad941b82c6
z7157778a310caf960bdb254bd2642c4909354fe345748f8d668597141a8077e2a85246ae85f9d7
ze57c21bf14ad705ead04f3e562a84e95a25db2bd775ef86dc427140f0eb22baa4908fc00aa8f8d
z84228a99c578d05aa8e191675106e57ebcab4b96d0f701b479331aa0fe35ccbd213d79a053c569
z0ab0f6c9132b01ea50cf9b5b5ea68a44ede42206a9bf770d89fc0072d4603417a4430dc23e4665
zd8d8d50513d3e8047aac11dfd9be7edd81b40341d2e52d14c9952d6517f49e8a46b76a826fe05f
z0d8d3a7586fe404130c3cb785564194015f790f7730c2646dbe58cee2a473425c184f4165a2acc
z84af89e76012cb2a9338a652f19a667f84f10aeb78bea115563a7db01df81d7bb0bbe0a252e393
zcfb4b179879c0a5bdcbb1f3c20cc06cdcdec9f0b8fea2c3ac2a710b49a72efc8e8bc2422769539
zf06c0a20993056fd787fa5c4da9a495ddff01ee8593095f6a56d2845d6b37c5995f05cc8e3782b
z4ece31b7668df523be29d2837d0dc2c76005947460a4fb4b878656cb3b8c7df0086831228ed8a4
z5f9ccf497427ecfd0fd5b751e59d035059c0f26440930a2fcc554eeb7e9148526acd844ee988fc
z329011eeed4871a908b709bc5750afe6d665aac3ccd2afd3969fc9598725f8a7fd0920b3313a36
z1205cc0c948b9205e53ce74cad0526878c58424cba0cea0297c7cd2624619843ac173e8496e971
zd7fd2ee816ee3b1a38dc7b2cd50197e3f2b8c06bd4a1669fdf07705497f41cf26e011da7fa5705
zb5e4291d9a02501e2a55062c152a0f97bb24b4b70fea925513c5b53488aec051703d78dbbd3448
z9c5ab522a287c80aa7385a7b169ca4b1c9674e59fd052e3731318ef09a1b86438f20c6567c7075
z8fae1f33fbad888abc96713224934838c20a43f1458fb79032f1621c4d8cf3d5683447824ced5b
zb17d1473f66a58815decf7c1f50dbfc3b17f738e78da6588cb28675cc81457c546e77fc60eceb2
z928309a409ec8bcd4940008e277a724db1c058621eaca2acd1b359bf192ec70e43f5d550b3cac2
z02d35d3e45ca2f02e92a542c794067a2fb23d703e021b9fc3b52ed46d2de0ea88b67e52b1a96d6
zeddb4b70d5e0ddeb09361e8e09c1d18f371db64d754a599b2f4ca84b75318a1b5ae43dbfce09ba
z35939948cc100bc395ffcff1d8e4dbbc1b48ee6195274b65abb2526886a022dc12f4e370ee7588
z95919c77f0d580e9f3ea6969f110de7bf0c327314075a5896b8344407567b00f2ab9a20d7a9c58
zf2f5261f146c455bac55b140cbf77d47ad58f6320337d48c68fd00889f7159a87d12d18fcfc569
zdda6adce497b87402dd38e9e59e5e15e6fae254e341731d9d6e1b25621b3d4131c87e2e0e4e035
z971406918c85d745dae0ea54f18a4cd4926f535dadcaf315fb3a087d6b52c95b0866ccf47ef0eb
z9678aed8c86db1e649c50796c1006471c6327d66878debf4bb0f860efadf6f433fad4ad2efc633
z7094bb52057b5a5458481868ea258ccc0e01b7ecf77b610cac9303af5f6df79e08099061c08fba
z7d382f1a27f861b4cad283c1d1eacc774fb3fd932fca29314f69c4f684b0a5dd6d777d5a7762cb
z249aafd0ffb2ca29c0af040e8f9e23fc5ceffb8f103d41e8fef38e5d88a30f405dbf983dbab99a
z94d22cd5918d2cbefa20d3c6ce82d600b8edddcad8ecf78ce675e8eb574ab207aed4cc2c3cb31f
z93a64d60bdecad87dbe0bc00881bb71fc4388adbad05dfad62f4c9c6cdbb10b121260bd21d32ac
zb936349fbf98438d8f3ac342b584162bdcd40d56baf8b3fe25136530c0d2d0e6d60ea0e2ac277d
z8a4207e892fce131206a0b5423b059a1d25c93b27a6afe7e3d4a794837c5dacff4af788807bb69
z41b01819bb6f09a67a8b6fb10b27b07e6773e1522438482a56199f013cefb18170f17b983a1f45
z3c22b59cd54cee3cb46e80eca997a9f237ab8a582821e05e2803d54cfffd175b27d0d68723c86c
z4d6e90d2d317b380d13513a5d3a8fc8bbe24fdbac90e1c628e9a9892b65a656af77d41f26cf99d
z1387d554345dd1f0fb766b94f7e81af2100da90d2dd48a2138626de11638a508e1221f45f2697d
zdd0907f9ce1532327a01720e12e9a95641ea429f1391fa91dc537f01b3c764ff7c08c5772560a2
z01c9823b46400b47ced3396a048bc3812642c1152b5570c96fbc99ca421899c1c355a4eb2132cd
z3808c6a1cfc4af87f6cbfebe6a83a21da844a2ecf125307cb4753a1e07f14ed1f268c44786d9af
zdfe8299cdf43c75904520d7d443a6e27bf85dc0d53670c8a2bc1456811268225ea024ad3eed012
zca876d61f3c773710f2bb8b8c1e46f72ee4d02fbf78a85ba35974fad31b706cdc9eae71c4e3244
z51c608ef8e8502e79a4ddbfcccf5dd32c8ed8010aead425c75159eea6ad3c6abc5dbb67d222b47
z4d26abe6f736d5c35143a7f23f7227c6b42e730fa7f391b9f9019d724bd318fd113340a45fe7eb
ze7632237f2926472cf75d9560c810a6c1968aa3a99e053e45489235e8379f566b8596a9803b521
zb96021f12524ab8dcb4430594711a931e99f6f6450ad61ca7839dff7fee427a37c6c2d88874539
z1e3ae3272cc78058a9a329a5494ccf57b6cf3e7103f436cc8f62db77eaf099cdc9aab108f239b5
zb4ef99312f2f6027e2b97f70554a52bc8d027a318346512bad228a0017702256607399e7af3117
z55a199c93d10c5c03787f168bd9471c2e8ffcebbbd2e915d506b2d9e1367e0af656f0c4f13a4bb
z1639f9250b268e6fc96a53768aa37eacbd0176f1c674e703c2e68fbba164cc1e9b2b39958945d1
z4ebd8f275bbbbc0aa871b3750fb9e84b46145ae958ff7b8b4ed78af6ec14c95f0d33063362b12a
z11f03a878ebeef937bf89afb1258e926d9ca703ca15546ca3ce73b9ee08e6633534a2f237e0e0a
z659f4fa809a7c082bf8c975f9caaf553ff852f8d3c0264faf876dc99da0010079c118f7eea7fb1
z527f525482a7a25ac3f58402914dc302de0b690221984fe6f68214f21a04b21941b6703fe623ae
z4c1c6219dc2daebab73bab02e76aa33c90ea69d901687d0dfd7f80c6ca0f8b579c36fdfe812351
zd3e7e7d40962e98481d5d7e69f80b2bc302fe4a68b5aa5ef26fcaa398e150e0c0044f570aba773
z61beafb32cdc075627a943b5e9fb99161ec19a01bbc3829da53ddde13eb5438e730845cb543429
z6b7e1d6f8fd7cdffaea71434de8f649d989b87bed4b9cfb8a49e94a612ae60174a8a05d5358eb0
zf3a5ff7d74db586d43404ab2c1bc01139ed946f7f5e4df7cada51bd442886d66ed2d3e9135daab
z6ab5da625d3604bd6c6113f941360b629f79d38626686e62f5a1240a61570be28ba7ccb4921231
z56e4b29c76b5bc06c45217d2b77c54b6f7aa2b451134ae63aff47bba86b99e7731e8471115c245
za40a4d73ce77675ceb3310413f7366cf1c0e1c4e88e909ce7be68565cb3bdfd6235ca9e2b8ec90
zc054a9f9a6b0c3fa6a906369234c1499ed38990e6cb80759ddf2e779c305ebd86d26ceabe8e435
z940530ad3535fb55ce3616286caeeab40e863a1839526ddd7b79362f032b8e2850a6541e273a28
z25ea982dabee868ef93cca2d0cda12c090f39d2affe39bf5abded34c51d66e57b951f9d3c6194a
zc9da15122e36d21a1d7e9c214fa9d2c837689dd233ace153918a4b4dd8a13a5dcf358451000d36
z98fa577481545bdc05526c61c35fa7909b627e91a52658b54cd79aaa794699b9fce48ab598c1a2
z478ae4f8dcf17640c217e05ad0388b8ec464093b6cbff34c52594fd61e5bd393eddc29e9f1e5fe
z94a0d317135e57304bfe0ba7f2f3fa49b600da605d5aee2140ea81a69f8555f55ebb7c5eb575e8
z6e81f99ced8785e9c09d61e2a29e709b2227d6cc33dcbbc6b91b4b95b12c82ccbc41c05caa3f37
zc2b4144d1409e737d9a1a2322123c64dee22d5d4f092f5bcf5c5c3f7e06b9280cc45cab1ab198a
z02d155108e8d4ed10155481afbde1f0c7e138e6f05c4eee5fb07094e860be43170358143fda838
z284c6e55f805b146ffa89f71ecca7630ea9d9b62d66c6392853fdf9641a35445291e2732850625
z5222ed312bb974bbec6f5f9cdacabf7fec6bb414b7313c0e537b666fef3c21d40db3b809aeb3aa
zc5d97dd807b2ea5aca11a558459808bf0e1c1c11c4c68fa13f2501af285a2eeacdbe035d1d1af3
z6fbbf6caf4fb357fa4867121336b3d9eec0af71dc24f4a4ad5ec5adf2b232853f8ca48ac9602fa
z6850e445afc1143f72f535bebe344b3876b51de60d114abc868565a31126813ce472698dfd7a69
zaa4371b92c3485f9298265892210a1034813ba6bd2676616500c071fdb079309c966301caba867
z7f8e2170578a9e2cefe3a6e6e8de6f0669cc9effec1ef604599f5e5c4a99877aac6d9e69ffdd92
z53335ca06c2255befb34cf2e83d74f4027aa244ab2af9d831ad52daaa63105151acc8dd7f30dd6
ze1e5e34ba1ec991a8894d231d0897b9a3c99d05d78831517f6061e6aa266875526660108f14f0e
zf03a87cdb4bf20ca8550cd5faf2e4be056bf18fb3b0eb0f344cbe1ae7d7da5f719e34366acccec
z745acfbd0cbfc407bac873c75af063898fd907cfc8ba9fbce184768498b1bfd40b2989f3f4f5c2
z96e6ff4550818515804bd9ed800f8247cc0e60f83ddf7bf85d42db913f60740bb1882e7112376e
z98c7d752048a535712d52c2ee8ee3664c0a286989760ac955fdaa46ee9a4755ba02fd221109d0e
z2088e972ad09137c772dfbfcab1494917693340f33d7e94059ce24f8e83b49e91bf88c50d4c343
zdf1cb5a960d458d6a8079d8a71287ae8655d994a989182bb9e9b4428c5f73d9306defde51c8707
z19bc1df785b8a8bacbb94774442606a5632fb7cbec27ad875510857430d09e514f56de1468d8a7
z77744ed8cb94d7c0a3b815a5f5bb835bebe51c08ce19a78a6d67114527f423169548a9a998f45d
zd5e684a22db7481228aafa5b8280c58b5eac173c51d95562b16d3ca059833121686248a0295825
zf1ea9a696cc031fc1a6d102afbad0425732c4a1f485488d00cefc9ba14f7cb6873196580436b7a
z7fb7f8e702ff5475d2076e59253369fd82dd29adf1f47a03a71a4d3f47ed1d40eee217c0444103
z15bbaaf6fef0a0177626ef09ec97195128b94012ce9b3afa0079b0c0585d0ba50a828154a12469
z3c5e1dc8c378b4a95c4898bd0fefcc1b1bad29fd25d128a1f0bcbe3dffea6b1c9f8e1929cd2f85
z430cdf55560edc69fdb109c4d4410824024b52d6924611514cea71a9230e51c1c2b350520e59b4
z4ec7fc18f35232fbac559a9aada07ca13272ffef1b94415b01afbf14d114d6c5adb7890ea81e7f
z57d48991dd9a8797da4d6702792df468dfd379f264ce2c6bad8c7f0c9e319c0298fc7c0adef4b9
z31746991d7a5d56380cdd44f905da7162f7573175996e01b170143da1ee4a7e796d754783f0531
z8e0c3ae7a7a47d1b70ff83fea4939f85057c68a28edc58d7ecfbf1eebf22477b6daf2b73093275
ze540e14d32795541588ffaca7aace0020427c08af42dcb8be9a3209a8085e9b91da44f42043f19
z1c7f190210eb37097c2b4432b41e5d453b2efa0b0bc250d90c01bce0a60d801593f9b09ce2a4b2
zf80b22d122fdb7ecf9bcf89d6122a477d69a78eead8b01dc57014354134d9ca5d3744c68901e91
zf774e39bc799ae70b1d6658e34fbd71356f0bcba1b728fab3e78e8cfb01161c66b3498c3c01d6d
z2b2212ca0f870148fd4fa15e6becd1efe50540b49225f1fc9a3802e6d0227cfbcfe7cdecdeec54
z412afa2ed934bbd17a11125d2772f422e272c8441f84a521416a0b8b6f8dba311631bce973264f
z673c71f763312aaf88ec9d1a48027dc9ce2596d0fed5543e41d1e15b7e77b00d4732841521b84b
za43029d4b3e947684062e96d968ff31c6d479a830562c1aa910f14f06d45d9f4cedfee2c8dbc28
z1a343ed8c9962dca18f2618e1351a96076ecae2d5fbe044f6e7854bd23c4822c04e50e5b5601a6
z09b5fbd05c0618ef93814df56ca424f769fbea9d51982a47b231713a81e449a1777e71b24a1b87
za138a7fd2dff60ab66249f51beb0dfb7875ea00e22da09fc40ef5d81a0512862e7b318afcb91eb
ze721c7a01e864410fef8503f7bf3c6ae9197ceabc69a2dff9dfe67527cd65a1e8f7f893669c4c2
zda6031e25255d6a2a2f7073806479493a22e8bda06c1e07cc35778d7d32d0ca0507e45a23d84de
ze1a39a5d89e40278c14fd74c49197123c1abd1f3f0b99d871031f4259a28a7fd7a525e141c3986
zcbe2af37dca2deacdbc483fd86c4424cb158d8c4967d78a963efba7d1ef9e16763b62643fb7e76
z8e30e25846064a131b74eb98af2c4611fc14cca0d6809d1258b517b68277fff503294cd04f8043
z5b5091189d478d7fbd63d857c13774f4870fea344cf0784f53d9d6f3e8fbd46de18cb5932ecabe
z14ccf35e94c7be07f6c8e95d2d18a1585f88c93edadc926ce75a93ca5eff628bb00537fb7380eb
z8cbf45193944652c7b998fd3f40acf26a99b8d052278c1ac494f2d8054e8efbd00cbcc049d92c1
zf2597ccc82e8c8febd78947b887508f4fe51847729e2788d80d9cb8ff7500af76e8b147474c3e8
z31b8ae24b8679960fb68706471b6ad97aed023eb0e2ebc888e8e7bae7240f80efa1283b360fbd1
z64d3ad705a5d4b0243bc64a2fffda2c3d72ba8a2cd060a4170e0e1c40ec02ac5cafee3406affb1
zbdd078bcd3eac2b6a749b99828888d4c72df2f0f680249ce48b84dbfa224d2c131b2f8e26eaf92
zd32ca621cb99a708c2033c0df1e5efb6873d26a1fec6310385114d2bcc4aab130ff5caa0226205
zbacc1c33f6bb3f4b22473486565b2c5b5164fa805d7e2c3525352f55a54cad6afe4f850d377d21
zbe87f0f8e0db529a139cd8ecf764fbe3ac2a67ae00b620e5b5e51c886fb4e530d4b6e690a9f7a3
z137c280ce7b58f39d418be2a11555a9ea809ca21f6fdfdc361f7a3c2144db157521b3ac32deda8
z2e4b1f356a4bef7895a9f714f09d94fcd7ec8c8db0c558081964a165365a78d1d3326ccf9f9e9a
z32e5a9b396020b4c84fec6c0ffb4bf639115b48615f880f8380d39736625f0d77be6ff190b7541
z674afacd33463f222be3264deaf7781a23e72ed7d5223d07d953b3b2e5e10a5ffd80f84deb4248
z6bec405b4f90f11e9bac6eb6b6307f74b5d3284fbdad7c68f0cd430ef3f63e16f37ce2c976bc14
z3efe5f26b91417ffad16f932d34ebee7de82119bfada18bdee0dae1526406b4e6c4076e27da8e7
z3b28f6e22d87c1c2b0653da83bb5bd27420080e98bc1121c32340fedd86fd49ea8fe5a13d46b6c
zb6d7581b10b9b0f6eb70297f3178310a15c2a6fa4fe484f22d4d054e819e7be1d97356ed529094
zc448cbc915bd1002127169573e50a8c76c55ce60f5fb8ec3d556ae9b66a6c373f5487af9886f8b
zb0c78f6d8534faa8704037fe3323ed34f5ad309a316c9e881d67c8653242d725b002ade94cae86
zca1c8cbba0ffdc2e2a0f882babcbeff4b32ee3706433438570b2adc9357cbb06165ccd0dd2fade
z14c7c3a1295b470cc452176c380647a810c4752345149f1ff62990e891d880f25db70f0ca2e3e2
zb2be81c98b48bb1e6cb5fac4cca35c39fd16a52b669e9a77eb971ee1560844dc8ba606f1bf3cd3
z64c4fb845a7c4445e081b865e81862ae9e8270bdf61de5cefbbb263dfbe7d17c416a3e19daf5b1
z4cc910626dd95740598ba5c984abfb964dc77cdf4903a2a7ea92f920c7dd146d376998b884d52c
z3aa2fa3733b8008bb4a13ed52b312b53710e34f7cfe5d4f2b7827c0b19193ac4eb38afcd980717
ze5de80c1eda9484e82f51b5e57307b90757090723bebf03e9fb179a44185ff61266be0427d3623
z640c3a7b1e405b74bb393cae801b42f1146bb5b9a0ed84c51b6e5205a55831c58b2f274bfa98b5
z9d6603fe372ae265f0b26ee122b97cb50675172f30598f97aa1bfb20508b8780443e34c508a23f
z02817fb2f6f471012cba1b7f42b3a4426b7318211f3a8f64d232065d4b550bf72b00328dad485f
z728c6196516d741b42fd69b0e70e4321cd3ea267187e54d10d8f0d7ee0028cab64f4290cd3e48d
z694a7aa03df6a0fad6950e26e4090018983aac232bd24ec579d38e32aa33bf4d8d16d97965f150
z5e06305761ca179cbfae2e04a7e0296eac176dc902ac73c9a54ca3e5a791d0ed5940cf2a811ef8
z7a5c63413954aac5ed9d1467930a7e82cafe120587a128f1b92e06030986e1a22a6955b2c0fb1d
zb342571ce6332d66448ab9b6a6872b4e617c14d9ec8f0ffef47e9571c4344af20d7794cdb9b31e
z6b5cd9d518b26a157d206dade535471e4e7269a310d7a2f861dea6b73d75164b44718b367c8408
z8211320ea2af1ee1581fbd21089829d35d49d70aa8f48fec0c6eb602dac325acd397b4f89fc91c
z2fee96949bc8b0f9b1413a748444b33568d4ab0b0a0954624b3d6ea9078625f7bf42ab040768a2
z0ff141ce42d787ec4dc6eb5f58c4b39569d9ab3f222789361a75d37b37a21654df71bf3957f404
zfb05c193c5e0f4c9f58293d2da27767e00514cc1dd580a994d22533c0c999338d9d24076caeb7a
z8a579616b8503c3be67c90f33c2bc063b1e056437eff6b9beccedf9125b7fadab7bb0dc370b9ba
z145518349b17d7d37dc39e87a3fcc655f82541b1f16694b7f1ceebd5156dffd5008fc6c1fb9e5e
z3070773d1492222733b5f319fa66b6265792051fb56a165918bb6d0d64b0d5c9af66d9dff2b67b
z80819bf4e11e2ee4f353fea6849fc026ba110bd5f3493a09222ae3961a771f954efda7be1f6583
z3c3e4ed53ef6e5192e109e9a4011b5eb5430dc8f4aff18340b949bae0fe02a373176f223dbaa5c
z083ac4796bc0160ab64663b75939e9db10b89e90658a2426051bf8b3191adde4fc74dc23ae92aa
z387cd22bce80e4ee839f1dc9c36193d1d66a1984aba2a0d60bf46d96d6cc5509b3584a0a5e6265
z93a669dfa5daa132bfe582871e3d4ab9577114e9298429b7268c5fdd8cbf731373128bc87b930f
zcada122a1607f9b850dc151b012a160d7e522554ac6dae71fe82e381ad37fa90477925583e3466
z97c533b5cffafb7928f6010a0364d3a27ece232d769fa3ac1df44aa12e6471aabaa3c6afdb9147
zabc916f7a4580deb4f7dfbf56569fbdb0a5b21c0934e4b101bb2d95125ef9d672e8776e4f1d051
z79285365dc2f330e46c267c021b5469a9cf7c5ecfa11d05a9be109e034e06b2959c281894b338c
zfb78a794033e890e8d8886d89f7e46959f98824221969218e7cf2fc9033f46c3cdd3b80edadcfe
z3d4556abcd055c4c8dfd139452512d1b5c6ba62e4a5fc98c905b7ae81e0c3a18b47adfa97dd45c
z5bab82611b2887f2e870e40ce44b524308e1350a6818c6ab70af52444b71c18dfa8597fe80abc6
z169f678e65c0fb8f7df6eabd355f4902139eaf7913f6cfe3e563f1b47b407aa38680c2b417e009
z8ce5ddb6f30da5f4511b161712f081e9a9a2003e01a814a1106d56801c75829c51e52bffede69e
z990fc25465527b4d65efb58c32a1ec20fd5b42f579d2de5446bf9c0a5144d90a2406f0d911f8ea
zc6acb980e2828a65434d460938fcbbe8dea646d3ea0b68fee350a1bfd54d92e09a63a31e8725eb
z86a772c5d7744306113f35da1a3a071c77977bcfee758ff4229e06a781887aea1c42b09155077d
zfac41e050f49458afec2b4e1d965a64c0537978d80c0ee71653dd02de82ee184412d1c653ed0df
z2c6c030ef8327bf80ae007d6cf61fc8d471f7046d57f416b409353ecd306c1f9330f2c90a30e83
z806de0fc001bd5ae2df89625efa2da4cb8011e12040e3142741cc3046f98dbcf33d8e6c991b510
z4cf8742ebe1b30df00221960fd7c1efd37be3d005f02e3a63abfb37a80bbd657475344db5c07a9
zdb58526ed5b3af088bc7c27eb3c3691a023fe92e854965c67f59ccfe82f3ade9bc6239a3b135fb
z7698004ea7a84466dfc4c24b4731246d7edafb02eae390a7639b4fdc765465762477240146d3bb
zf34a0796b4478d104319ff54e876509a96ff2cfe89654ea83184d8b4bf0342765b94255a71b464
z434bdabc2c53c2ab84d255cfb16a6d7d0a9b0f92c932925503087a02cd783b36ae73cb7867e91b
za7ace482a02cc70e9134a881bc2ebbeb58d002df3f3eaf08714135d83406268366775d0121fb87
ze2631ae89815d7864d65bc268fdadb04ae503233cdff15b21619e494a2ca2181319c170438a961
z22d2996121f93251d189b231453d3b0d1e256fe23d7c1475b3324eb41d18839b6e5c54387ac7d7
z5e7c610b9d6e367c959a89741f0dc99d4c574c8eb00c07b8244c7d61f9fb64fc3495eb2a76ae3b
z3578536be23589371fab8462aad658e1ddfd13ba085152f9c4ce19bb4716f5bbeb1628a16d344e
z24e471221e0c74fb8a4c3bb2892097e50bbebc33fdf0b66b31927da4058f02e8b4efa8ca0c2c45
ze2f77412df708521b33b812700cd83095010fa0f0f1ca2dc03952e510bd756e6259dd0e8fbf0b9
za63b1d46501c12f8bb94abac656caa92a0873387552ffbd9649f51ffdcd222a6a29bc85f5d3408
za7e09d0191499c8b1901dc2075c1b4519f7812816efbb12ab129d9a123c31edf1e0dc0dbda7300
zb2b965cb72bfd202c9720579f8fc56a7564f5792801f0d6baa12bb7d5ae796d0f4f56b1bf7ddeb
ze0587e6cd76862077112f75ddfc9fe5fdac257fcc9c04623b9bc11a7ec2db1c5c82df081b96571
z7cbf4163d69c92173fa04feb69d4fd0f048cc59f6d9879a5888371f159d184d50ab72774567713
z1a3d5bbc35afe3e86e8bc003db20f30309ab080bada8b2dcf49325ccf4ef0e8cebd7800a44d744
zbafb84bb62057324179b1b452a33950f38ae024af73611c514a4264ffcb8f16c34b5ada55d3eba
z47b55220d671a9f1b277c5164a68c448ceb9d19e82fd7601cdcc2768a8c60b40822ebffcae301f
z86b54e5fd4390db18bb8e325dbfc54dffe69fb0540f5668bbef911ef71d96208cd3791ae5b6887
zfe7ae7d49452ba7f525106f1327bd42ae3d51cd6fec830b2c97683bb0f36e5d5d349f9e07ff471
z85295f35222626ad35bf143fef5d4cfc5c13e0edb11d8e6d20adbba1643a6de26b37a98d2b8a5f
z6f7bb0092884e9f4ff5bc45d33db280d081b0e12a0b2da6c6b62a1f40d4c0c0fb2b6ec3462f90d
zfbd19c8bb276c5e8e5a0e5e5fb913e87efda09be0df10cc49f5f96dd4d50a80a11657a10118f83
z433c0943c4a90960a3b10908cb72092db5765c8cbe05c6727b3a21bfbd09c48b8bda77e2232655
ze896b750dbbc1e7d463c0c026d224c5b7d2223b5d9c6df633f28e21909807d51f0cec8a9c7e027
z58312d5b125797a972afef04bcf73c4fef1d83d93e285a6cfa5cf28531baa845b05936e6f9ae72
zc431ce04f7e1adab2989830044188f7b8e835df4c261dcca67c0acdd3e445d94fa733dd65b9023
z7d1c53f3bfc5346749538f0b83e1cfb8fc08d4028e182c4e6b7140b51089472b216eee1e61200f
zacbb2955f152653395378583bc15a8ba3d9eb29adf27db56e0b6aaad05c1317ec9c3ad790b1f30
ze28a73179704852b54ca58410feb5fffe8cb7f511e5af912a73cbafe1cd0633ac06651bf037300
z53c141d8bb68e66751d087c44a675896cff0449df4268284aecdce7c38aa3c2d0bf4772638d76a
zd53c6715fb07b4ddd11a883f9b75ab9dcd66ebe9c9d75b58a68a85aef53c8e2d8e171c2d470e08
zfc79dc884e61a2a195ae982f94ce301adcb7b415c53d92aa5bc970f00776094cc0751cca47715f
z4c6f08f8226c311fc6b52b247a14e5def0b784143ba9c8b3ba0ffa9f8197c7d4d1d2bacc650dcd
z6e5108e4de7a98a9039b2755254d16683c32b49765efdc9b5eed435edb93e21bf660d7ea2ddda7
z03485e0372310ecb1003e5c666d38c71efa3afcfe76e8ccdad15d00cc366b66ec36cc6a17ae676
z6a96cd336175ae56bb91fffd9dff012f1b1878f43b271c927ccda69f0d7ae9c00f7098623d22a5
zf6fe6e899777c7294bc04de0d9b0b92eaf31c2386aa24ade9bd62d9af967076c994efe4ebe04a6
zbfb6d28f7824df145fce02546b491eae8c3b9011952a4b124ce8516f31a2b9b9cee311f3e12aa0
z823c0d1749f266bfb2536c1ac34ec731593faadb23f5e6eed11319a0f7a603bdb77789c3bdbfeb
z675330014d2e9b847ceffe69ebd1cabb6e06d5f7bb5223a336f4cbebcc7cad5d9b72ee2abfcd55
z264f4c8777e9d8c807f77547132d3a8509dfc0ca575ae70000c1e27f38a14c1972b001703686b0
z4b19f89cf3bc2d42bc53f2c445542413b65b48ff3a23e7547bd15d2100bb3853d78cebf1625398
zc68248026293755935c1398f8776ba7b5749188bc6371f6789b1dd60c90380d9cf6f5792667f91
zdd966925341cd4eb99f6bd635a56eb311c2242c3473cb1cf0eb2821792938bef6e835d7d2dc84c
z41c00bacb0c0e0c4258560c2173b2577183e91475846b65f780e2288a722b3df55613373a6125c
z8a4356bdbc95ecfa8fc03a48dc77ab067f0ad13fb740bfb6529123fd2418a7e3f87b15f465f329
zaf50a424933ca0f3a2a9e906899e3053aad23c28ba49e29b185d846c6b07470d48ceeedbac5fb4
z90e7d87023459c559a8dea90c938d68db5594a14e2980c52ce1ace6bb25039b7904af8f0a44bbd
zdfbe0b5f8758639c20baeaab46e41a2f892f5c00a8f81d1b95f4b8a6aa71a9039251c7f90824a0
z02702b5cc307e539eb2cb4951b24f03643172cfe9cd98888b62aae80214ba4e603da0b3b2bd018
zb9ad22241aaa6b50d16fdd0e5df688b9896ce038fb6d7a2cb2df2084487e78170e37f84a31b3a2
z07e012972d18fbd08a98720920d497f101c622a8c66579fe5715900fdb827627ed2590a0cd7b2e
z5a99999494b524b0a9505f7395f1b216986e9ff6ad8f7a05d05903e7317e73bded3a8e418d4e47
ze2fd0c4e5f4da06bbbb7d9e3ceceb4157ffa57813936a47c8f4e8f3c99f20abc096b7fd4323fba
z6c8327c6adbf0f75a4eb71ce1ffedaf7d9bf3fee359c085d4f535201bc95a7820ac4456ac7cbab
z7be2b5e46df65ed90535d6fb1ee7f31e30aa21fcc7ede25fd4c631cdac50fbd6d9ef6dce846265
z8a10cc0a82317cee34eadf365a1b6cee8ebb329c28e293a5c5e3db428c5d5513196b85546152b4
zcbc57999ddfc7c373fbb4acad27a7526b7cede915a81a9a1b16d328800089e6715e31493e0d1f2
zc2a8be3ceb367eef6f5ee12a3f24488fc633b911c35d768b80efb58979cec118f5038e1c2f9a73
zbb77467cf2fb3be3396eb0ea951825cab418c44a4d9360cfec6583471e0e4843907885e6f9b6e8
za76570d1362c7ee82650ab788e7647ccf717b2cfc6acff821ec2e4508541fed1350d40d171da53
z9be7bf36d1207353c09a1b5ff559654b2ca0c3a1b894ab47efb5b295044b076881e1037946c802
z36bb68ba6e99e219885ba2b5c01a999bb1465506ed6c6b5766074fdec5e98f8b00d7d784d2a996
z715d06895296098fd66ce6b3544b2bc2a299bff8a24233af4066083589fac97cb1a55608b523cc
z5bc28b07db126882ac93fc50ff91c69f82780463e5e3f6a3c27b95835cc35e43d3c4948152ff93
z3eeea70bcd727681720f183657d060314e4e1b39b340055d31e9defa5f72e378a6b82caa091b6d
z8fcd13bd911a059c5a569dc446dbaeae20eb08403342c6d15ca1add97a5c22034d55c42a963bde
zb21f2d9c16d1dcf578c67014e4120f2c844db1915b8c6ae715a78231010f077b6df8097679fb53
z7c4674b018a6b1f6714639faa57ebfffcf8ae54a765ceb192bc726b1051b4cb4b3fd72ada9ca43
z03547f62d4d12930fa4a058165ec2c1c38da662a203c1d73778d82af7ad0604fc1abdd018f2278
zbcb9016e6d6de5e8eedbd4aedb770f15ce94c9127fdab4c90590ccd310b3d2530a1f8b3d1697f0
z3e65d286a2a7fc2a3717faafc41e59b164c6bedfe1d95da1d55672c5a2c4e327e9ec9fe36c926e
z7e30cb0d84181d5442981b6f69f90c315abb1f90a27892b01db49b88ffcf60cc941eae38e75068
ze93f71801aa7f52732d39fb68f54417d64774bca69d1d8323c6f301d2cfc6f1add0e1632b48ba0
z80de490d9b6609a4877ca5eeb1fbda724e414e68c9e87fb696c7aa677ce52463bbd910c02e5fd1
zb47d0ce774a677029207e20f286ecc1c236949472ffc64d6876368cbdc9ce7a483794a92528efa
zb9fcde8fd5666376e3dd79d92a9fcc3fd6da11fb3ad8f11842df77ef393423bea6b5ada3e4d722
z992399a815c8f1184b3ac5f1cd2d462ea4e59388625f856f01ae4bfa34e55ab4dc856c91a4c18f
z2cdf739c3ee58b0b10b9cb211523b400649e7f63d61fa23addeb809e465890dde4563512b27145
z5300d3b613a3284918c8b40564ed848f4e946070780097126c82e6f381059a1a89aebb1f7ae1f7
z68e37e6e013f889e1a8ec4ca610e97bd451939f700de8c3d8bf6e52369235451431b9a77525b59
zab68874395cf402cb7644ca99617bb89b62a11c1d0d5f475f36fe18210b57e4c9d734e7e551ec8
z763ae571ee97377d45d6d1852be418303de664d8c403c8a680b17e2d5bfc2c08e9daeb39fa71e1
z0d66099784c55bdd8dc486697b6c357fc335ecaf22eb7059af6ceb587c6ba0473e29474f9d4e31
z9c76e72e745e75ed391b4f0a13749da5c1773cb137ccb9cf20f49dfced56d82f076282d3811275
zf3aa8f589c7b1fdbda4000df31946dfa7cbbade22eb6807214d384b9e63dd5c9b80b81875133e6
z05d63f9d2535db3153368e07b8de6af8cf72bcce4a26d23573a1ac7ab013ec77a9231bee041c3a
zff9cd1d8bd0691b3297673fe43a05ab4f7436762ff176fe985eb8e4b56a23da19e0eed4412b0b2
z1989e7af10c5279a6b7abe2b8afede0f0ed5f6f1a019406e2a2d32e68b0da9eaed388b71978e78
zd05b4b2f8b57916ffed5e1348d32f2d72eae55dc64be00210662feefbec6b0050043aa321b9703
z3962aa0b9ecc6190449f4d1b29d656957a3a6fc681ba182c311a8040f17934de572d6d75764738
zd25d406d662690c2bd183742edd4456713b1e1ec1b20e5a1aab94183c6945ce0969d69dbea8f1a
z1ee48c918232bcafa568f201751161e17b0bfe6d04803e016974058a0758b5d4e9305bc9bf9c2b
zf79e2bb8a8edcbacbe234fd06e779744ceebd209eb28ccca22a872be57c3aa771787f6f87fafd5
z34ef5fac808f3dd09c873a5f372ed8242bc58ffa460238fc30a76fa9a8a412f6e711c470a8dce5
zc3113a36411fc601d180b417a2c0983336f8b1d1315d8340fda3ca97a1b744343aa30609448c83
z9ac4f0103033bd0f982715971ae8ee7fc0ab6e78f929950df6f374dd3b4a68577ba303b190b560
zb004fb7cad7e5e654205911065f9a233d83f405ddd2d2a7a841351536414194609a09028da686b
zec40538a2d264ba687041fd3d1d44a59e7ddd5d593365462bfaa9a403e8eb01447cf30504f6a10
ze9500133a8cf305f00377ce1119962c7bc4c1e44af1ec36771dbf7e5cfd18286997dc80eda9433
zecc42d182f0338995bde5b821067879c57db51d7cce5425424c1ddc18cd58f699b32a573fdf60a
z1d150e47b7489527b89f69b1a1f5e2447e7f21b382fce701ec3c943358f77228b93529139bad87
zaf7b790115e3f0b2b123fb8ffd6d68d928678c12b924e7ecf8dd96f32b99df00537553fbcf2e59
z84c15bb909620fa5ea650d95fbdb1e310078b90e5cd9d65339783661b5f92370e5abc4c6dc2b14
z5a9b91cea14b6c67cd771e60b5c6e134758df44a19770366fbfb04a7cd7cb42ef9da44eadefc17
zb4cd9109ea66092361ee3e8ecc4d69264aeac291988ce4cf65cd1a079d094c26843ca5f80414f8
z3654afc3095f65efd526db984172c7d788866c5d80d7e78cae9ab73b5138ba5881d0a21c33fc47
z37b7cf02f167520c65876971b2b0b774f3d2f6efabcb2aaadbbd80927b3ad5771076396670bea4
z73ddb47eba1e478a8611a83f301e906a6ac0d64b024efa308ae6646ca41290c635179f73d8e26c
z52abf5818cd0cf74a87319aa9b842fd7cca93fed16577aed374baa6d8dd567fe55344ab13b0092
z958d21d60f1b37d7daccdffa3f7dae47b6e2bea69305fcdadaf189916a025b8f910a2f773e45e3
z25be327b0e80a8bd8da8322db49b558d92704f5f7bd4bf7d9020d9c4baac80b0d1bf487e96f60d
zfab05c4948074e3b1f6b39cb884d9953158ed2afe22547519ee0df52934a53fd912076a2cb2822
z1ecccd330adbf4894194eefec0419459610918a419bf976ef1dc50a4d8d796becec816a96b64b6
ze5c5e91ca62fe07368c1d0ac40cfcbadb718f0dc5060958b96272d154b4d94bbce10e0a57285f8
zac37c01e3510dc68db9099191b78ac484186a6ab87eff93aae22ec315e7722a6bfeaf040b5dc2b
zc34a9ddca01feb2c950a8659ae874d385c6456b8b65076bfede79d701d976081f70c14b7b4c9ed
zc4153d8623b2f8c049bde0774271db46d039af1f7179aa8e787385e6eed347c17c5a7f6ba03c59
z51bb44ee955b2e7b07407aa2541e1473c186e8e9feabfee5ae143afb04ca447948e3c93a4f1824
z8ae78557a60c2fdeb27907db720fe075f04302ba67d89b9beea67979f91fe34efe6a5cb4d04505
zb3a634039c15fb582ac78a03e11db0bd0ba7caa78315053f7fa1173a355576e3e6ffb0f1ade227
zffb085e59207e4d615a5637fae14dab35f76be402d6845ece9fa2872641fed080f82d93834f807
z58f30a040a500691785000508826d70fa8e763daa548fa048bf0f7b16eddc950621e786f194c8b
z963830c46884bef4a4bc56fbe16848d2c5ff7536badec347366b339142a8c30093d5a30e95d0c3
z96dce1cea2baed99c86e31a805474d461e8358276a4696872315ac6bf23ba271ae8bc34f5fab53
z372c479d94dda31f49ccce50178c0ef24e262c779a48539fc3f16afe23eb4c71326195447cafbb
z1dfb95ec23bfb345c6f80ef63fcf1251686430db74e5fd38afaeb66612b54bd7a0bc995cfd7bba
z100d09d53170763f30936f31c28aa26d2c95fb7db74c59fda21e3796fb132c084559ffa4b90cae
z03ae977a4cb1ce08bdaef95b5b27637fc1161eada7fb8d96538b85b2e92d0addd634882cd687e5
z88260341c5d0ed1c45036ee7c3e0fdb94a8a43c855b3bf08c0812e6e3f3fa18a77e93a55c3eaa9
z2a0f41128185144c4dd0c4a6c1b249b3877cfd1e0898e81b69469dfc3638749e6ee1d3dd4fe333
z0ac0531749fa86571a0cf500030487359f94d55029c2f9ef835eb8f2f68054ff4b2d6671206a5e
z542ed5408be0077129b5d06627a9cb6d671e0cecfd0d9e8062b0ce059ce509d46b594159ef6013
z673f833c5abf7846270eadb30d7d90fb648769f1fcf936a016e048e0e7fec17f18cd6dabe88f9a
zd0fcde1b77d1686fcc41da943fdca9df6625dcb8d926dbc1bdec4a04331a7e16196747fe7856f0
za8d56866bf280386c1b8c2e84a96e95b29b26714cb4775b645b9f59cd9c2700ba0279c8703ed5f
z4615f2454441d66b0e15c59dff3e2d26725a856f6ce66fd9e77ceac92708d19bbd49e8a4a01aa8
zad3d02b66d4f942e43bc29bd5fe52c86a0f85793f0edd75ceee6f6a8b245ae89043af283a2b98c
z36ac7ce4482683ed139bc77c98d34af30648b5270da9022e6ef893d7b4c9ca72df75b237eb4a00
zf6186a8f69aa61f864bfaa7b2138306fb3fb067b8f9a573cf7bf228605a39ea4b7f5b53991676b
zfacc32788950097a59767d1e97c80b380b251f82447e173e803271b73249e15046b162de95589c
zde6ab18b835b7161983e29eb48cf44cf2e2055d795ab2027077d64369a12db3d5fc33c19dd0a78
z9b520a1bea5c98f6dd7723de10dce32a0ab5360f775905d5c0d873007008862ffc2f5de0262da5
z9e5e6d0ec628dba10b4b564c7865d03f2b2f778f5dd493ccde0e2cf361a6626602e7564a9fcafa
z6d00c436b94d34722317bbd66b943ebb71f910a38085a5879484a870faf59b481bfb9ccd9261b9
zad84413f24c6b87e113051fcdb0f7c07138352fbe39a9b555841545adb741daa0cd77af1eb3d3d
z86a1db76f53b822ae3c10e4bd90c28d6e0541245f8eab4c3fcc256f884844e93a03d19a5cc9a81
z881c415b98e58a80c2136a8a1031ae0d9e0ba34e119856fe67b83cb53d7a89664e70326c6cc580
zad57f1375c640b4c1443c4bab2ec2bf614f0f48fc43fb6e29e49eb1c58aff4eb5ef165ade5ac30
zefc5065c007bab1712bf8fb283dc8107efed9cb0a054c7ba340e1095f1bd5cd059df22b1c0866c
zfb63dd911a3fd1c3674088fb6d15f8b9f4b6de61188c3a87e6fe6711de95f144956907bf28d01d
z5831a92fe05aa7444af443d1eebef0036c8ff668049ba622dec821a2310032396363ae499d4866
z93a9766b3ab1d34a74e6619b2b21e5e2efdadda3d622ed728a4ed3685f0a9863b9f59bf1a88edb
z09000e1f6f451ebddbc340f6ec9310895a9b4c0a8042fcdde3689f7b7e0e2931f88b5adb40cad1
zc16a546026423b8563dfea54cf7a68bc44cc1ea21eccaaf3d274585114a3e0f62ce4cb0a9bff73
z029f1061dc1baf75ebe8c2cb6c115288fa215e6dcbe657043a6ae8a37840320d34e66f3150f2ea
z52cc97c8fd0f4c4d625a4079263586637f4bd84a44e8a3efd5a23f12ef110af07e1fb6ee4a9028
z31521274c2ab5f589fe0b527bb44663e6ae750dd576557205072dad2b0d816343d04c2b62543c1
z79193462fc96c17240fd81eb82eb3ffbc09fed30051f01c8ed5d34df2418a1cf11afccfcc73b25
z624549a4350b293f16274d94c9a2dd9c73ef56d0ef358803b761466728343cd4810c1fe257157f
zccdf984b5e0bd9032fce3268a3a0d0369770b38e46b232ef27dacf17fc43c7006e955550b821b6
zb9380a4a0b1be8f0574547ecd8c454f159d0510c60a2b378178d0f964ef67053af769a3c8360b5
z37a8ba94c0844f24acf844d321a9074a0557d4629038f4b882fb052132c11e9bb9942203db66e7
zbbddf08e7f33a249731a615c67b2994eadccf3aeff8faeb1193eb4d4b1c03b64fcc1bf761f56c0
z0cec93c86980c845cf156dd933f28adc1fb27700ea61f3cb74b5f3a2f017c89def8750499a0471
z0cafadfc51d86bd7d03236a5a417b6ba5b8874bca7bd7c1839ea26474ecea3a9ce27a814404486
z8613533c7d168f8ea2172c1d64c4c1b62d6c29a5048c930e330a4146fd32bfb84ad2c4ef7905d7
zfe574169e192be0c0afc9213ed9965cad91ed163355de36ca95a29411d5340eb206033a87a59f2
z99eee9a03e52397f0696549be60755eecc9b061ad06a5943f9aeffff280669ccf5ba7517f2bc84
zde8ca851eb7ebc06f9c9468d37566244fedc13ab2aa3bf332d90a51573edb4d12ff6074e94789c
z7236b77522ed2a3839a96b5de79a9b38552340d3d9dd7f828cc95ad4a8989cbffbc46b9434fb9c
zd5706dced01504edfa194fa85f051d05ff456149af446e1da82740234bdf7325f93b1b6a93d933
z46cfc3b34a20af456f9a83dce829dd5a4f2cd9ff34ac46e159ace104dfdf06b2e7d13ac4cf39d1
z8bc92a7722898d889c20bac38de299ebad99ff738295e6ed8dae3f95036f359352214b5bc7dfe0
za542338b78055d31bcf2f1d0073864dc262cdd2e3b048342cc68a96064706cf4780f4cbc0eb6bd
z38f80f4684d697c856d3398f5a4f891f1769df5157eb6a94b9d57f52a9e62c9950c48d3454ece1
z076c87225c8913144ab4c61191e5a9c89e8c1b855ff1d5f0d4698f330a84035d32500955dc3f36
z9ffbe0768baf29f64673dbb457943792aaa513b8e9043e18ab2de8b2ad6c839387cb8d51104013
zafb187c630ee25611c5bc0478a032b3080fcffffde4c6e41892d305b46abaf75005027d442c3dc
z8c2d744045a745ff743a0bba6f04a94713dc26761fc1df21a647085f703832b7d5e7184b226b63
z32e1795809e33a7e91f6177ecb33d13c2f89db83d2524b743d15556aea57a26748e390b1ef949d
ze3138f17ebfd19afa414cf98c2033bc590b633da95ed5ddd1a0843e4a952f5f9cfbfb3410ae841
z62fff11572bb6f8d539b43fdf281a5018fdcb01ebf6258462980db003d602e9ea92026f278e4f3
z38020eb10e452cd143b3679897c5bc551c55b6777b3ed9b1f7d2c9c742bd2813a8953441a16854
zeef533dd1150706d69a6530bc793a24f20aae1521b9c045c6eef0493d5feaa46769d56726d7383
z0a8951db406458cfcc8fd5732a32bbe8c40bbf81109235ad7e663bc760163978a384f6dadcd4d0
zcd5cd026387d9766d0ec509df3170aa5ef2cfda2c3cd4a1b5016576c40efd35d4853f37f59fe66
z6a3aecdecef6fe7ea54ecbcd52478f9b402061bce97ba75cdca5dfa2f2280be189561585248667
z9bcac13e7d9a40a09d6c66483857f545be223ce7b2f5af9b1f4d119bbaa22d21ac7399704ec041
z7e94c2bddf0b620829df67b180fd5eeded4ebc6fef013bacd580671564a5272d8e278118f07456
z807ff7009a1572dd335511f5f9cf542338fbd2693fdcb9b968d3be2d6369251598e56a3c869742
z60038d8ef7f15b7a38f2d56fef3c148cfd899d9ec749dbc1724289d369b16c077293750fba87b2
ze573473944fb84a69c668b458f55037e8d3a867f40d7b5a04e2ee213efcf5702350c4de36d177f
zc14db38bbc1a301ed8f7c9c2bb8ff878596c96f5d65370ec8aed701ae5a146e7b36d42b4a1aab1
zc8838df49a06504db6d6f4868bdd2cae1cbbd5798287fda6d20740537b7448465e752b4cdd970f
za9dad12a0ab867af51124e7023c7cb2dea4ba70cd12833ee911331230d6ad071241c46ec121f13
zb73c8fcd69ce7001326be8f216936b910ee2cc1b7842fca18f0d5e524e8b99b5df20702db59725
z1337a123f9e76d1b07eea1a40cb8ff5ee451c9ca9e2d004100c43fe5b0dd0559bdf226e352a606
zee8e2b7db490c5c5742c5b45a3f3a3eddd062336bbeef38916b62013935ff481c2ed60c8c4f41b
zf9d5b862e118267a8924edfe4260fc4da0c4b13689f56589b737c433ad6e4e01f27e698ed176c5
zeffe7277792fe7b153b2a50a5604f660eb1c5d9a39dd518d64ea14ca115f46d03ff28839c39087
zd4a63a82f5c1798cdedcbea24e8ee9d26cbde307d5b118da28b9f92cffab6dc0dbe785718dee89
zbc42c83bbb789063a2f6e9c43f253583b5319daba793b489bc3a3d7afbd84261d7b8a910e39533
zbbdf1917b387a9201259784c94fa49910d1b58ad54a0e7a1798355d69aaa2c4f59c5c01fd66303
zc0d5fccb2fcd5febd3b7ce38f7e2690774c4716ee7add4213f75374934e1c15c1297b825a146bb
z189842cfae64589f348fced858d245e8d93566fbdf427d8cdd31b5409a75d967919fa11ef26944
zfad2b1fe8a79df02f80e05280e69aa607703a962f1f21b49997f55347bafee413c6da864b23c2d
z244b29b276e994498d695ea64efd0110e63a8865bc3bb421aff0da6f1f74e5ae90d745bb3be5d4
z423656c07a1d3c91a9f1a1c9770c007506cf2a144a05c6614ea9158743c2fe40aebc5bc117a2a3
z7ebadc99bed909188ebccb500578a2c68215db46660aa0b65ac4a776e2278102f96cd099d17831
zba2e04681a66f2ccb1963c87ce46b32c84381f9d47617911540dac108826f7372c697a152cd43b
z65342394d70a0aae5ca884113312dd4b7e4592bf96171d9b1df547d115e785fb29c4c134e9e2c3
z95e3bff6ef6f9addc725ab292c21e7008916d8cb6bb21099934a3d49d94b9d677b2696e9789188
za0f76e060f5143b79f662b5cbba981f966d6c99c055d01c8db91e9bda511aa4f90992a558cc646
z96f297fa5e83ddd2d54c5f63295dd700cc2fe45ac55e9d330c2d796eeb1f13777d676b38a26fc5
z664d9ba7d227a0133da52e34878549a132ecdebcf56d727f404d26eca35b02bc4e960c415443d8
zeeb2b1c56ef1520e20f1d28f4531e5b340c07b8530476dfdde5c8789045b141509a0e54772c60e
z031309ece60aa2e3eed79ab950c22a7bcbea76034acef12ad5220eef5baed59f7eea4ce8e7e0f6
z6df0e63da14015e364f07263289f28309536fbf802ed0aff3b65330a6a332a7f540dbc0c83a54e
ze76713e54397f79d7452d234ba27a7506394c8a496094ade6cded5545309e0b2d154e796ca6ee6
z5136c9ba8b2a16a041f49dc795985f29a833693c24906d8020ad42acd349c42e46283c3c4e7239
ze796a842d47b086d2fac6f2d638e899b06bb998ddd5d51d96fdda4a41621c639a62fe6f3af255e
z88b01b1b36822642c4e879692db81cae6cd11ba3c1f4faee9df501d915e55898dd35a2e5123d5d
z3c90281cb74b5bd05ef59b31abea42072716cedac042a221f6b1bc8c0d8f120c24762422d79cf3
z0a45f2de1c876fdbafb54a6c9b2974ceafa3cc09864d6935da55d9ba6ea59f04a4ad1f414cc933
zb2e7d4ca1169c6001df420ba8bfb87ac18b4344af7b0dc5e5328b6ef9b7f5ecbe2f0f455f11ee9
z49b08306d6b90cf82c816de6ba56b27df152788ea02eb27a8743f62ee619dac4f91a937ffc4f8b
zcbb32902933ce13b5c977f92bc5cf27514773b91cd012645409a6430db3308ccda88db8e84bef7
z66909ff527612fb4b598505a46da99362a665089314320645e23b9148fc4499bdec877ba12b7b2
z056b4fa5907cb9ab85b4cddeb3d1a48280dced51681f1a5fe6b323d715af0716275b61339b698c
z7d5829a1888d4972120a6985ff0e978508b05bd6758bdae9bb41422cfbe939b971f3cef08215b2
z977d7fa3b5eb1dad8777378296bbb297ec06ed4e6f3a0ed67bc7932cee00b5495559caff93835a
z1164ec578baffbcae20a9bdbd3d3fff653b326f1de4d3f03b2ffca9eb906fff13ee03f58989a07
z977d23957f8f7c6371d218beeb6b7f5c06ea3cd448ddbab5a2207312b24e6caa15935260bbf7fd
z804a5a790c94a89c6b9fc532afef7924dfb58e3d907a5960a1f1c77b1a4779583fb2a47377da27
z9f78e4d267774806d4dfbb2bb419a6282b6231f54dec273f4f5156f360764e9b9f2ea7e853d6fa
zaf973c484e98df489823c4b31558e1e7a1a4335027189240c48bebebadd535179497296014a752
zcecc727705efcbcf05f216acad8380ec8b68b254a5a56d9d481a4ae36ddb00838402ad293b843b
z6f57d5882c4cec66756583057f71a595a7bed41e93aabb88ccec3065e9475823dff630ae1a2154
z23149dc045de3dbd988e76980d2c4d5c79ee421820d6d9ab54ce76adcef68a588e83b0ab253bf4
z0cc704eafd3941ac02458137a47270076d3140dde5d4c218efffb01674f0057a348167b55bb4dd
zd5e6c4026380b9acbcd3be43e89f48271c7cbbb2ab60472bd384584693af0f873991a651815f95
zae0500d90499b2562028971eb52e763b726f5cde3cf5256ab3d3840ec4ef81f3a268fa8ac8e5ff
z050493fcc26edcf924f2a0aa98993e43c15a180a4689cfd951880533e2176e39db98df22a54992
z43cb700d00f439c93508419ef78b3d07dd11f3cf11e5e0752b6ff0accbc9dbd6677c13ceab42d3
z4d500c85f1802d65189e140f6749e5024a0e8008f5c54bf08dd5123ac55933d6577afd0acf0c26
z60b3bd36b30c6e45c70ca8d31b8802b8330bef3b2b35737476be135945ac058b8438340520c109
zf031358f17ce8dcfb1c5ea4411f9b3e3b32ca570abf80b431f16889fec4f48b860966a4b2020a8
z57c28a3c972c870d10eb1ceccece0a9ba54b9f4414d25029b0e69a791f71abd9f617c384677c84
z471876d39114bde9b288d81c65c4d92a295c1b12214b90d57872dfb7de5fd198be1851f822a36d
z3bda4749b730bd3e8c234ccf3110191ff2f042627b533655f50c440b3456770386f476b829b5e6
zb1844ce56f759d12967323d737c580380a6341fb23533e8821132f32cf5847d3693ec42c802966
zf36cba3b1d6367bb74beafa5d6a19043b2ecac65dd6ff9567cc353758e3ff42cbaf9df19e206ae
zb82c468a58c36e5be08537c80100cd43e970fb1e9bb8e2cb230bb59e4ae3e10d973fa631caa2c6
zccddde353e574e6593f4aff333424c1ca24c1f1688a22292e015b19163078f9ade42cb0fc394e4
z0deefbbb3226533559c12971eecbf9031d8e2f586a7e867d27e6247a25e612340d0fca86f181bd
z9badd9d29f9577490b8c09dd73ac1682ff8f0c3eeaa9cb83abea9f614012511ae3d2f3d6fe0ba5
z793020452a106976d7b1ff62f471644f1be04bb417d4758b643152fb06c761f89afd41f9664ffd
zb1b266d88a0116f24fdf5126dd73cdae278ee3bd849638c00b79274e9c08d144bc89072a155a6d
z0d18a7cb005de63aa353f8fa80f820d849977d8644806124e1178de1de3126c61053ec7558b031
z03e42a090606a7a3ff99e1821a0baa7fa54c9b7f64e158a037edae2b329e01e2d8ab8e3bf5019e
z75b94d36f0dd0b0bea6c54d61201479838a879c6cad4f7f2291e868f96873eab6f739622acf627
zfcb97179eec673a8873ed3bc6789565781fe6ada482f1c8171d584c9f41dce276be167b28cab0b
zb728185a84ea07638788be4ca5eae47665693b7ff14398338c13df6f184bd68b22dbf980a752f3
z4cdf79c3c8d8e3ea9c0cb6a1e407167e84482de3bb0284eb026ec50a4e6abf4bc678e333bdf0e2
z82949932c3818186033e70c311e91597d3da8f627673561024c3ab41d4ae6d75fc5a39d571418b
z5ff84b474310723bf2cfa1ec9406192721fb8992300736fc9d75bb33d52ab82a5eea22dac948e2
z81b12c2aac2186347416ad38d8bc5822b94e93cceba7ed6c30125b5b20c2b9a68c98b2fdf4b3a3
z3a6dd19bde98f4b251b4012cab068a776b4ae05fd7c159bd099adbf004b07647d266a3eabe62d8
z5f929acf3052f6d798152b5dbb329044337e21cf3f7fafadeac4fb1b4d8c1d9c3cb8f62e800ac5
z12699cccdd7511eaaaefe171aa1d2aaea9fcd17c26adf38ec81220f59eac908ed218dac139ad01
z90d4f095e2aaefd236dde79c4af885223fa8c9e19c91c9417a7070b46a0b3ef89f1a96955e26ad
zbcdb333b4debff795ea588855ea7975d1a37bf9c55d66856ff58f07d1fd57b5d2f2dc5af57d79f
zafd5db81f492b45a2a9447d57460678c1af0db7d18af9e6935ca1cd944235619923f5bde5ebfde
z4a33d56e1ddaa22716866461eefbd384a04bd4083cca85c2814d5227222bc5de055dd20aa9a1e8
z7945f6f5fcbd27dc0546910fe0bfe5d6bc73e4cf80fb7701573a01359c3a9ad46da863fc669180
z339b29442b595dcabe564dc69dfc1ddb2fde01159dbf7045ceacbc68fc8594707c14223d2d12c1
ze25407fc01a9bebd0d52ad691f501a2b2d869523b70d56818154311005ccf68e60c061e8ed6b96
z9cc57e9cb171773da84eb97b8e54c9d7c779c2e4e6b5cb892732da5f40aa0209c55320d49294fb
z1b2f9b3c79e214026e002b733696f5c290bb1cc7a66fa4a9a0b533d74a7bcb1bca97d5690ca8ee
zbc7972ba017836d5d3bdfe7b6c60cb5c8915d24660678a08555513614df5ebfdee862a2c669eb6
z5f21d02e12676c77adffdcb729101d60539315312adcdf548b0c729e3954aad7a5f237f850ee02
zcfa28e012b82989cc59db813bdbab74a18776a42b355c7cc878730d748966e2469592cadfbb58e
z1a2e34134c23570aec10af28e19d0de01516320d9534996cf9410ecf3e81361bdea78d428fc08f
z732475b24c08ddadccdb1a77263760d53d44ce13d602767230415e5b4e1bac9dfe771dad94b992
z9eb399c53af59889dd5233e1a08187834daa079ca5a7d8df0b6fc6c3c199cacf59121819536ee7
zd4e14ce6d5cdfb99572ab78f54146befb53f0dcf351036cad3477cc702c84aff909d63b3aa3b2d
z3e79321278692eaa53ac0b7b9ea8e7a83f1428786371e517b6dd1e681d277961d1aa8dbd59620f
z65246d2d7ea801ef42b53c1dfc67a26dc4c59a93aa31d06d69d1409fa7d5d8277affcf1e8e5952
zdda108750f8e523855ba96b7f0fab4083c4c6e2f848d3bff4990c0d7f039a2689227532f8ec949
z8a57717ee62f3c807b5ab32588e2ac59c0083c7c85ba2efab9560fa56776e15fea93bc4f2f1c25
zdc9f86a8979a368394e06436394fc3a986ffe619fc2482a6ba68e0419d504a0382aef3b322d0e7
z958d80af3ef6cb24f8d64cdca93a42f79c0f151b6a9f94f7035535366aa86e4c442757c5a7538c
z010dc6e2d11bcd2ea6318ef6fd66a97c73d28f6045d19aaf33f8881ad708b67f1a609470de6ad7
ze02d7a96a5d08c07eb4d3bd331fe492eb8fe6592e4ced18b227ff8d6b971b0508aa3e428de4681
z652585839a4c4109beb0dc525818ee4054b778004cb0a7d71327c53634c5916b4023e3ebfd7279
z9dd13887f3d8e49d4b6cf36f803147de0fb8c851dc00d1d674edb5bcf7660c50e5bb6367a3cb94
z54bdf415fc664ddd1abe373e299a153347c264994a6c664d1757a287eca1ee331913b5b2276a8d
z820e0b149fe093f5d0dcc4142c7f55240b1f63f92f61b39b2d196e5a0d2003ca650cde0c09f5df
z54f35bb29cf388fb7cd61ad9ca560c3120a30205899b8606a5d46a46bdef58a49ff5c12623d817
zfcd1de26474fc729af051ac739f7bd65dd043e49483e8f5985aceaaaa8b3ada473192f097a0a1e
z822a996253aa40cd1916dd131fd44b2e5b892be8c0c02d76d8db6be5ba2eac3be20ca1603b93da
zd89be716edeb00535806acd0abbd8b347253d945acd361095e6780e8506e1ec63dc6f8d618fca8
zcf5df575d6e8c08a2015b5bb4741e1076fb11b32545509e3c6667326b54611e1062472359e2756
z29480053fc7eaff701cbef2e15eb55908991d2a4efb7af45b4c0f21120413db6bf61ccefd5cc27
z6937b45eb21f150e50f21b7085e9f0a157b06b66eaaf14f3661bf674eac4829f515ea48366e6db
z1fc41622c39ed4fd30ff3018432185a98133bf907e123eff5bbb0b1065ab639afb5e37ab1a7c30
z1eeaab5818d7dc33b02d66efbca7ac3dab4cdad329aff87ee1550b4ce2c6ee14f1cd2c0048fb33
z63f93b665bd27109164a655f8b6d01c3a1c7a96256b04229d70f70e358ab59da20bd1ee5f4f770
z56779a8244fb218471247bc51935b74cdd3daa7b0d15e2320c23eee65e7809246186063d7ba380
z351b906e89f97f1edeeda27806d188756146c0111a2d48ce20efb9fb0c1e0b715ddb3d7ec96b50
ze90b3ba9080b1d19ced68b700a71f11eb17b02d6d2223cffb5d6775e763dce27362066b9e75e77
zb89c26ae20dfb590c9bc1fdbe2148963f761761f92f13730edf98aeadf8f81f282d8dad79e6648
z22b85a185ef99459ebb604863f181a92bb82dbaa3781d00cfe382799b28875161c1fb3be018807
zb7cb991575a44ff7ce187de4b5076705575316d0bf27efc2400f5f26b756c0812faed954b85b3c
z87e4eb278e568a81c559971db99ced1fc9f46e56336323c87c926028b45ff9e3591d43b5c2134d
ze6310bd4d4734ede3df894c1f48ed741990adf804baae249d1a700ee2e1819f47c2cbe5b6c37d2
z9cbdbc800ffb4130b623d4f914b1a159040824d3e588131c9112e26df671d134e35f8cc5f6e443
z54f6a5edb9ee30c6d19602e2061a28beccdd3cd5fec53e5538691d06ee06261b9226a0e53aa3ef
z45a2634938e2327adb947428d436501834bb53058a0320b113a0fac8c0f4e76dccfa75bff9b497
z323294bb4d63ccdf7a87067f18c925d78fa1f74eaf48c7e2bf799f26099546324d66991aef409b
zdb54f38340fb860ee910cd9b364fe10aa688e48250151a44e0b8f1d5d5ffae34ff604f6bca900a
z21d2f4dfc5dcab60dde899f798ace1ef08a19de5d797ecfaae01745b9a659c6e23e700b96c18e3
zc567a4ce78495aae3f218fb51f7dac0d223b17df57dc671a99fe4d819185c8c728b7e64941ab17
zfb80ad29922a83f5420623c00cb9abdcebee740ddc2500716d0c7c343cb0075df2155fd513abe5
zb95331de7de64f181c39fcc5ff213d2b2a885775f9dd4d3d5ac696df3b9568f319601d6d841030
z54f2fe27f939fac4ba1238ade0a061b2bd07a481c29792faf99977799efec390675e6aaa9895c5
z922e2008c6be72cafb95dd5d79b51ccc35e754ae18274e23ec38ef6bf2e77f7b8738b669485acc
zd7268ff789bad96df8cc238d9d370ead70873d595b3a899ed0c10f6dcf76b604bfea53e7379e5c
zb6ddfdf17989e009cd4ab916f1efdabc17b7d4a259d7521c7754f040b262781db15b87b902a824
zc584e0e88825f8da2b4677b303ab7f72dd3e5c9343bb17e853f4ed615346d04a38f7a779f3c3e5
z1c406bb99bf2250631d36d0d509264a82ed424f8908c870f785c588131393362d82634ef155cab
zc6d89452bf9f7e9b6ee7cc1c6f9acf6b4a27e60ecf27c4b378b37f4f1b8a92d88ebb54b84bb8c5
z4880e2adbd804d90baf4bdebb6ed6cee140dfb224b62f45f1c7ca60d13dfb81a50f7632959f393
z2cc5075eea28c5f7574d0d2bbf2be326d71d498a4c04df6f400a3310417fbe546f56f87e5f91c6
z4955aaabd879391798e154b7fd7da7117430342a1059e3939ab40f53a911f14bf1af39c1b3cb06
z741070c646743de88716110cd3f1a9bb58bf55c0eadc1c08443e38859faef1cb89510b72ccaf52
zbde2ad7481eaee74354f8e284fa964776c76fdc81cdab14c684a323517e0af48ad05180a72ef9f
z45bf016c9d04702774b3f9b3047c21afa5f82c41ab289607b5742b814b6d8a726f010d59f1c23d
zc278bf0eda24f595c79748969f01c10be6b0192c5839878fdfaeb87c48e12080066036340689f4
zb276378040fa703f5a8d61fd2670d1dde3447ce8133b376e779918f365a21061668a5ede958370
z522dcd7e67f860caae8f9accf7e2b4ed67814d4357109880fd38ee5b0dd93cfeb69c3ebd9d30e8
z25da89a47986b4fd9c5c7656922867df90dba012dfaffd927adec8edf80aa83760968a639e6008
z493c3bdba4aee4913ef6512e7d6921e1133b29673a659c7d265f158f4d7932c1b58e80620543b8
zad27993d49265b42c1e1dc821d89d3299e0021b2610cb01c7f45b987026ee5b0735aa615456ea5
z8935b421377ea65e5d9dabf6f2ab8f5ab78047a292a8410ef38e2fb7711377323162535107677c
z51c442650f08e8db81bdece8f500a041cd5906535a7b50eb5f75c6b293c2cd099c51fc84913e79
z75a073470509d3e669fa2f39e56d82afeb529bacfed9524958223b6454e638d521b09a3e2ecf45
zf5484266532819a932150ac4579d546dd2b0c722e8c1e6b58ad910f009133c62f89b8b5737409d
z292fe151b18d2c1fd7cc7479487ca555458bb38e01597765dc8c97d5f48c10f5f4ae85bedd0fab
z2cd1ac3fa83de8b51b4b8aba799b1fa8c82815f4ec6d8da853ee3f8e7f48fff7841fe41ad837c5
z4971973eb71e1275666ba5a3ac859c9ac53e2ccdfcbdf88c7e6b7296a7e9e60915af4fa978440e
z361b2993ae9881cc0e7e95858f9f27875e55d1b124241dab3f3c4b06195685b84b69cf85770a42
zea45ba3091c21a941271c0fbc9c7b118e7860300001891891ee7ca604771d49d7d23db224799aa
z9de0cee5bdc42098ef9234ce12787d5f759269e6137564c66260e6c57de59f93e95f69004c9084
z32a206d932d1dc0dda0af7e6cb695016cdfa978829e2863dd02a89fc1e90d68dfa2123b221f9fe
z74b419d618cedef382ab75276f30c81bc5b64c66247320a82a40ca6966a30b6306bc3c8a678472
z9b44b2f8f3cfc59c796014781931a8cd3058c51a83ebf2a37ea50de13cb9c5f1e4cd8107efe9a2
zd389ad2f249d632afa79d70704e760dacf3ad3dd85a4053809d36278648b37df4172ca3ae4b7eb
za3708b40eb2d4aedeb76ee77bce3ceda92860cb1c923e74d2526c92dc27c7382d3b612faf7ce77
z69f859b2a0b9ff5978b879ccf1908aed84740c147d9c1a3ddc2894df9ba05ab734905c7ef22a5c
z4f73ba9feb746a319e12a71ad0c03bd65f04e573514664e9339f36df06a366b16dc083d17adbee
z6f8bbc4aa19df4bfe1ccf6971124549735fe00eecec800fafb0d7ddaef4f938928ee9a4bfdb4a6
zf1f071f715a94bd09f57491f1207c7dda84b27e0b41152ff20296c81e18bd452c9011a13e60c24
z7c490422739aa36e908a46f0238f3637778ee9bed38561ebe0d6907d3896f1332f691c711190f5
z8e0b3b7576af3cd37d9dbb795c95db4b491ca686b48ac7c15f0d97f9275f3529a0d877430508fa
z57d5d814bc5755d6dc63126f215fa5cff9c4504b9bb5771c305be5ef88b8ff9b9e70cbe5d2ea27
z14ebb706e943ffd21160d3c4708d960c9796ccaf6349ae52e1a780a3a6f162816036dc8f42f9aa
ze26aa2e6a338e3ee3d4019269ae4e16c00a0694c3af17a3a7890734908074403576a0e53312815
zfd0106368d4c77567c12bc26df8cca63706bee7cfdd77b3e35aa82e67daa792df177cabcd93d0c
zb511b1a7c4691aeab44a3c061c4f5ff68f8d6ed2961f523012cff20d333fc42bbd7b8640ac9285
za0de4b52363342e88f434de19965492e02e93845301e7681da29b9a0019b1845dd226b2efc6d9f
zb04b16c3ae24b3fe7accc7ad28c2767c09c19ffa66a9f9f8b690d6add0ba06423ce8d4ee5a1012
z1dc4b2c07e8ba5019e407701d941aa5d60c5fb0d18b473ad38eb8b0c954a10d03da08c1156f52b
z7c76c0dbd52727517e6cb5aaeecbc784d729e8eb35143bbe1641f977e00d1a6e76f770c0a869c3
zda8ecd327997f75ff31c3433ab1005ec4514a2141c2216e07c6c29c0df1187a42afcc65c3c630d
ze936bbdf6ba1a30e1dc6c0a5309c77a50636e130277141b1e5179db093564bbce90e48e81b9711
ze49ce7eb6d9463884a3250f13398c385a1fa5bab104ce95f8fec425ad0474ab76dbdde58728d83
zf9950f18055b53b3b16ec06178f387578f223a7d256d778130e4ee822e39585e2c7a960c0e8a9c
zad54cb55835dc9dae586b9f6d18b4c8c8c8577c86101823a670c63ecb61a5108d4e7f435f9f900
z3509830834b7c5a0f2b3d881a9a1b5ea90676fbc5dfb194f40ef58f011450e8520d105ed428de2
z933badaae5c103c63058ff6075d21956746c31fe430a161b6742d050e57b99e503bae15dd21f19
ze9deb232bd0f846ec15b4e441de7fc82272c05d3e4db3d14762bd3f20ce5d1ab05bac5d676f3a5
zeee256e09694d5c0f2d1818f8983b244cb1e25e3d86ae41229577ae938dedafa8bc1a45a9b65bf
z1ddd4b3122aca3f7c0fd1828035320b658829fb58ef0be38fc96ea20416f8f3359c16497006db8
zc0038f593c5b7c5d88344e025d0c2a10996123c0a4e75177c931ba18b38c18041bea9e166b07ff
ze5a320c8c7e4e35e01b52d9b13b040fbf0d93a2a024ecb067ff52043f9bdb039aae05ca16e47c4
z8e665b1281d3fa4a4a321d1d7c914bcb0b3725ed8471dce33af1bab4b7a059df8e859a34251d3c
z989dab83cee7ceeafc2ea342f682ea503eefbe4131ff44ba1938d5c8f418a774e94d31cf1a07a8
z12c6fd10bebc1caf55d7034dd4a11ffc1dbf1343dd9bfb23e2cd8474d9e280cd2b33425dc76f3d
zc4d5a734d32fedf6ca17e7e8fae18293df5bde227ad56fd54661bf954be605b96eff46d263cbf4
z82e2c97ba3ceab5c853938b59e2d95780f2f447213dd098321d474827fb6415a6023fdba6835ac
zaf817bf0e3502465ab6b6ab65aba0f972e80d1716116ff8d96657651e2dd41d23a4db977524b72
z809cd63b073960cbff5a9ea351c9174258e8f1af0f5bd2637b439bcd98c6841b7b6c15edbd0bc9
z6ed5a707bb375029ee2dfdd40ef0a57ee5aba48f4a4eb4d6e37f5e490403ee442e400bacf74c85
z831058dc58c80b257cf2ac2387757027528c5e2f17dd7dbba32c82b2c28d3b4409f54dc4b78ff6
z6837fbd420b3fc3b3fc362052bb4cee2873ac4b49bb897b19707e13923cc434444a9a223e6dc62
zf6233fc4c22ced1f294aa3009b5634d9145f6c1f102dba746da5875a72f243d7816881e14212d6
zbe99e0d3a59d8a489673a19ca8735229262874e354c6a40124a14e4bf2cbb5c93d9486e56d9c2f
zf892f168fa3f02c0e0411296ed94a1b1af67071f03a6b66649609ba92c739e05b1d77910bcb20d
z92248ea80801e72db44b4dad2139e121e86b6cb5bd564db89a9d4574f8c19736744168fffe26b1
z4bc58d07744d9c00ffbb0f328f1c788fa9fdd3d3a903a7aac74d7bbc384842c370cef400832845
z3e5610ea0a341a858d57c8d23e97a724804e5792cbd7e55dd34bf3787de8628e4e03ef20cb697d
zeabbddc787cb985a905fa61448271849808cf53d961591152cc5560abd21e8954a05ace786f790
zff40299d01c47b91b5e8107d8c290732c93fde2317daa1851fd9f16c2f61820e5151c25c316b64
z456ae2d1be677d0f0552335ed6732a860680ac1037ea0fcceed0a2900265364f0ae35d4048de67
z726134523dcba2c39dd79d7aeec00631441ce894ae97977694fbb0d533c34db8f560f32a58aa94
z8e00a0e80e5953d71814d4874134097d3074df9fa2edecbc5657ef8d53a7b321fa44863361c8fd
zff72f6a6caedf8457c5ce7b9d999730242915b0b9a9c2fd6e906287c8bc9de6781e894278f2178
zaa9202f81e259ec0bb3c7168a8f286f7505e94e0a30c5ac09478c62629a8f37e163102aa197c2b
zf9d4109efc79505088a3c22b8a26f81e582ad3d0f2bac76e7986db4d326d06abaa655cbec531e5
z19442dbb2c2336114631daec6898ce952e7582d3c751cc28b07c34b1d7be8aa92ed8fdb3c10d65
z67900a5aad298c4f4239d1a55d8d4fae1bf731e1ffc178af90d31e3ae6c3644be8c84c5a3fdc13
z0d24cc65f06436542de3d16f5f3db34e8b8a49a4befd9257f1fd33cfc3482c4ad7cac1652439bb
z7cf708376f6024d7ec8d5d0df2ec10132daf4a3cf51bbe1be6697eb6ac3f664b660986bb2c0ed5
z016f258d925cbd0e0934f11f8094a472c27802382e9bc73852a223133e839dc5769105be711c63
zb2a3c2ae98f2f759f2a8b45fc963b1af1f4767705fb5d06108dd0a7d5287a92bd21a8804c4989b
z30b1b97e6b5f07f56da1e0bc7f9ade7bf30199f32a90d48f1d314834599be30a7fe33761520e59
z75e4ff3c6ceaa3caf408f8b00d64bc30a845929705d3f1cd12673560cbaddcbb70533da8f24db2
za86c3216d1935cac1ca608f1da38900238784314be12d1a5274a4a5fc9e8b44ea6e0af78af007f
zc4a2026e8c2df096a19502c39d63f2c94720754fa6aa8effb43726de3ca2218eee032be15b0a1e
zd55c3c192f21bc6efdd149cfa0bbbaa828b1f517eb42b71f6999a19c69280857c8c58569031f86
z2feb4e3966b76da4536d7d5bb96fd324898032531e7edd161e6baee85a18a28bf3444c8c1e9d86
zd1a150795229d7bbad1bc52353c231af3135cb3a9312fda18c69b5992d3c9809db494032978ac6
zdf4ed4bed736c9d0d4b59bfbf27306603167772cfd8fb11090fc6b7e376ff614f2a66395750f92
zcf8ef388faf260424d82ea338533536d3b139b76d558c96e041c82e1738949a2fd30b4bc54aee7
zb04e9f9d296f4a26413bfdf02964b78876bc8d8da5b3ed1c019c7eb5661e5266f796bbda4cb59f
z6442116765c9cc778bf92788827a4183432a27c9f80485d450cb2087c2e336aec15f8d937e8bf8
zbcc1dbc7c35739a409c4743a7d072f8efc8a7ee9ad842a3b0bfa34c82a8ef863081f19b637683f
zd84a50482551e3f70f7f125595637bb3eb5fc286f6e9438ad31a298f7e51247c75accdc716e22b
z5f35e3a907c5877040dcf158d460768cadd5d69da7d58931e7dafa465b3647c39280b6c72f92d4
zfeaf8d31ff16bd141dd1ce46cc810f1779dd6217ff5c713f9ad8af82870d1c4fd0db9df3f2c335
z9965dcf51ca62b464074dc25e179add7e200fabee332de8542a955711e35a91eeb2a6d71dd7c75
z287ccb861390669ff34f6f6fe41c29f3e6028e8a84aef02586c0388f1e69e2feffc164130b64d0
z555d0e4f990d0743279ca5c9208880c620493a01be26a37b272045b50a08123d7d9c17e79a52ae
zf6c6ffd5cae4579f61472f1d74c1699ef31d483068b98854c7617a8cd4eee66e58160122cf8844
zaf5277a29da2b4631b181bfbcbfaf9a67f1020fa0166e8703cb8409a0da678bc4116a13eb5538f
zaaa9e52da0580d339f3452501132d41ef6d4a35db9619a17843dc4bf52cfc6ab57ccd528e45d19
zef579daab7ee9fc7bb44267842f702a619465c127ea7dce04944722ba61e50ad1d020c0e94ca46
z96944644801d01f80f015f523df0e379bc3f51ecbf58b3ac44c42c04ba038ca64074bb816e2e1a
z285394b1f56f93e0b6b7e06b0326439c62af25c209a49b5de3a121e0cb549fbbe47f06b1edb980
zd8a64fa917403381d1eb17d1cd2e37a96fe63c08caf94c921e10fe64655e6d675bc5b989cbf342
zf5dff18419dfe8da1923c52d30a7e5cc8fd6960a51a137ff82b95c142b8d1280c77cc9204f7d66
z6864eb04a9147a3db3c774de8c6493af91e6596969f4a30696578574d5685a24e834e80fe3b914
za211636e8df6b4f808a7f2f3686cfcf2775ef1926923106b34e0db87e8a2d828776c30f346fbfe
z9f32096a4f17ef9b9feb767914d09ba6cdb5d879fdfa9d5b41d5b5f8b7e75e0cb0156cea38ea3f
zb8ddb228b280a19b17a0552d5e747456eb130531a95da803b889990ae15df6ee51fca2a2f0efa7
z030197a4db01a0e5c6536173d9e11d412ebb2b0cc2217248c8b14cc38f30a8c30a34f81f831477
z8d6ea2895338d967c887348c69e164174bcaeede6a80fc6fb24f8324e41952d4ded4b90a6e1b8c
z31effabe0532fed51cc790c7c4135fe1a1f51b35fa9a5118342a74691e3c7ddf14c71794c195dc
zdbd62efdf80c6a77c0e805ea0d88712175c05f89e7ea69023d5c74e313a3bd5e25d3e498cb72a2
zb10353ac65d786bfb99d5a4fcb3ab53beeb01d15f190dc6ed681750cc9fe71b2dc7e7f73a5953c
z2628f5f84c01c27cb94e5eabe9da717991f1608b7480dad9cfdcd6c9f509c6c1120db2ea681266
zb8e4c31e52f7b6fff9c03f00cd7bb36da3a5f05f64006537cb61e83dd892b3e2b7eb85bcc39025
z3af719402354a708c98854f25f9d8c66c9cdeb097b2b7f03f13d52d0a736560267af54796cc861
zc987de46652729c4b5c646d0e260fba7cb75b3a467e3427a6e653ccea52d48e631c349f3708f3c
zc54d6e2de4701eb5536c108746ca6c0bc82ed9e4dd0ec94a3a254c14ca1e7547532890ec656860
z5c61e85b766a2b2125c716adf9c19af0849175d03fe8f1b2487dfa71ba5f0e8a245c4e573b8fdb
zc9a87a2c4b448052a0d10b15343bcf5cb76b4b2eae5d08ad5f7fb6add00fa7ec6b0aaf3a5425aa
zd972efa79373dd5686fa6723ee3ca37d21b6f4078f999d697b22d0aa03983f5d6f522c509b9c0a
za90854eadcd5900748afb3263476dbe9122e5b93742543e798ae73ca6acd3cf08f5c48ad3618cd
z65269945029ff8ace8b5329bf586e0965aefb69d3aff322bcbb5690275214c3bf58645d9b24ee4
z723a559f04a92d578e66be501a345878830fd62c993f0d2a24ae10a9824cf9ff1e74587580ac24
z45f4eb0a2f0275efd646f67a32e3cd748e4e94a428538bc25e1bc6c20050a1aecd4f26d8b25707
z519942ecf7b6f707e4f2735546d1d8e50c7efa6f90999eb7cff0e3724ada723cf9ac2202e29d1a
z402a6a34605d4f10856adde6bdefd83d5df62885b264e6e65e652d557a3dcbb1a5fb4c30181158
z0249c8c5d8151e32bf43fbfe29157d2a129b6c91c8fd8d42f5ba1d8b95508e16cdc02fdd32a883
z1ccec17ef1cc63885924843bfbbfcdae334732ea4240cd42ec24f2b21348b2bd79f28d970fc2b4
zcb61f4fdb15e5a46e015596c83a13a160402b507d9c6fcf720fe8bb7dde5f11a983093a09de5d1
z3c98c16d61283dae9f4dc3ff7b293ba9b087f5e2ed347974f229a5176cbaa25cbd43ae35c6c9a7
z0ce442bc135809c7f0f0a6f2a017362f31942a9ca3196f98c8eb68c62edcadfcea3f8b37ffcf72
z8faaf7241d2efc37ff8ec45a4fab2e6859243686a3247758b8c63b1fdf6e2f7ffa5210fb682c8a
z9d4cf1dedc66d8f893c419b42faafa74618f7347df4c137ca161e39203e75d1477fc627432d6f4
z4ae8f03e564102930d2f4237a4b74752f045a783ca606b2325e76056cb821163f70887d7d18660
z7ed007e1afe05978efa52edcf645956e44e75c898220f308bbeb326055171238826711c9a4cadb
z92aafa9099354510624fe6c8aefbf183860d148e55ad3ceedcdf3bfc016a6972b4c085ccca74ac
zdaf7dc8c36f32bc424fd88dff03e60de2f65cb9aa95f6bebf9e399557d6eac93d9ea1477444f9c
zc5e280d7f4076e3b029fbcd4a507115032d05281ee13bb14acbc0506b0155b210af1e46edefc7c
z1df14afd93497870929c36c7b769ea04ece53dbadf9296f566a4337ef26232e7c8589ce3784c17
z8bb4ca5f1705fc590962775236322316af22d78c8617f752bac8ac1df42e4f0a1a0e3eb6e2341e
ze834aea074cbba2fc52917083a05b5a812215dba7b21979371d3e8b5aa0ca85bffb25c3d37bc08
z81604329e4e798ffcc196e649e1fc4e80f3b063fc5c55206746e05a969a39a99577b1276e32289
z6c5bf09d5ca08060a0b06ed986debdf811ee4b5cd8412267284ba3c7e8f8ff9132e41959c2f6c6
z3de897f1fe02e4aa1d114016b93329af383a55e5cef998aa2eec4ae9b7a67650633d27dfbd42be
z79b354eac74a20b90f9ece4b8247911b20c4c76702efc1a5de63f999b69fb0bc5fd0f4fb946a64
z2018e14282225cd4e7954b5e1240794db9710df24c4d434e5781c61d3fb90f40233b95a1ca01a6
z988e93d4ee36449a1c9ca7ac9064c3b391a1517769af2db3bc7be330b427ae0de50ba517989432
z602264413dd94086ad9264e9a68e9fe1cd62dc114d27d93596d6d1a638766ab84e648d27966753
ze3788c3d7bda4f2ec82bc97ec81287ffa2a4ba07603004e5f2beff7ee250f1db78e99bc565a0a8
z4de02600b39518b1c211af580efac97f6f304816ff122505a0081d4c31d08e79f46ff067cf56b7
z7d25cd1304e6bd7a4baeddf0b0415dcbcca898e40251e35b6522b265aa068daf542cc1a4e4e774
z28dce916070b06bdc709052a6bd1ee27fc25e6671e7cfcc1d8e45205a0341fd3900b270340cae9
zd8cc39c2392bc1c6dd6b46266a8d204210df6eed3ebfa480501a6d482d474fce5a7f9da9c9eafd
z1a92f17ee953b43df4a72a1c41c5924aaf6ff3946f581c2b7721b1317f13e8f7be0a26af97fc14
zdb4bbacd384a352e1f9ec705efbd61cac8a74eb92892a249ddc17a8f2c5d4ebd231db177fc6715
z4e079a1cf7be5a2b9294e5777d4a563c52a836e0ed9f4217412d9728a1ac953286892ec4cd92c2
z3e37e2b150358ac763b47467f91b58710107e08e5ecd0874d119599e023d7f8873d90227f52d0e
z3a5548a3a04fe933bb66dc0053b708163ef228a0adc9dee75f993d1df0bfc2945e2e87ae03ac6b
zfed169286e74a354de278383d26df8442528c32376ca23d173b752bd7f1ec8206e2c0a2f24c9d8
z3e2159e728be5bec124cef2b29e5ac10b5782c0f212df6b17ff18659476a6570c129fedeb39666
z198e62eb175f9f527b227735fd93f52f826d02522687d9ba3fe1f5474cb43ced058e4a6981cde8
z64b61b45344abdfee387de781dc54d9e4ff41b5c71da19ad6828e47247fa6808e87751bccceb60
z3324808aa2a0090feb5eeedb1dcf504c8ed5c735df4c2358614a53da6f13b99094a26fa8fb9047
z4d0e64227431cef6f064193caaa3675d72bad1cbaabf65bb4616e4dd25e9a3b1359693f21264a9
z9ada14b2dcaff595db0f384a115e0087eff70cbbbebe7e2b4f93b29fc7bda5d7ccf5be2ab67c29
z0a6a9434f7dd551c08694a233577b97def4496d9559ae6c15a503f24eb147d3312773e3fd42a10
z1420053516c46ba8cbf2092129ae7286509def5814d8406e052389df5d88e549348d09927e42c0
z78ed39cb2851bffd4fb26d81bbf0732eba0ad646252a9531a3da2f0fc9fd84d179eab84232ebf4
zb061fe6fa14e0542ed1c7dabab3c604e4239a03d45e9c5dff684acfdd14dc0fe6cb9787b92dc42
za0ab154ed43fd98409d2cd7efe9bdef6a282c86337a628f18b3bb3cbd3ccd70ab6e40cb6b53a8d
z766ea827e47705d1323cfcb7501e9c9542527384f7876e06ab53075c1925087d9b4f7feadef1f8
z9368bfdb14e073eb8e8ff59e9f97c7edf3f2012bf849cfe52b581460bc86aba731d81eda1d9455
z71836eb5676a04d6df7c70133c219d3a3455d2064861cc21890cbd75383ccea289a182df439b94
z03541d9763b22948619aa7fc3be4ee25d2ec6b1d600a382cc2f41737272f47146db2b4610f6f78
z27449094be449bc55176d8ac42e26efa2cf157c0f8bb383302f8453fb48f4fc7cc799b4377a4ae
z0965295c2299a2fc8d47ac66ebad3e1c13e58c14e55af7f5201b332f4341a1376e928212b5d981
z7a666cffdf2b5fec1f0425c1d220f478d8d4860172626ee56fa0e83bd04247ac397f0d419ac801
z4ab5739cb8cd1cc845deab11c2e0bc571f7ca85fdf828c92702a92c0bad558c6a74dbfaccf6897
z260848f8dda726b8047dd4afe4e96670ac136ef0d3b6c3241a145bc73c77e4f58911ed8b8e775d
z8eb63f92ebc9f9f55bdae629ef131a56d37bbf4da2b640d3dec8c159caffaa107cdbf8a84b5a29
zf5b34cef928298994580e89bd304e6c067ddaab439df3a0a3865039473295a86b3c5111ad34186
zbe82a5dae387d174ea4641df58db3052d19239043dc6ec8c1126078611e8d534333aa801bfca6a
z902fc552f19b61b1983801832f6484fa680018a30015bbfcdf4174563b9b79ddb5d31061fda503
zf4aa8d47b6be3def7db581d58978b56d68b6711fa5ac2dae2e11f0987373c0f551d02d7bdd3704
zfcd57cda1c79d58c2c56e9ef0eda9c90d355c3492e214672b439a7b16b6c5fbe84bc9babcd6f1c
z4f16ab3fbd7c302ee8066c116b7a722a206ea2a7687f19ca44bff3e7f7da34cdbbe10feffc663e
zded44c55d2e43fe65cee1f764e2f2f8b93ea707531616c63f227c556a8f59cbd9542f115a71b34
zcd90628f98661024d5589259d3dfd500ce236f923ae62e14dcbbef20ea96ab13a29fa6679d284a
z31e2157a2aa42e880dba23fabbdebfd0d87f3044644fe1dcbd984f11d4b9893d7ced1d6a95a02c
zaaa0f13c459ded9baede55a25145ca8c3dbda265db329aaa8b6196eb8918156f2f6f3aedee0e37
z2cb2bd9495633ecd59b00416055fc6ae6ea0a32f2bcd283fe498b3a97c2ee6ce2f03768cba3ab1
z4a042549978297f2dee98b43e48b9aef6cfb5c52accdca3161f278d5bd87a61d257fb2ee5d09e3
zf53c381589f043687b0bfe479c17e2fe33c9f7e21953a35d6f23bdcceaff2f8bf7d518bc7ec578
zef0bfd5064faf7c224c84d425cb4fcd88c90a23196574487ac62487e1e41f1cd8a4c1af0ade193
zae81858b052cb503d7ee5f7baf81b9f1f80f096cb771601fb4bfe4db17a16f54bc1d8ef3fb8627
z964bf9620628270ad1c59bafcbec3088755c530ada81692d5c942a90c2db0bb56d8de9ba2551cb
z2b1f1ade6fcf30405a144934bcf5c7ab5f3626884b05f51c627f61c265a873ed8b5eec43300697
zbb0c5c09174a05efc098f7599deab1bb8476b69a3db3a4fbea8e6bc6a45dd6b3c7aec1bffa55f8
z8718ddbb1061eca7a4aafaf3719a33ea56f0c43f42929eb694cd7ad39649415bf994e44e293cfd
z556f477e8e5b1e957a972121a77d8b33845c6beb9c4fe9cac94fc638bf4966cf50ba69f57ab4c7
z11010b0ef5070daefea1744e283b516df15ff8fdba63eceeedf0ec2f9017a05ec537be8021715e
z98812ba47210cce2027717195580b22746c5f7153e97251c978f3a4b2f05b3bba0cfde3d7e0315
z69584a7b6fa0f888a00eab83ed1fb956fd25de78f204a1b0d5143b364dea87f26051821a44aa32
za10ba179e60c8d2469fca5204874051a1bfd683dc6e8e12629dec71ce70d4426fbf18689d3f089
z8fb411ff14cf0f84e4fd7336c04f6c97d44807fca651229a7fee70a07c80815bd75a98564e8fba
zf5758c27865f929daab084ce8c8e678c37694480265383e8d541acd11b2e884cb51d838bc04bb7
z1a8b39e473f70449aa441bf1b0945631359f7c17ff21bacf90d9348305463b8f155199eac94b06
zc02e1d3a74cc6b61d624aa2146b2576cdd6ffa7f7810817918b034f3e4be0a2aac5a3035e4e7d7
z433aa88ae2e97b0666342468809425a35d3c73897062c949815fe7a7d98724171548e7dc0efadb
z9dd409950f68c4c51b51f87872a36b85bea0746387246ef1e0bb143ad15bada456847f570d0422
zab73d6e3c11f05af091f1acf97af5d89016ec086b6438647a3683e7847fe9f71ae19cb2d115875
zca737ccbbbf6ab8237a8591b3fc28f3764825303c5c6075e89b432752a65d1c565874c040a1976
z8d05ebc4ba96589b09fc6d614640ad592c25fb362472a7a31566c8e2457a7524efb5f84aadec05
z51faa569c88a207ffa6567f0ad2f6d34d7964113591f8af3293b5a73c43ed5eae16e30ba2c4011
ze451268fa6c4b85cc482c320c9116613a1214a19907aa92d13cc66eba308a1675bf1a8cef97a53
z6983e40604531527abaebe2e6fdc41c0ed5d3f67105f34ae129d0fbce71d9f41b29f78865b3b06
z344714b8dc5735945f4323c408041e4c5e0ab434f0ae5d99c8981aac4186e337d3ad03607480d3
zffefe53e4e2b1983516d6599cee81e3c4dc1ccd79c249bc49e12405cd2e95c0b0b88a258dd3ec1
z508091bdacf5a495b8dfd9a4acee21752eb536fd2485da75492b62e082d1b15699d84783bcf792
z2d3a7248a7bc809cf40de64420f8fa3ac872359e0366894ca795c478a590ae71b99a9e652fe8d6
z16df231c041fa6fe17a305199719acd35b7a8f96efb997c43a45b153cf2d9832ef1462d03f2c5e
ze82b296a3e1c09f1d6c94ec1b1912978b218f24b591577b7f5be5712bf45a50d474229b85a1f0b
zb6b64be6114cb2602b42e68cce08de9e88b0f4c69f9c455ebe0b252553cacfdbd299c3a976a6a2
zb995484358afbb9526da6d9a164534663a1fb0c2918a02b9b04665bd195a96a0adcb291f00c53e
zb7d3455854028858c3327eda9471e12b8031b005707558a0465024ec4e89cb742dd0080f0b161b
z67a6cbc9209a0e0a9130a41677496b4f0d32ad8a6be00c724a4a8b5ff91e7102b61fe32c387966
z17cf1889bbc22ce66ea632e81684b5ce7749d1548bbd3c134c99d6f2c4a27813236213722d2d0b
z1b56c4db38df89a464696a934aaad5eec90369d474b4d75f33de344b10f14ac072c7e984b0944d
z72e221682511123fb457970b5c84a770edfd1e86ddbd37dd88d1234ddebf9b04b782ab5e71a6c6
z19657b6aecf69c020564ac02ced1c7cf1236ceaaf5444559e0d604810dff32e9ded33cd8d1a175
z441d3321b5eb14fb48694f22d5022ae00d9f4b302905393fbc59665b760768365fb36cfb57d2e5
z1aad3eac5cbc2a75a43b038e33b9de130a2fb2c7fa2f0fc1b8eef2b3258640378adf34445bb88e
z2f76deee43156e170586ee5d082c953c1779fd1667387dc11ed26e26cf04cf9472721bd189062f
z16c0d02e92fe187e5a9090536b5638ed88ca9939b70bb7120fee7e954aee4ec189850ed69aa291
z9e5e4543653957f8da1285743ce80c453516d90b795f4bc539d304c0b980035fc2ce73a5504525
z2926a79df1531a81d0a198f35b5b4e5b9cb34d250b3bb71d6a06600e89a2e1f7a0e46fdb540101
z3a7178be4b6f045ba42a5ffb0bc84fdd3fb0f11560a36677b2202bc6453edc7e2cad5b2fd8b68e
z3343e6e5dd5dec820793d9e6e98d37a864dabc9f5adb0dcd2a3f28e4dca70da36a1e0375464053
zc1598e9a0ace1346dc7d76ea0789f882c9247c10ebb9def316fa58c0b07be50b5d4f528c098544
zc12c9660088a2845c7763af419793175ca31f20487ab75c69e650ea7d8997b59c6231b633d7fd0
z12277b28f55973bdc389bc8b337c3d119eedadef01c53f827351c24124eb06d832d4b447f9e1fd
zc4dfe2ab77b21dbabb9314a774381a5e740cb6c72e7c08a7c90a7470e4074d29cee9013192b102
z16651cec22dec9124ed655805331123c2d976c5ab0ad7b64e0a0eaf2172889703d2be0f9fa23bd
z3ef396fdf6c3cdacdf8b9fbbbcdca6c0393102b126c1e696cfa22a785f37b445b01e680eea941f
z51e90e4823b91b084aefc16813fad0fdb7df7526e90e0c1ba2703165c528b6730ab8c3f25b4cbd
z8044034b3290d80c646bc87a026e9d19d81b8c693be5c263f04831b6a1042327f8a999b3d63eba
ze6aa6daf39475c7667c1858e0035a9c321e7083c89b171f69447422e7a96b034dc53fecc704d8c
zc6fd9ae42db38a4eaa7fd1ffb2035149db871de1dcf925b5142f73245668d698547ded1fbd886b
z3821a6b45383d1e85817fbca314068b747d31e49ef3ded7c7138d4d285a09b57c01243862c1cb7
zda6a3639608532346368f110c27767a2467a7993e6ef90863d561c7cf8ea04ca7bddc02562dca1
zd94bca883ca21d86a07ac9023e9f06a65044d129bc500ad429264fc3be3249f1cca7b7b85d10ff
zac219d9fe6a5c39425ed76d7b315f4d556e606f1fa11ef4c6712757c71362f36b13ae1fd3c6af1
zf569989e6152c794c9ca909f2652e27492b7a4571d4b1209e3c5613c231afab32870823f325b84
zbde360b52f8fa8e52928c9182926de395085b0f4dbb5522d0d9de7596567c1c1d21dba18210e50
z0516a0724f99a33dd798c8b24a6d0d98a7ac9275e8a46912977ff06bb02f50c119b141d1f97943
zeab5495de0a0be7b669c1cd59da0bd16ecaaf9c140c57cb064cbcb27a1b8c43be1d67c94d1981a
z88c7a38341c7ce306370a7021632160a724565c19b33e5ad68e4c66fabb636e4c9cc5876a65295
ze40c94ab5002a3ae986f3ae765089a2fac33e5b5e651883caa7dbc9e681dab823cbba08627e070
z869cbc56752b87da7cc1ce8f1845e30891a7b3bce0933599224f0a5fbedb8080ba6b3f7e113cf9
z7d319ab93fceaefc4043ec9b0b18be79a280eb0020065b268ea16fe82d05681516268269d87311
za80a0bfab2c3ee2c93fb51526357c1106bfc4a132a5b7c4417422fef68cf7ab168a03ef577e2f5
z5981fa1b9af7c047bd47f5f82b815ef2d14ae6a675d509c75f7dbcab618170be903b56ac7b76d1
z6a838c2f54b9beba18acd19a0ff560cd46d974fd2bd279ea3654b15212d0a8853895c11934cfd2
z1d95114343d015d1bb81b1065028840aa8cb7c2dc36a43ae68a1f2af2a1d3d475b2d1e1f29150a
z5736e05f19b3a59a683965a0119085bb3861baeb8e2b0702f7e0b92df5077f8ef82c37f8bd6388
zc7ddb758a058725f0355a2740452809b2588921265646b6f442a0d80e1004c7caf0ef2c24372dd
zd6190a96350378d98dc406277ebc365703e81c19d3e4ced899401565e3ea972c7468570c13bef9
z1fc951ecebe4e2cabdb5ca5bef984bc4d8353f817cf2e9b7d487eba5f8a18917c3911d0ac6f9b3
z54292a4cc2b726d211b2d57b7a61e9082ea85c29fad8f2636064812b7df170d26d136ff3e64929
zc69836a597ba330086d7475dbd951ca590f6851e96dcf435a473d150401b08ea9a0bfa9e224e26
zd97d642d48b40d967f3546704afcbee786425535ed1f34ef5ea02d42a8de1798cf1fb03bf498b3
z0f66f06c06e18d992709c865f9412b081780460e5cfa7d17b17a34d706a5251b2fdda2988b11de
zaa5723e178bc6e5b712b9ef405cb9d3bc2d704010910468cd6d2234332b89f6ab6050379ffdfb8
zbcc3cbe82e41b96442697be91ab1e0b53520c0c236a65f813351e697272ad6813204133569498e
zefc90367c86cd9475b8ecdff8bdfa942f3e3d0e0e9b6ec7602127f4935e3718a8bee998cef2d23
zd6830759912189c42f6528fe0f7d40b173aefa99300b2d46c0d47ba57277b8d9a2743313aea616
z386a3ad71cdcb73a3c353817ac4f08e4619111121580196a267fdbc59b60c578628c3ffb52c4f3
z61bc69ff461e40677232597c02944be002d373b163126dbb5e82c2d48742ec82ccbbe6c981171b
z804cee97adbd95645162b27afb335e8a9182e4d3b85700b2155fc5b93dfef52846e4524abb112d
zf91a3589563bbd48fced65f3837369cf03132ad1d8fef7709a2618a0c3c0af547449331762dd2d
z083b1027e13148921d0bac6398f19720e6ac6ba71569d21cd984040e5b19f42b307820a8afa8b4
z17bb70f9be04e41a5146ba072771907d760143bda2c9c37d66ecb900fe6605129ac23340ea7d4f
zebe1df5e3d63474cc8b4e12bc87640488065021ef5cb340b8cb531667eddcdd12e444aaa9a144f
zc04ddaff0c4273580ad760f99a5fe53b405b5604d86a17202cb2ff5eb539fcdb2a8e8d64424aa1
zec709da971821943ca61bdbdba7bbac740239a20682d765f988d4afdbbd77e49e6a158992fa284
zfd9263b67a1a340e6ec466621446318945e0dad136f7aca5cdc3596a538d84ef93cfe16ac63c72
zfa02cf66ca7bca210e697f9f6e234dfff10e0c85752918c1dd49c4fba620f521fc1885434f11ca
z8b7fa1a7f8974a4df97b705e7bd4f7dcebc0512dbbe82a962aaaae81dd4af8c263c003100d837a
z8e0965404304424064c97bfa86a68d9b235698081957960df3d966bfd6ccf1d3c743e9010ba5f0
z0b7da2ff2fcd723b49057288e6f55b974f6ae829149a78fefcfc83459b7111921776a5f68fae6b
z037e8a8baf54c73d3b04346bc3009161bfd247dfedeb9c414360cf61b3faf093e2216cf8e8098d
z3f76a54055dddda77ea82b09032ca81ac82f8bbf9f770eb49538dcb5a4be8e8bb2d60f27b3aeaa
ze34b9bacbd4c4b9f9ad8f81eebee1e05dbce893e952f1dd22ea27c177263bb2dd72878ae670a21
ze46de04f60494f666f340bbdbb1b5ce33e43e6482ef5ea67475dc8dec6edbde3956f1b2842b06a
z0fa6edc6a5a5066a06c92e685361c23674e742c14bca6f1d04bed741ae5beeac2f9af5a9af7e53
z4f40b2f86473627c50a173b6313730644c7d88fe1317acb73138234d61f987158bb969cfc6afdb
z46e984fec01e361c53afa9348c027e01139071a438e7ba44ca0f2e3d2be5dff993e20cca76fe8a
z18055799ecd6d4fb132331057966ddce743ac62ff59054acf9f5dad8639d53675d6abc96a1d84d
z8cbe599cec1ecb5367cccdb3eb73115004a8885fcd9f7c0520a0496c992fd4a4afe3f2b5eb62a4
z6c23e7916c53fadd0b7da1b78f5854ab67328e07c0f209b7fa8941ce033d82c2ddd1fbb3695f22
zd6edc89aa6aaf58c7c9a27e467148d6155d7c9d4dd43d90c4f0d2107f9c698bcc9c56e46c09256
zf292d9adac5a515b39b05fc395c36a1f1608228a3f0ef10084fb85a6e4fb6e23f17c131a3847a5
zf5653a92f3829c05a5cba0d8944cad40d1e89feb32c0c75bc93d5b093ced6ccbdb3f1962d185e3
zaf9ff76d69f168bcca374a3000c1d213bc3edc1e2ccc3310e7363f163522914082879a027acf00
z83b42735244a840884a7ee47e39f9ea602fdf37ad42b660127d65fdfadca90eb4df40f50f1e333
z4ef69202dcc660b43f97345aed954693c2f53ba3686d14cd30313a9629940f4ad2f1fd07748bb7
zd3ca6b6aa96d575976b449303efed1092b02ab4cfb0b3d77b79f7070b863cf5a82c66f8d017390
z9ea348c3a3d7aba2f6cc04134e3719bdea2fab13b44bf20e4887c9a8680f4990b73857cf68102d
zb9cd6950b31d699c4996e577be08d3a8dc5cea30031653877c7e8436a733387b5de7a2c135677c
zf3b0b732ba0279582ce0621e13ca1721c1949708aa59e55773c02a2733f3c2e68e52b4b9216eb7
z13323fcdb92a8fe0d1fc3e91fda1f489a89db2cdb6a4386e3a4a27899469c431fb1649d71ba884
z5621e54011c763557db8cd0b2cf5e42535289f870466c405ed56937a21e8e1cd3c50f61fb7f5ac
z95eaba8fc20faebb9a6b529d112d1301160292e869a7cc684dc6e137ac37075ab4f7bf2630935c
z93cc24b480340a18301a111fd081300c399a664ec6ecb93fc410bb8a7202f6d45d14279929ee66
zabf99d68a97275e17e5e4a3b1cf0ed125ca9346fde109275ee67b768f108254be1b61e6678b6f8
z4000b02eeda4b27bdd0e74d161ded4321742618f8db5a076df5136334b78520614267762128b3a
zc3173bd8733774538ae81c239bf8453f1b53c0c1c9ad0ba38b737e2f8398261ee0c6bb0150c5ae
z7cdecf3ac4c3b765d6b4e2474b5465598acf84490e908ad304bc8975cabf54f7ffc0475103f43a
z9b08cefdf7a2ec11ac98d8887c026eb1c63973253a9f2320798906342b8f666a988e4cb9ff8d86
ze96fd4ebd76ae4dea5519067bdf4e8f27c5471f85ce5ba443a54a79de1a4b213b28de1f42c7e21
z722b26e9e7c5e01c97686205002d0dfe87f38d0749bcae293cc3714a1955097a5ce432c09c43bd
z5919468873017d95583b353c976c71185ff2738d867863080e68caf678f24f23c13094b2b2c88d
zaeaf835fb872321e15a41b75116f42d20c797afa5e835182414584d57581081cbe4e3897663cf9
z763299f666e3e9a0dcbcc12be047b9eca0e4e1f7e41895603516ab2c5e5cc05b5bd2c8b16f46e2
zfb4a730ea0b3b4ef25e46c19115688eaccb6382f5376d6b142840ce738b90fb05c362e743f2545
zcf6b0ac64983baff5eebefd730a85867ec2c0442c5e76fe829a08c72556e2c5a03a54832cfbf63
z5627dd616ba149b6fb0d1b88a74a668a0652b877544a2a2ad4ab068aa98a5f2539a1cbaf51499d
z5c463383c8953a1a18963be47e8ba1921355546de92ca42c8ab092e598310861e83d22a50a4a93
zcf6b92be095ce1bf15bb48b2f76621f8710fb6e2a6845a185a7446334445055f6f8cc9beae67a3
z9b1a901ea6ca268cc69c60027936bc3ef206d5e4587a3c6db8fd370bf6bbee917a5d46391e6caa
z5e6681fb03467e729b641f643fcef18f09c7b8139c3c93cab024ab09f48ad0c3e47bd9fef5551e
z13472fd2942ace34f1a13d1909c573b415a241264a2b4d4a5c016dacd72b79c5f4fa1dcd0c45b5
z938feb0b8c4b149f0157dc87375f8e09e5f587662ecfed27395b706f853fdc491817d66c72cc55
z029ce12a868d2f814553726922aa7e0fad2498073b9f9f64de8c4587e00bdec458a76cdc314fb7
zf5438af62aedc57a2d011055cfd44fce26d2113c9433516f180542ead3fd7e349713e60721070b
z9d67e5cdc807e4dc3ac6069a3ac25f26cf6b60aa424479b96585d34fa6f37297ea924afeaf9d76
z7a30687a62be6cbd840dfb079c8add16c82ad06bd3f90f8f9ab5505ec607a8ac9ac226a4727dfa
z3ba28265d403b447bf90c5c2c53c3c27ccfc0a28604ed4b8b80c194d630c41528edaff9e39741f
z151a2cc60dea5fccede1827ecbe30f41f9fb97808dc5859b3fee63afa1341f9d2e463a12672bcb
ze9aaf4606c8a3dd44a4c8ea6cd166555e0d76c55c916bc04247413ea1c6dedd5b755f49d1df289
zb623dce782087eb05237bd1045aa279b3a85795cf97b97e0b9142c565a214e9eebb04f04f57202
za937a678f9bbb3535562d00a174b38957b617fd1fd45e04d053ccaf674a5c6c0d3dc35d9dd3f8a
z008b27a6f061e1cb43bf27bb890f8489e8013749131fbe41d03136172802033a0e95313b9e0e4e
z5b5aed80a31617f3d457bbd67ca5aadc6c96aafd57b01664ddea1618e9ac2554c31f2e65e9d56c
z87e528d4873c99a8af6af85aff2646c6174fe9c6cdf0b087bbb5d86f72ab5422ae2f6a881c1cdd
z5d74c51f695f03e941772308ef0db16f3bfe87f8b7a625ab9f68a314ce46458ecc75ecac8eff48
zdf0e4ff63a978ae541997edb20fcca5642446d99fd01ac7a78239ee8897dfe1e7cf9876ac6e3ae
z871b470adbac674e9ea71210f2996e545da8debc07a18bd999d0a5ca82687330bdf2e49a3c14b7
zdc77ac0395ff5c1851549b1b421ef1257bb50408deb98889e87099ab3644cefc2047abbb8539da
z8dda0850876494368ef5175d37f7aca4f76d92d05c212370f50328858f5f70a21521e07cb23507
zd9f6ddf21c851f64109cac85eb3f3bf3fdc8af68b83015ca7eeb1f62686a10e54a1a71c0349768
z8dc630f461264c458c5700a406dbc2496e2777553b8d34bb60b26fcca72d0e41ce0cddbc16abd9
z93a6ee06d3011f7d0a09b077bff1ba56ed1d17ee62c4eaa879bc695a16ce1a47c781974a7117b0
zf15e74b7b8ff0eb04a12c749038bdacbf7109109f65db6504d89e4c4a3ab5a0375ae6d826a2b14
z51f41aaa8ad281cd57c7b71853e7752d574a07571616f166a85fbf3e87f85dac8aaac053723d84
zfee0030f4bbdf54294d19c14bf89a4485031d7deb76782e725d5f9c2e36d6d8bc8a12e5591d135
zd2b83dad93301eb44a3a9be537300e0fce37b0b4096d42b5b6da14ae203f2923426da24d73667c
z8620f70735d1f65719929382b8639c2ea3180bf0e7a09e21f7e0943d92b5c706e0a1d306002ba5
z5f2e3288956c02df1666859e79ebb26f46737dfdd40d30669c3c3e7b646accfc77a04bca2fdd20
zac9dcc295e4f790d2595ff412175f0725f30b94baafc9b54bf11800da118fb14261f4f3afd85f1
z2d54897eaa7280a228c21515e1bcb9518457fedf483a96c4b6f635c65d1f1a33b8c7ab156f0b79
z817a07d9ef69e3d2562b5d112f2a799f8cc30fa803fc617b8d9dafa6c9a324f3b0cce4fb030a44
z5a4a4c2c37040db47b303f0b55096871afff55369ca626bcfa463ba87841f9442d07b8a7d37aed
z902f64611126b353854df63a306979f8c4e1a51847a514a83169a11c737cf88e6f8f4d521630a2
z3ab2de94a89c0aadb10f82e34f52a487bdbfb7ed0d53a1235b3ef57b9ab1bfd7b7b641d327fac7
z36bfd76fb96e24eadff7159fde90523c14f553564b0d73eedddac73c7f88bc38c1bc591e5c7dc3
zb21c06103487768ceed0144d3ad40eeeea6306cd3bb5e7ca95e1bf612d44f139a919b950c28841
z58b395df739085673786775c8ed02b9f477554c421548134f5e9e550da46c0521c335673087329
za0ba777e33202713e6b448b906318db7397d3599b62a2037a487ea1558cb0f5ccd2979f7959706
zdcb8031b4b9c08e32b6711a68e2e9ee9a622b923a238c33b94253dba01c3f925011cbb6de9e7e6
z95d8b0c04e28c594a1b3ef8c458f461406b25981868a4b0d9743e63e07783fa5fd7859f007bc30
zab5f5945ebd09a12fcec131d678fc5c130c3fe6112449ba6a875f47034a9e750e07a793f0f7f35
z7fb08ade778f7afe980c19a6aa7c367217901e82a019c664c553706034750fdb72798f2f2645fa
zfb5e6c29f94d840e2296424c93ee8d7944e0a4f97c53c87489aa6edc713ceb8ed0d1f32b9dc3db
zb2aa86bbfbf69ae0800cb23c7d1647f20563610a54e66ff6341fcb88ae07a3bf1cc9ce77944e3c
z002201f776a6f64a25cfbf9af5729f1da2dcd100043a7d2a2f14307736d0fa6f225adccce724e1
z161a067cea0a7a7d44ba724eef17ef2b0de3211eb02f9a4a1796bde067a15708ba950b787a16d2
zf2e1139d5a370685a928eaff8dacd014a80c92039df65012a129d204e623c200b8d3078219940f
z8cfa8635e4bedd94961dec5cc03896e61a6df6d2f5038c0f4474742404757dca1910a20e5f7bc0
zb80be97f6fce1e781bea9197c83c8c56bf0b4674989cb27cb7a1af551cd6a5560f622ee609ab05
zb3ca5de3b8d118f8ef7d8cfdf598e01a371d051e5b4dea480dec68b74f064c84e3f34d6dba149a
zd73d93a0145c8efa3a6510d7f127c91dd06a109147bad37fd270387cc133f95003f1c8c37f2111
za4e6a627c5f9e673521fe0445f9d397ea4e020c37c006e13e1d04949bf3b48918fa5021b83dd4f
z9836035c5ff264797a6930303093132c627b03da88edb15f87039a7599116da664bc2402593faa
z1aa0a2fff5cfa272007e152b360246f423f740f5eb4cf7c0172731ce5c9221eca91700cdfa0c71
zf5793f9dae868654aba7b4c67a21b8073a6a2d54dfb394b99f2c7072dcd27afa1d60256a5f694f
z619d453489be83d7733ee31b39dbb1f7fde465b99643275471a25d0d181ebc26806d7d3322641c
zfbbdbedbb3f7ea129733395d1e5e2d3fb7f48bba5a3bb027d82eae93f5d607aba38e3a5e871f3b
z510bd4820e309d0720d77e77a9827611bfe7e0db719459c974a83d09f547c7376fec493dcdaced
zda3f224664d20e0c1d274854489b734f5dc7472a043d3ba216b0ebb945ee59ee6eb902c725a18e
zf8d6b9b992eddd8b4cd678af39f26978a820111609d57cc0d6bda7193164bc27f02ab586e17648
zac83dca05fbbbb9ff1dffe9ae9c04a0af777ddacf6086965b71743f372691e84ce04fef57ab078
zb26566f86c7d8530bc30916e695b1bd9664a5ab3e38d31e75f4a097b0011f680aee00d0e7c58e3
z4651ecd37039103fa0de996328897a012aa25114b39d00d021015519aa924cde231f29a5f0190e
zc5bbdbd0f59a0448f6410c818088c9a19d72b6d5d7e01952c4b5e1ada46aa64efb3c1a18128fe0
z6da61c29660e3bb01f02f65fd66de0f9b03ec74170fa1c884fd60c2d937bbd341fb5c34f62499a
z62979a78706bdcafc5372e078fdc539f66c97c19d5fc6400884522053821310ef0da12225f2d7e
za449cf929c388da966fd69d73e731c23eb6952a3f7d195400f4f8a23de85eefda52abc6d4bafc0
z489baf075e803753ba899b834f40c0aed7fad13e967aea4614429276958d46a39f7251f7978656
z36ec738441393256f7d2c3c6dc4086783db5718a4b42df3f138d97364cbc960721c51ede49fe8d
z725519acf7f2ffdb0cda8810abcee27a09ba7481c3d81007f36d69c8eb79a0e5f39e1c4258c9fd
z52b3aad7b4762111248a967707a72fa100b662fe9ffdea4137d81fa2573d809f21ca253de52937
zeb0d9d27f4258c9863ea3f67d1658041cb99fd21469fffcb1ae070b4382ce0831c6551485d291b
ze0a45649fe0ce873cab347387ed0e021cc9f60adabe4f1a16622963b78b233bb77a3ec087545fe
zcafb3b59fdb2904f150f69e15074c3c5a586509f43b189e1acd742e07ec5d3f204d5865a44bb4a
za4c96d03e003e6553c9b93a76e1f38c4588c37fdf662c4a7d8fd98b52571062beb8fea19ee4c93
zcf0aad3efb6b6f2f9dd10474c35a23c037cc4c688f5435810689a09fb35eccf5a8f2d6e89f0bab
z2b1d52e50c05fe9f73c9ebddf390898a163f58ef96d2504f7fe608b3a14c9605c5c700c3f8411c
z86f4faa4d7bf69f6f160ae3595a6795b384dd2bdda98961444cd19d27dcfe6a7c7ece74d50b13f
z0afc4a01d626edffa1cc081dfc615ab6ea2d4c0a18d09b3df50ca4524bbaddca22aa4817671ec3
z192c2bf943ebf3c5c31233a332cf8589e80174662319bd67e0b6a199afac41cfb5896a1c63cf0b
z04a3cb0889ec86db78dfdcece627992019c66aae834f1f33d368b99b1b844e854b8ad09f96271c
zf9e8a2c66c7632d480f9d1974e3c6e93306dee3e574a464e1f20f3b5a1e0ed2e423d5f874925fd
za74e20feeb97b442e6cfddab48795999c84c480744774f60f5b3b0c09975984576f7f2574446f7
z1d5a47745f5994ad161aff25a0eb0fac1d55c44e8fa1cc5df13457681a3ce86e45dd8ec7d57c34
ze87fef55f400d5c495b5b489ad53f740a73375c01fa8ae6418152a9c3aa099d877d9a1da9a2c92
z6678e75d862e59c8e7104ab0c043e5e0e957fbc383351006a987a8f061dd053d73b5768ad18b3e
z91716beb2d88fac339332ff33da03234d3192663340857115e226653f2200e55fcd2dfa881ec60
zf6ffc3152928b491957317f63f3dd663a18ba4baa6ab3f9f47e7b5466ee6ea4e7386b48fce121c
z914e1fc4cdf62002709ab8d922560790620b01ec0f4d59ba49150fb94fccef8cb9c41deecebf7c
z57db46b9aca81516ab5531be64b076904bb5e627641b78fa28e026dfe06889e6eb166622a41e6f
z8a3e3206cea24e4f4be9fcf5f17ebecfaf10d9cfafad85bab1431c420e5fe2d6f75f1a0b066279
zd43df4ec9323babb43d4d128becf1969757db0984e2f071b72dd2037478af47b0d6ce9da3b1632
zd13d8112845099b59b02e20df7e17aac601aad7cfaf5e792f4b9f312cf299beac97e6c366b42fb
zf47f12e4f3e454416e4d309b30c934a5abc1cce03125f5fe6ba2c57dac73756dea33abb77cabc9
z45407aa1a9c3f26f16fd7cbe799740a6acaa11e1897bfe20c47146230c6c6caf9829c65e45ee36
zc2d29a61129874012fed3c50d9b8780c7f5136dd39a10334fb671e6650d68bc187c352ed156eb6
z1f351a82955e81de00a06998d979891a05d674d6bebbd40c0ef870520e22336d69aaf5a39e6293
z3f66f702bf9e155a1856a2e5d8babfd5212765d8fa20146d0fc0b9e63c20c0e89eaa6ce6e6907f
z37eada6cb071458b5509575ee476a73893a24b01e31b539e9e6a9e858697574ceeffac41b9d6dc
z80b55412b1f18b41cc8a07ab600b94ef8af4c3b8aacc45787eaae380df13e2c169d6a5bd59b9af
z1ce2b53c819717116056189370c938c26af591668ab3d6458b8dd6f24d9a74c3fc7dabb8c58401
z3014d5690a57052431248c974258b0fdfc242b13353e250f3093c0ed2ff077261ffd8337a45f9e
z2d9567f4db74406cf6d274039858577687b6aa355ca2bcd3ae0c83bda2aec3e9d53e87effe55ec
z5414b16765418b9f838cc642ee6fc12e935d9d122cfe149cb5b4865b48648cc6ed2c5686b91c64
z6cb6b48f0361f1310cdd760f28a7716e818f45c61d71bdef46655caed04f125f23e1f325698117
zc39b1228d16e2c24e41ee35044ca793ad91ff705e2ebd88e10825833c9acc7056f5af8d4a6a684
z7e102451bb0d420237aea59b110acde01a6e409eba044a078a7545b76fa02478ae1b4d6c774a2b
zafee14814823cf27157071cd448cbb23410c9a249b5001b688a69e16b5d079ecb290a08f635387
z1e2167c0a17fe4b2e22fbcd4245047fabbd5ad41ade4318a9258c8af6585c4c674b4b7c8fd90b2
z4f39958d8f5aa8a134817725f20d857cf496d405479f496eeab6f62fc0bd9ed0e3080796e40a8e
zb94c295fdf4665b747fdd4b75064ad20089fc01ed1401c2251b2b9a4271cf777e683af75245bd6
z77a8d3129478ca885c07195cb02538231de641dc3a7a5ca1ac91177ac56b23debb9df6877a93f8
zdab496c76500957e75cbabb8b0e0adfad23156cc63738bf1305feda3b1462ba267066fff48b0c4
z3dbb4732919b27335e0eb217ff2626e3a088a93b005709903d9efaf8af24ffec5429550712de01
zc5b1efb583836be5a4eb585bcd6913a4e295d9ca3ec80de82b78e61a205778731fe4ec02d91c4d
zc600c8bade59052a32b47fa346e6ed74c390b9069e70124f8349824715b8e5da195d5a6cb2235a
zd0650d80c9aa05d0c698f4016eadd06bacae4a41b5287472a996b68f1d41fe06e52618f2e52dfa
zee38b5fca457e3bd1e5bf32cd365ecc8993c4a834f5130a0f4d70fdcc02717b1ec972bf4f623f4
z201d9c91545921da6e2f49186c1b2d498a24abaffbd21a286359c0aca0b69e54ccca40d6928f8e
z9a5c9e455dba2ebcd06319dafcd8c009c350e1a9a539623633716978440cfc3962affae54aeba9
z7a7272f02faffdf2036dd4eb3674d1487d6c793a5005ed4a9bb7628e62d2022c7d8f68d84dfbca
zad44c0ec610e324b93aa3dd0ef079a18a82d6a5dbaa3d4d181eab710eb62d589170ff6d28829d0
z143f80745bb58e8982a040bd4c458edd2a54d7e032048b11d444f389655468ff6ab64f3f528106
zee7ba8e149ad979853af9d9b0e2a294165f5f681113bfbd0b3cca7e959a468ec2f1fb130a78fe6
zece9aa7876110aa6ae855748296978d4e6a477de5082aed2386abf8303c454a4a9b6ce69a02d8e
ze40d5d67f1eef1b2653d17a3486817dc3f238c7d97f5c4c81ec5e33e304c2150ee96c4f759dbe2
z28eb2bd0341e33e299292bdc9e93be9bb9b2d5bffb203b5bd6c186d1e503d1716cfa33822a8f1a
za34e1617feb56d214939392c996d11c22ec2f56ea1373634cca3e4cc2e2f253ae85d6a1cef9802
z0b1b36af14e03aae7032b9ddc80f6e8972782eb275d813f6821c2fd45bc544d8c9107b42e0ee81
zc80c3c8cdd8e99e11eff0f66b758b6778b14cc202e118847a15b60870c3fa9c127715a0fd1eb78
zecdf53eaeef6c54e2f88d410ba83d1679c8e8d943b884b2a1d748948c8f02eecea1000c473a4ea
z57cbbd91d8344bc6e5f4048def33e3a020510aebe3659e9397b4cbabf1295a32226aea1b632398
z79a701dfc4aef9de84f05e9466d5d202fd04fb225af50dac3af5c22cd57f4856eda13b958063d1
z3223ea67b3d4289877d5e923f62ea5eb128e6231f1f02745bd2f531dcd9306e18a9d2aa1f6ec1a
z221b9afa09dd38099f6c6e67ee68ed0879372f999ac65783b84435f93bc27865ca55f9c267e6e4
z1530b023e0253571de6440e88d9d5e13098dcd87835531da6d2b1327923c11387b0099dfad3d84
z81d510b67b7db9eeadbbf646b5d3f5618b94ea64ed84377bb49842644236ef3b838a1127256cb6
zaa6e1f9904422bef9460abbe324bd38c78fe970e65692f9ed6b67f37c2a1dc9c0dc62b490d0621
za5363f7536da104c6d9dbbd575ad8849b276b1bdb735af13049290667c0f6f9ee8e821318d4ead
z3456737e957a8ffd8dd8ebfe3807f8557f7aa9f1db4343a9db6c52e4b1a7c301312c098353cbdd
ze08d09922f9c1914f59fe5cc8bf803a9c7654db0c670af14ea1eb9f1481f2bf3985ffa8e3e537b
z7d418e8309f07a5eb526824bdbb54c6fdc5caee1edf4f13e6ee26dc9c1e0764e668c717ae670d9
zb87b2a600b56a36c02372de7ca9fff42061eb5628670738e8b2bb72e7dfd723e37ae984d1fc700
z33aa4fe8f39f49c734802fcc09b935e0220de39730732e16fb4ef0ad57ab4c63f9b6f0a23063da
za934e498681eee3ed9fa652c9c52f01a2aa4dfd17dd48d0c9f2b15e4f342f11d3f631f2639bd3a
z468730b9d8a778749c028deec14bb861aa048de7d5fd8dab805a555f13db8a18199d1064dd9235
z65d6094b500cb2a586b5a5bf1aad9a52f8e95b7b3f97b92be552394af8bf30b3cca8f6fbe8b9c9
zb3fdbcda7eb2f039ab0ec47b79f2509afe312da7d8248996c95fbb5a27cc70bb701a6d4baf95ae
z4f44de9e165225dab701271a28457249ec7a3cfe2037c4ce5c04184e4c03e7c9f16f5a7a35d492
z7c7a9f35d8a912c5ec04b2192c97eaedee6db2acd1c334a9bfe9c81481f046437099da99b9adea
zf92aeb491d3a674786c491cca4da65a34451052fbef05519a1941cca7797c512f773a7f5dbc29f
zb5a9871c06958919e18d2da5ae9c5ba552b43ffd71298de12fd3f8ef8763cd8eb0bba5b3f744f5
z7a6bc1d898d7b170abf1e34df741ffa0fa7f233ab5dddbc0cac93d131ff31d0256e3b20af9abf2
ze601430df3430b220919c044d4217cba5cdd0a01a7d3323a796728120655ccb13262ec7f720b37
zdbd968491f76ef7ef996e2dd48dd244a75a438973eabe7bc80d9132676f9fad93e74afaa5c22cd
z71b9b2f3ac5daf44ddf30729fc93e7a84c95c7bddabb8b135ebdb0f1180b6e03fd6da55a6095f7
z0b0d27653bdd15a47453d7dcd41e1d8bdc1beaab14d07bf401d5940894cef1e2a6d1b0bf833423
zd972334e5894a59abd74b774707ab6ccde796224034dec729c5a2b1de6f42d2a86958c143648f0
z8c7d482c67c1d2c5e687cfddd9957725a88e60acfc592da2be7188e3102a53fad0852cff79ba3f
zf0f8b3e5f09aac31bc5757f608a95f636fe1535035568246b7e86228fd7fe8fc173cf83881f64b
ze4e8c42365a498e9f6f8191a7af62c4054c4cca292912001523411946554795ec1063a58e9ca9a
z73124f2312a42781379e57aa51f5611a7f832772487e6d8e497c6c9d7583d935ad0490cc403172
z1e99f276cc2453fd4c3527019a134556f4463a9aa9aac453ae890fe7885a588bc182d38f2e7932
z256f765a468bbb4c577a91f46e0f97b237264fdda0d25be71ebd17606595798e92299baf73fa7e
z64436b676141fbaafe80ec3d190830ea699165a043003e0dc91101812e0640e75ca9f002eb6ef4
zb0358aed66c028ae6d6b8bfcfe8f9e9eb94cad8d564034c9a0de75d779c9e0cbd1cf054858bc3e
ze103ed631f8fee607287bea78f3658b50979ee5126a7d49aec453b4201174b1a1ee8ee21bc56f3
z7df6a5facdfe79bc3f474d5a43a74dde0c91d4e09753c6eebdd6f1c0efa414f1fbd0f2fc62eb29
z157dd54e9d51d2f49e485d24b2fa0499aaf03ebcba486b41e10a0b5e3bcff34883010716eae454
z38420d9da47a594970787462406cdbe05f6808ccc43fdb28cfe21b48dd1e3a14cd38dc933f7832
z96adfc55a106dcab2da7af149a7ce5ab14a0c3999c3afd04fee0e9c9d8b70dfe4ef2ad57271e47
zb538fd3f4929a9f665bb63be04ed4cc3756c4b3bc242e5b251274451d9c61ab0e763c81952fafe
ze2247f4edee7a0f4bebdc5eb0328e126a5823ecb92c7d23db130179987d4bc274688fe4f708944
z9086d33d5714853ff55da8030a1ecf1313b916437c8c4ab6f4e85364b8abc1a6d6134f7897e557
z4adbc3a52474eb10717f8d68c859bb1465be8d4dfdae2a79a952a459049f04c5964d5a86427c74
za584550c92d60726a6206f74f823e0460f0c2570d49fa2ce3e40836415091955bbc5f478e37186
z0bc122d6cc88b95b2b8763580bb97b49c03311968b57d9dc94f8609e98095c3718c1e3699c3207
zd819f9a417e52660a008c09441a3ce4872e8cf76acf954f25fcc9566faff254b78717ad8beea28
zf09e5e1968739630baa1704e5cbc02c1355e008cb9245c2a5455d36ffd5e8f045bc236a50d7547
zf8e5938ba53c3d99d6afa3f65198882bf2516e3e227166078c74b3fb87a3bd6e3b6b3d9cde1a60
z334b6d9f1a6023d46a9d86cb9e468b65491068d745d1b9068f28311e4d1e8a8c85d7744263dc0d
z808323ce1506ab51a724e27aac20922f241fbee25559181c2477f16cc9d86c809927b0c315831d
z6e1ab1e7524f31e563e21adfe9d262386491210f720cf275969bdd5ecaabf1d1e75831dfc525a1
z7b4a0d10901dd3e8d746d02d724bc9fcd31f2d215bd69425234436e35c013e59d0c42e7c75e69e
zcb9d66650967eb3b5dce9b5e2803b9f25a1b5f3f576793ff948c312f46d677c0b058011c47ef24
z551a3b6424e01c2bab2f86c50813c7874aac2a9a2972c74559b1f06f557ca93c9de8c194357b64
z0f69b1f0a6842cca6127c019ce565373afc1fc829483faef1b88d75b87a61ad1abe444888abe8f
z25fc3e7a0b6d660ca64def557db1d960575d3d55bb8e9c7be2dcc6832f2f04cdb388038ca13c1b
z19ab0512be0ff7b5be206ecce394c8516437b0f12704de5370e2500ec0be2ed05438a6be736e1a
za106c3e3cbce6c956c7ee0a7d09ad16918719145ce6b2636be3423fe8bce2fdbd4de7c9b9556fc
z7a69912c167615eff3a46d840be891e95bd806c22b857213356a5bc791db4251f44205cbe60143
z072570bce14957c59ecd5e1954b0bd9678b10fe514dd0b797e1a0a72c4ff532d4a858834f728a3
z30ed9e55524438fd67a15a9b2a94ac4e513d829f41fc4117df1aaa6b1e8ea652f59a467f94954f
z3b0511236c9a3bfdde7c868746ed5c11257a115e21a881ea9a90fec19407f9dc5dc1556df72812
z76237a0f60dbe06a434c019aa974183189ca63db9b5b364c79b69b91b3b429ec5849fd500626cb
z4093907fd2cb98993b08cbc97866fd4329a32ff0855fd2e13fb9c0b54beec2a3a6b53d4c03754d
z66b28c7437dc2eb50f5b26db7806ec2527fa29add4f4735af6127d4f5730da9388e4d321136367
z24540dc100c391da4caddf9718434ece614598f5f2e20bb3d02f09f3713558ff0dfed595eb7f23
z1917862292efd83a252b7620b2f659c0b2c1c218a1ed166672557f007eafe87687c08976ebefd3
z14cbea72c1085f7ea331a06323d999be3c6b86a2d27ad3865db8c6543f6d9307fddb1c6b732cf0
z9685b3a60b6d0692cd0aa1b8affe789da0de52f3020cb7a2321743e285ab0bb3cd6f58f11af7b5
z525e1e2163af9b6a74beae384cc0b8241d36a1739a311e82138c497fa704f8912cab12f1f9a389
zc2014c0a95350e4d5acf571959761baf88b40706c02d389844f0c34c48414b19f6a2ee5b029c54
z80f6c6910aa47616a23f672be184d2be4f4ab8bbb2df4c3beb90ca8cfc7998b1bc99d418d62b96
z64d23099a4dbba4f634d4b47ea147f71f3c404093c708cc1c5eb95803c6cd0f02524236b1ff187
z3e9b187c6369a4a80617d02a411de7efb732a047aeaefe7e79599ac5d43ebeb5685e58148db836
z074d0151724bd798c24c86b32b266df4d6ae5bd8822110ba4002f65eb7585425c278ae3cc4a85d
z1704cc753f8980b5e00633730bba15f82ea8809d9ce30e0524c11cc626ac0f6a68cd013754bbf7
z5184b1736031874ad722d76e535a597bfd42e9589c988549b40eedcdb8a0533e622bca52314ba7
zb0ddb886f2c6749c13959357560a8c0e61ec55cf4390ef3def06e0fe9831774a9135df13533c66
zfb38dd22b45c029c45c54f2802ad175ab5bbe6adeabf4eb8703dde1d3a3e2d4a6f6667029f93f3
zf4c012006b9acf3b5b08a6a96b9baa853cff69a8af3c76ee71aad824bc138d54e3506953661a7e
zc8296d6569701a176ba01aec9d76e1e4ce033a298a067e096d7e33324846ba0e34a10c0ab680f9
z0899fdcaba7fea44cca3dff99c63d6e21da79109e8f72fbffc0569db8bf55c9167d76a5fc2a28a
z4d1ce772f806926699c9443781af2ecf75b14b6e9e7573ef8297a537a20168c596c4707662b04a
zf378760a9aa241d2238f4f3d99247a65cbff3b716968c1b6b4faa7f387ec7726a23391967412e8
zd6bfa4930acaf62a922f593ba1cc21b20bdb22fda5231b8f03c181dcf1befb292bebac989242aa
z74e355d8356e402287bf13da875856e05101efb1be701c0fee19042ffbfeda8799ff2ad2842587
zdc2b120317cde1b97093c95a91513eac1bbf642b3f9d1038017f29a934820193e29a6b56980a76
zf474e98e0580f95c4851c0bd772841ae12f63b75a7157e5e694722fac14acd473e72968cee304b
ze4d49e26c24ee614cc27dd56baa2837bd48e13a78a7f7c278ba2a5a68e5b4e346305d376f16c4d
z5865411d3568c821773902a22ca84b5647f41fa6eadb61f4b397dd57b8cbc76c5a7697f4d24c02
z7acb4c74b429af7dd3316bcb3df80bdb3dd9b2ecb55cf22182429aba8a8e0f55fffdae4af81176
zb2a63bbacce41a44d9f89d6ecd5463978eed8871b351f4ad1bea9541539fdb02432879c9aae57c
zcbc67459f2289da034c0607083a9323167f6fb3cb4ef8f4395c7e0d5c605e6ab17c23f9cf0ecda
z5990400414bc6d105ec8583958e60cf0258f31c8eb14719e55bafe685ac3a13ac7038915f27879
zbf6f275f7717481f7faaeea30b24adb8d66643e115acc1421a46f0d93668f012a57dd9557443b0
zff3488a12508c43cd8ee901dd503ac16114d90ff299e535a251e6987811e32c64aa6fdf070439e
zdf40026e5fb7f4c7628ff8a1bd2d591665be0dfb9e3d03ab3eb263999f3d6e0e9acaae0c49ee8d
zdbed6d88008e413791d838c531e30636e6691a0824c6d1c5b3d96a90bca3853e70fb1f43ad1f0f
z6e9acd5b6a6dfa29b6da7a442c75856933fac520db519414f8760e027c6ddcc026204fc653f276
z3656e6a26b77aced4f1c2f49b4c381d69d1faac506f4559a1e696237f9a1347dbc66520aa687d0
z3c4a853d3c9af5268176f5555a2b505a3d94657c29c74bcbda2901f79d9332142619008713edbf
zd18080f633bef990efded33d2c24d594eac11e14e516a1d28fb0cd92fd4fde503d5aad30c28971
z986caabb163642901603d03536b400872a27ce62ec99ff3f6bbc2d0e3ee34a054c543521dadc65
z56877f55a1170e24309d144aba66f5a1d52cea1052d9321c6defc8b68a84390abdc298a01559d0
ze9f40ebe34da2e2a3b31ba6af09fc51e608a8cfa148fb8e5b021a06d6b3cb3dcc848b80090311c
zd3f59e2a16417b665919fb6c97e7c927b8d357d477b69ecd639a266d9ac00123b50b7ff583a291
z5d1b823545799293ed4dc95d949c38a5e8cf982c0851d51bb92b7462508bb7233273a72bb77344
zc6bc29d82652a23d3259fcf609718687ea8cd994954977b3708efe09ae9c63a645f741b27c5524
z1287b0f0227132eb04fdfa41ec05597aa039b8dfa2d12b3bd24e2feb9bb721a979ef22d7d58a15
zda94e13c15ae00b8085c383f4932b40c46ff0a838c133926a17e463e5870af44bcd64ecee058ef
z7efb020a2d0726520660e3e67b98e0ed537dddac19669e6b58e51147a557c8978e88493f80c405
zdaa0162a4c05678bea45a3242eed75fd097feb8817e1401c8224557d8c61b527ef5c4ade5d0512
z3f36c91436b87ec5ab7d1f1892f0a06e41b77201733f29d09b7019debd08dddf0e0323fd8050b5
z3bfb1e16dc6a69a534242c74ebfddfa560af6755879047accd1b91355646e81ff871b3c5a43708
z3554da998534d9686e6cec1d6b42a886ee663f34c15bd1cd21fb4d7275623154210a397fc8a172
ze4ea423d0b360b7be01a63fa88e2cd18398e8d68a6e9a8b4dac2924de986bd093c7c667957c270
zf5f930aa53783371884948c729f0ee3200230ff79ca827293f0e242d37ce307bafe90b8cacd032
z9b21bdf3b64970a2007f7f046c961a34c77b22ff920bfce2aa8508faefde23bf51e9abd9cb4e7d
z640464c3dbbbc721fe0bde8791c701aefd8d7b067085832486f6f54e48c93b16057ea2deceada1
zc7775d642c4a5be86fb66dd7123c4d79d3d9bc2987e323f4f89f42b489c1ab4df9b1522462a1e8
zffdfbf952cccac324aabcd4410080b56b72f55865144d4f6311195f15f0fb14872f3fba3e15db4
zf7ae6ade8c445bc95861f49b8396ffe24d4785467435a8decb05792387aea00fe166d921184925
z189bf2076b78a7e5bfbb9d643bffb5e20c6d3fdbb1b15b852aff9577328ca3504d145684298d6b
z5872d921bb98169ca390df94a32b7f06048ea90e0d367eb7770ea242ebd8badeaa5177b52960dc
z1d37a9868acef0443e74b19ce80e22522f857b7e1d049146c1d0fcf61981cb7b89679767541f7a
zcf1c1bca9ef7cf5592013b82d9dd84809ca545c7bb0cf01894182cd56319c6b3d04cd11d071992
z021064daefda8b635a1f6b7e68a2979aaf6c5d4b38dfa4b57ee06d779f78e8bccdbcc8a02c8b3f
z0a1dd9f156ea23f0283a27cb907df08e2733ab127328df38769d26e4867bcd543a9faaa687bcd5
ze3b0ce352705a8d34907c59780e478c678a401812dde8eec46792fdc9d01c6c3490b101a907ad2
z0ca7a5acbf4752edf911022b99bd49b5b67383ff98a9fed2644028dc70d6631e6af8dabeec8ba3
z39dfb29565d10522307f19bc71921b13e5459a5bacd267202413489c1071451382ccffa1bd82cd
z0ae7ad9f2ca83a7ad2cea12f84f5cea8fa5af870dc31a737f898c06a867ab99e325d3d3d1d2838
zddae552cd1b94ee1ad5afef056505fa52a74763cc6b5212d7fea57c3c2b162b9439e6ce6ce200a
z91042c2e9a0ea4a2542bbc58620d3ed03478d75d8d588bbdade01c49416ccbd38d04c0e2d690e9
ze9810f0acfa8649e4d6c510886e03f55397de5d1b9d6c00255419a8865ce636462133e0572d47b
z01117d8785bd824dbfc5fffaf2fe87002566730c3f77dd5f72fdc81d9612b548f0f71da38d477f
za2237eb3b217ae5ea0988d9db627ecaa5f6825c3a28f795f1b1e136c3ce64a6d42b27bace2d639
zc4e0c75be8db517f37bb9d0cb9385516a5e5b6729b37c10e9712b44988c05426141c02dec97495
z182be4a2ddf7b327b03ab4c924643bcc49d76ff0cbcd506c7abd638d0f075bfcbbce781c99c255
zbe8a96c3a7e510a4ce5e279f57a62d798fd882ab62866533fec62b959a01bd3d89fcce60231c8f
z0706f83e85df931e2beab19c9b6bbeadbbe14c18f9652fb53c944e922792a6e4da939a71d18bb7
zfcf79cca9a07929c42ed7c48c60728331c409551bf39cf68f04cf102cc0dace318c227ce37a5ef
zce349b38892b7b58164970ac82b5d9285b799fa3e73ca93155f3b6eafb6095c74507328bbc5835
z90ad94c6d6badb5de401a7e0046516568c1ccc7d67b7884fefd42ad72ac38dd05e3d0d3c6258a5
z2c75eec373a829ba2c521b30236b44eedb1f1791c129dd95cd66e2dac8bd64a90d749ffc15d454
zdd9c711120cb19b3a41ea21b5517aafea8d5952e1c53245ed1415639274c3d24e69f6d84bd2712
z8399200c6c70ba5edb2b57b05bae4bf1331457f0a95a42a0423e4d0f623cb54a98b1485c2fdb69
z171f956f2ce6399e3f06be16d9f1b0c9bbc315c52443a97c8dca031eaf7eee9ef46902ab78bffc
z86b0fc33dd809117aaf8df57a848c39e258249d1ed51d2df347b5500af4c9c04166a23f3d22dc6
zb4a5adcb0154c3d1ad0450c4fa5c39f4f7c4e1299fd8310b5c99036bd4e65a5d68774f427cb1cb
z05a0ddba4ee8860390a02577223a31b1618408386e89fcd23b6aa80131f70a7b1535aeac55f922
z780dcaf074ea6e36d303afb6b5785a08f15d3c6223ea42d1e3984132924aaf98a99e66c3d209fb
z755523afb7807e4298fe408490ef8e38ac1bff34de1f4e8b80d086bb1bd09b331813d230ed4871
zd5f6f26c692d777e8900e9d68b010d7423d234023bbb97338009767020b59af504e8d6e6a076bf
za822faac57098b79d40d9d0d642cfd2fb3307527a194e37c5e48a38bac46171c980c50059136fb
z21d0eabfd8bc5f8b75250aa00a3a374b26711036934cc725b7f07a9283c137043a85d1833c45dd
z544598aef39d6bad5beb3eaa9d57c3ac608b85bdc019bc106504d0aadbcc9118f20538af67c215
zff271a9043dea4185f2f63d3613ccd2efcf3d7eed5e667314c2ef6b3c928aa7895ac5bdee292dc
zb6dba11b0e5576fc32e80916c757eeaffe5b09c2857262b73edecca9943395f8e6483c1fa4c27e
z31162c5e881c03e9ad97fd6fd4d96515eb4c95d20a5a1729aad5850ef38afb10d1e3f3d4b32608
zd9f04ab956d7359dafb1b3a78029afb80aa39abed47e5ada5ba8b826e7533d5914de302a459669
z9fe7a653c8aeaeaf839d42b609e2d9de3c7a1015d8d38b69c7066b28bed03bd80a6bc749240d0b
z3f3c7eed9ee0d180f8f3820fe26566bb82dab2ff93d0fe6b0f81145d99aa47ca086a2e702b2b61
z56ddd19fc07e164fbc2610424534d133ddf6224cc8c3686eaa16819b2610e7e88d01abfcc1de6c
zf9813b34801edfbec2e90722da2b7530cc455c73b2ed8d342f2312fa9dd4e2b7bea3c376862b9a
z70debe859298ded422f4b03e6dd8cfa142959c48b6656cfadb296941745b00c87c2ebdbbda8796
zddfb220d84a9546d24d9e5802a27dfa51c7cd0a578ba360c9981f93256bcb8230c2238297d945b
za6b1ee7fbbb349ff4b6388d58f7b1d2358e449b8a2a0f30b3505ebbccf9c4a2e4b3ede30bef6aa
z01d10b5b1f1df6e1a219de0d3014e9e979b74155e34829c81caf069a5f2ed57ec96ed7dc171b77
z0a7c55742667e38372f33c21bf298b70f82efbdba8f24463d271000d45602c71fc63e2b61ac985
z6d0dd81a8b1bf427fbc326154eb07c4d4f06b1bbc6f88655c137b634ec3b2cc10b2ff2ea794614
z5ade4e120a5f5f194d26ac511f4ec5beb19cd735f945eb947705b8d6337532d86a2a17ae9ce707
zd90766e42a31401d860aefc78ce8e114d2f632c523a09251df3d8c4cc735ecbb7419d223f768e1
z4b52100b979c2eba17cca1700a96615c8c3c70a227c091072dd146377c76ab55b45948dc137299
zd0e2191e85179b0633c617642179fcb93484f1a59dc88b9510c48815433e35acc8fae25eb459f2
z96f6f5edc42032247dde8475508377ef1442bec63597c83403f817ab98d485a1f1ddec2675e3ec
z64dd299db748d3aa859c6d40b904be44440a443d4e9905b3bb0a0e3e84f7f11735b6c777913a6c
zadf9047a220d230abf9258ec84fb81bfa6977d29e4df9180f47b1ce9f3722a35e595faacf55f09
z06de0eb076b958d6d63de3a78b913dab117b66e1bf83616aaa194dbd31b25ddfeb359a6d837f46
z2c8a851ac237fa8e6b1001d8483ad61491cc1256c3bc0338c396eec4fb365dae4ecdbdc1423402
z2933adff607e22340d0dc25e2ea83767cbabca2d1b55a2c50b79266daecc306a34c7beb5b52bc8
zf7964bd28872c2b8fadfa8cac24da9572f32eae4b31b8dcf5a24d9ed5550ae3e5229bcdaf73da4
z7bef11d669841908061f649bc6a7ed24b1a6938261073497b8e7c6a3225611ba36dca6a0bef245
z439d3f9421d6c98d194788cacf0b4c413f85e0256908a570a531b6861c8d0cc26fccfb33796371
zfde49ce8dc8217fdfa0f0016ebc040de23cc6254150eaf60b06c24f3ef70816d45f8f6a33d98e5
z2e6ca8f4b3247a243541bffa759ab20911467c1ff9e24ce86be25d7864e39eb3d7b1e47b16df1c
z35f66c74d75760085bebdc8bc24248fa87bfe615f365fde5eb0877356c1e747ae7e845b1ba66d3
zff52aefd57b0b97e0e709af458d48197a509ed1146c67f0b21450ac8d2dcfb83003b40a7510b19
z48ad1fd9b5aa6f8d5e2da5716f86c88d11e80827f5433fa3e8efcae6f08952ef03cae0552d8a13
z42192c4331fb80bf2f7365036fa0b7866379b92cc6ebe8f05e0198394d0cafd736b4d681f7a164
z6fecbbe816c6fc7c65205650997cddd0accfc2f9d8af42bc39066a9c1d37d2bc2e427c4ce66010
zc812248dd0fe0ac935476338f82a5ebb071e8670f07868a7da585f5bbad9d3b49db2a39d4de118
zf248fe05f71e67c1c09843a42594436026a8ee856a79b8e2e84f8fa0878bb07c4b6c3bb4335168
z769bf2f6c607efa1df011fa0b9548a846d2628baa554612219619b9740511ef8498f2d78d0b4ed
z2c792d2cc376616a3a9890574d479a57711764195a896579e1e5e29880e5aec64f35a81ad396db
ze4bb2b58e6a96d1a2f507b5ca6fa5f5bbcabaa851dec4c2bec7f648e3b20667362396105fb208a
z1b6cec72c56a5a7e4a24114822653b0ec6cfae0f59341fe028fe7373588fcee11c46e9b0c2159d
z6cba2eee37f402161f0ef5e682bd25c3c726cd5392ad18aead9e7dc16cebb7fa9bd7229247be70
z0fd9af218a94f6cf126f7947a41ee2e998c5ad9351476953aafd3930ab8466f6b8e7557563a6ca
z426289d5baedbe8448d21c1f0fff0fdfbf987c6bc06e9a5f4ad1dc87823b919f2e7ba60848b4c9
zbc14a2fbda871d238e182bf851e2ad0cf39a9440cf218d8a1137b51f1ecb540ea7c09455f5d4db
zae8ea89822e4fb117b2afd8a5ff9ca9e8d2b3953ec3a82d6ac81b7fb7667824cd9ca327996c00d
z77282af9e69d1df9877a680af2419f77bf4074e495c127dab7132117c9c30ea104e98c170eed27
z889cdf801fc3b4742641336c3b94b31db38781ac95245fdd9981707e66fa063dc9f7502a8e247a
zc9f1bebee9830e78de59cc0cd030b4c4e2c28999ddef0cfc4e484be6c8b8dd2aed3584b882d988
za3c0efbc48ec5b6f0c38311dbf34f211e3355465666e3e75d2bbbe1056f67ccca3f6a53287d40a
z0b4997d07d5b724ee3e0ecc643ab9b45667e23e87295d3b73d125016bafe03e5cb18937a173293
z3d9b7d94c2d29c6959504d12567e7652055900d5e7588e7bb0a99f7f2a26c446ce15b54bfb9d0a
z25ea0040483c96757b31f5a920b57264b634021581dd314039def26b3df77ac66921bb8795b89b
z166f9e3b9807b20bb43e58977329eb356df56b258b43db7bf65b4379e99a0cba8bfa6f2b0e9efb
zc07aa109c4b37e9b76b73622baf7bed2aa73f931813af749a79356e28f5fdb57487d8f614d8d3e
ze2e02064a6c5f28f39aff124199fedb63ad297f39ffde59fed59828b15cd03c80d7493e5e0a11c
zf6e9a4dda429dcded84c89e85927c05c617afcf92956da27d3360ab8f9b99babec943d28e0dc54
z2e3f63ea590a78e826782293ab624e2935ed92f93333ed2338c85f595991f4bda670ecea1eb5d6
z30e9f174df8a93839be68b3f606fee2f4bebb08c6b95ed09f5a570694280a3121faa9d0e309f61
ze4781f426ed1ff7129473e319a01321b3ec110062c1da850dfee4b6669245045df35089ee46c7c
z190fc8db6bf3314f89f2bb9dd9b0966c6342c1af9dd473ac9516098211830523c5e0a520961375
z3cd4e0d1405995a8f0a18df7dfdd3f339dea22b2a9e661806824aa062d66a486ed3e26297f27a3
z2f3ff9434cceb7746ae740e8230ba2d146b4a8a52a575211919547aeecc45328ddda1846bb8242
z6801882e754dfda95c9a1bf0387f4b0e53b4755fe45fd6be9c687e7f060b8961e14d7e181ff241
zb1ca393e1e7a051874971bba46bb20e5906575edd29f188074d7d07eda031304e81305e10cf0b9
z5b967565b599a7486ec65f430e86dc68f23a128915f7be76e74b57183c8ed91d382083d63a9268
zf8d073fb7e9e3b8b3184a258865cfec4d438f7d5b11169da4464ab27204663987e08ca39fc5853
z5821d6215af7f4929da76323a4626e343f0c8e22162e81052e81496cda3f4bfbd78a3c2c9f4ed6
za5b7672f818cdb7c5af471138b702ef6d893677718c3e331af9db6cd0da0f334a8ddad9e6a78a4
zf26c0ead393819b4158071f0b65c21e51f2eea83adfc22dddec690bc31dae00916c5272bf7ec65
ze5dc715feac22528c0b2988d163df1320139de02f15f6b82e73e6e51c3a68c996f38b3618230ab
zf220537d3b6afacda3e2ba15388da427d238cb7133df489a4881217fbaf19957bc2d4c96072e45
z33e7b6ea58c6b0d70cdd873df4a82c16d10e9bde012390c19e3fb8fde4fc275c1f474ba8690c91
z55fb3af086470a57fee94d0b7fd5a45b1c5680ccb7c86def2c81e8ac0a38a2338a4e07a619d283
zcc27d6db5b5c3feec470e73da9ccd5df7057f5b2f3b113b5d51066fd076b35b5d1a7fc6f4c818e
zf34f4900141248eafc035c2c2a2e24094e78f43db6454910e08860ee5872be3bf5a311f5c30f09
z6d0f22ae83f8ef8788ffad864e7ee8a3b9a70a21b8eca7cae29912a271dfbd562882f6e80a57a9
z5a804d420bb2235280bc25a4423f601e573345217495209f1848d20282dce947e1a1c364f80c7e
z1a5f8c614962605796696235f9d4fa08203c4ace05b6bbc46e5adbeeb86658d004fc563401c3a0
zbe9a0f634beb6a94fcc49f7248025ac8bb31342a38b419e12bf68c35160e0527d3b321361c1a69
zf0f2bf5392bcf4d0b27f218c943466fd8b1763257c55e19862ef96c704ea9e89aab30febcb9387
z61cdc66611bed01e0a6b0960a7f727704e976e407ae324b751fd17a6a18aab54e7ecfa43befdc9
zaa63051f4c70021a803b20ccda548a8e21137f912e9e6ec3c89f7a862574e5aad2930f9e190fbc
zb114a28c79a8c3ed79a17a5198b91e2061bdbfac76fffba8e7441a10efe318a664c84a49f63fd6
z47a1c00b755fd2821d55d004b8a113bbb76a148470a1086def97578246652894b0b4333da4ccfc
z41b83ad2ad8132eaad963f1e8320b632e768d8c9cda7ed6f02e16c61ce0cd4efbaab13369aaa71
z311b5f79824a283626cabfb4eab3f2d52122e386483e31f4baba633dd692f7d25095759feabda2
z81f538607b98470f34f26324526ceb39f045775aa01d4a4d7b2e192992a6f87fe1cf23cc40564a
z92337742b714a37c841dfe09bd76de551795603bef2143c9e2f22448765e7a6542ac7bcdcd02ae
z61fb68c053674b5e6aa2aa48528008a040720094dddfe976ae0b944ffcbacbc833282c1266de07
z01f95bdca8a92672f4c4ae649d994ff352325cd7b2e229175ec7900f302261e1e3c2163855cc6e
z544fee6aea79959d744eb188cc1e0841685e4541af88a426546ad7b204dcd138fbe95b084a234d
zbddcb14afb3b2ab5cb60959710aa558c3de51263b5338f18f5ed4a8b464c207d9404f41523caca
z0ff556b0a79eba0e7510f40b4594b4e4f1d051f21e5f058075982d208a85f4dbeb1197b6ea2809
z29a0e90a1ae348fdef3f0b8ef4d6e736177b6c67dd98c84f87ad4b418ec805a1fa93cdf4a786cf
z07819d20bd5e6406766c3e483fdb9290c90a72a6388b28c9d6b8617f4304cdfdbb1e12f0c43187
zea88a41da2173bcf1cd4d68ae2c2e195e394d990499a36282aa253d7ab38bff88bcef36941aec1
z7ed6d952a5b66cd91203856027fabecbf71c1208a58f05040922541d84046a56fa6629a6504c49
zee82828df45e7faeecb97ac990824d0ddc49b0f240c21290ff9dca8176662d97990d782c0ba77c
z011f6c453398bc4c1ae0210f7d263f9e1da497e8472fcea7ff14c015431c4d99f59f11ec1294f6
z98341d4ca5b0992c341d401bc35d192620dec75b3cac6f88a356161115e6832032b1742756f2e5
z0fd997d72642c138096dd8b4114b8acf6c52096314b134a64efaf3e3ef2e7eabd72c3a5dc152cf
z9579ffd2fb7445b38643a54236847d7de6f4a0e404adb47b41615a908aaa34fdfb2b42e320f351
z515352b9c6b0588af028d62946eefc2372d88db8aab6f3227a58890e70812699ee079f1dce7a7e
z345f5742ec1b3db78397134216e6c52a4b28c6fa55bb75291c6bae54b48b2af61864ab07c1d10b
z166143ef01683a3446bbb8da3034d22c90524af64ff2eaa6fb2862f6c2b0b4559499830a79fd25
z26d07f3272edb33139e197369197601e4b451b5db0d341761c1ad009d748ec43b00b293bf7de00
zfb52ceb44dd6b9b55211006320809c2024af0178bbaca8a113ee96ce288b4d9702b13391f589cc
zb01f6ee023bfdc50484fa4920c6ea07884b21b019b34505026bb401b555eb6c7c9e472b476029e
zac8bea71ca3836fcf5d019f1296dc0c827edc992a427d6a5dd7d73b06b088d073cd7cc99eb23b5
z4da86189b0e61ddaa55c87798597d23ed7f41b66c8daf7b2a057e3e827a391acee27b1fdb4cad5
z0391dba56c28100bd803b7d4ad506480d5e8977128dd76b5c4492d0b2efab4130327870bf4470a
z348f40ff63893729d3942015bda8746d318bc7c97403de6e88cba61931af6e1b68feae6980c8ed
zb3381863dd49c4c78af86f5bb97cba146f1f33bc880ff40fd08db63623e6591385371ed44f6639
z68a3fe1bacb9d0d0ee2962e86a0d9e5801f3a2bbd9aa82017b7f1d7048a42f4aeb76620fae2cc6
zb4d8a90d16cf6851f475d062fe5411fc24c20e230f9f2d5f7597ff8bade4f7e2e7adf792a49330
zd66452c3b4a9a43373098bf2161f8017f59484fd2ead25df1a2ab65466c501657b7081b5e333b6
z42481d088f738c9030ed39c8e0fcb182fd1945b11f9c445954bd8d25126869584bcb27d0adef61
z6619876cf0fb43ebf0dff9aa17c6e2b5379334026b1bb4b8084216e68e9b941072b9e270738a61
zff0359549774a30c3c07598189e54e141ace0624b42292391800702ebce2c847389efc5528140d
z35d3235a7cc7768c768e68eedd714558b3305af99506619df5ba5170043f425174ce8117ae54bc
z9718e95b74f520d51bd230085dcf5943d6cd3df5c9266b9e8df3bb78f73a2398386303727e505a
z89789e7ba89e9c38c606e45ad2a4d698c597b8a5d5282a6df63d34b5f82d91be4efea223fb5076
z246492b1f050ea195255443103ee45bb57f1f46f2c8a029c88a4c77f0768e7fa2ab9b102601448
zd375c6933b69b72053fabdcc6ee032f337a22de0ce9fef2afeb73d5872d2ddeba0ff461611d2fe
z6943f4d71c56f095d01811ad5c11f1c70d0121d96d28013fe2cd8ab8100d81e9c3891abe7254ec
zdb7a35d1e01b6798222be8ecd836dcff10f4c9eacf40961b62ab55c4658dd9c37e16f11ec6e3f3
z2982c657194059c3a3da598959e58412849b17be6f7d3ce2abdcd7ab944b879b5e84bf9b507e64
z5c4247bac973e1996abac5d8b2d791eef13e58d59f4a10b879a0c2280db6259d357168ad3b683e
zf19884f45c0e4786006b6afb8572dabcfa163ed2bdac69e6ad9bb4dc9757e7639c1e4ad771a36f
z1d1540a50210a5daff346fd53c519a843968a45f1261d633e15c04f03968d63ec596a468a8cb40
zbbb148724fe6458f762b12a5d7a5b674d545dc093f232db278a4f04d9bdb88bd486243073dfe4e
zc4f18cf655b5a8b3f6f3eb522784e293ca5645bf391755dc788cfdc948283732cf3f14660ee5ba
za83e5ecdf0982fee0ccc9a03a45aaf2e47ac1a12f6e5e265d665dfdb28c48d13d82fb69bb52bd4
z1cb690f1f7645386b1e04e5617918040fa222298cc2ffb4c6448d6a326ca2a36be865bb12bbfb2
z103d3f557422e6a6acce3548a671dae75b6433a6c3a410282eb3526093645aac891ec49906a0bb
z1d43dd2659cc17e804d3a52cc5ce505c79a4c737db2c030ca91ca8e5d2193ac6aa83c572fa5897
z9aa6b5f8a60ea2d62ad01e732c937c5ee612bd967cab8352259532fc59190f19bb42dfb0529710
zd119a93ac04871afc5d78fb52be9439f806c642fa1f1a30f6f35eb1e88e0268f2dfcb4a9c25554
zd631e9652d94daf53f4e1c4add407832597cb8abcec0c757e430a36a77b72de54d4c0f32339b02
z61e1f86b4b9e5463d196eb8854110b5c11b5e8385b994d8554db7a7449c6709c367c88c84e3652
z0b12fc108753d84d2647c4bf4ff4c62daba6936f7672586b01a67823d59d45366a296f88303187
z7e49d61840da286105f1237965532b170baae1dbb8cc30582afc6e1076120cdba03bb8ca55b53e
z2422acb2c7084a58ab48a219224bc21937cd631e5a6f8c2450629378465e75c93f6e77ffcb013b
z4971df7ddb818a417d897ed68b6ab567e7b84d01d357434ad2bc0747307222d511587acd41daa3
z72d271d3d97bd717e69c017317ef91daa6cc26cf03d58bbfadfa1eb32251cfcfef9a8c5a368201
z652a3b246acd91096cc809132e338f6c210ff4f71d86469f74e7b99eb8c7646bb7f2ed3c76fe8b
za5f063492e70d4037c201777e22caa30c77efb520dd0b4b83823bbae32721d08cb459d7c625ca2
zbbeee38ff3b487f8f2f18c737ea94c37efefe1bc76965926bf9712921f35c0a72e69cb3879d9ab
z921b8a613566cd9a7049809c9c5ace97f351c634d0bbe57ac817ef6f84ad3d3fdd9b10cac211df
z3b20cd92e3ad4d8f56087332ba369d849f5e865bfde11bfb7f4558e9e8f82918b1db9cd33c1490
z293a81da4ac5de47477884d85575fb6d10583ecb42758c1c717945725feb0a278ca5aaf8a7f0cc
z65e2edccc51f90191a653768418507c84921e0c1c7822ba37cd32f0f8e9087b5840f6798e0a758
zc5aca772c78d17804a29be8623bd537d47f62268361e38b87efc575ca41749d1af7835e7d48d6a
z48f761684f24858d0df09c96be3b24fd3f2e00f47ca70f03d0630eafaadb2dc5c86beb6cfb604a
z9aa365cf50018c78de59a52ef0f003acd5be89cf8526e7a82e93f233e852fe4813f18ab7b2ea4c
z1c64feeede7f7d338423a1149c7fb304844924cb9f48ae99bb1378dec119c013c5fd551b79298b
z30a136839c0d30814dd5808415853ed133a5748e8f609c6637320d635df67ea9090e86e4abf2d4
zec902420bb20ef4e39da19bc2c0c0776c1cef960d0b51fc19faed8f57cee9a68f0e0d8bf6e0961
zc4cdf45ad2be3077a2476a38dd756699ef698a0e594d33666f909f67f82e17eaef415ff4d14768
za075b10738ae945653c17715479851dbaa77128811de55a2d357a87465a45e99b439535c19d980
zaf02eb9688ee74f9c97940766cbe059edadac00482f10de0256a10c52c0a2be8318a73e2a2cde2
zcb3da63616e59e8af7c2a1c64ad09b7361d106bd063a8698212c86b6c5898d128bae7317f8632d
zc437f061d0c21be0f97b72a70efaa5a15485c1740f8f0399f709c254250a7dbcbee30c71ba7e4d
z73833c22dbe03def2ae80c416b76c2ce0ab6bb531c2d4eb811c6db66a8b2dbc9357ae93aba08b4
z3b8ec1624684e46c75cb1c9fc76d14a339954da95d859f245ece0c8c4eb8b8ac2022fd67fb848d
z2ad5c388b0951d6c9c96e51d5745bdc974a5bda1f6d8066fa70e79c8d6a756a3a48e74b915c954
z2aa01301616cfa208ce1562774d9c84d11046b0b556a7a5480d099fb05a0b312c787953406a37f
z423a2b5a44331ab874d5f018b630523c4d13e469bcce9f49d8f0e5308a9ba4cbee5370da99d401
zeb48110d995ffd61f9ce5403310f7669e774f03ac0fe6fc630d6e61ef634bd8dc98a9dbcf8d649
z48b2cdfd53cfc727df6b07fae24a2e7f99087efed4a6ed62307b8d1be2e5024908fab7ba5686a1
zdfd3c3f0df896a6114707c04795ed87b27df51565310865d22b4f0f456d068624ead40a13e7e8e
zd294971872a1030d370cfd618663b237d7c16ef3092cb69f932005348135900a656f77ce41cef6
zfda8edae84184eb7f63993864cfee33cef4efac5c2f7c2da1c83300ecd6a1d11d43b549927dc38
zbb14e8ca047d5935c79747bff3dd68aa421eac7446f928e9bdf3d9a4d977d860e90c61c79e1003
z6bc1b9770a50e6b76c226e2751ab0ff1a34b17b17769921a5b01aa316dfe4d335bae4ca028088a
z2a09ceb4779ed946a96e988a75ded7a27882e275c5b8daa1eeaa4ab019fcc6ec37fa06e17ec0ea
z5ce4e1a009224dd6915a3a70671d944098e2c2464bfb5a7f824808ce0a6703d40bb09bc9ed53b3
z6111c1e92a6b1d40f08b7ce9d5d60a48ae84575c93f4898e7e1d64fd9ddfb9ccdaadb6a3fc245a
za3c5b2854dfbdc3b3ad0028b19711605801eea1280a104b5c91f79fc9367c14f6e8cb8525693a1
zf4a6001a16406fd28f15a096b557d88dba550e936aebca89236d027f2d17824fb93b203da44218
z01a04ce8aff9fceedabb0faf49182c08c4a24065784d8c81ea6e881c97803593cba18be6d41b92
z3481af4287b9a4d693400e960f75dd0541deb73c069c8cfaa97950bab6ebef5c48225c9843b44c
zb67f5136d65590a7e6f0bb9eb26399a4c9db7997cb77bdfb014bea0bca909e12e7a4f24d719898
z5aaa27b72ad9fc9a6e93245ecc793c2cce42d7024a740a6e1f4891d4e7bcaa96dfa6a1285cc43f
z8f36c17552423418c7e4fa9c9ee604279a4a1c86b5aab5a44c9e8b1883486402ed3fb3e6a8c488
z5342efc2005f52a3bb197fca9f3b5d7cd3930b5026fb8c61d0afa37b39a921c6b3ee1b3a7c787c
zf55faa00b0525780f8ad5f6d496ebd12e70d21ea25defad55b2d3e3ebb673f70b9b10bd1f0dc82
z3fc01bf82f53d1a6bf9800ba484c560ae399059d69ec433f863db4fac933ca917c7383eb189b36
z056c9a791f31e1f390c9b6e115fd896f9d96630269dff909da4967eaf73231f20ea5ed3b6ad99b
zf57acd5e081f99b9bec043fdc1b423a60cc0d3f4d126b464dac832e635a2becb76aff502542e54
zae57fad7c6443480fe7694198edbdc6be3da1e823a873bb755faa8ebbb1a1d8c47594a7fb217ad
ze23d6e4a6f52600c8ad1453991f2b22214cbf20017c048c0aabf0770e03e33c129d18672fbfc92
zcb7e0466b10b5fcbeb58ebb7e29fd054c45aa479848ebeaeff47b77891ccd03d0271217fd71f8d
z9edb8512fa998706402ef37166f117f7fdde0e8b5d1a572a43bff45d631ffd67e97ab4f97adc3f
zc2f5556199abaa0b17f6580acb0efdee432a7b0dd2e6bc680aae5e892fb64805c9d85d8a4453a2
zff96eccde1e139de4167a5dd8280f0788264ba78540d254625469d112d528762f2d81d9362073f
z8e27cd58bc79d3c4b1eabd244488a1fa7fd7715d52fdcb859aa55fe06428d975020ba17b0d2c31
z1938d001bc3018ad0ce72e0669eff1a9c1f0f45582404156ec05bfb9a716119d8ca5149a72412c
z030abd724ffd427bfbb4a322c5e4874f3f8b5fe2ed8a598b96857ab18bf2289c166f537c92c932
z3edebd37418c2a5b21afe525029359d96bfcab5e70123b4f1324c504f53c998a349eefc3619eb0
z7009adf3bc2d670dc0e74105aa30bb63772f785740c816787d0626c08b032315f671cba218a65b
z9ca33166df3d7f4d395f4e9106a109eede34e983fab770ca7e64bbaefdc0d5d4c2ca872f2fe593
z385406fc7ef76cc82d5f7c8abbf0b297247000fc452722abcecc9f342a8848e5ed839d20a5c7eb
zf20943aa9d7c975ac68dfa62bccc8b2c690dd9b3b3b9d051fc8dc893e8ee0207f08a22951b427c
zc73708993fae9d2125e958137efb6529fd8f3dda072d283139d42612d4fd3d2c970f011887fe04
z74bf8d9a3950a08bb3c0e0425bd564220be52b93e01e6ff5107d149c0d4c18354089c6c98e4f28
z8839934ca610aa5a08630c6f8040c5279c13735bd4001447cd532ff3e0f100af48c6b34b82f8a0
z3937f1d37a70b07b816e4da65d021e4be242e485c58e2a3ff816fa896162f0e086539212b32961
z876bf4e51f855a2c6df60c56912f565a632bc043d31cf30c1a785b273d995500c819602daecfb2
ze65a278b425f79221a3b4da8cc7d7ff5eb5058b7fd95cfd47ed4e0c6832480a6fda9b369f5df26
z4aa946dde00f8ed5960466a19c7ae7567f40a143687cd251916a5f45c23524927d4b30be16b8f2
z2fc9faf4288c8d252e93ceea49f30b9a1503029a4d65b28853bff3d3916d6a0858ebf01f8ab36a
z7c605fa46f425f7e8dd90dddf97b2a33d579721cb9136a4059248d4a7a3b4aea49acc11e668a96
zc91cb7bdc47c41ccce4e066e49296ab86d925b9108171ef1d6ae8e6be03fd27cc5376634c199db
z397e021942e10fc8423bf0132239691d55787c4b7af44da8c09f42d619ad37771ab63bd4222624
z31cb595f67633a356aea2f2c8b4452f13526e9e963d51e8489b662a81205568b2354a7edb4ef22
z4df51c840c6985cee9bb2c5720f9be21900f6be3a14dd1c2755760e6c94f92e0e8deb99837c256
zdb3cc52083051d69f5daa253000a0ab934aa42fec5d991ae52fca3c162d2c1ea2a001a5177cb54
z92f140b8a0ef9ae5688297854ad0976d3a676a13e2b085dfc472fd88367e1b3895f50f10fd93f3
z08ad38478a5e125ce759468dbf1ecd5b80c4c47ae0efbc2085cfc0a49fb75af6b98393bc7c5a16
z9057dfea2daa7251e1358b0b3f14668bade6bebeac03201629e16037f65577feb1e4bb888d1d52
z41d503335d43cd661684fbb5e881bd627e8927fb2bd7007cd233921ee74fe9bad24c7490f93538
z1b6afe0b9d02ed0dbe3cc2dccc95036863544b1d6a1a8dc81bf95c115b8b3bcf880087c8b89b76
zbfd8f4e2ded2f27893a70dcea9ef92f6506363655d571fb0df72324425108b712edd406e6f1bf5
z8ad308c1715205ca78e50699f4787eab5939889fc00920149de58ec54d4e22bf1f92d5bbf68f98
z4295b9be37f655fa0934d87f8b0eb9f5904cfcd03278992bd19358557aa19a1880a8c05d54cd06
zec6f0117fb971bd90fed9b12dd5bd774c972cd2d070345f82c2020b4d7d9f254ef9692928f6017
z1f859384fa94dff7f65ebfa073ca46c9f81faef0c4843351914c1c562c4d0f27ea640b663c79e5
zd7128a696c53fd5e8c359f1414575fd9fab47e33504d941a5ffc5db55a7c1132e9f697749fd8fa
zd0a33b6535de63d022a00094a59e734d878d59a0ae2af29a300514b3e666d8a74d6aaaa0863ba0
z0595cc2a7e08776002ec3d2cb83e7beace5890ec38972c3498b0419c3adfd0020483c443b07c01
z0a394d26f772b773b708392fbf4d33df4a35a5223997ea8c4881350e3cceec623475cdd813d6f2
zeb804964b9378aae9333e12e0b755fd234e1f5b3bcd0990e478f7a87e68bd1850c483464266499
zc625f9e724a3a3cf39804523eef79d22cf2360bc88569913cc5dfe63c675a64598ba48465df5e8
zfa017f708dcf45417758463cfdedca90179868331210a1f50e7e8466e4f645f13d627980c6088d
z7d885c182e7fb0f5d97ccb6719e5e40d386541eec554787e31a535e8afcdd581c737fbbbf4c88b
z7d1e89f794ec093dd91103317517cb999ed675191552f4e8a2d52ca679f4299a70592e91d4a27f
z980ca47b451ed3bf4a0992f8a49a7ed02868624b9c93defc4b82fc75f0467fd73c7671cd410d48
z265c1b6d1a3bfa28232e3529fd99431e473f6e2e95b0fbf9bfb695146befbcbb1684997107af6b
z90b4924904e227797841bb81f647149c30bf70fd3f39c2f551cb8c18a6c6e7cf9e7397a1141e11
z431a0eff1a9ae5c6fa2f23cb5a09bc51a79abc2d2fa062dcbc8fa677c5c5812400df69d5dda33b
z1a2f8f69ecbb3e91ed748a72ee09cbd67e6efcb9d1294b01ad4c8124d70a012f2fdd08d86def81
z8321ffb1257badc4d19d57f19a94ec5836fb039d290c789986afd2580ec773e7a8331f1ef2bc7b
z197219f6391cf267989bb1f8a5b65267551e8eaedd859403d36a6c5a1dd74502f7539b7dcdfb87
z88a2d06110fc02a3a5d79d3325be9c773bfc371a6e04ead11437c770122a7dbabe434f2ba6fcdb
zd5b053b7efaf007626cdabaedeb9fcd8a7eda0506acc37e6ac876105f4ed2899bf68b255fdcffb
z010f2a6323353b90889dd22d68ac6fd0cbba71fbeff937b0f369e5f6efcb2e00b546eb03990b27
ze81546dec22d22657d6877f4ba64411da12251299e71583d6924c09af660518f77a290f0d26120
z6edec99c7c8ef00a7c8ce73d7d07e1f820dcfb307453c95ebccd5d615b1daea41adcd4fec4ae57
z42660d43e81b26196dc3c9039a9f099f2d0a25ef628b8a8cd98aa82ed2f81f3165ac4b15ba4f27
z4b165f5bca32945e9735cfd4b4b07afcd387b7823c4035b4d4c67ad34e51a893cfa99a0cdc33ad
z047d2d84b2e92f7fbaee5d743cf3c510a1eb73e4f25c7ccf9f4ad0030ccf2afb07b0814862d9d4
z6dad69c8a5c5181831f08bc591f46c2d186b0e19392e574713be369d35e71eddcd9ad1736f4beb
z1bc37f2e8b0f4157f0a22dd818bc49c8c2c553b29990e83153edbaa88c116548dcc318e89bd5d6
zaad852156785f43bff721b26235c0f692bc5fbc82de8cf7bc92475b7f1c08ef8b43f23655c265b
z4946f9c635782f8d6d9048593b6148d33ff19563e4fab41333983041c23ebddb213cfe09888a8d
zac5669274b305dc8de0dfcd48e60b4d56069910039b430b863c65500e933304477ece1ef57b0d0
zef37825c77437e5b3eeded82056f7323ba85fdcf66fd3585c2a24013a7cc8946beb31473ab4b05
za42509d789d74d78a1686a7b6a1b5fc79039d76678e163fe18531ad714bc3dbaf6d05119d305b6
z4069645377e52922ef8d732d936ea0975106806dfe39a2c90befb833e20d11655f74375609ce30
z021969f1d5c59fc9a47f4aa50dd9a3980171600ceb047e422babd4144132ec5c665259f448fc5f
z83a8f731d7f8f43bb035585a0d3bfc1cc7167eadddae5b4ac0da944dbcf9d3c07f3f6c3cb14203
zdd74bf36f75a1c62e4ca226e8463cce78f3ae5a53f29850eb52d5a479abd2509d5e82d2841770a
zd1290c83783e16b71ad25401ba75e5015fdb979a955c010951c7d6d25d95cfae38001f8d4adfc2
zabe6821ebab2f9ba59289a904ae31139f5d4760c9f2b263b9ae3bed1afe3e0a3d2ba7289e08332
zc7338ffad0cae1bea41f7d2c7daacc8a3a247e33dd1cda1a3a36793fa52ec9d02971e6ee14e198
z983bcd3591de31bdb4db48fd08a65352ff70d92447a6d552659d8c7348dc09ed1f6ddcdea6edd8
z48fa9f0229f655b329a230ef7ae7c1a8217f764b769156bd78ec4dda92b3396dbbe40aca440002
zfbe05cfe522c3c6deaf193a41c9a21bb0da63b0adcd05eadc8c23714c093082e2a4cd956f833a6
z611834b936a482c88bb9fcc2af6f56754803f630cd301e6f7488d2482891bdb4e060737966666c
z75eed6c124a053a4f99fb993863ce642fb613b5c3ce4f84e3efa04ea3c15e76ded1b888594a927
z7daaabf6c580c4be2077fc59121ed1f39640ec30ad20564f094a701651c6e8eba7d8be1d486cfa
z4e9561b74f2cbf4861610bf947a45c13774ef073d50fa4cd41cd4465834529b6139fff28a6b576
zaad296e391c3ce2191ab7358f5b28e18469ee8492a8783c077982de8a01e3f70f5f01e67d248fb
z0aa5715515447c0bd9cfbd51dcd308d69b7bd0b704d1fb181d4aae685cdb5fe85806d438c8deae
z29ab6e8792cfedb2d860c87a921cf94fa58111e5db542e66f41836652862bb039e8a238611fca6
z92b019b5c1afd5ac9506e8c692da53f2202166c555e86d8f2bbe1f2bdb5353d2d242a9e7f228bd
ze1cdefadb1c6e566f7822de7a9cc831573eeac30e2dd543b8edf1ceb2138bad7360aa30ee2e704
z8c1a3ace39afdb9b671705943f4deb6480698b8023de2046601b281ff8fd0b45ccb3566fd12b84
za80810b1065d02e3cefa4e2e9878a30da3bb57d77b71e2afdad49bc5b1dad01cd09a4d69ec5069
z7eb96abd5a098d3c9468921d1617f2d1ff5c54caff4f728561e1cb64475bf90ec438a72e7f3e9d
z81389ff81d111ffcc5078ebd0ff47d930313c0501427e233c66165e4d6907a5def9d44901f5f17
z7bac2a7aa838d4606ed310939217a3d58c800897454403e292270210309d0499ce295923532ba2
zdafa99274b108e0e2b3f9c5fe868c97e59bbde44d9f44c830f10e37f0318c23c4be05c51d4fce3
zeb4316548c7ec9cbdaf6cf372d91553c869b010e44d231a09ffbb56d9a99c5ac92500f9f0189f7
zca4a165e3202092090b872c45b1336a6fa23263795ead7b7185f8bbd0366ccd8ef72674c83108c
zd8a44ec1be9292eee3444c8bced94c1718173ce7103e22153a74056cd8f1e9a20ac1ef8fb88d3a
za70d9826fc5ef7cef8c3e59c35770c3e3f8fd8cd7d76a482aabaf4ba9142d553539739e7d0b4b2
zed9589d9c2cd91286e2bd0bd5cf8c08092c341a5fc34e688afb2cd30f74d9b543d9d34c1adda7a
z7735dad6f7b6b84e04ae01a0acb4aa40f1f3280423f6b489fbb4ca8892741409958853a7b1290a
zff8b8ae81a348f166f9eeaee56dae92d3ca2b51adfe1bbfc727a60da509db96bf0b8d5319612e3
z9757a9df2548cd2efe0e59f5a92ea3dc6b9d08abc340e857c2fb22580857fabd52d84cc76a2046
z0349e4df974dafa558738f6e21badc3f782239575536545fa2c863658c2e248788b26ade4bdcaa
z7e83e21655bfbc7ec4145e23974435a0d2215987ef6ccdcfb448d433c36b1766c23aceb1fae3b1
z05f6e2c6db941c48bf5eafee3a530c6da9a8f44df8614962801e98984ee9eb48d41050c5adbaa9
z13105bcf22a9046be238190985ac1282f7c4d46577b1120be1d4f2c9385239e1e772fe09ffc9e9
z9e9dafe210176cc4f825d6fa2928e00af1ce7835e76ba964682bbd73c19a3ead84874abc09199b
zf5fdc1e6f7ed70fe9022782a4fa653d9fb67781d3f33159410b0f420b91643418e228288e61809
z450f632c4373bcac6007a93e4a60663a1917a1f54ba478dc540855e02c0ccf24a83dcdd5b7b28f
z91667622cd85590108f9a4cdcbdd1a1265d11600bb98d729b46136f3c900fba3474c189dc06fcc
z3a5818966ace4c433c2ff43256c0ba91e4cd18066cfd4fd35b91bc3536bc73030bf2b331af98ce
za3cc3e6846183c5875feac0da789bc310c1f0439243d1132a58f6c119e52df59775ee111a65f1c
z6c51f031ad23a05b3fc356c13023b4e119c9cb496a9e295840a675f4456881a4d825c9e31365dd
z6dea0853fec9d3f6e43f4679994dd9e5c82f6ff9e905e83016e52bdca5fee0ad43373e84c6b16e
zdcf5ef9ba455baa1a370a2a6cbd7c2903588144a45be254f97194ae01de1d5cd1e5197f1d36391
za82ec804f2b434f6f9e79c5db85c2d372598f911e385798ae3848a25ea600e48798ed3a8c45753
z77f2c355d0312b7e09d979345f4848ce5316828b88e709214132c29bca5fe22d4a10ce475dcc27
zbeb22f6cbc9211b70b57f1b76ff4f83b87e0f365f552a88ecd9da4e3daa11e5a95fd48f7428af0
zf94f2492c7fd767e6c9a8697b8b0e1a5cd429bf4ca3e6bb0c783306667561c2b4ca3d785ab0440
z859f4564e2440bf4cf5e2618b51e19a44813d2b2ed0014207395470d82952513b710b22220e40d
za5231c57410c0ce0de17c4d228ab522430c0cba9f75b3ea537f9a5cb4b1afe0f7c8860fe532143
z507c006f7774babe9e98ca500c5345c760e8852f11c210aba06f177989ab620f861d617e18c10c
zaa97e60bd5bc5dd972fca7fbf0a1380449809aacaaf7bc957ad102ab990c18e181ff35d07ffdf2
z1bc375c3e4b3d80bac0124c72e07451b79fa4814edb9a4b44a14edd0f1c7de91c84dc838fa67aa
zda3698d1f4c2451208e2d4670d6c81923add30ee219275120909fd8d5aa5c64ededff9816ada35
zb6891b0a7909e772d105a8e27e6835b1b16fde15a04c2922cd13aaf2e9691ed18bf111c8df0402
z0e759741e6dd39d7ea58f6dba8f7d20a5b97b54d78180f2d398ef718dded809d34a5c0a5075f81
z1e2d607182fe6dbbaa061d1a3ff97fe3d5037462148db99717f8103f017d0dbba57f7e2bc5e060
zd15d80ae2a78bbb375efc939839c4a7c6a3e229f253d60b3ad216672fb8f43e61547a004487d9a
z50e3fe535c9e5735bc70ae84333cf51821cf2a4c07c8115dac8712dd456a8105ca413088be7802
z3a5a244911a7e0356b4a8eaa10e5b2a9ef836ca68fe5c17e335ff233a1ef189bcc64f3eb82d3c6
ze4add172d93cfa55fcd9cc0cc16e72aa5989ea5819645e6e198abc93b71d18e456094874331b85
za75aab5a73667b2f3b2c61e3c7f57f73c388ad3478c54be68580517d0e644f61e428ec37543d17
z1fc0c304073bca7ca5f242ba183fdf8ee4c5ba5a28906eaeb8328756fc00f8f6533af86d22ef41
z9d63afb8e77c6ac3a8a27f3dac72cd4de73d84a3b5094833e0dbbe620195939c789f1704bd20a0
ze2a12109613736f13a2d093d7af584aca223b7467471826f19d1d6ea103e8b12ddfa60e99abc67
zabd0c4d86ad985d949ea19b4540369aab68cd17e5df2d85bfb1a6c8e4a6430e2330e557f8fc0e5
zf75c4163fd36699472896b988c554313fb41fb9644af5a448543ce743a4ceff409acefe624be03
z4a9c6172e7056b08164830121f46be2e5aa1ef285d7d418e2a4fa5e35440d757ca33776edaa980
zd1c559e6ddedd449c7c5229f350e60eb08f438807d13ae9eacf9e11c292c6f34f49a9b47c00e21
z5a865ae5f90633e2b8a1b78a685a329260a37ea30c5f21a9cd536daf2376608f4b83afb22a7baf
zfc1b616dd33c59e71a8a95187fdb249acc190b5c82373dbe6af4d0bb794df6c990a0dbe54e7b85
z0ba90374765f4b74f7693c4935d3ef9a46d1d0df253d49cd7fafe20a93cf2fded2b548a0a55315
z295f421fe0752b1c5f1a92d18723916844424e33077cd8315146c624f5c8e7ef9f5587c7963d66
z5c95bcb6564e688fe53d999a69506f28a3f0efbed73eca4705c85a089b205d650121f0e7e218f1
zcb88e2cf2a8b52f687571a78c6d634e9810ea6c87c2c5f5d4dedec810e9b30aff9ac2139678d53
z882baebd802698573ccaaccee8f243d676c2980eaec39256b83ac547f1162a5d1e426006badc31
z77325b7c72afc58cbf9bba9a5b2270323043d6f44637fc2349e43814967098e56bba5897cfd68a
zce493e5c4472fd718cc7932673ada0d508e186375075e80913a3173523ec9f0ea56cfb40a6fa3e
ze212c3cf768965bf98772287d0d51e4dc5f8925383eeb776459b36b9c0be8e1e4b244c59d4ad4c
z8a0bf2958976c6f3940b71bc8d3747e56d75f960098cfc56633a248dea8822bae5b7539a8afb95
z28ec6f661a380beab87f42536ed9eb212608bb5735e302ed8cd55f51456bb0f875e048036f6f10
z4837a2a48136c84fd1be41f79cd0d2d7a2c05e9af134c03000ef8de548f868a0197ca4618e1b77
zd3d76ceb5c2cc2feefa88959f6297575125998c0c229a368e47e1568364eb00eac2e7b6b677b0c
z203434f73604b6e436eb21c09f94e8bd6a72ae165f643d41db9fe99cc42dacc24bade2b6ca1698
zf930fd2684ed988380747c620ae9e3c58fc670df107069048c8f3a43c18745925ac3d84ee79ee1
ze2a62ff2ccd94fc5cabe440c28447274ba66e343ddba0478a418fa76232922c31f01c31d4217d6
z31b5b94124495a28d631bc805e13b46e9c2492339c1307d54bdc69fd8a177658b569f515902bcf
z28254840ee1a5aae13332985a63db7cdbaee4014585a15718ea9cddb3264a8e9ccd6a5bb606495
z0d260596c8633514f40223684c089e4698017185dce58f479f9c3aac897e24ebf3db0ef5aa6976
z91834fd9681fad402b377097cdca52ae7123d62caec42b76e8d7e876a550c4fa11cfe6bb1bf673
ze4e23911d16599a7103dd3072bc61a458b88dcf65c63712e694a409899374dd857063f1fed6dd6
z2b8958adfdcd942e1a462bd8dbf47d83748b86b49bdcdc7ed920079876bc62b6f38f241b76915c
zd30f0b58b61ba296f7443fe4941bdab3aa5ae16aaca86f21aa57f4ea5ed72c33332f2ee49a3a0a
z99e54561599636d67134730e9f15a8413e054da2014580d4a3d47516ef18f157a27e7793409cea
z99d14d3f5d9206414e1246dcfce8cbaf14948863709a6967f29c0b23bfa0ec812dec24efcf6067
z600205697c9f6b4d0a00177293654bd571036df29af204510a345e7f23a5ffb491ba805f574c13
zab7a1f4a04a3d5747f490e0da0308244d7afe7cfd573583459ac511472dd508717c61ec4502363
z12a5a8db07e952f8defc41775afd31c125af6f905f457468cfc8c66a5fa1e62f87dc334b7fb3d4
zd112b9e6c6a5319ccf512d4587ac365ab4b7d7a4b32d6178a48c888b057b9c5d17898ab198b707
z3da954dd2de42ce84cd65c7cf71da2a580d297141ef31e9829ac54ced3a93fcd18915819c2492b
z354fc6df601514713b390af38c304f263b549c9a548804f160a0bfc36ab0a397efaa56267a22f0
ze721fe857ff1fe083e111a3000307d4f5a563c8c6cd6ffcaf3c9e9e062d7d37481a4445fc02042
z11e39462dbce262bc88638c3af66e29c2519ad688fa7a385a030b49be12b64adf149b6fa77752b
z672b5ce10d6d756b89789b892e3306bf1367f7d925ab440157d83488dc616832c248fc76f60c2e
zd3347034665083e5557d36eb52e4c204b361e7c199bfcae0b957c0ffa8827b36e03cd95501b5af
z686207d9cfd6304583f5598a8c2e300be0cf99d915fc0df8686d4a9bb31ea36191ec1f3a9c3e8c
z89235239853800032790d87f81d6961b395994de1d3fbc96d9659ce52452b20bcb29d7d7f1a54a
zc4127c8e865c48f3c9129105f2bbcb0a90c518cdcc0d7b3eef0cd70b55a01ab9a7adbb446e24c2
z154bcf8f2cb40587886520145b5f264f0673e1ce200b1427fb5ac755471f64562076ab2e62451d
z83b2211e00a8a8015e7c5ec177e875c34f3c9adb7216e7b93a0b2e17b89c09f6ae0cdcf7988d4e
z0827c622346db9a08e86fea75ae416d8ab8b31a9e12de56b225ea2ee047be7b022ae3fc569509d
z3635ebd0b6399403f0158d6f52cea586e2685892b075d6e4289348c5be5050e916f31ca1514c17
z8ca18472612c227fca0a4fe517276c39624263b7ffccfd7586a2f0c3788bd2e57611d6013c6d77
zafe81d183c958e95d84b746a6b3037c36b1512829db26387370a580d919c5c66491e361ed8588f
zf02aab81c2753b734508fae98a671a1839232c8887f898124b981c25f37ba2accda0430a30ab6c
za49c0d7301831ba3825b437e69c96fdca2e0c25e8816819aa3532cbb167ce413a2047386e9f4a2
z55f4c9396c47b2c257785f7bcf4bbf383e9e3ebe00968848fe44d433dfcd3a83dd571ae335513e
zd44f7e6ce9babda1c47f8edc49f7caff56c13a2cb1093409fb7a1866fd50b1d549cacee664b4a2
z25af1ff65ed536ca4c436c1d539afb9013e39fffa1462ae8660b54d07c9ceac441c62dc8600622
z4cebf29e415573622fe16d1ecefc0f264b53f9e00acf9d1ad927579383c1e7f47e38896dabeb0e
z2af8ae41b9dd30726be9f5a45412f690a32e401afbbcf52887de95537ee96bd3d99547a689305d
z12b3f78c5787bf4a51bfc86075dc0955f1a6e3fa0288457902a23240aa618e9d647ea3cbc07995
zbdcc6e679f9d8f2442b78d2c84face38820b19d27f204f394cc29e6ca27cedeedac04d2eeab556
z933c800f29bd46e47c5267cb147d37b41ee29bcacc55d7ec708a1fe0c14c7481fe243af11fae53
za32a556afc2a46c7defe3ceff53db19fe632ccb13b685d689805a20efac28a871a4056f545fea0
z1559f18399a79089e0968829872d776112b5288674257a8ca1e286e79a959425126a1f9d77c080
ze0d99a4ced18f42493ec69300447692513e9f89ba48f09d0bf38eff39933835a7db6341408cf06
z1c5a549e89727fc590e30fae19f4debb57ede660bdf48bde02d62c4b04da0d1c00d145019bb6a6
zf9603288a0afb3d0b8956c5965fc41b268fdb412b7f5d78129a4537a53f0cff80c437f46ed3df9
zc9c0f313444dc08cbc9ed696191d81f9b23162b90383eb509ef338aa95b0a713b605d7771859ae
z68945896af9c3ddff52aa456d886d81c8cc640a1fb07a6c5ef7f143a11d598add23ccc57154178
z076d2d6a96aec1de359e09bb5cfe89d2611b4c86dbecc3b6d7a3afa10d7162d094db70bac3656c
zcdde8ac6182e28dfc1b92d02b36f460e17e5bad336167b9d0b5974122a3d0b5303fc83db5623a2
zb0a93784861eaa92df3aeb3944d93dc796b4f49469fd735bc2cd0aebf3fbd7fe69ed656cbfe5c9
zd6827664c6c54f2053f8b623d73e9d45b30d954d5dee8dfe90b32047534c311b4c695ac7124eaa
z4aca79e925be1c54225d17632899b7dc8785d2e2aa7183fcb991989649851d4b9447518d694b72
za985654bce3f09a59d5ba1a538b27966f8cb6ae2e7d005a42558d7ba0910ae4b89f0205887c0de
zd60f52eee05e20e19692d61a9362475f45478e8df48b2d651305a9419e481393e1858031f0e4fa
z4c6314a84963f11c88c4f5d8a2496ad71463c1f7bcf1b3d7d5cce5d0006b9af79af00e17b3885e
z50a4843920fca215ff93dec61c36068d5a73b51aec972f6c72a40c7e381b141b8ad6cde352de1c
z958b283e91237402e4c7c49909f05bf1c01d00405d8332132e644efc83177464abb68f8b195da1
ze5b7e8786b31b8a741630ae328d211e449a606dc754b7513231515a80cdcb1f9a0f330c62fd64e
z64023cf510c80599ccdbef5269c9bc9dcec9fbfbea9e43913cafd5f32808dbda0647e9855cfbd9
zfdd61feda97dab8e1a54901fed307ba7d56565c778897604e8551d253a697f99135c38c7925c07
z5f78c9f1ee4637706a8c1cba356630b45e0349927226caaa291444dd40919851f35bd71bfd29e4
zbde56d10d238871ce23197ef01616b6632e392cba9f69a62fe2950468e4febe172cbb1671fd096
z25b712b7c895a360b2299219d204c12bb4ac8241204914def575dba519b0e0be2fd4a695f102f8
z5feac41ccf36157ab8957c162fcc601bc7d0c90334e83468a66b8a74163240ebe8e55044a36bdb
z6055468035d976469a87c5bf02008bdd68052cd0b54cffbcf9b1f7bd4727cf91b990affd125509
za037c9dee9aeadac7a08b359927a2a549c1d4a793143ab7d99300256e02b621303f03e4033fb79
zf155d055c00cdd5fc29d88391021f55e4ed1ebc99056b4fafc3fd1b92ce1349a3034f751131981
z669e082f93767872ab65b3173acbebf8e9954c91535cc3765a268b55415db7744d0d057aa0ad38
zad64b5c3332455de44ef67a7db47a65d97c1ddfc602c6647ce1a41bace782dc61d393f6112ba92
z925d17cf16c093567c97e41f0c31b1fd4a3577051ea7cf8d197e035dd0d94f27a9323da244e9b2
z6d006d1e0df9a6458ba756e6fcadf9f430255ad0a13713be0aece7b4adde65d8775bb3c30175b0
z35af4ea5a7bd6a6cde850aff427edac4c30ad2a0e972593505f94a9af648bf9382d60bbe160a31
z865f6cfca18a875cbb85b2ec0f69bce61142e9559ea950065fa45b37463d3df12131199f73ea4e
z687cc946f1f9b8c1425733218153ed330615d82261fd7bd7ca2e02cd9c28361a311065b3207beb
zf70ab6c1f3fc1290629393dc6278187cac00a31660c43ba08aeee7bdbba0b6b19e14c6dfbfae85
z568a71cb9a9efba4072a77c52124de223287391ea9a224ce6645ef5603f487c7b4d75c619c1e90
zd56d70f87b95bbfa4d2429edaf1864e4910853ee8b0291a297ae688a20c822ccdb782f67af37c3
zd221efb7b4570508fdf314d4b12114f458a030215c2f11f216442a42b1c165abed2b5fc004702b
z6248cf086011d9e95784c9dded4e2c8eafed967b457a383116990c445467d4c035378bd4547298
z088d7078b185300e95b2be31d4adf9be8869f0e228c92fbc9ed0af721c2ee5871b48d6b7b1d0fb
z950d5bdeb9a0a6b7c5ebc0694a7aeee1f3caff74260e21d6d32803f8d94c692c5e2584c67f1615
z74731018241dff60b359ab7dd6a3d59ba1e19690aa8edd82fa1e8686ed165c232d259db80100ad
z9d333e2b5aa4bf070d0d96ac0d16f5204096841645b3d356a628faab7678660ec88353cc30137f
zecace0dce6ca0c8050532860d4063fb3d643d37b74300c54ab959f5984209274cbb82d9d6b2c4a
z8d7253f018134575d80630f35b747129daaefe6604529b3b409abf8419a5c763da6a8cb5f8f5c6
z063777ddfd757451e5e9e1fe9c12b5a032a4af9aa5ce2de00c504ba8f3313a7a89941bcc98d906
z0f471c0c083019690099504fb5c6ded72253725f1e7199fb2e1ed8f5a801ca20798c160a0fcbec
z311a8dff40c8c51e77a6aa9090c80d0ccdebe6c296cc99d5d71d5e2ec0c17622d631383bc8a17d
z213c8b380e8abe94c94dc845f15ab70cacc8bea82b841f6b98af0919ff3cd9ffaf2b796b9f956f
ze0f1194a603aff26260d8b19b44adcacb981373a5ea8d08e98a2975f1a33116d06d412dac9873d
ze6ef7c402142bc203187e235459fe26dffe20a9f689ef7d7d50491935130290c9b53be44dacfed
z54ebe3f914f809a4b79d6067220f7f49856362702d3e7102bf73ecc05ce854e6b77f9e5e69004d
z2f80370be274b7617ca62a025425be34480a50bd288b9685c54c5c352a8a388ee17ec47ace05f7
z2af6ce70c3d7aa51fdbb3efc3ae9f821b6826a6cbff37efbc7e7c3a52f58ed57fd96c6af507875
zce6605a53180d7fc22162f3bd4357873990bbd9331ad8bfe5e2d962c91fc737e29508ebf631ee6
z19c8bec939ab4b366f6374f10d6a0c2e6fb3cc19f20100f515f6c67a8b003e51f15b236181a1c2
zee23c6435c3a371ba9f756857a15c2d603a8923ffa1d9e9908625430fc80c6d69feb211ee85080
zf8df52f22c6870dcb4e3ae9059a625f8b06215e99dab9cced6c192a479a151781c9fc07fa77d3b
z2551ed5ff776a7bd74dc27b5755b3b97122743a5cbe1c4e76760a2de79c289172aa1be84484939
z1127dd2f42330ed2721e8a0c161c4b5649b1fc8489b2cd5263c45c22e1388c0b9402c8ee4a30e5
z7b79f4a01544123e63658f7a0b00d642424355365aaef83db9fbae88d829ef2155adf4896e559d
z10b33ded3a1d14f5fe7c7c6df446dc984765141c0175f82298653067319d9890b75415c89eff94
zdd4fad9c8b05b5073e1cd6d03e5c2865cc78f98693f1c3141d1fa0ede95c0d4e012536aa8e6254
z359ba3a20feb6854a4bb2572aecf7d68f2b63b886e5b8354727310c8e0d7dc8421f1c0bd351417
z681f66e3e455887ea024e20a9b595ce4acbd5e5e83da45cf43d4a99669e51b0be517bff1dbf01d
z53acad37144aa49ea24e4adf0a920d8e4c2f9fbc82c8fc81f9eed6d4bf1517e3df59d7009be3a7
z0c3b40bb5279324a2a811f964118455d2046cfd4e76cb7625a62464a35bd5b6ba3dd91595fa776
zc3447244290ddf3f1fb45d2596b5f02edee9683aa4d00df574010e83dcef155e0a04272d283ef2
z85a61f7b82e349ad0023c8390695e10642bae84cc8e7f8d6596049c403bf9b647d3da6948e203c
z6498f3c9ccff326ea74dc45c082cd44c5f0fe1e9de11d260bc759f5063be28a3eee6832db3c22d
z8c9acb9f3d2ecdb5f29465259fb97207d4ed978d2d5c3040625320c13423222709b620c677d350
z5cbdb43aa850111ee0d5cbc81d35ce4b9a5fbc16a00eebd66a374b30fef1f8f34f85ed22f45f67
zb3ddbafe0fee5d7b20c746d3fe94af6d1d8e1dd60ddbd305c53d6c9b2a09924d3fef3c45bd0cc3
z32feae62771169c17e1c8f1e5d5d92b5009dd8ef3563b736ff672f243c888f7cc63f36195b9a9c
z21a9e51ba961f28e8671f451a5859d221db9044295ac74b82c08bc8672c773f07b8bebb7911ec9
z4b93e4232bf52a254d0db6e1011d2702e7aaced887336464297cc6d7c5ac539844309316506184
z983faf7ad3d72c42086be8226683927a2ac81cd9b277ba53286cdcafc32919568181dd7523f1a2
zf6e15b5a6e1a82477ca792382fc535be5dad5292788badd308a756c220388d838241ec848e2a31
z2fdcfe1421c0bae28643c9e521c08c48179d33b992bbddb00788709099c83e73c8f18586bf9bf0
ze10694662b9ee9bbd113e6b7a33c3adef82403a956da2c9a1c6ab1ce81bb79b668091a857b9b85
za0c46fb611b1d3abc94f0e4d47b097a4d1d3328f1400df534215646f8e5063ee2056690be62fdf
zb746dc9a26d6f8bf43c7d3770d5207fcc8ae9db4e13204d027db8400b4ceb2fcffb7fadb1a89a9
z31a45a50024e2a0ffaa51657557bbf38c7a07c5580e526982f819ebc33a109f9def5b1b62a257c
z2efc09c1049f4033203f84909676fd7f89493d832af966af0e344da855b97852f6b9303996c402
zc79d51ebd0d151deb30bdf5fef977f9ef20edd39383dac1b514fc934758ff4f8568523a5d858dc
z0bd773a1e45af4eff05789178542cc55b4fc7322681be9a1765da60503d7255ddf34396e2674d5
zd8cb7023f5567c99fc5c10776a3063ee3ebbff46cfeb6841e6c9fab22a98e5bee11213d94cfbf6
zb3bd25b1858eae71bc0487a5d0a3bd3516dc85c5110d7a0cd73b29a62dabb203e364520ddeabc1
z6603419808cb2f322bc0f47827a78a545c680233f181212a2db418239687fd765637d89295ab45
z6e5aad40a37ede7aa5f612d017dbf0c95e966f57c7056e0ec83815dfc104f842775c4f81ccc33f
zbf8ec5d08505a189ce9a6d86e125636fa944c9d70c2335d33cb8f91844947d89d53d4aaf70c3fb
z0d7e13fc732a8434f97739285ae55509fd81e8b5613dd5c4cdf258e1c66554e347515889893ced
z6acda08b0b7a2ba30a0de01f0e968702169b6a644610cdb9b5a26836dfafe5ea62dbcf2d28efaa
z3d21d79d02c3555a4877707e155211f880629e1deaa38552d0f4d50e28dcbeb816ff9605ba980d
z92e210dd54b6867275aaa2f5af85d63884945038e252689422df34aaa3b108fe6760cecaa55204
z482a04db4181e985725b768cff26b481357982d29b8fd66cf604f1c61e0d8461be7392b77e491a
z09f064b3fa6c3ed2bd8d7ce92d457ee7b1d73ed7c4e0c4a5099c072a29e608ba8b9124852136c4
z46d4cb2ab7584a14ce633c4cdf62862139ce4b385e0b89d8c0c7294cf1fd029ee2d73c9612462e
zb71f42741402d1aa62f12c6d1d6703498e5fa29497661ace29e73d8d50140b3a2f36dcf4515c00
z732bdd7587dca075993f906fd7fde7ec3b0f373aa1c729658abdddfc79a1cf29da0b1896c6bf6e
zb9f1f6b1adaaf139580de0079b261d1b52a639ec8a75df30efc578da57556f3508fdc35d2a03a8
z6fce7807a07728701b1e1cd4fd92ce34ae1b950a55432f56c731d8e9c93dae1fb155780cfb8fea
z6043621711c7f71f066f31c1e37996d9966173fe03227eb5dcd8173dfac61b6a1e3674bc6e06d8
z3f7c4e8fb8a6a5f36f61377e4674c09b1f475f5ea95783d35cd8ae8f935c520e300f9264dbac1b
z601e9c8baeee24f352ee4405924936b113a91484e4706680f80cb8eee53390c5b9250b38b654a6
z1915c73d5b7acdfbce1c21db5521ca5982b248bc98ea157478cf00038a3bddd0b49728ff5cc168
z82edf5ddfc9e60e385c6920c0b7999dabad11e0d53ba8de49fb8016e776b9a0186cedbd5bee397
z6892c86048df484d4704be86b3890296e945cab5902efb2dc302e94fe8d12a8b8f8754a413eb6f
zb5a0e388fbd0bb085de97b1efae6ccedc506ddea03bb31db697cbae61b01d6e1d34a9cfaf790de
z5a232aa18dc0984a791dd7560141318a9d4bdf7d73b03156f7ba91e4a6226f2dbc2710b5190bcb
zcc4f4973db5418d8dd022c0a72975482492a003c54f19576f6eab8ecd7ee14a15676890af7dbc4
zae3fae7da902a53ec5eb41d03f714f1d04a79ed0404020774f67e239f6eea2988d1689a6484c3f
z015338b2724bb15e05d286f63bee73d3afa1de1dac202f2136bd9a6288307a21507d3b34c6ca2c
ze8b8a249a46cc778e8b82b67b5d3de07ae7b43f4d0798fc74f486dc941f8e465ec773f7a007a13
zd569992a7624e2889574f88c5d9290a31d826826036ab66150338b5aa61233ccd9491874fa206d
z5c347f53f171451ef52ed4a9f767b73e58921c9b96eb8b5454e497e06187ce7f954c35a683a47d
zee6679208e9d7e8814aff3eb2d60ba756bdd02e1bb60b6c8aae9c1accab1ff29da234b019e0848
zd480d3900023176d8185ae1dd9428f40bd2413fc379fc98be575e8e90cd06b4f27dc8e35f49b75
z2a00649d547e907b0a17e2e298f693c4e54e669e88233941c35ede697e2c6d1af3ef17767a2de0
zc74af4a8f9a7d0582d965eabb04cd07776d01e3804d119be2c6948a782cd63379e2ed65710fdea
ze40311f0b3c5933267395c5acf8d17f4d8ee039b216493835530954617922682ac12ba57eb169c
z49a1582c145eab9f3df11cca044193b38d489bd267a2b43cdc85825a664031ab6f81d69db3133a
ze70e703ea6dbd73ba39acf88359fb3d9a8628334b40bbc3c5daab88bcb0bf5cb5fbe4402e13f32
z5c3e6edd9c1ee3100e52806c11573e3c19311910542ffa4b5563cc1b369c56148c335be85c7edd
z6694893eaa2f340a4e0e7b67fe24cf00e4df6c19fcd3a21f5d8286dbdae67f1dd83deebbcb20a2
z71037b706c94f9ad7779f4e93e5b9b14b5594ca062861b627335eb6950b9e58216fe152868649f
zffd07c206ec23734e95e32840f13a6abcb7b1ec1f6d0be471ba6a9cbe8e262aa17167d851dbc42
z9d326aa5614fa51e589074e1541fa1fd0bded9af35e824da14fbed5c002008034d180682384782
z483f14422b6439e5982ca31f1b2f31286ae7e972afa47906dfbf59a86316c3a79025a4284845ab
z740bd46f2cff5edce13794c36150d810d3f0b9ca85f5a94229828bca7afc89f2a73fabe1134ed2
zf982ff1c9595fe8202915d75ecb1d9826d7e0779f5ec50217073f7082588bc53c9ae00b847d0b2
zd16b7c8c55a6cee54437db59d7cd01803432c3115ca28e1e49a7cfa682fc3401b7b72f3766af64
ze2333e8499f9f0a74da3e81606cd4cd764049cad2c83e4c5d4e403433512c73434818a672c8c27
z7c4b631bb3baf8b8023d24ba2e67ba672444d2e2cbec20ec254cc780c1f947ec4843aa611bd144
z6ff126c01b6734c828f141a6a8e18f627836856e2a333012d221ab4538f2be02470769a907b778
ze32dc9babe91e9f37a6711e670d203fde569f5af99e160f1b1a233c6713e12e99b48e89fe2d113
zb4506e674d5075a636509115ef7132863b7bc0582ee88354675a370156439fdb9d0d75f750b7cd
zc166fc903678ffad0dbfd4c21781b215936868a8ca1fd2c82e004bf2cb48b8e6aeae9cad47b858
zc467e8a9e1d50aee1e8ced1604acc1c8cbd50ab7e13b7bef7283d5f147baedcfe91643ead45b03
za6131c3ccd679d17ea92c8a4f688e8a97ba9c3f5ac0001779a30f4a6fa566f185f4d221e17315f
zd4578545dd9189ee7262601bed0a8c7798ecc598b9213644d16ee73c6b2d3db0b35975f9e49634
z384b851dccf1bb678feb7a93b7d3e8d3ff16f8201ce4ea07515734b62cade434577a26dbc52ba1
z2f2756bb62c7f0f77726f0d9cfc0414a2cf8de511bdd335e9b4ae560cff1cf43d6ced1b7b4a59a
z5caad0999be97713af663d2be1934d2851cabcfa16218080476e4906f46775a023fa04f5ded44e
z0b9630dd7dc45c3994cdf8b59a0bd02c4da52f346ec6f7049f9afffdfab546281f72573607ec4b
z5356bed6349e48aad92c8f677c45a853dcf495da8f691214679ea3ab40e6404fa1a8212a5acf92
zc22ab694dac203061479844450e7413aef5137354f806a9a0247d0bb310a5849ecb88e85017905
z76bda0ded89497f074f041fa218d2d0697c045a817d8b862638ea73833a706a80cfa2e3b99a718
zba38f3bea895823066eb13f93d6dfaacde0b600787e985734f25c420f644c17bf8978ab1c80c30
z580310a3837137853e733c52001548d59f9221cf18d496b4e8aba995262be2187fe0c41e347911
zc94fc846e750dec1813a4c66dc129a6dbc271737fae5ef43403a927112e0996c93c4e4afc02f22
za1ef07aee561ae0e118f7dfd372121678d0279fc3faf00f4df8a6da713ae089c5b6986038f9332
zb776e2190ffb7e85a765cd1d04e2bad9f857e72a8ac4f7d0acd51bf6622b50be1fe9e3e0e2d2b5
zc0c783fc3769810e08e1488792ed1c4ad370ba8ff85fb6f34bdb0a2b7ad32a699adcff57cb7984
zc2d24dd4b99d2574eae0950f2bf3b3179e8d66e532245bcbd4e611497f8e1f5a223d1ad2c93267
z167af3f9b3df2521c294ca9b9eb28739f81cb5e60c3a224975c0bdc405b75989b865a89b0fb35d
z38b7b9f84679e0bd9f8b5c2cb396597d1b8b2267b9d957e5a782a3b230cb93b8849ea8a9a711d4
z90d4c9c1e7defb5852f07af57113ef44de3f40f9bf900aeab9cb471c4cc26cc5e149b4f920c9d7
z4242e3a3bb0b56b91de0efec1d55fcc945a65904f0cf38efd2fc1ca676bf9ad5d220cbd89f09db
zb97765efd46bffd798e550ef970c59b898b402e5d8c472d39368d6f2005c1b044c20bfddba9ae9
z995d4c90d3b37c927a8dccd0c599c99b1410072ea9a19fa953d4d5dd47d8d1713fc73b346cb462
z203d153ccfd3c8d22dbc0c2344d6ed519a3dcf1f84f39b680740987efad7fcdc2be966149eff2d
ze123f0bca5173840822a6991351a9ab7952a936873b1b04bcf18aaf855f145bc63efed9f77dd43
z7aa66cc80837b1d64e4635de61b9e7afb7a21dd12f481f5ad1994b8fdf8aa8458d6395aed552ae
z6314688767644d5bd6b3b807d2cb18a3063d8249834847ac832dab60e8e99134c8ea9be2b5b0cd
ze52cbd259ac18268e792560c64578b96f9096bdbe9db9b2fa734ab2a184ee4b4eed75ada610381
zee3c37b4218faca407b24cf556f7fd51d5935a9765010cf2aedfe1e2eb27f27d414b53bab026d7
zb9bd000d142e31578aec2acc0110a201909eeb093808aca25108fc26afbab8ca65690bacf501dd
z0b7a7d82fd79e34f471a8cf6870226dc340966ceff75c9c0501debc74ac51b6c6f8b8264be70ca
zad03a2615fe611b0d3e3c683c86e27c8e5e0a389b1d5d73a3f3f075d715d4db7ad4b35b1db228c
z82304009662f7beb73cec3694eea837f8535b354ae7562b57b3b6d144a0041274c2ae3c49e1d38
z5db6447591c06c509d261d4f27ea05e5ff410f31f38fb08f137510558011e24c2ec6bcd66566a8
zb4f7e6b0ace147814fd07b27d51dc14be05a4971b7e4deb9f05e32cd571b2d006674c690329290
zb865fcf2c510df0b87b9d98e24f18b4832771440f91940d1be21c055539b81923e5e4563e07d3b
z87b2e8da3a68b97c416f0d7a59a16eec69a9774ceef7556f1d6f5eb63e5e1fd3cc7cbd46a5f4f5
z83457611d93050d38b1bd3701a7ba824dd7de45f8bec1c50691cd781f867b94189cc9067c2500e
z10a3b4e324c1cca4697394147379a132c29613cadbb26c69ad15d91c67c2dba0a2153a2e347433
z656657a2f15f0cc1ce4a047974b7d301044fa78c2f1c735620901acc1c59f97352fe2103619657
z1b379441e634eb9823897ef12422227a465d4430b2f4bcdcc465bf0e731c9efc6f8b368cb97ca0
zdc1f66fcb4e562fb0dbd0943422c7f70a3ff2b4c80f25bb30bdf513bc2cd99486e7bbdfb6be34d
z8bbf4b8d1faaff0a9ddebce016ea86aaf8f689f2849fd04364b61e681de7e359cb7673ffb18093
z4692bb1f6a03c46e48339328484d05ba60084501e19ea6144e6ab1997d15ef43bc36dd91990fe2
za134a4c949218bcd86eb065a6a156faff7361f3dc5a6a15703da9958b7b8e2f2e049ac24c65fdd
zf551f2dd69a7eeabb9341421ab805ad5db2fb92ddc127016754fadcfecbeeb314d6812a63087ee
zeb7815a6cdaab2153486f80675d7edc2ed182953232ae63d5a680b60ceb3b5c1d10d45fcb86a79
z11297e735b3a71b5896a7b8d6dde50fb1b0b7a2662795a7a47f982f19e28e59e84589687bc2906
z8ce9e1e5cff60fb540e12169c999dbdf976df8fd9c6d14b556bb5b08b3231d177da9d69716fa94
z728698d4278b9f10d4f1eca318c312a1a5b2b5b1fc3665d3b7b530bafefd6cc992a3a79d3b261b
z821230966861c69527f1b280a7ef83d2611fd613b7cef45cb57d14e3fb7d129359ca65a032236f
z5112094a7758ecac49b45016544752d4bc6fb0c5a401e05dc3c121dd27e4776ec7844d3dee06e6
z3a5f6e04d9eacd4c584147787391018c5173ea0466445253d8cac006e7c3add66ed06b8841707c
z330228a6ddffb3f87625bf5bd31ac0f11b4bbec2831898afad07e2d606140c0f4e0db6f0cfc7e0
z56c744a8d7de6406a5526c754a29bfedcf3fa721d327eced05fa3a5e0dc99439beddff88364aac
zc0b45faad5f04124d92d9615a1f3077a3d691b39d929d5a7a62ade27e45fd79e4a6ce3363c0163
zb19ef7826828fd0cf34c42077b86c0a2db08c052acc751730d6ba23435f1704aa48bebaa304b89
zcacf0e1ddcae82fd8dbeb9ca394e0d8843644328effacc8b17fab5910016511c1a2b37e4731c1b
zf47cabd1574fa2355dce36a1ee66fa5d2a0ac821660f1487915a8be427860285c9d570369357e6
z96985ffb3c71f219a5dba7ceca58a71e68f671a89bf18a8bb3be41e571d8cea17a62c347ae7721
z3105617c15d4017c3b143959914bb9aee433ebee7c970156bef4c01f195d5430206257ef4e6d25
z97cd78b294952be82d385537cc2d168034a27fb50c3e6ed1874375e8cebd2a945a213a4f96803f
z3a710aab6ff31c4780dfc70d69e2a9140e84b2a910148f3842a0f7c19f53cd42056997b46623de
zc61265d17ff506ac162469002dac53f1a425d796b54a3b8febb206c04138da5e1015f3bdc19ac8
z7de0f8d1ce63a470613f0131c91ddbbcfa785b7f7d46088c2a0b8a296383df57b4c99e1324a188
z45c52276f8e90a18ecb26119cf0d3aa4817437c0bbfb3d9bcfcb06b147ae8852913a1fc4d21f75
zedcc4bdfce7068d516186d5b3dc2f699ee7a1a79bf15b2710ea0a2453d9bd36094cb61f36db376
zdb75d28eaa8e2380aea53338bfc945f109ec87b82285af17fa6791e58aa4d24c82a59bdd6865d2
z0825df62cc66f485907da178c91519311241eba4f735f0c19e8c8adb7a8423bf380ee986ddbd01
z1626826677e051300767c500a2d7dc3cda46a1087c952bee967304a436529811456f2b589403f0
za00d05b9d7be174c0ccfd166c058deb3aceae813ec3e4d83ae2dd31744586c77fcb4c5e6d843c7
za58ef04088140ece4abff68084bbd2cc35997555361873f6d9cf90ab7dd600945723ba95100393
z3e4980998f143a1ff703efc64e5d62ee291b077daf331c8b7a6266fc4bb3f29d28a2a53c7b75d4
z0b5ced8e90fcd40ba23d0907c103b0ffdc7d6f4a9426695f276ccd73373a50939d90a0520469ce
zfd19af8673ca8f3ee1b70482ff32a54590eb57ff61251497b83ac234376547a34828176a97a752
z19695c7c20995763711adc44ed4685cd88d959559bce48a34a10188aff3f60e6905e9b9cc0a618
z2a38bbc4f85814e6d1762d543cc37dc163868630aec6edf767332cb4f8264f85ae08fcc0a334b5
z2d74def36f2cfef76f7f41d70e183b05a823a28c065134cab2add679f4e1dca1655fb44f5f3a80
zab03790ac2885940c62e91abb27bb386ebe7af037ce9f87364bc2dfbefdaa4d94eb40091c111ab
z777d7e3b7a95368abbd02665cf52574274f9b98188251126d54eb906b7a8ffc2c4253e842d64e5
za63c21a3dca42b3825f2e505537343e7c6d5c3d3be74c83d142f613296192f2b0b41e5ccee61cd
z51de6cd6bb49831ee9aa5acbd2897ae178eadee3925b4db9f6dab88bc8e49e612e0cb5ed537fa0
z32aca8920c9150a23f49306bf0f37a1c96b7e24304793d887ec4f9633a47c90baa30d75981eb46
zb92cc44ac622936cf7e98253dbb0520c40a000c9d6938653b30d6532c8fb956c669a7df17c2a8b
z0afb796fb348f84ad16c83a1f50a6c7b6290581ab56069173331ce23f1b5ed708f8146078c3ca8
za94caebcd6b4503684041bd3497304787ccbe11341b5cc244b56809443961705dc7f36de0db1af
zcd8074ebb97ca9153b48887a4cb3bdef19eb879a392dba6244782ef5fdf77f0143afcbd665d8a2
zf5e0a9d1dbf12ef0cd2e1abe4e24cfd99a81488942ff758a5f1405d7ee163b71e3295cbd125b42
z5d70f0e0e047ef675d1c6ccd3134350ae2c8452b75559f271f5795b0f4c362c62eb30a56dd2be8
zc56115441e68a460a316a433c252b36aab4b6866ae8dc624de51b1678883a159d5212325022044
zab3ab8b69d7deeb96970d9e5f385353330bd4588f3acf348bc17e29ef78bfdee0dfe1fc3e3bd7f
z80a197986d0dfe0763a08dad6d1b9269e7e0125e9bb853d643f08c18706d210c382fd41397b409
z6c37873ad76f41392db456cdfbc18dcbaa8efbfaf10c30f01012f4f2bc132823d49657819e8940
zd4463b4dadcfd347d92d766443b04b740c233da7710350f08e862e895ebb8c395cde4947ab5b2c
z57a0b964da4553364f5885372aa8520f8cefe19f3a587d67a867985586318f0be6cd3b58919138
z78d57a0be6b11abd65a574d9e12fbee44ce7c3771cc22208b6f6af9ab0bcde96474e6e4e15a56e
zdc817b1bede66f07e080aed9038aa03e75274ff46670fe18054d8fc64fdee961cb11f49a8e93f0
z0bbe7692d45788b31daee735e1ae9e388082fb737fe92c4ad4184391e2b25a5836012881d97139
z86e98c947f01ca488a103cba233bf09199783c9dd7aaf54c1275060c7a302c83350a70c0385101
z4cf154916576f6070756b2d631405108c419d190dbf288f0307e050f22c2986ddfd9a3c59b654f
zaa9d15f7fa7460c75bf5a0e48d4b3264f76191c0665be21e3e7c5308ac30497b23e09d1e0e3c61
z1efe4c7264de76168670988837d92fada172884d983ba40800b2964277fd33bd36e9fe4dbcf8ff
z24c073c1fed32eff9f3c767f1a6702a6cf5a05ed6abff7ebe2f6a255392124119ac7ea2df718eb
ze7c04b9111dd76ac6f67357887ca23151759fb4aa955134f5582247221a8d04a8bce3145422c45
ze567b9961dcd20311a6cbe502587c79fd22dbb0243e85c43f671a3de00f593548e49368477b982
zdb6e2377495efdc9db9224b6ce22f9089513e6d3cdff23fc6cf45eece9cb77781b57ae8f4197e4
z8aa0acc6a7308c681724219d2201a0a730124618a84d17020f2b43632309cce7bb186e4b2aea04
zc397c579659b147dc4d5ee0d93734c7d7febe583e29cf69a3aad847156eb6d93f81dc428db90b4
z03bf893186213572456651919ec2435558ca51ed2d54444d3745c3ce697616b768968c604c5fe9
z0a540eb7c8ca304dcc2ee3030f2bface671aeb366d596fcf1366a8dbcbcb9abd7998707253e787
zc8ddb03e29993d21180ccc51c313e1e60e3f5f2acb05d1ab01ffc1e437665d523f87dce26d1df8
z2b52bf269c8083899365786ae0faebb1a69fb0938c557776c6b0b9e74034c443676320eb720b5f
zce21a5298ea5d1409e210c31b0e76efa485a71b3381a96bedd144e2bfaba01fa9087cdd0e48fc3
z19ada8b1fa40e5d73c004419468833fef956ceeca64700367f6d4e16afb49739f87f6c26979994
z27c6aa2d18e9e23c42b83bde826cfac1cc523f11c954d7fcf542d947f9fbcbffb1c33a42921e1e
zd9c20d20d56adc8dab300b1d428ab31a4ad73ba68636f088a00f4813bef8a369a99583a899e9b1
z39a37777c676acf94fb67e7a5262e7860a8cda604159245e3f5b134ca63bdb2e65f96e3e1bb366
z51a7cbfe43b950895267482c4417ed95cf752bbe8a3452e5aee852b976ce79a8d5a9c1759b061f
z38a9bb7a430e574c208e84ae9a57b45fc233af53f1bb98dd50ce05e9a6e4f4c0efa9d33bad9674
z57571b5b07d25da681eff8be61a9e79afaa71bd1f695e5805465d21f520c22f52c55a9352c4448
zbbee921a92628bc81ab1132ee0d30e627ae8fd4102d3bf570199336cd39cf9385a969639fa4937
z5b309e81c43198fd693619543cf52f09df5420730f80b5778e9ae8284d0e8061e93db92f6ec6f7
z84b62505391eaf10a11b2ff7cc6f7df4535ae28b915186370cfaacdbff1331837d97f49f7b0079
z8b94f2d102a2466ea11d29cef4ce4b8cb48bb63f71e68a534bf114748456b39560a3c1594db179
zaf89f42ca4cfda3650bbccdf87fcc6f18a2d69dbb186c1248a6a13468d55d5a158afc0b42e3966
z9957f3da9134e3dc54250322e3902d1cc18c6f7c824c084ba1b42944b45bd268b0c1c58241495c
z54c5e589ac21a2cb4c3a70bd19a61fecf95d57addb9b400588f38bf42596ef77dd62f8002611c5
zc6bc7ae20b15cbab0ccd96b1bff1e20f71b95bde3ea4e2b1d3402e75c020a3b73d1ad1fd34b4a4
z40892fc355b8d70c05ff28940cff3bf3e8c37468a19be50bd6858bc1bb3af62bdc3b37321e216e
z7183af48cf013ffdd89b20951ca0751bbc29e271ae2a24eff2c660d151486b2a9cc86537bb25bf
zb8058051a89820c4e5c10e0c037afb7bcecf780786714bb86707ab840587cccf05b7f38fb894a8
z7ea40de918651a281c4197f038b9739056d1596c448d6491739582179e6cd62e590f11cf8e983f
ze20a02459439a4e46fb18d34ee9380d94c1a5e24db8c5374f6a1dd20bebab21b3fff7b38590a94
z72b0ca0c6601070488d18cff5907735cbeac37351ba428dd911d64455a0c6ff2eac28ac430b17a
z8eddd94cf88647baf1177268c157c954173c2e239abeb9556acb8d32fb16aa5e2d738ef569c5c5
z4a74f791f5a019f486f7df99aa38081fd2faec4219a66d8b31de96dac35caeee40d1560dacb74a
z59ed3ad0184f438c9472036be4370672beabd7bab05975b2b520def1ed2413af0e8cf5a31aae01
zb3ea096201b8ab3abb36779c9b20be8131df72f2aa95170aeb1f4ad05bc0c48f600c8b1a043326
z9c112a1cf8ed98795eba00b63d6a7175591444b67f31c9f47e6e48a7e1fb20cd5ecbe0567549aa
z5ee82dd86b574068e0868306f5c80d50fd9a9410ffddca2a01ec182a9dcb1013d6c120c2ef6c97
za08058408d2b8239f32a39e6e85522f8544eb496037ca268e17a693f7c18e53bde7c01fe20d59f
zfa3e184e85be41ad7e5ef74601c6d1557ae0beb7a0352f41ac8e948d639d944c5e201b8b20417c
zf3cbae82601092d6d6777d92699483dbf13f839b442c86b011ad9a134802e88eeb26891eb286e6
zd57c8ee56fc9bc0f07448c09ac42885b0f3abc93dc5d85bc3ea3464edc52127acb3ea6b6c983ae
z0795a37da7299f0cfdda958a0659a4b644407b5d3baabdded4cfd58b4a7e824ba9805d387f6727
zda45312eaeec23d043093da29a752ba1f89cda881bc86d6bca027acaf8d11194e31bfca848aade
z49925496872eed47764e2b00185beded029b69a316bfaa8bfbe8449723332332042a8b139722a9
zce306671ed9ea03e1d60d443007dfa84dce611bfb331bd31ddd831d246d599f3a5f6c94d51ba44
z56d92eb4249ff9da07146a392c1db32dbc9f603521a7c1581f363ccfe1c2eaa3a8ccc0572483cf
ze1145fd853b6e1525f8f7c84f0c090258ab55c0c264edc230ab8cb5d1487ea28758ea638815e28
z070f6f8bc6f2e383aeb64d0460964901988a2155ed0c67a322def379b6ddeff536b9554406d23a
z786b07e8fcb97fc24cd563405e643b3ebca1918c0df285e9a8c50508ae60e08270a31d8273e463
zda02c73acfb833eea80ca7273d1ba228c878084319577cfbb750ae42453b7f5ec0eb702fd610bf
z6e86b00418aa4c869bca084dc9d303931489884ef181e45d2792e5a0e972a3305084cf13e6b0be
zffb28e04d6b4ed3ebf5195829e89ce41cd0c9c288429824ee6b3695e616fc3ce93956aaa462e20
zfa6ac0d5fd3789c9c023b5b31e02e330f17b9e520dc2c080bca255d4b4dd3bf1d6ba33cf0198eb
zf71091bcde4ec3071d7bbb667f2d148dd261c524674b656f46c82f6317daea81151b8b51ec22aa
zebb96b67cb59e74a7b52e03c12c1d4cdf4554415626188006879c516b21b846d25adc8b378adce
zc90820c03248b83407d7a8f1114512e955661f1a4176b6553894656e803d29f8d77c6b4c0c3106
z7ad0139cfcdf322efb70b13975eab2a8767ccc51b5e6a87e5aef51670248a63a7bedc2235d0cf0
zf0b44588a1459c5c3ef34577afae277fd981c103101ea5b7c2d77d3093080265f9fd87d09e1c1d
z782bf392e5dc4233d91d4c91dbd5bd983a9b6be098938cc6078f8d3b67ff485dc263732198d2cf
z9330d252e51f737c8137c5b6dce908f2302f20ab4938d7b68bf32fe38a3f7859ef7b6bab697274
z218b00e647d823dceaa2afbb3066e6ca91a14c76ff37314c774be613b0a045f60a11913515ae55
z9d813d7bf44012ec1c86dc503004ff414480704f4a09f7b4b2b029a9ebc192713e7a761243ac57
z991effd5fbb18dfaad7ef66f1ea51eee94bf0a1c3c7e21d233d9373efe66e2d5d397e7a77567af
z9f243ddfaa96ec686ff0dbe0ee55e2cbc4a53c79e6e0cc71f937f76fe82538779ab8fd488defda
z199d3f23d9a94cd61edfd82db32854279c4bb06336bcef7ed5d7b2c8f0fa6804bfb71b3ce75c52
z5227675d582713696ae77093f92f4dc80ccbcf7af3e4b9eba96c08e9f4e0ea41bfc4808fe08a64
zc352e845e7a7a1520e2f3182fa964e088c2763fb9f6f585809db6cec437702672b479ba7ff9ac0
zf72273a57c29119262c4c1b7230fcf08a99819d72a0157e367b22a1691562cf66f78d570c0f6a8
zcbd5a1b2309dec689afa4be29e8b520f7d00c4927da6a057ca0116565daebe79f7fd89e28b8de4
zb3dbbb1cce7e7bae5f1f836e3451a6d9dbf6a5dbba2c700a1be8b74b041faa5446304c964c9723
z06109905b558a0c758ebf386dedb82a92764b631c8f638ebd17af9011a697ccb2b24862f3590a7
z5b5290ca7735f48fc4c99177f3956384a9ed285e6c477ace4ffcdf34b6eccae624c93680670d92
zea0342f812cd0658f38c0a71edaddbdd8fe489642cf3a0530566f4d2e352391703eaf7d4e7b7f2
z920bdcc2b866e6f56b35110c4379e7e7b4e02313856e4475c4c2bbd17608389488867d087bc478
z035b84f618954584686b07b3c80903e10b596980ebb070043ed2c1fe481df52db3005078c57d31
zffb4152c2f88fb8b58f0b7f33f35e89c6cd77ebaf64b8e75dae60016edbafe988e751276ccfdbf
z8c4967021d34d852d73e65ffa30cc1141e8face6d3f8fb958d499440a168d729455c39cbe1a56e
z835308ba1097d26d90dc619b1e7d22c246dfc7ac20097cf4b73bb5a76bfc7c2945edaa8c506379
z467bd9d24fc304c9a62701d90f70a3dd7e6ef48626867cc223df40aa19faac1f42e7a6cd53ec7b
zacb1d52989c82e8abfe126199b514eb4943a8c0446dae15d48a7c93d40871ade414d99cd3e6989
z26568f0e139a7c8731fa7b2f9a09fc193e1dceb16ae452367f80308317ec2f1a7cebc0f3428179
z62c2784ff32dfbb73b27f83cffc2f869e1116d2df46cd3b546861da07b77b8c19a1456161ae9ac
ze6db87b1f8909004ed475e91cb273c8a2044534105f0ca3788cd7b884522b40fc5857e9584d078
z05028e7b14973fa1112652844cb86619dce35d66a0aa77a5f61668e64980512d426ff81ec48c15
z46052fb8ea20bcaa0a7be4307d4acedba011c2e78a3610d7dc99e342a9634fd3e23f4a04f5573e
z2614a80de0a4dc25ebb32110bcced17e6ffe49e2c5f234a45034792f8019056e20497ba480fd0f
zdacd441c68c33b8e431a9a48f07e390a82e2cfeb7e0efee81e771bdddd02d8d8eef6526f1f9822
zc509d8509cf472a5b7f2446d5141e06efc689519d17241ad07c4f226655d3ef45524ebf664bd78
zb59ab1ff42052e2ac77b62550048633a30d05b8fd685d3cbc01bc6381a1609fcfa6bfea21fc2ad
zfb5eebc85d0bad688c27f39776fc25467bbc0f9a5c4a0da3f345fa2976a144c8c9418cdcbd7841
z40b440ad2fc24335dacf8ca1b366411bad39ce7b7f8a240f4e047a67121985e9702401961f6c02
z9be86e3199bf8559a29f3c7810b98cb41ec8e31eb382df3c4085d80b4a745b54188a02dc6d53ce
zfcf4fe5cafda2ed2e121b22b679b338fa58a8579aa643b025ced309022ef6c23247791e2362177
zdb5be687fe86c2e8608d0c6bac3ef9925f680cdee084a05adf5f7c64557c24e5c3c7025b110ec7
z2cfc6857752f4b4911c5e1947b5f2050f0156b27d264ccc34ae6986a76dbcbbf9d535bd7897934
zde9d7970ecafa14acb390592a7596dbcec30e6b7e4d2ba3b389b82227f15460183ef83c7f71a68
z1403a55cf4ff14c55d10365c9451dc4732ef2cfd474ebdb034788090afcfa49cee9c04a8f5fbcf
z038adc1855025f8ac0e4ea825ac3f2146073ed5fc886845c6c7158f2074799de5616be9be43430
zd79e5da0966527789aee5b432202ed49eaac1ac1c6baf9a9c42653af5af6a8512c2dcc1444873e
zb4a7b032c0b71c4769d5b6bf139c6de2e2a6d7f603a12ff62cc16d4145b00a28846be1056ca054
z22baa0f90815e94ae14549285e061491137e3fd8d68880fad46fa6846b08f905314f9746daa626
z33647d3db24c2d25d67fa09c8420556b433c77b9feec2bb70bb57a17b6b9be1775a10a31a228b4
z1df7ca05632ad2c334bceade55e4b85855ad6d149aa897895e791989ef3847e5d03f7cd78acf94
z28ec406b997e0ff8693976de881dd5705e4c30264551996648f6dd50e9f98ad7baccd69e3cb2c3
zdc138bb2e5d8b72633e9e063edd76d8bb34d33677cfe46c906319206d8a5090a5d797027e74918
zf4a5e697a8f2ca2c18d7f48c97b79583b2a30d95291e8b69d82dc9207330ed4fd49d3a13367585
za444e9f55c957cc0b24e273479b26f5c7be516fa03411b7a3d69a8652201cbf5af9c61895ea87b
z8c8540e4346f9e246e81064e1f11896f8e0a26807b539dfdfb5ce3c337094de7d0ce88ab8d88c9
zbcd39d6bf8189fad435c72a68fb68d111fd02a893b6d0945f48d2e7f16a405bff3b31e37e0d2ab
z6cbd756b7f43f49aad1cad88f75ca9aa069e8d288a7942883a5c6208c8c30adab8a44077825013
z4f2d3dbadc94c01504736904dc8d5921a941bd7d8057e4f8f1ddcbea081e93fd403f7f5ba6657b
z75cd19fdf0590c3534b93667604831b94681a2182c9e6d619c54c0eec702e3bc0a3d8793d79340
zf9b69e1334f1c58732224ae08bc042b914fff7223edad2a1bc185d64496c4d2a741e4eb91261b0
z145f46b0c76ce09e3690de6f3598902df28d159ff7eda96ac4960a671e0f4db779e42bf05fde4e
zdce9b54d07e173f300a4aaaa810f5c69138ba682cc23a03e67d30537084262bf07c5024378b652
zd7ac15c5bedc6a5ebc9a170db4f0d02a2ef5c48b4d458311a82a89867d442211d8cdd0121feccc
z1b49fe74793c17d113ed13566721998df6017062e489fb7a6b3be7eb97645180aa22264ab7c566
ze2cffed26bf82d9403a04ca5e59513336802a7680ad505e3bf9527c201948a703aea6185a307f3
z1fa57d3cf6c6c1b1a82295720d805284dd0bbabfa4ca01b53169bef91d58e2bdc4d0f867090b97
zfa02ffdae8c1972df4c2f9ea48f961a106d9136be3546b02de306ac40110c32e7bcd098a89b4da
za216828bb24db9f92336b1128567f530e9cbbcd14afc5471695bd51d42f0f988bf0050cae925ce
z95060129e083b192e87721d6752fe73aaeccc6a66a831a987bafa2cb54b09ae70fc745c9fd88b1
z2a4e15eb764c3d708cf04b4c691e8cb4c56ff3b5cdd9f8ae8618dee22ea433e042609e34c61332
z4217c65537ffb6d8ab9a3fe5e2f0943af3335324bf2dc6cee4941219600c1eb71cbde8634a9cb8
z75d50e070471cf21d38c38722bce9d6ea4108d922c5dda91dd00ba154059e3172ec40cc59d933c
zfa231425d629fe8c89247491661d2c3fbcd0b04302f3d264550c7d9c0126eda295fee7077860bf
zd78f118b8b38870b3878639f850973ee4c33ae367811e733b447bd5c17ce5186007c306bb2206d
z07e9c32cc74c40e404d15bc2900c1ebf901b8c33606ee490b56abec317f0e06315de93b5fed046
z912fe07b9e08c224ef571ac65a42fa937f5dbb901ce33cc923f00ccc10c2acff0b9631f1f59a04
zea9ba7cfc4d1206718e76b47e893bfd8fedf1463da1fcc2d7bcc5b6e40c4efd30d4802639d0e46
zbcb00163f2ebde80bb707b3e908db0d88b7121233e78da7a76147e3ab64d3b7dae42f81fec1fc3
z74147de3ac1366fe82ed3303018f46fa566bf49f3df885babdeee27d660a325b57be23bee11fbc
zad457b18b01859aba7ed1a69cce3b7ad04598ab11eb43e0750a185ff0e8d97e42513b515f709c1
zabc6d472bf1f5916a3847b2b7d371830758c4ff6bd2737940f04a98bebcfc52bf9b180b6147bf5
z43ed4f237ef3e7c85c1d06672d7eccc449a8c133554249a72074314951a7c9eeaeb1f18fa9902d
zc340dd9cbb4a8b0b2ab0953f36a41e61b756488f66db7ab1e6d62c2c3cf7ee6c5054c994605967
z9eee36a3c39a271fb476addbbfa12d640c11c32798d103d5d258160b3174f39f7ba31b073e7ce9
z4972c30d482c55b469c3f7d43eda0b933120eba0145bb68a12d6bce47c3867054c4cc3d172ee85
zb4f562956728b20d203bae139b37daafe3f946668f50de43ab7e8ff9091780b9f623b6aa1a360c
z454f03617ff732a06243c1d14023af78fcc6710f53d90cbf37c394ab381fc553eba6846ee889c5
z5cf0c7903521f683a4d71459670903ca504be14343ef210a1f85ee074c13bd7debb4365f5bfe1b
z0def85a2423addcf7b093b7ead94827050f7f2b0e389fe76b8f1fb7044a42e3c3ed1a0e17345bb
z563c749de176b09415ad67491a6daab5b6a995b8db7b5efe7e46b7ebd877ade2634402fba56fdb
z476e48d90d21cda441adbce7ddb2a8cb40ced71498da9c44a6be48fcfe88f3adfa7d48fe3b4fd2
z474bfc6e9157582864dc0d7cc551c245340894c311bb9bddfa6538dde4796ece8588ed0c1eabd6
z46a5c6cd95efec12a56f5b2227ff293a8681acd5453be7651bab5a90310ba032ebcb2dbf87cd6d
z1d18fd34b85274a595810e917e79945a4544cf46f14ec5d05a5669e94dabb6a3dbeee3d96e6455
z89f838a060f6d58207c0f9926c6c3984303bd61a082a2a44bc4ec94b2f0397fffe75e29e0aa6d1
za076906e03bc73c5c6282cd5725794b64aa6e7ef922b44af3d5180f455e504b1304203d142a044
z506fa3e3674522b72ab981bf421d87aa1552cf58fd8365868c3a37dd329aa177f2fed209feb409
z9ab25fa6d622d77ea787c07e2e8d999d12b25ee5e4971cc65f6302f7befbd3586e7349ec72c63e
z3a179e9e7962fa0e84b638ab76f7c3d8c16f87865575958a5c489e0858788dcd7d619a571787e5
z2b618dc0063d144a9ec31340309c964be86bd1b99d8e4db37419d1de9b6198df8c36ef602c9abe
zde0ecab5e97c2160211c1a75ff72f78c78cc5b5c27a09dc90f8487b411ee047c15e37f3d150797
z5c47b2268ede3331371f93797a453ee33ae380e1bb9c4c91943dfeb6d4b411313bece85cdd28ab
z56cefa5a337af7699fe1d6478cdcd20ba8bde684d6c2fbd1bfa6daf5bcc23fae5ea5e424310841
z07b0e7dd6ca3fa9bcb0ad0a7e31e04f3d2b0b157cd368ca0c1d23727a55859875604cecc739e42
z2f17bc2f921d59426e19d73ad7216ed63c06d5d943fb1e9f93d2fb6a520c3cfa65478b128f47eb
z0886d4b06ae435b6a4694c4a8a9d2a9a8409a3b2c2efbe06b3b8c427b67c8862d6ac9200d24a4f
z332af0a379e2de76e1bc2f906d6f5c1d7526b6b200c2379badc4416623d15e8d21d3e8efb96c2c
zede5e321dc4ced5a0b8bbeff8a74dd3e0ae729f0dc17d8885ebc214f31033f15490a2bdcd31d5c
z5a56e759c6d1cfeed466e776a032107693334977d63124b0f1e271e7f2474db470f931f05b8496
z94b5dfe63eb66c23b328b57895b6adfc2dfdfa73c4eb2168b3d26eca9a587bc9c039660ce7152a
z7f00af07222801d15b426994565eb3ea29754608a02ca46b59238e144a6e1c85eee0a1b5b5494a
z5df51e88534ac7d0974531b831d0bf93f794d2fae8f72ae3671bb3e5585aeed7d6fb39706369d2
za8e6b6cc700fa517f879140672e26a604710f6385bb8a4757b9564d5d7ad4f517631085ef76b09
z9b4901251c6310e1b72a31592089898a59bb6b97c63ff970131648c1b0d62c6c2afddf7be3c5fa
z974374d9b3a11cd172fee0b7931392496d909b202fb1f2c0da56d4ab6a26dda3a92cc108f3dba5
zc1c4dd83408da4b25cd16956d5e50a92ec52d2e61ff62689d4fc4513c6ed5e69cb3ba231a6d222
za5c52bbfb45a1d62455e3f25738b24edbbf277910370930a2e5a90a79838328c023db16a4bd92d
zd89e5352f67b135369ea453f5bc37942173fd096a126694cf8ab0b1b8c1d4d9683ccfe71933119
z88226cc2609a41b4704ea33f2af472ff3e71b8857cf63e3679452d775d4ac4541fe851d4fa781c
z948da69e5bb8b0c6c6bd375ee315be839046552d7be0a9f0905df853d3b01b73bc897900b61c1a
zf49212bb29fdd09e3987d3cad9ed3efd7b0c938a123eed91b7af70239ed27d607cfda29f820ba8
z248967944982169cbe96b5bf70c1fe1b5bbb1113e61488c4708f3c9ce6d099160d6457e4349b02
z3864b8309eacbd66bebca05c0b71179f5f53eb8ae1b3ecc6f9b2d808ac65e1b9e736a9a099ca82
z9400d916c968f550cce271523b454a1415ce348d07a4716ca565f41eeef4e2b1cd8a8e1020555d
z4050f429a848de28db3955c6481ff5ec5fb5ce44fead4fd8421b1d3827d96910cbac2982241fe2
z459709c0252bcab55c66fa028d87fc96893a0e629efc5567fccf69b232d11227987de86ca2743e
zef0c93c673c1e0692f24faa5c3a613bbe79cfaffa6cf31450c48f9ab7b3d3746ee48da4882db4a
zd0370ba37fa232d1cf26c6dda32e7c0a61138e624fb5d4677379507af535848b9534e58b8a2109
z351237704f20b60101584a77fa73db6842a94591af15bdb9046bafb37985a034401b8ab933a8a7
z94815d261ba4ac0840354afc3ae9208102834b882dd0f6e86d3c771a0dce81ab196bd7e2c7f0d9
z60a2e0c088cc3e937e93ff8fce1e1535af3804679141da758018163867d2caca6fa0cf448c0c01
z417977b62df7713be659862b416389359f4b0a0304d5ae024f20a173b32831e82fca18f0b3856e
ze7337650a9625d65643d015dec368c89af4708080b66d5a0e849565cbdc19099a3133a17891c07
ze49075bf079a59c222babd07c3dd9333478d5226e9a5821973926dc8238a81b85a575c6642bc1f
z0dc87458bfdfaa37d5b5a393e53a4810b39dd4ca4256cfdc5546b3ae52b8a64eeb30fbb11aa96c
zbb8ea12e89dfaa178b28eae87533497067dbbc4593410572e4cb6d9acfd0b5f64c159fe6404731
z81e9cc5f5a01a48f92afbd0c889cca0e6bba9cb5753bbcb8b3193d5c62f4a6cc2590e1729d216d
z2602dac86d97a64f8377d3fc49f216988bd411a6f1cd1b08cfa1cd4f069ccb852d0520f34269fe
zadcf8a0b1faf66ab1c59221249491a2271db1fdff8ccf1769f79ccfcf1b82373413497ede3d5ba
z101450f1c782028e5a9ed64ee245b464936e7447705a4bbd39d5a08203010a598e404a1e75f17a
z6b87ae909f238b50e848bdd90d07d5ae0defe565438da84a2ec131fc88848b23539b6595a8c295
z2b7a1f8dd2fb2b23533a425e2463ba99aaa24097ed20a2e0179671a0c06298918f1da5378a418f
z24ceed0f154f95c5ca0360cb458a6561d5091124971ad5a334c56b8bdd4064daa85ce388781273
z18ceeb8c88952c41f39c51f8657b5fef60987e13869b671e94e1a652c5702a6d1a2e90a55513c5
z092f1140eed9fc2ef8dbc048a64db91f5a3def43ce9ea4fb3006c68e43ca294c436dfdc12932c0
zaff0cf61cac6e95fe1ec4d5553d43c5896ffba50d94939082b5cde7564a22b3c7c86e36e122301
zd837024dd002e30a12210eb18f8a3be5c30a19a07052a19d7335639e8b49118ba47f73224aa1ee
z9efea1a1e93f56914d33ee274791fb174c0467b891ca7ecbd8f0c025a44b1815e6b61f6f9ae239
zbe57bed741aa7307c56f41233d322d4d6c8bc163799b0f5731bf0c563fb83d35def43d4202260b
z4138484bd7bfdb007fa893eb8afff317d500e3e68d44b2fcd762f1e2c45a8373cc780a4e49fd27
z9b68d1f2ffbd739974945a0c7c065594f0063cc0522c4cf5850b516c7f4ec561112145276d2c98
z995f92e764b66df39410896954d41376beaf2e37d55c42d2e49cb85fe260a5281083ca53271a5c
zafa9931fa39c3ba939130c41419e412f9139aa38ddb94529cd4f0df7492cf459383c5d5522062c
z9642688d4624759c93f611b7e73c6e137d3a35267d5197dd07685b1e7307851c11676266404319
zf86d2e22dccde5b87da308ed40a59ab080c1f41371acf202af2066a14a6ae4946ca13a2e5721e2
z9811dcb9cda43205d5e45951a05b2d84dd07d3624ab26d687ebdb2b7467332d2a64cc264717270
z36b7efa8395300e9eeb9dccd3436f95f9d2bfbcf94fd22da0ef33e431ffbf344bf6fad14dbdb49
z07baef5ec188e34c05534e8511b96655dbfa9bb768c6d447325fbd3b29948e3f3bde954daa8487
z184a871a82b32c83fdcd751ecfcaf97c2dd5016f5efb7a3f71b4f130be4776927142286cee0121
z31898e0a707b969f9a5cae7f9e6ab0ee74a3eca5f1acf548b2958c4217c78cd1294031a68ad095
zac6f3f49b1484c20ef85bcec0eb4cdd2058028d8ee88d3d053f28068dd609607be0b4fcef469ef
z6cf7a7bb3d876a14498febf8f77e928857069b386c6f02880db58989d6a057771268fb16cf5892
z449eceff1c6f40f6a35e310ea2f5fa0a34d8d64387d93bd4d363e3cb47e9a246bc39661d96650c
za78865d276920fea1b1a7e1007fe72b8250268194be922aedd92fcfa96843dcdb5c473c697c665
za514619e36c668523b16146e3d03b64ed401d82109f2e97b0ff64d96315df2a06ea04fd9a92104
zecdce0087079251935480e3dbe9d9b3dd6fa6588668113e31c4ee1ea9f27e15e10aa36c6e1afc0
zd9a4c81fbb9b3b60d18f8aeebba5e077d757f209a6580d5242150a0718c07296ffa3d1c0afc466
zf93f857c71f3e361e348727bc6472029eda9f769d7d723c0397a9e34ed1a2a45064ddf8d0778e6
z171696bd4f2ab18b137589aff09fc52340df2adf3df3630e9e3a543339c9066dba8673b34e2ebd
z5a40dc79a5a3dc267e39ef3f70bcd8055e88bb40a414957d3a9f87a3aa15688762de7d645b01a3
zdfab0d8a36f13d8a07c77fe3cca2f15b46eefc2a9b2e572e4afabb59837014d1e508dd512754b8
z1850b4833085943c9febb9c498065e30456e3726880b5316b6824af05118a20484e86fb13689fa
zea5f0a38c7159152275cec3b154c5e954151a694918e39fdfc1553ffbdf5aadf79223c022e85e6
z74b8321c8194d6da24d21f04d674c605bece52569ade51272061ccfb8c0b2a5de8cbc941cfd770
za2144998a488e7b4fcfdeeed58dfd70205e23c48d0fb96529fc8e3b8a115a2e1bbb43e01f07721
z126a84a1e62429a48f1ba0e33fd464a8bf77c3ab89bc9159d446affbfcb961a0fe9287bec1137d
z90460d1e105290b20f743e4cb2a595bb643eb48b52d468fcbddbb5f344a73d46be3162f2f7decd
ze1fed0e40ecb20320df7b8b93c470c89c187a8c8b11d037cf565ee1a26f5900b5e592252e3c173
zb4ac48f7c1c6ca3b25f27349a6bc402b76f9d07d8133efa23a7e6dc22dd2dc9d06628fd025905d
zb7947ab274158289f966b26092223d9a25353d5503758165b6d58afb51706f6316afa74dd36af6
zbe1e79295eaf80f18c489bc172eb855eb5756964e46add9a664b3c53427f4604d0f80a83c13ff0
z8871ba20a8a781d20f5817bd3bdae5adbf2dacad06ec06843534b9c8f43863685a58f4d9f85013
z26739abba561a2c810d259a465cfea9bb767db91d253db8c6c67ff7fe7f3472f5babfc7495c618
z4a19bc163a3773ff43196d0c128834b7d57c39fe8116f75dc08c26390e74cffe3cbdc4d7300e88
zc9677fd87ef310b74a00ea56220a7255c91c08ce4de49774e568cc057de612f5124095f1aec7a1
z627c7c1179d3c83217247decb12ffe29f1dbcece4354ed5f42160d32b526fe0b542e79524612c5
z8341e92abb3cedd978987fbf02c252819d2c43f498140446e1c7f3ec8adb48b98d15e1b7f160fb
z633a9c0c9dccca7f23c5b7df31f22c35dee1f4ad080c363ed29d8043af745c4b7b89668a6659e5
z7d5578a4ac1f4e448428a6001a2f2dc1d4d979510b05bcdfd73ba630312dd4cc0792a6a080f5be
z0557fe3a88c0ad2f7fe86e38db29794ebfdde3b009d8f67ec582e604dab6fe5a4cd21827c46619
ze1501e79502916c0a0303fe1f52e25cc578f98e36bae0534a409406b3edcd53ef9ff4e7ae9899d
z7b4cb720bd1ca8c6055e858701612fd3e7def6e2b1b88ddd96a931fdf7c2764dfe73eeae795d18
z6e31c10b630eda7b7858c14fd68d988a895a32a544327c65c783e09d587d56f590d1c18a6f791e
zfa90d49e38357384275a73d1d63476925515a2c35cfef9f52a1d0cbccb7ef4af1105fbf799a59a
zd9272b6b450e2d2c267a747a2affd1e3d6d22abf5b8fe8f666491932fd88a3649877ae7fdecaa6
zb5eaab636c70662db21638e6701b653900e86750c2646969babb5f626df2641fbe29960ddbb70b
z4d56d27a6561fc2d7a829ef73c6adf66f3f18555e5ac14448b039fd4c3f9348276e7275e65c57c
zdc08594a858cbb0fe3270030209ae279cffdab060822359b126ff4cc34e511de87063c4de85108
z6c6808d9bc99a526b4c60d2f87a60d0dcaac3e81c65b8443823581bf948601fecf8ccb46cc1a9f
z1fb8b6a4e0655c0f26334955fa9c501db9d98d9f736609bb86ea331aa246e827b23b37eb1cf8a5
z2231b9da4ca9ec815b5ab8f10e9056330b7c79f4268ef2478e77d466a5df8040bac4421c29091b
zeebf51e6f3c09632f12810f8e91cde8f1fd27b6fb550430f8c5162de62de1558b92345d0566fc1
zf7afa5446286ac35037df4ef6cd14c5278f74175bf2c419532cac10a5c9a5e6e07d78d64dcd58a
z7964c277fade65f5dd07f04b042e46f022af6d1231933815c3b6d0554f438fb7a074a7bbb35496
zddde18cc102967d34d3b696fd5459256fa6dd0cfb48308592e4ff82d6a38f3115b1523a9e5c74c
z3932d1d31bca7786c98878f889337396a7fffee6ec2e91024718cc3bb9f0a049bddc383f09a9fd
zb9970f074bc17c156c00510f4ff3e2be34d702253bddc99034e6c150aaad960903f381a74637a0
zb105d43ba1419a3fe39e78afe86c09b8fa8e48c260549adb39417533d7e0fa58563928b5a5d6db
z442ca1e0a2f1894cdc27903340e577609213be33c699ae7fc864ee180b6d3ece0d3a3280480974
z815548ff76d6ca70cf204f28edf1f71e0d24d24a0a053d7b4ca58bfe63d7d1a226cc208afabfbf
z3b7118b179c1bb6db34c26003e67f24bfc16ef61e8d4de002f22592c2c844cd90d4cfdaace9ce2
zb95c4e08b5a3d63a78ab9929ce549d3962a1ab3da2f2ba7ecd2adfe3094f66b4b3a13fde5d1fe2
z3712cc162bbb3dd08cb74bab1ede29c4070c2d3ec3121375e1122700bce28cb3c32ab9ce7fa97e
z6a3e4cad346393555589c1fe51f3046368f5b3a62502e2a111c7017cded850a6de573f26806edb
zb7c073a189f2d37a473decec4fd68c44a08077de4c08689dcb114d0c13b8bc91f91c6a00c1ba14
zb20b2da08e9473023e60400b32ba6b891e1620fb72e1b31ea6999d29cb04ba488c7f6e42c3a662
z9cc536d305ff577e176d7382e80c5f707dcc068bf00919b58dd3205276ffbe19b009d04b44aab1
z123228e28cc859c39b6b7f58ec695cc33418f01800f6712a60b15e441e2244baa1257bedaca859
z8231643029f216e5feae76feb0fa11142847bd0a39e48ad2e36a345a3e59e19881d2d0681fd9e9
z009cac4b3db3ebfa3d7cda7e0f93dbf1d3491e8535f0896f794fcbef314d0d27363e6a3fe19c9c
z45feae14b31eeab6f040e5a85de53274edec51d72f8a79603ccbede957178d6c5e69b97fafd7db
ze12b9ae5a3b5dba15fd7f896b9400b02943f788766684e5f48d86af7e8f65098853fcefe1b8db3
zb2a224219b12bf77036907126303eca5d56807bb8741cee45909ec44170d685fc6b67292c960e7
z4e7299a5421db42efae1f61fd3c3dccd411fbe4c3cbaa2b36b608354e892d629a0605e46f8f5ce
z473c5b07eedbdac138f122773769d0fb8379b4679ec76ae20f273ce29eafaa49e00aba6541498d
z8ba8c48b9ded1523e1df3bf8fb77538be3d65dcc847a7c130d8c431a855357f9de8167859ef3ac
z77789025fcf5880037c1bbe3227d3d374d31688e3c712edff3f14c5623af3ec62b06a231cb750d
z24ae6ec38dfdb0f0336313dcc751420a93b87eb972bbe169506bc968612fbab9879c66d13e7d73
z0fe164463c2342ed52ceb8ebed00e9faff4307d20a2576f40621df12079cd20893d6d08266d7ba
z2f957cff72decc9601efb6ea36e489d16e1e9ed6af07225faf1a4c933d6e8f416a09200c8527c1
z92934c38ae8c8bbcad26bd1da92c3843bf8adc8984de5f6f2cce4459a55487c8636b98e9d29542
z47b294270fc905a6d6724f19db3aa9cbcc2151710abb2b99a216c115f41e449715081298d7120e
zb781ac9d25e910a3c6bdf9221308efb5a781eab72cb5f51d9b3bf061ede8f05f559e14ab18d0e6
zaa9c916fa12ec38f65c931c9649ec6811d80e1b7f2f6585cdf1753ca16aedd1df98d929c9760ee
z7272dbd0385f9e897f080ae960640117749b63e9db0c5d59e52c1553b592ff46eef9153cf50361
z202d1b80c5d0e50ad01a9b952fc605c8041ff1c8cd9aa7ca0a939646a960f92e745833ab92ab75
za2d3d57178d14ebd357c1c93027caa642b84324c31759c0148fb908b378c42777f44405d23ab88
za52b825a1e9210c1649a258b857b6710b87af7b48918b4be3bf790cd10983654f94daee55ce17b
zbdc20c0b7059b31c940e257135f238fc1a5208777d9307d6933cc65dada9e39bf33848ae7283b8
zc514b931c37532289992c42c30aaaadba2bf1a591f26eead1a3e3b0511bf8a3a10a38088674ac0
z234c6563839d0815ba9ee62ca5ffa88b1883c3d0047a526923fa451428a03ed75b73a3a541e9d0
zf6158c6f2121a615ebf5d00f380c3970bfd793ca8dd7da6d32e6811f72b288ff2d513aa47805df
z73aec87000d2d0496d0a905c01c3659a49a5dc6b122a8018e69a3bba1cc37cdee83fd2f041a7e0
zf70f9f70953c3eb37faf20ca8f2c103d2c1ce9f0d72908147c6695fb966f43aafbcbf7a96ca21d
zc32bdd4986d45a2a9bd3b483fa5d9d3b5a07cd65c37b7ab35594090b46e9ab8a4323da4c0ef4be
z45a2328d988a1d4db944b2f4b1af6c8ae5cc5ebef1e30ebb85e5b1672fb68281c245103c09ff88
z8a587edf29eac30b4e7761bebca68b897c573f763462809b367912a30cb2f6799ec32898c7e5b1
za78342a9c67fc90f60479877c9784f3b8cbbf14978971ba2a8fb9b1bdfbe1da9524fb4dc49c784
za9140dd7a44e304a39329676ad6d8335d7a7fe3221a441bcf7b1d887c961fcf971ca919a02c99a
zeb5f6c15b9f7fd2478563e6bded8439ca20d7b630d454aa27b9401a72bed1244e7e4f46da3edab
z904f07b38c9c1b60a270dfda9a12cd297825a7d79005118dbf9a30fd9e42b902c323f1e6cb283a
zfaf574844737d4c56d0cc67a52e5ab3b0623241217c5aa4e99bee05325b37233d513824a01346f
za96ef69384141333979d62dfca5cb7be5a234edcb1318cd88af251626f52987c3d6bbea883ba84
z9077420d335161cf45211d0622841010471db246d690dc1fd7f60615084ea3b196fb6d0f29b3cc
z223134110c6ccfbd2a52db5e204b9e8942ec1ef4488f448263c5ead16a89f1214fed7d78951157
zb024b7451281a52bbe3390d83880c5ceda863ff7a8c4784e74fb317adca2bf83f0c0ca14b50c05
za4743bbe2dfbeeba7a9fba37baa0196ebd090cb7a627b5956e7368f9d4908b09eab13ce8b4191e
z13847264a46cceb107bf887bfc521863e4f8686f863e05dadcd4e3c0c19e543772cabf34722581
z5ecf4c4ebae7020e00a12258588f54db1e50cd9f72939555f78770c686f045375c9f19670bfe98
zeae622d7cbe669c3f7ba56165a206e45715e092fe0d9fb8de5375e9900b31b148b878c937b2c16
z48411f36582d17c3dd410351b442be51773bbc69c8008b9bb1654457e3dd8953907e26a8e030d5
z91cac3dada79a0351ad98458a0021020c2df33c41d06d3787e6aa54f8a29de49a83a32d295ce01
z76f8db1f8ce086ba1927fd19fbb6eff4d5ca657e9cbc90298c9de4fbc3a25cacf77fa410771b27
z3738b1ea6fe97935e3fee6f040fb3ae474f609049847f6dca6f6cbb780ff0bebcb533ba7c37789
z94342dc2a3f914a96bb99e6d8add9c0203e94c3c972c684d25e30e6d123511088020dc1a9e4bda
z0121e62d04879818508cf2e5a3d8660f06e44b56f4cbb36a55880ec66663360f2a694e16554f29
z4f7b22a604bd8c04a04ea701f992a624ac6e67af30bcf12a78257470563ddcb30cb47114624e37
ze07de7114bb6552249786a33717599e8e76dba414fa8ccfec0caa37fbf1c679b8726f86e2ba694
zfbaf435045977da4b3097d9cb0a0d696ee15232b3c0bbe8d4ba801742f1bfc88911041c968ebd0
z581b0dcb938d44bbe0cef50ca39f5fbc89db245d0af703b8b360a31001ca5fd8a53eed55619daa
z086b14a767516a3d220d0da6064554b47c580fb98a23c62e54533736a7ff22f5918e19e4159403
z06d2356280bde0dc7a903c337673e9d2cb0b573e5f5277c82e61a61d27e47932688c86bd4a9288
z22af44db091622b50c4d5ee298a3e93cd4498e086a1643ae944ad4a31234e6c9ad757b1a2246f7
z19f6c8b744033671bea888cae90007a2a28c9917818839efd3dbb28b46109f4f61a9fe3f054896
zec58570e79545886a3d0a0aa113dc2a785440d823bdbbbe2d67b5c282317078f9e79425b04347b
z1b9eb487b091ba94dfaf1c94eddd3f4847f6d646cade229d8b6edaa891ac21e7d5354c0e8db695
z99d1e04aba6371cfc8586d11363b6316259c9b19b1957caa10ba174874ffed208c87345b01fb90
zb049e1363df25f91e32c3881f2c263b0144a653ff5bd6334c0d25801169df0ab3c5c08e76619ce
z6d92275633b3912d928e82a18a697e248843b760f86786cccbb07549b0578d06ea8679651cdad3
z1e0a2c34f28572050033a9430b189754eeaf3c0adb41d8bb17a8bb55670aac3ddf451676dd7a18
z8d0e788ba554509b9770760ef29395a75d30a87ccffb4eb434d32d697e480787a0774ca8ba7917
z3617b483fdc7f5d01b9a101723e4db79fa504cd5b5a49da5b09b4ebefb4d3567dbe46ed2955eaf
z3f69b3cb56060b1994f0bb918ff8002df9e1f3a232702c7e48656ada635158acdc212948b7024e
zd4e674d2098e77a02d66fe8bba1c1ef21777812f829e66360071b4957745bacedd6187350ae02b
z867ef4ebff4c1558c4d8909e169c6d8318015b3ac0dc3a56596bfba603262d11863df5e56de0c2
zf5046e4d292be0e0fe968968c573e7d5a1786e2ecbdc687802f576fbe098a93970bf7e480e2af1
z9b4a5a51e3e865d6b03615521dd28fe178177145db571720656f37f0c22a0cb2285e9ce9596a7b
z1a9413bab288e27855236cf2e17794b3c2315a98ca4116e6d5f27498e3086f5c2b6703b3df30e2
z393093941777d56d38b1af693ebd92746fd7d8d76c5dee960fcdc7235f0ccb0894d21d91d1e6f5
z88ee5243b928779ab6a4263860f30a5b5d8f76ca23f112e2f304c80df3dd0a1f19dd490027eb54
z945db5a2314fd8ca3cafb02ae38e0b4dc941f3338ef6cf3aedaa22ead0317d4ac6b94b47d9f24a
zfa90f933f22cd19cdb07c9323be2b23548ea760bc39b3b9cfdde5f552ab8f81c9f13851b8673b8
z16de04e97cd34a91006c0009d220a455f39d0a61fa8059a8715903ad173aee1f377cdda54b0e7c
z862b22ff326ea8360027a1aecc652b7a3520fe4a07045e2c2f2746fc2dbbc5b5dffb6f53482eed
z4e10189d80dffc951c68d9f1b50c2c9c8299fd03052acb462f8e20275bf294d45363bb73b867a0
z8d17d5398f932ea5a539c7e425524dd521d2f924572fa947ab5d58d3a72ca16c9308c60d538e80
zf214dab9ef7a47d1aeb8b7d8eb735b14495493609635ae66970b7a75873943d0cdb86ec5b62b56
z03aaf833f1f73022a74dcefaed0edf209c5b46b8eb8c8a3b9766c1484fcba147571584f27e9982
z45d8bb354936d10cc7293a2bf6327ac7f28de797fbd50c33134e9fe87bdda5ce51a3e3bcde29e7
z5586cc3becb191ec7c5c0d34947f03a90be0e4e50a0324e8affa9212c1f8e9ce0adf314b2069db
zf607c29bbca7ebe04e7330a2497c73bb22c30db68d0ecb888c7bff3e77cbe8ba2b018d4a7d1422
zc3de7826ce3a05d08f37bdd508b27fe181e86737aa168f009c84a8c5eddf14afeef6cbbc87aae1
z80bc5711fa70ef051264525921d443e12211d3f3456d2061c741239630a752b7566e6df3f31ed8
z936862eaa26132b42caa5c99218df6e9f577abf9782f0cf14a59e7acc3f55cb95631edd7c5654b
z231394208a32ad70d92e69fed6533fa19a91e6e9c14c76fca0634babb7a84edbab35d94342bf06
z1d663dba4ced56a49e2a97d2f22fcd924791454b9cb8e59b4d5d028160ce9c4b7c4d3d10c3828c
z024470cd5f84b9a83382ecf8e6c0b2592d797ab947c04e1ea90a7a0e15fdd84ca3ee783bb5dcc4
zc5b7b2b92765e8a0b77c0b221b5a8ca7f86335f30fc05e07e42eb3e4da7fb752bd53c178676458
z53c2a022a15e038737003e97e5e5ee3071d4bb1f5b1a3877b0f70fd8afee3d3d611db28851cdc9
z7f5077e4d986e6c404f924a1b89862b3cb32589960c6a7ec521ffb74f336c58c0777ae3a662e62
zdfae834c8e043125af87c6b7dd16f4a731836e035d043980f287f3016a37d2fb1351813ca261da
zd433834008836e9d366042213edc42895aa9852360d3c67a42fb0fbbc29b5cce5bf6c3558c0684
zb7fbe6a0b5e887b20d8a94b4f9f4cddd52fe1b568bfceb2321cae4bc1c8b7075bb29b69bd36b52
z40f4c7296fc61f36a57e13bd1460becad5ab60bb146d268280748c4e97d78c4e54489da5b3b02d
z1f483697f96e049b4b6b890a4a6b9d7b3fb82bc043a290d41cd0f3f3140b231d70a34a0ee5392f
zfe2e84397c656bc29da3f6d295bece02721c53507d0a40e627b0602bdb23dc58db2f9a1d16a3a0
zb9cd4ad8b4084897481ccfc54497bc8b9d3b922b03a576c3fdcd8349e81a1a486f96f8626863c3
z9f731725f8f054720bb8ba62cf73b58200f5c3069b74e03a71fb5a4884df8df1afe48150ce4d15
zf3fb926ce5a777909ce84d75cb5e4c9cd308784b08e81b8b4fce3a77025370ab4abfdbb62286ab
zc001ad3c55a11fef362cb3760b90d2bf95d9a8cc529dd0bef6fcdba3bfb9771de495aef75a5a21
zf64019a406f61940c05ac2b576af351eaeb9ff22e19a9979ab32c36e84c4fdd90c2ead860ba970
z4c42cd091de0c30b3077302882dd49373df28c6dce20f60b51502286d7be66f54c21610122cae3
z92b3df711825d8870a4e246350b1ae34edceb546aa162c199dd4881b4eca2d23fab3f74c8289ca
z4a621c73d7c1eb6b7d10a45b45ee6ecf1ff8a3bcae6c9b9418a5365288b70d066ff25b89f50f1c
z61167fe18a09fb0f097b3cc7ffde799120c6038f344a68d4279027066e2e730cc46db1ea1c78f3
z598ee37f7a71f2ef90895f9f12b243b0ccf710acc95a44debf882f2a8e1fa83aaa07fd36591a93
z919ee7c41dafce29c975609be854a9a8efd2dc4e0b8ff8f906733506e75d8855804cfbcb868cc8
z02d76c90836810bf18989417e698f6dea6974bf45adf5d0380b2dec8c18b5e72a38fd116b88cb8
zd316b2f22a65086d4cde44658fc86b8aa5e4477950f892dd6a01ba7a8bbfc3ee090eea674e5f8b
z89f12d704a6d73d8e47099ada66644b002e31008a587450abded3d92037a7a08eda64f8ed55520
z1d2cadc9915d9331197b6630470235dcf831f31a8641f4f0dc7e72bfc8b7bdedd315970417d535
z255b1ea36bf2e6316328b665be6358653b2146db6aa3a5212e1950064f1f93f3c3e4a8bc6ae8a6
z02ebce2df9ab0d4289119268f6b7e7336aef4ccea09154a3c606e6b89b44619adc17262576c064
zfb4bf4651c81b23cb5e7470e71c56ad86820e3f1be57cfc2ee5b0983754f9ead110488d8c585f9
z97987c800da06bbeeb76af583e6d22a15686beee3d336b94afb618eec1fba85da8ad95f79824f8
zf803b8dd989a1fc2830bfa177504e03860ac4ef9aff25865d464847e19e370d93b693f9d9f881b
z1c0681c8709a11704565e9d2d3fde1566e09e0d348542dd1c702a35fa1159c6aa8fee6b584f7c7
zb689c992d0d7478dac2947d81ba58cde6e4bd4d9370e89ef29395194048480456e1811ad8cb715
z81ecade8bcaacb9c3a3190ee6dc71d943d608bc1b52cf1787475b18f68738da518fafc556684cb
z9373124891ec7e42f8f718c96d6876f8d53ee5381d6c9660d3865551037f1f5133a710f12182a9
z222c9a0da463f43291656189a46a332907a586cce167f549fd9820b307b7b2abc8663bf84702cc
zdf454c4d499986b5c12885be4e15535bff8290cb34c4138806e83dba313ad965d06ed4b342e9d1
z4298368b9ab07ba9abcbb22d2efe7312c24a8bcbd0cb02bc57e3d96de476a161558e9c38b166a0
z562d6e0748bff513d4a7e3f311fae767fc3cf001ee4eabd186f8f6d907ceeeba0996691f6c8b28
z136379b2fa427a49df448f3462fb5be8f4760eff350cb19898e871954b187dbcb04da76db1e0b5
z79f2eb2ba032dab67bff5e5f56b62689561ff6ca2e844d7010882492c9bbd801fbb8145b1a5a18
z53b99c032b08fa0b9d276c45d7db18a14ee4cce97fa99775a14d84ca8202d64d2432739d6c0ba0
zcd0111f366eab2bb98f09e019ae1e165e62c6619c6d46b3a0944a7d3f82ec88ecfd6538ace6bbb
zc605b81829fc5f766e85eebedd30843b37ff5df98c5a6ed8e59d6cbd48203d75dd54fcbf3a8047
z8a436ba2e12ba12b05ff7d490faa0d33fdbd83f916690788d2d0ef41bc4c5d723ce75964658654
ze440298937df8546e104acd43fd8928631725c2813e7044b7a948517bb484fbfc8df4c47844186
z2d49c0f2dc4578fb179f0f2c53634b91c0fa3727365bcafac427031160ea347a5eaadac558df8e
z151d3b2ca8b7fcbad810c79b0e5f1fd74587cc6620b0d865f1441a0e01265cd1894fed705c1dd3
z5c11e4d508fddf27da7c51b1146ccd2bb6bf1e34e0b2211015fc6e8c472bf64b2ece0bbd78398e
z72882401e1bfd608fa1cd842835fa484bf97c10b98318f058d560fd2f23c3698acf4163ac6b579
z57815677ee2ff1e58634ea51a1b105d570d45700561d88399323620d6afd43fdab93efe696f1ae
zcd16e966fd39c795eddc8f7f04441efc0c18b5102e051b155f67b8150667ba6af3c0583a5e1c90
zbb55f8625c22f7cf8677c5ef734da8370d56e97b430a64d4004bb460443b89f7f6ceb917213b84
z189a0419ff05b0b1b99703b57b2b03c1ff113d6fbe530e6c494067499dfcc7f21ec12b98967fb2
z9ff23df8c339b64fe272ce9cc6f10c3418a00844b06c2b0c9ee3667dba81549cceed544536875c
zc19badb84b9d80c20f55c991046451f5faa01cf91bb98eb18e3c5d3db71dca4c99ca604ffedc39
z984db49497c8cffa7996c2c0c84560aed1a3d9e3cc629f60f244354bda598bc9df42b7d7e80de5
z48d90a1d1c3fc6ce69897257a6f2380db578e35eabd072761889ae02206cab373114836e10d142
z34675801473145572600881f5aa2a6e759e651a12ae7ab1f72ee32ed287d6babe2f7080983c5ce
z0ecfeea063cfc56e2034f1118d92cb0aaeef1076907945baffae75a34e3ee3370386a570286041
z8bf58d1597f4701f634cb86f87368aaec6596015e09fb44a06dcae9cb62b573808b9b6a8de23a2
z82909d4289358fee4d117a3a354ea87e5d74f54a76aba3b1f0e5d9c4cbd974a3ade17c54b495aa
ze17e13a47902e5b7b4e62d2624b4564a3879f2b7ad72c487925b5ef03d6a77326493226732c63f
zcb4d4a1c6b9e0e0f7f75687d71a3e025870e280652424048a30b0dfc45e34aad1386dbc7e1352b
z67f58bb8f5b018a9316c3fbc183aff1d856ab350b0745971734fe9135233c5fdc7c4d05c6fc420
z31282509e2acf29637cb9e0f074b41eaa31690f294e7396548d22d335619a86d9561ba2e6c7cec
zfba758f17e60780197d6f7bd5819ee4899dda5a99db526c9fd14b98381bdeeb7378eb6aa307159
zb9815daf1dd119beab7b4b64e286bdd980c5a8d9e0eca49997a73157733afdf3ffd850f6597b40
z39f2e1c99c04109a736d20707c969e8dc7fc614510c3a8497212acb835194b60126f90514d08f6
zd2c52b34365661d47d5c5e771bc2c5d9ab70f2704c9199323d7e25ea5af52762a930536c439712
zb00e7e3e5a34da35d6f7eaa63ba537a37b552b770ad29706a4f5d6b343283e109454d501afed95
ze0d8aae42a378db8d128a61fa19130206e5671681baf479c7f8469e69ba85b25400cf89ce30ec2
zd26f26b5a956ea8e1bdd2eabf0d4da5593ef2868c496c8cddb0471b2c3619d83b29f6fa59c67c3
z2795a1e3537a074842c08a0add8ac4b029ce40e6c136c386d2b87bc456945163f60fd306084c09
zffb3f45426105e73302a64ae7c44033f9c38536c27c40d1b6d04101da9907454cef9f2c43d4929
zc164ebde43127a9fc16ce83a7c6299c88d4a30da29abd6dbaa48e7728c503052a5d05d8fafef89
z72913de9087b17dc7fa4c701c690775ef3a3fca376190bcdda6065d26e417273af6b3f71dacf13
z3a4f72c0307c271b89c0f048865d8467d6008eab9dd25c29371406f450efc2dcbe15f27373e874
zb344bbed8750bbaff755dfed17b940fb578aee8a7b113edd219d61ff9121fa84dd488f778ff298
z2a2774d67a0f1969e64c1c88028b74f6af363a989b909215a65711278322d8abee44efb658a193
z99bd0a1a826a8718d3c0255ec9086f7b1611524e7821055249da5507f96f4b6b4074ee3aaf4ee0
z28f0b8fb19fe94a0fc5c18116d690f06d2419c1f53e3fa08d06112d7d5138a4094226694f3921c
za6fba97a98f8cbdc760ba2a749f84a08e6a27bc823b85561cca678029d22b4e72ec04c9f00937d
z06460ef19bf4865350fb97f06440bcee8c14d6d6a976402be52fec0bc8a2b441fe821bfdb00012
z41678fbe17eb0a7b6a6138efa45cfca4b0cb96fd6d156692d8ee3438dc95c73f5520d9ed69e4f7
zd3adfba63fdb57a71cc7fd5d30b82268dcd2b217edae6b1f121bea33ca1a4f8d3d137655e0a301
z7f44a43bc271d9b867fcd9e3a0db9feca4e21a549112c1e8d52bd2f734e5cb7cf1be386ffbd71e
z1b3c3d781956a4c491022c860960a8be43ab8d79b0009a5ab2f748d111cdc978a325fadde04eea
zb0bc859048018d8996915dc59bba9d4726aa21f37903a6e97fcf751f2f29c8427fd77187c751fd
zdf8780b6f325cb0ab631edfbe05f2664b282f666178d1284bd215dfa26f4f88d620cc82f6e35ce
za96ad375e48883826bcf4b1d7c0f890581c2850a5b16facb21834968deb2c6077060ffee2f85e5
z893f13338cf19716c30273d240372fa936dccf47bf90aa56750464fe30c99ff452923f0acdb7f6
za47e96c346fe0a26bb5b02328f11fdee90d5a18e96f45c47aa48a7d602ea02fa0c3243fa848fc5
za2c8fec4e5443a2ac428017093fd177d0228f721030b03e17ad49b3c993e72261a221f55015817
z74cab94f8abc471d2ebbdba13c39e9d74473c5619816f6eba33a612de19227f31c3eec3c1652c2
z36e4285efe0f0b6e3106bff820a631335e0cb28300bef53049b18dbdc742edeedc00b59ed3996e
zef1804fa74eadb610c20f5f62ed753816dcccc8b479558d0a33860567e5caea4f8cdce94fdd396
zb99e86981f3c29a2e1805740a0c4dacd9bf05904b1a7b631009e611c45af3666bb2db5304c3ea2
z754b458a87be0d36be68c9693ea332f35d0bee842a0ba07a14ae672999b11ca2b8209669e82f37
z9fe4d6390898b4088ac88580a01e4e5f2a40fb485561f447a2001aef73106acb2f553ab41c8ed6
z788fb8f31c66b3643d1451ab8ddd55a8639d5a04f469ec06db3d7c0ec84aa55bc261c804485b9e
z5de683738f9df32570be211187f7245bc79a929f9c6dcccff90e7b9bd8e615f9dd3fb97b471694
zcd6b9c3b889385508edffcdbdebc1e1e2a995a521fe51471178d5ed33d1dcd8e40653436a1317f
za81561cb93ac5cf27313b30103b485368126162f6a474a474c2a831b4104a3de7e0533fa3a5094
z8dc391c3169f18bf98f2ff5c1454c6308755a67665e1e75abd4bbdbdfd32fb91c8caf774139b8d
zb6c035e77328ac5fb129d68ff7ca8c686bd827937d5e698d905ba006a021ba3763d7641fecdc8b
z0b56601bcea530202e4ee9dd6b69e2763534b5a194c8d7989441abace53bd9660117fd9c5b7853
z90dcef1d0c06eed34bcd8ab7dd9a021ce3762f9e9c70d19ee93a894bec9734ecb2aff62652e5d9
z10fe287521b422d9c7c5786ad5b085c949fa7d8ab60a123ab398a2c6cb5f30c476f4e8f92b3afb
za66345cfb4f2a995d0a3bf76282f03bc639c0d83dda19c1cd0ceb9e4bbca3bcc0ed3f66673ffb0
z9e080d79f9b2ed336f28372d73173b8c6342ac1f87c7ec6107dc3bac085c2fa9df5151f32d9962
zd356e8e2a1428b379c4ee9855ffcae7dbe70183a79baa1098cec1058a8eed6606b6fb808e71d36
z95199a8aa1936252bf4616dd28ec3e6c387251747d6b4e5e5dbb5beb216fb4d155e98261ff5977
z7a097776ac1a1d3193f050e93568e9ac3d94cfcd8a148aff3309f86bd92990dc9ef83c46099a98
z911f4008794ee40a5731247f7fd650f9861471646f604f4d6c605658c78745c0c03431c6065747
zac5a4da865f81ab85b2ef701c43376c69535bdd9a91ff1da9082084a49ed8fdc01523e37cc24f1
zea75f53a3b6434c4f8408305dc559107bca02dec9db34436fea167cd58105127fd0dde4071f1c5
z7ecde2be26374f9b08ed3e9e9634fa6db17bdf118da09540aaa03008aca3605fae0abd8007b449
zc430ec4ac55c8d622b5d96824ce065db54577b669a38ab8d8d3d9a03b9ac0ccaba283b6994e93a
z3aef72bf9fb2ea62abedd0e7ebdc391045cd26ce547458bc083438f1f7d1489028bb49ca64f46d
z5b22d5c2f0a0c3f1d5836b058ec51145a4b262d4554ac3fb151941924c977e6dc1209875db6ae5
zf4d24015e4bccc1a416c449932fa9d3aec9fb38179d0e0d0004a08767146fae6dd5178ee5fb695
zc3897e8cd5fefd2960c777d65608c4a3a4e890a1f241f81376c37ca0f7a039f4f038c7e1029867
za9d09fc1805ed617d264d6f58bc846dbe62dc0a972532d650813a9378b43b1a91ed13efa7d139b
zdbb0158a9014dbfbe59e36420326e33f70eeda0a68d83348f8f21f7adb3eef0e5ca15fc613daba
zac6b85cc9322c854d4769cd2887576a4f306929e04c6f408be071972c56ec64e286955e4e66b94
ze60490114f752d65b35b382d5c9500020a15e17efff6c9f1bb5ac6319e6f8470d61b35c4c66271
zff030cf7d3f80ca570358e37c160d91025b158a932d5febb0a86947a175f87b421dba880e762e1
z565fbe4aa70635984b14063453a67ed221d74f4952c5c66c034ea73f3c336beb453091bd76174b
ze31d982a8dbe5dcc6e80d87ef514078dfba47a106beab14ab2299c25706aeaf4512ff9e02be472
z1f469c52e588124f07f4aab92827413a3b6d1aa76660d1020eca0c9c231a850238b98ecbf78922
zfb87782e125b429cf32d891795b4be1462566273facbff46e5b7310cebb7e4785a4ee4d17ca7d2
z5695917307ce63331359a6409d2abec88d29ce7bc24531f38dd172c7ee9b97d5a9c82f859d5623
z3064ae6bdc8553d95508d8f99e4ddaf2aa65380f13d6441903a539a11e81e30e91e9f8814c522e
zf9e9c53fb18dfe63fe4b5e06440ecb0dc9be72d1ebaa8bfd2f61c9fa97284f2434d677baa20206
z0afec9f0511f955dbc8b526757c71819d808f89808058d706756237dfcef5bca902d1365f5f61e
zbbe0a88e7f3bcb3eb162a7e1bdafd2a51a1e924b06214915685275d63032c2f45f444879494426
zc531341c0b5eceaef819f5e0eb51890cf1e46be4f34f4e6e1d79918bce36a6ef35f44cc42d5704
ze428ed912ba1236b8b271a30c0c62ffe129fa2748c963acb668214b5cbe610fc828b2b7adb1a49
z0dd1cd5529c1228e0ea679a34899e75f853c868f871c2e17a01edfd3d52dab695b6942d8076f70
z9c956a395222950c9926de5c016552f85d258cc794cdfcb8fd65e92c91cd8eae471d35ffe683e9
z7aa8dffa507c68775071689bb198dc5ae3ee9c4841db35f5bfcbfdb37bdf8e06b484f01609aedf
z5c7023b0bf032842ecfd8db8b22ddeaf75b4f2b88ec433ace1d324f5fbfa81708acb74fea90a01
z4e01290723c47cff7af25fb3e34782f645776556294dd8a577bf4abcd01c58acb2687ddad6ab2a
zdd53eb4e823b42bc5e2b5d89d2f4deedd47fa9d2548d9a72fb3aff8ca26c920e6bcf5b31bc67ff
z7845f22510ad734785f81a4675bf79a64bf49ae5285506152ee749f860ca55f34835d38ccb62d4
zd8688e734f352d113fcf154d2807f02e112b03585adbee7a814353a6d8c98069eb84171d75e177
z534ba765d8238703c3fc5cf5f9951adf6adc330b9653c0e3dbceab9964ef1a6a201fbdb42322f5
z391c205dd17ce8debdde7d7b8ca083dd01fdad4355b25799f5e4f3d591bd47794365c410282b73
z37c35a107ba9fff8721fea2bc4d11024a1fb4574d632eccfb8bf2377682a06c49883cee787b0a7
zf702fe66704e61a50e0bb5fa0eef89f4521db0e8e2ddf43a5f08d8162a639aff81548ef32c92fc
z58e42c6fc37a50b27e9a91f176f6e4da9b7725ea0916d74afa3cbe9ff96bfc821f81873ab93068
z596112cc983a05103712ba7d7471a838e6782766c35e5cf3fa741a97983bc0b3be0f70ff22eb72
z9549176be1329114b109f4fb6cdee61c9fb34016f13652c03d84a80e6f3c8e4727182239b3e56d
z1b8003af644bfeedd5ad28daaca0505675375903b2df1936947298cd85b667ba5ac5acee6131f9
z7bfc9f4bbd14ec5bd90c62f6bc3533ea844c748e4272689a7a1a81c686c4e2ed2bc6be0b1b3323
z0693f98a39bb31f45efc6a46a0469ee9e098389f0fc1a39e8bdf18898fb911ff97dc725f194f53
zd15fbc85ba83ec628ff40791bf481edee84fc60865b62d569cf858984ad26fed9f28436774ba4a
z37811dcfece7d27cc894385fadb1dc5d85744f48ba93be9d70c4808016c3c7cd68f27bac6162a9
z45468670cf61e39b6311934f9f4440e02ac26e3ab3e1e7a8181cd7305d64be141588d95994bd64
zdfb40041685c68ac102532cc889d3b1ae9f0bdc7de6841cb35b5dca624bd33ce0d02f85fb317d2
z6491fd4754d87639173c006bca288d9683f7207a9b0ca17b5f561cf08b825369e49f5d67514591
z6016a6302227e42e816403b2d0f7f3b796b032dd6856d9bb48b622a505f427eda23c4b7d87d10b
z24fa4061af05609be223e307dbd5beed7091a5c45174fdaf30a092580b37829b32bd5cfd3417e5
z47f055e745fd34f67a8d298244f47e671a0baec2440e8f1b8bfd674dfd76d795f9af458c4b62af
z7bc9100a31fb3f436e39bfc5a080b539f4967cc9c27fdd559d8ea26444c5353f794ff6b8cdc1a4
z80d8a523c7dad9fe5ff36dd64bfb6293a57e74f9ed7e95cb080612b9ca7bf9681fe5505f5de7bc
z9b2d36d087711b5ed88c860ee8269134317d4d736584e9fbe7a9d52e007ddb815c0e9ddeef98e7
z2682923ba23cc0144edc030b3055c470ee9f45b866b1d5dec17e84d291b42a254ff45d1c12bd9e
z6dcbd52d95e15fff1516c6eda58b7d056cd409c0400fbd112aaa222af0b0d8fde8a3fd4c9914b4
z992b29c22ca3198b6d7d93971dbd748dca642b298c50a37190540dd560f40f53c2a6176704fd6f
zb3a2c976476bee479a0b386b7676410d15b7401acee21569d256429049c0fb65d6146d54b4a066
za43aa474f6daa7ddcbc0cf3dd584441f23fc452154d75d173689d58354fae713586c6e1a8b2e83
z16db3a8be134441fd9ccf810f9ad443f6577dbd4606f504f0eb16dfd78f564a76105174aaabc81
z93f04b09f2cc0ff2dbbe3a8c64169d6870ef84f74fa34605045986de74562d040bc75d031a02f5
zb146df35f85df4fba40df8342094ce92f3901fb6115f55adda1490a60c3686472e67a9d7834fb3
zc83dcf69391fa3bfd13374c6fd4ab3c8c928282c8c89dd1d9842ab4a2299fa1ba4d38ba71a22b6
zf8b971e8960ece1012b03c285d08d824e73611c6e7dcf002e8281758e6730491845358138250ef
z00404518bfed910aa85598de39824e7e5fe5b23f4c1ad730b922103ade594f2115a8dc00bef6b9
zd7b20907a79be1341f8dc7345e6ec52f52542df15220ee3845ea09b966ea4e7ae802561247fae9
zaea56164a334d5793f6923d79c49965ac0baea0b1287b36a446f5b7f5d8975b92f8a5f570bdb13
z2cd62fa14f1bf6a23aa48e5be4bffa7146b3b7c45430ca91b1042ef4670175658c824b8f611a52
z69236aa342ff509b4ae40456411336a7fb38436a2baedb9fd6a6d857386d893d7e0013504efd1c
z622be0383b3925e9d5eb793959227705be6cd8bead3797da71c125920c567761312e4f2d6b372b
z9e1ea5e9bc2bf8f8fea070a5f8fb9dd37b27a24624868f69324e1c305655472cd1f221fee8a6bf
z0bd73ef46bc2aae583cbe971b4c8f47f7322cca8786e6ce8c097c549f0858e06dcaacd0f5c7191
z61a01138e2f403c41048d8c5b75f3dc389f3ee913a81ee0a87b785fcedde65f936461904f946ce
z94983555d04a72ea44b6dc149d93d48221a210ddc5d71607bd1788b6e29cdcbcd6c07222619019
z65a78a89c765ac13e51f5ebda3b11550c6b5a6f994393082c96f0e804f1e70cc77cf2dfb57fc8a
z1e44889abb2762ca9effcd889c10d1f62f323ccc8cbfbf7d9499df997ca1f2e2a9c51882dd101b
z0c1372641bd68e976b0ba5e72e32df81e6d70bfa72137cccabc186352b1adf4c86baa30a362a7d
z6896208fcc5dfadfc31d9e717ddd2a032fd641f0c0febf7fc665be278252fd94eb84c556e54435
ze1d5949ed254af3f24dcf3e1496a39ac1e131dd3cfa311e64ce40fb20550e11592edbd84cc7ebb
zf30acdce473c41f1665f494ca2027716d1177be775215eb1c48c1dc4547af511648e1fe70582c8
z92c26aa68649f50b796e4cc4a9c9279bf5f91344b60bb15a8b5b821c10f1d8f49272a17a2e7c7f
z4b39d6871fd21a7a267a5b7754795df0f20aaa22398d4327763dad181d042a4adf557a5b33a956
z488855bb74bdf19f26c2fdd73787e9fb899f556e2514e3a5c50487ec210551ccd03b415252470d
z7d31fc8720423ecff4ab07ffc6f972dda5034215a6d67e1ff7ac7650b066fb506a67bcbc5e4054
zdf3fc02a9136c8045ceb5627986ea5c583f0ef19fa0cb4b218f10c1a74c34f7d6daab3500fa91a
z854c9b3bfe7e12d47ae0a4dfd1a15ec8a7e02fb57481ed05f34360cba612a22f3d96880b8a9779
ze880aa6f6b111f4df8c791f159a884a0fe14535f39fed95ec66dce98c5dda4543b75a5dca43932
z3ccf07996b3ebda7789dac5154c985687b52d06cc30b0e6f99cf94eb6f5cf3b297d5e115a538ba
zac58822de480efbbd3ff806558728907347338bc18dab0911cc87b5c4d2f80313c6fdb909a844e
z2d268115fe67ff958c881117fd0e14d872c983b4e482c392915ebed1857eaae0dc6c594f1d0d5a
z40b9d20118e3cd527955551c86a652f0929e1e7cb4228de47fba5f5eadb38f3ab7511a83af5b7e
z2580e1185f86b1f7cb8993e4fcea4ba35d735a78e14e69b0dfc0c67da95d6cc6b6c072b61e8826
zf35e24da8107d789ae096c45b0c1fe0f9c87290e4f8edf70efb424f6419f92259fa35758bfde2d
z5bc16f2235b02ad015f8998153e8606a0897b4d5ea51478f32886b6701983121c10ccf5fcbd0d1
z35aaebcfc082e33f60699d3e7ceca92b352276040481a454d7a4a56c1eb1c08a7ee2da2566b5eb
z6f867a25196186feb6a09b4e591c5f99b736c0dcbf3652184fe09b07748b96beba26b8339ba9a5
z224db60ab12cbef41e0c3481dd864acc5669ccbc1fe7f38d157ef0635810422d898ad47253afd0
z6643013943f747d03074c18cdb2e2b1e6908b1065ed9d822b52bc140037b8783065a579dec86f7
z39348a36e2825832c19060eac0da8ab1a4e896f595f2227d5084842c9b7ec7846750433c571379
z216638b8a42bec6b7f66eaaa0308b958f4be7d85434eceb363ec596de29427c584efaf212e5c29
z64c53a44e334c34f922b27513b784f864ac53d51b551c436d4bbd2ba97d6bc53be78e95591d847
z8a6bb9fd090484f9e47afe153ef0532a44cff43f7b5a922f1b8e78f31304e419e6cbce16cfadf5
z1f78be34aa9a4a42d0255999b6eb68987034fb2ac8941382f0b64385ce0822c8a6de4fa9fe4c4a
zf3f9aac812022317617eeafe2bf3dc951d778018be8bffb9f560e77de7722b1d6aeb91043228c3
z7f253cfd4fcf4fa25122265e7c38c1be6ce9cc452571a7a1897b73d6594061e7a5114162099037
zcbaa9825026b0b0100594e7f88613db5efe2aedbbbd158e038bd3411fd56be6645a12e3c055e6b
z1529179c01b1ea2aa16f2616f6285c4d49d67ac7a76a2e1325338974591b1718dad7d4daa6d174
z92de84a5466c7999ae3edca66f9d875abab3dd6fc87433fe94e86e8ca89085d1fa99eb1e1c7710
z041fe157d5956e5221ab5df01e1977d8b161d3bc8b50703bbb9338c3ff75267586df5fe29d89bd
zbd6ca1663c9c8e5d585d9055d95b360669fdc8fc441bee0c9f8c5f094265ea3fc536c413885af0
zeefb66b3e0a9084c338b29a1da2081841ab6b2a9a6ea9f69de4723ac85e1757e753c4328c71304
zf7f6391577bb307deb02bbd8d7ac795981b06a9d2f6005e76e12286fde292a0550ad2f66382f6a
zf96f028794a2e72c83068e64793cfab2676fe23d03fc528467a1bacd4890da78aa070bf3c7a360
z7b583f30f73033f585b90db20caf61b296265877f8b1e539b3f58ed6fe52991eae878f7c0da8f8
z2a669fc7892254e6c48a53e3480b527a9b919ba6487ad5da5f140271d049cda9d793c1e06b7534
z5c4413f7e8d4dde13bfb667aa4a724733635d8cafb848e1a14dc80ce0f5e2149f1f91d42d5d863
z0906a693de59b06d6cf04baddc8aa5836fd9108b56f5f5986fda47edb1deaabe33b860145b4614
z51a1fa42c182d43a6b1d8f2934358fed5cd7c08379935502f96ffd7ebdad89cae2cd065786a274
zce74a4cf00454bf41ae3fb5aa3f32717057c8b4af3e3e47318969f698f4d44a8c0eef2623196bd
zafa69dcc6de54131b90c176de13ffcd2ca704e8ca7c1f3a964b8d3599a9d60f7bed94712d6b2a8
z506c146fbdf18cdfed571c8a86748bb5f4e3f5d97213623692447e292522b8c49abefa09fd5112
z0988a1ec8b82f8702a4a2c11277c9f8cd745df69eb12f8c79b8526a45dcfe5ae8faaaef8855e12
z8365ed50e2c61bc20615c571daa7b9553adc2e3ffb692780b42640273f459f07c2964088a667ca
z3c981b709babb90364d3a21334625d9a712e49de5f4c731648ce4763cb7dee00b32ff7ef5810f4
z87f8862010f64f86f35626638825774c56f8c8f5539d866e10904490cd6ed65f9cfb231b6dc3d3
z5bf686379b6fbbbdf5000ec586f8b06c3392dd7769e08eb21a5062d6990e3c1e630f95b054c054
z117b7cf50136aca8f1058c5f7b54ae89af7e0abf1512b4f054d1a975741b3789462f3823b842ee
z8145846460d19a858d883c17b80070e01dd8c9f7027b865545f56095e4926b4ca616150611663e
zecd82bace2e8eed876440d5cf462c42ddff36a9a4e187634961d9620afe235a06891ae92d81040
z513e60fc7f10a7e313110c05594ee3c1941835311c7a2c7dffc09abcd6fd8cd04734caad143639
z7455db9e9e0d2397a9ac359ce71e6f5ae888d4c72315c95a826ee9533c8c9ae84f0daf0e9fc509
z42ebdf64c7a9fcea096a575c6e717e41b113e6d1e1d6a8ba52bf64e0b53f62c8a78354a3294881
z22ff1da3dc4fe7fbb9e17f00ac78c762bb81ea0162cd9ee5ac84fe493fe5f37010078c1069980b
za96821e99b4a4c7b731c82590afd9be45725ca62fb332f89b156c3bffa79570e045b8982bbfe16
zaedbd7e5673a85e85b4181773d627b73dacee2ec4b1c1f6935094d0f0d4b3d8b3affe34fa1c28f
z0a6faf5e7fcf5dbf876feb3fa379ba2926147eaf3c8d1f61179334aa45e0574038f1748aadc2c6
zd357eb7f3e60df53a7f0189cfc759226624437c0be349362b9eca8c839bda087c76ee7c71edeca
z78e347aa8812317222a693cf506068fa6e25470a4408ec8c000ed602602469c41d33d76c39a382
ze14ccb0156659760fc246a0165560c95bff633d9ebd812d7317b074717f4093ee72aa45284431e
z379b2a45fd766362343703ae2b0f5b6763938c5b14f29e6a066c69527c4a01adf4ce209ceccda2
z106442d52d4483de3e7210ff553e46a10f25596d96db0d7887061e8ee7c8ea90c26cce81628fb4
z2c9a2389c3e7c4fcdc135aed22bd2cfbff83550d394400fcfdc50de18160edc28a453e05fe11ea
zb3c999adc99d23a332625848d3143ecf6698f0e25f566b2748bdacb23bce64f47fdd711e4753fe
z1d66774139749c73b276eebbbf3039e79d42f482dbd47c06de43ee4fea3f6853287bb9869d48a5
zc6004566cc9bea61e61fd4c01402ac0ca440acd6b0014f302a00a69c9dc43732e4b0107157ffd7
zca891890f01cb05576b184ea0dbbf4a5c1f7be55df9da328b1a3b7a893101cd265a98712bb1ef7
z33611ded09ea331055d44e708a654a59ba728020d62bb63e2e4d031b2458b41e3c3fbba1517b2a
z778e03ca9777827572a44d2ea168e0d7c4cae13ed11f8fdd47dca2113539150f22c0708796dde9
zc067cf6fe7d3792509260b72b61a6dcd3756a32b64fb184d0e0ad0a9564940e7d69204ab91ed1a
z6ecd799cffc66c345c2bb9caccc5783f15d93c99ab3ba57a95bcb5a56e23709adb82d5e2dacd81
z81e9fc0d340b32e9fe27989671fdda1840c6a07d4ef864963bbd4d2f3d000c96876b09bec5d91a
z0802e18398065354d9730331b9dabac8bb90987391088d63dc79e678b716fd5aa53b9e09d0e7fd
z0470811ac6bfdfce4371a32b23f4d6f74a8f0525ad8f2e73bd982569d3c80c46bed4f4371fae67
zb864182985b7ab99debd0ec221c129b4d661ed14ed229ca6b8729bb366b3c997c1e8f692d41aa2
z368419e1d13adcaa2a61108a2d668d7c7bc8a5585f9533c6042dd8b57917cd20fdd612c193aa57
z4acf39b9c00af7823d712da19ecc57be120277117ae38d2d6128e96138b6195767a4bbb87c8b5d
zef8f3eee0345bf5c58b749984f02381d4ad6e101f1c388ff0f9a5b52a1c4f24d10e7a69216b297
z9b843bf333aaaed956ec9b32c090c12d85cadd1845149e9150fab42817cae49eaaacbf716b9db5
z9c7da2efd1718b5a877ee52422d210250969126defc6369aa391ef2c251ebcd69747a71a996292
zf1d188ce9b893d7b6e0ee5df0ecf228aa8cbf019e42112350f75b7475178584a90f51060a41a81
z84dd91f37704dc114bf30cd62129a134e0d46ea6b33a8e7bb3d1a1bb2273dd620b7502eed05f3f
z65711e13745fdbe86b9e71c5080ef5e85e7e5c103ec6ee7090950326252d742bc7cc295f4d80f0
z8d36781991ad10631a89ad0e8d948f727527edad3fe8a885a8404a0d3f67c32185b7286ced960c
ze371afd06d561226d88ebdd8e2ab78b76fb3411fc87da8f72dc61e03ba38251bec94ef2846a679
z8ffaf310acf60bfa0a6e4a519b83b8935dd535c06e9c5058bf83ddb3c1d00c04cec2fbff10814e
zb97d20e17bfe63c6c91ff26ac07611277d5e8a846a0ad3b5ecc1ae5c234605c164bd72e54bf435
za439daee0ac010efbae824b146f4426f8da921a77d30ee2a957c9fa3056a0e3661895e6ebb3de6
ze14cec02bc247737b8a6cbbb0193df7e9aae7e184bf6bde595aeee3083e7c849b660474519027a
z6bdbc943cc45617da428aa04fbd1993cbc4532cedead9c1a2d5bb11be6738bdc8e43c5e56a6a00
z5817be3080a77e1336f3b27b4c67f36057893b5998ec611c4828b37d8d916d1c37be139a8a3218
zc1591536e9c661ce13473eeb60d3757cdbfe7c3d9d89c64c4f04832db3d9c427a4f9897db5e120
z46c9e12929f424d39f383b9bcc191f8c10ec9f019cb4fcabded1eea85342ef53152efe85ae5d5b
za7e3fdb22c06753a680d5976c226348cffbbc937a3761c09249275a6a6c5ac39fb3915019df239
z48c1830f41c1baa5cc7d05b184cdbad3afb085e156384bd9c80e9f33e76b9a53e65a83d0ed5a48
z080fcd9e69ba28fcce4dd823aaaa80bdc018d7e1829ede901e65dcee646225feab6c5b245d73e0
z561e3303cce2ee0fcc01bb03d35ea7145d2fcbf0c16fefd37e0a136476ad26fbbe3fb812a304fc
ze7b769f9680a764a5d5178e977c6dcba8299324a751e7e27bae222db15b2488748a971d2026e04
z56d83cb225b7c45f29ae8dcb3c42a4bf2bbc61be8dbcd76ceb1970746f42cf5f9d2fdca22a10da
z80cfd2b2a2496d598a55f153d063775609a70e87588da7beb5364b9c7399be94626511e563fa83
zbb0853329dc68f30dff27047a6378b555ad80ed820af25da84ed705e611f1789d3389dc5bfb204
z30dfb2416cb25e6225d1e1de84d41d85965cdc09855bb318df12ec34c26aab313707efc6f12aca
z1d20ef2c2a37f530d3c31d01661a53588bff70067c65cfc8fc8b1bc2eeecd27aaa91a487e017fc
z94227eaff0bb7bd67bf39c0edbd149a68b703d5110deeb7c54cce0e82f722a89fcb3e506fd896c
z9d641d432e4c28412eec57ac8dd839620d6d0f13275053145226ee879ab5328683d98ffc358278
z7fa60f3a730c7a51a6956477d162f5e20de6046187c20422a4a2cbfebc3cfe4a3d2cac21127db8
z69b93a5ea24890865e846eb4353e435819b521df4c7cf1441ba19c13cb37431a9284e0bde3f658
z549f752f67146d30a4745f211042e550396af57d3afcddcdb62097ad32b69b7d59932c4243f87a
z575934c05145e6b9962f59e9c845ace44c92552097517f595b3437ecad3d2eb428e99fc429727f
zd6b12bc5e1a60601002bdd7febb28c2864bad4265ec910b60592fd52c92a1040f5e07169fe71ff
zbaa174915e5948d1b1c8d5c6563adc49737c83c1709941f5db39b604fc4935bfaab7c03f4e326c
z09d0f0aaca31b34698edc9e92d3be392c68022226b9192730058cfeb167b0cea2702c9a668f9c8
z8e0488b8263b386024fd59174bd727677d30bf860a3b9fa2a2b6500174a1dccfdd23a7ade9e8e7
zea12b9f9608fa76f4e4848f2708987bc966eedfdaa528f31f422c1178685cb25b1dc04a7c1733b
z99ee2e014831612a3800fa190c1bab71f92d1227cd24ab2c4905e8efb84427b5fd4f1cd8076df1
z05247cec170591297394666b86e9a8df4544f420c0e5f4f54de26c6081d5d62c2464d5dbc03f08
zd80769189ee615fd66ac02375b6b69ff8f5fe4818d6998fde16555fd8644c0d0d570f05b77126f
zca2ab5226b81ae76be31afe49d8f5eca5927caa49f7f7d79311684b427ba4cee0490004a2f200e
z881ce32653ba56cb40d77272160fbc085df869e62f4f280b85c805d6750fdbebc0ac58cf0a18a9
za28bd423621496dc8f4b970ba11bd48ab3b4e460195f0c13f8e26584180f86172651822752abb4
z3867fdd3edb333a0e05845cf9b4d69e23de7818f6baf77bd6c93f227bbdeabe145fb904d1ca931
z58e91545302b52c49cbbaba442a76190d3a83641c843f08959240e681bf41caa2f9e27917f900c
za557bcdbbe6ac40b4259708effcda577a920f0f6681f3d314639cd620d0a455e9fa2af029aad45
zde7f214acb06bc3c14312ded438352a334b3917855640773c47d9f056f5c0ceb7ba147431d7a9c
ze1d6daaf6fedcc01391696eb5b22fba0e97604b08449d305634bbc3d38752d994f28cf867a9d71
z156c587d379eb62079010722b43eaca48520aea3793f7adbdb6f4a3a54b7c073b0d86a14f59556
z1f50d7a2cc866be38df4550f2e52f760bb0058378ca4b575fa6b379bc2f571188352b8067892bf
z7fdfa25c4f42b38d21d78e99325c4a04047df13d4413777d43ae93710bceb50f035f6b6ba0f8eb
zb63e9945a2a35c80c3ef5d1127cd77d74ce6e20bc2c5255e8c70b116baee6f6b9694454f72ee01
z9de1d8521f82cbf598f633cd7fad44436ef10ffe3a89ca70adc9529bfb572ef1e9573d9ea13cfc
z8f77f092e106dbdb0d9d52f3bc9c7e9a4cdc4e7ddde720b55f97b418e9b368ffa7af99d2ce8708
zc3f597e1b61e9500788aff254e89ce4dead87afcac5033b84fa894db7f4d3c0159cc8a7fb79d0d
zd6178d4a1955be9cec7035861f5c227ac933a1d708b3fab53761931252697e58e379b2d6b35933
z4b437559c6a0c2170a3ab07bce23edad9afac71f082b030275f6ca8bc23b4387984f9e524f8f71
z950c92f14678c27c7473ba979634936666931bde0cde1cdf4458b6026e8cfaebb2a0c76a4f5886
z230c95365e13360fd4cf986336ccf98a124e2a19468da59a0573f62048d4089ff7b5f0772c5b94
za97030414af088f7f09117e0fc9fa918fc8b8f418e7d9e8600605f3dce697074853bf454f01a35
z8fd597f5612fdb1f13bf98b66306b9e2792c307ba6a868efc23384f3e103ddcd4bc1a2574c704b
zcb304a712c621f1813a6c37f75755dbd73686a88ad37e2b72be72dca181b6d3dd6a460955dd1d3
zc22b6884d3d3a63cb3116b61623e5402fcbe268bf9b43406d3c6e43d69559117bdc11dde983035
z1f38570020dc41dbbeca774543f0a5c58fc7cf0e74726c2c3327c3b094bddea38ed399896871e5
zecaf1780c82ff620124414557979dd2e151f04f824fdf4e32c9e6a3ce774c76db857a115008ecd
zf82ddcee3e249845209ac54cc0726420b227eaa5128a85dfed8323fb266eebb2cf47e0c96e4955
zb5bd8fddec9ca5d5d12ab17a46d78238f3d04892314a790144a3452fae00f09ff5fbaf4f5b368d
z3f7f62955f409060c1f67c70f476200db1885568c9154ced7d6e5edc7362b80dd8df43d169fbd1
z6325e89e720993d6df5e4ccc1ddb2cc50334d5ee4f8c6ae9d0dc8521434b8423b2be763e69f169
z6436d6408b9fbae3d9dc568aa56163b48b77266efe49576e92a252d8f8acd016aa41cbef3e8fab
z3689117f3707a10ce4e3a0b786a8f880dcf51305e1bc527dd7f38d4143486da5978473f4ec0361
z5fd9feb2adebdfc11f1f7cfaa3c838c88dd06e9b94912096e4a4f6b9c9ecbf5de854926c5ace2c
z489b715a20128b4983998ebc07a78d2909286841db6589dcaf32588f096e53f4654e4833baac89
za6ef1068248d72c30c896887be1169f280245868ef9203b2022aa21335bf89d8f2bef95448866c
z7b977bed8d075e8db689bbaff878c8f583daf9cc37235799e3b8180b04545fab35bf6c0b76a4df
z6021376b165599e64a041357f4d7412472023d4c0b4a8d083ef6ec5574031ec6e8c276fe65009b
z2d9b0658b39d1b044106065b6e926d12328bdd94b4e877aefea83c496902cc87fd6f9b3028561d
z07f5d6a87d84f620b95b0ef436aed3ad697cccff4de512a9aee72f603ac2ec502e5878d8cac51b
zc6328247e0c88d6b1991cc3aa50c52670eb6b139fe8d2541c1f636eb5d2dace1339c1b0f784b21
zaaee87834d2be137635ca38a89e0f21df7f1b159b59b97fad7eafdd4e3acae86e9fb583f422aac
z3ea6c4a486874f174390b185b7fee31c7a8056781cb2ed50b2e2b1b5e3d74638e04520611c8d43
z70a5bb0bf177ca506a8258c87ae067ffa3fc8ab73808e5c2d7528bc058588390004b072a1ab8c8
z7c605918b92a6f320745f68c4e2b5ea053ddb2e72d8350e2dec78b9b1312183d4d8e259d8c98d5
z617df96356dd1fe42e158ff86c1e6af84b247db72d5a372f65bd8829bb50bd40d771c46d9c34c7
z80d55f2c36dd1c2d25304a2693916981be91184380824c5e66ab65436e60701425a61d63d15568
z0a73d8291fc2fd4b47bceff48496b2f39c3fd3b6c2ca8127d6ca57801441c0693c211c53d68db7
zda0c38d2dc483ea979499618dda81ad625f3839e1357bafd0c567fb6c877cdde1554361fd1f34d
z922701b08abf2e7a261db9e124d59f08c74cd7fee4c41a5dec1f87576c9e51fae6eb91ce736743
z43cb64206729a5e4d0f44a86f48e8865cf5180a74debf7094d36dc4179fbab8d6cd20463ebc8c3
zfa49b4d9c9d7b75389709594841ce542626555aa4412e2d4d9acb14d79336b5121b2f258c9aeeb
z1d54fa927c40f2381848abd99e8a3b6d656153c92ffc2fcd06bddd42cd836abd9ca4159fe5725d
z08682fb4dee6cce87e5eb513b1b3cc20c229ac7c3e89d482f55632a7cea015a997589f89dc0ccc
z4f27d00234492fb427368827f8e949f68ae90446407ac70ed7e950fe7d21036a3166b372897579
z6811b5580f8fa88eb1f7f130635d43effb2e210204dfb5a2e034048f2670ae62b3b35b83f55545
z44f2858b06c439b812b82a7ab1eba4106f1915615a3df7c12bbdfb5ce104018713e10beac14a7c
zc8c5c356b2159433640f429364b7425cda28a3c54d88aba31959266cae98c66b8fbd8b44192ae5
z94a2f243b73c2a59e9178fb479949b1189f16863a327b0470ed907d26b1ff0acb8dda1b01cbd18
z082f7e96d3495a5b024d57e5e9c63a5c229a5da96333b785e75f168f5fb4c3be3e2703a4ade90e
z404c9074ab6536b043ccaf4e5333f663a5bb03796703487e6eb1c2ee6e290ea2370ca060442974
z012dcfac85f4d3dff419df29d7850e3927588e15f04b2f3f93747051a15a593f5676480fafb97f
z8371496c416b5fcaf44a9abefcbd3a5b1914a2ead5eb57fe032dc556534ec9a3a3f64d3482c37d
ze7e5b675da78ea76a11a384b879dae13dc2d1cea83b718084f6469ba4f8dd5cc006e0c9179fd1b
zaf896520f1bb1dd50cc3562a8476a9aaba59a9e976a0aa12193f755680181142b6be4aed969437
z19cbff5f2e5b1da9b37087c33c52616b7933deeeca8e0f5731819091b4583b075f0a03c050b092
z9ca5db42c1647098f5463d119eff36e5b0809689ee97aa43dd3c27731a8ca76389c159651ef1df
z799ef009157ed44a0eda9abc8c29bce4775e32a6970405ff0316f1aaeb79e5a05aa2f7724035e7
zc4eaca9768b75f100e1fc28cb8b6af0e3addbd824834907a4457dc900885510943eae89a527b4b
z906f0ed2c6eadc91ac897bd5dc35c3947d6c747028459b0b77176265ee3edc482e6753bcdcdc2d
zce6d5e37ab9f66be82a8beffa1fa0a78ee48128488d4454a2168822d03f07b4a2f5dce84ee40f1
z95b479aead82ef9f45b70468b3f8b39cd350695cfe58c7c8c0403f199bcc883770830b35f6ad33
zde5b0f4ab067ad709bf4abbbf263a6a8d42e3a5c098732f667ee3d136781930ac7a203202efa90
z8a5ab56da1e22bd79e2176d911c669e36d209f4bc2d71d433a897946042525c8498610bd0f2ca3
zca26bc2a88a9acc9d78ddc9244a966a44f62a2f2876f3742534d94506b8d8fd3feeb27c01c9961
z2d4c03371fd75b86de6763fe0585b37770f9e43ca0bbd62b6448ba1ff581f1be2af30b6acbd132
zbebad0d0a5e5da7685d0efcadb7fcf288bfbc15827c67f863f9fd1e4192b68ee083ff3dad876a8
ze6aae068c698d3030fe62378de095454d55b548d3397738e0b607e23f9c26b542858c6516b1b7b
z0149d4fb314b28fe8db9b8c322286b4b6997e52226315e6a24f1350225e1814043aed3541fca3a
z0d4f3a5b459227637f6d8c73557688d1e160fe9a5a62eccc6538b9fe83819a27e679d8ff91e0e7
z153f079dacf144f12e3fbc70aa78ca8b4f33c031fa043a03ea15c053c007a922deff184ae9a40a
zfb9066227ceda98e9d49ecd43c0743308ed80eab1197faef59c741faff54d63ed3dde75a0673b5
zd84cbc9f024ca59a9a4fbb04aa6b56724f280a5c59354eef242726899c022467b95f1cb6e8d053
z603f2b2164225f9c0eab53bb159e31e781106a00081374890dae47576b45a8f046239b9e17f823
z10877820c557d12f20e9bd105f4ad3d6ba265b96e4860e04e3628d387d827c2b3a7e7a5e435ab8
z76f9389a7cc54eec34ea3975b5f7176718b719a09283faf6dbc585f3171ce628933b85b53086fa
z6d06946fa67cd6920d8b5ea4d2db4bdbb28e28bf5e0f10d4fb6a79785b51d00336cb919b18153c
z5fe3bb2d33bf1320626e021d93c82b0a927cdd8f726eee1e643422da2abf4b0d9212b788f78650
z1f2809be3cf77c2e4b1009dff283b02a59ef512bd8c10c1cc5ff960417203a156350040fe8b351
z42bb681b39c9310b7b00b10c4d580e1a9cb92f2a9b6fb1340df12e0ab5d2fcdd9be4f0ec834a2b
z14f82ba3e377e4b18b0dfbf8026e4ecbf260601adabbc0cad4d4f96e49f52fd8522c83a67f4a9f
z9744c50e69f72dee05f475048352843baa4eae5b7ec67b48ea8bc8053192a1b113f555b3848b8b
z768c69861c489b441351ae2d0cce362b0b33d3b46e28cb1cc6069068e2bdf4536b12dac62cb735
zf10edb1269ce78183d5df16d59966d3e6ecf3c120793ba094bafb222e5a3af322eeea7039d98b6
zab250659c0e53b9ed53163eecad9eebbb62602d0c35bfc638e100e730c9e53262e5e590195f898
z3303118091d945a194289b892ef0a5478d8acb80e4aa6596e7e0b1d57225197a0339abc455dc66
za9f5fee2e0c84f6ed4db6a4536c5c32b8c873c026c7cb71f1ff22e8a732a227305281819594d0a
z1d8e3016344e35b4a05cfdb2fde422518f4b92f6f00b54c63b22877114f8c4784192e85b467c9e
zf3612c826793ed23a981afbc1306849d794bd05b85192cabe5b07b57378c8839e92d866c47e52c
zd70b2a7c0295ac061ae09dfbf95df9f3db1e382e8da0439855acedc45910c9b7c9e83d217249be
z02152f60794a5154aa0a49f4596514d072a157a878a65bd4a342fab69002cf639815f50fe98301
z38c624723798b3ba3f868e3e83d92d76a5c2a9821df9162ea8cf8c9416a133ca456c466de9acc7
z2e485751809e314f77368a60646d82af39efefe02b07f4fe9d98f19e02f26094443d4773c2912a
z93bac02cc0ed8a1ef5720c3b3fb0f8ea8f493f3217705fd3d44f0bae048c67935abad67bdb35e2
z38ca87e28a4c29f519787a2075cdefd7f5b6219b545a15e2cec2bb8c183dfbffb1fa2d3f6206a6
z89426bddc2fa3b86ae9f91f2ba8d5f004613b7c49790075a951e365af940fa5c4fa692bf4f113f
z5362e948ebe364195802db34d6cc3a04ccca110c9ef79588b76f7d9b2634d4bb6dcefb147077ef
z4d91f235e3145b1a48fe485c1bfe77c8c17891013bc6af1b69f0646358eed2b32145665e926cff
z827985953d29e4d5f045e37e128b4b5697f3203e4508f44cb302fd470c3f8adb6c4ee97869f08d
zfa763dc0bc89d50c25c8e4f2b266faf1fbc830e5565b611ae7ebfa9e9ec832e7277b4244ee8753
ze167bc8ea20aa7edcff9567d974071247ae152c1003827fa4465020740d94e3d3714ae398152d4
z680cf11920dc32cfad06d844cd5a66e1f32d0a7f5285f7fdc45cf0ce8d432c2a03fd1daf3a3b09
z50d6ef81f89900d7e583c55e994ad101e142c9214d8bc63d7c5a852dbd9dde6775bfce1bd405a8
z0581f3c3749b4cea21a9232197491d3da3377da374768817c59e5fa10082a5d63d17def57afb08
z3a9d86a8030c451832122f09faa6253280104b1e36906fb1835c3fc2b8c619534d55fda4ec1863
z74c17857fdbd0afa80d4dbf6f6edf5ca6658e8a6d56b550249a3eb649c22561f8c41c39a0cbdfa
z6733db7f29331f6d630677a1cb05b68ce5236e762ec63d0abfa8aec0fbbc9f761ed68a5ce2844a
zd005520231bc781133ec5790e7ffcab65f7a52195b49dcbf97ace1c35095ef9f223dfc2bd59a4d
z2d6aa4f1576df59f277b04cc68ed4df4208b51fcb76b7de3bab41e209c11f6f873b0c7878c8fff
z9d35587d13ed94d9cbdbebb608ea20206b7e4b53f19b14725980ff605f49720ad0782c82656b89
z7006c6420bf95c02c21606170c7cadee2b3e13d952b0b28e0a3d45a2ae27dc8e9591b625fe9f50
zf325bd7d81ec5acb9244da75c2c8357f8595c131c697322fe14d9ae3147ba24a7bd093f54bbbde
ze34ae6a75680ca35f9c498e67128894627cf83e420c2d7ac6d108b131d5c33fdaae543390d140f
zc95e7125afa06489b16ba07f5e5f683cbc966db4389d0a431678fc6ea8f8675e0c61e2c36c72a1
z6a516ce6ce3b672fb2751bc73fbf8ebe270a0ff0a7a70d1245c8433d333cd0dec7b6ff9a56098f
z9690928523dcf2233105f739204a7c8746f65ed53ea91689e4503127ef81bdba7dadcb4cc83a35
zefa51e0ad12744dfd5dda4af09b25cf2917fd475400d4b973fb6e7715434fced9b7f3e1cfc6da7
z18d9faeb67a7d1ef2ac287de84bb438d2ef2db19962a965e6b934130a314e77521f3adf718ce78
z451d7511b03174fe71a7c8eb8e7b2f43ba4e4bb150587f53aaa42bb4471fdf12dd75f5f976f53a
z078dd4d9481aacfd3fd32a2da2d8e9e5bf2d48464178222a6922195240c6c8ec3a2b6bda2b2bad
zd9d2cca7b0817969b617a45265c2b1d71100dc5f783a0e6b5790b13e902d844bf64182f6236b31
z34a3626a1d754cf8ebe98b9993ace0065f82e117e00814d1a6c6bccc5784e4e88cde84224af1b4
z0d78a8a9778fba01ccd64c1ecacecf2dcbf3fbba5394b1355dd88b8a6ae47412607e8a993a2d12
zdf8bec843f74547a8d4d10843ac633fec312e2eae0650404e041d56cf75f6a6c41c0d238d90829
zbd29bd31f3c256bf9c49a9372c2469f4476172a11d52510888f46a2e8b9395db4000ade1a7fcde
ze21137cd3710a2a93e87ae7f90cb3039cbd0fd6a7938d39c093fec6ae850d36cc9d83bf437db3c
zfed197d99ee238ebddbae8df914dbeb491ef07102ec2200da1276d8ececd71eb1cc4a69394ddcb
zb64ef06ec12ca6ba8a08d72014720b7f69ba3dbf2cadf357c93697857519e72fcfdb6e5ee92e2d
z067aa5ea1698c07b78d6b8296cf272a30e2a47317821a7319420b2f664394b19671018c44be1d0
z591164dc00034e5e4e2685d6017aa3ec866e8e9d5dd8c0317dc3c7e82c542db3b16524e9286791
z22767399f57e23d798c47d3043117c821a01674ff721ca96f151228fd6ba73503cdea00df5adb9
z7d45d41a385fb6be0306312930685dc3623e076fc41aa9433207d7f7b9065adbf7c7206d5197e0
z5a7adc505e44c1e7ad4b5241b18a0e040aa141bcc72d91db917b6f3065ba36d2d0e50d3ca51362
z54d32fd9ec95ee5fe19ff98214d3c06ee9eb8fdbb9ad7c87a7dfddd3741c7934ce793b1b6c3064
z26116771f9eabed8f59f2b2a2627232db80936f36224399554a2962f997eef485153056df84235
z594b11a292e7bafc88bbfd377f69abec56c2f5568ab15987c0c4063b56d85785609f6770816afb
ze63a065a6e3d07e7998cd30ba1880b5e7b132cb92c95cf0b32d8b90379e649cb24ff3b4463db8f
z1c5e7d265f65bf68cc2287f310e1493b054f4b6a73493c376c6a823d653966cafaba1b4af1b767
zb2d001c8ecb751a10fb0810c63b7cd0b7c119cdac42bd38597a66b0c7aa61da7dc6efdc0e5a8da
zf3adfeb57c3590ef55e96e6f1e17e1527f370a3505cf0f56191715d00e146b613f68bfbd649150
zb110066b96662556600af7d65263daa74ab3c90697d65179cf5b806b50bb2005ec227fdd3b3c8a
zc4619d19787fe97cf1d09e538a1d47beef402610f5b59c3c199cec6a71c3b3f2d29f17025426a1
z04385d458cf9d10f1f911f2ac9f51b9b399bd8c36c77806c9ddbc837c7127de84231b2378b3bcd
za02c6d7ca4a168f95fa6a9d039690ed8caf6fbdc06080da676ba3a334aa370352f664d66af34e4
z113eeb1841a588a791a00630952d73d9de9350927c31dd01961e1047672c8e7f8f1cd23023cde3
z0e5a1b610fe76c1cd9f6d5624ce6b92010473e5dbf6fa711eafbf0636c6016367d851079f983e5
z766b39001caec66df8ae7c9cfeb5f850264184bfab5faeb0530d2cd26c15c333621508492d5d65
z45654d37ea5b3915e2f31ad2851cec8fae4c942c959fb31891f35e0c8233a1e913538a7581cfd6
z2b15a7e71f1b043903b6d7db8f21271c094e3a93ad4f7a7ea7957417015942f71b3c9c91f94541
z9a229725f53baee3adedba65c5e5a85bdfebcaaefd53247fd00a033fc44f5e0580674b4e3b7d81
z173b15709c0f1004d8fe959d66cb1cb81c42d32accdf5964728ff987bd83b520aa40c26bbe4053
za6de2ab3d5f8d17095a41edb0d2b2d5225ef63c1d67b0206dc4a72af0dc985814e5b13d99c3dde
z7302f983faa1153bc9ec7f47fdb028ee6eecab074604417e88add17b206a19cb144a37fc7dbed1
ze941f806bd2fdc11881f1c7c53b6635df1332f11b4eb6b65cb027e5ee0aeedb55435be7a68069d
z2fac91db3ae269a6fc52510c725863a09faf7896185716a15eb8be3904b6559fde1130cba1358b
z0f6d172d14e5a26752029e32f650fb0d6015733e15ed4935ebd7ad944efe71e8029557ea9709ac
zdce8da12a4c1d3ca42f7ca673916584db4e7af08cf69a228f3da9f1a638fb48f6fec4d10fda85f
zf7d1ecd0e23eab6f4d45b82b3b612ca63a069eb59a4bc85af3ee7d1772d062757dead53bc5f8de
z52a51d1ed2507e0998c5d95776880a424bd044006e590a1ada982372ba417abc80e9978a5580c3
z6119788da9a35221d85f55fd30a1b0c203a56b1966b25f35803b96e7d1acc11df202991c38683b
zc5bedfff9d82036fc6d1e9924495669f89243a0599dac9ac8f56e970aa9ab1c0871772db1a6d3f
z7889baadfb016007074ac7c82961222c9e4528cdecfab0369c52bfa57ef97bedf38841240f2a64
zaffe57e674c675c2b6f3664d1a9c16fecc7133780467f7c6473e06114aec1985b6bc8adcea6b39
z42cc0428a68ca88350d4f399a37f23bb949b4a4a5790cb4f7b88566ff979d13d144d42feb524a9
zfbaa539c4d9031e63d50b6ef9d50f26859c31a404dadcde6b8acd143eec45b03e75b01b4904b6e
ze269c63aa21ce080b11effe66ec59a96bc840860a1fd39a8a1200a7066599c6bff99566127fff3
z1442ca1cf82cf85877f5456a71605f99ef78cfab05f9c920d63c10270e84f4e7db530f62be95fa
z02e666a718dfdfe217b1acda2a797bbf8ced39a0316d328d57b7bd1075b07932a773222f3cc57d
z1a5fe96ed5c61c04e84a3b3b50d9ca1f6607f26b4f3c24e4f7c96f7de1dab7e7db75e34a1d80e4
z7dde65b596e8bbf2100288bbceda2e6d3fc0dae4d78e04d659458076a753b6b06d67782401ae3f
ze9c559ba0d99e904fe66c9ec923024e7d23a9f2b8b01deef58a55d7ecb41dcdea38259d14efc40
z4c8bc77cb6eaeb909e2bcde2b6a32d6f168e04307d338bcc78c1c1694f7c85e6ce9528dd56819a
z884b9f45960c4c3de15a21c8e0edfbb27640265b62547bb7e4d2c7bb9274656055081acfdc2281
z8e0773ccfd546061a5d5cbca6c9d958fb359135c187a1df835f613b169a789173a87deb1a3d3d7
z7059ee317b37a3b9ae96c12e41ec78ffa433e4b42b9a2c54b9558cf6ca5dffc5b85b46232672a5
z6f2eee7643a460d38780290a2af70f1e67db6111639cb34442623864adf5d571f131e2f073a0d5
z5ce9206a5eca0b362e07b00fd63481d40c9178c7ec0580021990895622d2de19230a291af9dbc0
z00d4882d9eba3a324821f2ee4692e5d883190c2c2e78cac06d0a3f575b746e436f612ec4487467
z161d25b6487781b57b4683f0791b09affde5fadbbcbdced2e94948e1ef49e1d50dfae6aae2b9bf
za98b6b0045233f5d1522fe95ff2baa8a363742db1c4dfdeb8bcb15d5d0d2619f1d0029a8ce7485
z0c8ae88e430212f303adf115c5e2ece95a393bdfd34d7f5d9ffa2c722f1a8ff18ad7de14305f60
z949e1ad992d0be2989701d9cf779d4637ec48fb15ceae8f124a07b6fdbc312617c9d9a315f3e08
z1899292728fa4d17f872b80633d875c4df7ec6c9ba5890534b12a5d6181b4c4116052ca499f902
za0aead4a903c289a5dbfd2bd07079a9e39f815d3f37d96863faa12b44800cf7cf1ef13cbe5b2fa
zf1e201b012a60e701645df067b57081ec84aad0551821af6d944c29e2e8f5f1e6fda71f5724bb7
z81a7e03f95c544ef2536770e56e4696f262def3e4a6be9af73a94b59f8385aad729e50a1cb6eef
z3cde0664ca5f170d7de735bacc9bb856da888d6bed7ae167f2d72ec73f7db0ccd3a42e055b60e3
z60f360ba40ec65defb0af4deb49e37dd5364539e981d096e5a2f719ce531b82f84ad28fd34231f
z1b7757e6a4004cb7d04765a0d7d10b6f0796047e8802e69ac224419a9b02d87bda6290431e2420
z6dec7a7c0167b2806bbda6e55f0e1ad2c9190e976aaa25b0f571490e8f4100acb31e15db87e791
z804052a881e3a4ea9ce03915eba4c33158c7ba0c311e1ee321242613de3a408c390c92f20e4bd8
zb8c20c64d613a4aa2b4db1c5a70951db0c53e741a8a33c2653e36ed1d0869e86ce31a461e1a98b
z26526727db5747f1deacd572e14f9cd73ef611336d2fcc8087dd4cc24aaf364269405407c2ea42
z6f3f20283d8c3d33d8ed8fe2c4cfb7c5c404d4c7cd59fa51adf95352de3d938800be83a7709c98
z58f0a5ff21f342579a7e563e2ed7c74b1e7927cc8d1a829a2be1248a9e7ee575cd802d777eb844
zc5bce139835774fb4c1c2e6423fd772401e3bc0f8b7fdfc0e458bae099e4421bab2d3bcd987eba
z5992c9dec81178b63cdf9ab7e47ca775adeeaab6dbce1f710c2d8d277d6a8350ca50b88f29f26c
z563dbf61822e115d7ea4ca3dc2281dc75662f18b405cfade84a71f704ea6d81fad519b8b551f6a
z02fc26ea44df05720ccfd1a833abf536e108188c63164a1e0fa634d589aa01a271d291ebc3d345
z96e093205bf2180493d28bb82f96cbdd3ffdcf3d399c8dfdb6f05828b2d995b2e7c96902e151b9
z89f35bea4d38c34df9a7299a74dc102208b09471cf3ef55d247d1ad20e75ec3620169ecbce58ea
z743c686bbc9471931f2ac7ee8d6d6c299ddc2c1d65474df50b6d87522e94ffb56fe83a214e0925
za88482c2f10b1aeaa6683874834b52f7cb271b0fbb21c96dd40b53409ee2ecc5cb986f686f3766
zf44bc0f7dbf8a919189db84c90595dc250d84010e7daf5b1c525ed697bf2ae5ef01881b216036e
zcd4bd40f4da4e5429b757cf32e78916f3b0568389aef6bbef9e85b6f25c708b943889d20ad5cb6
zd876daa478c68f8f12db1ad1962ac9855c81f05e8e01aa669a5184b1d23548fdce0ced8e689998
z178f3982648a96e3180e6e208a965dc4fdd27bd862c3b01266bde8a14dc4a32189cc43027a6c65
zfb5d50fe47a577a8827994d7f628d6c4dd3d58cce18c7452b05ec588d457de425d75f0947464a4
z60531635c1832e6679aa1dde2ab9b913163fde8ec27d5c6a6acdc793628ef5c13d23f72d100313
z9a2499aca036f86d3237c336dc64fe7fa27ff483db69c92da2e427f4f1af79a42501c61c06f148
za027cba6b4bf33ff6d99f4dcac9a045b6186536db0d8ab39fd4a7d58d39307712539835034357b
za39dbb342c8d072162b85a443f6738681c6f089f7c3f41ba3fd5167332f548d4c9c79d5c65ca29
zed51bd9a531a33b2beea08e6bb0293bdf2e44e33449ef2004764ce4dd886ccd39596d31fd015be
z364d8477a2796c40ef24d3fd5af2bca030d77be4aabd9d89e0a235edaa29085560066306ae9c1a
zd14e6ca1f64f891bda46c392500d4539b2353c0d10c00f8eae4437f2ea6201b75e9c6e7ccc8912
z065e083eadcab57ee4ecd4fc45d35d459ec3579ae6186126e4ab07cf3941f3b53348ca0922b214
z90b6c5166926617173388ec2bc6900c52fd8b5f2571507b861a63fe58c20ec4ce8ff76be70c679
z406bbe92cfd138f0ec6065cc137e1111bf2282c55696bb33a36d03e721260457371c5b8eaef3a7
z29aeaffa10019dd8865e22bac9e9773c5aa865d3cbfb5385f2f93d040ce8c8521794cfc326cb5d
zc8f63860afc27601fbdf354714d4e06b51cbebf7bfb82f961005824793d4822d7f7a1bcbd922ae
z97eecf38b40ea13bdf723ba201b592ab513cf7f2abd2e630af56000def023342c0cd0da273275b
z150f9db0c8a15ff5514aa8d5cac94ca77d6894d44a1e568ca8e1f90a56f4b2076a9e9fa1d69296
zd967f059812d84546142ae1429d65d13bf6dce846282a957ababa23968201d160ff84a605f52fd
z93f0ef907ae5db1dec49aca8de6d912d17bcf1af2f2f2e67a18a56c7c2eb9e8fd54d79677ebbd4
zecea843ada134872c5458a40911adc930cd2528f3548edf7fbea380207f43a81e77ea75d60e103
za9f009b50b548fdf86337c615cb3b6ef59a3b8b2b9e33a277d1c71dc7c371be4fae14630fbaab7
z9eb85f96ad9b732e30abc91f545b2e6868036c8316e1132fe3c6cf3d13f525ce121f54e99ade85
z1a02c6a6fe876bf9a8dbdf899fa2c5ddff0bb52812e94e6ee60a1134e25e8900bf752a45f2d0b8
z34c30c057e0bcaa95d5b2435dccc1a46e2b4ee16a2e309a078243ad0413c8bddaaa898912b1664
z55f87fd8e4a9f5e0924c4f5071c6dcd5cf690d5c20f5969cc2248200bae866c5077e65c93457ea
zae302c54c726f93ac894ec6202a7fde8647fa97824f0b3ee20ea128594d21f3f84cc0fc03919eb
z36ef8f1983b270485c798edba3f86d7313d81c7540962f6a490b4f394ff6965ab375cfe2e23261
za025515f63957e132d6d83c38e1baa790a17880fce7be436388effe046cff2025d6407dfa9347c
zace21db7a54a3191d0350d5885f943c8ee8a169347b371cd34593352cda4c4170839374a668647
zffaa4e0774c143d5e0eaa0782cfa9b7ed8bd9f216a91c4098944a89669e533cfa8d92d374d6e90
z7c3033720cd95cc6e1934c63a35fa452047cbf9b7b1523fce71cbd1597da76560f0cfb4d5da8e6
z791fda24747304121ac7c81ffae8dfcca70ce343105d13285be5826ffd0641163d319b496db2a6
z4ba6f97057f0249e3cd15216b757b03fc0404f45aef93f265c046f4f5f8a59380181f435edbafd
z914f3753462efbbb67ebce42907f80b502ec1b72c8327cb16ca5d946a6d62e35d2b062206198ac
zae3c8a4095b5b6739b4c0087f725f2ae10b093863fd4b0e5381f752774da48913d9ad3a26d3e78
z677db2d2e934c81dbf1ca1cd8b3368765a237eb0dd7a4331e244e9828048d708acd8e938f4ae56
z7eeac44672fe4a6fac137fa58a73e53033c7b88f26c0e3a9ce02a771c83358cb7e849140c1e884
z727d77d30748b032c49f194c920d87687b9dbdb50e259b1b314b6aba2b7eb56e468440ea43c07e
z7e61e054714343130cdafb5a3743b298434acfc1f14d0c59bfc576bbba9873f671255b5686d66e
z0b6c995cb8bfbd54102153b80ed2b9f58e867e4884427703fd0c365f413d593348cd604eaaa878
z9962a4ef0fd53e5e6931e00f389447a5276e388f7601297fed94e00aa3210fe81ac79bbb3694c9
z23e6aac7a1219bd0de7c74cd7cf6a4b0e11a6921de6f5e1967ddc964a7801c70b7fe7fa80dd0a8
zaea20f60c24379eaa4833ea6d5df4b25d24c31e1aaef828f56dc110cea15f47327096cd7731474
zcde069d62f646eed52e48fdd8e56d8e2d6a2df62228959ea6b610a71ae3cbb5ccdcb321bfdbcf7
za00d974a35cf54f5ce9dbe6be71b96f4cacc7aed17427dd60318f359abc47083d15cbc6694a613
zb9109646c641950cfedb6b803c53bf57081695450f228eb019b709dfa2046e9db68d307314cd5b
zf35027fc4312e31318a2404e20af381432a578db3be2a7f7ad579c30eb6a1c73ef19404e96ff55
zc061e5cee8d45ddad0f50ede10bb03ea62a1d09720b5f1e32e50eabcab40f8c05617c529bdb3f6
z4b73edcf978d1c9f7f0dddb970042ec424c15b3ab704c710a768a7ed815225f25ac95362ba7d6b
z87aba8b349bf1d9d9375e4460fed0a25c38fba5bff2ea1ad93723f21a61ebe47cfbf5913fbd9f9
zceacbb2d513d1be87f993591b424e133cbc5ce7686008ef0fa431fa0091ea5a557818389d27719
zd8f535ae43781bd68e4751b51dac779c6252558657e97bd3147381f2a5961790da5114b8619dbc
zbf10b926e981073936376389651287eb13b0d12c3d1ea8dc383d2f9acf87cf3d65f28be3c3d354
z283d115279b8929e24b0eb6a0d7e905ba32a2be68fe6506a82a41197defa7b9c759e0353e6ecab
z9e85b683ed198c7cde8882be216c0178d74ddc898b68e2a9fefea495707f5470a87a40b4cf0e86
zccec9921feac0fdaafc2d9ca60c64c11f335686836e086fa9c9a21a7d88d9ebd634227a794cd6a
z604517e673c2f628c04acbd127b09723749e3f10e4871ea0efd9d0471e9d2c33b82cf20ad27a30
zfcba368a03be29a798cb1c4011be3125543e7adcceb340ae5a7bbedac04b2581d85734c60d8e15
z81ab670a5136cd460151b7a3f2cd277874ef65c8a86a33d26dc07ad3f3817f7a7603c296c486a3
z43b7001097ccb3b5f52b26146ebf1007a2149ec31d875e04d8cf0946b64efbf11413dbcaee003d
zb2728420d10f0e4e5da2cec042e2aaa7df515a7b67c91205b61b0b9ed97bb8dc6dee2e4792a6fd
zd24b6111c4cefa35bc5610fc1c896032e615eef7ed8edfaaafa636edc542fab668908ed49c2618
zedae82d787e68786a3191b56def2f1a8d87519d13092c274e53bf6ab052055ee5efd22ace5226d
z455735b4a8b48ed094e096f1224ad7174cdf0b3236f2529a5b0c5ff431a1336e4c0be841219b52
z371daff2da99623b0a74d2e47d728b51d49b6ad9a892a1d3138b2cdd083a462b32a2ccafaa045f
z4b64dac1d3566b325aebda8f6b2903285b352ff80b827ee474a309c1969c262c38ac172e00ec66
z6a69fedea0ee7dbe1223cac85900f944dd1962ae181b5554abde50d2524d4333bfe6ba9ede28da
z2fbcaa9c4352e70f0d9d049765eebeac8bf09c679973d1be70a16b516275ec5b8469e3f0e2705c
zd872b42fd4ec33513218d84548e0d8b3788034963a6135f76556d69a43f4fb7f67d65b9d1a6578
z0b47fd2d9147caa33d7063b4cdb45781017833332693986f74a32ddeddb72fb9ea97c80883cacf
zb9ad4abcb6af57f990f565b41e64c030833362e1595f0c15179ab12a72cf84f240cb55b078eb5a
z30a9c698375a3512d654f76b0d8ef1afde3aaac5de700230ee0e736bf18f1a1a821edcc302d897
z14870471c9590a884a3e77c7acf90445b5966670ce55a646dbd2003e3f47b54e3255be9940b8a0
z120bd3a9086c88bac3ffaced1b4a4a8a4718b06d0df55012ae21047240144a5bbb74899c734bb6
z4b2709ddeb94ab32de298653b3635ae549e71eb767fbe13b01531000cc5198fd7c5a203d998063
ze441771fd2e274fe464bc55706693904d3e0f9bd387950a20659c8ded7066134fc5ff2fe7732b6
z96517e630064b45cb8f170664ae80e86e3515089f88d2d85c74d83b04f1d96f80c30ff387c1c9d
z4e2c8b062d7754e097cd250821da33a962c75b53e76df3a1e561ed9b4ecce57b17cfa5ece2b708
z0170fed3263535a14900954937bb604517713c38e9f018da4536b155931bfcc34c0b6632b05422
z65f89b0e6b4f62fa7d54c86008135443a0a6fd9557e6980ae6fa580d7dc553e7f6be60b13fad2f
zd3d1de5da443e50bb25520c6a6c9eb5ecc03237029b4c63f03dae1502876623af7d0d5cdf2af05
zfa4efd593a6cda594052ef9c202f9bf8ad638c993e4774b7a54d81985c146cf3cc7d53bae46389
za0571bf436e741af8c488e440b6d6cd70a5c02080b90351a1c238f55ccdcf5326310fe4bccdff4
z573fa2f75ba586b3613ab11038edaf48f6e0df8247c77d31623d795e992904f2cb9b8a979bf031
z189e7b6bddbc130994ed7f029e636a9d2980aecb60a9256eb28e9b93fcebd26fcc106709124706
z4839e2d3624e481c1627b842546ecadf94d462e9ee00b836542366bb70ea513027fb8b06e555f3
z5f66c6b3ec63cb0716574561b5972b39dbda306c9b6df276c1fd48323d86986d7936e9bf8ad70c
zb24b3fa64715e77c34e093dcbd9cd0acbb3346dcfb35890ed7720e3681c97e2dde1c7aa3eb83a3
z4544a9de80af0b9b19eb27449f8e7b12ed92742a976964036dbbad66f1f0cf217d867179b7abb1
z7c9113f69f71c81bbff68fdeb5c5e78c852db98a420461c4009f651b822388a6bc76af9e529554
zcdd61fcb003bde154724bee25adbb46ea098528b7e19bb67213c38d2cf8b5c4440f5261a665a1a
z588ec74a5130e138f53f1b69adb6e651373df64d87bd88992c4a63a774a0946221530d407a08f8
zd61765a1f64aa35ba5681cb6a2f3bce00d1f91b8b7a2837fd689b1771c203302ede8aa788cb4ec
z6ce9731d56155876159abeeaff200f046ba4b0afd081f477b7e6bb2f53e3b57b00786b7743323b
z118aa467b10498edbea9ae000116db642c78505051d84a14061559acb6b5f32e177b869ee9eb40
z8ed7c7e7042cd5f532c17748539ab102fee4a4bce4589b853a31cbe3e0a4ea3cef40a02f5837fa
z728a2276bdc0df1de4ce9def6c070919516d75258067885eb09350ff14bf7380ce068106ae281d
z2dac062f65d271665a888e544ee86c4371f68d88938d78e5764971b2d0f650e84fec143f3bffdc
z145e90d52d895b446c2989965f0c0929109ffebae5775677f3b24bdd8a6567d0437da97d051f5e
ze4a23362e193e246910f7bbb81fad848ac21b71d544e598e6b55e2cd54788c934168fa0c512c85
z0b7efd544f001252403ea62172b1a5063b15fd0f214773af783f493d136c57bba9100756fa0e0d
zc24e21952516e1d7fecd08bdb032ae1a1b1a5c42efe1fc15eccdd43c1ba8d658d8b09e17d5e3af
zbae2a22ced9893614bcefd28ec62d4bcaa5c4c227ad24002ae05825c0ca211c0741eee6e44d4f8
zd67d0ff251a67d01ed8ee5fa944d995896241384e4f0dc867fd65cdb84768c9165132469a067a9
z85fce11269b9a243757429f63059e9f8ff66a4dc4e8087f602e239783a40e842b45681b7497c0c
zc27e0a63352cee89c59cfab30b7b6a91c2de36539eeb67437cbd43104112d1f208d803ee269c62
z277a978b0148497f5592b3fb63e5282bcebb436e73e5c6f6170de17442651e901834d7a0f1e2f3
zfed547f2da3de63778789f1d6c67af33c4627e4d1e21a3e28a59f6c8ee6ec4e72a162ec2034b02
z18cea2795e1c6436a283c31a471a2c996396cf3bac8e243d7d820b07df71cb767c7bd1d333ed51
zbc0fbbfe759839e4324dc6c2066a06c97fb9989bec62eda8531e9a7c6253c0f2aae3cedc894193
zf94a24becce96a0b5e00d06e013f2bc3f8d3ff2783124a9e3e5761a043341dde5cd86b729ce6cf
z8b094dd8e16ead9ad44c617770e8fdc3331e00a85b692e6420e829d0f9ecc1f4c6959c7509647e
z748537fa5206323ff67c21028978b00b6e4a034e8d22a1f2b23765f24ac26693ae305540e7a8e6
zac1873168f9f600091ee68c5ce2fbb61e56af783adfe96c912b43fe09b3d36d496e752245d10fc
z216a34d0d6dd0431654a721ce5be2fbae2e27b294fec3637f6ac2a1a0d4445e2369d20f2faf35e
zbc20c428b5916500c711975ac4e9814665abe93204b7965a35f7d96fc69c77692da4c383d4f227
z2e07dbc1d7b6c8136719a05e90df573f2bc42cfa5f65900d706460891d052ae24ee7ca46c980a1
z8ed525ca67c1389ec772d886466353ac4743838d695331d493ac48ba90bcf6e1e56cc8a38e0f8e
z18a728907f12735197828dc26453acd434c3ca7f7536f848b7465d84619b5f0ebb22d5c1e76d4a
z251a8ff5f0015bee42ff69301601e4320af1b68c2a9705b67139cc4d975ee65c567b3c9a22d76b
zf81ad6294e473158b614228746ac92662e532f07d37abd1dedcf5f694597714941dce0ff22e654
z23f60a74a2fd9760e53403f2ceb4e55c96271e6ec699b9086127e9a095a377654dd4b5634ac62b
z94c3c44d5ce86ddb168c6f5d4267f07c3c271d452f5dbb404d818bc3efb1f4b35d9305dbae6d50
zacd83d9f3a6af770a32e4629c4e342ce0223f2527950f5f54c3db3568512fb16665ce93a4df68f
z65cb6de86b3d7c29a3376326ef0eefc04d5c10a547155811b86eedea64e8989f39aa9fb96a1d15
zdecd2199c77a4a3af5d61457af9cd63d92772ed319384c47036d1c6c7906dd144fb83e370b3072
z2f6e9da3962a5e3a4e84f236e6d4d9749128b0a46fcb1d22ab30e7615c607149f2a8f8f9bca29a
z63432eeb93a2da82d4ce54d02fd4a9a86d0304ea30454f3707855a01de48a4f9aaac2e020add22
zea4ae4af821e051df13768870c5b4853ed10bc392cecc1c37222d623b834c3e2490cdc3973ce43
za9ba3b441b6c4d87bcb51993b8e22c5cecad0cc31ba3d398b2c282154a3f2bc7a039c0da49fadd
z4b913998c7d63baddf2ed584cff5ba5dc8f7e8bc460ae4610a3ad2c6e1c4bde82381b846d39278
zd11bb1f06c8028c97b54f79281a4facf3be0b96124f67ac36b52a64f9afba19b8b883834897644
z1bfa1d2d30f6ce36a14cff18e7b372bad4d7fd388a9b94bb3a1fbe8db3b1c348c456d66d392b2e
zb39c14c9cf4022426040517acefe82843a3b157e1a66e4267e8a3b20f3c2ef0981ccc8629b36b9
z896281f60eeb0ae0b6393e3d8aaca8361e4ce9551527ecdc8049e5681d9f1edd737181bffe2f95
zcefa34c9a123c356507f852922d0d2c6acd60569d476abf09d3f6ced12dd85ce7cefc8d75d324a
zab5facdb6bbcffd6e4971fc51d6065635417597c82194b9d0d65ba91d5b7fe6f6fcde91617bae4
z2e4470703aca38aef28a1fcd92b266049f4f5dff8150ff3434547dd51ce4e01c86f0516cd741c0
zbff7380da5cfcdc1532fb26e96859af715bac6c5527be9141ca9b3955de3d0094acd4f6ebbdd70
zbfec799bf8d1b708b1aeace9281cfdf75a944811480ef93f0b2bea55861d787452f010e88b7f68
zc497e7e37c6607acc7d6a0c8d696857332fdbf4ffc03f6fc33af37ecc54368bbf6e20049266d28
zd404f27f8e48543bb51f05734f941dd2acd04e9472282a5f76ba280e957ad7ec639a70d943121b
z6606d88bcac21bb2bf0074d0467f1abe9fc3aaa802d4833509e8eea70fa44cab5df22103ba5427
z6e651a5e609308b6dc1c4fe8fba3f1a7eae9ee1c9de46a9942efd6df177ad102f0cec2b34d3ebb
zc8fdc9986992a9c1a3fbbb180a5921f838aa52679e94572c7aaec3da4e3364a46785a6f9f6eee2
z5763429b26d1d21547b012547f847108a703143cdd56f70d8dd04a386e2679c97ca81ad1edad9f
z229da81a58097c50b44081a7eae24b3b5aa1ad98e23552f972a999e6987639e3d9205b73fd1b85
z096b22921e22fe53364ed859e88a37cb5a16f9b7cc04378849817da1d7bd4ba09a018c3f0c937e
z588b3c9e498fffde76c9603f741e0beed68e3e438a975312b246fe65c965dac1297350e6c0a34e
z66b4c137def2666bb0b66e34bb47e53a1b5d61a40313f15de3c66226826263bfbe780012aa0b53
z3d6def03e33208842cddf210d331d09e272d634c114ad4e1b2a631d313ed785301655cd2e9d686
z5ad3481c537b4e83300c51ff9a69d0ce8c0f81d7c8c74a5bb8a9d013ddb19796e7ddbd06467f80
z867ddd0a002766a5ed1844c34ed1a3cb0e17ab5e78a5b038db62ba9d011fd0a8ba106743dbc39e
z41d79d0103dc1207e711b0eead0086da9f5347df6459a29ba159465d9d799c869e868a1edb4041
z6a2426718116635fd3f9f2b506399bfaa3c7dfe7b492c5b4d908e0a32e0b1f7b2806d0ce638b1b
zd69474d9e5e96478d0d0264e2b0b127c8449b61ce38897260422f1690586d02fe9dcd372bd1c70
z082983d07eea7cdcf01c1573216db2c9b3e11da772a65e607c2426015494e174c6dc68a4039d78
zc3675a769de135cf5247e628cc1a42ef44bfeb5be333b0a0e5a40ce8c63aaa7b343c0124ba6461
z85eef2a1bc133dfab66702865dae1ac039ee68232e5c11734261746c7c09e3ce59b8790266fefe
z9698f94a68134648563117e7e6f7f34f15b9d2c202e4ad4f13020fb3199ae2a7fc40aefe1a6c92
z9c36337dfd5ad084d85b54076c0173ab8e766fe7a50ff1eb5c3cbb5622ee7b915a89e4e61275f1
z0e3bc255b0dee24323dbf73aec76126b8e14bec366b7f2031a15db8dfbae3e19dbc6152e49d91b
zaacb09fb9b9458135a0aaf244e9d6cf80bf3a8ade2f1a895d30ae8df5a0840c4ea446ab2b755b8
zc25879d0c3725f023b1d9be301f9b125afdb16e390e0f89028f62c2a32cf0cc9129c7f67feb2d1
z2f0c345d9d25b3797ec8a0d2279b3c81bb2fe53ad913475fa2146666770323fbad3a66aa0337e6
z2cf47de8cab47ec6178d8d259e0468d8a2b86e82174b3bd80550794ace416e4162d65a56508631
z63b42f7875f3897c776492bb6a0bbd8f31755aab3a4b82519ff86e17070a55bab2c6fba5c56939
z0f37c0e14031ee041ccbebb3bdfaeca2a0a94334559ce31e8ae0849ca975c14ab172d9a4b04ee3
ze3d1a62ca824d2019a8c27f43f744ce6317147f79390106500643cbae87ed3d8c63b3b64fd5864
z0ea318d7465abf36a9b2e7b0d223d528655d97eb4f0df65323e42404fbe23c180b3ee7e72a13a8
z6fc94a36658dd8d30cc9d532e3c7448f7427ccd9ccd1b74c258aa4f40d6610fbc81eb8578ca65c
z4937baf0460448e122d035a9a33580cfda5f31bcc2ebad95094c8324d97ce6d9fe8a9d25f7092a
z4893cc8355ffa716e056198e31f24189b3bf1bc9b15aedca16cdbf3f110ee6f007b94f4cdab21a
zf016981c510502f63d4d9d3edeb40d25307fccda137e2c4bc3a6925822585e18ed4a58d47f98bd
zf625c008e491c58de7467339394acb0078f373fb9edc01d8ede7f1d2ef145a5fbfdff761b193e6
z64a196c7ab09e1edb816819b52913ab52c7529fa71a97e83bc1dea451f9e67bc6586e61ffadc57
z7c5004e22041fe55d83ec9c10c56f99d476533f1b871c3f60114b042e4e2a094db528a98962ed5
z5e9d602cfe6914d5ad4ac7efe8550dce7d86960eb066a569459f71644154e9b171b42d3b726ff9
zeefec6a53791847d0f48e6d65fbd087beaf5c15db44a6dc7f4b190258857e31724ccd347ae1957
z59ef088e51e5df35309ef4fa11d880e0955cb19bda0a4557065cf5fea8522615c9a3578addbee2
za91a9f9c1f5ad7292e2300ea62228f4de436de15a01a2d115740f98cb14c87f7d1a0ae088c1aa0
z4e653d6e67451c9530fe9b2bc8df143e8061a5a167595f33e08d499541549a45ae67b1246d0c60
z5613348fd54c67601de63dc4d9103ee3d0905bda0829edf9573e849c8cfa4d8f8f2a50018c4f4f
z01aa10308fd29d2c22bd5c692e54457f02dce7d1c83f9bbd9e730b073714618cf5629f901afebf
z1bf39e5b3973080e7fb4271c8dd67c2f86563bfd0fc127dd4c49cc26809006fdd2c7456b0ce066
z94770cb5b46ff60e762877018f70c39fd4d29f90ea81a6896f35857423e4a613e7fc79abd22e9a
z4c34598b9bf890670327cf714567ebba7e133ab879b8d94b0b2df1f00e8753f64e2ff131ddd0a3
zd62d5854efd2936a80dea92156c04c8321a389a090a7665c862d09331a09c469ebe866c7653aec
z681675b34f305fd9c24ff185ae1e4f71f50ab1c399edae853a807bfea5362e7622523040f692c4
za527013e0ca08be730577a772477dcf2db5f612e58f6c8d4a49cce7e6885e16d6a5a51d4288f62
zd671d3d61e3d91688f4255b39a0f94c92358b6b19169da95cacf0da95d427eb9ae7af9b71f1ac4
z72aca40cbadc791c81c72121846c4f4b2e3a1fd1a1245fe1c4aa4d64b25c8b80a3dc451987a21d
z6a00b146b8c43a3e91aa6f2a77e5e7d23dbe4f596ce6c37cc36ed5b6b66138d56bb4e0d1a4f1de
z870f25e0e76fc0b85f81942f4cd9c337d3f3d7c5a6902fbc705c7e1751a741d1e30941b92b34de
zb33acb1870da9b7506411faaeaa338a8bd2c95277e6396bde0a3308c714e84dfbb8b599ccf4a37
z2e58e7cc99077ac84e9441e1089aa41bba250411dc1d5aadc50dd0690348bb417e1c9025c3282a
zc8a78909ef3ab70317d189c7264de5f2342b6ae2f4fd1b47ee4ae01e544368cffd44afa9c7d545
zff8c32f8e09ee5c8e9ba8073319dab3588cfb89131579c8a5705fbffe409f9f8290e6ab5e5b83e
z66864ee25c5baf7c5e317e1ebfbb6e9daf791df5769369dc85c6e2b719389f63e0c40b1c152689
z2926af0454249c7267cd525858322c4b48d6adffb213fb18cda23509960d577267e75e732e7076
zfef75cb4e4d96f7771dacc66b26b9dde2a2183a62a0100e622a9d08a67713f0189b59ad556dc17
z725dfb54ad7484f0fd6a1087fc1169e1b3dc652005466235879d84f471020a22d6fb373b133512
z7bcc48276f187c2dbd2f5d2821a717f4821f1570269e9f5a5f615e9de3c397ab251405965419c5
zd78da9b7af5e1d8500c35bca56e5a54e8bdfd6d68e54b0d16ccdd89167bf7a974a88b461d2dc56
z1482438281f0a4f32b62100f3d08e0353b6bc54afa4f6434d4def599d132d5b49817e70527315a
z8a974932f8cd02f7c4614881aedf0f0ff9362c7d9c3852c516e62635bcc2a9f387e6085d76bbb0
z0be4154e6b7d6ea892e3c5868b82287c609f37eccbe2535446723cc7c953e8ca353ab912b1363e
z3932032324dbc31e4f3258c2c1ce6c1d13991d16c5e4683a7f322142c3b7da66d8853b92feb873
z65f951560f8878507f5220d761a9c9da1413d9809d43af062bd6b5e26f61c17063391bcc9d30c0
zd6aa5eff3b8ae236359a3174e63295201747033d382dfb01b474667a198ab90e75289fd47eda4a
z699cbe74adea646ba0f55cf0d764d3f441d206b146491c354a5a1ce5f7584724f062c3d9cd26cb
zc3d68e9e9ec022441e904e3ee45a7751c9136d28cbac1c0161c07760aa7b3e0da11b316df9fb36
z91b1fb368da3f0c7c295d84cdaccebb2b0dec41e33ee8f79cb9831f021bde2f0e67427abe33b19
z15926bc4aadae386be757a55cd0c90ccfe35dd000fb3e720717dfebcb92707c585f0c638b8f45c
z2a140b88aaab9238c8d73cb534f9f155cf38dfe9280b3d819701a5f4f48afc1e0ca65ffe42497b
zf6a1c6bcb5aa4ad94a4939d0f9153a1a3a733b51958effde8fce299f09657776cbe3c6af73643c
z39b6eebffdeda2a42d992915275494fa830427e1bb4a209c89748699c3e3762f24d63205623d89
zff4ad97aa494564fdb83ac1335d1b063fb02f160ea420e5876d5f3fbf4a1d6ad3dc3702b247858
za646a4c1162d632dd18236ed835d8cd2b21db0b6b8c7134338de8be9a303b34a084e54214a569f
z678ae42feecfa548ff867f9bd1fa4624368af37b09d2d04de37d0c777fbd915aa4958966e39935
z7b3a1993443607981ad9e6dcadc9650f2ffd61b4681812d90f4f69d93b167b7072ee3325688987
zc099e04830057925ff7da5f399d2acb389ed2f34ba0eb67faed7c7d6343a4b480590683142b01c
z147996757f4295fc852a8cc3ee99990bceefaca76472410c6ad5276e73c10439650d43816103a2
z65d4427c4bd9f2040c6094c85166fcbd05b18732c3b20c28bb525bafa9ee9134830f1df9049a0c
z957d3cfc6f32ec8ec3ca5586fb25ac1485112e772ba281e1ca7ffffaef8a28e236b7049d12ab42
z419abb1af9b393959212693580ed1a59be920b52b9b7932325a7730cbbc910c24bc3b02672c23f
z5c3db3534b8bbba5af5fc52bb51941a0bee62020fe4d4c9b1e7712abea7627106713d155ef3b80
z0c41f842ee6621da7fe919d9eb0ce5ce9496c204c1ba4ef43f0c222729246ede8941546d0ad2de
z137ce07a6722f1d277f68dd408d6c581ddb90d06fdd8b6862a1e42b8836d33a3614c1a4f65b0d7
z77be3fc67fe403ecbb89309d5fc9a9a03ff490caaa9dcdd7da70a958898a7a14829cf38bfa7ee0
z99ec3ee2118db8366035618ae277173a5f3a5d0c35bb58cf94acd89b730c05b7ec74821db79c32
z3dcda2da39130737dc9b8858062ced0fbd0f261c80590d8ca6908a849c0ea94cdd1123a52d55e8
z8f1b763f142a77cfbe2c992ab87e5082ef117fba3a7a76423c1029b6be5810ac5d470b1043fc1c
z8aebf0057084900292b43aa1d31a008234cb02b5ed2269433f1e49df0101a705a07a3de789b322
z068aadfaddea6132c830999b0e564cc0e73952cf70a679cd6abdd133970ea2716c2321382c69bb
zeed951ea7f7ea411d703f897f910076cd74c7b512704f98569fcdfe034d1a664b26b5d9d6b697f
z46abf0ea77e5aee7eda59f5379c6a0db3eb566a0fd767d8db1e8bb34717a7512148c008ca213fb
z485b89221e1c6057be139b48ea1a20334791fd3ee82cde31a0d14214e8000d0be8aa403263b38c
z4908330cdc23b624214aec29af39ef788b6ab21e1ce1ebac548bc1b502633982bdd171209b0704
z38d7a068b69dc1484b231c0587a518ef38961d5254eb9d63f5bd7bfe90ac67788974a1aefea940
z984d3fa6d59901bd96308580d464d5b98bfb2519f9dc0e542cd60995b122532fce3e59de1986f6
z0344cca97c18fef3e3b8b1bdb463c378a2ad7e71a0b3bf9ff5a5c4f44fc0b4c633e51e34e78248
zac55c300a273c725e065234c29358555189845133a600396d8c6ddf34fcae6b9b57fa273766119
z2953cff65029424533ddfbe351a6f76eacdb1d3a608381723adeae4dde88b06c0aef37ec293697
zc9ae4a1d6f812a1c1b74fd127cc001afacd7ef50345563922cbd90edf3ed405a6ebe8ca824d8eb
zf96db6634e3a9e872fe383387b228ea5a28880d4af3c5b8e8cbcb051aba79682856b0c6c7cf5b9
z2304b04635265dbafb8f2aa6348ca29c0375141c898f13b1da759780e8a19c9107317dd3ee27f0
z331622e78284a8f65d5f5d6c9ebaa8ce6143613328e310b4fde2d51525314ff60776ada9d5dd8b
zd0786a4948802982f679d29e503388cdf2e6aa6accb99b076115691105aaacf4c1ce23dff676f6
z74ebd505fb84d0648da70f9ee53a91d5fa99ec9a65c529c69b28baede502dc2647796688ca4f9a
z0bc0657d4a897f937ae5cadcf3a450dd9bbc1a06ddb1bc5a9250a9086a88f686bcb3ff4530eab3
z272e1fb725cd99196bae6bcc90cebcf7628baef75213b951c72d95f621067fad3d1aca6bd489bc
zf311768f3e44e178185eaf7da9f3ceb44edeb35069d39d2b0bb24167ba7be9188210419f85acc1
z304fcd22143e1dde1b41c3f2008ba46dc72f797bba250b5cc76d6c68fb827d6cbcd3737e39ceb0
zff10b85cb8684c2af7fa7f53cd0b39b7e19d4cfc67be356bb4287b20f9ae2aa2e229d4bd202634
z2df65840824ca5c97c338f2ddb40000dc4c9d47c95982c80be47b752bf05c0a4aae71104151679
z8bef696110b15f663567a4ae32f274c53fd8d21c5e7c8b7c941c4094c4e8fc8b4d50c1b5c70dd4
z5830f80a9e533983c79103bcbba6a27ab780862e56d616c104f920c62bbae250a1716a7173f664
zc11589af3c43b540d5e0d4a769c49ffab6361c38133c5ad67d7e9de9a5c63d895f0edd24136100
ze72107682a8560a1d0cdf0a0459b1771b503792b5247e2a1ceb144d9e263b55bb3540456017061
z6fad4fe4edff0c806c8606d86fbfec17cb1b556ee20a11ea86daf446309ada6a4691bd23f6eacc
z3997c1ffe2b67b38dab8936203029b47c1ff122bfdfe59e232c2d82d6a1ff911e72cae76a677a3
z0dc1c2d73d322b9fc1ad12f07d025f73a7646780ae6881647980d64e61d048ce2d9817517dc534
z649a847ddbe811b0097aac9fae717648d492ab5b454f6eb8c3443bd3307ad72d62c476ea2e89a6
zd2a37cd8ce8f96b4888b1e05a012880cf444e5fc7ba016c9414fa2e9b992b823b126bf3bf5a584
z994fd1ab17ce8fe1820523ce062bb7c4ea42ea35d64f262e48cd1aad87c7d7d61d872904d08bad
z7ce17b41440721d8604faa9b34dfa12301a0bc2d19a8a8d7826a29df5f722821f6eb13ce19377e
z06532e88a6e2936d7680e9b1ab4cd8afff189e4da1d903ca31bc550e655aa67861a8dfdec4d4a4
z05484fa95422d11152c2cbc45704a9d4dd83fe94ad87c1ae2a723d019a58d03946a320189febe5
z0984a3832dae0cd40d1760310c7f49a6924034c12644e72ba22bebe2fd8778e4411d27e7f4ce03
z135576345debbd038824aa58995dbd61ef0d5de9120c73debebc65b3d528cf851cde8044e7dff4
z5150de3caa9ac8833a5c2d5a186a4b658693baeb4f13e40ee5f7744c70e0811b283ed100a10ddf
z8eab72f643fdefd45a3c305fe5964c9db8716485df648ea88753606d63a1abacf8d6c643d3b3b4
zfb3b59182a53ba964e32717976ebea982bfe512f7e7bb65e7d7c388bdb78dd01913c5204ae0e3d
z65cab8424cca66e983e2f6dd23200fe808d805ae64c6f0278667819aafe56ca23ab8a9533f587d
z77aff0779c904fe9e275fe2cbe2e69786a630b3d58bf80aaf064870fc2b6ff3fcb33e93aa74d4c
ze7eb8d90f60eb605923c9223fba61856b1698db2828f11acf113834636fb3246e6138ed3158e35
z1e1918da52d9c2351fb82adc858c81c7055b55cbecc026b90efb2cf9b93abf9c5654db3726406b
z267ea90ce54ad65cd59dbe64c98c0ff7b9de0deeb93e85e2a8e20fd29ef8f539862a9b854499b4
z9b5c33e5a09d4349b74f45779c8f2f6cc05abf0f26c342636d13fb9ab615e9c1a9df1c73fbef27
zcfd8086b84983842b8a6f5f98e76b144adea079eef3fc80fca8027cae3ab78d02afd9974932a35
zf8196e94a0569603078bebc67b21bf52fc2dddb80af2a14e9abcaa99fcef2e6190573ed3e9d715
zbcbcc80c9695afa8934ac45d66fd5497a7cd006b21ea789c680dad045a0cb1933d91d866e411b8
z699ea6d16c93e528be1717f40a17cfeab260cb4cb101475620db871a686c1a3f4265854faf38fe
z3b64c7a4fd4e9b74f925c63243c8b2a497ce2097d8562b24baf77797b658885d9793e8e87a865c
z34de4bf40e7be395198bf8c8934106a09a26ee09fb1593814e4fa158041bb8f7b55d8e944099fe
zb100a894717b34736d3c7c56f01ab23b4560c929222914f1267cfca8d489aec8f1f6b6c07a6783
zc44fddb75385f19a91f9cd44aebc648e603dc1df09a3dac0c64fec71f5e3b3e57c70e273f7593c
zd1deeed40106a7fd313ab13e636ac2e2c709833b99119894eba4d6a39ba9e8dcc20a060ee18e7b
z97935ff830df168f287acbbdb7e3d0619f677f917f6f2c0d5662dc80706d1dfbd2f1ace12a95ab
zff941f1831730971d1f0f87007e342357146d54f58f5b981a9504d1769cdd3c572c8f6430d3488
z4a928b0fceb99992945aa2e2bd6b9b2cd11a99cabee79621b9628f1b20d1c3a8f11f6a46aaf22c
zbc2221bef4435445508d43fbac353e7e30adaeffae7113b90f7326786548d28a9956e345d8d2c3
zb6ca6fc4a632fc249de5b7eff4d0335b4f37933a40bd637db8af41d6d5826955e414d52284e02c
z31de531778ff7582aa9a55487a88cef13d50f9c97ab10a5fcd9937daf0c5acebfb39dfdd1413e9
z3563fc166ac586eca169b09a3c7795aaaedd2dd4a315568f31b0d56793c9773400d1093472c6a9
z7e6487c67a4e880e0d46e56047231cf5036937ebd9bee3d77dd0c17811bf70e201b976a69dea64
z931793756a0aec6b6623d94ce31e35bb56b64fdedc291dbb143a887c6ba932f77919a7a05cdc7d
zaec84d10dac1a4a8a8e916f96af871a0067f604bbd0de85071ccb24b600932302dfc0877d81311
z9fc39ba95a3feb6bd90e5d2dceac77f7e4408553336ea578d1a88a186c52112fd5e4f7bfa8bcf0
zfdaea213a4b573f10a03852c9943c9a46752a79701bb84e59ee1f37273a7b68cf5678392bc42ea
z2920c940ba1e8891b2ae1eff2e24f925684d19d07ab67ec63ed7748bbebbc43217844227bfc1c5
zcd51b2321cf495bdf7381e61e8e613ec59820c61acf7fabd44dcc6eac882ef59d2f86bbeb43369
zfa46fc8d081aadcecbdbaaf3cf8c83cfdf8160978f663afe356d1f05ba5e7f3f306008972c0f0f
zf84dfcf73c3682d05733b45fb9111bebeaac5f7823c7fac649834e42eea8f146477ac5ea9a4aa5
z163d49e438bcc7e8fb892a658abb1fc35a0124c3d5ec8448e9c40ad261b9013af1298734e31e46
zd4e59ff1415eb70cc1af177e42022d39713263576b02dbebfd0d68e48dd95f2bd526f1ae28c5ca
zabf892a824d7857786d0824eb9467553d72b9d71f6f259848a65405725314489c641e820611eb1
z3286ce7d8da9888dbbb27e111234ec28f45c947e0194ad8e509d88276fa308908a0a8fa1f277e9
z216d47247e713aad3bd343934c6b7ee42816c187c6f5f4e7636074b391d4f63b4f4439ccefcd5b
zcfb31d97070b05e8932ac652b281a4fef75e771967062c4e337868aa0caabc55968c265fd08261
z15793bdd582bf847c2f5f01112d9e599c96133b9d82413c0b3a64b48d0f15791d71c14892d745b
z5ecca3ce785a67bfd753b2501a0f687f0553a2f91596945ab078d8ffd3f6a10507b734f1657442
z24712e2d9ecf5722a1d67f415f73d28ff0e3898d6ec31a81b19bfe1ec698955022d1f616a0b5ea
zda18b5748389f7c99838d6141a8c1e2a45ec68eca2b333a1c970d213e990f87446d6d96e82a1f6
zb2e9bf719eae57793bc394ebae27af8f3618c49cb460e097b13cd3fdf701395dcbcf6ffe38812c
zf333704c0b8e7d88d4a35f78b019c882d032f42da9d23517397aea9da2e83bd572574972f3f246
zc233fc52116d70334d10fdf65d230150e2ee43ad324ce38ed6c419c50cd42974586b044091db0e
z98452d1d731f3a603f75933ec94d6660563b44933e8f4d1ccb3bb5f98e31602b4bc03d0ee56900
zb5cf928ea541bce440ffe3ef28358b5a6a48b17d140c5b58555eb7bd3f36345064de5cc7560a9f
z67a3a660914397a154e5273112729787939bf3118c3aa4ebb7d822482d7a9d62d325ed3e5acb19
ze28c9f6d71aada49ee0fbdd8e049bc826122565f11312a3c09dc0d4ba50ad7c7562358150b2261
zdc23955677a2a2a1a366ac4d1bd72017e424052296ebf1ab63fd06805d6369f5de2e97b5998884
z179f78953dbb6d948086f223aa4ec6ea1c0f6bb1101be7e0107a1838178f3e7dbf5d5bcc4e7cd7
z8715d383dd5fdca0932dd377b9e4332ec8390b056471c097e3cca862e813a38a89fb76973b6fdf
z51a876dc00293536ecad491b1a3a8225d62dec977c8b564c1931d14cd01b01e742d279524889a0
zc1a050ba5e49e4729783804e9085cdc67a4470b998957095b89da91bf86506814ffcd5bbfd6def
zfe171011d4ca55caa2abe8b0add73e9103eeaa14f71a1d6de74786f72e50b74cf0b73e74b45d48
z6c041159df97f960b091007e0569bf548e6193aef195a2d4db0e62d228dd0cbd0f981564b27769
z39cba4d50b9319913302d0b7066e595e260f81d3a8e08253de08b0c1068ddbe7dac5ebd88a29f5
zfee53e06cdfa3aaa12c8e28a8f2c65b3f94789de364561ca94295c90562e0fd7bfb1fb92334a56
z8a74926b4dae17419f3b8272ee2a37a9cccfaa3de1703b3c501db4a8fd3887e360acd0b3aeba57
z12c27d2f1b1560c3072588cc6374e32eba029567bac73b3d2c1dd9a1ac3ce4699a518b927f0510
z6021ad0b0330b8036738337069f6495e1f3f5ce7382dcbfcf0a40ded406223823a0ee5882acc07
z04506c5b02b0284a4ccc5aefcc62fa116dbe22bc9e63c0fcb3b4d9deac24ac6e9b2b21adb4a250
z402594b751447dc8a7ddda66ef23dda6235552538d19e9ff791a008b29ae9912e5be97f3e1d0c7
zfec04d12307369b7e275d6520817b48de76f0ab88c085a34e9480e3f49495fa3cc7e185f5045c0
z3ccc507af83148778672606a4dd087aed94ca991ef274715bef1cde45abfd20c36e348742339d8
z84fa79f4644b5aa32a1c017cde95089f124f9455349d1ca60200c94ef7f771e9e8c42d13e4ce33
z6e411a07822b5ee9f7a3713bf94446f7fde11b56fb337f51f367814b2a2fcb62601f8464d789c8
zff0817914b37e840f64984fc5646f535520af9cca44a3d9037413bc7ba499f81edd27260f0c85d
z2bd687de2a1162b783ca341740f62cca8adf9b05f4714648a9cb51b6609106739ca2a13fde0890
z5ba5db9844852ecbbc012886cb5b76913193effc1ce4e49894d18a547aa7486b76a30bc41dd1f6
z6bafda1337adbc3a80c59d6ed6d4a256929485f3a46e3f25106950eaad8fc47dfe4c412cbeeed7
zff5740cd1d3f587aa902c376fcfda5b91d8723c5d5022058e8eeceb3bc2c4c81d18ab79178c010
zd4da09efd1c89aec87a5ba75ba69fc6a9bbc3b9cc097d235eb45c720b44586406d627f0be94f67
z808a04f60c04f917e0663bb2cdda26b40638b6040b1a11160c5a011dc668a2eedaeb69258330ff
zeb188c58e7695de03c513a9b7761ae16448699f8961ec44c5bca3bc67f36343ccb58cb14cabcdd
z4297bfaac9ac735d9b880d004313e97007d652d339e5595e0af58cb31aec1d24d290baf9b7d482
z06d7ba36beb0c29ca2df8ea2d214338e803952008a3892c65dd0e40235cd3228b03835abc40548
z5b1910f534ef27bb2189af17682848893e35be8636e48813f0588c892dab2e9474f4f61634d51f
zd5117df661f9ff310d647dc4077714d1addb6ef65e06e73e48d0351c120eb683cf4c7f13bd80fc
z814bc7ac369324065783b4285e2b34384662bdbd55398d1752409fbe5d0ccdd440e89e1e987cdb
zf4893c9a96f40e9f37295d423e7a21faf3c93e992af5ba512f8f696c892e7b6892dc1969232c8b
z5b21de11b13d4c2374495e38ae317914133582f682ad3ce0ccb160c0a924dfedec98b45a32fc57
z4ccabec01903661c0d40b5e8b55a7f1d6e932f0001594e807b6a744ee99f182c81628500992da0
zd02ec35055bec4179e6b200d4fb407a00828d600589353931327f02fd4c5340041376e2bf631fa
zf2b9fa28d26f8bec823a4185e41d4191519e1b4369e0915255c424c9533d68e018b68d5dd37c69
zd159ce3487a63afd04e22064c675a7996cae00eb5c5d869710801012f25bffe72706fa9fe18866
zcc6a1dc7424e80d5ba4b12bc37ec00ae2f5af054860d95908fc7311018d32c366be63c97db82f5
z7c2446fd2c417fa4df84d102fe9a806c638f73a6d67b27ff0ad2246e5236f2bd7d3514e9d4cde9
z40c08b2f9bf9695f553f2f51bf6a2ffb51cdd42421a9500e2a270dc1d6661bba75b14cfd4ffad3
z1ef133f4e03024ae5e24d2526102778f1c7be34e4a8a4b9bc790a39c8db4b4a33d472270284167
z93fd2e905dc81c9e33bedd1613ee24c25c9650f6181a059701e3feff1eb4c9fcf5e15019b77f24
z9c2f0b26e238575a6746ae6c2141944105b4d94646e35744f7ce0f25fb66dc3231ff6374e2cd25
zc6385878f96de960bf05e3514907e7e5b0cd87e8c73f058276b717656805e677d66cafceaab086
z93acf753b9b385558b89806f87ddc71b1b498ebf479d41231b7a960e715a4d5ba2cc6ae3106e88
z2c44c01525e62a4a4310646cb61970f33aa64a58714df0447c2e4ff56a60f1c302bcf557d802a2
z9b4a93b5c683ea5ac8c11c58bde717ca3181b8c2d46a0b95e079e2c5e6362c5103a1030723fcbb
zbcd88c249989e5595c40d7a56ea8b2b049711721d86e7e56d022f0015c53a447c2f4dc3afba8aa
z323f4595f20b4e6eff5e60826e8048bd341f52e36c49ced18ea6474da96de0837f2d72448469cb
z31c3091c5a28759f25446cca73d265e12ea5c3c58a00c4883878548dc930dd8c03c0657c429f37
zc6c452bc7efcc775f7557cb18046e22083b06ecabf21904aeb13a34d103eea317dab2e88a3a113
ze40f4eb3aac3fed04365d1c0828aae8d421ac710da01927541078067959141323d89ec1765bb3d
z62ba0b3b11e85696d1ac30cce0933c4b469ed773e10f31f4dfa44e5d951bba690e06a670080c1d
za717a5377d1bbb936749f84b5c73a49ce511812ea266c11c1ccc7c3597335f9ea6c09af3632735
zae8b37ff0572f8471438e4b4226f949bdd649c55adcab5eb7a00bada14f4fd1392c241cbf21dcd
z9c9e6ae219107d4951b7d663b9b7fb6b8a059add8bd36a6b3825077fe48a956b83cb011589a70b
za833ddab22bbd604afcb8728494126c3716848da2dfa8fdb8e17d224fe65d1f044d6272592195b
z4d09b91cbceff250457ee1551c0e7bdf12546b28e7e6d2ba9275d646b21ae403208efba2e6cf57
zf367aac26e490688948fecccb5dc76558aeda4d473ea1df729bd638ba1625d6edcedb086b1b8d9
zdcebf0b0c65b586ac22c181f57b0d49ef4fae1708f2598eb878ea55008be262f392b0b3f896655
z1789fb5741a40f3c164313cbbba9d0931f24a3ed3a13d2cb4283896109778833730d141ef189d7
z1bf9dae6e9d68b0e22b23e47863a8d4c9e5f5586e88d8e16e67af7f977bedb074fea2547ce305a
z6bab9f8193dd62b01ea046f9f362e5df7dc64a4a2e97db35fd738930d873493d128d58231796c5
z38dba7f4f1a7bd92986cedf0dc3ccbe8bef57d075a6289d0dc10a7a9ee63f71f903ae998c386b3
z7f0a8352e16fe053f18159e089e083ff787a757dd174703220d2c396afb6b565770d1589bd770f
z41515208882512d5c041098fc483da61fde07303cdd99bdcbe1d0f460f919486c034d1c61203e6
z7c6c7021a40089b17b7799bbb4549ad09a1a87da0359c3575559e399738fca23792e832c2da484
z7c5b42ca662c820cd5a36104e860ee65979e87c38e532c4550d2c5a397b58abc7f3c1a2b6b7aaa
z8e18db7db5d03f71f0af84b4a63eed3b19dbd198625055e77f0ff014f6eb47142063a8dc7910ca
z987a644d238c503dd9edf332af192f4dcef3fabee4ea1a34c06ae46f809bf18b06b7e682b62f31
zc0bc5ed771d12ecef9b1315174396ce41b859db813b322a4b8e3ca7d2fa142033ced03f97146da
z74878fef80418468aba542e08bd05638ebde4f0dd351a4882aade415e0bedbf0db01d36a343d07
z60111fed587d3ba31a990dc4a0790f02539cfa0c397660a0ce0ab920ca1583e1ca422bc61f2405
z43dda8d8d9d89a0295907bd9ce76822daeb39e6c0420aae20fdb0f8a799c80821f09b5bdb5c833
zeab807a903b3b5e82ef48a21ec4086232f3cad10f10997c777bd2e2624a0ebced7e422aeb8a4ed
zd50faba10c106a420aa6cde6fe7ea1b796879b146b02eac773d6725067f3ad38d87daabbf8c715
zb926abfe5a08dece49da1ec7bb5472ad68f51d48339d276d0835371f7db0eceaaa1a0a6b59207d
z17d9be122963f7166cb33b715790c244618cecfffe59eb1d471beb44588e6a415ad2d8dd8d0470
z01e1688efc5b1a337feed502d4b18c55ec06b75d04295754a38a416b621f18e96d8646a76df439
z60840742478853a358fcc370ead404b7511c755ff26b6c9a764737573496a34eeaa6325c2fe4a7
zf2462c1bf9cdc59e804202caae3239bfd16a23a5f5478b2afaa09dc1a5959856578d0aac12d248
z9c41d5366dcc85f04b3a7cca3709b090d29de35f5651f7c6a7fd256884cc3e7dfa36824bab6de2
z7990d0779a4513c228fd350fd44ab92e1f72b267fa6e4f297d40c8da7637feffc5f69908be812d
z665485525817042aa577c9eb228c5f69d49d1e5ea19e5a0308e5d95da7f8241d2a5f79cea57273
zbe2f1dbb7deea1ba1e2435b0230fe9d9de5fd7070cae9379548b33adff4f2d906c486687c8ca5b
z99bc828ecc0207f3f931698c69e24650e5de9de850f7fee72b4e535adde67b24b1c1b4d9667f46
z311a0ff332accffb19a2bb0a8abf0e045b549ac7847622cb38d00a528862a92805e147ce8ef9ef
z7028fe32cdb2e8ba4db3ecda23017904af23b9b82eaeee6f64bf435545e02798b6351167646d0b
z7e745dd645773bcd4d550913bdb87cccee6c0095162412aff6a6f6a34f6d123aaf2e5e6814b748
z6b45509dc1ae9a8e8cfc0fea420012ff4850288e6ea60a41176933c98d382c3dc8a27a7acbf89a
z1e7e41ce7b736c2cb9e3ec36503637389b025e4c65a80cd9ab3f6cb6263157ed7a76e7b17e2933
z50732b943e4d363a5e0d1a0bbaf4d2016157c29497023a17084b3ca5b0cc9c39ae4ceb6f86ef40
z09a6fcb9eea233b8cb9adbc5462c8bf09e39c7da2a2f4a5c0c45177b14a3d9a268d557dc2f4d1f
z8480abe62c85852370f5d189223a291a90498e653e99a948542e611d09b49581a5efafea8fa82e
z26ff6aa2331a5fdffa1f5931cb7ce6e535e008dc9067fa0a87c8b307e8045a2e20799229f5e820
za729722640edb7eba7e49aea7b7c365e52afcef3a68d3a58ef1d019ea7154d0d903f106adf24d4
z419d03f10fe0ca045558dee454f12b5edd173ca8953f6bbf8617b29a247df3fa7fff44e8da3a38
z8661e8bd5c2d3f3299e565b65c21c6e61bc80715a4e6b500100e2373c606cdbc258c7f62b3231e
z083f9cfdfc03069d872a5115d9f71c6ac502b082c70dbc8521df7614c218321e4bdc9589560e9c
z55a5bc92f7694d6ecd7770957a97514c4e5a43bbfab87f33dc2b69a5e7a28c93766f08d11a76f1
z5ac36af3dfa95aaf2d2e9091116e1590fc0a0241a506d0d3294d8435fb6e27a09bf35e7f5af6f5
z5f50f8f247280d79a85e55e08df7f34f527977e69c31ac5fd05abe50e1a89378d3d543e8381ad0
z7773a44678bb74dcf7b75fc06b9318fed56ea4ca5456de421653e26c17bcd79ffa11f95fcc7427
z6a450679de68b7969d79681eba870211f4b860c708d1280dce9b55bf577e9ef194249acc71e965
z652d4f99c740eefec25005c206092fb1e3c71f7baf2696c07b5512c19813c38fdaedd2afd2a7c5
z084a64628d767bc13604d663ca3af7725ebde792d2d66963417f773de0ba93fec43ae9b8aec45e
z892a0e9212471bcd88323e4d56b0f0f4e39fcbe75a114a01eef1beaafd301e337bdd975a2f34fa
z6934ff20da68145d4c3f50de1a6415f3ed6db80e246dbf0b5045db9e108bde55af3fa02806e52a
za3759e15fadd1a7123b7a00a0ee32709a7f4492efe6a78678a54419859fe448172c8d77768f05b
z34d7a9825b4a73351a50209b1d9310a21d34c0910797961d1dba7f78142802f6c38df248034ec8
z62118f93d12a1258e6031d374c6f28bdc6b0c6b48235a2c22f9266e6db9977a0f0b3f033614f0b
zb9234a3fa29cd3d0fab9eeab67b3dddf93070f9d3977fcd4c3784c632da38e08acacde97e63a17
zd9141014357a160461be31b0cc3e1d044d1018d2d351025379d2b93ee6834cc9ff575fdd2bed9b
zfe33c142ac4b93a5f72ecfa484f75587cc96be25da2a52995666c37997b2f5852a3d21d41d583e
zb0eb22c5e014c5b5b7a68c46281fb0ec7090f67807aa77b93148f39f9e65850fc8eeae0ecb71ce
z7d875112edf5d4f6ac846c51b68e04745debe8ccd5259003d4fde8d65b0df6349e586991b81045
z41bff76aa573b5f37d165bf270d0c1fa548d16b43194d3409512cf23a9ab8387672a5075a826d9
z449b922473abc908298a44b48fc77ac29dd9e3ebb19f16a9292498e52e7245192c65a02cb1162e
z04207a4803313f9e1edf13a21f17d1a747003b35620b9b33e099f8cc41f7297f116fd234111ba9
z44a5d1523e671c2b1813472ffafe1310f853e55e065c36f08389d855b6c6bc8a30f30f5bc7bac1
z4d3e3052d9448395d3f907d9484d5ca4ccaaeb1193825e30459ea6f9272c4e05ae8ed8dc227331
zac1076079709560d2b8f18411ebbfb7bdf2707db688a920b274a93d373f7afdaf1197e4a542cfd
z38845c10b6a50972f88e85227378c90d8dfd913ef2cb7d892fb679d401cb8e481853ac2e7f53aa
zb894a661a4d99d87c08419d6c6f6bab4ed3efc3bd5ee688ab141984098afa2a063ec8766260a27
z59ee9c71aabb1bd23870412208f6a8f667e94f9a82ce94e436b22ab8155579422cdfca04a65db1
z44abe25d6ee106b10ae7a425600a636d23a1a553870970888346c4f8d067d8e643dff1b28d6cc0
z2070e39df33ed7971eb38cf03632a19dea1688d780d6ce5bd5ab85adadd1c5e22b34efb8fc6010
z0b2a5f2df47b1bad976ffab49a3285e37d02428b3f25dab345c287a6ae67372226662dcf358383
z8583972799eea126e7958b738fd0dd51f6b8c9d5798a13a51ee7ed2712705203b601256cbc7a88
z336fd0d0d7d2344c6354cff15133489d26d182ffe9db6d41a1bfc59c3d745023ba68aa357b88f2
z16e5fda8553e8a2d212bf7348560b5585a652568f4a4beb09afe3263dc90ccc5606299ad8ff938
zfa34944cf68f17135872b873465587c70ed323f21e7a1773772e8e88b08d2900576d0d6b8117dc
zb3972fc33ad360a53b45ea9e3a64d51550f2cdfc3e915da0e81b146ce854a40f0cc69758cdea7a
z5edbf880e66c7111db5cb09541ba177efda1768c5f3e5e66233368aeae74fbcae975dfed3cbbe0
zb9134d05edc6c39dc0085193a7b318966abe3c4a16b5cb3cc0305570389d65e769c0904a97ce1d
z6a6837f64f65b55bc24d5bee605409a3f4d2abffc013fc1747ece33a91a9618b4f8b33f501bf74
z8317b378092b0a678764fc0834ba2654ce41e15e2a058a791b507d1e16624ba955dea8823b92d9
zafbe4b36f68b22be9d6f4efa80f241fe00560ee48f7070b329dd348a80f0385f9a8e11a5c23fd1
z8a040653a34d27dfa0cb682632bae6e3406a3da041e6866b1b24cb7e7865cde8f2c53f160cc83d
z5332ad6943391cbce11040ceb0c81546dbccae8615097548ff3c0b79a638a4f83b8a67412de1de
z0fa0c3f4776848c95d6c1b671e1778878858f3c4531ac15b9199e73e36a79458ec832797815f22
z631825ac91e077bcb9f4c56f6799082ec39899c5d28a53b114144b2a06f999820fb094c153d08c
zc7fc105efd48f33b1a47ebc0933f35ec88218406d91b056149adeac5b559e4c733d246a7148d5f
z6a2cfb797e669196c7b4b0a5581e55ab1725d8f9a4295f2ced4506c8c4c77a4ed53197a314fb0b
z2c4e97b9fbb526e6a496b06043d2bc166302eebbeed73ac71f189ca59190cb04c27e85cb85e2ea
z2018ae9e9746c86ae099ff55c8f8131b19d43b9b0ee87dd2c455a70f05849eb400683ce8bc999b
zd8b157dc178748b12e39d1cb0b427a87ed51bb038775d7d14da67d01775336d75e8ba1baee5c43
z73d3ab59944bcfe0f9b6fef9431adaaa6fa2cfb6ed49aa35a7c37e698e2fb8b2b1376d0fbf3a90
z24d1e2303b9e7c2832f997f79eb25a2aee4ecedc40f768791b8b0ec79a1b1e958e912144fa835d
z2107a96fbc9b389bf795a3d83fc5fb0cd9916c9f85fed412c529e0ee1fa87b362df996a3e68a9a
ze821497a99d3b4ac4d33cbaec8b5282e4b9e5ab27df3a178ec2c66006464e7864f6869a2f575c6
zca4f338fce34ad7b4c872f25f7f54be497a9d5a42cea6feb068d51788ac88d7614c0b9d8d1b8df
za9eaf5b7f7d101386c904b91a04e95df219a915207f239b1b8ddcc98fc8ed100de57c3f6fff718
z5bfef20c1a496c5354d10b06de64bcaac67b2b41a5610abf61cc251754c0e5607548dd4765a44d
z66678deac5acea04d1f6a62d7797a05db5ed84eaff03a0b8f53f61d8c6d19decee41a97e283c2f
zf2688ae48779147a7433434c0136bde256183e5a144cb2534bca72c7356c64cb22513c652eb81e
zf55d2773deb53b255d26ff7889da497a4e58167b6b08e6f8ca0cd21ada877ee72b1ea2a770ef12
z8af00da4ed67598487457bece56c4d915adca2da0831315ce67b37fbce1f22808e809cffe70ecf
zd63abcbd1468c7bd0ce8b83e41ca749cd5cac9a57f4843fac26050ae1d4e56b502b933707b47aa
z0f9d81a61806c426fa5dff335d0f949243abeb5b124efd89daf9ef59782f1d2c9e43fb6cba212a
z7a04790fccbf99568ba7017fa35630b3183581046865ef5e6187ef4f6cd3dfb78052f8e5c08fae
zbdfca2bd047d8c347797dafb29d2cf65872883c66e29148c3e74e87637b6bc0f7531f4d2b83d1d
zdd31b23bff7bf42ad8b19755383855e8fe253a9a2b17983f04e1eff58dfe3c8e4052e3fa59cbc6
zfc98876a8d9757224f4883d2fcc33fd843b0ff0fcb6939e5703278bf53d6a3c05d0ba9d4cbefca
z53b273d843097926cc273ff2035b924dbed0ce33d8b51a966f1ac04429461e3f739657e8278e90
z86ba06180ca954444b3ac84fda2fa931be0d4f4cb4472ab377ec94335632f428096b1697133e4a
za84223df35cd8d290c74a0a6cfc579415b14c6224d8507739b8aaec88ead1991fcdc79e468dd73
z7d87ef9f1b8d3cfaf3625877514533116e7fac4e56119a3edaacca434fd50c1d4616b0631f5af1
z4ecce1541ac7d8025f578d37bd1f64f8e5478176ffdb5afbc98d03998f27c48146eb8f26521520
z851d490dcd710ed26c47eb12057853e144b56748a3af34c43c6b3a9f6c4ec54f21cc9707d2e8b8
z1b6925403271fceba6a71a7dcb4f6c66ca4fae4b41a2b05a413b3890983fffa3e66c50afc6b6af
zf2b68907b427f367a7bc98619ceecc4acb6b31136bcbea85b1cdcad6852df43a6b58f5ebe0d553
z6ef5891706af14f7b2fe74b3e93d5c06a3e639c8d76b3282fcf4d330f16cafe8cd76200a75abfc
z8c9df38534965dd14cfb39f35db97cac7b8caa979a6a6639b4cc03b221c791587705d567c02ce3
z1ee3f3707cdf68fac590533b5e817698f5ae8b840362eff59d23fd5857a7fd50b5b340702c650c
zdce2b016fb2c3fe31c48af0af24015a8661061094618d5e967a3318d58e0a3c71e28c7a5481045
zfd5c63aa2fa9649a040a4e57adf6ff882c9e756e2f962942c61c44e9e44baa648aa4e3a35445d3
z972b7db736ccd4cf7390c9c05064c5508eb57922ec4da99273a05de699325292e4da63018cfd88
z853baf22f61affa37e3a1f054877b724888779045d9d6448261ebab2d39889c19fa422af4c4b14
zf0b8c26eb647e3893e482c927b407e7bb94cd65673a463b61aa22997b17eaa54c03d12174b3ec3
zd8a9b9c23d0a5f7d04054d421a1f0e83a1820269649c3dffd0856c78f775d4de7d5f766f04a78c
z4c6f168b69b6ccb5b86678b48018054f48cfab4947e0c183ff1d4ab37b9fd34b37cc37c285adfd
z1751e2a9415d82693697206e57c2af9c03bebfcacfe790016bfc3baffbcd86f4d79a7c3dee2c5e
z44da5773f7f2dbe8207e1987ca760f89a53d27f803f8439d2e12a70ef3f2e7cc4ca43809a05e88
z9e6aafe8ec8c7081e39f72655d3bb1a6d2464827345f13663e00712d4519a8c08b6e4e05ab1ff3
zd45f7dd8f0248e80b7555816f6eb47d2072ecc90088087e215b6406e13824fd78c78f54da91208
zc87fccf3060293531b95c27074f63dbea6621d30ae9c198c36a10bb93e7b6cb4155ba88683e123
zb2a0af253bbdffaa34778aac6f4ffc0e9ea8625c6a276f94e9dd3d4b6b7180be1ed2ced998bbbf
zd51e6ed8b17d1f674a725b43513195e9f2ea41ef4fd6bf18a791caf9f2761f0819eb916b68030e
z04e539fc2c79f818a56187a83da89865612f843489c7cfb503448cf12a0a3581cd75e7c328acac
z9a173c4b3913f44691156742ede7b9e4f0b5cfa456383f177894d362328f73d9158ca3257677c5
zb91eabcb248104db4f9e2fe3eb8fda7497ac5b751555f8f158c2454e6fef6dfb79fc6d6e69e794
z280a7211395297df495ccbeb07230e9a4593968cf9a1212705e5c31b861759af08e27934bdba73
z6fdb79054d624e75534bafc7f41a0de33a61bdaa05b2ed1593dd630ecd683caf45e3f68a23f930
z6df9e1e2baca0b4e77613d3bd5b3fe769747c9cecff9ebaa21d6da7c651d75cd0cc98591cc86af
z1e371b4a85b5b7de4ed22a5b3fdb406571a31e0ab43fbef4496244616d808ac5188db53bfc03f4
z1a0c43a5d37aa26e5dd3176c2131b3dd653a64ba8219e303ed5cbcb22e039ea7af873ccbf2b0ca
z4bb18a32e2ef16cd4a651dcf7340a7f4d390fc8762c7d083eac84727019519474365ea27dd3879
zab287f947479255632638e2852051ac225ef91663b616f4cdba5909621a7e5b7ddee038f822d5f
z203876005ea1f99553f3632d9ee775f3e3c61c72aca5003e44de5c6ae14d693119ffa479fcd1cf
za0a73e799a6aa28a3487ebd9e63c0d9a2225853e5d0510de495d96deb1acb8267be79592b9b521
z797130f956785db3fd44c9e2c701f02bedf0bc50c2ea98e7e4f5e73c72e7b87aba3c402dbeb607
z94122720e03767d99b90cf0e36dedd4a97a730e2d622da3ef4864e22fe4a95d3f43bf3dfd8deaa
z2ac4fa2fe18d178b7f745e4291e5d3cc601ae986e694296aa493986772b8bbe63a606124cfc3e9
zb77cfadc6ceee02892115821dadb964a7d55a84aa46b1f92dd9c25ee41a7637b98eadd72ed1cb9
z11733ba9e2026a4504e757b50865f51cb4f577bfdb79d93ac13792a0e2a8342c11c81ab1afe974
z201a54ac60550be5744e44c2ede27e05c7851b8d493ae6e16d12d483a3cc134a7187ac745b8368
z28e0897da6703624fd122e19314f3622530d68d32378b3a27dbb88399e1eae79016dfc814d962c
z2166f5a2ddf215e8ff53be3fe4b36eb85bb94124d1b27f38f94d1916ea464f1dd0d750b88d490f
z2a13a19c9687b789631b8072a6c2f5da4671becc0660e687e2d29aaeccb1cb18bb9df41af7a785
zfe00479f8ba440a5490591c4a5607da5cd42efc248973dea4d9d0fdd78cc84a56cfa2347508cb7
z0dbfa2ee1a2f9953bd93c62888d37883f528dc8b526a45e36a21ed8be70d5eaf370bfaf3f5ea3b
z95e58fbdc58b2579bb6f745b2410bc02c565a1c343842d3af51a1e8b5f523968e10163cb315f22
z3b1d2230ace497e098b07f7d98e016ec7c30ba636f54c558153db7578444edb0459a457bfcf074
zf30ec4727b929df3ed4e4548b949f99438929681f689576956a2f29f7211eb6e7dd2126734b504
z3eae887d6d20047fae4d9b98a39316c1eb3dd1c58c167b55bffc6ba6ea178d21472a115f641715
zb591fe8462d80c2fd5bddca700e68a7370aa975c678470ef193d31d099c2ae4b4b443eaac277eb
z6d865bbb1cced32e31eea823e0885a0f6d0f6ec4d4bbe81b6307e01d0697de281fcfd1e4f03aee
z13964d3dd81428e9682c6f18b07eb9dc72153e18f8c0ffa00671a2d50d31bb9c797940dfaaed02
zd9731002864a1f6c80b6614b50029ea03e081f647c86bc76a3fb8c5c4869eea45b96a15f850277
ze667c2072543c6576510113edb8c78393ec377c83ccf9f4f5f81fc18c7bc4a2de434369af2da13
z43a96f9fc0654d58b7cf3feb4616ad68fcc5dd11dfd4a28d8e09cbc69e412638cbce877eb724ec
z5ad2363cc74a68f5417876ca0aeec40ed2b796284719eb2c49bf7d72662bd87cea40c6ae7d4dec
z9227fb8aad93a5db0dcd0d007ba653925cb5841233352a655083d862e351c9a99f8d3ede3aec30
z4e900eb9f7dd2dc033920b22ac85d3fe6cc1f55c3f4ceb6cae05f8dcf08475127b1708e03a55a5
z5929da8c490af897dd9308c734918b899a9dab5480d75ba9472d13f3afee2f1b614aed0069f4d0
z02fad40ccb6b83e19f20d2a66899c335431c26184d6db35ac5368a060c39865f35b6fb53925c34
z408fa4720eba18caa7fdc6c0fd3d9691cf9adc4b512139a230c3778ccdd664b40116ebcdef30df
zfd703a3d1af79abd9d22cdd84a31e1e4e36e936c9755c965534fd7938a68f34f1f9f56be752757
z6c50c0c9cfb22ee03a5203090ab3162ef5362676f0e13c63a0332cb2a7eba8821b4bf5abab9171
zc30697a289e8858f8208b7ce0778cf6881376f546d0e383cb84abab902311893dbedbe96277b6f
zd923e5f33be9bfaf450e8cd0d62803b22d616b6ca706be6f68900cd473f5361e5e1d54e72be7fa
z50872301102a596f6c429cec3ea82824a0334beae8e2020eab5f4edc26379402b77dce7d916c1c
zaadcc00ba19926a3f0fe22b69e87154c3c3156434a24cb3236a664282fb6732958f23839852a36
z50f853b97987e4aae6c5704deea7e924d017e930e11e5879d0dc489684528605025c61b59a5c59
z6732db113a2b753a32fa0549f239553559963a8d4c7ebfa8a4ab214a472984ed5f3ff79b0c8e84
z0f35b01694abdfccbb094f7d4cf92d832f23d1c4d149517204b89805800013bd18515efde59a1b
z54c59e6b1438429bfef428bbef8173a1ba4fde18dc0748c7ac3826f9ce871ac77822baabe68a5f
z8f6eda337fb226b40550f0981b68455a42fbf8d4d21506115353e2d4cb1ec18f48a4bdf8e605e1
zd085f4baca7c57b4674d5395a099250167c08cb3a702064894e2961f6bd942c04f5f58d02511ce
z3309ac203b56b53a6b9559fd45284257734f79bc2b82f28ad8cc421b4436bd855e36ac0cfc1d2e
z0558adbe33f8fe56cd5e7159ac89930a29b90949bdab45008749acb6323f1e04d54ab5caa632c5
zf48c59798afbc5770ce954d633523bb59e0678a505ee21d9e22c8fcbe868202d0615ae4a72152b
z584897b8983acae4775eb4c76b263f5538974868022b327ad898740b92eea76bb919d919074a28
zeea4ddb7e64e87e9d7fbe3a088c3fc438c84ae226ed4b75b6365d5564fe60705fcc9b369378d56
z6f3c97c0367d40ad61247a6b657ba9834ca5aee2b69c6dbe8b72455dc43bd6f68c2b13a7793d00
z8ce6fe579a3a917b168a9aa3fb9d75979f35ec7400142a33c82dd547042ce0ceae54a9bb13721e
zb2b27d55297e0e07c66b1fd2c23e6e9edf85e3f9c4c1a2e72192a59ab63d1f455482a30736a13a
zb68a40226c5443ba74e8bf34c17026ba0b50957ca74b0c9f56bedc2abd1aaad5710f8765105680
z8607c0b7c80a72f43c13b2624ca26f8660b5246b2e0778c2c0f6f63fd3c9748e47b33c0ad85ce2
z9df66a5499836001c4025ac2a4ac60407b07ab69eac109cecd81a079c321f2b235d5328c5993de
zdf31964a0f801170d023b249375d2ec7c71aefce2ba35482459823f5f8e569cf60052de71212e8
z8d8b04ec5ac3dbd12c779ec7d2f78344347c181c49c1af1d9d3fef6f458b34348b667c016a6015
z0eae7391cbd8bda0758bd6d318e37763bf393340d56d6e178bd4a9e4505ae466ea39a0ce942313
zfa4b5303e6bbd746c533e2fc575f1907866f2a2594c66f4d7710ce5bbc2e17be53a3397c8738da
z4a950c93196078cd7e6e0253c3ac4eea2186c7249278047508479d748255d6585a05b9310b4eed
zebe013e06ca23dadbc0f387f78dcff1dee873b672d5f7fe39217b7e665d9ea19a36bfe29d8c36f
z6544682bf4fe4c993e93486013279ff2c25bda816613a3b3383b9f25afb727891261887dbe934d
z9951f454cca52aa0d2e09352dd452f043689a7a470b18230143753f94bb735fdc29ec7fb3dc9fc
z4b7a43a179f9df573394be44cfe460d0ca1576f48aaa2a1581193cbc77ea4ed7221f1730059e3c
z92c20c5473587ec5d9fa05b243b9c7f98c460b4a9b699e7e102281c88025d674189a34d2b7a03d
z008a9541dc84a437ed81b1b099e5a86651297873edab5a6fa9c19cd785f40a53ffd16ce084ae8c
z487a52f7c90668ac4f85198cd92269b1c39ef315c18020440a1ee5f0d95eb8f01bce75141e1b22
z29bf05d15db95d5f68464a1660fdc80aa5a0c5552f01f9aa2836d6b7e3ebc955fae529d9e0e29c
z917dbba16c7b8907cd0f21c7f7cb7123d032594c8cc0661994947f74275ea905f5698ceb8bc686
zb7768db3a2cc50530fdd8a4af216153204ea8be8264ddfac385756c994df266a91b932e880369f
z7febc818a6a56289d9ec91223edaabb2e479a7448bd488b8f4744e057672e9a925661b5fa99c5d
zb46b766b02a6a88c1bdb7bbd4a4878e4d2c1a0a231af2d5ffbd4efbda788b988bff4786c23e52a
z76e2bd861ce015df67c4b46838f90deaa80393e52aba7a9c0578521b7b1eaa4cfa1fc0bb275f96
z76d45eac6189a40cc59f4caa1f5107abb55d97581141592606fbc130454fd53cb413689a684bd5
zb603a4570e2798b1e1a1199cd10040df956199a794f2ca76406e75272a9e151a1534176d9f3c29
zd4a4e1712bbc5c741aa36dface0b4ab90801ea98db18c5bc287b4155b3824cfec342daa97df4aa
za30328acb993106e8031558e13e5cbd4e5273fc03733b9e7473b0d54613be51d2bf005a04e85c3
zea5448feb3cf2dcb7666ebdf220d4081b91e9c9b6b1db2328ad82e1a2f54b5ac2a7ad2e5175891
zd0d06e4c57a0e51bc91a62e1be037a7c9430455bed6afb0234f7e5d19bf8833631ac644ff95932
za4580414c88be02c09a1ad06ac9bd3d44df193f0d2e6d6b47cd80820a58b9ed24d448d9b785c9e
z11680b995ac023f9fbc4228305120f9da4f38f74d1d1d88ea2bc0017086ae4d42810b5e47f70eb
z97791bfe40a6ba28afa045640dafa1e79b5680ea96b27ccff9e0af843a42169fff13aa1d4b8594
z01168b25de1b74b6e124a957b7e6ec07cabecc7fd39306d1a7cc7c62e8131aaa2b1d8c772e69f3
z4025392e2daee38b358e768a64df0658a3f90e0fe8efc58943e7fe990092d710731fa2f23656e3
zb229ac9e72549b94515e14cf2515690383fe051362f47527b616f663bdfc99755988eacd22052a
z9a775d0b72c95be35248d29efcad755597c29d6c50b47b5f2a26484b40c84fec3c49fadfa8bd6b
zfc48e64c684c383e7b547a686597c673ffbbffd117ac7d886ab73a36f0f1ab003c3fa70a807a5e
z23213f14b361a1c6d4f8e2a68c0aae82ce985d62b9f45817ac17f6b891dc2fe8936b6a13fdeef3
zf699ac8a7974b871f1d7a3743cf949825db26af9d9ca5325255b4fe3a6e01d9d899cd98f93238f
z202d59c705d4489f7c99d32349c78a8f0a4f728bb05451744bc30fdab0d5bf6f6a7bb6d047b818
z2bbc5a51926fda2fd3017e3515f147b7b8459dbc4158a95884586f25f9a14980edf6c3fee1fb28
zfba27254cb8465ec7d58dc58850c67e8ad1e83ff5cc04a1e282da46d274914e695463b2a0cad42
z5c4f7a9d541d8915d943b306477d9ad6544dc11cbd350d7c40c121b328668e794c26685108a99b
z6b9c5cae6d791ff0f0f683d7053f41e79a4d7d419eaa0df7f4790c2a859d50125ddce89ffbb303
zf2c2a974de1896a5f29ab38cd47e3377deaebb1cb74d38ce3b59311b9eca1b984e5f984485139a
z75df58d191bd38167f44f318fcfb501dded10f173f2e214fd8a4056908406b411c66ef7cc886ed
z232fdac429e911bd15c1d7b003ee3768e4a591587042472cbf757e34d1d19deed3cfd0a634e2ae
z72769daa36b2434033b3602ed7629afeb0ce7b5e768e9cddcbd2838678992b7724f1ac05616ab6
z0a3c61783f89671cbbc927ce04edf5a944387da61bfff5169995df18ef1ac12e31328a3219da47
z89192aca22d84b386d94ac20759dfac4fe65dcc5f975020abd759c0d1fa3b65d8179366e2a0cab
zee90c1321361069a8e0dadfd25c45de138c7c2d31fe04a48bb0b6853c3b4f2f30e726633f29619
z10754ae5822f192a2c238d9bc110be402893592c71da214d3140a4248c070a8fe99991bdc6d6f3
z28301e5412ba92efd49db87f15f4df411d52459f5fcf5f405f620bc0766e42b2b8692bee080ea5
zb5e85c5c6480a1b160e7490b9cf57a7d3b42de662e034994201e1b25e6a672d69cac505a0e9b39
z9fbf75f339634dbae57543a82b8b81d221ec6c4ee5b2bb77a1387cc13408e2d076e1b25985e837
z876a337ac4883b1ced19af81469af313bdb237b31afd6afc1e1f03f10d75cf4fb23f0f76e75c88
z6c6ad5b617bf3a0a882a911f1aa8f5f471bada24e8d87a2df074ba59f43fc12b1cd2c55b8b4121
zac1986cd46bff67aa484a7f4dc85ad54a98b303492d05351404a7dd7286cbb906cf7e68d3c85fd
z31a766502ea64d624fe02b54226ef189a2d26799b45f160a116da5ff544f0c4d6fbe04f643128b
z8b8c1c3cd90efc4cf54154e10ac8a2260c4041bb5bcf5bff85d50aa1ecd47fddf047f1b8e1c73f
z8850050fb5f266d3a49d7c2993f9ce1e75dd3c9b9de999057b203696605e58994a7c4d450ed6eb
z5d1496a88fb3051df80a3954c972355b90937d0d25ccd388c3cf613836c0751360441cdd893496
zd77d459ffcac19465f860a130f6a59ecd9ab68d3513f39541f05225d8bf094ee6a80d065ef09e0
z89a4cd9e32b2959d09ef381d31f9301bd83405837310b7c60fc55fcfe9d5f720184ca9a2d7861b
z50baedd6b98c8f9dbee17db4625b96133c702e7375352912f2ba17a2877fd2ddc04a28fa282ed4
z5a40a9018330ef1a9b0f5355644759effca979b9659357d748bda57f355990aee76ba543fb3de7
z9273a01580a42b1a7d83ec2919e85ea62f71e3e96501b9545536d9df93722abbedce1f7229df52
zed63724e75024500ef167008a1a215be97d88f413ef2940873438f56a37538c7306e70e826989d
zd7067eb602ca265088ab54a788842e3db1ca5cb2c12947780b4182c219d27204408c092cb9f254
z140410041993ec68238b57d89607699b710a572e68a14947a430b6bb3e5f5bbd81334ad748b271
z62f335f150f1ec1d0d4197bf87e6169a3f219f414feb0c167b07cb7653e2b86d33f240b431455c
z0f5c39dca1d3ab01126388bcff18719746f178b3023b083330120578cec894316ef0a110d607a8
zfb3178f8da1900081652f727ebe2647cfb2641d807aff592d7001024e8931b20f69030b8683e94
z624c350ae633f627ff761493f3a289be0354ab7d11851b99a19a8f2476a245462564abb574ae3a
z882f33a31399b04e7039d1153b519c9925010ce3bebe4a2ff98f0ac4cbaecdf963731de421b5a5
zecbe906acb2be56ba678d8fdc105a88883cec3bf45ead0d01f018010725396318ad836de815086
z669416da04ebc684c5a052dbbc8ff8dc0ede7e5c2f61adf06006dc3619c42131bfeefa1351b3ca
z59d91ebd382daf88c1140aa29be3d8717458470000fc8603b892ee94c0db9095dc20d92d9c9252
z760a8f4f7516225205aed5bb8c261007bee32c21c425b71b6ced8e9f35c5c682269c2efdd18e05
z1191aa8d3bb1a18a30db99b4f1374f6bbb97633901d1586fddeed6121547073ddd99dbfff87db4
z03a6532478d03d6a1cc5d10ec72d2dfd3ca1ee44c9efe642b5558c85e79e8a2e11a6ad9681e3ba
z0720a507aa48fde61d2bcc6f1452a08e62c4cfa6771caa063da537df18aae39a6d9369adff7960
zfea301ba751d922e5738c07fa82b535d713e5c6228598b3bba2c5530d42f922f2b7e8605d10439
z3862af086ea4982003dfb0a64e29627144333f88618ece77f3411e2db10195f96003475fe4e580
zea970266370664708d6f2fbfbe1e9b93bc44b415e8ca5324508ec5f1b6543ae32ef373f183f071
z8fb27f2724d60cc2e62d5bd46660062155a89370729a6e3c11925d5a4841c6cc0e7e007f90743c
zfea9406c3ab8d14e2e0f790430f87598f6fcaf9e1f855cfe0f164fca758d22887adbe03f8ed245
z04e0555c4cc547c9b74895acac838d20bc6c749298fd9950833f7f843c160f4077e9716189b059
z724d3fb87d58aa2981e2daf48c4038b21f7eb45f6f9f9555bd5b8e024f3db515dd909bef1d4a3c
z3e3bf4f1cbe447dabc8d92db395e034ecdb14c54a82035a6c6baf826b4c65c38a7e9ae073aaaec
z9160a80f64190a950b66dddf163efb5de5e9c26ffbdaedc81092a003c6fd567ea372d37650ad23
z8e1a305299517954f20b8661b89fe2f4337e2c92c803419fe5919e5555f19e2e0eff6d79fd00c1
za01d604a99fff71122566e31ca73247510a721f45214f7a8cc73a2f97803efde672e0915f631dd
z64049ea6945a6089034b54796a6fafa242a275e07490a67c1c7206237874de53d3a510849c5205
z66a6d03cc7b77b6183ac382e85618a51c48e8fc1b48fc3e2a4e0a256df87af26daa4ad65433dde
zaf8fda6fc8b8b51bcecefd51d0148db3bb8abe49b817f5e8e3bf2650ee33d0c79e382857c1b86a
zfd2a640e57ace305be3210b3bb577c2a5c7670f4494463250c528453cbd155dfdc7b93b0122a4d
z5fd9158e04049aae8241621401b83ac8ce5de9c6223f3cea03583ab3dabd92b93bf80e0a45bc00
z2f56bc6844f9ff814cfc54bdfb78de3a4bb5976076988a20aa17610c28cb4e7fd84a173e4b8db1
ze923edff1e06fe464b795ffcefa9ab5121c114126c0c8479040fc2275fb6f7fd3a03be9e30d39a
z408e796efa4b246fd86bba2bc855ab1e12e8a0aa00688eb84169b7a76470ece7097922d7ce0f70
z047bb69a466c8a5abbf113814336fc2ffe88b076ec6affe692b5db83adb5ea99163810780b1f01
zd0ee4c8538821b78a6fe1e301bb7ed1bb3db924e3b1e0e7ef3a354a34d3b20e7aa5c6168974482
zfaf236d650b1a31943ce05b2cfece310dd069d9b0e3f75791b4d331fb1140b88905bdb3cf95bed
z37cadb112c9f952d274c9dada26569afa7787d946e6747c45bc9a746abe9625b22d4edc66a34cd
z173a220b414e29eb2cabd8d0ce52b5a8e48d8fca2ae486d8a91149638dcc90dca0131565460bf4
ze03270abb6bce5df1d1af048d5b2be8cd0a2c77bd351ded730d395ccc8164d2337807c36ffdefb
z0acf5f3e0826e779045814f954bdeba4a3d1d6f8b69458b0944056c01eb0c59418aab4f058e11e
zae95c73b686d740a8bd42f6b24c8528ca067f29a99880afc7183453e8efcfe5c7da8c1ef5e8529
z9370ccb7e321f188936b8e20dd525ed07a34e7864b278675b0d7e011e5515f42ea9864f5feafc7
z02f5ebc2d6455269f2cbd915d3a839f80dc5cc11986dcdf79ab4318355e583a446a166ccdde86e
z6578cd7cfab6820b96331c13c5a2fc5b495ae1ff5a2edd1ddc113e4d63d7dc7ddaf83375c7582c
zbd24d5b1d54fdc65632bea9da55198c9b8b7fa73e2dd3d733a875a0c231fd78e56b7fbcd556852
zab2c656665b391b7001cc385252ab7f5d03d1db0b1bc52639e2a1b75549985c3bfccec023531e9
zd801c9752887a243ba58d7d88b0fd67dfd7f3320041b11bb17a47a905e0e8d539ae5ad084d4836
z87a7c038c93b54b4a0b7bb91ef2cc9c53f7fd0ffa27f2e3050c0a403479093c5ad54578134305e
zada9ea84d141ab71140f7c8a6b3869d9aebd332e4f9fb778b073a600539f5fbb9da2658d7c05a5
zc506bbd4b92178679eba57860cdce4b73c7d09c5d7e22b5d40da55c79f75cf05ea3868a7b7de45
z16121ab952d77878cf5f4b040f302b5b8db218df859bd8ed549109497809001e75c3261e1df52a
z254f4e5a8013a317b30dad37fcbb8ce872e04acd5a01e29650e6263c793fe567501568ce70672a
z898d10bafb4aec15f244220e58dfa35a665f9a1fc7fe416f98b760aac101328fd08a0f988967c5
za589021bb07f6047850673eea544bd6a6dbe3962413854620f3ced55dd54a3aea784a94d47af75
z1a84a357ebe13999963c6483e30849ca940ffb7e65f2b72c06853ca6d6a2cb5dd19e0912c79932
z1909516d07a1589ae33cd87343218d15b58a95843302ab70e5cafca24e1624a8de2fcd95d5e69b
z47e98b0454da1d24274ac4647bf585e20f4917da8862fdfcc62cc1e8aeaf552b1d108f5c4823f1
z7b476fc584d133bc90a6a304921baf97d183f6234c9d333d181d3001496927ed2ebfbfc8ac302b
zb86e4385d42948103d6b8cea34c699538eb85165df24eef61a59e54d01b92e64459e419e22ded5
zc330368fa290a56f76b1d299fb6a36817104d651f8174b29772717b9955f5022e55204f6a060be
z11009ec6535e2ecde089e20b20ebf2577ac37629290891f854dc6339eb472206802e078aa73f37
z73e1c146166edce2ad7e639fc4012b3da51a4c695def67df2f741de80d358da30efb36034f868c
z8ba80c61364cbf52a6e404822e964958f23cb62d441f48d09a47d60b88b270b8beedb7940190db
z22ca82aab49eed835b09e0e5a72f3d7bf01a69df3950eba5dec52a13033449a9b4223dd0cf49b1
zc0f3bbce9b6573676b78b3cb5cceed2c19b740a6e9e52dfa72ac4a1ab6b3623a3564d341ec70d4
z3b2cdd3f5ac928496363ef3b383f4f910666f2aa6ff45c1b7a1a87a87001e2f4b2f1ed19942c49
zafb967e3bec4c622d79c5395e05905e087721dca7e6a66f84e346112bd61053b8798dd36649cf1
zcb1442ea368a3350bec61c89b780d5c8f9efc9cc72da3979ad8e2d7cb9ccc0cb8a918c6e8c710d
zb6d0fd648656623a64be4b7b91f3023b388baedcd089f2984cb42af2ec6432c9c9c63de2fa1646
z37c7531358108eac63ac613b7a2b927283f23fc12d5943e2d73ac6af1f0168c2ae9079d2949b49
z8c72b9e4250006b7ae44c7ce846aeaf181921bd39d00c73f0cb4e37b40b99c3e37935057b1de70
z33f290ffcc0993672db7c5d432be7fc7bee87119f5abe9b0e3ceea5b6c6e5d49e29d5e0b999bc2
za94855a82fe6b34d6e7a6ef1a824ad08ea305f0ce261892dbada9a0842414d4c4ba8a6f33b6e13
z28c35b22ffb00dc8cd3a07cfa40be2d5a07de2b9796010b1a34545e74c463a86045079ca8552c0
z87b92699b23ce21b6b88be72e36261d9acaacb35b98f9a65cb10e1509b93265f0a108798608d16
z3868b437266460abf80231f1af0010257be903a7f56f559f33f9a2959b2f65e1be4630309e91a5
zcf05478d839dfd3e432f33612bc497184920cae7e32b7d1fe0a78fb490bf98a3430b39556c7baf
za3efa3210812b29187f788eb430f3695f15850594881aa3f446d61cbfcb859a7a675997ac28a9e
zc06982ebd05b0019ef987e080e80f62498997052ea8464d9b678bcc93b5dec19b3f5924d770180
z5e4f5c0c7afeba892d09d9a7ef82831854dfa2ef735f149a4fa4e6c0c173051b0076be2f070236
z4384ab8258a4499939282fca4c921e1b38375b741280523ca5af6778fbda85fd8abcf6bd615c30
zb9133075550b109642be88c9006a3a97c83dd8b08c51a16511590af206e1e18865b86dbff69294
zb8127d398f37fa307b8edb91f540f0add5324574b548a19be138ea168f60ce37a1513fd82cb7a7
z590256144e65ad9b3d81a055e4743bf783e2d9ecc55f59ebeb669b745bd3318e699bbcf9a68d1b
z2eb0fd6649ff65e8b25e5559094fc30a667e44db52a4b3e9ff584760c4e0ac50e0afcbefbf522c
z349fb1575eaffaea8c09a3d6375ae0002cffac9d96ae693a85eb91a89521ecae6842965ebd35c6
z84e7b741fbe48cea7d2c42996954672ba933aed36e8eb8fe7ffcddc2068fa8ee2f28f3637e4718
zcec4258363b8071f55ed85d134f588de1e2e16e0167260105b73f551aaf1930f1a6d2507b1fe32
za659d2ebbbd803c01d7a1e18d4980c9a6860c9bdbc554b15b77ac8563ad04d9340b25e743a0f69
z19b37c5e4158144d36d714b63b8bf3c0d3f38a0f30e3048dc4e55e5d0d5a6fa229a09d1de117b2
zc7aed9ffc1ba4966ae021961cd42a91e64adf34b8fe7577d4a1dd321aeea70387ec7c52c52679d
z700d0ed0cb5a5cdbbddc7a6f43100bb4037b5ebe7956ec404b329cc4cc334ad03564d07881c2d5
z7ee837ab6bfc53a003d7a2a1aa261f70708e19d7d4ed9137fa40dec766a8848e2142bfdc4d7564
zc4387bebf90f82e46a858622abaf31defe115c211a1d167d4d9461e8255fe8432a0bde5538adae
z1fac325c48cfe88704eb8b8e472537f0d28067855b27dc7dfdf93add029c92ff168719fe432d54
z6c42e692e5073e5e2fe0989bf216c89428911cfdd5b13b48b2648b1b7305648d64be1670031b98
z95b61c5c812c4562efcfe8707829506f66571c89fa24b15572b60a3ddc60419f644540b95e6ee0
zeef9c8ea3ec8538c91ece30cac6ba81c800e30a1e34061afddf7e3fd18b90fe959a1cef688d953
z263fc0ea43796aa34f428ce3193fcbdd507d06b3a3161ce308f0eb384eea7020a69d1f3283315a
zddd538829ccb685f0c401410f3d4249a54a32ea97a26b08afbae14f87e7a32531068a8298d9dc3
z667088666a5b023c732543b16ac79bbdc1d19f21db9baf752089737fc4471cd0d670da03abede0
zf658d0a2aa2b12e074bff3caae89184ee9df16b5ccfd79db39bf73648c98b5b090f08c96c39485
z3f128d99db77cbfa03ed3951ea08318c59943cd71e018c346321fed418adb2ae20919464c07217
z395ce95f598bf906d8290eee98a8c64e76c5f97e015d2ce27fdfda6041164b4c8cdfcef1915111
zb5365d8ac94e49b5dd51281923867463d64ae135565cdac2bd65d9b25d6fd4795ff8cf941e28e6
zd5169b8eca66429b0b6c14455890320f1f9f0b2358c91bb395ebc18814b4b54cb05da48151b273
z1405577e6d99e6a5311a85dbf1f53d85c0afcaf07ae210708aa401e98f75a2d8bb270ef818ee02
z361783a74346a37ef75f99ba1c3d80e0ca66f23e2b070ca87b0fe02194aecb07753a342054b224
zde914ba5ab235b78ea4bfd3a80e2c3b41a6b8339694b52adfec11c868c0d59ffad922d480d369e
z963ea8a1711968703432732ba7716a65cf72f73c9261527d3b420712604fc3f219b1c8006a26f1
zdb8244dedd3872cb1b874be93c323c68b04fb51baf7a3b2f752a314ef7526da91ba8210c51f196
z7f5bbc7cb7d3cde579f794becb7f74f80d2c8168fc284ff6fafdd93e5ae920d61283a010701ae7
z11e1affa04d6c444fe3f6e1e215e3a87d0f44681d8b8d44f1fba82dfe0b0bf03f717a7def2c571
zb17726fb7cbbe5ea5361c9c123b85b9cd8eb68a5e17050486e3bc87fc24f973854ff7d6d58b060
z210ff580348708a9ccd4694d33c04bfc430ed9c7ca82b5a68cba2ae34d9933e8a8be8abc467a23
z3a0a407ea3d4653428d12ce7de72e3fe22a2fbb0f4ca4c589b61dcdaaffbc28347d59a99752ddb
zce003aaf1a0a332dde8bbd448901e8c3f0568cfe1e8097a81f82c2ae100311b1635764b890b9e4
z8b07ce3f8732ae3a147027704a6a324f206c79b72b11865d3a04ce14b8d9e992a2628c71a0ec0d
z1fb80f6f0c2240bd3e5f3fedff910ac3e805f09502ce707c6e899338684cbc4e865cea161ff4ca
z14272e796e6886ab667394392aeef22851757929c57f137e9adefc190139c3312ee7da0e0bdf82
z71f01f32ff972277a40528ca567f95aefa0aa0b15e3e1d47d9657780d39fd6dfc78a7da840832b
z0719d9dfa966d2aaa36af98e81b662b158b007700eba4321b3c211d7ea766ee79464ba782c36b2
z283261ea00d7d9c39c3e700fffa8ef0d336a8339822cdfec427dcd10338612d569c7811bbabb04
z8aa253afec3603e6f87e83130a35a6e4f2e934c0b0ecb3c5c214e2b056288ddf8d7fd5e91197ba
za972645611b8a602c291b846913ccbe96bb54e5cb0511d6ffed7462afa920d4be8c24f2197e366
z46a3d7234f56b4ccc1fb06e92bd806c89e407c95ad4a6b2bd2efd1d266263848df11af4a6d03ac
ze546100a725ea3cbe77d06095c419644c214cc6e15c838ee6fe2f76d66fd88331227b2c7b6ca0c
za3209dd0603f469950af7ee0bc9666e86395ee0cc9b9f6383dbecd87e05653f6a1d796ff6b36a9
zb26ef0899f8b45a079595060e026f6e4b56aef9c2420d819312f70314a038fb20207b2f90b59f1
z5589cd0b016f81bf36e46d2895d90df619a017151db37a2ccd49caf2e18b498b59fc869ebd0128
z78926c9ed74e30ca719c13c3b1fe1c70df97958d248d532dc890a6ffa344cc2deaf3e23b4dfeca
z62104516481ac409ad58bd93ea87d3fd78d86bd8b1491cf426680a109ae23d12417f24ef9410cb
ze38f8c7da6ec075c73cb46e5f6cb395685640dabede54a902ac4bb6c64c8f21a94a78a86cdcea2
z543694ec4a7cb401f85ea2e5802feffa174409d9c893a18e342170567d330933387b92d30da091
z4af37bfe9afb0b9baec5f3d5975af4abdc85e49196eb00c9c75278a19bbb0951d06b15e511ef5f
z98c7f1618bde34647ceb880eaed7e77732add7f291c39a971415f821f2cd8fd74fa02cd24e47ba
z08de8fa502b46375263eff3872bc48fc35c82b25a3eb3332f9c9c5b814aa3d6577ef5363b34cb4
z7b5c05c213c30def42e424fe5a9de7a64d73119892496676494c60d11580caf7b5e42d8e365cc0
z2a3fd3c83c6add072e7c1459b06d8f3e257d3f086e1b7d38008b82a431547898584ae2dacf6d66
z59d0fb903dfe704da501ec3520647f98f9406d5cdce15e34e6d0a2baf331aee6013b2573a2edd3
z15ec84bf3f2ae287070593077b5190d20116dee34761b94516d4d3af008eaef320ec83d8b807bc
za8b24647b06ff9bc5182f97453341f41af4475e33dc78281beffd2ee1fa25de2f009ae1044249a
zf86a95f10985100361f23809baf7ec3f0bb3c104cfdfca7c3115043d506d4915786fe35152b746
z95c911870998f1eb12867e24161563d3e23f3a8850a9be549e421952c11f4c3bc1b23cc3df560c
z710067a3357b7f9b4e848d0cec6328055a5ab3af0f004eff8985c41160f0ba10c55974b21ae8c9
z3c5caa6d4920e68477af59999eb9584a07b505e3ce8d62d7a35b9ffc9b0c0159b409dc4016f2d8
za8d7bc615ac5afa8eeab089eaf5c392c344174d197aeb5d86fce2b517a4ea4d10813f0a656fef5
zc7e098c85253a60a4f992cb38a4b973a58bcb56b0fd43afa8fc3617c2e5f2c70556e5c09ca112f
z90b37f9d1c85a929a6ec6e271f841e7883207782d5c7b3702ce165b46e08e588391f25c2cfd0b4
z8aa8217b14239e0cb78ff737cf0faa8d529c3dc0531f6776aad37aeae585b89f6f939554ff9c96
z7f3f49ca9dece162d7f9854bf5bbd373b1d1479a73eac3f2d16bcbf4ad8f09ddcbe965357c24d9
z58820e82ad7e9c26b6f70ec0ab09238a0198576a6a32f11dbc579010ffa5dd7102ee3cb94f735c
z24eef1a654655c37f30cb387b419185bbfd6fa695bfcca8e4fb63a5cf9f1685acb74866f17caca
z7f6c3bf4f69b6ca40f9b9598175056b7266ab082aa52012bce77829ed0e3c54a4ea719e4564373
zcc3f499010135eaae1e0efc856a03b682f50cd47ea3f144726560467e115219e89b0a40128c2c9
z7a467b22c00fcf631415f2a15e5e8da88e467d0e3f6083b93041baa8738d784d6cfad3dbedc019
z57007c15d30ae02e9b8cd6f9fa16668de93307fb9d63f856ebc3fb838ed4018f3b0524e62cf8ce
z40d33c76fdb9b80b2eeace4b0cb66584a2e7cc0fe159807d950e408b8b435eb9d19a3813588216
z4dec0a7185a127871125d32641971ba1880ef76d926f9f4e1dd7779740fb1447e75fdb7a3e988e
zbf1207f143b9c83f9da295ac51d6d115c6f4fb300bcf0b76d1867b348a67291082d1f2bb83c51e
z6f67b2159af8219960059e82a73c2bcb2e013d61cae9f31b9ab74428218a5211284993e4096c28
z6b53a934a0b48c80eb8eb81e9f7259cb9b8639315d823e7441de11c12533a2611bb76a316c7a98
z79141c5aa3102534e57a123b6bf65d2d5466eec8f18c18130fe5db50d35b4110efa3774bc1a8b6
z6e6e23a78d45015f40c0753841c63cbd5f647adbe19dc1a499d99bb0eb2b41c0cea4db72cdac51
z3a092173d1c6fb6370c8dc0f9ad4ecd301652ce87edb6301f9eb6ad1f4a46c951f1ef073e8d6c7
z8b114e1b0dcb3da1fdcc6cf075a651b6bcbb7e582fc2b80a29c8f95b326751d9b7e8d4b9f17b48
zf6338ffd7cdd6cc19da7a015e4c8ffc091159f044dd7777afea932944659e727ff94fc91e25a11
zf29551dd0a2caecbe2f289d7b5fecf970bbcf52587b46cbf90e8e541b3d084f5a61e8d07c694df
z0c837dbed38998b3156e610818f743c3839b64f43a22e54b5f527fd7b1ce759754ad7b89651f71
z19d200cce07f4b2b322d64a254fd34416c5ac57b0184634620033e80e73c4d4e9e794bfd1ac01d
za55fd78c87a43a165289bcc06e1b09bd2ca654807d6898ddec667744068c162b72ee3426c5131f
zc71f121ef6ec2afaf63056d42f1cf48b985cb118eaa8027f48deb0bd40407cf53460f5ce862230
z2b0d27e0d4c7a7b002053b00b26b1c680990e58c26fea665ac3357bfb5f84668916f647e9ddb25
z7b0c384488999e391d0aec2e1791841502d224a0325bf901ebcd4b9ca933e2640719825eecda66
za4708e9b9b9c7311808b02831585e37c46c132bf3d05ab9bcbb1be8c841f103f7169d7a8d309f1
zaa580212028c21c1a1e0b9f2d2adb86bca54b203e46df01f46feb659180ae00053f15ef91680c6
z0046e255710d1e821b08dd69976f9d67ff2d77eab341c02a037a2524dd8b1a880520a23209cc07
z040bc34f07f042e467cbef37ea9f07b72d5019887b87b237883c35ef0966313fdc97800fe4eb54
z24aa334b8061cff5ebc39953248d05afb2eff0940e9d051358f1f3fae18730a4e664199086d6e2
z8ed025c917f0982507f50dd1956267ce239aeb103286f2c10de953e1af0cbf27ff983e728ae949
zcda6c5bd9be5d3db3a006ac61e2c5ca724401e8bb25d23b0160ea3830dca1dbce6633ffe037429
z5e45830631c7dade99525375ccb169f206f5d3bdc267c164115cdb0eba8dfb7f3840df52897ceb
z2a1fafc87f57b7097432172076707d837dcfddd6118b6f5c39e97df0497c0fa78a213bd557bea9
zddc2671ed6019fef66482eab709bbe6e5e6061eeee90591836a2becf8cfb07b9086d878752c116
z8e1150ccf735152cd34399db4be420db
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_spi4_2_rx_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
