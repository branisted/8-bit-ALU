`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026201628cee5aae21fb892db766c4
zb5b1406e11aebfd6dfacc9da5ec03b70c276807a3eb15e28ec7ab1dddec42388b9424ea285623a
z248195c9f894b36317ca6e59c86f11031163f5f5bfdba36b10b435d36514783bc1c6e60eaff7f9
za2b8eba90f8fd9a9cd7c932ce34efca1757e6b2718aa68644ba032b1bdd74efc688b935cf38d81
zb1f311df3e5b8e4d46dbf459c824f309500192485674c175e61de609f1c94488da73614dd500c3
z680b7fbf510ef6c68927870992ed3376661d943d2a929d90faac51228c485cc4f90c0eee6be4a2
zce41f6565994f8c457ad3f059f0f75d13b595288a756e41a6033f636eea17dcdf0844c8e225d45
z55436586fc78f7c2c04155001676fa3f49b24d3beb3584c63daa43ed80ce015162ba22d33c9763
zba142d3955797e70f433f00a9ae14f9d776b76291d31153dd23eef201b698c8aa3a640b228a83f
z18eedf1d37da4b3680484605b10d0117d140a2fec482eb066a6b3e23701cd7a6c894de14b6b8d3
zb677e1f9bb4ca13228f369d9dddf6dbcd0b16acd11693c47e9f6c7357a4c391b34dad72e54c342
z6c4420cdc072d7580bc0e30a06dc17086f4da8431bf9c0272ccbac2389d86bf9ee28c7b319f937
z1b9d9426376c8955be3bfcf3aea1ddb252af3a0c6bbfd12a0c62f959b5f0739a7a8583034a7c89
zbf08a54c5a6a0ea9a33d5a67901c83473c176de06446bcac2486781935612bcbd39c561d12cd4f
zdc33270829443dc3cdaf8a7f6773058b1b03e073d5e2bb6faba53bc8f9b8860d92b24de0ec1505
z0cc0a215623d6029afc16c5d59cd085796ecab6ec90a709944d61cf60144977025609850f177f0
zbddc58fcf759603cb33727c802cced0874f2bb0d14f3435b7ee8b1a94b4ed366d39309710bba2c
z7b3aa24358b1cc35ff35c4739e2ff8ebe589fc18de7a3baefa6733ac3bb9a27d2f8935ffbfb69a
zc8ce9350d9caa3bcd5cfc85f55398f89cd4bb8df5da81d3917bdf8ca19247333308c8836cdfb81
z8efdcde75b57b442fbf0fcaa0c28e46a094a3f87e8c19c87b248cbf4452f9be38b939ec7d1b2cb
zcdf6f683148aebf2ec21795d29e484a0c2b9bc8cae9cfbebb9c18a525cfa743c170e7ccdb3335e
zf88753485831a82eb7eb7199222adddeff77b24309d204551af5c2be4de52aa49bcf7bceaa224c
ze9f6ba25f246221d581ef3476c31dc53f33a476ed160d1b8800c221ee04e30b5a4c89df248b4d4
z44b396e2e312bd35fd6e1f929b78bc3c029e50b8d141ee478485a87b7460da22ef0fab8e9ce177
ze9b8eda826b1a7b272fa489862a42a9d33e6983056a3c547aaee8202a704621e0ed1bf52b966d5
zb6cee30d888bc366da0fce8ae691df2a9061f88b7d397e7b0b3e6915da859fe915ee846f3607f9
zc9ed869b60213eba346e8b2542a7ae6ea818a1ac43baf4d3d32bd18a7fa8a86fc78a096ce4eb6a
z4704d56bf9a83343981ec9b43bcebf371fb54384ef934591e0363f6647d75464b398a34624706d
z0281b1c6453b5c46a89da6c62f671e2962f797b28b567789a14643e3c5151097e2fef776df5abb
z84ecf9c8a4afa4a7511b2adef0d6cae2882b0f7c599981dfae18a4ef35c1f3752abeb953847756
zddf15cd7b6e18f0dd6dd0426e652cd511acd2c55bf6bcefccc18d85694c2f614692874faba28e9
zb2d30c9dea3341ce9fdaa1ae5dc3881f1bcffcc3f41550863de7a7f01835b94fd71d35ba615cf0
z912e65961a2ff2b3ded95f89a06dea004ee0b6abcaf0339e9f9ae09ccbd546abce7b6571bdae63
z7f74c896e8d112a88d0ee07de3b43a36027cbb5d841295384154f9db2fb82661a52d69bfe3d278
z779db7ad53744158d84d6353f6a3f609a46702d2076d15eb6241bcc200cdfe1d1fd2be41512f36
z75adbb8eb3973b4407e22724396e09e851a3a12cdb55b3f52003272d793f06dc43a7d1928f9990
zd7c38f3b1fc63f1ada5f8e94c9260cf85322b83324d56cd542f3573d50d9dc9381a498874cb5c2
z26b67841a2fccce1ab7f72e0085c0d39b5741f6704a2b8e8cc39cc743f4a76755a0e45268aa9e0
zd172e0859ceede7da8dfe8d3c84c5b5f927880c1a54adeb6dddd9491f5513ab106805cedcbb3b0
zf755b3a658a6a00ab5d1b5c04c0078bd4120fafc726552b7fe807cb83bf7968f35e38d9afc829e
z2a90e3fed4ab6051d3c7a0e4a5d3068011b28b43d542cad7e49f1fb3b630e6456b343f0ee64693
z78e5c382a44f47f242fe659964e16e4bb5b913a7140b286e31c8a3005ec65ecb9d4b693c950337
z680ffbd21656a7135d73638e4b43d7b5dbeb1d9a50578b0e1a658b57076e607fcfdf85d214ef38
za657f0e6ca0abc091c7110131161c781e79b4da52869349018f640bb41eacfa12dd2491a776912
z81f9768a14e4bb37c6c8b4a8dc433177b58acf0cceb58a7dbc30733a060b7f4bc3877385031156
z7cd6612412c18cff80fa52315287dfb6ccba56ac17e8c78276e7b4d9068a3c8ecf4d1089577091
zff679968c60b0f1889eda96aa27a71c5b4ea6df33ab9aa80892a749f44865f81635414b793f717
zacac417323dcf1df989255ae5a7f1b0463dd026335c47ba6e9cb84976cca75101e0cb3f03e1531
z3f1e360d930b874c5ec0debcf4633731d27146eb09696b8e2e445a48becd70d0bb42dc857bd73b
z225a8cceefd715a799fd6105095a853d74e879bdb5c565c4f270d5ab1102ca291b4fbf3d9010ec
za479eb0c8e2ef231f74330af51e0d99498740b63dde5df270c9b9763de5ababf6961048b1b1576
z7146e8427fa1e97d53ff3fd8f22883a8ec89dcb32f9079a826349f667eecc9fd9713c23d56f08f
zdf681e6d6ff42b1c33e2ad3b36fde509379742eb8151f2d07d5a4b734d029e6dd3ddf5a8b8e452
zc28c9670ce207e355628aca50aad18f2be98f52609d46e9339466f846ea4f68bd7793428e9ba16
z53695a8d041f6da10327bc8e025120526f4d53eb165c3d74707d5c01c0da909169c06a12b604ee
z17e01b38de62d1c688493774ce1567a1353ec9245c0e8362a8d56aafcc3b51a023342b686458ca
z490703f6be4a820cd56c14e5c7af4d8bdcf36a95a28ba3f2f45a2a0e1e068e9655b209b75b49d9
z037edf3fcfdf0aa96a8c2f51f94cebb84271861f59132f9aef31ca0008b58c10831c6fbcf78935
zb5642b6969421d2a1ad6fd39127191f94c5b552ae009c54d234106a0593aa8365f86fb5e3ca16b
zd5430d2c27bc3073f21029b4ee572f7188cf958cd766a147d449218a60b95d258454bb26a694d4
z208a1937286b2dda4a9654cbf84765ff2d60b2ac7632ababa1f5d84e5e8621ff1b98ab804b1dbc
z0d92b1b985bfbee615bedcfd7839ad2555c7909645bc43879a0126a4cd13918d74610f58fc0074
z7aa5f97778b55e99bc23fb51454dc4f52319096bd8259be6126e1f3579f371195dfc0b26281117
z0dfa76240aad80aca1cb9e7509a85ab055dee348b4505211eaa598d1eb2c0ff2931a154757ecb8
z0cf35ef82076c66ff55957b2afbf5dda9a78d1ab7e4cf549766da49263ca028b9aff477c1be73a
zdb2c18668b9938f806c2465dfa821e2759a07e9665a8da380c2a51d169018a2cea24caadff27d4
z217985fb07cab81c651dc5521e37d83ddd16723527b6a03b23607a3a4a1774898d7bd01e6727f9
zbd443b102e770f76d9c2471bb76132e8f4c660d7d905d4ae1b13ea2cab0a05eea20622ffd48dc8
za7d5e75b41c9d33dc368fba8e7bf4701221093a47a72c14d6a9dfe7ee3c0dfef80c4e4756768f0
z5fc4633de26dbb0f0237dc08f716421564362f6a4d6aa925fd205e2b4e82f2414f48c056db5b78
z51c54235a495fc827b00b9b5348ff2847aec1241f5115fa32a7608489a4316b323c75f84111122
zae2a61192f279950fafb983baf16dddefd493f957bccec8066e9676ecc5ca8291c2a2c5cbd01e0
z91ee4c80c9c25fc51a031fefe39ece2f9ba49acd5f05d268a361ebb00546450c882355a88098d2
z891128c4ea305dedb0ad248aade730a5033bc44f318ba12c03982c1b1bb04d7578fec51607c042
z54681bfceb780a256d1c4570f48979d7d9117ed63bf827d065f1408382ec838abf030e2c7d1bc9
z6c804d129273627f8c7c9bbd68ac1d6ee87bfedaceb491c8dbf632985dd71d1ff96e234bdcc4b8
za4b2e52e6bcb12b5378f583e30a36efbee530b44d0a13fac53c8c7ea7830447e4ef6d669b1d916
z04b59c94369adbe4b97ad522666f686c4d1930cc15ee746b07e17e45aa09c3b24b5865c8a6f0d2
z905a4067df732e63ad2ab0469618942da830cc6e620c439ddbe61a07e076c8efebf40025c13b08
z81351d98a39033450a8667b071d4347cbdaf051a216083666d77f5a767568b54441a5d7d6e4a47
z9094a134b2aa92722e31bcb00463b6005994c277bef4747b00f11b388c2782ba10482e27f9b502
zdbecdfd12c20b9914fb91b5e8025a3ce40595320d460f8a325e06488b7b68638a1c37590fe88be
zfedc344e22b7ed97bf6b10e865f2a00e49f0974bcc9b508659d3f737d222bef93db484827a1692
z3fceded9639614544138d97131d6cf0a5d509373e581ab6a9ef954a65a90c554b08e907073b4cf
z030049c14dd3bab470883e3deb4704fec6a458a1d3c7d2cbfd6d7e095da7e9a1289a06150d635e
zeafcef4513c764d942ecf06563f3181c03d455ec5ac1c15109f5189037accf8fdd8fafe41a14c3
zb0109df97e927a0a0445410206fb1abf61881a779782504e67ebbb69e5c2790c8a1071a74c0d18
z682848aadfdb3f8000ddad3c7720d08f39314e7e954f4d1e6716129d6897f0a85e6b9d7a0487ab
zf03a8012a665a4fe3c479e479b75e5943f24029f74b5387d2b76b60c9eaac53a647903e978eca3
z0e5b06804626e8548333970ec9fbb6ea0f5d92017b5eba7c14f641f8c12a6757e31ec8bf7aba9d
z8d55f87a9f6899ab63deb97d231e55a161e31e3e4dd5f31f730b50db4326a2b685053780872e74
z317e0049c9e1f579bdcbb37ddcbdd0dbe440903a217f22e515c047c0addbc297f7723b97970026
z591cbc08c59ccaf275cb3766e43828306231f820f1219d174c2df01893af2c432181d7fba85df5
z002e25878eeaecba42eb7c72d9a18540991f91922e99cb34487dd5509c0732e4f15b2433504f6a
z15f2656f855a95617dbd344cf4444341d89bc0353c4a481ed9129cd1b41c1efa9ac4b487a5d296
z6b3e8bbe4797bef64b92a76d369be81c99ccbb25a0835a6bd898d2578d7527eb9bd4f9cf3e5856
zc2d0343e0b8aa787c4aa07fa7a02144af00192856cf86a83ebb87873c7a9cc831e1730f8b0dd85
z419bc03089e92e8e5609aebaf2d95ca5d9f3d94f2519e0b8d116159a11f9261ec8a83e8f293186
z0b512e513f75cffc2671463d6f9d060f63dd481e311eccd58548507291ba55f67af0027ee2dbdf
zbc29fe19745cc65f463b22221e369c0b75ee822f2c8969f24c52f2bd93f3561c6d1845c2d8800c
z6b9c4ddc8c5db61875aeb8fc0ad53b53ab77e87856f2854c5fad8f331d68d3533189b6e7441287
zbd7c1fe0e1fa655bf67732a855befe562ebdb54a2720420719a31650809b98dc63126e8a6b1656
z6a4946214fa172209328bc78d220b55729af35348e45b62b75fb14c30b2c9767800ea1fe990bbc
z22810e258a75d231963aff2c614dba704652ce753ac6a3b6a85f9ff1ac626548eca623afaa203c
z3c4ea4ba1985c2c8db39ca0ba3eb9a4459ddf37bf695e9805457d047e7acd84df454a40235a818
z0de2ec4db7092611cead6a778fd0848bb637503c7884503368446f17b40c93fb388f400fa16915
zdeb15a6815a89e5666a2a13e1e6ec0251301e0614aa5045fc3585b83c66dc0bb8333906cd8d5ca
zb262a696f7daa98e2e88de33934150108a79694e2b1d8d99403c13953eb3460a4aab3068052d6c
z255b56fa0dd726f7fdc8dbe25894eb7b5952f1c6d447fcd4ad345f6a02e7b26228a7df46777a67
z6aa7620ab8e4440c6a32aae4b85a3a6f5b76eaa942db3754cb98f924d4656ae44734bde9849b25
z9dcada7ee371ba9cae79458a213d451640be39cc51dd0e701b8e710caa11d99591535c2c50192a
z0871ac0aa00197ba9b1d6ffab8ef981a798f9f6fff0ba8a674eda5a0f7da9013e7d152eecfa4f7
za11291bbf6324d81b459d652806fe92956363f4f06c2bb5db078886b1316ead31d0ee1a92fca6b
zb08f6dad816c93cf3b11e59e1fd263cc64deb8e24d7d5409a22c9cecaa2765be9b77d711451063
zc2c8c5fc576db97e617539a772ae1407b06f4f2a403ed025af470fdf3e623bc9123970ea6eef38
z3d1315c98829b6da1a8ec8bbe4b23b75b61e6e489c5d67e61656ebbb5ec7fca625050036ce6b21
zea2896a8c3ed7f349cf2b5152cb2fc143fecd3cfa2740275bb5d490dac0c6e2bf142d311163416
zd2aec332aa8ea12811dcb2a207d507fff1eee0e950a17f09ac99008181441526e62171b5aef6d9
zbca48372bf78d9554cefc387db9644cb6dc53cd0f77f6926de110120354c842fae80569987b0cf
z57090e978a8ea4162e7d030050a15a24c1b918aa7f75dd58eeb8eb163a96eb89707189a76b667f
z45042c9114944e636f113d4af58340fc56573b534fb4f26bdc813060a1fc7026d3d7f79d3ae205
z5efd32c454fd1f5a87a3f129ce8d45b2432605dd02d2b934587f76cc8b653bc911b220206f8faf
z0d577f31421479fa9c6f50fcfa144101375b7854606587bc2697a7d320ec67028716d0e5a63c01
ze868e654b032ae1d51e11ad95dd7c5f212db34ba163e8420df22bba8b366e7af488e53ab647019
zaa0d6967972d386392f39980b8afa6278974173186434cf7b2a0b835942685585602195606493f
z12365eb16f988cfbc1bbcd0011e5a5b4c78cae3ca26dd575f7b3bf157679cc53cff3714fbbd31e
z930d1713fba663bcef8373f715509e7023507620090cd82667c251be19698ba222503e4f41e3de
z1e672dd737d7acedef5a3a398ece469373e176dcc69c60a57d0013d2673fc0d37762ea422af61f
z3f2fca06a985f74be143f38fbe42ab3d7d0b065c712d0159db2dbc54735c279f256af47171cdb8
zf3f3d2430726b4b212236db740f39157457637b96d0861ac6b7c872b2247edb3545339e32bf391
zd2e386255697d21f9ed26e470960f14b7284e616dc59a1cdf5acbb60e3b1bcf99b831a43f1901b
zab7fe74975498052861100efd431cd38bdd100bcfab508601f22849cbb6c17432ef80dcbae3ab3
z30bd3d5dd3a13d29815fc4eb9b49003a0b07f03cdf6a08e85d638f89af21d40af440a49697a341
z48117fc8347fe2e655a0a2cf4741087ddd93a0acfc29074e6271914ac48eb499cf53683e0b9f22
z9e35f2ffcaed038aa37f06be2b8261283af97bfaaac64770e9e65ad072c400f5cfa39768c5a911
zfcaa8cdb6a4901a1e6829b7e83e843ece935a391a02d18eaa047a7beae722a4564bd8b33c731d2
z3c7eee3eee2f2e2f73a6505fe1208192851d7471d22b003762d15bf968c38a4a5ba4aee2986c08
z66e3346d954318abbc9ee19758082b0108e2771dd6ca341be21950aa7d4ea382552cd5951db950
z1e40712545eead742a37cd97504c1ab9a210ac8ea770c86e4794204aa014fc79001a1e8625a6c6
z51267f5c7e0a85c3f7e9d0e0ce16df35afd9f135f95e5281b1c1eebbd89dcfb6dd32af05848fb2
zf56badf674111ef82f7a8ab34d23b18aee1c73b54c120a71944736b74f3ce96a4f5d9cab723cb1
z3818793459ddb648d3eac9076558d93ed78b54b10aa61d7c529008d62600f2c971afc8582fd567
zadb2583863fb31e12531f83f901753eebabcfd5f2cf0ef217c7c74081ac13e7975f2ab53adad30
z9d8bbf677c1be67a02571a484b620edc8e4b81895767478396c22b5dde5930347a966a458e0971
z4ce4ddbb9c08fc753335c0dc975c1ff431bdf905d27c8da17a691c4f2e927553fe1c9c3fd9348e
z5e5d402c3bce8d96d068acc4e3a10ec92f3e1291f30e23b7485e6e7492bc87db645a8959d66918
z6653bda2073e9b502f9a9b2637f3b08d063764ebc959f0e526bf237e5307dc30e274ed4f2a3ae4
z8cc11e065b8876630926224630fd6ff79fbe4f207083001e94e126ea0dbb9afec66ff354faf461
z2274fa0641ff0e0d769aa61028f01cf9ac019a4a0e974627a00e29002130326c5f269468e6490d
zada2ac4e9432418e4c0d7797a0ce072f4a8c920c5d492fd4402ad0c142b6d342f89a9db247aa7e
z859bc80cebaa371bb2ff54f96a70879195de7bc094e2f2d594bef2c9593a41f2886631de91af60
z13e3365773c369cd2dfb0d73c9620bfc1fbe0d1208ceb23bc73a765232426639de914efb7dcb32
z83944bff885548239568b5032cd11e307ad32210be5cfaf2dab3bc4614b222c9a40f5b94ccccb4
z917356fe4f0aaa39cf7d1edff3a1a15262f7bd113567c226ded7a6c3f5b13be6f4a39bf830b4c7
z3a005016e121083206d16b9d7507dea7c6f673d7c6ad050c09238fc95aa6875837a00ff2921cad
za3c9b4ca5f92f0e7bc41fb92eb54be03438bb5c38fc006a2ae5cea382bbbddefc48192ffa48e37
z51017a4c5421c540eb655fd4e49e6941686dc830a8169b2f121e1337dc71576d98bf962db904b2
zf4ee531a828a5c4475243c705753a4e8fbfc147566d77a6165802e688c550c8275ce43288463ca
ze4193680ac1d76fea1c1ece44fd4970b1867ee4e64540aa989e4a079409790895fd1e8de98bf05
z73d7f43e622332c8d57f7053fbc88796ee6f64f5e261445c0a0ed839227ebc25c9150ea16f9cec
z548dd280549a634068051177d34e91a773bb5624076a1e215ead9e80319f01cc68b59df071cd97
zd677a06ca9623317bc01797597a6aae828c508ba366cf8d634d330bc99a06ae11d88069591f6a4
zb7878f678148855d4cd50f466d20a5d14d9551581150a72f4e1a3da6413df43c5df746dd467fb8
z14c7ed3e2dec400e24cb1a64ada9f5e42634ee86212c7d14d57ca71f7e4712ae2d0ab05c006f91
za1d0f66ed7c438a4cdff6fbf3d69e97b55cd4a8e4789fd36e6f60e384a10701c76d3f104b3a019
z944b166941f14f471ce2eab59ccdfdf5761fd43219d45766ead1af0139d52a661a337e98ea0d0e
zb66ac748c4dd33723c78064fc68a65682b3d7082a4dbb82dec48940d59dad82d31ec9d99a2e568
z7da3c001791010efee0d92fb8e77c7abc200c56c48fe7306a4bdffa973e87bd06d7aa33a65668d
z4785c28dd5a6a8bf413f9bd32792c9151b784075f0122820b3c09b3fdde9e0819805626387de80
z410bfd3eef45b787602b38d360d898d7647777e8d375fe58161370305d2e70efbe7f4245f01d3b
z92404e66c46ccbcc885de2a2b859aa25675482acddce4ba83e58ec054c2a78820461eb0150f284
z6ed746f53cf6c645b10cf0ea35523842b7da2f88740374a95bfe9a500f40f0c5441ad44f13a25a
z639bf515efb1b1f8e6eccc19f41d47dc778c6db430d53fd673a64364dde42d498d9a984fefeddb
z04b77fad3c2e6895a861e5620752a97cb8ef485827d9e9d9f7b76c155cd4d286eaac311f365faa
z3c63fe890ab560ab29fefc90cbafed9cff798aae52238a956fd70acff1ab67a95d492c4fb2bf7c
z257036ed07bcf50c355eb978c9532e473fc11a955770516011beaa256e798f8da138530673db24
z1a9b07c31d4bd7adda99a429c5c6a64904b5fe5873f6137b1e87cfe2a9e6cb96bec3ed8b8cb116
z9468886267f28b6cfe6808d89853207d5eb1d2340044266e2e17769371778829f6e5f7111be7fd
z56feb9379553e8d31269b668d4b78e395e56971d9fdf09bccfb402ef60fa6407123fd42813fc27
z2b1b9f2064269b98d8fdc328b2fa010576c50ccaf33c5e0e7dc34cb1fd7a46f41cba27c2c6e934
z03e742cbd7d968f9f1c500b660ada8fa4a8b404a6e171bfe30bf0d3dcdc2f9fe5e7a47febb45f0
za9dab35de05ec5053abe8a9b414e81715edd0e94557a06c67cc801ae9550d972d2974aec166b3f
zc70d8e94bc24ccf71417888c30e5a4ffcf9fdbd7b156c8c1aa0a6ede4677cf7d820d49a731d312
z96b9a803c2067e2a929b5f650f3904205790ca7b8f221a9dd2ef1f7ef4779b3e9411d115b5141c
za17a60ee7f8e99a3e738e0402b7c369133de3a14ab6b28255e625127b62c1e296896cac846074b
z2221cffac2b719fc498e37b69ee066fbe8c0e89fe889fc95600a6df61884d11e26194621653273
z2de70974737600a9750b057163748c21e0c6ff59517f8a63b029c94e10c6a0e850cffb96c1e7e2
z72098bd05448e409e49983e885e8d693b87220a78801fa325b288bcfc383da1f878ec887bbee9e
zc7ff4f4541487967e3bb0e7b7ddf457b5d988c99eb680624cd490d593828e4596b4ff0e8d461b2
za18e844f59a665bd789069f3d5569e849e8c2e5ce858d0942d51620a976c1aad4f55a3cade9432
z54e47e772f290677397c9b1ce2b1dac56539e703194d511920ea32006297ffe1126a25d93e231b
z6de39b24fa25a98660ece01f88c7e77f9828b2c3dad52048c728dececae37d0764c1dc82e44215
zddaa89d1d5a32576afc025f79906994b676c9700c71464d1e3ef4cf309b730d2856fad8d0adb2d
zd214259850d129da9729392c9be5fe0ac9de4cec7cf403b35a25af67045c70258cb12e4110ead5
zd680118310b775664239dd591405e6fffb13eec077d1131c6fac663331b0f45cae2c7eb6bbd266
zd0f00ccd6106bf12fbb2a60fcc1ccd4a0dd0689788a3e94ca556c3e10e8757b9e8ce5678cad89e
z91162badd484e982acd9df07b47c70c583ee2069677bc4def6fc4a7150f855f924ad6f1dd502a9
z96c782ea8bf1094e486ca2d23ba993031c5a14f50db3a7e73ede199d887fc4f58daa6fcf1a75a4
z8b9f65d4fbebd966d3192e8573cd9c355099dd1be557eb3fb60272a6b98451339427628716432e
zb2bb3f002fbe21443336bd8edef238996d88de13134c6745c64c821b6dbfac7bfc2f289c8503d0
zdea4de00308764db34dd2e9c6b038102b0b28efa88130a40a91e6e1f210c3fa9721b137300231d
z05cb4c2d8ada9960d218fda20db01527da09b812ca94e69375afeebd206dbb8655ee1e0eefabff
z5b9ca40884b7fa2989ca9182b887d171eadad048b9eceddf97525d3fd684f229e4daddc64fd161
za1f633b497f1352cf05a0ef1dc98ffed80a3e905be39812d374dfddc63b9761149d133fa5b2b29
z9dca4d8fc7b89f83364898269c68baa2e05748c375db46a8e0cb8a972e7ed8920bf55b2ac716a9
z985b67b0cd73a95998f48d5edec4062fa47effc478addb4a83e1377c25e760fce7933b3c9069c1
zfb7a02a52db756eccfb9e6880c45a5775a86c04f29ff763713de8c578d78d4f13ce382d7079d04
z166a7c70e08a46a71d2d65fe2a5751bbc6fc78077c846b20ee4655f90dcc0512f08dcbeacbe5bd
z994b788cec543ca8fca3105a963e6e64aaba9e4270c6d9b2cfeefb2eaf737ef898bd5b93a1f47f
z667d507287ecc361506211f5dfd94a46009c4dae10ab68fd1f47d144ec0f241fe36b67491db9d5
zb6103e2f78e7c1b08497d1064a529b14efe120cbf621671ce45057d8bacdef1b584831eb21ff53
zb38e37a526b82ff9479877ca95916735fd1b0b0301db3d4f3682f8ea3a5c1ad14fda3f487f27fa
zcf294c2144220d9e81a08a8266574b6f556dcb8585cfa3ab6c17df226a89d6801b9a6bf89aa68a
z4f26cd8b9f2ce177080f4f678bdde299b317c9ffe7482f97c55e26a3c29bedde417411eecc45d8
z353d2c361576c03ac83d521e9002043b89a354f2777aedbcf1d2c48b2d6ebc35ffcad774b4242d
z06a2889b119620de8373e74c63fb8d5f7e937e289d71d8820af96878e403aa6c1003e329fb4f31
z4116118e497de189b5786ba39bc045a24eeee038747f4d58d130faba4e3d59206f90cc178ded98
z50ac0683307d2ca72da2b300888b400f0bca9216c856610ae9ed07e5315246290bc3056ee9944b
zdc31d3ff78b7d49a34df104211c00941641fbc57cb7e6ce6718fdd31a5402302611b33008c3001
z70e33ec07f3cbd023ced916934751cea259188821a8694bc74d33104e3afebda10c7955e95105b
z1bf9791127857d20a7886f255b647f9c7df88a844b7712d874eb9a9e5f412f10848f2cee283df1
z0b878ee0fc50511b83f8bce1c6dbbe0688637fdcc04c098359cd7f4cbd684dc699e25d49dce4b6
ze305409f839e958d9932a5aa3dc66a99d71c5f52eadb188f76f8ee30e6c79916d072ff4c1363e5
zb64b81ad2e4d10edc5982309f4299a0f0edc9b70c69b0b69856b72fa5dfd45edb0ad1d7637b36e
z896f693681003bf8b9e46c00a97206de5c23be78152e65c4558c3c33c1eeb7e389198266e69c81
z33622707767d26d00fb8403afe1c7a5956ca5e8c72f71ae50d9ceb8595b4186c4885b28b548bf1
ze8249ab6febc3a139a4b01dfc7c050bbd30b14051713ea50f1e7924ce4c440527265e7580900b6
za8f589aac339dea7ffcf476b8a0dfbe565c59fbb947863b35dd407cadba3a598fa9ca7faeacf60
zb0c82d1eb981a845ad5f1a158d5f5c48b46c7f8e5750142dcfb395c978f4e96656eda37525cd0a
z730a32dbce2057e3b2226853b5842734007fc0ee92e62ec6df3f19c24b71b18b1cca9512af87ff
zf50f1acaf1ccd8e08ee6841e5ec82126d632c42f89402d58dbef02bc577eb2a642a3f807e3dc08
z9c68213b2a16504a8e67175f092d8d0c012dd2df1a4dc391ef38b9cb2b72f64e79184da24402df
z00f32e28583ea06136fa69d41241516601bc46a9d11e3d4df175859d445881dee6ef2df9dc38e3
zcf267e7ad21c2e0084f55be36cc30125940cfd97a50fc86fca97191ddad88d63007d34918ee7f2
z4b1cf0d46335302a267ffd59e54704e1caee9396ea1e7eac2ffd5f2f9a8c031ccb248a2b055ea0
z9df985c1e2fe060e8bba9b919b34848fc560719b5c7f87ea3e63348b77c183fe76ae83015cc2b5
ze46cf07e0addba4b0a6bc5467b3ed09c93c8b8ef959f40179a59e86b5d882d0050469d38506560
z58f331aef3df9ae42877e8655065f3570dd5fec421ad21951aea22491fbcca0e0fdc29eb7cc09d
zb249dabcc9885c858840a03e93b78b82f261e8804f2ae17b959ab85890ade6b7f3a9e6657741c1
z7aa8be6bc325816d04ac749353d905532fa8d5d0019fc8b619f5f427e5d82c6272ea6f2cbe197f
z667febd6982651235694fc14805d764827f6038ed6e9744a419c94145882c07009da0293db5d85
z520ea8927d833d147badd4dd52222312016f6beeef2a2d213a78f4f74be9c06eaa1dc836cdfba4
z05e600ebb2b6c3fc52a417e024abb604b17356a281d3a87d7ab33b19ef854bcb194a613a048474
z02d81b9688f693797560cc7436f87e335a98877d0caa5ccb43e00d12db79911b7511315a7eb873
ze4dfcaf215ff685a7511c3a4832b61924181510be87fa6101998c0dff456c69b524e60e836379b
zeea14706df8c0c9a0ae699716604d4563260e09fbf6875b841ab1658b0c588da9ff0242e536583
z8a146d7ac97fb1f0b106839741bb0ff859518caaeb6cd0f9535c5ca5e64529e7b8a8861d89129c
za06273ef3522b169516ad0d177842a632c89908340568c0e16a4d0031591dd9333f18dc0833657
z94059f683733d59fea62d4f2ab6e8cb143e7a1cae5ada96393c79a377c809464d941d4dd239422
z768acfd93ab0ad3d51b9cdad0a6e48d1ec6f2da31c27f64fcd6e01aa38d6177f0784b76e31467c
z6c0bd79d68c3d51d6904ec08cb1510253b4339af2a6463598220c9bfdc0bd0ce3c2d89f26ed0a8
zd595bc175b8b921272cacb8e00655857ec1cded2f549e81b11a3395f87ae00757396703c067944
z0fd93156fe571bd5f1208c8d42d764cd7cc21cb9346e58e48fb70f270206fe423cf2d1cac06f6f
z5d4a6967b537a27c032aef74a06db0ba6986af14d73dd657ddf8246506a818cab219bd12a5522d
z2b7a0f643dbd4e8d8c4f86599096e6f9f3a4c323b3dd7ae513d134be7920fa914402214124f6c3
z450beb43da03f1a7e2128e41aae8aac3a90573aeec46f00b951a94bae2e4a0f0e8d9702f25d09e
z0bb49e78369d60f0e0731f68e4a2a51f87da6ded7900838eca36d776d139d77bc1cb683fd246ad
z554e113d46ed1282bd687b10293d15796490c7d2250e6cf4c2d01aa5edcee5e75760efbffb7cce
z0d31811023c75ebcdab332f9e0c9735ca452008c879aad069139759e9dcc1f7d5aabead0ec3d81
zcd25d6a843296944c1f6704dd7601427c1a10786a49642c18fe99a49da0eaf689d3557c235f6f8
z19673c7ec115ecc50ca050cabbf173de36c9503f02b2ee9f4c31557b5f97014d3608cdc174c99f
z0caef4b9dadaa80fb7d8462828a5321150fe296e93d62878b5706000fcb9ec74a55540aac82072
z64d40358d7001af36b0b72ea5127befacb0a475d885b40eadb97cf0f46b1aae577fe649472cd57
z83e75cdea7480a8cfeee051bb62df187ad1a2cd56d43d252013245d9010509528a65d86f6a7157
z4a4d40e9f57134730b7dad05772c1ba118a4505bb111c75a35190f94c94fb376fe2a3dc63d8467
z0511559a696a98f0706435e9edce03e286a5582078139ed19c0491c00fd49341b1d256cc6cc145
ze42531064855fa56285a214ebfb7ff97ef25b1e556caf8b694b3049a6a9919ebc82f794e9cc172
zfe1db529d1976980588b34816ecf06e6bd09209193758bbf1ff0380d15e462a7d4bf3cf984267f
z7b7fe259b1fc91424a743a805a88b71c4c1b3331a99ba2196d3bf679f2b5fb2fd763e667d6efe3
zc8c52bfe0f8fe999db86b9300580df4ea461cbc01709bf99536c770d00d69c6fc5ae22cb4879ad
zcfdf2c348302bff91ac65c28141ce58c84d3c18f35652825e4b2265f22d51e549dc07a58bd542e
z526b8dcdad7d75d00be95c010cc0dc85996dd8961c98f43b93f96ec10813872972900a6e3bd021
z9c3bd2fa6d943b164f2f60a0c63e551fe5bb817cfe5c0b5fa513fb29578430cd4c90d8d1f45a02
z5e20be8819f7864c2b8fc647d90c370206647ee4f04880eb861c1a968c8e97e070b05c44a03fd3
z29fe05255b338965786f8979df84651c03c3a04bc42e0bbffbcc93b8de2c4a8ffa9854f34e9cc1
z92f99647a869862b82d082633af7571a7f962f219c7cb3a226f2ee34a1d2b91a4f4c1a0a63fbff
zb67039d58b6c51bf1558fb788d8bce8a01f9ae9a307fbcde5718436b9611aeb01ae3c091194def
zab5c90f9da29a9e8f128ee545a0810e8eca7643e730fa63c7c2ed4b4b109723254f27cb23a772f
zc902fa1526caf4f828d856783c6273ba724a5d4f584fa8b4ec418dc1634c16b0c385d8a21c70b4
z68d443f16aac430d37830102dfc275e803e32b481955627a62063d3ca52ba8967e9e57be799ad1
z7744940ba4ba77365d1a7752182f94f4457fd2bcf34bebb7b0be82ec42bc0287a2c635756b1ced
z90c91eea813f2ae1734199514535a1eca26e9aa39e474c4515cd40aad5419596f93985d5180215
z5e9dd631e1a258c16b2d0226ba48af45fe07fdb775f0d8f18ee1e976292cd87e8bf48596e9e142
z388312808282a5b55ce148b1f72864ac124feacbf3073da4e0ef6a039bad0cb1a1c489bf921420
z26d1325b7d61fba8bf2c6c74babc40dfdd606f0870601045828489662f671900d9494ade96860c
z219fbed9903f3985f4ec1f1b947b2fd6129085a83e9834737a5fe84d50731838820dd9f92b2614
zd5626c7c56240783c50cb139d18f7c23db247f2b17369c597d5f03c7fc9d30903d8b87b5f0bdd5
z3fec26afca79c61ffc878d69104c645751166831688be2f113c3fa22667ab6de71dbb4dad272ba
z3ab7bf4cdb1d830c79e8479d1d9e04909a38da7065ee54ee1d0d0884a20580bd86f193439d1d19
z61f79defeab9046ce79f0cf9667cc23dd29dadca377a0ac2096ade7aaef747b79a87259317bcfd
z090a854efe6193ea2fe631b1c96164105a58bad499dcf6bab2fb3aec5f9188f540f4743ec0c89e
z3bae376227d945bea20f8be6791959abb15dc57ee8b39efaffdb9f469edda25b35782ecbd8aa07
za2c7f0b2eaafc698a0435974a368aab5ab9721ca4d3278118bc3a7b3dd7a4b1741bfac70debea7
zb3b7f3f1fecdd9d7a6659276c2840a49f7c04792804dc938fb330c805ad8487f88612150439884
z7c5e425847a5a122cea1899e642e05b662c703b512b17c1ee256539750c7957ede904a5bb64a1a
z46ef9037240af2d9f878e52041923946d142a9666bf419b702b8a960c643e076dbbea31745fd49
z10825bfed92b36b1a1f3ff51973d13ac89299e9aaba3e4671689bb2602217564b91d0d426e42cf
z50a64b15ba7eae4b848cb559632e09b6c271a3adc4670d64f3af64243e8316356afa8a4f338979
z50441e71e1599524c045a8ce39419ecad338caba3c11f2839b9daed5b8fecb588e384e3b3eecfa
ze7160e80c69078f74315111238023359d1e80401c2dee54a349216feb9628f5739e04f3a409818
z5f9f7dabf385308fb888d4dbdcabd59fcda24197480eb22f26f9c6da78289c032bfcf3ccda3371
z7daaeb6aa1bab1b872f9c8104c4ff12993058d8ca86fb9bd1b40d40442701a4e90a46d1c12bb6a
z9f63f36574f2c1d989c34a48283a10969a3ff8eb16e8c1d2862f126fee9d0eac414b8c3140b172
z1006d64f5d898a6e450dcc37355d6cebe83eb95548428c98c7630a442f8831cadf7ecfa67d2357
ze358f04158d860a83dbd5710bdecdc4bfe85af0e2686007fb04e9d8cef46d911bf2095f3af52f0
zed4dcb4e772945e4ada9006576581fd02840be1947084496457cdee1e5e29af79798479d0d464c
zbc81f87b45303a5fad7ad19ba88667b19e09589dc4591fb006ae3def917b5ec11e885c4540c793
za8ccc33137db1be2368beb6ee41f433e863f7631db78f457f51624c9e73a854d2934d06f3f7a6e
z7ebb4345270ab4817dc30fcae5558daf88b4df6943d93b05db43d4369acb21942b57addb942dde
zd9f2ee212a7687c4021d7f7417d0380fd49f17841762346049f8a6996b4b0caf4b74d6d376f8c3
z5f5ad4bc3dae50db4bd521125fcd5b4cfadd2a2dac3c4aff70b4d7f675c7e2600eda302f61fe07
z739a65654b5a15a5784d4e44d02b2b1b8cc79a5c0b68ff5e9afe863411fd77a034b4ac323cd2b7
z37c8c3d6d61df5128bcc5e0150ad4d8e7594ca74f2576db24561d5497f581aaedd473a072c9ca7
z0de66fe0bc4f12b6878cce7dde3811703c79868e06973703edd7476cc53262db38906462bffd93
z8e211652a9ce7379d7d2ccbcac867b0836e15bbb82b38b757ded13e1d290c547d001fbd9ccfde7
zce5546958141742bb6de27ca6020a2cbeeff2e6c9c731baee85a0f758fa5d8bbf2456d004c5c22
zc13f9236f09c526ccbadab732d2c8a6dc10f796bd4a736ff1fb6f722d592c70b33b65ce6fcf731
zed47509c5903f4280d740618534a1fba672e86a2398bd8b62ea386878de95b4374c08f7709946c
z8ec5a050be8637b847a1964d4c95c6878ea9bc3d308c15c7142098a7e456c32efbf0609bac5b7b
zf0f1ed2ce9d71dd83ddb4784aec9f83a77bea8a207020883308298fcc6dfd8151ffc23e874619e
z2ca59929e92f10e5ec950c00a8689242a3b6d69cd6160d23612bca606211a0088e22294da0092a
z3458096f8d620323985773635f10a5ceef2ff415ab548ec75d900decbf91efba1c45ade0a22c82
zb78445539dce1bfc0b57d8b2a87aa2a84a96ecbb2aa906d4b70e233472ea639ba57b6c6ea744db
zf9b09bd16f38af9adc37eea1e37c94ef1bff7dcb48119a9878a9cef26fb27a356c2b96b050f808
ze3375f832541b3672863097daeb8103f0c5b29abc05de6195229afba62fd025a420ee899ab9d30
z2846ed439ca6ca77f0c0499a4d18c5fe01b407be7fd2e41aea6e72e9797f4ec69df674d8fb5134
z8c1efc01676c1eab6fbf9a1a60ffda0ad40b4da15074189d7f5a42b1dee101d5b88ba7a3f565d1
z2a0f5d35afb821b6f7ffbabb206f36efbd10bfb977995dcb06eed36802a2bc44e47a84dd8d0ef0
z8aa95f8cab8f5d581f2fafc2980b8d2586e8240b06e432ee703d4a03910860865727d4c6f638e1
z3d8ac3d7a4bb09d3dece56ae794200ba4920c9821408f9539ccd3cebbf03a2cf237235f2c0444a
z8d84487bd779131f0eeef89b1434b7026771ec8d144eaeb41e5007cc495185cad59b6872609cfe
z2dda5608e639c0f4999a00e6d6c998e7bb4e9bb6058b50ec483dd0487ab2c1ee0183662c28bd74
z2b0da6c7a38c97ef96148ee28477d69dd4601a0a655e524e7bac3e0e361a2cfd5296b1bfc3b2bf
z131f1b92ce81d6dc7cf6ebc3021d50d5bd5a165f08a4e81a52b84d9a972f837ac76585ff543553
z53466e3d8bbf4457547dc5c9e8134aa7e72827a082610161e475560f9cdc853c64b8237ff5c551
z6064bdc535b5dd7a726c4b62e71b4a5715737a7799f3352f66f071be3a3e279e64dfb20b0695ad
z5697faacc47170df748990d315ca28d40332f6eebe892882860bbbe43c3a02df3e6d7dc5b88298
zed77bf34dc5de423373305b5d1d0a1d64e41126f80b6b52f063a570dd5e5f15bfee4953d5b0d69
zcc41e889675dbc9d60986a2f9078741afa320d7ede5d4d00fe36f9de0a23ef348da9050e8eea7f
z3feaa401e9fe54853603c07aabad1cf48cff6232c6ed4bfe9738b5243219debd6757edacc165be
z0e2f68951287a8fe8d105a5b8e174fa429d34c695d5c620c5d7daa735b91c225adef03f97888b5
ze66f2cac74d3eab3bfcadc229f7f1ea2cf873bb14d431065f564f65392bfbc4b4c6c371b1e73b5
z65260b998ef5347f19ebce8b68976a8a84421096bb74de7b068a003b5021502cfa9c57053582b1
z8acdd99add341175ace9f5f1f4410168df3fe75768d958fb1ffeb5e83a51d6f727d88db184b511
zdf13c1aa5db022586803ce6fcd4f34d059ad35c44f508ccb812eea8378df2d8c223a320b4ed2df
z5e074206edb238abad85ca0683117649949f47ac092e2d22a132da9c64cb25e7470d40a31c2e74
zc5bab4e8dd137c656f6f1a8109a840602e89aca426932b7f93c78b8d00f6ecd82fa57517420a13
z3baea7704d42b12ff31467f40cb7980f19c077310788a9f1fd5ba6820a05331b1c018d9f73c3a8
z552b9744de9e390e40fda93431b8a55f310611f52cda0420951a335813c67d560794e9152fe633
zec4097dca50fe4345445a2f714e2e9b7b155d15cb4f5a53c5267bf7dc5af4eceb1584d36a2b7cb
z0df671bd90cf362587e76446b9470034c6acac08ec72377a4d37d875befb3aa119512a99ea6154
z45a4e232d868a8f05658c20fcfea9787599621dbb21d3fd9657ff912b58491a6be87df3f85219e
zbc1447c5c997e65e22195886afa3744a74af4dc5974a4824296e546b46e3cc2ee5b5a5e08988ef
za518fae14a4944ccb3ce955967afd30f7538e874a748e605fede8e5130e0ef59159f8925d53c7b
z9726eb4ac3fed9daaa967e076e30b284392d561627fc7e9f1929de11eb6c0a6a03d1f57077dd11
z264ed06128132280ea317903f3cf622afc358088165daa659bbae510c74c712021a8a143a091e5
z2f0fb50fd37054be10221194c002256bea7c49085cd8641642b6d9921b2d0b0beef3c459b3ff2e
za0e8569c46beeb17222240925f50879e2b83350ff340b2e4a00592f100412387c75fd432f88dc0
z546be1204ccc94bdc45faad5b146a366d504be19bb68c63a5b1681c465087721e7916230a427c1
z51b9bd65e0f5dfee168faef5700348759f94c58505fff9210fcdbf9f79604b156d7ca009242386
zfa7e51503179575064f578831b1f1fd5c39b56c50728882a49e49991c788411dbefbdc01c9abc0
zd1b3b837eb6b3026001e37afeff3e28b511545198d288b85511026cafa031ddcc5100ffc55811d
zbd9f376a931a1943081ff438232b7885795ae8c850a5c24afebc78bd13c27520576d314f2f3241
z2a834245ad8bf09476ad60af293be2dac7238b7df82bcb2bd979329e7055e2e1e91d838655c89d
z4ef2e86ee84a255d230be8afa53b399f54eb5163796b8cdbbc2c0e4e3991f1efda0d9bad89508e
zc117bf9c65716bd90b710a59d84094bb0faa372ad1be6be3b1b17322392598dc33cf8976183fa4
zc7109e22f3582253336747665df3763865acb44307c4b7b4fd1e23b37f9c7c622949585a430c6d
zc57af757377f4ce75966b7715c8a5fba652d8bfbda2766620b78ca552143a180c085eae86b3965
ze4beb45415cb0c2c7117f37b860989d08a28e93220224a28128a1ceabffaa1b52794e58edc88c8
zcf54837857868627723b33790d8a3d694aa0056ff7d56abe886f02805ec1de33a106f7199a7b4d
z5df79b13eade1ef3d2e1ded9b7e09069b6df98f865632fa4ab693d6be51efb5499ce6ede072b99
z466db1ebfc8c00777756b777d06dbd214477fa03a3f996bb32db60042054f6541e41e2fce23e35
zab97f2f1e344b619a7ccc85e65bb6d0a87f422edcb4acdc79dff7f1023e2f2aa2c43989e3970d0
z1026d875b49c999810a7ad3edea8e6add76e221f9282a1f0d56f902a276e939718e7fb4671f874
zd4f7aee6dc3fd7e236498931bb355c212c42aa1ad8854c6b017ba01b9a08fd41242259993706e6
za685971c71ab389ad114f6c4f435512172fb0cd3c7407f3b114806d2a0b18aaa6ca8b376d35dec
z744ff13f700207f15c5535b31d3f722c966761ae9ab2cb8dc532a8c2ebcb9c9d1ee434e63f284b
z0b3ecb3450101c551a335a6695993ad4d63262f883e9d942e1a30de00d9a0e9a068fcbebfca353
z42d68d4d3436f2a90479279f3ea7a94ca19c5396bab3060a6fef3e16abf9bee8082204e3fdc46f
zfbc349667eca84bb8fb681081cdae7c75ef2ac6c64a9a0ed1fd7d74e52a934780a997c7c21d5ee
z08bb4b6efcc756715e2f1ad36e256a3c47de49751f57843ddfd08f90b1d860f2091123a671226e
zb8c810e04a5dd35b9adcea6e3a4ef87387116942ad893ad377502c7b16c0b56b4d5ef39e2824d0
zc65927ac9ba91f42d5849e26efe0e224ae95db57ebe7c13a22d0a9906d391a311fb6eac006233a
zcd2e2da9c671e79acd7306e7c982f43a55d33eefe0354fa00e1903e05945c92bf1ce2062b1ccba
ze7134357449f0a04401350934e0b7f511cba74fe69cb95c7fece50f2f6d9d70267529b7dee46d2
z84a1bb121a054ee2a4976e76ba3ae9d6c4d1d697e4b982b98b4d2b57e976e1eddf8c3ed6a13816
ze171232e93a7a17abe1998a86f4f59571f2ce410fdf08b2cdcbd0f0dc1dbdb1905a69502eb5aec
za89aeb5087df350d968f17dbe23af1799c89e1958f6de22ad98782dfac5258acda970b8fa906be
zb9631d9e207b3ce69d8197066826c7f483aa40c5bad5920ff39541e64b3ad4778061dc6c92805c
zaeecd02c465b1675deee2c70bc36cbb02c54990c631272178da298bdd643cc0d53a61cc8750c22
zdce22d8f32382d5c4c8f0ba71cc65fa1bcb8a4548dc0d8b1aeeab87ff1dea33904db7c7759f8b4
z5fbf17610edb38c448a0d9d92eb3f3c6a4ee116b6371107b075b7c7393d2debe9eec4aeb3865c2
z125d2a6430aefc36ebc9397d1e0f84ba69db25619d250c81eb6e74d715bc7a43c1c384de07f3ca
zfde083ef6b83288e191efa2f18ce19066ca8012b346c97338a7a40a3305a27a62c75c54ab17ffe
zb94f9eac2ca5474e6cde6df3f76cbd834c4ff52fdd547f2493a700e2ae3dc6f7120204e20a49c6
ze91afd5f22d48914628f5224058df2897f0f10dfcb90623de409002701d7693a5cfc878efed423
zea6987581a980a3c8a7e7f6f95cf43b0f7dcc31ac1e7755f050fde2417221c0caa87b77abf1240
zc52a14dd70434fa5f79f55b36447dd5c9b3ddd3f61ce912da161ad6c3e0cf16d2fbb978f2a2152
z1d9770f530ab67fe75f2d27b454c5bd619ad0b38e3f1876826af97623eaaa94c20df7aa0e8f0af
z30ac13941714f961bb73a1d28d18fc9d7973983e0551fe8d123d16c20b285f8de8a84c5db404cd
z0b5144809e40a347a7088cf71f10b224bb777e2dc1f68b531bf474273e909bcde0b60fe47fecec
z40086959303b5f62a75aa4be5eec96ab2589cc4a587689ade30cb4bb51ef3bd1fc45c240942b2b
z47b7c8f292060d7fac548aa71ea482a47d6c416cab1dd38c5f881e81711cd57e4e7a879be66de9
z8a8c41bdecbdecd08dbd9228bc5b849fe708e2415e3bf888f9ec7d2cdb1be15aafdeaefc4f47ba
z5d6b68c690896d281305f339da50e9b598408443b7fcfe27e3c60471abf8ee64b13c4e641bffce
zbf74f6ed32b010b100be9f35798976010189e1524241a66c15a8f4765380be1209fa1e25c5ca7d
zacc0a2d817d60af82c303f2e7e8cfa8ebee17afd4f152378e566ec4642295da40363c0c3ae728c
z8388f0343a72762ea6a3156f1328dfc65913cbb14ab5270711e68a2006b6f317ec3ea274e82382
zb8292b90ab5c02e951699ca5ddffe8b1869efa18a5359a03515959388da891d066f28a470dfb62
zb356cb475f5513e558b65e916adbfd101936ef702a8994465d933c82f019600607cb67cef38688
zf35a4d08e2dc10e574bc00de19ae6371e0e9a01fc46cc0b7efdad56be53e21fd6d713983784bcb
z2fb3050cb3d9d6fd3354f302121c6bf1d86eef8773f8e92253b80635466d45a02cba975d494612
z9ba8deab0aa3c8adf27066f474c77bdae60004b070b10c7055c31b020df3dbee458fe53b629ecb
z4c8af5993deed634f15362737ff31919a43121b11ace512f023567eb62324df37a505c58797499
za83aa2cb6d15ab03d1ce037181824e5099363363abcb258122fd00790558abd34dd4cef44fb975
zca29578db35a4b03975d88a8a8617ba39aed92271e65d9b17384f2f09cd1f1a0e898fd82d93348
z8075290443a57519f1bba8649beaf853bd9698aefb35dfdf380faeef6512e45a041d617ce76297
za55ae0db149be679399261eaf9264935a09ed7dc65d4b4cfada7bbc905d055207a27f72d2191cd
z550ad62fda49b7a9e79a4d4edeecfcb943f95732cc05cf99244162f404b45968295e24c06be7d8
z2667f87b96646066952f8808417869244e40b56f8ec470c64e839307ff938b3115642db0b5deb9
z62b91a038621f2c298ab311ae6b17ce1a0515fd69f257d3a566c721ca7597e858dd85a272b1c9d
zd98db3f23bbd4fff46a49df6cf78aa8e94897a5a8a3173fafb72bcdcf58318063a1d0d5f361457
z4282c5951995cd1f15091ce8f47dc5dbcdbc9528d11908753493cb2df559702e560cab50680784
z415c45ef6c20aa0b9162dac851d8265b656d05e2ae4825e34ba31e88c58ef459fa5dbce6d87444
zaaf1a20bfaa72834bfd0db7954151a64ccfe0ea82ba758a37b12d8c04c561d1f5c694d589b00f6
zcae59911313ca64744be7c2ba3d3eca6e5183fc6b67a804f467d4848ebe6029a7fbdd06a6e5faf
zccff299325b9620fafbd3377fe6104e4d6e62845135a7ac41773d6f663ac1a3778ad0be2f8aff9
z036be05dcdc46220f1ed0ae1103067ec96b5ef2f25900d00ab55473a6f40a755ad756f8d7439a5
za27f724eca502f2100d1cf63bf669af20797e21f9d4225e4ff955dda219242d0611fa6175ee197
zcb8a1c543c1e1f0561340e6828e21ae4f212ac1ec8b36850aa282a77857731bbb83dafab35f7d1
zfc170cd5f59b113afe814c293295cd225c64602a46e7a9956d1ae8fe6aa4e670e7cc23ad42cdd6
za17329e131d725b5f3a7453ec10f6ff2f0ce7844d69ec34d06f34d3350a7e3dc14a98c549bb86c
z91dd3c7479afc7ec67c33870bf2f220f2e3089d140ac92a2b1eca52cb749a2a9e3359c355d4c8d
z8474f5f223c923c714d1c3d0790b02a0cd2b719b142f91a2e5e413bcea3bae6bf1dd0f0bce403f
z9ad25d7a690882a78cf284e502a15d7e848473fd79638066813a1e8fa09ef52dfeb48f4ca92565
z156c02a7f79353699edbdf53839acacbf2c6ac2e21e49f491e0cb863c93393a012f4e328ddf746
zb484654cdfc63e564628ed7e59d866d7510b1311b32f49191b2c2260d2e4509d0ea96086443fd9
z99dfded00930b71b33473a00e4aa568b843dc6257e14c7ab4a161ab5422aee0374d5eee63b74db
zfd70ae951ad8cf90eff24fe65e30eec125822400264410ff25b1667c602e9d031ab5bb7015c99e
z2be106777d97555ccd88b1cb9bb0b7e491ef6c458c8eb3a177060aee53f287450fe65d6c54c604
z0be00c48abd693162d15c68901c2449f4663159f3891763e009bb5cf978e4ca8e9c59709505980
zebb1d4442a384eb1dc0bb38c17d4418654fe4e6618210b08ba91cc2f06ba9501f5b318acba52a7
z99b3ad28fb72e9a9828370299e8456f6d8c4a363f17f4818acf7f638bc94889abb544226a7215e
z2e9149bb00d5085da465a8c315d63e9687efadb1ee76565eb356e3ab7f4ad8dd06ca46047f5450
za2290609a6705f5debe40f7d338c0d7f8c9ed161372347fb2a94999740c40e6ed2e09b39dfd01e
z6ce6dc119a63fc2f7c84cf1941bfd7a9042233b45110fc76988f742b1ab64f0cf3ea69e9564967
z253768b6f016d5f019705dcc002f1b79fcce7c8fa3116fe9e724b6363168a389266f8c6b97d761
zf98abefb581e07bf85fa00fddd2d594eef3f27f22e7f4aac9ec6617736ac8180678d594761be10
z28df6d58247f20b4d140a2aa406cbd8a25cad483c9b09fd56cecd6dba74ed09e52e8c1b1551823
z8e22727d0bdf7ab0b7291339e7f1b0cddcb3d2ed8bda4d3b9e06907e66f6cdb201374cddd71dd1
z057a5737160666635b0cc0ae56be36ec9f29698710ef211da0970cd111905c34c3993515aa0723
zd687a51ae4a371d22f94155596192255f10e7f7768c1a1d9260e7c7b31042e77dd11c7bf204f12
z408206525c759bfcbca942229331a46cb6b3054985f022f1459e9fff052f351dca72cf8a009271
zd04850a5e7e66dc7fda90ba6b762c286e2efc2a48883bda36bc45cd9fd931f0dbfaeea21f61974
z41d208473ef188e132c66b2d087255b36fa2ecc02fb2d1436465b63902e7ca62b6cba2046cc6c9
z8163453b94c8d1ad4e81d358c8d1e4ab22bbec500ba779127a6f2edeb7560b7de7e2c30c9efbc2
zc76779d31a7650c8389fe2f53aecf8d2cf960d7f7bff8eb76507d193eeaae813d7848362401108
z7aeafc201a69e1daa77d45c7db3eba2e37e6c11c2adf8e45a671ce9bde4f30a01bfc7b34866758
z45a57eba67d45d742c0844ca49f49c976c1bbb9dbf9a9c83df1b3b184f2658951a90b0d3e6e928
zb17a75638bc209f3f4223c67467066f449d06bd38b08ac93160256987ea0e86b46c9c6d3b2a292
z0c7577685a00f082046712062b8db0614adf8d21cc8fc18ac1bfe21143ccb1a04b090c66587768
za8ac305bfff86c2f2ce93d10a2093996ee4237ff040f1ab5948e9d50a699ff63c4f55b9d38c8c2
z5a804aa1e37dd850aeb4cf1fe3382dc0d7a787c2eff58369e99da85059d793864389a74b1b0e1b
z98c55620f90d6d815cc63e64e5d5aef5d2cc554805384fb3e0bc93b30a0a8a8ad7b6fefb24cb82
z3f8888c3e50340484b48a1e92617ff2439f68ba4310dad5dac5203753453b668430815792c3fb5
z637ecb6a72edc0ea42e1ae2096fc66c8ece0f8a6410e7e4e77c43c20909d3190f2f2112b2b04b8
ze505598f09dad1ce340985e8a3828c592feeed943a4db6311c67464ce8ad91f8b1106c4011dd74
z4e77ea8d5460440b002986b09bda3534e91b5a534b6d61e303b1ffcd82c3a5c0189ee8b1d6232f
z1f73e510d4d8d24a609ae8d6907b0f5f82783d08236544f8aad9dfc9e110b6b1a5f4dc51ddf851
z1861a0659ff26b416651b8d620e5bf72f03b550cbf7e532284344015b18829f2ac8860673a377c
z8db2005d9469c20adb1276d9c29571e27053f267f9ae71f920651fc61b5472a8c6d870bb8eac31
ze4386e3ec2189d711b620f675d62799874bbfd9c0cbbb2baef0bd9e80ae70c7d434741b00d5596
z3c72fdf4f3b6a50727ad2c3e0c464b9dfde01a9fe4673b7e659f8afa3d4f55554359f1da08257f
z44dc40db2473ee2adf07a30c2857f0087a746df9ae144c83e8da496b1c837721582fd7d7c8b7b5
z99131ba9eb175db7b7507a36f5209327c8615f567d53d9481042fd32785acb4b95fd87859d2691
z58bcc596f9363d73adbcf85096b935be03734a4aa72394edd23942509c7bb25e6f84dd1a52af5d
z701acda3d30eeacea7a1d3cc83c450bd84a20cc1ce8a190cb3ec9de2ff8e2f17d90ec84aa06532
z43849b842eafdf629174d26c1d1d9364e8985c0550d220f9ea3ae1a9acbc94fc08fb702782b53a
zfbb3ccf2e0c86c0f9855034ed0a8d2da053b4195d295562ce86177e4f04539455121b5546f21b0
zd518d8b8c8a1ce30d6842ba409f120f83a3b41ff46457e4579ec925fd805f7565c9a7eadd3c01e
z62e465a0a1a6053c2068e25a39d1cd752fe3824b674f480d3a4062a74791a9e3ed8c7c38c02777
zc6323fed848be488dd49ba1886558a515563b44780934db104c5f1e6cc2241dae0c454d0a113c0
z92c04e56e02e06ef6a6bb2dc0b59a361d331d6a09f7fe9f221e7270fb44d75939a67fe411e0c21
zffef513b36e51cd8c43e62c7ddf0a542b4e5a3fe0a7644e6625116148df3d81908fc6145a1cfa2
zd773a2b5979389bedfe72c03636cc34e24245dbe180bed01ffd9ada73394d29d108fcad834850e
zcce8e3738c7dc37a2e8770e4d09d9f8a5ed4aa24d516a06112365d6015311160b7e49abec6e3c6
z066f0c4a92d1d0b346c79fe4b81f00cc0e33345fdb82245e3272b66564a353e7c49431ce781823
zccfa2679c09b40dae813405658f071bf96c10d4392ea5b1971e483b34cf08ff438f6c685643dba
z9fa3ce051eb7aa838bbde2d5bb12ac05644e1f0a7edca9a53403bf5ebabb019b847fbcfa0c4d01
z23d689201eff8f24650366e8a6b372bd58b0fbd8ee55d2454464d23298a8839099e0d34389c24e
z9911d31bb1c581d09a14aa49bf4e47b25eeb1194bec1e1bafc191c4cec45ea8aff8341b43e3439
zb2cbeedfee7a86956a959fe42b60fb6527e81cf58aec4b10e1adf3387743761298575e13fd0802
zf0b131cfa587e2c4b4a394c44b5deb03363fab1f41ee96e7dde80433dfc6dc90649cd9a8154326
z6c24772fecd1b4e6bce67b764b6ebb4628d57e5f28faff2295374b7e5c0cb9ffcc7cb94e768b2e
za93c42fd635685be6106ab81349a074fc2335c82d0585fcb542a307016fa325015dbe245978bc8
z883228a9cf209bfab938b7febf96987254093e1c51c89acae9b94c0586928166e086dd9aa83eb8
z80132b217f1c32a2421de009f964f1acf4be963e52083ecb8af96758cd5bf77482f84cb8c48f54
z5417aaad96941ad584d4832805329653f3411685ef3b58ef55adc46cfd189e3f2a519d57de9e5c
z469d990e4ac4d48c403a863d933b73b0378ab4285dac1695807db2101eb90421f9647b3c8e54ff
z7032d4a27ac011422f8b93386863ff041ba289980e43063c5ab6a85b47eff6a37ecfff1a82567f
za10d189129db2b2492f158b117affd8cd1789bcfaf8021f63f1a356d68756d388e73e984bb24b1
zedf894c3c272182c09f76303400559166ac83505f69cde6824af7df935d09f4bdb241e04b48487
z0df24ae641589c05fcc53ad2b641ca2f3873bd164e22df7bfab377a55bba005aa37d84500d49ac
z283e6eb0d82625ebac24d545f6aada2a797d95d78da397c8749fd31cfc35ff7454cf37770eae91
zf9d4d44cde7c86941d231e720f0a783b9feb41d27e609b475c914946e3b1de09e335ee7620ae40
zfd7457ebfdcfa7acca868e05d31d51df083f8519a88d6fc5e9a6b57287a8f09aad675f8fe025e9
z9294e3e614d752f7899d7a0751083ebec339c9ec97578257cc2f378e60a15a8508e7cd2ffccee7
zde4dfee0d77a88b6d6d5ce121a2e4385c2ef585a89dd2e330ca9cf4594be0c72cba24efd3ef355
zd19d965ca6a5f85413aa54005760b7fef5c56d9b8ae6905f384fd11dd9322aeaba7db917e7962a
za5d471477fdd4f25bd2abdb8450578538293675d28ddfda438980b91af679b6016636ff0edafa8
zd2342cd1734f2a43846c8367439e341b3135687614aa65167df7e57f20b1fa0c3fc3cd8d726c0b
z8a735f25e3c6b8e5c06163dfc302170664f32875eff8080be4ae7d98cfda1ec5551b31809477a9
zcd513c50761b32e659b2387729a85eb41f1bdf225720062fb092dbd2ed8baf5f82e34909711cfa
zc0f6595bb0e7b11427cb795baa7e71067c10cf115624b8b6ed4bf690a3e4eac11229ec28e33259
z96c373ce83867173e2ebd99e91479d4f0c0236d52aea0b17f269d8a0afb5794a296ba9f4f34632
z7e2bbbea1dcf63e70454e8e430f54956f0499b0c682ea7a762c8b3bafea8f937bb231462cf747f
z429fe3d9e8a35926d6a3540ecac52d9da73426c475cfe11af9920733602442740cf359218e33ed
zda1922ddfb9bd9907b757d9097460263bcf8200990796410d675d6b6a7e3d915e40f7317e450a3
ze41dab989a08c91bf1270fad7186d92241f790647716e7a4cd56f31da21a99a71891c926f48a5d
zb0a8b9cf8f6cb0dfe6bf7b52abab844c022371c3ec2510c03d2ccac8caac2e441fe5bf0afb2c69
z823fca2c1583ecf26533d1c42b3db8e5c911ce62ec387cb281bee5963249c9b30ef744f8025958
z4e97412e3048162312ef9e5188080a56938c18f68ee2884bd75fb0158f422571d0d69fb00d8fe9
zab068dacfaf33a9472660662b35ddf9001ca108026ecc79fb8fd3354638cc119df0c47017a141e
z395c59d1c06246c48412f73036c7c0703d9d54f9cf0ffefd817cfc17b288bd94b3fd9b8005f53f
z430d1c7f9d22e1b059f9f6a25fcba8d1342359e6b78d1eff315504f9ac21f13fb0f3abe193bbae
zba60506e186290ae20cafc9e40a6e0e474e73e3913bb601a1d75002330725a66a84b319aaec3a5
ze73d058fcbbe4d02ff1773576d7b2dde5301e3461af7586699f64a700ffa72646a56f0925a8069
za72518d9cec73121c1dc2f3c05080d9d9b570ba4ba8a0a36a69d860895a1edecbfb246a4e7ccc9
z099502826e8fe3f5001caea51b167e95eddcf6397d1dad090377cdf8227ffd56cde3f8d19e6eb4
zbcf3f0dbc83324d8c67fd3f521a50746c56baf9b1463070f4d23d0585bfe2aaa9da9789d61af3b
z35354bf6716787cc98794a1be08fddac58cd730ad4f914e1b08f5ca42df87825717129d6053712
z827ea80553ae277ab2c8453055daa36e9c831849e9688d5d6ae285a7aa615285025c02ebd97b68
z00925ecc1e2359dd62165bb62390c263a04c95ee8cad713e983e9fd867569ef5a6fc5d64097041
zf9c2a418cb7a90f5dfa96e268666a610ca241b14f8c4bf74e33df2b82901002588553e696c2e34
z7d91dbccd03c32a9b2b1e55590e514cc460b6e428dccc892ca3808b7511e3753252b4d276de8e9
zca544dd6579c7b1eab9894e9fe28986974d164992d86fab9ea04f88ba54a676ea58c33974c46d4
z7fe5812f0307d962d4b414074c11b5cf600d1f86591dd268767aab48735fea715b14c93941c0bd
zb6e7e7c65f08744943fa41829f8570ee369af5fefac28ad699bf72fd2fa756c99d672920f04f66
zb0007e126cc1349169d254b1f2f3c3fdc4c3a88e539bddee73773fe10d32f24d1e06c6d1bcc179
zbb109df2c1713f9d4d54821f1b1da3a4a930127f1cffaab96e1d804723a9bc6b1abd7293a6b5d5
za7ab1fb045415de92b00489203ffe1b8d97eeb8118ee4d4017494915eca9837adc900c2a31290f
zc31ec626e29b846fdea145595b55295642d8539551248d78033851a9cc2a9a5ba6371f13d555ff
zef0535d880de0d15cdc378e9d287e4235f7b627364f73c75a70efad79309601bf095fe2fdec424
z25ca002b7167170c1bcb0913a6f667962bafb9cb45079e81cb36df33e388139d606a9317269e9f
zdceb41fd2548d3d0348ef90e9e2d721bc684adfbbb32a404a232c8726da58c67f69f885904b3e3
zf3901f2b2579d76580695893c9e3144e5e672fcf9b521b3e908f5f4f187a6f927bfe184db51043
za5e01b29fa9525a0b9bb678e55ba44a46fe3f0e09aff18c1c0872c8d6adb41cb43556bd5a9d26c
z888c9e091ffd533c9a64ba30664d984b3dc4c099cf3c10e9343b75557189310920617734b47c53
z31880cc1d9fde93179a09101168165bc6ef3b724cfb9606ade62258a4dc7984239b13f6a5ee3d6
z1aa3a8707c44ae0976168e77c83c08fbd09b66c59b640b0dadbf5a2b0ffa52bdf54ae010846386
z93a0bc9f95077178b76bbdb466b741ff1834a4f6889a371039f09309e738de5bbe6ae237543b49
z75035300879edff4a9efb1b84615f2dd17c0137e459f8954f0b16f8ef1748d04673b17251fcee2
z0f659979f305d5cf196a260c19c190377dc6844396845be44ec5baf3c19a36ab0f5ba4375e3399
z26b9f7b3adffe80bfca267b00313d3e6d77eb222ce181528f8eb7f45206861d715159e25684f99
zbebeb9a3b0122b7996a10de5135dc0117c605ae890e3f046fd63223819fe15bcd9c497d6519805
zdb9b5486fc894cf6c4ae1ce132bec3eb96e9354dc3517231ca08930fc51075cfd24de46bba46e1
z4b83c1c67c77d07063a44d9f1a928ca5f17d6fed192c64daca54b51935a855e4461496c105ed3a
z3ef4dc37f64996dcb7f8774fcf049718b681cf8bf38b85a7c9eec79cad8a08ce38746be9c7636a
z5a32ab97a95dae90b7ca1a4bcffd4b711e613cd78d2d9cd11cd26a2d4ad1834c328bcec06cec2b
zc4b04fa44d8d6e3c8c85d74481f488c3084d2a7989f9182bea8794b7271fe002bfcd5faf689e57
zb27b5bdab18e912d1567ad7d828dd103a56e04b266d30688920f2ec7083588fe27fb912e90609e
zd0eb4213320172fe946ad24f053af060394b10f69303352be9f7da620878a3cbeb0055d1c6d8af
z4d5084ec2e81e2b2cede250b4d436bd6f9e5ab18139b49b579c701a191e51378162983686fb5ff
zf6c8150398cdf570e1dd886fa068effdd16726649e14a9715cbb8d7bf58b24b85ed46f31f51616
zbbb71b944fdfe29e1f978c64356b677665bdbcfe0feee019eeaf3d87a95047b77e6e30592e2ecd
z8fee7814afc6caac37c74d50b8c976707b4e1dbab9aab3951800684896af17793e9ffbcd83aaa9
z5f0f5d5a87d68014dafa17149c06aeeeaaf83ab1c486529d0d7e10563a23ce0800e4d4f5824e81
za73f24d4252f0cc42d1e17088f8f59e04d37e59a187553b7bed3e0c6322f24cad79bbf44802a33
zcf59700e098246ce69df7d46d4a3c7331e66b9d02dcf6e9b73cf7f555f72d83d320c18f5f8ede2
zd51fcd3c415693274b5095966f5993b2f8efa2edad7c3fd88634846ab7dbd63280a254c5f8e1fa
z0122b75ccf4389206923e8bc2d2d5fd8b3ba90909eae9c1fd331b0e929a05907a8c2671918f23e
zdc2229fb7870f42f3f6d43ac83b624d6ceb8bd432401c4382581f2c69078f605b9db99f8249e64
z673eab0b5930f83d7aa6ae7b834125689d5dad79586702cfec0b6023307113d82909b4573d18fb
zeac183719b43c13e764340a9d3b86ff69b2efd01ec55ad720ce475d029753ae230aebb7763bf7b
z627cf297c69868b7c9b9a252f9534ea48db436e7a8308d4a45b1f6f91fd52eb6c6a52af9a00e7c
zfddaf187ce59e1035b113dfdedf70f2bb19977dd8bee41a7a63f73fde6ffa08291397d171025db
z26b8cccc68374e0adcf6aca00d4441388ebee3ba754a2ac767134d602ccfb85dc22486f07b2e92
z85c862c07c31ffa75e264f5fcad7b74681e37d10c81c88c3c3155efbe1e4508112ca383f809036
zd83670e87f16b6f6880b929e870271a6ecc59e9ac8f5345e1739d23c4a2d89c415b9e10f36be54
zb0354fcd4c942886a5b007e07b80fbfd1949725815e2250a2aec315d3929d3cda25c112abd8c76
z17b58121abaada45f689c89b8d4a00220ea23146c285b1dc22e0b4e3361a07aa3cbcc1a896e36e
zdc5ac2df9259a1cb9a68a41a7727300e4d972bf993f81db53a055af1c201bf2e02409b797e2485
z44c6b35690532220867476afebcd1cd468940bf165d2cd79a6f237504c2a4a381fb6b01c59e3e4
zf0205c1b56769f19c454b2d2acd11fb0c7174d62e36cec4ac5a8b6f8ba8773adc513acc846380c
ze647b52c1b36ee6e590baca189aaf69602d2909cd8aaf81c0395df2e9290cf67752304c698bfe0
zeabf2cde5daeb7b49a92c4245825775826e14383f20c8b1bdcdf16fc3ac01f824e134edddc5fb8
z55cc252ee5260714cc21406bcbef8df3ab6da886cfc9f4e6f606e7979c36f53a76c62be811a3d5
zb0bec5243a310490bc34cfff30dd020304424f2a6af47de856f16c7df570e2dabad8176c032487
zeefca879bb34740312c7f655569f1f9fda32a508035ef42b394fc2f297a0666638d9b3263dc5f2
z5ddb02e9226263f4c064b014e9ec88975343b1396af8157fde522d198da193e78086c16a508950
zf92c0f3695456beca338ef1516f84b1daf8e39291f6929864777386fda79fe0a00b441362ded1d
z1b424694d35f586b4e39dc3d2480eaee90d95f9ebc08a7f746fb4fa80e181c4173ead0282badf6
zb2b56cb1b762cdc615e97b9ac3e2b594921b0b425a76cea031720e13188bdc4efa7e0303bdb620
zb01b8f2b2e14b66238cad052227a8c1c4a00b6c74e2fbe299d90467b137a779a28a9e2a98fae4b
ze04eec181cb91067bf4fa7c4685dc53fb4f52efd3974443969e5c3ac34d177385b535225344b85
z9222d36cbb833f4138d3d6e5e4385d294ec321e07ee51cfc4512c26f37d803982011ff122c3c01
z5bab8fae481db35f53da181e58c3af90a2b32f3945c221cb86b822564354f9bd09c38e8726405c
z740fdc3c782d7f9f4d48aa5a53c32e33254ef60423930e8644004b012ce4c06949398e1293d52c
z7828de4aea906ae3ac7bf087db38185ed8dc31431d66e85cf4cd983d823a7bedb614ee7975790d
z933a14ec8646fb2bfe3814fa94759a24cc80d6ac16a8a69edcd78fb2f33f8014b21e735c3060e9
z9dc501d4a34d455c5f9c8fc21dc996a14772bc9b9863fb1b71ab4dcd6f074d19edff4dad9f3f37
zc20eb667845152a9a93f97ce27dc8330177d5568603348359e45b3bdf5a05a6ff72349d1ce385e
z315d5103e3f1c0181611c1d8d2b5f4d57f5d24ab8fc5f12dffab112c83bc07b008f346b7faf0d9
z2b219d1f739a178bdb56eab62723ea0586cfa6d4d78eea7eb2a417047113079794cfebeaf0b16d
z7814902686011133f4998aa530cea733521f0300d7b9fda7ae6bfc0b1ab8062391d1ef481b6e04
zda6e76431a519b907b4398d4a3f657913bddbf6743c57c3029326b456e37e700f127752c608ad5
z68069f807d39e06fdabc39c359a6b59772ef7a4d2604d297184e51749b28153562848cfb8e6a93
z5bc4708e35ae038ba72aab03a200528063f7b416a3c7383c64560cdd89a03fcb668e01ccc602cc
z99a3d432396524daef94cb8c2c1d6f6e55f3d1efc83390b11e2f1d5a31d5e2b03d7fda9f3018bf
zdbd25e2ec6c4c598540d97576ebbee065764656a83e1947ff11d775e9b5a2cd1706fea9c29b02d
z8ca940a369f23c6467d3af7624d02dc5e3b548a2f68d1efda4da637655597605561f7750f85a57
zb75e39cb89431a8563fe273387812a9b5d861b869be42ebfb5bbd9289e917fd5379b800c0c2015
z4b8100f6f291824c8d9dcb6535c417bde6ba37b01667701f32380f0934f82a8fbd338207db320c
z04d43866c3b02af8b0b6f7f3f0034af191962478991937c7628bcd3cf39f4ea6dadb6160747118
z162fa898c056ae26bb2867a126cbc0164d8d350fc50b5e00dc07d8bffffb7f0347fbb2f35456c8
zd2141d36ce293df6e04c47c24781535a7e93dc8546a3f695f4289122b7da43c94c05e88afe2378
z898b57c11f2957a562133e109bd7fedac182844e82a013c9d6b3fe22590af7a7ab8f14062a4156
z0e7baadd45435ca5b8a5e78387cdc239cdeb0a49e9040dee6d82ccaec96d2db3bf5f6a799f54c7
zebf986746b1c35c8205685719632ea3793687e25712b3cc062c6745ee01cf006f5737a8dcebe15
z6face1048e704e0615b048bcee4507000e3d8fd9338c72d01455b6def8dc49d05d0c45b2af6834
z5881e53382cff5d5d4e2478ac193535ca05976952be6c95b51f786f6b812fb9204c2ffdf11e35c
z675f07299a19e7c799c474038e4f390637ad8ab8268d62e47429b749257fadb8b7b5319ad832af
ze4b152b054942614da668abd5d5bef383d6e4cba67c3e4b4de3afe2470814fbf47f15303578e35
z9e4da5e6a283f8c4963c48c2e7a2b709effe986eb0d7b35eb898b1458a9001ccd5ba0db9bf2476
z71c31f6843bb8ca6af8ed735a98ac0c4a5f9263969d4be93e8361fd688d984ba0741bd0006bd3e
z05e00bf4ad8a323660bbe791cc914f00a6bb14d36d461ae756dbbd5a6983f7d353fe161940cc57
zb22d9ca19da1a67f1fcbf0bfa033fc19d4d35d58d2153bdbc36aa8b1a6be66236848eb50efcfcd
ze2fd77d9114193f97de7c061152b0a8fc2bad5ecbd61f2c703c1ed3c2669b4fcb4635b7439a956
z25dadce20b89cdd71ebc8eefcb60e276dac93956acdda2053ffb09d77e09a6d6dfebd78e45fc40
z1615f425f224bf5b047dbeb4f2e2cd45bda775eab08d6464db9228cf9ad3714bc4b770c5eb77d6
z6b38daab354dcca296c08b497059eb7176e69a86eadd5bb2487342592a5e3ca9bf9ee33407547f
z11ad76508044627737235ab5476215b7f900ec9e5355e2b40ec2092985628e3528b55e6abe44ec
z26cb486887fa94ea751deb0aeb83b0c7533f3e7aa2b60f91e373ea04ff0c6476d758b1f33c1116
z54dc8abd3e93072a29ac8a0f092961e282c6a36efe505f80445123eea50d0c99a30d919ad0f308
z013aaf03dbe8b0e4aac3961def981f3a923a714a9f83d6a5ae5d858ad8b0c9d9f0f1723e3b0721
z18bb833cff6a0bc5bcbcaf4d7c5ed78b20ecfef77aa128df6732f0a681cea1466a8dd0779a91c3
zdb190972f596f6f6893f6514bdc9182b1c77a499a9741276aa2d2e02bd59d70238f1cf4fbac793
zf7b9c7514ff332d30c4e18c95b4aa102ceb606f717610eb66dde3c58ba46cb98fa8bc1af70e8b7
z1de836f33f484d032a80ebc67c613cb10be0ca7844561a4aa463fcf5b92b51c029a7fd5d58be3d
z07d2584c3e8d63ddc19402daba758a823ec67c0e660a311a49d41b222eff9a6109d68314450a09
z418ad7fb46101ce21a09573ff2fec80378b7a94c8cf6a9c17f623fbf17df68a32780c0412171b7
z983427d34184796c746cd37dcfa7f23be41db66741be037dedc095586270f138588e6cb2129d24
z6c843841e28576a2900a283a55a8204a12da6b5a9d03a1a559168a752c45f849c83f2b35023811
z69a05f39d8145a2ec23122b6a58109659dd1118d23d2b79cf149d1b96f76d98dcb7e2165f62ec0
ze21ca4df26d197656fcb1779e97f4fa4025d33bc01263bc224046e1cb68a0a6aaad3fcbd929f02
za2dd148498f577da23e9e2eb2cec50b818df3e9d8b64450363e9f0e6cedf64c4723082f354f7ea
zdbf364d35c613a8aae39f23a64707b47edcf2ae691b4ed0199fb9458cdd9196226be604591758b
z69ee7b5c68a726febdd34cf4cf319555c8801ab7ca992a4d97e644965de61800a5e371ade1ef05
z160812d9f1ce0ad60ed4fc8a27c2e314b9050f4254b6c6882dcb6e000df2f830718b7bb004dbf3
z88b0903ada27136cfd5b3b8d5a7af17c04f52524c547015621c1088c11fbdb8141ae74bba1d00f
z496d164da986acd4369f5e402bf4d14faf565d8ce82890a66a44cad0deacdb7002ff17a89c6839
z2c19376c2f7b61d44254c97524ef4b6db4b3d1445d7676239ea901686a8ccbb6e7bd806cacabfe
z855c60d2dfc51b6b4fe4ae9c12a102a45a843ab9a847a7555915f321c44f3664bf4b300ac7e941
zd1e7313615b148e11f74bfdb69a4f00d6d680d67f69690bf61625d6630d6a4eca091256d952272
z337fca650f7334b4df6f628bf1e1b2a845edd077ce17a1e6ced38f623f70febb1e295a250d32ce
zc0309659b4865ceeba31d30c6d57609788e58455d1558593b8f2d8b9f30a6772e63bc0cddaea5a
zefed3b47d490daf083fca8586c062b675c75a23ac9d9e049fcc389a7adcf362ce29a249b5e682a
zad85e1fedbad01a4a3c13d5da0931f3f86454d7e488e2fc6730201be446a9cff287478659adcd9
z9dd2fd496ff8789b1feb0a1d22c73ff573047f8ef0bc54910f923b8978af8519eb072aeaae7988
z48be75890a28536f6ed6e873d3571d8d4f2dfad03cdde354ad0a8f6dbefd4f4fb454120ce72763
ze77390bcbac941a8da3da44112328b0575fe70618c42f94dbd470d4a30b1c50a1257f445dbbcf9
z774ccff2e5ac0ab8c4bf89281bfc0a8bfff5b03e3f1ead32b0e645bc6a50c5eaaa9e2f9ac47499
z6426c1cf3cadb9cb0c7eef11f312f2247cffcb29299ed40f95e8e4d80078b910f900dc9232f795
z50a2fe258cdbc19079509b73bd1643974f919c53b66c8dda330ca618c8aa34721496e4a59b137a
z22c4ef6c00e719c4af9a2cab738959d2edc9115ca9aebf48578d3ede0efae1a331cb9687b4f3d7
z4bc22e7b477e013fbf37b7908de9fe76360492d81484f166fd8cdfb3ff1c03651372a5a96fb5c4
zff504482c136917cd7ad093e25a5d899d344ead5c382d94afec6968a23693d1e60da5b1d01efe6
z9d386ee3923da44ba278ed06039d994c84a2853638028fcc5d572977573845a4bb07de543d8c3a
z71dfa9d5ed53de171340d164e7c6557f655f61da2728f6322cf916c7e6eab0ba26d3c3ae865632
ze46c05669465ae3e2aab8e39d55ab4370517ead2a09a57cfa9bb521472846716184898e4565ee0
zf50d42120986f08a976966f01bfcbe2deb65fb5d51273474b98c5e619874b5f65ba8a63dfe6e43
zfac375e8cf676d6aadfebd48b6917a356630783b716fd36be2bfb3ceba532ea21acea5c853dddd
z52829775e5d09d9b7a4ff539995515dd72e4e792ce958483495109173f961a1ef7d993a4ed6a8d
z3b98e18d5cc216ed1998e1fbc746ba0d10666c731824729c1c1ce1ce235cee842329e4913487ba
z0a8c7108ee01dd245a2c4dfcf06edfe75bfc6611dba06c70a53a4dfdb99aa2b68e10c1d8e563f7
zd364bcadad6366266cc3f071bd67d59ba2e49ec065a58285ac228a338ddd55a04a1006e07ade96
z8eda2dd4435b773ce565e0c2812a7f4842322d251a786b96dd62189fdf4fd9c0c2420b369ae54d
zb1e05b58de419f2f943f75315520a5f7180baa128a0f8449c0ac3759191da8b97f19972cb29a4c
z25d48799daf7f6c04316b5e7575846485c921944c105eaa4d6de86ef2cef4aeb9686df6420206c
z2072425ca65499973e846e85637dc7397fbd6b53d29027ee140be796a5e428ade8722be6496d95
z034c46630a0803ab9a7f55992d18bef60ee3aa956a3982dcddeac9aa3dda1d5c25f0913209624c
z850c13d96d74bd672989f060d7f08ee87b4dc856b8f94d333780bec3dc529decda25a72ed120fb
zda6bc0c93e1bf1d403c2965094b5554cb84d57e2cef92a0bdc0b99506f4af4df37cec326957a19
z1792657732566e5ff008aa4ff3d5e89fe7ff8d797ea40479c3f3ed1a4c1ce67b8216c214c74305
zca8275d2138e3470176955d06b05862ba29655284c1fbf1d62c14c7b748b17f6002d0e86f516bc
za05c8fe0a2bd4b177384bc4c0a57a68e533ad6ae1dfc08cffbf665056d02067ea200d836995ab9
za36f627ad772432610cb2c209ef2ec13cc0a464967c3b43b426819ca234697add32a218b951428
z0943b2f8cb939089ad8a0dd10a1ea63f56613ad54d4b6dc4d5186c7bd842fe36f08b47c06f7135
z4ff5328c3b38a01b74fba0f88249f775fab29b971974974db9cc959cad1bc93472b617a21bec2f
zf7a8d9d4a7883f40886e536813f511977c6d5a7337810e9cb6c6b3f1ca2060310f393c4ef632ae
z5bea7cba808e7d6ac1d8f5b740d79e9fdacc09890e62ce992142ce9dd5900b3767e26d35c6bd3c
zbe19fea50c4c567e72b904b69d12f88ce887b0cced3ddcd99efed2e170efc632dc7a1a17d3f0ae
zc03e75254e3f7c1a66d6bba3385abcba7be2574647395b523baa7fa90e81612fa255ee1422f21a
zcea5a7b1a95eec736b981b5e6dca3ec008c057f0d2babde05bf107f7b47a4a60731e87de63a335
z0d506d8c47fb2c9fdfdc6a0267faf40af68446213b48be761d3d51f6e55a158e4fc60455b7be5a
ze44ee2bac8b1d57315bb7bb9c4e514dfb9efd14f8b41391393b13571003bbf17da458ce24a39db
z8ea6003bf49b715e4e2543c63115f4f8e3cfcef73f490ce6c4fb4ea8e241ab1d0150113d8d81bf
zac0e87464f941cc91ebe32c541582f10bc2e0172b2278098974843c228585adc4a5b5ef71bd57d
z34c7f02fbd49b825151f875fff7cdf76442116db20615ff6d275b978114aa96ab8e13dd2d36306
z1532ddbcceb80e2a631abf5a934b4397d90b9161bc8e05d351803c7346e9da909e5c7740a32910
zc13667b95b5a1f616042b9f5fe9577590127dd20c934925d232758493a3abac2bcc42f61227d4c
zbbdabbb899ab1bd3b1936d67fac20647283c59dd182b0fe061d6c57f254458da15ab516380c0e0
zd9b10e9d1a7f4089f09b9561f07ee9a66d4984e1a2e5f722e624ebc17487f634a7f9ecb2401d6a
za035381447dc14c6e868dcab1e4a031016178c98a996c614e8567613fc737b76f77b780582e1a7
z80dee7f1afb8e48d79e7257a9b05a223864bb4ec6ca98785c08efe3adeb153e11f566fee8e20c8
zaefb7ffddf6383ccfb0cdb7f088ca573cf6e65246bb02de4ea171b1d2fbe00e16470e77e220769
z0e84086f8ec1e12d96ade06ce9ab70839146658f17e7585059366cbb6582509b38d2258fa18ccf
zd719685f58419ccb50f254115620d1a8df80f6e073827bbcec14ade3029fbfbb1dd9b0a19172f8
z78dedee04c51c295a67ecb5cc2eb3c4d2da8f68b001a9b86f25b663811a4269c44335a1e8cdee8
zf384cbe0ee78f7f3281a61fa5e184222468c08577ab7c2d18c3a433455177116f6ca344e0e91d5
z618bffaea2d316b3e1eea9153206ea6408c642c3d75c3a34663ab457973613155e922cf9741110
z0fcbf3f71bd6da2cbae1b16765e0246d0279b7cb399fa042910d323f9b19693a996fea8cdc7a65
z826e205c21d69fab9cfcfedf8028993d4a95ca9de544d2a7cfd8e343b276139718f496c07d9b64
z05b0fea03ad11e71ae62a6538ed030c4c5dcb75b475e7e6340bc0093cbb602ce056618534fdb34
z4f4f0ff1997ae92521c2e546651cf277e0454f5f48923712902ea8802d856631c736d886b0c18d
zfebd6e95b26db1b6b14a68182b008849193493cdfb7723de13d71995d4a2c973261e5e3b235a83
z96c88b5e50bbb67e71e29e4c7e32e0a486ce4b2228bcdea63fa8cf318248d8a9157eabbad80b8d
z6bf68bb76aae72e2a96e6e2d70609602595407ebc008554d6f75ac1ef645dbcf3899b46505943a
z6b6397bbcc2c49f4d22dfccf29e2f7fd2717b26b4bb3893c5d5eab5def3504282ebf4fcfba5a2c
zd7da22cbea76857b06c7d6e77119c6d80062e63df7189b789919b6e71d5a7a78caec7e2b2b7cb5
zf59a6eff2d9e9e4bd974fc571b03dd5fecbaac8f841f9cbda736a34482e320bf0f51858a01793c
z82e4abec82073ac8fa5e56eda2375753c67ae61504ec315f3cc6daf80a15752d57f8d7a715ea1f
z35aefe8a752ed5091b4e2d9a2d4c7e817f15ae641c0e429b65cc3da182c4d3e33732b15b48da96
z04d41c4a3aece138c1c22cd4664d716264b019b932a63aeb36956860b109762823d35091595775
z7bdfc88cf0de523328f7f214e9237abc13d1ff2840d97b2217097de45c4a6716c3113ea99e0e38
z17e2ff2fe1933956c3817890048020fa9bc563cff0a58853b2a240e036d4fd14bdeaf169858964
zdfef3899bb3b29e13d8a3c65e19f80048cbf80a057bf80c71487742acf3619cfb937ac1423d916
z7db338815d67030e24bd292deac4bdd8e97c6ccc7584b026ea990d132023fb3fe7be7d1a7e7f33
z0729ed3ad06703a9976d63b67f8876c98b4a9518b2bb4b6c1324154a81b7eabadda37d61db33b9
z7f736d8cc57eaef63ac8ba978672ce13f329d65557a7c7b2f18ca4006630dc4311311966b72270
z119fd82ccf6b2e96849977232498b5d37c0b401c928662cf029c0ed014b06702c3898d3778eb41
z2308e30cd96c29f69821b5c253a0cdeab7b8afd05820c24087846156e901d09ec6931d5d7cec25
z3346963ade3e16e21aef681077b8e0571310faa02512619ce12301246d69808a4eb3969e2c1b03
z1f0d3597a294af587cdf301200c46c9501ee75d17d39965b175b5b62ee3a18ec6e6bcadecd6090
z45cd03ee3fb7f45ee40165005f5dd3815c717d9ea580a60496048c6eb1c8a08fe53332eea93ddc
z217763ffe9981cdad6fc5f05ab5d1feae5d4b67cde0490df7043d32c4e243289589a1938d80c0c
z8590ae78a2a0fc4a3b0e9f72e2198949bae5a3215f1193c543628a33460306b2fcbd6f1ac5c685
z4e810cc191a2e768f6656f1d97521589cc3dc10c2be34042a27b87b87ba52e0b21be5303e03a84
zec9a14dba6ab50d35084cec3d7697c2e2c09d8ce98d6955a785490a56755c574bb23554c7c8607
z931c82c4ece4342411517e7a0d3b78191ea234edf780593fde72020ee2a0e1c160dd9a05cf147d
zabcbbc7f213c51b58e9dec31596877dbad2eb72df89a39531cefb563523cb97f0d73ffcc2fbb72
z9e74baae8d5536c06133b13e7e504cdd4f507bc8f684ecca19782ca4c725b38ca7b954a089a423
z4925ae5be3d061259fc192ff41ba46858310acde6ea581a3d82a3b221e86e60684916e08bc2e71
zaf41809686ccafabda6c5b8e8d1de241c43d1a16d6bbd971361be9acec2cb426aaa2831773b837
z47a42363facc0f52c448d0f60bcc71f2a7c7fc171041750dcf21b9c9368153e87589c73138ddc3
zdcaf2f1bfa5434eefca8cc1a103969d36f73ab49f3e3ad846959fd6f101e7a35dc9a03d35e2826
z87d3de810fa6698354ee80a9f7b7f53fe20572bc98286fc05f2287691030e2699ac42f4796db44
z8bc4b2b07770093fce2dc66648c38045e19b94e2e2333ebc7fc5831059b0546b6517a5f32e4b0a
z54ec72e1b963a081b28e92b743a8dadfd139fe3a73e89562e68d68d21614d3d4c3ac7c5a6a6863
zf85b1eb7458be52581a8e5b06444f30966038162a5f80f04216a99b9d969d259383adf4d9512cf
z98ae14e8e2c17f01022e5c2e02632ddb3fa4f65b5ee81932f6fb0c7908d6859c1bde06c53ecc2d
z9c7efb6f91e5405d0c8f7a51e537241747d5a81543ef0b5b4b6134ede85e5967993888be14c4ea
z6681a7e1c8127229ef54ff0e9f246a8a83d8548a8bbccfdc62da9313fe9bb6324ba869e717a1f0
z170370b116b4ba9bab610219c0f6bd15ea9d0ff43486102af48188c40de31e1000d970f2693ec1
zccea902ee2b94b285469d4d163f03bc937bfa201922b024f3e547023782a0a1cbb49c22bc4e3b0
z504e6926fa3fd04c04066e0871b3534469b2a8d5f9794ed21e4b6c4de66e2ac94ed979d08e725b
zeed55cb87a3b9bccbc1ae42861428fd79bc55790603564798fcb34741fb9e9b51a6f1561380d0c
z755f634f0c1be0a130d751a855e1dd42334a6671946f31b4c81d503c1dd07c0001b28c29009188
z7ca0ccd4057ca0619f9b7525843f14e8f64ee726f913e9c6b9d0fefd54a17bda5a003ea3742bdd
za66fb0b7d2ec3a07411dd615a2f580bec6fd8f74c85b450e394b1f2e57fd297b07fc157a409c3e
z69def9043e6a4fc9280a45b4f32f97a7abff09f482c89aaeae33a76e5f512586edfdada777febc
ze9f9465aafb56130cb21c32f076a4afb6a6a03c481cc0b11dea45665bf73038b8ebd1e188def33
z863cb8a1a8277c98dbfad1d40989918f23f7a6a068de723c0b4d3cfe0072987e657d082b19c7f8
z41c94f918c560420c7c552273441d92afbbf7643c8153718d38ea0fd7351870360ae180d265551
z33ac353c785df66f8da8f61ec767107304fae69cfa8b60bae44f1f86dc44cc5c46a797a5f068b0
z51334102e63d557302c228fb996a768ac05903bfa7d6921b82645ff1240f19b4596456de465182
zf164fdd262a72025424ed5bb06fcac71073d5c115fd3aef2545857b074a92910ed35e2b5d95228
z325bb7e27e5b0f78a4cfaf40c62802f52b08424e3c74e7750e79bdf968b3d002c258ebc4063c39
zaa8cca2ff108cc024316f2747f74cdcc84aab74b256450a6922dc891a7380ae35316661ee2126d
z31dad89b7d59170d784143ee84344181cb3ed859a1228a127edb835ecb1fb20d7ebd0bf2620b07
z03e6d34589529f531864cdfbfa250c0874ec95eba52df789d4d5b7c80c985d53073bdff897d614
z95d285033212793cbd624ff2d0a15bf9623565235dca31d08e4ffdc292bb602d1efa0858f74028
z2dce16286d645d4c1e375b8739baf623c39daaf6041e0986f22abe8459c7f4717b971faebeb1f6
zbe62e3287012dea230eae3c6e63eeb6a52158e89817a4b940417bc10e4521550ef0001eeed500b
z930c7ff84217c91dbc5bde591933fd57b5b8de5740059e198cfefa84a840b720d6ecf735c5db04
zd2d689e96945375bdfa59d79ff5464dc0b93712f6246095e4957f5889eba62ca21f816fc0870d4
z332d4634e7b711e533a4c120d5f187f2f24d6519a0960a2d355bdd01818c3388a038a5fe68fc3a
z447a3e3cde3395803bec70c17c26b0c48d56f111a34a1b989cf008cab967b44d96a5bfbaa0a298
z7d9a659005b98da777c7eaf4ab69912aad5e0b1c7275b41e791aa8909374fb0e40d27b8dbe7c81
z438700db7f39aae0d0af161e3d3746179cd2ff2d3772c92ec6bd6dff3cb7b6eff1ffc527cb5e9b
za9b8570e786022d77ca41d8f6ceab597baaabbfdeb9300d4ee1588fff7358e13a5fc430553f50d
z51e382e2a7f9bbac34d9120110a01f8d58d9e13c708b5f62beacc5849df012f49be8d4b7f0a4f3
z19f295ffba0d7a8212b50cb74017d4330eae047b4d77f5db290ba3b62eb64df30cc6f44abf947a
z0eb8c6feca2a9656f0402344254ba8458830d2e9f661267c0464a5050d1eb2d6446b9ff0519487
z5454c2bda3fb79319e11a6b991b68e08e4470ad78c239230072a7d87d4a1bf3c7028d7f81fb895
zbec62f36b35779b5355565173b2ec5b99cf979d16120e87c700cc075dccfb78eb6649dad45ee4f
z5b943c753444f2de60408ddb26ce13e97d035a091286803ba7c10b4f5f86fe9d4231c9adb0c265
z0a7073dcb7762a3ee75c6d37ab33c4ad2e6d56fceacefff069024a34e2cdbebf866646381d0d8a
z784672674d8c49f14757fe897dfb86ac8e683fb70ed9bc0dc1a0b4e591a72687bcf7b9506acb3e
zeb705ee63b98c8d62d8f49e9033e7fd64b98e27db11eeafd522d2ce7c6c15a7e8c18c45e4dec8d
z47b82c42fb4599706fa737a23e6f1572d007e83248d16697ce267fb24c55ebe9aefeb9dc988e30
zc6f22b2782cc47589011a6864177ee35d80040c9cfc9f9ee1cb4b75d6832cfd0e42fd22e342fd5
ze60dd4520f48a338a9d3ecdd0960784fb76f2407826ff530cc7672033aa68856f19de42ccc75bb
z1b01d289abd691474804ff57ba2461397c37fb28a7f2ac67622b1e4e5826dbf5924aa35082a3b9
z06fbde51ecaba152d143a86677e64eb9c8f8729e0bb14d972cb99985a239d9548c9bb83c55840a
z59400b87f50e56636e8632d6ae723215ce8bd4c5cfa4f8ef83e31a438b165bdef658b8b01515e8
z7c1f5d1baa40e459b9fcb2de862aeee2c09193630b38b7885051d2745461047eedc9de7aaf2d72
z88dc791533d455ce1949c35d2a521139c457d7dcffbd442058f26d83a6685e07a2cb7450b132ee
z80fe72da400ba0e840c899de2dd654ccd02abc6e6ebfffd025ee1a719592c5601ede4bd85590a0
z42657530fac3836d85144af4852350e152fc88eb9803006ad9f80953e140fe2a364c154c913851
z2a34900cf38a124e6755f66e1493e7a3c5c1ff436d9f862d115a5d73482e0640b0c2e70a5dac42
zb34c62a64efc1131d55a2590ff80e8c701901d40528b833001614495d5a377c1bc76802ddc5242
z635ba1011d183861b6e57e54efbd9b584aacb53a2fb02bfca3e6e9abb64f023675e494521c366c
zf95898c3d078aca80d37bd4a2081cdf4e3ee4779744173d48a57f328bad0d4ad2be464ce96c939
z8e2eee55f9f06c7894139a41e3b532af139716abf71589c80c47c6091ce8399d3b224657e55ae4
ze122db3cf7cb67c86a3089800f4f025149fb282faac79a9f4046ff505b207812b40f5fea98dd6f
zbc76f57ebe5f3fa32ef4b57b29e6e789db97df4941038815729477c516960cd5e96335b965edd5
zb4b3ccbc4e70d90bf86c3cb6795cc05bbd8133d5a025e6c94a7156fb3b3371fb5ea69e91bd6af1
z131d36764eb30cecdeb92c83c50caf576176457970d3dcd574cf35b370ac8a7182c8ca318f6a67
ze9b03dd541d09d1acb0fbe9f649ca24bb7c176d3a4b9a0b7ba3ebb5119f8a5bce3cc621c696d21
ze4f20ccff0b999ad77b9359b62a74590617f65a6837fd4a1464e5a20de456e2eba9dd5c2b46c84
zb0fc32c3eccae9b0c37f16592a17e237c35339b9c2f21e69d9147afb8f33dc9a2b2d2e0766e315
z3d8c85df44926740dd620ccecabe46a7bf73d9f352661f97e8ac5f7bb325b62c7effdefd6f1305
z839ec0e95183c31f7f4f8b296e1a5d5f87e9fd8a8dc75b425340899a778dbf3ff8516728b1642c
z69e5aa830168197a761cc0ce6abc0f05ca6ecaa682eed3f754e5f2ad8c4bdc3f9119ec79ee6a36
z942238ed461ce04df792bf576c4c5a956806a8f5a764e4add4c43ee98a5f4a68a6c5d94a033b69
z37b2e3f2b4fb27c2e83312b7e96b8ecf4837ca2a8a76c6d90be484e0ca0330a658d733d6788b86
zaf872f55543a23103b3ab26721fd89ea03ab153e5945e6807cf2473e28c1f4c82beb3351d8db1f
zad9e60cc8f238fb7742d7fd571e74b579bef2e6221949c83cd40e53e9945b18ab73d0e7f0f2a06
zc8d3353c2f7b63a09904eaaf52921f617162c095d69e8262928a7ccc0c219917df2a2d275ec3c9
ze8ad69d8440aa610be77f9f7cf28e57a1d590ba552fc75ec3a1969eb5513171aa65b2d99ef98a2
z27d22db4ae95bf21ad1cd5083af98dda7984906dc4722c2880ce18c26e801b05e27d83703ce99a
zd5d74e9b55e327eb62aeba4898aa7498a581444d83df1d5ba6158b689b39f1683bab1592ed6b80
z2c7ff4cb6622d954ba37e79f1a63db3febc8138c7c92bb4d71f159b5526cb8e4fe917c1fbf6c2a
z61d9d194a11b1973a907d30e4a0329e1e30140677e8f641e275ee75103e5bf753b184a8d94da93
z019f15d3105f6b3498970bc6415b194c825593ae861089b0b6863fd8646546bff33de41d966790
z3d8196eb6255168941ac911013cb1a58b2e0e474f28fe08345d2b59c057c9a22d825f744417ede
zd7c38eeaf26f03ecd1639daaf96f3e59ec1b65b4fa9d79575e8609ef3e325ba7aa7bc3b9931b4f
zb27421bbc16ce64bab808035fe6bc1fd7f129b8bfb67210372bbb69ff0e715bc42672b46cc2866
z7e705516766191639bf74080c35252132c26bfe2e0e09ed3725db45bdb6f88cacb2d2a3981af6f
zec4d2b79e3bc7259731d1deda503c550312ee7d0179e1e627656599beda31d7624d86bfefba08c
z2e8457813b519ff5fd89c5566de26913311dd495153f9c7bc6661a45524ce3cf469731a3a2a5e5
zafb6aeb9538633a7254482c20098a75b3077a4fd4512309c1f461fa25e21d09b74a6ef0ace52df
z93c1eba1cd2d42f29d59e9bc7233831ca8e42e53c3f90cdded5eeaed7ab5ea7da3c692ed5b9e0b
z1937acab579730b8419b4807658741f2c170fe728a464f7f8d9ed37b76745984c1c739c3df1da5
z8e6c0d7a7ad43471f02b9dbe063aced63d4462445646c6ed78ce2b658a398b46212badb2977628
z9d471fa14e7e5e0911185f0b75732cccb45a7ac9c05b15677bb254c596cf4398122a62e86a0c40
z66dc46057598ba588d119bbfa7e633943356dbc813f20dd83cce6fe6bff6bdf23d6f4935cd73f3
zeba0cf754bcb2c00af4536f960bf17d24e4d92bff403ae48584da46b2109226dcf98a0594d4238
z38e2cc0fec350c17389263bda44e3a91feb83a54e64662856fc84b76b58d666a4548ae7baeb509
za41ed5685034f365bbf474bd5f78bfe285b0457c1e601b9ac47bf620fa852df02acd5fc2a034fb
z287acd723f32ec5554357ae568603967c398d3f1c7dda3f6b879c2d8a82da27b84dc15c8a3601e
zeff22fa68318a583549ba6ef67763a0a5ffc736ac1aa0bb43f58478273b7ee40ac33fc70f75ffd
zba6720ddcb4887d6c034a23f2fd0d5f73ae18a00503aa241742fab5cf7ed1c8409d02d40534ae1
z226efd321f6b35e51b0f3576ca4ecb219493528fb67d0185c68542e796c435fdf90310a925910d
z34353241b654bd632283818652b79dd346f7b6e006190e1a61e2c9d64b9e2fcf98e9121812a7a3
ze0cf40f129b41fcdcebcfc89ed25e6794dd6fec06780ef53519c88f93f88214dfc76d963416f86
z60fb028d16762773aa12c35abb05f01b69e075d3a18b98a2b73f6ff7e04d91424f225198d328d4
zf053a97fb06f83888a9cba78831b1dc9af93ae8ce29510601712bb1e5a935550550a632bbd7ef0
z46330c541311f13396bd62bae3e904024a6980d5dcf0162aab8e586d0fcb5201079954dc32af62
z20a08c96a813c82b7d5fa18e9cd4485002d0233c8b2bd2a862ff8c217c9daa24af6e855d150be0
z4fb35b522f82f6900a346927a98246047bbf597d08dd83fb02e2eb1aaf0326e362fb360056beba
z2fb26c308c352ab69620d7f61da73e4cb01f0a8d381a60306feb2d8202cd23b012b5aaeee78386
zeda560046594cece5fcf5c871f9154bdd01a01a969713f633fc0c03b70009b8a15c63661b65cef
z2cb59133bb8de517f7af55e1b712be04ee818ec153d0da297ee0c4af2920ad19735882f3eb9c09
z3d08a6376bed3ff937bdfe3fc79efbc850cb00abe83f8aaec9260891b833bff78f0df92e0f067c
z07ecfcf9ad152c9739d56029c07fb50f0e63a64aa116e41485d9c35f4f4ecd1f4852e2734f79f9
z9ccf84d270a1b56a76388348e5e7243d5296b00031700a6bac430906d2cf0e9fb1be39e79b6108
z224b0e91c6cf9dbb4a96bb6866a8c7a23cd58504a335bfc2bc34002c167130dd6548c030376a46
z91de047dddd033a8c2fe781f6f2280dc8fd30da5dc3863b6fdfd23f21d574f4ae133c0b9d53d4a
z0115b382d7dc6cb8d4f2fcd3e886750c332ba49077158bb981925ee668b71921c061cd5441618f
z206e8a40489cc06ec76430b7f1cf3254dec248de38c7057e7d54cf886a29a8ee5c80867b5981fc
z7a45a474c3c98193765ee59a9c4343afad52312e3edd46dce88aa1dd201c74a4cb156877542116
z69575065c5524faf4ccf447de1e0ad5ad3b05c827cf66cfb3d72396c80a2c9dad0e50effda7505
z14b84fc59b6e10d848779c1082198f4c5a3a1d2df57752060b1f90d372171f31d6664bb1f37932
z2ec33c2eefc9049152cc3d8df5f7bb3e4585039f17e58d6133c8436b08883adcd847636d637ab1
z376ae8e2fc84135cd68f3a7d97546ffc22f2e87d3ab96b9af119bfbc567b35606f5ad0c27c5061
z8c11b65d0e221ce78583b61050cb1f8af34642d4e0e7438fabe50537fa715483ccf73b0d877233
z2d5549f026e8b626b46b49f917eca773daa2be241692a4b434baf26226dffcd45c9a3e90ed022d
zb9311ea848258c0ae14d204f0d421cb65aae945b608ae421023085b32f58d363dda1d729ec6413
zba25b30d34b325b85a4ea9b295b1a81d881925975a6124b8428f0b7ee2093ba965b7278a36f9d1
z74b0fdfd94d2c862e88cdb49ffda89c65be229d4b77dcb453727ce9fcb6c22cb5d3fcca0dcc514
z9c41ca9aa6746147dc7daa3f610ec006ff9d3503d0cbec84a99f1c940ec7d539986adb42474df2
zdab711e7ca88fd0745b908b38cb8a5b6c0e8a1cafdffc50ddabdb26c7268f11f9f5aebaa6be73f
z8fa992c05d090327f8605013644c9ea3b851a9fcf2bfd5c60798211aa83a54cd5e442f5621ad2e
z4360ee6b7ab97d3b6a33979306da33e3241b022c185ffe062d710f0df581ff12165b1c31e1d744
z493ca5a3f8d7d69633a134528d0f476082e7ef3a5d19d50017deeab4b419df9940238555e29937
z3879a71523f32de373c93eda7affe3b73b1c16aa8633b893426652e5b948502e340e1c4cb47ef3
z166ceb729bcfc6267965f0f06e1909ae53cfa6e581a1b8c2db3c88e3c3a885901f60411747477e
z05979046fb8ab55114d12847be0a5df899e99589613771f7c2bced58d2fe87d06c45069cf6454c
z1c1241ed8c7447ea7d406934d51dbbcd71e51e18712c19abdfe41291d872daa7215aa73e115b72
ze6d5c62a0be53bea267a0f8425cf856c51a8466910f9d926cb5b564c6c5833bdae7ba719e1c474
z94d3cf5fe3900831b27eb69bfe4e4154f366620646d3d329c8239eabb0cc81d255e985d38b73b8
z40d9afab8d6292985a45759491920dfa17a2aaf11aaaf4a40fa95dc8c20e194b7c0b8b2d94085c
z0d90012e491bb28767e3b810b961dbe6adb3bbee1a3cab1da1f2f2c7bbae78e6f20ee98e1ba584
z2a3fbd708008ccca42304b4f6858bcab7621c4fa9f3953bdefc66469c44428bf3e3757dfe05b2c
z48f358db38f02859177db2b6b722133d8c9ba340bb36cf32c61c49ec127f179ae695a6bc942e40
z6f3dcbf439e145ff1ea6520eaf5aef1a85bbbfaa01ddfbe253d4c5f64ac80c9c3f9a07247b9ab0
zfd81c7f1fa92692000487a8faf348e48461268f66ff50c0aa358a249cfde770900023b1a7b0c81
z28d28932981ffcc360b799a5ea7f18f3357fc3751925086e4b1b936313b7fdd875dab57417b9af
za81fb2bc9cafca6b02b1ebf0b63390367f7948a70f24d33de7ab2039a059155a2f343439a275fb
z6461fa6b32a9eb03db81a10a3954753cffbfdb8117597e2411fcfbf2e56984467170507dee1868
z091077097ef4e48200fc7604e11a73fa471bedcb2c610105656f26a310f192a4d6d64329b2e779
z36f2bf65dd406c7559044691662076064c9ae29e743d50c84b84d70fba7e34728a40411271526a
zc5f6e37686e2a81c7a9660a290e650cd60e2a649be99a4cc36324db1bc5a35574937cf5f5ba379
za76c2f99504ef1a149248725d9aa6ec990f9e8cdb42bc487f261405cdb9420adee11e7c5b83ee6
za8f0334283c1053e61515bdaf8d09a88e107751db9c3bbd0c4805390a815f443ae4fec9b590bff
zb9a40dddd870bf1b4c8e20392141b72cb57667c9bec35b385fb68824e8e187d587fc4a75a20b2e
za43f2eb2963932282912a8d4e52d7d7fa2f539e7f62128a80ad1e6d5febec40efef705eca99a8a
zcb2adf7b4ac46c94564ce83eb9c0fe58d1faedc44e04adf695b045811a0566082ef7b271d9cc90
z703a11710e0547fb534320122c7cefdd83f3d79b69aa54b2e8f69e743a92e114b3bd70a7abe027
z35aeacb176545aba2cec574e78725bc1a3ab4e2e43d3c32ef61a317db2f28aff698126791fa38a
zfd27d4dce78c9d40fe4e6b686082414783a1c411827e3142419d4e3b580020610edc119167a40b
z0b5e5c81d08f16cc0c8fca19dc56cbae5901d33fc6be232495219a8b5614c3dcc5da796cd94966
z2a01f9030f2d7ed1baa5fb75844253f8f9ec7ec90f26a1b03df4970652b6f47f3befee06e7cb8f
z2a478e76b0dee4344487a0b33731a34f77428046f9ce9af4feadbe146ce8cea94716bdb9332c35
z55ec06ff6e2fa15f8810858cd821b551d26668047c2bdd08fa836bd9714fda9733fe9d91ee2f75
z0473e7d017674886db3632f33237673fa92cb1b563f79b7425f7583d3a9e24f90be405ca001f4a
z13e6b83e5b1c63ba06b4206abc4ba81aef67185fa8df05fa32c5203ae7023d7b16c13effed45c6
za678d2a4093e30c907aa7146c8db48cf696623fcaf4b1eea39408cd145282756565c1bf4fa2066
z3d492fc39555dcdac92854e3e0e57b6a9657828873061c62bf501e1df2d65aa1601b0a854dc79b
z1a721d0acc3e4bf71d7324e128586929fa106b8cebfb7d4bca8aea0ae737393f9017947dd61b0a
z3a58b152cadfd77a3354c2247ee580097826c506d56dd5175e28a05a2cbf5d723c5d3ad1468c4f
z24539237a16345901b6f3cac450b515655501a01c12c88e151ff0f6e553f84fd860bb29b8e9b93
zb32229f828ff73091f70cb076fb98d11b73052f4500829777af161d9656e39811003ee15917f4e
zfed342958e103fb78b136a0024295355d3adcab7d65ef0e5b66a517c1f15e2d464df712fdc4e74
zc51cf1c9e4c68b6ca95e01f82cb658639f828da83c8aa7b6896c0f9d259fd916e181643b5b3a55
zf9b1ff3a5b6c3f9935ce2dfe49d5e37830e97c33bd249ec888a358e616eea88caa50509c3a7f48
z0752e22e197cc169cfe42186d8ad2deb453d70b38549cab3f142beeac30defa8989a16c804ba30
z9af485f2fcd5434b04b650bb3a5812edcc160a90c166048a5884adc6a4109bebb149b5b1f088b4
zbb8cf49c3de363a7e94ef8d989cda5fc8b9c08775c7ac8fe3b0def2571d7d052cfe4f4daa8dbdd
z5f76a0ae7f7ff71970fb899e776e936495d5b6e6096a57b696e92304595c25986251fdc14144e7
z84c17d1f05a29d43db77dda137ebcb59796b3f8e5b870dfa10ea71f8258221429e357d2b9c9846
zccd2b63f88b192430101dcdaeebe66c4015ad6d7ad46eeb24c9447214a288765a757af4cd76308
z56d0fb073d3c01243f4efa8481b5042d1f7b26f5978509c49f1d2c218aefdd11681353603a3572
z92363c0d00ca923089acf5f319984d952a30e263c13d2012348e25820ddfee07482a51c3e96e57
z90f4b003f0399e2d6fc53fed198cb7934be50657dd8fcf4b28fe72a483b65f12bfd503acdf1100
z1956225b1c75ea5d080a16f176a48678aed087b45ee79e2e1c8e5296e227afe48893bd70c90402
zeefc2aed0da40a11e088f8500dad5141c5dd8dd845569b60e4c56873fe627f8cca186afca339db
zb0602f84e04c17749e0a1b92936f4f07598ce45a6bc1895a9fd076379707b301b2744b14cdcd59
z8e56df5ecd4e386f18280556510f2233107c94506c77c48a721260a1f4a6681c67a38a9ddb9227
z4e1f5c280451a166e9feafc06f11508c3d19b7bc3779b9b57f06e618ef17a06899ab0793972ed0
z83f7917707fc5653e06fca5f3ecff18118059e6e772c23f3225da8e7bb7fe40198fe84cfa3583e
z373e86c4852f46abecec892870e728bb32f8475cce5169e6ea656d7fa83cb7a2b93bad5dc2ce54
zca75e12355ea645fd94bac473691ec3581009ff1d496572352a079605bb4c4ebf0584314927a2e
z0535289e1cac5c8673cc55f352e3ea1b12fd87588e03a1103c2b1f2dd155ca80b7f19c3c4983ea
zaec48cc189e9f4c70309863157cfbff02881388471df1fc66dbbd65d8fb0b21c2878d8fbf9cf7e
z47f8a292a31d1b5c4167fcad36e38d9a09dc236cb46d3461a397c881d2e6c3fb69666a5ed94808
z0a18a92736aee408184fa9eabe78a4fab020b0754dbfdc105665c2e05afb44ac2f69684b78e678
z98723d819a467494123cf0a3a8d55dfdb8d6cad146815175444b1e1affb4f2ee7e7266a41a1b5b
z696d53663a0276517dc9e4bfebd8535ebb790b7d715c110e249e3b9208584a769dc495b3101b89
z56a8f0894b59266cae60ee381770ee9beb5f45822e6c99d1962871bf37500dc1bc9d7729943ed3
z68102b25ce32a426faeb25877dce135e978c1c57c4ba206b9ea7de5aa654803bae75890b6b12fe
z0ed7036978079281bddbbdd408938f6678064334e81da835576f92219babffabbb22a73f785934
z69b3f088ba111f5d4af933351078558e9819d513b9212c3485680500152b4fd6bf3926098ac2cb
z84af535f72f3e1fb96708359a6990da5af5db40c97334cb7318067b8fcf4c0d1977856504eab7e
zb383d5353dce4290c569d5204a2017201bc6cacbf076e0ec8e65253715deca7d9a65cee3fba784
z6705b0da3656410f0d871e4c2f9c9a21e56b04e782172ccc85563c37a5de778b30bf3cab539630
zfba76940cf731d5fd96b7394f9975aa04d89093c952bfc3f4d35361bab341c2b691a7a626871d3
zd09e0f20910e4ad630bbe8e798b9acb1b0711f9a36bc064948d46c7022c81c968b1d466c4c031e
z69c728f822679ff3f65a451793a334e439bf9d59b5ec65574d27c8b2be6051631953e9e2ca2c4a
z4438d960735c9c0ff5ff991f95317640b80bf87dddfcfca32099c08d89abf54675c25a92c10b77
z067a133a68eac8a5e1f18aeb6cc6e561f86d3821e38f9b6c857b37543f9bc499e0286c293a0d98
zbb05dacaea898869e98cde563379e17653dd685e07b5cc3c5ab82da969110f03dfb8c7063cd00f
zabcbf7663ac7170950803b4c0b0376c5551780f9c0f79819a4447e5d0daa702fd0847712320744
z7995ed4b2107dca5628ce04870c6bae27dc65aac588120f9c337b45a295e23d7f1fc4b239fd03a
z1a5409a5d3f0ea77fd18b3f8ba678a475a3b857f295d34a72e26de9971ac50dcd2b7b7b2427855
z677afaffee912af359e0a3218459b1897434211d843786bc9e9b79cbb371cbc253689bad540bf0
zca3914baa699f6182fcab6d0870c99ddb41944d319fe8d21e8de6c8ff8446224c0192c4b2c651e
z1aeb2967503db7f7ee76e69c86f8f35d0b0f1cd3ae278b7f836530051ea655208f25a775eb9554
z05aa7b85fce56808f36977714dd5319ebc627bc3f8db564f024249e8fb13ad82bbed0156d2b615
z0c3c9ca0383b85ee8feaf38bce3d6b6b5134ce490f9b5ce5ba74f44d1de26e8201e4da49368065
z526beadd2208054a81312f5a05bcb2f555e3dbba7b5570fb04de1070adda9f46a4e6ef2edd3b2a
z69e420657c72151159934e164021377a7e9f7adc3fa0cde81859c91cd0def11d6afdad0ed6c389
z262b27670ef5a1183df598290de6191bc55affb66bde0fef773e904ce099f100871bebdccce69a
z811b346ae129fe0f3191737464de484c5e9482279ebae0e7a65dd5cb91fc880be6be81f9bdb91f
z7c726b99207f6facb7e2266f7a5d21579fb69b65e3c372ee37b6e32334d55addb79fa4793bfdf0
z334d3e863a5365b0be48f096a1dfe113d6f8e847c32b1e02e341ad8c4a239b50fee23f71a7d595
z726c129080881fbc504553efbf1638f999a349973eee5f6b43acfe21f50865e5c2471fdd7a8acd
zf06aae00b52d9d8f520163ede76fbfc1fe645f576f57cdb5dd29e90cc1878fe867995f14126868
z7a1876cd4c486713a8d654c5b2abb421ed768e29072da1dc9f75d49bb34f1761e39307b3310007
za9066574b86dafc71453b793a09e5727d57101d94a22e2937b2170ff69abf214c1d1d49f5d0fb8
z74b8f47c58ac47bda45f70a6284ec34dc8ca79a43d7e1f35ef9fe7701dbd8a15bbef7d589aa20d
z53efd5ad9aec820e78e161de9462e20ec5610d6e12d90382f34dc6a2820bb65f13117942879528
zc17f954be54002a5b9fd99740ebd1b49959468bdc514e401a335b906986dfe7015742555b1b46e
z4cfc38cc57db9e72b0d782e61e3e202be3f176801d7612af100598972233e1e859da2abfb7e4c7
z6c2566b99d19a511ed73431b19d9a860dda858ba67a1c6ab490978109cff0969adebcd8c6607d1
z7fb531da800d8d6378d485ed737b5ae8cb3994041508810c6bb05f2fd1133cb2e4590ba9e211ac
z7d605e5ebd455673e5ee3301ed32c9be39b3c44d77aad54d7eeb4e2b229a8d46bbef3fa5dc07d4
z8c1480f5272df40c694ffda2df7f1d2b41a660a0f8777962e37105430a743ad5ca79f5889f603d
z10353c51003d893266323af30b66db3a9a5f7b9c1158b2bee6ba669afa83bb4ea439fc52949de3
zd5d01753187bcd58eeb338c855e92fef9aec17fea712ba1570649aa1aa48205738eb0eddb0763b
zc0771b75d3cf2506fddf9f3927666ccd4b9a8ca7204075425282919414ec98493609421371b7e3
zc5af223691bd0cc5b964b42b850fd467d66bbabb8ba35d230021049f79713401d1e3423eb304a6
z7caf99fd22a00d4e12adf163597198dae336ec091c87d937c929ca75f9e245d6b86523f7392b61
z32c626164fc2f5a75ced36b6f7f360773d60999e3cab2b74f2c1b2549e428447846a122150e755
z67ada46c9c455f7891dc4637e3a55c539865c12ef69d52324daf2db96e7ea1bb73d4c802d81c6a
zd5b7c5ee6de6cbe511f67b97c937119fe8ffc043ac4b6b1f2c2efc1d2262e61fb0641e040c466d
z94146e84cfdb7c60003edbcf25a28bc4301408bf1273809c6fe0faed2c26fdadf671506b92d970
za3dba0597505757301ed846ae09c2ead7f30909a8c80624cd5e6f98aee8dd55a23b3aa6b454ad0
za608b3f78065c10dd1a83cde2edec1bbda2ee8f5caa11681c9471663c104890a8b51d8311e1c3d
zdabe017db913448ce6d6ad31847e5a5b863b379e6ba157d3e77ec37096a3f937be238bd65813b6
zba822899f67a9a98d535fc1a61d8584218cda623df5f1a80ffc8dd1b1cdeca0a1cd41095228850
z8606e5911f91f642e686841a7ca1bc1029fa57c04cea13f5f2550b5f39367070928dcaee2246f7
zd0535ec2578a395613db2ee06a6181ac61e248e7b5b3fb51ed804f26465949174e621a2cbf40ef
zd46ff82518f9374b04f202dc35a048ebd3e26c03500945e8478842676ad059c183e1fd53d60970
zfa2808953725c8a963e759b3a22ed64d5edfa6cfac3c8e8fefdf3e3367f4168ffd2fc622d4c45e
zdafa73d586422506697dbc62c3b5ee0309111f6b021a659717c7f6352ce026573511c45720933a
z110d3aea8071703b097a4df55badd8e48a798001a0b9fbc29bc0ab32a0cc5cbae96cebf6398997
z141bb092fb7fb504292cae107e5e5713a8244fb7afe068682ea15228753d6a54abcc6c8a5dd3bf
zdb3fe68c6f10452426c3d104c5a3cec05c5f226c6412deab278154ab1563b568a18ff9c5e78d9c
z79f1e543de44da47ec63d8b23296204de06782d8e30035608feccc86a78fad568a5ef7d4073790
z9f3f6b485535e689c42cd95e8b9d2b1cc2cf2c43827d11e8a51186dbcd13e64310fba920161c37
z667a133e04e11fc435caa93b0abdd255b92679ae1516b01e3866bf403384dc84f6f0d14a0c7713
z57b1569ce3310b450207d4d0093828518dc3ab420cbe7291689f7deb3f7b47ce31515aa773263b
z5bdfa64489d088ea965164a7c71602d169c93b1044b4b2f0ce97e121d6f0d0f5bd7cf45791d99b
za8bb2c88d4158512e5def487a109e41a6072f271d4a478e52cae0fa8959a4f765ea81003a509c2
z6ac4e08fd5004cfb3c531985049a9bff531f063743866fb012d283b5edcdc0295a9222262b5793
zf06a6730d772a1fa420386d3561dc6b991f8a63f480069d5247383ef3a132cb785aa706b3d7f62
zb8c73e2ab88c8d5ea79dedca68516de02ae5e7d6f677a2b91ba31267387608a6d6557b8a16ab24
za5d02f7c9f980966801741a318138b1a6def3dc14f95625f32d030ca958628445126f11d654ab0
zae145984573b7e60736be63a543f13838f69b40cf00aea376605cc5eba55221e519032be9ed110
zcaecd510d83a155114460acb12251e870f5e119a5039aa905e4138e848761cb684f31f8a9d9052
zb202b89d25a8c21d695a13fcce4256f13fe9cbe53d6a5bf62965384faa76e60a04fa8646f01e95
zd26c4fde26d52a1de40085bcf4134c1dfbcecb981649e05f08ba1052f4b69af4600ae4d6005710
z8dce3efb88a08622472ee4b103fc7e3f02471bab5fddb2551a9475e1256af6d280a9e712f81cee
z0c2a476921d224137af4c5c69755da5d23190f56b2a6e7dfbcf4c16132bc517f9507829380ab42
z732e1cde33942ea033de077ece93edb56e8b75602d7a6b820e3dfeb4d31a7b84b2c74bf0aa08cd
z2b0c6e324c1973dba0041554198d01b4d5182cb814852f8d8d6aad3ea6e513b511e23e16e05598
z2a933677144743ca5d06cd37f2cc29cc831a8f2484d5413308728d60bbb901c68ae3ce4dc2dd06
z6fd0c9837f88b230ade1a12e6fd054e57a754b5022c06a6f80f232e4a24d543aabb257d17612fe
z0ea339327576c97931405e93393c5e3be3a16d3d0c170687ccec0303d8d32446f4ab750f32412d
zb30617e4fa7eec7895580e4bb933bbffb133548bfbed8402c226e8a83d0c85999bb46b1e7d3b35
z50c3d7760b38a32d1a12b023c28c0cbcfed468072c6b5c64e3e7649f5b4ae22bcfaa90b229e75a
z4752b36b1e9553ac4a5e4fe8d45e2ab052d5c426e8704c46fafe6e9c0bccb8d8f24b6b200c8dea
zc56e05182281c3b86178d1d400173e410393ae641a136dd5e813cff6f0f3e98bc0519d98dff0cb
z8550937195bce846d0d29ac78c5cd39d7b90b482b86200f82c77f7bde8b3d1474a90c5730a3e4e
zc88e66b88f76398ed30d880f3167595f9f8e9cf3e55664e8c091273c7b8ebb1d008d4a5fcb4f6c
z06857116ecdbc1d5bb961e84b0791b5e7e74363a1a79cf3b1a83c23c8a135b99f79150aff23d60
z288796fd691c14355013fe98feabc7df8c54ef4f0a77cf082fd1b94b60c990889cc9618689c25b
zc128c6622ff8efc2e9a7e3a3f9e91136f600cc384397ddc368c0113c05623a27ed5ef8797a3b82
zf1e7ea6a84bd377e22d7a9762219722f0a8c213607d06e8b72ed1873ffe9eeeb25881d280ff64b
zf95defefeff817ab118fdb928ae97e0193a9745a0d42759fba6d7681dfa47db320d158ad3e5132
z8794d3e752a28e963c1158f232e4326847840df6c2134cf7a5fffb8a02174aa2169e8fc0ea4b5b
z7faf435d2ac31b1219c2a9e3224a6ca46582d049a091cb674e7498c848882f930ef9c194c11da4
z4d56ef2efe0b9dfc9c12227a0ef4c1beae47715d2950f36c192249e9af4f7e2f325c2f53716096
z52414f61aea6f8edafb8b4367a80861344943a45b75588023e05e1233a2d5566e96b802126b30c
zc5fa43c9bd766bb379bb947f45cd47089200906ab6d2c1166d29b34b3c879d512163cf15a67f93
z4b06225104b8a2ec6e1c8c43dad6278810f26d8f096a3263dafd8d4bf64143be0fe9b52ab3ccbb
z582c49910b6fd31785e180f78b81fc1e2d7e3739e6be792649500e9f559d4c3c211f3e58df9769
z091867eaf4e49d37d73856522ec210bf2646468f62fa288e36ef3ae2a1cd0af99db1638239e3c5
zbc65f2ed8dab2128765a38e530a900d746ec8a7b9126bac19ea52f5a945b6a6c45b6ad94b4ab51
z6d561de982ef036542b581042bb6b3e3417d6cd619b69e96bf5759aac1054b5dce8d9555748137
zae6cdfa4b970e0e755a2dc823e206dc68e6698ace5ef0807b567f0c8aefc743625df1e7b52d7cc
z475bb6cfd4caf5ace3790a471ae8ad16a641ba50557122f5998c9a669acbb96ac81e13c0bbb423
zb8d0b0aa43c86e3c601f489c0aa88d65dc5ef504755ac4cd8459183cf4303d0d02cd46b93e84d1
z0b8820a18f3e8526f8ab74cac545f3c015221016c9f5c542b4db63df2171213d7ba3ba59396917
z967395484f0c34395b859414f77f9e01be257279494d3d36b2e70dff378c79289e5b292fac295b
zb0336af00c66d9f808e921c5a1f71830f896fed16e2a847853755476118a8765e123fc62283d05
z43542d71d1ab6e2b3bece15335f2850b885f4d92bdd7174528f8275fcd7d245da541f5c0b92fa6
z600e610762ba2514072159f96e29ba0629ff776989beb009ccb99d8e217a3a6d5f097537f2d8c0
z82344391fefaf50957b78366d0d5c854a59c99180b06bfd2d0dc55637c02b86864e70fbf0471e0
z4e1212c5e25cffd3c36d9eb5d59b78f1d2733c2573199e78b136f946d39186d078c54b34318aa8
z2f7884825464a9f0a7e72f00c96284011e202a58b3965bfed0f6bd29ccc4e41f0506785acac29a
ze9e5ea73ef6967466b39e8a196105d89bafbfea3da18a47453c68a017ba591ed5bce8858831ee1
z70412251b4c582a58a962ac2a2c5ade3cacece79ddf5fb992f3abe8102afd59c5702974a515230
zb7d4013a7137439ce857998b7e12cf527f461353d15a4dadcb319ca7f2743453555ba9a43dd951
z76fa23d22594b01e74b32e1381f8d50afd9036bc8c1d609e0dd157b48bcf13171b05a368338192
ze8236e1559941deeda8dbf340367aeac136aee8b656c32e605e3b5c7bac364176bf0fd8ef12f19
z57d844c460c1eb89ee5c1400e99f5ef6e92479c20d15cb88b148bee937a6be141cd94f94d3a0cf
zbcaf7349f11ae35de9ef33f70eb92eff7d055448bdeaa09f4b77379ac62fe1a6a68ea00d1910c8
zdd1972ab445dae5d4afcbabc8365c40d53233b357457322f2e8fbbe959b3da43a5222c0bc1c8f9
z4f64fba0de932eb9c479d2bdfe2679069dd0aca62aadd94bcb8f4fb712598ebf05af978f1dc47a
z322ac2abc1876c152cc4e3513a1b26cd23188d103701bad1a47b4551a87f5dae5816f4092dd313
z2f91670d2ef46c36a544617195fc2ce0888a9111a91a984b21a767a57846234047a3188491bd15
zc3e70d26e449dea3df6191dcff482e5fd1c38a6a2713084e0017c719acc22e715842b70c3a31e1
ze4f3fc2a1ee4665d9d68544d36edfd557631895f5d024f468d67404160b2f8c156893a93be1086
z72b0c42310932fa3b3f54a9826ef28bb9c728e2f75fef6f8915cedd5039e40e7505c961a3476ff
z99aaa8c3bdbc1e2fe6b315ad4a21dc8f31ce6b37331e5194a50c8dfd43c079e1b78ef02e48b59e
zfbca13c64c8c892d6ed2d729fff2d47a389625913ba354f95080064acb4ff922321ede9c4a888b
z4c066ec891b36385223f8a6f791906b82d1ddb87b188414cbd67f8bf6d418989413e4128ec302b
z60907ced3573c6318d0180dde3a62c817aa4f487597579d98971742fb741a1fdf7a79899b2658d
z10289e1bf80630b5c201be4d3027d3df3cb700ee67d00585a2cd69ae879d32c80f831bc21b3d05
zf7030d5dbf71d5a719b5b20ffbe04c6c79c50c9ad571a8ac94f4e995dd487d5e9b26fc95c95942
zf74fe0668490f107d5b3483087638920d406d286716ff6bb9932322fd4bef2996729d81a1e7255
z20596e0e823c8d714f46a2e71b3cd08c461f9c309882944415e5f8c1950bb7c129b77e6fe9e35d
zdba3e9f55a6fffb15d2048c4ee9a207584d0308d6c859b97f02588396d92929787fef664df8128
zcb69b1b9e8403b9dcddd98135296ab1d7e46f62ed5367dce3df1876a13bbe33de57defec59cbad
z548230564cd2f5e1f494a5ae08648db750e18b19b718608f1e845ea26b0a1c56f7173b2fb0918c
z5c9604755fe509f439de21f9bc4cddca15c94af64e246d02d58d5551327eac3d69e32b3010efe2
z0ce25aef962ff1b323126f92917095fbad6ae917df7a6ac4c90ef78c763c3f1e12b7ba1998c8e2
z5cf782c680310b73fc5ea64c264fd2975c90c25525e394daeb381d8b65a8e40303e5385ebee043
ze47bc55b9757a402b3b539654431dd93aafac1324e7507d2dfce208b3fdc10ab80596942034de2
z7fc739307e27c36f364ae4d1188596ee26faf11eedf3f73aa274d0ce4a812210e542ba44328698
z271fde88be969314af2d42f35c8c9829d9c4dc6c7fd656cef34cc1625d42a7cff9149e5127750e
zea45f3e8effd5e696bede143f9f5d924dbf6fb587dd2d5c536821aa7ad30ec654b7d9fed552f93
z240fe1424ea4651f35878f1fc70edc0081952f828222f4cfdfdda8ebd77f6e25e465c595c359e8
z9d4bf41a411f77d4242a8750cec0a102b109a1b9bbf2bd7581bf960a537a1035964b9f7b3dfca4
z1a848b9b59dff1538c02eee1f77fb75600b390f283e618b987201efe1a9ffe3708e774d68ede35
zfda7e17a1141c2df72a1613083ecb844d33c854ade4113d04a69d7151259e995eb269f415c4b40
zf6dc013a218626a5ae38bbd76397acc6176ff20af9cd399732b47676d65c153df8adf218daab0a
z94876b4c1cf36a6dc5d7e180351dc04d32c091812d7c646411e1981c18e79bc5bbf00241f975f4
z7a7ec0df1b7fed55552d46e72517a023c268855f1150e67533a220902ebaa02d4ff705a359afc4
zda7dab8d2118df48a89ada5fc1558a96e2ec94afa001bd5729d7a993be069f54bef41e1c57a251
z2df4e9db89e7f57c59f3423b211d6899a6b3fcdb9bdd17911c7a1a024ae3a779996784c1bec93b
zfff60ec3d16b85b2b406422d59e6dbf71885ecbee4d731619d0cd45f48ffa57b209e0e1bc8948d
zdfcf3861e984abcc87ae7bfc1605712c761177f41a3f30c42558b97cbe57d9f0c0a8d0749727d0
z84187cb958f9182dca606a5ab3aae1418218519487ba099aacde23e2dcaf9bba3e308bc76f8fdd
z833f914a9a921d7455c977595ca3f38fb7e2be65688b1e845bdcb3045ca1f8bd358fc00071befa
z06a926b32684d9a3ef51541699cc6d82125275eb377c7855b2e7daa4499ac07163ff104eb574b7
zd5c12296723b27eaff9e20766220c6a95af505a814f9bc10b30c48523fc45f6386a8fd5f661b26
za6afc6ad2effbfa35ec19ecce3cea221fd78f3bc0165ed2f74730f106d6fefcd4ab566a15cf28b
zb8d93bffecefddbb7d5b752dda03c45ecc6fa2d147f92b35caa5ca5eccddb1579c45ded52efcbd
z15ba661793b8c428761c21fec637a4526a006433af3961a6a44ee6c5d7050cf596d18a67c3ec98
z241242ca3ba83a1675b6218961e1716b74fa5388946f5323c43db41040152e026dac96056ded8f
z36e25f8f0be169ef67d9d70169749f3e818ba282ca7a01fbd6538f09022022f7ed0c0cdb952e7f
z72d8e371e5d3fc62766e4444eb0184df3f4223e569b406a6b17b530c082bb045f4b91221aa6c99
z2020d1d352826577d41d19c70a8ca07c630eeb504d6f1591451b15df3b16657617919e2ac9ce0a
ze23c0500f3bdd16a33438791aff2982a2bc76e2246b052e447c4ec4bda084c0e7f4713ff393d14
zcd509378873faebe3db862f61d3d4fb4a2f3283b57209cf8ab9e6f1f8e0d3e78fe3a5f74c5fb25
z48e54d35667c6a5ce46eb1d274454180d5cb9752e25b80c8590038eb5cafbf27ecec1d85cb85fe
zdc27a5c6e94ed114b5a0c757ef1a5941790e84c49104990d66fd926d8a971e1143e3fa13f3250a
z8ea9e6e9c55af13fbc9da12ed7d4f2ccf3c22698772e3f47719d2622368bdc4a841f133d8bb997
z2d1190747ab3673b3c8042cca4a6815ab3aa8a6680f7b12eb2df63b6e61587f62bb9b117c1bfca
z1882f2ed091feb2c74ff2cf31a6e82c7764904544a239f92741bd8272a597df7afcee2cf91157d
z43e47d265b9a4350d48c9c28aebc0701637a7c7176d1a1d0bf94d09d746f9a91e73626b52abe2b
za227b9a8422083cadc8e27b7f28b742a12e9a8845ffcae4d7f4c0e2f28f5f6dea797dafb0f3828
z29472093c3508c7b0d9afd40df65bf08352dd8adde95aa04c5f4903538a0ad7b3030f9354db081
z4db7a34d6df9498d0d291b8ce3f476be272f9d1e5763249ab52496e1290f165c0ecc7afd8121cc
z3387170bc5a173f0be51833aef712f1db1fd6680bd7e131c9031714c23621c4f01e9609cb29f78
z8adf44581ae6ea36a5b4889e68a16a3fda9843f5f0a25108283500ce702c06bbce89d73db3f30e
z7251a906da7f637c749cd5f889df5f427e686fe98511af4ae680b80597d96ff615b0fe76b7c3d5
zb150c41060df61b431351131cf9e819bfea1ead5e047de4714f89dbc06881873a56c53b1aeb8da
zb35438cd4545c8caf2cc08f18deb3f07a8746af3b880ef9fb2d78a49995a45a5a643c47a8036d0
z843f359efd0383bf904151dcd3dbe001a1d69f57e42851b71c3cb713eb00c657fa643ae8a3259c
zb9f62e9b4d17616d8467363d3b67b5fb7b5a58a921fb8d3005cdb25f0541d69d9e0a812b9090b2
zf749b6c4080fa518aa72ab10da6ffb2d69d1401a3ac75fe5babe7720d5712ea3e54ab699e85069
zb6127fab3faa42b1d5c68e3da7248d082e6a5f70daebfdc93228a0f400dfac32c14692463e5878
zb095e73e1a3a4be0e695a049a72ea093daba57106a3f21bc05253683e657defd163dd2a1ae9396
z7f1381e1446a7b8a4cc1f455efd479355ec0b33d650540b3b3f0b07c0a69a6cc5d1c87e9d7e949
zf4e24ff79b3f0ee2cf9920578e1e5a1af7ee1c63061e1ce6709d65e6483cbd364825af601b51d6
z238be7e7bcaf3b22812f1e8ccf69fcd5e58bffbf5db9815832bd585ce611b500621affd5cd8294
za391c4e13dc079568ad94f5da188e6d3404242a858dbaa467257efca26a6cbb3764a6c44e8b231
z3b9042789ec8f647f7b724bef758f9376d49d7c0eafa73e54c94a16d4e75d753a16a7b97ec8dad
z9dbc3082be0da026f4274e8a3b2fedc5366c4a7be14552539686a383aa26a455ddd1f6c8e95389
za73e1fffac968c4a54ef7fd422bc751eac335f461b1dfe7f00477aa9cdb22b743519203d4aca05
z0d1655e7a6b8ba667378c52709da3b70d7d8b153cf8be277fff50d785b5543d737424ece5fab8d
z55bff4ba8e3676ff97ea8caec28aa37cbad3188f84f762dbcd9a9a4a9d8fa0c399fbaf7ebc4101
z84fb0a126878200f9ea4a965a8934487e6c46d49351bb170f58f1b761abb6cf9b0e3f98448dc15
za3ffb3728d8d83fdb6c68438c923a7d8923e6f86b956ad76320881fa3e233279df927a92272bec
z806d982a3f9c0bddd44047543705030c35b1960115f763fe5d9518b6d58f51bb3b1a0d2d2d2def
zbf0d48e9d70b53d336b4b0c7d708e743501d62e63b419726a101e69d91815f5b2f149f9177b040
zd2b25c3c2f4df510cc6487471963aa2de9b8918878c9cb251db34c5bf7759b2f0e231412ca7ce4
zf5e77042534871cb714c69b381eb47bd363f0e0519fbd49238252949270c4718388d5c42cbd513
z4c705ab5cc0ba8db1dea9a9a9d47b6f536e01860477fd1245465d799a29346d71ed2e5955f6278
z85e99075d11309051d07f6fcb69f12806d293bf0123620b8321e889ae94dfd52e19e0288c078b8
z518c9bfe344012bef7233d5c7d5fe1a1bd417938c22f03b9889fd1102b88848623be5b55d00bae
z16079bdc5f56460b5dd84240332fa5e6bbc4ca1a2493567c7a7a6f7cbb8f734ed332ccdaeb77f2
ze7dd476a09b7c6c534232c21fd42ae2d8f9e2c620e514a03c3961d5f25b5af5d12878ebff4f276
zb5b0597d122080d7b462937ed7df7041db13681bc379f67180b192cd6278aad176f970e679cc52
z400923e0971e18553f4ed7bf53642769439c99fcd5d22fd8713c82f2fa42baae1988e846635487
z640a00d3b55e8eec760b66217901c98ebdfa36105a205f7b5a87bed85263697eeecc01c69087cd
z49c0e23df32fd27be39ebbc60d4374ee6f598f81db356287142ced675f4289620e63def816eef5
z93f75a7b4f9391a2cefec014128146c6295a00692aeb5960ce519452052fffc36a668c7f406e2f
zade5e1632762205812a18766a2246c98123145d16f52bb91dfd5f2575cea57346a57c0cac36722
z437571807e73157f6d593d652e1fccdf304eb5917a6acaf2c1845f6e9d39bdabd4a02290a0b005
zd9c24a68d6fdfc9524c5769d23e961d12206f11b7c8f1a078dcc72b11d5978300c540cdc4df532
z466b55ccb2d652b2d7479c5041e27c685967b6f3edae3941d89529e9c0692f36080aaccfc25507
z60969ccd45e31170e58574c6d8d1c46056a8c3f40fd927f695ca572f3dbf73ac4fe9d94c0bf8fe
z8aa9bf67e0157b8285bd04beea1ab8c15db58c436ee840a5e217743af5acb677ee930d94415c64
zd58039604df392f9decebc4f5688c5dfdbd905cd44ec960d20412d44f56e2af23834e7535d0d07
zb96de7bd7ab2f72f4a804e6518251638339d2acf307fe3b319ea66c5244451926c34b4bd8072ab
zd768af800a5831dcf4d48584f3043443f32238c696c762bdba1156a4a64c77756072ff6e28d382
zeba9cda034b663a2a69ae318a3f87d88946af68840d730f25d204feebf355da37f72f6c41bee1a
za1bc3efcd837246122c53db997ba6165c92d4914c4fac5327313ef9b2fb0e9b23b029514492f04
z501006ec172624acd86fc39faaf07278e5f35f577f1cb0cebc2315b3313845015c9efc5538fc14
za896b2273ddbd691406fc22c1e1fa919c7be231462119e07b228a57fe94e7cda2dbd30e47a86b9
zbf90acd0f173443a7e1b43ec7ef688a870fc0888c44ea4a0de5e290a0e1b2c47135f58c9b33418
zfdee4ca745792eaece64dacf73b4d1aad5267cfa985052822dedcab5529c2fadb1a4a48f24199d
z8af1af4cff6fe104d4b0efab1de36655313972a2b9974a039e28fe158b2e293542fc4052c6d7dc
zfd0ab408cb9cae0d04dbd92b7222622de3284472956390aa81a5bfc543bd1a3e170b2fd79f80b6
zaacf6d9b8d791224609eb22377d08b0bd66503730fb4412aa6a96682c010555e49b33df93e08a0
z69c3f0a2dd2f24aa2cf95928b1a5de6d2551a30189ebf2cfb48ae5f4c782b203670d0769c21786
zdd00d2b6777cacc1e644191f8f17f2187510f72425663e6d00f246309cceef7d751fcfc8d0a124
z95f50e1a1fcb65b38c0ede8454161b27794158a4484a54a6846b0397b34f74a47349873473e774
z378b6a37126ee38dac5a4021530a5cd97b45f137ad45f062da8856f41f32c2a8f50a7febdccb35
z8d1e032d5acb0f65200631c2c7028de93e8e1f16ef71ec02a98b42f86774a89918e3364030244c
z5e15018eec64f094d68c0c7a28d17ef7576bed9a2b5b692557504e2fff4bafa3b7313d865586a9
ze74c3997cf7921474bd0e47d4f68d847cfd78c9f4ef10846f4d4922b93c02dd5581aef61c60d06
z4254dbd3ceb19997d678ee297740e57f8167221d622cc79de85b9cddddfe43588fa6a4a6511149
zb2f950ef623acd403db1e97303558f1a0badb3f1b13f5c0ab20aafa29a5e688e01188400dfc484
zaa9694f7a913a0fc4d8d85818c19e6ad2d7bc9b81c808dc0defd327bf9f362b06ba75a4a6b545a
z2a7ea4c0e49540f82f34929f84d4cfe082a5ee54fc9057f8fdf8d9a6223387102e5e5e94be54f4
z1826bc43698e29d89cb35c17549c9ea160462b4b6a883531b76959fb29ac26ec8a5b6129334a5e
z78d9f9e960e740bcd9a6d7a3d6931ed2c06075e92bba1ff1c0c245085b12d0edf5add04b56f6a7
ze6c21a29e75f3dd0d2929821d4209c15faa0197c5816035abcf841c64f7da046179bc3a05e83c1
z814a748f3e76020e3c0ca9d4a176c3c212dea687a29a41708127909eb046e5395c36c6a19fc4d5
z67d61f5ce7fc71cabe8d6bf87f55760feee2fd5c0713b889e4f94eaf787b1a244de7e79b984ef7
zcb162996c490e7216245f48ef1b70b92bf9922cb68104eb978701d1bcc345f06ec70023314a005
z60b0544747f60bc69b9f79793f54a216716b3dfdcb6ecc37ce1bbb0b1cc5dd8a6eb67052a33e9e
z96a4ffeb07c903e4d8199751fcc12a33dfaf635941d40c1a899cefd9da0ef93aa221c8b37bee39
z976b056ccd51d31e8a2605f99d102bee4d6e7ae5e29932781b6bdd5e1471f1bd488678efca6d3e
zfd9558a1dfe666b0df5fa73ad8c838d35284c8b068133bb863f3d519baed8b2ce52225ef546f49
z6bd5df304630fdcaeb00fe14c5c07648a0b566d7193cb5983880e7e0b56ed981b97ed372868dfb
z0b10d20712395bd9af3e6c2f95419c089a0a14a1d13b7610d898d2072817f39878e01fbd6b1444
z209007cf1ef36ea4d8908b8f86c594c9db82f2de485bfbb88c160bbe873cc54b77d53fad32f0d8
z8ff00a282b4ea6c731314e55c76bc3890e4db2c6859fb87145045c09bdcc63ce35eb09f8088216
zc2b53f5b98181fdcaf43b0dc59e145f90ff6ebacd21a2fe515b0c788957fe05d58aaa53a4725ac
zbd86b553d8849b68e65618f12fdfc140ce9c212dc021a3532f06ae564eebedf4af30b1e0b4c8c5
z41cb931ebc947c10bdef291e7064b8d38a840190701e0263827a66ae7cd2e22abc7322d293c944
zf473384048533cfa6f63c02a38277a9f901b07954f84dbd0943e9b96f407e0479271030d1607b0
zebed932dd9c7d572c4cd5fa349ab2256ef77dd42a2829656c6ba6033f97070e2e1cd858a69ab42
z920d990ea4efb2caae3520cce31c777b960447ff9c071b87d53c06d13f1c400b1512fa8f2a8129
z1afa5c57195a52e7c9618ad6bc7f2332b8b1d39526b9f9c5c815d33decef3ce980aa5bddb1d725
z63c78940361c0b62f362cb83b29506f8bf877d85ed9b33e4b207cbc9baa288c97e2d5bf2b85c39
z5737f384e2bddc4658873e46d5178e2c6f01a8b076356c12c479ddd206645d35d9026f7813463b
zc18db9d0f604a2260346f91e8afb322de922184c0ef312db81933bfb65280a660b0a59e660e1e4
z14e52087b38b55ba4b79efd5bcb6d93d8841443c7524fc1fc12c91a19591a34ad5b684d798634f
z8a7afc701831f4891a73c10a8e4ac0ce0fdc66d4d5963aae834f625a797a193626a4a89c527fe6
z904d6e428d30e81fcd8702a30c835fdfccf4dd400f24e09ffb5a4d8e84fae367b037235599709f
z3669894666f4f08994e5ef06328f14b7d6da610ad84b9adcb9dc6997a510350e8e9e9ef16fd407
z51ef102824e8fe7502b05a5f82053123fd694e860d253a438e1e916035affe0666ed1e347dd71b
ze13e5f743baf66f5a40c1ac8ea93c1fd36060cde19bf6dc27fb2b190c8d68e47c0f212b40c73eb
zd0c9e0ec501d4f60d89b1120fcd739cd22fc975d03b6b27b1218c6df56127dac7e8854b54ec0ed
z620c705fc8c791572645c7e70704dba00d7421a73bc5aab4da6068fbdda6f7502da83385057157
z9b9e975ccdae4288ebd3eb8edc3a29264a667e65991724d90fc88129c100d4ca62eb89eb8425dd
zfbb7dea89ca5fa236098cf39c340cbbdec4b40ae8b060c36ee6210c2d68a51942346f4a7731207
z68065bd6f7925f8211ae454abe5588c3da939dc4f9af2c37bf17dd36390a1216e4f0818ee64687
zad3b83be12a10f8998646e36fa9ee9adc6cc49a444905fdf2ca0affa077d10a07286f1bbd9addd
z8eaeb6f7941c559851bff11c99b17816a306e2160bd20a0e3fdb849d64b0a04da1377a3d97df25
zcd41b5ba4a5576ae7ea620a880eb8d67ffe877c87c7fbe6ca1cddff6eccc826bb6657970650a51
za3f7044ece5e71d49a6d92936886d752f2c038d388978599eee74fffbf96809d360d3bf69e7c29
zd0328b615d0c8704d97a8e8bfc615fe8a832169f66acd202e9add1d4096f465115fa949d23d129
zf1871bc182841203773c88db845ceb2e6d60c6a5e0e61a5162f34755f8029ec06da5729c324f51
z85febf304ee873d233a3f508ebdeefc3cdfc5064aaf6cd81103a0133500765ae3c306ec86fe3c7
zcf74aa9cebb4d600f635052a6b183e0e6eb158224f12e41083cc30f12b2950095c1ccd8d360b15
z0b8e16d1f18ec4f92cd4bf94d32a38f751bc2e99efe07781673b0a4f7526ba429dfbaddeab8b30
z98674ca85e62faa978a79a0b0f12d18ee22fa6a41bf82ac8794c29421de5dc289e189c3f8cfd86
zd7388b6df5966bf3f58b34abe7e0fed94dc2f3bfca29353dc2b2b2f88d3d44bbd9c4b778f81c8a
zb5f2f28a6d6592d31fa0f026eaf5f4c6b2768c6c3e015aef0a252fbf453d3149c20a2f5605fb26
ze597493499a3caa9cc09cbfdd0f3b001a2b4252d1ac98e0a3dbab5a89cdea289055dc62004587c
zcf66c7955fb4e1f39cbd688043895a13782e0ba5e8f56e924363ac1950ade6b900d8e2c8a23190
z1edb8d83d82ca0577b6691887c7232cf2edc64736b0a3aeff11a024ab337156ae3e1687916951a
zb1e2c9af62ab3df9ed5b1358e7c9b3063918c7c26ca8bf10d67df6cd657846da1740c1bc89c2b6
z63d65c0d7cb0bdadd497a13be21071118636b4b527e9d023dd47bf9207a2bec9701c993c0c44f6
zd56c9e1a6077078a40fe9387f76cc49d8c106731dd894349c71f337343013d26ff6bed6d79fa35
z0d2efdb4ff4ffc210800c52f2b6b86d6dbfc97951d6720eca5814c14bf1881e57183318646d646
z1ba0ea30444edbda033843ef19b00775620c988f973a8041b67f92bbfe226494760f4aa0c1d149
z8c927596622324c4efd9081f4b5569fac0459e9992502cdd283aca5f86d12e60984438c9ab6184
z286a59bd8fc8705181ccddbae6b578365033cb1f5a19e3513f3147f28b100a99a4892293aecf1c
z2836fe7c62036f34747c2fa9cde356374bd9834c10b994212a056a35b63f4d995aad1e0a8fa14a
zf85b39b53be09778ce717e6e386c3961d6bd45c6e35ce127c6fda12e4759c5878cc8bb35ec7193
z8afa649578b98d91ffea7c30f776d28046d25ca7ebaf25279f8a9c05b1c3082cfe7488d47702f2
z03f1f3235a47bbd655d33aba1c47e268e426e31785b19b9c84f95d1216189e10be4190fb749a0b
zf16347561d84bb536358caf13d3c95e8692268df4cb6e32dffe875a59084a00140b57d18dc4af2
z75e3008d983cb334c0fa03d8c6f403c6b8c4609c8248ef24e446f812ec61a50695cdfe85301582
z41a6314529add4d5e4454f76a62d7564c1e691a919e9683bcf2d92f0767793c874a899271ee5c6
z7c41702cbcd839bf3f962150597e3e1e576c4e94754c29ac92e30116b0b27c6f2657914a4090ff
z6d3ea32f78b0309b6909576e4609d92201ae1d9dc5e604b191f737a71d3fcff3ba5323a7bea698
z1f1609afc07cffcaeb3bd8f5fb53d89212783da2360b1d353302aab576dbdff384b75ccc9be5c5
z62152568b11dbbe986f3d16f48d0e0748cdefd2dd32d8bba19e5ff6998175b38437a28a73ec706
ze9549ec4c05eafcfd6c7ba18c6e3fdcc4877e399bd1713402fa01ed141cc92a1157306f570b0eb
zf23743f018f70687c7caac78fea3afeed5bc1d00206282c7bd0e5c9817a0f9739490bc76aec2aa
zfa6fab60e38ace616ff023b84b990cd3cd9902ce48aff3642a97bb975401bc76df2b83856db07a
zcedcc9fe57eb9d1bd0bb02912a0576d4036250e6ce17ff01cb179423bb54f5af811cbd3d2decac
z3b82b918a3d27b83126563c6d65330f23ff4a9cd495acf9912b85e07ccefeb96aa0cabcddf52a8
z5cc900e1258ff928aa37a16dde7c7fd2f462bc6cdf133d0e97df8dee60b9cd30219bd9acc10208
zed09d80c8fa97aedb86d5be363e38af107a678e9e2cf7ea2f4d9da40ee62f90dc18f05dad74698
z6f7b5419b9b3c78ac8dc47a1a86af0a2e4ec5ada7b09fe7b6678dc7129bfdd283f4e5959c5ff96
zd8771274f53337c2803ce1e9ff2ccf0d8da3b0431a13ab5ca2c4acf127d7f35aa16b466fcbc7a0
zafc72a7d284f0a3718b00022473d5e5bbab300fce6539d629270e70646e05dfd06acc0931ae0a5
z8cb25afd9951e120a9583c64dc29efa1cffab7887b6da23c378e1fe99b44501a2f27015662e4af
zf0e6397d42817ee550e19e16166519bfdef605ce4e735435a7a24ecd3cf4eeffdecc719492a054
zb23f15c90afe0ef875f0be8fd0073894b6eef04f818457eb7f046d84a159ca0156d947a34f252b
z2e7c86ec8c56553f89d136f4f75e14bb258307b1d425e44e2d43cb3ea43778b586b377dddea140
z1afaceb829679607f4fc0236b98ca030fe59b6a21fa0aa529266cee73c4fea3f1cf0e7007cf824
z6492e2e35f2b7ab869f3327208408c829c30c3a6e27924129fe735313cbc14d4cc8362d8dd6577
z718a6c462b12d59f8270e7342e5529ccb0f1cdbd85bcd71a2c88b9c285907df50473871ba69eb6
z4024ef2a9932fe8e143058bd442b567971560ab3a7a2a9e71265ac5ca558101ef101d93791485b
z8904478b488de683aa1e178b0427e32af87097dfe16b18d7c48c3d72c408d165290bff33d4bb7e
z1499470c79bcf518bd4b5cc6f28c2bc5aca5570af4d19d9df6bae8b36d0dd65079d37795df7016
z72e3ba241b5285304a9bef6f314c34d69a0599aba71ca9c7c0443498b8cac0d43b9f6749348388
zf7aae52079f946d0fe81a44a0476d7b185a2e42ef789067f1c9353d982b0ecb80c004a27e62ee0
ze3b62369fd4df3fe4ed2dbd64a84b90eacd5f88ab5efc3b0a56ea78bf2a95d2125677be20075c0
zf5672d6a97b33a44935852dd0e23ef5e62733fb71b2a05ec207ed6b2259846026bec0fda1740d2
zfe03592396ac480dc48455a07eea7653dbb25dd2b6eac9c4aee3145c01623204e78042f84fb25c
z9634e130d1e95b1c04722e15750b3543aacd4e6d3790339756602e26a662c04e9b3e5763bee81d
zbb3e71d9a0b291e997ac8c395e2f1af492a61b31f66827d1814b2416216ea9d582c5cc481a6217
z5f7e665f3db0aa78e0d804860b92c97e450ce83e3e7f6565ac98b6d55425ce61cf777d05c9c906
za94a74850ed850cdfeb481bb46a6d1a6ad4d0377e7664f26600434a4ba299b8fb0fecef76b52d7
z35825d2f50eb8973398a25859dd65240f3e20303854fb2c1261c9bd5224083021c1154b6110e56
z76d6d0fe1124ea709a7d8fa2df75fdbf8774b350591c3084ca714062f815913701553ff6aa2bfe
z9dbb42523620a034036acaebba40e2b9a2da1dcb7318f93f9fa0a0abdced9a9a38e49b661fd4db
z0051424cdf92ec94a4382b80c5d8603777d1a52a0ffd1578a2032fd9ea9ca3a2d8d9845c799325
z1aceb6243cc35e4a25b369b8322206cf3e783c0d64d236e325aad67d77cf27e6c48241af1050a3
zbaee6ce2d23c523a13b94f3cd7aa5463d32b5389129306cd895c1a7338cd97de0c31674a3b8c84
z8edef39fcd84fbe4013c29ac61ceb2a49ac6d1ee52c83a7aaf7e85dab59ae671e70a7ca321cb70
zdd2fe3e5919a5ad57a93356c9b48a073423a711dad988c32145a76c55b35f9d5aa3d7002766cbf
z2f5a0e28f1d265946a8325a3a4f3db7a3d0bc812d8c0b97b23506aeb52ee8f15f4836e2f684e97
zb68ebcf5e22c5d6073b586134d830756934b168801dbc2ad6ba74cda54a9d1824e095cdac811f3
z9e5302b83910b96df3b54d4655295eee54b25989b3428348a0cd41f9a32dbf8b6add886cc0e2b1
z1d2d77ec2ebc4d8ea6023f576e72d00f19fbf3fc1c6353231390c532ebd50ae67d22f9c8cb8ec3
z7f53c56344d3d3623d425c9b35dfe496bbdb48bd76baffe7e92cc27041243c06f74f739f64e9c4
za0c24ae75cb280b01355bac1557e1af15befe965b4815a8c57f4d72fb1ef194345be66ff8106be
z656347cc4e8475914d3e42a5a1dbc9e6073bf9a5d5052bdb692d2d73ecdcdd8b1f135b07a85024
zec0587b434844e0315a93ad60d23e1152dc6b2786d5d038c0d5fb07e748e86d38c9d565af57c88
zf05d0dec6cbe4803b8ad3e7c769c0aea048d94a74f0c2c4ab4a00071ce6c1ce7ddfea4fac680cb
z48de28d9b37a66ca79ebb2bd4c7d0971cdde734e64462f20e0d1326121a43020ef7c1b37335a6e
z7361d085016794dcee884943e8bef2e7636d0122d639ac0c5de90eb73c66d894d6fe80cf9de397
z0cf301a481cffb4cd16db33378db385576a232869ce63970ececbdfba194606dfdbba8d6c14970
zc8d328b42f258b05d9f0bf3dc632b6fcc0f641ce8b1ebfc1ddb8513b0b29dd7ddbc76712c195ff
zfc28e3e2affe0dce57fbdbd08ba78a7c0121aef18046e1e3540cccc066b9d1c444e714b89a7969
z54baef30fe97419290b0cd247da25f69acb474c6615cf667c1827a851271ff70d6c9fc236d223c
z89f61eee93bbcf1a4189d367e9b35e35f57907f7fe8302a932c899f683e4ebda135f3afb461ce3
z467f62d375cef8e867e2c7958c5da17acc4e078e440bdb43d4d808fbead41279c2f6efac3097a8
z417b334d9040fc82bdd31e8d7a0c9417957105432d14390d5e91f56b673650d08e6140d1fef8ea
z1e582b34aa149decb4ac3982de6aa93dcefd218d72626ede68685965932244d1e83a3afbd6d09e
z9c420fa25522aa45fc5aa06c7dcc1997b0c51d5aa556f9fb9ba61ae886ed0c1d5002556ea7f77d
zedd060a568852c1de46dff5022a17b90eedbbac45763f577d163ad4bc4c2ea4e371ae2d98560af
zf34d3e056929a541b03979f4f38cb284c22f4d5d109f3d85edf5cb8b6e6cfa259026abdca727f0
zaac2054c7937d459836624a63833b56376fd7674da3ed3c907e0242c60a32a7b628cb6e9bd4265
z34f6255d07dde5247b3840aa5732d1fe504e2bd122aa3eebc283d5626b2258b94f65568e0f3385
zc8f21e4cd15a7c16d8591ea87f8a6fab2edbeb7fbcdfd18529e67b77c143a43725306b7825fe24
z460988100581fe2faef17d0ea58363fe797b25724dca40964145d626d37cb509464a3546a17db5
z96abcb0319534a8e05c25b0c79ae6748fec2138636bc0676450d5d741f19bf12b4a5636d08f061
z8dbef2573fc1afdd6e5cc4d582c7d3f549aaf85b6a94a3efdd291c235bf474a81bf8b357987314
z69b83b4914e7274e1f96a2786d1da850b1038c6d8a3684ffa30adc9849411a2abd5dc81818ea4a
z0bbd42912a3f8645ef74b23975861bc3b5c0271c9284631a5f7933c4194253ed2fd21900151e15
z8d9a4c9bbbd9571e9c6d56be03b81a35912d8891ff41ea9419beb1d42454818f4cbf7a9280a3d0
z8a0fd3307e5b5f6f5e2e3990eb20c23795c4df531ebc1f672ea1fbdb5325238676ee661ec70ee5
z46dfcfa6cadbf4d9efc3ef6e8a89bc089f8ccfd7c17be0abb1cea1bf102be74f44a26d4467da42
zaed56c6d46d65f66d25bdb45db8a1ae67ca48fe7e47494c8f7ad99e080338e72f9656604c9e261
z1ea4763a66c47a8c04cfd8a57178e820fbb78916802cd7e7bc0e2b629fd874417e5c41e25707c6
z15449272b97500979b46f0c9c2cbb5bcb3b3ccddb23cdad7fb0cb94e37ec744036e9487e48b271
z15b16a26dba00cbc9a3bf7f473eed734fdd7c30deeaaf4c47906e2499094b946df97edbc4685ca
z98e1209aa1bd9aa48cf7c175cfd4ac012402ce9cb4fb43568b105101c42d9d8125fd5a55b59567
z3b6944747eb5f1a388d0c85bdc5b3c183359003db17d2f24efae92372f31aedbb26419587a2b57
z7ecdd553ee22d3fb7ed801d1d890fd3e9553dc089d3b0d4cc47902193f1253fcad8ebaef10c890
zba3e0b24cba66b4753c644c2ceafef53dfe341dd002ff360c0dd9ca0d8e95d736493655a2613d7
zc0798e52eec50db9bb6f7de0bcd9c39ed4ba518ccc0248a2e6a49320470dbf117ef19fc5e21383
zcda7af1053c4094d52413859b859700487cecf2ff7dbec1a63128bcc622d19833c318bb647cbe4
z6b6a18ec50a6bd157db37f8a738622b5024b7d6e08d855374bfd0422a2bc99625a3eb7e2061b6b
z955ade6b3801fc874bd07ff79aaaf327f8d305c1c48b2ea5404f8629dde0a02e44d63a8a24f9d8
z9ed698150a4f6cc9e9a9bd37ef9fb54050aa1283a078b205db1ccfcfe0e6c4a10442b381d8ba82
z5bc46d5ae6d86b516ef7c48434dabfb9b7062d4f647845c556eab56c8455f664e6afc097a5367d
zf0615047d5fd9674cdf9993164d2d6ff45a30e652b357fbbeedb7f2db36b280dcfa1644bbe8536
zdb05cd69e1220bc20a1e2f3460f1ab956c4b2b9a296f65034d4608d0467d4efafbb89391e76221
z2d6ad390f2f815ce291e81f1f901d3ff594aecee67a28cbc052d56e78b0bfa76119cfb7be8a363
z65565ac46d2fa17bcc756baa87b27f0658b7d06feba9b21db85e1306806338341a2df4d25b4f0f
z0b078850a7644338ab59f142a05945b52f96c7db1239ae9aaaabd1ea98c6934c890b6130624769
z14882cfe82983707294e5c681631be2acff2541b251c796d0a7bc37ef45f7051969d1139b9598f
z9b8521efe902a1aeb55f038daa16dbcbad606ee6411bbbf8d92a171d25eaf9b1b38b9cdfb80b70
za42b8496d868281460bb0bf0d0cf83523e4411900e66829b2a7fe3f0fcbc062ae58345aa61cc19
zb90c517719241e96540f9840b159868a3447f3751b9ed946474f0b03b6f64c890b8ca5ee3df55b
z9c7c18485f7065a9118a7f812e2f49c80147b2c3e0808f8139aa2521e7ac861600f294cac33be9
za92f91007df1d335b25a9fdd91d52819a96d60320ee087df62ef1a6f5f3018503a84bfa0d0ab5f
z4fbfabaaf0bfe264bf82f236aa4a7209359b178cfbf36c476b34000a081791e9b459d35c3d81b6
z6eacebb6ce0e5e4b9607384f394d2d8b38bac9660122d0916ab3df12eab2747be3aec7b4428fb1
z4048a7398a49ced7cf83dcb79e23735ae35b8adbb06ac274a70cc976c2209d663f4e2d07047cb8
zba374e54e76667a600043f1e689b22f9001dc97ed3aada4be31ae4af9fb6de6dc2229fca2db6ce
zefe783c191d8ec8c847192ea1092ff7bdc7bd584526203c61e3aeca2fad8d0c977698be6f4237e
za49b3b7d9401a63cfa4d38e7a0cdbe81502a7023238eeeadf0672767b79961cf662882bdaf2961
zf4548ea7579a03c9972bd5f5ef3728e2b5c75351efccdac92c6b3c3803fd9fa5db7deaa903037c
z6764af9454d7decb97d9087cd89799a07d5848f0d843fc2a8dee061274d4142af01b5586ec31ea
za3694a30095bae9b818f49c45d5e347e17be89755870ceee29b86c7d2338a48a2ff320b2fd8476
z4259f3004fbcae370da405cb4eb383e4f2efbe0b32545a076560740e25b42fb5657d06b616b516
zda737da9d203d8d2c4bb36b2b079b19ad18e0c34fff9f6907116e4cac868df47ba415b5048c641
z888e4e22550c63ca5b1917938fa7c930774cbf685ab79b1dd459dbe9f7ba8b2a8c6be2f4ccc571
zd40aad5b88310920760f265d4a8abce8628d857f564b4c05ccbfa49e9857b4d698087beb1eac73
z24e914a337fbd7e9ba05ad07d20bd3d35f05dc787113b7290baada1dec28eb063ef9d9d1d450ad
z7d9147ebe0fc2a2bb6e909c76f0e0c1aa4a97b1ac960ae7c20373618bbe88bd4d32b533670c833
z71e6e85ac6b63038e695192754919ef30c64c054a2c8cca354f591c651d11300ba1e9010d50b61
z6cbb8f4a055498cb70998bdbe2fe92d6c86bf4fe16cf17deb286a31490ed23e4964d44b5a7d6d5
z2a75158cf9e2424df78d293f8a1a434a2a21f8673facd2c7abefe0d564497b551a677904d12651
z21949c7f3fb5b7ecffaa384c065fe0141770699f779e2049c7cc3762af986d291b57a37a718742
zfb203beb2157c4b45ab426aaf5ffce8951eb5bd3ca69f4c898402e8915bb549fe3a83a6b5c1c9b
zec7f5dda2a32b99de4d599cb51281b421303ab9570b4ede6399a0aa24b383e483a5126f4c56c34
zb4443057cd4b9380f7fefa37295b92761b45bad55b014b18c43d40bde8d7d761a3f67a75cce3c9
zf00d8d61f847e681f8e3d08d2840d96d6016eabf745cbfc9d09d403023068f6f3f6f9250fd75be
z1ce0c231ad200b0f66b62d4c3a9c37de19c603dfa9cdc67bcaa868db89f92a35cb4154481d4acf
z53d9758f5a33c40c59d7aadfefbad71170aaf179d7abfd0f1715df54de849b2146a78ab07198da
z25452a644602f29ae455e9abc7ef21128260d6c2cc28c191e6b836474b01b0afb29332e94bbe26
z4cf0d61fba9d499a7aa5e2a3ef76cba894b236d65543c140be0d7761bcb006a141300733152e0e
zc5e370dc88efbb6de4d2e5643e4a9e15df0bf91030f19e2e9df4125b0bb15bb73edfbc891fcc1d
z3da29f72dd5e148ebece04ca3842b6e2bb6aa6644356223133c2a0c2d887ff6344e9248c95fe3e
z84918cb23d17e235a9015fc9ebddc611a5f2a0dbc19a6bd4387e64862ba9b48512a54ea085b64e
z8a9b44172cead58babe237b22eef4e73f847545652d7a85c0c5018e273e7265c458ffff11c05f4
zf25165a036bc82436d0c092266c29e981ae7bc47fe0a899015ee4a9fb4c357a390647215d5f814
z8b67592a01098cac519223972b3f1897705753b52d352f54dddcd522515c4442ddb6cb97f77cea
zda4bc9dbb8ad7e31e3d429c941c46a9d05ac717aedb7241fcc762071d94823561a204284d9c504
z22efa1c121301b82df1d3a3f1d5602d4579443a3594d67e1b8df99c6402da3404b4cf06426c4ef
zb821f9d67ced4b53c94b5f01109bac49fa5285311d50fa27c02e94f638f664f7b8fc712228f840
z942bb07c2b9ed5a4c3b5e6b951a4f52ec54cd0d1e5494421e2feeed259521224c928bd8fed6f99
z23c952a6e1a89965ba9eaba0bccffa33424d4233d724afed2e5293558e9418a37ad447a4fa4da6
zc0b66948850eccae347b054059ec4236826b1230760b296a19187e8168ca4f763adeef5a756a6f
zb7edf6abd700c8c4d56730710a9eee0f0579f76477640e50fc5953f8d8635d5f1386dd43651546
zb33a93c922390e7cebaa84ee7d86fabff152b36dd14c65d2dd22d37cf36c7fb2b15ec798256b65
z7fa5635c0c6c828e5102d505fc4ab6de32ec327996c3548c7638edaa453c668925a91a26bef67f
z61a4da3ae94f93921703c59fef0aa3607cc36a577b45f8e8c4a526636d1661d13239e7ba4ff24c
zaf50e8cc252663ca5cea5a3208eaa1c9bb895f75ea45930f9261159ee8c18b23daf743a8fdcf01
z1d1077bbdde2fb7fd36abd9e7e1710046ccb7a2132269c8fefa30b593e6c422ebd9a49498fa2f6
zc88fc085eb6fbfbf90b6354b81c7054d7c0ff93805bf43085fb113bd374de98155ed2a4cd72a7e
z6cec63040b9c23226f0800d948045e5f9d6189453701e1a28d157358208605d6727c3e964d1517
z7af3a9a245f0e225b9a1624c48278c22ec3311a7ff4e5a95f14e5a4e933fc94629ff66c80c3485
z4877dd445431ae5e9231c6e5e24fcf89c54f861a0471c5120d343820eacc24d5102c8375aabd9b
z3d782d62860f94dde1700a623bd74ba46266d5b458ac472b75c387c50b03e29c3824426a0605a9
z3ea8046234857744dd86d6113d0bb66c3c97f71b969d5b2f1d66a0dfa1ccfea26f07bb951552fc
z8ca8f6e6e9e66e93fe0abe3b64fd578aac2946c9bf8414dd2e97ae9713b0a70671878dad27db8f
z2d32668067c37db8b3705392994bb6b251315fb9dea3e66d45ae1b48eace4f6bfa886e52acb686
zf204355781954b82b60e554d83c687d553f5eda1681c05a3b94e7f5b98c52af2ef5c0d2c012fc6
zde49685dda30ff051c287d78db5f4aa3b8da67e2b2a27e30b1627f1d04693b958e81255c4ee2bd
z281fe5d5b401e50051b2e2ef9ce599cd70d279acd780a4f3c5cd6b0559879d478ba605513fd7c9
zb6835975dd26f996fb73fabd28e24a5943bca887e13a8e2479c80517a17ddc9cef9b6e8d692444
z17e6126a5862450071eb91776c1f765961b096998b62ce6f9ed4531d0c08351a53b94a5eb242de
z5e911a62d366ed472637226a142ac142ba36337f8e7dcf029e438ed6f81a8865d0f72bb58ef44e
z1b9835104ec5a8d9a308f26c2e52e65ebdc18aae3f6b2b553ed1f324a9bb8612542bcced451461
zad146717856be8f51c00279f1185cdf66e10de56dc0a9e2d0e49f202efc0c3d801cd14d8d96bf2
zffd7478f0b3f72d5d986d7e676654e5c2832d83dbb4ccde9e26d631bdac0b3082419289a13b766
z8a23d6357b939b75f6bbb34d8af2a526cb65b577339e9daec5d78dea4e65d68216491a8300f517
z509311fba5739e3c07620b943e1f7116548a0017a325108d006adf0576b080ba02743d0e375991
z9c345e37052ce008a5f69100a7dba26911eb5baa12ba9b483634cd4c526a32531a480e72b173e6
z2985c7b3b39ff417ff7f7ee8acf5c55286c60983f1142dc1826ee3ba3af3d1b6a0625045327dc6
z1b5e8a194000a124822ab81ac5b5a6bcbf18e5180c3e598893851f36fe3bc0c8e0aa10e49a7191
zece54193fdec4897cedd5bafc21168a57a633054a3bcb7a44188a2878f8026f6a0bf46efd60bfe
z5e7925e9cd99cc60b8335298da76f661d6963b9ce525272ace4f2e7281e7d54189f38f6ff0e7e0
zfc51fcc566c47409667abd1327199e6a7c7325c5b3728685aeab8c7d631c631443dc636a26a2b2
z76af13fe8cdd5150ca5c898cdfa158cecbb13036b03303c3ec3538ed6691af29e56da4e6c5393e
z18e1a3a64a68b5339a71d07526c0e77aaaf0c0ce8f4f5fa1f8bce7924d91c05337785dbb1e4e8e
z71484eeb9ff01f1bd7c81d5a4a2401fea25209224974c2cb762a4222b5777e978237b9364b8072
z4b5206f322c742ad2882768e189367e017b572d16ebb2ab8a8c6533fb89135a7db0758a65b8a49
z052cddd976be43fb90106ab8fdfb38d253b10417f799406954c34193bb9aff8d60d4b6e7af2d10
zccd7b55a05d0af0aaf146b77fe340c1f906a9520988b2ea95affe8019bd738d915575635f93ef1
z57ee7e1445ef60d42719ccf80df6512982036478fd55eff8e83a2d9954f283d58899bb5d778edb
z2f60afd135da20bf8cda7b619abaf31dd1a9985112e65b9b4f472ba43bec3cde8c9e15faedecfb
zbc9128b42088c833e99ba34efb00fe065f79dcca2033800e931970989ebadf829ac3253ca49bad
z24a6b3c5a84e174a0f49cd71e95b565e72db3d7715b5075401904383ffe7d701899858ca6b218f
zaaa65640809a3556069736fb339f8cf7d45a65c528eb6e6a5d4a50ebc082f487abfbc04418cd1a
zfa45e0a2e40ccdf53d01ce1e58e5288b78fac9129a5f9bb0e198e44c9f7d4c0859d7c78e9e2cbf
z282ffd56accd24f5298d6663d861b69aea0606e3dd5b14d93a6097b0c3933d97b29a2648edbe5a
z0c92be4344d5d8bae68f3a82c8d0061af65a9e09c59c23623187e64f8e3c8152e7a0fffe979045
zb163acbdc1074fbc2aa9975545ba1fe128b458402183c51c10e563be2060b66f8ee68068c31aeb
zc2bd3dff5e26c9dc0c24cdec1dd019d1960cc75594a192f157b71399489d3a434affb54f339b9d
zbdf72bab4b19ac938769ddc24cd81cda316da87a2d8fa22a07299bfada8f40efd30df8b3c045a5
z0ed8c70aa2e7285aa839f9a1f8d251418b3241765b4b3213b1c72f5d8d193a8e9825cc28a2ce75
zedd4b54320dbb35e217f8fbee32e85c30c24fad1ab621437768170c5a0a91aba4e72555cd65dbf
z95b49958e03a8679dcfa659fdeb3a216496ca7aaa1738ad31d87f397378323fd79efc4dfc05cf6
za45dda6affa6512c537d45bf5643a23d4fb2db82d2c612fe48bf77b9a3d487e864dbf842731f8f
zabc11c15ca9515858f3c9ce9f6ed325c200672726b36ca08d8b426b551a27bee1596ed0e7d0489
zb89b82a4bb79dcf6f3f4cf00f74bc46e1e04434b724f885936b8e6e549c7c7ae8ef2bcd43f5d6d
z614df645cbe3afe72af78a5f57e9c689854b30773dfe67e58aba6d813d0b2b3fa690612e8b548a
z88cb3fa1da42910dc2cd913fb64df7820ef7bb5369455a52516f5371d73bbf145b8f8684407e3f
z8030578daf53f4f056829336e1d508d5e17430c6b3bf5e63936416d25f742896ca68783d1d275c
z38ed7f9a5048702bc2accd37aad26fdf31573b350768187a36684168429c20311347111a29b13b
zaddb804eec3a1a783353e5f81a766499cb70bc3e087d947d36eeb1495eb901e4fc952869cc4631
zc62b9131892b4c7df39b26e92d04f5ad73372b3171d2d6d68d9dc9ad949ff4a702efe1870b3b98
z7b58560bcfc04537835a6fd3a06bf3a1f35d2b51754c7640a796911c00bdd28005861a94861e13
zfc739357aec35d9ab020cb2f51baa8e3b329aa2be6e4268e55a9a0cf144cc9446f8303c3a81938
z257c7fd34a669345ad708ffee1d31eb7660510c23b5295cd3a48ebf95aafba66121370c7ee9271
zc6e0c7e57a14ada9290a2e39df53fe7e80e97d3d45176a7b029df9ebef0f550bbb04d916b2c7f6
z0652425cfd437f1fcbf8ee17443c5144d7516652d8718e2615059b9c7d9f2bbbd37192fdf532f1
z39e55204568986688d7064ed28e1d36959da47cefd83f471d2c12028363aa2deeebbf56dbfbba8
ze3d34750e90fdcede9aa7acb5ae1297387f699746fcaac79c260edce92c000dbe732130bedf2b8
z40468bbbc4d765036ac5bb8b3237698b2f248aff285682fb9567aca7cd9328782031d0cdeef165
z8e06186b41a3a52397d337d9117d818d730bb0a4f3fe09ec3dfd7aa9fa039b42b4e12309ff065e
z2763f38cd5b54e44431251c1de02c33720c27ac8a18a4a92692665be9821075d35a8626f5a3b06
zbf9f819ea30625c976711efbc84b1ecdeead77b8b8140cb2c571816e2038534403baf00fb8603e
z060c8fa96e04a9ad6a958ee588bc6e3be7c78f65d748f706f77277599eba7008fc4c4fd82583fd
z0df8b039cd72a438407a381715772548dfc20da4ca1cb612809de8d26c0172ccc8fb52a9dd7d3f
zb25d8d0cdb8b314655e79ba784b7c41252473b861677d58fac4e687598770a8c3bcb74d9813101
zfbf327fb8194dfb4df2dc97cf0959cbcec1555f2b3f6f04c2a611e9101c998575a767950fb750f
z5b486776af9e61d3e07cf99cac6a1cf0ab6d16a40286f2ae5b37eeac2dbef80b784f01ce4be447
zaca5d35de5c0c2d2fe19c0edecbba62cafd2d5fb40cb5bb4bf356baac55df0a8d1b9fc9bd35ef4
z7553ed4b292637ca7a97157ea2cfa1fb4bfa55bb360081b566b604bc585cb8af44d49f06380827
z10e3dd0feeb90ea6aad22267500803d1c026ec425d24171c006ddf53a7f6a5c01ad26e342813d2
z2f972954e923b05ed3310ff318f3517900de965a1523a3b4f11bba3cdd27f1398e758894d71b33
zc44c753da63f4ee201820661a2c971812983f7bd72c00c9adfa428072bba22880b7c9139fc3259
z66d6ef8bb96ebc95587d8d04a8527bae03b952458935c2ad2ffe14543eb913f4d069aea88906a1
z4ba5e0e7d1667a619bbcaada7d62a90a74f760d4d0700bdec50b602347eec53b9e2ab149786165
z415a9e1a584f4a5839a0599bece6f7961603a42b50e01874e7fc19373a33d7446f94dc4994fa0d
z824d58ade465a226c8c45b5d23643928223846181a546eb619deefb91f42832385bd13b3d8fb94
ze59ceee1a1932a19a6ded9d6f4687bce14f2cfa236326338f370d02d8d9e5f9c81e7d393b2a35c
z1c09187c5b82f4d7d10fea4f3f8f57bc29c3142f18739cd30dfb714e31bbfa19e0ddeda7073513
zd3fdda20cb4e52533a2e2409fc97758e80c4e0d4cdaabfa6aefef8f9ad149ec87fbc45ee23bdfc
z97ed53da44c479647d2efef225050c8473b6b672b883bef82c82f25915b34b4c99ada7c87107ec
z4ab73a1ec1c96b8c3bf004bef3a3f150f8000fc6d7e48c252001de0c878c1f006ff248cb76865c
za8c29c29ced348e61f6f29052e64328f67f4c4e18bda85f88152be105adf11a4b75d6905ad3cd7
z36a58ada4a196d1b42207af3295e1404f52dd9dcb3d8922c8c1e7eca8c280d746c7ab0c4b13fcb
zc862288dac9edad8a6671e1c290af358a33b8847fdba99f2f69235a432146873fdc97f6b8ebcc8
za1c25df04e9b7a5d96e07ff66c380ca5c97e41a0b2d2c72d9d431fcedb2fbbf4da5b75e4fa94b4
z56127b68c61254e30c805d121d51d78d695d91734fe56d39c23e8dacd16224549ec5b990745513
z53596bf54fd07998508525e861d8e4cefaa0dfb2267041add6cbe995e5d032880b92578e1a42b5
z5ccacdeb7b83920eb23ebc5b070d5bd2bb115456b02efb5325dab65cd514c35508ae33ae7cbf98
z71a7adc8c3606719ead6792fde7e1315a185c5b73d09d4a6aae45158c166f9874cd20591888fc3
zd92c28c612d1252fad891cac009b25777f2691cf1b5b857d8a2fa5a0b82212bad61b7f64c9c212
zb141c8ffb3f803e1bd00ebb51e67a783323269740eef9b998d14cb3db85b1c34c6c11720f634cf
z626049b7fcf958524177e7ce0fd34a5b41fb056867b089aa95b2e8354cecdab45cc87c6524cf4f
z991403dc5068127010f57657b41d7eb81d0d9854fe4f522d781e40f9ab364c25b49a2ff50fed14
zc57ac54ec41120115a487eb0c8cf3d53e88e305f5e160500505fefbed799ff076e426377114839
z92924b63c4365de7ea0d110bf96bb173d995788d290375ddeadb87d369eb34bd35bffbcf0ef583
z7922ea378b96e36be003f41b60f24c99ed925befab57ac21c1b1eaa52f85486945b69ec731218d
z4dee0009b55990501fff146a5baad48427d0d2c55efe152ae3d980921b225597a09ad0c0b5c3e6
ze502cf268c9f62fa8f34012ce1537c66956546c7b5e6547f6cb241a80931a9445b9e3291ac6c7b
ze6736cae3d67f7045291d9216393ee474918195a94e5d484b121c3eedcc00dbe34bc936216a480
z23d0a7c3b7515ba4047ec3794140893151fb22a8a3cc8316bf49c5ef68aaf2464a4d3a95233395
z07f2763e346832510ac51156156774827237ccfcdf48d9e4f6294496e711f56e3fb78aa5997eb5
z2666738176e9030565e917e64d9ff35fefdcd052c2c193281ebbd9273ec112c2c18aed41d759fa
z2eef863a90bc154c3a2f23d2febbecf1cff627ace46fa97ccb422fdd449b80c309e7ed18706599
z81b69219d3d50cd169c148c11298a89a46bee2d08b4f4f8323db568349510c464788d37825ed5a
z6d75c62c043ccb939d717e31e467bdeb069687ff4320b27e5d40d9202e927efd1c8d8030d2ce07
z7fcafbb184e96888597895c423ec6e1c54fc5432faa0e8c6c147031753c1b769fa4e280b58ad4c
zc0930c4e3fdb348df9809abda3a04981091a74724a7c554c86dd1b672c74e1f7c6dca6f9b659f3
z3b67c8d9b8363f76d4b1dd9100aebce502a239293fa2ec8c0523ff2f9fe15c87ef1de8287c4ea7
z46cc5c4c6ff9b169055a21906401e888f5931ab73a48fa40a14131f9d4ca7e52a08550f06c1125
zd6ae16938bc9bcaf078601acb42c3dca70335acdbb5da717f774e3502458bee9111188793ab9d2
zc170b7066345c940473f2c5e6db9f80d179c6578f3f2c8737d77fd348815effea39349d1ac9f5d
zf9173a3274dc0fedb89c8881492f65ce6c87e5f2fcb31b164bede359afeb636f8917071e8875cf
z78c910447fc87aa197a81250837e359282395410f137b7833ca1e3a04fce4560948019f2185fbc
z84ac3c6bdd3f227ce639d24d35f974c877f49a352b6d09f36dc500d65f8a124bd21ec4a9ea7c04
zbf87f5db1eb9bec64a17f17858aca9585edd2af633eebcd4631e00d901818c9e6af3753424f16e
zaaebb4269dc9e852fb6561ee7946d89f128d703088f32b0367d24e08a83ae2cc9a2b995657273d
z28939f3e0dbb798eaa8c9e20c5b248319ab13c77597a1ccd1bff894669c01ef22d0b0a380d6a3e
z75f8867fff9e3e2884aee58578169f527d5555319b752462bcc651c5b38cac9c67c3667997a7bd
z7709e57c39dffb442f38e6262bc5d426704d15a0b83f043cd62cdee598fb5b69c7e255debbe568
zfd0393d466960b7813db54077c4da545958e7c2243767cf4c015639a53245ed9cfd21ff35b8e6d
z574505c4981a5a7aa9b12cdc4eedb579a9f8a28fa541dc034033e4aab14060b04e6c01e979a20b
za6591aefcb0c2f49c4de727d56e35843b68035af505c51a1c8bdee0660dec0d76d32223625fea4
za266f83785a54424929d42e9da8c3c48ba47e697e0a746aed6bc06f2f486cb3baee9d680caa749
z2c7ce210f12fe672e7a208c38bc10418bdb9584f696843c60df2d99b5877903e293597e344cd18
zabb0f7b9b95eb22466612d1f98388d12d32bd576f03b439e9db1fd277c1648325065df44c0cb5d
z590cbe7ac3941cbdc68f44ac7a685bfd6796ddd18670f6fb1439a7ad6ba924a33730cd8381d9d3
z17fc6e9761dd7b8dc1dc7e6bde7d45d0e44e2704bd2a63991cf12997914ea38c37dcd80d2fefa7
z13b4e76c2e6eac7f9c107eaca0b307c101692a099ce9ff0f3931bbf06c5c90e7afafe1d998b40a
za60f3d57ab050c23ab5cbe55898c8ec55b60e4e337a04e5ab30787446819311c041215de7c4786
z2a71ef1ed333d082e376f5026be84d682e98bdac74cdb93b39369d06796d094aa8aca6c2f40ae7
z1092d4f1c7c6b649e2986ff9cea03b797e2f0d9c5b7caf9cb89c0c51103bfc0b5b22e5d472e347
z7bd7fd38b411945d839431b77633759f95a4023bb469427f7ad82869d1452bc29ac1a6273f69c7
z57cb3e3549be920b973e807262259245890024561c20f0bcf2992e79ed6818cb6625ca494bf54b
z8be134743d325e6d8ab81ec950fe9a986a2ea20d8511d782132873f6d7daf39d9380767c17d715
zc5091bffc61f852a15cd032d279be97a9b3f032319ea7eb12dfd3f78d154c0dcb8bd8b8959a4a9
z25800896d30bc9ad84aa346b61f1b8a2a66fd73bf66eb978b7153a6a9a7c8bcba0083ddc3bf869
z799d9567622417268505c19d700fdaad93e606c317db3f57c8414addd219082341383d2ceb6509
zc6153b82bb35b3a9664b566b4b7ef34e0394d97afeac342cd343f926d1dae5825fca7624364f1d
zf06fe9d81f4f88b5b4cf6f7bdb901e12cf1f87e151516631c623d24f1488b5d796419ed851bf18
zd359bd9c1a7afd8d1c87dac40081fa772f60106bdc37ae0fd70bb8b9420d70713e1f898fd67c7e
z0f6f0083260d4aaa301cc9451848a9787ce3c48a78c9f0b8e3bd6619b3359b4c1353dbabfc7e68
z8499e838c871ca40a8f998714a495e6f47bc1faff6a4ae22b58e774b496a8117d7a138aec92caa
z56b69c97d98315c72305def9c02dd58aa6f460040ed5fe0ca9edd1b6fec5b0f055f4d7cb4e5c4b
z79107a19744ae4132597d6d70f64e000641043da0ad0a86ac681897166234ab32d3752d4e98f3e
z7178c4a69fd6ee1d6f68e25c6a0134ff318ab32d9bcbc359ee4a687cf1a52a137a2678142ebdb2
zb3f58644cbd0d2e4873cf6abb7ea4b1c29797ef30916c120149f389a8f460ca26d00fa44036525
zc96bf4b0020bcda3c120abf434e6d58fd7cdd083abbec3ac15e1987a93099d9f08b1ccb02ef427
z2386543887a02050dadf7292161a7df533e1beec748402a0b412f8ff36b9f3d247258dbabaf402
z042aaed65ca0bbd9b20ead21e9ef507c285098589f2547217836e0677c28ef305f000bcdd419be
zea429155d413b21664b796e449c5beb98d38a375eeb758e826386b0ddc1c2e01820b977f5fbbc3
z71c05a49f67945432f01da0c5e489689aaffb9701313141e3f0ea1cfd494118a95c267a90e1d59
z265348ad3c865642d4c3c3bb78825148bc1bd5798b04428d625438ba407a6dacb42b0504dea183
z7fd1b1407b56ef84b48b9b4269578e2b60d2437af5400244595be5faf44515586a8891517253a0
z51887b4d2a7381362bf6852d77aed7b9be2cb69a9508eb110b5858329ed8b6afc3f8ae9e5c7ffa
z9b6e12d56653fe0a651cc40fbf72371e78847e7a4511275bb76509f527a67b4d2a37bdf2483d07
z537aaee187f7f8c526f8c78045070e228c09cd7f9894896379ceba6fbb8f3a9ab678e600b1aeba
z68308d1894c66ba16dac12fd74ad68427276ac2d0971a7fa7cc891c8fbd500c2ac08a25c858006
z4a0ee3e7ed5b71f7c369e7b97e4a657a77bae439108cce1426aa42be95fa25e383bcf2ac5f459c
zeb8ca956f89677b4b72a1fcce10c6f3e84272cd96a42297dee14b5d70ff6d9435f398fabe14bdb
z8ed99070441bdc843a7cc39943ca8dd6202f06b38ae2109166a454ad7789fbf251a1f2f9651fc4
zf45854e74a7d22f1ba7405c662a5f8df577b20debc4a6158a7519284ae4b0e2bc6c32963a788c5
z651ef12bf585d541bb86087710f09f62ac21aade561657953fe9b7964ebe584ccd61fc853ed15e
z76a1c57fef7358206f77baf2cfa351c623f715c8c02892438ec60b2d4f9f48ec8d418233f03d70
z4602f5abf7ef56d446d4f72db598038ad662821d69532d613e59ad0691052864afcfde1642f90e
z04fed22a084a99f7d1581e6948bb55dd66cdeef5409b80b54ff9a7460f04fd6e0b87014e1a6ae5
zc871b6c01356f2fd6bcb2550d3a11a7d6118452d2b241453787e991e96ee89199208a561528668
za36f19bc29dc6240b76039d3ad203884169e49aacfe3d833fab873181a0487749d1f86486001e1
zd2b296735cc24902613cc1b37704e79c9a399ab39f4b66f4140fb3e74b653258bb45e0f4e1ad26
z1e28ef8fb77b704ff8bcbc9e24ea0a84f4a93bbd11fd34fcf2b23d7f851b31312b7471eeda9219
z00ba7ecb8de27d8c87fab42ff8f889f5c1a3c723f2fa49f1ddb241c66112866ba5f87a809a1e3e
zdac864065b12fbe6583b46bf92bf53a8d7acb12698bed4e7b0c50f23afaa222044f92b4772da33
z6b63717eb07189b7325302591c3549697723171ab17571e4321d1d475ffa8ba96c1ed47445d913
z5d12a19c09e47ff1ba14763c223f52988f5b3c0845c3823c7810d7fa8eb1364df11a07add77ec2
z9d480775cd44b4e035628991d9e8fd7ac245abfd1ecbcfcff9a6fb02f22d39f9996aa5e388da9f
zbbd7b1492aa7e63ce1a8fd03a2082ba1a6d68553096d0b4acb1716cfc740b2c32fa548664605fb
z321e20d39d84f56898fe2ad5bcb7588488a6981dfe7330697cba616d9f0d06b034ec60ea54f82c
z6b46757b2d157b757a155b6d2d6b19db023fb872ac39b9437ba32eca3f6f1a9e018714fc76edc3
zb86b8d06166401b194c9e27ae430fde172f10c0fb55cff0260929cf289428c753240050212e991
z95d498bc8e39de1dfb8ac1c49fba0be21d2d5265675563161d23b652ea5f37aad12a83ebded4ce
z772d6b36b5d2e9fc269c0ee93b82c2b24130bb50e15fb4c62f780b5c82731f3c82801461867d98
z90f5093fb6a498f53c3dde6344eb4273a7d4194ea15c2d5773ce8f60d190ce2e1449f1f3fcc99e
zb2bf42affd3e5fcc2dfe18dd0831cfa019c255bb1900ae3c34dbeb687fde4a5144d9310c48a00d
zab18b0e87726e1f9d286cd13ea7344c89bc0a7c05a4aad18598744e0834f840043509a0a11a88f
za1894269f3112aa69bb0e4e3236a483a14a0b18ef3cdf6983833fcbfa2bb4f50758892329c52bb
z6cf7e90b4969e9fd5b4b2fd2ec69c433dc62d7634e5a4a0103b6f942c6f2cc7be4015fd881d6f1
zfcf3b9a0c204691c5b3ea1cc4f6e156af29a6c98e816e250d6bdf39aecab268a408ff41492132f
zcf05ce541a8006daed4a878091c272293535bb9f58dd826d13a4e6dbca1c55bb451f8f905a6902
zd62c347d717c79729a57756f6cb4fd085a5429b142435a75999962f1229d6923e4567859545a36
z5f4f7ded30c7ff3e5ac697880711a1e7fa427853d57ef0be8a8c52a072a44125c8918ebfc94034
z33accd35adee574e87645dd88ee6889145467221f878feb5549ad8124645c8570393c75310a156
z0b788245b91a89dd9cb04cc363bd7765a237446c224ab025112ebf4bdd82fe05880a79de3def2b
zdb24aeba95d5bb45456ec03bfc78b6e81583db4c4dee3afc24dbeaa88ac76fd26c1681f1b3a0c4
z373c7c41ef0751c74177f5abb11984a1f1974efe518785914a709bf4ada240117a5b957dc85d7d
z8a9628e842504a07144dd7d25d094f2b57aebb2687fbb4c4a9072ae753f7a27133fddb97dceafc
zbffad1efc83da8948d0f1e62077c9d2ac0b1b7b50bdb57fadd79912e241c3637c1ea53a3542c54
zf1f6762ed7222e824fe4b393a50af99148d4c608ad947f73188abad36a818a39ebfec65ac907ee
z12a6a36ddfef14c32128b4d47bbeeb6cd5926e7566a36f0e7b5007d9a09920403d5b4beb739b38
zf25b44ee594de5a53fead87435bb30d9e1bee9a32c906052b732dd94e618ecd6c27532680b0890
zeccef0f4fb7be9c0e46dd4363f663dbcc62bf186d079b4a0dd2e0c84af4da500d413b3d707467b
z98b34245d296cd61e52edba258e2e48be2c069143206997c7624f840a69551dc7ee28251009a32
z8b0faf17d103efffd2e6d49b7ce6b5fdccd1fc58ca3b7fcf4ad77102e891ccbd9dbff8cbe3d1fb
zd9120a3c5a9bf9a60e915b1218ddca685766e731165cac4a99b2e24913d899ffdd86ec5d788894
z2f63aa0b18531608b0bec5c8fb7e36e74a6bcb44b03f5119c909f79ab14e02489b2157dad8df23
zfffde7422f707ee9ecb5096c9bb99a4db199623fd68b922cd74eb55414df6cf0cf15d735793388
z266b50e7cede1a7c62bf7d39ace81061b6adf9c78e9cac3c867b40b39ffc342cc5b24e06de3530
z51a280082aef380e212bdc80f65e8b595e67b846f027f195883ec13b7a8c547fbae7b341ffc4e2
z9d05a622503afeb55b0266db4f25705b898bf1b65e6b09ce43a338c2e555fa4239815fe6073124
ze1969a98412ad1897ac032a7cc54c5eb203cfbf1b3514666cdd1601277e219ef83f9ee575eb506
z26efae1bc101fb8351b9c88ffbbf89d44c8e16d4066f7a4cc4e3d58966896d984deb1cd362bc62
z9fd8f02563244a26ad24649b06dcae5ee5d2bbb3618f81f01f02c652cd0e735b7378969dc9e7fb
z3e5149e703ce5a7f8c05736830c71fa0e025173ec3b987cb352cc588285387fbe54cd569aed807
z77230e65213dec939c7cf4ae1ea3e3e340b3b8118bd3ec3703fb6676113c459b373c07925871f3
zbcb5b70af9a22bb497b6e9db446cd444c6ac5fcb6ddccd7627f10870ba170b88867b84c807ad04
z33885817eeef8d40f27eeff78cfc2d51fbe885b65ed7fa575580fb0817b59b2b4ebcdb0073e309
zd0e25542bd8e1475684fc5574be24ad1a249e5e74dfd264ba747ef24d970e3fc6364b4a101e18b
z52198d7fb5f460cf64861afa087b6d85245c5e8ba9de89d9fb7d7476069016199e4fee0c210a4f
zc248d735befd6adcd50ba1ed04282aa02a3dc42110bf761f7ff226512ccb390bee9aec80bd0329
za485078a650223df3f3cca47b83cee51db84cd46159875d820f80ad8b090c8ff8d9080f130b4f8
zb786b201ae39e52edb952cb6e17a88c44f6a0ab937d88afd4613d8382e2b4de846cf9f8b4ac9ed
z6961957a1ccde4b2d33fbacd357f951ce0338074df50d85381cd57d5b3ca9046288496ef5d7326
z9e49d2b893b2a3a4492e59a487e8147f7ea389c33b2546049763eb8016647046530259003101c3
zd5972b708c38297ca496317d964ea27643b4e17287eb0be9f7872b68657883d7f201780dd235b8
z74a95ff1d4ee4f8518c8f50cb72996415e9c6bfff54278bcb12078687f801221b954340edcb51a
z6b466a93a45bf5c3ea70f0070c5ff62de0bde48a9503298642ccf49d9b756f657a7bdc59b89acb
zbfdeabb4686427de58991037cc335bca79576a59c98304d01365dd432eb3a5c8ead9b9feb0b6e6
z000da47bb6b2caaf90848f3c2b69e05ddd48f2841837e8a160c65f09f238f6e75adfa47dd0925e
z9b05bc1a89ce2a647e9a47d6a13364e7603d7abe3f8af9e94ac8bb76479b410b6e099ab7916031
zf95376d27514922b2c5000f5c47c280874a054efad50c4225b52e2a5f985fef38e8f2ab6bf7d22
zbc9f878398f39681442b08f122fff0fa5b678502b02443b6cb23fcd546bfffced7356d3692e2d0
z5709e65e4e5adc9f96106735144cbf3df97cfa04c69dede6f7d09afd21004ec6c6fabbe672e83e
z2add7099d4b80b5578cdce0e29ecc9e4e9bcecf35c5c6a9ea7b08eb0c92b73d5a329d62fd88e38
z041625248054cf38940012658be56ecd0010d7a7948e3fddacba3d5d306557d0c8d0bd91b9a33d
z4c8f512041b7f27e00b615e1e34396b10c8b8f6c0f07868bcc505b3681a7d6218ed548f8623eec
zdbd57c3ac71babb96ed92d9b1acbb7380c34215d47913dc1649113fcbeeb09328a1d00b0efda12
zc3cef1de9367d6e4eb123286d20d85e6c77ffffb89b3af2dac74ba6a2da104e663ff0d77a17cbd
z78933a0aae4b0b37fbf01781371aafbac8e40a6a98652621695c095308a40d48e0d72a9c770184
zbe6319ece37a8b93e97c19f8119c35ce0c1e600938b45f418dd2ad377545c9ce5bd8d00d8cb10d
zf72ac0d7f842624fa619e426906847c1e2f9570500405bb61942fb8dce83453b7f7f8a823c9630
z023596c53f2adcc5efb496132760e2585c30b2716cfe812930ccbcaf2e6da1490e456e131f30c4
zd205cae696e35ce4288204d7a151dbf89b6ddd637fdb4a6ddcf68f4fd8110d74b32abb7394fc27
zba63a3ff81b1508bd6e138bfc97d5f03642e20b48092b6df6db7a2383c7db49bf82954f2d620fa
z309cc4abeaa98fb6b46d92fb69cdaa9145a47cc9ae292e56354978659c9bac6c19c2af0c46265f
z859d9c6cfc260dfd4f71c5660bddde34b7691be2512e8ba4b7fc47c715883c6e7609500c5bfb8b
zb525651c9b8b0ec48bdbbe537acde7620d07eab47900bfb4f6d3fa034777572d0d4a311beb10af
zfcdc497bc054db6c15cbb76e29273fe8ec6a3c187dbb6ce4d89873efa2fa515970228de2bd2e93
z59c08e26191a47bd5b3590dedb6c0d9b88d03c5fdd30ecd0c5005ebfe865b942ec435d193d621f
zb8de71be11780fb47eb99ef9bc97064e1bd6aa7c8e445842cb46f0cf5a4e7071cd70ec0c0f3964
z978d20e10d9441b07352fdcd8c6c61216fb6123b7668554d19148c8df16ea350c2cb4f5adc3043
zbdfde5ee8f721f32114697a13317474ab9e653c3410e51d2450d0ccb725fc37275a19bfb246923
z9ae1466ad8689bf01202405a4e96e165a38a84e7d8c06d48ae7c7a81e89fe71601c1fa0b5a5158
z815a5248f69584157cc210051f07fff860e15ae0720d20c82af97757710931d8d648ea59286cab
za4fc2e83df11a6d64f6aa912d290f0aad6dd2476c5c8681653da78ca2c606a9b9b6238c6fec374
z7ec42086e9e4f2e4ef2c8e4ff10268febd7fc87d81201e4cc3cd39c597f078acd9c3b85e331d2c
zc414482e5a354bbbb571c3e171a9f5180030a3a20b9bc1535bc8e7d2c622e330e9a0f81042cdee
zb9a91c6223b02a7ff2879241da006ecba9c770834fb880a021a692c007850ff50df12ff7889a95
z40d3065dcaead5cf6ac05f23abf39659554feebeb8c99914815c6e3d2a1128d8d656d6e1ff5b3c
z237ad8eb164d87a753e078ac467d263790280497015f14263f097cea27ba0e622dac5ccd8446b0
zf59076c3ddd8934f1f4bdfccf6137d6c5fd2a13d8d8399f00252c117c67c26e889d1ffe53d3a0f
z65ae1e4edfc0fc797ff6e1afce46d1677632e2780eb0560d238c44076b90a31f6d9a398b13dcc2
z93f45484d7ebd2db6f57fcea60c976503e8a97023e5fa7df0950ad430864850792b47517598a8a
z0abaaf7a148ac79079125355bcb49743235f3449c984f951ba4cfc5c3aa368ed26ebde20c431eb
z9c6c7335775a7fc05747f76cb1265e34db1492b0590d10765765558ef8817a5dca1ebbd2cb8546
zd616d1f63c5e5a643b1f15c10e97d5b981d60b4a08941aa6c1c99148813eea8e2866c03c5ba2a6
zbf873d477cfdecb5668804784e2df64cbed802cee4d66c7e158559922c2f1e4aca5478f258e756
z5e968b1d631af68f6046eae1b54c31c916813e0182c6640dc49fc0e0536c3216892a8570c586b9
z62620bd537f73989c8064a6e889330c07e7f43ab28a86ad28789714bef07d1465691caa9933444
ze05f84f82cbac9940fe4fed6e3ee3f34ea0bec176732dd4a77df3832e87f7b40b8987ff30f3f7f
zaeda3e903afbb85a582075ba59773e017d0d50ae55fc5ab02fe26bb481b46e08315cef501e0699
z39fbc06694ce3a9494ec8a13953e31e6ada017fc7e1cf19f78d02a59273e58ca555d4c8e62ecfc
zd9fb8ef914e355119916ebb53336d2776b84b9b06b0964876b8c656f86de7ed285f64914c97ebe
z7c5a612e70da9af9af6f12bfe83e574565f96fa972a453173819177ad481bc6f6a211946db2c06
z1254b6b977da33b832d9933ec2a42c7bcd1ef91b5b89b8235b800476e8b0016ecc98bcb61f9f18
z982438ca34c3150c30df20eed03d026a09e156bf62fcc9eebc3cdb50db00f575f56e801f2fa085
z2d60eda58878e5bac7960511272769e56a99b1dd0682b3c0c6f4cd3cf54a8392a13a59d3718726
z6edd9ae657458345cf7cfbd0f4e3cc22609dfb60a9c92965601edf41fa2e890603107f5d377c26
z0aa175977082122bbeca18b7c66082ea0080c8c0eb16433276dc8c1be220a5ee3adebee641403b
z38d214a0ec53a3ec065eac9aece3aa2c74cb145e4931d6a870c105039097c7021051ef4c884f6b
z008f6a65ef283f940278ebd33ca6c889b1bf3e73f4e6bebeee154d3b04fa6418b6851dffc35227
zb67da07061665e2857099c17a292b8c22c42adcf06da420f99ed108fa9a98cbaf6c5d1a88ff59c
z4e588501782263bba1c57a73f49167c3b474514efecdc69a760da354da8f978e0901a87c39b911
z2758d6a9ac57fa4884114e5758e7a3a3b12bc373927f98098fe00b97029f188074f423bed80948
z8c409a7bd998db3f2eb915b826cb4b23cd080ad1e2fb5df8ac50a05d8113255ba466efb847690a
zee284e0cccbc7ffef9c736474bd91a4d01defe48b4a1452ca070517b3eb1427b7c88de3e01a28b
zfba58fedd3d90787c9ba4ad33b34ea5693af7426b1ac96de52088f8c5195d172231a4aa9d65913
zda30555853b8eb206084a8baef911dfd2e0cbaa09bb207b6e282505c629f07ead6c2a1de625754
z78daa6e2ec2f7024a1bae56637fa3523ba32717733777b0ac2036de15463f7023d41d2ea97f192
zec6cbb67aa267df1d80b905eca95787600b00a5436a358d970758d869db61973b489bc0f80616a
zb7e86b9ecf401fdccaa501e20be220e5c1466dcd3cfafdf5b92eb037a926007ea09f94f8c8f596
zf4443c4012a849f1d08b8cb3baae4f0b15292131d3db6c6fd3d713ff7dc1e750287caa731fd44b
z5bb9e999cd5232326673ed70547bcbcea10b0c82dc22c2d63995ee5d5d948a91d7e0138198b8e3
z4c00616fa908475798e2bef6940751223577ecc345ccce0c3303dfd2a52972cf5ac8e7b1d5ef5a
z24d6c3adbe373c75db1d8084241730f2a126af419d30935f9138566b3cb078e27452402243822b
z9bd041ee43aa2364497e3a2794eb43f41cf2cbb47686e5eafd804557329f689f8f08e61fd6b91c
z61bbcdae9b4021916e8cc384c3386c300ee059fe1adc8b4f6ee36b0a58ef646ca53c09e6f6dd97
z1a469b772dc62e2461ad42aac09b449b8f2f7da67e6087c928e5212533d0f91a32a14e447e6688
zc8af6e68c1ad6d83b4d089315f2e5b1e87069e6bea12c67f1e62f30029e287e25fb7fe3f786bf0
zdd9f5c4776a7caa89f7fc4feb84d3715be5239469f67a823de14c7d09edda76a8f3d597717020f
ze47ea0477ee36ba0cc945eb0edceceb81cafdab01ae1876bb5c21c69ba220db5ee383c5765ce68
z14ce83dd0078bf4b04ee0cae78b15df7f2ab32de71bbf08b7f1a8d8d7cbec5ae998c6d3d0eef2d
zd6c28cb97fbf5a0cbae52bc1fc945d549029bc617f576a2fc5cc89fc7b5b66cab4e29874d6aae4
z23086e1ae6ce1f1e5bd0fe10e077346122d0e2fda2612b3422760c6abce85199865126bab32f54
zc78599bbf34329b7cad69a708b61cc232b0d868bb8aee833bc0e4332e49f820916d55d69982e8d
zc4bf757a51b8d33bf9ddc1ff16bc6deff8e4048f8bbe776dfe5a67d149da2a590a0401894e96dd
z0765c845d923c3780e2a12f125ca2dec37d84856400adf85ac000f42b190a2020461bf23220080
z01f41049f44926e7ff88259a8e20ae498c5ef17d12e395743043840789dfb6663f064d451beed3
z5b7f3a8a69feb594c0d96019819ea02e6f5d0c8f353be52395e3611cdee22747ba1653a4b99ea6
ze585b56d84c20482bdb6b929ccc7b036e695e92e6196e4c2b0c91a1cf9081895f0225abd324739
zdd516888e6c6276025b983c59dc2a82a27a8407f4f9440af707570ef4122986fadb21563c44cac
ze65313a7d0187d2cde6bc49f4710f6f662e7f041ee779358aed46b4d701cccb72d1b98d82e0e5f
z960a0b6e4bc86a022b0bce03e006b28dc84e002e4ab80b78f2bfee3d2e857613e84c46037584f5
ze157eaaf683997f133c8c22b7e721e4a6812d05153d51d840f8d0d15b2ba48acfbc307c5b7625e
zc8e782b522bdb7b0fc6f56668eac952ff6974eea33037aa7f467ea09dd46850b07320cbd2d4bb5
z85e8e8fc3440fcd7fcef70df925e3529cba71083b1e9f2b218cbc332f612abc571b9b8ccdb1022
zd862a263c5ace98b2f6d0fbdf46ab31d1b6b04410fa0015178c50cb1cf1d16fcaec36f744d63b0
z50c68a0f3707613e1d8905bf51e1316532e9a344e88192cf6e47b6be5b8335c3581824aba9c438
z403cc88d24f94e7e47bbf1ce70d5180d128c6d7aecd04b208957ebe283c6045df344b1a3edbe76
za5e044917397903bb901e3a2ebf89ecd72f02622b2f4d401d0d7ce8c40487de31c3936875f6dc3
z32091cde8dac8de1df1466e511a6d50b4d848ce73cf13ef4d0492ec0b2d04781e41fdc0b0aab5c
z1cb1a6543af69d21f4ec320ea6814fd90a9f12ef4f7b0be060691e8e1df8a5f0d78ee95ec12a73
zbcd97160132cab4a3585bab48e89032f4b0877b5416d562624ba98da4be164e3c1559c533fd268
z86afb67d0745f8e9a54dd3776219e3d783d22c43bddd32da7aadf0ebbb77d590ae94f5fc34599e
z63a24b0587a1d3f16df979f3267e9061dd5f653cf05912d4d7f2bf1973ac6bc4cef40d0d965120
za8d38b583343cc0c055f26013d21af3cbc3bb76a34e642e8f42a2a91aaa5541450136f3146d88a
z545e1c961406d13d17a901ad603e769bbfb633858d280485eff504911710afeb708d903f701beb
z1ff24a46d6e06ecb1e6e93429f10631bf918e989d89a410cbcbeaaef94a10b30098a770d15270f
z821f949059f7cd291b5eaca5709acfdb71770c4ac835c6231259113fe42dce8a9950bfeb5c98ac
z245b5a2843b5ff2ca2305948162eab4c24c3ef6748a8b3945fb654450260f13476bb4f400b3479
z5e0bf468eac5bafd49b9b55752d22cdae31e3041cd47721fd46a340895eb1caa040464e2c2062b
zd37bc316cd7fa68baefaf5a597d77a98359a5b4cfb5e9b7bf236b9297552fefae5cc20ba86b2ac
z4f6dc573f607d41cb49c6e6efa4aa16eb72cae9a96798b628b25bc035f51021276f6c86306c6ea
z48b5254f9ab5aba8490b1657cd19835c42187768f42553ef2d79407691daf5fba1a86c482eab77
zf3326578f31a0beb431141271f590484933710552723dc8cf0dfa3f743969ed2312aa5015387f3
z17da702363ed3d6b3909b26050a37d716e2261e9e75496b4fb5c817e8bffadcf192adc961be076
z92f28a13caa12db27d067370794eb1d6dde78b4628bdb54d7c7cc262df7262c9dd1df5b90948af
zf46aec70b7fb8179ba6469d85872130eb25d99e7b5081bf0a00aa157a12fb76eb01101930bfebe
z79c5b64c15fa18030c41ec54cad8bb26ef1fe90a4bd58868fee771bdb288b53d5ff9074684c6ff
z44546adca6b7a3119fe767cea997295168eb26110fefe50a2fca454918dc30a1f6655e1624d1ba
zde7c9bb5f03034f1e25c2892796736efd311208fc8a04693ef99df1dc37611fdd0bb25143e61e0
z02ec0efdfc2a0ad09f9bca197e3d2cfc08ab5c4e796c1fc73b2e7985bc89625e709edc9d8d870a
zd9826aaa3c32f0de6eeb0599f6255f96716a43269fbb49e2c24a33bd5bcdc3dedba9cbd9ab703c
z156ed24fa4e593a775929850d84f49fc0a81caa3c6afdab5acd71e068c6ad99ac7171767313125
za1dc44d4a9c3aea2309f6def85463dba092c3556672d4781f7f54bd1b40a65dd5226296e8ca201
z16c99a41e0d8f207d823cbf92416129d33c12eaa7e4cc305652952b67f9a5db93cfb9121f9b6fa
zf0d294bcecece0e61439cca05148b23d8d9234feaf28feee9044ee0b4abef57ae6963d94b8904f
zcbd60c093e221ac6c33e68bca4f5c1e6f3419c4d00134e9bb21cc9377e5a1892cbf35f0a375008
z530e3c0b14f5e92311a0be9200abb2d036f78d5e310dbffe7a61344067aef75a6cc5189ca96e47
z2936493aea169f22e605350cd4f96971299f26e048df8165269146381d7b33057f90b787373e51
z54389a00533db6522de549c52f2ce51b2f496612cfe3fe883b5abeb7bc6d7d8764924c881748d8
zb812acabea47ee55038d57971d33fd27e65bb0ba2ac25cf6e2bebf40e1dfaf8e39c495eeaa4bdf
z37e03fe2d1c65b37e0a91997193d24af3dba4b308260c251e5797be9697292dabd697a84b12e55
zc65c3551d6aee8132d4a3d0f8a30ea5a8da73ec95d3d611eaace56ca05009a3e67a802af62cd99
zb81502bbb3080ce3d59a6aafd1a99613220914f5ee31db5266ebbf349609b7ebe6874036327618
z25b1b008c02a28ae8e8ab1da7dee66322ced182ea4edf5043d093039346ec142b0b7c2a4fd405f
z60588a1cb31f29e152a1af7f248138bbdaaee07286142c8c23ffed368186ecc7677ecca5962f2d
ze611a0d9d7a0f58a68e5b4f7ada4287b4e4e464fae427913f0da94894ab965c0ac4dc27f5b11f4
z039258c36d23ebcc50a51847a0d23a8a7a2058496f787f6a9e1241199ffc6d11bf303551518a75
z03af57b5539f26233a8bcdd31fb6a8ff20c2aa98eeb7ab8979b82df7e6b6036453f0032c8c0375
z7e2351d76496585de35661ac48e9a47505f20139bcc2fa9d29880e4acb986bd021d9ad2599a2b6
z32a1a2968a4f3bba352881d8c0da464780cd6f49b89f3873aa1aab25e51fb28acc27dd9942fc82
z487c2fec7a09012de0de317787cf2f91b082338535a6d7861501ad74e65cbe52a6bc05e8919d75
z502e7b51bbe4cd1bc5ce32ac55f153fa144ed3cb87892fe84c991bc8a023742c4c7d3f43fad44a
zfa66f63b586b6481a3070afbbdd3a93db1c8e677eea24e274675c9685cbdc4a4f5bdb79496320e
z8c9d7c1db8f62d599a23504f255924f55e5c66cbf1033d2b3ba83ad20a06db9dc2723922115be3
z4cc40a7cbcac62ecddd8dd00bcb500b1750ef9fe101073e7ce7f454f4ddd59c9c6a0c2174e880d
z256ed343ebf2bceeb016836c8d28e1dd66ee83090a81202f599be8cecac463ecc10bd3a1379de9
z037abf2c0cf2721593b6482587adef174a97a64a111dee41311c911b18b0662a8473001a024227
z371f34d25c832225af47ccdfdc2d738e9791e7cf2ce824f902af22b3d51a48928e84226b677b1a
zd383a4ddc8fa48aceea3477d8ec14aad7427a04f0f27965bb4a63cd0f87adfa1d73617465da780
z4ccd7ff96c7c7bd589ce671e76e4d09c3ed134d805977e693cbbc4e2470e14af531e39bd9a5a0a
zc4dc8a18ffa52f8c74b91c23e4b6df13f44b8886b50cf597cd35b30d468693a74d0822c185cddd
zc877a48acc51147c8837f97bcbf3af4952aa6ebcb0974f6c12b9286c36cfbb2f7d83ad5a7639cd
z869365336e2a2304346a0c127d403f5b8f031b1b7a8372d32e18678e8b17e22f986249af1a9293
z1544e60151648e763b60412d8e4fa40e38d33f85e852fd3b714d88aa729d2e66cf59ee1b890209
ze2b7891faa73d5eca0203b6b17a0170395087f4a3e9abee466b6d5da42dbb2464a2a76775769f9
zb978c5b8e1f9f0840aa1188a15208a4269c9250120acfa87621cfda64d2d31afce372758badbb7
z63ae3f2f35c3323e8c67d3db782d0692a54bd395213737c3a7a88ac134d2aed24f479181b8a9a3
z8813b96d1d5645f2d9ff47ea1bc962a9745abf3738cfab3272095642bd8ff3f8bcd9a56250db6e
zd464857b8e29109b777f05b7ea3dab064fefe11b45f20fd183e5edcfb3ead4bd23fe6aa092e5fa
z213952a024f89a4b4596b773e550d949b66c26df9cd57cd264f015d6dcfb580ac2bc64990107b9
z976a0367b2b0117dc5705bc62a6a0fa9609105d375cf5f4ee56a9f5a10fb4c98902ff05f87c643
z27d9232721fc4fd1dd01ed614fdff384a16d3dda7374643b3b425537f92a816cb761e9d77a3542
z68ccebe29a703af30b362832b8dbe541841c92dd37221cfe44d9ef15d5612eb75b7b19e9aa6eff
z2175055362a3b7bf67bb0c1a75ca27e0cf816d957b473dbd363d77fce88aa22a67cd273466abb6
z92daf248fde15da64314065fc919d96df44aa0f648b5b9b90766e4ac6776afc9ee7e84e9c77ad1
z395789a8f2bb0ce7039ec8b4482f51ec9c13de23f9fb3bf1376da3a7493f1c7e1b2e98dcf075ce
z4325577a6651da4cbf66e482cff5f775482067eae50980bb0947404fdf78d75519e0ac459d0288
za66cdff69fa79e8513674409881cf20383414eaca1f791e47521f295454e0710f6b36fdff85a85
z1b0e6dafd4c9a1b3ad5737a67c6f1465fc7bb99fa88ec304f3c7d5773dbda2105df90bf6bb24f3
z3133d60978cc643848b2bfb638b5847eb688eb10881ea2030a58d1d541fa2cb2a6ae99df299211
z5aa26e89f3d77af8b178b6fe1ce18628f79ecd1061c79149258a1c443105a17868d884642d014d
z5a0fd7f3d0fc24ddb9b5b17ec4680c16e0675a8c2ddb245d366d31d7495ff91a490e6f645307d6
z821236a6758c7f2c08c350ffe2d96b19596b4febbefca77cd02204c94af822508fe25598338f83
zcd6d8e12f2383b53abb0e7674bb9cb7cd3c015024f35c0c14d2f199adcd1ded38e0c3e3e100ec9
zdf924535f5b562a91be8b80ae17b6af41294b133ee7b3cfc4e9c71de6d6b3046da0d4c2ccbc809
z434932751834fe1897fe2db8feefc2c226bfd8bc104979a88dd9dfd3f7bb800a8a83ee6e338f6f
z751547a358e38734d88f82d114c454aeb0534437da535f7836cf9434741c3a86107d7c5a4bd081
z2ba811468894e8157a9fcb72e2f8c155a8d6e9d92173f1138adfdd2821ce8cc6e42a9f5f9d61c8
zd37393283679ec79df4755ed457058bdd14caa6f545b7be33b089e560e2da84b195f38aa28ac76
z173cb21a89c657920d6538772ec602f5bc06859f2bcee7073fe956cb7fe1789d2c0ee7175df93b
ze1d500364aa5d5b1bee5b2e02621f51545fd61780c3d6fe874bb1f27a50de9b70d0d28a541e795
z54193fbdc0ec5728cdb0f35fabb780edb84e9d12ade6276d497b1f489e94eb58f2274347d4e272
z545cc1e27abf5c7e03575e5a01b6526f353835033e0e704d740e70ab60876da68f0f9999ad4d33
zeed219e1c53e4a7a314cb20b5a86937a3f6d60a0e96b745adc26c789e69ce2ce0844d6ef00fd1e
zf0df9ef4e52e99daf0a72c5c028ecce8e496f9399ac05bab0259f053c14c4afff15da479981dc3
z4717780f14c575657cb6ff9e6c35b59f8552df53cbf83829bd6a6061b1af7457a0874a8a89937b
z96d3ba93aaff8c67bd08c5ddaad9e856d21c0f4e99c105b64f257f8cafdfa9bf0948015d5ed57c
z4910dab03f56d5369909a213b12470ba39279754e142932aa04161132eda05fb1ff744f45cd6d8
z37f75d6c1fb77e9a3e2a877a6f3364552006f4e3c20b705d13aedecd51af08f3f2b7949e02334b
z90467cc93deff2ee9f55be70a010f0fe1e4f0d9e3e788341bde6ab4e90038939d615df93a8e221
zfdb806179953f2607bca913c424e2da94da091d831a7e66c59ae8074d254a2893626ca18551bba
ze117f6d2a0c7c29dba7b151837d27e889a06b286b4e93c3030683998ba8204e6a19a4a6c2c943a
z3bf7db22db8c955f482e3da0afcbc2cd5abc181c0988e381646b0d45da6c8d4c4460fec07cc724
z07e0d58a68f8bd7e373d3607c8e4af32b82b64a018fa3dff51298407f828ee15af96da06e457cc
z9296a67eb546f0d6d1e719fb89de6708715ea5e4362b1da74a5c4dfd7976f420ae27288c5624bf
z0f0f6ffbae4721becd5393adb7b5a4cebda852c1568c967a868c8bedc4b7d00e71169903fa4f39
z09fe9d9bf7280911ea1f7dab9e5197e75cb112978466cc86e0f9f48446ccd25fdab57fd3ecfea2
z477881b69e2c97869e474974691f1b097c31e5f311f074ba8a35223c317a2850f7ce9803264564
z72b58e3c07c50f0404ceefc74fc560c7ce6ea98895004ffa119354c7bee9f06d2fe8c0138fe94b
z130a1d834bf3dc1424b3e771e9f75c831bd726a26c730129bfd8058baa87f92fe042ba274d368f
z85f305aaf339b3a36c0d5ca778b2832f59db3e55233f297cf0392fa694baf245c99dd795649a00
zabee2fffb245891d6fb962d496f980f54bd121cf0125a5f2d5bb2cd16b3eeb6c2b34624e7b0c0b
zb8004278a75b36818584dea3f39eb042048fcae2d49681514cc7fb47e27ebd9d14ff45b71b7fd0
z2ec5d9ab1c538ad308720fd17f3200b4caf8062c3309f62cd5a12d40cb6f178f226ab616af5e56
z5b3244d2461c5de40d844bb4887824b73ee21efd324bc3cd5c7292791ae960c92246d4762ed914
z9f98c547d8f1d7795253efaebfc378f7188074deb6f9636364f043b4d3598b3b7c98effc20a6f8
z0e75eac7c31bbf66bf671e4fd3e8a7125e22f2ed131297cd7afbba27ba3d3730308226b44f8ef9
z46f95bd6e3e43599b596ff41c4d98df0b4d7c52f26817692be4d53a347bfb4c0bae623264b77f3
zea8ced486df617ac7f5deba4d4bb10a2d5ffca6366080ee373dc6024d60c4e898ab0089fe8df96
z78588b352a67e3507541d160b553cb9fc517f6474018a25bf9a388d41dd118e83e29b0d670f7bb
zf7bb2494f255f8f89cf4928236f6314336741583397e1bef5444a21e96c85f0d3799f619d3e180
zfcdf355a2d3597a7e203839d54440938696dba13ad5cc09f75dacb9cc9faa6bcb2a37715e4f4ff
z866f71f0cd760020bf07100b02a93ba6894ff7a8f4ddffcad6714918353f1baad995adb9266059
zf2e7b9fb9e9cd53a5144159305f2c428acfa7bbde1cb678de5cbc66191e05c48c9f889cea1cf15
z9a451d90f0cac9af8c68ea97565a00f0137ccf2fdc485f0e15d6112d5733ebdb07ab91646ebe56
zea761f7b9bcefe9d620bb3dfac9eb6f4f9367066365703a100debe3e502b504622f2a89bdb3cf3
zcad20da807b3ed481f911797820e4bb40aabec2650f672948397f768d4f79feab44088ea5c68c6
z690cd73515ea4ed82f0f7ed650e61bbec2a5341b8a4367638e2cbcc3a71177f386159828875012
zf5d87580083d2912afeda5afdc9382cdb35de385398cb72a5d8d5a440f1e15a61abdb931eed369
z2823251dd7c13c8543b4ff1da3e62c1861311dd5feedc243432b8bed8600b30f18492087491b6c
zb54859922a4cd229427f1a4e1e0b62418e2dc5e2a637dfcdb1d3e812a0bad9a8d974e8a3d4a82e
z99d7f7346f00d8dbff06d53887b733ea28f601f197f3be9e6de982f7ba8b15ba0d943c490b012e
z74bfa0a29a7f47ce692cd70c15ab97d737652708459d96ec48367c1aeb22e387d9071d04030926
z81504377400da46a19c3f6972a505b486afd3b74db25af3ad22e18449bc9aa359ce853858ff54e
z79f0e779d327e968a483511badc509c0012670897e4e97540698f32cef2d3116a6c1d73bc08eeb
zafafa889a8e824fa6a231c6f84579a13af860d163e30bc99728ad9df0acc52fc7b63e9548263ac
zb564d210424c3ce18abaf5021699646bec9c65d72d4e0adba096dc88bd37c840727a9ddf8b0d04
z935a8f06a0ede53cbbdcd638dc0cccfcda617f54072d1fcce6b0bf017b30902396389c209f4679
z57ddff8aee5c8257e7fd0d80f72398bdaab8e8584c38033a4b7dd718b6b8b9ff7f7170865298c2
z5e89c05b28e860089e38c6dc85f3c696e03ce746418d7d3c74a260f13a1e3ea77774af7adf21c8
z5220989b1838d2360df8b17da3627a17d7f90f31f4c3d939b331bb6a104b7999df71621b5c50ad
zeb6741b706e39b54101d82395e8f56e623fa78809952d0518d4a0b644615649b49dd26df5c3735
zc9e5d3482ac3ec88d0648c515d3448f46e57cb11aba3debbb3799af52304840300d5dced514a34
zad3e20817d70a8f42f3995f5cc28423efdbe96f43be21a938d8b02734911be933182c9410414a0
z5362c693d7083c468e12e215fc09f23b450e0e79b1bc73c56e8104a136b08fb24d3d6ac6824bfc
za493f2da6d5d375aec94aafcea0c823d7e39a8520a16d8c374a3efa7fa5fe95f9c3420792b8b69
z8d9b71944e61221f40fe8038d1e3bfcd0e5279b82d3f28f4da2ccf2170cae1d1ff41fc6eec478b
ze5ca8bd4a736e1844e129dd14f6a523275fd32f41439e3cbad4ca135485005cd60a5bde793af27
ze54ce4a0b1a7c1965d349e794ca3c315bca4fba528d6bae243859673f4e3c0b8dc5d738541e0f1
z21ebccac16e46ae8ccb2f61a40a7d121bed36d9044169db88238adf07455b2ace50e0b420db283
z825759da4e6ccac6ce2e58db4c81c19ae3f0782a8d071bd503c5b64cce75bec499ecec76155ad7
z41c86d01b1e316b1cc056f5097cb7ae485de81cbb1d3f8be62f949925d08a11561c86c323ab65f
zf742bbded60858729088e0469a68cbe4f0f052f2b7ebd06fdf4d4120026e1c96a6f9fda5ac76b2
zdcefaf3dcfd72153cb9e6f6983539993b6bb0d4820c61600f8ba19b60f6d355980b67509a55729
z5201be79a45070e346d2dac9d6b01444eb2ead1c5e451da3a2cabae649ff6e2d2a414f34cc0b6f
z0df790f63d73adbde7e1a3d8db71d105fa3046ab4acbdd19bb6bcf2f7f46e4927817856ded2693
z57d69fb30aca753b3e8490e19db983e52c59733171794e891061bd76e434b22443c4cb666f4d8b
z29a649be1afeb22f16f2e672d35b64114815bd3594922144769c228a9c349a826e221f5c988ff1
z33dea6886392177cae7085d87c7afb77f8cddd4936b2e15724f0355196ff4e5441ce63f81dc287
zbcf4ae5ed30397d34f3ac7d3eb87a0a058f720ea2dbe69b68c983af4b0ab01b28907330350ef67
zaede4b6cc54f0246e5a1df1650c30223d9aa552876d3bb648ed1dd80297b9a73e115646415be60
z37189def579d85a0511f1f1f6fe11a3a81c2edbbadc418ecaa715db3df4e98856e919aff9a122c
za300379c0427aae31b495870a512027f40a2794eeb0f4b4044cf77c450a138d7c9f8f1f11361f1
zaaa9744c4e0012fda9beb95d83fbec4d4df1edebfe005ad385063ac6a20c34a874974dacd05b74
z9e1f730125ae98a7f0250d4affdbd39d4fb3dc17bab9e265110f17f59741222c649f4a8755a114
z9059d8972b40dbc13cd17e7ebcbf5c6d7a1dfce8b90c1393304e31cf07e37c2cd9416018a882e1
zf3f658d108dd8e7c8841f49f97e19d2116534967ca4204221a4ec46bb9eb80ad1923aa56176481
z23be93e37b91435a84d005db11483e52ba267ed57ee3271aa857c6af74f6004afc16ec4d31c26d
z181a74b32ec463accda81c3700102d523902ab2235154bf3729dd134611b69ec7849ab9a59eafd
za54fe603c6612990bcd37495b3b67272dceecaa5481e6b5a15a0e9fd67005054fd1480ee868013
zf20ebc37316a1501dca1e37f5b586b443edf7ad881adbcba8107420c5f3437fbc95c5827b63a56
z306408e976b3a2867f331edd6b9f9bd67d5e69d543a1755a0252ae915e5045fc913e6caa9571a4
zf4409ce77fd469c75f6e503969b8e933856b71ce9de1a1159510c086793abda51b9944d8e96d01
z77d44eff79846b0b5a9612e7addb4098786b5fde1aa71ed24a6bce18e9739d16f29b3f4e87b8bc
zc4f1fd599c18b4ab730dcd72c617dddc74a93be3bb4f7093dab74d9fbea907a5436c9b843813a5
z7aa84346e2360a3f9bdc5a7b0a12b2e0d787d654a4e42c5a65876fd0c3cb05e0aef506593bf4d6
z51eb3d442fcf1746b6a16b7b7031b58ab1a36bdf2e214fd25dbd99ee122bf60cd51f0f9d7a94eb
z115ad8e23ba96a1d93b50439dae820de75db87a88dfb190113dee5bc126b0f2d0c7eb934835df1
zbbdd03afcd42fb16c16658c71d82a2881ea0f357d736879cd9f9f90906592b82dc575a19177909
z94b64f876fd952711ca7cb964cc3aa9a395117715793b3ae41cb1081f532e99036dd0a2312fa06
z837cf8e160c39e9b9413fc8fcfbb120c25fa740f6d6effa72e8a1294b5ddc1c4731f5f17267cea
z0a04b44cd1d4d00c48926c709ae6f5e8c53f62650a514139d527469b61800d4a8be583715bf1ad
z7fbb737967e46f053d51c8717ef6ba9b3daee93f5dfff750b4ca85e7a64085e3c85b7595f800cc
z3368df43a0e714fac16e741de9f28b106dc66d12f37fdc7cf3f3d37ad48287b3dc4c8f6ea379cd
z560c9eebc08bda94e408a86da373023941edbfb37ce09acfcd182815e5b0739a7b2c0147834afb
z80b957584583f30db78d619d7f8c7013a32ac0fb5d5393c6209953310c4fd73b9a09c5b6490229
ze9136099ee97179c3fd2cf32a535c18a9450e226b7498e10e4e7ba89d2e709af33bfc47df759c4
z10b78e8c41c9aeb6589204379a22d45c4e29f64f7705ce3e4f5635c6f3d4a411fe1eacb31a66bc
za049d0c2badcd60ab458ba24530ca53a15674a5e39bb788d54bdfdc2828a4a5f4972afc5c3da17
zde90ce09561c090a8f4a4046df19a9a018c5381dbbb533e085e818d3f6777e5e2f0eaef6857634
z78b1e557a530eb1a3f3bbbba0c5192aa0b2a339deff3665058ac86b6f70fa55c308601dfb1d7aa
z6555218f4a35a423ea26d89392df7d6442839c70a084a728b1007ca8a34aa5275b0065ead0da96
z4d0ee81ec76d5bfe13b3b36c2ba5bacdc9a336ba5a2916c915a41b8fa8c04d4ca65a31e902a6ca
z94ba838e14abaedbff776dd17a8e3105af777fb1841ec23b1dde5c2a0e0152a25cb69ee0c73321
zff56e919f9101dca5d429f3fcee78313bfe9d0fc2c9013e8c406bd4f5be4150caed80847cf924f
zedb509e8fbe63f6eee4f3c5496a98020699e984c65d8968d5efd7bdc012978da46629d5e5c49cf
z2cee81b556a02cbb3d478ef69328df07591deec3c256c03e28114a5e1ee5b5581167b7e582562b
z84304c1cc7f4c3f7d4651e645d12f282ebe49e8a590640f0d30551c7926c3880ae55457403e48c
zbb02e425cefaaa035ab07c834d34d4b493f790d09599f8b58597f6a6cbcab0a27e3acb9719fcad
z5c89f08e2c4fd536926a8c8695bc0048daf4d17d7b3f6b687a3af53ebf3a2c230e93e55e95116c
zf81d20c01982f148c9ac56ef0ca620d7c6a0732fd65073c9a1214501ec655cff3dd7b9a6ede8c0
zd72d359bca0f3c3f4302ff245c0fd1784842c7d5f1968650b36a5a67c598b98e05ea7441bca4fe
z182e0c88e79fd1247c1dc07c136f15780b1fd30868dfc3b23118aa3eb524b419c53b788f96cdb2
z8be671fffcece1f2f04af532e0dac910112c3bc124cf85081921ce8671ae086a7f8515f9a1ce8b
zffeb72d40ee83dba6b7351ba42321fea1c028bfe4d32f1729b6f3749563a14a9dad3923d843de0
z669ee62f6b7d36b37536c07f9b4e870b900859be272cef37150baed6ccc4878bd5ebf26d4cd2af
z4ac40d5975fce0e6e27b25244647081578069e5d78740374eb97a61282809176d390d93eb8f5ee
zb1e83d25a3d277da579d8e202e2d8bd1ed9a0b36eff5f4c3fdfac275461bfefbfe1d0c3330bcc8
z8fd267574338d67fefb5ad3e2ccc7d98f9e0c806d0baf6ca787594360339b5f7136e9bd210d3f9
z77d8495bdbe6cdee177bea9bee3a0fbe6cc14736dab67dbd84d28dc824d7624d2a112eeb36ce22
zb1697616a353c9d4a8256c33fd657101d91b40a99834fe6189baa2fa8942394612e37b9d2299b9
z0ae91a8720e41cb4f5bb67b1d4ec3263fba2e29b7171f0e6206e77f2fa78b3c912a36f07ca2478
z0a37c6ac09a4a7833dbddce91939905d099b3d3ed38ec043dc7068e627397a773d772768940ea1
za2fe3b22638fdd5ef9a0b4a8922d51414638d739656c841cc0b8c6190c0a9b309d1634e53131a7
zdddb1645f3778dbb093ac802777939e197cdd8534e34bc29051a0ba3c28353f44b55b3c69d2ab3
z8c7a4d9e10fab9477b274da4f012d01579f940060a7e768244709dcf8f60327ff678468750e9f3
zb951d3c867752774e94d7ec8e3448d59922b7ef29985c686c524d413f718ff29de5e7f3033dbc1
z27e363df87238a0891d7c5d71fdd4b7b033574c68a4516771079f5412ce2f610eb38780f289a7b
z8dd6c82c6b465371c07a180e6dc2876fb4a3e52beaa6a5d3139240d744068e675cdbe3f03a1cad
z79d71aa158051a4d1560aa25a96d7d181c4290e8b49e6ddaf6de760d0e77a6e30b224108f80c69
z556a3978ceecbbfb2ec5e288ca7aeaf71299ff920120366153cea2c115f4fb9897b031473f32fd
z2228a1bbc287d6062c810d464f04ba7840ab138b65d0373eebd1d3dcc7198b303d14dfc85b06c7
z16e9605b8ca783af5793ffcdb5b49c6c9094aa25cb4e27970f94dd0401141e167e7c6126cb15c9
z4968dedfd0d36a1213481d420ed0e39f44afe5f5ed8bcd47d12e895fc64247177f5950c077d5fb
z2bc39620c62482f0fd0bd9c0242202657821c94ebe3c5502c8d65f91c38c752151c942281cd265
z25d395bb37b7373435e612c9dd7afae2d14a3e78b6c630a95941390a5422c9de35b5662accc9d6
zf25204d7843cb3a7e38164fd21557ac33b65d8a289f683afe978860e209c6ea0fed1d084d10b41
z5a1c9a4db74f6d49167fb01bd956348918158bf24ce65f5c6161f10520e70965f7fa0e3b7ecb54
z3abad8aea120394849adb64fd13263294f4e735e52faed18da04e1acd885ca06be142f67a182be
zcb0c163211ff71ad87b58043115339a89a6dfe72d0d3ca340216f841b414703dc7a0e4e3c0a68c
zda7cb9795ddf38633804d3ad5c19fa1324a73e8b6caca7064fbf506dd525b87575c36727181640
z2647d1bd8d8785de15d90290794bc05a0af3fea30f391cf4cdac9df209c48bf57d28e865b7e2d1
z107098c28f1a6b63b2fef8514372a3b345a48ce10a18296ae8406a252f5cd7f6b2ccc4f1acf946
zb8b609617bfbcb0cd50c1a3b34991faba5c19bd2d3df5d9d8f4e052a169a41e17a41c131f6e347
zff16387111a01acc7e520ad8cba8d0176107d7b3686273eca5259e97c861cb8f43f5c81df65287
z38e18f250133fd4aa3a01b683a51b1e75c9d5291358e2239fe4473af26d8c3577b8e3562520a99
z964ed3e734ea0b8de00152ebf3d610ec70d9e91a14863b853e8af29fc0fea46fdb17637534baaf
zbaa4f97fabd0b22c90bae47a621d79873c07b2151bd13b365f87f25edca3ddfac4758288198e47
zd391e90f977a8e35c7d278b1fa4c15c0c0cfb5735622c21b724a29f2cf4b921e26c6a0810b4502
z7eb1f994d7fff9fd42f74f79f6bd418f10aaba06d0527033d69acf9de0cc1a5996f9e53169f474
z50324fa26b0d0efd1ced7a75a8bafe31ac42b17fcac51c4e198a1abbd3cb85d113517629749fd5
z3e523c5b36c8d7a77021f9f6e7030ea85fcdf2f2a925b3618b1a9f6266ba2aae7850bf5dd65cf4
z7d857bd8b18c482650c41b03d473325c208f791e4b958f544149970afe6444739c0541f37537e3
zfbf850b187c07a4dd473784ffa478902bd559f68f38f52880a4f857e3868fdb672aa8cf089c011
zf42bee58541e041192d8dd2da8f112eabd2c2739e09af8abd38ca6a3c4918894ac1d6d8f98f45a
zf29e3a1b655ad2861d0ba02207d537b2374e7e0694d9fb4b979089986ad70b84d1b5cc34632178
z84ea609675b1ed875f3414f896fa23e5d147405dcbb4c8e0eff790361cc2179a231fd4817ae316
zba9fcb0491d8dc212911b23e2802c5a80d0af00049a30d96a2128b927dfad743b8599a622efb13
z07fce7a7385614d2a65510e07c48660df05859d94bfbc86889ffcac78b984a50d5b53a247ac5d8
z1292a252ff13a3a06f6c3fcd9befa3dd406927faefb6349a14f78a5c6b8b8654d737223a4ce29d
z4c0f60efccef80e314f2f3c77b3e527efac947cf258a76bc6533ffaba9e03ec6814fbfcc6be0d9
zf32dcab8159d9972a90158b9b719427c8592db006aa7d8ebb381ca2948009604d7ebb226de970c
z9dca481838fb85c8b88a2eca2731d00958add4d72566479389fd289a4f9821a434e9105d3af384
z93a15dd6ffe93e78984b6eddd980eb0de04a9d57dce03d47c215544d81c39a0e308e67bb03e42c
zaad8e25c477f0227d1b2cc46598531cc01467649ae08d4de1a450c23777e0dbc71597f405c60f0
zc2a47ecbdcdcd891fd8c3acfa19c0efe0d681d897d0a1e8452fe341bb6d0787453161cb04ba804
z0b5703e854bcad709f7a758ffc50f38e3b1aa33545fdefacd4e51efc817b28437d3a8535cece2d
z9d555326aae3d9b025605ddcbf09089f03385d21be44ce2310e361b57dbcce40a438b8c16eab1a
z206f6df201369c04e06cbaf56c8de608bcda825822d5aeac129f361fde898bc341306f1be102f1
z6bfb8518866858fd029e9c54ac58aae1e631aa12760f14bad765ac7484c41a7ac1b06252eeb0fc
z629a47d5f28489007695003814fc09d0c5eb32d82b3f776a3cd7b0010afd7b8a3481a17232a343
z96ecc02e1d000d8d267214aa91074915f47190333cdb980f517d33f72a5df8e9826c46985f4940
z25712a1919a3211529a4b0dc89b7e2db279dc33853b8ee3d29397ccb8b4df0cf3da689f554ded6
ze2e272f0ce37806e18e06720a4e4e57fff9dac21962c572b2727a4c2db60ed4219228ae7e8e0c2
zdb80a5ed3ce7f9bbb99317dbff867db9dfa6857d3ad32745b494de2713a1730f8b7e115bc57ba3
z19838f58f4e79cbe2b089e6c73859d365d41c2791fb9bd1f24cb70a4041ee6074d506da28b986a
zfdfd6fcffd5bb848cf9fb12a49c10eef38e1c9f592fa06a9196945b364d7446fdc81e5dea465cb
zfa7e920a23c19e2de25637138fc69d69b302a4fb5435bd97d6c8b0c20b32e97e31ca157a92f1a8
z401fa69a6689004d8d85a64a80a91b9720999eca9083505bb89bd48eb846f6c5ddc09badfb482f
z4097d86ddfe68b1daa1109411a07dc39b2b9e6d5ad6db32d0796627093953af5c69a978723aab3
z7329724861e47697decf922eb88e4092563e70681623fed1e9a30fe748623bc08291f3181ad2b6
z965bc848fa43a16cffbc59812f5fbf662097924bf9b47fc2f689f9894a07ff98d788a59414d389
z0d4856a759d69bc6a20d5c2f65fb03d68313d7cadec5afc780abb385471c672f41a2d15397ce8c
z410ff2603b3ea019d8a02e950f8ddd540f7fc95ea728043ba2c7ffaa42bd9da3c2af26b2cad5b7
z3211ea07c0ca8299da810a8faaefeca26000d9bb0630cc0d8df9cb69331f88073aeba11224ee4e
z3c8fc10dc0535c37860ba175520eccbdbce07e637c136bf640aeabcec9903093714085d4cf9f86
z46223f5eafd317f1831980f4f05ce05824d955c0c8a44a788eaa76a8413c36a17f85dc0c7e2faf
zeda2030217dc83699698fd531e01b0823475908c0dab2c9c953a028838c9326b0139281a567cea
zf27b45ea4937beb5c2e14214b40aedd844d583cf87ac39c80fcbf40f0248f88aa49d25d586d01d
zd2c0005e8622af0a2fb8f03d63ae663d2b20a48be517b61c646294b86fa8fbbec3bb0a7eacf7c9
z4ad50d46c71ef98ef0d55756cd7ff227144604e64ba707373ef18cb8ef2846f1fab09e4f815739
zfc1cd065ec7bea0beae200f970dcb9ad35fa86745c1b284b581b646cd742eb968fc5f61d6e9371
z9fdf5de459afa1ae4da7595715c457d6f0d7b67b20aa3953942bfb1598c5250d5233c44f3f311a
z870517b180ecbfd9697d59d2ee9d59de3d0a54afbe0df875674d66978d7029ac8cbacbc64ab4b9
zfb5e4f9976beebefcb372ca4727ad3c35d413bedfdb8ee8f88538eb2907a0ba83f7bf8517014ad
z7a74b2de2b7878e54eaadab6e041c59a2b52b571a69047149ca649a133e2f1a03bf73baab46aea
z4a303844759922163fd8d1af8b6487ceb855bb048bb849f0b1cca3cd39d8b596d5f0e1070e2c1f
zffd1b6e72134c975dce4a3b6d43793bf6f251d4bb8a1220a2873ed0d75038b57932c89e8d03a31
z78d86b2ed3a1b9d9c59e9e252f8b588e7a77922b24428fcf3a74539092d31cefc85ed60e20a80b
z5f81a4533967868b3f438a033ea6447c1ea68c0c4bdc4a5027dc6389f13e7218d966f5e5594bb1
z210fa5602a46ef4b06dbcf2838492a7ea92929531fcb9d43ebcdbaba4fb346cd399c184255373a
z70e1c07d4caa09de5faea2225f4ab91fee822beaa8426e4c8ab341ae608350a9b56703691354af
z2bf1013ae18a4dfc51dbcf39fba5dee63ffbf5f73369671c6127e9e7b857cdd7940b53d091aad1
zd5d2a8f2752bc1631636a5bc210a878413561130409a17ca13e6b91d55d99dea22bbb782293a4e
zc1087c36ef1c73807f33eb59bb6072358c39d8b76a984b74e7a25cf8219bf94e813eafaab66012
z4155d792e4d34ed2a111349af56f04167fc1488308908b9c4e311298b60b7c302795f023169f07
z1923c9c5b3b7546508bb9e87d337cf4bdb486eeb67c1ca539382f2cab12fbfacc78712fa6d6508
z3e4a9d4d66876979d1495c1b0875c2f9053f946f2ca1280fffcc5bd3576357bb4c540e6216c388
zfaeaa4682b176fbcb1d01ce06412b564513ddd6dd4839fbcaca9a204fee6670510e1ed53a5c939
z519f1d8a383eb192eb7b98e94e995452aa886077cec3a5cb79632bcf08b850e65c513c448f2e0c
z98923b4828ccb11b6d35f1fa3a0b32c94294622a36ecb96c2f04590fe6d6eefcadafd0e2aaf0cb
z151f80f5d271ae12acad1072c6f4df7d89748b6662372519d9e68a329deb411583b71bda162e87
zd6dbd1e2b557be0483c38540500875b25abbf67484d9ef3f8758174ee2185e26ae5a6bf0c681d8
zba1d717792ef89624254e2abee080d84043043c87018df1a2c9fb9c5bcc72554c7b78facb3e118
z597ed39e3643b12b625ae225700b19c61aaed465b88ccae2412a09fa561d41a4bbdf8478d3339b
zeceb2b54f91e9c218e15469d55e78731df3ac8907fde26b68b2071f41fa2678b89919e278a007d
zd0d8c544c8d5cfa7485458f24250f19b26b5825dfeaf990842c737ea5c2d61d0ad92b8cc473f9e
z51a9d2026246ccf57f129769ebd5b0f1a842626f07ab4c4f168483dff94f819f115e3a78a42073
z0b5ba9eeecaca3e994b74bf7eb1a6c3d8f20bd0ffc41c714b99e4a88458fd4cac357d016304951
z0446ae859b0333e83711a9b4699ab5893f3a830ee308c3e37e74f083f86fe440411edf119ace8e
z91215669e3370fcbba7c1fa9032fe799d919d5339565eda6aff25cd829df8d34b9c1148b184c7f
za0218f50557af2d3bcc24bcd2f9c0c5378408b4fedf6300f854a30f93b11fb549aa8c1c71b6db0
z2f3f418211757c76bab4f66f0ac3396c0235846f1be308fdcac42a25c8280cef1a15d4b1396fc2
z0930714c7a2516a70558c8fb301f873998ecfee928fbd806a838ca3cc3c5df6a1d1c7af26c033b
zbaf5c693d780eba3b65ce381527c25d7d4d10c067f9ce6ad344fd9cd96ca764717fcd41c2e4de9
zce2b547c10b246455fbb36c2cfec93a19e1d06a9d143490ea384e42bd160de4d7d007a0f6e8179
za704ce705a0ed953634ad8a4a4834344590e3c94e107c78dc020d3459c01e185952dde38c5a84f
z7703755df9ff463a8c04e4b219152c60aefcf767a32e8d31f2af9e73fdbf57eb8b1c99d8581183
z244c0c99dd3e51ce5f020d9b4ab675a4cfb76955d149278fcc35776f6f8f33a65585de27f74f9e
z402b2dcde9ec10071c067074b1825ff14909756551d6a23b0a18ef34cfde98e2cfb7737afd1e21
z086ab67f1e9f640a7c2c24095eaeeee01b03f65226b4635f191f76f1f7633ae27c118f9cd133b9
za3dc25050639c8ccaf0f02af6ffbc9e30abad9b7e890f19ea92f444fd9746377d15c7ae173e312
z42c11edb7715bea326f1c635d60b004d1ac245b729bee33290e22781db02704cbf532aaf0c7df8
zdf5df0b25f2a50181c496ac3b8feb316ebdc384584e3f02935610378d23f5c853dbaffde7bb137
zf0e15364231bbc75dae4bf1051a9d88967a38f391f2ceab9efa199e2746482816b8404de581e42
z97419da8f216a761d3756e738fafc8f81201dcd15118075b3d07bde27480a1633f56bdf023522d
z1003cf12f1dabd7950543311f3d7f695d513ee365312ccda65884ea285f5c327d4ad7bedf37243
z1c94fb7d89ef3e00a63b1e2c4ca69da37546c66f6ddc3630e570f7d917cfc6fec84fd9a8101bfd
z94ded2d44d8a2d9a39609b99f24f17efe95ebc486c0dacf6a9b8f7fc09c0ed252dd833106dbc1a
z78769bd93982d8ed1cf26e5e502d034d5cc19cc71603a6b6bc09781588ed9b784265c4962b506d
za1c01a77926e319dee107a69b2e7c7a6498714c03f145775cd7bca67745ab2f643d0f04ca7a547
za25cd4ea108cea27f3ff8ec95d795f8b9737793d34a52dfcb24fed6c310f2bafe13d303e47eaec
z60eb04ec9970ebd83efcd91803ab5c9f1fd6a1f68b6d432c9c82619abb6543592cd65b67ba3683
zd47149cf713245c4f0363435b41ad83619eceb049dd730a829fbd47fe743ea5089611324e60894
z527c1c2dc31b57ad885ae4d921233d4bc9b42075c3e8173e3d6169801f5f69d1eb1cafdc213d7f
zc57688941595d389fb09c379599711cfb0ff0d8d9cc8c83b5f862b0529ab3962501ab8baa4670a
z34a3f8dc19d9a6e86d163d507920acef33ab954206e78db7664f688b16ee8e65fa1566aae4f646
z5a9d545247b706b3e5e696d631b86a625f6befe777cc5c1344802f9e4aa05027e3e4c7a2c29e78
z9cc94fa20802add258ec0e565e23019f8725e35eada38b538388d7d37c81502c100405edf7db6a
za851b76ed1465328ea4bbda8111f3862c789bf18a815993b8135c8601c371e4f74e55c5d463b82
z5148f975758c7217f20fbd85124b9ff6441efbda41abb7382c7cd0441a49eda45002bc28f6b0d4
z31077959ef4bef0b942b4171e6a8d744496d94cde80db95ae6dcfb13306fa17351777faf2119e5
z9cce0b985234b7734ad47e56c9604ef226695ef4345649fadf6602f88600078a988b17b993b1f7
zfc8db10ba8f2f7a541f5051a1b0c298d6faf94b063f380f32607dda725a29f6143ee164e224e24
zcc941ff034b6280889b8df0bf5c77c7253c9966544a3c29da27af307244e3051dfb0d11350a055
zac7073c27a973985e6fa736a7e660fe3f30d241fe70b4bd50a4e1f43e37535a843d78e5fca3032
zdf88dde0b8eb23f6ffa5ee47b2ec0e3edb92bee18643ec23cbc8881c23b61b2228a6b931543d52
z36a0753c5987006e827f9a57d957d508ddf2d8705b49843035402330acf205a60bad091c465826
ze7ce162d9429d420d549d3fbfd3a4aebb2adcad90484a63acb22cbf7eb15f6c766b2fbf728ebc2
z7b61f903c692c711a1d6f8c3cddc0e8edd54831a9bbd5b914bc5e6e1c7f4efdb3e23699fdf9917
zbf3cfc91dae0a6e569380d5d02951960ccae5e7174ab70ed1cb5877e399d3f42e822566d9d36ec
zefb51194516f9d702fb821679cdcc47c44f38a3c63182397b49b3133a9073ad642a361fc4594b9
z8cf14cb618b5dc918fe1a5f13db2db3bbd36d7aabb7fc0e1c4f8345527e5a75098eb4994dd3e84
zccca30067cf029881abe8476dce1b6f3a5f2b1d16be0a02f8d100337d6bbfd4eab1a6aff930365
zfa8f556c3e3b492f20838337e7fae098b26734c12bb5610cae606df3babdc1aaa0db3220cd456b
ze5fda67f8f4bd2b23b65f0d927cbc280cf34237db83ac0c9296041a40c2b1968d2e23fae14a292
z11b201f3b74c1336eb5e6ebeeb00351ac30a789852156aa07c157cee304cba70a3c1e699b25ba5
z4817abc86a03f5fa30047cafda1a6708764c06f713e37b0aa94a4ea186fb4e3b5a6f3564c7f1af
z7f3f6bc039e6cd5b21602f0255ef6bc2b079eb87356f4aad9c92c818e3d932e88aeb880bcb9acd
z20a4f306ccaf861357d5e3b3631354a05f9bfef82b4f3e433cc25e3c980ee2e0bfddc8d44d3d53
z3e92c14a770c9ff0ff5d966aa85134ecce7891d4fd9d55dd7e0e88e6ca49e3c58d602bf66ac584
zeb012607836df96119befa8167901d0e9b5981264e0934db7a82e78622addac934f48650733248
z0d0e487c66587765a5db8ebbdb006a9f85fe1e22b6ebb683e363b042cec8d63134392095d72cb1
z90bae18ff564d887301c09c011fe69b89358da1e952cecd0fc617d8b19009f66ad30cd9c37fdc7
z35d7a9512fd24f38b904e01bf0df3156781235f3ae3b5bc909d4262fa04f9a6f9175230e3516c3
z4d93437e03b3f1d22f2a56dc86e8d4fc9952c2d2c0c7abb4c27cae7b77c12ad153fca08f6ece3f
z88ba242601cc47082edbdebe9586cdbd4e0127e88a9a97ffac07032362fd05774aa41011f491c1
z923740e8f299e4ea5c085b8bc6e17c9122fc597a888a707cd4dde52a6420641894d756d521334e
zd480e9d3f520e5cc248f6b685d5c5b5d60b3f5044486a1039943e6dbc3aad0f11872b3394249be
zd7af453d920e89b6d6c2574c9d425c3f5d896c80171b9d29e239887da439523282fd617f7be8f1
za667580af1bfe288f64fc6b0e9648076bf34cb394239ad9934e90d9f092813402336ed94333ebd
z52ddedfba2488eea0a478a4dcd041d4d324296776a3d06d037b7066f9a465f0122b00b18376aee
zdd8317e0075789293c6a52a0ad03ec41991bea1acc79fcaf44a8fdcde3e10a1365ec07dd48063a
z23e2c02dfb311157e0000b5bc197b3de6e1de283e3e251445e1bcc651f85102263c7062688b827
zfcf4f59f7f40fdd06724001ac31e32648d61ae858155bac36fe1b0021b9f8fa9eef2cddb1e24f0
z56b7681dfdd8634164897b71daaa7cd0f8fa1cc65e23a66b06a9b61781e77c808120e998aa1b03
zdb41b7a338d5be02757c18b6d0dd3dfc1016fe115f9392324ca41c5c8ca44e6b59d8cfe202a171
z8e060c5b980f2cdbf74c03403762bbb0aa1011c2dbbc42dbad966f78bbcb117d7a1c785c65077c
z0bff95c924fb632103eb66798b4e99409f5deaa5508362ee144c47e755a2dfbd4ea081bb9153e5
z3c1197d5d8f4d9105d7043779b85d6151624006be43bbe35ada2cbf1297949734221b04fd8d62a
z5c8c29e3a0e1104e6c96fe914be5b7dba2bb4b25cb46be25c81b68b85b83a400cfa13dc8d09597
z180aa988f906dfbef59a2cd22d5c2d514139e09d5fb1787985b72cae47f687dca74b2e8f6a482d
zb1e03680ac7700058a7e3b338c3db65d1444d70f828f450e2a13b83aead7f8944bc6def0ebba45
z2af00374ed935ec0054831d05cc000d24adbdf900c28f463f0fffc98429e738e8c04981ab14508
z33be18651651ddc8f66ab39fadfba5e07700d667af8c704e1f5a7ec2784ef58b475410f9bb80f6
z7e9dacc14454921d3f707ec0e58abae704606bc6b56339b24d832b08153643ae1902101c2c4cfe
z76bb34c4baadb48d76f4523e32cd9e0b517b145024165d78d5264e40e70bbde7a06c70ab286c3e
z08027b529e5a0b8163ff1def6e65c426b368a0ce9b338cdec0407864f5b5c9fd084781497f13a1
za60f959b830d2758d8dc07dbbff6d477b819aecfa9cd7a106c5a18a317d0e6bcdbe3118a907c2f
z786bdd6af86b1f5a765c4b9e253743e09ce730e4554313305641ed00a5dccbeb3a7934cae2db7e
zf97b71979dec7cf950fbb8702dded69d53646c2c2ed13d914c1874c09b0086e0b9ce1137dce128
z380ec7d1be9510ff001c95f8c510f7c9e0d9e7f5d9e1d39e0361e3fb3749e39ebb9b561c74b527
z82def620c94581a96c5cfef5e59d8e56c4f8bcf8677713c5fc9476141f928924da811a76e45e80
ze356ef6a03ccf0583583e8d0d4a24c8a1f6d842b8c49cb0d8b15ccfbbd975da66a07cb6c329774
z87805d7d9a44b68d4f4684e467f5ccecac32d81434815536c06f664ea18a84c6579e16df0af9cc
z86df47c215a012fede998914f93f22255aabb945fe07a9ab79f30f8d86362ae353938495ad9d21
zf0f4154b056e2d0a686c03986c83b7367e20d48cdd24bbbf63868d85a38097c0f7d4d2279615b9
zd0c298d17a64bdc0b75ca29ccb5eec74f3c860c2a82f5c5bf87d688b93c40e08378825bb404456
z5581a2db96edf2eb03ff2d848dc150dd072e32a9e121e119c83c48a5314dc9336e4fa1283fe7a9
ze26d041f0d48fc3ba939e5d0849429ef5bf198ff489e9128d1e6a85512765b5fc846cbbdeea3d9
z7f29a6ea36f96a811500a8b34d28c637ca26283de9630c7ba6e9a2d8e4cd7550a6862f1892af92
zb062245e55fe5f13d439495268321af8d7c55f17025a74b363b80680850c29efbd9029563cef26
zf04ab57f33a7c72fd6f2f82335280ec5bf17aed08ad46c9f592131d6833aa7505f3af2f79c723c
zdd8dffc4ae36bdca18c69e35656324ec817fbb61e08a2dab2535252b5b92ad35aec7faf45c3a8c
zcc72b5c177e23361e3d0e9696cbd07f089afb714c4630ca53555cce61f980901830b2a637a4175
zc7826914e5fc1b2644a7a9c02d3ecce5ec740e57a6eaf186465191545297ad9b829204406ffe83
ze2151107af69f14260a32c42c961f98710cb01503a2b524a2893940a3d39e9a1381005d469c30f
zb5f251c51f81b683e810ea76ac3e951cbbb9bd620df1a0e6fb85bb9e84824de0ed9c5d3dd9c40f
z33f51f237c7eda01b95e71a4fc556ad59c09eb5d774fc6b0cb235951b0c2a7101b3424e7e004b7
zce46745561ad3c457624df56d1cdbe95949b9d335305ff0efc1665c674bb811d87eea06cae3d2a
zc764be0050be5d6fbb85188edb50fcfdc1fedcffa493b3c9c9176ceae5435d408922f17f7c8802
zb807eb21b1e672e777ba5ef1fd576a0b1d26da04be57b7be6b96116542549e4a76511315d52dc6
zd070400be44654fcb961aef54a245a1ac7412622f142d03b56fac242b096f63ad2b96d525f23c4
zb8d7857ec766a3954d5c083bcf160b6b4954b5762bc587501794e84b5ca03026a235fbe56d1bf0
zbd0e1b97a630c4eb616b83084ea06f01d14c29945dd4f5d6b7fa549ef46d4ea2b431862a0de1a2
zff126de7cb4c55f93087bafb7b6d12156b7d0417607b38b558d743dcc2fbb3fcb87fcd4f754661
z879954d144480538a0dc5f592c9108a169fef61c4a8bcae3298d1dd64b5dbbb5d4b4034c8b521d
zc0de0b2808f0f838abcd1076eb2959267c821d766b5eca0bf423161da798290e7183245a245bcd
zca8eed59d9ce95bca68d9f7934098898b57532c2b6f25dd4678f7f61342e1de2c4ba4f51054e90
zd3e15679d68701e4e0446c0c9465c4f4e5821afaaa4054a973f94f17a1f18802b0306007f8c0d3
z097b0af8eb390fc5c86a38dcca845c71326d5d0562a168d49e23a1e4cbb57cbc348e1f56ef1a54
zde3883fd65a6e4ea05fed625b0c7a56c5741d42d54a3d1ed9f137350313e5f09edd3bf756d6cae
zcbcaf7429ba0b3970d30a552fa3ec94c288bd9e464a67121621b32e14a48025e7f155706c88133
z0607b7657973ece09fff3316669680cd3cd29f0e1e4c22cab1bff52a95d8d1055c7a236565affb
zd21b31bf0d74ef802166f390b4c774ca1c997fba9959efeb52dd36e41cec06bf465bf708b92f31
z80f83310c8a458e6a93a09e7c7b8c9956557a35e818d1f6958f140998735d161bdad4cb87ff267
zcd6ca839078d0b2e789bcce7ea75db6c9f4dc726dc191c0e16732edebe4418adbe4f140c9d1920
z6ccccd9be26f1e9a14544488c87cde62db3dd8d9be5d4e59c4924c416889e9848bbdc1c3cee9c2
zc98d7dcdebb4e9f479ee88cc7f8469506a34253a33f5129aeab8d989d399543e5a3632d6add824
z976c3b43e36ab2007b2444566ec4747a62730aa828d4f09f179bfad5640f326142afc551ee1a08
z68f0eacb7ab114620cbcc2a251b3944ea4a7cf1ab8314eb13663ad4d581365eb9cfbca069cd72f
z83670cb2170105822ef16beccea8fe863226f2c5308dc3b06d147bf669071454ae4ff4a7964ee2
zef74564c157510c5e6e07a9b1de40e8860e65e35eebc538559c5589e3300d5b644d48bd06ba5ec
z5d5b846f1471e55df6db741096dfd8e1a67bba9d5307a8fc89a854eab2e3550d01ef55a279e258
z24efc3a242e7eb0661add7062fa6e77eac15374c2439e37249bc241f0fb23e22f9aeb42b7ed7e2
zca7cd2a5617ae5d23c8d655da4ccbd610e0f4b3a0f66e84870ed80e3b57708222a74f69347c333
z6f5fd4cd68afb9639300a037823fc96c9eb9476cd61ac508094dfa9a33b78e43616a08952b9fca
z94833fcea34d2963bfe60330fc978412d54db1d4459c51702548da7f6f5311dd7c0474314e23e2
zb4b98f2e7987ada119f3560d79bd886bf1ee1feda8a031567c717d188697f2725dfc8eed789940
z6c940a90d0b13c0c721922637fd90e40d64147484dab1717c5e2238c6350e29ecc51c3edced0d3
z181be8f279be875df3e13bad470ee3233bc01f5a9832c828c49add0b07c10d11251306ca45fd86
z52da21b51882522bb2c1c3e0fc9c4c6ee4ede9f616e3511efdc1269a6c672fe3a12e92f6635795
zcc2669a7e2a8caa8bbe58a4d61b1d14891af0c7813d0a885ea51abf9c010fe67e25a7ae550df25
z85219713eaca6090a7022420b7b3424a4e210b51bde36974e4d53c8f98a25be9c6dc72eece38d9
z1741c54cf4c0bf6873c6ad3c7057b2908d9a0a089b29401360e95f9ef02a5a8bec441737e68c5c
z2538757fae34f5de55be86d111e209da2022b98c19bcc6f0fa4b73fb5bb755a4f88ae6de4a8791
zf8ff217ef374b7d6bcd875cb72403120a83dd671184311cf35f5b095ab4711c10fe819a536e71b
zee81ff76bb67cd68e2d1d22ac4743f092b00e0f689a57b3e3ac990564e902e4f217ddb299a0812
z2426c11a2d976c6b398ed007ac39e50f94093283b75a8bdd05a6920275b90460fec0c1d3e96afa
zcb17d277f59621efe4ab5619dbfbab4299e046c0009e71fa0688ed7e95c83baf78d1dc2039aa9e
zc722a8a96168f44d5325c6f9e7318f23b49f6299f105123bcbd2b24d8f69124dabf77a89106d99
z4dec8e2f19a89e267077563f8253b482e0c88204570723e9c8099cff71c007650468df5d5ae08a
z4a95ed07e4b2842c7af84c776019aca4653bf59bb41a1373ac66d7faf88b026551875b58fad8e7
zdcb3d8a675fe939039d4676b58c4f6fb8a3717934e0af71a97abde388d3c8a4dfdaf1c51afb71b
z8f861195b97b27a119f48dacc1a9fdf7df65299a94fb499c5a7da08fb2014d3ef6410a575150ce
zbb132800f0cd77b29806290b04695f7b73665e8af312c8bc15b2beda6129f64986b736a324300b
zc0a1bc8e17f248c18eba2c462873d8cbb61cad8793b785ab5de29a78979d15cae92cc2e63a9eab
z06afbbad159012265e9d5c538f369a68da8d28294a730eeaabd64787fc0324aee2f002b0687074
z68e3a9167d7f13b64b661c5e644151d0495e89635aa50e28832dd2f68a5400c1b3e94b992cea21
zc780b944282a212f57db29191919b30c4aab3d8316058bf4f0cd32d346180677c1ae50047fb8af
zd5b917d1c2bf7087b2a06b3139d6a406a18ecea366e9fbbafe3be0d42053fcc7a3593cda9d677c
za2f82a435e15dc40ff725a109d64a8d5d734548d2d20c7cd55a828abe0911238b2f50093442339
zd1109415437a8b88b21fcbde098653ae938f1ab428fd14acf833568c63e2f56bc5b9ae1633b154
z8fcacaff76a88cfe9e5d85ec79c501ffbd60589ff332af15b719ae92b1b8cdac232a540f437a3a
z5e0c0d762f30013161534cfea3c652ac036a87b35e9ecd83e8f61a5ee59a5db270424aa0875427
z29ac72643b8bd22ecce4eab09e90ff0afa4d9a66083bc4fb9d7df2efa995d9f76a6ae6fce399a8
z4a771c5887ae1991578cbae993e732532851054f565bc13d3746c839a777944336b6dc6bf2a93e
z8d84b6cd58b9d3c33a2191f472ded109350b3714fceabddc63a82cd80e017bd97d23167021df01
z933718cad155d315ccf7b242b457e6a5d153a0ad921d02f45a2a9bda97e8bb2c409b9d18847840
z86133a05f7e90e1544a393f3debaabf98414c2aded26706fd8f46c862675b691dd3218db1293c3
z77dd8c0e864f1064a5cfc6d249912f41902c4271e6b00a6afe2134849fe250931580cb1580459c
z7394b8741d791f7ed2742351c4c96728998e1463ccfb4d7d44ab9206c0a9ae9ef1d6cdaeffb22d
zca58fe05095c23766b39a07815ab7a654d19b8cb26ed3eef5e0135b141dadcb0079b2b480422dd
z4ed1242326544f3038f940bef64cf2c5b87526cdc5203629bfbb84daaa6d360ff31d0c1f4815c4
z27fee4e6565faeee0952d844d1fb56847de04f6579cbeade15230239a9d1e8be192cf0e2bf05ca
z522d79eaf71d7216ead57ad3cac80e84ff34f51fd6a902b0c05c0b9f44c425a06e53f0a2742bd3
ze0597cbc3c322c9783257cfeb61536f5b0ff90b83ca1f18b8c8cf17cecaf65368b42a44916fd68
z99cd1479ca5b3d56990af8759b193b08dcc82aee991cb645ba9030a5bfb0ec021ab359aac4ba12
zc6ab3e1090b290c1ef93d7c132080773850ba77f4ae0d4ce47256f95f4a20fe4a08648c28f03af
z02626447c426cbec507e281515f2b660f844f08004eea12d15ecad5fe4b31fe5cde09fcad8188f
z24522a8f246bb93d7ddcbdcc77ca85f45b6ea0ee78b24eb4f3f4f6f0896a6aa223ab27be3a5200
z5d6eee5cc3ac3fbf79e0210c4f4bc863359ee1eaccb3e9d38c9cf992adeb390db821e248d29b94
z36275310a429b69d8454fcde81c8391fc6374d77357b73a1dc815ac0a4f4f5252ddc7526508cad
z7880ee3763669c840256831dc80925e36e43a55281934d73a329c0623ab29929b93c688ac8ea12
z816fecd0868ad34dd00f57251aa839b648bc29150fca142f9437accf5109d543701863157e44ce
z9d8d9db32547ad99ad33e42febbb7122542fa41579332bc5d9a06c5d6af5082fcc9e57a64f4090
z8fc48d9860031087d0b87da205bfa80345ae30762972acd69149387b93dfd2df003f2f7497e82a
z3246dab75d0b5efd7080e162eecc9e0b1ef6aea39a3e79e93ec6e595feb1b06a161df8214ce334
za306a624e2d24dc002e6ce9bacf437fdffbd5801db3eb3b6749ee5470b722e110f856cf6ae1ef3
z28f69b08fa01126d974675e315840a18a9b56dfc199666b99cb418c493f13dda4a6e5243c6004b
z013c663f9280c06e359388bfea8998012ecbf1559ea635aab5c2432bb59b30e532de865cf56d46
z1819eac9080037820407ebd02f120c00048a365c702eabb34a12a34281a503b2e54e26bdcc686e
z46f3587b3307e2005a76a3c2d94f03148c1541af356e27254f63e3be4719617637475bd09ac760
z826c79695bc94720cf2e1770606fd87b685e5540f936e84486f6dbed5828b4dfeb9ce0dca61ac3
z0dd73dfa44814718fcb02b5e199338becafe3957676d53eb9e23e0f0746be91edbecdbd479dfb2
z766523eb1b7a950d1a2c8728994dab832f859d5a1fb4ebfd7998facc40f21aca23a22916f9b52b
z9da828675f74a004bdab9b3d71fde0af812e134e05456d0593662f9eaa23291ce1b13bd5993d2b
z97c078d73efaf821754c42be29030ce4f0c83293e43433259eae374a5809068c54eb5b32615c84
ze7678cf869f98d2514f6576f6765fa1c6c485510a103f5ba8a4a258200aa1857bba072e224d49a
z6488bed104be7c91fd980ed9c327f074a66ace0539200b795b655f78393497ebfa16863aee051e
zaad4faebaef58d56edc768c7827e80f86cdae35522190ca28f328594b973b530cf98ec5e71ce36
zc7b386a9153022ff798d0b6dd4df32e0c2b9c1e31053b1bc923fc0a09db5706fb03d866ac1e35a
za544502f68999d8c598fd1522e66170cae18300f912b6e0c9c786d6c0b6d881f89093b578b60a8
z4a3047a5318e8d73ff5d0fcad89e132cc1f22cd4a1d411e145a8155aa1d013976f25a6027fd91a
z4b6270d340c3939b6c2762a179dee8cb9a16f6a53631a896d50bf3061d6b9af8389f9b28a635c2
z0e86420253bd6f750575189ccb22767ff648d062d19f54843d02cc1937d7bfaa4c9da99bc39345
z04e8ce4400a0bc39a01deccd2c318ecbee8e3e72d06ca4ffb5a5002047c4ece279d9ef9a0ec7ef
zb2148168c27928149797b8baf31c40770b342e0f5be9cef65a8f4142606878d087716449669d8c
z87a5fd989fa79802c95aedb7b348d870c51600ce3d42cc878740d4aeb8575baa1f26ebcef8abdf
za94be68459b12343cae0a509d37a06bdaae914e7340f2609805eb54078f4f8288d5edceeab54cf
z3997f48482f765a0bfe50857b44e5a12af6f545906ff9514df32d8f03a37cac5628df0d9621b51
z0f4672acaadb031186835ec2eaa85815b3bb9a48bea74266ef09c1bbc69c0b21643c1488903bab
zc819b92ed887c363ab01d1c8306edbcef4e524de8c938ba95b89752ad4c28a44ab175e758fe5cd
z07d08abd78b05b0de80840cf9a6bc20a79d2b4b337e1cdb70209567423c040163e6e00d384d076
zd98560ff4498fc11b79cad0335bc37cbe74d567f2f43850ac3ff32b175b6b8ab1a09caae4702e5
zfcd9857616046116f30bde0357198b39cbeabfc0048f5d33b3df2dab5a61aa2c57277764392a50
zb71b7c73c8c4546e1e16c8d9d563cdd1024b3bd7b1618098456ada2834eb0ba679094822cf1814
zf9923ab7fbe49e8c3c05274a13d836339d12ef5db5eca7da14526d6af9d1f1167a16c097fbceeb
z43aa019c5b9c1e58a4aa58ace2b5cb59d30b5f3108e7200419afe98f794ce30ba6a891ae87c13c
zbf4381e657edb071a99b630c11a9fb770201d05555d478f6c982f9f76943d7f5c5d946b930be2c
ze8d9e65485b8e678604a5db51111cf412bc36a0495b0ae0182decc1adbe471405fb8fc3c9cfe35
z4c2b6a9ca386d79dbcc2113ac755fcc387ee0d8bc67038787898a9e0b590a5990d0d36cf3fefca
zc7651115f2a93ecd2638d56102c71b241099ca83dede6c70fe70f525c8002a408a5a488c0ce265
zddf822924dcd900f308af696563cbc427a082b1c12cd23aad1b002e2c3f6c77d3aeeefaf3197d6
z6ef212560c704bbdf43c1c3f3a9ed7a4a30bf75750aa31ef440210d9573c05d01dba4fea277243
z649b0fb5ba50193e1e19406435768f5c407c2eba1a5a3cc5171ec62122bea77f7123d425c6d633
z2927aeb7fc96a4fd74f0f90c2afe1b2c7ce46c0921a83a1e605698a47f5645b3caadb798356a10
z0496e227e3ec6e6978888379bb81fef4f27c672f5269d46fb71a4b4417fa3c0b9e185f6cf92321
z831389481f0c5995beed43d22ef7d139141a361021b067b37e161004e24cded472990f73f26ca6
za0a8ea5ebc5be26520a260dc1849f7288dfcc1118c1dcdf1757f1118f84f7d232f96b3220197e6
z6388a68c2082f4a5e2cce79874746bb39c70d90b186fe85635d54b706ca4fd1adb01eb5773387b
z9973ca452ccd0d975f1a08ab5310ccdd2a5398603f4cdc39eea35ce710d1b054e49d1db5811777
z55c12ebf360137cc1a18faaff3f9bb87c083bc0ecc62d0e04b248f71872362b89127d9c485cf16
z33a533a94be3af1c2a9f81ba80168e4b45368ded4d01541e3d4af25caf9afadb4015f98962eeba
z82d85db569b3105a87059253f4f52352245be2492cddd765a46693bac15e7b8b84fa41573bf461
zecb7ff323e20748e86b9e846a1cfc399deb1f81820f9462bd44baccd629858d84e658405e020fc
za2cfe057fb20e6e6f80da5ba48b6be7a345f6561fcb3454cfa28e7a9b3e478907b936b25be17a3
z63cbb385aee5e5b6490c344260297d8358f09a27af714c343f1824d05929fdf45c0fac3092ecfd
z757d024736577ed3949c4de29c36ea43958b86a10e817684bdb6b3f5c6ffd7f359cfe0edcda9af
za472605521824ef522157ddd49b2ea796d94677deeee5218e1c0a4a289a8428103586b08a8184e
z3c772d099e256b566338e63f5188a4cdc3325347ee513345e7ca4560d29dbedc11ff9e431d273f
zd40a53e8a0c571804657e2bea14028a93e157e1a0c4d4a5b1e4c502b2bf542bc714842efe2d83c
zff3d5679f8ab8098ff3e55384a9f70cf5b96a69902f1fca26758dfac7831fc5e6c3a5f121732c0
z9015bc85c94153a9a5704bfebcda0a91e64b3ef7408aeb439f13ecb9c174893efeecc953040d54
zd0e850116fdf3e5a9035c0328405d6917f86646e46a8da3909955ed2d0ec74176f0a4256857ab7
z4e7d0def6419803a50a959f8e1b63ee819861a0bb6d5866b35684e28fc91057d4d288c317c8eef
z40c2b84767bd61ce6f604c79c1d69d5aecc0062ff263b450ea8780db780fd595a1fd92dc4c009b
zc2b30e2b85158491b4a96bd03f2ad04f82292fa89acb8eb97abedb11e90a7b7dc173f1752421f6
z50d905d782336fb05e19b2142d7e4c32993334cdd396d019567d11063aca27d2eb1a4d07492a28
z6342341ee00bf35e39b0c6d09b486cf9540f7277bed9368bac10d7163963c6ef08f1549388d18e
z580753060373c476f563d6db934bef999e2cf87b05189bb6549e9362b5de4e5e125f55e177cab0
zd59e440a626e0ba82fe91bb908f37fe10a65e913dd17ec0a30790fd3c7237a7a4eac764948c03c
z4cb7086cafb84a0e3318107cd479ee577ef468a67c27aad1c3908f475ed2c78dcfce6a9eee8c13
zeb294f98dee2b0f0bfb8fb7d865b5ec128dc7fd6fd51e33ab5231ea8c8896c6fab2d145808f46f
z1563a19c3b49f9dc117461fc8a771dd9b843dcf598b8dbc38ce19432e5745e470bdf0461d76213
z869b68d4baabaf97f0b980bd11b83cb0cb7c5f136a06f294d8cf8cb76f2b9851a2f661fe2f4747
zc2dc44db1ce94c04fa74702c1a545190c33605f79ce667018f18890cc8908126831348c089362f
zf30adef09e7f6a00039e8ea454eba4f83f51930d67936f4edcea68e020859aca9cd2767b8df8b2
z973ec640bb994fd3c632d1f48c5efa12fcae151f83f5c2397e4345fb96d71d565d960deaf6a46f
z442235599c03e7673e2426b661fff4f14312c99c0cf92c4a923b85a2c2b56c3f0726ee434ff9e6
za77a392b6c06bde42a2a3c324e66742c971fbdf6aaa8d0737fa37ff0176813a3b74f5b32ee9bde
z6ed42bac419c390f6f49d28dd21ff8d3260b1c7ec7d7371db615bcd4f42c56fa4c9f6b55ef8393
z01bb14ddb52836abfb12e694026ec751ac7db061b32efe7ef002271353bc4bb74bc27e483671cf
z0b9be5a9f2f5ed39f903cb49c082fd9ae7754f9225c8b3e01c95655e2d75bf5295c9b9c3d46877
z85a6f9f741942213b066013002a3913850db52f3a54b27390a1cb94552c808f56f7b4c5c034d87
z67f53e5f266122da4fccf1a650fbbda1aceef42e246868e00acc20ca1a7b81409f4bcd16704d02
z10b165e733990361753b242ff2b71b3eac7e5ac11357555f7a48dee0a3280ecac9a7340ed8ab60
zd5eb3bb6d27506359cf5281c1973b72031bab1506a4af6b6cce27ca2ee25ca7098e7d397220e12
z5d4db0f723f18d2d5ec5faf1b225ef5ca71d879a6b6ff8c7d66bbd40eb3d4e1cc19d41a97f95cd
z3f18f6450570e494fc40f6e9a384329feff8258d0e08d90016e9629a3767d991c713f22bd5ffef
z4348475b678f8f101399ba334dea4a1b425d902e86090c45a88d1c065fcac96e3e9de033d2bb21
z843937de8171fe5e1420690dfb00fce1ce63ba1b46a37af1e4d656854e9250ad0ad5c6a47ed29d
z59911693e5a623d48f09cad3a0f29629ffa7c8ba3e999d618da379e803d7a48bc07e20e2d6b6e5
z03c29d81007bc9947cc5bae0adf0ffe908c342e47d60508a12f2de2328ac77ea825c6e650d0cb9
zd626d00f361e22948d26482a7ff39f12f646b4320ca2f8d320eabbaf77c384640ecbf9336ff166
zb72c60a9d32be288ff3e880f3aefeea414125acc9f01409e946efca7eaa818ce732e482d858a2a
zcf3add0ee547060cade779e92c9e5ce3590d09124a655185883de1369deffc9c9fecc93a2afceb
z893154621e49eba5758d971030cac8995e52fe1d76bd2786877dc0b703dc23c5c78575cbe23297
z6f4b51e370c2e1e4d982c48c934de65747822f0c7be22cd501c15ba40e28c475c6c345eda31203
z7265e9b582ddb095a1cccd2064726f146218efc95b34d8dcd63b1c670e341acf1917a00c31feee
z767ebc387a6fc9de5eb68617aa1a2004eff1912da0d55cb206717205a5945a82e21244116b8197
z876193f5b75349a20dede18342fb3216e07d24c4b38c8a828413b742aac67057f1dd12251b27b2
zf21e85baa7541c319a53701e6d41e5ca31b90663feee1ac4e88a28dd5da4363003a336c09626f3
zb6ee836d1812aae592b631b35e0756f66f1e883ba19e876553874e99cb7c4045a554cd891c8dd2
zd78ddd14823a51a67e2b43f8e39fc43d578f2be12da453ba28f6af2ab8b3acba9cc8128159a8d0
z87974c65f2fd81bb8de8eb8367bcea2c2dac3f7744c9d9842d3959ff1d55cfb13b03e1b4e33865
zed3b82f21378c567ac2766da00aef66dd17b7d78daea985e07efd85f391760ece18b84e4e3f776
zb01bd023e5c3ce832e89992f9d2221ebd1538eb306d102b6c5c7962cdeb734f199322f9271d1d0
z9fc8e68e22a704a479300f9abf55c4e4aac86c16ceb9d35b482a76ccbf75ba8bb2af5b7f8cd829
z7834b531a28d75af893f29fe9c4181749c1f985c392178b222a8768ea6d346a9ebb9faa07571f5
z1ded9a87f877ea87c1e342b678fddbb8e274a76ab99bc8a80fd1e6ad27c21f94251f43c8a0b896
z1b6541decb42cd1a8c7a0a0c897a782a3193954cd47ea341b1525131f3a40258ccf9a41d2f9ee1
z625e167299ad4260274484eb96cd6aba09ea7a8cf9c2dbec47f10184e69512d775bb036871ff4f
zcfd3df53189f9475c66e8bd8456799f839a1f280b3d5c72dbdf230aeff4f8369eaf2be2455334d
z2a48c8dcb28808e75729c876980940c0662574c09969dda28c63a0477fb4438bdbeda43edd8920
zfd3becc6723995c372ae23bb6272cde2e41976c219bc62c3611e9e2926274a15730169852f0948
zdfb35c27569ef8055bf6cb63a73de17ae3d853caa014c58045ead71a5b7a81bd0c587922e89694
z08024c8978ad90569be838b24eee24da97df7fc6085dc0e6ba3b2f65984c300671214baefe24f1
z66c520c83659ae0280bc45f77cbf37767b5993f94f32a11d54270514e6a0657ef1909c02cc73f6
z6a50338c1268a34365ab3be05125017ec0237b765daa2515271f7e2763daffbf8b84c28687d8ca
zabc6c2e58bf3e2a34757fdbfd09b6ac65d89cbe981f7a531c68d74792c6c24f59cfae1c945d3e4
z7ef4b96bc454630a3c92ae6f295bd48a4d06755d7275d6ba1b1c67866b1dfbeaa5abdf226b0a19
z9d2ac2210694baa977521eb997904615ff9a93141e0a480a68e3d471cdb791c2a43964e64f4cf1
zc38effa1a88070ecfc7639ef41f755619d8efaf7b352def6d8a95e804db61c6ec79f6a261cc258
zfc235c52e9e82bacc1c8de1d9d79044517212f3d3e8ce0712b316975a200067cbf3550bd1b22ea
zc14f8078d3e8452c4bf9d8659bbe90f11f2ea177752d2d32aa4e451e47a69431247bfee47c629c
z92e7987534f6bf9490ce1a6f4f217357e826255d92bd0b1b15406c17c2b169aa2c4ce1fd4d8ca9
zdaddc6249b250b2a76c9382f1b47e82f33ddc777af2ceb0910a045d5bb538c31a9b59526d17bd1
ze908c5a791aab5320d3f91ae04f0a6a4c56541e30ff5d8cfc7b0ceaa49657fe4ce57701a130634
z55812c36ebc6c442cbd2a5ee6da62917fd758249fcd5b588caada9b7cc980da2754319af9ea256
z596402fc128f0e9aca46e73c299e1dfa149218ae64f76cafe9aae4a31e0b1c884b7c1da0a33952
z41f89283365f54d5d55663262f4ed6ee70ab6bdfcdba480b4f0e076a6615a72de10e5567c3df14
z426554b10c2499894a49e0643913f8a6091751a7b2f1e4599874ac0f508fc77dae6fef3985cebb
z8497888e97a9b56206cad45160fd371775f1741760a9ea4918d30f30767db1688bdc0066d31b99
z3fb59b49112f349d06fd59d13b34514d68328308a05383edbfadc868fe4c9991df9b40beda446e
zfdb55791c3f816a4bb3d8f34b1eb6a0fba0bbece49d51292402e09a068582ad5f8bc98baf2e584
z202bace8de371602f8d12186705ec6cf769dcc07a8eb9a3942126f0affe0984d0f06d3c60609cf
z87d56aa64629e2528288364ba20ed810e173e690187c1ccf4669c2ad1ab40f342625243add6fa8
z780cca9fd80f3be5e3610186df108fe105288ff957d0bee8b51e3eda5a42aec0ecd81f2e7c770a
zcc3b1d3e999cf3043e2735bc0645353c37f55f4192d0ad45c8521f6a4d2796a2bf92b22234684a
ze7d514917b2aaaf998e2a170653880db47a81943e0e97f7451bc39d309ff15f73a88b048f83caf
zfb4bdf5fd4f1b47853c0deb8fdaac424ecb7cc30d31c79846c9271d08964e0c07350fb8de384bd
z559643b5645cc583b120c010b39cd38cd97097602ccacb1f725ee7561126b8c3302a60d2691b8b
z1d54e52549df42d833eb23def57da9279070d4e3d765212a216085e3c89a48453136f259a4a6bb
z9855738db2ee995fed06bcf3f80cf398b307bfb0abe4e3304c0cfc23ea80d6b0aa5ff4063b6e59
z2fbf23affd994792ca9c724e8474d145bc6aee1e209722b7d9764f295cf79b235723a7e70348f4
z95106c2f5f2ade8c17025183564b6def14880ed345849b43745971e1bbaf5037df2e465970dc5f
ze4190b2de6c48d9bc68fec7a26fe1a83155ddeb20576d90d5a36013c65277cdfab0e80a27cc132
z1f6fee52985ffd92e9b0d1914b75cf81a0906fd1681e753b71c221219646086df3a186cab5d607
z91d58705c8aa4c153c7a0f3c00daf8e783ea7e58786d35db055b2c47e6679718433c1fbbd1fd14
zb92bc34a656e2721e05162e5058b3eef571f3df181f1d1bb8e7512afb38b0eb5d4916061abd6d2
zd3492480657c938e4668431b447f26d1d40d0103426713ae89f7430fe914e865abe28ce9715e6b
z85ec454a8b7564c7f022086fe4cb447410a5b2cfcc7dd848b3e93120f49ecbc25ed9f10c34f29f
z1e06e7c5e5b9f3270916a506c9c76677dcc2a13a1b6fbb39d752057803f6bbd9e283ad5b31c81e
z9f452f0d8365dec9ec0867a0fae62e15ca5bc8447c46bb9c53985085794b16eea1c80237372fe7
z355444cc190cf10ede404d62b4b1adfa07944556b4c9008c8dfa2b6681b8845d4e73731f0c13dd
ze9648e55cce198eb10fc78bd8c94d53485ee7203467e90606fb407ebb7ab12e73295e7373ed2c0
z50f074b50540f9b96fdd38af9a5589c12cabf782dfa989b15eec3ce95f1bcad4740d1c5ae29c9e
z7988b079deb51c314c84835158c99c2d69375c55689d8db2ec886b6b0ebbef5c458d3c2f15ee3f
zda417b8edbbfbb10f25af3d81c0fa6cb16428e293c5fafb2c3e5cc128caa09ed0989fdf62afc20
z0d879780dac2ed319db4e065e75232c0411366d05acc581d62d49c52beb7798b49d657a673f9f5
z37b6eb62fa02fd0ce0df8ae8cc2e959deede30f957017d0cd63ee304d0724b1683e98a110e2ff9
zf1cf500163b413870c10b88d01500aa85796c99f3569abb7bc523b20dd40d04822b4f57988e74d
z65878a7aa78c17da6f14b21539f0fb37403e38b7698aea396e076c18ab47345161f6ae9e03d516
z18bfd23f6e697661e1774b3fa9be05e80c36da75ff523fbc9d5e7edd5e1d34bba51f9b660e5c0a
zfebdd721816bbc1e294a02b2d12d8b0e8d90f7b51eb800efba6ce00ac15493f54b4b0097bc06e8
z1b6578592fbbee1aee9dda98ac6aa517c8f0e8f6ba64fea1cf28729580fa70f167cc217b20e9f0
z601033bf2bcbc5a3432fa6ec9541d15e440a5dcf4f84c63e403fbc3c9a9f2934eec8186de3e2b0
z357b541c52023ffdf8e1ad794badae67e640d46b6b0a4374c0a3c747e9e7fd946cddc7d2e84585
z2df5a66dec8abbc50aac9024f04ca949134611f448f816b04ca593c9168f8e1741fc5e7b479804
z802c0f6f75c2e9c49ab536b76524cef738eedbd64da7530dba8925c5d5c1c19a069b06bee41dac
z5af5505f35b13c4fba64c8925c7b7cf9d13369e4691048df283abb676f1bb7af96a5f0a9aad10a
z74255d67ce5467b2d141df6eb17a56f2e997b371cfe3dce648e856ed4b15e49d0d8d7ced90a4d0
z67b53d2bf8a0662ff98ec2c491aa1853a028300811977ddfdc06ce633dbb382beea814df3c9e20
zd82030b4f56e3456960d2241021bb820a53dfe547a5286d8450ed70f3e4341200854efb2ae1194
z833edc0f42352de0480870e23fca74cd0756c6e9619a2f2892771a24d6c5c67342d4607ce91886
zbc9a93271d849bf850d52015396f80cd7cd54b2e3226afd3cff53f17428800629f02f8fe289c97
zad0eaacd48d2e862b03a25378debc7e25c29099c37f3d19311c261b069acf8a32fa1d162327202
za9058f8c9b9e6fbd8db098de79a553e8642f137e8de0035f72a7786ce14224eed386927ed3c3a5
zbac2e2215024ec5e6e97b36e062c972ab3e9e797c679693071a1501f65b7d9c40c1c4d73acb79f
z853db1a5e7aafe1b418af4ce5e5cd974447a3cd3da0acfcd5b0200b49f1d21cbdf1abde6198b1c
z0542fdef8dc59d48fa1c7d4a375914f2183091ccde37b6371c5c894b4de93bd19b1ec4fd998ab5
z3b41765ecc93da45416685f9301eeafddb1dad975ff2eb7808b4eac170b73cc72d735268ae4030
za113082ac3a35223ff565f7c12353a9ace44e334d10708f9a1ef9caa3809bafddb007b3ebfadf5
z944f5371a0d590e12c04f46913269a6236126888b05b75315366091c399a5ec246748b163de33a
z92c39654b9f422ce35f37e2a0b1f0bb10cbd5a8c46c7557cc963e4db9a319bf8a2c057feaa665e
z392316457c57c934af20ebe31a366689e7882964f5ae0f76666075eab3d480ec6191f57e355758
zfc0f68e4fb50547532cd345d1ddf04c1b0c43ffb65e7d92b03cae633128010e86328fd77fa2228
zb859a47c53b1818a284a4e58728cef969be0412e28ce4a02ef4df7f4bf3e8f68402038ed4e711c
zf3ee72c7fd56bd01c2a36d4d2c33b31e65293dc83572632b8312d27d671c164739e281aa64f74e
z747fcfe7fb6827067cd6d969d02b60bdcf54c516698524f8b8808bd72514bc034da259e85ef718
z1b1463a204c578521a759e5ee360352ba7c6a2593894b6e0a60b4b40449e4e10ef10f9d683dfc3
z2ecc85a743d0835ff0c87d7eb1b946e81bcebda13affc877d737568bc61818b81e2eab591a1ff3
z2099fc85e04e60f68f3096233e1fd119d07b45a72d00299c08cb444fd6963993d77d756508c4fc
z97749550cb11e1784606dc3852b3b3d18f3b792ebaf9fe899c2792af10d109123beb437e1c2e42
z7a713132cadbbeca58dfaf6bba4e1f5e828139f7312c964e72305e87baf7d3a55e0316ba92e067
z63be942fb3c96cbfac14971524125957ca9dbc10837b75db8797f4362c210dcb278571bc60646b
z30366267cf382b48dabd282e229eef3c80aed3c51dcdf181e68058b0588e8cf35d8028e870d19b
zec3ae4271ef964685e1bfab366b8400c82fb5ea2444bb9bc9cb2280a1d63d8baaa0ac4b4a00efc
z9fe1bf4780a6b9b3755427c3f2cf1ef89db29d99a115622df4b5e05a2b23b2dfe3aac7d9074a3f
z82180429f4038ae82634b69861df7860f6208dcefa36232f7fe34938d5cb56b3a2511372d1306e
z5bab08cc9c6461ccf3d65c2ca522215578a5f3197330f364275e75ea0e9fb326ad60a618f3c34e
z1bff75fcb2fcd2e71ceae690bacaffdf5127a0f0396e51c61c07da8593033ea9a30dfd32cfb17b
z734f6b9fd2efb9e728fedf3020c13ae8d29acd78ba661a6f4d913273ab6b695b6af73e227fd561
z7319e04ce467c598bee5c8a2f00b8b21ce58f86938eb16116e70b38947e0d54891ee8fd4fa7c05
ze58a9346f232ab0a685c0169e7f49a80df340773252901761be74f1c7d8fb3199b6963b2ef1d2e
z4fb45b3a35de7effac56d2fb2d22b119f1a5d4e737d8b347a01c55274a1a713a69167b0b0c1c86
zfd2218b943dcac99ac1a5eef6403fba560e897387bd0ca50a26cdfb2e87a4443461f4fb58fca22
z48693fe7759fddca1b2aff681794a2b78a1ffcb536937a10e4b88ada247471711fe7d6e27d8f73
zd02a3eb211217232222751c8a6f5216c4ebf15dcd050739d706f663769366d3b1b234f931224a9
z748dff6612307674c59afa3bb1fa165ffd2ce1c89f2b97b18df93e66d69aad70ba663fca12c63f
z586aee11ea123b806e5a11c9a103625644a1140cbb4d31ce06b2a975541e4c269daab8eb89569c
z81ea2562e03d2c42f7734a83eccc64fe898c1020a76a9975528958ac6eb17c916af95c452da2f5
z85a8d97f811ac2c5b2ce4cdf3bdc2bbbe213153bff527c466edb9eb030400e339203e76f09ce69
z59318319e9a9f762ec9bded5aa85499d90d7e4b5b02ea03381b32f8e36539ae17280adbd7e9243
zb48e6cfa14572edfed90fe70e53d66b7054c7b3951d22d5465e84816ab85b6b28eab2e1846c4a5
z3e03e199431ee4c60b1276502839bb6dd31d486e05aa6ace43cba0a463bbe270f125c3c65950ee
z49f6eb486848e2663c4f51b5b3abc8811afc166eaeed840d85fc579bee94959fdfbd4081b6e720
zc68e8aac219b47b1f3b9f30dbc4abb8d99d392be152bf4015b02c0e6574167d66951afa319b44b
zcd4db8ca2ffc599440276844d364caa0bf030304239bb0ac255d65c939fd931eee20271cd75def
z064ee07d49dc96453ed8ab57016c0233d743b101614a1662c00623f539629b8d04e5bd118626c8
za8fd24f118914d350049408e73f59c77877c4a12eb4a0c9d05de8ac1d7c059ba0eb339c38b5e31
z5ef3c72735098e6f71b01d4110c0fd58cff52f434c3ec9f992e6ef7ca2d6f67a93608a51a86872
z635a2bbbc62ca281e3a5bb0bc1d0f52ac26bb1b47dd7f4ffa293d74f37996d5cdfdcab98f27e03
z0039f70d8e1b32c8c0343f0d83f3fd3769a2a885fa9e0527fdd81cb57b85c29807c9e7380be0d4
zaf39352268bb574ae89f1a5ffb8b7ddb98bcde0626fd12c745b08d1d00784fb5c9f545bfa29463
zdf053a385fca1f74114f8db8b223296fe44ee97df0132e923c584b29e07b9da168e70784e17a4c
zf8e6f2fa049c86b0340db9a0d7c27d54c3bb0c56113ab30438c5eef13832342f9aeb55ba2fb611
za7843099cebc1e1a245f826dcbae571a6e4fb7c084deae52513387036b7e027b8e607e74b8c252
z29dae992a1d4fac3929585ef13aea08145bca3ace078eb5e97a4677ee697ad5e7ee459374bd91c
z37203b2f95906170ed33243140d3987e4ff9a6bbe29cd64fcb6bb82f1ec04cdab08d32ea690d27
zcccc1d793c9fc52f772769f886a22d069ad18987ef7f4004bc5a48ab9097fea6ac78b288c088f3
z9403f6397ff200fe53db9b6a387bc3a2985436890194f89e28562c7b5251c59777cf4a910d2851
z5a0c1903af5e909198172d154e8d70f64c54dbeb86cee949da0ba125cdf50e2339a4ae213d486e
z4c84c9ec7b9aaca51d0f0dde907b26a7e7a563b5820fefbd85933cf133f0896ea1d39fa60a1f8c
z86377b60bc874f23d4f8e472b24cf66102e48bec16433f1421b9c10c17ac9d590de31e70b2e220
z7974765082723588f5cda7bb2248b6826f7a19ab348fa6309f383a7e0c0383959efae044d30736
z3c104fee9a3c1b7b65d7e6d1ae3fd6aeba29ddfc8afa63ba88dec60a3d91a47121a57255f966d6
ze263dc28fa9530c547595e0c1b718c21372f1c93e7efb31cc2ff51d9fc7a9a08076b3255871201
z7a596fe87635b51a98ab53e7ae35235f82b921a9b34bdb558050b2ca96fdee427377a14a1fccbc
ze269a9cb6551aa9dcd4bff46802eee044db33245c5dabf25b54b46a7113f276c44ea4ce872a557
z6bf81167d46d985f82a04bda089733a30a53cbab43765c908974edf5b3350a5e6ceb5fb24d2de0
z85ed18aa09ebee4f79ae642d6f1e938d6448a3c104a27d4cf853e7b0d5d9b7b8f14fae602d93d7
z7c1b4216e7628eb6a115e6d6eaaf928de52d5f8005241d79ec73bc12c0733c521e8b14d78d9f47
z52811070e0e325e65a2b9bd5af8cd7bc90290cc002533609d440f6033ba7ab0abd30c6a9b94fd2
z2f36ce915abf02012c9f6d2caef5221928a84a1194c3a16abc54c13214c438c52d63c155ef299a
z9acc127745b627b5026f27a60699ffb7fc7789d437e80f751089d641464dbfe5cc836504a8cac6
zce4b776796a4b494c5acd007a960045b75e1be9e1ce9f6422e726341dcce8f5925cf3f0c4060d3
z76f7f2ee18fcce7b908a53844be63d2bf20567d46020cd3241c2d272af0440337d09206afa3ad5
z95e6b21eb6c0cc212611ad72baa2ff48303e31c9be8e209be83ebebfa183757cb6b6dbfccb49db
zf0c9a8d9251af4813eff58e5035212c70a6e5c8f5edb55daa11ee2563f73733b9ab479a84099ec
z22a656c319f68ec5090214eb3c0943a33329926ef0b8c05d70515c01a3009ddcdce664c683569c
z4a193cdaf34320883f5c6964f6c103158403fc5280be83c4849e0ad3865e0da164639089d0ebbe
za2ac73f7e4174046f359f258a930946b90914ab3c20b9a8372dd212602d7d187c19feb8b9f630b
zc299be5c7612e67adcf0150c17549cb9ff7e7b0098de12cbcc263dca9338d39c93f57f45239c6a
z40c52714d6dd7f49cc0817d4304f9c62bc1e237d0207dce211609588d0c0fd44d542210713e5f5
zae0d43abfe2d835c36bab5837a78d7bc3eba15d3ba682233cb92655fb4b664bdcc93798459d96a
z899e7bd77ed29f343d8fb0ff339a4deba23e4ae101a6a7874019dd7b1c8d623a531f3c619c66c0
zb32a9100f4d07252d2e183e41ae7e6d754f2a3a1f3440a7b9ad410ff8c69d6de0e33339e005267
zf7e98306c1c2bd18312a42099d223698be958e10ca24e6118eaa036cbdf9f06276fad966c39df7
zcf35d2326558851ab49564dcb27eaa9d4d607f0bf887903876ee0f334dad160397300643eae6b5
z563f049ad0c439f13be562a6a447d7f1b2bb0cefb1aa5b71535941154d3cd96f2a4f450411e03d
z28c7535059552bbbad7ab90a3e5cc1cc971fdddb34fed795a18349b49eebd5323409dc9e3aced2
zd4179de8fe3d1f4b2edf5e83f7cc5ac7fc356e8778d2889f6a0060dfac04099fb102c7e8252314
z1679bd8ec296178e9fce562b717eb854b19aa04806c6e5e7b60e8670b17ef018a2e940f0662c8e
z3c5bec2e6ab73ca30d1416e1c1ddd84fe884e7215368462c81ddf0573aec617156073ca3faa4cb
z39d15ade84088a94d3806b95344c0c02775aa14e4f2f3ed71c430fddfbe3cfa1cf04452ff41af9
zb966a34fe2ee983aa978e0876f237b8b5274b5a1f12141d460845e0501364d6053222f9e2fede5
z6e1c97d6efa0ee27433b918415e6bc56cb3739089e9c789bdc05128d600637ecdb06d39543fea1
zf308919fc0935efca3239421d4296fb97ced96fc2e13ccf317616d9a707dbee00c9895292a9f70
z2449b14b59c7b2c3504b711a9b7a839f0f0635a2b0df8b7083464f68184efa58de6e3530fe849f
zc8e4e6319c7c925c2481ef2d33d936e24868fe27c2b7f2689a5320ad5c8a762f0d68f2c8c7f84d
z8720dd5d6f0c292d4a46da0d97408c41f325d663ee8bf28a425eed202c6a00c5dca31437510afe
z4091b7f561fc5effacebb4e4fd8cbcdfb8bb3a605b6922af7766a1bbe8de6e51ce2c34deea714d
zce885fad9d5347e1725a89671526d0f99b950ca8c8c502737756372634cfe73af850d56ffaac93
zb69d72ece4ab6b61d4127b18e4e0a0e7ecdbda8aac0c973e35e601dc95146464210aa9f3cb5aab
z67a19649aaee13f90bb31b15bfd748927dabaa5960b5ddaca3faa3057b18086b575745f019d870
z8623b9bcd808093686492f3b71645b86d7041e4af7942e848647dfb78610744350bec4d18797fc
zad2423f4658f791357fe1103d3893ff5d368dae815a494a7f416e7a71f6e2cabe167e16bcf789c
za1739ab559718af85d050d53a2b4b90ac88a3cab5a8ab71c2971e92d1abdbd00869fff993a9fe3
zf10c8ef94c335cb0604bf01133aa5e789581454b95e6f7a7efe9abfbbeb98d0566e4372d7d1083
zae705989b6f1cea6386d8c9065a7410f08908827c70023a67590aad62fbdbfb75c4fa47c87794f
z7769aa9451694f43528f6ecccfbedeebcf2532d1fc2cd3d833193e9d2978a7239176f0d71a5f7a
z13a2caa9d02137363aa41689c7e8abb695032d3d5346e61a3fa8170a7290c169b06fdae24b8405
zc63ed6dca53656edd9402f8d03f9cb0c40aa835fca1cab1303ec8f255d836d8b434821b5556920
z5c11416c4e20d3b7f62af335baf8c7de2ee2c21b14b598804fa8ec9593fadb53e27b8c8deb593a
z54c3b553343ec0e5bdd5bc118fe8b975dc5ac177e0e309f251589defa301fdf7e8436a3bfca326
zd87a9a89d0402d04b897fee03779e1504b75470fe0c8dc5d02cc898a4a0ef4dd53ac0c649c6d39
z437f538964efdc435066d59aa84e45a199c8c54c9d5b92ee4a2281abece5023182b1785c7447ab
z50329149d2e5db8439a2613eb2b26adff3d9b5bfe7f71694c5370a29070433302223719c9a1fba
z22aee3ec892195c2ed054de1f87368dfc6c4b3ccc5e408f10c24154e3af8e39079b5049fd4cbef
z9aaeb0672b2917a50848903cd82bc66000c7a6bc834372c04066c96e136e800f4b95194f65b417
z33d81d7fb4f009be567c06495505a218679ed02c86cc418ed82fc845c50eea2e101104c205c429
z7da347570327085847627254791ab8029d86f2980053e669bc401e09ebaba6f9151cb15bf6bdb0
zcd2ee89b0e34206afcb77a12022b8bd219224497d8cbaffb4185f22316c470374962e74197598c
z2764823431545be4c14b8e5d2484aba03ba80657d55d195e05360795e1cea61579de253f781572
zbb7272969274124a5cd31194d0794af13f8ff93457da8a26bd313d3f5d7a8c77b4a4dd4a743d98
z2afa7285460feae6b10fd69a8a84fba410cd676691537097a7db9115992b51c9c1471622e4f275
z6263e1085b82a63ef7abb114d16f15f0cb9a4fd808703a67383ccef3835995c4a56896e22bd550
z6fa1123458969beb21fdf3da358ebacd4d099b95e266a59b702b688f961086ed8329d4bb804a25
z27e0fd4d404619d0afed4ff8ebb11516696193b972b62d6fdc3ecd246ccc67f3b3dd6ae82529c0
zb1e6b26668610f20578602269c5f9d921ad60b96e92ec1d6b0b4afa59aef5673a54e090e4b2506
zb1259cc201b38b55ec1f028424c824295e9e02e756eed1ce35d57a121619e72c738081226a3148
z2e819a42bc2e007e1bd5dec827306da92a1ddfd58894f7954248bd197f3a3e415fcf9843ada16b
z635c1b20144b7afe6304baeb20f73fd57626bb010e50c91dabb089c0d42d9685d9c32c3f9e993d
z13d4452d5f369bbe288f949f1c89a28c0f093c902cdf5a7e199fac08ee19725c7565ccd7a1881b
z5308a6e125e9285a3a684f1d97eddd59138baff986744eee77fbbcb4af20a0dbd5450a371430ea
z786f1d6f10cf47a9ac8fbf71be3da96dd4b4c96732fefa63ba5f88870d1a133a7c25964328f462
z04ed281e0196ac017767ccbdaf29e6595ede5d45066efbe762351aa663ebb77474e379cd97d3ce
zc201571e5c757e68c02de34ec5f2ef9735a76403ad72de35cf39ec7fdcb78207b329129713f1a8
z544f705ccd81290187026facae23db0e1215273fbbcbc78ecd411223842fe76f10525a25ef8c09
z30d970819047e05c559beec37cf900faebf910b2c43aea96cdfe372c444306e048dab09c76034c
z434fff80120bcf5ddd84a37d775731ceef54c76671099debf8df530de377e39bf85bc7890f14c6
zc2713e99462071ab1b2aabcf8c09ae682615948d5147755dc11caaf1f9716ec038014ee108868a
zb5b397d93ce2a9327e5ca04f19843a75b5c88248173be5c1b6c12fdd6f4c16105e35b140ee6f58
zec16d32f8934c8d0fc9d210a6abe3a2038695d5eac2c72b2ccabfd4534b8cbc8a0b0fd3afc0ce6
z5c3036952f330bb1c579e4c79885e7741b796db3e0447c01ba4f49d4c316b219dceea2dd332943
z9c3be6280878d0d7aed3140bfa787391bc36003cc3041c8210cbe3b401652b4bc6ec61957c391c
zdab3c0cc262dfc46300c432f6c08da3c3323e0d342ba5d1a08f95eccb17174694474c3d708eebc
z8be64c66d0852632bec72232074065422d911f6e7c7c6e1d1a1734de9353cc67d97416a0de1ab4
z2498ee19c941eda751f5af93609e5bdcda1d6d56d34edde196ca4414d124f4d06d588ab2b96d99
zcdf55480e5adf5952d1285942b7f842e9ce02f50971cc09b0e84e0464521f0cfd95ff4efd36e03
zea3002ca2849016b9340f72455896cbbb3d642f7e4da140300e98c08de0d98d3eb781c3ef9c0a2
z65c0a78f3a7453efdd5d9d709ef35e9e2d3dedd872990353570c3c9ffb50d7e984605d6760423d
za6740c341a4fd72f12bec8f4e0172c6a8c39ffd552477478c192d5e51216dc138a2d4c2b1c6ccb
zc09ea6633d0142524087b05cc958d47310a8b1ee2fd6446b09ac7b92e0c8541e3cbe710446f592
zce735b4a554fa8bf2b2f97d27383a2545f72302f9ba3642df180f27fb717a0e5514267493d4ae6
z261a7b32b16900525c68c7e6aab531faab44975eaed7182323b309a2f7ee5b23e3126606540912
z843eb95dfcefb1961c09614d876f1adf873966cef464f25fa442904d03a233048b2cc4a606027c
z84fe35c873f15711bcc74e921152807385092c5c029c1274e5539fdb8c51fc55a33a49a96577da
z586b455b41a25990e8ddb5d87e5fbb1e5d9139a9896c486d583e4be0b2a3941f2f22ef3a11978c
zfa552a01c36ee8e815d9a8f179bc42fb63a84379d34529cd3053d6ec6bc21732ea91fe7c2a01f0
zdc4d5e867c70cd0c27a044e12952193f2d1234d018f9e45b472f050acc8f5431c4c88c2dcff910
zcb0cd378cc5a193046441b3329f663822465b74833b291f332547b86e0f030a61e606ee5d8df53
z0d6ff0337dccbc2cf4695c49517e743cd4c3a42e6820940909af76da4e404fe9bdf051b7ae7b97
zb9e5a62f355f9b4c3bfda768ddbee13adcbc79381dc86430b0a7f6e2dd5d65a806ea718e2381b4
zfcda3f838c6e17b061c537c79905aa54c8bb42633040e483c2d8fa52763a8a0d2a9b03c6973b1c
z14f3c5f01ea719b62066ebd6f84fd710b244491db26afda63999119173b102004525e81eaa8936
zae038a8f4bf59ac0c547803b0743283a9250b97c178bf2f9809b2a3ba1e4271880f89d840cbef3
za86fd374c38a6165da4e7e90ec51e440c821e78f604ad39c1814410149a813eb2b05c139942d9f
z31bf70516e92308d7c42a72314d0b44f7ec26b804b1ed867087fb056251e0e06b0c0f4974ab741
z07bd8beafa3818491eaea1b701c4f70410256f6a0cbf06676deb39f0ec6ee31d0b8e768e0fc651
z8478dc2fcb5cd62da85ba8b5341e8d8c1b6b34fccac60aedd3d3ea5a22dd651f565997f4b6429a
z62cebeff53d42b4bbac7cf10bac682d87fdc8229de89240bff7236c75c278ecd6361bb743e7249
z4cd76e46165b5563ce195843d6d82973efe7faaeb666faa014e1b064be775f93605ab47874cc19
z626e3e31278e68e353067fad32e5837e5adf1b4c23818ab8559ba69808c8f4dcc3e5b12a0c04df
zb2b862437a2ce3d112e78b49b568b9cc587bd54554c827034784c799931696e20ef3177963d123
ze8dcf5f8b6b75311904c21b4a6b3604364948c9f2183fd7bf8c3b8d56959f9e89da4d9426e4365
ze84b1d07bc484c48b8f223542f8feb2e2340c86c217204b4b54971bf46ca84100d707f9f568155
zda798a4c1d7654df96ee151a52ff3b452612f8f5df0a5f8e675ffddffa9f94b45d20527b17ca48
z6729aeeb15a57ba89d93a0cb5db6b5f872bb81980ebe83ba2e1ad52b6efcf6a7fda87d3e9454f2
z4d6ffba33767637b6dd7bbb206a137dd567d1e922f0afd3abae35337d846ecb352701505bb7ba2
z1ff89cbacc91fd24fc694accac09a238ba7aadc30c73aa7eec28ef802105975873cfaba76248b3
zd771180fceda9db863fc3296e3251898baf3a34d85e7d2d2674edd630dfcb09fe10fa74ab09789
z689c447e631ad693b9a6c4761a37208b78697f2dae8add5fb4bcc540ac75c988dc71b470ab26a6
z54d836c0d3be5f9f9345bd48bc4867f5f40eea7650fdc1a9bc61c1ef26209ca887df44e72b11a0
za9202ee09714f6ddf7f802faf5d26096a3551ba374f569f70c3ec5382cbac2beaa69e9c445e6f0
z774b642c652a23b1bfdd74c8e2d4f4e5653205a6d76972df36f59de8806868988e362db796098d
z8cd0dcdad0b8ee90682374d5114513426abf6e6147a063c26f9366e4005c8cc58fd1b34e9ea74e
z1845ea5cb9d5cbb028023e69ce564989735931ab673c33085457ba34fc16c7c96bf92310d245d3
za784932e86944e2cd72c708404432525c81d2718e85c8db28aef4586db4df192d17c48608cc45d
z3aec68d421fe57a430ba32bcfb079a7a71f57976ec192daa091f46aa80b7d3c3b714f632a90626
z72c51cf409dc38d932071d6215e9b3d326f39be1b45a3f5c43b3abb91dd96eb93aace922086e7b
z9bc70ac1b4a88e795148564b84fea8adcc7a76a38ac2ce80edcbbf4edc9e4f411bac5ab82126e3
z3f64d41a4fe7504dfa04a5a58a86d1d9615b55974a5f68ed7fa03e6cca191f8d6eb1252ca2779a
z51f4a4afb8b2fce0d50db6e8a2f26f409921c4ef59013c2adbf3514fc732deb38efcadc15d93b2
z1a92086d3e9f16735dd26bcb5a8dd275d3d1d5dbbe020fc6b4ba7f4531768690b40753488c854c
z62481c0b8f29ef377b2a0cd1f8ddcf5b289e897cca8d4d7e7323aedb0d25002a5eddbe5298824c
z3b04f5226a29e44a6937887c39c8343ba4af32d6d594f2b74f8a13475f29e086195527651d8bcf
z5ae12adfe2384c22749a5fb1b8701fb5ace9072ca239b3fbc3e3dd31aca5046bf163f55dc2bdb5
z7d04b30a18de48bec6f51dc97f009cb840cf84ae680d6532a531d71da97a6f9888554e654a22be
zbe8c3032459d2c94efaf00a13da8eed873e49e6d7c382ead40cca0270429514e2e4d6fd40bd3d6
z99eecd6f47df145b30b439cba3585090b4c0327483c2a71bff41d93f662a17731d21da8eb72c54
z804baaa14386662121285402d22f8526a8d39e162f5894855f772b7c438fdd2e0e95cf6398b0cb
z25e0f509a0f5698f865a2fb9dc7db579545503fa74afe9909868a15f29f6007f3ed602b6d67852
zd853dade1a922c364a23b0369deb2e437cc8fbc80e227d37218f241531d4773f588674e9a7b6f8
zd322feaafe8ac93fa3ecb54048771c163f64e4ebe6da4cfd88f3d0003f6cd20b6a224899a218ca
z58e301b836189ea90610a3751e9568b84e36ab1bbd7be2b9d25050d9fc95e96b6fd597cf590db5
z290395c4942d8be00ded17dfa5ad3132f9854daad995ff11acc6425e3516493c29fb06ac68f254
za86ba417f3e76271ff8cc03c86b094367f136496a15cc256ab9a078b68fb5c7af2c7c666152657
z6e2ba144ad75aadace48eb3e94554962685b2e6488d79f308db12a614a85a5ec3768ad6caa6259
z22b4c311fc8c5abaff19f4eb72e7ea523f81c3f051b452dba02813635a8cc1290c869f53af9267
z64fc3443bea8bed777bfeb403f75de0919cbb1b583390b55508bcd1ff0eff38a3f990617a45d2f
z6d51c744119a054c9d3f9986153b4cdf14914007ce0a5c006cf0ccab6466da5414fcdea00d3acd
z252c648f8a46984395fa53dea23175b51991dde4e4526022690886760f17789af2a0f269c058c2
z93cea3bdd4bd6e102a2ed986d8c6acd3f9bd117cec9063eef175cd99dfc06d97d376c76fdbe5da
z810a01d010b63cc3016f76d194c51c806e35630eb6a54f3bb4b0fffe36061559359165f2043477
z9bbbf53d26673ad1907a4b13d2cba4728a1c937152feb0beb34da03200e34e66d4f7890f72c76c
z579341943ff26636afd07a0b08cefe8530e9be48bbf82804a4aeb6b9f864a39db520ba51371d0d
z9e9614fbb3e01b4f37f52691016bdd76a241a623831da2badb543af3b7160eb56571a5e78170d4
ze9c140c6a35061afd04f987d53785e3938540d1d867181a04b476f00659acc5d05844e67fe00db
z867984eb6b3208e6afa800f3429103ad8a643317d3770332c6ce4b44350ae0a5e7644bf240caef
z07f4f362bf3c06d6e51f96d70c8d6508170b3bc4d1c375e9a1c8d0a4ae9ba1dc7ed153a080db4b
z4101775cf1bd4ffe9e493d467fd07d9312fdcbb878aaf89eca92f662bbb753d0673b7ecc468706
z76e205536c5d7b8bd1a57811032e4fbf02bab386abb13e697c26162e77f64e42bbbf9c78779a77
zacc148bd691660ccdf8c4638770caf9017f75312928793bc2d88a48967e6335ccb021fe492b40b
z2df43534c4059ac3a778ef366bcd0a4158b4ec8c97d29c5ce0479f666f798b5da20eedcbfcbc8f
zb5ed7b332f9c483c65f9ddf7ce5f0759e6bf2b74857bc08b02f678490f0dec078c6078cadc00cb
z26eaba606106f3e96bfb0b4b14f4fc95f6c53e631daf86d6398c1cfd03762d159912e7c70c56cb
ze2b9e7b3df956c27d9f88dd69bf0fa417def14c4c6d71eeb7462e020fcbd9ff12db6c25795a726
z70ec708523a63d3a1ca7a37bc46c2a73f6daaabc0e2ab1ad185ba3578470aa306194bb5ba127ca
z197638fab9c21b907c0a46d200b4f2c8e5bbc0b02cfb7927d43e22074459df571533a53012fccb
zc0c3d4cbbe23dab001a9376dffa17da1a50c160db1bb775a9c4ca325217d4ee560dd92ce968739
zf4a5bd9acbde3b5abb0eb79f4ff184f917c679a0fe0a3ec489127ee56b76267701ad2fb5e1fba8
z99b784616989eee8f64fd7029d741254752990d7e54333b9f23dbdbc59ee54a383a9e75ee1c271
zfd5cbdf15a7930a2ff9307a80cc4e3c0025218feb92d25a2c3626849d2128b98bc776878757838
zf075ec1cb0f85d89ec11947215f2d64ffa56c236bcc911e33621c3b7fc5e6d3c8688708127ced6
z27a5613c8dfe6cdae4a5106b6981bc2099e60e65c24319ac7624ca3b198085b04b1b452e7e9dce
zf1a1265917e85c4f2e4765cfcb5501e11f41d1363a3cc127321dbf38969049d076a3da88c52bf1
z1b4a5f41a0a2576706b535b555f50309ea579ae24aea257c62fa4c05b539acf8fdc9e8333bbad0
z91fc8681aa17a102ab3fe1dac954cc67106f5abf366ea98d644ec25ffaaa28189bec6e548c7837
z79faa090c6e7f018afbd19b80679932d3a12e16a42cee85fac79e23f8b163a5386a3a7bb017e45
z73674b38bc2664d6ca6a43b5e8de963c68de6a8b88f85d9d3c0b90e650444c9438bdbd3478e810
zb5ba5a5adad285225cc279350eb856f793dbbcc4a4b0a53e0c9eabfafc00a512e5d6c11672cba2
z0830f1e8f6c7ee67713e4948edfe7706ae31bdd239dadaa2ad02d1c13194a05163507fe962b743
zec5a8ad0ed20326984f9bb757e0d2fa679b79ea420fea103e620de880af512207383dd60d46d11
zffff390857e9b3afdfa5a997ea85be055611be3df40dbe59bb19b77c6c4e810601971be01e0d57
zdbecc75232075df203429e99a4c59cb1f1c35e3a6eb6466e2951e655b9f08f8d9a6df8f073dbdb
zb55a988050a25a689f02b419190fe44d4c78cbe6062f36e332325a6df36f7b828e2a361abae982
z76700e8d1aa880bab35789e4cb4c36667500bd1921331edcdedf5a5b0403e4d7accd1ea9157b23
z9e2b9ce47c074bf0fdd0a7dc8631fcbda8327ea3122bd349e6284bdf5929c317e9c5e53cf8e61c
z9200d0e2e785b620d5591430ae57864611d0b7264a165c970e866c1d513bc399b2580fd9bff3aa
zd4a3de27f513281a405c6c22275c9c00fc2f35decc938450e5c9226d7daeadf47bd8a73a4726c5
zdb7bda76c326e3835197f14f565ac7854ffc5bbc8f9343abf8f15bebf9305d85c9d0f01db411db
z78af2f72b0c0ae6653b255053b818b5ddd462b2eeab198271a885903216926dcaec17b44971a39
zf8a279c1329a7544237ff3d4eb70854356378815dab409f4089448938a41e8dd1f499967f2b856
zff1d49d35e26283a0fda7b6c90c2325c85c3197cddb87ed17fc16b303a3ea840f47e1afc53ddcf
z4756c7e94c4f7740b26fa426c23e562fbd254b6079d6631dd003dfed8f2c1665f7ad0131af9f37
z5b47226057f9cd530766a4ba8dd52a429d08e4b1f85527d41d98522066581beec1a3130f8af506
z4271be7066f2a2a1226569cd3a6ef06bd9c5d2167ff15d61b1b7eb5d1821a07d0c3dc6602575df
ze569990713aed43226ec04714c53c1e583d7a6e6ac549ccadf41d3abca915664e6131bd31bb63a
z31dbe2de594f15800afc5fb66fbf8f9f3422fc3527acbe54e9b62ca8d0b59b88499fddba7a5fe4
zf7360918cbb1706f3b1dfaaf6eb61a9181ac4783d6a0c3f91b7fae8f07d647c05176c826568e2f
z666b0e7b5bc2159b6d5bd038c836297394e0f7b95a7ed4a27f0e61c16e32945c6dff9582a6b737
zf19387878970263420308f7d61feea7492c7ceafc5f3ce02acb75e55aeb92026e4399a5fc4bf3a
z4823dd7cbdd53911364421e6398e821f9ec1157cd944d5ec586d130ce9188c234173c5326783e5
z24020da2869fa4da32b7b992cd85806993582a51e5c6b0ff0bb4c1c2368ceac5024b982e2c0db1
zbccebf26c3ae7682c1c2d80c0419f384781bfa23da25ed3b40bff94d49d54c723148e2e18d1099
zc40a02a32be6a0fab2bc429e3a3cb862825e05a726665f0c86e3654298db89a970ace124b61b83
z057c536717be8a08f10da89f98895dc34f758424e95f3f5c201bf0b41d72b947fe7e783f0ba3fa
z10df25302d076853477efd1d3313935a1f7849281b3678628f73aa519c15750d42fc3ef1e2bb9b
ze60d9cf3f31f5dd0ed6959bc636036b5e40b92e2a5413b7f10e0c6b21b9b5d2c0e2082f0aed1d5
z5c89eded66e589e36a3e4537c0a621d3d6115ebb88095f253d9f7d9b28cf9420312a0b6f5d2e8a
ze04b5ca935e7632830980218aacf6056f73341eb1db5617184512000f7b24b010439740c55ceda
z6896b819f9de75835291859214648e70f701db90897ac889d0a715be95bb75a2b413dccde51398
zc2a6dbc2482ca96ae321555f05c8e4839047dd3b75c67d40a5f823b193ff9d5f99bc12a3ca3c5f
z46972cffffd0c1a2440dbde2bc020fe8d2b561b84d94a63906831cf2d1dfd066e9dcffb097ada2
z3857a259266731997a3ea2325cfc621f31fcd6777cd3f203c14baef4fe0487d1a51b971b2b1b10
zcd9a81f804b66bd14575fb9bbf6a2cd14128477f8018965c525d243d5fd3ac77f1139af001b72a
z9c78ccb71e0d9347af5dbdbb604770e2927a24a1ea43bd87064bcf505c690cd498fc80f0d988ae
zd23d178cbe95ac4bedd5247968e5a59e17882fe7a973f9cf0ec1bf379f5e58153a0465dd9036ef
ze6646f399130256cf66dcb9e56d090ba5b09dea66fc502eb08f88b773aa6eb6da27ab966bdcd3a
z770d9009e3faf7afbf951b03304b56f6178752df82922c14090c191ddbc89de53f24a593d407be
z229f3df4d174c0513328dfc2575865d21917fa3f0218346569e6920df852e5cd773559190cb961
zf31873950851aa13568f69cdd249e4d8ed2cf15fc0f8f1e4c173593e107597cc085fe29cc6d83d
z1600457d40bb408f9d0ada5eb21a303cbdc5e62b77fe8be6938ad71d81811098303b29e741e122
zb69ea1eca0fbcc77385b82a90e26a8e322fd970bcd53be7c5d66a9ea5adf0ea2f2954b9abf0e90
za3bf10afdbd3f328535e5490f50b14fe7ab84d39da8c60ea1f4a690ed758650644590b9b10ade8
z7204b5d5b4647230e2dfca6bd404a9c2828a0f692d6fe26dab8555791b3798afbea82427c44f7a
z29620106d80ccead611ea94b4127bec4e59818d9a295f8b39c9f54aa00c125d05faffa748a3646
z9f708d87fa19d1680261c17263fbfc2dfa22e1db0046f7cfe8f4b0fc7cf167d886c6635b3e9cd2
z9da64d42cb4e2f307c8647dcb7c263bfac7eeed8d72157b72bccf18a13efe8663c50af70e2c5f8
z81ab1849148e724e5550aaf4a99dbc98c0a48a018b18c50363799597bd622b48a1bcd1936899ca
z7e95b69f1dc7d620f60e64088f0a49412cd2722e3b7edaebff099f8219a1a456a9b5e8f3097533
zd5ad82c5fde8fc918e60455eb81a0a691f979d33856176146d1c8d3053bca1e0f785c4abb40bc4
z601246d6630d4d1bd52c9a8f20e35ee20616b0dafb859fc7842ed4422e096b49d4387fa6aed20e
z87a266133159efa11e66cec0665471bca1d723e5c0fac07b30dcf317b1553862e4b2582013a9d1
z904ce7aada30bf47027615c26fe5e94faf20e16dbdf1cb6dbc2d842bd3fca185d1ca0efe8a7dd9
z7d84ef9a68248ae92685461c102345f08041a7e337b959be4b911d37bc8aaf295c007d313c2e98
zbeef7ffb2a21ec005b378ea65ee8144fc5aaf996d289a259feb4a35ebcb26afc5da12067ee7e0c
z046c4abd9678ea78c9e2811e3247779045d4fd18fee6ac795b08b4ff72b779ac8a29a6e7de8236
z8226c1a9a035197d4edbca1b78d6e4de7b1fd62e24f4ceee73e88fa0db793ef2822ce52d7d735b
z1902a17dda4d534c5e9bf1e35af60b7d95a39746871a8be0e7f4c8b3a698dbb0b1a925b770314a
z55e03a3ccf311a3001c18a34a50cd56e02c09608034ae23b82ab96fd2273ce7b0ef0347e2f63bf
z9e26a89ffaaeb2b31fe8e8178ca74480d161773bea01f6997b5bb1f2cf339d5a2f8563bdfa2bdb
zd4e34a209dc1e517807ffca40a85f22a396b68675e73ae695fbd29ec8aed83b67a3a35b1779b07
zb52b5d0229ccaa48123cb4a85fbefd3527a913d2c9e74278c023bb637597a9cbedc299ecd6293d
z03a66de51b4eed0e859bc69ed088bfdd01c70a1a8cba02a006e5aee99b5644f544d47917aa6092
za4d612b9c7be0462f9b6524d218551fa45a329f4551944a4cd3903ba4968f29532cf89ac5c614a
zb69ded990388e3abdf42016bfb1e83259db91c73dc145b28ca12ab194f382601252c343191b551
zcbeb66551010e547b4d325428a8e0bcdd056f1f2ec7d2c4c952981a561c1f85852d1e5662250b8
z4e703c7f3ff694421068673fa449469112db87ba53042b4a9818d2efb5ae144084bd87aa663d75
zf4514c0d973263e21b9bcdf5fc0c0ae232fadc1732d9675700079e134af94473bddcd97646ce29
z2f30d38928ba6cd8d6c4759e02ae383bf2d023801578fcaf302dd5b0c69f4906c6e37cb1f9c15d
z6a79461d2e35c2e0c30f86d9986437cef894c5fe122486705aca12fef48404ebdfeb6b1acab088
z1b5cba60dc819d10ca8ed58e2a17466d748e1644611f301550d4d325f1dd16f38ad8d706967ae9
z31d2738ca09ef02240ed8debb0f0289074170988e8a1bf3be6a02a70f378913f1124ad2fc6181c
z919ebfc28b4604e9223bc9005359566ba86a26627da755a6884596c1056311bff9205a7d7843ac
ze66167ff8ad6c3f4250287a8768f289352c7b58e4d4dcf1fa79caf9b70256c75319be8194a01bf
zc5bd1c6c666461acf0aaa0cb053e295338bcb4280f3b2917fdb9a0f0a85724334cfc3cd26e0a05
ze95795b377210da9c4e8dcf0041845893fa2b1ab4c64091d411ef1676c1f78491886d01a97106c
z0c1a2b5127de352815cc12b106f086bf6b9d25e36df798532487d4780ae476387e5e7d02c79b35
z7c23a1213b7eebbd4856d4da096ecf05f736aa9a33039d71b3611e2fc993689931c999a4b5a472
z902bb402f1cb4e0eb564cc4b6445ee8aa0e5021fadf8f33011a81fd5b76e3a5f9fd87cdddb8115
z7eebd96859a57c413836d915ca86a3f75c6faf22394d716b57ab1c18ebb7fb47de52103acd0267
z1e2d3f280654fe6f83068d3d61fd7657bb234d1c25d0d7621c03fda42b22e039801f1ed25e3c80
z9918c250d0b14b621bd74303937720208f4188f98a97342ba1bc0e18b716ba2713c644e207ac1d
zc8bc6cc23c06e2b767aa3d3cd89d87cf797db0822ad4fca98efe353282444fd533017506718033
z671ef5b2190657a633c29f9e2c04fe8d06825ba8d535d536f9cea1fea7455486d71576675cc8e5
z5560749ca71b19b25b62eed93feccb3c504cb3089fd39136fb7afc361a481c6e7380267dec42f4
z5a9ee2a411bf9307d5fb2c33faaaafa0bb6860da8ee0ca8762a28882ec78557a9d09333f004e5b
z80cdc2b3357fe721735fb08b12d4a51e3c07e270b06363a2d7ec1c1c9f7a9a71b21ae52ad7d56a
ze2d21c5a4dcd7d13190e51dab8d9749be7e68e5d372486440bd7e3e9b789efd37fec8eb8ae3e66
z7b3b496dc7f13d8026e495613fe88f4e9bbeaa33a5f2e49620c1ae0653449dab0bb1472debe6f8
z6b93ef94e6f2670f575cb294fe6f336d51a3bbf9574a3f4fc25c15c389249634f271b97c517516
zdaf4d2ece90589010294dbec3342e41faf51e9ace26622643ff50d740499ce9b59fd168608f2f9
zf17e560085b7d7c45e75b74c913dd39834322869646d6482bbaba767d7042ecb5f85ffaa3bd1ad
z1d38e5a56bb2fb4d9d4ede12e76ec00c4d3875372e81e14b6379ecb5dfe9a3cab1de76c8b17931
zab8d4e66ce904f99ffe8cf5b46c4ea2dd7fc8133a1d2bf02cd3ea29748dcb7bf2bafe960787d87
zecfeceb72dc50a57a527dbe47603b4a954ae82192e040c9020e512e6852e39a0bf59e4c80047ec
z19be1095df4fc34cab30190a04d9195907ba8f8cdf2f88a5df4ab7b440f8cb5af6eafddd5a6e77
z7699ab9785475ee9f2e36636a09e63c1653a61d4155fe1cd09ba7d111b07469a91b3efc200e5c9
z12d614704396ca5d036fe9f96b4b2e939b71903b2ad9f527dc36a4ec759bba1f62999de9d27a72
z415aa620d528bafb630442ad0c5af7f1e5a83f51e4c2ca72ccf09b3e91db10a8940873adbc198c
zf8dc41ae626c03c59cbb5dc6a85def1d8c19f6010bff2643e8512faadc4ef82328bd044d9c20de
z8204fad4458c585e8f38e19784f7187189289933e5e642c3e10943beab001b557900570bb8282e
z29ba47199abb3936474cd6937d9e3faa09f28021678aac0c722e873213ed84e6496afbe8c93e05
z6fac71ea06d72405db3f01e1134f6bd6c36a6b7637768638e26a8425faaa1227abd1817e733a18
z1aae2f3ea65453bd51c5451c06cf44acd9121a0fd246c10017a9b76a8d53ab8ed4bb38f7ff1ffb
z057f287f1e2fcb5fec3b47750abe496686d22ed6b945ef8ecf54501b711e51ddaa623c3a01511a
zc30a865c787c635f321cccde84ff28513d0f02cf3a629ec2542f7aebea31f562de42892510a177
zb4b475e02715472e619557945c4bd9ae75302e27f8760880f95e7866843b9904746ff2b801c1b8
z02c63d3404a86e6a0c9d657fbcf024886b6777da0d4ae0d30aa999052cd716e40e5d8a65ec2582
z44b76cee37e10f40bf5f75d010d110862ca568420176e33344ea9a1130b38a37ce0573ea423f72
z031f2d2da8930569bafb0ce661ea64a749a20e804fdcdcbb1139879579477a1970522c03740f17
z4d9d1eab7aaf15f2f1357d263aa8480353999ad13f6281b0e2ef06b5a7cb40dae365664b4b8bf3
z95849aa57d38bdff1df55d3056cc3b917234b04052726c6118fe8a6359f8d9962973bc3229bdda
z876f7b51b85d6a4784605fadddf87e898b9e52056deab1e3af4b5b3e1a5ef31ea6dd839344ea11
z0db8f55be5d3be14c72a5b03ff6fc044e9a866dbdd8fead0bceb65737b9608ef3aec9c4f45df9d
z791b0c7aa9db03019841a50337d3dd657404fdebe12d789c2941878e7e7b5b573b1b53707f6efd
zb46da63009f23f7d4e6bfcb9e4819a2b80a4fa17e3d8a699ed24120fb60a45d3aa98901053400b
z347981e0b790cb4d4418ba9cb91e6127d1fee9070882ac14d609b69e794d188cd41b42bed13892
zf35b7ae3b75960f15155916267d80f940f0d8439fc5e775c16f1c6bba920d1f03d00f205fceb62
z1f1e0b23d8172dfbffe2d854b771d8693a3639f82ac2c27d06ba841dc7d40a7b09e824adb9dd30
z1923f9545023efff7aefdcf4b1def735c81f822a46daaca168f02f5f9ad6abb412a0663e807be0
zea4dd368c7c30226d30077927696b7cd947e710994ced92b575a95521d679f987e3d5c4272295f
z056c515da80c92fe941403dfef5890997f7a0f8ccaaea450d2518aa6b99bb1adbe53849cc07697
zd9e57614b5a0b213efd0d57984b0a54d5e298f26cd951708ba14c6205236a44a315057b3926f5f
z4282e2910979478ad411ac7bbf293beb74c9c3b26cae8116c00e3bdf31ff21f1d587572bec3582
zbf563f615cd028566c0feea3317a8276a3221416b12a8dc397adf6b0ca6d67822628b0c5366dd2
z43d8d1315af12f5d1d5df80a43af55ffb94fe3b222da01d4fc28858fb767f315c314fb4530c0a6
zab9355fbddc2857afecd03e8a08065202cb0c62608f713b123c1e30d043d76f044afd6c7cb0928
z68629bd7547c55bfac09c2e4391bd1fbdbc4a7f7d5ad8e19ba8f6d9956c0b462ff906bf02f61e3
z00575705089067efce6bc1ba16d2effe3f1a2c566192b574b8d059657c93a9715a76f11cecdd26
z371d15a4f48321938e2615ff60bc5acf871ad33b8ceca3b877bc81dcda896cfcc78316150394c7
z83c2056104240fe37a4553019ae34f52c750e7927823ccb2867cc6b349e88ff96e4e8623db2a61
z36b1a6c3d95f31797ef69210b468600dadbd0a83a755307731ebc51776f60337946120ea3d2113
z9bf4858169c059867e5469e1cc22c1a629fa8b06c14904f0f7d701443ec067acad2d39fc77773b
zf9019ae950742045178ff90bcb65ab4affc797794cda236aecf343b1e74e45337c41cb3cc9f86c
ze5f484f92655c52b43faecdfba18d7c5883d3c0d82969ae847c8d9e5725de1deef96c1bf7e38f4
z9863ace326aff8960ceeaadc424976114b47b642d3c6a591327e2209f16edc8caed88fe94c749a
z416f901ac056df48227e193832fce66699b04746880a6f61f9021aff02ad98c2e5bcad12dd35fc
zd7d99cc5d9646ee0eef776832be1b243e0baaad03d3187b95b7ba0055ea9f37cc71f64b330657b
z2ddce547f50e1be0c2f8ff7a22c53017be58ce811c2dd6fec27c219ce85c06cefb2057d00a0b0b
zc5ed82ba46de3ea711e5decfb0d79335aa8db15bd006dd930ea35f0df5b41585f699b8387b8d4a
z1eb93e623c50afc7a0f23245fcdeccc3fbe02cb7e24add4ee040719d500db04188ed132f88ae7f
z5a6034a14c423ce0484b28a08a89f39be1ed0d436c5ded117a8be51b89ed030d942d5771ab42b0
z354c4d2084191324deade330ce1b0cf741b0652eade05c01d60c6050ab029c660ef76ce57af093
zb7f0d970c098c6cd219db35c010f2d5811f63759bff9737505e351d7840015557bffa8913e149e
zd89188464df1bad796164685d7a21fff37a9c9e82b5860928f8886e5c68ef48c631c1bddc08465
z043a7f8cdbe4d26d92145b9916706bddae28c3459aba92bb5637b2e1654c4e6c07c4138941ea53
zf79aac65d5e5ee6bfa0f8f6ba41c99d4330fec69ce5e67f603dddb5ad0d8150847d4e9159a1027
zdd5ccd8fdb5acead9b44e3139a8d155f43211c9eb712a465dda9c84ecfe47224a1408c33e7e853
zfc9d171ec2b59752f935918bd9ad05e7a893eaeed5350be8bd59c9a7ca6f0d0a7c2ecf85f70372
zef5264274699cf5859e5886d8c3ff33cdfcf9fda2d9cf6794aaa093429215c67a9cc77e2187941
zc0dd26d3a2c6ca19384aba52885dbc524dbe82b8346cc60a9b129274126a8d42f232f15c6ffd19
zf96363ce3a3e3630949b9b0c55d42bba376f46c76ba9441f3428cf0cfffc410f78355f2998a7d8
z5a007595bb605df3826d4ea3a69ccd69b88155ec3322e4e3ca5e3b9c223326d9f1a5381fbdc4ab
z1b87b6cc51b98674611bfe917c286a037372e78a48327111cddd5f1ddbd82b186c07fabac408b5
z3dd82f834439138dce1b2b2d0a21c067e99ed642755759f21e9c6a6bfc906e0c5c4bdde4737dbe
za650a9e5e154223313121e2561635f1c2dff57675d3b97c9d5a308ab6a64790c9e236d43d42acc
z1b244d29637e7fbd58b061e0103ff8b7044a0829e65e00735bb7ebc6b72186435e6d2d6c13e7e5
zb1d0c475a0e479f476f6b1ebbf3f8ea43d146d0d2f9a933f05f32eda3e1ad2b4e00c3200b5aeeb
z27b69dd49dafa2eb8ec24f2d2c8e0271174ee615302e8dc1c3f2a726bdd3d9210e1d4217bdf4b8
z9485d34103061859920fc64b0bff5b1161aa4deb3c8a25afd8f4452b28ea2a9b2d690d28e4a36d
z68174965f742d4f21250e48a9e24602369e12bb2782d70adb702db3e489310a4cb62c71a4b1dc9
z9caa4b7dcc9133bc3d43dce36ecc0582135537ad49f36b0bc1dd63e27e3d8ba71a57b27b120fd4
zcc2b83e69c60fa9ed699f1ec94c0c17e5cfafc4f3d63d68eb206d52d9a5e8d6115e6ce4a9783fb
ze9e1dbb5ff7a76decb58ce57124e6fbd1fcc5093f25a8b93cb70b4a4dc8cf9782428d3af8cf5bb
zd7efbc1b2096ae1b519b2692f8242c5f21f7aa161f5a053cdab8827485760edd7ca7413930e428
z27df060bb8737ca875ef81305fcb4f299e3c0f57e00c651f8fcef7f771d9178894404a9ed36772
z0e81c0c91a054d0e29b1407f5b419b8e9a15d911fa2b33a4499482addbe165ebf80a8e6a132728
ze689bcfa6d9950636d5817dc03ca01deddd621a76157f18a3fa075087289abdd3360dc48b1c7c8
zbf147665d335982549bab7663ae2442e55ab3e59f19d1d405d54396fb307d55db8f8ced3dd3261
z58983e10c68fc04ff1d2536b3d7f6b3010e8838f7444551bf06d7620efeb26eaaf207f2d9b92d6
z282025f02b17d7b2a2624f1e150365368761b5a7cb988fb468e8650beaef3136ad34f5d9daf44b
z0c81827eddecbf20f73bf5938c8c579a8ac9914471d5f9873d056fe091b5a17596cf4e933301cb
zd457a159c70c1573ace06463f5520b621bcc5c0df0b71b2c068daa1ff09b5b42a8d6dc63d2aacd
z3f0896555c937df16c8746d38ff92cab782338c48c76c4ba270c2d628d60419b1cf5e789f8d8a8
z5cbd852302b9c11428c7204a4fb0da6919fa1581acc725c4be5da0ee2c5a581eb20246b6fb0e95
z65448e777b15a61da0d5b1205f9cc35952d1e7038388bb2421e86212dd00e2135109a5c6d0554b
z846574c39521dab6d922d4ad24cc1ad61ccf55745c547e65dc2469f244ef739e088d8ca06bef87
zd5c5423cf75c0517e4b200ad2dd681fa9591ccf7b6f8889a47afcf65767e18fd319613f0f0a6c3
z2f27c1b98b8dfa0d4a090b6a9282318a0033517c44320049ce7fa14275416fda5393b77e82bfaa
z2ddc8f15e74b751984e4df30bb5b3005f01f82b9fe17c33f1d95d17777c5f1b40c12500efccd2e
z06343b1a020c6eb048f52ed01aa7c63c59fc16c281267a40ee6abc39999aa8a09e80cb737707d9
z20708dd389322a98d7a32d9e47d18f7562b904e401131d1e5d6431c91a4ef91a36de14a02a2357
z7f66f86a83c6a9ab39de2dedf7f2eea4dcbe296c96c5c64b534f09636c6ae9de5bc87362eafb72
z41dad33f93b55f26ec2266b575cf3eaeafd77a86b7ab5da4752899e6b14a1802f9a5a0439a5059
z7b760045a190dbb618ce546690e845230aa017b5f7d92652fb745b6f997761f55530623a978741
zf45cca9f0fed2afedf90302a02addf8ed3bf2b2b083c686c75fbb7f4df027b7f652bd436e3596c
zf11c2bff154d29010f914e0808ca04ebd2954465dad9b1a0f088cab5a4a3b767d138634348ab58
zef9417f01064d9c9d4c75fbdd0fd89dc548acb6b3b80f0081cf555989299b5abea187b96ad9b20
zdc6cb69df6e34a1e66be36ab0d9b91d41b2e21499271e7f30907530569072881b746ef43b0ce1b
zdb1b02b615f6b7aecd1ec6addf439cab5f3edc61ea8158c6b2e1066a87c51027696dd44395ebbb
zb74faa5ed93397cbf60eb0115b483adc9b4c916fd05e879b00b6616ba38c27e7591438d9e90eeb
z6d1f8b2cb4aa17df5e573805d9a8736ff5b80224cfb5d0b204370ae17dd69dd325122e8c58fd89
z70fbfad3a0aa408e5f087dc50612822054f977d884aa9f722afddcab43dde38aa17915fe7583bb
z1cb3784a90b29f16030c9de56bbf1f7b2e800e56606f328480dd4dad28d757459c8c4b8f578a66
z0cd2feba0e2f3b2c677f8bad395d65838b6a13f255bff62dd104765acba37dd30c37caa8e21a9e
zfbc9d67d9e154053eded7058443c9db6a2d7b20f476d0a2f32d0fe53e08e164d466e544fac1e77
z31c193d94d3bb1768c30205709f36fd7160643056f869529bbbe062307d558c5952a1250a20deb
z65b09ecae26b7b2682fa2866fcad93eeb198b15de02da97bf284eaf5e41f8d62465863db3ca93a
z5dd6813bdbf6eab331139ef2e839ae4b45a3ca6d633870f61ee946bff7630eb8d3977b548e648e
z020ec6e107349e1f74fe9c1a9d62c84534abe72dbd6c3cbffda4037f64415a5d10be5f91104916
z0f5f406dca4ad971e6e4b0390ace376424f35eff8c5a3db45effbfcb74df4142d1c9a2c1aea4d5
zc7dd7d0dfdeaf15ed295c1ebcb636299feb625bf9f44c844e98a6a9b0056a8efc1596bf73ec24d
z493d1936f94fcae03513d12241afb0d04413158bfe67962a7addccb052e27e3fa22cb452bf7abf
z9b66780840249c4122078785a01ce4cf9e683e1b42082f23229b3d04dbff76a7f780c3d54b680f
z4e33832a49ec048144b90bb790ced6c1528370bd81a05b000e49affcc5484674dfe91e202a614e
zca71f99d37e5963e1ba755629c682ea893612a2d36003ba0ef571067eba867fe8d4cae491aa7de
z066a5ceac76490cad1198637e5ab058da310b4d09683f6835a595159d54181a8717e01b223f459
zbdfd07a77597642f1d04397b42d6f52f85f80f464137f4717d83f3060a35cd5629be261bfe72b9
z5d8e6a053a51aa1ff1b6e30005f875b912aa4057b60b9b031e3b66421a1df4d4bc9295aee01f36
z757f69e19ad719288f620a2d079389e97e1ec0eca816ed06b466a7e0cd5d94504d1ef0d2e9b4f2
zd92e100faa94b57215a56db3b2f8e68ad28d995caa3bec06e1f4bda72b46475c75b6a792642712
z83b77772555229df4ef0688d45f7e6267982961d2589457bb9c96c5b159ec7df987b850253ed0c
z80db9f36e13a0bc6dcf1a97a931ed7287c07a95ee0db2b085a4f66e2aa42a582d3527e7fd208b5
ze64c18593b3941c65e7e5cf0cda5b3d7d69140ab1796f2f0b99c6b430d1a23f8dce713976ac97a
zff0d880c07baf43a5ccd77a0a3d84587e8d6817b7625a0315750973e896ba0936153f64b43d325
z0690aab82d1a0810e5865b8012db542e49b3b030ae41596e6fcf2dd30f22e928eb4f6c19f1010d
zede9d611cf807b0e63592c3908e114a8ea861a6e84a2ba56a9550bc6f73a991d97729f8754f1bd
zc82c47d52f5341a29f51eed76bcacb06716058174716fe2879d156f55a8b87714a0fffbfb0aca9
za23add234d07f3df1f3a4525e50b530baff3c1d3bc4d212f20c499c476d9534a33f746524e8305
zfa290ee07e75ddbacbe70f7543002698c28eba900c7d7bebb2de0044f58beafd70328ffe7efa63
z53aa666e885ed73cd07fa6acee36b1fbca79405407e01e92d605bbf6fb6ec34e5ef279ac2957b8
z71176f88fcdda8004e49b18cf2951314fee96c8a5b14d3d03b517fdbb794e885dc185cbde3229d
z19f9b1803c844d75dedb9a33d373c9070fc6713145b728be7961e224465a6f2d7396c06922dabb
z73d3b5009f3ea721ed5a23861a9dce52fe9a3c679d3bded831c999457989aa2837d831fc40c9c0
z6c9d52320ce00c1984d3471ae7de340836fe339c19398e4b6d932be46e9aacd0f2c37b33bbf903
za479b915a96f137b5192c6c93b4ded6ad4ea88995fd5ded8232d2bd540a106ae2e0af104fcb79c
zf22398b98cf2af4e2900cb8a9fc0d9341943e4fbfe24a9b5de507aa4f68a8d3369fe40a8335e31
zef0bebdf3c95f041e02ece3ed04933441de6ac7f0a37f8e69ef9d099c149ffab4e050f1ca680b1
zd9f11cdd9995338b3b4020c335cbe666cf297ae22447f9565be1998fd9bb6572757109e15e40e8
zc4a6ee8d97eba5a64f48b2cf0e5f139274760fbea4a6369302fd4b95ed281ea7fda04c6d3f6447
z15d91b1417e628ed006080578486d24e284d3ad2c58ee88842c1c054966f6493b1bd4783a695e0
zcb420693b26858144bfa77148610aeaa788d8d40b2d7c1a954d22d70adc6fc2401a876698c62f2
z8694489a3b734a33e0bbed8b1bf76b821a69def45b983ff9f81dd293240f8e3d8fc892796c6731
z7b4e758387f612a3f12488680432a87a63f55ca2ac675430db989ef1c9ed860efd9703ffe00b45
z1553a9a00ee812e4c29a9f6df4826e3f9caa9da5f8b16d986302fcf4d3785e7f8d4292087f6b46
zbf38d213712d31083bf6541e5935ec04f7efe2f0744ecbe2df941ada6aa8bec743e5953d35bfa4
z1f0149d7ee470f38319d28e65ed01ec54e98756b6a5b0cc2a0da4daa697a7cb0102baa419586a0
z25fdbec51c20940497b0def03628bd2faf548c8a98792f8a07930e10f095d1e17adc8e5575c270
ze475fb87431d838aeee8dfb0740756daa1873eac54ec9d9685e6db429ca8bb5debd474a04fb161
z7f7441c5f452e06ab018cd11342d871dac15a1bb8bd49a6f51ba7228afbf1f37988a0897ce3ef3
z0248afbc0cd2aab05940c05a0654de2c55605796cdb0577973d9022365bb7c87c7062ca9271836
z8281e292bc93c0a92e682059566d91a44788468a73aa3e607b48bb7e15bf99bf098304eb913204
zb9da61ad66e573605debdb96256b2693d9c3710b08ea715fe51377c56cc08c29b3b0a8a09a20cf
z7baffa18be401cc92e6e62e02e8d6ad8b6d07a693db025078de4374ed7ded1b6048b1831bad22a
z27658d4653e2df0e4f74295aed6c5d5bc7d7d60176051a5eb1c2f9056ff25591bef247550ded70
z9f9c30515ee13081ab09c71a02a00e538b829c666b1b1f989e417c4eb57aa2ff76624c3d7f0fa0
z4d75d851515775eadc5552c89fc695abadfdc611de75c843bd65dff229e5987c551973c88a04ff
z2d6f7990384c71fba8791194f0882f830e257a66e55febdbc7e7c554719ed698ba2436bf3f7447
z790061dfb1ff6db5ace49e85f7711e05a86e32d9c677310b317459aff703c0fbed7f5dc2aef047
z61ddea8e986c4b1ea4ef908d4909a994c184bb449dab996cd4713acba9fabdb9c68a4d93efc9e3
z09f6f3be051b5457e41fd574512e768d2244853935c43d654921ee9d28fc9eb00a13c5e6df00d5
z66358a9bcea420917b730dcc598ec9e7024ebe006463591f9b8d74d26cf0a1ea227bec5af43991
zbffb6d0c403e62bb668a324a10fe19ce7a466c47a9e45874cc2dcbe257d4a3046cb207ac0cc4d6
z718a2388360b4809ac24c145d3740843ecd44ed77fae8114ed8e2803199479dc271421dfc78c0d
z4d19751223514a581f0c97be2db9c6507ee13bef90b8ae6ab55c8a6669bf3e35ff7a2e942d7c13
zbff04f22889bbe8c64b31e45d474025b28c9dc54d2e483a7bb64dde09355f097fd9b2d21915e6a
zefa1f406c8056a0eff74bb861f4ab518e7d27918f15a0c9bd3e068d3c442e25f1b37d3fdd520d3
zd2fdd720012b739e74fb23e10a6229261e4bb07210d8977b20e0e1eaf9275bc13036dd20159a58
z1a9d2bb8d8f167af0362137306a761e2b49f7e7bac832ab7b1733ba5420da97b9fe58799d71f68
z41c417383cccfdcce3b302732ac96c904100910c74f72642572162003d0c3eb19c1984a84120a7
z2347274b52207b7cb10e80d0d93a63cf95be04099cfa9f9092f8c918ef77d59b88691c8ffe3ffd
z709a39f21e5e5f6937e4f05676221af06cc2a4d08652a0cb5a2e0db200fab643f0e782ee30f317
z39563491dad535243e2c7774ab77c9e0e383ad66040215ccac8e02ae7660645194bb60d6da9cda
zb9da44591fffeec36e103ba4e0f2a958095667df86456752458d27a6fc03df14375a5ee87abc14
z5f68b92a820aa96995da530e83c7ac17d9de321d6c2857e1c44775bb4f6df0fddd4792fb6d1b5a
z5992fe9d4086243319eeff8405144c0d1b158b104e57c66cca0dbdfd35225a15317dcfc5d69c96
z5bf97f7d0dbda0559cf6942de60ff30d6c80f073a711425a9e696cef6cf6960b223f7f8002102a
ze19e4fc4359b31eb85aee54088f1d15039d73e6e56c3ca45596173f8f608f6f4a182280ce02180
zb057893de55170d042226ee255c86063298487b477de6b229b9df5688a9b027e92dafa4d837729
z14edd2b892810b23455c2bb8b42ef89e1cbaa47b4a9f513b54afbfdfde70411a442c5f49f889d0
z51d00ab3a038cac8bf871596056cb2f59feb52375ce43d48298180689f47e985a28bb04cd0c4bd
zc18ab424cf90acf894a86ccfb121b0f2c7db61797efee69d4232fad02820ed948f81026d16bbc8
z8e6a9dca5d46de78d299ede6b42c17703913c186be7ecd6ab311f00a57adae9c26bdc2af58b97c
z4ff680b138fb884cb0165da8379808246170033970a66ab7207f733397be043172535834106ad8
z8867081548adc99f1ba005b8a76d6039c084ab515909975f3dbd6fbe8037cdd757860f4d867a44
z33889f338a5e2c02a41825ed66929ce59b6db4af79e9ab0870ad719d5456caaf25e68457574da7
ze29cd46a191e9eebae91625b3447d1cac9231b9916dacde6a691b865d3b7bebd5fa76628e35b67
zecda4ebfd89a8739dd12466b6872c1fe5ebeb7523cb2021c9bcbeb34ba8b26c2d85bffb8d917f6
zaabb2eb0ce065a40c9122eaaffa9557be520b804df91aaa07fdf1bfc9ac1a94cc51bc82ee1cf70
zb32e5f5de394a981b9c64197650082ab9f13a39be6c2d94a21119a4e8e09410247cb344afdc99f
z8c7539f0759ceea122f528b3f502aadda0c31513e957e26936a64ec4437056d431bcfdaef4192f
zef2084658d114a3df0f0e728ac54565b6e5cfedd6359cf4b62afea3a36ef5a0c2b9fd5a99384de
z3680e8e2347e65d9b7d4140f277720cdfc83b1bf1c79d93057600e5e9fd40db3c54173ec68a08d
z8f025e21235607f86e40a666071edbe82f665a67ca3dcec075493a1e04d60795948e0267843299
z0eb988678ed241b1a5344d7ec54e5fd244547740a01476e5c65ab5e415a0adde2971fa97d29749
z52bf17f03b4337d389e1c726a82e18a5238ca872e1fa0bf4dcb6d86cc2958a82b749f1ca7e4045
z9d6ebd23117fcd4fb7f4a21730f01730f2fd95c1da79bedbe4c6d86d1846eb000c73b4f445664b
z206cd3b40743b9fa0176649c94b8e96ebdec8e6ec52937a2f2c7386ac485de16a2267c826ca11c
z4a7046bb2ddb3c7ea74266998b651be81cd64be968a8f76fc974e5956c22334ad6b6c894bac05d
z507b757735443dd6ae0581cbfee5e252ca4496f0402f328a83c9992d80b4cd41bf369171209079
z7fc4ecd034a73807789c9426d67427eccb3b129daa00670c91232fff8ce5379d827d64cff67593
zef5e9a9830f6aa5d5317fa104a391f01753da204e9d6b82d822b22fe89ecdd67cb3a072761c000
z2a0da0e859d5d8d66313f2a8075bd4c2062e400a0dcbf1c0d7615c57a1eecd1e5ab97fe8f9349d
z80495136125f2996840ed0d137b5396c1431e6679c16f1f91e2401af648ef598cb835086f0206f
z71249c10ed9cd2ef7205c40507b6bd503e58f81ec826744e2e401471be2069dd1510efb95c9ac6
z7cd3b05be74b0dd140c32bd565bfd3263f8a82abf11a15fa20f105ac62dd3945ea640ff9371582
zfe1b7b2efaa7496b1e6dde5eda2694869cb9fb7caa877d8ddc8f71e778bb7fe39a9e24685404f1
zf96b69a13eeea428e17fc2d558fa17516ffe64ffbb6a9434324dc4967cf1036f269d4a8f5332bc
za4005604dc1a92e584167f65ee8172e938ee048340194f174eaf24a369cc74fedf2d80136d0368
ze3ec877aaf32d4bee865226e40f711426a7a9fe4dd66f72456d79e07de80a7002504a878834cda
z5fed91155255f6f002cfae5d376e2181c5ef1e3733f162ed798ccc5322486b4210fa8f458dd0f6
za9cc37a2305d7940de5237f715e223a3ba857dc8acbb46c5a4f16f2452a403681a9e9422277b0f
z84845cb1747dfc9ccf05e90a4a66d27441e05bfbb53c27e36ab276bfec93e2965b80de5c9b57f0
z6819d45d3bab0518ce0626e9c97f4334b3d5052878ed627a7fff2acd598101d597632c8276b443
z13dd86a4d5bf5ab2d7b4a7509dbd0884fc6beb4377fcbae695c99c66bc2c17798641845c14e916
z2c17e40ee26eeab2398c9dcc9e944f81e57a38726c2cf7d713a64d25d8ebdb1175d6479655e9f3
z00b4d6bfab6dcef20cf9b2577d89291bbdce5bb2e014d760e616b37ba597d34ad21436ab0e65f1
z6c3c09c4e2bfdb0cadc7abcce08cc4b68536a56a7ba1143a7ec6bb94a07d4afbd6445e8ef8268c
z7a93bc84d94342013eb9cada7b2f3649c17c64455b0438c55ce720f2411759c455b58cdfe49c63
zad155c975aaaab8a08a03b81efaf41c3af288ac0808acd8910d4e27d20a651c8e6237a7f779199
z8c9c7809481baf3bf675935b11b6fc485b7e854a9bf62c386cb2dcda268cf086471eb4e35a8ca2
zee9505ad8e8f8c4c29f7a4290f3fbe963d64c4ccf90fc94c4d03468eb9ccf1dadef02abc073ecf
z64b8e481d70556b1b55992bb5861be7b9316add0fffffa444c3631b54b04945b2eb4666aeb78b1
zc5550207c936800cc2b708272567937453b8ce8363658fed1407afc4327d23f0bd4b840771f444
ze6e5010bc2b47dd04c83f1731073c04b4a346d2e8879db104148239eef59f1f3dead3411e030bc
z7d67f784a9bf50d7eaf4653e93477364a1decb2c168179352be0df1267e7f13300ff9c3c1109a2
z9fc84d344dd65c451bb13d1b589947b0d02d1d2d60adbef2161e92395c61d6c4f2c14f8d2dee5a
zf7e7e979ecb145c323230bedcbe65e1f584d7ba92c552e2cfc3e05cb9205d570f9b9076e0e0f15
z03b006a9520a628d78e225a154ea596d38a58b17f3744a67e8cc018bf9100ab10757810590684d
z4c4803a294a9bb8050a3a30980ef2b2f51785930b3ea21124ca7dd1b3b3df964caba21a70d2f9b
z795f79d6635bba7f49bd385c25f4414afd083ba893feef284c65ff578d6bc0d2dd79a6a4746bb5
z6bc1bd7c10f6a331301156e3051a2445229197cb293518cdceb6bc1659f94d3b94099ca466084b
zca7391f1602d213512a3ecff3ad2876eab93b8121985bf9b7cafd18923e5e6d037b9bb4b27a78e
z40b74bd6c2712e557e4e855c65f61619d03ad8aeb03a40cf8e8341bd406ad5779e52576d5acb86
z4b4fc573213926638aa58b30399e09f8d696eff51b794ec3e93076a6e227b1dd6b2005a54baa37
z8489d579f591153871d19f163c393e60c75839df45e81760ed1ff628f33599155d7fb5ca1c758a
za25d2b3d8a03c69c5fcb489db0357cc6f5755daf01f34f2c40ffb8ae062f16a5926c9b4984ccd4
z9a6627b37d6eb17b2046c4fcc40a783e91b7405376c8fa62dadc2ff9cf7f5e9e2d1b809f8b70bf
z7dedf413072d0aca1adc5801608f3109ec5f853bcb1b269d3143440a257e1b67cf135e193ecdc6
z506db71988198d2170183c856827ec9c5918b5f07dbccbccf4894eea5a60512b1a907202225a4a
z0d11f461644b6fd0fda54ea7de0348fe396a48ec2c7231f92f16ee530413cdfe68026774cd2773
zc00dd1382eb25b58a706009243f505baacf66af235ab09d39c93581591eb5cdc63c5c7317960ff
z8f2c5999151506c3a9db0206702733b5832c9fb3acf50685e7a8ec9340b7d15282c5795b4f9876
z48c06d62332c8c75a25ac7a3b8ad39b268562943bba533571423b11892d6d04680fb940f68773d
zae3a7b1495daae44e1c3f9800db8b69991860aec494d6180d29712a2f24e00f21341947d4ca5b2
z93a8565667675ca635c121ed2228c330ce8ca005ec0f8c64a370fc4850552601fa88dbb8626bdf
z362dd8dcfd50ae1a52349daf620aba40eaea2b0f8b8bea2ca3362b24b60e524ffe7d40f99b8a43
zee56fface62e323968ec29bc34447574d9380d6d3c1b8917f0c3ebb3b772f05552bdb631f55870
zf40e207c11ff54fe7556fa3cd17ed69d820370dbd744ea4fa1a158b57129b3057899609d0f0396
zfb0a2b39be70114773e3de9e3b40b9592763989a5241a36589c90b2df4f8f4032f5186fb7be4df
zf7e2406bbfe779285de253a5aa09a39c0fc678e7df32992c3ced147e8ed4a8d92cccceaca1e5d9
zb1c443b1793f272a0c646eac491acf609e5af83531522401613740b2e2b6d8244aceae6548609e
z62470fdc7b4b66ff9a3d024be4fe49ebdaa556ff7b2aa5971653a20a5e4ba6fad47d6784647163
z6bde9b874d668d577fb9c980c00be14d8a888f12feabeabe11db332c3e855b5c2f86a77b454059
ze6b0e616ef30f080e32000e266f5af6d59b5447baaf93ea29188c5641948762bdf227b94217178
zbc44f9119e3e47f36b0ef294120bbf2ad5c681bccd913bbf1079badf1f6c24914ede33c2a15d2d
ze501dd61360a03d05eeb8f7923080941d6bad0259c40ab53adead28d178a85001de905bedad73b
z87e9f63ed8c18f41b10a8e91247ddc1f18963ce6ab9aca7d1936e4309fbe7e258ea27f9b10b246
z57b820967d86921c6b09a093c848f41903d9116847cb2888eb3446ab307ba15d04468671e71010
zf48065cd45d60241b474e628e6d553f8f74db1946a5cf1a362f573f5b56d1e395d825215f9c7a5
zd926cd2f7b75a695d0859434b83fd3c84e30329226e90e329ec100a97807def5dd1bb61fa22f82
zc9e1f74df2781946a9bd960b990a2a979b0e23c968fb204e25a2a1decf19e3d1b1590299d06ee0
z7370eb5dd805c3a2e46c47676c6dfb2d3839fd8625e51653135fcd70498d4f433fa5e2112ec21c
z2cd9b106445aa499fc2aa5a70a2a23ebbe561a1462b31bcd13ed3b2f5882c4779b38a8c51174a3
z5eb276012b729efc0cca4b1674876acd4c282bba3e71c8339195465342be380d43bda9058e9df9
z415f92b233456ee9f04ed18b74632fdb6bb960829d48160ba47e3346594e70baf847df98f8be97
z8f73526df01c8c29200563e2a6e58a36aedf8cb944c9ed5d6548902378b78174fc781c3d746504
z97911d8cd69106c2b94bf9928afa6f31dbf739a9c3959e147c8fb964c327f20ad85e0b66859b5b
zb2ab137bf1fa3bc50a4e4fd7ced0ef65a294dfead06e11d5246923ec0ec0b8953c344792fe1dce
zec27445e9eafde7f10c4333403c945095f70d02ab0ad81c4c8d6dfc1be64f4d938855d50ef0e8f
zc78df2f559883298cf6008f1431ed9c12af3927152e1b73746c1b63b1f87f0516de5cfdc321af3
z3020dcf764f10cc5137b9f1ac91061eb6e863e1033d7e74b3a0e8b2ca5ba32ace25211853b3199
z3dafbf62496f7b0c19eb483f9e676b0bf10876758e1249ab88dccbdf287ff2c1fe10ba0247518c
z6e13826138b274a8acd17368357b5929039e163c1bc93ec930edf94aa513d4552b0f2316f0e397
z66c5a095c0572ffbfae9bdf0cbbca20efafc73b4c76437b596bf5cc9b4a06c787e510e930962ed
z0d5371e133d610541f83086df62dc73cba0fe0f2719ea3e3183c4c3bd1e2f92c5b639be12c368a
z72ceb952f6e76940188886d9bdbb710ee4859d324569d89e5a1843042752d3cc433e7a220dbb21
zf7dea307284d87975d46508f6f0cfd1b3bfbb0d4638b4a932a500a072cb0228f590611ee3ad45a
z7fc454f53ef959389267eeb3164ff9a15379c3aaf226f649e088c0cceb748445f03130cb1171b5
z51542c7d193157a09b03b334adfd6f23babc216e55d1bd41f06c815847ca0272b9e43c0bda8e9e
z7f9cfc1edca5927a01cb2918f8af8763c2236c591f6cc639f29b16c8bec6931650e933175afb52
zfab087e6788b4cde085964a43fe8aa9b31149ba5a3530040565b7ccb54bf897e0e664ffbad5f78
zb39454ec3a5a7636436e8d711e188621766eea9766133b0208931045eb84eb778d8a949a87c8a2
zdd8f31f9350c825725a1ae18db3da45435b8733f2dd77315cb6657f88252ec01d9fd5ce408819c
z8df7d827f8bf2a34072d44e15fa979c667ae65f1d9bace813a7fdfed370194105c9a0a37dc15c4
zd55d1b9f0cf22a523dfa6f135d2ae26c2242b93e3d20e04b651e556802e83dc546ab7ed52d534c
za22922ba4ab9a534d39ad36f35035b146311406cb12bdc6ba3202a35adfc799853d684d295726e
z0ed75c09940a901c711cd994e0a47b022f47d79488650b572a3e8f5ebd323a416ffb6bfdec78e1
zd9be0d6b4f183ccb75d1c06bbd9df952d699c5291a80deb9ce05269222235f91bd1b543f1c3729
zbaaed60805325e392ea8ac8505d735948d3736b758a32af14de313ec76de3ddb2c96c41be33a66
zef66124a5f2964d7805d732e5424597ef50eb15698414b9b96f7b91e0aca4f391ca9a1ba2624f8
z1cace5ce514b876253714ad4f2c0e6e72a15c3e0df6806693e64fa8965b5cb656738a992bd135c
z9e9323b01c3248c3c6a642a8963d15f415df411d21b6ee9f175c76fe8cfb682f112cd56c27db67
z3cb5f65002034fe73ec626e6518a216f812478fe4e3a5aa8af5eda0fb14a998d6b8dad19d677df
z9d5dd177711fe2ac60296c18ecdfd09db67da228056f375d1e1c65116e3577ab9e1e76e2371e23
ze45aef7b4bb1aad7a0c68288f37d50f1e0301ca997d5cb6c37692ef215c7f1096bf36b6a08c306
z94f829b318d1f4e31008d7fbad50311566c83d6c1936f7b4002328dff405677ccb68dc5cfa9057
zf2e727e3fe2dc18dcd98ae4f9d3a6f9d6db2de7f615d16d59f87c832f678fd556a6666dd16f370
z827b791e996033ab73a1e87a21c6037631de8db7044a805c9882492c33324aa53ba4ae59e341ab
zc186fc8c7633639d16a42cd296a4ca921959fafb3ae6dfcd9f9d79db1c65177cc78172aed422a5
z8f9765d69ac455e5f79a36e86bf2fbe64537cfd9e1751ae15dfda2d51a46d24399bbd5bb82bf67
za02e7a9be10e2acafc2e1c7eb5047fe473c78ad0a05e640351c9787f50dab02cbb2e3932764da1
zfb50dc7990b8006ff6e725a7e27838c9b3df124378eff48ee667aadeeac69dc285f7e3b69678ad
za2fc20d6258d8a8ebfb4a8836d1c3235d5d8066cdbe6c1bfeab611c141977a90f5d64454a50887
z1628f1eee5d0e35e5f78ba602c7ee4f51d4cb34c21be36f799b81161df0daafb00db82d5f4c614
zecc8d575c1de9b7b11d8f4b24070f3cbf9c66cac49e42b19a38ae697d994a2178d5e27e9fd5f55
zd53ca383d367c0de02d0c54b08a6d9cb98de0125dea1212b89596413bd0a4ddc3dde831d538aba
z9a2a76c3c411545f5ebc61f52b946a9ad19d3fd77399bd439f54267f8ad55362c2f272dfd40405
z4072285030335c45792b1748f7bcefffc4141ebdd7a90a6fa60cea98954f7e04c0542ae290987f
z78a32d00203ef26dfcb2dd978c78d550aa63acf28d889493eed6cfb57bc5fbdceafa9e08fbabfb
zdd6d032e3052cc31e89f77c0d58cec32ec5ffbb84eda4edda236c23019eecb6bfaf241a8f002ff
zd41ca9c7381d85644bb4040c62a4eb96e283babdf8ed6f99f7cc34e3f1c0dbd54f698953ec2d26
z114762cba5d059c90cdea1f276d9e19b75a68fc64ada4016725a2e807606f3fac1392aa66c5e59
zbb4b6c2ef3c682bb56983d058c95363122cddd0b9c931a002f9117948b01c8ddea9177d07288e1
z587eea70af83c710cbcb844ba75912a306fe9e437a15802c13b781bdbdfcea77f324822a3a3b44
za5e8678421a3b0298caa3b9f6a97027dca7a0f3033b0bbefbc7033d409a4b3010646e4f7a6a678
z7b4a211e1baf693f2d56d0911c90388bdffe2a2d423fa7606d53de3b9954e3aec14ca367557682
zcf56381debc759cbde5754cf993f79dae871e8dfbba0a4169f85b8ee3d71d03dfab42b260cd0b2
z2b5d12510e2b834b531ce5ca17b3eb37a297ea5448615ccd45a47444f1107442164a5a5f802558
z801c78b1a222bd38d73c40eb1ab0714a6102a1778b4cef4a174c49e549f86aab5f17e4889945f6
z5590fa534b638d2f3b508fd50ae58c26571608c7fa0f409bc487098e5bdca6b2859040c8705415
ze3af6bc5be2db53fadeac664ddf88f5b90966b0872d27626a6a5143502918b40717ca8c3d977e0
ze89571fe0895981d2cb698daddfb5355d29ed98227f0446dcdfa7c3e6f8f235658243bc1f15bb2
z74ae452a80bf0dc20238200e4821b91b9c271bd952d45dc3c067965fec2557fb872bc5a4b5d193
z00b24800dabaa6c4d3bc5d3a8dcf8e84db1f442fc715f6d43b846e1f6ef0d6e7db4cfca5820a1a
z9750053d940312dcc78c7227463cfccebac01ebacdf5412ff957915ec9253bd0a0d7dffed22861
z536cf8885738a40f5a26d015577b582db8161e37fd643f392e69e9d23518564103330362f49e57
z15ccb3a533f8712c444cdc9e72e79e17f42318192099d6bdeb2058ae1d13565a0b719c6ea99c25
ze123004852a8f4031968a18b727e82bfc78e9e7a561be6363f5a5934c3029712075b3735639d8d
zf734fa22460f644f2db4a7fefda547a05bc15b45ed213326679c7cbc156bdd30ea6eb030900872
z4bad36417f532dc7273c7328f40154ee321b9f4a63c39193831aadbd076e01ad000bcdc10b0915
zd8ae6818c00e3bb1c13065d0343893b8b766dde2e4513165c1c7c525e83f6e166b16002991d0e1
z706be81d959ab77edb0f7a482bbfb4802a0021d155e3d5bca08e5d5eeb1bc988cb940297bf869a
z82ac3726070c8006b21bfca0be369db909a2a5c60c5154a3b5a67a8ff5b52218460c75893a362b
zd54f20b21cbd774a7f48732040b88ecb4024c722755f5eb418b64a9285505f49e50baa60d98257
z0a781ed2d178edc93561f931bb586ca796bb7d8cd99287df42f9ea0dc624a39b420a2c79918cf3
z091ed15b165a2d052d2e372fa0f5234d4f42f5e3874a379ab1345e8f08cd8988ab23c5e1f0ce16
zf8ebdab37aa4a1264527e1d471bb1400cbbed9f23fa92c1e32343f3696af6bb7278e44980e3d57
z6efdc27fb9148228209191245c8585f993aae9a85fd3b1c107ca7ddfd60a3e311933814260fb9e
zd78613eb216c9fa73cde635b76761864e1daf643641ff6bcaed8ebfdf3694bf1bf15193ccccb00
z1fce2308b3149e7af83f6a51f887d57fc3d0e0879717af12010e3fb24b42fbe724fb82ccac9f7b
zcff0719bdf8c86704221a31be42a7f20d72f0fd67f0769f6c844e4bab4c9c18b3392faec0573af
z30242f2ca90212d3a5f64157ae63d9c2bc5203ce86259d5cbf87fb91e6b0055e9faa0b15634a14
zffecec54a008542603374bb7c983cbb3f27fb0af4b2dcb5364d34867a3ee36064665b98f1b4c8a
zec6949d1ed0c8283598bff226c4ccb2c3fddc4ead5710a3c0cb2381d2160ed9af822e182029a2c
z1bd76da89f3d0e23ded5dec2b9a3f3536d6dfd1f9b6c3487b82282fddd684f2390ea29c93409d3
z46bf575b949a7e828188e342ed7c3a99c399f96c2d9124dfb719bf61d0969e2fa8e88bf47ec5fd
z799fff25ee08d0f372c93cb07b6b5fdd92acfbf28689db9fb047e0d5da020d7b275777632bea61
zac7f6fc3df544cf0e15b4be5d2b2f4605df534832c3b7698305b02e3f7afbfb8fa69ea4923061f
z73346661568f5e6d800eaedfc61ecbecf96d7721d487b14dcb494a4b0aa11d9a4b3cca5a36cdae
za445bbf7b5ce27875bcf957e97bc1160cefd3b480304208cc062617bde7fec9c293fec0cb2b1a1
z59e0888a593703b44207c0bd42c8095fd42b66f5adbfbf7cb3b3c931195f213a3fc8abc79b44d0
ze8fe21e9db9f5dc775a314f78e7ed2345ffdf446a5ea63350901550b7adfb168858b54cb0ae650
z572f6e4c9a015d65156f87fb7a2040d819ca2913e8c7882e13d70d827ae1d3a5c045057b66f0a9
z4a3bc58aae39b11e02759b8fae5f58f109b939c5a6c9c4bad7274281ed2ee00e73672e880f73e1
zea5aca2da5420ffa579bef57961a980668e0abdca3ed058c2729ebc617d89a51703f7c7e5ee2dc
z0a434ae4c88b75e71f4fc22a7c2407216a2e702ed3271c9de08e02c6fb15c9d2a9ee4e303bf0d9
zcbeef6c43e02429e23054c57d68018775a0ff64efee5bb0f593ac8093271872d3a1abdcc1243b5
z7b7d8cc759654b2d18b2837d4781385f1bda088f19cdecf859a5039b1057b8790bb613821554e3
z0057712e09240ea84f8a7ffcb963d266f84ffda5f341b777d04f08520bb036df5b1305575da825
z00ca0b3f19741cbd71dceab27fec1481ae18d423ffea1fc235e0a78288df9fb4c80cfe4a28a40b
z4b30368d98b682265614b5acec5500ad3c921f62745e03d95295dac5d5efaf7a8a28d49a8ee164
z23e1fac8a0e25759e43449509eb642f3de97eae40cbd9708c3330158e7213e902a548b6a346384
z3538377cad08da4b43a0a7b0363f23cc310302b5996b7531392570095ff47c79292bf45958383e
zea0a6e00ddc9f4ab2b8c9ab54b2ce95b4cc48531c0a419b097309b7ecb179033470fe75ecda2bd
z02d4979e326b1733907eae5b7a135a4f7956949438b77532990a928e9ba7b948db629974618866
ze50b83e6f03199a01878e6dd72cb81e1522c8b80dad031227288fadb463f064db6027c144b7b59
zff14e64945b7d5730069b06a3b5af0046ba1294028dd59c73ceb30410d608898e92bd9fb317186
z9fcb5fdb708e4c15fa1fdd301a342703574f06344bd77cece1da81fae80d7f675b76438e613115
z70f2f080f679243fd26cd481f6bd3d47d7d1aa9590987e96a74a0e6872f23465d6f5379916c5ee
z9d8b4932cd8e869b03eede860646a701402aaf2840b2c1d1defaf57d785e0fd3f9b352d029e7f8
zb18bcb06b5e9629fc71a085c62ee12417d0c32fa0605ef7288a46c72c8422673bf9280c8054926
z12169b1e2577bf66df8ff7c7afb9ef6dcc09794042cacc3b502730dbf1bafe16f40d39f4857a04
zd0b9f3fb07cce1682b33667ee3ba3a4fee9970f05b2e78d6ceb150777858db0ce49e4a03374fe5
zd21e92de71316ca738aef9d097edd1ad8cd0cd52a868a6f09fba322aaa1d77e61419f175594004
z1f933216e0ae4eb83e9fe09e6e2cc5fd92972f21c19026e9e89236488e0e458f5ca57f145e4b43
z423e556cb0f76ae1c9c77548f6e1bad942cf5445f6f933984d6e1a9ebc39e2f0973c83f6193185
z47cd44d5ef15a9ecc132f9a1fb1da5c963b24c4b07f576790d3a00c1bc585b83cbcad5560f964f
ze9c409f252db7f57ab46633940a3ab0dcbbe6045ed266e6856c1e7bc5c8b8a4efbc6bd9368a170
z209afc485eae4764d201e70d7a779a5af6333f404dca557c0fcf99c26dded62a0085fc6588a895
zdc77577f4d3e962cf54d1243fdfb5e4ca80ca5cecf00fd05661bf46c544cf14a9ba9600e356a23
zdff7b518a0d904f9b20ccc69536d1bbcb2dfa50c67d0f5524340fa7d206de0c10d53ebf6754724
ze607f9a75c2beae57a569dfffc95127203e82a6daad2379e6d510db8471a1b64c69418d20a03c8
z0c9f7941ad4c6dae2656e03fc3db409ac059414a5d5179adb266cfacf1469d74b77389402a8ff4
z77f64a33c5b91afe8e7572bd9bac267776f29e1d81e8dc0c8ac27d8b56f8690990ef6d706e8906
zb99624425005a1342b7d7c758141e228df6300c53caaafaacb0e1c0c2cb75ce31d78f15c8743d3
z324cba1ac47b16a513012839c6339dfe696b7f5155753c10c91a1bb15285b628fcc06febfaf838
z6f1b8bc5ac72cbfc66a8fefe9c233a4fda7c9708391a4ed6b14017a3eb32567ed7d146239cc078
z231f9f809ec8ae97fe3aeaf3ef372364d2e79783a5313f3ef8bb874220ae3bdc8ce3ccffec4931
zcaf98442b90f7e8a6f707b5ead5227bc493e807936bf5c352e028b4a448b38634e31dde99146ec
za0fb511458240dc772d746c218794ad66037805d217c3ceb456301b8df29ff1d145648709ccd00
z09191f20b8c16bdbf02e360b32b7160c5a90a1990c4e02b5a6a74e0b24a988682b3c770e673d21
zcc7d5bf22206763296c78507c4b733ee362dae2765cec0288c676814d2ad2a1d115fcafcffb57f
za2e238c311f1a5912e4e051a3a7fdb49ee81f2966c2bcbaf2eff62147f99465920ab0f6dec117e
z5a139833b88445be7d1a44e1b78c3ac3a6e4b3238df576201d916f3562add16f1aca890a19fc14
zd1b6c8f2ddb40b41b5bca12f1f277c5f0d4969fe70b7b46e00e716aa81463b9ca9a5540535cda6
z189547ab0dc0665107def4a23d9931648bb43175293d4982862b2f60acc40834d58be90e78ed6d
z01130a005a8fcbde5bff07413764998a9b0b97662cfad589f37be9395a85c49c6d86a538bfa8c2
z52d461fd3d5ae679195f0bb6281f1cfae91f0da1070110c5d5a87f8f4e1308873915927673b4b5
z333017944e309a1f70806ded5b14330c57e561fe96613d0ed0e8645b58cafef8f64c9a19518028
zd4e68f2c4fd30c7a699271ea5d545d44fc311f935670a3fffb5c179f1b1d5c69197bc083a5d76a
zed3b217f6b62e150910ca8d8f405dc11dbda431e8ddcb7497103d42830ce7500c8240806137a38
zfc3ad8f03a9e87652c29f02d4e09704ba419401aa4883699735b1814febd1a1a54fb7856f1d236
z8195ea3f66f9fae77398df5f06e1468aa1e40715badfddfb9294e88bbb8f6ccb63a96f982f69fa
z10f7d4c6d68f87688c7ae373b0f77b7f71f4b7edb4ae64f819236ddf747e8f90ff3b9a71aaef3b
zb545acf785fabe18c6fb2471db667e7f542386407d360ec955f9f0b328e6875a51fdc83b4e2f8e
z98b38e6c5c7fa5dfc557151bdacbc038b6a5697b0070a76fa761ac927eb5156909183f3aca4a54
z152348af6323c098a5a2e136ee66728bd16b14fdc7e8900dd3102010fbfbb2aa6f92a0b32b78c4
zc18318aa92f0d3a6b2b939588f498043da28b1cbff51d28a8e9da721a2046c661b8c23dcaf3554
z5acde388f45417af9fd773cf0da251c2ad887151f0e1841c7337d68f74f3b3021311e10a567beb
ze89bd327843dd4d1be047ec0a3a3d897510e904878f89a28866a956d48305d923d9015ff785d81
z4f8a89bbc846fdd5e7bf348124b01d1d845a0200c61191ffef94d2a2bff1d7da68dfeca671c7b8
z3c5fc5467c4d599e05832c2adca0410e7216e26323fa068b318abf95413bf042ef08deab4cc491
zfdb45019bb713510ec234ce537acc067870b043da8ab8833957d0f85335051ac058cce277c19c6
zaa1bf903243b383b712d76f7a2c67957efdfc2b8fba29a328839a9a90af640f73b817ffe290900
z8a1050a77b1d2a42064069cde135d566273458f0d0cea07e5b08a6f3d2dcc862df04dd1b56f72d
z327f7922f9094f75e4debf747f0bb90744c71da1ef5de98a4ae51ae609539b04e034fd42f0648c
z7d395f5d9c4e5b57c3cfddf6c22eaeefbd5e22d9d3b9f8b3b6cdfeb019864751f78c6838c02652
zef61d6aa9f360d9840a63368b2b70d1c7828356c766d83b12a1305277d93a5b34ff5de966e4857
z68dd63f62aa7bf563e2846fec2688b2e9920fb7f2d1d212bbc3cfb10100da1f2f67fdcb0f1fde7
zf0aa97ea30d4043f5accbfcf21f214a1e6b84e03dc08583feb0623cc743d9ac36325baab731d99
z60eef1565b44daa8527318df09686614e7852f632a707f3e24f0004a941a5cfd65a8de85ec9369
z67c878faa0bac24edb1adeed4928f38eecbba60e0661fc9f637fb173763aa1962dc52b56ab7f1d
z18f9b7fd5843105ee840672f41b5f9d20f6052c0d9bb1422fe8d49eae586395cd3add53ef6fdb7
z23a7b5d99114f486b4b1508fa522a80ea54bd9f26771cdc85a7a413b3d6945005def6397c8552f
z5c38f7cbe4d4169934bdd95e326c29865fdac3258952864c5381960272522648cec154cb235c17
z2e92726c7d761016f86333d88d64729c65cd5896f67d08c4a04849b9d55ff40277f97fea40932d
zcdae605711d62612cbd6725586c70b97b481afbbc4ad4be17e8c0b6cb4fa9a727b13648505d341
z5e2952cb926ab02316cf34467320a5162635579c02eb32c647563e3853eaeaac8a343d71f0ee41
z284e345a1a507798980c28ef3a7c83f0e97494ae53cfa7eedb5715ffb14b70d61cbc31e2dfa05d
za66cc3204df6f48c21d9fb7ec727b99119857387ff4ce3ea2baf6417f3d2615e18e82abcc712dd
z52eefef382eeac10ca9ed44a8507c88b0274357f484c211b9354f12b6c850ffc8debf9a590e76d
z05fb32d65dd02e97e57347986e72953107d1410c4e0461dcdbd99c12a1d9c54e87ca814f945244
zcf1045b3a545d72d791f844ae4da8a0eab22cf883bfae0450c518a2d6c07d5876c63853da87764
zfa156cb17dda32e5e34ed1e23dd39f14fbd200071e35caea4bf9a5be6a71193972d26609058a9f
zbc841dec0b5702b9b8464b2bdef222603648c26ad2de9ec0bafb9f7365321b5945a6c59d1ef7aa
za5b8f7a43df9b1242977be00c5660b937a938597ed772c6bf2ecec1b473d35a963da5057328df1
zfc019bca557be5bb02322a67a24fcb4a30c0dc829751511f07e59839cc83cb93e4a014c379cda9
za87c93e837109b539d58772faabadff100ee021aad33ef60f0eca149854db31f31f5e798a53676
ze2f85ad9baf595f76bbc400e7588172be9c15edc9c13d0ab9235c68a8d6077d76ba8726357349b
ze146bc6dbb0ebfc20b3a2b8dea1aea9d02aa2ac671e5f22996fd3a4f1bcbc3336384baf2925506
z1f0b9563d3cb1578b550f22b68ee5604d8569a9669129d912f6e5c32a57c44327bc30feaa868f7
z4421e0cdfd785468317bd1acb0d6bcf1eab32a8194611bb92bbfd52c9e3516dd8533633215b6de
za8e01cbe54c2e4f1892c9e85375760c4be1609b8292d16aa40f00f04eab2f6935bedbb53b45241
z3eeac401624c51315b99f0298e4f71bd9a78d54330efb1162ae11f1b5167fd8a5cbbac0fcad2dc
z2de47893e2ab8579cddcf8955fc0bc938b46c412efd7c587451740ade3e0dabc94adb48960f207
z0688a34f0118d3fbf91255ee10f1ef96990de790c2577eb37e46ee015747de021dae68c627021a
zf1d3a9b83e425da5b4869ce95d66ed0746393ad8005a39b6167fe27230a093b1810b7cb974d0a8
z1e78e83f7becec3a1679394a53297b185df06f214673512395db59e4e57dc99db932855d21c03f
z711d6deca0c5ee9ff625bcea5a4632b7f25a42b6983e3e97b0607a66ea663cd0f0fc6c28c9b1c6
zb6cd2b457b5a6b4834e4ca308cfdd233c382f1105986554d139e8a0ef0ced132abcb4c68e76c2f
z31670c48d27308bba63f91e8054f40219735f51e5cdb0739dfa661dd884b061d912675338f78fc
z4049aa4df87c109bf8f707b27014d2056d7fde7ad9a5c57d672ccdd847856f89bbbd0578f1f80d
z6cfd04b0267b843b4be5cf0d5bd30f8c0d367de2e8afa9a6758000aba87254ef0ba62a9fd9e325
z2497850992d313836cbf7b78730c6c7f5d72c0462972a34af927208438c27b88f94c0aaf89ed98
zbf644d8de029bb998b8bf60f3447e9c196b855f51f376f49652eaa317af64069713db3934bd202
z62cdb02e984ac371cd4a579e446808a08408ba3250469e422721885766469abfd89f41ecd169dd
z93074623ada17e6b0cf03452b5544697fec923d78399ab85fde14b2b2f5ba94fb24700532c28a1
z6f72fcd07b4d74d7217180c76fe0e711c2bcc28d11e07dd7f6eebf58112fc4da32c7801abf086d
z1d0af127dce38678cbcab16d0433e6a42f839c2f120bf41bb94812735bab44673f89dd099a287b
z6fc6693d0da2feae92da301c0910bee312098a54b7d6139d51e3c5ebda205480aa859fc6d0ebf3
z639f7d948b1647157fda293ad97924e4e612ba93cf23037d74a9e8858d00b5624d4077911d002a
z1a4a48ef5036427e184a5d303b2d9ba15f7ae1c4ab9bd77e337feb9916b198eaa16d652fc045ca
z6e1158d4d4d8c1e99c1a249700deeef9bb07e1b15395c302a6e0c9b7f2b83682517e412888a5cf
z1e3a5c065a008fd50a860ab620f9fe3801417fcbf8ad2313faa37ab8d7161ee8190226f8dcc021
z8910bf78b05804a9b087f1a0f021351e7f0c2dba42d9161dce296ff8bc34d98417c91900736aeb
z03a92ca961ed29b5225821356c9eefdaeace44139441027f61a5193243f856133eb03990413350
z58c867495e397ab2bfa45f175774c082c40f485eba4ccff3b324f3209cfb962a38ae19be2bad5a
z3a196a3c77a4c284d8f07533d0297e97bba29c725e5eaaa9a4a0bfd3367b01284095222e5425d9
z7175124d4be4f90117ceaedc78e4101161053227908d089f57f89255139e483a3bfaa93bede219
za93599d890076e01a0f3357db0846bb543114fe308ad6831f2f7f2f558c3dd024367a8d2c0893d
z349963e78fb7595832f690560df0aa95d188620792ab94f8ce3fa1b75ecd0fd962c4f63993e9c1
z9df99dca9dc8cb78f573f19af115caeacd966735468583812c32b7b4bae05addb85906e08d075d
zb3343912ec5c1a3cbde886c41b935f53c83d59fbf9ef7c0ee8781180ce7ac56e9eedc8d6afc624
z95dae8c7cfac6d734258bee2007bb9961fa00f9b6d6a5d26a0b5454c0b76edb705afcf2b9a7b89
za668b77f5d01dc9af6300d4bd3a93668d154da487d891a6b966c97163528a6f7938e2abcdba4db
z0a61e1e596659cb8f095d412d66aa22d41cae4ee8f321222ab0260efee32ae3c102fa32d64c6ff
zb5c502ae32708d6af96692a6f6ca961f610f317e3e1bb7eb9d8d76515223b81d1e1bfa51384b4c
z881cf8e1eff9a801aa4279d1c5a0f2572bbbacd2c9ae17c4efd13fd83a27ef9ee0c96e479a2a23
z8908e0937b02a6120c6f5fad7f01a33d1d13893fbf44da153a8b865b6b6254b85441bbf30ac7a6
z37a35fc08fc03042ba62d5b77f275408237236a004aaf9a9b88deacbc060e9ca75b0165b67f8fc
z42c1f0c023607fbb9eb2cfe5b9cfb1bd30f76280e616e69d0ee0090b0c0a2d9c75af637112acb3
z4023a20a06c53e92a0843343ad6141433478c7f97f14e14f754fe11dd60ea0fb1b068065cee4aa
z41e6340a8c7735716b135f83318fa9b56aa5446d725d166f020a60c71a32786a681a5811ed52a4
z79d4ae187c40ba440ba65dd75f7b49315f7afe5b7dc637a997968a930e11ed4d8b08641e36bacc
z18d8ce48ddbda0fd8256326b44cb65bc2f0a8d8ed7ab848e81c80d98be5327de745f2e1cdd18e8
zfc3f712371fff3d0489ac1834ca40dbd14af7b6b30a3a371fa759218553a981113d4eb86715a51
za58e9e333b1fcd5f3275609b0d3a920819242dd1adbaba8e856a15e82f969d12df22680694ea65
zad8b8fb57e497f594b1e431b8988e417c19c7a1eb02bbb144a8ae716d2f4a75f0d8b8332905449
zbda3173f0958a87285710cd2a614a34386b902f21191495ed6f7c76c064875e4b68881ddc25c0c
z2904253c7d9ba6027937ffaa66fc577b469351687e54a7a88d0dfcbf0d0f437623117638a2d3db
z42dd56d8f81108ac8ad243de1251dbc1c60050ce44933f93ef25bca093f2c665d995e6b80ac5da
z4ca2804e16bce3fa8f0e48a7da16bf9e15b3c1566bb4a27087058802afd44e54d2c2908d4e6c05
zc60de11937256bcbfc24f34ccdc0324c585742839b7e35699b9d7a3a1bee07035457a9714285e5
z822c77aa314a69e045b79040e326470c47bc91eed609a520e84fb52c254a6ae1d1b737ef82b9ac
z431065dbc6bfcb813ceeed6bcd8b0eda0985cc0825a7218908668ad8a3af58773f87573ee3b074
za3f28b932068170e107b3ece181343fdd5728f86bbd5fc10a0b7e6444a104677ae0cc357efdaf5
zcbb1620befe8e037dfb76d9445de8b37a3f3b8be726a4b90dab8dc90ec2235ef67da3603dcf7a7
za6b42f9add492f95977f3651860110fb02857148a01b6460b977ab1994b6a50f88f6e59c23838b
z892b56cf182beb63fa18da994213c04fc07416ffaf920d9890fe37e9b09c76df1f16d54924f21e
zb1027ad54522728593d57e34065111b49d2b97531c872a11b075dffaaab749c65cb4f365640cf2
ze8d20816ce87df44bb5871cf97385a90591cda06b1824d0290d46c7c4f8f806b24bc70500fc677
z23b737f5ab3e264bbce858b1686eae6f0895cb6f62c468e9ec763896edf572e82a081cfe08e079
z37201f379c5b256caa4455e63c361b37595a6d7268aa544ca42419da4199d975564a6fa0d41f6a
z0f4406ff61b978643bf0053891780fce21005bd6686b2a92102630f7a5af6feb7a471350402aa2
z949c49efd4a7df832036a766924fc912eaf37cb12a614fbc7594436043252438c1fad9c99fce21
zb5e3910863af3180987cf75fd81723fc67fc7702ff518460230799a6dd7ffc034ed47ab38bdf59
z4e6acba68eb8364e7653dcc36de4a434b904340d0442ec39dcf155a5e19603906028063492c53f
za64a3f864861993499cdb93ae73e33db8cdafa96807354dad62750ae78f6e9e20f18e6dd695e25
z08cbd4609ff74f4a99c254b37a302c453b3f47e0240a8e8f40d57043e372e8b4469f51d308b7c3
z23809794b1bfe85e37b8dc773f2af4fa90a6707bf35d8f8be89c5681e7d332bc20b526e23bae19
z625aadf434827b647b609ec3b44d0285a439f429875e952f0da410d5a1ee99201c22e9c7c6fbe6
z9e82f92691a7a2f29dc2e81236e108a2f2043267ca6240d7f7ca9ae403e9eadb86ede72345afb5
z403e155152ca1f41528e893ea9f6b4144f085f28510bcefebf0da884b701ac55b31421f06fab5d
z8b2f3d98b05b3246e2807deceed2b2c15b39e8dd3a877f116dca3db821c4baa442a26c1019c6ba
z4307b6b749831281b2babf9059839ce8f57a263bcd0de336dcc8ca92e40ffbf92c8948c0bd398d
zb1a32573d642fbf979cc8be7e0928dd5e12c5dccbe0b294359129ddf30682b27a566f5db7ff2aa
z6624ed28df3949192c92bc463a322aa9140ae0c5c51fbd43fdb90f9fd5cd26b0715500b33b5743
za9c8d170ad44bd28a1854547aaf638fb0c7da952872b2e61f3a16958bf6e74e8ae8e08eea97b84
zd4c7e9b0f526f9fae03862c1751e20495bd109d3de23352fa2f918a1bce42851a0fcb81756ab67
zc4d0fb98c6a6873422ff66b3fc661b7d847d1740b24fa0fcb444be0550d6aab6aac6aca926e6ec
zcea26149a7e5670ebc6686fa757c1db253dcc6c7e414b0daab3b776afd4567fc5ac2507306c152
z8df5a58b2f3f9fc70045068c0a0097bc24fc00476ff8a45e711567f24f07a659eac0fa22cca432
z58687d3362750fe4ec383a4b1438bfc3d1d27182bd8c093a2c69403be2be3e9c7746822eb85ed5
zee2a833a4546110e9e210e370862a7f9910ba2d0d44ef6d7e97593da128539e620c21cdda33c23
z8204d827d7ceca3aa1b43667d9a9edfa64c18b7148d58fae614e249fa63e87e0cbde2b3386d26d
za59fc8cc62fba9acd6336711c4359ce4ce6b86a18da063610076e40553f2146581138555bc4801
z2e2ac04056661c8e0c89b61a5e9f95995c385c934290e6caf6cae7bc3231caa4cd467be485ac9b
z0a1bfb4872421f92c6cb1d525150585b44b23f255ce71c9e18594881f48ac00fa2868cdf860de7
z30bb7e7f0e19f43eaf5d77701905b491b2d5e5be0806662a185018ef88acc13e98592496e9c4c8
z70de5133985252eba523266cde8dd0773844df7cb1d55ee285608a4da13af368953a617d364944
zc304dbb4710dd72fe89df05dbe6bfd256ca4a6734fc09379889578045afe4e6d77370934b0fe5a
z3a903933893d45473b7b4d754f8374ad368a18ccbcc5fb2df2e390231a415c0823000258005120
z5b3557989d08b98e83709a1ecffb31ed58f7fde59ef2e9e3a3bdf7de2560f9deceee80d80fdc26
z2be8379a8743009933a5ae1e860e304d201f70fba8eb23ab603b7d9d7cd6805c724e470f0a924d
z6c8077ba1f781027f6cd213306676ef7a9f06239af625280a4f94784e89f8e0973eed300259aab
z2ed5147a8f50d692982c1c30fa2a7343ba735067994ebbd8f086569008b8f0284bbffc42abd191
z4f4eb193f484b8335f8fec113b8348dce00794db78b8293cdc37665a2c45ad0f77e54b270a8fda
z830bc43253be6315e847bfc748a0d03302cf3197d2f0c8f26802d952086c1e9fd034add5a88679
z88a56dcc6504c2722e44b112578102898bb152b109f1367ddbe8941aea759fd4537bd779eb4f25
z89acd742fa654c5ebf43d2dff287e9ecdc52cb6c254ffecbf8c2bb7207b0de55762f61da046b88
z3fc5fcaa6f96b2f0353e107802dbea4491482dd1f43cf65f8d500775979fdd0ba1c38d83ab3285
z8bed0dfd48ed61728da24bdfafef49eca149bcd46a180e9e03ab2ebba9d426639570acfa67815c
za518a3db0eb9dbb831b99143324c4b763fffd0b9a141d05099e3170af6418f7c87fdc9fea64fd2
z57115edd21296c146f78a57d3d78ba94fe1d87ca2b50243210036184e0fb2212acfc8e9d4aae5c
zbe7f894b43aeb4bed413aaa19a9eedee32fdfcfae7265dfc5d40bbd555d6d0a81ce22a86cef3c2
z8dba0a28e617b74e93c034f3c69d42b88cb06b64e1cad858a106169672ce4c80dd971ee220d6dd
z8d44e63e686e9aa0c07aa7c002eebdd26e89e1ae6b2ffd96233110cb26c7be901735bfa3b407d1
z093639703c53f712dfea9602ca037574dd851911e69ee897328fc8132e681d959e14b493e77a95
z9c529fc62b286925d4c7d821c5bcaccef96720b0875e4d5f28cb914a63574990375ab0874b034f
ze9af607122224339eac985aa128e92e41aa8b288d63f57ed077e33cf077f5da514004e059512de
z50e2c27008ad4b737bbbb22f591d0ac193f0427f60456d995e1ad1084aa249c8a6c8b8ea333426
z99eabda832704b17b9694796669c16f6b36495fcb7c469891cf5e2c9b2fbc35a53c772627a26c8
z2ece2d187a16d33bf5ffb7279dd200d455e66b0085e0e0479c7f5931327f8a04f899d94209ebc3
z7ed8787d9e40ca8c71c04b094cc6ab45dcb796a4b64fda12131f3cb658cac6bfa1125914a9bb07
zbf561fe68bedd9c9e1fd51b1524c3b3164f8c2a83c4b15079109991fdc7664783ec95a00834d02
z66cb387e038b819dbda6973ca07089273327a515a542abca33c9a0b65fa4e3eaa071a4e1346566
zc562a97676cb0b2f64cb9b1350f5b1fe733254475df67949963983fc7f4f296ebaab82bdbbca66
zf2b4ae509ffb3d9fe1f4c5b5a9d160402ab8a389883c677a52c2cd255f3ae279a411c01e892ff1
z6be66f3c807fa6664658fbbe7067d627dd628a0c6790c7b45f55b0e4a645afaafa915a155a9a00
zce0ab18a3a2efb7e1174c13b017692f7d2a4d14862d4daddc1aa2bf9bfe6a2109d0e9e46e2a1c0
z1d186b97056945c271eca56a7d04b907519c6c15b01b9437914e21f9964a51a8fa2f77922569ae
z61d5a512083d875f3f994039d1986e98c7a230fa7611b7d9a9088ecc750829d85370343b71641a
z4f6c022bba31344fac6f1c7b244eaed38e521a0d2171dcc533a8f2bbf82df318aadba3325a8586
z71556846547166f0e79b3ff41ef8ab3146827f089a22fdd250fae453296fe7c73b0e109904c641
z4d6ac000004f2a7f4c233f472d20ce36d88d6d7ebd8a76205cfea58df70dccdc666ca19b32a842
z0a026c24a16dc71ea2f5ccc0f806350450200ae56c52ba6b230999bfddfbc4b481a620481403ce
z8634b58927e43ac3b7f5f366039a03ba215efad7e8c506e466ea0a2c5d223e0c86aa7c29939e7b
zbc71f2d5ee169439ba1d4a0d8498f41f9a3e9d1b06dad082360756c4fe31dc29d075b340278bfe
zbe3d953a61e545ab290d9db76890c5d349ad737de64095c4ba897dfed7dae9a62b28d227a0d5c9
za2fad935e71677e40d23d8e01a77a8e85fcc13bcf7d5da87e20761e7fb2ce6601479fb7541d2dd
zd035dcbd701fc38190221d18761bd0ac12c564c9e450505673c93762985a76c9c021f3eb224c6c
za16c016992d0041803a75dff52e477aa2fdb41a08463d74ce2150dc6b423c40732a4b7da9a3945
zb0fd76f4ceb9a198567fa5dc98143230da1880e5b7c28100786ea0ec00b12c52ab783754fec840
z81e3d191a34db99004d3d79678e73a0c84c89cf127d8aae4bc31ccb0047612b96288e4bbe09819
z467f09104bef4ef96961096aa441a1f59fa14974cc980dbf55dde0d2b37b4be15661509cab564f
zb65fc2813c1b66f0c48eb24fcc4cd0fcb5560db18cc56d2d52729c9f6f3dde65ab348508c42682
z0584a12d69894f8057eb06ff9c3690669b5723a3bad411c2f9849c9d24a6ecd882659f0d34dd99
zabd887408decb955b37bc8e2af44ae00ff04d5d2a137f7df597bccfbf90edc6e26efc60d0d21a7
z98c59c376e63b7a3bfe34842ccddcd9af00228fe6eb0e38b9b625fbee3cabb66df3ab0c2a9c610
z0d15fe45d31c79d646e28d6222f24547681c81775739e5fdcfa6aa2777825808374de99c3d7712
z1ed46dbf45c6d90359144c6a60c9825a12062b5cee60cd453f1900a26f6cb12e9d0ade10979c6a
z92897f0d27faef376ddbc39ca2838579d9f1dc731f0df3c56f5de2d451b38e349aa307859cf722
z5d5194eef6393f732f38cc9d3363fc738b1308c9bb16e2cadfc896bee236ce236ba00f2aac560d
zc42addcb5011bcbd320b56c5ca6b30d9efb69bc9437bbd7ff3f922b7154c793bb7b5677d63ccc2
z65c125f7e191b3cd57c0d997dc30d2a88652560b345ddaf43e84da1be84f399cd262792055099d
zdd6654ba9479ec80ef8a00f4d9d7ee4e9a0168c8c5272e045f1b6f1944a37703fe9a1154b3fd58
z68b06a1fd668ac1a034e2b8f522e3f1c59c14639f3ff372fbbdbf07fbf55ea1b1152233c52e0e3
z223ec0fec6651fb067d86e2abc450ea8ad9a6a21c90d69b904bfb3290ef27dd95426e294973a6c
z9d8e8a31f6a10a9a0035b813d306fb4bc5f67eb3ca06c77f5eb2bf07dc81eb3ed98a92cff089fd
zf7c69d07e8d95d91176e9692dc224e4138584667aa1c6165f9fd8fc195e1d50e48f50b1d204739
zf21ea533465cb8f906fa81ec45c332697a7467239bab01bf3f9fe4c8012ce628e532e796c62c36
z5f2d5404343e7ee932db5211b505a947a4ce341bf22e50a96ce13dc2a3147365bde1d6c096ed3f
z7060075aec54952ad9d50ef870cbe784e56a256ce44c7feb0b9cc29aca0054329ac1b10759dd57
z12fdb763546b8a7f825478d0e5c7452b21989819ad4115b2a50cb1c488e01ea7890f3205b79696
z6bd298da56146ec15f2bb3acc86bfa81c2a3d9bd0ff4bd9c22d61eb1a15effbca60b2c694b26ac
z8edbec1fd599914e6e1f6a97fa34fc26ae0693d446622bce0bf852880b6df902f72dd54cb8d2f7
zf8f4422722ae503a043eae02470404fbbf821bce78326ed302e0e6abc4c547ddf2158771426e7b
zdb2057f464ae8b74df77cf304fb6d9c35449c92230ae70ae20ec2546bcca60baf0b5b59fd210c0
z15edeee4df042b807e860f154a71622bb619ccf0738f7d871085eb6ce3dde96b51aadf3ca3cf47
z0f25db0af5c119e2afefdce97ad9b1b0d781e7ee6a709d40c38fc29d5ac3671e5a9f6722792e00
z4a6380704203d16a1ba88dddb1b6ef76902e412d3f320d40573e7fd21dd5d0400bb34e96159ade
z7634845607527d2798b78ab36664766aa5cdff877846f504710c79be0e5afac4da8704feeb62e2
z617242de89a907887982e798232346416644436e120b5328f65a75cd1d7d6f00e7b1152d8b9749
zfd500be5b7252ae37e0ff16b8cf35f34890ea38b1884156aad0a3c1a41ef443e1742a52d73bd31
zb6489ba8768278b7951dfb2dcbd2282f7b027085ec6e0515fa8abcec7ed0f11e2959583cd4d885
za13424b6d3713e2d998ca8d054a92ad78b18b055474eb210dd7592ccbdca4d885853657e27aad3
zf83a513c8ebb92c8c83164af53126fc9777ec13dfbbc602ec911949b538a1a0fbd1648f55c573c
zc43a811fdbd3b62ba2634a836965560219efd288a98974f9f1fc0b4f7b5bdabcff78e750ea2eb2
z0084c40dca65b0bac45cfd7402d61c6d0f9613533dd2afd1625355d4ee44665e79ed4d32b40de7
zd7b1d0c5339e768d8fff5078ba87a8cddd58b53f541ff7689682ae77d841897585a42aa8cf4e6a
z7f395a82b808486fdef4159ec44a0dbb89897fe70f117de7e1d16e483ff77d04a55c796b22c778
z5f6c7a40af24406609db3e4e245431fb79a723c92ddab409bf40dd51b6b631c8ad335a8fff0424
z91015a0a7d6a88efc9526b09a93dbe3738a8f04aeda3cedbae9edda5a92589a8f2e6c026868a7d
zfc22a32d1a70f1664f36f5e83e1932942fcd09321c6d0774e3aa945d197cb60276641bcfc3aae3
z0361740cf9c6c94fa3dffedd15e2ce9d5e81909dce2df8d579b0fc7ad60a2db8da4f6232b99291
z1b9822025cfd94018c9ea284ea90a1e471cc49da31fac113706cd8d0a7d9b3821afc839ddcecaa
z90d720d67eafacb2a508f6a4b3720e9349173a633f45be1621e4a8b915d39cf209a5560ef2d364
z4e186aeaf0a2a73150538797c4ec149eafc2707d002b26a545c910fcf3525f2ff53053ec99f81c
z1a3ff2f07393b6a2ab991e93971ed28c2ced3245aad5a5b7f2f4f46add2f8f345cf26d3cd23901
z1e5ae975e5463311a67d6fd6bbde890d1d488b7d0e13b0ffd88986fb29d9781e060fb1ef5ca080
zeadf960d32a51599aa3faa2daada3942f11e6f99dd5a25df168119988a7ea4d329df777bc9e915
z6c42e467e0f478e43eab02620377831679054f8fa7fffda20eeefd0675e66af2e58b86a27280f8
zf8284de8ad41ce820d1d52acfec433eee2cf4eef2de35fc1803dfc480551eb487cbdeee9f3995b
z25997d63ae184eb58f4929555dfa68fbe769625714769d09cd4f1afed53e8984de371d1c3ac540
ze3e2e3e515a8656aed054720fa2e8e2007214359ab91f29ca697a36a45a1f8d5fcdf61ad8b4d96
z67dcf04a47162a3fdf4d37a149c11e15226307be8fe8c009b17040f703f3aa80fa9d5e7eb15b67
zdd3c0ce46082fa39b3d1411c41feb27dfc75ba72b1b06bb6ee499c2410266046e9199ddbb4681a
z04d470f4a2ddf0ce991663a91c612eca82d1088f67e6a16e1af1f4c938b92c38d08c43b597b8a2
zcf62abb49541897417bf61315af0c4841f32042ff15d6d17d143ae4ea2a1b330f42f9e6a47e0e2
zf4818dd4c8084629937c215b71015b125ab753b81bb84310542cba8fe7ca3d5f6b9c343849b68a
z1441bdeee08540285934538a5c6c5746d2cb81818534ceed9d6e498b72256673d288fe28abe8e7
z2e46cbacb791d655eb1ed10cb79e32b77978ad962fc3b5846f6986720f6de5121de724c7e20229
z44f920751b35ed416e99bd5d3b052d7f1b4442b41e3e8956980040b3fe3093e24369766e23aa52
zb588ca992e2acbec9294dca05ac55feb30d0c2b819fa682ea62451f6602735699c6958f68b25ef
zbe78a681fef76728c0d15b939c952f4cb7eb98d90c0bed2cfcaea837f5022aa2d5244bdebec6d2
z2552ee98eee282a3e21e58b055ae5632cdac57ce41d42ae5a540411c3a0e271c2b8518be408c49
zfe208e6f9999e517b6057fd875aee3702bc8016b04fc5888b0bb525e0c90732517de96b4672fa5
z69db6525b717a39f95eb057868571cf5ec251830c4c24241c4f59be5ea701224b7c8ae8407bf70
z6487ce325a06810f992248710b608cc9fc064cf6b930b1e73dd24f3c91eeaf4a945c574a0bd7c3
zc60c6b60c4fd2b3de74e70cd7c1557c31f1b3051edd55f4e77f7024719733f424027c4564b0fbb
zdc9c99c248594fdbcb6f7f1d68346ce8605506788db696151b09f004808799d5152bba80538e6f
z906cc2b0aaacdc12081cd67c79e2b1d00de2c43fddcb4def5d368f445e4591125c65df69af070c
zf730f179b743ee1b8e10d79149aa69e11f11262a4f2b73c44e7d4bfb1d35ee6bf2d060f2b71366
z16f91391c44e1adf5d497e01b820261c9ddef2d985bedfa5898cedf381c7438a4ea095cbdfc32f
z461e38d4b243059c7fbcd8d73b9da095ea336ca0b2011ff7495c56738c1e4f066d44f2c2435a62
za47b601be8e4478eaea56dd81429d1e3c22fe9d0af5f3e7e911ec67caf683e8fee287586e27b3d
zfb44f749a0920c26bccac98058fb96fa4a0f92fd7d0baf24725723daede44aa8b59b111b024eb1
zf5c2ee5a01a37a1598e3c75eb2f7cdfc365c0545f62f12f0e75bf20b54c135a33d14131fdb7318
z6023fce0a061a433f23c216c6d6fab42d5606035bc5fce5afed56f33b624af652959c557e92195
z5981039690380b8711ad97bb46fe5b762babccedcb71e252ff1b06d71b0be2b557552a56603968
zc0cb8cc1019e2aa6f404b0bcea6a552eb72f435cffeacbb85e3c2a814115ba2b3785cc9fa71cfb
z0aa8c9ff7bba206b4b9323f22de3f5cd1e2b49683a6866d06107f75d86006c968aad0da8a43c7f
zb2e7452bbd49dc63a9e662de0e63828ce37be2f6c5f8af9311954596d4da3706ac3d3755aba72b
zf881cdd54f9248acfb419df44fb247762066c9c96b9b7284362e3378c6b54f904bd9f7c990da4f
z0f83744cde58757603464b9bef9bdd011a8d1e503961e37a240e9ba3ff1041de5373974ce93b33
z09f14d5ff2413d98b85cb7d5318559130d089158fb1aa6679cd647f7db5023a9b5ed6e8afa97b9
zd4df5adf7bc9bae97411f27fa31de07236f2dbfed4a2bf090a924f88a27e3cbde7f5611ce9eb2d
z7fb0f67f4df92506957219e747c6e67869512ee6198f2549c332c2d29462df0c5327b08fae3030
za364bfc428711f11931889fc6bde560ee8852775673ef8b71e758125d22f804939773472f685e8
z9f53159184842f04f52fea3550b7c7b4cbfd86b62dbca7a29880fd92f5b275778123bde3c9848f
z494c6e42b81955bd1068ee72069548b5dd21d26de759fdb6283645d44346eb01115e5349fcd302
zc11369bddd1b3fdcdf8d0b792e97d8404fe16863f06100900b8f15073b8c003e494816da479471
zc87114e0de2537201c5c38c8c47dcecceceace1c8a104226d20c1bee59fde7d9aacbef041e7dbd
zfce700c911d12ad9da428fa86e24c8c10c3cb54b5953797a054b308494c57e47cba465cf3a600d
zbb1c3239c42a9e95c62acff8f20736b67059ee00a41500014756c32b150d3e1f98cc7f4ffdee1c
z02a49343745664c3a6cb39adea92c38f85d2b3274f272758bbaff5b4e4292141924c6eb957628b
zfdf9191239dfc52cd146ec6fdbf575c7096ed84d761b3264881e0875afd643f35fb8ddc91ebc14
z315d40775e2a907dfb516c69030f85bf5703c1d457ea7080c82429441e503f77a9f22cd59c85af
z18cff5a68bcc708fc067041bfc68dd3491a11ee66b362605f8b794fa92d7aa067e225cd1c34a96
z08b36790fcf5b625907e740cab3a6af042c1ac236962e2068556e53efc3e8f9ec671964e93b0c0
z1a5e7a00595b9683d8e5afde3ebf4255da198bb64cf3c65d0742c8d4cf66f8445646dc76f93e0d
z7a887494a6f0e388513a028098f40b5dbf1ac2f11aa18b7c8fc11a8ae20a5230807664ab02240b
z1a393dd8a3c3bd2ca4ec25ca527baabc976b23017c82ee67f92c5a5198e72a4ea85e2eadf9e533
zde1db831bda1b9f39f87281e20993f0ed26431b14712b7211d96dae8f6533f39d984b0f918c3eb
zf80e80384642bb08194f8102f815a36b20c8183bab889888c3961593586ce8d5250f40d2379cda
zb7cbe5298e2ce53874b8e936425ec8500eaba138d9187dd614fa5b7038c4e921fbd5395aa8a816
zc72057a62bde8ef45618b4e41c69dcb0c5172d35811735b6aa0c11f1699f3ded18cc3e65645db8
ze9f5a167d196858b735d07ddeef9df56bea5d73428444466f87886b9ece3fb8c09117c48e72d6a
z52c82d66e4ef59d88fa98082ad4e400857e7c1c5f96ff106e185fc83eaf1f1a11825637d794931
zc8bd56d1ef30e995acc715270b43f9af5ef03c984310eff23be17ad0d69ae17760d73686866cbd
z72d96bcad8205a1c927284760f46150df2cc0880101563d6e145b435f9eb19ef4744636b9d467b
zd2addba1209a9b9e578d118aa926c506869d6d909d95a71eb229a6d5fa69ec35ee4e8da65b4a07
z2acd4ad7278344df7e58a72fed29c7cc0846bceb6a40220928c6d9a79b86e4a40391695cbede89
z4fca3c5a23dd1f8aaa6858a7786c7efc60bab5d77ecafbe93c0d00efd421d9edcacf8138b483f8
zcd6d0ba659f73bf4f423fe484f41a619f5e5abf3d15ed1ebefec3b368c7293a88406e8216e9d0a
zded384f18f128e2d95d738a8a07fe9cb9e23ca494bceff35153cb5f1fd086a7443a20bbdb59039
z794bb0d61af097b9ea8a722d11a6542eb4e8b633a143900b6d9a0a242312e751a71c8842468f28
z7f527297f665355012465454291276b9554c6d7b905e7d436ff7fbccbd2483267b19ee0a375afc
z736ef14adb1e2e175577177d048cc6e60425eb5db7433e1b22663a339ff1af97481330799c4e1d
z2231ffca1594ef0b3484379d3d3b79b79283f671f6ea38774bdea453bc24d923767a3ee276bbcd
z17decfbc54be39745d1ec9f7e2d21e9c36e4f9046ce79737d93eac0a24badb872d44f00224b04c
za8b3118cde545f30ec21840cb6511c252f149ad8f29fa433a5a95f887f4ba469ceb54195d7a9c1
zb57efe7a23c349e28d9a30e9eb7ba0e83706bd6eafcf2bcd933fed88181c8d5dd5477cee5a8a47
z02e9ee20b6f2daca4f8b10f8d9eaacbda7a8a7c8947502e067a611e3e562e45cb9ffb253729ead
zbbf1407b2a3e9898a6463dc71c095bfa8ef11648842971669760f394b0865f35b16d6d36ce122f
z19ff211f4e5cbac8c1cd82ca4eda1fcfad875b2ed389afd9308198f54897bc59b4e2e7539b6bd1
zdecc8d2050118f68ffa2268dba0ce283b6ae591e8bdaa3acdb1936c98524ceab6f2c34c5484331
z04c90e5d4820d186ba490cd9d489e1412eb60225951f1fb964faaa371c92a87f59a3318349a194
z94ac9bf0b7909cd817ac2e838a94fc1fcf19532ebd5c6634ddd0d14e2de59a79c0178446b49496
z1f6c7e059d25caa672a59a10006946af53eae75281b4265d7ef52901c3c06be0107d27e0fb2e79
z4d0cf6c35909440855b746ac69e6e3293a4a480ee6eafb84c5c1e251e34f698a739594b3796df1
zfaa927c472a186e7fe4de0de148cd172a047ed6aa3905c00ae3f04ce80cf14eaecc594962b7ef3
zb3ad7ceaa6ef92181c4909356bbe468bf11894961f7f43119ff6974e66ae16b838eb60a268ecc0
z05f26ca41b221d9742dc9abf7590ba9867103f92ad4e9e645d41518d0af2771a90c26dea37ec29
z8d47793202250a772cc4f873d97118bc7cde295c27eaafd8575e9a29bc727c72b2104d56dbafc8
zac7a454f2cb92a50c475d2e196e2079c97b9bd587028d6b88d45a923ec10e7904cda3fc5dcc824
z26c7f04d60a6c1b5c2726087a270b8e6307bed96aa323e4e85e42c7b2f1a790ad747d7dbf0f8ef
z951011ddc2d3a758a10ac03987da7e4ae4d8a0f3d4a1e5a4117d4481bf48841a3c505ba81d9a0a
ze15e5ce038415b81fbb8b06a19207dfffc7d80659fb0308b7576a6cc710fe609a5b2eef7c70191
zf232ece96f7745d1c898c01803cb50e99089483a2fd1114dc242a623070148b858664b83a11abb
z4d0c5d6aa4d34e028e0d6933c2cbc33d2141af2150078c5f8731d85c5c2188c89248c9c21cbbef
z1d7468f6ea9529227248ba85815aa729940c355a6a1438a4255625ef5046ba952b7760e5e7b72c
z4d384632d307f01fe6be3a04a44a24f3f4d746496a3894d80a7c449fd6d8f2f33ab16b61895d1f
zf925654cd1b7e29dbd3185f63ec6aa34a18aea974569ad6029ee4e4f00b65535f1d25860d91699
z500255c8993c2e22a2b1d014013f5a3a63f283fae0bf17251d216a2c6d0d75a4474bfdfdb89f78
z33d33750fc3ad4e793dfe655fe1d0a792271cf5c3cab4d073f6ee768ff16b1ae7a76a7bb361fe1
za01836568dce0ff2c4204055c1cf996325c77272ba72ce1d9a9496e9c460480d8d688e93d90eb5
zcc3fba25222074cf68c17a3f610e8f52fc7b098630a5438796d6491ba3374495aa416c2e10aa38
z4674289cdbc1382d3c9fdc7b23a06fb06c6cc3b27c5160299502494bf11d355c5499518fe2801c
za23b538deb2758be6f6f54e7229c883f5c63908b01a881c1bce9e0edc6119acb4887fadb69cc10
zec485a6e14cde952a9ee042093a5fcb4f84057e7b322dc0296c3374f92531e230c1273256219f4
za8b2aecf94689d70081b9cfbb650976a765caaba26cd9317a00b56a767e890c0d716714350be78
zd9dbfebb59bcaca442ac090682b1a83eb7479883bce015e3c08096a59a27d1d59225bb9aae68ca
z11e94ed1f10e07cf2c101caa9b3ac19cc50b82175beb6f2454e9d27088020f3bf954599f23165f
z7e2eb3b02c4c4d70eb58555931b57986ccad89b4934573449a822eac5151d4f01c1ac5b109cf74
z6a203662d724312ebaffc80cbb4e0229dfdbbc77991887616756451041005dc931f16107ad21ad
z59ae0061ae13aae10075f937c97a23059fbea5c0ca265c7c85247090d243645e3b245d4cb6aa0a
zc71f30d706694e087ffc15a80906823860ed157ed61b771f938a2f77cf240ef4ea9cb6a39f359e
zd7c4b786c21174ca24577ec5e62915582e9957290c913e7bf339b22d8a4a3eb1c00fd087daf401
z1a9cdc52270b4949d5d8f230c2d4107f5f681bda8a824e32623ceb397e0194f4f46cf2df7948ea
ze2f505e020beaec60d095dd27ae037eed48cafa4017191beaf7ba0659ce4286fd077d65b48b617
zc6f9c9837976c1a0f84b0027593e0d6b6ede104b10061104b1750530444c8b6fda836732abd561
z17fbae55ab277dafcceaeb30b44f9c75e4ea6fab6cf691eabb56dd0ee7e497160a3b5cd7d4e295
z10a1fecf44205d2f0e1d56b9b0e324f98f85a32fb574c94d61ba6a9b49eced17a194b6799c0b1a
z73cff44b7e8171a075a32b4781a2b9c9f356279073b43702a8be63b767be526fc277025e250add
z1570fd0310efa67dfdeaf8138cc7526d0702c81a2e570e27a724a2b94c050a42118a9cb5bbaba2
z13b9472de809529cf30c80e510ba2ef88a671da807934062deea02b08a546f3ae688c9659806d8
zec846c865f8ab3dbd84e04ffd408ba216c70411274c179879386d2ad34f4839909169fd4f7c52d
z5f61a8e04eefa88e57a553e3e90743cb77f7245283ee6cb272ea3c4d864a9e594afd7443af0474
z52bdc016dafe9083d7e42d44c0f42966862e6428b74322d150c9229998505539c44755afee4580
z57fb5586fb900c1b95d5a41b3e30844e883ec446099cb573ba59be93ade45edc9760a85c66e73a
zf792fea68048d421adfd0245862199c0a004f10ae87cbe1789a9a85a5be813532bea798e063158
z89ddc9132ec5328f65611b3877261675e129a4e95d68fcb157fce6496bbe3d034c0d48ef782d25
z0378ed2f40c22279a09a1ece40e97dfd0d0f3a91055e1f930305e32f7fece4bd4bdd2b8aeba56c
z26e98b1f00fb35ed0ded7b49914bab25217e25af532cbf8f07135108b5b30a59911b0ea04eb288
z69251500eb19639f8eabb359629c60f4b930e487dccd1cf2e95432fcb777ea427ec11090b619f9
z217c3dfe03a350411d1bde77b104b7135cae9cd51db662a29894c8f430aa7188eb631d4ed34da2
zf3f7bd831a788ffffe951cb67c7aab752b88dc629f3001c518c48860ce02530b7bf975167ae4ab
z32fb9a71f488472f3591a6695070dc77aa79cb5b16e5dd46e6f5c720212f1a55d9b8305f65b568
z481a353de2567a0f39be275c3f31dcda619523526c80fdc3bf16398fab7781ccc613195989cf25
z2a774af77c99b89eeae91fcc282661a60411218b30be7e7b1d24a7624285ce19c32e56541d0fe1
z8b07c20b54d44bda9d8f5b28473d38547e8ae675fc7103d857acc7dc3ba0cc7231783791a4a5b7
zeb947640da816be8c92b1c816d79d3a542fc350feb7da72ffd1234636232fada85b8dda859fae7
z024ba81c5614ffea08dde58e63be323a2e519ce2140e79fbe892864cbc033df7b5c327a79545d7
zb60abc2f54e7608bce46421d7cfde2cc33d3e40fb464e85b9ec954a43ee238834a739ac7e95555
ze21fc43023f2d1a19ae9fe30b335a186cdc96c428887e40cc02c2e6286a259607509ff22148c44
z54c7b5695ed871b13b8bd6ae033566d9fd3bbaaebb71e789ee310bda5dafc7dafe4dde7100da84
z36f83ed5afd90da9ca190d45d979ad4392f0f002d8ed834dd00580736a3997e3262bf45348ace9
z364e16754b62a9e024191042dbe2d6f86dc0115b470d9d849a6c69f6e4032807ed8e7107a92d52
ze8e970989da47c0ea4b1ec1a2c9fe452fcb0f9046057c7717a101b6281ddb35b52cb6031d1ab5d
zd119c563af7f3d9f5fafda2fabbeedaa448f6aa7d486d21225395f21f0db11f765efde95524733
z29587da73bf40592505b211a3cb877147773e982ff6102b65c89ea77dd403b8f297ff588e26594
z6642869302b2573ce1f1dbefdc2fe5e0e82624fe11904a146acedf3946f5ede500eec4034d430d
z92c54943e22fe3b0d225870f441c341352764997133e2e58de932924a9aae2b44e9caa6c7efb4c
z9cc47ad6c9e9339b55d46f72957ffd9d46301f8ac781c4f45908b99f97aac562c385378e50651d
z3ecab954b03ed0cf79942e3c1b3333396dd09ab637fb3e757307509cb20c889f0e621619399b8b
z1c66a88c357874511bcda34cef485afc2c658532d7df2b59328ad06c96411a82cc8930d0c8a1bc
z4ec97c18152f82062316f6755949fdf784ddb11a78f0c189465f97f6a156e234409aff836c3747
z2ee76fe9c97fbdae3d1929bd1cdfb6c7dc5a1d75d910e6ee494480c81151c4fc81377eda12f33c
z08471203550438c739b3c6449d22f546f0ab913f23e3ce05463785773c6e2f3372d42f3a666a3d
z10b443d3deb7106146a241909e5f4412af50117d2614694c4054151419569f7a0253315dc3ed86
z52f71edb0e507e049634c1363a142c2bada477e40a9b0ead1a8b8f8a8aac92fd8c3faa7d0a75e2
zd05d38a30f61e5bba6594f19f453a744526725a55d93f88542d907cc84add4b642f2062ce62e45
z6652ae3a72c9039b6552ca185c7879562d99e9276826ac798c1c5aee95aef83452ea92b7e32bfe
z594cd622f6838ae5eecadabfd296f7afeee15a1c539a9a974716c38fbde3860c47887ba464ac9d
zd3c9dbefd0d6645a467628da98ca8e29463007ce34ddc8657d60017cef7a2fa497e151d8a69fd3
z334a83516d345f4d2ea9fd790090df4fe6090237758690f7d0281459ffd326c76f9c8b4610c2ef
z755bd3fcdfe363dc9eebeae2f303a8503f0078dfa499987f86f01bb7894515bb9acbb717bfc002
z7617c3a0dbdc496e32517ac5841ffa080d6f5d34f464c9ef4af41b4e50acb8c3d83ff1d33a0d5d
z96aa16e3e13adc1b21cb4c8afbe414e683703efc0c1b696de2f6d6000c24c94a452ff7b7fef775
z7cce186eae45cb86993be0a04c72a99cb6ee4a98ab3554148efd6ac4f24b3d89faf1182c345223
z09443c899eae74caa3306ddb41a0297f2b0e695346fd083ac3cc965fc95f7af3b35858ba7283e5
z5e0270d209495d2f5070bb2f0542a60bafed965423c217ef26e751db6db405ce1caa4569e37cf1
zd2e8d26c5d58ecc7706f7125e23ab89813f4633b23caf113abfbfa32ae50c7fddc432c09b228c6
z43ad4e915d8bcc93462e1a2272c533d9047e6a4a7977daa749213f795a6203050727bd04687508
z4cf9a484eeef99b2eca347ee073c6f8572c228ad6930c229a850bb90f53e4061915790e36b3956
zd304a832a606b52d96747a4153045bf17d2e1a9f1dd36072d2a4c39c67256e997404e74a9950a4
zc8d64eb20e29ba68df68081437456353b34ebeebc15af1aa2c7680c0df08a1efcf26ad7a8a3897
z4bc1d13f359bc9dcedee09c922aa3f38cb9d013d00a6060fbed9b496edf363361295c1b3c88ceb
z6be557e9de5edfb35b6274a175256714c4b73b170fcca9df731a3c297491db50fa045bfc97c685
zfb812e9853c8960a5d62818154a2d44cd78df57d793363cc6476cdc6e324d80fa35aaa72dbc7b3
z563e0e14af331b994ca26723e923eff4d553782f9e97535e2ec90428373d44aee0990277b1296a
z5ee548c0669153b8edc44540dc3624894b625e45f2dd467b8ebe542305dbb8b06436dff80faa84
z2bc2f3ffb04c7e69ddd047306b3d08c9d548f1f506fc3e7ed4d8a4dd1044984900b78c81293aa9
z133975f4bb2661a7c7812affb06d1baafc54ae0943b24c85bdab6e77994afd699c5d532c49f843
z7f7306113d450fd25e19e72b077c2fe5cabd5ca86bfc5db8eb636e23460e4e1325f7fe2353f027
z9eb5e5a98dba3ee367be1c3208e962ac25889f6c6ea1dd7dc3468ceb5d671182d12bf1e8bd0290
zbd705b9d1c12e1638eee1a445aea15bfd6abbdee0565f54899b37da8c9682656072dd539fc892c
zbbd6544a39a266a47dd17c15cecf369c6b54871d51e4b458794998805181eb860b5fea1a819aff
z1bd4f1223fc3bc67a6e5930329d4bb1fdd3de848e1df31f79793d9a1069202c806e0beba3455b3
z02324e92aa23ba248b30f0cb28a5234727eea0e5af65f76aa495da7b3b401ff7fef04bb99f0090
ze5c0da9a5fabbcf7bd798d8d787abaf41d671565d67db42bafeff75445c6ce467bcd06bd49df01
z6bfc22cf76d508bf9eef4858f011d076cc443862471c942d1dc57f953ccdbacd992d80ce033e8c
za06e55e17d63a6696d067322ebda7f6a7665c2426ca1ba65d11d5d86c17944e681027729adb40d
z71d45098137655bf84b4761eea97c8107d90fa1e862588816c5ce37453529549f5d4557b57cec8
z08c37519d4f15d082d30e387392c1ef27b626e5f1860d008e083acf87f19f371be06234b83868a
z388f16e3d7fd23c3c56fce8d1b749e0b3d2528c31efbe2173e8f9d41fcb55165bc7f140f38e1ee
z143c4781755fe84df0eef4bf365dca32f6e6b785a0bf20ee701691f0c609f6061fe24a1e0e9180
z4f687940c546a7735243b16cce4c662b8d91d95f9daffa708ec5bc35722f72b6e188c0450edf09
zfeca7c02befaeb378ffcdd67690fbefc55de1f2b89616e0694da4b536496c433931aedbe9a2f25
z2bd83e12583874b31d145a8d80fb37943661e4f247e893849c03800be4a8d8aef2561c2e6fcdab
z1f8d9e41fee36303372eaf12c47ccf02fb7cee0512dbccdce58380f3e0d1d6690eece944e4b455
z27f0ed6115425b45454d936ecb9ed9f4e59b80a4758c471b4acbfe4b54707cb0cc9df41fc2e538
z8763bb2c281d41592c5923176066103071ad3a731be59ebcb92b5d60b5cad5ff38f39cc9eed361
z5cc1cec206a39f7bb54c4e7f404c7f04ae1683a9b0184d790a144052ec2a9714d56e2f31000cfe
z4dcc6455b0dc65401c41114e81bb32d51b7a1af590e472298bcc02b3dc306794402433f27777b1
zb46a0a0034bc1e1971f4bf4fe60805e7e845d3a74063b37e19bb8465ec66da70f2d96478785b37
zbc33f8a895da80a7978763167d01781aa8d151d5c24172f689e202674efc47565c06dfc8b155ed
za7b80064e33f87c785531b95173db40c121b44b2964a6e2941d4863ba728bcc5bc3ee959fed3fe
z53f658fdecfd368d19cd2f6c44d557bafd933634975cd6b4f2aa0947635927ef5128a93cfe3adf
z824c2499362a9ee9198c479476489839c9f7f408df4b6cecdb92168e87943162809f83823b437b
z3b1ed0a408b65d9301bd00f4db762271fb496e16dc1b1f01558a5b39d8c007e8e7f68570889cd6
z26a5a6ce22c99007907519d724f6c7e1ca7a3058e050871fb9bf6a27f346280296a60078adb8b0
za08a312665ccc0240b6876d043b36eada9aa33f29510e4e4fb0b377b83cdb64e155c26f887b23d
za1a1f54c33ec4be2749e5121fe70b38fcf3fccb1df298755849309b8117ae81b283d4d630e4d4e
zfed2b548f4223fa0b202082aa5ee5bfa06e6739f6e5eaa2dfb85b26a97b9b391533c333bdb7fc2
z9fcdac5487f9cb2e3e7efd7c0fedfe3d9088fc21ee8ef999886dea7d40d6e392d108797e244506
zeec6965bd1025910470ab0695c046e1fe7d881f5c1bc817a7a77a3ff037e3b3033ebcf326df197
z1a790d41c59e32a245ca99801579002c9f9dcb0f3d60757455ae50bb24206c215abade6c8e4768
z92b58f722901ae2b1f423dccde09a2aa86e0ff8c059a44b9fd111527f9755c93f2b57bdbfd3165
za092d40f08fe57f298e795a855c429890fe4323d9bb006bd947225482c3de05a8f7ed7ddf4b724
z84a0508648be49d1acd909683798060bc9bd0f2700492ef541c2f6843d3538a04d0d8274217873
zcccb8c98970c31ebc57ee6f72eb6f90a63cce5ca487fe6ab4e50f110f82f94b0e76c90b0624deb
z1b4a7d7d56574a4c0dd847614ebcae91a9d16ebf5255d90f595a341bd2d9e149470e4e68cd0137
z53cc21f1f7588e5956ab76e3238612e01187a771bd3331b3060b5d0e515fc5b957fe178f421724
zd4972f557ae99bbe9ecc426fa57d5f17a34691ba54cc8b88fe2c41d7adf10d08b0196d65cc1a0a
zf7058c313b8234931a12fa92ccbfc3e398a02ff1d407e51c3209ceea00436e302fb56b4146bb0c
ze7af81759fabaf3eb46da91edfc3c535c015da7d7a514ec4a318fa9cb44875f2d2f36127334948
z4a5f22f0da08a7530bdc4bed2cecd2e67f8274f185366d937e799a2645a035bb6126772d5b1885
z92df1ba75839300be7151a8d5030be661f12d7b0f523d004192fa5c2f1754ae718d0328606a225
z21b383a602049b0cb591934b8b1d6096f8ddbfa0596ac9366e84a290bbf69f2c5a0ed99406029c
zbfff345734e8504035963712313e76317fdc246619e7dee6209a59f7259904bf61c3e5a5bc16d8
z44182b5356382ac952828ccca15ef34c920937d22dc1acac2bb7febe4eea7a9d731b0e909068f7
z9a9dded1c19768f350c83898ac6b687b0c42e416a9af9efdff3e460bfc3a150ebe9ec95c16e635
z2d673a577792f6a15506af55ba424810e5dbd223af29d30ea02a528c6d13fdf99abb14dfc4fb66
ze86441376627fb9c5234bf5622f6a6691f7ec96a3fce570787d529c06593f22dcfe4d9592821a9
za4371ae1b8583e679d4c3ce0655b75b1757a076011035f30d88b6296b3cc25f3ef1f1d179df540
zf14c0c5ffc2cfe78c73cd0ba4503e24f71444200001e5935b293b0dead277385946a2f91b416e5
zcb01e30ef5cd9bd041c1c49c0d77e8328f1d1bbd2096994483022c86eddfd20674e4b2842a8acb
zad057f45508385380aa940ec69e70e5b0ec2ed76e5962b60f177d274b1516352341f170f189cba
zec6a6e1a10d952a285901377de1b25bcf0bacd51227758f58bb8c8ae818461d040bfb8f57f0644
za15bd5e9797162a0714bfd6719872452d983ed9522631611d86e7b00116ad8c7848a4f53f72cc8
zd350c5187af92e2d38add1eca24c151091e978b4d8d7e098be611977cef913e6c6f8c62be015ba
z72ced687bbb497430a0899c705dd4121f9b34d266f386fd5e5adcaee8691cfe4da547563318138
z8765f68956e80066b6c2df164343dd23703ace788f7179c4ee17cbb79314865da9e1668b4a1c06
z28eb1d62f8928e8d972a4e309c7ed5dc74b21acb93b23ab634aa262b69502890b74df0616899f2
zdbfff85a722c54e4ae64f8aa19e2e67a2fa4086d2096a1246635026434946da742d8feabda53bb
z07e058ecb59c9721862ee6757f38739e3e37dccc330b13802ff3517a11128c3916a81bc1d47f48
z8df1ea1a600b54d5ebe78d592100c083162e6eb07a2cf589db812d2dcf88e11b7060e2b5d07c96
z2cfee44fdca74af0c62f2f7b4f7cf37570117ac16a6eddb32948ef181cfcfadd957e0b0bf4a830
zb8780c8e9540daa0e9560a2d3a3c05b30ca1cf5c568e6b4fffa830bd80b4be27c7ef4a97b85b1f
z4fbb44e772ff768902a735ec105447c7aeeb40901349dd289f90b20e00e81900b1080d06b05623
z53cab727dcf9afa7fc897e9b78c97aaa1c8d030702cd5cdd780e179553f5f30a67c223221c659f
z1b3f18342fd4413dccb37d435b1a3b689b6c5e8ca0ebf5cae8c38717ab8aa39a8bbd7262097c51
z8c5e54819719eba0f4bec25c05080587f604c5d17000807cbb19ad0f05210b813b490d5fcf72c1
z77acd086102e8ea432656ddf76c2a9d3e6ca2dba893de28ddca177eb707f952441597778397c60
z0292edb857b750330907623219ea198afb8dc3bb4d5bf5cb9d780c5d2d44704f1321e57d93cb07
ze3bb951ca4d0550930b65f19f2ef35e43e5e87a4efeda7aed8e4b51cc4e1ec6508d1c563877068
ze514e2d5973ad4223366f9d3f1c818b26e8a8f413d87fea2e6cc128a0dc8da1555315fd4ebb822
z6ab89512fd7128f6702b6220251c054e4650a0601ab766f2b110a6ee93e6fc2d89dd3c4567dbe5
z2764b48a0860f9138c600305603e44c40f18e9999d4bea3abd102a539c0cb012503afb82555591
z5f96807cb43385d879b06f06654d5d328d219e866a693b1922252f857ab9076e10f4c58c84ee8d
zfc9fa74e0cfd72703d5f33e5f05445da8a7f1c09e2ec6b20bae62e5ee3f114a9ead11dcaac9a16
z24476fb284d65342b8561578c3aa11e905c60a0092523ef143759f4feabb2c71e5fa17ea472888
za09423f7eb2d153ed9c3bc1561d2b2d610dc75b596e6994826ab0090ae7f9f71d476bd046cc6d0
z981138dacf28de88f2a245045cded2b1c2ecf7871abf16201b0c96cb2302beee14172d8770b035
z921bfc2e57db5b05298716ac043535efaeb2adc303c0ca7e16757039c53a5b128db8104adbafeb
z480279e1689051a53082b6e0250647d7008831280ef82acd64f7ac0c42609f097f4314ca752464
z337443fc01b7d17206680eb0c80bb4c901a6a57d0893ebbab065a844dcb74e78cc3a26aa088c45
z20f58ceaafc3cbb0788fcd0146493fc42b4ddfc1b65a7313fdbb0c390e37cb507cc187a7c3cdcd
z2e91233695fbf30ca5e3d803ffe714898d3f6babbfb9730009420313334a89e64464c475805f41
z7e61cbd51f4bcb02c12dc5a8a192b9175954a283a0cfd76ce8a06d586b99fa292b22804325407d
z1af367209f01461c2ec5a0162e01cbbfcce18084c30437d96eaa34e4bd393da56dee1325699f44
zb3b1f40f8c2b3db57d4c864a0a3921d9c90879c7c8156bdc5587169853e8835a23c37d987c095a
z1955a49034621ee630c9f1a9b11d7d56155bfa72cdfab8ccf8972809d455260340dbce45200a8b
ze6b858ebbdd2d52b3b71ae54e1b9016a7a1c58825e8ebd397f16ba34c5218631c7f5b319502118
zf2bf292fb69f4a1afd34c49dc6ea8c6e315ac30ae9092b101a9a7a1009cad27006006ca2aba296
z6a3606dda1e43274993f01dbc9d7c9c0e5d82d25281e360647796a670be9db048918a96b895c7d
zf4b6fe3d9d6afd9d7a17ecd31b055642ee6947c734afb981b8d78056131054d79c678d16690003
z534641546e9e6481f093f1d56c75125a65088c4352ef416e4989d6f4f08d1a1d92b221a051294a
z9ccce8128a6f39ab0c841f20d41cce5f960ac98e07e53ab5d12b22211b211a76e5f050bc81d796
z193ff3bd9907f2cbe17fea098e6f2cb9a010daaf79e1d55bf2e44e8749f769b967226561fcc7e5
z083f757a30d54ddbb808263bfe3cb1e0a4254ebed701571e8be85ab8b812d972707e171394e1b5
zfcc6cb5cdddec1e7e2d865bc9df4cec318e389f5fb5bebbee42f5dece697661dd679846586b470
zb468fd4c93346b2bb03aafbe543afd21af259eff6289f38952171e509922583eb171908db77f9f
za8d83fa245d50316ea5403e1a5320c7cd17a5aee85834330c35a8d5643dab8384211a77a98a536
z554a18e746442160e808619061cc85d6b81e1caeca268f0ad7a7b02e56d3a0d69ca12b303db46e
z421258b9b4e464abb3e120031a4dae13cbcc7cc1993f540063e5add9f57375cbb8bbfd64bb9042
z47fcdbab604f7afcf96578e82c538260234a7f670010397a88bf1b2743273d92fc560df6dccc5a
zd770e559909ffdbc65818f7a8e060dc0fc9f9d5a0d1ba31ad432054aaf190475634059e2306642
z5e1f3e7494f29f5e9518ff91078805ac184e83ad82b7fc602476bf3548a2adbab701a26b08a50f
z50244a293dc1fc20bf550ff2dabb6ad857b6c178de60eddaf063034c08e88e80c2236972f868f7
zf2e2ad7522138e9c1dbb430c14f3059163b5761ade24b3ff9942a02fac6e332c0e0a30617975a0
zf64b64c66604e9e96090ff516459ecf622767dbd4958077fb40581bdb9e8792c9c3a9fd279523b
zab7c5ab62ab6506866566ec5b7915183e8a3d45e02041ff7e546b6399305f083bee255f3156882
zc9ae8e9466b438d2eb8b84aebe5a900bc3df200e761e5b32b83043489ffbc8313b2c2adad4678f
z320677b21676043933b824f3c49c5d6a5211946b6b36d71f77b34c7e324ac17931e548493e58b9
z9b2cc5071f38c43c1cb34b07385d188aa1dc62f60a153d6092254beaed4ce2021a62f73a71e47d
zeb8b6dae34e100e53ad4cc7836c1f12c253545146af7a27fce3c8ed81599fe01e552e3d7fefea5
zf0f963aa6bb02eaeb29c0bee9ff7bd174faf35e72c890a18fbfff5e68540a4125087fdf004c411
z588384cda4df0b051591beb809111f601196aa917c370b7107914307a3081a6d78ba31cca3fc29
z27fbae4e42e7ed00148da81b4cdbb31a9bf8133c92c8ec5ef8bdb338cc0ea9771a522a06705ab2
zf13b3ba5b57b5b0239e9c0471561ac470995f506ea819eee79dbe45be8280ea99d715b967a2b19
z0545537e59477a6ae66357186730edf3bbede0730de6fd9ae79b765a2eeb5fdf8bc82cf1d9a5ed
z8665a74c5e33056e999b450c9733420968e77fb8e5efa80ae0fb8ea699facf71e9c551e85212a3
z017e7d822f5ffc8efcac60013c0386495d8fc2ddce3d23e8c8b1bc2ed98ca21f6f205e55917288
z78ad3b8c87c3d5998e85bf9f2371fe29240c7736760df7a4ee402121cde2f31af05f2519f74486
z19f6bbc897050ec3b6eb2114cff1fc65f5e1acfa2f817c3ac88af85b47f77ed546b4384fd482dc
z3d1700c3ebee8dfd5bd4305d93176d2f228db73e88a243f093bec6eb3cfd2d5c7170f28344571d
z387f3d1db480266bd0109f61541d7cc9456babf5cc3290a36329bbe21271220cb88fb5d6486831
z6e8a6415260b3963124fa89a3ca154fe6f1df0684c7daf0d92c46b86ef1faf44439540c3f2eb8e
zae199e01bd3dc95194fde60e444e9d1df38dd7c17bce39810bddd0773ca8213f8b4f668586b42d
zf1e68dfda6ab64da224a41f1ec37b26a269a9a413ea44ad20b91d0c2e1d7329adddd64562c5ca1
zd095a2f840864a18884225b81a9daba59cc5a32c19cb956bc98185aefc128eae0ce9a4d7d04be1
z23bcf7fcc47aacad6c81ede544bbfe1cf400aca823eb524f2bc012014ec785b34864c3d3791065
z83efb5025905e991e5c092e791cdb2ff6438504bf6e67355d316df24a80ec8fe72f5af73b68b40
z6ecdbd35b04f5f93228df9632d3952bde8acbedd35898bc78672fb9dcc5fd0e22c06c210da4fd9
zcdbba622dca720065fe24c9095c68263027214c82f7c81678b1dcfef15426fca19a827888e10a8
z744874847da0ace162bcf823ab9f6edbb5f691c0ba6d38a7106da6fffd7ef62c3078dcfff8e488
z2df4050d8d9837dfbc23dc121e129d0e660f58a2fdff8317bac6fa9656b8e0073ea8e75e5fd4b8
zfd76f9fb0377e0d0b591247a4152fa784968504feb0512103816b74a8bee66508d378f7cc0aa3b
z4bcda4bf1ac1050b5b091d129d700af02729ffb129008e3dd1638351919027ba2ea81ac5ee594f
zaaf48996136345839ba8aaa4b90c00ece3d3504d579fbcc8dd66ad91dd76189c0ed527ed982400
z5f3a011969e479aa3e17690a3cf65b4cd4c0e10e23188d982343f7eb05666414bfaf53b5be475b
zd5915a9ba95c487b0f4581049627d072fcaa6c5de5b902cb43d1ce3c8a66b72ad80efd465cd208
z05c6d41ab247397138e71bd0cedc0820769800ce8def1853ec93f245931c6b93067af7c5a9aacd
zec187b94a46094eb7a6515c9b64a76263b7ccf815d75a5e5017862eccbadf755de3b2199507234
z72cd6bec7c1b98e64f8146f36f2e26cbb0c48458267ccd3c660df439cf7319a79c69731f989e6d
z83bc2fff53277d6b59e1807d2bb3ff925f77ef79b62b1217683978c07863ad3a928d850d34f417
z7c7433fe3cc47e54cd8a697a57a3dcf3fcef715751039788d657a5bc5601fad2219c50320fa901
z89df99c621797b1b2656d29db527a07900e369284438040c3f970313c4ab825a39de3ebdd2f43f
zedd91f8b0c56c084bce0a7b82e0dd9e1ec9513eeb3f25235d0c02cf0edf01b47002e18d2c1324c
z79ff20392fb77592a070a96376b445120d3d57756b51f8f49330e6b145ea6f7df9a350b662348a
z9cce9a574de06707ad31a94a50ebb0e40535102218a80405cb060dfba04e4f829802a4eb2b728a
zb3c92a9d98a76f310585282e78c2c9d8197b5a07c1ef9a7530524438f83c6f97fcced80d352bbc
z24715152ed499683d6f6f29c7313fa21163a3cce1a65d9f6f7bd126d30c3996e2a90b9934b31d7
zc06cdee9e8c7fa420fcb8d78a11adc26d556d7624804ce432c83434fc2c1d99d30327307e7bbb4
z69941f0e525fa2bd1d9a8f0896a6d9bfe5b31d5b3484816e95bd66e47afc3a48324f4c1637c5e9
z541daede133d8b47160e91af638be710a2c1c4417ddf7413983676a1e4b0e48223adf3fbc70202
za772e242ad97aad8b918f5b03798276b91fa1ecac36032642fb782514aef17203fdd00a834df2b
zcd2e39db3fa601074cea2267ebdcb623b391dccb958177d8c563aa3e42bc699d491a0a79a36b92
z9506bb891bd605a0d20ebabf12d3c15dfe7026e1977a067b524b990fbb117b93f74ea55828a076
zfbfc2d9e3f76e7f9e768c778189cfc49f48f93585672e5e6e0b22108c504a6322d0a3e096ab6c9
z43f68d98c6f23fe8cc8cbe9baae366c6bce00190cbb61e79422092780c6640463512084733eb02
z9eb597797dc2201315e1184fc09425b53262360ac09bb3cec273b40093241c4b47a6061cce002c
z45093e16c96bf5f4d556f98a02daa9249e9e5227dfa99a088ea6dc45fd4953c6e94b10d9b24688
z96087995df2ea984135b993b596baec9796198dc90b37f45bca3921e3e888a68ed8cbbddbda7de
zc3ccef1106bb5b2b2270e54a7bb89ba28cb7d07d4e29132e2aab1c486341bbd234a733db7257b1
z94e273664ebe983137adab9a108e30f7f8b48265ba669cf8bc7f2724a61f58062990554a14efa5
z7ccfd068570713e81330b234a3c8303a481b113ab9a0996c1b26d4f8cc8b4cd0acd8f2278aff22
za1ba613a0b19f80888e2ee89e558762b2973655a0e21e85eaf92bee7581bf09ec74c70bcdbbcc8
z1440394ff53bb46f80134e897e99042c667d98196fc90ac66f729003ce39db34ad59de5dbdd3c8
z4bc488bf7ff923804600ed2903179880c95fc56d00f1d588dbcb465a4e3d40003ba08bf8dd43d5
zbdf92b88acff74a4011f70063ddef5af887a9da41fd3e481cce49b8e85c79ff672b68493dd3221
zed282c0b17abc17b8eec6609b4739aee68c600417b24dbacfef330eacece2a99063ccb3f1896e5
z2c1f5d3aa569a48fe1144dc950f12c03b46ac6d4dd1d89c0c747c794836696ad491bbf2b4d304c
z29004c6edaf48275c3e25707cb19d6358f523902be2a139ce7bf9e909d7276430d54c7e3e59ae3
zdb4a1cb7148da8f93088078554128a45325d0a60561c7e76e224ee6c7f7ebc251b9a896832216e
z195b7e4e9f0abc095503a77409c51e0d1d76f6f0e7b3e885c14f9adaf2382ca570f8bb78d430f6
z9d2c03a2b7c0049bd04d090297cd64ca9087d482c2ae6f7b4c23fa477dd583df8b0a5710799a05
z27700dfe80ba77a5afc01d4460d8b2cb3642005c1725eddb83ae684f0dcd5527aa6b59786b52c5
z461a3f8c8acfe326b0e49a8e8663d33dee0854270e9daf38aaa1a845c359c8c2aaee0927119e0f
zb5b9becb3fa025adb4438b534158773fd31bafe4026c242ae81cfbd13f1130af5dddef826406c8
zcda6e6ad95b10f1494b1bad5a67cf5fbd1ee062b471713f423c754d5e6ee318256073025c1c7f7
z675391f4638a129c493a8b81ad3ba3b611c2936b2e8a671dc0d4f5f99a7609c6b57125fb10672d
z3f9c8fe6047915f928267e3b96fedcef6f938472471bdab4207385e25ab07dfef2bfae921e64fc
z4425b70ce2ab654edb4472c70c7aa734c7a6b27c65e5b95b6ae303f4f65e7cc63c29a5c55386df
z71e1e9a0a52c26991309f64c08bd85a86f5637b7f75f62ab9730eacb3f97e4399844370ee72340
z44225dc40128756ba1a7030e50e571091f515f337ea049d6becb041be61609beeb08f4807757fb
z394e18854248d9d6d57e3622d33d5e925e68b66f56ad3064424a4231e6eb0dbe789a8007575554
z7c4e97123f3d5b66df39724415aa9daca53f0a78eade25d65062aea8f977cb796761493a77af53
z59f2133d595229fa117de999519b75d582ce22d9d5acf964fea075cf8d9af2bb247bf8b8f47b5e
z2a3024e90f20c14fb551f0f714a50b7a398932ce90a956c8d3f06a76b4b5dbab4361f399ae3b8a
zee48
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_sas_dynamic_timer_values_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
