`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da33099ba6084c0bafded292dc1
z85dd2e3925edc8b79302536c5a94d857dfab42a4b162c335c207c17b63516c48d4fb6098b4cbe1
z1bab4deb91641b63c1c6e839880afb896158ee4b6eec5adb8df2c114bfd3f7cb263585ce6a864e
zae293f3ac9985727ab847f7a79b7b29fb626d39f45e0ce29ff4021627c694e4ef5c99b33052480
z8015184f0dc497671bf47c11d83ce545041ad326d4311d2d807fb87ee6d058fa5ac515c2ee5318
zca562c1ca11f575425f802d9e52ec735032b5a86bb5a7db41ab5ec1f347a1607d7dcb17bd50450
zab9033e30dacd5e238e3e7a1281ce4a6f699c7e3c9afa79c5fdc746ded6e7d656cbb3f4f2429c9
z27762690787cfcad1928893e7d25f20f58c5c232033c75f373e7a1d68c6ee2ad58f8327aa4432e
z4646672dcd71c503278e37160615aa56398ba0d43fdfea9fd4f9d15e8aa1ac4cf4355fbc7b4335
z4fd6ab2b66839b8b103d329d206410266a8fc22318b1c7bbd4015dfa803622f48fec4fcc7c7cb8
ze9c39c31e012ffb04d7753fdaf3d78d82b495280977b255190cb116c172f202803a25479ed81ee
z1e590cdbaa4a2167b27712dc53800a9b76e91a2fcfaf2acd086fee2bbe0ee456949eacfb03fb38
z9b982c7bc21a9e6510f6fe4bae36848468aec77657f54e0fe96e11aa20b58846380ba7c0d5cdd4
zbcafaf760875c52927b865cf8af8f9de9df431a2663649712e662a7e535697ca2285653404012e
z05901e50fef3cd078f09163ff97659875ae44140f761cb9b6cb800375c7ac3b07f4dddebb12fbb
z80e1a1ddf744a6cd27579920c4620f470e649fdb262c3a546887fe0108641e85dfba4212c447bf
zd43aea17fca82132a7a7f48e0bc5da660d71e9517edad07e9a9d01a1a3f5f760457a1fc3b3d442
z5afd98a3811e7f91d54eb7e8e95fd6c9b607944014c6285f67957d84515c0e52cb7d7245ea9c2a
z0ec8dfa2ef524c9e562839d90a1a656454b91c7ef56add4001410477d31f56c9b32e87f8b52c1c
z2863e7fd274b1c293e1fc4993817338ff1a6bcd28f2329ab26c42fa9e87afa2f2f10f8f281a459
z894e6c3705eb6c40252ccdb351247f3ad4b30631ebd3925622c18b7427f01e127bba6311452d58
zaf2615f545bde959bc0374d97818332ca5336738d400d02a326b30e4fce9c7c18cc395daf15cb6
z6f3a58474240a64d6a0144c83b97fd13644a251bf5efe25d8c5f131c3f8bdb4c697893150fea2d
z8da66b9ac2df45f4755f176eaba14978a17e19d21a5a42581c0c68d7a350bba8307a63c9f400ae
z22584561a1928d35a0e649dc441b988024c7ce9808c247f3d80918492da00861cc687f1d9aaad4
z64c62f81c4ba36c39f060954793f850b33e964e990a63ad2e2560f5e18c794caf7fbcef7ff4677
zb9ce4c633c6676a4f29efaa923c4f1bc3c0b6aa8f54ded80657acfbb2146eb109178ed423e242c
zd8fcdffd4ec9092f2a83f349a1f3cde077eb17b2bbfac76a32d60a294a94fec7a7e9c70d4fbb4c
z410732d662db6984fb92c192876534d1eae12de1b7274d30669cb5d7157edfd64cf571a7f846ad
z809e3b68228c05bcd606f4fb29a7d41b8281098ebedcb73e941029df0572818cff6c3a3ad7f6d5
z403d94650344039ab8382e3074964f7c50eeba2b591c78429dbac184e06b20fb5191cfe0597112
ze95ba0b2dbc54ded947a9e0563e5b3121dffce90e371531d3373bc97741135d4eaa145b3ed2a03
z0ff6ce3f1adeb332f9d46e4c7c618eff27dae481e36f6f7b31d295adcf0b72570898cb652fe771
zd1a19e03a4acb5ee06be8b9dd03c4e569fc6e787992373a274dce20be03d849b1ba6f84bd73363
z8e5fa79734143d86a05977dad84c7500635b2358d43e5c34b0b770290b07255d2b172903d045dc
zf9267286b629c446932a829cab3330f0361677ff1a3c431dcd77de96f529a7cf2f6a8d14d0b5ca
zf62283922c7a386100ddcce414ed64724fab6da0a70edf9a05c9079add9e2299e4534719f4ff94
ze095b97be0df53856d7834868629589b744a1fc2a3f753441314508cc603add7a2c921be4f8241
z908d9a3157eb4fa7d31b80f476fab40f38e2791087504d3f7e6f27d03415aecfcf4b41aacd45e5
z39e3e5031250dfb0cdf35fad84bbe005003084d57f0d9a212646f3befb6bf1b43693101d565aa7
zf76c1a26d5837eaf67c6e03f9611068518563fef9d9a73d75d96958de3292a2b9fc90320e31458
za82c25cecb8c7d2da5d306a07aeb047f065a4e38cdba93a74f623579a2e834bd3b0761226b625a
z30084c554ff25010e7a08c2745cf0549d6ad757b9e40e77c6692ada447351e9ced5b3c789e03d3
zacfe3e8c15e0591b4bdbb310c4bfc1eed6fb431ac46521aea89a06caf9a79140d9644d7ccff71f
z5e0b08186e7a4aa9bc37a5f92cab9960ed61e53d898cc2a3bedde2bd0a67ba7b02c8b3d10749fb
ze8b18b47843053c51197923a97b3992c637ae97703be7a438c869de59531efab1079383be75dcf
zf7ae8403f5dbc4dbd826bf2b2c709f4d67ae05d78ee1844b8e8c8bd30dc4a8729d8c3379634b1c
z3881d5f79a7d634e78d33cb6396826204d5f4fda36e375bef565f7680933a31e4a5bbe563a86ff
z546d34f090b66613318281c1f2ece591cab6461a6697818871d494fbbb1628da908c53a355642e
z091700c47c5d9502140e9b0cca5a2cce5455f83e3a3cff4128cadb3a0411ed639608a519b0dd29
zb36e9c3c1bbea1507c24f2d186fc3452258b4a3a773d44f992667a27c4eab92fe19e72481dd215
z48145ff1c7e8297f4aabdb8333527bbd1aa4955ad9eacd8744f8350a0317d3e476a9119fc8bc89
z06105f586a7f8a4d2ee5b8c0731a8a4d1f4f63a20b0fd172fbd8777174842b5286f66ab182d170
z8c82c26633a5ce4a5ac2bb39e6ebb03f57c634e084f1c4e47dcadbf4689aa1f923963dda77403c
z4df833514b518aef0310dab14f9260ba6690f5339a096b488288ae5d20d1b9613929711f8b916b
zfe43f99579031f8b0f77eee391d018470a109785c73ab49071c89d5972600fe9af27cd9da34af2
zb595d3e85f168e392014ddd859660a8c1c121c2cebd9ab0283fbebd19996af4bbea15720e5179d
zc78027c0d88343b920956d61eec792de932e1d81cceb233facf66d9b0188166b7e51cf059a6a3c
zb4c5607090e6d75969f544e5661619f73eb785ae5ab02df9b456c730923eefcace195724f9e6a6
z216324fb8e1621f7b9d8db4d0e97befaeaf4ffcfc0bcd16e1b5c0e1da7b234d3aeb6353e231c8d
z147ea648046072085c0013d7a4c8d7b418c4d19613755c70dd8d247b45879b7148a56eb30eb2c6
z9ae711c320423358a4d38e69dc82e3b0eb27d86297056ad807f284648cfa1a19c5703972963eca
zb7275550a604f252559014144063d577d78eaddd5bd11f9af34e60924dd2e496bd04ba731ef4f1
zbd215816b51a1e316ab7bdd95820358105bb7ba495d62ed4083f003d61ea57ff2fc52b37a057e7
z52d68cf1ce0cffb37bf35a897e833391ab346f33a5bfe808f27e153b8a89050966531a6d6e0f07
z801736b06529856357bd5d08ee893ea4c3c658b296033291f62b78aa613790a7d5945762a5eed6
z3328e090b2c6c3cd7feeb4a213173a73a62e7e72249b1ce530ad734354c2d79fa79e47c0ad7fe8
z774155494e83e76e8dd1f639c45a940f8c0483ea7a0524dd95ee7e19e789df54353e80a1162f47
z2d4fbb0c69518f612a3309030aede992b40d28e8cca9be32c54b7d364fd22b97b01af0a11740ce
z467d2805d95a61f24f25d97a1f9d922f4d71629971908faaf3e6ece6cec2bf485cb179a936da63
z2a0c31b8b8aa45f78b06d68866accd2e772e9435736db5d112bfd4d3699fb23f4dbbab2343eade
z6aba91c78480e6273bc32c7a55a464561cf951331b903f83415816253a1fa1bf150b74649c9a22
z18e1301deb6e30dbd46b4c97bff637b9281d232cf844945a861d38fd613ebe37cdb1b02060a227
zf90e85a0dacb51d15c02898b6d8ebd2f41f7bb8a673456dd2a35b4908244c108f909f07a889c12
z578eeaace5ea14407d3d4d58f5058cd4c194a0554e5bcd02a2cb0db59e67af8ad7f5a3432e18fe
z5c80bb56c02750cc270b25500e7f2fc82a70fbb68c441feb785e753a17b60c686169f10f42a279
zc07341bc286a0c6011d11bffe9f980f3c3c718d43911bfa877a01e979602fa1dc60a319ea70fd0
z8e03a15572a9f819478bb52f835c2f4cc105eb15b8f37d8850dd1179a98a0562fe23e7b0d66f10
z1db9eb913d41f08635db26ad000848ddf51507ea0e979c7f895e53033c1245aec30483acb1fe81
ze645728ee3975debbd00fd89294393cd13938832820c95dd0be500fd9e8d752d09a358a68d881c
zaf30ddfce79686ca424bb0060114fca6aa4df4ae203df31aee190304502c0115a4061a42226a29
zc6c9d8c8f1a2db99635788c5bde39819e9d83a0464217bea916ea836736281e267adc8dd084941
ze10f493194ccb942d7192bed3905f51b7f28dec564e350e6fbfd24a5cd363cea5fc8696e44425e
za8e79a4007bc76bc5d5cb8031e789fb49e9fb7ba8f8915ed31f1cb4a421b298284ef602b838b0e
za546782fa1e663a3181cd0c20388a4ad9e579de726d1d9451d0cca63b2e00e66811cbd540fc9df
z1b66705b2fa15502a30670d5bddd6cd21363cc1ef759748aad12947a547065fc4a2ad3aaf4aeb9
z6d3886b10570a372f061d99236a389669588421070ddd96a5af33986537ff9c2947f649e14bee6
z161a7fa3cdd9859e42f5f184c56875a2fdeb9ce35b12f6fb577f5cace6144e2262d137a707f74c
z096e9d041682e03332505ba080bf364e79733e184735030aeae0714bd7d211d6fc051082dd976e
z27c372a6a3cdd69a94e8b40462d71953062993426faff760c68ada70aa7e64990b879be7b935bb
za8451a72a8ad8552b136fd5a69f9586af28d4f74ffa550c3e613ce082627755badfa4e9f48dfbf
z1d4354ebd010b3861b121270528738fce5cc29662b81c4d2b23e536ee7482e17cbff9f0934a171
zae43cacae8ef23e3175b792cc13f8b1fcdd79e11a050c10a67e1bda3abacb6b3eef5250d624243
z291dc8104862362f698344735f6b58e1628509a04745cccf4a65de07a3a827ae3c91f412f5c810
zdf9218efe0c4179ad52a9a6018169e33df4dcd8d85fc5f6306dab68ae8af635093131ae4a5e199
zd806b5fe0315c23664913c4e81a1dada0b8e785fb1bd1bce20d47f8e4f38dc8775e1e5767ee99d
z08eb10746944432c36c666a8c6769d2d4e2a2750f2b50a9026209c8148478b97187323747425a3
z7fdc62cbd30b171a77745fad11f007da2f456aea2d4f9274f03e7879de5c60a3b71c0421a5ca62
z7f5fea69031e0e02d3233ac59ea69c31a3e500b3270c8089f8cdc477b93e1c7e0fa8039ec18ea4
ze1287edd10fafddc0ddfa1cdc6d525d21ac90119b8b69f4ca9d3f90853fcef952659b2283103a4
z1dda58e502127c19e5b57633cec06510ff18d485f226f45ee3fc566d16bfb3964e0dd14eabf45e
z657a2d3f803e97f567dd252fca03ca3574f63a1a77e5374a4162043f5924bb5af136a987fe9261
z88e8f91ec152a39f97e525c78cfbacddbb5edff5f9d4a8debb490cca18e87941feb03a9501113e
z6d2eaf37f220cdd5bce58196025e5fcee6b4395271a827e53466a91ea32fc8ae52af22e0dac816
zb8c570dd89c7e398650d1ed7ddbd06922691669b3daa2f460bbced2f354f114c70efad31b416ab
z7d72aec10010565eeccf426b9b202e494f9b82fd44a0e28d95ade7ab0bd6e771cf421d0cd8f724
z7863e5d2e7e87868eab62a5231d3b3df3a764f592826a2becba55928844f9cd41d184887d79371
z27b764ee88615fef527616b691d8f00f8a654206eb0295014e223388a8996b42bdfda407e8d56e
z44c8c5367054b58860e9886416b3f57a11b0d82bc31f183f0373f63d8d2b4be1848f38f233cef0
z2a17a40c540d8e5e7abdd562d938cc29b5cb75ef881599b7d4687aff442833dd8a5da7868337fa
zc6a9af1d5454689b341f8a7846904cfd9ac5219ff6306fcdc4151e14521fa10a1b057afb4d4e91
z9e492dc320b161d6738a5b4cfa2a5133c6a8a77bc1f7ba4c8fdb5ea51cccfd199eddb6f1169fef
zf2502c2c93c6122b0e705b211e545ea2b4f5b2d227f5e109b017629320f107d8e43c50d9814d5b
z868e93167a8a615966749be2bf49466752ede392dd55ea5f20c94ba1452d7d9b89ce64081c6bca
z1719a9246fa13ad5b8600aa05fedd3256e5fe6c4fad03837a94d84a49b160816a6b5f4e9d1136c
z57dc768cceb39e84c2c3ca12d7abeb4885504ce946111ac393ef18766ba332c6cda9594da64cef
zb3b542379859a09afcdebcb1ed5250ae1acf51f13936ace71f9e8b5c6c7b0cbe040cbe8498be76
z89dbe340751a7d1884e1f2abea508332f57e527209c5c73a6b9c892b7013c4a61bec0e6353b27a
z2b39df3a31948104f1993f1b8b2f216c91199f9ca62b9ceb6ba23ae12082eebdc6b92d67fff1c9
z505bcc26612f0e33e84ad8a677e6279356c10bdbaaa345a3b030f9ea92b0f24a9dada0c5ba71e2
z80c850154e0fef3f4f579ef5403cc2f04b1c3c84d84974108ac3ead93487f5517cc7b8506f2e3a
zea7e9d5d39834d841d7d6a8660131d4a0f980b64c78c232d4f5c550a7bef382895e3802e2503a2
z245e051e47a29cb969ab730299834fc3b843e05f0123c877b18a7567c292305ee99fcb70db88eb
zdcfd1b32724c529d339d5ad4c1a3203796c421aae041085616fd61aa128c9a00850fc6f102e8df
zbf2832b1361422bb4ae7148f4465ed7cc9831d378a18b465597b4efc4547993b7e713dcc78e7d3
z3d2e8785c65ea7c845efca13a3491948efa449013cd9cf9f3f1ce71bcaff2f58dbeb19f6ca6e18
z04c7fc916be0a1c460ec0abf269064282e099a63b5ec6379a8ed82dd8826f0acc2b39db8ca53be
z9296f7a087d41e9d7b8139f4f96451ba2b1afc8a49acbaf7787372d1d501e87a99e84ac1ae85bb
z8be828e29116be7312892e66988c6419b07f19ae4d54979bf6d496788dd9b3c74033af0708daeb
ze8b1b6ccc3078da697d079acc219002d5b50c28ddb805f7d0f944bda977e47380f838b54019336
z08331a74231c787c4d80c3c5c79c3e691e9542e91338ee1fa17e90ee98c957499e7889c5d3b558
z0ec07e44a1c2876c0d4c62a2d45a377b883aa4e58a9b059700f11909dcf4dd7daef7a76f336136
zeecd48c9606f84fa3a28ab94ada42a8dafdeb0ef9d530780e1d1ce7ce4b8892a28609d7ebfb42d
z8e4ba2ed43094206e94bc2311496fe730458c3aafdf0c8b01d04b70f9a99e409859865ed5143d4
zd20b6fa89aec5cfae86d5c7b957ff57da96e0f013cec25061b761dd9559c8023e9e4eec074e28e
zd1422728b371594e0a69ba3aa0b7ef1c43a659bc0386eaa8af5a3175df64ac16e6d91b65c7127d
z8cf9ee46877653e1574b4082012dd574f9a371f83abb50b2bdcfb9ba7ed2a7e1662a76b4ae45a6
zbfbe3793dc5fed84a8e4cd88d9a3bc6ef3936888e5bd9773154c6489d4dfabc86bbf581e95b379
z70c8b2979d2001d3dde7157662908e04c8056bfff6d75352a99e25cf8a20468f4438976d93a2dd
z69c0d0f4a71fa20b6fae69d3f5818e41e0a8c6b29c8e1b572261c5099b50eb11a3cf3922aedab6
zbd6c67da723a2c78a09d32b73e91b52dbc24f7d7de75a73e6e2e30e82dec997282ec2a3159ccbc
zcd37dfed975fa2abc5db7dff8b7a394eccd133a76fedbb765450f4206c2c8db80e36c50a5654ee
zfdad5444209275d41173a381e295ed9469d836df97f133d367977749b3e462ecfee7fd2379233c
zc526c9a7cf2b40de83b470ac25bec39349d3d169b34fb82074b2d69b9a71cc930228ad9c53ea5d
z2c8cade48b0bf70299a2dd1ecb874cbceeb142e78575a46e12a44b309a0ddabd856d310123fe3e
z315b6d3d399cb106c13b2d50a19f03bbb7e12dca6f09cfd6aaa45bf5d5c0e742df091536111838
zb9bec2e12309ede99a372f1c20845b19d7408af2564380835bcb51a3ade48d1a2444b6ed205c01
zd0d3d3d77930f720bfc18569544e24e3960bf468fa075b638c342e54e3b7d8a74a0ca77b31d53c
z23910ef475388cc4ba82a91215c3d105ed76c5e2354c1a28ecb51ad64c192a0267ee438078c213
zfb84052774239ba45affad4bf0b0231dd1295691d7665035153ccf368adad371c33f02ea2872f2
zdae9fcd70bc78665d4da3b85832f8acd156b48ddd4ecf53a0b0eef4b2a269c4230285494bbd1a0
z702c883f7d827c83b659084d88215da8b5a9f12b8bca56157b677dcfe1a90643b5eefa92c69b93
z71755d0757635a0cb0433e4d2cbe49990ee46176cc08eb972cd7273e0a5e0e6dcfc3b932f10578
zd8606a1940aa0a3f2d07924e6449083684f7efb43d1b9577a109ce10d6d587392df2b34b4a40d0
z38d4361a4c21f99f970ff678429ea74a26702e5ad1b603cc4c5ff38390a7e9e9764c37df2def06
z0d82493d6e57930e7503b9b0f9f50273235581291a42085b92f6bb052642210c2cbfd871d54a3e
zecae4a18c4697b4ac1ce08e7efff350428bcfa32d6c730e4f1ba57447ecc5f223bf8f493b0d437
z11ea0b4ee5c7235f135cb516d7f72ff68d70072aaf696ecccb9ad13b1287d74f8b108be8e85bb1
z801b134401f72204a75c91d79215b7132e3a930f1edbfe8068a3cbe3f1137db8b28507cdde986a
z5829bcb7e97545658c1a6fc01e425c2115f1ef554e5f5733dfd0ff6d1ccb775ec248077b088e67
zfcbffccc25b39c32b5f0814761548baf086c0b51d0b4c0748248203a7ca4d2bec605c3104eb381
z68bcb8b295ec82267b782cabd387f403fe0a628779ed4ad8c98f917354e911c62f822409a64510
zc90159e530a02e5d24db442a587f28f2e7a7b07538e7235d26b9831863cfab83d770896bbbdb6b
za718f30e8188a4145222095c46624ef7a8ec1d18cdb344a57130da10218d4c4252dd802a5fdfd7
zde094cf17e878863c3138bd2d34bbaae64042afab9e5397c5ba9b14a45c9d43c8ae23f0f20daa1
zd9ebd844d150bc913f55e22ec5239daec837bd1160f4152ceaf2ae8027778dc28b94b83f2946a3
z3e7ba8a27060ebf692c8e2562ccd21467256f308ac56b1e96efef342464caa59f4ad956c429e9a
z63893ce96d015c027b568b24f2337e76defe04c34b47849304f3a002ca3dc254e4afc45fd52d83
z95b52503bff0c77f193ea6b84ee83d313ce6e99398ed27a9c3e9e839ef1e9bcbf76d69162874ba
z80955c6d2f8bd1cd3e05427f83c56f51c3ba079e39a8a4e585bab36d1be87a0d83a105dc46c4fc
z2446980e37a1932306635228a94c44f716b6623a8e4895183097a5bf4c9323a3fc0c815b6ec3bc
z4ec038740ff47aaaf99341187b01a66717b85da1b10e0797120dcf55c282afa0b0d8b3e32d74af
zd5696eda3d3b2d9883e49287385ac8f0cde919cf9d05a01a4e846d521f7daaf4d9bbda49074e19
z007d70bea9506584a7ee912a3bee52db92f17d5c186dfa7cb28868a6a869dd4efd2db1a8fd13f9
z5f9d394700440eba73b10384b8482f324332d7a29daf7e4962939878c2d10359d835c3baecb044
zcb4b637de72c8c82eaa6970887caa5ed00db114e2a1e3de117659c11cfb1bd2161c45885bbd264
z33ab0afdcf2d9a5121f942e3e09349e0df7e6c4a372256019b33085006f52401ba0902b341749f
zfeed12df954af74e3c7f361025c209087539b058c235a757775e9deb5c29ab273e67624ef69ac0
z26736e077547010914f082ec24d20fbdeb4428d7d8d904c0e794492626f231331654d148d22628
z4830cd34cdbf37639458e5a007bad91a4fdc301ae587e0eb14c58134bc045b13830cab44287bc0
z087e1005666fcb475feeba93b3fe00542a34a094308cb0e6ce56227ea1a1834963b88c69790454
zd0c211e80cb1a6fcb6815a6732e38f5cb225daeb2e6435e291e74eba1788dd40696f823e724a6b
z14640c3c1b211bb205e32b93c787849db7eb5f3b59c51eb6b70c53fa6cd439f3ad13e36f2ce534
z8adc0c201afd8a9e0c16a30c176b41e5731f4732d87e04bea8779acd097bfc16b0c0158ce118e3
z0137f8403327aa3bb2cdaadc3a21c01355e47d221c21d1ea6acc544b2fe420d3f01aebfc9a4930
ze486f23b565901ebf53ef249b2f3c2fd9affd107e145b912004b081c82f8ebd173d011acf7a65d
zfbe8d123d6029f7652d99709808adc3a4c6d0cfdc8970f4731f5a8dcddabb2e05c7ffe7a1d29ac
z9632a947a491f53188d25ec6e6e1ebb2a9a01bd632b4ff3f313b758cc5cb2c32b3510861fdbc42
zf8c86f39f87f2fb176ff5c921b185f5cbb1a7b12a583df8af79af1c44e5b37906324313f4a7764
z45bb76dc270f776a34b49d8be37b9c7c29d41f890817519dfbe5ae0eec5958b034bc5473e82462
z99a05ed2fdb1d078e3d1c822a665874631af292554471db3c11300f96be68456b09e55018dcaaa
z67e693f3cf889db94b17e2bdbaacee847e7663f4b4ae8e921cbb6e96efc0c8acd1ff3e49453690
z5c22d32c4f7df2abf67ec3523f1f428238d5a632bcd3fcbea1a42ac92aac9f77f72901db4c1250
z8f2e47bd137174d82d705601df8811e1a8ead9f558e4b3d62b5633d4dd3696d5d08290efb3983a
zcf3fcd3db5285c9bc938439a4742ca457276cf37f9aca73cc381dffbff6b607c121307c677594d
z98fb8ae9806802c812a686d89a92655bb58d805e2aebe5de3b30d4053b6d137825fbf357e08085
zad55d772c52a6016cc757439527fd257075fe020667a793413d38130314a23b86799462520b1bb
zccae5584fccc09e7807aecfdc08afe15899822a82ea5805ae06215bb6c753bdf0d36412e8349be
zf2ffc959c726042890e9d8b213c9317698b23e1ae6988e93656d7d6e99d422cf880f3de7586bfe
z4e929492d452615d19a615c21bda66f5f59614a09f805af8eee97c2725f45d6843e57303cf10f4
z1846be9379c80470fde189b4a4501505c7d65d64724e77dd39feab66d38457c20790e61b19a037
z6b1742c16a5b1b819a1021bdaa0080d3d236a2a37f8bc9f1ef3cec432c945b40b085123e1ad50d
z850f37609c980c5108982f973e36d178749c41bad146582f2e8930efb2ff328549dbbca3f62b0e
z4bfc099ce2516da594a25870a8eec51857a7d680f008e8cc5eb36e4edb49a00ce393470081ec17
zd743e80ee7d5639cd747a79e8f3a57391aa76fce62a047251e273479306390e43c5f72688114dc
zc4d6eecb8cbf82f60f9cd358647a3aa5d52714fccfafe984bf4b9376d4f977fe1b20ea51ee70f8
zcdd7e37ee2bbb71f210c489dab5c724591c72d0a830e9be6c1cdfc64b81c5b2bdc28eb5692fdeb
z0c39047807226528c853df3ff02f995351b69335e8fc91de93617d3218eb730b295b29579dadac
zaebaf354310dc195544b4d20a3a984ba0e79925bdbf15f9c782eb1a5977b6341ffd6e4c9da031a
zaf24c07914f30143f9cbced9ba8ad67d9912f96e2567cb298991070c74f2a876c8c7ef5da7ba15
z9f89ec7def43d766096f55d4eb786f3547da2c0ddbaa53fae28175ffd896834c4967b9ee7b733d
zdf07594e893c239e753b1f36e9390e92cea1616f27f6d084b805acaf51febdbacd36c277db8eca
z693a99c3f91f1a262e901def50b98fd4886c1e357c9a7695a5b9c861dc47d6b9dc67d941942dd8
z4d18cbb92dbec9a92258093e7e56cb382becb20ff3d80edfc79369af02d5ffaf3f61cdfdb22ff9
z787103a2a14170e7d8155124b94f5e8130e2eb04a6a82c640f2e01b6e6dc7c278cd194658b6ecd
z7e456602e7dea0cf82c8b81e5e48d817fd1445420dc4389e0c9f4cf196785e7ea88df55ae55940
z849bb79a4485a0e6cdebc65d72a2c605c9db40f8d654cd2052ebc69e2156b6e67c6fb2d3cf5121
z5b461b6b6c0b83478dede712ac7492ac2e17e369a69ae9eb74292210fdb48d761fdbe9d7a06037
z3fefef34af2d49b5f4630252956be65c434244d508308108433d186c011b113565333817cca2f9
z2b5366b48f1e9d39dc27a1b10ca85d7a4d56e88c551ceaeb7392618494b0b4811fa2a0dfeb8e3b
z820e2168a58ec7e82ad54100a0bbbaf218202698ceb70b748c54c7845e84bc9997a8378a3acde1
za749336ab9634f6e2eb916a401e08c6fde4f1b8bc4d67957d30d44b7d75ad0ec7f4b7902f35113
z6c52cffae970ff125797329158bd3892686425d07ffc0ff884e2293699336af4bc72db1c802573
zfe2328902f37c42345e61fcb4b6352efa0dfb04fd27625597248a3e4f966f8e94582f6a073e1bb
z5203b9942c335d9d8259750e5bd939c898daa7649638a14ae87b9955db40d917c48d625abb582c
z7f35cdd1041cc3be66b0c0a7165d6ac6af823bbe901133908616227d984f1f7a45d981b4992633
z445257c0c6bcfea99c0bf19634caf61c533da81d45c0f23ec44a6d5761ee369813b9d4451e2b7a
z658e872458ec73defbbbac319f3d2937744b03b63c29e239c7905cf643b640befbf8244f25c990
z4ef0c9df8af2cdff06ef57c1d057bb294619559ae8aee316d035f97b1f5817e9cb762b229c72fb
z0d26282a75065e42e37bd3a8ba0c347d6ba7ad2a4a700bc8e877d62adaed38547f4bd2c5bc5575
za4013be0d2aa67019b155dea222c23bc9352f03ca0cbd826f40a8e83405c80f6b9b72b1af4703a
z8ce29736ff93c6a4da8327fbc6e57bf099298b0e80a80620fbaa87e0c03902e765edc20e176ded
zd92558b590c61ff44d8e231b280afd97d75e4b782d35084b86d56694247922e768c89276eb8f26
z520397130567291a7ef3bdfd0137e5aad5f13fe6c19b3b654cdd08024e300b321eadd33a060bce
z231620601d3608ddb381a20a8cdc20f47a4de06d5808921bac64cf6147ac201a2dacffbf4cc4fa
z2b490d8ca883c0e300f5b1e0bce3b523f891437ba5222985ea16e33856aeb0bfe8417ee0b7c4b2
z7eef9fefc001c682777c03349a46f3c065e96d3001eeb70ed6660cad9b8de0ee60200f48604623
z0df951da39790ff8e2b6544df246e10003db6fe3e8d1e6057463232194fbb496eef462f43b32a9
z0aeada5481245b944ffc7ca6666e92701799dcdd4210a5be3627f7bb0356430446ba8605cff183
zcbad8deda1b651eeb0d92c5acde74bc181400c2c11f593037f33ac6b7b0ab33e68dad89e9fdd2c
z8d8879857326566389bd5f68a553b56c8911e9d08ab22951eb16bdd0f8913f19000dd4ec9adfc6
z5f04f6e3f00853533b7098d1f3b32f7bbbc764328929df97f6a8dea8d7732a0fb98860f0859b65
zd7ca7e240221933fdc0d26c2382b57c2e3201b866788c081599baf43b34fc273dc21f9ed4963b0
z11ecb0035a8929080815c2b26e9d9c2e15fa2d0f561db3451a6c7d2f9f0d15540a873a9dbc72f4
zff7eb5d09ad162298a674a3a5052c8d20646d8b80fd68526a3df53a9cb149f9b8f20a8cd7d0ed9
za901738f3a589a95fe6e697e6d442861d594facc5cf87c8ff003e0d70a909a429ce4d0b3e25607
z131716c7e36e1739173dd64746f4f8085747b2f6adfb6aca0c5bb824e54e8c84de8fb27a8c900d
z7f42b0bed1a096c149971fa3e5250b8d0eb1ab3492d7ae4bd02fad546232d8c9768fecef8502a1
zaa137e3207f36d120614dae999be1e04b20f96367924614a7225a306b4e9b0d74a8cc27731c6d2
z2fe51b35902532a6696f28450ee1fc6691e6029ab52d2bbbb7d9cae47eb547ed9fd385d093b0d4
zdf910095a6660fc52472344c4c9ce77ace64ad160f2b12093ce5609c66e433ef8741637591e066
z802707c8e4a23e92125aa872f0e2b3710c922b4d87e54a2d611e55043897851a2b6183980d2eb9
z0b1889841d0f574245a4ca12a44e482ffe0e8e0fae9dc0ab3264497d89e33d6655dc2bd78d03e4
zeb8c99844c8190ba82f01d820215edf41e6e68e6c571eaf1a53dc45ccdcf9c7fb8ea6f5c001386
z0c59181e977a512dae9d659a8c2ff81bae12bb6cd611c30b8f548b807672e5746133c23da3f795
z95ab24b29e6059cc550d5365fa4a8be149ea84b857243ff678b68b2dc689a3b1b879a35fd21d8a
z87483318216ff0b8da5cdcca8f57f772c7e69f869f52f44a6888809dd7200161fa4e0136e26f09
z9f524981f5eb637ec325ecfd378401f6affe178a78824a06290c548586a8233213613f60972d20
zd2daee12ad00f176bb893b5b7176d2ce52585cbdd4ddf6a80c7ea8d18131b0c0817b95f1f89527
z2c78be5676074c7058e64b6f236d415d5025b4857b20e865a4000319d0421a238514ff02d8e280
z70b65fc354b7c94e1607e13d023ad4095531e4486da9935d352363431a9b602789582e69a4ddfc
z60802ff295a7aebf0f89e7efe76e0e1f27865ca539002d481beeeb4c0594f05cb36cc76f32ed22
ze0c2b0ef4a291581d07b276382d17cb0863be2b77913a2ea1eadb8233733751105e7489ccf1287
za9591e93cb5e40bccad6f5e9c8948c6e69a0392b99cb3a0036b6176a72123fb180bc2158927624
zd69b1ff362068579637f0cd2db7889c817235550e4ff29a02948120964754e89f5ebce322a13ac
z3356d3af168abd6075234ef4f5e87457b38b06bab84ff210d6ea285434d48a87d57c1bd5c96a6c
z92a29bee8de39b9ad8c1d910ac0c5a7f67b825ccfeeeedfa91735f9ac95bae1b9a23aceeb4847d
z13d53fbb7b3951ed97ca8d93ab754b45b1474bd859fb7a723671ace60fedb83a4015b891c9880c
z4e952c94940a359d48fce4cca001760052fe756a9553e33244cd6b59ef25f16552586cf20b19ce
za1eb70fd565af675b333410d75070e0babc913fa51eb727c40ecb99330fd7721f6b20e98bcec22
z778fc1ea19392ae3948e324963b7a77948b007c78caa8eb8c9b15fee0faa281b0ccb2d5405a5c7
zf8f45fae2a61fbf01f031aee07ce04661b75f871cd54d074b11b53d1594c6c6b5513244d6a64d8
zace258852bb553c1256ecc153c8189760a984e288232ebe8eca9b852f35aaf140c77c096987ac3
zd2fbd83121e5879c53d66c16ec07103044f181fd99362c5b7bfe5a8e3d074ddc0f805eaa1b9ff8
z25c5c704dab44fceacbb594d271420dc5407042f76c89aa5c75fd9f1fc9a4fb75741ebc649a1f7
z718a439f2c5ba2c847900336686a9849a6b001e33d5aefe142d7d961b6b68ad1daa1f804084e07
z32bc2203918f0b68fddc063a748f59083415ec61da148e25a56610c912d3dff98c299bc2cd6d4a
z4e608152965058896441fc609c33ce9cc82dffbb80eb684ead12d1266c86b7c949d02fdab671fd
zb666f0b0c85151bdcf93979289d4b44b8ff08a666e725b961b61b56725a5065a9fb729b1f0c454
zdaa4b4008044f6929f3caf04a3d71d8da231f5333f6bcaaf14c50be75bccce4cd2c2e3b2c41b4c
zf227f3ad54b60656ffa616b1ce0e25449529c6cb83d98e8d1a591fe56d792d5e737982d0c7de5c
z323ab9335fa6797eda84b803c184d08e07276099b83ddc853255c97a6dce9e2c2c6cdc98ebc70d
zfe024cf7550a72bb2613718151a74e56cdc05122e5a1acce5f95d86fa1720bc2af5df18effb8ff
z804a85c24d48dc2943540bdfc32c37e947f90b17abcb38440de4311a906faecf57475951bc1c0e
z82e8058053ee8f0180f994a9fd040b822e9d3c1354ff013e0829921bb2c7f56e6c5b7d842862a1
zc1c5a479bf925144afdb2f4a21227d1f8c8e973a4817d4b6d4872b77a06a801908ac845d43cb67
z31158233f947b25deb68028a2dac1474eec0706858941599aa7fe9d6a0926f350c655ffb5b3d4c
z44d4abf769715947317d64f45e58952fcdce0c868e0a05b100aeb42bc9d9ad55200cff1fa88ab9
z7fd842a5391d7d9c388efb17081dc68de6149061a12dc98c55c295fcd653aea0803876128c07ed
zc4007d8c594f253dfacdb6e9a6dd5603714491b533bfc814f203b51ef2d3e086fc9a163593c094
zd4fd48e37c73a264f5cbeb683f7189f939ae513fe300d5db5a56b3623e66707bc6cd90405c74ba
z39d2554249681c5ba0e3ccf3bbcc9bf92a98025070e242582b5424e4c6dfd54ff6f16f0f3511a0
zfd228bbcf626dcb097e7806407478afccdeb46558e84ec8f0d523dc63873221164ba0dfafb8c08
zecd82525021467737668988b63fb0df73be2d13352a7440740e2db0ae7defcc1d6e1f6486df1b5
z2f88cf05b1d0f491eb98fc49ca6d0f398f835d29b8e24ccc921b0805076162e4e55423eb0de791
z7cbab8f834146d5e64f560bff651c7e1835471b17bbe48823195a146047d543299c10877233dde
z0de0ab64e8b26b5feb7b93e8a351a934d5975b0bfc2f9a8692e72d6c3eba926128b5a770eda5d5
zafa574ee5397f51dcf680bedc48f4b5d6a2fedfaac2da2ed9f4a286b791750f5013c5a59f0b369
zd5161e782400f019e5722e4ae47556d37a570e937b7acb532c61088988865c958af8c3d0150fb4
z824747d9e969a5f0d220bedcec4e9252d4b81cb53d606f19c21e34f45d270d2f04535d37470674
zc5e55fb548efe21fbd8101f71f2af5b9b1a563a8a7fb0920b361fc28a5495b6435e71c0714f071
z67813aa2a77c6bed834b8001f520ab5e273858e28dd78045047d5a9f1e16ca52dd1daa9ab3cbe0
z9855a4b5e433c98a606c5d54d2900a3a1d9ced810b18a1ea72aec303dae12ca3151f507949270a
ze61830d0029a887d900fd4017c31130050204af019782014df6296aeee4ccf7e90af241ae9200b
zd6d60105ecf5b7108f05fc0d4f82ee52562aece01d5e31116a80136e996286b5aeb04d7950aa1c
z71d41997cea75abd4f606bc2269f4922128e94472849019502632623c2dbad853bfdf7415ab78b
z8db9d7f967424e676b1d07789126167de779d7334e31fbff587daac93cd86eb9e8814004ac53b0
z5a27b20d40c0b8f6a72bde4aa5ce62abf117ba5a1c1039b70ddd6d8539b8e6aca099b26a64c14d
zeb75b5388560259fca13e85de4649a2c4f2648e5f97ced66665840c27883bc1b9f5457294221d9
zee1a2cc35a7a8fd5027035c823cb83ed1b3e5accf784b71e2d6d91783a4863034e7e66e9d7db56
z62591891c3cad4cbbb16eaf8b574d3622bc4c11d1dbd36ec8f9e363adc8fcece92addd3e5eb9eb
z1596a7172f14783e837662767441b49256fdfd0dba882f9df9c4ad1736d39adbb50fe5f1d3a4e9
z1053a9d479dc93527a217393a28ff204720dceb58cbaf54d64b3d7aa2e7ca172aacf784a3caa4b
z2624539cdfb909ccbb188850e5e380366861503d197af6cafb62c6448292275969d294355640d3
z7fb81069bdd0e42499cd7e0229074e9721729f1a5b30173544dfdb1187a88dc0d81b23d0a46cd6
z4f816c7176170982f9006954bdf0f2c8fab7c7a7b93cfa23913653a8746f67966f456bb8c1aebb
z049ddc7fe48635b455a7f75046b988afcf743debb3d613f5beae06a1ef7b6e2c06f6dc2ec5de6a
za034b4f2c1bc8414b89bb0a31d5a68b8124ff14928a7e22fb5150dd305e0f749040e10aedf311f
z4f08d3b8a60b11dd0cbcecb2c399077f88dbb9de1e898a1365025ef1924575f52a34d3f373cfad
zac339a407d5a5fc99208bc36720aee98b164f65efcb80f5700b716159cacb8dddc8f5cd7886bca
z613fc755ee39c5e61e33c681a41bca8f63ed006eb19185c7bd0389f4878dc5d01df0da70237394
zb7a57a19751d66b5ac9357f5de6d28fbbc284719e75f42b6747459a2afbdfcd57e2e108d9d1726
za05153c1c222d8119df64427076f5398814759b279c4433219cb3d67d015e7d25b63bf609b203f
z880337801356d6af90ddbf1a90744d0aed87cac6d103d6404466b5df1f547b80667ac3089b9e51
zba088a4ffb803e30bbdbbb0eab2599f85b0d4e79e69d251da72b5800e24b4e4cb7d3f88a3a1d8a
z8e882a17251041fd586543e0ddabdec767419943f0d0383288db8bb4fc979dd5ce9fcdc48c634d
z879d9eb91fdc78c21b9039c7d81dbdf74e42ec2d59c1aa6d6b4efede2fa15f66c4f3e0bcec0f01
z544c875cb2d3f1e70eeaab1f625d28f748cede4c8f2ebf080998f41d1b11d0b0eaac74872e63f1
ze9c0bd0d741d8fbc06aa9aaeefd34f5c5b3f966f92c40ac856d90b92eb66e3e5c019f32c3b2188
zd83ff7b4b12b023683a9b125b4c58d2d3d1c50f1d402bc3f813752189dd780224a5522f879f721
ze21a8cdcc76dfd16464a6c0e597f11a1d7946ce86a94a89d1c3d4daae47ab5e4276d41666eaa87
zef0c3dfab2f31067688a08db4c86fc8fb0af1fc21177920512df05c7b937cdd3613d752259cb56
zb225893cc03397689cc4c072518014d79593b77fa8ddca38c7ac711b626621ab28262b10d9cfc7
z94e9d7ac2f7b5da61ca350eb472c3aede97be7890fe7750dd6343c089fcef81fee9cda87cef0fe
z7d2d24b605281136eaf3d46230320dc0e6ae2f7af33057c1de13a35d73cdfd2684df18d2ebfc21
z022142696a3be57d8a3f773a33fa8a45cdaddc04797d687951d65138f4174243095efb64b2fa83
zc123cf20aa7a70c4999f28c8e10bbf0046afdb0ba25cf788c94e002009edea2548306f9b333490
z986babab7910023fea82aa8b41d789258a5f39c7bf0871d07535637e4ae61be19c9ab071c14a02
zd83b8a977d736e70c0224304d4ec8571d438a63795fcbe9188b6d8c501b1b28c08c937e50f5321
z77855ed00bf2f45bb5b09293671151951a1b725038dbdad7209bd426240369d632d00aa1988b8b
z86b85c4f270d3a7ca6072169a4722ffcef20134a1d39fff7aafcb6fd2d1b2cb9b602f7fb36717c
z3db07539db67a32a93f35c73842358afb77d9f358eb1dba9b57a33bdde05b40b3f507a0bf61c5f
zed32a6c3d329a823dfb94a383c0c561c03c74cec8fbbaca9b1824fd58acc08a861514e00e6b00e
zfc38ab1046af7b19fe098caa8916e0b6c803b42107df559f851b293418a7840d65970b22c8a6a0
z70e80cc406bf04e93322dfcd57d9a35794b8f1aae3ec6b0d10684c19fad9abcbf30c7bdf85b670
z50c105baa7355444e459e6616d2d40d70b57febf0069ccc3a9ef768cd92f842ea9b440f1b01005
zf7db15af1d6dd320f27abdfbdcbf1d6e9dfbfa90367f83ad2b63619d1491b20a79d0fd150f5351
z448ab35df008677ae90b0a415e646d1baf866990123f80244875928ebf2232ee05e8cbda6dc417
ze385e614117175f1d8546511cb0e724a1a4bb26888f59ef59df40cb92e63198d1394bc0fb91097
z42d91b735208813e3ae5894f441449e7c4d748aa05125809eaa377e10a01b05dcee57dfb2a44a7
z2b3034f7ee585d9c653094d4c461e86ddb7135991cf49e026472263a4d11624d4e7bd1eded18a4
z44d0b82b0ccbd7b5a48e6f039484d1bbb2d9ec1cd91c016c1b089e4c3318e6d51594ea0b967fe0
z2a1c1d030e25853d30a79bc29b19c927a4e91ad0747a1463bd8194ee5cc970abbac0da53fbf47b
z966fac6212abaf6dce3869802175f7465a94c020ed17d7a51ee5fbcaccd686ead9143979802156
z2fd5410a2ac3400d9beea8cbb3608b2421471e3827afcece63c06bc90cf70232783547a918f348
zd6270d60dbe79e8cfb07ee2349a142ab8216282dea61dd3a81676fa53544e405cbcfb2215c4c55
z7b1e192293f8dbcc4d5276f5e5502742fbed5dfdd81eee37d7d03eaaeffe4fbafabc6cd952f186
z94d49c82d6fbf65874fa5df97a2c37fa29698b09e2d6647339fc607385412135fb38086f79f93b
z3b211968f14fc679d7d760299bb0d3ef12f5cf58fbdc1718aaa99534d37a47c5b2ab95580886eb
zd334cbf9f17096af53f326ffa1a462ef080155cca77cc3be0c340e470982a5dedf9e79c2825e99
z68e06b0d0c26e64985ed050468cfcef0799a53985be532484827530dd7e9f3a5dc28d7d38eb099
zfe681a8d130a2f8273e3a7cc90c7646301e75466c6d327a95ba87ed69511dfc0c7f58a693175f7
zed2c7d0d120b30143b23346f0c75982dfe4cd2ebe9c7696b95604630460fff0773948d741a36ad
z3d5ccc7efca52fde9a59075c8e78ac96261320f7a650a96cd437867734c626227da3d3fc981271
ze103cf58c40da290da97a1b47566d4e5dfa42c52453251de8bee10786b2de541d5070ebc9ac1c9
z83e79854f3e78e22e3e2f22d4ed8a1afe8e57e9f9e61b767c1202c9c05c8079ca9e586e1cd9916
zcdc53abacf4b091e29d56dfdc184a7d56ff2d709870c34705c6538cce6914549e121ce93b7719a
zb61931728efe3c4c704fd0101a14c9e3cfc2ab5b755dc46fb584cc8b1eb03423076cadffd2916d
zebc297b371450881502d1a2c827c3e6ec36836ba276ad830e0733cb4314aba596f04c494395957
zb722087293ce1619c377358b4982b7c8b97d502e0875addd975842f11e2da09fcc021ba0dfb001
zc50ee3c9308cabe85769f16c125764439348db1137acdcf825c738d8aa3528742555b4b0911ad5
zb8ec388e54c808cbdf83dccc7ed76672fe211cdb0738f08cc3be6bf19b21708e691af8ee043992
z3b15a097ad72531df18141eb26f0bd48cfb6a9b0a0b9042b121ab785f759651cc63cc30f876489
z9e6de1d6f15b4a0d40e82176477959b16e6630abeebb0088f3a3fea9cb0554f889267a1ae567eb
zf251255735ba6b8c10210587e1fa04c4db57987bcb7b3010d22e3472f2fbc77717a7ff5a39e8ea
z527458a4d0055c9eda8f83227ff48dfb55434002a8fb1c5baf231ebebfb7d04029ccadcbb12eea
z2eda5d26c29c3f49bbb3bfac05416083a724ea099810705242d0011c09bf11146f3ae24b508285
zc539b1be10e5eb4404d40604712e6ba12cacdd746b7c1ec530c85dd356b6ffbf1223f6c9167da1
z06a0871e13bda4163f76334fa5cbdc6dda3bbeff2de4017332a59b312890e053dc81b2838bf45e
z6461d6a72cb33332c322494cb2b3941773572b38306b9ed965f2c45a857adc4c952fcf18fa6359
z1661b2be7874a7b0d7f92039eb413daa2e37dd4357fcf108f151ebee6ccbca2e246f87776fa0db
z4575188ea1c3956939f1f768ba7361be80008d6df6b4db34d496adea82ab2420c7e1152d840858
z62266025619e5bbcc5dfea997e1a020942f5ceedf6ac7498c4a9553b451f64da0d7168761613bc
z0b3b0004d46c517c687d41b3f51b7d98e910b3b7b0bea0438780f716ba7a411c5350f7f8140703
z2955e0b10bab35a0f0a151980732bbf8076e60807f431e48f41812eae91780d60f6899cbfb5218
ze0cf60d2b3d37a0dfd0a8ec0f4666691eac6da7a0c2f8e367499cff275ce369afce1c5ae44a480
z8a5fe9c5355ae83a50fcd0f4f2f32c2e66ab93b83c49b78cb341d8967f645971333012cd687e4a
zd6778bca35bafb3cabf4ae371969583d5898d1cd19d1560b77834f7f483a24380447ea45fc68f2
z486cb0ce68e338de9c29cd015d49c490443195500bda8035ad34403500a0a678bdba0c92b0d902
zd660042a930d342a44ac832c0ed15346ca97e4e1b30422f73939a429317709d2caa61b9e2b0b39
z1635b884806d54871cde793df33196b793713318c8b3ed3f51e28529f3aea692b759e4901014cb
z1f46db6115255acc5d386d683e6bfaadea41c713d9d404cde752c545b4e48003079cc17036d2b2
zf8cd19beed84e43331855705f273884afce17808a4e90b3965581f2fd9b7996500913847b66221
z6c3a741f76f6a31c7129c4f974489c102fbf317974442882c87d7e6c2e21fb81b03797eba7f2bb
z16fe4f05c34087fa3682c123d4e19e085b61424081e09b1dbb7725f8813dd662c9faa17902b3f3
za5c6a4edc22c6dbf341774b93adaae87ad3fcb99e89a917ebba476c762c191ce740a5cb3938cc8
z72d1d19d49f0c3271e98489dff93df163a710c8069cad8d21d71ce3a8c6eb6999dcaf0a7959831
z1373150bbf4b34670d455eaaff01f397c2545d91133cfd644ce159d18c348cbcd1cea7842dea01
za4fef799fb5ae2181032e5fd347289389ea5a06002eb36c9998df3a9409a676854b873ca0b304c
z09fa4db47a6a058d17883617c0db2c400f739745c8b95d868e7d63c8fc69f4ac48847d99221b7d
z26fc6436dc158c969b08d1b5bea1d00137f7e8f513c60db9bab53954f74507ec15dc61eb1bb06c
z2fa0640cab6fa886a12b45eaf5967e89ea80aff46bd35c1bf51d143d8aea9a52ca5f275a41df7b
z19aba5ce145fb5bee09028050d401250f2a7e251abb1c64c576eb53572cb2735f205a4af3f61a1
z6e432b48a19c8f8262dc43e22d2217d6fd03068c2c36df2efc59294a2a803bce1ac2d32c62b2cb
z1b72e7aae718fc379e0cbb5a08ce790ae04972d4b3dd4b25677f347507754736c1d858d06b8c05
z632e016eaf0afc4cfd2f72c09583a20b0c606bcca55662824da2fd5203ec598528294bcead2d43
z3431c420cbb75be36954be193a228b8ac6f05eb60e3cfac6f6a12d965b0fcbb86983d407c34369
z5b54d0c50cf754e6cd82f078bf77d2eb9fd3ad6446107391a257d3ffa2222e8563b233ed47fd02
zad33af669ae294034ab5dfdd3d4db3d38265b1e9ea64f95a6c802df9702e8d4a8bffdce861966c
zf7bd53b097b1e97f5473719cfee3755947e44eb62a9c7af6d7acb5345f7cc30d405b31b731e8c8
z00c235dda6071ffecab579508556d1dda512f78e73bb572441b91027f87b4d2e4acc55fd71cdbf
zd87631da853a45b449c7fe2f972e31f464ef0a82de5535654bca44aa50b63d8178a4e9af2572b8
z7c62cf59eb84bf6df557f4135a152934b2d5ca0ad489a9fb05677f6ecf9e15700bac9e4a5ceb05
z43cdb4d3704fee122d98dc91bb25a1f362fa2ba4eb9670ab5d032e10aa88b5dd6ba148b081c11b
z73a85ad5f5e63a57ff18731d47329d8af26652b775a66634242b58e5f6fcabe3d293ee5e1d6b77
z73444a14ee22733797e45cb765286869c86d5a2491489f311aeac9857bc0a076c7a28912f0fae2
ze537952e8da9e4b6487e3afeef50ad55f4e0dcc3db49a8f18145e9d3375260eb867c4f67ba2387
z13fdddcc46111dae4f97a44b24769b3f0ceb0c5f9e63b4a95940031719113e21ad7b89660b0672
z33c4887a5bb1ae0273c3dc41184a00a83bfc918064d9ebefd8769376c3cb928a88ba70f5849cdc
z4808e391c6e1374b448f34390c10dcaf00798c6714da7a0d8cc71f4ea183a54e5b65b75aa48b7b
zf8c727c66bfecbddd203e86437cdb0bf8cc0859f00a5df326466d55a802ff8a3f0e862eb308893
z741d8ac4d69dd18457c3d4a9b012d04b7b23ca46d37b1a840406a7ecb4d043c9e4bf5ea6bc6e67
z0e598ef8bd70c1678388ba23f3446b0822df936176acaf6e8d76d20b278cb56573b36503233ab7
z9807af132caf5acffc6c1d6529f674793e08a76cca107f50d50fcf762df8822cb91f669400bef5
zf7923a08d5a27c6abbd9e793d0009655468be9fd67340a801cffa2f7ec588ebf51984a88be9e1c
z9f5eaa6a672f4e7fb260532a2e483cab6a66bc8971fb83b7129ba96bb2801352f3aa1e9a5a385a
za886e35da561dc6c8d81d5203b0c524600e4902e2c3129519dbbb8d5aba5e56e11a43c9c4d1dc8
za23eb56d98011c766cc9f100e70d9f05ca98b5f7f98ec34f1f348066ac14586cbb9bc5f93ef038
zb588107a4c4b788e66ecc84682f5238ecf8e7417a9e16c75fa19fadf8e11cd59b057b597bf3189
z48cdfaadd0fb4f2eda5bcad45390232ca43b917940236da8f2b49cb5a4d7efee145a73f9402c44
z210b1b0710523a85cbf81e14b8d9d30c4b18c4f8b2e7fcf2e12b4de5b73e4746091f91a1c2d9fa
zc25e789f15a94ddbc969831fc552a1b97d484d9f4f59a34c8acd868a7ca020342953a2be5cc894
z9ff486cc0d64f080ba661cd7cb1ab5613dd132f5474721c63f7ee1c47734a69719494234f4dc30
z72a552263a94016ef5dfe6805bf74ba3783c4293283ca531d1a110ad3e1f795fe1480b52704f4d
zead19604668e48004344d36502578663ce83dfe9a8813372e6b684255ba8394558ec31efd1ec4b
zdb7e05be9d5a2a82b3cb716c4c8dadaf015787ab16471dc495fb199caafabb60b4a229b68623b4
z0ee2bd8fbb35e549309b9670d941ce6dd8df3181ee6b974cf61795e74f77172a65e5b544ac6716
z477adf943c15ddd1a8c7445a6b5bb5f6d7b2055c09d1fb2420d958ef3c414d61b016402dc41d5e
zb9f3eb069da640aebb14469970e61d0b91d0d78cdf6b64c9eff04332bb4c1402f8422b43e5baeb
z95d2fe5355e4477d1b35f3e7cb6bf0d7744baaf248b3e8d0769fcf2680fb57402728460b97c6cf
z98d3c25b54b5e441d208c2e7f0bfca49bca5f2e67abb71f3808ae1b2c1db4089937e280dbd90af
z8c6cf818ca836df4bc851e3393cd617598eb35bf0b9a3ef617f4da7ed8aa9c94f03952ce3370fc
z2ea0e996ce5a25e1383a161b0313749e645762d8c3b45f66b3e4f20da3e62b7078a563f9e953fb
zd01ecb1ebb71b6085f1cf7ef4cda7e61ca7a2972569b68cdd3bd93cc6c4b03a171c6a881bac7aa
z36a32b3a71a90ae1940d2eead45495eeee9be6ae97c797396089d7bd0884c6f88e2e03ce850baf
zfcdc26ecf298c24a68d398ebe8b95608b494a49c57b9eb8ffab2846893def87d6108ddfb339554
zc56fcc1c4b1709d74c3781499fa61dfadb931d220bc469b24aff64b0535a0bd801b47a61f82a57
z5449b6be6a6d99ae06108e7fecd551384fe4b1548e744dac72027b39497c207d45e9d980fdabea
zfc0ebf114100189584e53353d7d8d98804ecdcaff427c924a4d5b160eacc2e147cdfd9e95f8622
ze334088384ad5f17a0fe57fd863193d94757a3695fcfe26f448d142427948dbaaf445cba9f86bc
ze5a309cd3d1ca9955cbea4cc2e5dfb37bd5b8aee39a04f5f1223e3f8c9ddec9d50e1dae6507cd2
z6f6320207e83ac018830c8e07dc25c013c367a52e0986d83b34b5266194e701f5e1f62f53a3606
zff859b79aa747afbcb3ff0dd13fe8c43d9256a3428e1c4e7762dafb934a1c9ffd4891c3866a0e3
z5b11180af1ccfcf003d511b5cbf734520b1c648cd0209919e8874c32d01936fe2135fca2361d2a
z5e8a3d992ed76dc22a003e97f27391b2dfa09d87e443afb0a37055127944123b6cee0c06c6b6ae
z72a7350134f8436363059404d4da1da4cefcc9cdd4a136e0813de06ed9454d2c61ab78aba75c84
z8abfe9e18390446f65c4b8916f90831dadaf37e19f54c23ba5de6609daade2a79a896a2c5f55cf
z67902543ff71af5c962343e55c4b754b38121ac8e49da74fdedde55739a527e3843ca0916d9fb5
z8cc6bf768d6a78620cf1119f998f563adfa8f486893b13e88d4341e21ca93286783cb22f1de3bd
z40789002f7cce17c200e3d12a4aeab18e75180c86391991ff98dc9fa9f86985f5cb15a2f5da263
z18f1d83b9e15cc2a147400caa84fc4344082606bf90e58b00bc60d27f04719d32d8e7dc22006e9
z5c42b301ac88352da9ed5393a7f3e62b129850f0be6a2cd065fca4a2dd5a2263084b613845e6f6
z4b033f1f244f0904e537fff146d8fbfb50d3c99b824b0092cdaf1dafcb550cf80ea94a72583b7a
z87f248de24c286cd3163a0ece88e1200820357707f112d84f76dcdc21264d3ff4d43987095a751
z71499dbc8304dcfb1254b87b7665f56f4b7ae04ce0472734f13af345004f7e97179e8126948be8
z4c4f795e8568d8b6acba2212a3baeebfe9254c187f2573cf7f07b6f5ddbbdfef93dd5dc5c9af02
z81c9e31de41c29d0abb6a6fe2edebb1cff8166cb9d0d8fd4b8671d5015414d9257e3d97c2f0b28
zda5d71649a7617fcf25b7cebd5dc75c883418ecd4efe369fecd5abb80acd7c62ac58f88e4fdbfa
z77740485234b9764852da747236f2be8f12584ffe591b9179f146bee6333be30a0864f1fd66ea1
z3690d64145c0f7c0783211aab4fe377739e2db44fd6856d46f00adf448083efcf672f4397b66c6
z17d1a99c52e4234d0e0a7a8879a496854c58dca7e13003a3513b8d31067a0da5774da711c1ff71
zb2223878e4bca3c2ae004b22c40306fa43f99a32c56dc5f397ee11546af0f1ad582807f4b92419
zd10b1c98b13f51867e58ffb0fa5f0cd6b6962acc1660b8f6a9db9260eaf37b643b0e037b4c6c3b
z2ce2ffeb14074972170b43ed5f233535692aaea84f34db50d8bcc0ae359189d55001d053695fb8
z9b58a3d6fe17ae798f36cea3d207b9950fd99fbb9f90ddc0f2011464e5ae6ef9521a2ef755f4cc
zbbe1c101a6f9a1580214642a41c332ffe52c8a456e01d7e57464d816919d55bc6499b0381c88da
z347a5ce5c3d70709d3387ca6ef4c8917db953b05c14ff65663912ac300acfa3357af2f203f3ba8
z5d872e155e077ae23473597280b9b2e1ae53072f33ee61bea8ac3119438ae1dc57042c28be5ed8
za05ec22450ca89cc99ec3d58d269d9491c265e8acdf4e4409f4392d338fe3d751cbf2034ce251e
zcd6d0cfb2214f7aec583ea65c790ae8bfbe584c7dd6ac6f78ce0caaa25a5cd6c28f2f7e21a239d
z63337eb762e932684dca00ba2de8c47e70305f7745a76792027941462a045cfc18a877f2a77d68
z71f968a19336cc3bb78d83380bf5ab4a1fa0502b82b92d43c129b1e8be74c709c9f87a5edc50ac
z723a8b04e6da859b4b96bae2ea5f95bd8c36ad08bf9540aa94964062c011ecadf430a29efa6a59
z4b1b14840073ce83e299bd8ea2d44f734f61572c4de110b0e3a16508641a24dc9fd7cec636faa2
z931fe89caadce0d76b95c74dbb8ec73e437546ab28893f2888df192811fba5fbbd688e843a1f18
z5631feddc54febab847a7fbd45160f40d8c0b0234ba6d4c258c46b320824e32c3cbe6579ac7ac7
z72457ec35df641f93fc84f35f8f60686d67ae26e223a30af4af4435d60fd5206abf9e0a765a54a
zfe3097da9bf429c79751f11952d0c0fc9de47ab2c83178b805e8d05c885a7aa340ab6f2d35949d
zcdbd9a4b6daad692570a8eac829a6db781c4e7108a4513981e92f12ef460569d9c8078f3a094d0
z0d8dfcff6022b88336023084b60af0a9f8d826e2d7f078ff9cba939c99f0b59cc9a0744a0e251f
z268e1bd82d3ff36e54de7f2529eb951e3e2527aa527d8733f6ea1b2d744597ac30dd18e56b6525
z0f35eedd9558ab6b11a7aba52a0f01e1f85da8312d1baae3f43aac4a4f06da239fe20ba509fec4
zc5f4566051ba978fb31c07b13a78e31780a1eb8f60fa29bce47bc3e10c6913bf68c7dc8053ee71
z9e4f73df950a459c5d49326a0632f384a427bef0df1311acf3a692eb20b5e0d5964724314f41a7
z86e98cea2e18874606c76a17aa83f313ee93edd937b3b415bd8d4c835dc61f53aba675b6df4ac3
z1a7610924c9e062a282a61d2d911dfdfa5fb60e1dff13bcbdf858aeb73a191df6b006a1c1887e0
zfbb7e9ffa707cfa9204992cba8e8743449d4b3067f639569e1db7b751a4e8938395b8020f31404
zea2e786ed491b5e0e00bbc449ae0ac4b9b7fb944399fbd7316994dc81bb18ae65dc90ae9d0f421
z05b2a9641521488ce85cfba38d0ce969a57073f4a64d59a2cdd0b74a608946298350ebd20d823e
zca70a36e8cf59c429fa8163fa45b7a43df1fbfcb83f9264af88983ceb2d3769e1b962eb55470e7
zcf34fb1e4a7da0683db3fe24f8a81b6139484c0b0e2ec678a7afa544a3c9f40c6764cd6b928130
z6cb7526b7ba2c54c893d0c5194c12ae28f39949b1e07cf9210fa92ffc85355ed87f895c953e500
z22af2c38172c107687da0299d3d504149982f69e66f657a55fe46f36bf23754b18d4e68e3cd870
z8fc69bcc6860e931f055f83adcd4ce8c6e8f7cb65a376072eeff72a0178e92dd58c27fca558daa
z2bdfbd05a82a4866c1143fedc962ae0018910f065046e08c638c0abd489b18c16bb29ba84544db
z3d488a6da68ed4e9552ccd252e47e7f1252f0f6123f89ee4763df1f1a8fa71c6553c5c5b86cc13
z32f4150c91825235ceb5907486b4a2484f96ce4cc25b32ac8361e25d9aafe5aeb6bbb2d6cda9ef
z71019976d531d61eb1ce5f51c763221675ab618ed46dc21fe8a3b8b60ed32b79c2ae0fcb5db939
z27bb2a6ce769fda4328d3de50d9b4d8b3a45c8ed5539fb2e47ef7684d2b1ef37157f9f40bb1299
z72a807a1a8502912a62a728e40a2d8b7932843ef451f7e6e92631a1036977fa45c630bf51935e2
z9b453be08c59b542a609a78281fefd2d9fae871033117804727b7a1cf24e5da6981a793c47dbc2
zc64686faa1ebf7b22d50ba7d6a2653836a3c825c1340ae722a68fdbdb74e6d2a6088c0cd9b5822
z7945af218c5cac6cb8e77e35bf3617143cbd3bf5d4f0d2f4b8635e8112c532c5157fbe5f205d5d
z1dc4e5c4ceabcfd8f9776f2a68d68a3abe88495b45bd4d3c4dacbb92940a7b075511899ea920f2
zc7e5c2938e0774c69378bd8238b1b299122f66e480682f4e0e2fd90a6199b206c696d67a395420
zd128fce473efd0f45c70f81bf71d5eea81df0c4a07ad1ddb01d7c91c7367657f29d99a3fc6e9d8
z1256d5bc332a9745dab8152ebcdd2cc2c7ea14eac6fede37f2db04bc25f05a3d6907fcb571c54d
z0d4414b36809041617cc57a64f73350082feed9e34e86514f690aa8c145a0b813eccc64cf27f73
z9b4c42119ba98ca34eee1f88129ddec4ff0941e4dc0b2a0277f760ceae805a83bf47c78d324c1e
ze51473abca2df0e6a332a8bb64724cb7b6277e5776974e3a6f6f8543299263e88b865e3b2c2454
z1ea3a7221c17e79ce46f4deca649062abf664fe26ce8e47e615608739111b6c19fb669622ac0c2
z8769506c06cbae66a276381241c80b2990e42d140056698254c0a453f004a51e518c9f00e76dea
z0b7f8e7f7ba85cf4d97bc0800cb02c8e41352d29321dfa098bc375b95fbfd1a913cb56ea10d500
z720f6d7049614a36369c1c70b4228b790ea068cb73e97199877c1fbb4e3444c8ba13a5a6b03153
zbb41f2cfd13970f4a5f9991da88841a6d362bb9dbbdc0a9f85a7a9ead446ba612453cdff66a46e
zf5de49e424d2c89172aff7ff7c8857555c5ea9abb7bc7f08ab01498388305fd7cdf98294343301
z83541ce9cbe77a80adbf00e61462389acf0bd044d90ba3e573a28bfd9f2ca213477270cda106b6
zdb87ddc08bf0be14d5ebe589095937ea49329f49505484a02db78eeaa71ee51c91243780db9a75
z632d8abd632223046ef000658a0f3974497d5d50097ed5f19ec11ba5a4c10e5460eca4ea22cb31
z4ef771987ecb60d403426271edfc75c3d2c71ae560b59df29f626d3ca720ef16af59c6ab27d492
zf14f31216fec1bd3c48c654ddef3b774e043b91a7eee6ef8ccfd40609e36c66929627f97632a92
z78b4e5ae2a7567f8c83b66449902b3620a99477d3d47ceff5c19f079498dad93410f6cb3eaec1c
z97e10958effeb5518d2e0c48014547b7ceb057ad80ca10fb481c592d27aed0eed4f36511947ec2
z9252821504daf78f11223a93e3936cd22080a7519dbc5701a861c32575ac80256f7b9dad79821d
z8735e297b334e745bb44fa680ece22203154e763b7d9c4f5e66f3f940f98d3ccb354ac77e5fd8a
z97d0517a24e6954940d27a72d21372439249cb1d5fbe4367c8496a0923361472d39c67ad26c31b
z1209966f252de4a8c706d8b68d36b8881c5417cc41fe084ef8556ce6d2734dc7031e7ae7d0c32d
zbc9ce81f3a89c4351ceb231664d04c38e9878435079f115d596bc499e065b0a519f62dc30289b3
z2cc6b7bb359e620ed4dd6e1bebd11e45f0ad967715666ff5baae7bc20d8ec75f20af1968e276b6
z422e3cf5052f8ed34991d6262e68a2f6d7e25922936a0f7b8488b63029ac3bb59a9a168ffc18ce
z98e3f244d0ac86fd87340b8fc41c10a44857665d1e1aa3a7f99e1a01863c7b44bcdb9cdb2c3984
z04a52486860695bd4b7cfd3ec67922d2b7ee76510740e59ab0ba8c260838155912ed26c6e2a94c
z5ab72965e9a9965293f45eaf78a3d37db6d89149dfaaadf9a4bc11333e9069c3ff9cf654e299cc
z4ad426ab21eb97cff2475f5e5ff308e0169fc344790121e4a41bb60ac2e77a94fd931996e0b49a
z8164c8fc1735bab9c6f109f8d1276008eb1fc14b7e60928395fbc4006efa7efe465075f7d94610
ze19891b642f26e2a3b070793d21f7832c324bb4f7055f43f2972a549fba13d6652731f62d17008
z881bb05799b20eb3b9be235ed693b70f235f89172761d2035dedc42cac7e1ab5abca7891be6040
zce87fedd870ad5071f623b138a30e35ed96164bbcf566245ae00b303f63eca24b577f40a251976
z320da7850da00b22317c4d25b49f633982d8eb21cc7323c244dfe3fc5326ffc428eecbb1e8528a
z610c4d2f5d96d752dda83186b6ef2870200c6e61eefc0f9b5cca81882e9a2f2bd1c5ebe1f703dc
zd62360563b5260634d20c0002db0de9787bdde3d8b60ef24a56bd1d847d0e2c150bf0c32706a10
zd8f25b1d27a705991509e311927fa56c910edbc29004929b73d8636a85df61755d93725b43537f
zc9cb82178ef9fd9e58ec604ff12bffae9f678c50092a87db7b56ea88a423eebc1e4dca525b2dc4
zbca809e475f012ec80b617984cca9c923db087ecf3ff05adf311f56a7d8914b19f7652f7567abb
z988f10c8a41c8b8e04c0128418de94273692203208e17768e143ef447f4ca715619833232418a9
zb7502db0d85915cb6119ff7f2f4c26a6f3530cb220087894ce72499d2803b512ebe3d48f7ff32a
z31382abb8eb796325a2a48a07f528e343759868a71c714c18f8326946cd07af2ecff6c99e0e782
ze8986120258e3ab9eabfd3fbe77bf44b3d871e6f82b5298b6291804118dc595e3f7bdf781c7040
zfb3cfc86a176732efbc5dd60ca5ec3288cc5ba8373eaaa9250394e94451bad423ae2c1ac410b37
zff0089cec1e46351683753ba38d98266f88170f6476122069bdd195022e4cd65a597c95f3f3d57
z23541d6064dc1f8ef054b9e827882567966144414cb550f9692158e774550b3c9e227e1d73e80a
zc95e0b22c8d760d572c819dd32ac33b9905563026053424ecca30318affec99c19b9b561cebaba
z786c0398c006ff1e14cb290cd84d9a0af0601b9552b5e7c5ea08d8efb217b0e08e5a93f66a12b0
zd26608e22ad935a0fa0af8e114e1ff1ddd829c4a14607912d3be8673a97f62eeda969714d1a9e5
z1f453fa05b334f43c2bf11524b5054c4004d5487b414c6932c5d7140432186dde2110e4ca24e63
z2779d7c2cf80149a2a44b9acee7671dfa2cd4264928e8876fe3739eb6da5706a106167902bc70b
z11245a368de1936207db9c2b09e6cea8e7ffc7457310c494b4af27420898c0da4301f01a5fc43a
z26e64844cf87aa4492b19b14b250b9092f49e3a3736313e31e6fb53c55f18a7b75faf6124cf0d4
z93b34b7cab61ae966638023a3056c352f84443f00049974d92d2ee3a93bb7f1e5c664793851a76
zaed37d4a65f484e4ccb4887f0e487bb42f40ffd4f7f65c61dca690487230c361e412ee5005fc06
z4205043e323f5b9a49434a2fa9e854dc73aa7e30ef09b5c29d340a3de543e82b732f6ba89f1dcc
z5ca2fc06fce3af2d933ab4b75ebc86a31d987cd8862e11023ba0b9ac4cb1d63a3133e4ce15cc3e
z59d07b28e353da14014f1234197171b46f4ec3a9392f0293d79316f0e873b5069bc34c7515fa17
z7194f50d356252d82093872e8db172325f1bd36f85a2f612bc4133cec2f04bd8431143257177fc
z6743e21a53d35c874fb7b1a4267a52632e6c802d7d6e2af4e2dfa565824e98a031c5af8f0a87f4
za89db6f9105b9ae5f69d9aa281016983be611e19828b4959fcea48a633a03a3469e5175b4eefce
z6240e590eceed103ca41603826969b34ddfddb90694a491ba64dd91cd159e52bcd037e3187dcd8
z0d6a717387cb225b685ad26cfbb52acb2e26c38013ef33e0741f5a5b809ab5bc29e338e9cda384
z0a6bf72aa234ce8c1ef791b871c56cfc5abe80543b1bc10b20ebcbb0b0420d51d70981541e1b76
z82a88306f99e80fa55fab9a02cf26b1d095736fbe7b86de3da6c6567a6670134832a8c03c000a6
z6af2c58360f9fc8491867e74fee4ac9c39a1563f87ae8028d906bb406128bff001184b35ba9324
zd0c19811dbf06b97f935c3876f7577265637a4e103b21ab3e089ce2e137e2bdf170d62eb22cc41
z81772d149764d5146e1a7ae9b0ea23a822d5a175bdf043581b874ac818df1d43e87903a285281d
zf5f2478b946c13474a43992d94efa3249a9bd95cd31d12996d1d71ab31a1fea31e3f9406e6c8d4
zdeed70d4f6dd5a6352fd43c327d283470f58308bc46276144bf29250aa0aefad66f5b14d1a1fba
z160a0837a44c05080c56e362445a94feb96ae7581a854428a25d84602c957d283d6c2679cfeae8
z866719e0a02f6dd81b27d829db39180dae5d1b4005e9bd8d39bc81489b27c86c0e07c722b3efcc
z95e5ac1232d823789dc28b67d12334972f056bf0e049a7283179a901d4f1d87293c63eb76463d5
zf24d35d583c5bd7c8907d0e1c84fbb3843afa2d52b08bdd7398b9b6842a42caa3896183b130376
z2dd628dc5607806d79d2f7509e87e9899e5cf484ae887af9b2cc132c0d69a4714e14358a18c1cc
z1bd1201af51b76e8d544502d68416d2330fda1e7f83aacb7b11dbd5f08e085dc9aa077a9cdd359
z6f7e010595a3590112d51e45dcfd66d525f2c6ce39e280da3ee7a27eee6c0e2b7c9912ff4c2b30
ze6e5f1e111d5e1514f8d21bd8bc671077f5ec93eb2170d79b43509bbd06876faf4b971a0f35880
z84dfe6c9e7bea95c97fca1d483d3a46883efd767739c6b0cfa26503aa5a8f51a96eb827cda527b
z944b0d90c85f7dfa692f94e75b9465c950aa44840062c58976d813554ad120a0a158139eb54a63
z3497cfb2650b1331265e824008e90ea09d2fd957133a54d522d93e8f6b960423f3a301b9383e8d
zaa86b8e414be62fa0797e8ec2295a4c5566617eea9d14e2af14956a91b97c32943dd2baa9b8857
zfaea9f96504545e80535932eedbd095b1ee8c419aa8f73b79ec6245312bc2ad82f79a646f5d3ed
z9744ee33ce43abdf5b7d32ee10f7ff5de8f558b257503546edf3e2372eddddbb4c2bb2c9df57a0
z33ef9e533d3499fc35dcb5fb9c43f29057aba553f86c9eeafbb71102494fbb52c8381926c63e7f
z9b85d68c343b1afa7bc835817efec5029d0a33138a7569570323fe1fe38b0df0ec0e2a2f16f023
z7517c0dd587760fd122ba766b4bce2e72447000101a87d8b883dab577b2da935e43cbf56d495f1
z06cc1dccb87b955d763089ed7ccef94cef556a15b1680778aff8cd55f91da40d15af0c9ebf4e41
z854635a562850ee1cb979b97e7d82525ecbad40b783646cb698ec4caa6c74acbb84cc84ddca108
z33c2b1074498345f8ea3fc73ab8077df3c3a99adfd425f054c51190e6c6ec99ef7356fb790d368
zb253660816d2b1e4d4454da8025408e7a52e08683e9f3e4ac0998faae0a70ad5847a5a720c1c28
za0a50b694dd6f02e3965187fc24a4078995e3454420df22e5bb277b14bf1aff674df812ff081a6
z6b482c0cc30ddefa27c73826244b853b319223bbca537a169ea4da88d389b2a12f8472eff0b3b0
z792c4976762f94e49b7f1da84a8a14ec1a289b1f9bbcd6e2cc42aaa869c8f7023955309dc937cd
z4df39f99b33d2b0dfdf936c327558e886122bd321107c7fbd76bef3966a1cdd3537548b4d6a466
ze4bd1b97f254c9143bc90f11f245c9ae5efc7b11a7a28186af79a2782fbf50d37b5403e39c065d
z3fee364fbcad20858780b63ca17e9198a0959ed569b9d8e8a62b9b1774f90f63d04a87847d4236
z96cab741f391d7ce4c25d2e9d1f9803d8e7602852bd335a74d7ae827d599aa6016296f2db16123
z74fa3897ac635493ebe25d0af93f58c5e53d8f65540225b504147f48a2f753f568a60109d46df4
za96b7e409701c2a35d4aa9c171b5b05271a6a6925bfdf2cd3f91471250a8bdaba79f5fa2c623c5
z7b66375057aa36913637b74cc3e14657e10089d1cb669bd9a3ff7c519066a6a2a53964067bea6b
z979f452c4e176cb5a5e2ae04e390b66835e8b96df53dfe6851b8921dc85fae408f8a195aba015a
z1dcb5547b4932c84ccc16a78cdf586297547fffc946558f969239033dbd502f3f9b896f5e2bfbc
z2e71c10b627c3fa7c4b1d7783e4db54a1bacaf4e5df1e75db224a0999a04da3192633b5f1d168b
zaddfb3dd44e6a48bdb272a3be9fb27739703cdadaee06e34217eb203ad36666119bc7f1e53f713
z2bd533bb4f67efd08c68e9cab39dd0681447970147c8a287ca7c260e7bc9b4e5f2bab33d8ab85c
zb9efd7f1ca6e87f6877afc61971721f03fce87d6d447469effa3441cdb39dc256f783939d79cd4
z5ca773829f0911120a2367d88a81e916b35782112cc3d69f5fbcd4f1e1055a98a39bf2fecedad7
z191a5d50050e6e86b2799e81b7aeebf01a86cb1bb23ca3c06b34db88087e692dfb726d457df95a
zf10380939583eda958009486fcde838df4f2e4740577191a3c025416fc22f487544151c0c2efb0
z786b47602c41f7e8f9bbf88c611f03ec5cda81e1f680bc57ea2784d94353bdc7d273096d9acf14
zbdf1ca0ead58814dabc150140d73ef3e63832b608cbcbfe096f4c69c8e1068af7b81fa186d3405
z832a9668199fc975fa56ec505347c115120aca7c199b87e188f8b6e0ace9377c459776309293e2
z52e514de1d72b3d8967be85aaea5f2e1047669f926a3a05382c2fdd5ba5c4d3c3c1d27642ac952
z1679be433ebdea936823136ce3f35b94b82eac1f51faaf539da7bad59f72bbe3c36bc817c79094
zfdb1d6da3b2830a8110b088d5fb538156fbb69b95860256d84755a23dc57b353791478968fec74
z6728b5595f9cb2f1ae324efbe86b92e636ee20a505e72b47f8cbc7b157475480b412364ff8b745
zfa863dd7afc11ab86273250c4405032ee8af06f6e35f4a64a203f69701442276c21bded2af2ebd
z66126f0aaaad0ed3076890ca0c62cab610378c47fe8d022fd61dcb7909aef7932d01033bd02ca0
z9456e9487a37f369a827eb3588e95f08bc5c404fba973ea3d74697ac8e364865e958805fcbd0e5
z59287f4d78915733ebe79d728097311bcd61c5729b707bda65ad0e86038323d74c4ec98239525c
z3bd6a3ad80342b5b42a282b94daceeb8f37e53f0ca3afb735054ac0efb24ac2b7f77bc87ec9cb7
z150ea96b7ec03c73071d825ae82d8445bc82b5ff427692403976b521f4c2e4e81d9100e20d4082
zc7ce10d22e064356ad6b7ea2c1bef913117e41344238e5e8db9d79de890b19a7601a6e9f7d7f72
z61bba0840084cb2c1dbb27a9c9d250490850b1f2ee9f977b37141d98269acc2f24ce1fd63aca77
z282dfcabeddf89dbdcaf1d82961b2842348d8e9d0674daf7117d19d5b955f117c3d25332549dc1
zc73121f8880c706d8ff7da64403697331a5843fb6dd3ec4fa38db97cd682fc327b4dbbb927fd5f
ze96860d850d7f5eed1502d207c32c6b41498388e9a3ac2b50ba1c0baad62629f4f7cfada0abb8e
z0322f7946a635f760f4c863fbab8dc52b3b4eca49f4f044213112ddc5b4c09972b9552abe6ae55
z90a682fdafe1f4ccafb8e7b702498d3a65b765ffd7a16e4b8e1cadb090e0b8e849c0bce440fd64
z52687967ca2dc780fa95d03953bf5e81abdad9a2028b8146fcc4dc4d3f8b298fd817a5302ed8ea
z787e442ee65a70931ef17c9f5a29b1a00735a462fe7bef9197800c41e35b5c2a72bd5ebb6be6fb
zf658f9a26d51b1a22807817d53d05424e2949b51d0dda3996a258a5e689e34c056b88df6304e8c
zef50ceff1069e713b4cdbb15c12b38889e5506702f44492cceacf125be52cf987b629796d0d80d
zc03008fc68b4f6076225b4f6ffb4dd92ab244183c4d753ff303db6cf351469128b14155725231d
z5bc9b0e8532dd1a260da3cf6e56dc3aa480158fece14f2063dad9fafd2c100c3a57221f82057e5
za9a652145f0ec649a7295a856ee762df128b0e494959b4530978b14de08afeefbd592add165130
z8dbfe68734193361926c51c6cf3c825b4441e26b94f7d6f244c362eeccd37dd289428c3cbff6c6
z007e1ea488e44d584812d601725bcfb1c7bbb762034e1e2292c8f420c464ccb84268195fa1a4cb
zb2ff8b5dce4fe0f24f8b5e1a8485bfaa430ab5fcb88f3278aa599eb71add7b1069311225d823fd
zd180c8276e17acdce1568b1f8376794d1f827cde0f4a624301ece2281cc82d388e44f52a342f6f
z1fc9535ffe3a4af537418370f8ac51269c452e8d717f10e9361c72b2f57cb92f3dea489f0ccea3
z7a86b64c0c79f632a5b73f2accebeeaac6b3aa67729f00c78822dc382df2722a2f574f74641728
zf9bdd3a02965a623fd97f224d2f942e1a462a0e21c7f71f8a364b56947b133c0ab8284daa7fefb
z8d6d1466ec3d9e934bbd5590cf2b4d64615b874645f4a378be9043df353f3ba63278c785f61ef8
z829bf4b7c6edfab3921dfc5f9eb57babae6ecabf3099569c9c9c7647d7cef33e554f4ee1ff3af4
z254c233bfcc32dc4caa4f92fb6c526bec8d1883457edd99e6c1173b66d6a0325c56e6dc5709a0b
z02e2d177f3979717410c7406bd33c9839f2a6c5ea8c2ed6bc8a130404f335602ffb2ae3cc48109
z774b753a173b58080d15e456e343495986a806fbaaad92afe2cd36273730aab20874c4bad3d3b0
zb3a8e67ad935925cc17351c99a76e0b99ce1d4542a51db394781b96926d99862587307bf01f9b7
z31b0ee9d5a31bcbcc2baacec081b928241da1f561f1efdc90efa551ed3ca873bf590111d33be3b
z47c8f25c3665308a5ec83da31843118997862a7c60e78837d3cf122107b32eb573d51765d30a13
z5a5c9349204152307b47959088b017a95789172b855c4fea318b4d45843af3d46dcf72570e69ab
zcdbcc43a1a34b7c0c25b6ab2740a647929150bdb914dde4303808cf2c4d3b6facd9af9a3724729
za68a0d2c0eb2d4d7af0794fcfea730107cdcbe725672b2579a3457ec5cb13dc43c4fc4477f8ba6
z6672c8b012a23ef3af2be5703060f1dad672a74be805bd0e177d1181ede1392b988d7895882377
z15aeeca1156edf5d8e391a8309f961d3f940ea5b78d5c3e4e64f57344ca937a66a2302b856d706
zf4b0c514c21b44d385d8f7db1629a58ec725029e7a04356df1cbe373f1a875d55c901aa0dcbc96
z471f7328cb13b96306c7e81a7f511598f13a5153e684f5a0e4491d277d594365e024d5fffb3b84
zb8da9ec6c1caab1207357f2b5bb2d8c9e115f371eea45615a08cfcfbd892dfc911c0a6227613ab
z838a46c55351d8bc685d4f83abdeeb616b2011f6277d1777ab82622675072cd6766713c522f4b5
ze207b910480a727fbe51c656c9356665db23483f200bbe6ab9bb4b753d6c807cee8b7128bb3c03
zd604dbae0e16d704008ba94f454bcb76dd45523cc6375e3573d1eb8ce26311ba3deb22dabf67fb
z7cc71a03e6f1dbffa815cc0fdbe39cb187e7b2b36ce35147b9093279a8e9dd815740760516c2ff
z1694ed99bdac7b5cbe5b502a0ce834e2230bd01f0ed212f6b02603ab17744abd94982a33035b40
z58b29b8088f631c1e5800c0dd8d9127a99782366010d170efa21e5083b19e18c6a30466481b414
z40f254fe5134a778ccb46af557cd398d0111601b2c77f2cdbf83a678c34a1f25a929dab08283cc
z6db4f554daaf7ffbdd1f1bebb4ab86e9cbe17a2a203b0138eaea1a65d7dce40423f74b6babc1ee
z9b9cea58909ea61181baaf423a745da1ea9392e2a0424b452b120f08de184a20f0f031417dabf7
z817ecb644d81bed159f1282fc91c1448177316227cef8fece631edd63f62ec1225d0ff410aad12
z32e055939de4027be7f3343ac7e77abc6a3cf1fd737163669a9e0fbb9415f4084d1dfa15173e95
z4920b1aebe7099f53a4d9fe794dd7c231b9954183c9a6eb9653fa897a7e6f3293efd03f987868d
zef4e23e281703fae9ab05a82c5d4e7642f319a46b5f35510b8e999878b5356265bec8a4285ee41
z855d620d83c44b96e8230e31cec5e1c4c28478f491adacecb469ab6caec93bf35c46552351a597
z07c026bf08949afa5bd04a8c8fde7bbacb860c560dbc970f2e2ad95c4f7fb28d75ca4557d5f017
z424b6dbb744aca774af2421284e7348ae887cc100056e096f10b8ad025a5e26918f7b9b10f59ca
z1a462cd970829aa1801f78577a5350e2ff7b3e9ce9fa38fdad71a0eaf63741effb4e13f962bc18
z414de2e2e9aa556312d80be20ddc3ca85e11a0a7e37089be2682656348b44a9cd37c17186b51b1
z7233298e22be775cc045ce2af6d733f59914539a07dc001769c32aafc84fc331807b4836b66a0c
z0683a3b71110a0c1f59f2235413c3a27f5f408967a026842cc390530ae3013eef0ffb404761e40
z5ce01036416c02b1cd9ca5fb3268c80aee4651bac2bdd0fdfe9b45cb4b3a2f2cb79536803921a3
z3f16f18831dc3dae2b64015e20ee0c5b94a7069f83472919969468740af048600b5c9a7113a0bc
z698d0586062565aa652c91d4550a1a1f0d29d75696e614facbd6b3bf87f8a0aff2edb425f0b860
z43e27543e39aed821010bab34cf5cc9f4ff418429c134540f3b20a593e441f68cbd777f3761754
z93b4f5be84a42f4c2e6a5755fe3f063ca4c31d4d3a197dda7074ff560c5bdd30530bcf13afde87
z53665be58bfe5dce955098bc39407ac58cec148c57a654066d6aff7b1dc8998cc1c56274443d66
zdd866f9859cb51231177dc4b438d8a0badf3963b6554313067dd85e7157b6ef9dc9616a68cd91a
z092709ec4d649b6f6404018e4f5ee7f6da9749372c84d97d004c5cc44b04341a63dff087d8a80f
z46d73190e16478020cd8cc315293a8e4e873c06189a1f912797edb7623864f8c6924a4574316bc
z073f9c91bc487e78173ea69a7033ae9af61492ea8683b3d36bcb0f39c81afc59116893cfc327c9
z48d028bf7b451b63aad82afbc35e609fc83d10edcc87f86278cecd5a14479ac9b494d0ead7209c
z467bc09e66c8d84cee2661469dcf6b0f184c20f08cf753aff50e3cb00b4757eaa46e22d4295d47
za87104ac3f0ed8c7505c055344b1e52268ab23c4b12f632e3ae97585557b9c9a34206ed6827ba3
z8d145376b1d6186cb2717a11ad0e463c401ad1063ae6b3ff8f0e4ede9b7ddb4250b7ccd0af8911
zff6c34fd6d8cc3a3746b1401ecc8271eb430aa177d64c9d34ea737feef6c681ffc22f417173990
zb8ee0db829b062da81c1f5f177cae352ddd252076d32938f541dd701152c31fba5ba7fa75b1711
zec31195d18dbbe3b3dca179ec7d884bdd6d435898339710515fe002069cf4afea1cbb8bb744540
z5d37605299e7572d8f63881e619125cb93932b0575a18231af5984b2a748ab49058d6385045ce9
z4b0f8f11fe8ef34ce6449db0a91246547885ca3a522ef1f57331d3c78f3dce2dfad9b8fc56e7de
za388ab075e384d4e61e7e0fca3352a24f6b95f2d30e55a55befbfbeeebb39bd896b85c5aa16c39
zf1fa4f66ca576a27e7684b365990086bb5998f78c1a0fd89837bc3e036cbe0b97143667006f842
zd37298363fe2d8aeb768f1d9f521e7c13e47c0f2fe05eae521710941ca09d1ff3efa980f0db042
z01bac149b94f4f174328b3b25f609e181b44296e105e67ae261f357a9f6e8cce209e4ceb88ac05
z9dcfec295525aeb559e77b283396f6ece057a79e9448a43e677df704e80d587a6842f58aca4ff6
z80cc6b90cfe402fd129ad66201cf0ce08a90fd8ab927e13242ad1807a01e89a27354aae5491b30
zc6706f209a5858a3f60ee1d80d5d3d4b6ca04314007e6580b13da9230f8a4d7f472d89dabb9492
zddb2a81e85c67787637131451640627c44172e33c7af2c6bf93fd846f6a90180c97b9f87b93b16
zd75d35ed4e51908977f5c52193c89eb63f7be765450bccdb34ca74daaacc45b8cae0d409863ba3
z40a1bfa95e12aff510fcaf8a793c8314aff18c5925497a66eb656c86db8344e7e93b6c76dbfe8c
zcc88a52e7b2bbb89daa409af61848946182c58ed38b906b132826906105f8ad30417fe4911e245
z1394240b41c4c7ece0a71580dba0addd0fe58cb9451ce8bfb75cb8d70dc21cb23bda8ef9167468
z61b936c944c3252929f09d0d85b81283532b78a14657e6229077b4a81dc9e2d89541443e28d4eb
zb2187e5c66c4da3c0ef56ba132f589e11a8567158d031540f3193099dc564ebd33b9753cc5b04e
za00916bf446ade6885f0cb82c497813611f731a88f276e53952f98f46b56b91a292384843ad3e7
zf7b5e2b2afbfe9bb5d1a6abb6d21d97f1aac63d9d3e9dbdc8c1a7731a31b36096824949c1c651b
zd4ca26b707ee5f6acaf31f7250dee39873f8b27eccaccc85cd1fd789df3916807b5ca74af04a0d
z2d1e9f5928a1297a8eebab5ac3f46d0268e26ee4fcbbf52bb51cf5dd0a477daeabc886b3fa4065
ze57afb53fce486c3d80dbcdbda4e6d331b9f859e2d2cf37751ab045f15470bc7dd14a016bd876a
z9ebd8fc23f0af9955a75d5f6c7d3213cfc9695cc52fe2b0417e76127cdbff0712e2da65e13a3ac
z112d0644c21a086cc4b28b607422a5113401ec609c9226613e72dbee28c09aa0838d52451e6c9a
z134226afebc4090f8bef99bec4cce415842229fe67a288f680e5e96c3dab7271a5321fa0e3d3e7
zaef1fe68eef38d82a5713f5fea6443ff8241d770c3fecdc32e216a77e029ec78ff437869d1e260
zed0be0c7cdec358f493928cdb6320fd4a0d994c5842dd23c8fd8d36b8ffe3f0ae47172edb47b60
z0e38a28690cb6637e65857717c39b12df621dd6d395348c941da8153727be37ea416c3f6219549
z9b835e16b44251837ac78b89190e62bf335fe53d0622dc4ce42b543cc38c69be656eb4dab50249
zaeaab6ef690423af9c6798f4a3a0032041751abb119935713f245a6477a98d3bfbabe869aa7ed4
zc9dee2e17c79a2421ef602a7e01f913719ffe62f303fcd0c3dc0f8a46bcfe796a33bfbf1679f8d
z4a8c17cf196ba1f3f11cb9b761aca44fb38301795d0310508342efae01bcbcd5e8cb3769322b04
z565f39e86fc7dc505c841daa8e156ea0fd4a95db73bb4287e4014627f7b03aa1acc690acad8db5
zbc972a735a2a32a431ba617d28e6576b6c3ced3222ad7cedeb2f3fdd5e4bf80dff910a79f70462
z3fca2b92625ad82d5333601be07c69b897c63752eb0a37d141e98ba54ac3b073313c385e5bc892
z13703248df8ab1eafae2a9ae65ce5ba7f386183bd312c603d4c1fc93e71b67d0ab6a7c7ea8b929
zece567f028d93d86f44e361621008d7046d4cd8b5cad783b7d1512f3ece7f8d77ef3430608ab5f
z9f825bf933a5fa2037a979a301446440b24493138b7e7fa9e1a9929963eb90e1a5563112b2d244
z0d4c5933cd2b2b4883c08bb0db5d81768c1aeeca5585c12415197bf416bed0fad90a1db79c876a
z74c14af67454ef6d483f2c9dcfcdd31ffcf18dc9a5481b18ef0ed12d5b47498f72df7186e68027
z4d33f5e26522fdade3445d0af69487b49abbd664a54a884943fb78ea4613503ee50114f8433f37
zd1fd586175ef8f2f1dc912729b5c46c80b31bbc2c1d7d1cfa2f4483d6c8fc98ce18159ea5e6709
z2570349fd9a1612ef0c08266685295e04e4ca669c630e3bd6a4f8a4258f1ad3a48a76277bdf36e
z325413e3b4111f4ed9509e8ea2424df2a97f3a67876d5fbe3001ce669f0019d494532224ea23cd
zc8cdb675c0ba6979571b5ee4795e92f7e3eca635c972de06c91ccff994de3abd3b71352edd4c94
z32e198e738754cd8b4257d23a36bb9fd441835e240ba4023dbc7b8042fbd014c2aae2eb8e29112
zc55c10ba958eee052e3329965a33b91f39b66e6633ad105b4c60b1cad91d60874a2ca3a0576f4c
zb47780709edb84a8ef6967d71656c67d0b0527299bb642818c404e51bd29c0cfc5762d8b48cb5b
z7491f510d15662fc91fd1185659621339a69866602e628ad0c8b3de324ad046735677955a87a45
zf739910a6b2621af76566ba38d13379b94bc858044eb298116b4442dc7b2161bc173a832c22532
z297140a5275ad5bb3b191dbc4da12eaaf4159ca77bf4e9799c7f60d35f237fa43b21aa47a1ff2a
z00bb655b7dbd374144c1d1f53429bfb1f6019d17d149b154670c03118af5deb052a8fe2716da13
z40a474fbee43aa969cd02c919f9297bc3ae8751a4468ba2410c8d201cb59a55c45f963978ea9ff
z7ecf0216e05251309e15a69e412afc7fc193aba92734373588a4b1375a1055811daaaeddb7a960
zfeb5c4debf8985d2959fbbc826612a5870fed4445f41446632610f2a1bd37ff951aac782272377
z0061592f69783f89314085aa3433d5473147fdcadb567314385aea045f119674e0a236adae3f86
z0971bf04f306f4b0517e22920dbacf32d9c8f1cbd5ca39c7cf7e32b23c570503d8662db7807827
z58c93df698a0b8bfbdd69b6c461da0c013a0dc95d6619252a5f7f1224b24c4ccac94c17526873c
zaae07a7f53bf1622de6e7b2851d8204fb09a9759ca048736af2e4727100a82a9a42ba7d1ac7843
z0480d23dc478ef02e87cba5f4fdce6b678bdb810b38b96fa79d03a972e16971127b5b40848b473
z090ed40f9f327803161151ec77b459866416fdeaca0fcdecd3e02ee646c5fd0abaac94dfa7be7c
z07ad719035ddb26c752e8c3c229636942b81245e761cb10997f0cd4ff7a9b0d2af17eac4f8bc15
z2008f1f5634a4db03162344ca320fae0da6b0ade062a3b3d348a41210612ea058353bd72817d1a
z56ad648d9efd2dd8b821f8579edbffaf42b2c0e201de9f60ced350eb99ec8522fb7c6ab66f53a9
zac31fbbdc542feade98b336484c5b380ae8204462dbf8adde42cc517ba17625166ffd408d4f518
z4713e3cd3804c806fb6f6e9586e858a45b52269a9ae98b794e5f52b8fc4b08901df2b1e89601e8
z9652e7047628859f57db228f93eb199788831a12e6c28f1c7cace79936fbd836bf5afbfc19f79d
z70db9a8b074ba742adc185ea8f0b18183e540b90d441fa583f9c4adb125542662c5514fc5ec1aa
z73574e4449b1ecb49a19099bc6f377e2fa5b9a7471779b8d72877cef6d8fd9e64677fb64bfe0fe
z180750b55776789622aa27368f09c263a7bc697f4a9cbdaee9e165643bd719164be839ec7d8d26
z53a548c14575435b35cb7651b58b3de4dc87873826bec4d6532268918115a2dd3656e444c7dc06
z719ea089100739c57b8073e387e67e5765fd7f9dcebfcf936c3581a22172ab77974a4ab959d312
zb796c40739c513206970c00f8b13270249771b58c61f11ccb2daf55649e9329600bb569cdf0c1b
zde2f21ba0b293a8fe04bd657372eedbf693df3c2c81e018b66472379e4c931cb2731cd68b6282e
z3aaec8cf5e33754b69503f347a4d0964a0798bf90538c780652ec84d305cb8dd471f3cb0cacf4d
za0300167e935780cb40fd4968080a7633575b6d5fe45465cd20db0d6e665f77f8786f6489f665e
z4f1f7c03b6ccb456583729a322ae624aed64c90dca8abc191d0c42203e5c56f7303080e76a5919
z4913830e90b255a6b169bcdf47b2cf316dff83d08ee27a06caf216c32fe986a2b8e8d14d76652e
ze907952ca7f806a91f32480ff10839dfcced21eba3972956b159e48b3db1acf2f5476bd26f36d2
zb3cafb30420b073e8f42be6db312b25a3018226e47fe8f97d1b74a8b07c12b01247e81e3a22bbe
z7a02553564b55a0def48a358132dd6fe229e68d7d8af886e617e48027ad6057aa9f8493cff1c26
zbb65dce22f021385c3caee4894619fbe75b099c85071b602820be310f431bc73dc359f4f20cd31
z9a32d95124fc0c8f1eea6b173e2fdebf2351af31f21f28671f076d6a2960558b6d0e97847111bb
zf79a876714b3eb41ccc130b0f39666fef1b7c152fb56187bae82f978d3396866fc80a159c4f874
z1edf00f161cc827429b0710bc5cad6c8d1416e35aaba11fd4f83be43c8aaf84cb5e22ac6e8456b
z8c831fddf870b00fc061e56a85082d95cf3953772496b4b3966417753807b264dc052245a1320f
z9099dfb97e45c961b7bc094fd87a01b93ead4e420e8b2dc7574c69859c2a04ef804f7a45da465d
zfacaf503805503da0b37d25b7a9c6fb7c57eb23c1a187f6bf009c06c57d0e24bed2656817ca1ec
z94383144e4fe7e6bc24baf9c53c64cfdde987dcde0280e6654a03f10cf00192e8b1ebf7007b4fe
z4238d0c053d4ff1d1ded40552c8ac9e10813c62470d52410994ca9cea9c9fdbf3ef84028f9c8d1
z2826e685ab565ea83f06451403795322efc33245bf365ec2ba230843515f47882978642053c719
zb9b8fb0c55c2f1d249209376e56e08166817429735e4ff564f820c02bd861467daa4782b787d06
zb704cc26d52e9dd2f910bc2f47bd197330cfa38a4050776ff5a6989a88b2005f648ee9e8c7bb09
zd0f6618021d34021d3c99e7cc2102c07ba75db6e405ba235960f8ea1fb38c48c8947a8afcdd5d3
zef13f51d220b964785bd3f4afcd3988e239ffdd33a27bf13d726a9f5497557b9b4e612b8007731
z9822803e13c0b16fac84f08d6b4fc29e2c2604df14c2de612e52dc4433761cbbed79902bfb30bb
z0e95546739721320498302a5081a6e2847ad065d1e4645d9d36d321fa5508ed8874a941ca62b2f
z92eadf218c37873b3784dacc328b2d062dcdb8505a10633ed65b5204a4d6b568c7260eb192aada
z2c5fbf1e2f0ecb5f7cb6db80dabe85504c43c29fd56524a4b4e8fccbfd48c82ad96d309f8c0b75
zb38a57622309c9784f4510f159331d61d1a6805cc6c9751879237cd10de77c60c92d24cb08d049
zcf673cd6c7285b59f55b22c9697fc0e071e0dbe0bf02f8f5fa8b0bf8520d47543645bbe1a515d1
z0faf9792210e8a83708644e29390cdcc28ac85c9ba6cec97e6afdbc60904e90eff6beab46e3389
z0448a8c50f084887bf77f5fa2f8e9a1527d97f4dea2fded96c4c47308e324b8549d15e0c593577
zce9ce32e42ad9782f9468fc661e25dd4030f2b9ea97caa09e3ec561993fe1ea56f6c70a2cf5884
z1f454fe351ab02596ffd3de72024bcddff225f79d0e111fa3a3942f77c80baee637e7ce5599c96
z56d1467a935c4ebf60ad4a887c3390323d3154599d3a848fd497b79a1e6bc6c328378fda4a4828
z89d29ca8a5b0acb85a97b4477dfe754505670c22341da85b9fa662c47ecb6dd238a09cb5b5823e
z699bc616d681855205ce3e7e94a3cdd398ede9e48fe636d9abfda00703d977333d1aab5330b57a
za1f2b7a51215307af9caf53e146bd9fdf5f324fd397ed958787250bdab5db962ef066b92f01866
z98db2b6d044b829bb341e9bf9d4531a60755d1e1c1f4490e92cc17394d68e65b5d1b1580dbba51
ze3d57af774059895c78ee46acc86618ecc72e367387dd52cfaffc65762defa2f2ae37f50172b76
z2d090f33bbf4198e7950d7d086234526dcfdc7cbd3b2204a04c0aee92228bda227a667f7c71092
z21ab46a4d974664bc7093662ff260cb86da7523451aceb73ff0765eafd2f12f295492c8d699318
z6c6fb3b3753db1db1ee5d2924f04374b774543f20ae1f09b2c2a225a4b63cf8c07e5cb0f2959d3
z1868497addb8e1471ceaaa6748d209835c0920c6bfebea99b4449650f76948590227791a561af8
z3ae827ab8d6d3c9c0f0e917dc37481f7d683937207c465d820984c5a8199545ad4417a23f5346d
zadfb3c61e8a935ada95d214334aadf41b645eed66b0a048ccaa1a0d681798d8235b8d886cb6670
z4dc8bb14f0fd7e1e545b3047b4eaa5dc95b5ba5458742ee4b8dae431a62c83320c46a2a6018da6
zab902e9948ab59e83fbe7aae8e92d463786861041dc60f899b30e7e8e9f3fed113f35e2b2651ca
z194da4b28baf2873329f3e9fb5a74ba02eca84e4090749e15c18de9312875b54cc67edab2629ac
z89e91b1dbf9297ca09812943b2733bf571b6a2ac4166e6b19cbb45643bd51a08c5f566d00acdcd
z89a1b7a088af1313cb19f3f135dd69f1683773e8629907753c548a115bcfa3798c7cba96961951
z9850905bb4e047e52bcff2b85f0afb02d5289d652aa8c86b1ad413228643087e3af16d749cae01
z7757eea015303536df8f41f770527094961d00ddd5665d211772f7c52c4e79d78a9eb29e64208d
za132cc3fd5105d171b583794b9bb4deaea302ac055ba3e9b7000759edafb2cb45d0f35862a4d74
z1b0b59718b0417fed518ba5f9e5a8142e90f994a39ee9a7cae15dba045918b9ef98db0fa0444da
z2cb723ebe361003d00b641939372d090a0c561a166fd6f41210bdd3a4251bd63fada70a672c323
zaf02674330895a58bfdbb9de8f7281309583326a6a993dbd957601e63e1a9e181751703f46aeae
zfd9eb10705db1dd36ff6626c68071ee68b488ae538d9a2f68dfd6448f9f58a0c9a9ac0c9615243
z017a3ab8c9440e9fa56294cb5ff16161f8de9abb635985baff5befbafb1071c0f3a4124be04e49
zf784c7b97034d4836212afb3b1ade77477bc751d7d8ae9bf375dd023798ea152ba93e3f71ff9fb
za05d85aaf6a57d351a12aa272d2007e92159be26dde656af6df921573e0954fefcc94e5f104048
z9e126af0cc47c42b5020b7830d5073c1e14a6cd96ca50d250c63f1dc2ee4378c2a218af9504fad
z8dc261f6679916528f96693ec2045a5482c85f28c2e06beacd6de1310642087850349b1908682c
zedae810e8f028dbb206b0f37c1320c23bcf23e0a157c11a5a410fb94a1e5ee54bbb35ab424849d
zc960d6e3c4e1352d6497da35c0d64bffc484de568087b023a46001a952c99f62e01b4b060a64c2
za5c9a5f58c7ef3584b27ea9118bfdeb3f0c072f8e09bb0d92da0cb154788fcbf979245a66f4aa7
z224274c9b7a332a11f5f1c2b3174ca3f9924f7fe3255c2c4dd0c9a7b936f85b6a26369f8fbea54
zc8e3fae3a6f91c931db1a5f5ad676141f6c6fbfb33dfe86683717cd3308f415819c9b221c65df6
za07d4d6e907a2bf6062b255254fb0f61b8ef67309b02eb0854b9d9906580b6e5324357c49eb146
z8887b1ed5a27c95114e89628e87a96b89c0ac06d60930f966113931dd352c448768cada98fa9f2
z9294d8077236f9c4ed00f843f544984dd28ae4d6abf24f5ce1d7a68a662373f9bab9461a8040b5
zb057008e1932d64e511901f4e3bd9426260f084ca30557a183b369b006a7d38ff64063c34c9f1a
zcc55b4ff60c508d9139dd35624339b4c72cf2f1aeda33c55e3496c732e7d2be4d10fc1177c840d
z45579af497aef2ba678992ba7c99182eea36f68d3302ac350bd06df1871d49b9a62560f644dcf1
z9fc9ddbe4422dde678300507cc66dafc01668d3387ecf74e0ad0eb06e9a49080133cf4cbaf4e6b
zdcd48e3c79bfb5d211b1508702121cbadfe775dbea38e88bfbb7d5c6765d026e69f82314c41120
zec9b0cd665ce5d7d8c982feebd37c95ad54bf3d75877c4613ad1f92ae6b0b38f83306dd772ff8d
z8c02ebd67077fd7325e2e780c7d76d6c98f2a3d9f803ab0aa4c3b68a5d629ac98c5c3dfe7cb610
z5fe7a68f955717e507ed4ae1083fe1e75e13acf46a1ce934c619dc287705da13d5c89117b11b66
z4a83ae46c41518fafe6997e5cbd85c80902ea10cf351974c3ddfa2c52c169c2bf3b9e1e02b73c0
zb5bb235997e4421b36fdd32823cd3c4381e59d97ba0c7029b1e2d7873c32e212203dc35f35951f
zfaf06bb41df09dd9a527e2ff3508fcc9ed67de700dee0eca87f6d569d96b7c5aeec9e47af73377
z055581f921b6848b844bc79af36cd3120d94c16fd91f3b88377d44031c15cffac7e6b9962df0df
z554440533160caf0a45307b6309a04ba521fab2d560441376c5c3bca4ddd394f37592840d29b4e
z5e63c410b84955cfd44c7c0d0c20ef9e8d0394355c20069ced69e008aaf50ec5322772ecf06a07
z7415f5f5370f2c346b900fd0b5e5dfba055d348aa639b662b2f64ecbcd955a9f7e643d1e407472
z741d84e3ef4d315e8be9986b0d37a8f8206ce851fcec2b562af4fa4cf9262b5f8d6e641f0f2eff
za4c6136a746ecc245b9ff2d94c60f7ee574de7aaddfc7e6443511870ea4cbf63bb805056a54ad5
z5dd3a65881076639d1ecc744879b239890f67cdacf18e2577e79abe0426ef4db77e1183ba76e3c
z7942f1c0bfab3ae2d1943b6bef8320b4170b9df17cd68e62c53ce6c4050ca5d370db182ffc1321
zdde1e5210a106aacf4cb833e795d449c788a89a0be546d0d905512a62ff1e33bed2d5f4ffa0551
zf4152422c4f9a200cda3488c7f1632ae2eb5681d68f5ea22fb12927b292b996567502ece48475c
z4a81e0ed95254fc90631de57af133e855dc1d71d09b33b6291fe1e8b8fd9f04545de9f00cab98e
zc6e86cc0edcfaca6a0d074dc5faa834741d4b52cc38ee85fceffae687d722a8a5c03af13e6e7fd
z0e3e707e94e63f6a02a9bc3d8ec445cd8f8c9adfe01e83fc67bd39b6e5610468212bf39eb8eb75
zf1c95184a666f5d33214f34b953eec760baa35b669e911e85c2c019dd6346eed6b60b401d6d320
zc17d7f0116348cf9853aaf49c3093112058b794849bf172c44005b045184755a18a715473c3c85
zd5fb34e0cb0efa610db0d729b9ecdceca2a517098fbee82301a55042e70c3327986a171e99e02e
z2843311692f743d7ec092e5103b2a44907bd76223833ece6a009b3e8e89ebe395955bccc3dd1ac
zcb5590e86006b612882d453d82d10b73feaf52288bd04e48ed3577dc8434b1933415faf219cf15
z52dc34652bf6d2186b484e8cde7288f39e6c573df02f8f6b6b68360d987216209bd3fed7db1636
z9c0f3a39656594094ea12bf8b4f8f9c1157e08cd3afae3d8387f7d0aab27e5ce88c90157cc3cbb
z633d46e4c9c2a55371f1eb09bd3524b4e339e8fc198bd9f0b3a6c6b889b8acd451bc857bc2355d
zd98c7c54255f344ef69440decc94e90577cecc994c6eacdbdc251606f728e46124f43c5b289728
za0646fc42e06d346e488b02c7ad0fd4696bd8148baaee6b73cd80905b8402b108f4e5e51f70762
z298e2e0d391c4664a7c073dce65f686de3496abe1ab807c741a39c8f22b62f56c0c56426a439bf
z922fd2a6ad91db5150ebfcfe615ca72fbddb850d78a3e5d091f8288f26159983614406adf0df01
zf0117d0614c4a2cd25c17ee4655873a70138a1e16081d31c9943fab804e8b33f97cbd16f65c763
z3712512209310820677f9a4569b3e56fe6a24f3919c19c9a4de53b338297c3bf0069ff216fdb21
z1e6e5b8cc6d282d1792a3760cee31ca5852de1044f4aa800c40ce94a6691a300eca36396f817b9
zde96a18cd9ba54870b87233b3013e214dc09d274fe4a7da46596d87dfe032be7f8d6e895797e67
z316ea991d7fb0181b4ed5512a7f9bdb1a387f186ce81e8121fb4b8787ee1711d73bb13a6dda502
zf1173fd735d9409d7849f3f1fcfdc092fb67c79b37215eb66f2516e689cb47a01172c080d649cf
zc5de71f74e9f2d03b17b03252eb56c502df566f26b73d8d3b19330be6bf0ec49762575c5409e99
z0d6e33e07774623472bab3a212b2bb6010cad507332222853528534cbbf15d9ede9594bd8f3647
z9e491420449ac34fec571cbaa64e9296dace842b88ce9131740bd047d3693ed50a11da2b026263
zc9ed230ab6df409b34ca762fc76fc1302c98b04f5a2d28cb25a3887450472a07fb0fa8b632f1a0
z68c1dd07aae66c568ff4100651389ac42041b3c2e333eb2829e2e5997b28bd3db3c753712770fb
z12ab94eebb2291e0d6dddbdb6ad537baaecd7683c9e6ce1068d14828b7c20cf63fd1fe87bc9670
z2697347bd6586a7aae47b81c25f90fb5dc06ae034823b8e259616a18aacd61a1542cdfca048fde
zcb19b12d97ce9a17b2f25af3f9c319fb7d002196d055ff58e9b396884b5d1627d4d222a781f41a
z2af6177eef1668c4ce96ec04ab5b34af592da05091fa12f19e6cacae687a969c887f370891d1f0
z3c37511ebaa3bed39f96e62282ce85292386f7ce7eb0b17f6cd65d39c8a11ed42dbf6c58b09450
z534ab79532b01453f8a6784cc0b74d6f9374db5ea3385753ba38f7d55b03a3799147405dfa84bb
zbb71766b717bf46700bebe5f1308cbd8595d0d33ad9804d08d46622ac1f9ce3de91e45f8a69af6
zfd3cfd514941b31a3a201cc92d351bfc9067f3098f308b5dbc2af64ecb034c35b79725c3fdb05b
z3f2dd3cb9cc71d421a5f4af619939e3a9f8b0e03558e0fc44e3a758368f0d01e0a46fb88d6ce3e
z0b0aac3cd48200d76471ca63ee0a9b7e713dd38382204bdce5c2effbafc59b2ce5cb0b4de56f9b
z2ebb6222e48ad5ad52e3407be8a2c008dfd40c6438c16839b460c0ef14b8aa43fede123f4ca284
z641056ab13c010f87f70619c8f4d1587540b5666373f9681db277547d6cbef1b2de4fa7ec9c405
z84a6a49ccc3fbe54caabfdb02231eb61a9984d925b66a5c3adfde3628c951e80fa90482c263576
z839b7c2cd02c64f2cefb94f86b867a62625acff22cab413a93e60226872ef0f36af55e45e158ba
z9ada2d8306e74d0919e544bd850009de533d7c2122efb5815b81940e0daab6565b27886228335c
ze98e479584008495c389954fa4389eecc9793682313212fbc17015acfa5ce4229d986983cad151
za1d017725561428f754b3b187808dc172e8a18f3398c2076a973e5fbc800d36029416ef03178d5
z587a006fbea292c7857a9efddf0f5d3a44f316b66925f5352b788e95ef2e3d149cbc356763c201
zcdb65bda2367e079ab67edb6496f9fbb72f58a0ce41437fdc5512afd2639c1dfc0f6fe52c375a6
z6110152b6a454fc35d45869380ed38ed3fe036748c4d22a34be049d4c35850d3bb7345c3860b41
zb02689a67ebf81db6afbb4f19bb9dc44d8a948d3aa1eca900035cc50368a3bbd4e712325337a3d
z7bfe0348ed48269180e7ff23e21705484da96981e6314023054b6ee9b28725da921beaa01d58bf
z1b45d0b8f6e4cf08c73e09bbe76b9ae4bb0e012c17c8fbdbf0a37c14cce5caaab5e032796f3a8c
zb6d7930edc936656aa182a904db915b523eb1946e5867ef775f532673220d442460f22c0f6e300
z9f64e5ade495224438aae5f7a2578a04f27d30155cd0362385e6a0fb4fe6f65fffc94217af6218
zcb55ecccfa3bcca3e176924a3ab41d2feab5c6c86d925255762f9435e767a105f8594f8dc46151
zc5b816bc9e7789e5bcca9694fe3456cb204100e0d8d74393f5a50618f8bfb067ed0d98628ac0b3
zf8dce229f813de1125ab4f4c0c7d5c016791dc6681fbee7bd1e221026817dc949ad92bf249630f
z11178ce825cd4f61a677bd088595fc8a5845f50b50b996d563e1d58d3b21e576c3e9d8de28ef1b
zb958378090af09507cfa0cbb10b7a6dd782ddd65d37f616271fac6e659c1919cf2a96c70d775e4
zfc737694a1ade222b60b06d3e66af725a0a57f41b9b9b29650023bac490d0b4721f7a8bfe2aa53
zede2d631e55633d144dff1b2dd6541cb627a7b873855b3ab1797f51735c2877a82496542cafafa
z1b47c8fd7f7079cc5f95b4b6e2a796b9e409a55438333f654f6e6d6e00782ceb31217921611f06
z103eb76b9645a60d06d213ea520390e5ccf2def9756a1d4384e638b2dc501ec50e1276741e8d22
z244f2012b6522315d884bed1209e5573accdde805e13ddf484b5e5ad790a6d2941e24207cfcf94
z0e9a52baee896c635d1be94dc95442bece5d65da0e69b8d4db697a479fa7cefed5b6a36fcc45c2
zbd3f41fc06f9deb726cc37e4b9c3145f2460d24ed515b42fda8239108812e3a59458fe50a56aac
ze6ff7e4b8a2b051bbff5e9d15781e899d095c5c6fdadb01dcb1d38ef2e24d4329e8e09b6160d06
zaad94b58d6c21118ab0197a49c8772a7763ef83b085db1b3e028d13e8f29b9887826ebbe16f109
z401fa82aac69269ecfd08088810f3b0e68532e09fa7d89730fac299e4456c43ac54dfc519fca45
z3d7e8f7abe9049d9ef7483df3ab006e38da2d60298644516df8d3a15b3aca740703c4a51177570
z26967625bf6f389cd328ebe1c715b3aaf31521b939637c294d1b52d3b6072c20bbb5a9c0c0652f
z4d3d1af05efc1f49c3ea86e48cd96bcac01dde23a613811f84059becc7ed5d490d4e7f0a2dfc2f
zb9019721d7395d408af5c1618f6461458354a0a88dec257f8355cc3e2a3ad0f01e02ea82e8e8cb
zd5d173f6416aab694863bfa701a543a1c7ee7a14da5b701adcf8ab35db5a4d437906295bc655e8
z2bbce527163104334f94de62381dc5ddc838ac0910464c6fcfdc20bbf29e7a4818188beafec0dd
z86fe050f86cb2e291124c693308e44cc8587f7ae0070e71282c2d11fa11e645cfc41c8ccb4924d
z2b509558498a0f8d961aa74901298bab5e8d18cb7d6c4d28f6ba5712d6c8ba573c3890de67b5c6
z9ea3d1acec4258005832f0143ef4ab4e20715816eed301b8769ade166f6ac8d6845f71bfa366f2
z1ecd5ccacbd9240129c9cb7b76a576869b4ca1e3d1ea026da117baef7f375a54f6f24bcae9966e
z31a732398a4099a4ab0f4189af48728e6b91fbcd2f0c7d60c70015d16c657fc4a8106d75e41699
z62bee0e3ed80fc6265ee6c8aa379b4360405322699f069c7f418e03e6dcc0adde226ac95bc7fc5
zdc66bfbeb23c0ac4a6faa74c855b27cd10304697197a626ec8defcfa47b4cd2860eb7213f6c90b
zeb3cda0ef458dc7d4899cc6b9938e62eb493fb2fbb0da909656d6de82dea7d9b1164a9ba85813b
z1a3c428e836f4af829e58952e5337e2060469449642c397a852eb4da46ca074ec7ed7ab2440f84
z2e7783f33f4bbbe274a128902033a47d9cce95a7c2105a91c1077caca87db6a80f97725d0b0870
z2981a0a105d0283e2313ec59e4bffdf84acf4ff703a7fbbea32c0ae0d727f303ab76fce07804ba
zd68c47e393a6ac7cf978bc713f794e24d3e9ed1a14685b396cdf7bd45034e79334f3703bcf25c9
zbf8e557539b76d7635adc0ecaa4a9d48c8121cc824c35014d7d5482f47b2b3c73901ddfec59e05
z6829a3eea27ee0e5942dfcca31ffea1a8d30dcaff96505910d5ed37a883e6c6581a258d7632b44
z085fe180fcc829527fc1d931ee6c727fe48b023f0c55bae94691ebb9402f37e1c3d719579bb584
z31e534c000c32b08f77ffdee6d9b23ecdf8f0dff4f059107e7c2600289ff36c0c458f77cda1646
zc7ae90aa57df3630e3611af4ff96df4fbb3d3547e883c4e58e2492dc47e69b34aa9e8eb1da71ac
z6ebedefb55bd91e622ea76bf13d9994d48297b3d7bec3d5e8fc15c6535ea016743aa536ef84f8c
ze736482d14afefe50199d8c9a3a2e5f66c6eee00663c478f98663bd5c6e89963b83e56373eaf6f
z6261249fdec4517f6eda597234aea32745aff66e8d7c5e1bda033929600419996b3b9ecfef3cc4
z5944fe9b800046185efdbbc00ce57a72c9337859f8fa688e162943e249eda143863913c34e1c85
z4f91c66ffca93f28d3c648dc4ffad33f924d5a1eb0982112e7d758b707add635aaca6b8500a3be
z694785dd003bf7cb4d4eb75c60a6f66ea54f41eaebffb07699918004c8b68772f36133dd8f0c55
ze44f25c177eff332dc6717f24315b72e2f5ab0e3090f728772c361b80c56d60eabbd1fd1a5b640
z89b22ac526868517cef61d18210c43863963bca0dcdeb32d1668b467deb28ed2190e62e44d890e
z836e3b9386aca7640443e88d86050e0d5fb5314d8bd4b3cf977c9e2ee298e3607329669e61965d
z6708b98570e55bf6daf50d972ba2f09b4e05bd064550f0227c4dab49c861a01fe569efbe1f8fe2
zb776b9c3dc2d97845c6d053e1a89878ac0f3f1379f04c87bbcfa5470207f1cbb29519aecfaf29d
zb3210f76756f15078dc810d98e5b8b936203e006b115ba8824f6892d0e272883b83f5a36aaa836
z2dc59aeb80a24cb2813633714de7a4f8507f86735cf5744d0db9beb364f4c90ceb83b4b28013aa
z7e7d034c57a0fa7689ff44e585d3fc4a357ab581b501528355c911979a1d88522d7ceb35a02ff7
z52fd4119e7acaa60ebd154273b5c23626e2f81bc76ae27b2fc779771ab01c108fdd12e3203bf21
zed114cc402b341edf93c59a77691320a0b0a68d807cb1a816af90813ba22b1d0c295fb08bd30ee
z695483f070a11a5207e776f4401abbe38bb3782205257ecd7a6732cdfb4ed0f3735e88cfc67419
z53089ee53571521426f1062a8a5c8359c128037d57e61f61c5d4cc27dc017bfafdd07a8cceee8a
z4e9eaedf76d74cd384a8ee4709056cb4c8163d93577daf2f1e018ad22cedda103dd6c939541356
z0105a0ed9b37db68f1e24b5686c9e6f32e149f674bc2feb4d8c064329c25b7cadf0823da1cfbc9
ze2f9d48eb9a41e45d7b5cf0ebacf840e30714ab9111b8a0ec01dedd95f51a14f89be1a7c15bf1f
z780b53e53df2e8ccb0625013bb6c0d2940cb7056eff210ef34f79a68a4772e2b27fcc24e3f4fd3
z1e183329baee05db91e3dc5c5a3863fa4c5b964c59f7ca5f41ac1d226ed0ef6abf0c20db90319e
z052924c838afbdb151609310c8093c11f470fcf20a4c8f95d10929ce32769b1f7ed7ff3a06dc32
zd78790e2d115ae457cb136104f21971cbfcbdb491ceab8bfbb9fc400264781b10b671513680a9b
z96d26129c7631985a169f51eb68b76d333c75161ee41b9bd37332ab5866b77d145147ef9e99bb8
ze358fd9e4ff86b06f2b740b3f53248f1b4876b4e8c91fa968d879b64bbd9043507cd808a919511
z987bee782b3236c4d30f171a5521b93d93830d7b3b9d407c7cf6a50711a6529222afb66aa43b11
z91496a8fdb5510028f9136d2d749a17fe24285363ff4b324e03effd30c3c163d0ca174bd362c3d
zcaecce9091983ae5211bdc28e21b3fa1ae3daf8647539bf645458dbaab26dffddb9e9ecb08c438
z78b63f1851947597df35d6628ec30abdd7ba54c0755979163a8d92480f06b74b2bb0bbd720a27b
zad148167c898b5975ba91451109ca56af9809733f92899458160638de54fae4108167662d83ceb
z91b227b827dd935586c6769ca50da9b172b6a87fede589e672cdd048bdcd3e9d1cafaead23aeb7
z794a08af16b6741631ff7bea031b74c300c2c68bab0e38cd23f475948e2cd9aab1a2cc058b7431
z3d3321e701c2c5821c78ec200a17a2c0a69beb1701ad41068dfe7268e480a3b2a6acc8af72bc55
z764a8824d14dd33adb50130b522a2b3be6490eb164a2bb8d63a7c6f967e7919cedc69634ce6bc0
zf802bab38fdbdc91f8564d7a087422b5b31af8c7a2d378ca06943ef559ca3cd6c466d1fb4d3537
zf67adb7336df7778dc98b97fd12ba19c52dae1c902ea436950c773b0edc28907e69a6273033958
z2c0c7be537cbcc55d09d81d9d6f7ed48e07fcb6b6de91c50035fbb7ce3433efddb05da9a35e924
z43d0c79c9371556a6a9e958c0c6cdc2a9b15b5f47322d405f483f7a3763cb90d9174c3013350c8
z96f72ce4936801ca567e771bb4cf72ce74d1754bdddbbe6e0e61ee4808003e33d4a25a3964e859
zab04813c4b82075fc90ed2597b43b9d6809adf8191052c85c0dfaadc070f22746242549b6f5dbe
z0e75afc0ad08e2436849d9b3b51bb0485b5275bef8ac2d0a9d9162761cad92767a62c8b2770965
z39bffa1e7ed81835e0644f4e0d27d387ebcd26427ae395c73954544d4670a5eeb7f032816862df
zec61a162b6898273fc3f0a17d65da850c29d31b81e3cb446507c2f97f93f9240e1d435992f864e
z01b2f9335ffc6f325b84f74c4dd9b6d99c9aa8c30c7739c0a5874060facffd67fd5e1f38db95bd
z4e6b14c5ab7540b4c8aa288659ffbee7deb9fd92c695bf325251abb93fbe6e1270af69cbf2814f
zc37004211c2ef50591dd70f7d8294f477f3e5cee9059eae3764f0f612762cd8ab540be44df540b
z1c8ff45124b50f8a8f1b273dab042941b4eab72f4d94550fa6f93348d7df1231c1103885881699
zfc78947cc766aef6b19974cdd100aff05dbb7e7c03b1a0f187f7fb18e77cc4d7ba4b3e01905fd3
zbc61e27e03d2a94279017a1e60de1a221603cb2586d4dd488f202767776711cbc0436b016f46e7
zc7bcedec0780f10e798288c179fbf6c11b68c145fb96b843c3e67e80cfcd196ea6fc290c93c945
z004aa8c3284863275ac47a83031f8009bdb515d8656eedcad76e6a491c9694f96235b4ffa622ea
z20872e792e69798bc4d9767604a34a1846a0482cbf260ff8a55335139c07ece34fb78d705ab31b
z3e67901c4d104f135f568334c153f6b18646a501cecaa595d62866f116fffb512d3ab5877570ff
zc0c1e6d1d544d9d2a968633faf1773ccd95ba6bf492899fab853ab3e364a82bbbd30a09567e8a1
zb6644edcf1211d8f9240c29b03461e2d8e47ef39386875fbb8a37ec877ee55addaadbbed62c5ed
z3ae6f39e63420c0666f15beca4f79894dafcfc75247782c0f656ed834187dbb73edf87162d51a1
z0397f66e8ee8b436aa92641c6e95180673c0f04f96f645c6e64194101980c623b03675ac7a20c4
z9391a9e5f9b850cc2bbcedb9cdf69bddd0ddc525f16e1dc3830ce8be6336eb5febebe36a7a755b
z83878dacb0688236f2a5f3d06633723a52ca9a71354c64a4ec6a982fcd9aad61c3e2587ac5bca1
z567d5971a3eddcb28a710ca2ad5bbf973d2ed075624796b26a6a1d6cc0aa1d96028a4bcbfbdd1b
zfae15fe581a0dc3cafe2ae4afcb424511a11112ea26901cb7547ec350e453a4349c1a0754f7292
z2399ad4f196f110a282a45bbc3366d934db052d7e8a1a8b167d68ad7080d83c90e4880c9369c4e
z9e8fa09a3022401a73639b03731e1923578c062928e699b98ef5d44a47ab371c1b74f2ffb7887a
zcfa9c05cd158fb48c8a3d29c9bbc9cae89dafbd3c07ee3a71094c3184739a52267fda5aa847677
zf0ce2ba0e64fd9277fa2d8774056abeb51e7b3a6214a8d27f2a6f547bbcaa7d493fbb951623c85
z17fe86687de9dc4ed91fcfa484c740022bcb969ee2b538dd20e62f8e26b8ff52336a309c60542d
z56eada0a37cf19b5783e1fedd63fc9b78e34c7acf72519d5a9d70b9d41af0bbc54fa420b4902bf
z32286fc103cbe4cda2c5e03c403cad040f8afd3b37d6e4313994dcacf832a6ae73a9a73cc6aa00
z170bbfcf0bbe7ac7bc57ab69deaad2b6cbb5535a926dc7da437c382e3ef21b572596a597bccf8b
z8276165ccd9f398612bd30e946dfd978883152e83457af7216734d62ed9a2f90e887d236469879
z7ee02f8977c56fcf02434f64323b8ca48ce87f98cbdcec5623c3f60f5979dc7aef9d2a17e26174
z2695f4d2ae47596a8f0b184fe938ae012114779b64362ce78703e3083517eed3c3a2caf44e0308
z26d429d2eae638d633473e3888c9c01fa7320a3546ecbad9748a5429fff45d5b85eaf07b23f15d
zf8e4d53054546c0406d0a4d9521c811ba111728239d44abb6f1603f6d9034751a5d0c87bbbdbe6
z844b60e474335403c5f20128368f54f0ed548efcdff11178d2a07589b96b8f1595e35cd2cb64b1
z25303c5adc980992294482b453a3970bad37b4a8bfd4f3ebbb3b7d561002715baa75175dfa069b
zd1e8621554311f6ab6f19c7760c8fc15cc1e9d4dc643ccac039ef7dea8a65cb1e02200017bca17
z21263b64777a22dee727366c29befd4abe2bc4a63a36f91365b02c4629dd983632168188ce3e08
zd02daaa350bbe1b82c0869b63461429894fd28bdec4a2be3043eb85237f4a5009e14eef9bcf759
zc1a2bb1490b40d09937d2ca8a787ea82c546621d12ffe656d9bef7b73a3aebf0d174411f12cc4b
z950fc32560a7145adca24046f9c8c2a4368028ba1fe867ea16a0eaf7c49730c6cae93a7058b4ef
zee83983ca65a16a35c3f314d3efe004a76068d3f8079330274853afde96ae3de0c0cac9a8df458
z75b5fce19f33af5cf62320e7b7154703f158e7d8c1986d8f37d3117c549a625d7f525e13d26680
z5725b5e2e2fc2847ee22e27a8b8e445f8b40852f2f9f03dcf3f60c298889e2a8472b64815c0216
z3f4c843444a28cbad5ab87448f7e74cfac260290f460130403fe552d8d9ce95da6db9b9438bdad
zba07aa29d10d05247c148091d86b582210b7caf78d1205daf8e5b344eeb32eab85875ca1dbf9d3
z24b3c472e6c197e1c3ef9fabbccc2f42e16d83f633e240b3fc05361ebb079b77124aa5d433c2b8
zc2e2615739cf6efee86d8a7b93a63a18d0283cdebbdf01163d7b30fd31e909bbf5fd7e495cc91b
z960c6c7f3d2cdf0be8d25182d4f1a4e5b06f33ad9882928eca252646a17bc027f957fcf958579e
zc1d39c3333a546e059d87fc46497fb161a9b2233cebbfc84615f6a7297f852c3b6058aef37034c
zcc6b577530dec2ea39c4db48fb2a437005987e5d85f45a0707932b7a2f208a14b2a6cc472baad5
z8fef4f7e14fa076e94943ef6fcebc1cd1192caef5af659fe24bb90c03175d4e398eca08efc8c3a
zdcf0a5bf2661114e80181e9b4cf5c3af80bcf13ffb5da4945ce4c24be781af877f66d59966e1b5
z29f5b6565ca03559a2387f73d1475f71e9cf86df3e7f3685100af9efae55385dea8244575916e1
zc317cecbcc188cc6139bfd90024911c0e5e5118412ab402f8f2eaf64df236a32415399d48b3887
z9e27f184efc971dc199de4bc06052b6c9c5931c72882be0b03b74b023416baa51ff6d46af408f8
z9a7a3271504926435084eab2e497e2ff3c0a60d65a9a0c83150c652ed1e90642d9663c3e32ba02
z9d12c6b794a3f00e6d4f78f762144923615c6484a66dcc1fe6a91837006e18c23da6c42532d6fa
zb674dc853690655d6b41fb10270e748eeff68c26d7326bc21a609182f34a101dd3f4d6ed01a945
z5ce099ea172ddd270d504b7730b11ab50d063779f3c6e217cda7bf8e690b06a20a1646c18ef72c
zeba718ce00b1fd46fda180ef796f5944acc862e142f6104e2b06b0c1d01ccfd2cd8028fb7a6f12
zfbb8506e8e60df5190834062cf2708794cd451a54e85f61bb1df610672f59d66c5263a1513c605
zab5edb145bdd68b50aeb6634a7041746fe51934e2773ee3641f1850f4924f0bc1f8d3efb766604
z1d4302adcffdfe90e35ccaedba80c4dcba8e095e0a3370c879da4f3f684ef84db2edad34488c83
zd1e3bdab5b9a3d382841ff9974de77bdd707f77dc36d8accc4ad28846676b5cb78705846976f2c
z0e09b5119897ef384ff8e223856f9e10e3e3f57b37ce3ea26bb7c71e18d80b429ba3e56775c425
zd68a7d48e1b461b5e6c79500e4487560cc7dccdb477fd81054b6e96416afd5c95f204a62e497ae
z3b42d20f70055c007a9ceb92664e51dfddd1a9de93bf886513526b37a662a5e127ecf2c18607d5
z8a7ffdf5a9fdc69f192ce979d447dc5fd3714dbafae7301f78f61eca9982b20bfc5cdccef7a3ad
z897bfc14d3fb9db160e890b2669c67e8e40fe6157a9e1a722d87b7336ce9447928e480c1f26620
zb115f57acb93c48059b4f8da1ca2aee3677d14cfb4ccd8c60fa46c0545616687777cdddbdd1e6d
z04c325966ab30b35ab845e786b2e830f09793b23d40bb381f5ac61eb9fed886389f1eee5d970e1
z911685282545d5fa89adb6ce1d8d3235a4c6f696f08eeb1e9746909d22989cbb15549441a64633
zf05be5f0eaac4f5ccdf4d699326c1cf8b6f8460c9cb7ad415f002de6993584a391ccbf7d81c3c3
z1dc445a0d84cf50b6c54304af2feb2af85385187f2bb579271cfb62ff7b3bd50d3b2c48276c983
z189a11c79c7b2cedb480d70be8d592fad727d43640fa6ca2e7f420b506041f400fd4f7176116ac
zbdca440cc047c3cdd7386bf57a1833fb2ad02b20dae6c3b6c14edd025ed69b174625291298cb9b
z10aa1063c1b6e4bddaabec69eda3406cba08ee1b460179cb28583df2b64353c90dd29342b28f72
z0cf5b8a31a1637a4502c8b0e418c4472c40dc3badc23dd7df10ef130eeef40582caac3963f46e1
z887d836504739b1e3a58965133541e8163e85adac8ece6084c7907d804b16c3a569a657643673d
ze04598f7760dc1252fe04647ed5c838da85d53170f0d7dd307e60aa94fa7707ed906cc2b5af234
z22e5b49688b9354d8bd082511a60bcb04bc36c12580334f99ec835f64a046b3bb767d5bed651f5
z493c7ad2ba035418644d67a497173658227feba6ab1da327568994897b2bb8fd2af5c6f6a60bdf
zcf39ce18a3a39b3b88618575d6cb926085d8e71020e7788cb9ef4df78c09c6483997be7301fbed
z883e9bfd5f065ccdf7b46ff7649c5af3a31c6daeb94c0b9bbbaa74854bd13380a04b0e8266ff9e
zcf9e16a044adef12c32a0ca58419e1da31caa1205804f5ec55352fa215c5c1fb37d78e830ce728
zf180aad566d575489d42cdf2eed9ede2d2e585df12013826f6e9ec70cdedcdf67ca61e1d896e70
zc49dfb0ec07b8e375131f0849ad3ac9270d260d55b8fd04999a708640b0781625e38ebb4deb824
z303728636924926023d3e3a6281fc00c545abd051d7685f1bdeb89ed3a1b0bd58042aca7a5f193
z92e2160c157256ce660239e2907159393d3261246e2cc39edde2336e0d019db70c9f6cc460647a
z15a44103465d260bfbc7a14bbe24c18d1fc6a085cf34620992451abafbac502bcc5434b407697b
za0610a035a261a104d35d405b61754388ecc772b337c4bfff04ff2b3260c17d597549ecf4950e9
z0a1093998850468db88df3447181e75b5f6ca3d39953d1a22c40177a94970cf19488c4332285bb
z26dcbffc9070732cf808f36859bb8df2f3f0fda5af15c3ccd19d76351523f9885ff53e726d2b1f
zd0e02cc800ab0a827f4431b991e94225e7d85101742377636276764985267d80f80d45c4b73a80
z5041e1b653f8daa5bf50185c8d1b1ad230bb4581c6fe92acd5feeee9ca365d0a4c5ad1215a673e
zf1556ba820e21a33751cc8215a5186849e42f40bbda5c1a05b2246556c7a9f610e53d9ca682c49
zccf3c3d114a75a943f8a650a868dbc402b8cb9282381cb43adb5963ce12773f5899c25f986667c
zbc98fa9e608de4a8a163bbef00ef3c319b03ed309c191f10ed194194b20b84beb4fb7e22690629
z37f5564e8b805c1384a78382a3b7c95c9cd99c2624c9f5344b84eac83cebd23cf8ccb10c961b2c
z7453f4d741b418fdf1c48452b3f9d148a8f88a64dbbd653af765b7b9efb184d4e6ce554836a0e0
z2565a4107d6b2a7d1e0892967126302e1c8b3157ddab2f4be2c01d6c99d0ac94405470518b7dd0
z40927f306bfc299f255d431abcf4d5110e4f79f09da265d5895fe81e73211bfb820f038f236054
zcdcf6348e0c0bc8e1a07e3e9205709791161549bd81dc1310b0cfe499d4dab8d3dc86bb9e6027a
z4883d465484471d0bab1b9513d2bfc0b9c826e47f84036d3140527aae9e50317cf77554b0e7ab1
ze2e11f6b155aa872441c750d780ad7a662f2ea0d4636482be14c2df7a6d37e12a9896cb2bf5688
z13bcb23ffeb5c7f44e8173d84d21a029d5ad0292e9362dc6f25e93ae06eaad116cab11c1c9f729
z37e021ed1dca7e7baf512146db1115a951c38205843bbde9cdf7b2074b5716bcca06c174418c6e
zcadba7fcedf34fef69544c81364a7d39d066ae785d9d541246913cb28e8c080a371ec5cc65d372
z494c2a2adc0790f0a2951833d42137e1250ebe6b1f323b132d310a37964030c4f99c130358ee53
z6057ac5d55b890c20e764be6faa1cad7195cd416d00982fa753b61fd2da32cd33eebe1c21a43e4
z96f37c0ce07c6e65c323fa385beaee34275cfe7ba1a7d2965f3ed66e2cacf42dbae0c78ea63910
zaac92294d92b745b266176589c485dd5526ca7ad132ec32c35f3c5e59fdaab519acb5d85f5c9c0
z41b37543526dffebf6ad6fc610ff65de5699416cca1940946afa8cbe4f7f050998e28aafb25a1c
z013fbd3aa3e5c11ff881a94c17037428820477d5274ca3c4317ce1fbe92ad71831ca61b336c938
zd3f79c554bed06a3e0927f3f3ab1be14ac60be7d473dcfcc18c65502aef6dd54f3633c16592ad1
zfda88f245edc7d650306d2e3553dfd80de5dc12a55b504d572cd61bb3f14489622474c404d0f8c
z2a419742255055836c731a6f60dca6db6284b206aac3d6978add44f38ddee5b2e87fd760b6cf4b
z517b79b771c6f13ec47f5c040a86e5a0a7787550d641f150d24c3669b9110337373775bb9f0f89
z9f0e248b0f008205080636e363e76ec8f7c8be08d89c6815f9bd188c10edba7008a216b8b83896
zea72a8cb697c1893870ccde5ef64e838474d666b3b9282091b4868c6f68a516f644d493a1e4b9e
z395edf6c1d17ef9241d22a68b1d0e3b5701e1ca5e4972a8bb494238c8b7a7b3f7c260b6e0d612c
zd719fe179644e0d39b494bb212e95838f610211fe277683ef3a53ca73fb5070ccd9ada8bc0af6e
z636675e724c97de7bc7fc77357f48168c758483216bd193042bf7eaec6cc34d04c49f456c2b126
z0ac1b243e3bbc92c41e23a129e32c94c0801b9059761ece135105e36bfc7056243e00f06e76d8e
z74a92d30b52512cf5123a1b9ac26f01c2eed5484eeefe643d9801ce900a1db770c78c4c5429b7c
zcdd2d831712ab5709954a9f7fe906ae925cca96007754470521b6509c1023f0226aff16a2861b3
zb25830ebd7c0f0a3cc1dbf4387519cc6e9f226c16a1464c907573e4777d013be65301e27ab51f6
z766512689911208dc45c5a553fe809bba72452e0a0ee3fe267c51a450c1c1930c1457ba7789af7
z865123764252a5cc7a0eb3909a8164890157c86c193f888bdc34da3fd8b3d369dcd13ee1fd8ce2
zed05253a00642c9139c447005de981894f12cc375dc83079387f030e10fdf7786c7669adad7bfe
z5f1edcec270165a0dc3818552d17abe54d205313cf537da3049bf4693a99a7f36d046db24af008
z3ba2267770fd5ce5f48e7b541d97581ac587ac33e8ead18e242f21da9021823232e36577bd14c0
z29d97932e9b02aa92cff631d7ed9796e0afd4655955cd75d5fd3b235f8734260f726583418042c
z6994d161588edad1b8cffe837a29019078d9374eed126d665e7d07720af6a2f0df89253f3d2d94
z459412d6a09ab32d171e9d5c5b83292a92413ffee3bc567a00052e40bebb6888333af4c076e4ed
z3c1309c0e9e76e6b83af8cd2e540dc3c17a3c5c7decdb18d43e6c0bbe384a6ee70dfafe8deeb99
zeb67da69eddb86b76b3d66ff17f5551a995b57840a977c1910303a42b46216b1d42dbc71b39788
z9bd1d54fb2438b9bbc14e2963c86bd038c91193466bb99b1325524caf8a64912fc40520dd7856a
z042cda19c0466d9410f66fc8d28d8dab274d2b27c4b5ca798c2db170adf8b3fe3872ca40afed58
z056db425c96b5e9489f847d5885e942784293e40ba82ba2d54d2fb7a13626239b55379b14e6142
zf5164150e41d37c88aec6d2f1b26e1a63903925fcccecfa37d72433fdcafdd8fe047a5b8a598b2
z1609a2528bdb9dfa92f9f968dcc782c847eb7be78f898e90cba02e1da8d0864ee1c12b1fd8259b
zd03a1e9cc926ffb2a987cd2849a48c239466ec6fb66bbb768feb8c63777d5c24480f40eb8ecf8b
z2fe3b8afd3693841b8f83965d4b94dcfc29eaf8b56e3c25f8ae52fec05ed413955411d8706b340
z65def1f022b41acf084bdc463cebdfffc139a1416a67b3c665160ad34551ee5ba10950977326e1
z6ee7d0b333f489f6323a3557c4bcd898da9e5c173ba5db3d7b3477c9bea290776b10884f0937d9
z69a1f3cc63ec10cebe1d08fc78856e04a140ac630f19702696cbb3890b27042ad03d8fa8a2eabf
z8b186fc8e6c3ddcf3dbdd48611d45471e14b1c130d8d8cfde95f6107dad21f2b918967011ea7d0
zf4399f16c948a79234e3cc0362c0b2697459cf773bea6cb364989e5b8b5f4cf20797626485b60f
z5e909daffc1ed423dccb36833dc51d447f1b9a83b2090271aa37578558eaea4ad3674a6c181983
z3f2298eb0259337e175df82598c6002c878cc6931c955ef9ffbc2fa22f37b4f13021afbdc4bd13
z1c73732bfb8b37c4fdfdf04f6a0a0505854d5bfc1731e63ae311aea2862d1f05c2b8598cbd39a7
za021ce954fa8f9b3259fc5733eaeba56b646150d2e4bf3816e01066d3b09e18ef16888953b8b63
z711767fdba4a39c2d834023b23cabbeee6f29c67145a341bbf90434b97efa784dce0e0d2eec267
zbabfae1b23392e185426433f09cd5df3b14cba016657be0e388080bc3dbf361a77ae4238525e3d
zf4cc211096d491c14e0f1b014039b8dba5c5351b1cdae1b3d3277b3b849e9bddc7b6e26f33daf8
z0064e86d295b4791de909dc6947c124e81ccd18a268cfc6740777131108d2ff0449ae37e9c8921
z00b644a5dca8ee34fb46a2aec799bf089d74395b9dce17800fb63640e0cf031e80e7f73a039fc8
z03b041a63714f7671f60bf7bacc810ca355768aa8eee36732dcb0969cfb38499459178e665c31d
z85d270772e5fe5d87706a8e709919927345df27eec880d02bfcbcd3a5754181707643469f67d14
z7475f23c086b8e2f19f934e500b5c6488a9dee289bd67bfb088345bbe7f02ae32ddb3326a4b9aa
z59cb70d58c70a83fbba58e9aa864399f3d21402becc4c687e2646f98ef7193192fabc60539d3f5
z2c0c2b597326d490940957b25a03014a641f0fb46f72bb02d1df533619150f8e44d9ab385c9aa3
zd654f5a37a6f50d02ab123b677155c172d93d25b89196e67581b04935a5f4a4ecf448e07db5234
z3a980c106c09ca4db27839865eab7874dd2aaa98242f27e0dbf023a87ae27be3e1dea5bedf97ca
z7a6d38f3ca44701cd959613289cbf09737bbdf4268870b5ed8c5cfe677f739e4bf50fcb7038937
z8925b44fd590011e35d2757134a6565f62206468e895add8ea582f81eb746ac77ccc28fed08cd0
zbad0ed6de1c4fa45830e278e0bb5780a0350ae3d2a4fa1c1c797ff1d42d5568396e9ad187fc1f5
z878c0a4c79ea5a3051fbfa39b9d63f892606895deca43a80d8c2e78c73ffb6c183c840d9a0b1c2
zbfc22cae9ac26fc85c6e24cf406780a37f2af6fddecbcff391090c995c3432e71bcaae1a45c0d1
za496ce425718a799d7570966973415651cec8e2f4a861987e0108c20cdf92aced01b863fba33d3
z371c27df065aaaf2acd5dd305cd3fff1ab413e7f1087faf8f746ed8c228554ccb6fd0edb38714b
z86f21d2239a867f556b715c1a9a6471134985e7ea32183fec9310fb19a9f6ae3a98dcf6b596af2
za0f0331c67b6fe895b3842b74beb53d627edc06d095949633ac21a53cc52d68da752e54f1fa265
z3f1fe7ad55c783548f2beb00fd54044ba221a0d284428e58d02bf1634ae95a17c8c9bfe6833d7e
zc8c00958e420b22e4cfe21d5c9e8dfe6d3de91bda15b30b636493aedbd7faba115e13d5f6909c1
z15599f3ff8636ce4760b47fe17c5c4b1beade4194919e839de21f489e770b36f9b20c1b27e5d48
ze34815990273191b4d342fd8a4712041449303783ff26f723fff372490bff4343f5ff324db881d
z34aa9f227a683b5ce84f3e4fe9e1d087fa71481d9911c9957057e95522831c77abbe8584b495b0
zcc1d616fe096f7d9bf9a6474cda036483ab90af15cb5f15c0b968b8217bb83c7be7b7ab7aea91d
z35b21ab3d3ba112f74827d28d80bd27b85396c15de18d5ab9aee6c4773c51fceac38ed5e2a7e68
z9a3061cdf9107aaa8134d3834bdb37945cb37e1c146a06cb1505e70bf2f30ee27b1522dcaf6138
z62b80e7bf965e172aae7ac960b989dbd9eb752b55b7e81c935f4a85f4bacd58effaae47d31d5e2
zc39c2c8ed0cbe1dc3acb07869eb125563f4183ab84b6b48b69924bfc331fb2953eb7f533749153
z65692bea7b455b60851e37003a242d2fb9c56ba09efb2b130d2dacdec3ab3e95976ffd75e24dd2
z38971a80875d35bcc5ae33107bd14275ffe218446f81f17b75699b940d852420969c6a8a9fa920
z65e96c4b27996aa9872b00bb687806e6f80a3e690bc0f448b18f5e76ca12c969545abdaf48a804
zbb885bb7d51eb10a05aff9fa94e693e6d24e5f6856e13c0033186d176a7963fbde85a0a8f72a61
z92a1414eaa2ad3ed093174eb8d8ebf15b035d550097620f045b2461e3bf1087ec885875aedd5d1
z839b8602be10e5aacb9536f8b91cfd1f9c94c0a427b4b43c6238f7284a8fb546b07f3e33ca609c
z2aed855b7ca2d415eca663758b189b4441be2c7fb0366ff828764f9e9390aeb9f598f461d2f832
zc209607b8a470a2ecb30117dc0db0f1ed27a2ddb7723ddd31ad2981f52d753cc27fa9836505e5c
z283c29ed6d03ea3a89074985bddb0c7e09f3f967b94521292b517e92a370ebc22705f0dea7a276
ze15d25cbbeaf543200a19bcd6c0a6d96873a6d80410a016ffa7010522f3a633befc5bfa99f25d2
zebfc4d0da664413a3b2c9aa392f8d957cb6b0169fab66c82e742b8c4f6a401f580f626bda755dc
zdffa8bb1764e45d09a2c846888b7be1ad8a176bb439ef7d50dd5ea550c5629b47d9905ed10cdc2
z6f684ea2f3225bda59af0218d0aff16efe82ea32987a35f513a114ec9429a42aea22fc5b7fc4b1
zc3bb9e702fe2befd0b51b51bd681f4f95e4e683ee74bcf508171b5026b609d53bb31c0bd5dbfc2
z55766817b566a54e35b87a0eda6c8eb294ee2f4cb90b956e9cbe6b241d54c76c37ed9e70506d3f
z218a42647ebd0ea68a6586f8e7ca7e5d1e61fa32a717b73ee5be6e2291c13cd13239870869c503
z40d877a035c42ffb042991a3442af9711e067c045254ad3870c9639db9433d9ad0d64b9b7e846d
zd91b2fb18f18765de3615fd280c891890de9f7f443b1cd8a512b18c07453062817f230a10ddf67
z7b2d323cc5b5222ead85d0701c2101275d4f0275f71b2ad1390e3d83ef40acefe6a872b25285eb
zfe30c2a9f5cedbfed0519ec6b3d153f65cba70c2dc9c94ff9e5d7628af992597f8dfac5cdb77ce
zd8055b9a80cd1aa22cfb49409bec497455ee150c55c4290ddba543fb9e25114a11c28090017634
z9b57522af0099c5adde74751504a65c82a57b795cc9bdf0a45cceeb5d560b5e22da307ed558088
zed6b7425badc11c45505d02ae0a099025de8e6da5354ff3dee44dc01374a3fbbcf11687b1a097a
z9c5e4fa20f9c13b443fe69bcf3230bc8766014c2bee0a87cc5d9ff0c287f9c7122ca9be76ae44f
z4e2ab6fa6d163ca501505baf39da96fea9d4944dc777c5df898bde4f7f299f6ddca7a9e5221a1d
zf599e7a6363737ca828e3716eae6c02c3f4fa7c3adc86129625ed57138fb4ea7386b48b8a2181c
z0fae8f00c241e212b5aa917045d9b571dc19217018eebb4604153aa56c48bd6e61dfd07c5248c9
z21c4c4061744650c4b28745bc8b539c6106d01eae8f06bf903a5b228cbc9d510120c1b75083653
z205115bdd0a25fd6109273e2f8a817bf32fb0c676cfccc9a9e6246a7407713412289a4acf09254
z146f3c0f10ecdfeca88b7d4b6cfd72ca4a2eb909185c076e574e9612560bf2134b9ffd14a743ed
z5ba9d491f0c1dab33a9f24e808fe5a6e60961497c1a9c717802b7182310ab68b24d6c12f7fc043
z695dbd7967144f70b7b2dfc3147de823be2766183a1497e747925a2b205c9106468eb17b45e0c4
z237cacbcdeca5cf4d530a05c4aa9760d56291011320273206f2c01feeb6e68b65717540afc39fb
z8cbcc9acfba49039457cd9008f0bcdab71ddd49570850aadf3b65a268dc2142359530c29e06806
z7862c4e362ac4e9994b11e9ae68005a144aae629a29000472b27c8e159322ce4d3a7f855a3a1a0
z8718c874dfa1770bb058f56c2d1a60647cf8dff64f96469e2b7ae3190b825367f0d1aa060c45e3
z1ffd7ea61f00002876d57345ff0e4b631084d90c7ce3d9f798dda47699005407ec3df948358367
ze853ddaba3993dff896a3c2865e4f318f97164da42dd355701ea764bc6786802854a1f4de5975e
z2f8389a7243bfd625b2ce219bdf69465cabdb2111fbeddfdf754666a2d25420831782f00a214c2
z1b62f56e14236a580613c4719e3a6216e0a0e4a87e5de5100cd837d76e6ac3eec0fa2fd41f4acd
z3d8e08e29c2d1732237a21e0953f24c6d3e30ffd1822e0127c2e3f965d3ce8af6046b36220f832
z4e53897e464027fed69975fb069b7441542b934e3f21ba45b5a47cf0ff81e668fa05dc8db575b7
zc1427bb29911f9e49fe0b647433c982068c874c1c68072dd8ab020f57223781faa682f9e75e8db
ze98ec7eb1086d17a8fda3f3c0410068715fc0c4a6bf6667b7d4f13c96252eaa255c2e9c7828043
z1504e8b01478240b3d73cadadbcf8d118cf412173b3b5255e16ef7bdefd88dc3e950250938f224
z426e693814b79d8c420c4b6f2fb0ac859accf2bd1d1db51343185263316f8770901b50ba4a04df
z0ecacfc295deb8ec2f526270160a79c066b8d358f95f4e49519953a700c4b24c6df2a43085fa4f
z69c321cdc3ff59fa4919ca10eb65e3e91d154160ccfe7d060dbcbd97425a46c71cb28f4222b53f
zc800c9bdca497b2f781e4c678919e9e7ed2a05266721a91bcf62fb9d7d9d6aa41d27e24324c0d1
zb1b37bda65bb3c3e8fc167e7c5ff78469635a4c10ec18d5273f91545253d13879be909c251f0c6
z5034887b305b8cbceeccb71f48070356535a3bfdb512c5cedff50eab9e614e958e538bbd84af79
z416dfa4641b6fe6a720274570552d75fdce701d720cb956787352f4840b13113b48a8e6cd68032
z888b912dd73f6f34a83801cadf534d2b6d3851df0c41aa9a7049ae22a49b21cfb224f50fc211ac
zea521c7ba9b134ae4d1b149712b6b550a730e9f3d5f75d32a1f8b7e80d60bc46a30051ae3dde73
za63bfbd5bf6a06e764a202846889c058e0d497dd2f1cd627a6cafc00c540dae9a6b57bfa099ef8
z5c0e27d22ee15fa88b3fb739a71334e3e15abffc47636751e9d2a94f6c188cd4c50f9e3d3326d7
zf163352684303b6d0fb429d23b95ef39d21c353da88e7c9db24dec1b3a4a5606dd91be7b3281f5
z30bec13be51e0c8a82c507ce1de94b9e3c8991e39a6686ebabae413f5e36e3032b5c49f1214d12
z7c10e15519f1ae8784571250219b27748703e4a7a8cccc3d9be7e7dc1ac1f2f8201e0e6f2a6caa
z3e1611766bafd92bc05eaefbe8a1df3cb302cd5f91413dc67bcdbb700621b8692ad99c6817877e
zea5315bd5ea49dcc95c429db718d9ea3e530fe71ed811ff1becd09b0ecd7e31165376ecef53d46
z4b8ea003fd2d7fc5546c13c2981610d2f658627f28d8bcd85e342fd3559f4e80dc8316505f67b0
z0d284353d1fa4316c2c17547b295b35a6b2f2124444bef1e4d7a6dddbdfd03eafd590641ea5998
z4f112edf3737e595eac4a1c29b89b9cd147075d14f6a35338e792849ba7a1f1f2858a50b8890d1
za1507bbc40a97aec890427d3c76a0410017d5ea39180f546e0d6242f016fe8d64a650e3565dea0
z871fade0defdeec5a517021a6a7876e251c06a6711090333a516965b83b20797c6cc2943741c18
zd59b841b364533fb4ba6a5c8b4e937c3b6a38fe75b530f99b15acbc959acfb5457edc0f25e90fc
z9cf2362daa058117e946be0968756c9251f152b849a18fba80b0541a11c4ef2d76672e431bddf3
za7419d32a5b5456679e4124c7374c74dc2bd3485f772ceb42dc2c89c7bdc32af86a52f0727074b
z0ec3f583237a102086c32603a47ffb718c9e1c268cea6251f960a9f9d1a6ff58379bc2726b5a8b
zf7257a9d5ab6c63c580442997af2d5febb5770bedd4fdd8a4f80c84b52798263891dd5f98cf461
zbeafc16784d19124085daa454924241501f798e45e4384ce83675868641ce81060bfa065fbe6df
zc53296fa66576a39f60a5730d2e077d0427c6678f31dadaf563d4a7822dd1fbab96360a1c530f8
zbadc756699b779e5e736f05ff780bfe1c340fd5152eea62496caa4253dc7bae2755314215f9268
z0d3cf0579b974c078fb825aabd63866c1a9f52de7c098a5ec75f2e103b1d0321bf0aab7b30d072
z227b0b86e38d36bcc6d637c914f246f43a45f541853b8876f204ed7825f4baac018af88c257dd1
ze675903bb687898b812d9f54c76e210fa80141f76a19f32545ee6c62120ce52d0e2e508920c435
zf5f9f39c7aef17418f2f6474d43a0a408414b1e33a4ba9f61795936dea44e005b9a786c52fdf67
z0513194fc93948ec2d4e469f70df9911855eaebf1927ba3770bea13f5a2d55aff03ac139c7dc09
z6decbec4befc6cb9a8245e9c4dbce9ae6b3d3702669e0e975f27776c71d87cb5412a307462dcc9
zf7cd574263fa230156f42aba314dcceac0e0c4d5c5977ef2138a536987bc118ccb41ea701044a8
z7da5e47b2d17ecd8a24a3bc0e2e2d27711b20f16a27787a67d4b5040f0559d7134d18db7951976
z6dc95978a866ad7805309156f32a2d60cb235f00fdcbc394f3fb3a420da29393ee0ef270788b14
zd0f4e639281ef0cbb286dcfe1e38ab3c80a69f9bfac53a79faaf83ae2b0fa1e83b4374f0a6d2e9
z9d182b5f03a300a95db01784e5a3818698687143cd5945301a5c450177a737e371608d01cbe3be
z3d13c268536f3e1ad4d90301b2c419dace017ebbb66d4ab374cede3cfc60a09af7d99749f41373
z12107a316a666e3086127000744e7667ddd5e2ac7f031e72da449ec574cfd3defbf4b7f9726b9b
zd3bbfeb4ea996b663e5cc4a4ad194bbd62925635f95f275e497d555e1300fa4ba72912968c7b51
z71871000b43e84f3c68969a0750098aaa098b11e3f3306e1dbdbe979cb157584622650360b69d4
z92551f728dec22c791f78629f929e115acfac472748b0c5f99c3593efb7e7a384c1165037572ef
zae694bdfd7b200494318dd09901abd750ed66c48d0761aa0cc1c7b444af1cdc2922713abf07213
z4fe46c877a9deecf5ae3f05a0e52259025753ad74fd79c2f4792e7b106a9294beb56108211a2eb
zb698ee120af40543f54a08f3935dcf6911e48fbf4aa2a49112deab43f0bc9487367d31394d3839
zc096c9302c4c3152e3e0a8ad5eed63f8b8c371527aa7f2e9db084915982030921b6b3dba880816
z4776e793177f730830bd8447b5ee8b1b4bf1f310f4bf5b639a6fe98ac5a64dbb77fcae1e26edfb
z4168460afb9cdbf26e401aa493e5805240090c2033d87e4af832b3e71424344ae0ac3f7884d14b
zeadf089d361578f47c494ca1a6c1ff1392d6c8b1874e5088eb91249b2cdd7a79acf701428976fc
zb58b5df4e8e2f59a0dda4cbda2943075532d18930b4183b41c71562b1c84f2001b30cfac566c35
z6ad5bec67319cf8b5c9e00b2c908d8b487fc20b49521c2b6636ae44a18dae90c67f3ec925b7ece
zf3ce59355a51ddc48eb5865691e399d165dda1ab2d4a56902ad15150431ba426d21d9dc6afe8c9
za49b928a002d9aa748c63799bd3e0b9fcc6ba838ed6cddc08350d30e838d42f667aa33d417fc2f
ze1d3c8b07fc063c495159175c36987c963f43f377def17a22de0eec7a80744a0c315e4c56913d9
zb8303dfb9f36c789e87e4eba82c932984d5adf693295554942affc4d5c1bba3d94a0e56c6da0e8
zf4832c61fa93b46fbbda48913d3f03508ca5ebe5786bdb2267363009d8f6e368a1d032d81d6f95
zfa80367004a13a3f0b6fa1c4a5bb001fcff6617c76d5d5633502c2c49ebe8c5269f9cd450a0290
zf78c91f71533db32478f1d8979890e30a9d9aaf76fdfa465447bf067a8d7e86e1f75b917801336
z2c20ada53613e9a2ae6f728bbc1519fb96fe2c02752c973335b1bfb82dcd135cb21eed011b4912
z4528c54c4da1b3d3ec515771ead5c605fa24e8a2a97f7c80e4e1c8867bee9c5700fc7b547b5223
z39e1edf4a99b4c137d1c6dcc8a84c658c9c8be0ea14d67e2775f9c7772dfb04c5c5c2729a7059a
z5af83fbc23aa174379fd4497594d646d783c2c34a1d53d75a61eb4fbc4146bff5ddbb2845a46fa
z272a8e10939e868a9a35f2a5dbc73fd90a0c776e2b5bacae139603301e8b6db91320e1a0cdfacb
zd70a1a5c6c94d43e8ce924f036d7c34211c8665d77bd324a63dc9f03d334bc6f90d77d210fb619
z9e5065a00afec9979c387fbe3e8b2b2df639458e227ff578a939df0e8d7264336d158f1512b90b
z13a599bb723154204d8df3b67264e9f9eeb2d33a125223d03f2ce6713983fa4513956aee99ca7e
z0d632c45d2ddae612569e0c9259753666b4497b46f846b266d745a4f7b065a0d783ff972809b1b
z7016da7d430c9973cd1d02d2d21023ab422e4380d19c5bf38c8d0fa8bb9a60548b897917575404
zd1e8a8309e1c8d29470e962c1574f83816970717f3cbbc6bb3fe1b2144cb382d3062f285c8e2c0
zd2069b377ffe8096a6773765f36d4e3d56022f8bfcc5e539d57bb1240b4a4381b7d05867ec762a
zfc1e0c551f1a184d7cad66f4ba217369da733f471955d6c8ed02502d242f7a6c85cda6d9835bc2
z92bd6aa01000409e2ea6d4bf1a309ea4bfe7ca5516c176c7f0483a0de2d7405b5868041ad32955
zc95ef6f704f899f62d92769d2af2c0a4af456f0709f72b7f12097cad7d925d63bcbd2aef2ed868
zb424f1e35454a09ca219568f089643c922aa0adf7055b834adb209b56ee5c9d8398a8841598edc
z800415a69328fe2031b12487efbba03c10ba7537adc98042ef5785b9ff4fb51487f1daa0e67281
za61380e492abf0496961d841c378bd8a92548008a2a79324be3365c504acb3e39d9608c6ff4089
zb2bff6ae3515ccde14d59e130fd286fec593863d80b2a00e925299cd757724c9c34f917bd83633
z6811a82327a385101944159d6d9839e6d25af7a0934010e6701d5d28327befb9aee406e75750ab
z7cfafca04aa66adaf8b15ef05d2518021ad80faa8e2dc826bd5b5403af94ccd780a818ef1f35df
z34323e6981b94ecaf0782c55990b74db6422f8acd6208e2be9d18234bf94d237e7ee0f5f793e90
z6cb8a511443e7fcc12b89fe387f3708c26b665073ba862c868903d57a90d483951b0bc0dee1884
z7b98bbca3aaedf6d0b571cba99c96a6bdc905ad04165e2bb2a0e1350bac7a917a58c682bf87d1e
z4f2414ba31038c04db56beff25a4c944d34c503c1a9098822590bce7a3a7a401b3138c89e35ce2
ze61f40b071426c004bf9ecc29f06509cb27e5355565c5bb70f78282bbdd4bb5acb43b25367f859
zedfb711abc28ef7e7c4523fed9a23b471410d5ba7999e6f964226c347a3a12b7bcc9cdc8ffa1c7
z398d0edbb1f760566f63566aa606961a589327bfb941a21eae48601740a0af4e8af7ec22c15e24
z833beef0015d5576cb60d183b88914316eec830b66dabc92f750cd7c40513de535a71f407b2589
z26e92783300d4c734c3149e3c9384e0cdbff060513e05864c590dafccb7b8e1288c7510c95a35a
ze00e14ddfa3e50f92066eb441cc6ba7afece8bb394a57bb3f5c08514412eb815ceecbacc5bff42
za51615d54c534be8c960fb06d6ea83db2be587b757eca1946719731ab894ba01fca0552d35c4bd
z06ec6ce843ba6379f95e9af81f6a745fb0ccf5ff53acad59b1ea4e2ffd6f06bb421202896ba7b6
z79b21533bad0bc6681e921378a2af38e3484f657bc7b97f1d1d73273bbc12b5b3540f54bfbc838
ze9702640e38f2d870b70992606ce9319ae70dcbb3513bb6079b22826f06b4734c3a78fdcf0c14a
zbf34df20ffb5ac8df5d83e2c5834ffa83b866f71dceeb5cad53682e39c29d9f1a8f803632cfa20
zb514a773685bb49a458e9855497e0a24f90f3e669501f09038e9817da4f2b95624f32224567c0c
z5d6649527cca5fe048b4865607efa1b85230611486577b2f9c943b1e9696f3d62bd207f5bfdbf3
za2c7069f4412e568afa7e91377299998a6f4f686825933733898ab3d6001ce3ae2e9b540f0c759
z4adcc656f2aedc5068d7942473ee7f238d7e54096dd02495056e9dd9c3a5242525dfdf8a4d60ca
zae4db965f1903add80a57837a3558eeb0f758154d180035696c9898cc27254559e6293d4827a35
zf3f85b2d76de10c34884b7f98fbdfc7493385cf73f8d4da0726308d75048c4d2999601516ce9b2
zd7afc5814f189c42c442737bcdff1a9e90c471257575b1744f477d4a458f8eb236f44e6ea1fa33
zbeb93f2b3568dbc8f8ce929d580054fb1c67a1ead8ba62f3448f2b9ab0f98ac82b8d04ebdaebf0
ze19ea12d53e8523721a8e15b2f0fd7b8bd9dae7fa0511cf74a071ebfb35b6da950c93756dd7488
zd12fc8dc33f543ca337f7ab03cc285ad127bf4ca803855e089aabb6f32bbd8322e0035dde66281
z3b7bcb3b3d7e81b5ae9dcbfcda12b5375dc8d542c4322366102512b2ff46049cd3d9d9a00ae617
z5f194e7ad4064fcf4fda1d8432328603a14610bbfa3e8c1c1516d3b9fc61d9ee8740bcc908947f
zf8558aa17a3dbede6ced99d49a227dc2dbb81a55529b7d27bfa8f0caeb9513bb6df29fdc7d28f0
z15362fea533d70592009e4320f4cb8488d22422b2a2f39ff5f6c2bc765866429c1ebd2e1293444
zab975f92e0713429a7fef2fa6c0ac88c30444be095074ca6f2c4c5451dad2578a4eebb147874b1
z315d709d8c304cc43e509ff9aed4f6a8b90e1aa74dcece76ddb2234ef04e63f11924c6bb0d451f
z278d38c06ae9a07022cdae00f23890b08b9029cf50769cbfba61978995db145f44fcdb258a157b
z7c8d8aadb4315d81ea082d0b9db374f39ce2ec24af09237df49bf6066087f62e57c177549d3829
zec74ae0681789b1de508580d005bdaed1ade6cd377059cdd73744a340844a16d9948908285df7a
z4febee7bdf84da44f8759df690a0256739cc8668601e7f8338c2bd45ea9a7eb35212886fde293b
zfd9e22ca77352f6ce1d16018302bad868b9b6a9c185db2d9bfa492fe95444960b057a628016a9d
z9bb1ede6a24024bedfe0a39ef50d9b761b6782de76d0973b725b76106de274e44a442376d21d52
z8bb22d4041b0792ce1cba4e8276e674a49215620aca9cbc3f102c184dd24d01fb7d39a99c2ce76
z9ed1a169907e8ea75f859244f808a61d30594d2a09387a038fe0ba7e027aa9778077b40dc95a19
zd05fc153e5b46f81c6ca474e4c50868b5e33c06f78fcbd4123c7a6440d8d441237916fa05477b9
z682cd3852d4f7ddfe4af7e869fbd5ce0ba40394523f8882dd7c2fe26332d73a105618ebb34bcdb
z164c4de139cd446283d00f679c8e9683f70aea81a42a38b278111a81e47e16c0e673ef10176701
zb5b1e90bcb19914cd936aafad13540c03f7b8c2f2901091d760adcff6ea511be9145a4e2db8e91
za9ac92fd5f12fbc6c086283dcf2525f39efd8829f89592e8d45c00fddb4eaf76f15aeb63305378
z2909a2132078393c950cc8b3fae2d5a30aaa770b76e423d942fc91d69bf84365e380f69f43d63f
z54d0307484e983ad4a25546ae828da6a41748f9edeff8f115834ce70981e547af56ce516124d6a
z8ae1b684248128bcf86d514b8e8f01e67673fd1c6e23ec3a08ff32b458549bb5f8f64c98bf8903
z0a42ce6cfae08e22ddd05cae6db146dbd504a8c1cbf8db795ca3cc88ce177fb168899c08ac48b0
z29d2cd096ffd2ce517fc1903b0ebc99a856407ec4d07164f4b1b4c44544f4ce82dc6fb198bbff6
z98e4a7d27afb92b0f12f726701e1614d1f5a7c7768e397f03d10e733f7d4175a4badb1301bd2b7
z357b512f20a97b5256e58432eb2342cef14849868d7299cdbdcfe03a8a47ac9e7ff702cfd1bcdc
z3fd247fcd6a0257cf7d8ef07e89dbfb86bca2095db4024b34c6a3269e528955f6207b9d94f3652
z38e1e19ba7490bcd94f0eefb32a348e7bffffdb575f9b5c3504b11e2b9463f0710c3b723c238fd
z29d15f2347a6d8667d0963d77ec24689cf7a8ceb5417a50a9977ff544354c803f4b9a1968b1871
z0376e65a75470491a832e04ec5653adae607dc4159c3c10cc6515695985f40eda3b0929e59dd2c
z9e9786f9fe6f3ac568fddb71807fab6bc618d336c791f94139b8f4366577cc4905a7e7ef0a4fd1
zc21b1b1f750c372128aa6b7e759436ffc79fa1c7839c36d0029e470514e3ea9a37e3d3a8c127d8
z21e3c4a572b4e4733de028360f311e2d1ae70157a101b9b02127566e2c05d7fa36334f9d46e477
z28ebda2849195c0b30041737039ce510b3e67c81b694717c3e6adbf20ba9bf239a829025bc8f91
z75602a843b1018740e1e490eebfc87adee5bb740d8e6b2d25073667e38c6817b6cec99d6ad481c
z06cac5a34247bfd2a72208f39ba9308a67d57416d91e2be641d47baadea4b387d2f36aa51d45ba
z1756089a398487674ba89b8fb944c6da650a7a6b195dc09be70d5c4e2072e042d75cfb9916fea3
za94fc98f90cf6ab6456e58985f5f9c140a4334359367572b119db64814e69f2b29304560293cc5
zb933c3ba2dc1221cd54ab29ed6e8ef8f502fa198c1418d396051980d3eb43a0370e778a386f918
z3aca5dc328549026fbb91ed1c991b04bea1e792945c7ae67f9dbd6fcbc2d54b6f0d1682315f0f0
z710437211b208585bb84673c1e1577374b2b0fe5f76219682f5ef4b05ac1cd75be575a4bfcaf62
z1e24f128167eb3cb0ec2c872485f2b3f566bc6b76e8ae02397c9b25567bc67db3c2d2d426a3806
zed59e68993acb7c56fc48b1ce1478c6d6ac22802d14ba2f390f7f1e2a3ab332dc20405f8c23d99
z252ff9b5c50e39129f7ff30138ec28769feea5647f2a8614e7f911982c864fcd4a30f30174ab45
z03f674c1e06a59d788b2b4c645aaefcfba6bf9dab1d38ebc614c11908178233fe216a17a4b07f9
zaed810807f2d0fcb5b843a77383b97ca91dfbe2642702c68b150e9007f31300c7ee09624696b24
z1b442ce80effb1be8855e44763746f81f5cd9f067f1a601a50a6abbac86d705c8073e5033da476
z069c804496ad646d62a87005d59f46a36d92c80e9acaea305d391244ee264f9f11535d95f3b6bc
zb3d4fe6bd98d39e18fd6eaec5f75a397eb52b3348c2819073229e31c9a7bba6dcb393e483a51a0
z0e34bfbba234cb46068380c9594f023de3d9ccadd95a4eda94c3b97bbcec06b814381ac74baacd
zaed6aea036c32a397d479f8c764f59a98a43d77e9ab402bca12dcbe4b3566de53657274120bd96
zf4d2ecd8c145202ac70cc5c7956c45666a1c1777d34b0fe8387fc70423746400921530729da3b3
z32a6bfbde78e706c82ca96343e4d3903a8e19fe52b8bce442e054e621d026192d93f4993d96397
za5ed4d229b2184bbed7c098af66a323fe91f4767ea8eaaf5981a212a0788793b3bef9bee9f446a
zc9218929defafdae00cecc88048cc9a8abe14cc8f8df8d3b3888c8a5ea114d3214aa44a2987b5a
z9fe5193a1e7b4a5cfb753db9d8ee297a7bd62fa1461a2c30c541555ea94a9599686e1ebdffeeab
zcff71e2727b3606e7d0d4d30755b503a592a7c6c6edcaf0be08cddd08bcfd1110dd7a3cd5314f4
zab9e6be8b8f4726f31f2f158db13e78334143a347e407d44ffb9330ac8223e03489390f06dfd7c
z1ee41e7c3ac569fda2551ba1548e9fd25217dd0f0b2d2ff8ef423c99cef812738d730d59a5e82e
z0e02be436f8756d7c4efb1a83bdffad51d322299c49fdc04217506e605cce7f28489c0dab17216
z97c765d046814f426c2118d5306dff9c7761a5e3333cdf67a7811df483ea062f278c03a63de632
z5041e8d3a9fb0e2250906326a211fbed52c1aa82277c5c0ad347a58ff8838755a322768ee45810
z4a96dfddff4de043c26fcc550887a2eff90cfcef9fdcf032d433dc8d6caca9980fcaaeb234408b
z0182582a0d062f71d0a9c45291bd8cc9e11b1b6f4cb56b88c5ece3f5ef967a45ab858a920ab351
zf2d7637b73f05886dd7fe3fce5a9657a26a3538a330b7a4076c3394011639f58ca3b7e5292638c
z6187d53ea2b39ab88f84234b17736409a6fc6e32e8c63e5a763327141a8cf77a36da844dbacbda
ze837938b93345a4bb8b18871ac30eb3469eee4ae2c811984ea18aa6d2cf32e4fbf9e3293bfa669
zaebaa600f950ac129bc1635573af0834a6d09f59864b382d00819397e5fa98c398045a89a3a9db
z5e9112c0410074b00ea1c416c26f3a23487f68bc1ec7e8ce650af7553e1bafadf8d3d083a96641
z3a1e36b72f5a73e29e793be8571652e36539c036b57786d1c0d2108ef77ba066813c32b4f74f87
z728cf69699b62b53d06f6bb3687d9c9b07a807288426e8289964b23a3f08e26196420113cf316a
z39a4f2d73c13e6ededf64fc04c67ebfb89bff3d529d922ed247ad35c8b52f3e6c036d46919cd84
z96bd53e5147d6fa453fd861600c546eec1319abb3d3bd10b71bbc2d40bcb04b844707c80375fc5
z18b428b7f2bcbed32c003dcc7b97473af9adc839dfa74adfc43ecbcd413addd844990f7200b484
za799419cd76194b2a387eda9c3e9c63e8a01990964a4530c2569c1cdbab79ac3dc57a00c923f26
z50d6f4e88f4d21ef44e01437d5b8e59fc1bf802a3bead79453977a54e14da03531ca6238711375
z4f25e2bec8e34e898d613cea161bedad87beebd8d54ec97394b34682c7db5b2bb84ecf886dad23
z207056c7309b70518bf1fe3348ed279ebf4200e358eb2db1ac00709b559e4c70637b7a7cc4ae46
zbf48bd85342a45603d56baad2f2af68b66143bd0d26c2728f2ad652d258f35437eed42911b644d
ze30d07e08fe9e053794b4fd6948fa0d71f30f632b55a560693fff2c00fa00e09c2f8aa3eabb671
z85d82dfd60c64985854d601dc87b66f84b3313d03a1a4d34cdf30438a9eea5216d0768d59b0267
zb1c09944e236ce1d9858e87a8a1928d481b2e1404e922838e4d897a49c80e2d613237823b5fc95
zbd9e80042d30ef0de79894dee1356c5b6f396793fcc7c37860d0e9358b0ea5a86dee6654871528
z35c19ec2fdf7cae21d274ebe0068facbc7354b4b5096125a6c87cdb4dd22b96a4a64c1adefa160
ze5770a3bee556be89489040b68f9b8114da6d6807111155c4348ea478143d2bbc84fa770ac2cda
z0d73ebc53324e91afd6eb6a5c505c7af3f4ad9fa2abb7e85bbde1e590cb28e8b4f8190c1efb09d
z709208006045c39ca8e81da37f51ff774eb1f7729c54d713b8eaa1b5fde05602b9ef857188620b
z51f63b24021edeed0b67811b015ac8741669ab545dcb3ea0204602f35a423fd0cfb73a27aeef91
z25f41656e8673ecdfc62fd710cbf932c243dcc14801e5ab08a54962234948edf8511ab9533d303
z730f65f479110374e7b657dc1148dcd64f36a96fb50ef0cc49adc0919be4a882fc014e112fb865
z3c573441d6c6c957b37c20e05e398d23fba3b0f88f8a0497384a65692fa70f6985bbba9c4e7c0b
zf23236f5b0b8d8ba83632e759721dd3c68375e9397b06ae47c25430468553feaf6f2b6691513a6
za9ddea10e836b47790f91a526d45010a9e17051f0cde2d17784c7b6dd37a82b729bff1dd98c8a1
z91f8a7c77f1f08e07dd90844523059f225344dfe67e7b4468e15f1694395e19b23be0b04e39e05
z2b38a55b1719abed10f0468d6525ad37c73fda7287f6146f656dfda46e5aff8f934192076711dc
z47d340d9dbcad107446d1d32aacb5bbfa2d804c6406068228a46c5bb1c22542f84155aa271b600
z3e3a971b9017eef302ae52ee51ca47c244d9cd9ba3d95755b25bece846515fe6b5c0072e8afd2d
z1ae1af3f47368fe70728d9b50a177e53b26e3632d02aad7b609c1a8a10e5f7bf5ec6c3212fb103
z9fe76aeac9597ceea12e5f959b66130f495fca9fa7bb181b9c3a440432ea8ea98265cbcdb72346
zd717c1078edc9caa84384cb754b94806699b761176380e03c614891e4b90dd75001f04f100736a
z924bbea2fd1bddf31309c014dda89b94df7720b4d8bd8fbc2de38f8e2c21edcbfe2d06b2890db7
z4032f1f17d8ca1dd239e779a903e1d85f969c9e637ef5b6637f927d3718ed9b77b450cbe52a345
zf6abf1b684cf7174e00cfb4a6ca4c5312ec07e361382e395992a853e317629499c67f7d5fb8771
z3c09721ee5008fbe5320ea9c1d1a0a89f0c8176f9857cca6e65124bac4f9f5fc14b96e02507146
z66e436b7baa83b4070094d89bea460f6ee12a3707622ddcce4e0aae9f0cb3924f11f48d688c93f
zab5201828e59a356c61fcce5e2335e6a27f55ee5a9c85410d43aea725a273d5d28c18e9a8bd91e
z2596fe6f3541aadd1975b7145bae599d09d9f265e79eb9eae0d004f55203ebd7b2429eb26f7e7d
zeb1402ae9c0bcc81ab96c21655b4f8273686dd64d151c548bbbd581b4d13b51c01926969d22b49
z2e473fc056998a0d75650b29dce6144ea9761bd5facdfe5a37e98af95d989b662b92770eeadab4
z4a1cdc2f6581d8713fba81621b5c6a9126917fc0423f260246a6de029bdd27a77883426867067b
zbd43ed5c55169a7711895c8f6b00315295d9e7d1e6646db2325e616262e570611256a0a62a0aa2
z2e6cb1ee73513d694bf91c8fd38cfb8d2038ae14745e3a4eca405df77105851d7c0a1cbcbadde5
zfe0a999c4ff995c1dc0a56e0803cf724e1ed9a7d40db266177d037b330a34277fccce4fa720aed
zb63268b11fc8c3dd436db2e7e0f8711914f549c86e30ac51b05a59ada43b2bf1244ed3e2fc91d8
z239ba068c448b7f7a960cb0e946fbaf3440e86ddc7dbb0b87a0bc65b43fa5d32766b6a58999017
ze695e15c844ad02be44490598e4fc9cc8ef6766b540880d61cd0f59b97917edfc893c2834e266f
z34ef7892508e76f4b53485bc4a475b83343a1f9b8106af38e776e306b9e453c47b58d8cadca085
z8658e9ab41dd88cfe88cf0a669cd2d85818a1aaebc18fee6b62bab10f47034d6d0062450d1924a
z74cafdc367a782c018c0ad0279de2e4aeaed9dab77d9546ff9e2585bd0bdbd5c7e645a04427ed3
z896318956b135f75f8f0cc1ab0fd715bdd4a544466b0d1595f5932c2b4c1130d521336eb6d8cbb
z3b6596728be6b262b3701cca93a66656f5a02fce24460bcc6d1ad6541ade8fd58a298139e195cf
z2809f5623f1f2311e54eb32affe647be8adac9aae985863865ed2d919e16ed4f103612ff81ebd1
zcf9979650d70ff4db6f8ac4c1760746db40daf0f906ee3348666c799b7c987c438c659e4b1fd5d
z3c02f3728693ee1ef8b3b29b2271306d9a11477387869b086b2cefc802bca0386918283c0a5a73
z3ca844fc73bf3b0462ed1d3f84e271f9ffa86ddf92c25d76d7fae6c972300946005ce76acc9c9a
za36a234bf06083e2d272a7f284ca8f216e646781e3700f9057cea977cc02394c3e986c8bdd678d
zcb67163a426ed43789f5db4d2d8e39db257d8014401ee9c85c1d70144935617d852028621c5165
z7a68491b2ce6c1104511f200712dce6cb7a324206a2f305a450674afc994a355e9adadee421295
z742878f52b5e80aad4a6517fdb1eaefe3b37d6c728e7c03b62705076bb31cf93bd3efb28cba3a0
z56e898b837d54189bada825a06636185997db3a7b40801e375f88aabd44c3a0c378273d1fb5602
zf6a5fbe1452b8388c595ff828f99f56950dd88193aefcfa0014db0ab85975189a811957a801d3d
z0d300ec3d27004be19833386a995dd6886d1f6393c5b3b7fe9e54d0028655a6d1d927d6be5189d
z078036624fa198cee3b82818d49b2e27b7040284dd83399b33c15e6fc537f51c2f79a1e8d402d5
z4cbac16c69326a81207cfeb5493881ab014d5037adcb5c9a872096cd2f6d9268f6300feacb21eb
z93d468e796a5975e7f905586270fc43420c893a222310b1fad3bf615d8da2b3037cef66d59acba
z59f2f4c05997b6522b0b4bfb130ad3aaa21207cb29af7c1690d5c7b0c849f9252b07b6b6b26835
z60ad3752532cf8234645501902271a1afeeef40c6d4fd1a7099c556cc7a9ec6df4d1c85cb21244
zd1281191d3549f5824ff54db4fd881a161ff00b3f3bddb4ad480f8cff07ffdffdb7d0f21bfbbd7
z61550ccd67321ebc1d2f3f31df570b832e1682e31a7f2c42ed89fc2f086035ca03df6e551e52d0
z695351e2b4c1b565c9b9a47ccb98827d1701321a3672e455555c936b640a8803359369fc07db07
z23ee16e0263694780a85c0bc46a3028a3b10410b2ac4c553cc0defc2fbd7819480558d884f5ab1
zcf69de346ed74468dbb2e80e79842eb8e1eeb00aa0c4578fc985af587b3c34f7c192f8feae2b3b
za535dc98c153d7f68d921c59b372432a755ae450ecdd1a58af5dc0d0dd73f2cb1d18940268b316
zbcff3d4fefd42cec44ec20b8092cbdaba6754c074af4f052e7909d9d6077f09b37b1a953b0177b
z5cec1e61114e167b9884727b859b8938e45775d5d8bc32b7ee5347ff246329b6cd255b0239dfac
z5e7e9a048ba344be347a8e3ce563555de2f189646dc68bee6e244549ebbdd5595d3fcfe9362759
z09b437ce85d839455f21f0ab984c5629a86798577130827e1514c7ea0a4e5b722daa362b357550
zf2e741d01523372caabac1b765707a57dc8c9369abf6c0fa6e2f3c590dc9a9c50c50fb6bd20c6b
z7a40f4e4b1e2a269b1b31560be8566f42c17000986017f20806aad76814a5de2263fe15cdc4e91
zd1a2ca6132a5191dec397fd8a35d4d5e9c3ef3d3481cf91223e8072e142d2c53e0106e2b996ec4
z5f94062882896ba5b98ef378e0c8a74c6ecb61c73b6b151694824e4ae85610f0941746bd178fa7
zcfeb54c2c9539b267aaab8f4dc55a06a1c24960666738715e12ea4727e1893e548f83345210835
zcca7336c7079dcf5b80d7440611fd01e44430517bc96519aedec74e22515cbb55790003a33875d
zac7cd311bfd2cdb36181c6eb264618f7e6f47d54d03060a31153c7455bc8b98b6681bf9ce59669
z17510761cd0934a89675b88b093b1d965e3043003a46bc70f808ff99d5cdf96ea47689f97054e5
z9a5422747e4329f1685b5ed3678fd1807b3996ca28cb28d1955cbb5f8144aee4a59e1109e6f74c
zd4f7a9eb083325ee44feeaebd3bdcbb84a08bc7929b7e80221faffa0138f192251ba88811b928b
z7615c5a504c2e2b22e2d0883421c2624fcc269430f275cfad1076a440e7a391e2777e9370120d3
z6ee7dd2a00e1b1fd36e04e2466a5940b2f4191e6558e0c4b7906c37510753b9275220da1436463
z8de32ebc2744b6a38cd8947ff9b8db57c9c7930ee4a27c4291f5e240aa0b6374c1c72fad875218
zc59536262c5404fbb8c4aeb9f9759d5ddbb9485ecfb9378efc7ab0266a4adddd3ec7d9381a48d8
zeecbbca6ef5e59b7b8660c55297c37887d1db3bffee469311b1f8aa3fa6a86565c6c210647908c
zd0d012339d06b763e2fd071b402635b589bccef0b20555174d805fe88f79d6a93085eb741a5f54
zb712f5a28d2e6358bc38d008d0444ad97e0b2ef445f22905fa73d76d083c964da689d036662378
zadf599411407da63d8380b293dda5266e25a4bb6d2ece823e44dc6de3ea72d5fbec2ce2fd1033e
z6880a48e46c5fc02b3c9402f148a926a4397340588940e67b792dda48d1845876c9d3ed0672626
z1e58c239c8cf5ec3413975bd4bf1cd109d61fb1d9ad705c5059b3dc8cc527d23dfccaed5be6df8
z15d3e10e1b3637cb7c85333861cd735595fe64ad9798b2e3ffdeccaf98cd37a99f326882bae793
z5fb4ea8b2a55fa475c6cfe2b91d6928acb3bb355f3f68ecb140d3bd5ea90c3bdcb0d8b37eb6adb
za97c303889a55102a10d6d660f7aff85e63a1197a919f5cd157308e21ab58d920bd3648a45f00b
z467e020058ba8b6c9cc522805cde0bb17e8ca038ffe33d654312c3af9e8bb11f6ff157a1e10785
z5bf748c409fa282340290e49f0de855dd820dafa77db8d27e198ab197526f57f106dbfd231d4aa
zdef8e344f58f8df262e12e6a383f3f1da7b9500c10b3e80ea732afe6ca0bf281c9469d551c70bc
zf2f45269f4c8becb7be604ee6f4a18efe1d5c0048e567fd329283a39d0d53bcd376271f5d46b34
zfd16b0ea8fbefb8b79e7441fc8c00be2f46267f743c5e0d29400d7ccc45c20acb6d706219cf2bc
z9753c4eb69f10dec88a40a14ef968a7969e2d6d0801aec90bd8a7a053741c39f778a0a571907a1
z3c129558f9607400e87213395b815c1a0cb13da3d4b488c099565601a37bf37b006bbbd5393e64
z075f8adfd183c0fa4ca948ac89607f8296a9fd62244c78fa35c296d52c45e090143e6d651878b7
z2c8b1bc8f52d46408a2728abd19bff974c20333ee55944feb08281064fb2d53f4a9302040b2f4d
ze129a5313ce495cb71789382cd908effc87faf6952b12f5a3954cd63cd604f226be75fc560c1e4
z24f9298e5ad3316855ec6b47abb5a4ad292f2c20a61597d1345c9f866e545859446bf3ba31cdc2
z03351a647e62dbf6bfff8c9f541e97a693558c308fcf331e7cf56a5595698204bca80a2a460cd5
z6d9930be1b00bce89c2701d065791198e2ab571a8ff87f7f1d6677b890d6f460d3d41057f1f432
zd2ee1f8cffdb314c9756345f88234e68b59b142895e76c1e1993d34613601fed3a4c0f7910fbf8
z132bb4c87d5242cb82870d8d34799fe4afe5fde23527d0bb611064e80bf82f8e5cd624fe9e65d6
z8c04c18708da9d7addbba5c60b64d9e5771dd4df8a566add2db12cdbdeb87f6273206c28fd097b
z53750749150c698f3503c666f8294f62a956db71d59c4a9ccf4cbad2163e4032254e16ed5dc465
zac9dc4c4036d5fe6eb7722ef4d260b30c53f9f2daeedb927285078ce6dcfa39d7a958619bdfbf7
z85fb70add2dcf6d2058f94f0cec7c94ce9f8887aa8f1ef051a2b618b454f639c2e3de0b23ab0f8
z0298db0f140af4606505d0a1e0337fea84ffbb3bc5bdcda841f17634c4ed15ec756107743700a9
z768ea5b76cd232820e52ee52ff123d92dcdf95dd92889db546753c1a1d4bd7466a323ceb5a5bff
zc9ca796a6bd5e347ad93a1d764d65bf89649a0ccd1c3de2dc735cae6d2177cac3f210afc96c4c9
z3405c37e9cab681080d8e118b989b8e6369082a278213ab2934fbfa50cced51b2a987c563e27a4
z9387944f5bd7ef08615c27e94a131214775c962b0a137e116e0b6268cf5be996cd18568069ad09
z9961358ca8c8b33948ba41304bec449aa985a502b80354d0a1f83c79ac3215f3d9877226a07e7c
z57b633c6139bf4dfff5c442572532e74c927f847e2466c2860653fe10f32d71e849b261d6f9357
z1d245e0e82015dee48f40dbe63dd816a4098950903175957d5c6a93c405817838da41141d46b34
z0ce526cf46f383c0aa4f74875752b53d23652837e46b4e65d93f2bd8fc5c4c13cdfa0d7b1b576a
zcae6991f0dc6af0b10960b1c401256fab366695118198bcd58cb5990c20b84065b033deb9c9d64
z3c105b33a624da31bf73d0ba0b6175506e0ffcf4a1bc26535f2ef1e13f12df0df9cc2a2dbb4394
za0023bfeb95d755636d1d46cdd09e3dec24d1ea9abf5189184cf152669651475b4c98cbb7b5f9a
ze8691cb205352dfac2b2d7f22b0f9a77484cdb912393c618cab9bc4111e76edd27b2d1ad64ad27
z763626af991f6f5cf9b27e8758897e36845136e11f406cb3b30da87e7ef591f8f5d5d8283154bd
z4548cefb5f4a45742c3456cfa916e1f0c9a7c702d63bb8f104a4ed30dcdd14278ebff87b532762
ze8f7737695377f549a5e7c7174218c0238bdc20dd2f789ac55cc8b5d800f82e0a98cb79fa0afef
zd68bbb3d7785a71c9b22069a50b8ef9553788d30d826c4d74efdf13aff16b8eda511e04deae496
z1b36091145fc083140c34d23e5fc112b1d54a8a58dff51b0bc56b388ee3becda722836ca6eb747
z5cb370a9c6a650a50e9e8531c68e2cd89a9a551b499a2ef5497052ef250b6c9eb2f2f2fd05ab2f
zf7ace87e174bfbd52137b7febe5353ba6cc56478cf9f7c48258a160791941e45207b813064292f
z6b944fc0f986cccf39610cdf0a9b145b1e308b58248a73a1fcaf924316a7a22c9d8132e4214b9f
zfbf933351f27283c5b56ec3da30908d7ac21af8161d7eabef98bf7f080399a8f0c53dbed9ab78d
ze4cc7f534cfa94fdb3ebb49e8e723df8ca465d2205d5e40846fdefec23c29a5ed217f58b5ed61a
z603f3df0ed79e24b99db483488cbe43c57893f45357b534796c1e81a503314a618a2b5c12c3b9a
zaac32d2637934b96d1d743bc627e1501ac176fe553b153f03ccb033fe32308e476f01cf9243b6c
z8947cadd66d23f6b5206dbafe3420dcd67f82960d8af9d2898ec537165e975725f7640627e9af5
ze7a1646798f84eb4a0a388ae8549747cef194960d403bec9a17f32639c101f4127069e1d3604a8
zf472bd28820276766d291ac7ba7f1c5f1058d9ef22a228f0cf5cc9e3521e3306ca084788f8021b
z3ae60b71bc6674eb0842059fdbba8d9fd0688f3813abcead7ec5f7d9ebc0d852c9bb6bb86ea445
z353644a62a7a647d522b5cad69fb857a2525371050a0e97363acd32ae053aea22dacf246189109
zd243dc8ceb7d1566def94963da27c805474955e69f8e4a74511f41d9f49dcd49a8aad5250384b4
z613ca3006f53a861580cde6d4b33231283e063140377f9a6fa50e72ef0310cabed30436c754bfc
ze0762268b2aa5f9a4370a80a97d80bb5a8c4d738223cc5df7d7de81cb44736d000360b5d7b169c
zca6980512c854f35b02221e7912f0797968e2978675e126fb9048d6cb1254cde8450371de305b0
zf7e542188a6998db2f788ef11302362c15d0cde6170a4bcbf076c276e5b076b0dba0960157b7c9
zd4c517694e12fbfc4fa596274d1ab10d17e734da046eac58ff4ce34027ad9da479d3754b3796b0
z3c1595379659279f1cf8c2335e6c37ca3d966f3d12232c150a27b5b42e2c0a40086b0d9b04af94
z417b0171fe7a0d70b4106929942f0ce0f9213dcbfdadb0a723948e98990e854594dd3aaefa5312
z74664d13a50ed89fd1e4ce8d28d139b17eb59cf386492d0950371cb0f0883e1b716d6fd38ef7e7
z66df4fa7bda7b14d92e0d3a13fc294f7cbc2a946bf0589315e40f37a2692dc4c87c14c7e161018
z7593015d4f25761ac647003213023aeac20c90ad88d8ec99a0baba22b17cf32d0b7a338acb009d
z1d662d0141643231fe37831f2a3ad27af8513693dff34555b3cbe3fc40eabcaf8a251bd3dde84d
z2b2bf3258746ee7b4d02b9b1b188ea3b433ca563c3630000b664327fce4b09f55d8455267df291
zc723bef18dbff34d5bce6301af64032590c1f52131be5920878ecef9f54fb8fddab5a2c1271571
zc24c4b89a08994ec2acd4a7586bd8be0251c5de456c79de5ffbd525a5b19e54205a83f5afab67d
zf13defa87cd45db37c6eab579b8e4816a9dd925c708264713edbb227a4d54e7568c21c76d54078
zc40a32ce5b28871b2f1cc89ce3d2015c59483e96971916f2498db7fa6f3c26ae3ed0e6f4214da0
z3cdc44ab086da00bf9363c3a738eef48e17b3638b6c257c59bae0c3a9578cfdfd76aec2bc8920a
z81787877af38c7ff493717c5dbd6d545b47592ecf05d6620b698666b81ef2109adcf1f3f7799db
z3b46c59c80bb68d78b5854b31b0de92391d44b9b0e012101b4227778afc8cb3221310297f6e1d8
z7de46e9d85e33407fd1a2b157c659aa0188010da95d74737c48a0193e54119bbc84b0d4b943bad
z2e8dff88e3de8d246e4f6466a1835f4a350660dce641bce31f03487e5a4962c259cc59e1c2fe75
zea66b783d6c4da8c536238ce1a28dbeae4073caf12fa3882bceb636871164835039a97f4e0c80d
z7e061c17fefe8504b0cbda3f65d10bce4cd731131f7cdaaa26c997dc93d7f178c3c6040db3ee83
z670f386c69ab50d3cc0a45676fc9ddebcbbaf6cfdf693c40df23c078f1d1c9fc9a52de2ee848c0
z1405c70e02d8218d6c3d19e8d96e525776cd76f5204bc7debe9e736709a4d596a6bcb5e969dbf3
z617144787bd6740e755cabcb2ee8cce20c5cea2debc565f1b85fb999b34f943fa5f97f3a1e160f
z044ffb61ddacb9cc6ae25b06f6fa7dfe5d800807356e281d981abea3628a89659959e22195c97e
ze514922fefff230a136c9bcc09551fba998ef6af5b82e267b8d8524e4c9bfb1667fde5e9ea53f0
z499002b156795d5ae7d6fc67daae3a37a4e2ec1ed672c2b94a15f889249de11b75db99f05a0e9f
z5bde13a4fa7b0278b5947718ef4b7a65483046158ac862b7e680b2d90012b7c1f5966ba2a88b59
z92638b44286dd73392d4483ed28e688a82eee7434d2f858f1622c41d5f382badb0537178097de6
z923557d510c737a477d4d106089cfd4104c263f43ff3d42bc0b78ce480016f25ff95245434f0f5
z6e1988c4ca3a66b3d03ca8288ffc383b1fb950e41c044f568d4181fd231e29d8de31cd0fb274fc
zf337329d97a6b8595b123f09189050e6726401a557dd85afdf96bbe18f044cd8a7d069255a0259
z6d5562c167fb54d20da06a6a0ad16efcfc4d3123f2a1c827821f0e18cab9dbd4a812bfb58c7d15
z4519ac1c8c09ff6bc492b58cb458f421ec14e2b44fae7e16b17b4a43c4e5555a750a18668e9601
z3f4a227cb107322853f0a1284eadd4e50b13508367446b461c2cfa5b271d00b38aae5eba4e1946
zb4e4f5ca57befe9f059d2b255340d0689e59e97e131759faa73cf6feb1a3294af93c4133bd502b
z09c3c33cf61e7c475d253c3a6ba775cd1b0aeb8ed019a8ace0d300ff72011231fa4cd55d5431df
z0153743931dc206f1e156f57bcc485a1792a8a09d5aefbbad37ad1c13d80e832cde75ef865452c
zfebb39d200d9ac8919e315ff66cd875d37d221e32e81b4dd3a1b0f9a45491d7a5e2321d8adf7a3
za95545e71d18e934741fe61542bbe98fc9d1167aafc991d1f4366ae21f4646c38ec6a6ffc9a940
z7b1988f0f98b456e7aae4bd57df928d70b357ae0a5fc46f07e0dd6b8bc3625aff247eeac892f46
z5100fc1965d28dcb5e2ec508f11c6c2c72a5199900b4d1e831d4643945a88a6ccdd3cf10d15dd1
z3da9f599c52a1993efcd99f0f41eea72a29a0cbba34d705990e07d7885853609dea00d069385fb
zbcd466de4219cf92e63946b318c5984c1c6d8d652ab1e0e04c025799cb0d1cd3652306c1259276
z710885431941a6eaa316d929f0550fe854f1f70127a0f925886054b376c12b9b94662b8b9c13a6
z5b03e148522f5b32db098292bc0a670cf5b2415f7c3eaa1b5d51e40da0510045e92b0201287a3f
zd46c2fe1c3db16814d9f13d029a1bdf31850e5741747174d4fd061dc2e81e336f5aaf1ba5a4426
z1739cdacb1b80dc51f94a9899e09fdf0d5db5f693b2a75f74a239ca192993fb7b379f8a4806e97
z5b3ed2e2daffd578735d67875003a2e10e2be28f71de2d9880c940ec7d55dfc7c7496220954d8f
z1e3b3e608835c92154a32635a8cfb41b52b9a7dee487afd9f65687ea6b1d6157242b2171d646d3
z368fa5f53181b3d591650c636a30284ce1f5423c21277bf44bbfe537955e6215150e644d8253e6
z61b72ea7b4ca9ab601c08aa94aa23ca1c6786e76b6ce9188efee1183f2331e785ad2b8ccb49ab1
z0f8b0952f49b059a42a48a6cd37f24ae31e094b560e4f6c15f4ee70c97ffa688d3e91f67bf4a81
zf6e6560680a339f83ba641c773608bbd126d049d0440fc59bd1058acdd9029dffd80ed7ca6bd43
z4d97e998c23d8a9a53975711105802ccff2f087bdb6e35aabc8b69c5aaaed507c7f7c2608f91fe
z3fb21b1d3fd73dff11ce2f525a42d19b62d4c7587cacd902c27ac233b0b6fea1d63d87d201c6a4
z93c11afe04a9fce40294efa49dd570e2f9d93d950476a079215af2a328858516fd732610e8fea9
z0fddb2e2b4e40565bcd85fbcab5a033981fa926be3d6cff56215a111c9113094cebf08c23cc907
zab3ab9e082a07bf681cc47c7ebfff86320a1e4c0ac3cfcfed89e637d116b88e47ae20a4a56ab7f
z12f8af535fd8e0a8c5a4691d29c05843337aa90ee2ed001dbe4eedc010ac67b69d6658660a9cc9
zdb14c13716e3b76a1db4b9223d31e019c24ae64b36c951131bf169f273640c75931039b064686a
zf3f7ef298afb7e642510b0938495033d8d1f28c0dea44653c5e077ce20e60cd7d80c99c21f84ab
zd8446cc4d82006c48560cfe7a8d961fc26ff67369d6b86121b1ba24e1e1289b756c2de3fffdd90
z6f8435d72cd901b4ba8c0965f0a4e9fd63f0798936b0aa608fd21d8deb582ab438f64774d81d92
z4f1e087ef554d0fe7983ba2f0aa9b37429127e9f8ce17fcfb03fae64bd9c0ea8769f4e1da7c7c3
z8f85066386f3b2c71033c17b0e07bd2d85743b0f62bb8c2ca4157668a031899b44681fe543a7ec
zd62ce67e464dee1c03e8d7f02f07ece75a2a032a0253f4b98376f9a40927e9e418b1a5fc4901cc
zbc00ce150d983e8502e441fd470b120c67dee55fd5837246a84240ff8d877f5d75a90240a73a44
zf964daa7a4c595fa304015c2c7cda94c2d22f80d64fe01b5357461fd382576d35f449daa76db31
z373d732764e11532a4b5c813afb377dcacdfbb19c7c2aba250a094bf954b5d77427e5c236c5d19
z7ccdbf7bea1ac2c52daafee0afb4ec4618b70115d9e77400c5fb133348a05174ab632bbfc44e69
zc4d4e256fc8c62a650df0e9c7e46fc003c5638fbd1b833bdf7b88b8f26e512eb1b434eaaf34e57
z90cb9df3f280f205750a0da6d7ecf1464bcaab16516abcfbaee076df76b5e6629daed52dfbfba4
z878f76c858a467bc2f1038a0b69a335f274affab56c0eaa2f6abb13f7724623201a1fdc1ff4f99
z88a9a5b1ec5ea55964af00816eecc11ebf108a7471e3d92bb334f4f5c49dc6251c71d7e986dbbf
zc280312553a7ed1138f320b818009f8fde3c3c56e810f84f1d80be5a04e2e30c0d888ccef1de17
zb1a01d801582bf5cc25d420744db34daddb93b81cfbf5de8919fa1e7ec5204b90d8a29a57f8b97
zf22ddbec82629b131dc48370c67bff1e64c7312826b2a787ccc2acf2de0e11aad5d90d289b632b
ze9cf9242176392431f7a55f73567e369604c8b95b5f7f0a84b519fd6e6cba8c41064c2bbadca66
zaf64fbbaa65219dc2059f1c45c0b80a79a7f4b0f473f1604b8cc5d8dbba03dc269cbf197207294
z0fc4253eadc3085037b3250837b9a694cc747ddb0367fd0d6cd70a90a02439436e3236aa617368
z2af1267b1251b6720fa6fa7f2f01a95d318ef7d64d25f78d8cd4ba26fa8860ba0c2c02cc1d1b8b
z4f1d16eeae0750900f2be792ed4d590ddb9ff71129403cea8c4cae4c150d6a255a9420fc90af28
za9e4a69bc49f24d7aabee0fad5ce57546b3b6fa7f52362135e6f75da262e46ae0c712e19ae81b4
z6395083e117bcb76b101bd468c83783c84b64312e3af1b585e0e8765467036e54b68eb284618f8
ze3f7affa5afd444a6b15716ed3bab48c90f60fb7cf49d78b6a67cb7d08433e6f35ff23db7593bc
zd7d7870293abab18b7d7a6896dd377640179f58a0e1d10a8f2e030cceccfce236bf1695a1e1857
z2b95b87289edc82fca3e6644b10cd2dfda6e3c36012d0eef24d97e160e667fe72490c80bd19ebf
z7636c1e0a4ad9e12c492f4639e4443c63b30984ddbfd9374c6a9885bd8a5c10762839fd69551b7
z477eeec87223e681b5c9dc1d4c3f08aee8fb8d9110aa6c1823fb5ddfd36ae0403432a3f369897b
zb9d56668c5695b7c5fb169a9d155342dbfea091772443e8b17191fe38de39b0dd41e7d0815cdad
z631acd8c08bbe0f5ea75a6c8091a7930e622387beffa1ef5b814402ae62920eb1a5ebfe4e9fc1f
z70f927ca473ed60c55ee3f6b6fe526d8cc91c9edf399fa00e6c934313da7956bafa3bfd29f6f74
zfca26f2bf1253af3fbdeb6bb72ad8c8248c3a3159046a393bbed88f20395519fe0c86286b4d309
z91f0c3c58150e74db1198092fb894aa136b6d78bc7d6dbfe2529099d922e7f68a0b469a91410d8
z86fcebc6b23318f8a8eb889516741c5d164fe5c06aef1a04f93ae2fb87e8a9a012de5ba0ccbeda
ze5bc58cb16acf26c4a846ec695c90cc3cd93ca81cea07dd4651a7f6f508467ea35a574ca97e8be
z6a8e913ced07f1c8fe1ca71e37adbf52471809655fcabf77a98118c297dc9491ca616fbc33876f
z7c8ff2701046eedc4480237aa0a4a9b1e1094ff3065b8ec949eb0a6533ce960729df1661958ce8
z66f506f21d2b197f08e0b014ad8ca5fd40d779fd871a53e31cee04a26d97cff81e15c2ce1a1761
z8851dc5ed1708ffd9fb09cbc81234f5f70974e26760374bd30b23f9e3f60a5b7fa7dad1ee69f24
z5997cb91d11f9b4a151059d33cc3cb5f779531efbef7e17863d688f41d8ce2f8728ccff977ef97
zcc06a3011ccf607b70c641bc1c03763da038350c93300f9470a7bd04daa1eb3547a07a53a36bad
z3278ba5fc6b3487302c2400419cf076c295607289e7a429ebb4d372c7f6ccc79b88d64d66db381
z0109620b6ef9c7bf3fc85999a89059ea6add4d836d73d4b04c80de20b0a3c0e1ebc673e43f578f
z66526a4ad5e700110848e81407483381c30bcbd0451c4a07366cf5afd090b5e6a2ae9fb29ccd75
zed00ccb0a653872b8b9e1bc29948244f6ed57b6657bc6228b2d4370da545c590751ccb9282018f
zb023fb8c2d8f381c32529481f601601e0fce6eb3e7cb49f72e0a2971d8c45aab57941f02ed75c8
z755da3cef6f4268dc442b6b25d956ecc6539ea24683215aea34b32a87e3b5af64d5d6f545160c9
zde3a3385de4dca2cfe1fc9b6b63fef0277e421959934d91f720bdfcba759999e1e1673b5a54983
zba763595ef6d536c0011c265002c5e2bef4f1edbc29de5d303c0f96b1b87033970dec5f4599746
zf99be2414dcd568a05a502ceddb9216de6767573e662bd6b42a6308553ec0d5c8b085113f7d58a
z8fc1d15105ce09d1c356de60121d272f426644ed74790038279dd03eafd1901eeac7d7f13c3b96
zc8472f6c7efb2f09aa7683a43968d6a60bb632de2e2a5deff09279cc787fb155b9b94b4a2089fe
z668f4bef3b424a387f610988a39cc5cfe8df8b7e5efc249a81fda457d8b974a3d39f6d727c8112
z42a5c422ad3c0394f75631661cfa58d1bf6c427cdd039205a390ede58bcb4bdc82d071a995f263
za6b1902da4c94c48d10c9480f616e0a81e6ad968bac1314ef6cedaaba35de82d28296a0e8cdeea
z4f9dfd5026a38bb975d911b3903b9e373446ae3b5e5a412ebb9d4f45f1222bd37a4ac67e17ac05
z6bad1e31f977418b4aec556cdb1b56347d82af0604def29ab0b190770330757e553d47c0327e1f
zd0d4931a285f6417efd0af435c9617f23af157c8a04b0838d42c29ffa9e6ee6ca07da8f9a52923
ze6d810f49970a348c047991c090029e9c9fbdf2b94a1cb0431d769050b7315a04747c13fca1b2c
za7e55c803df61bfabb0e85330611de9b60fdb376c9a9fca8ad59c9897c9de7c6a60d91a09cfcbf
zdc1203199f2fff5dd1a3a82d33bd78724702fad6b177e0a87e2b988beaf202015f3bfa2b19b17d
z34f9a0d512a0ee6a6c2d382dca37b2f30d7ffdc3a3fe38e431bfda2fe060de10cfe92a8d22e50a
zebe4b08487a14365d803bfcc7349d9b4d6ed721ad7a81543b6edbffafa71291e93889b3306eb79
z1c5c99e9edbf528cc31ea216f2952b644ec5eb74252486cfbecf5db5ee5155f6fcc9a8b18543c9
zc457e5f0659207abf6271d416e11c3862fb36efec96149f6e65fe39496ff8fe06e10e3b96da152
z785854f1a70b1bfa80087079dd71f3c0526c071da15910f286eb0221a97c70b2fc58ae2e2dbf92
z7bb7ad9a01bfcb792b84f78ab9f00287090655deb2477b0bd430e1034abe186f081454a8c47be7
z5212974df28e2a46ea602b612b55664a7c84b834747ed57af8c38318a2e7ca4a8877e084f090d6
z92674f314596a11120d3c423df7e09fc121b6f6fd23d766e6a5d412ba1b0dcf777297711bf4b86
zd904ac8401bbeef54059b299ca8e8271683a519f0b823d55f493a34a44284bfcdd84abcf1de0e6
z1e6bc55ababa7e2aa7ea6d20aec13edef3f094b04d227c52b6b231372bdc7265eb970382a384d2
z386ee8310b6ebdcc1e7460284590ab38e5ac2668981ead1c255363bf22d229be07d552b5309641
zce4f36cd4473bc1e68e6a0b2fccb8359d03c33a34ed1998039db19ff8bb6e7b6b692850e7af6e3
z2d8f2081cf63615afbc00807b69500b454a1abd2c3dbe6b87a0a882dde1840b165c274a43d5bc3
zdc303540444ae1c6574a0df9ab05ecd2e237b8c5d6f3d4ffe868f7f50cab30d583e14853b38af3
ze0a4b1779f221a0beaffdae59c9b6eb2937c263b0af1459eafce671607ed6601a2428ac9d4fcde
z19dd1d5c3ebba2e8d9998f0ddb50f84693601f06752faa025cde4b37dac86bb354ff9a63a6795b
z9b9c52d25f80a68a2dba8a75168a359d0dba7dd125de0eb01a3dd444dcd14bf5c300ba1c0e9d84
z9971b450c2fc73d9ebdeed040db235abb5da0ac4170867b3841f15acc395f8af91c87a15c8c657
zbb7f73c7ecb7ff9a526a27cfd5895f099a938d03d44d519b51ad7f67a30a2d273cda7fbc1de2ec
z23a7f4b6467ba41ec830c36732b55105895747bbe2a2f2e2fe32ebf22dcc6dcd455708f9ea6f72
z8da9306af2e1c84162c19281c2540b206e8d40415c9f79d41fd1babaee0fcf4fa2db230e3e1a35
z570801a6d5de4d0e8cf4e8b819321eaaf1c75b13c95f218419f582e059c1ecccabdececa35bb12
z4f9f86ea092eb4a6929e763efe5ac05916de8908635b142372643fd753e511b93a66e78df70e74
ze511038a5b8f8a8f85a9bfa5fc7287dfac071aefe894229ec2e881fdcfaaff0b395a9b5d68d2d6
zd5215ee58ef6eb3f1f9afc6f642a4b22b45d23f3b72d9677f3e4a4bbb5a2b1be1e881732ca992c
zfc1656b82b89c01255cc9db4828b577d72b4b096fe22d6dffe029c7251097242858f9b585f5cf9
z91a2070c347ab6ca9936fef7eb4ef54796dacad030ed0f3c0e67cc066202df14307a035c93c4bd
zc5d567906d5488e4b8ae96596627f52dc41dcd8786422da5bdfaba21acd747382aeb055eb1a980
zd9c41a8d679dcaac60076844560d7df5c1288e43b10c2ebcf086f25b822416ac085bd92a03a356
zbd332570a4c613b795fd79cabe3093568adead46a0df962c0c6e8dacd59c97ce25fd59c0c4176d
z6ba0183b0c7fd2cd3f72166ad8ea8c78f139a4dd3ed8855fa540d531c4dd0a601df908e66ef3ce
zab94667c650d0468a35643621ad8cc8131e182bbc0ce5f07d9bb018c469eaf32a33bec995fe25a
zd3992e8efc6b93704967c534e2b4fb2a9cb3c6765c24d6cc923f3f7bcfc3eeaa8ec4229e8ed5cc
zc42e05174c780a07ee75e7a4e4406c7aae4c73922d6bbc3fd5123b614c05a07213841abb85cc99
za7f7626c7b0f584058033b58d7509cd095244b14618900c2a2a15d45030ab71c2fbfe5bce28597
z134d14a1b2d71e3de27fa2c20f68b4b6fed528c474657bca5eb0deaf0e0e0bd67d3b2e36674694
z5ba30a5c76b80261f21857b9eef6f7c14d1ef6f2cc24299fbaa49319d2c5f219b27422cfc80761
z3f80191e8e3083139592d3b547cb482587e7d5ed34c0cc7ecbdd4f75afd42144526f3a193f588d
zf9b97d0b1878e8ea54e494ce8690bca9bebd3869e2329781a6ea5048e3cbcff3f85a21024087fc
z8cbe7746c727bdb0305d044dfbaf64c33f7443c84d2b6e89e1bc83949ec7e21ad17d5ea26cf9e4
z853b44fe231eed896125e7e8035b7c7d3caa533eafed16a8d5b32b4658f181bc49bedd2519457b
z1da8057fc5cb8dc9af8dd056d5e8e71bc0d296713be72f23352ad2542cb4acac52c4257a856372
z9f2f1d1fbf762c7360af6deb7d37847355110e9c83bb50ddd06846a8abf7d5521a4f8e52bba109
z4df8520cce3a90caf319aeb79e461f6a7837fe22f4ef3e0d6e7d8a5c60f7aa75cd8a46a77573d4
z4d1fbafbc540fe02f00645da3ab81761e22ecb64b72b5aa54e9a8684c75052be5491c25ea2987b
zf5a5dfdf967b385fa1121dcd57bc6ce6858df02a5d2f9ce51a39fd9cac4b72266c9043a0b00f0e
zbea0f20a258485c2629905476974d5f569478c882e850a4ac64b0749827aae84a2dcff437a262b
z1b1c5f36a806b7e432e73451c3dc937ac4c4d7e8e3c2eb378ef053c315b814b2c099b4c502b7c3
zc593e4ce4a4b4696229555b2f51a9b13795fe97c58fc7c95fabce98f909aacdb5444ef26338ce4
z96d25da1681ebd14db29cb345dde0f6cdc4cfef8a8acc18ae3a7233af620b80337d0f44eed9181
zb56604f3b14d84e755850df709e7e2ced16996e6c8c5c17309f53c24596b3766de707e927cc734
zf5f03b378c8483b9f283ff04dbc5dcf3f3035643f2f004f58f8552a52569a7aaf8bbdbc1cbadc6
za050fcb811802aa1e8db960191aadaaa39e6d87b887cef10e3857db7c884114007a48f3e05b119
zd9923e4ec75c1d4391f4b051a6aa4f91c60854c85867f625c1133c3a821393416b214a2299b54a
zf5b95e1a325c474747aec3b08527937fbf0a9e97aa1aa132d710750ed04d6b4b114d58292c0239
z787e3e9a279dcbad8877748a47754d27320bfcd528d580ef539f3cdd8ba015130541701db69556
z4909f593eb63ad47d3dc5f1f67145345d996118e6e2cede8a5ede6466c35fa4db7c2ce8bcae31e
ze72ba3d5c23a17417aa19d0c7c833422ed8fa3a40a64c56d28a06966b1969fd002513b6a91ab5c
zaccd3fe0f9dadf15cef00c8e043eac384b1b7317dba8a42b37fe75c5e10bbf88a3f91fd6907d16
z1ea8251528584c11c6abbf1bf339db9c8772a8b046ecfea6c64f5b191b283b670792e70a9ce3fb
z3b6bbcc3bff049bb20d694f3d373338fec483b27d1151b0e356bf952e493589c620384a8fbe99a
za432c358a4457bd8dd31065c23943d14e0a8542cac239587bd21d0fdf40468a1e4a014a6b9b8f4
z16c96f4d98249755ef92eedb1cba8d94826ceca01bf788175fca3b95b6fd66a399dc7ebf42ed39
z544d505e96eba982adda1ec480ca6d7cd6c497e197701013f06c51713bd5857c6a0f3e24227652
z492a4f832e2f208e155399ade5929b97792a8e953bb952acf500cbf8b0167ed5573714c7137dbb
z03efda036c14b9c277941e6b76c3f2949d6338878868c81e5f2ae4be1e8987719b95886337895a
zab41daccd8a2103eb39626574e0e7ab70c4b3601ac579795063b3caceb01b0b6d91d61e8c5452b
z0e2e9f323d6c8cb0e97b3e1593f1473f686157d147184fcb563c7c6a41d0907dec706f3621921c
z05c3882ec3b2c87f495237bede8c8119c63ab09c154a3f8c057a3a26b2fc8bd471d083f12831ef
z31a79db55fd936b667e90fa0d4fb23da3e0b79975e2210cdee6155efb267523d08688ae0b91745
z900e20dd369074e91549035a9e30d4b699dfc56820302815dc9c7bafc710cf0f7c11f34788f7e9
z0e48839c3aeb01f194b83f0d9ac44c6c4b1e420b946e7615bb786233bc5fb925f6cd056c3c1d7f
z55c3e64ec9eb2a4fa88e5e7232501471535ec015fb78fd0987ad91425e50ae61ba70964dd010ab
z62fb7081e9cbb9911d14febf4bd100700947542cf71e2c58364dab9fc90ef21ec3d2f5b1e8c380
z727aad1197fa05eb0c406c670c5443658db9524f3829d6d65f8688fb0e02788ddd344aadc97de4
z639c5a192f35d54b2fab62ce4d457e7a591f9e64771cb1109a4c34d7b201d88bded81690185e06
z63811251d61b3a291704e72a916092facf31cc4e451b607d3fe8f0e1a60a7a08012d2799cdc6f9
z6f1c338bfde94f7d006f2d691a020149395540353dd545c836cc3688c87ec7e1418ae0e7ee159a
z28e513c496ca9ee14958645d44638772c58e153a808d46a61ab5339ddecb2d9c3422f9102ab1f1
z7c87a70278646ffa08a706ed8a2c61e657b9a3a0454f6840fa179f98ff2fad69121c2039b6e3dc
z1acc480461e9710853dff20016047a601e0e57e6851d4c9d0e0c4a224d801857c7c3f372da2ee4
zd447cff5b84440f4d20278a0151c6cba8f7e5b432550843615cdfe267ea5d8c42862bf353de840
z033125030e91524b32efc83b53f0e2718a078b73e4722bc21539e3f790f206ac701989e17e7ad0
zdb5f0af9ceb012d1e2de0376794d38dfe357072416446e52933ff6c3e82f1051efe684d7af8df4
z0fb0ffcb5e0b5580839b5b653c1258c32128f0183dc9f104860fe56f1328c357f21fae880ed48f
zfb4e62f41530dad10ad94254dd9e63f7534e10961f2e51a70ff7bf6209848c0e748a2b56cf302a
zb08c75bba4d01b91bcfb6266e150012a2d72903b3ecf401cfd205ffe6827fe33dca16c8d18a7ff
za8fe91b777c433ae05261cdc0210ea54e9acf572899764a15616c57c8ab5132534080ce3b16cf0
zcd58d8b093890a87ad77a4cdf6b43503edf25c7860fc6c9f731cfda25d6a01188f918ffe4a6a48
z99b9c954a9397ed9adae3fec9f77eee96c6ef101427673633340e4c484f792de09b19dbb547b30
z4f8326edb820d46b80694e1704ee2ffc632af80a540b8b9f4c408a35d068626ba4dc23b997b126
za78a3770551118282e5023fe333d8b935871ea836b99a4d1df3c2f732a49267903162e48c48cfd
z7ec5001b13a3912b6904ee4fabbef2d83f8fe916bf256a1556dbb65110382c53f453858c7447f4
za71ad7623283a9ca22a47fcbdb5712d5cdb8bc1da598d36585dc026e8032c02fd00e0be6658a1d
ze2ea84037113fff6b648579ebd49a2a72b2bb80b550534d59703644f7d31af161da37876557045
zcb1689b627c016c2c011f950ee0ca573ed84755547eb8dcda8439d62a25da1a45c44b3c68d6d47
zc8040965cc59ef121eecbc4b08f98bcf50e3a12467414a4a87705c94d189de6a44e0676664c467
zd66497a84d287b6e4ceb14a3e1dfc2dda3ff88b8d99e174c0c1710adbe49658b5f4227265dffe9
z1374f12d01c03c1b229e3262e0039ff2cdeb59d3c63dd57652ab342155edd63de22265f839a3a8
z38d08efe60b3eaa8c3433d94098df1ea617fadfaa66c51cfeb724c82657598931d92eb906c7a88
z5aa47fd92eb16586cab5800fb060c9d653dfb1526dea917d5b6fd45277c4e524c8754b85f430c6
z79cccf4eca78eca53771d2695cc1e7904ad4c75216428dc49919e2e255aada1987b26de66a7c2e
zb191267a8686514dc0b7d1903670d4f3e7c0598065def4596f75b3765217047ba49bf9ee6f7b17
zdb1359483951f3726f1de55445a0621c1d8923c51f7d0d0165738d2667935b6723b237dc1d93c6
z1884fcacadad740b1c3cdd6687d43e7f31672128caad12975909eb9c2cf9bda16113adce54c67d
ze12c62a09338aa321afccedc4613d6fa0e966d1898e440fe12855c858ba65f4828dc3ca7cc7f25
zb8a17859e65fd994987e0b953b209334b3158fbf7bc28df12de80b7d798cb2455ec5d9c35774c2
za8e875577af554c60e830ee6fa60452c13a57887234cd308902857d34e844157fb7d913441340e
z0c4c19339e76a82f2fe8acd22c6ca937b4c49f031483afc2878d3f66997e3e912d1571776cca80
zd525bdaf8ab234e9bbf3cea79761960ae4d266e94df530bc0084d763b16f379556744fcec27b37
za8cc95542d1b3a4fa99fe93fa226b989c3151b2ba00399f5942f15971f3dd3d8113de0708d4ae4
z5adb356bfe43203eff509919fefe5d3d910628c0ea2604fb568de8405bbd617af7c33306775a8d
z969dac73eb94ad8f6da3ec6e062f3e132a31ebc35765c88a1531a447dc0ea202b1f99be4b1b1fe
zb7d7faa8a57ed40adbdb90e4892dbb2baa202a96813957a70cc4b7e77b78e9f48aad56db4cd44a
zf3314254b02c0e10728b82819fd46f8854b0cc6f5c0bed0a2f815fab4e4b46e59918547f2fb5b2
z23875ccded98180c349f9e440d5407734cab2552293aad654f3d74f7eaa714cda18a01d00247d5
z88be1a8a43db7163300a82a050313a88354e66c8351184349e160cbbced554cd2ede4bf33034dd
z43b4a81bf936fd578d413c5c9279ebe6a62690c92f01e26e2e0b4277604a9071b7c1d7e6a410e1
ze2d316ad7589aa142cedd5a103dc9912e320522d3ec4cb7c7ac0814e6a8dca758f6718d3b09de2
z0a843c61f4809aa8cf92a41e1fdfcf38f5fad77452c27bd999a4bb3f2e0aca540d63c70f8b9b4c
zc57d2426b2a809e509e92c209d5c5b612ed96bdf1a15fbecc6d0367cb11a27080978895cb1bda9
zbc2f9cdab580bd0ad2320f3c0c73f821f990139fd6194be4e234de1ae9e30d74dec871594ff802
z975261a56ef7ed35937667b08d0c2720635295643193ba1ebb079ed3c7c1bc18237e3e343f7f63
z854602aefcb7487bad9e0c476fc603f69f7518008bc5972f0c9668538d4fd656bf487efcb87ccd
zfcb2a7bf6b8799c49749bcadc88c446626f589aa391abd73367f4d845b950d4bf8507101610652
za7998eec9edcdbcf8429f1be91e6510eb8f1719a33077c9a40a0030a79fd8c269ca9542b719200
z546b5fd0b53210ed8e29bd82f63a2c100e1f33fe10cee0ce7c821d1b80f1f40726d99195128f3a
zf8ecc716f2ec922d30130f5e66d62088312934fb9bd4b16731182055621b0eae995c4a16d62408
zacb301ee0a00bd670f7e122b12d3489f1aefd4326685d5e17a78feec516e3d8f0680997e8bf8b1
ze7236a102d0dd107ea21a098c0d419b5c03a3a6971751ec1d17ecc49d0c8ad155fb0f173d28b40
z4df6a7d5bedeb07aba3bc12766ff096002e72b555f4682315e5f913b31911bf1f1b43f8e492755
z0afa9ce66f150926299f4676ec6331511a4918ce00c7109d8b41a5cfcb20e3efc7510f7401ebcf
zcee96f733361106cd5806714b16c29bcd8dbda25d4d181a35eaba8d3bfa1c23c0bdc5fdc77a457
z74e0e550b46a06c57a43d591ed52c37e3ab8ace94061420994d6b873560544f5af0180bead8836
zf7a05522cb7d6334ac3f3a46a12b027d24236122563d416ebef4030eff83c863579109a2a2bd89
zfac8a2c1ed8a2f9cb6f3b0c5d5fef85b0d3c3200408bd6b529ff098a6dd03d86fd2bce42da6944
z68fb47af44dcaf62eaf70f687f6a31fa4a7e87c65d64645363abda95ef62601c64d9e274fdd887
zf8ef9298974ad1eccbb2187321b71a83f6f5dad366621306a2eadda19e2fe00389384b48cbe4be
z560fd97fa8532a28a3039e398488184cc0b8b9fd2a77911e7f11a63ced881210979ddfd80b9e1f
za36da86ebd2aca8c661a0e83f5ab20798d6b25f5573eed402dafaa2b26d15b76d7780539fc200e
zfc20dbf4df220b839e95d3a95029e60ca4a3cec124228ad851241e9f08fd6daa881883ac8347ee
z6016adef3acd728684def0549a953d916aafb37d29d9f7d00b318e01cd02d10aa82a9ab85e341a
zd1abbe31830749318f8f8d5a0306cdcbe4a215967d8ca75b8749dff01792b79a9617c43f9f8c46
z95ce6d56f673960c1136eb9aed95e6f4ff2aa3c4962436c9daa6e3e2428f43717533a2c010fbc3
zd2e365ff9c51bc53b757ed64fede5e83a79df9f2aea39e7a983f9139cb57e70044a5502d2c838e
z4601736226ec2c1075235ee9d315269a16e4263ace4699bd36fd8974566d25ff029090ff63373b
z99c6695728dc6f4a6aaad0c7246acf30ac42ef1e6ce2230d302f2ccfeef48514eb66068d057943
z8468b8a0c894967385e29b6f618e5dff0684e7814815c0c206693a357e04ed0b5a866ccc9df1e0
z31c86881effc588caa20d1290dbea7bb50e001f42a4c12a7f86ff45e88cd0f333ee886d99d1f0a
z433044c3542a70d90e9bfcfd909bb5f51305c74e5536c95c860013f780d8359bf9f27dc0dad97d
zc9956a55f0b824868f554162802b1a39feef83ff158471e72a5f9675aea080e90ffe4f9c3ee14a
z85d12cd6631f0b22f3700d7336dff96bf650c4094c85601e782f9c668598fcacd08db9612759c1
z3c384a5f32740ed439d48d3d35f144fe8cf946387860ca7a5f185ded62ec74ccd7615635553ccf
z825b574dc3b3f2dc87eff0c4118d474d302736da45c3a43297ef169ff50627ae832c6b53809622
z7de84f555d5a81ff4eb9b39e6e17e149dfb6693a92e52397c909e7333500fea921579c7cba3c8a
zd09ba5b8e520716cda278fa7aa015da5032e29816ead3653d4bda38d745ab9c69da277e094c845
z8d0c530047c927a24adb124798e37b3341732c92d83648c3b1869d18d8973377728315277385d6
zff84b393be5378ab87c84ab5763c4563f0fcc63e76ad028fd9b5e36e52404bda5b8085d5397ad6
z0ae85bd573bdcefca09b6f5a483bbe860127a54b645f0a40d05935637d285f35f317c67e4d6753
z5858740a8c9d0a5b019220c4b2ff9d1685bc9d99febe9dcb87ef9acf6f6279ecd945beff0180f7
z65f469318a7e2c103b7d85137e7acebb37f3fb8f4c0a5b511a9b49f91b2991b45f6bed7cd0e5e4
z9a9e66202bf0ed45c9e53e86da27bfb4d79b812891c5fae0b46f1d7d5c2aaea27a8afe24abf88f
z7f2b0b95b3071f7a07227b5bcbe8bda31c69e5a8814f49a2311b5051133b754be3eda9eafbf2a6
z33b07ed8e796f703f1af26ff221336aca057ffea1a844260d3fb99bc651ba7454c0ec12551d539
ze1a127c51beb359aa7cf00b1b1004fca5a8463ca8b894cafd840136f56baf3f27bd43a4deed239
zd166b0fd3cda77ad580d8a697b2e6dcfe528bf1274625e16c71dcecb5d5e988bd4f08bbeda5526
z43f7bc9036476dc274cc92d6bee70c51f2a603a0c2064e545960b8d9b01d6adface5144190b734
za66abe9fafce8d29dd8a888b074d788438008e4a183e7e92f50c07093a9f40c1ebf06167e0709f
z3bcd486aee3e2ee3135df2bef5bdfea46b568fca5c47e671596e9a2a16e3b9fbc3cf55af19c768
zadefcaf2c89b81af16719464de02a763cc6a6c530e6e0d2f27765d8e2081aca008691950b3ef9e
z1391c92a2f22009ddc3bd048941dd872ca2199ca6e6a155fc796d0ee8de16a8199e75d479c8ef2
zd30adf88509a786a277daa5f70068847c939e918cd0841d41d58a6b1b83fa221b0b409a8e48f56
ze346425b102e3a290e63a739d220f98fa6e3d661978908b870393ce60e6180984c683b12eafc5b
z547673ae0604e905536827c548ad9c7bf71bad579ce8813de31f767c1c252157f468ba9c47d47c
z0946b5c06a01307d585e0d8c54634aa47ee836c6dbbb35e66e1fb3ca389490c9d235f2d16d654e
zefd560a10f99b0980993d327a06f86ad6b8ee273c2bdbaa699c8959802f1ec36f37b26847ea054
z80b4e183818e66be9675dcfdcabcaa0e8ef13564fd45f122ebbef6563b02e52cf8122ac5bd63c3
z1897372ee59000574f758b2a5091d0195166b3956e576f6ee2f39bc7addd4e503658e965fc8463
z0655e7c8049fa884ca92d279d5dc0495487f3f94542492224aa1dfa8af3365ed0aac51e2ae817c
z852941375ff97d6004c201941edfe31ac0d52ec1e967554b09f84fd568d5e17a7523dd3f064c87
z429d371de2f8a20d628606aedc77677ede245a1e050df07b5cbdf52e0518bd9038c34c7370c2a2
z6426df04af253267ffee56ed6b4d7e47a3ea18907f0f8f73583ae34ca7f9640c77c11d9361acc9
zeda42ec71f449b6b83ff877133fea3b9ccb567a996ea96c57a552171e2253ccb37c9355869c96e
z6e87a80fa2c3cf6c5335d6762edf5fc2a074f2ffae489db69e96c5209301474e41476d41093bd0
z65d1a0fe6c3015cf5ed737a07aabab61253a8054494b7baea78c8e01aa54ad8435862105e4fa5c
z803de1a69fe9193669f02773ac9dd42e7dfe00a027a51f9c44dea597f8155c2899e956cd0a6da6
z7bfdc0f8bd2a330dfcdd598ac19a04e1e3faa10d3888ad29184c2b6b6f717bd02afe4ed5bba480
z47cb30ba93b523f9d21360b60acfbb21a3f9002b45738374d2e98d8773d66ec369bf9641374845
z845964f243f01ff5ac32de266e1238ea6d1ce65b252546df48123b29a0e156f4cd10b09d64ca1c
z79aa05a580af08046595016b8b6fd141378325dcc7f2d059009da64a290614ed85d2c12beacc1a
zf32e8b6e5f4a616d5054ffdbd3b831c1f554ba02040a4d3d2b68d77e9ffc6591492e42829bd2b0
z7d1817dde3c4fc61fb3568d61a934bcba39f9a05a4b11bc9b968119c93d3654c1ae21838f85ab0
zbdcdc8e0cbae782690d4be7cffec26544172932fb9d90c8b4c23474c665f8adc838607ee753bc1
zce207eb94556dda13d5ecedc3ca7d0b073f5e5fb956c7b0a40996e27956040e238fbc29b858d0a
z0b1434c61013569ff28259ce5430e7c221560e78c8144860aa6e301b6803871f4f5a078b677fd3
zad7925e36829553540f930650216bb9e69aa6ad06fc36e6074b2c8aece24fea77d5693e6b6395c
z0e3136c74e060a5ecc4f7f1b973c121ecc907d58546b5778896c3341ff1f672db3ac5faa6bc329
z462498e15e823ffe411114bca09d4ae1e1496a5a45231d126b1d1400b0b28f8cb16bf39c3494ea
z56430a50be4915d6e601d0f93dad3173ef5d25234fe66e67733ece70d8d18822eb31d4289fc115
zbe54038f51beed2f4812dd8e4e4c6759542dbf19e96983e863cc89d669371d513d51e60e6835b7
zb734367f937e2fe01cfa51e9a18a2697d6b885eb64332951921c136942db4ef7b0509d35dccd17
ze1708077dfe76972094d2836f5a000879ab127a3939280e1cf9a1be938ee3b5da4ce4081f97203
zbf23be7171bebc489449309e50341a331667f099e39bd091648e4b7f37e3b081e19580e1b76387
z5233439871f44c73eff1d131ca56433d42ed01a8f22227a1838e9d59ce3a532f9e09deab396d2e
z6dac742c8e1368274fb476a732c0c151e1d4448abdaa309183a186756f0635edda22cee73a8e09
z95faa9b50484cfd16ffd17db39bffec43482868ccac7d24066eae272b3de0b9337f69350e0fd03
zb617bb5ba7db4415d8883a387e46b0f05566a2e4cadf6549e01434b4a3d5c486270c1f698be4b6
z4c6157c5b7b62f4a8f6bda2e1a643f2c06becdb70d80c9e4c27450cd34953ab464d836fa646abc
z85467bb8a618335602cf2fc9ac320cc42d341ccfc914fde070a3a8012b1ff6ac0ecc5dd24d4072
z8f4f4f7ee7eba9c267cdb7b50a50b3033c71c3214be1f10c4f9b88077dc0c5bc44ce4e93d23b4c
z1539e8424ab3081ae5e776a9b6533ed7f9e161f36800e873e2142ea7bc2df8263c31572b19aba3
zdfa8ae78d2052129b21fff0319587d5ae347751f2fd1269d61837b3d2d6f59f867d5d913c2e225
z6a86bcc0dfc173bd9def291161db308feacd00fa30ff05a5b69223f6860b6eea5b4bd5a82baf6d
z0f6826fe45aa956879c86ef79a1378bfde2f0bd32537c12ebe592e699216d84b5d0d259d78f63b
z4df8b94d3a4062821dfa65132e23bf99b9b16460f054d7dfa40840fb288d74f60272a6a849de98
z7c9f750d267fe115d67e7a0c64f9c797a2236c18d430fc925f753fcae7cb95d6911bc942d9ed0d
zdb46b2f48c8f1bad547d43825a671db32a3cce074508e8aac61618bc585abce7bd37437bc4b75b
zbe382f4163f2d33e4fb57e1e46720cd0973e74fd2be6d12776df4748a0a1fe3b8dc99da6efcbc6
z061a5e4651b6e398c5a6122f4b16e7d5a930689e99524e1b417cf854640ecb528465937e9e7f3b
z7c2c1a1effc5928ebc3bff1bfb1a828863d2e47ac4d5dbebcb1b6d95d85a93983e6d5b2c18f75d
z90d647d6d26cd880aa14b255923d25117fd50eb7ea03c97e62483dce6b8a78d2b9d3360e8f4245
zab5ea52f9e51615ad88f1628e77cd8ea3e389a8d51e72c45a85611d40653861b5943ec76115535
z639a5a801d79036160680ac98c197a427eb4b0439979d7b5d510ab874b05ee5b704f2d1b688174
z88a0469e51957a770005802950647b93e6bb4a340041a46459c31392a313375f52dc649ae15b44
z7eeb07977dbe2fcfcbb3e0664b413a1c82a8e5cf04d5bf696c9e79826cdebc2dce2558804e2c55
zf5680cd597c17ba3bc1bd08556b43911e96c4facf2296a76d993ead29bc5f39efe89ab009f1689
z82af2744608fbd2cfca2c125e778205da460d755d6d6fea42fc9347eaa1488f031c55175e86907
z64ede876e3fb9fbeda9f7608e35313639010aa3448e7497fad6d2fc11ab65454e3c5fa4055fe5f
z5ee78902f51c71e00bd8b9fb023b340a55f421dee9c343f6461925769704bb2c89d7f826499a37
ze98239f2bb96faec4b888f76b4ecaf2dd1cdac705549d89d02db03f8c8872952a429f28a6a5180
z6b90b31c831393b23ccfc05d4de05fee7b3959a3ed10051030540b6e73f880c159246cc67d9c35
zb49b866625cd159bd4c1737fe4119f20c3dfcc5be3b0e958f083e704ea226d76f7b8627624d57e
z10b74603f929230bc3f1e8fde00af57b489604bc9f098acf49c8574df21f7c9912c49e028978f1
zb6f6950fb1f72d8f4fd1e1608569b130e8c69c32376873880617add7ca874a8510f0853e8327e8
z25fac2faef04a747f801bc88a5d3c86750ccf0c851f8d5a9a6cecf7d035d6f43683a198a817506
zf1d85f43b8188e9697d1f601e2ff4f76def52d82ed2b4315a53500599e7927132b17dd9c4ac2f7
z4cebe37773c295b1340cb8d45cce1941dd1b02f451bbcbed73e63457b9fbe41eebf5e393d6f185
z1e287619a5cc29bedc0975c1dd27e881112b2b9ac535251eebc48917d87ef5b5a7ecf2d718edc6
z63e096a7bd0119d25f1f9d4a7bc15639047b714612c7b21689443f81e81dc04a9df33f9abd2e4d
z6e2955fdc9174ff9cd7a2217d3d76d177093c15f57273ac52e9d5a35f193fb00be88f5cfbdbf18
z5d2105a193b1b6e8a9de044e810c4f42e3e4a82e17c050a320721fbd55442c718f631ac47b9b6f
z4107495e8d501a8172ee07f948509450363f916ade790911f9d4c4e9c9fcadb70f46d7a24be9db
za466cb8fce35e638af571e28bd1e32b2a44437786656052e260b0c6b1cc68152d3828823e027df
z34a27946a05d9d779fec76187b76c66f79aff39c4d00bc49f730a7fe42633a936fcb9781e6ec5c
z3d45982986b230c3d7ffddbd6a2d4d72ef98e17781bcd3852c677df66d605ff91fa4bc713b7aae
zc0ffbaca7a8b4c59f2da876a2058443cf562addc80ee208de1c699d7f38a6520904a7103a1aadf
z78731760e6f924da3659821216f6d1bcaa63f666c80b4b2327fdfd75c355ffd4df35e1b47a451a
z642e3e6a583c63dda8f7541a3cfea53f55f6ac1d73d2964f73f183dfc98bf126f29c724613b3f4
z34439e3156980871309ce870a622d799ad9149208222c0f19900b54e983a0c746e2bc09e51ede0
zf1dd040c26c0ffe6e6c2d861b11ec92d3d0940fa8866696bca45cf7cc7ffa7a123253ede42f1f3
zf0a88d0b97f49520bf222d64b2f50fa98c78e1e696df123dcae06360beaf1ccab59fea925eb43f
z2e9752ad7ee1085d070a9b949757edbde54722aa91affbf828903d8630f64eda36e2d2aeeec4f8
z323b595970d20f6d4077471bd9c45ced0505bf4d84e57e32af04d163dda71b069c33c5413396d1
z58624aad264ee9c2cdfbea48c5d04c75d60bebd2760f0910949ed50758b867d0654c567235b161
z55a8f67e9c0f44e099ce8b410688b066a8b6a9a81143026dc8ec3109c0bb8bada0d7942de075f3
z1d39eaf274b5f731a745a991c07999436409ac9f6940cd73398ef30bd0de0508b4701ab78e1ecd
z3def3192a0687d1fd2cafae3a02963ed083f9a22eead8c67de9a195f440f475f0fa7353737ec46
z190c682de52ee0620f8ac65c95b0789110a29e737a83562a9c5d2d90f2f01fa4e9209d38167b6e
za06212dd72bbc7c0f86fad0314477b148d30668f1b6dc4b6c768ade508b969b0119d1b57bced1d
zd2dcaf24b71c21904fa780c48fdce5662b08b52365e09dff4a1b68954ef1cfd891ddac48eda094
z888610fc56fee9e434eccdab5767e6dddc08ee85d294b9f8bc95bd9ee8a005011fba06df3bf5db
z56ef041b2f4ed14027d8cd1e5fa06f191d7d9a34111eb6a9f28b7603efede9d5766128b3aa18a8
ze04683adcf18a622369fa12a6d3bd8c853769f13081b31717463b37cff2e4e8a726c50392ffed8
z0b2f5bdedf7bd440ccf76008b384cf5b96546f6c2ec983a1bf4e77dff832916e20dd9e5e9a1452
z3fb91ccb86a9296c2bd39e0ffb04b000dce74f38ccbd63d85fb1487d9c1bfcf63e667f960cea87
za15aa95731111e2d19c035cf77fd03bb34cca6cc4e3fce30e84149268ad672d1dcc2cfbccec8e0
zbe2671dd9b7fa1e9cfa260915ca9a072c92fea80f8e425d059a098e0295604d05310ec8ada98c2
za487992e45ffe4880472db6228237fe2aaabaa9fcb6f64077e3d88c9eed9770a68725e9061a4d1
z9d10aaa93f60a334abac49d32f93c0ca522a4e6737989c89bace5dcecb573652e7fc37b173715f
z3ba0484eec4709323b6a6e6d83a8fc4b19f264e19cb6d649923a2542216f6e872da3e3b3409800
z03ea45496e493698af465182f19a73514d19f20f1044602d64d45fd671ec2743e96e03e2c5f8e7
zb575b3f6c8384bf1b8e1f54dcababfa488846a2d005865d19578c2056e74fd0e7f92fd1cab1c85
z185514199a6a9b2c03e2e16950c8196702bf145d80a086e35563e9f149171966c25b2e1ac3d014
za3e4f5b21183f4cb83d829f31e58a7cd74b744882bdd0342d7a11bca164ccb41a5383d284493cc
z9ffe69d6a911a20a7837b17cd4d701806095ea0820bb50b1e7ae63d2a5633369e7aff207a66f73
z423f13eb2f2f1e376f1d207d2df10ae1822732ae5543cc76061abb3fb850d51943403c7459a6a1
zff14e2d8ee76410529e42076fb3663710798a58c5842bde4bf73a4f4c76c5ccbfcecb00a92c033
z4ddf313d817eb330d0c435753de6aaad19ca2ad0469f017a4fcba9d0dee4c282bf4e2805a44583
z04cfc25c4386d227506d7b6a7c843a18d3c9d9d64c0ebf187075f80e503a0296306759f63b6725
z63ca885a266d410176d4603b02b8c8a54f6c4af362c7b5615005529da7cad7e008bdc84f7ae85d
zf4b4092457d733c41fa85429643fdf9c8e9d90c12841456cb2d8186c486bd428fb8f6cab1697c6
zb51b47837a4cff0db046258d18f9349a251d31b3257b31d64a8ac387b0c4d1d596c44a8142fe22
zc5cbc7a8e392470a34df81ad762664d08474eae0391dcd94dfc7f3c517635b001ebcf881adca1d
z8c42153748c3b979d83df62177394732ad12c64a772475c9f53e61f12dda64feb5c14c6960fb28
zc9f86c147b3c924163cf5c97086e09dbe9e50a7190c3b20a6862ff4418e85aaa83615b9e04c80a
z05880fbd22ee952db9614e63ed53b4979e9a079792aa6e65a81835c6102c59585721f4e7c3bd81
z3b4994ddb4efe8d2f06363af789b413ff229760a2fe9353f2c507ca39448c57aeba33bbaa4f019
z59c24c359bad096cbd36c898b6a4dc4c94bea65ad6e3bdc78b6786da0b7c65ef0c620643ef68c4
z4c058681db7f3930ec91b10d154a9831f909c95eac76561e2b01b96ae2dfb401bb9e437e678da4
z75b204c2371d2f15a6cbb123554d14200273d512dfdfbc13fa7de47e1e5d9845742c6656f358f5
z5418d00101003a3eb13a5c16ee62f0138fa93f72ebbbf7239bd6ba71b9f58ef875dd0ddab5b5b8
z8b8a23261e8ca94209f63c65555ba7234a08f84acf2ca70e5ee6c92063cb96562abc72d60c25d1
zc6a2ddcd459b288118f1e311453b992d9d31a729e92a90db9764745f6d635076811103ae11738d
zf134cafb108cd2a47822db5083261bfa5f70b6c1b2b16f501086726dbcad5f67aa8ddb16b90b3f
z3415657f4b976249fd6765c86907c306685283a69c7b1b73f5987432b34f5261dcb8d6fbfb02aa
zb185defad1edeef15aa05374f700a024fb895e8580698bbcd76c9f094b1f67de910f0c171bf236
z373514fab877754b255809a07ca709f3cd95e1362591346791697b4e4bee37bf5158082f2d9c34
zcb006d83358aec2c9a13d82566f38c8ca1c8015b021ef15c77a9ebf570e4b87c153565877cb809
za274f1f40a160a7a335a480bb8d94442ae1917598575dd24b3a36905a153bfc218a22bc753b09d
z3407a77032b43bc79785a2e14b27e7b1ba50413119323612791d2815011cfcb68c360f353ea4fe
z37c5db77dcb68dc0255b73f56d2b8f5046e61f8b8efbaa639e5c253c566d90a000f4be65bee5fe
zb3c4bc00132b5c60bd7a4e61a1423fb47c949d076804dc7fe87190079c047b964f4348ca977610
z01cb5979fc243a69fd1c2aeb83b1f20606bfbf70e4cbf0a411df700ae296cca04eda0b973992b6
z9a112ce56c08d8079841efc7420695c175b9e1e0d4dafd5a56aeee8d1050a4ff103b7850953bf5
zdcd4a840af22c180a34b34ecda2630625d66ca1feca30450950c9d4a0c8dca20279f4d70e235f0
z82d328076b1786f2db2ecf0cea145144237b27020a4e27da904ece2039fcc52ea7007b72bfb441
zf6750cd7e06c2566c418ee22469aae801d02d87a3462417666b67b461ea22b160fc0dac5acc1a7
z7c02e89034e472fc59f570fb4e16d37648b7568c36da08b9aef6a82bdae838bc157310be19dae6
z36f9fa8012c91ee5f7022c91efc8f4c146c0c1bdd8ae43609c131d2f86c66494f96a4b3f45fdc9
za64a17e829ec7551728212a1cc2b8751e1d79873900b6a008ed3f62c46c5f9622f31ae1528c39c
z956fa823677a98659fea9fb20e650a8431a9994f4730dd06716eb5559b6e46587a407cad35894d
z53fa2ef149732e9d4d8e2ede261f3cd28c68abcbdac536ba3b8acb78b7a29f55922a445ff64bed
z0027b2700ac9f0a5aaee84637070fabb863aa815de49a32dca6e02d79e4c1c2260936ef785e978
z9c2ca76e18045a25478c9a459cd031d5d7b2651d6f03797a262ee8dd5ba2e97378447a4aac6ee4
za78b2fb954701ce55b79d757942c264335a1f8dd2cf00277a02bbcf23a3540e0c4ded0c66865a7
z157c01121fda82ef7daae2442f85c5761eca7342c85de7ea2aff7a3a1cda39fb7a16ec7bcaa5db
z98b0170e53e708d65f5bfce715407a72476d14278e0754159ae288ad6f6c040a1732ebae5bb8a4
zecc1770deaca1070534a0e742a7e62ad0bb82bcdf2bcb3d94c519f74809bdbc482829a892ba16b
zb9b9fd3ac3c9cd4b32dc40d91ad8fef6cdc4230e28b528fee36ad059048e0768d76d9c57d572bb
z936a86810dc956f43155f8bb5811ba56861d911b300538c633116265f36ec6c7814978eeefcec0
z86ce205749cd1abb9447207a01e57e811c5d727f045b74da2dc94450b715d809ffb1189a9c524d
z7eae0183020e13ee0488777ccc37dde265d0b9a55449bee2b832c5ba628b85ce9b4b25ee3e876d
z2adecb46f22c1788f92b74f3aff3b1f5347bbe0b2f7217d0809c32f543f86356aa61150503a62e
z4c35b62357d36cdc79a3944036625267e694cecb20d0820c0fe3161d9781a3a14b446fd2a94db7
zfaa7dca1e8c18179ead6c0dd4ecef541746d57d08326fe5cf9ca5c1f19442d9b41300c5b0bd617
zd682440cbaa047f4bb10341741c00d9193aa8e1ca5062586831fe1d83518ef0c2da1664cc515f1
z02a9365992ab95daecd6da3aff664e7c007225be227b168bffbbd0832fde5bafa4e52669c8a6bf
zfa928af020514bd436f8f49503ae8de40c98c1dda1abc500dc2db65381ab97bf704c73c8e00397
zde1699a2aed48825e27ce43241fdad43c7ee52ea1c340247f95598dca86424e5bd066e6b466e2e
z6d5aa4e36a2a43c56d72de6c0ec612cb8cb8a1adf34285051245df893b9f0acf055521fd11ed5b
zb69f2380c74d06c9b15f55483371722cd1eb3c32fb334744ac0fb52d897b51bf7f5ccf07c24eba
z420539bcd0559f7f501ba8a14b86e0e4f8374e9ad7b4ff1c720b8b2dcc93a42e47f0587f14bfd2
zd4e56f0eee854e92d89308a124a5a9a82c6f556b019837e617f2df13f27eb329f0b77a0d9e274f
zc93e3136fc15f32ae95b0941e0b7e792fb1d6d5580048950408b157cd2ae806931d75365ecbcc7
z9b785d3c78da8eea2206592939017042a1abee58576f7ad62e1d5763fe2d4db6043ee7cd00f465
z88bc3769bd55a97410d055f567c77de5f527d938cc126cef4fd942ede19e7488598eff789539cf
z143aab44995a7c878cb2ff4c77df245575c58fe42acb3a424795594ec493f44401182a79c4eaf1
z87c45b11010c96541d5023ae4eb2544e1bb8110cf51c89593ba8487da53a8ba7a65aa10bd6534e
z7febb960e5d917815e9f1909c122b5c6b07da00a29ad06f9d056945ccc8e12bb99ede75fe3979e
zf34050a0335bb10be6695c3389ed6eb2d1815c85fa52551661b6329bbd34912a78a45ca2183866
zc950d8562343c0275720d88790cf3c046c695edcdc4ab9325964401428ceca88ecb6edfcc47d90
z7d0ea58724dcec8a030cdc8ab2c5ee2ff28a0d37ced009c5007c989089c5e0d94e5638bf8f21e5
ze1110280a052b884c543c21f693fb30ecb634e70e894979ec961bc48e703773e8ba6319a921679
z160bf51e171ec074e8ad891ef55670b9764a08bd859b4296f5a9a4fea43e0af8bc009cedc4cd1b
zf3f81f21650b2cabb49547f1da8591c49bb8d7f3daa834cf444b5cee86a023ceed65c51695e7b8
z1a8ffbc62944f7ff946b10e8b1e87efa6f40a429f4ec8a0ad4a3e01edd1983f5cdeb5dc805e9a3
z1fe22d78ef7a060ef8a8983daa751d95b357967de691bbe8dd0ff6395ba1891132bec04abcd17e
zcffdfb949b21a37ac1408f17db2dd25089b66e02fbe37069629e4ca5883a6144fc846fb2aee6d7
z8e39e1ebb68b66b1f729225a33f100d1752728f68fa36d4e6ad8b86f984fae942e8d3f14098b23
zc66749ef91889b2db99eb2d95b6b52bb40fdbfb79961464ebf22a29312972c4a04dbeb1a8bc119
z4447977f783a77a07c9930c02b9f5504710dff416ff3e0ef927b7f513e62de085dbaaee44fcefe
z3d9a15c3057da7afa85119fbf44bf20932d6f9735dcd63a93aba9b9f6198aa60b3a651fd184b6f
zc3450f9ddf91d2fe3fa1d6aaec6a5a26d478e73b2771890d61cbaba1b5c27e6bf4a65b24c6df3b
z65fe621c8f61500582ce2a30c3ee20f3b6419ba2fef3ae1a25926d0b5e7078f4d73b074051565b
z0fc19cece68ea8c10a0d9d4c16bf3cb676be7690c1f7e5b228729e8a8c4dc56972f88630aff002
z71007f9f24c890f21b77e7c70319a069f1fbf746b44371debd2746dbcfc535f25242e162521332
zeadae26d20339819b26c7ef135986d24e3db549eda9206b981b616c5e2a7ea30266378091a0455
zfad7362217c48a8cf275a5e87d8d41f07a5a4be057958af4d0fee627e9a95123c9c57a6812c249
z66a15c57e84b9bc81072af63e85d6cc13d3a6e386d89cb1f72eab1ad559f160506eb7ac1fd9f14
z425512aa04e56449892b78174b6c283795b6dad393cc1b5f279a6988d2ae8e4125fb5ff68602fe
z511dc8d77543347f0187e90a81902ffaad9f98923bf064925c8602bb28820b5260e62fec7cf032
z7e421c421f56d18e7a3666d31bd0ef5701f48d014fdbc493a0dc11cd66db7898f6158ece81f0b0
z3e3ebe2c444bdea3164788c0b851aea5439e097cd45989c166d3058f721cb961146f1799900178
z793a08bf6494e09cf27f557423fa48e410007c771a5b1740fec82022bf4634f214664e92d625be
z830cf967e852db874492dde3ab330922628c9195e016448365e763968719cee5aae1fa91796d6e
zc87dcc79802e0e68015cb415d01208dce90a24ed6d8a120b4b1b9c96d387a576dd410e82d5a478
z39754824d1b83468b11f03ca3c9d0d6e34ea69dccb63205350e44744a1c2df39d62f2a4cb32192
za9bac6fdccf5f6c4f147672aac46a9362b0ba122e6dbeeefe5fc7b82fee15667d94ad9fbe67ecd
zf6c4b9e59b40f2a41ada3fdf25fca1509ddf5376ccbfb5438834ac65c0706e27d122ceddbc9ee2
zc7d887fc32e55d07e77d42d28a9eea99dbe7a85f6d5634c724be58a9fbacef1a966e4a8a47d18c
zcf1adc037d05403240e0db2a30b850c4d7492e1e061fb4866f4cbc06a268aa3f8f083593d99c1e
z4acce947ccd74ed0fdb13cdf0329b2061ebf95b72f95599de19c33e313879b915b17dc90e1f85b
zf4013d1da1f26c8fc9cc5977c507a69517ab2844993e24793cfdf8129b73ef3ea0be6706a3d89c
z819f8c263f1fb042b10a156b90fd0f5522723c83b1210c4cb76584bb7928b5c1779a0a3b3c68c5
z5c6cbe65130762935d6e77fe6702a9c2017ec81ba36d96f22ae4208c9b9abec070e77aace7eacc
z6603767df17ed7d0085fae9d3d691c8d734ea74fd0f7c00a7f666f975b88cc7bf4504268c42ef3
zb2945d0808b72137f1221350917cb503a6ade68619c6bd6de9c15cdaee3e61b005ca43705e42e8
z7d850041c33c79fa5c809e19093eea920052eb1cfbf615ff3e8e3a964cf29196eca988968f9c09
z2c91a4fbaba768bdd26653ab8058b7380f0fe6cb23ce745ece633c2187819929d11c1bca000f44
zcf6582e47fb624c0a00803ce18a0042b107142bf2f7b4976ab84770e20afa012b439b92f14ff50
zaa504aaea81b64fe58f5c8e31d5565d9752310b294fc33f4826d2006d9d8c3c51ff69aa1f6c305
zf9a0ddaf380467df44202207b53921a08271826f944372324882be024a03bbdbd8d07415a73c42
z3704fe772f88dac3f26d071bb88fb4b19d3cf7bb1297c1f8df58e8d6bd0a461a16d4d072ea8da9
z3360c30cee9cfd0c8b57b4e7eacea53619c5bc138a046c484f4ab1cb6effb5bb8cfc37a2e6be02
zf8668fe3c516cb06d72297cc9a9b6f656a313f4e59c6a540a235770d533c9a81e27439a167d594
z24176bab41b946083653b189d1bc8d25489d404f2685835447c273bab584b233bddb14d8a3fa00
zc62d9fbf7746fa5d1446463b43d13cfe5d7283f5843268962d2ff74310a2ee8548154de80d5cbe
za32e06db56d1075ff5ffbdb93d2b174c99f536c1766a43276af02f80cd0cfcfa870cf8af24d13e
z770656c217638ca9bdbc289741c54fee74fadd2f4361bb3c938525880410792f815b3f1938455e
ze03caae2e6aff0221e77e8636c14359f4d3727ce8e6207ab5459f775d194c1783bd9b2bdcfdd42
z4737b30330482382563c88ebae35a0ae8b8cb87f41e684948428ead578df0b0a8bef5d69a210a2
zd33916efdbca928e16b3422be271405df43ecf0b9b9207551b262ac47f9e3912dc1bd084bbcde8
z4f49f2910efd02c3221099b36a407522137a6b77515eff0ed35a1a6f32b237d4bf699a1e64e6ef
z5ead2887969f801e39c3df0d3b59a7bd5f5c1fe7c772cc956e21fbdf10300eea2b9beeef07e364
z2c63c11a1bc6f7b731d52b198e73ac39aebfca0f4d3718e632e5e7274d934ddb0285cfb954ea53
z7020df7468029c5157c3d5dbb758486311abd336d0c8b44cccb8c711c91f69210eb15664f4ed48
z8ad2c93e2efe42951bc5f3a2db7d426eef3289d089a1610c7135ea7f9d616d85b1e4f4f4bd5add
z1fe28c788f680642344bd87cde8b5c2fbc7addd04bb99cc3bbe2329e4d8fcd72347b16b34472a9
z62be9c7a9cfb3a131807c09cc243cd224c877c62b97569d92a0eeb6990c94e5aab4f9a958aeb9a
z482efa0692466184db36d4899ae2fd30c4ae631a942549952b79c6ddcaa339f23c26c1da148b4a
z3c17f7ccba5fa63cc854bc9cc815bc057a5479a88a09afd3974b97fd2229f37c1e7387539b271e
z21c6fabe75dbb972bbf6d0384b8f6c48ec5704b41acbd469201ac75b9c2420b49aff7715d682b0
zaed39acc9d00304e74bbfed72b8355a7eeaccd003cbf42e497d07b88ec1ec1a6d10675ff205510
z6af1dadea69fa8bc74f87bbe396e0f8ab159333470907cfb0fed634bb85719dc2ba3ecc10c6957
z4b1dde4dbd9f56213ea387a79e437502ee97da6a6bd1d2ea41a8a97210882478252f682633dbc1
z82a4567b06c8112ed1ab61358cb9ca9fbc7658d5e3e913b79a121358dea9310fe1105d8c09f497
zbe165e1414dba90d54f437c6bbfa021b9f8d1583e9d99b7f815b255a68ebb4f27190aee7246337
z28129cf1868d348b1c3e2000f7bf8153f9d4d069b6c1b89102708ad2215302bdd1428fb73b6fa1
z8efd0d9ea2488bcae3a5d18e95a75ccdf910c3149ed0089187cf03ecab1c688a50a69f761d8f4f
z3d8540d4ccf23b671b4a4dbe7b3fde0ac842c3e8b0a92b0c4ccae122ce743b235acd2aa39efaa2
z50aa916742b7b0e146bc9322f355d2f6b8cab0c7c370063e97afb2d0434d9982333ba08942c1e2
zd5dcc661e35e1755e572752aae070d93d9758a07202d713fb41b7515b1ffaf37819571c0c3e552
z38bbfd93d7b25db6da48df699fb067545c6d576ebfa584b69d841f5bb8bbd70bf91c6453b4286b
z91260e83cf4a3640ba4ec8dc9294bf4c71af4d1f92ffcc59153177ebfa0346828eb03d1ea4654e
z3311f64a06962a1a340b0c82d6f5dbd8b5aa16ef6780a367f65ec757207ff854f05564b5c9ed81
za021a7613e588c124a8365c236811d21089a4e24d9d4b6902f7e3b651c9d2a0d72558f3ef0175c
z0dc25da017d6644951fc0a3e4602caea47a47f88d29b3a3d40b1f3b7072a783b4b38af9d9d0193
z770f7d692a6e1e47c13048b4059ce7aca77f4c026f12c50d848ca5c63ee444e8400e113229f971
z27ddcde81e197f688e96a6ab5b1c4d3eb7cc1b997b33929a919fe4986defbaf57dcdad9d8a62f7
z01897b8843808f63d10571f0b8239af5ef2e9c6bb5aca913a5c173d34661f9c4b1f929b8e8a689
z1ff830b17b69158efd0c8884d73cd1944663dfea0f4bf379fbd508430355ff59d5bcd73b3a6fa4
z9e4cd1e7125f44ee220c758fe5929b2306ceb586f81d5d008c27146bcedf23eee59601b8f5654a
zfee6dc5b4d8a0dab11c192c45524796ae2ca194e0c95c537883cfe8ac1acce04429eea39d4c77f
ze88a68c65c1cc43dde2de9aba92d0209ef3a2d061a4564fd6c570fb0a6e572184b9bdff7a362fb
zfd06aed9f7e54d1aed3011c93e848756843697bd60014fdb1eaf5615708e5a88c231cab7615c65
zde0dec9d1f8e9eee4409e1b5731a2c7b50115bba007a2ab2f0b9eddf8da909c154d4e0a8d5043c
z0800e3beb1a88fef7c41a12760ae5121303f5ad919ce91109a50706e4f189b352a673e35468185
z268af691786e7a41a4d3ff2ab02317aba4cb35e7bc0323b03c0087ae4e6135224ea6083cd9b458
z15d89335aec594c2614e53926a930eda51b72ce534a7c2423e52feb8ecd16c06514bc0bb13f07e
z6e3654ec51d05467acd0153ca6d7b1a6aeb4a890590ea8ca3b2bbc323a528d2ca2117919646fc5
ze5779ae8d2a5943a3cedc24c1d77b0fb20dae364fdf6d82e796c8c019604dbbb94ff439c68f0fe
z7aa223890a57b3372c14c60d311e4211ec53e998e6b0c3d8ee0ddd0edc3e23b7d13895af64d288
zdffd64abe40d50b5cee0dd7a8f2ccde61572907da3cacf2aa296e1797b33deb82f871483a429e5
z3eae898f3aeb8f863289c1be118fb6342f3a30bbdefe30c6fa5a27ad73b8ab5c82e63b81e0a159
z47d62bc350fcf0dea556b1f09cbcc8ec02450c276fb6b921077f380d5b14d93f60012497c66b23
zcdf40e7f29e967b660b82d05550c70139c6730707967ea9e143afa81df4377b67146715815e61f
z5a8a7cf0c8555a608aecff810cf17202cf5d0fc0967b6b3304fe721a68da0edef882fabfc7dcab
zc5b2c30f1e1e2141c339db610a0ed998c6bbda805bda21ee2f3dec781a44ffe587cbca71535367
z025b76bd6d298649764b2fac0135034e517bfd7d0f6cce965951abea67d019a2f20e9d05a080a4
z6ef571612012be6d1a8f8c4026bff6be34d851a170cc427e0c7ba298509af82710f252367535d9
z2e28316fbafeb51e0a9664f2efa0af5336cf6822019b463357d8fad3a54bd62c5102039ec3f4f7
z8b0ec6ee5628d7d78b0a5dd79697cca783261c778a1e7e570e889332e75a51d4fcf29d77be5f68
ze4cd29a03d409638ea44c23b77ac7b250e043ef177eaf3ceed2fb78a5a2469d7ef4f923ca0c72b
z56fac56a1b8fe0900c69487a5308064585ec1da15dfa63aa0b1ca656103ca9eaa2179a10deef5c
z06ea8027b3546d154a82398a919f955c5e24293a42bcc3f693edb6257683d23d1118f00e0649c6
z7eb17d93e775d0944cb51bf842b1afd47fcf87ac98e6b3ebe591e897021e25ba969527d3ce56d3
zd0e79066a4a77aeda6c3262eb0146000d672d614e72d79ee4ef89178d5acac5af042c2e439e42f
z2e55d934560fcae7676e30d8655c3c63942767b95c95f832345600916167ab48d98f0c30d7dfc0
z66034618cff151a5baf11a8e11247b425e2b5a5cd3885c79a7596bcabdcf146c6b4e587514394e
z7b65c9b2464323971eda24bfa4164deb184b2b22683c798eb6d1c24e93d5f70eee37e5228b25ab
zc1fad60f992a2bbaa64841d83da90eda688153ffd8f15f1816781f4e2b6c989dd215434410ff3f
z1f360dc524a90f3c9a636f330f350ba6aecfa7824a143af82f2ddad9158a12fa4314fc3f748ffb
z1adc604eff2b7e06f5439e152cc3d6d6e7bce7d180cf55aab160c95516ab5e9b88288bd520b3e5
z7208bbc5c6c475db5aefa489a7d8b20b799316167835d7d2d25712c2dbf8ddc42d92fd150f801c
z37b280fefa9c63128731e2af8e91e6f1034e06481d2911e0aa0e2747d3c07e04ac6efe456e6a17
zbb78b3cdc53e82e2ca6d8af0d6ceb3cea0d59e973e1885d603e9f73231aae13ecd2384b9ccccee
z8bb3b03e18c762ef3a1f4ddaa685c5f7f7c23c980058c1be51262fec5b62023fbf5bda19a5749d
z3b3e3ed1fc2e8f897d70c0877af9a7cff4fffef26ddbaec1255323d33ddf5d27e5a52f249ecdca
z50d3fc554b24f76fb46ef82f4cff0f590849ab8dc190bd519725fd5960d4b4c8168f935fc85519
z3603b43695f4bf3a81096f65d44c1f4a0b31c31eb45d693e73fd43682e28bbdce490a2dc138955
za12de6853dd582f1d2aba42e100aa062545de53aca819f3b681d0f75c1219c1b7fdca4a70c7f0c
z488156cacd9e8b2686a4d48f699624d124356c0b5e5395dbca7c7a933fe7e37ca85fabbb3953eb
ze10870907e39debb6466e09ef48fd0265661b1441f190a97849fac093b5ef17e26e0f24ec35654
z99c51e0964ecd2d3f3fc3199f19308bc87c2b2ef1fe3615e2d8f29a322b906cda685f2980affe6
z7df767af0b97bc9a7b0f01ec87a59e2717a4edfc5be9d4258c82c33d7bb5d3e57e384995b9adc2
z9bf2980d0310494015236d54dc1f112352a57788606afdf26eed57d1cbe1639befbf57a1e4a92c
zd0f13ee5859b59749a2fa37b54541520e583ea4e1c2c50ffcfece05c60d5ebf79c8da3f0fa4bf1
zcfc6eb7b035d69f61cd930a32449b6984ec4ad4bb6d41c0f589d628f111315ca04d68f060c7646
z866f9c23539e678469c7ee1cd45ed259ec25e6c56a2c52adef0cbdde29ecd801aa79c997b97695
z5e97eb24c6986fbc73ed39630ed8f29a3c35c0709b065f6b68783a21f920086f0b3743bde5cf96
z0f796b327ef1f135e290742312704bd68c13d34dcfc6287206c5a0367dddf8d016cb5af67c5a4a
z7a9df73aa81377334610f250529b892e2f26e00526674b3b0482f630bfcad7c17893632366db6d
zc40cf1151a7e64f5c35eb2c2ab5ac0cb60870b6a93f475838a44c2d0903151f4d8c2d0987fe032
zd44aafe86bc01f1e3c7ec4749f7c8e3ff31c1aec8992d7ecf9dc96cfab77b79a443faf8602a985
zc57e60f562d590b604f8e32329cb28f8a1a08050ee4e320f472a91fe672c0c53b31881cdfb8784
z15c94a16d3b1fd0120536c2e18db49d1087e2c289b852f4bad51330815a57001d088a278092b1b
z0069d750bf876931b52d6e7c5e09ac7bfd4b8b0772d4b44351eb8226ec7ddbdf36a26923c276fa
z62094279e3bdd9288b0941283cd874ececc5b7757ffe3e76fb47f64c150a2c14a59461fb82be59
z3aedf6b3975e533cd0f2206bf7e480ce92812da55be2738a0b7a2e27a018bed799288ff149f132
z34df09c8b1087fa4f867f5336a2a674222ab3a22347cfecd689a2676b247faee9d8386e6d192f5
z8ffbae1336e0a30e489018b5fe89d5c268255a0676606f19358295feb02ddf37a77fa9a8eed2ca
zda57363330f09ee012f2692b4f253e35db2b98a6b66c64aaa7ff8063fcaa176f9bbde0361ed276
za96404a21d10b485688e84932689cdb1d4e4165f36a839ca36b3afb5c82cb9bbb3b30c550f319d
z1d406f6b08ca9de06ee29dab71a6a3335dfe6913b9f7aa1ec4be34a6ffd5d49c9075119e1735ef
z84f8f7e006b237b2653a81f394e3e13c295988d57f99bc5bfe4d0df5cf225cc266567b08a81b9e
z78a878f6aafe369d5873115ceeb880ace5a807726e3ef54948656e3be5a1421572a33aef4c9342
zff95b06193c923b7b7ca16437ec335e933b4f0a70d22357caaf25e7f38433fdfb6a6813d3b3027
zc0f5be896b399db13107b45a691361008964864cab0c7cc0af0d208fbc32a642b191da7b3cc890
zc8ad2ccffdb53c15f772aac113a44a008b17a22f733dd0b481847a71e77f00fbbb5dc4eb39b9fb
ze7d6ff4e06eee4eb64becc0e632a9a387e1a27ba4ffb4ee9c0ba487fcc9482f926fc7173ae61e0
z5468ecd072c026994ef296a4d14f5ad5dea76008dce9ca3dca3979fb71ddf6ebcab959e83aa88c
z26cc5e99f24c2324fca64a26dfe7251cd3ae02c6a946b197dd626904b6d80e8141c06596827b2a
z7923e11264eefdce1998cc92a4bd8d0a1099527a694dd9a753904f09e3b5e32a8ac2e9ef06d0cf
z862dc83e33a5fa37ad773a77b145dc37da7fbcb93656037cc72d30cdadfdc02c1034362a98c477
z39ab3ae6a2949fb2aadffaeb779f2b38e5572d0e8e4b4cd52afe3fdf61cfe161ac9d8dd6a434df
z2c9a5fd7df6d082c7db4d915ec7f155105e7cd554a0e216e1a90f9e88906dd8bfe64931dd60ba7
z81152407bf3e00e70ee1bb2d1d5484a5b8fcbe340e621c550d5612cfe4e90067656698ce39b20c
za3dc6a2bc6c29686d1581b741a2298f5df6d418e23992fe04960ca1f8d332da33192af88e657bb
z593c91ea18ce39deced8178b7a8ddefa6b19fb8e737b89b5b5eabdb74f5a6e181954cd382324f9
zd418fe3e7296b4e9922db019347571150ffe39afb449cefb708966a343d6f0a7090f3f29548866
z1dd687b95fa298090e87c4f3ac7477562377d44b61570f7e4c550792042674d420f2dd182f6aac
z25c132e997259d61817716a3f14f6047e51af3682c05ada0d3a53da53ef74901d65dea5d5c3955
zfca3c08bbac6750f36674e521e873914e80034d9e28d6f1c771d472a5c2e62afa83b3e826e14ed
zf1e90bc6e10425667d6d6065affe203987c08d3b386960319c716e1d1eb5c1c050c0979d1c8cb9
z7aa80eab66bed6ee24d3cd84b1650b7baac5892d60c9e44babbfc7a489cfadfff68c0dc2b90cb8
z622d10cd71f9b963bcf12d6fc46e093c5b488f625babc4df78570e8a12cee2620f8dff1cebbb8e
z0569e8619404ccba1b99dd44e9ac29521900aa7e4f33e8e369d70f56c522c7b732cbff3cae4e04
z6dcdf83f3c2e268f8995bee91e88443d358a143f0042ef2ce5aec3c4dc121a1bbe90c827ee39a5
z87cb4c7f7326ee78cc256b2b59745ad5c3427b9e8875fa93518f7fcfcfcac4cf07e35f5cc3ad4a
z2acb35123e918f0b4987534653528560fbe2b46584542401e36eea522e499b4e5f715e6cbf8941
zdadd38e450ac32c08af10bb5c1b6d6b94791ebc2f1ee2faf1c69260d772bfaf0d75b2703d05d06
zfb3330a7f535cc92deb28c7407b0091423fbc80bc8bc295f7e3758838f54902b9a2bd6b8c083df
zc6a0ca0a16a21c87ca7854d50c289d4120186e279539b05aa921bc4b29a59ba7689008560eab1e
zbffa9f05ed734aba2d68986206e58186e2ed1d124434c042f7c03f9ea0e7ba75a0877786ff0819
z570e2b78ad9a670e872af56ae87970f56050beb61e71f6d58a8eb317aabd4b995cb16dc075ed38
zf93ed4361dd8bb550d4597d54706b2ba43cdbc71fed38a30d311b9d6c5ecad26f2345217fa9877
zaa0155f348d358b405208e168dc7f1ab05e19672062c0749eb9f5424901dba28e0fa9eb6cafa04
za46808244f2a838eb837c50e35b2095714c052d2133dc6fd24b74983d22cf3f413e2ff8e8a9b5f
z675b9cd61e05a613b95734ef90546e689cdbbd34246c3e5c9af5ec369e9d2f38bf92a2a5a74da6
z7169018a07f26ff19b7a2b9f57f57eceac32a3e8119e08c0497709877cd125b3508e1709421421
zc035e868fe18a729bcc120dfd8b91db10e37c0c0864f2d3c34186fb6df34766e2f6779f9f40a0c
z849cf0bb5be782f07f85fb372f5456a384adb8235a038ac106e94befbc2e4d72f4b9dc4a7c888e
z8452c4c133a746772866c798ecfdd05192319a28566572e801bba1bb55acb614d817949513b2be
z6a7e6098795ff94900940c9ef0c07853b6f1c02c67a494a4e67c34b4d8834b4d0dfcf6294af715
zfd3b6dabc44b4997c9df01b993b8f8cb14f3aaa12bd16995fea8482f58697e81686bbbd7d6af82
zbd96709c9b91984399954cce545a50722d8e25120a83559dd16aefb3caf5764a7c8e54d40d3e1a
zfa52298e9f9884924807acd6e19f6dcae49f797c22107caeff2a3635b70fc4fee44e81e86bc849
z8384d3c4d11d4a2adeeacdf13124e7d7f82f36d673e4daa68bd5f243a6bd3b374e70bcc7e4e486
z8f58caab2aef99514e6ef95f4bd3fa08bb2c7a345cddd8b831c166fc9956f27cc07bad1fa9a0b5
z4c57545bc6a6abeebb6eb0377194ef6b96310e2bceb17693c5c3dc81aea910a366693155be9386
zcc4e0cc5f7bd974082bc3350b7d1b625a0c19ed3264054d58235d147a53e24155fdb426c9955e6
z98bddb24cc6050ed5b701d7cb55d32cad037ae3768e8d4b239cad63e392e9fbcd459f1c6bfd68e
za99cbc2928f87650aaf8e55b846ec68e068154bb5f828036c9b3cf7bc2f2e4470586f028494dbc
z817b15da941cebdd88e3e53c7b62c0e88cc303036a71ab1ac62854d0f025dcf088dfa668eb280b
z79b85ce64164cd692b8e43697ca2c1ef0512aee093e88770a44a602765044618dc31f0a6d6856b
zbbfd6f0958cba7a3cb95daf8599932e57f0a3f7dd87dc0fa4a34798e477cb05e83bff9fb666f04
z7b946c1fafc8db7fc7d752f11f20877d70f38641d79d9579e0a6b2c21c9cec233176d46a0d9c91
z4b3f2fe978909cc3b314febc116977e7813972d2ff19eef639aadfab026ef92c157b020cd239e1
zbf513c2d915b3c1566356e05280bb073d766ea48dacdbf646193ae67e62b8ee33accd147fd6f65
z74771ed0713b0150cf2bec7aaec665fcb485d09b457d295a20468f16473c6648ae1e05b7998b33
zfaea92b1c64f07fac9aa9b643f6983c50d4fe52e71184b473e01149fb1982f561c0fec09a59a5d
z4ac1c526e499545142c62ea0f082bad44552c780da9da39a16fa88a53617bc472639320d0e0ae1
zf99edfc978b05f6f20ac6d61aa16c6495c148bffc44321bc9a9bfe799b170fd1983d5364e499d9
zadfad0384657141c7de3e91780a475ff6a91a396f0434dbf6f5e8a976f0f6455fc229ec64ee1a9
z9de32822d3a3950e236664d5b8ff7fa634ed331b1eb68b9a2358fad1210621451da66073819040
z77d68bf937879ec0325c16c67b25c0a00fc262fa90782b3e1e26bbfef506d445c1bb77eb58e16c
z776f3257b5671a3d20e10a132f400fabf8dc5c498708144ead0e88a411cf47f92eb409e02d9205
za2eccdf18c2ba363c8ac3edd17246d42eeef0fc4b1642853fe5ffc38c65cd8cfe1b16be442f6aa
z8fa9c1ce48b4bcb6a8c55b7506d087be4911466e48152b373aefda445ccff519dde5c01a9a100d
zbe21e095233423affa17ab9bcb81166d391d364d88bd8771ce7937241b52445f7052023969ae28
zaeba198750555c61ec386e368101af590736151ef72e27173e2b4ea7f8b994082b65010b7fd322
z3f2c7b240ccd6ef712f7a2eef242b1a2298e3b807487c2b4060b897990521b9df09c5549b59197
z0dc81028bbb176008d28e1a0cee8af0c24eed7074d645a4ee7d955574f4c00ff07dc3256396452
z0017c0d9dad9b16a07a3d7ceb9376311b7367a24dd3b550af9aebac4c52bf8b62a5215b86d93f5
z8606afc60a5ea9823da56be3af17307800e20f8cfd9f9856ed67c78db6172b498c0d74fa377f79
z3bd4f3aa0740cf2d8cc9379bcfd69735b36b59d6a4bebb002ebbd373a360289a28681ff375708f
z55ea187f5faceaefd63d0c5fb806edb93f1c4045457423395b1474ff3e215518f1fe958a3416dd
zc8d1898e2eeb33c3e61c10658e114f47e997ab8a80830786a6e14d229d339e0942074f677bb4cb
za115db9dca24f5676678f2d0947a4f9349b5a8e4c8277caddcf61521a35decec32566030b7b003
zc2217d80e0de65dd6905f283fdaaaad305350fe35970bbcdd0e02b34d1f149d7c01939217c6760
ze31d2a8cba1ca684ae654005337b91dd711b68b0cc69fbb2b5bd202d932abc6d44b83393a865a6
zaf9d2f5d9c03e5679567fa5cddf2afdb573d566e633b68f18bedb410da1ee40412b81dca975ca5
z6dc406af107491740dba7b580f95d6c5fe9cdf804f2fd9907f57f456562381b92295d767ec5d10
z027bbb84afe57e9958feb2152c62a07207d22f8b60d1c7891c55ed9012ba4aa571313acab03815
zd2f6c855ae7d5575c7958eeef3ed1f7446a6be08ed4d050096130a3e884c3a734b68eb6187c6d4
zf16eacf0526f7727303666e8e72896cb9154489521149635d5dd7f89f2ebd544185f5601bb4c91
z0c5a4ba351f0936ad02d13595e0a055e15c20a639cf983222bf482bf6bdc2994a04f02f410be54
z949bf4a4e74798ec6370a9bd7d266bb0f6eee9d8053448bb4cb2bc6a46e8f454b4f9270e131126
z34a17787384be25644353574a89eb77f49624d9bed989fae65596219211c21e6a82a14630ea26f
z8b5a5757fbcb653c706945670e269ce96737b759b17fd43ab228781cc388dea2437c334a8de28a
zb8b5588d93e1fc307607a099f5c39abaf9c1bec5560eb3bd2df3939a9e1d2d31b6404238a7df8d
z6756de2e28f5eb0c6a592ef4f5c0e18b20f541bd2fed5956e4f3e812c13a6034be7a6c03507a7b
z716fa70392ea9b2d9793c36012b74e9d28d9974ff1b70e6bc3f27f23e3303d6b0449ea71dadd70
z06d3808dbb7b1811714e75dc0c49af3792ca97469958e8578555fff35adbdf7787000739f1df7e
zbd0e1703df793c25a0710a80e84d0155afdbd3b59a856b6f43d3239dfcad62f850853cd895ad7c
z759edeecf7d50a948257424112781713690418e1444da289d0264a9c0d34e6cdebe04625a2b251
z4f360bf8b81e411642cf7a1f2598afb8fd9bd101c9c9dc8744148c23398f6f991b44c412284ab8
z899468e38c5ff7647ab8e9870eff62eb873f1264c49bca5a7e396737894fe830b1c361da8263a9
zf1e0dba4a2aa4c0ec4c925e4d1da0df9faa775293c8dd0c88b7b8d0f9f6b36c143261cccf8a624
z4846619469348b3fed3ce8c1fe5d86efbb3615bd92b9a80e0845b7edb9e746227398319b2d0532
z677736c6887c9f342d9c5cdac960ffebcbd9eefc577e0668ff4a47bc0600469415a5a78d9ab4f2
z7cac677d78656fd91b292101d994f17d1ae84b2458150143a81ae144ad60851034362fb4a08c14
z64fd3f7d77bc5c5cb4393e099af48b39b6ae4f3d192be698284194189ad0803a96f19dcdfe5b99
zf8af66cf535e4b4c3c6c998a6f836dc26483de71304d3e9abc71b2f2b5d579ce34e503f6791e32
z7ef8de790b3c94c12f6648354626926fbcb42c211a0bed5842e327f601ad14476d352cf4d2a328
zc0e43d5f0412ec5c9dd674868c4b73b10d7dee6f6d6dbf29a8440e52bd045d74862da62286e6a6
z63348c40a59485c550797e512a3e96950c9132632ce1d58dca2831a8f5904b7c69746280cd215d
z07262fc6a08080b8f0d46cef4fb6883216cae22c565a83d01c4ae9614b8292662d3c5ed83fef48
z3a22717bf1063667b98e91343d6e7414ce8b3077446d011708803978f06ad51f1b445be47d4425
z1d5c9a67d151769fb89e71019d44dbfbf9c8218033e4d32c432b3a5eefc53c1a529f18595c2840
zc25aed2912db7239b6ace0759b49e35e018af685ff75f2edcf464776ad9bde3322350f6ebdc872
z637dc7326faef02f7778f38c45865a95a1992b0fcbaab627359cee5eb18c929403bd804d74dfaf
ze62c1c1505c089c79b06f7025cf2c65158df24e268af3743473369ae7d082edea03c26d896b9af
z457ad91724f62947fab5fa8e79d89aa4ef81889b0fe01c0b2e17668bb21e1ee68ca25847373afb
zae55df4fc11b8e9599305b5a0d35e38b08f51e3439c504118ed783c819b8993b74d9fb2a203380
zfd7b09509ce5463cddf4e5786db7c0ee255d69f820d564980c47af1274331039df7bb12ca06bbd
z81a93e9f19119a489cb385d92b1974db120ac1ff15b755f7adf2ac0634a288c1ebb8e6cfc46a8b
zafe0eb3dfe356b38ee3a3cf24764db1e62e566c2fc7986d83045e52e2f45af7bbd09d9c2e3d7ae
zdf466446d98f20538232245c8b42e582c678562f364ed4e88fd3b02c82bcfaed9e1facd479cd93
z179f6d113ad122c09caad923e43b9ac87719221d2979802ff5614e6a556a8b7957bf64cf8b91fb
zc0427c1b8faed5b19340ff4136b77834bc874007c7b390ce74d521659ef14a4430d3f4de5efc41
z52f480cb91cd5686026c0da0918279882cc1c92a0ace67cdec86b681724eda15730f64f8106d6a
zf4d47ec4ddc898d4a1fec597929dd963b9737a99e1a8c6caff51365f8b48a631e2dfd62bb494b4
zc918d73f203aad59bcf371c564d07a94266b4db50a061f475fddae4766572a84f1990c5427c56a
z743893a37cc012153a0543283e7eba01074751cbc732d510f5eb88a049242a87792ba46ad7da46
z17882101276d387a85d5600bc9bd52c594657f7d1ac76c3543ebddd8431234df173a923bb8cf80
z0aa96ef2f172bfa51d281439539c2bdc38c6402c7ebd20cc190fd69969d8a91653eddbb2ebdc01
zc507b4829e314a78a3b07ef75f533ff0bc40702411d64842a8ea2b6302eab333c89d96dfe242b8
za9feab6d1b86aa6384bcfa6b7a551bdcda5d64bd25d315359a5edd5cbaabdc86682f63cbf4c905
zd8258ee69557446fbdf58be7a354cbf59669d67a0fddad9bde7e88c474f0fc63e23c886fffceca
z9a310226a819f8287d67faff452c623a027f4768c01084215a5fdf64bc3877d0d4487eb5716d14
z060a8990745727aeec7ef2b704c768f74541d1419c22e75ae31f8d59d5674148e537a3e6913d7d
zbbb7350160ef1074bf3395430be6bef384d601d9b712000ec056283f2c23ca8b77353098597008
ze4d24a37e0505414a4b0f4b4c19425d69e10773f9e5a5671119f719b583f93b8f71c5f42ed073e
zd71a0f1cb3a609705a17d0d72b7c6c1229f61bd3244f1cc0bcd5df73a12aba38a1bcf1b3c572f4
z39affde848f3be020a640d75193b8f5f6a490103418e3278181a8a173f0762ba08abd9542b0176
zcb1cc45c40e9325068ffd839479b71d83cc5369bc086052ad6e45e5f094d23117c906d298c3dfe
z76f72a0cf6f03a92322b7eae0747b44da0dbeb353f869c98790a5869ed92c91f7ecfe443b5127a
z897c83ea22bcedd74a78c3d5d6a3d884f1a1d3f7cd766ddc25d5b1a19a5d0b47ae8273c005e37a
z11e7185c45ea64bf5449260cb9464347c3ea732944c5fa345ea574289e540e419a224cc74d0153
z87c8ed22b5f78d425a97d345b731619d00cf61b68a68134e19cd26350a22556663cb13a401850b
z70a124ef4e9a7dd729ed328a38f0e72b0dad3d3d74e8eee6ff6c09b37652eeef12c210660820b7
zb56d6d8930ccacaf5401778dd474f24989e167c204ef71b12ee5c466ce36ca97fb46d05609cf48
z9fd7c456d8e6324362a4ebd5db6057fae18ce40eef7edc958e9ebd34ab0ad78f33fde1be8c2c49
z60a039a69f08842dac6b573dc526536598969a0c6ee1ab6b77b2270e78d9861d42104aba3ad91d
z8eb19c4c797392161a47a2652c397abab699c7a0c997414f06e8fe860a1d5d75b12a1d9a489dc2
z0dbd68f6706066823bec8e5f5d35268a08610e683e4240bf0c1bb583e8fc12124e4c3f5501e4ce
zcb424c2b214e2c67e6740678bc62d8fb804290fc7970e320e64606e7930d4e4e015d673fde5f46
z97b7a2c85e3cfc2b56e047e4aa4a5583fbe3ab248a60959bc1afefab345ec33c4ca74805ed64f4
zd46fe52ba7606392efa07c8aab4b035d3190e1ecf61ed35d06a7c6555cbcadca7d789a00f88763
ze765e89dedf9fe498b46a00fd121ad12b950836e335b23aa260add6b0a5619b0cb121f60371405
z679db5b1f25f6430938b0a1c769f27d26976d22a0a091ff787d50fb1165b49ca987b0a1677e51c
za69c22514a9d365a17ad237f73f49b6db1bee31d4dabf409c5d262f5b443ba6438b39037f5a8e4
z69e3ff072b6a4a4719ced492e6a45ba860c1380d60d8c27499aab1cfbbc82b62233faffebe8256
z26b272ca31e81352cb69656ab1eb2635e153ee85dd0b754abc908b93efb4c3061c2ab52af2afc6
zadcc85f0b22fabbf5554c45c9fa961608c93fdc69b62427a9e5938706b71b12d3fe7c9ad879038
zce98b417900a59cdffde45852c71edcb2c37c8a4f5da9da842b09805e1a3b86a948e2b33a70b48
z6ce5343ddbee7c67358b34afd8aa78298aba858d081bd7819d2de252667ca5b2a948e28ffe9f81
z96a65c14ddf5d5b891e13703d967797f134eb305b69b23a2153cf70a22b57bbaacfb1ac165f6c4
z08fb19e45000fe9254938a34f84f60de42288f6293f6a320da04c1c0248fe8f0b15d2a497ad817
z55a71e3d4e5f6d27b018268dc6e6dcf8b97f0e540285f09aa8970f16c776bd5201cec687d09d06
z90f57c836f9c2ee51059fcd5e77e105d8d24f5cee6075aff28ce7dc839dd307dd2df3103c0851a
zb0c6bae239cee77aff74f195eb292d4422384cdb6a071c21f87a73b899ca994631d828ff1b675b
zfbb7be75b8c348bda3a9f65f412e71a2f43704b138f93bace73d97fec9b6926c6c0b4245d93990
z7ee2dfda28c9d1340d898f7c844f99fee62a9855081097c7853c979fd6a7a0babd2bfc4847d8f5
zf94887fe4e3c0f2ecb0134f1b18bcc838c19c8991f43595470602cca09ec50e23d0613cd3d5267
z754c79d74312c51e65b7cf7c86e616cdd442e7345405b2064fb1682abad1348136385e89a1dc4d
z8021605efe7bb1cce67b78d0acad85eaa7d38d59d5ea25c650cb432ef18ac41d887923f7af536f
z5a133ee624987f0f21a897f5bf8c6369f14bb489e46c038f546951d1343fe0ee2386b77647a93b
z5737eee27fc3a764f512e9961870ac6d757ef51e23aa5ae9d7f9b3f73b25303340a8eb49cca285
zc5666ea9f84ed198d2becd21c2e3f051b8ef169b476801fa5f5fc7adb494d9de0787ab12bdd40b
zf024abd9e82898cda62247f38c6c845f78ebc214cf58fb6211f0d509992b1554d20941ebbd413d
z976f71c486344877d8f12c40934bae1d70519ba080a141ea0063ea6c6510646e1894f5ce7c65cd
z8e3807a1d725371ffdf14c57d25165fc056d0743e0e3762cdea79ac46c271ac93ea195f4b293e0
z76cb58ddfa08e963a4584cf0e51b1d832175f141181ccbe1c275eb4ffecc7b4d26a7806a9cf7ad
z76032accff3f8659f0e0682333fe380f56db816aa4897a572704eadcd3138a7abe59bffe79402c
zf226c52d519626208e061603473b3bc909fa959be8f065656374c41ef195524ba68273a31660a0
z09e7022a3fee93f4df3c59550c91d2c3267c3fa07321aaeb50d107d6c45d3ac45f87cae90cb976
z13f575ddc7491c7b11f6fc3f247fd184b50bc2d9589b9f68a3f4b355e2e4047ca30d2c61bfa505
z23b49e0922bee6173f4a269e05fcbb371dc51f5dbec7519223c7c7058bb3db49c48e6e4d467451
z0494e64894f35ac9601e57329be37f7e1ac6437b783702aed721c5ea6fc2cb020168646e047e97
ze338f35bcc3c7a931250c320b5c79d8e518e242fe48ae8911643b167e86c1247746e8ee4c02f35
z3bd60965b4bd074ea27c1ded3567160c32af2597dfe6ebdebf3168edcdc789ff899ec6f97f2570
zc74d6b739c488b19a6af4106466fe0112feb21e6ad9216196e613eda9e6425d736ad26df0f2594
z6a421ae7651959b5bb040ecbeb719ed90e80d736b5f24395f31d36c08fa5c6b44587f0224a882e
ze54d2d0c48cb65e2ea27b0cf1d4b06fc610211f7ee6b55af86832e45407f7e598157c947b92f07
z81bfe5bc76f98093481f0d81e1b0bd766313c55dfcb2d304de4e2c4009041530fdc96f1f70974e
z782c0143ee038559d89f132569bb0bcb3c3bbb2004f9f38fd408ad90f5f11e76ee19efc090ef04
z574a81ed0e6ef24fc5e839f69bb7ca5e01cb3fcb438010941b71951317603ebf9e32d82914388e
z8a97c891768dcd3d4d7ccd424e44ee55a8d9378e6b73a87d81552d1c1356551970fe980091d4cd
zfae2219e2037458eab61844f0e9b15e0a0eb83139134f3a20b764b52a728cbb065c5c58a52de9e
z1fd930273e23c5c457ec489e4611318f3c657fcc361d776f8f609ac7da56ae2f25e3e0ca0a2503
z347d1bc4813076232eb3eaecbe3a3cdd452319cd757c06d52e950736832615f8e0423015609fc0
za0f74245b3d103bdae60de8ce569b25959dfef10d213ea4314cc888e49af83c41cfbf225e64d6e
zd5fd2cd6f67b82ccd32d1196cd096c82c66972ba987652921aa656118637420f02040ee54acb70
zcd42ad8139151e85eb97c2a9236a282ddb6a9b5b0385e2d684a0b1ad91223a98cfe2866fdb7f96
z10d6f795cb765d4f052ad34a7f04b082b2931f131180148f14ed4996bff9a02299a41e7168ac62
z7e22bc2759b7902002af5e19a23154d65501a3c9a038e641dd9a4bd4732870f4dfade8a4e5551f
z4817080f2cc1bd2f308399e506a22ae6d16f79efc203c4bec22063be334983c92840a93b35888e
zb48746ea64afce311084aac08aebd7f9739127da608c20467239a9d7740676bc9575cb2091eaab
z8cd8b8bbf8abdc9b66600419c9b5a27825bd30a803ed2e41e4bc5487e79a81f511ac9ea122c419
z90d5380dee28a4e7e8b2b81a984b4f48c9b34c85b56756a112a2b5e7cad7be2a54a0edcc43a5ab
ze1eab7649019e7bb1afa58facaab007df2e166ca3283e8862faada0ca2c8428da9bb9925826f41
z9115cb30ee7f804a1e92f7bf18af5223a0fcc7e994b85c220d5d8f392d4e8523053c42a035ceab
zd26a7c8c5539256453af46d59da391d2ff62eb30f76ff7ba07ed7f3b4860d7d6e9905fbcc66795
ze8389c8968df458738b2c87923e61828aadfa06b86891c8b27ea68aedc8974b0bd01465fd8e8e6
z390d9ea2bb8f7e06e7c47e6d2ae4f6daa0d30f58cdb9a19d9b39f7cabc75e02c855d4bef80ebb4
z9d3a7a1ceb0322132ccb555516c77ef7b207c78b2628e38ace2c627bcc9cc8ec8e9b8ee3f686e8
zab6c6cd3150c996a284050eee7cfaa6f3a6071eac4487f514bf78b13503c4a39b45cdf2eac7cd3
zf941eeb697fcb31f2547dc3cbdf84f0041187514140b2815e345873888a8cbc7d7f1d09a16ba33
z6bfc2faea5efffed4683b39f6e60ea5bbaf4544c64256c5c6020522ea36a105259028e5898be80
z6b7e844c384027581f654352d8daba67da4475a9eb0b93fccaf2beda34168b18df2cd552c7f06d
za97b9cbb290904ce25ff2eafd04b765a65e1fb3ed6286cabad8c3b16c2cacd3c87709714552964
z31bf8433a47ee35857d3d6e1103b69bea113dbf804754022707fc8244e873cf6f8354db1da306f
zbb39b0fa5cf63ea34cb59b414b4b5df672e936c5a55cfa46d7d1c680678db07b4e12bd58fe4e9f
z03b3bc762f5fff798a0c7eac548ac8cbdd999e1ce5779c9cbd7f42419f3d8554b948988dad2c24
zd802b6b2d7302b8f89c5ea32390a0c51a6da47897cb7b04dabc5d73027f56c54aad6fbd22f63f9
z20a6f10355e9f3430ae68ce2e95a1c43686a9d2c54b5110f84c3d69f72490d9fd0f796bade4921
z079ad5a94b7d71f4619d07d1eb334c96ec485c3dedf9c440f0d9c32c904bebc00572195deb1ba6
z7096bf5fbead5776b17effdd2e8ad3529e1da533ccae1b93969bf3b6f88ed6d02e8e55b51b8aa1
z14c8ea3cea4bb34e7ebfe3687f9e5aaa11425dc50598c3471a7ef348d4c70c208e77e392ce76a3
za16f8fffeff939c8150f80804c07b5751d0d2613a23e81a4e289e7c12e6846a88d0d993c56ee15
zddf015b7ac1fc4190cc8f3518b323909083282d1f91c8ce4e339e6e82bd3e51febff2bd94ee600
z6a412b07471023cbfcb5cf3c473d0a72107c2b5e4a912a08b894aa28015b2077c13214c44e48dc
z0c1e94c31b332d961cf9a5d6871e6407d49ef6126b98637cc3fdd900ea8e68880c07140dc06f36
z0904abe48ddbad823fb0cc69086402d1cfdd21b4de0991d36d92842ab73b6bdf13166a4f79dd45
z21c6a46089624fd74d050c4a4fd1318c179581c53ef52af3139236b8f8e80660a706f3b85ff13a
zea108e0118b58ae2b2ed4bd832f023a367547f7bcbe2f212fa7de09284cccdfa4acbfcc400838a
zc1a603939fecba7640288fa83042a0e8f29756d91e4f547fecf0dc6241773ab722e7754be47ff2
z7cde067231c72750c57d896effdeec2663a8e46d9bbea60cf1ea7029690aada9f7d90cb608c677
z734ec79699e0324917215e5d641804667454da86bda0329beea5ddae072dc54a61f1247e6ed647
z11e12fc916357529ef51ccbbdd955fac98117f72671d8cdede2bd5f9446602f8c2df2fb6c486d1
z0514c5a2b92d0560fe5f77ec671f183cd8bf5351b8e07f304f5e3a2bf78bb5b605c40175d0bb41
zd2ff804a782ed1b2f779a1c3468f5e7e7fce6fc5df74cb63670265f5387fecee8a4611ea7ed68a
z491a9ecf80b46e2fb898e2bed639cda88f588d7a512d0f52cd53f375498c054b8d64261850d311
zbe0f92993a131a4c457b1107706de77f2ca87a9c62ed1c0d3bc18e53bb1e249e8b5913675fc9ff
zd81693ad8538d6a59d6a10399bfba88833b36082c5342c5b85c4cfdee8bce1e5d20d465ccdca44
zcda9108448333d49451bb69eae6e0af16ab2046f697bf12076852b749fd130f539def12cc06c69
z424832133af0639c8361597146a2602f5a937952346a6e81bdfc6b23f5356112ff520a83d62b74
zc5c55e6ed6cf1010a8eae0c628ef4c6ba4f3ae0c9fab357517cbe46af640fd53125867686521a8
zc7ca4de36870f16f3b16a30d597b25edb283a0b5736c0dbeee9587927bad45e63e0c6ea848b8c7
zcba8eb802c76b2f37ab8c4a6e87920b39c47d0b5a5ce06c6b264cf3e1aa05549b5ea37d6ea85c5
z6bf52fb58f0dbf0112daf660357d1f925626cb395aeaaa0d00ac373608758c375b2d724a77e769
z6816a5775c8cea8d2461d7265f4558a247f54dea6134584e01bbc90be3427d445088313f8166b8
zd6e6400725bd5739b954f9b62437efa8c9b1c92ef0abbc46a91c184c341b988ec9f6b7349c5b2d
zb5b0e70ff50a979f49d08098a155b63632fc475d61cfa7a5fd3d646c607fd0ae2f31ada90b3a24
z49e3f611a75606d8f8980d431d1e2886a3fc9dbf435199a5958107769fceef41736830eb2740e2
ze21badbc26c5ebc97a70229d28f074ba7c8b3e5e0f53386052f871972842784ee0eeaf94fbb534
z266eedd7843fe687bbaf10134e53b5b2f8480fa4ff050ca7638a6898b1269f85c9f053902328de
z3e6cc78e2dca86bd51f43d82fc756c6936ca7f8d4ca7f642ef5711e64fa1b50d8fbcfac7426db7
za37e77451551d4608e05450097e6254b6e517be70491159381d49a61e4a4c906b0882b0a670cf3
z738c79e35506d931885df94a7ca2b4861964d57c8cd2550fc9bbab9a670998585fc230e0910993
ze2ae7bab6d5c69cb65df8e161d036c6186f14295bb66f8b33a891876562d48f67fc62449089a84
z1626576ebf2dea5a2bfcef67edc472bd717cdbd64cd583256d9da9fbabf069c883d0caa1ada1b0
z2a4e1a3559ed00a28cafa2723fef40e8d8a995ee57a08d37761cb848ab7d6590c731b0d32bdb47
z8a8fc30c59b8f0f889daf1fc73fc89da33bfaa998dda77622d1265175e3fea15e6e438943f3ca0
za7e82364633bb9abb42cde2fd13b72de3f0e937627c49a2be717ef99a5dcd17d5fc40719b5c571
z5caa0924997d53818e91e360da2e04f6496d23353140bb6ec5fa8fcd757a277bea2e37bf633c83
ze1da7f50b9e101df1f598ce4f04b78125986d3010c99eb6931f8c54ea8a6867a17eae455e86362
z1910fe814d29f1605e2e9594b09a5d0b4f36876c06ad9043482874ae76aca0bc75e34a9bda444f
za8c154d33487435e3f2c411757066a4e0f0fff1ed1c1b0694afa7ef80685526663273d579e3c3b
z3d1369eb62ebccc5c92639dc303b6f6b4b2d4e78824d613151168b59b9738871bc60e86079f3ba
z5a6ceeb0f4c595386bed414460e27d8f1f6223d380b8c4123ad9aaa8799ddc16fc7759cedcd550
zce77a132888415d047ea9ad7cc38a1e01cf7b0cc55f3b96d252ada67b30887ecab7d6d4f1d811e
z8194c004249ad04a7e860427f3af11ded05b375b3d9b178c1e9e775f8ac470eeaa163e102ba051
z5ccaa879070c400862cc95d35253a3d9f155c6882638f6fb54bbf57be8ffe0208f2e3b8e548bbe
ze3f02e341d6f0ebf501010508ddb4da6db83d6e12056a8588dffd03c1e5b31c2becd6b792cde6a
z113d1d7c97b34320d42f53859fb44fc8b553e4336f221830da51b07f1b46c9646d39000273f9dc
z6384c831d4789027a6416b67b19d9fc45a02472210b7d80559397119590a6038a976d6cabd1eb7
z408f3180d58e5b51180c31cf19eb5ac533661d4ab908799358f5e7e9451b48d9c239a40eb28536
zc35bd5d26cd5fa4c504df263c99942fe338b1495e5a0696c0a88cf53702a8473fec1d6892ae744
z84296d9117bba3b4a4909a19779484892964dec25c08453e9577366c441373a1560ca3af4e8b30
z491f6724e7f7921135ffee9a5a4c1a4d8983be85d946e6e26ebec225ad245b92f819378456aaeb
z48d61602f60cd0c0318cd43aa371638e420092f1c8eef4ad71befc04a29fa775fb8e1915a10305
z85200eb9968bdd3eedff4205c521a78c973b58fb82f8e414ebac5305d37c49c15d557757006df0
zeb9fe0ad0d23bb49d1ff1779efc5d151e43bed7e7f164b40764745f1b83c6c9ff3c05e9084761e
z01a5a83b6dda854d8daa6e6f3d5883c57ae10a36d7376d2273a95efaf8464e9722b88b70cd0a72
za2e6ce9f8803e04bc53c9dc4b243a7eb2f67591736cf67a1bb99b765cc933a0f19451a3a143db6
ze551edca8ca5886897226d77b1a488f5ef1abaf6543bb23c07b8b225ae3e212e3cb6b7c4e32528
z6e656fe30508a60a19dacc80539ac2723083f721793d92ba51da8131eb9f9604714715109f1337
z16064303d99f5861f1214a0f51842ac015750dc4c71908d0040b3ffa415ce39b17fd1518196288
z15a8eecf92133f6942ed0fe65d8cf47a2aa1965adcac481a605a9bd23f7dd868e89147bd5a2d15
zd2e31905aa9a5c2fd91664d3383d583b0826df89675379d75b19f95fab64177f4f19e3d917990d
z04d503d48b53e556883b170b277097d2178fcfccc5669c9afb76e73bac7fd42379cd0f69ec301f
z17135518dc5e0db412a30b5fbaeda966e2c84c190d6e231d864185c4d73393d7feda1ea902ce39
z72de6cb7f7d40ce0345d8cca019a8421a189378ce35c79a551b5d44021a425492c596456348f55
z7f63210dc401c929350c08378179ed6b2eba7ecde1b91804c377ed677268776fd8b08a490a8cfa
z1777cb7b615ca212b13e3ec9643a70e9ac078545c927fcaf37b4e2a1038b9aa38e275abd652ece
z6dc813bf7fc1bb0988db5aef773a0297ae20d747954b07dd793bc8bea4d018d294fd45f9e31416
z83b0acc656bfcfab412e73e26c630a231055d5d689d92eb33267f4eb7c8df3c5242ae7544a341a
zd9acce8ba2fb668b7bf789299f141195a9e23345c6e96015caa8e48fefd1134f78d0554c4e2fb5
zcf527721f736790a2e7e7cd3136f06c7c3603a06c7758262f690659b12338ba692f276c06ccedd
z4238a4da3f4cf8b44efde0e0d8be481d53db8668447b1707e57bc9c17b292c488da8ffc17c1b88
zbd683bd883e852c774064608e861defcc1d245e55ffb8bffdeaef4fceb8dfa23585293eebe50b7
zc82fdc5a4de1ce52c1bb259ee883fd90f833d74259127b2f2fb39075533390a29f9ee5d3fe6034
z4abe650916a519dbaeef80705b67a0863329a01eb2df54a16186023d1c88349bc0d32227371d46
z6a1f7e484bb879a3ce3be734ed06876339fbb646c5767dbb73d5e21e2c30cbe90f345c0c0e3a29
z601147f796500b3c34e5318906d130eb1e0bfe164a3c69c19848c45ad3f0897695e0b774fb0a55
z80232e00e33045e2779efe256fbc1f5c03a57f6f8358cea72eafe70ddfba07861faadeabf8754f
z43718ef33976bf368f99751cffaa9d919283035a9d6cb0eba4774469c33da2fbbfdd32635ab8b6
zba2c0facc2098bda4287ed01f4941ccb94b4a1afd503e8eb640751e6174683a5bc5e823e2c44a2
zefea359c4543b18fce94015225fedeaad40776b15be08693999e1ff23adddfcd7a01fe28e83e68
z79f7d34af5736b68eaaf152afbd5dcaa78fdad3e8e28762131c3bf32ba7d44e7558e7cb78e9c01
zceab6549b37beecb670f6e8d240ab3a353bd0c49b086b21229219690ce7e32f6d06d519ece97f6
z8e4a87a03f84e15369a07ec057de74056ef51ce65f483a2de5b413e492261a718fa935f3715583
zb645544eedb4c47a676e636a51fc8338ae4a95a8d5e04915fd43b04bfb314b6e3c7acce653f369
zc4a5ffd8e98247df7c7812fcb5c915947f9df0e2b70f891b639aaa2252a81ecbf8fa94fdd0ce78
z53c28205a08368ca90cae36f46c724e35673c163ba99d40ddc5bf37daa7e81ea09b55d8623072e
z8a3c7e1363360490372f5692a695a2de2ddd8944a4b7a1c6243f2f5e8f0c0c0dc58dcb510dbfea
z3810f3e3c8918bd5263f1c1f61456d50665edc639fd810a2c3e7f725561511947418120ffce2fb
z450c212df70f9ad9a07dddd4690e39340c81898198e70d575571eccb4aaf6003b451c6e47aae28
zfeb4396e5caef4612984dc1652e0d5cc7c37f1fe8f0056ae5cb89d00706acbf6ca847c94178233
z994450fe2802b93dfbc2b183ee85a689a1b46e53b9bf9100d391b32fb859a19f2230533061326b
zeb42426a7e49fcc299568e3dae4e62f81aeb0b0271647ada4c8ce70a567bb44e9d7c94cf59e043
z3e4b9f258c96c5546cd6c03dd9ff9294299af315390f9350c31d5f6b1e45964c1f2c76d204df62
z519901b72a99ff7c4b61f372d629594fd99d3829b173d62ed7d549c42fded5f23d9d8caa4f03ef
z0428fa019fa7d707ea7d8d87330319e67c47512bdea6e2db2a2045d14a6d62da6b0b526b0e0c97
zc3cea01d0e4ca6d0c72f7b912b9ac00c785f79de350d482b7d4ebd7c5bf405bffe1c1d71315df1
z7d39b41042390a3c8e4c03cb56b119650cf0a9449fd5c0acb36a347595c464c175990f0b40a046
z79d23bc4deadc6fca312c47ea0d65ccda4663483049c264165f79ac071b033f7e1de0b999c3ba8
zdfe6be75ca53089b61525e977337b112fb40060cbc8095a031552390c516b91f4d799e43fb7120
z97d5ba7b0e65079a22410d237ef33a11d0cb0a2b838df5d06a6d45641b5193c407d22d95935b90
z1ba19c587c3131e801716027229909e579f440b5625a122e2dabe6936471c11d43b482a993676b
zc812485bbe6632a978e8bfc0f8371155ea179089ce059dd55a31160504a009ad14a52eaba98d78
z539ce557873c076763ee769547ff27c495db3d00792074a1a7447a1eeb5c045d86eb5e7ad46e74
z6fbdc96cc8db9f1354ade351b5435d4d75973e8a8276b42a3184dddc206c494bf2e69fb49b312a
zf4f80b463c2079a5d57a16c4877bad99a7396cd1218c6b69dbd7aa357be985c2320c8a45289a0f
z667d74e4484370ac3c73475f6bf32facaffd904dfd5e3a2721dcd9e09f691a28286e7dec27a980
ze121aa0b97af92653df0397d36481036bd03766a2fd43227ee94a13cd199d931a9bab19608d046
z2f6debb5aca9fa9d2369544f9993933b08f3e2d5995d3dd2ad90015f4bacc54df9ab7262cafe0d
z7ff1abc7c63ad7fff7b213f64b579805820cc3f550525231d122db3f7a6307573f4c4cd8347dc8
z5ca62192423d858752c25a7409d829a17ba70a2811e7f05ff0d967698087a6b259a211a516eca9
zeb90e0acd364bf4937b30ec69821f9ff3058bac1ddd49a04d52ecde87008910ffb3b19232e8ba2
z24a86a8365d3ef77910431725b9b3ba46fc513a7432bcc7c1bdbb91167c1096b1835578958d602
z85d722184f3f348135a83f2687a7575c8fedde5a58662d0b969a301405e0dece252a2793d99490
z45f6ac8e54cb4ce190501343992293d70728c62376a4c14d210b66ed51f29ccbf018c5ab3dc00e
z765055c591fcf286ea8e66907a047b9d33729e4de6ed36b6cd2475b70f1fe11a23df94c199848a
z9ff987af4df6a81fbfc6353b054e0fdc1fe89f02a1bf0c83c39e20c2ecc939f96382c418eefd75
ze8a59f19d1eb4a2caf42054ed3eb3e89c8c411479b13c4105efe174a4866f1a2184a3655cfc16c
z5d1358610b64640f2693a99f3411c2cf406223d6f96a7ed0384dc838fdc6fa5a148b520bd2914a
z5eba4415d4613f6e1c7af239c6665c0749641f4941e078c9e30c697971451f1dc06c46dbba542b
z6de268d76d9b63cd1f14d339e4ba7530ad385020292077191a12cc83cf38907ea96dd4eddbc572
ze076b41b385628f6c8dc714f190b506d0fcb50b1c3e911e9116b40615c80729a6fc16bce3ae2c5
z6ef11371fc7bd0e4247e037c6130f95ba5da4cc647f8e6573fbb49451ca3f971f814033860d12e
zb5dd6e1bc6e6bd35ab2c667eadaf5bf0d541b44670d0ae763b802001240bd8694197493e5479fd
z4af86a45a713000f84cf3ea6ad865277aca286b916d5ed6d10067f615a48f2a0aa62c21c581622
z73669b5a9f36ab4a97dccc1611f0ba6410045e504c0aed32279685ad09afe43ec614c734c51fa2
z9fd017899ee4e286f3dc15580a2d1e353b88c151e9b4a31c3c725f72d7571577b5b375627ebee4
zd0385fb1df032a26556ed567d84653cf7d773d89de3e200905d8c74d07eb29aafe5e332acd0525
z46222200bbf752ab783cae2f2d3fa28a9455d04abe6c76d2bbd8df60cd99b2baef1b91b5021021
zaf670910b7e5909aec4b00c0e3aa772a8e33d2865db6847ef0c4ccd5c6c38b322c311109813af2
z2a085ef15bbd13c0be262c9ac41a29597e6da498f4ccc9e6252309098fbb1a4b1d275a700ab80b
z0dc240904de4600604e2f97bb09601fb303cdf15ebadcdfa5143f16dd23599905a5004d6032cfd
z3ffdd85861191778d3f23fd2fb32ee7cc1e81941eeecad7508055f7abc136683bfcddc251d56d9
z56c7cd64654139870cc51597be07742f15275cafe6b931e0fcc6692a8c385c9e969d4bb66d91c4
zdd211dd6078dbac3666f470c692d10bc409f9b0542788508037b64e78a2414ec3b458aa48d8826
ze9a5bdc30f297ccf193937ffe5e4ddc96cb7892d758625f38a1ddf33c50707c0d0aa2371f31120
zbf73478e91a50faaee1c5c0e845860a07ae261d8d6e9527630680ef4bf63bf4c6aafa904eb4284
z7dbffda91e1dd70cd90d074e9bc1e016e6df838c7b887b3aa3bcd6dea67c45cc5ee43ffc4286a2
za3bbee9a6231ecb00fb890481f99a04b985d852656fb0860a10deb929a58405dcacb7621b7294d
zcbd465820f9b7776f7ff24022122f56a60440a1995987142bc188a599057f3fdc407712d8a8bd9
zfe3085f7671e44893c4e87844d8389964fc821bcf2324212634cff4fba26a983f644250b4062b4
z7e3e7b5c540b5e00e36064257334dd48ae261ac1a609efc20800ebfcc71ab5c85d13e5105ecf3c
z5725e3e0752d8456e49ad86df59f1aa47c2abec0b0d3cac9dc0084ab098ce5c9d2f36ff1d41b0a
zc6779d1987d93454e46db8372c76441c407daa65f315595cf74435fd877b50f26f34465fa54b6d
z8a78e6a8d411cd7bdcd85f84dbd628d54d49a76743bfa791bb1a8485babeaba21aafba9bb3b3b1
zfcaac3d9d64af1bce62ead6e5762a2e8727e743de8d355e3c291e530616ef3b8e43f1a091dc80b
z83521b8b812e40c669217d8c6a52aaf9a2d4669468cb83664c51f20a57c6589c68459cd08bf3d9
za64171832b9ad0981db016d298545282b1ac8aa55dd6f1bc4ecc1b3b306ac94e2eb2915357a1fc
ze54cc5575a7fc3aee607c66628913b2405889d63dd3405598e4c06be7a70966d762fc7d9ff76a4
zfeb74e44ab9457f443493d9b1052d7dc272175ead20a098132c4e8e383b2b87b6f364e5e250f96
zfedf74c517c0ec03734be05ded8b0d7d32e9b439386b37827bb6648972005deb6341fd696d8d26
z1d492958e702261869c9d5049dfae09af87433046bce1d562fab9f13e109635e50795f6ad0c847
zebd7a35d8af12ab4d3a8cf3251773d8c300d3794e50fd82ed38c834556b3bea24006f522d66b06
zc8409834691652928635d831e4cd412f0be705c8c3c1a915ce1e213ec3b055e5e68ea7033b4175
ze3751137b881a2f5dba7b25a44610aa8db435d336109354e79642efde031479f29f71fad0ee1e8
z583e4ebd6d4b837af9389fcf9e1a402b046386eb889e5c2627fb2a7fa7595267e18fa2c95b58b1
z61f4f6fd61e471be6f0b9662bfa592ee31060564821cb81cf926918d1c5cb68a9f98a863832e69
zc669771d04708a1e4db66f6177421f47a97cd751738494ded51b0d3c647acfa386556dfa7a6aaf
zea33ecdb372977c2a29ce3e545d2fddaded6b1aa746793529e89d365f3b5659be4772ec57b0ed0
z858841ebee7e768d25182babd36dfda080451a068239e1506af81e5c688b819f88a0c8c81c94e9
zb9131bb93c37dc322bb4d47396cb349eb37718fd44f32cc88b75df431ba089870cde0b9dc36c89
z1eb4dbe63d5b7a9903a40fa4fca85a59049ab157f40285f8d4256246bbef9189f90f9240c41cac
z1f5e0c209e89f7c5c8e83855e72246e99eda548572e57746e1fbc156857a9c8828d3f098b69fab
z00b10108e6b334c10250a07df8494438dc484774d015d9707fcac86eb16474ecd749602d55a0cd
z25b2556949aa8edd7e0998527d4657f39ef1db9bf417af20dc8b5c507844f708184680da819493
z84de7d30bb21fd693bd04ec377dd4f08c63bf05140e5e15ff2a06eb4a6f0ffa8256bdf9bbaba8d
z30c60424c049b916390056accd9e60f1866cff175764650103a3ad1bd119fb9a312b70a0e08321
z4935cf615e7bbbad2b3bf4aa0133e9560d1ab7910007432ba9a0a7bec60fd370fe54780681a4b3
za9f1c31a2f8b8841b4a9a4304293e2e22572e16e29aff0c0a50cb23b09f109bd027e3c50b2e668
z26641a4ea1e579e0fa163c80daed33742d4e81b3c1ccebd35f691b8280f9b14c1a4c1aa77e0152
z6ea7b89d95d217f9066b74ad17397e8b2543aedcf98206b319f493397f8cf8e91fcb1fc7afe9ff
z78e04567bbd2d4beab5ac8b3d72d46f6fe77b07c2764b3c7bd83f291a835a5fc655b7ea5a86484
ze52e00a336d1c3bb3e771f82d237fe4c37db07abc4e3a85d7e4fa07714b8719765789fa607bcde
z6e377074d520803e25ec772057e2e767aeda246d3890efc1c00b72f3e4de0b529bf6baaf5f90ca
z1fe4ae55f644b464fa27c33828f1cb2c47a48fc0f7bb96febbc40e401d637e27d8c4f317f2e1f8
z72d4d38fd718da22e9e5a0c3d7bb2d8632bc23605001b5171e8fbef8119656b2b4f52d49e6035d
z3247571c4e6bff6871acd819daffe63922bb9c9be17e94c762805a764bc65e93425b8140d0f5e0
zb623aa0fc396046b4d5ab2749b2d38fba740b7310f851bc0d4f7e4619c27384ce623e6ebacd8c2
zbd32182df22263bbd4852e508150e6be44270d2bec781441b507947a62a2e51a6849fa12b0c454
z1e9ed2c7313eb0d7ee5999d7461374291eb57317586a1e4d0f5b5ce8be4f3e83c43af2df3681a7
za6d9a0155be733e6f89f27f2b628c3bad97cf83d08274fc4bb2d6af8f990c017f7d404552ab875
zc73669eda4a16feaf8c1bac45c3e7f992510ed1b221ad6c7c951390c1eb5f2421af500c72e4ed5
z586d24b844cb00a1fef8e5c360665060723dc67f00c7a50af947d43341378ac48618c31ce766ab
ze9e8ed4a60cf95eb803f76b3d1b273009976145fa6cd782ca659e84ff5ea0b2230ddbbc0c82b74
zcc3f630f35f51cbf4edea27eabe2b29f43b94968c0ed3126e0c20f317fd2fb5da58a3a4f845d72
zfa8d4da0b4a5b53a52321bd5d6d89684ef2ece3b4361d42de942a6d8509fa458aa66988bf52196
z8e69fc2675a13fdbc8d020118a03af5ef278b801b8afc2c297bb9f430b0e19ce6d85ac4b42681b
z65112ca4788f4ff1d169b708c785eef73af4c654f7c66e5cb6a15904dfe5e663195a9eb40faa73
za36a35b72f95baf0e38e8a1cd405e108af7c907ff573079485f8815f8cbdf1cfb2eec28aa27b37
z14b7b5de765e2e59be0a9c019f47a109018fc74d56fd860f1709c0c0dccef6bf31f38a3afa2863
z49ced8aff34d032da10673ce842149182c785782deb5b2ecaa515787bed9c00f1e9cdbc4e8a0fe
z9a232f296cac816ddf1e233aafc9e814908e61ef9461e6d59730d0bcad58224220d27b723344dd
z9959bf1198522500d0f4c2418d599513c5e962deee4258db4c58d6311954c3f7d666737b01bd4c
ze00715fd60d7aaaedc61f1fdb2a385ead8d09a927b28fa79ac82f1a2620fbb7b983a83e2417b3a
z736cab84937329d432f9f697b060fb055b6146636a366f19e8d427e1bab5818772e3157bfbd433
za71476f572da1f2853b2ddb5ccdd3e262fa2a72edaf4faa08381083852d01bc364250461d88e7d
zf91421dad734a98ab85f3b17ab06c29d754d20490a0fc3a4651616d2f58dd7190170736e1337f6
zdf6dd491d6614f113012a844dca497ac409e48ed96df067b6f14bdee4de5f29c87f3d4ea717a7a
z0e015a2375d44c0debd3a8a704de2a0279dde419369a0b3addf1ad893e9f665841bdcea5401616
zecd71f1737e035dff312b881c23e6888e05c89197b0d993357dfa548415b779bc7b815aa5e738e
z15e126c15aebfbdf08c74500426b554be85ca7aa4cc3246c08e9315d31a999dce3007694ceee93
z257f7cd5f7b8c1125dbf2e302efd3dcd10632071c99b31df76cbb77c40df1b3da6e8a1ae20e1db
zb409a0f39ca257cc48377c9e4b80c120e39b0c179dba569f51c490abe898cd3cea081c05836616
z13ee9c0c57e7ac47aab79f7166a091cf1b50be228dc3435f2e5be59386640dde08259b226ee4b2
ze47ea94e516799cbaab5eeefe8963e6438b4966017eada2d38045550edd9b2b0370897c4fd0b99
za86b17969105486a97a7b0c199ec538d15838289e0055188a3734978b7c9024b41c1578516b89f
z8b38572a94a20fe3122fc10d8f569b871b819cac55dda5c22d2cf86c708865c82bf529b9a1bb25
z0e487f782119982cced81ed9e4fb4c9ac54e5331add7607a960084749a7b80d9b785ad6c5059f6
z2d1ee87abf0fbbec43d65d1c204b38f4d83bcaade4e81b7922655da74388ffa5a15e5657a6d624
zbed042bb7d45d332f2a1cce78e9580b3a1ea90405db6be4d79203a1c32e6abf4b534c5c50ddb33
zff47e4517c4f6ca1cfae06f2d762db302ca9c6a2bcf05394ee64dbb9d34526e37fe68a93172289
z453ad8a0fec489b373ffd1acaa396881286925278d44d498e863302e394df37191ffa18e8348f4
z1c07c580914a29a4a750213991ef09c86f602fa9c99076d53c926ab0e44797c1448fcf7e57b5be
z40a078d225206465e7a39074b286c0f1e13518390cce8e05d8f6393837d06182d68e327b7a8a7e
z041bc9bfa6d46471923336ab562b1aba9bed85c124841ebb1356a0c34fe7414e1bfa727a874828
z4712d6988e7ed41a7c089be4537534729bb81a11cfd26b4d0c0ca144a33b10cbff7322558e1949
z55f0f2012dadfd52c4e932c4972331f555eb028b42f536e219ac1501ff9ec1d8d722b39bdb2ea8
z6a90d46aa8a41a3dc218f0c680debc7bb2fc31e087c8842de16e77199c444ea927cf239c7f955e
zeb3371bf5d9e60ede2ea10c0696ec5f330fda2a20b4d50168402a8eee12238a822fa8d377f1287
z3ed5f149bdffd61f59584ac72e76a71fc07276177536a6223a016cfa4880b62dcd47c1974e553e
z933a1d0ecfc34b13be7e79a0a79f104abf6f1dac634b57d9b5e2d0b040b4e055cd57888118c6a0
z03d16bdd1ae2bff5a855d4724c6f7891cb2afe3019e21db7454bad8b71d34956ba6cabef727df8
z940850416fda5bf0f84a37852335dfe6eb3217a28f298adc343ead128d37ad382efa53f58ab8d1
z06c7c5c9154f9b9255184e8da5dcd509c5dc3cf858b1bf8ac124ddc6c98b04c5c6056c1f35fe38
zf2c9d9957d6d703363aa55715cf93750b52a87ebee7253e788e7191fb20eaaf28deece283c2d4a
ze12ab0362b19ff0c1fd1abdd0193fac02fb0bd87c3f999e0df5278532281b3fc6a7f5972e7e42a
z00d6fa2de22f5cf784f56db10206c1057a0638ce90c944c084e6dae660aee84b6d43ed0e4e1815
z1023b5e3622493ed97eb1ed9fc5dd381904945e90a7f68f40566c74647b53404320b2c45f29866
zd36862d25a3bfc833e01e8bef2ccf992c0823eae67a8bcdfad23655d7eb57b60c6f3c4daadce52
za2281062beefbdff0a5d8facd8633b6f9f71e7125cfce07d70c3ed2f88a5cf316c26271fa3e1f5
zab2b189420f6c684d2b533d1fd49e63aac3e3eb8089357e04583ea2238b938a46879d9c7c443cb
z8712416948b5d3b18b321c05d842d29bac06b4d29d7fe03274e7e951a562a0260ab431a97e757e
zac72baec9a13586af0f8d5a288ff4af46e0261d945a843cb6fe58ec0f8c5d437e814fc89b513fe
z561cf8bb9e829a3017ffe415335407a2cc44ea9a57eaed38e1187313bebf123a895374cca63fac
z1863763d88db8d26e3de77db49f0421432d1603a7828cf3bbe4ac43cc513e06fac5c94cc3079b8
z6aa1e075845b938bf4a8dcad0324d9752aba83e4cdcc71511b240bb61d6135675ba8d66a0f94c0
z15fdd2bf93d82d832c356f3238eea47e0ad94c5fb4e30651b4ea0d3988e69387cbfea979f8e0df
z9e5686866d75aa09e9b8663c7c79407df0a2fb60177362a5485a0e02a8e2344a6edf59b19b7250
z5f7084dbb5d1a38dd01221a0e6db5a3ccc4e1bf3112ae97f1c2a7e7f6cdbca7c38e19a8b08f415
z3c8e2b95ee4ab06375eb3fca532b580c4ee5940f5cd62b898023538b33ddb264a06bd224fc6ed7
z3fb7a708fd37d09d6506ed4d071114e87bc2c8e4bb7310eb84ec3ec5a2588f3a6cb32cc99c758e
z0f195e99f4b621b3b4ba15fd6962def3d3c6bac25983790ddb21d8af55a5a6e0c6e1f6fdf6c276
z8924150aba0f1fcc5040e842d5fbbd8d87005aeace2d0afab4a6596e48efbbfd472ed32bd79564
z9e7b49411713a7f05a50b221d819153f77f8358c9bf986b6fabba349498a74bb61857359dc3a91
zc9ee62ba8a2f00d7de61c08855801f96b969efb49b64bb6dcbc36f78e6ce28e5a64704e0902f14
z27a9ae4a7d1a80fa803425d385e6cfa7e3b92d70ab9662a7413a3e3d431c56f2f3fcf4dbb098d8
z4d5973c34f0b10561da34168d28a395cf0088f78cbf10b4afa88924949b08dd51a95c9a35269f0
z7686e3a7e0bd24833e2f2d4997c272ab9bae6f3d824f8c5f3cf0585cb3ca2d9f718768ab524c53
zf1a21b3cfb91d521b4d06b4715529328488e57fdc97df65c48ae6663f1906f141f9fd6d3f0f596
z00dd6bf5750f355ac178223b5ff9b039dd4a526c9c12b0eae2d4c9c8592d142997f3805b308d24
z780b40ad158fb3e65bf12a36354145bcacaf380caffa8516fd4dca9fa074317a0310307642822e
z80d8d5bcc5adc0895f8389344309d80a0797cbea8926682850d106db7fff075e03b6c3aa0239a8
z333cc2d21e59fbe8bdd3bcdcd53d6ac5c9561b05550e58d18ef6b1612ef8b69e972fbc334553d6
zcfc3fa92c88fc1aa2b22b3f353d54f90a3d37537758db6739107408d1152f8007f80d62f5bbbdd
z843fc11950717cae0c0fd7fbbeea32e1b6acf0a4304ab0b16fd325d3a896301cd5977ae51348d8
zb904c2dd50fb4aa751e4b923a9d881572449ce02a1029dd99f6b99e830c806435f2f4e30bbecaf
z1ab7a21917759b6a4a3f40f886927bb79b788e33dfb3935df2185e1f748f5f9e192fe40bddafa8
ze1a3c12c19283ff0844e2e3b9ddb0f3798c0121b67157d4005c2c13cb9337e19ce7f323f4e9599
z7e594a5c28e7b83361e044ddf08a1c1981c94933479f9e34f873015f96780c7593acdf0019df71
z07382c555e9c2c45ea4ede113e927b6dbbc742c14697e002f84747a64e86ab2d0d6c694172aec0
z59b3b46c132d3eea00e970bc9ab068522cfa76789a47132b145c3cb6ef71a587052060f0e25d65
z2388253691c55c82ee6d081de5f450444b8d7444de0f19687c5416539c1bedfaee156fab602c3a
z8c42b72e5a1bcda52ac9b998cd3dd222be2ff7d6df19e953606e388d655490545e224e6c1fea90
z513a9fcef1d2c586805d5ac27437b7ce88178567a9b869e8410e998999d6b28aa4f4de30b7e2a1
z47e683714c1b29b618b1de1c5dc9a8599cae4b4142dfc71cee56429c490e9f23d199cd8c75682d
zcde7c5327ed48d34d9ac1e765e7960c9842d8ecc8f440c0dd376b467bea11c4c4a0c9eeed94370
z13298522af9653c57461a1ca3969a78f483af0579512c5ad52db13efbf0b0ecec5b9da66e9510c
z947ed61136a8813b2a8a0d16da95f0685b384d0cf0d297aeea5993924a1fd49d66ce8cffc39b3f
z3a202aa48d8d3ca028ded8354a96c5e626a5cd7941ac0994c22983c5e87eb04335d0517f444fea
z130de6a47796fe78d83bfee870d68f02bc8a3204d491f0f20723b584676904f8325d51840e472b
zcee4f1159e1066fb350b7e854519a2b4a8bf62c02a994c4f60a63c3fc10329330448e7b3aa6ce9
z9c574c36ce743ab3ebfd4d21a54fd2eea1cd8c8379613d6a581c9ac02de86758767268b717f4a9
z598d3b91970a521390978e7bdb75b9f69b028262e9e5a4fb34d97f2bfce7d2b1bc3e55401f124e
z2fd0171bb496e101492e8807e7c92c6a93fad11182972b423818475bea0e140709392086389ae0
zf2bc6085315bf4c25a9d3f5936de207f5eeee4583d7076d2d85ec0b8c9ad676c674af4ea5b9a21
z95c8034f4f6eb2a9becf8fa74a05d509a7e691043b1bf6b2896e956590356362dd9440c24e8b6a
z94a4dbe3db8412eae4e76e8b82f6047080e2afbaf0316f483675f4f4d8d7e0154a5b616193a45c
z42b8698046955683c42a3def37942e7e0bf1578c5c6350972b50148042f39c2161822bc383536c
zc5d0e4fe1af691bc62d3c7d3faf0f25c60499f66b2d32c24859afc1867a3917fc65649c05ad54c
za1622068239b7f017dc3ef7d64c9fb5c70c6b7e5b3d0c9fcb2951b47e0bb3e336cedb23c117183
z6ebbd2a9fd0eb5766c4ce93adbd7ae9f9a4aecaf7e35e341c0f04696256788b217a89b885f7e33
zca23679f9800fa0591fbccbbbb9dd4c06b591567475b975b263ecd338464768eb17fe58f0b398c
z6032efe50bc6a1b035a9a3c2b0f83802d2d555a0461d42e43b5b448db250d720af6dcbb0c975b0
z702b4c9803c41d3c763ca9e2a619937f1ca58cf724f4d5267b9a8fd1066ab0f8df34f96cb68f9a
z42027cfad7855b0cb2440a009db9751435c611a11c3dbe45298bcbc459a5fb6f74c3f2481ae3ec
z6cb2894db4a660cae276f62e8f8e9e67dcc53b6240682bee7fe4430d0567513dff83ab9c74cde3
z2726e94f8e4e79ef1cd27ba0e1da5231d18637798408ca8061e740a4fb6bd76871c50c61a37917
zfe667bc3f5185b23beebb00284aad6ba5350ea1cb0748bb1a6bb815972d1ca7c029103068e1709
z412f665b45352819ee4fbcc2223f6de50efc10af5957ff9a8c611cbaae45fa1c8e01d18d22d529
z2abf2e5143827eb0638659bdc33992a3102b2c18bab70a7023c6845a6064b50e63a65b46dd0f1d
z82aee8bde45598e1717b3e8502f917c912721c334a2aa6a7cc1d334b6f8a7e7b3e0bf4182e597a
zcfa7226a53fe23b8bb86965faed49f7b73f902b20e16b96126cf32626f734f21edc28dc51e8e36
z04a01a7834df0cd26eda0345efe13ce5d202a2ef00aed5e5e3bca209f222c2f40dd84468d3d843
za01773af9a6ab06bc4b93d4f738ae3112b13d5043eb3821bf3e2f7464ac22e5cec86fae9091553
z7ca02c454f962f2b86b223fcc2240893be3d1cca86e418d42f3549a43e8b93c74c61aaf7649177
z17a415de288226914ef85775157d28da1b3ce99e2c05a8fb4812b3d58238878c1103e21f5fcdbd
z0e60afc066a2488f977ee8d9d9ba86b13ec7d779e19edc6ddad359a8d350421c2cc3b9fd9193d0
za65f2bfb7dc559540363e3c9e7c5b8ac776cd2a8c9c4380767756dd39bed11d982aad5e58b6f6e
z920218d06d3d72b87cb949816679b7313f97a87ddf7dc9a90468430a86c188e1e71ecab35ca24c
zeba37a2fd18eefff3286f09bee9eba2adda4543eeb35deb5733034895602ccc9c01dc262d17676
z5aaaacc56602d71a247d72c5a93f07e1b521ed7c0fceb6055f930b493a83a5a6dd2706116dc874
zd47ed239c37ac7af59947bf019a32e68e54786e105bc74c5f7923f6511d65612576e9cd5b47b3a
z8fdf9feccbad17138e1a184e07eb76585a5897e4a994bab3c4b06d894b7d13b8c8e6df939585f1
z9e207ebb9202625a17ac8929522a893a39307cf86042943c232bd435d6144edb54b82f1854c948
zce668c08a37c50c7aec130739f2cd8791d432d867b31f1e44bb038c39bff0780a6983eaaf7bf96
z2819eb7154b30f3e8e4b71a09c61e808afd9538e9f450308116baaacc869ee07559f2b851ebaa3
zab578738fc56be6ad438e6253caabd9090cec98f88ce7d5ee1038fea12133c4cfa55b4ce7ee405
z3d3842db259423e2f04b3c3c65ae5b974dd9d8425c5b77bb339361c93b699ebe64eb9e5abdfaf1
z084ea919a7477f7af9abd211ce8a2530881d1f0d4a4a636414abfe7cf66e43b7f680ccea765081
z9d7663d0bd6168e03c065fd235973d0f6c9e520b86f4be5eb50c23208e75267da5d8358ab3ac82
z5cecca5457dc2ab6e7dd2d02f9c05bb16a396128645b17d2c52362980e00730fa92f142b884ef3
z8102356f231b17922e8ddffa965293f7179729d45625f073597f64782013e0f89e5956eb2f20b1
zd7fc4a84b470d9ad306301c2822816f1df951c15c19e9131ff7c7f6d56b4ba58aa5e854ed949c0
z483b7352acb44a8fb91ce353380fb6e16f7625803a47ccbef852e2a466345f9abad9654c54046b
z9e553875f9a83b0b4dafede21f8be2ba737e2bb20920a93093d0437021ed765fc2e1610d30843e
ze99eac0bf7d5ed26dcb3226232179fa26a196fc7475c8337bde87bd789d31e0b8a6b20a33ca4ee
z8f860281faa541173a056d25a0edbacee5d03f58ab3f67e34ca5435ed0d51352cad46771e7ca73
z30b52f97806bad5c581bf7e18db7a10f346c3daaa6d579ef971893789b9fb20e6cbd7123aacd6d
z4cd6c47ecbaf097a8c9232f979e8071177cec5897c711ec8b0ea203017cfb72d65e4491081a156
z828a9ea940bc042549bac1a79f88ad42b20e004357caf993aa3db4c433ecd09bdd1febcce1044d
z7096312094412925a52521d340e19ecbe5986e20e17722abc2dea9f30cfff3a9d2af6de18257c8
zb73ff14bcbcd36075b12cd57bef7dae4f6757edcfeba7d65ca6dd4e13b4356d24725fe21858bfc
z141d6cfd9fe9be0082be7b7b7f43a3b1f3b383074f5a9e0d2133e6089ac81a79a970b7a61d518a
z452b7bf4d551ebacc2afb0df9595c7008045ce3ead72fc4aa904d7835b37cfaf662e8c57504c73
zce96d652d176fe261af7c90c0028387adc021357fa6c3e81d725c07aebf9443559c943f121f5ba
z70592a1bf0451a7d7e7b57d427d1398524e1f9cdf153729a066db11c7b8d76d8c8078f5fb84e5e
zc705892eca14ab8d5fc0f7efac41557949c568ccfe616d356ec92a89fd2a288ce1e698f18a2343
z77fef5d899daafd956aa1d7ec601e147fffdfad8156b18366e149d7b213019b1d42af38eaeeafc
zf01b96ff10bf3164f081a6fe893ef31e9a7737f381ecf9da6c2819f12510f1934d7180d2ea2b1c
z0e515ff6980e3755e70ddf048befca33f2924a91a9b59b6db945476b6088901e449dcac05740c6
z2795eca511232cf0d740cf9af9ad25e0daa4fa95f138162e8bb73ca5fc45deb70507845e523361
z4b999bbf0e48c9e087678cfe0b5d1f017e765360fa2d0460a451fa4620f79bf47f085826b0b16d
z2f989392184bfafbc27a840cf5dc8eace7f8f4a7f3989eee27d102928bfdfb1666ba6268892c38
z389bff1cfbd6fb0543199bc34d93e842f3383d65f24ea134f264cfd67c363707836fedaff5323f
z06da75b319adde740ff3b1b10fd0e7988d4fa1ea24877cd98cdc32a8b578771e4f867d96a6c164
zd887770b775a9af17815a54c03e7d9d375d85be6eba1ec6400dcc24c8b74fbab40b0bba9343ad8
z00945e6beb3c88ba8dbee8dc47980ce29d433c6bee9b9f05832f7dd57f9da17ac2c1fc89f00b39
ze2343ebcb55ef1c5617ac3dbbdd1df79beae01431c29d882a2056249ea73ddeaf0f78f22caf78f
ze469a0fc59aeb0600e2c7aac59380e92c6f50c9d63f26f1dee44770769302b34db416eee4e1a25
zd2fa5e58cd59da353622117654e8709ecc98592bfe835d4c382b1216719600b2624824cbc03511
zfd02093bfb869030bf2ac09563b43c8d4c40fba82d150677566263c05de7c02c1216709bc391b6
zec8fa4c1fd8fb6b32d7f0811541bafd78d52f776ae136a91d1ce350dcbb1e019ddd08fb89b55f1
zce796bb165a0fc9b84238cb9e9dabdf65d324ef482c81f1afada548e5aa04ab09b833f98ecf3b6
z8c93512130f758dcc939b490556da78255dc415af8425d1058b6270981745112532741387fbb12
z746844f3a330b38ea8e402f0e52f69a7478f6c9a507dea6f5e39037fd46186ff3c8f980032acc0
z8adf6c7b9b1091972b4f93d0c0b4cd366e6af3843fa3699bae50b2eac54779e9c62c724a46597c
z236772d94be9cebe9c802f1fde13eb3b5d3ce070536824385d5fe300896add7ad48003538233f7
ze08c8a88b3ce348aed2621ba358b0b25715bc7895d0d330e77b1e7e71fed9d1afe67e1197874ec
z5dcb77e993b69786e2e53be906b9a662a391fbad4adb646a3b54d55f6c9a63f188152342f0268d
zcaaa64e5f75ac5c1dd11462a030a0c3703999a148a87b4de449747fad35c575ab0a518f8bc2095
z58f27ca28e06712e3da466db822e8b889eaeb3d70789f35904b9b257418d99497e88406c6b240e
ze499299d4e5637ae6398c99a6dcd9b0ee4c11286b13c86d644a063f83b525ccef12f77e859f029
z89f84661c909a2835df559e657ac973f4f7f3091b91cd0455f69d923c67662738f41e49cafedb3
zf1c4c6c2df68af891b86c31a27e629d07c82b1f5e1b14b6b3a772388dc30486aea5a7a3c7d93ed
zb20d9cd18f7c332af4c0787f34c467ae4405248f092fcd4e2b2054c66eab5781ee9a69c002b25f
z5ccc9b742663062390a07cabe26ec0a457370798f0ffa26f3f89a38eef279dd38d2ebb7513596b
z71c0ab1e51f34015ab3eb722b5e3bd13874af2a42e4575fef229c6fbf888b8b3f82efac8bbd439
z56c59322755bedc8d7b4cb7f8596b116b8e20f5fc71a5c6d54e340e9ed3ba2f0d008292af6a832
z8632decb1accaacc7d4367c955a6df37e0920e9dec734cb720954d2b931ee0ba5392cdfa04dbf4
zd24c1a927c22eb9c0fda1b0739d9f1e3456d0267df12ab8179e7c3daa3152246e84795fa7f157d
z17db1cfe83d9dcb9e8d0f90a9851e214270077bd7714b655e0ef27422d67b493c042cf71cb6077
z30ecfceab02b60ff6bd43d4df2b819c8576e4be2e5687da996582b5f0718f7673b1b0d39044b71
z740d4edb718c8923079aa63a17ffe180de369e422a5386587ea43c36a03ae8aedc9d01ece30399
zfc25ab401da0032737b5d7bb3b62b459065e111c0de792ae1bcf45a38cd9c70bd2332ef14d7ad3
z2f7f7a57e38025b7134eeed69f16ae7fe72b0e66c2f1f5b07ee32c8bc84503ac18af92a7b419c3
zf1dfcd7a6fa682fd8e9af41754a4bde0e1e0ad672d20f5712ea01a34e3a55c458d8b3e96bc5d7a
z9e2c04f53894aba1bf5a6d5f33e92b25d9ae32d6286dc78e91c2f129be1d27716bbe6c1b6ac280
z737a042a97b9ac721335f1614b7885cd7ccf146ccc72b420a3f0f362c8cb4baea0938c5e38646e
z692d8f3146081333ea2f3fd8fef90c66148c1fcd64ed39c5829f636cb8c2df432869cf1857c627
z71013de17e7f3f0eff14c9b1b9b9611d03ef24c876e609cb47b47d1e0b4740f1b19431b891442b
z3de6f86a38f57839d44dab77f009379d447e9730a660a49d113fff3dc8c5900bd99442e30b0a20
z9d2329f1305c5a320fa5e4950c41b4ad97824c987e3d1da39afc1e3a1cefad887dbfdf1073ccee
zdc5dfa874c56003be065f5ba02fd3d6daa4b2a57d690b68e3133cab16fafd4a4613c291ed53c2e
zb77c88212a06baad7ec03cffb97dcad0af893900447787b2e8101c01726844e65b8d993c5a9f40
zec5bf14d6cfb50b3d0d4913cf2aeba750727ab5b6c850431ccd7fbd22cf668d60ecd879be5c598
za51f0aadef5bbe74bbfe5a08816726df2d1c7e8532b56dc58acbfc8635eebb47cbef2e38b264e1
zf0a92817dfcbc2bf07528cfec5b46b0d1b1db69b244105b49609040bfccbddfcff6ab3dec5c5c1
z079c756814a20e422a2bab40ba753e2e8dd049851b1c89e4630c0e7bdeeecb1b2153116eb4499a
z441a5315ce7bf4be08eb8a5a0058d730e288ee5ea1bb30745deb9b8a2e3c867358737f6760c152
z427139ffbda69d9ea844ab64f55cc42ad67492c7e52c2b41e797678e5a339f25403247b3a6a1e5
z3f767e2a2fb16f175e1568dbbade6957caf33e5d59873b9d66e2b084f15281b52088170d0a1152
z112c9f19998e78b99ad581da7f4f482da3767a91e75f3448b40fa8ab765ff344535681aa001276
z5fa843519822bfdff5a40064185bcca8eadaca948a326734c42271e77117e20758c9a3bb1f5e61
z7500dd5aeec25ea180ca6cbd43ffb5e1ffcf401540f30a24177f9490565c0aa51ff2444b4d75cd
ze5d36b53d301076c3ced8ebb46de0fb799ef368ffb4bd39df4b38adb823bea46da2dbce123dde8
z22cd14fa091d4da30d2dd5dcbbeb43ddd7f4a1df871990d7302e128a7883bcaf2e6ec794561aaa
z1233a978c0780447100967ee96fb08a172d83fdd79b4517e5b81daa75926426296a04f0ebb0e6c
z4cbe175af0691e73d50a3f2caacc4a26ac4067cbdaa646120a49252e4bba52891ee6a93017e9dc
z6668e572485e29d4a2e264bb8507bd892d9ae237f319c466c40080324583a1d0cc32fcac13901b
z3932a483adfda5ad6902c4b86ed52d90ec5dfdb94ef374c58ddde72aac684154d27b1dac6fdfae
z9681d450b5b15ba0cd4cfdb4ae2c573f12441c769efc8cc6c8e3259b996d4ce8b1c3c1c2acae9b
zefbef6196ff34427677051d2aa2c4222b37d139ad14a3235602b8dbb9ca130fe7abd0d47909911
z6e674a649ce19547263c0000f11d21e9e0e75ecab9bb76aa3765eb6e5cc2805a873766ca09d421
z659b2d5a82e2473c8f7c7ff26612f32e982f64e61e38b8824b4b89a21a527837dd1922585e5eb3
za6bb0dc0cdba961d5da8e20d75e8f073d1eb08bc3a253ed1a534d5b7a83abcac23d4ce667ccd1d
z1092f83abd1ef6e961cc2921d0d121dbb6f44ee07d3b93532ae1721da939bd7eab3f1f54a7bafe
zb8d4d95f8a234aa2c8c4fc01607b3235a1539eb962068f62bdf63f585b36dc26ef31977dd72221
z6019b637bed5618f753a1a1cd627e0addea7e6f59ae507adb744574013e6c7c518dec357ebe495
z3bd96e36766aa11b5dbb63155c2ea639b05dcf78bee9c9e06ff288b384b946d6c6772223a5457f
z25c13ca025a2b0b56c7ff43cfb00fe1ab6331044e5ab76043f23f7b81f00166a8e352fab6bed56
z40f5d33391132c3babadd3913a7a502e4f271e133295b13f57aafaa20bcbd9b5d9d761a5ff9a4c
z24a82810618a0de3972aa1ab89f6b1543f5a710fe6d4e06b53f8930c785383e876cc7df2cc0bdc
zd49789b109b2ebebdc55bea89be4806c062a048c04d9e06ac6483b8e165941dc746f90c5cfe70d
zd72140f6688510a657a7e8d3c458380ad27d40d4b2c41a38487ee4bcd05411810fffc36e86237a
z47e5e91ff81fffe91e42da750a249d02dbca86545367bcf03d1947f700a4ed1a6894d725959349
z829d2f655caf230550126bb3459d1556ac1010d1cf52e848bb912c155e922e2dab3e807dd6843d
za9f50b34b743172e3ccf0bd4d262a093ac7770e6d73ce546de0c7c015e9f1b766281216988be5b
zf8c7f843baa3f0db719e355d8f2025997704439a0c5bdcf5230b5f03cccbeb95db13009cc9c7fa
z6d44f3ee0ddc9c985f05c4ba3581b219583a8e82af368c3d74f3826d276d1999be8b71ada02136
z1954d03a80cf41021c4b99047ece6267622b4f7cab9e730857fd2a6736fa54ebcb5c912cdde837
za6877c96c423ac0fed7c1b91b8d64c2356f5c86b81429f5c409a8837db27fdf2a34d8cf07c6627
z60214eb4c0c465d24fc9cf6010a6f7cbc6859924becc279064f4be240dc57f32116559521a4643
zab95f9bcc4d063ebff1d5459764e3caff0ef2b2607c6fae9fe7860393dda60cea6092fcad2acaf
z53169771cbb4b6decb44bcff91d3fda381949006400224c3b9dc1139bed943b42c63783268e70c
z7550d8569911c0861ecb0a61fe617afd8bd279269d4a09bd02667a1365b610dcb5af4bd479719a
z8e0ef684d6be608059fdef9fb71dd13a49bf7272676297ca85977a0787d71494e58903746e877b
z5ed1ed07b7ee30dd1a42400ae3b2fe004839157e0f941c2ae3c1a11dcc23d8fe9fcb9751e9989f
z0f441c96f570e7643ceca84c3702d347188a503f68872d7d180d7e4c9339ee018216ab3478cf72
z357d9851127bf94faf7322f9570c760341fae853500ba8a685074570d8f632836b3ec82a997853
z9334512925f714522375823347e8899b8738cf5d08d101eb4f9d3e24caf21ad7de1c8ecffc9e90
zf4f3fc2636d0300396654e0b883d7f62f046aa9b6817a39def7da6270832b04924e03300c467eb
z28a0723efaf890499921d1343e00b068142597aaf2ccf2728c5330a87ce1cc8bd3680bffc04e72
zed7af84e738db19164d383b5459a2689f07113cc4c7a78ce73900f07e3d627cb93d7f08d344d65
z2be49209db95789f048e23431126846dccdd665ea7504f4e13329659a170698254c70d686bce6b
z964abca5cfa6e2006b6556ffcd46fed7abf4c70aba5588da5b2d23c0722cc5f0fed9fbf0225638
zc37dadad469e123cd9b67d620bcfc4c0c1e53a36b5edd2965508f98229aef5be89bd10acf91fea
z08425d96db58894a18810ac1368dd31513bf3607d6df501536702d596628d36cbc37cdacb07df3
z869ed2351f38384a5e431b91cab29f8beb3b6d212aa638ac5e2cdb40e96bbc94c086ef2d4fb690
z2052eb4982b00bb47e235382469bc946762e0f7d6c5989bf66bbcfdd0c69a5e74a7ddfd41299a2
z5d69775cbd100a88c7884b23b87f16a7c5e16793a86a526c92c3405edff4c97d0ef4fa5be580a4
z7c8ccf46fb2277182a1bc646e8cdb63f4940f7010b268302970341d1147adee79f64e10eeaebbb
zfe48af594ed41ee3c02576e76d7c88eaee7b99677fb10cbacbe537fe5c17fe215d7ae2a018dffa
za7dee5ca43de156e06c14e971754f8e2487606144039012371f988a6af975eb5a030c94a8abdc5
zfee5e21a09f32deb0f353a7f60cdb71ad128912a1bc8d990753eb19ca4e1c741d6f617cfe3be29
za7b665015dc8b4a5cb074b110cf8947cdc9172e0c60064a121c484592ffac4c6616d0353332eeb
z3f51f0a479c8fb47f1e18510aa931d061102611b7cfed9f0e45761dbbb477ea9d2a91b2bc09e85
zba0a171ba8d62073c47afeb65f190f7b97c1b7df571155ac124ac96d655e3160094e313c3a5197
z7056d21cdfc0dfef9776bad45262cb71960c70b51227704facb4cb7a701c93dab51912f1703988
zfea690cc361992a9d08e2e3a6c6f66c5ef757f94d86566174ef18e9f685eea3a45d70788b81914
z865ffd6ada977e3e3f99436cec5474cd45d5fc210179260a23e8fb7c42b106617164096b0e67dd
z0a17448de4484056a0fc044ba41d730cb2f3e9df4e35ddb8409f8cd45206fa7823070909bd1246
z59709c5154e50d0e564fc596dc879c3a20ce2fe801050e780d8098b273a0083d3b3e7159f16bdb
zb52b6d68ee8d1f0535cb6d4c22192431396903c33d38b72a0fd79797a57d7bdf10df9ab6801eec
z253d8dd35d3b43eb8e5ebd44ef25195341846467f9be587bdc2977a60a2350404fa053eff43e34
z32004d79ef2a41835afee5bfcf2de18583f86002afb55b4d83b563d389c545f5b08a21e29b477d
z42e89e52ac9514795dcad8b4390dcb736945135733bfa8d1abd3be11cf96121497ad43407444ec
zc41b73bc9868fd007d6544ce683e837141c32ceaacf42ae1b7d1468f3d43c0647976e32e5fdb4e
z3d77bb3f85e318b9c972eb7b37b3d91f88c53fc70591fc1f85cee2eb30dde50f89992c98ef3320
zeb118fcfce3d004b9442add0a5af6507ae671576d2b14ca5000331a713b966947d965407fa13bd
z1b2cbcc3f89f21f77904db63ed072c64d2f2b78ee4ff4fa6ef9369656940fd8f6e85001af41593
z9c552f3eb9f683cc2e94080f58fdadefe6df0c8c0ba32a119b93b6bf0dd90839e873a2c9fad69a
z85edbd4f0313d3c359e73578efb1df9c6df83ab6d2fa9ef3680c49d114f341500972c51404d816
z64fab0ff233cd54173e2fc07ec52bd8006ca860148abfae1d144bcbcc6b29a0b84913f74bae39c
z9b137d12201c95eff6ef5ffbc415ee8842d7062c7f69c832ebc562c9714ad3a68faf6077d04f79
z0b5948ca6de0063efd0f484daa15a228bc074a16f9b7438ba4dbbf84b0954be316061461b463ea
za96c62701a61593546a933c765941d63922ca3493a52d55af9e75537ad8da0c0a7ab2b108d8cf4
z384937883c14690db3e5af41c3b33b9ea33a9f21a8a8ead89264960259f967aa447ed8bcc3efc0
z3267c7189eaab68370e2244d14f63240d7f7fc45d61ab632dc291d6663b510017c2f1cd40dc7f6
zb46db985355428ece53f6c2cbe43edec351c2e172103d2b134fdb27d52773debbada30851f30f9
zfe0b89383368b945e677ac7c5a7ae0c9fbcbdfac2989b86b095e00265a61708f1ba42404b10eb8
z53f38e961ad23b3e6d99a2fbe836b884fbdb81c07062f525858bf29d537e56cda622cd41f4e532
z8df11dcf3f9184b1262cfa369ed523bb8141daf650451df83d4ba47795f4ba0ffbc9dea09263ed
zdb1a82e8e2796181032462c96be8d548949acab3c16a21edd4eb5081017bf7a02108419b516ad4
z8119fc70bc9929f48f4ae5c747f432595a10d06d9624b8e7ca00b6239fb6ee1f3ec69f988ecf48
zc5da6c1decdfa786e6b6ca48687eea02bcecd9202da9f2410e2a6b625c749fe42328cc4447c1f4
z4acebb1fb64554432e5047bcda2a2b42f1743e794d625c6f85cba3d51d84a36e9b2166cd54f446
z09364f076f54b45cde3c9fd07c2e8c078b02259f74edda6fb130bf8bc9e90fd477f212b727af3e
zeb25929f75cebecf98572416781714ef328ba9fc8805f80c24e64b53b3f7512077b6951f8f2fd0
z4308e04ceb23b7629aeae820956c7696744a99b0bda21344b9f951ce9fa990375b0c3d0b1497e5
z899baea23973a4bdcb3b1cc87c9d23bab8b7ce5b45774956ace27dd8e135e61a338953b76cc416
zc24f226716b6725691b52f75237e3ab632559df1e3b6023a1dc3f91a617b93eb5f2084dc8a294a
z30cf320c5d7693593b2de4475699b7ad3c828603649b58066237d1b8f8fa086cf6010cf7d93d36
z2eb9460a9a14023708db216685ba99998a750c7d82c0f1f1e4672a89e6b5057894a3ff5a3f6d92
z3ff4a6ec919a2d27b318962f7d6ed157c848cfe831964e098bc550016dd6361b2af5adb3864ae7
zf6da518248dfade465e1cbc1db44211d2497bb7e8b738015154071d4989241dc1c14ca66065b97
z3060d2313824ca85ffea5c7542d9498f174d74bda4474ea598c6a913799a8310069b6c91de6eef
zc5dda06414db18328f768d8598efa825fafffb9f26ea678ac9f2c0fcb8d4dea03f82d041b5f254
z08c0e6c89884bc77d623924d0bcab8e5b51d3be4b2de40d32253a33cbf2ad25dd3f1ab793d58d7
zf1f2ddf2f9ad5f8a937059a3687aa9fac1999b279b2c3d79bca5b9f331f7f293c55f8a5969af7a
zf29cc7a777164623d0670a3ab1f8a8bb78987f4a5b0bf4e942668f41ce6426b893aee9fe943077
z3c88024e26a91698faa2d8bc20809e9221e69254f29c57818075e72133fe769a8efa11e332ee7b
z8edf00269fd2bca3e0b04f18b0a61d1bb7dc8d080a3ab59118cabccc5e8cb957c85126c141564a
z46dfea57788f692edb9d80752f5aa5f5e3115f70e274f9169ed311f3a62f60d0802d8a52998994
z0bc31ee887d965cfbfdc74189ed679fbade87b96c285d5be0605aaf0e13be396bd974d7f633222
zd4053e61010d6914bffe6c56751d3ccca559849023934ab048c65cae92ca5123ac18fdee176af0
z763342460aacc31082a410f7cb21c4ede6f291c0cf7627b1696d02a35d9b0c69e07312d37ff6a1
z2327e8c029eaa840ccd121e9853edb0f94422a561fb6b20f6883cba7d68e33e451adfa8b7ae0e7
z11645dc955291fd7622293300f150e670b436c7ce4593156f2b272f79ad66349d52d255bac5455
ze74107ee881705f34158f3f3b9695dc74794ee5a0395e1cb87d764f367da6e3ddd2ef1d51fab9b
zf6969cdefc7cf479dc414a268fcae769a5a9e4538cf0449a671c150ab5dcea886139a7d5dc9843
ze3f01391d7aeba79a9c87735c14de4d3b42165c39fb5a35a80a5344573f139c9203f22fe4f9a9d
z0546ec08c68d01be18e7a9aa9dd17123ebbe46b08fe6837fcc172f2784a74bcebfc494b79b7eab
zb5e9fc2519dcb43b5befa4431af007a0634a413c6c28f6688a8a3dab119c616fa8d30cd0977398
zf6ff06e6df46061d12e675208028207e570ad1244fdde4b60d5230570ee70f53c1271aee26f61e
zd8bc085ac7577a5672b4bf48ff82371eedb8b1276ed8553136b87dbb8069e33254d994743ae4fc
z499ce749856db75e72544e3c58e375da966bf22bfb143b06ebaabe5cf5ce429759f198642dec0a
zefae649c0877227c35e4e1f27ccd15015f9268fc04adba1c330595e256e03a4850a9aa0d3c5162
z9c0b2d8e424891667bb4876df504447c584e2788887f4270568e39c085241f81d4a91a66d677ee
z95f5c30b6aa2e030de437d339271cef72b0ae69d5facd8515d056e429ab33108d5f4c8ec028c4c
z660f3dd1ec1aa37de49e071f62b66409bb13a1fac187084e6991d6ac52997a39b5d58262a3d6d2
ze6912cabc09c04c059cb0021c2ab6f25b6f25b04263f136bbb3ef3e013802aae98c54495f5e611
zfe775f2b6f04c7f5adb640d7a77ea30c84e968fb91cc520b05d0301f0dfe553e0793e8d34ade48
zfdf3f3d0f59b14049203847c95ff73a25a54a6998cafa4214489e946295b48d2abcfeaef9e5d85
z5376469a91468961b85c301841e8d93ac2462ccc240c5661db7900e31dd054717a78728553308c
z34373aac88cb8370b3929af5cd90d1d8093885bb4e8d748412df2d1e0969a08b8fb01c214eb0b8
z2f2a5c372790e3cd94f110239416f033786f42e3f687b8ccffaa092404a620edbe48b2bb978f05
z47f197066db9dde2a7ee040ffcfb7635f6ff11594ef3dc8c8c9f55fcb23ca0e4983f3e459ee6dd
z15db3c14bfc8ed85848ba4e0c16c0184a7680cad15201be2a1de3e86d3b1f9743a397ba9e6c87c
zfe505b6529b29801a66c73ae1a7925dd594d12bdccd6284594e00c55fda23a2c873b1590784153
zc3df3085246062c4a430897d94d671c7ddabdf252877419578a51085440e2b7d9ed2d7f59467c3
z4a66d480e982dbfd46aab50d9f1b38b43bb9078bf8d005f075190e2877fbcc9e3daca4eb08c2ca
z5081deceb544b7d7fd51f286725c96b46639cde9ef176d412595f3a0dd1ba7c2d8f577a4651100
z6913c6b575d06911e333cd0d72db9f551b3c743df6ad2e2acdfb091912b0cbc7e3a63b2f2e22da
z57332142a443e10d5a0e3c3cdc87600b6dda1b04e2f0558f470d116b262ff2dfb43590e4f3cf03
zd5616c15b7bf7b0f77e62784bfee97d51e03e1dd6bcbd2dd1fc6f71cd6194f4bead320bdc568fb
z2c9237b0008037719b252930b11547497b36a48a74291e29953f8faf0db751f2e2771ad9052a92
zbf0b39ba7e134110b49270f8d090f17ec439141cc5d6ae60af5113669090da37d645ed291b6edf
z64cdee5b2ef912a50113dec66f215c8ea97440e31f3f63ed47364ced70f2ed6a16e17c8d28040a
z7831c4fcf8770294dd072ff0d67f6bcb331795ffa1e95e02cfc7c03ae6b9dc862ec21ee10bd72d
z58da5a7d9da2d03ecf5b83f7b34712c5df0e965b2a74601512067de9874b69d53d56c20eba41f3
z5e69d04622e1f7464c5b6970153e00bf9196c12bf8401a7779c3bdbb7009f3bcdc6f05708c5856
z7e82c963e71ae2cf4b39f7748cd7efca9783039548d2b7b438807782a61e91f961105ff09fe74c
z7b502fc7294b62cf6321ce4e30572be68da687e18d9ec2baf018e7861fd3c64e2da38c876ea399
z6687cdc39abf9e5764d9a3e547ec141fcab5d2a6aba62827c33cbcd38a2f4bd0ea53972ac14df5
zeab9cf8d90c888d549131347fbc7b03dd4429ceafdd5af4283d82d3e3e0311a00ffaf8986e297e
z0e3a84d89bffb9b951829d383243433a1f34087db07642c474c80bde1bc24f3023f69c4c000b00
z1a0f341e734adc881c5cb7f7b1ebf867550e798afb0d57b6661ab7e53a4a5bb10c5caf5be38ac2
z8e25d315783fb4b57acfe44932b6660bf29861ab0a7fdc2f8de5288a0ca95e73b082d34d4dba72
z50cedcabf8910789326944e43635565df254b2644e11b99ef9fdddab3bb5b916d3866e6c991a73
zb0b72de214cd7a609b3511db278071337262fdcb452839bb31bf069676b611de0c5e981b73fd88
ze9083bd8f6f6c48e3dc1ec4346f3d1e4472573d13c8c61f68c1e8e4ac0ac5b743308e11bb2a59d
z5d2cbff54f5554585daae56582c638d83e373a2625aca9e0fbc7a0148a3e9da197cc3ee92b9f62
z28d965d25d61bb1ce74e91eac07a28ed207d117d1a146910707184ad07c5a60a450cc36fa2d2bf
z687eab3ce73e99f14270692b8587b632b1b64bd0c5a64157327a8242342eec71fa9ac6aa5fac50
zc05321ba4dba6059469955603fd31d97bec9c95ae821bd7b0f5b609b40d4ee4cfa586adf375c80
z1d1652124d26bc9b4d27b85f3b874aec4ee9f6ad7ec91585a098bab194c6a9f3aafd214209f553
za679d99c6fa11739e2c8231e7c9286bc884df0e42f44154e53d62cf85da8d0a67e782303122d95
zb6225d06d40ffd000044a45d4015e3bf317cbc0e63492b8f9f2bd0e6774292510e31d9838272dd
z56d3af383e96fb03b1c82d89031f7c5a531904f6f60eebc11cc5fd447e83b813a6493c11680885
zbd1af7b5bc6cba6368ac324f544e8dd5e2fdd6a9145e8ce558f45378a239b9e2bb5139c190c28b
z5deecdf89f986b5b0e000c608756109e86c22f44a2e0bc22e33a6b347a5ab76ae77774e77b66de
ze6eb63f7a458c167bf0b960bfd6606c09abb67428897f856fd8e67372d34e5bb7e144a8510c229
zc06dd80e752b84726b84891a1183ff18e7376285ef8c7569a8961b41dee5c76257d9c6beaaf822
ze33c51641f489d4e800f26e54ac4a3b39fbd3bc1fc68187c80c1d89cd98bd723de7b45475236cb
z36ea9607abb71e4633756351142f22c3c0c413ece11b3aa6c834dde2e1144ffb9b2e029382e67b
z1bce9fa8251a3a5a726dec95744c0ca9f0335c24d8cf8ce65f7016523c9656a8be75ffada6a01c
zc84a384c026a43d7c60feef0e4fb94623a6588c5dc531c61d09988e44d59180f6bcd1bc5dfd526
zadda732a9494da9f831e6d61d46c6747342a96180f25bc771744d91368659e52a2929db81e5512
z044544819b2d3b4d571f6a3f9cdc37bfe646c8d3cf2dc2a290c47777ae7d07f2c63c4596dcfd9d
z7bd2f821089bfaaba0db2d2ce399cbd70739617761beaeb6f617690dc6afb0fb0a5eccaed2b5ec
ze4f7f6e1490344f2cd88c41d641ca96b3a9f667fa750a142d3a62452bc8096d28036e8d3b92fb8
zb7d0ef6140925b3d3ce47a4b388b2c3cfba72ff6f686f9c1a4d9710fc5ea0c0facf328ee152443
z6ae05b33d7d3a60e6cc91f4dc43bed3aea85aa3df66d7305642fedced7ab7dffd0a1189181298e
z2b4525f065a00363d519ded443225863e02970de3616bb93408df8a68d713ee5784280625ba792
z69d718d8e164903a01a635bf684de945418dfc6152ca191b47da4da2a66314e8d7567f40d04db0
z9bf9001788c75e8dff1594b6414c42a998df1bdaef53a2e7c20d3bc86458ac862ca1d9fe95e85e
z421fc62c16a1e699f4cd34a500f4793d43b828febbea146c6bd62dfebc2a74a109d9bcc7c8ac60
zfa65298171c4075568ae2b69c7ef547fe74681aaf16750fd3890a9e6a197c49cf5d75f1d6b5afc
ze82a3c51eba519a96e5aa7a43de5788285aa7f0c32ca6fb9c94ddd22cf234e8df9f2287141a17b
z9a667dc4f824dd3805b5b66eb2280355096792650f07d97db91b6d254e3a41d97a576f2ae0ead2
z6c6f804cede52912cc11a3be826e7134fffd26fbff4f419c09042acd33445fff9f08de8531552e
z233cb383a07089dd5b67a59e48bbe0e5852b9171631d3ce5e1a0cb305e3757af05fd66a77b14ca
z90f8dc8c1f7ed80a43ccd38d5e4271f61802a48ee16d156b11e4bda5c00b81fb5893732887f437
zd17e50c900f180cd7aee8d786b1185e49c7f736973ee272dd6c783d432abbe1687b1e88cecd673
z14a088b5ecb77e622f6821c4c2ef52aae08999f63a78ebf693ed1159eab091324baf076951e14f
z2768bcb3cbf8397d5959a70b0f0d0c96aac6466f52a3e0ff6041e2a95e386404b5badb6b5c5dc8
z1d354a188d199d197ee492ac2808fd7535e837bd1a79ba27d359fe78cc34d215aff8443c808e46
z156b06615dbe40e0b97c3e5e0607c969897f6194c61efb3394f63effd31337dfa378aac186bed6
z07cf0ce0d7835936c891399e03dbcc52cd0d03bb5980b38c697c54808d8a4f41fd3fc9d7fa4c98
zc5726498aa1c80874cd1a3559103e6032ea3cb042d149c48aeeca36cf50fe7e652d13e368bb720
zc433e8024d92c1aa6ed1264bdf2aa52f1cddd98bdef61d8e03ae21385cee84883c2c1c46daf53e
z89e3e16943d41006b18c2b0651f7309ee89ce4408eab7bd766ff992d46733ec5b7645a0b958066
zd55a235327caeb334270fac154fd4f146366f15292378d667d614fb1cc7bdcf902e1bfa0b28c06
z678f6a572300f381c858cda37c2f4835cd03bef0e27760233ce80e6729f68fa004490a90e75b60
z1a863dcf135e3ca7bab46469be1acc40a90946c5a02a873b8826f8ec83350131fad63246e0b5ea
ze67ecf034e6d91637a79228872f49190e3e47d6015a20042fcd46d26fbeee28b88147c6de64611
z56b661fb049c473b556d7969de3ac492ff33c97ef57b99b93f61ad1ff5ec2eb1d0bca1314b2aa7
z3d0fb93276a96f058b3460c30d392317dff22eefcff85d60af66341fb48f400a6e751d31d86746
z4f549259f52a364e4bf444aa183bf79fdd3698f6c83bb93ea179f6d63d672782c4308aed01f550
z250a15a96485df30c09437a3564a568b1e0bc0811341657a08e94a48dd14c37bc4ca2c3ad58ca6
z4ddef005c5f3a0f17c5c7913f1fbf192a3b46c8d54bc1340910c9f7b20160345f9ca47b8e0914a
z5f9a7a88f98aa3303f52ff2d9a87e73c7a34b64985b51c337e7603015b9b2ce5e2fdde83f3c61b
z61d00426e7868f9a52d85ff0ff0bddbb79452ad75358d0d529459c4d4b9cdd38509e119bf1a00b
zf83a16428457783dfcd6bbbbff9d12b8a33c7acc9a862d786244a275c6548c278347c2befed9f9
zc56c247b01c6d861c963020d95d785bc88be278ac2b3de41b9430cf16b13a2eb5adfe2ad612d4f
z273b43d2425d414d83e85b4393d44d620cbf4b71e8f27423ad71b982bfbf0f4a2f0efddb4a8678
zc26d72ed5d517df340f17d4bd695b9f9ceb7c03bd221506c30086148bf3aa0d07c590015af1731
z5379ba8bd908af58f84a5c0efb4ecca7ca4c83a1fec9a7e80535d9c5d6d1220fb661cbc863d943
z9b5f7618d6b08d04f9fca26f33373e911c1b02baa74d598041ba8a49b4bd777a99cda53d97c4af
z24688da3a863cb181754a27921bf6508becd955e097360e668772293c13b0f781e5e4695078a3d
zfeddaa3ac7b2812fbc3dc58d2485404a6037031f8155b0d0060f0460f959615de151da493b367f
z07727b2a68b53dd9bbc795a63a67a048f0001b3ed9eeaea5167f8df33fa7f6a06b40e2ef5abf62
z169e2b2012672b0beb07241042d404fcd083c8550140836b296025988c40f52a0cf59bc3a65ced
z8e06c87d584802e690899cfbdfa3651448772b2244aa3b160388b0d37b81545776a45aba0fea38
z5179525735a35f55748dcc4ea3e945aaa2cfd2ce53838af7957a990e8a2944d16c90ab4288c617
zdb61cf3deb8e86e708da04ea4a1bae045f6484c988e579015477a30d9d8696253a9718e06a31ad
z0cf4b968269f843f4f2e82980fb08832b4ed84e4dc57a52be143e5712443526682805a695c3b55
z0bce14fdfddef12e08a201e6cca896df151f348cf2db8e80303a7a81735534e82655fd73333948
z6c0f0abe707ee7a0c105baeaee8e17e61c0bfee51e13153a8c5e36935421347df37e47194fa75d
zf6caae43e10b6db973316688091b99612eb2e7fb7a780a190b20e31f617c2c3dd4036acb7c4f4c
z11d7e4beeefa3d11d06afc6c3c978ca704ddecd26d907d8c2b2abec9cd571d1e8e7efe5a254410
z58fa1eca3e4fc8eea385fc243a6623b0d6099c935d4ac05eeab35cf1715156c46355eb94514422
z486c4b830b20ec2754ecbba071387002135a81058a480a4a59c344591ab2ae60cc0ef93d1427e6
zf1cbb96acac610b465c5607431c91464e2c875ce2f39fec7a749699af55ef6872fbc8462dc3463
zae0e29155d8bd3eaef1ea13e66b1d3052c5b314edee3e10567d2ab21b0559977a5381c55adc25e
zef95dd6fed97aa2a3bcc13aaa89d06d5aa6579eb3e28a6c747e682f7378ac93f843a56265ad6ed
z205b7622208746c79508dc71de7be80284b86ec2ab4b940006dfd2fa936f63a8ff802374a844f8
z9017886c4a9c9f0d4989e3dbf06c8cc73f229979f6c4969ba0b0b8cc760f017ef19cb77c42a046
z41ee2797f0a53d162af61b889ee46e964b2169b47bfbd28d970f7eb4c36e0eef7bb1c3893b29bd
z2bd26b95c168f18c08cb6815198bc32b5858f89d16a7e1da1d0bbae873264d596356b115bdfac3
zc76770298725ea7cd5f80175fbd34cd8de16a1a7ba39029eb9f30fc765d7da181332f5514e4f99
zba6133547adf773dbdd2fdb1f8bdb32f0a7f95c0a6303be43b13e55a5ef7dd6fbcb16ae9f77995
z02fcea295d404498320aa4feebc721ac35a24cdfab0b10ebc45bc45fcfc70ccaa29e6ac8a2be46
z1813fd4c244a68e81144479242e137fe88346ded2f5c9fe74c1483adc3913bead82b8357a69cd6
zc215e89191202c1a720de9cee390dc931184f4db12ffdd5329dbe4bc0dee842fe75d94c00b2830
z35a07b1f17cc8f5cbed97a3c58f57bd58e785e2fdaa725238eb2728c5867aae1d62bd2eed97586
zcddb4cb8cab4e4b7c36e173444fd0fc188eba40d9b6da41c85fc64e61fc6ba02d2b110caf37d1f
zbcf85cf53a96bb1e8833b4a4f61a6bccd5d8e79c2dfc04e2af5a81774dbbad9323b588437b120c
z492cf9a4607152d92d764323ba41d767bbb997e23fd3437106041315b5af2b323138e56f839536
zcc36065e1ff345ba63d6c8a8055390a10dd7c8cf354946c88a9a287c15d925bc72ea6a3962eaff
z2ec88f923b2c7de81533c9085ec0c56289b9cd219f85d002fc783b7812765f8b4eb4927c8f3ab6
z5763cfd2c59ded4ae5d9272d274d35f79665210222d12fa8c4a14274ca2e5df34c27e83df6e049
z60757eff27be636b5290e2e3b0bfb4fa997adb7de9b300e236217b428492a1f8df918dcb199580
z051b326c9623a7e6c9b63b4eab487a382868454ff7b41d21089558de1f4a0137fea83d571562f0
zb19269fbd68b19501907bcb313f42758cda9a3d388125741028ea6508e056695d1149d368ad9a1
z23762301d7923929981dd0facc23d104cc82dfb4404d1ec14f5063eac0d88f2f5582af5981cf01
z13e790e27e174bff76b9c31a2e56e0aad54f5f18a73315637cd47863641cf8025da4c90b01686c
z37174f7a485f3e1294833f5c4237b38d6493e2aeff03c237cccc7bc927f23c5cc03baf4fd03db5
zdc913e6dda2867343ee8ea5d03078f437918d0a6b1a06413769be888bb2278855b534543d36b18
z2a5d0f31fe687aee8e932d367766f6b72335e356e1ebcd89e60b839a6369621f63819f8ff650f7
z12234f2a37e0105d15de4902472ba566e68c0cd8c93812475cebee0141d7c4827d4bd1a35dec3e
zf36617700478f43ed13a075b5a2ff8760d07a002e24ecf489c50a1abba1b34d08cf138774f7e80
z4cd557e7f69a1005dffb12bf8e28c4da45c17f4633392769b73a41412bf1022cbe1f9d735197d6
z630e1c53a25dfc1d50751406b8ac0737a1b0119a3a31e6fec7dabd8414ce179a631a8e1957ae09
z88e1e61b1f87d9444b0d50efb7ef5b92724dee3cd879f5522f2c3c233a027e7996296f88ebeef4
z7747b3c3f265a96be7f4e0e5a2f3491707a7009e7ba65960c46634e6a6f16c4470cf7674643b77
zf1c57f80c113212917d8715f2dd1bf712cef8e2360f170734f59042fc0a2d29f6d463303798349
z28247d67ffe1e54bf69c08e5f0fd9473881e92f9d752ae4a885b8135fbb3c49fb0c541078a9eb6
z0e53e892956f81a71a3e4dae00d6a09c2aac023df298ddb671b99726850b6284b85905a922a74a
zef23856ba68893ad5b308cb68d851b9a3a9472a8e5ce7bf8d493aae38dab2f6e21e3d708b9d29a
z327b69414eba7ac22dff2f3da025e0f072ba9a335f189828572315818976fec91a02ab6e2226f0
z6f2cd195289e2a442ff44bc108ccd854c2770b8d41f95ed0d3d3c60919387be93e83133cdb27b2
zf6d5fc472d63fec7341ce04550564543a21d0ac9abc4be765cd09e46ffd90af2a364d879b6faec
z172dd55f5f8f4cbff388d86b73e7a995143d9e95f857095d48a2233bf9f58942bf08d3659760c8
z9db6d8b98b7699ba83bb00092144db2f58944f7c201158d42a03e2be62bc22efb7ac1faf8dace6
z77ffb847c0418402747524bf8517b0859bbc000a9965d6914d5f3fe0443d0b7cfeb50967ec1c02
z90af8e296489b0d31502fd2fc17c2255fadb582710c9305cc0db54bec45f73b1897980b2e1d1cb
z2ddceaf70c6f42d7668770e794b65e0f3ffcb1b5a8e18e9f9b22834c8ef9ab89f4ecd939a16057
z7b1c07a8cf9b46588936d92b45a914b75e3eba3cd3b16ce6778d872554bc73841792933ab70119
z3f2730b2e9740f389d342b3f0380cbf8b6442b13bc6c0c875c6da7a7f5ae8acd6cfaee5acfc149
z01a13852520072d1e56385f7a58b6c236762266e47b3f6e0db1d610b6a1974c45614396ff69c4f
z36d784774f83ebf20ffd8b084530e9f7dba2a61251da5e35356ca2628e72f23996b960094cfca2
zfa1de02fdc613c43a78735e8c235b1491dc06d57b929735d59f49d1503999acb50ddbf7310e57d
zb40a80658386bc18e64de88fce2245b0509f260e1c7bee5cb71876dfb82f483967af2ec9844ddd
z280d0125d5ade12ff7d38e4504839c0028ad8fbae6a3775a6b466dd6bc50f42a9913f54fb75ecf
z63b619546ab2ea05b88bbc618f03786ca26606ee62d58f28f6768d6cc2327e5daf899993ce535a
zdda527ee981bbc28364f8c96854b495a999dc2075ef7c9b2a584c04bc59c928f690589a7c3b58b
zd6c550630d4426d33f969348062c6eb2018e56424dbd40d04ecea16f0d23ac502a3947b3d208cc
z6d3c7cab5a36671d5089f4b858dcba5634a7797ea205b1066530b6a61b5d693555fd619dcbcaf8
zf1a059c54900cc0aabdcf673563974ecf7bf3ec37efeca880b839aa9fd5a055a6c50c36080defa
zabebb8651afca1abea57bc539111470f76c465078a5b7e6f75328d4f1dc263c26fc9ae16af84d2
z4d963e3f832a3677966f5c03a2d2fcaea8f60143175344f8bc54eb8b79c610c597e4095c3f977d
z0942c2e53d81ef35aab9cf5877c9bae8246156ff7c8b3d44db4dcaf9109d5e450c31d575bf50ca
z170c3dbb047e7ff9b34515e075dec2efb3a3d85cd99d71018d198f5d1026aa2df26c5f930031b5
zfcf9e30512a579e733afc53b620f613d8a3c0a31a6a67b1d33d422deaefc7ff983298b454e1fec
zf6a9e9c62ac9c1949f526a5daec1d313a0c1257813a6f04fd161afdd8539867b75b4e493778bb0
z351c182a034564042917add4afe4661560dd3ff873dc0a5acc3ff600ed8f6270ab03b62d6f9cf0
z67c43dc70baf33c32909ee7cdd34aa7df6d3ef3ecb31f0d71753d073ab84667f49709df7bed478
z8ab6e37d05c62154bb757725f2e4565e39cb05997a3d87cac451a987c3265023754ba769c95d4d
zd00b23b048b68f203bb6eab37dbc02fcbcf9ca99a953fee2cd6343a9f836fa8ac9c1b36a1f0b29
zdf88097fa8495061655fd27cc494a914ded2d1320cbbcb711742b96e56dff8a709731b40229dbf
zb4cd37e020cec0d07dc0123c39a9756a128b847d660b161dea64215a9e91f54f7ad2e5a18df2ce
zd8402b0fd231a139187d2174bb85ce2793ae2e768d2af4c6c610ec0dd0e5f2e0d3a3b5f74803b9
z10a9099ea1c1571fd1dfd3fe2e73036f6c4326bdbbb1788aebf564441b94dab789ec94b85b0979
zd1d688ec574c2ed55478f23ac6aeb39e947789d0be82bdff1208593297418fdd7949529326fdc2
zeda02bad1b937de37fddd8eace174d5c0f4b1bafd2af0cd429801e7bbe3cb0d511058354cdd070
zca24add2e1506bf2a77d8a0edaea21e6a9c0d89e801ba997ee2ceaae3391ab4c59cbd7fb328c0e
zcb32c3c19ca944db0f2abfe63390a71e950e16814dc3b3bd002cf295b926f7f8e278189e408c29
zabb22528e5ed3e04ed35df82691f9be71a39a7c0d94775d26978cf6af0dfac055d5bd4de3206ed
z8106e706acb7f9d574cdedb5a79e1b07cb203d3acac00923f48fb49df28c8571a7ed28f2b0bbc9
z90a954202fd89ca35bad9a3f055fd47fac15f6154ec7bccbbbec641fda7e424445c2c31c94a140
z2261f521c8e964c539f555594c919227169f2d43f60d2242082472d61b26ace647d9ce308b7c9f
zc7ed4a9d781deb1b30abebad5a45286a1beab2fdb76e7a9805b5f06ccd9ee695d57d184b51b8ed
z7c0d4aa2d0c47a4d2507fd8c62dd1a794b03ecc3b2140b5fa487abf92ede98de035d9c1f6c0486
za0a796cae99e60a6c13aeb3420cee186ff1bd30038061e5d40b6af27591cf30a6e06d7371d573b
z040bb53c8e046cb4699b8d0ef278388a3933db8e1f7544c4b12f25194e717ab1a6dc98554d762c
zee2e25b9cbf220550cc38492d169d383e4dff782f3b2a7f4dd2c71d37dccc793df29fe22072a97
za218b2bb679be9ebe52d24a77da0685ec9ed3bc4976ef5b4196c3f26db5800c944401b905665eb
zedc183053b5670902c9a7ac934ac82682aeebd4ec301503d435a541fce504863d17363dba28c8f
z0b87896b942cad036447937e26444d90c7c619fd4349d3fc261368e6b0d2fb5bd3406f9ab5d6b4
zb91dbe90f60e8696406a61833af358ef55e2995b0c79924cdbeb8263a383294ddbbcf1c55ce390
z3d6bb86e15809a41ec060d893457b1e121281bf2cb6d2ddf7a88877878423e4282b71a9d8e9100
za48290bb05b12af0b3514e0c685430ac79c42da94831607ae75436ab16161653d7a84dabf9fdb3
z1fcb376430619c603c65e078554c5ea9d7a1af35b64a110d090ecda590845b2ecc3eb205de513b
zf07e61d75ca416c8bc922978b4a35c16bd06bb0eccce5e2bcf43f8af211eeb95cbff22311d6978
z8889a7938b8626a0a98959a1ea892e578455c520e3018158fa9cadd9b895f25f38d6b050dcbbc2
z81614838c8f19f877f9987cec3b8e7f5d987d8602605960d1afc6fbd6c653acb12db9fc8c32f6f
z81dec5ed6d48238fb86f2337cce1df1180a449c765ee32362dce48dd2aff4bf08123fd1daddd73
z4e0764700258f284ea5bc719e429e18f89b660f1c0e45ea16cfb3f83cc5f6aa7d094f727dfdcfe
zac29e9a9c74e073923197220cac0055d7f7d1451973146dba8c79db11c2722bd5ee62ebc5a4ebe
zf1a7879a7659ffbf410dee36679337bff08f4b8b73b77b4618ae738959db3d1914120f998bb0b8
z68ae89432ee579b927e80af411bd8d5543ec42ee917ce37be2169264279536ddfd66ead9a56b89
z35f08e4c8e9cf658fb7898727584246f688796b5577c36dce180aa2dd6ff9e47057ae980155855
z51954544af22775104d0be4b98f3493b7905a169e9befd092a12eae1025e194f4f4914f9426bf7
z8de12646d604046e712c985df07adc18fff50c868a9bd005039254e2e804d61d72c2f7cee0bb38
z56d214c0a538541198758af06dca17a6e2b693318aabda13dc7cb582f03a3db7427b7511c5efad
zf526567258748a501d1497bf480ae88cebd55a8a7ea8cf8606b1e2ca291fd7215cca13398407f1
zc7840df88f0306f52a009691f31cc5346a81bb70190e42f4add485593c8da76ec2c0341f64bbe3
z02e2f5d871b34193deaac99ac481e2a8f727d443bc137573634accb467b47319effdf76dfcb4d7
z35b43c3825972db33d0ee8ae23cb89488e2c7b75fbb58df740c10f6f3d65047f60897c0a097773
z53fe0b23b81974be52a00a20058a1471cf51b5b3165fe17037c51cb2b53497e8e3038e0e665d01
z4d676dca30de7a946c871144ef878b01f62ab4c25b2fe202d20600719ec9f998dfa9a176970ca6
zf4433cf58e4e9cb1d989d777eb9a2655c57631d385f15ce134a56c2638af7be367f9fe97e3739a
z0d6200b65ab1a91549886fc56337fd5c1eb1c2cce2672194632f95857481239010322d48017536
z0561fb16c6c7e488ce03fb7f233e1cfb8e51df29b8adcc3355c55297c731456572e7220aac286f
z77e1fd30231b435f7c33f5117ee78f77ede951018e6ee64f1ebe72d769f8f0a20ed6128d7af986
zfd738266aab3ff50bd8fea90e8cca266e6e2a858bfeabb29fde276869d5ec0d1e1723cf6871213
z921751f5312e2d4871048b28468997e95387deab7814e153e01ab21e15eb36ed2ad7bebf339e46
z3d92a124a7abd781f9e1bbc830d6e6a7909a7f6963ef45fa8afbb12a5d1824959701c17dbcbfa2
zaa29b1301b79c1ed43b99b13ca8466d1588d032e0a062218519da347aa0820a35f79a07df397d0
z50545829c9090503f215a36f1acbb34a44b05db795b7db52464bf6f0d8b497714529cd99e2b2a8
zc7cea02fe3fdfac5ce75199276dc36d22b55635b2342304a051a14403cd6c5a5ed2dfafb889f64
zfc8263164aa60ca9890e6988ed71e9ea08022ddfe91d1e8678a6d35f87836573339f2ae3f6c390
zb1a580a1f84f57f30856c709c65097962b9e90ccb53b72949779856238db4b32bb06e729542053
z1e840c6d029390d3ea658325ab463101711bd12273377dfe4e8f6a0dc54911d70ad6d750f80132
z1fc60dea6c75369efa3ae439ca58e84384eeba3912e0f5d645c6c55cfb548ede3bfbf125d7149f
z37550a232b95fca4e9e6f248fe8dfdf0100e1d009f271259233c5234d34403ca63740e029b3705
z90227afacfeebf6052a2cf6ebd7ca3ca2d8608992480ed9c9dd5932a764b91b4f4146cf5660374
z5e69b02e08cabb86d4deeec6dcae66ff289b6c549ec6492bd676c3dbaa2204254880b8f6fa42ca
zc6cb7f2b22e2cdb6fee4230c0ebd09c71d1c3a82e8b32ceb3b158feb79e5ce2f5764bf2c9add7b
zc827a786afbcaa62664d8a76d32923dbba0bc8130ca435a99e325f652634408a8459a487aaa72a
z4e765e21ffd740f11d2c16f21d37dd4ef8ba98234d2d80a4e446f71db819e1c165b2b5e3d60b89
z61e50afd57f5f78310a674a22058a46a55941648d8ebef8b5ae3b0e17e8d87ed3a842dd97a997e
zf4e1e3145600c1d9c26844ce78ed20250bcfd996b8b427d885ffe9bae9fff2831c7452ea275783
zf3fb2da32a5b5f9dee643247152cfdba3087088d56c8da08fa2ec0ce68129805cc551cb17fee50
z90c0f5eadb99b775880c8083cd76be618010a320353f082423d9d9a87697f5424a001c555a9af6
zff68ee6b0891ef3d1660141fdcf9abd0dca86ade9739bb42675cae55e76f740847fa58e9b104b9
ze46ce2d97a9f890f3d529b9a2f6caaf721354485469f047ee7ca9b14c0ab84f3f33826ef9be07c
z60148330dd78f0a47b76c5d6b6bfb15f473963e07ed519f404c1f064d202dcb420e853bf5ebca6
zd0aeea804766eae4661675d01097de6adba5cfbbefdc4e341f8605c0bd3f1132f7f6593d4346f9
z48b29b09a8ecaeef170adf06801b6f449883322c35b3dbca9ff0d5cd7135216e2846412e64cbda
z2e961e6b1c564c2cdd5ae15daec9613888083a41e5b80b7b819207aefe5299fe4a2ee33c4af153
z72dfb17ff040cb601d2cc785dfa08a064fa2641f151b1e6c37dc17e0cdd5333b6ba9e7dbad1ecc
ze78baddc1ffcf024e5549c9e5b31cd139e986dd4d19f37fe8a62d4e84f8d5e7c504d6eb99b3ba3
zc9bd4bbd51a85b3f0dd052b1a8e9d7dd5609e39502e7dbdd55ace3e2314a3de966c94ebe7c9ba5
z2bddb90e630762974922dccf3ed9bd665896dac698e89360bab54e11a468736dc63408607b784b
z1592bc2d21218ed1905b44ebee2d881a030515c5a8642d30961ee8e712937d9344f0ec2d41e92b
z98b9b90f36aba8b21e473e9b26c5b26ea85752318cb3a385cbf93f4974a01fcd9220135a1ba226
z0acd54c7e554cefd5ff961553ff73e52c095dc4624d329c727aca97c18df38d5d05bca229315f9
z5eb2d682eef5e9cef54d38cdf2edf67f42595a1a6dc223d216c6f942db03dc94bf8f59f905b983
z3c73737301bafd2b614c7b29b0bff25482f80703c1742e4091d5d6c9ce4db6683114de6a6c973b
z4a15ab8e26a6693c8699df10f78e4a33cad895f6391a04640150d86e55b2ae48a94df67db0d572
zc54bf5ccc82de1d723ee8a5c57346110ac84751db57927ff60517690173e17a52c667c0e062ef0
z5c7b9713ea12e460fb0bdb9b1e50d22f3394c0bbc4a0541df722e86c6f124df6f9d098c8611091
z3ea57454bd4c51cd3d4f1447a32fb2f635a13035d3bee81f1159a6a49ebcfcaae39c23f94526e3
z66eba4b2daf2fb3b7e3e8d94d1eec3b49e2395b1b9f29a87c0590ac832f81635a0ffda07be1461
zb527da9a0c9e550961a79f4c623ee5320be68bcb5f6e7b920812cb44cf64983e217cc0a7abadb5
z3297f02d0b602e7e4b4e6bc60d66df37e890091b2ffc2a8afc878724643b420e7712e010d08473
z878f218525db752e4fc0f3427c666c532dc3885003596a0bb202809e642555c310d3c765b94ec5
z58319f315392d34509c79dd45df84181b1f7a0e77a043a7c17b86760ac4b0b07c311afd7a79172
z879ef4f47de594ffe84f9fca5bf9f491b8c98dc2e352a83d15b4684a3c93ade6b3c89f56349440
z88f06d2e263aad3db206172762fdd1369dfc34e967dbff9cc89d36312a08ca223613e36a77168d
z0ab9ae4f848d1a8e47f14f8e822ffd91af5fa6448b9847dbf00434b299b9791e47376b25ea2a6d
z22e059e4b5bb6ca6d3daa6ac2d2f0b9c74d081cd02b68c7fede62a3599a5fd5f7302a8721c8d7c
z502adbd374b30b65601e7b4bc603af11cd28fe0bebbb3eb070eec2b1583ac38b9816485c42e286
ze17b3db1dc3bae383627b36284fa244e8895738656a7d197a482050d960a3331121e65a6e0cff9
z0f963cd6065b16da7aa5e3d6d4bce85eb26a217bf005cacb4874c81a115a6cb099910869465f1d
z0d196e581f36597614784c8a4f2498bda3f8820a6b44dbba2292f21fe4bd750ca23624ff4d9512
zb7d031bb119ddec9bd94a3121da2f60e5695833ce0e9488ded6db5c1ca3b3d1d714ce8722b0c37
za01f26773e0c3140b51eb44de0336f9c3da5ae204478a24369631b65672494e2b91fee4fb9a46a
zc9789a2ac9141ba12d451b475474a7f8a9e11fb07afe2edf810c74273bb14f4300259fc849d5d3
zbcf8f070433af0c93218a1dcf1cda1885ecaf5790049985dfeb98082110a2f4279fcf5278dfc27
zfcc825e5172a876438d824d10ab7fd5c5f7c5a653376938a2ce103a8de738ecdfd93bb95f0cb00
z15130ba800fe23181be87f9f287925a6c950e93e7a225a52428b9f96243ab81666e5781951a6c7
z56f1fa424a7364c3f1a8933c693511594a18db77370b5a90c44c933b4a1a97fca50c04f57158b7
z9fe5f8c76806d4b716216a5a4adf4e969ed1a98cbf1f2d12065a65380ef64cecdd5f43c3f4d2dd
z2b6ad4edaadd38097a0a80d28ea2505722f172f9e2b7490410aaea66c35963e628ab881a9c2053
z7a3cf1e2072f3b3876f233ef11119697ef480ac851f1dad8b8e4cf8f4dcd32be3a761943529418
zdc5fe2c7394bb306df273ad3fc4427c86a1b14872628e1200dcaa3ec93b51161172a50ececd446
ze46e31a79797b2db0c994802bed07595d3be300f85c143dfffc3c4eb5ad77000e170595d5b748c
zbb059fd4bd5fdc17807863e2ce7422794c2dec3d2bc6af46f8b390603bfe8a7e42cb8f774a2e54
zd5abfea8ffa35ce0e5a60ea1f1b97a362f43e7d23838d8c5658dd1ef06a6b8a0704bef4209c73c
zc97ec1b9b275936f552b58d347d4147ffa6e3d26665312a4f4ebbd26afc9eb7c4285503656fc4e
z6738d9ad76fa621f761f6e71465ea920f2a96a571e0dce8663feb74a2fb5dbff2663d3ecd75bfe
z286abd6e455c25ad32ef0252dac7410bb910b078e571888359401f0dca1bc9eb4b906cfa0f3fc6
z304e5cc526e9bf100fd88b880d666f95809241ba2b2ccc9833492de75e18e317d9af77bbeb4145
z22eab6f8ab37d7c6ada434974f15a2156622052aedc64d88c338fc0604cdaf9b9c064db9f2a8bc
zeb594f81185b717eb2c86f2868286c455083232ff6c1ae93eda03700deed7cb1261fbfcb6edfe8
zf52fe18f78127cfc68be822a2fdebb83ba4f07f8dec80345db40b40c842f38ba4a674044760b0f
z38f3b808bb1b2fd6e5619931c9f545101717bd4f2e2327e11576f482038584966248ba0b67c0ad
za7ed7535ac0ffe34e879f42b546d10558805f0b4660bb06e557e81673bee16bf355f4ed7461558
z77a596ecdf3d688129797d0e9b9a91c73a78b3e3cf35c25216e211e6bb6102454a22e0035749ac
z0fd70cbb894417746e11a7aaf939cfd010e9525d30dc58a32958f9a7a0d6b3d0cae05ead3daf43
z3ff52570f5663cdff8b705af6c1bcfc6d6bfcf2448e38f95c4ce0d8bb2504799da23d8eb74f50c
z05c53dc36ef5fdaf69835c8d65dffe379f4c0a1356e0a6bc962214b567f8bde59f60d1a1a1d34e
ze1bbfd49083436ad72c7c79ca7687d976810a36db415381cd2ad44e1a2f950b1f671470c364e8e
zd32d6240b208bb76e0d54bc3d4b249aee15ef08622312357ecf058bec371967541ad415ac157a9
zd4589979e76b9cca4085e950560abef24512241cf6b47b2a358dae2890c1146bf033b746f55281
z671b3ca5b9b9275ed9cc3bb230def5a763207376489240e761c19aa181f570fdd860e67b8997d3
z1ad4c2a468b56ad79698b2d98db8afff49964a7c979567dd9f06a6ce251c0ebafff0ad9d31b978
z2d42952c436b59e076c3e0e89ccf6548c618a0ab9056d186d0a83fdabcfd9d73473d320342374f
z3a300469a0f7d8b67f2b4d340383f2b704ed046b431d76d19a16358d30605c22415a1e7882a57f
z5afe2cf2dedd8b57b02598fde6a63add114c7879fae27c1b7d90d94195433311eadcde08670821
z513ee83c3cc9bd07644ec6af2f855efe8eb05bf9241be994cc7154ea06fe4ca9aa08925b12401e
zf8f3eb949143b5fa0f336ff1c77f767c6416922c82782cf509d3bcac3f6a7d0e32670af452beee
zd172b32155e8923d0ef95853299f258aa44684ee448b32000e282260d13e7e50314dc7d8c47d5b
za33760595cb08b63b544637d797a69bef72f032aff61f8f1a6fba24980d21f710ac02d7eb87804
zf75b0a47df4e5c5c8f577bec9fd036558fe12ec1715534b0f28d9092d23eee733a520c37bbaec0
z26bbc70c5f8ded07ad24671230b6688abd6e42c8be7b0c920fb984d2eb08606e7e64db3d542487
z8a92833ea326a667fff95be47e92e37e33451677d662ca7d2dbccccb40837652d7bff4988b1e82
z664bac854b682b10c3136f78eda24196e3a5a25a899ca9e34671431b6ad893f1749c9d71028b60
z20cf1350b97e8dc50c61c82c0986ee9928bf8dfe3cafcc409af122eab28f12248f212dd721467d
ze358e3374d2157a45e46e1377c3ee26c8d8aaa24b7d74701e18ed2ad484e467b6fbc24e58e9fae
z6642a980af4110ed56646b2a950d51e57f5da37905461cf2692e3f7a6f906de7d92228ccc29e36
ze454875daeab874cb2ab64ceae9114f4bd8771c3a5aa9fe020f2cb535fb6d2a62efe6cce2bd50a
z78a07aba5fdf1c9636076441bbdfeccaaaef739507229f09fa676be7d3e49e68fbb37fdc90d9c0
z24b65c70115740eefe496514839b0dd0ad85210c20de35ec998758b7030700fb42505dc64b290d
z2e6fdf5f870f2bb1096f7ddfcd460768f1f0378d076c0cd068322d893970550d46e05542622c6b
z797e33aeb1b092866e2629a47b82ba9b46dd6ce45e8396b383acbe12ab2c9520b763e90b03f067
z4e4204a43f0d5eb7fa121d6972f5439a6f619abe2e3498704107021af7db0e84dffc8494d83b55
zfe17d43bbda66e62c3a7d038f7a55cb25747b8e966dc573141f7257b3ba5d27a0a19183c638dd2
z73b1595e5a971d823a3baa0b4d4ed0c773feff89a0c6ba4266502319e7f7f06bc5387a05421192
za5cd717fe682671f605b13ee4dcf19ea0855de6bfae745629b2cdb079b7b21a226df010ced3f55
ze9c9c86bd834e6c185703e6484f5dddb3a4a92e55f32516b159ec1397d324f32a3da1088e3b918
z038c2728493d234879f2a1d752a4983c3764c290faaeb2d05e967e95424d06731899620098fef7
z17cb4397789dbe2d6d8bc4f39a386e422b633e6c24ab2cddbd67ee6d22ed925e75527a6f5b908b
zb0c0c2c6c9d5295bba663d4e189d16674fe7d176200210011e110e7c09c04dbea8113bb7c2c539
z6b0e05f3e585c2a100c1e161477b66fdf1f7541c5faf1c4291fde1451560613c930c32941b00c1
z8709987b4cc3ee57b443a5ae7ab8cefef93d55469df656f78eb425f6889de6aed719619747652c
z4a2e47a1d0ff5af745a3d4474377d35cd3be3fe5034fa8c7598bd7af7b4c601ce41e11c1d0c6be
z22582767cd90d8fb0007e3ceafd8c125ad15e50231363602c81c00a81b82a8e50036360ddffe94
zcebdd3843ab56a1cbefce60519cfeef2caca06bb8fd2a4790c3bb9bf8e9a42fbfaddfd880d1295
z29b2b6a68d8b2fb85de7314608890e099ceca8ec1044e9033276166da0e0859c4835464676a24b
zcffaa19705c5130ead817781955b3312130dc53ace7dc986957116170a2dd1ec4c74116daacb44
z91554a9deafd1efacd01874bba87803dfb9f978056dcd7a2ae63dc5310f2d1262c35a930026692
zfc5a5b7bfdecd8155aca82e523a80c36256b95ec0efefa2a4081c35469c9e02943a683e5ddeae9
z3316b810d32b641f15b0f0455288b402ebdebbf0dff2da70f194879ae7b57024633bb52bff1cac
z35861299d96158ec21abe074462231f33fd0cbcd7de34f5a19b718f9570ea2b9f132f4e57da506
z46edac31e3236c45fc7df4a7f60c7d90a97f22fa3559239b80b86f00e340231a6393ad2c66065b
zf92647cbb63802733e11847e6f7ede1392282164c8262011af5df085f93e282801320ff763727d
zeceb18f4ba2588aea7a97c5a6f0ce634302e783604091bbbf3e8d120cfde0abf143297a14571bf
z0b8b752ca2e2d47af6a7b4e01030de99f7328d2098e168f5b24cb7a6bbb1bcfd98cebbe627ba13
z13733b0430ce2745b5bcb6450b59569fcf983d1406ee4feda4d42f5e9d2db1c52c70ff8b229ad3
z629a722a0073a8cccbe768b6d73af110c785c61d591442418b3457df7a90cca31924d1265e7928
zb0997a7a984c167b9b0d97293653ef26c5e780e3a662615e10c7e42379005390a3be2d4ba7a4b1
z0222a5683718c67d35239e3711d178885f1e2feb2056b77bab7c9ab6312af84213ba6efa0ebbaa
z7643ef405f5fc1ade0621b5f81f34bc5c48ac879764f0111fac748db0242ab6b6cc750d1ed882f
ze82e784e0774dcfae3bfd037352b306be030a753624b798dcd99dce3265ec23dab6e95196dc2c3
z48c984c59ab6972c3c93712f1a1f836ea818f70449c72f4fac3d57d353ba80bbe8a99dae8946fe
zbf90707c5be6769e6b6a0fa522c2dd26a8e3567308c17686c200d8a7fbfdbdcf9bf11c3f82be1d
ze9bb471b73d4690430299b5997cb823176d3c1c08d4aecc0775a28b8aaa3c38f6ab7dfe7a976ee
z7906999d4f53a4c5f2f79071d44e3628db591a7b086296d2e4ffd4d9227a3f0236c50cffbcb7fa
z01b6cd0529498ab07d985c489435f225588b0f01a1dc4ebac049707b04306079cd13287716ff6e
z6e9274d9dcfec4c412d3f11a52cd09c316f0a632c76737178689519f2b
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_ddr2_sdram_bank_module.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
