`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab30857016fc53a
za25afc8341302f0c829d94450c399b8ff9b0386c187cb854ee330605b7b59da379b1f26f488e1d
z36e675f0b1336408b3a1ad87d0723054f952fbefc8d5a33eaca6ef5be8f42bc59870a29a5cc9dd
z4fec09ce6e44cac279651402e7e1f590df88ce49ec26ab39f12b4a02855703c6f03b1e85c797d7
za357087d98e5b1f45502e45892e5823d6fa4b762932009620038c05d74efcea7c3fdb38901d620
z36515d0824367e48d1bc182335f158c262d396cada6b0ad58add4f945eee634c2dceadbfb5118e
z14969c29a743830a07124bfa78707f3952b96b0db7af7c9ff36f77137d8c490c4f79328328069e
zd7d5280e4f95742c9841340368b9764f0f80413adb175ecfbdf3c40716abca7b8cef6f7fe92ab9
z6bd2453f1aef7f7899c5365c5c83793cacc7795c269413f6cf0dabad14d40e9285afde8c01a47e
zb61893788ec5060288cabde8fb553f21b02eac61ab0b48ad3d54f4d1d76508b22f0c600861b5ce
zcb30ba708be817b1f50f59c0f6fce449203e7355c1be55b662fef3f92ba58243d81537761af8d6
ze27d7864d2dae99372b2b75bacdc0437a4f7e011d68c3487a89759e3625548fcc920ad06471ee7
z2d701aabf726859343208b0a543c73eeff8406febf277e3babff437ec820fb49d6b78e73bc2353
z884917487d35a6cd06d7d73ccff5f05355122888b886d1b7ae29679db6c9d2d7f218ac9728369e
z0ba3297b105b1781345d5dadc1077db50a0833d4730649f7637b2138ee147e4486fe0551f541b8
z43cb1f566ce4a86a39651786521e6c831c0a7a8984a034633d4209a41890c86668029516983a5a
z2a2918caecb85c3a38d21805a4b7e2da92879621bc299fa7b4555f7e1319c222d5509f48164b83
z9f45f9b9fd8b57ff2290408ba1dbf726ff7b13b8cbfde6de453a22cf49001d87d40be9d1294fea
zf8a4e779eeb3a77fd351f4e30844995b607c86e83ed23c87f1e3e643cd626a797a57229093c8a8
zb49b28c85dc6a1ed8378a68ece4f75f7bc8bb425df5a97e4918abebe960a92a0cf021afadd210d
z740e80f431452ce69f128befc87baa75ec9d83b23a4686f48b2cf323daa0a59a3e38084755a631
z92d4a951a4d8b256132c71155014cc2a9019d87ecfa9868729fa4d25d8d39ac022b19fdcef26ac
z69ce6af9f588b6bab976bb0deea06990aa19b72d2e4297065a463f37e0a0daed85d3f8ca9d9451
z2c46eb108943fcefca599bc3959a63f8f70f69179d930e368daa26f925c9f1dc337a3df12f0fe6
zc6262ea9f96c6110b734e8b9ea9098d3e016a1ecaf2f54445121c3414056e47fb627c9fca22d98
z199446dc00bcd92c6dd56e1da7c21f7310990a18c094290dee990858306ca1643f488deee62eac
z343cf038f0817bf0e7212c929b927c0b3217fde6af48ddb57b883811b066a939536769ecb25deb
zaf964ff94302fe8dd7e399d60bf802ed3fd9eb7ea4025a06eb854182e5fa6f23b6f44381afd46c
zcf9d05ba4cf08e04f37e3b792cb917451401320b190658b9aa84de62a4f3852b56daca27233083
z9042b64454ed7b83677b2581cd07d466033ff3592df15c67cfbcdca5092f7ef4d3cddf7356d15a
z2bd4f6945ba3ab9d24c8a03c4042b3bed6687e6aea2fe6b74dd3d430370f2574d84216aad60d2e
z1bca40940d1bd0d45f17c32bef5af22c011f1ddf8a069d46b688fa7f948dfcfc666d91e33cd339
z0999f1780a8a0655da57ca178cec0289d0551c9e0ca7e2720134077a4edd450a113645345bb585
za7ecb61a96cae8cdaac4b43d3a8a6b746beea798181c9a5ffeedc750a90e51df7017ff9e0f828f
zbe4ec278f553e1c90788c72264525783d070ac748baf9b31bb2184c4730ff8d50209dc28b0dfc5
z6166f410bd9cf591a80eaedd150b997b9fb690241eb0a39aad892016ae37f588c0d6e3eb1a4435
z466eb465ec5990b52ce8c40f7dc8fc88b3ea8a8279380fc19934e98d267038906899a79d9da68b
z4f8319af725ee534ca5543173f6a2f8ad351ad1791adc21eb276e2ed21723892b3f1ce1e2879bd
z3c80be845e0868e6a3d8e8a6c3997eaa813ebecec87f708000c27aeda899ffe02cbbe532af0b21
z7e8cc679ea3ff08fbc149b3ac81da554d45f9ae372b1757a9b751dc9ec911fa6d837dad94a5252
z6383a8c4fe5aae2a1889e014166b382b649133bc6ccf53d2b9b96fff7dc8d80e3102d14f763a1f
z889128f49778ef9d5c3b328b310f14ac7038ca689aa9343df145a7f7a22617a5a3e5f853931b1d
z0bc50e0997c71c0074ad9172855a8d62593562f06cd1ca788f52fd7d3c1e2b32c9fd78be060c31
z2afbace0eb9ac9aaa22d8a1bb86a5c5d097eeba68a5db669dd6416bbd9c0cbecaacc22052c8e16
z5129386f49d41955f240fea81526be7ba1b8fe4cd4f430914c6d85814b888177b709a32cc8db27
z3a74478bfe39a3adef38fd5a13bf1a8458ed41bb4d115111edd87282a70d0b3fc66ef6aa1e42bd
zd8c175abcee42350906c48938a0e388acb3950d5cd7961a394befaecb51953b63d6a72d558ca49
zc96fe81afeb694ebeafe916f3970b3803ee454a74f5cdc9a5a91de18e316dfb39301e1f4d154f3
z1c212273906d802c128776a8296a0f6fe47378def4bace96337b579859c1d26decc31ec90d69dd
z397253f245aa85d5a1bf5d9ba596625a0a1bf1c1cfc30e5cf727646123f169894e30abe71dfea1
z8e61ff0831690fd7ba08edee737afc63c01f3957b140ffbe0316156a09784d2956964cd98a3318
z4bbc063575bc71557b498d9996868912ec2d6dfb3716b24e2d0f01c23af2fad2c56ff1ec89b90f
zd61e602ab83c7e5b73ad081520831e88c973490135986676d23a1d9cc937c44bc581ff6d758ca5
zbf876d349546aaf49691bf41a4b666c8f70ec7af3f74e9e864256e8d77ab941758800965e8fb07
z91f7b6a4f9cbc41133d8cb5ef9454e1dc3235922eb4a28a0a6fd8200f0dc0028beaf4efbe66d10
z373c0e8af8bd80869c0ac1ad07251447550b23c7cc4a9ea233a5e8b7478eb9b64ab396550c4162
zcded83722c13fe66a19b9dff719a07008e566d9526f56857e88d8a66dd1d121f1370079dc21f70
zd4f29d6c43958ad6a0cd49b274f42062f33770ddf18820297720b0ae79b9d7e68d086b487e5ba1
z683d1839ac56673ba1f94019dd6a81a4b818a2dd9f6e7cc0761fe2de1fd3ef09f9cc2fb4e15869
z1c6ceba0166945e38f422be2ac1a4d9d7af091cfe9c2380a16dba0ab7c8006efe048f8490c49d3
zc389655c25ba6689f421a66b03b08fe0f370aca35a1f2f1585c09a5495683fedc4ad5b030cfe54
z2088f73db2c383f3044f75c106bce4d4196c3a6e63f8b49a48490b08d501beafde5358342eb3f4
zde7b69c6ce0896dfc5645eecd0d79ed84e68e0254a5e0c38b5715eeb393188b9b2731ad7e1556e
zf740c451b2ebc86f5ae6321766496d063c18fcf22bf78d49896f365850a2fcb237a8b3aadc055e
zbee2a19b6846f469db9829bb67f8dab80966dae3074c374418f660b3de5827d11c12241655c9b2
za03ff915c1b4b16c065b3c65a88d3641c808756a1c04d763caee3204815fb0d0df1f6c2f34abaa
z479a1b20f8c50b163c3cd0fa2b80b6200548bb4c32d977bc0a6cd0496cd9a1babfd8a405a021a9
zbdfe1c518b0e6bee802cb8970e790a18a7c6ea207a90092f9c1af116977c08195e58502980b5d5
zde8e4ec34a379c67c48dcbb189ccd4b69d3646f6065f5c2e09ac449a161f3ff568afb852e14513
zfe36e6e15403d3becdfa185da1f401b9e7053a6f72296f4801af9f51b527dc260dbd19d39137bc
z51b27ed86d26bbb063ce40870320e8fddb3db46217f1c59ae6ff2291e1c567b69ff2d3ba54bbbc
zc50ebe0629962d555791e3d5d534b9ebc3e1dee32d1120b381a8a24005f693ffee866400376ea4
zec20a2ea7b25d370a907f1c3a9dba033bbf32fd6f8103a0cc3ac2b2afb95b56075d6760942a962
zfcb0701181f7109cc41ca55099a8b57ef6b860be5dc3ba19df3c3c1d00453300b7e04cf58897f6
z51d9ed5e3f5adf2fbe5be7c4301c303adc8ad670c8277ec316489d6de8006bba548f55fa74227c
z0c04ae8c57fd52875bb2d98193ceed87dd69d1f44423facfcc24fbadbb318e08870c73c9c492ee
zd058f74b7df2cf020cd50ce343c6b78602a64843e40afd74bf0785b5399988c1ce7a6786912513
zc4f5afad12a835028a9645700bfbe1e688d920d062c2b4d888a8f41cc4c6cf96bfac55080e6cf0
zeb811a6467c81fd790d2318007244300d0551a291ddba414ab843f232b8b3cc3f9cdec5a19984b
zd5f07c26ead028b6a1b3a2c07c1e9c34a1420646c6270c57e8fc5efef3cdc28cc25a9c4b792ecc
z1320b16c486d2e59da6e7ca9f529b854893d846a3d0ac0d5a1050819a866f69d2237806c157f91
z4c51064bbb090f907a4e62717ff8324c98fce35fa7b448ce97737937eceaabdbbabb32ab4f9dcb
z6a114b8b63830ec0535de639c516c684725dfd84c50cfc0fb4309fa1112fe180cc6060af764d81
z1b3f3109c59e344cc0fcaa8a228678c28c59967d952beb4305e74991ef76e301aee5e90c042bb7
z0dee1a6ea94b810ff927fd952adcf8d6f1bee4f2dfc5ac37056308d38abea7806d4ade171e0303
z18ffe0d5f8c743112516bc57e4fda57015bc7420f4389a22e937c230678db4f3665e2b0514402b
z55a9ecdb75b0fe7fd896756491fdeb83460d58b310194b01dc520de76b2ceb24202406be4357a8
z8a812004f3daca743a3868ebdcb0817434e75acc24c3fab3da4fd3d46db5b5f1c766df5c5b49fb
z68fa2172bd180a9b137878c9f80671b47dabe05185a5c497255fd5d4d91e37e833d0a0efcda6fa
z349d9a682d069b174c79d7497e460715df0f6f5abbb1eb8156b826694cd86d9483d7fe146bebb1
z8787f7ff027ec46306210e4d24e91c1f6f210802a7a2e511dfd4b1de7b4528c0d1e50a28ae8fac
z5168b4b41195a3ef70037f52a5d3c38fbafa833eafd35a012f9ec74851351ab7678207a0f4448f
zd31a4a91c6fe256abb7286d12becf3ce651e49048697cc4e87f15a1de90c960bd4424c037b5668
z65a85da29e5af3479832901f32a87fac2a29214f8ea08eecbc278d685b1005c6d28dfc3374a7a9
zfcf75e9e7f820c651c18d31f425aa4047719b5daac474ea39f56d49d0ee6815d3bdeb5226d2113
z3b96fdf1da4b826772cae6cde3379c87db08993b1227b18d6ccc6fdf178d33b198e3abbcd11895
zc48a59ba03556f9fe18f2dea178279d4e695355bc56af627de673e1fea6e9ae3e068167e2d2470
zde07bade38accd7b1a3361b7b17cd254d2dd9fc936cfcc9c7f8176659a522d58162fb0126d1b3f
z78b800e8e2ce94eb7dd3575aa893a75e43dd2136fea77691aee47c076af2fe47dd1b08d9789504
z493439742ac9b500859eab12867f486fc52b1d3c31a17f55709505f8ae847c0a6097a1dcb3abf7
z42338064f61a8a7a4728da48b4296da2bd3ab981ae2b79c67b51bce164e6d258d0ab43c4a0d21d
z10da37928f1eac029840856426f8ba9b71b2f2f2f71588f94607996626c990f89a03114a4bbf62
ze410f21567c6d96d7da7117be709043f695e6cc18174a9d047d15c2f3083f7c4fd2bd4fda99a60
zbfd20d81c87896446486236614d84811b8bf97198bebf033af53bc6dbe214156a5b0b242affef8
zff5d3db8f29c4979cbd6f3a00ec6d6403aecc5b5150d2df1b177fe421b61d4a9075f15ef5cc059
ze52e84a616d42973dcbfb31a676f5a496ae5067f69f3058044885e9726b919281237c9db66a05e
za1256e599678cb7d79ccbfa8714c91c2181dc5d0c5bb98421e7f62b30ad3b21442797c3abe2456
z106d133cf48e5231a2d060307ff4cf05cb4829007e24805c77af222c2a0287001921683814ffd1
zf9542d8022cd2f37ed60aa456b1bf460caef67535b99fbe2692b48b72c3f0792fb9872b38ba451
z905ce9a6589d8ab8fae59448a5fe71e8c42a9eae3510235707e4eeced4e3fc8c113fe4dbd9af02
zfe64dd34ade144e809b685d8f4cef44e2faae54ced30f027b0d07dcede35593776e937c9a31b21
z51ee642c5481d5295debcd99586ee6ba17c3f8f1b52b784fdc9c22571c00ae9d15a1c11187ff20
z59d1fafafa2f2f26a554338dde2f9704957d209923d4a8ebac73f595f969ed6a443d831ec62b50
za8e49751a9222fd680350036d0adea8500b22878ea3a27632a08e293b09c9ee2989d3169334380
z417c53355c0d25819faf419d2a78e0147125eba2d94c89d2619ca83d1b9a21bea7ed4146d04bae
zcd9092649484c727c16603b9abd27b2ec6c8e4fd42a27716fb441a3d924103ca995d452eff6499
z299ec0946b2a99220a295f41728f77e563cbe1893538f2f2486e416f1a222bce18df76072e6ce3
z94afa1c8c92f5da9187a47b84a67519d9879150c58e01597039c670459b5ee3e146652b552fc67
z3de95240d7f77c799a6d90a714c76cf96475857ed9f87f8875441da64aadf1cd6056924406fee1
z7117d60b7ea1595b13706e36b71d3a232bc3771e486d84a2ede38644cd538233c67f9384d9fc7f
zc698ce1606e98823f2b5edd67dad5cfb67b2421f6b2d0680e7fdae7d1a5dbcad57985793afdfe2
z09795b7ca8606baee9a0fbed82936a3dd83e1f0d8b41368999ab5c2f375cddfd9920d1fdc9f3b6
z6a981cc759b04cd73d4f35a160b8770dea83439d7ad2a5ebf511154a1b2b2a5d5c9ed3d1db0c41
z8a9e248bf1aae8df83548d84c7f5bc2ca1f99ce65805ed52938758a0ee8ecfcc61539df82cabca
z2d12b334edd44e12fa3798700e7c536ee29307cb6255ff6e8098e64af530c84c8e5947ab06f892
zf18ee6b80de7dabc01bf07b96dc33e2f25d0ab4f03cc7fa8ac4deb1ae0e22debbc594657e01451
z06550df53e94e33358608fe93237b85c9e4e67f97026c92a0b0f91f61eebf710ad45db5c47252b
zb61f7c137694bdb7c508583de584e46fe8fa921cf2004bcfd1b6c0bd42fdca6c8a7733ad87b2ce
z6d99a34a5a3d0b29279a58b1dcb8eb78a33eef7bed72ffd970000e98ac0d773033eb63cfe1dab2
za75e762743a3cdbeb8413026bd4e43169a822994a691c2c4c7a75ee0d9ba88c47b90050c4dd827
z0219fd3cf48121a4718f28e3ec508f8fd484d2e7fa6bb6764e4d0e8e7820c6ec8d6de9960ae65e
zb40dfc7033de9d48a9a56b568f5f027cd3ec2e4a6f98ad4f39eb6069cab5c747097b9795e63922
z58e3de7c603c824d85d384ac48d3143290349131cc6eb9776d6524ad2ae8fc14f2613b5741e700
zc8e6f612375a22218912326e1070795b7a61d97ffc0ac2e1eb98a408b004f83eed9768646f5b3e
z844bce1c3488c0fc57dfa271a64bec0361420eb3e9b7a69baca353f8ea8b676951208a1def7c44
zf7c614db72e0b84699e1065ff385937f2b8a54bf3e2ac3d46b43572d6d62d3ea92094f293a5370
z47b6533a44c9e5394c12e7374a9abfdc016f4b66a0463446e20d163aa72019969f22cea430a2a6
z83eb1d3a0067a3d01e380a02235b85ea07af175c123827986ae2c3563da12ca113199ecabfa599
z549a5635bcdf75c288ae13eeee30d53c93e575324e358b9c68eade3ef3fc18fd34ede773839588
z4af681c2aa6ba54aff090030fc6d5c2ddfeb46caa47020186157f4507a8401fb33d197b18215f1
z69a79ce1612a13d0b581493e675bc962b8351a74887954ed37e8b9ca01f1ec0e1ad8837df15339
z73c2a55aa263b739705b63085590c040e5947e9bbcbe81668b6dae2a508e382cb466c0b7016a0f
z5ea6780a22ff4081c0cbc011e93a1e4807bb3aaed0d6692116d4a6464f0621257c1e20617dee4d
zace0e6850fdffc4a3468f066f40f2f034f92e73e6d4442e99ee958bd335d01005f01e6c1959009
z56e914e2ec81b95dbf5bb02434c88c6f2688aac2d8aeec729887b876e0e2794b6ed0a9d89ef7bc
z55e2bfd44e2499d51bac6569a43b4333b4ac13d62c223a553ffeb5d9ff3857b300ba219e027f56
zf55580349dbbe94d6e0e3a7eab61d4896d7a3fc123cdf3ff7d2fe9b286e8b9e3a3b75bdb13db9d
z140b0c367b4fb00a4485ce183a735bb72fba22b5a4c36df0987024cbf3156105c1d7736d048fa6
zfe83e954c7439e5e63e79b992022c3f256cb4e44bcc1a6bd817e9c4ca0d017d9cf4cbdd1f08ad7
z833f6d658cf7968bd999eedbfbdd6e8fc5b8a59ca4d2bc176b2474bd7880f7cc447eedde09f958
za897f811293dacb8f0a910cb4b5e6ceec8139005440897c7bb773b53ec04f6f669568d04f55398
ze76316a74480192e04c753f6d328d1fb106a8f08d8ee3f3ea35a6e5aa2491f015a0a630a0a2888
z12aedec5147b74d5b728881d6f7de858513f19bc648634f53c450b54512840f41827f738552047
za7e1d8b85af7f7dac450c5b98951fe1acf948d3f2d841bf3b3c753cd106ba0d7935f31d2943215
z44140f152dcd244aeba28e595950084f7d6196d44428b5a25175355ca79fe19b4f7131389cb36d
z326fe9d92657fdd3b574e15689f7d8ff9ca5d281fb184d2fcb88145d887099e8030a835547933c
z6c0c0b07c0d5c6f88fe243acec4a24ed5bf7f7e23cc82eeb8f68af21e1de8c2a75e0d33b855ef3
z6fe16c6c219007063e28763bc8d44f38aa45549829c9a629078b7dc323b199612fe115527059c6
zd8af586efdf2be5e9211eafa6447e224a2c5c17d77e888d06d1a3d61d7586025b5d98902fa1e22
z42e9462a00c3af38d5537a28b33cb6242c425adaba2cd5fcea7658b4e6bf8c121fcaafd3bf4b1e
zd9f59da31bec2366ccc01db14dc25d0033060cacbd01d32d447301086218eff6f39b9e53d6fa9f
zdeed3cb7af3f6f8b07523a90bc98d8aa776722b03158f9e849e827509fff892b1f9ed353998da2
z3df3862ad803c9615e3bad608ab24835f26ae8331e4e66b0b647d1933e84a259c768bbf98fd64c
z825c8b70ea5088e219565cc90adda6d2a9214c97ec33caecab41328ff00cf68b792a3c9c983c05
zea3c845ac60b9727e8ba22ad883a2b709457a4b8b3ac663f9200331a92162a2047fe0c820b057e
z29db09e422e7ce667f7fcec3b9c18d066e27a58ac25fbbd4c30602ce7473d15d22552da904b904
zb273cb1b77935e7d3270b98053868a80bf11e438ff42dc871206c18c825b2c8aae9796bc99aab1
z6458dc5ab05f1b864c89fd7f8ebf4142db36504caf36eafa6421ada88e535ddc5c35104c2c2969
z80c753d8b9c9341ba632fde9a91451125b45258e59e6cb4a471a1fb6473d1d1ac8addcbc9d7e8c
z555d3d50b6daf69c8cab906c3509bf5a9b17af4d157dcdbddbbe140ea0a00c40ac04e02254f9ff
z76f60bbed3df1cd766e818074eee25b060ff17899d346b52f6333b530c16c4868b91be3f258335
zac601867852025eb7ef2680ef6e328fdecf783f9e3d78c728078851869dc805798131287b6d6fc
z84e7644e5b478936413b0be00889fa381a51c5350c85261a44ba9dda951d3cbad7bda004dbcb34
zcdd6decaab712002ed0a34ec4616623c7a5d2ab1e2440c140157fab865f26251a46ea18ad7c878
z6826270ef4dc749baa03fba6f5d20dde5413928d5c3fb2e7c17199fbcb431cda6dda827e248520
zde1fcf97af040df8d6fc0de6339ff404765f753249595dbb45d09f971429f46f4b6cdf58d92736
z5bceaf4e4343faa8e008b8ce2fc942c276ea62535092ce7b47f6a7209b7e952a0cb4bf71d47d90
zc098577125d8a9630b191ad9c324343c0c969a1cac99a60445eb93901466bb601e704b81cb1190
zbf5df50e4b76cb7e41907f3a326aaa3db5cb0b7dcfe0b1268fb6464d1eb75f71b1704e8107fc96
z86307234ebcae826b9457ce214568ae89e7d9dd6415a7e0378f15e4b2ebed5286f632786297135
z8666569ce6c20cbf7dee24444f6734e5b4e63d656703f268e769e74d91f8de2b3efe27b3656d98
z1c43825b529934fd7d64efad5a2aa4f7f5d4f9c2a0d9e181df72da93b8ca1037e376b99bd6417c
zf5b988da0f41df32d9ae088d64391ba99c3f78bab05ce0113a1e2ba59e47ffbd47014e64669cb0
zd9bb6a0ee7f887974af0c67d715ceb243f5fccf6fa11922832b5a171bdcc69c45f19e4ca2a90d5
z9b34b4c892200a211d3e6c4518ab087671158bf93744282eaf7aaf47c573e0c46ac411b64b0539
z11a9c17e5420472c1b98506fe8cebac60ccf9701f5038ca2ea4e249b723452f1e3057ac6399b57
zf77048cf584b0ee7378d95a0ecdb1deacc14b98011456e60c50acd4f4d827b2b53a9dda72379e3
z7ab5356b27ecf3df376d0c3531342750b5d97802fdaba8510b1f4715f78b4b26427fb2bda58526
za91b7a6e33804ade29e88122803431fedabd1d24e0695666caf9e36d83fe31cafff0126c2df0f1
z17d2384fd34a2422e645a46b1e94ab4c119efc667e1c677fad1294fe377f1a3be29c005d607bba
zd9ceb8982f3aa4a2a48554aaff821f800041b576f04e4f42d93ce2c4ba07807e4f8189a12bd98a
z40b74a9c156469bf3718a486ed426539b531b4278eab6d0636fc650e7bbf6532a2d87198cae021
z75a862a7e7b9d95a64e37cae10eb7d31e171f73f474894a084ceca0d7680ed107b862fdc67d043
z781cb54b1b77f331703f27cab48c4ccc7d8cebf5577946ce68481ee2a3eb59f3b1224c3389525f
z35e60cc6e01a8ff9a2571355f579585b7d89e06c97571f761979edc759eba4c9976aa61afb391a
z7f525107a92d03cab8b87ff0aba2c1117992abf59ac66e811ba8023c139aea26df40b2bc5a518d
z26728f3a42c38e6d569baaac83f4bb12fdad25c5b831f5993e810da2b021018f57679c880737ac
z914d2a30e4ada5b377fd07d35690a996fb3bf199bc46b3186ed46cb111bd630a48dccb6045ea40
z03c53f1998b1b71b5e900976a7a593eebacf93e5bd49536e2b31d4449eeeb620c80067d373f489
z10e6b1aceeb4599332a65521b210f00c26cdbeb46403e12c97b3d4739721401eed1376abc758fe
z6932f063234b17dffb17b87c4fa708f89ef7f1043b4feef002731d68c3381d221f1beba18236cf
zdfade1ea85733fd1dee145d8c6964d9e797d58540641048d5447827f4a8523675d4da2b95484a4
zd492a847ffe038a8129009ce476cea3b000f5759cbc8e3516b0006d2aa6edfd40f45fde09c5ef9
z3a07ce42dcb0d4f077af3b7f0c709998c341287be09bddbd242d3b633278508127050ed85fc294
zee7f12b71dace6771ea74296563736df918b243f96f52e054a862499f7988f5b6253f4a33a67a2
z768e77c8e5e1470b2283d630eb4e5e6f1a3300832561b0847ae119bc3a55770a0fff8fa6a6373e
z45b4c2b379add1e965f4251559fa0aa58f2728d38122c6873859be9c1c16bdfb653b18c54ff6a0
z7560190c23dda3db412af60ad2151ed93c5508d826a07e4a5d0937ceea624a30e7477d37205492
zc58d1f51130b9d1d0d0e7aeec7eb0a5459f86d200046756773c71ad6da0a91dcb45dcfcb581588
zcac57c06e8cbbad75ee64925b7981f031cea63e64836d256ecac0c68b85d985475d5c66a74d433
z62667a4daf2f1e5e538d18255e26f288238f64ccf56a4366a95f9d1c3e0beda884393d3712a819
zbd1b4cc05b098e7a1f9871f476698f1f408407212bd62b8a35d7f6bbe188011dbc59277c46b35f
z87c840d46c4ca5d93011de5205cbe1fedf03e7e545564f078989a7ff58a5d6504d5e4c61de2de9
za8594eec797b83a6eaef4f67ad3a651dad1c962a31c6e1a3db61c6c6a44cde883e35007acf8cc8
z55228a1fd75c553f7eaefdb5d25592d5976ed8f35e434b9028ecd9b048bec5de62232e0302ff63
z0e39796a9ac301a48760e6fc784c915b793f1f8aaa485a662d39c24c874741c6f92717e81e008c
z348bc201fd1d3347fbce05dc3372416681ec03f26778be573a73c1ce99dac79685182f8f00c5bc
z12cfd9e5ab3723ee7f2ba2672eac0c6e4569eacf968ec1f2f7755d7cb26ce56ce0bcc989ad382f
z61e0c44e54c16bc238841bf4876d23920091193e83361a5bfb5d305eeb6a1710be284ea9b5d7de
z7a3ec232866464898f3c20c96eef2f317bb5ef2ac84712348264f4709ec2c3ac5e4f143ebe2d39
z05f7235ce7ee8a072507445850051578e2e0abbf62f28f4db3b35f93dc71f584ac0ef889ebcee9
z7e448137ad14d069e8cc8b4fe9eb3ecda28fb09c9badf397ef3d7601718f7633df4ad47cd25dd9
zcea265f32679920404ff31ed562863e65239bdb9a6d0d5655d694ecde47a4fdba83724ced337d6
z5969344e4fbe3a1609b0e047c56634a9566966ea5d091fb4e5f3f414c5d216c14b8173a6ef73f8
z67129307741120248ff61a0b36eb428a0c7ce9899b82927fd028271e06537fcf1b3d76b18a8461
zab3944a775c973465dbe940e52bf5d412ff22e9e3aaace7d2daf3db66001598ccccc5a61b17f74
zb642b58105fc8445c61752152a122e085fbad843ddc4d49ac9d830708e431a0814973d09e6cbd7
z92e5ba328b161e92236d81cbfbda409fa59fcceef5d9567119a6600d6a32b631e4b1f0e11254e6
z62de33b544949967f8a382f28d2f68684023f88dbc29e791d4385a3c00bcf927ad6bb196713b4d
z075b3f3710e578002ad35ec69d9acedb69236d5142faa4b1053a51af89cffe9c7d917c9e902425
zf5ade9a88ee406a365ebe408211f4a88e2500ec6ecaccaf9825304c537d89979c72fa0101cca71
z9fd33bfe70d88737bf07e19d8ab52e94c2ba7d12b73af3589b4939ebeca457114830e6ea21493e
zcc39019144321f404c08c9abea217e371e1e03bb8964ba0c014ce132e12160bacf8b1f83d1772d
z7de61db9b794d28077ae691a0efb1fe6068843e9bbecdd1e9d563e85abe4b0b2fe92084e02cbf7
z48a3dd2ed360b01e7889778819292f55b7e101322bddb9bd7e50ec80b0793e9b740617b553202a
z95bbe64e2d35ef5db729e4ef58f2bbf0fa5a603463022559d6eded3291b1aa1497c8ec70595115
z73010b1ad7b35b5b9bdb851e67817af89ed414886e24c13f434319daba9b6bad2021d7b96d81c8
z6855988eef769b28b22fe1f28973bb1edf97525d3e6c9b834cdcd880a8a858f6d02ce229a1d139
z4dbbb0f1e41b2882a375286d4b1e088741131ed5af40cf013d34c291992d70ddb9ca8607ff6e71
zb3c66748dbb8a8cb72a467ab9904329ca1c1de3b8a96b7f14745540e99ba49a8336b04550919ec
z92188e0f47c5f361dc011271a6ee5696f54af3b23bbaddd706d046135f6901f33ebde52a02dcc6
z42a31331ca1f158c5c1597286dfbe42a7309dc42cf390985478468236624e20cd5c7e237ba8cd1
z816ffbebdabaf08dfcc5d67b20eee75ca0a1ce4ff2083011ff199866cfe35ef90902fbd724e38b
z8048311327710f10dd98fccc1a91115619d2aff3912cfba96662ad0920b6fec726677fce992bdf
z11c307b99d4cc7e34340757755da1b663547fc0bdfcef2904e2a457b924a244de9cfc7e5d87e54
z9250b5dd5055bbead52208b24dfc0746a354f7f6cce7c0bcba2761885ce8fe220f27dedc59c05f
z0d87105291c9468be553e82ad1fa3e073acf22726bfb217eb18415c5b6f5f8b7d72f8cad5fa5ef
z8020f3431c27eb25f0f4cb9723b9b47e2f9593095fe5a49c5762479d6bd960a9a1a58fd395a1a4
z0d84031746bc162d854683d79aac6900a347404cad89a63bc3b1f4e36b027d6c7effa98ba54d2d
z375ff0f45edbe19843b0e0425180a2e532c1acf9ea239f9ee1a2b2d751e781522aff7e437513d1
zce6b0f384cceb549799610e61f4e25b18c74f20ffc20b66ea4da55affa04b9196e2806f43de267
zec46a6816e6391c59d78679aa24bb4dd0c7dc3971fbe84217fa086d922f51b64062fcd4d1a3df4
z7d43ba57bf653fd6706b6b886c611c18e1e71e4d38f16ac2fb05fd63d965c33b3710302bceed2c
z30a410ea18db98fb11d9a4e89d7302091dc450983b5c233efb296fc2708fa2b5b816febaefc9b6
z8c7820cd1d62eb96c41dd2139d225f5417e32bede172f4aef58573a118a9f67768a13d0f4cc131
z06fb1fab1b5ce43c858a0f4c4f5483eb08d58b7685ca79a2a0f9dce564688a94697ccb96a00cf8
z39475e62a06a95ee6adb019d7ee5e8c793f6b6169384c9b4243b7db7f397ae8bdbc8ee4f31b23d
zfdfb2e272047d92e8ff2c78fd46949e12af6f82985895a1a34603acc8ddb76713453a52a156b17
zae6da84f3ad74c3a482b37cd3394c31fd7e6c6a2e8e8b029336ad5905ae7c16a2a375450cba0af
z6bad209fd3b8c352a98781cf793a410cd1c6a54662e0dfda1890068881329a1c8937ceded0a5a9
ze3523ca9bcfe4b287f3594a52760bb377c22127017009810d69207c932f64e6378742538c0fab5
z27145cb2990a22934eaccd60cc603098089be8c37d385b5ade64dd76accd12e0637c176ab8cce5
z9162c0a508e31996059066963360b30b7a16c9441aaba2675631347b97e826a9150f50fbbb78ad
z5c7cc35b3630b2354411ba233ce2c8dbe08f5752de0a66382293dae74ff59699bc27b9f879e491
zf0004b4080a637c61ad25dff87ca590eea0c2c620f353ddba7aef1685b157ae462b8e89db2bf16
z6b5547b6c9b4fc125c04f01f930b27da9b4723c5335804160c467aeef1aad343ceac0a3c768d1d
za8c28b0a20dff5d28074f1492816c85d8ef2042fb96545e2702f5d5adc6c1acd5f046f61c6e809
z4c28861fb4071f618fecfca3acf288289b43c6e67fb0e1117d357d282513d5eb1ae7f5cfe52b0d
z5ef61d3f24fcf720192cd5c29601286cb8eb4420f78e70ca9d5a97a681aa9f61f6fad1105713cb
zb0d9189c16dcdae93e21bf06b1ff4c3b27ab3ec53bfc107b50c613dc5d4a938452d7e64c0c4451
zef9b357febb6af48a83061f321e5a0df385faf1fdc2d2e351bd4f01515c4284b3e137bc0c1739b
zd45e861846e65675309ac7757c8fb4fbec09fa2522c7f443d5d08ec53c373abfabb8f961b33f1b
z4eed4f5cd13c640325550827526b80aa89a32e60235a6e6cdce3b180d6ecd6775d702cb41773a5
zba1a707c47b39a2706c5f91f6e8248d0077c3749671e9ab072dfbad59d444a161e7a51fb4a4664
zee8e31a5ce36d432fc0048b0889816588f87b0880e0861b874575cbf1d5c4fe4900b1797a0a965
zf7537262823a53e9f73e1b00a1863b149477277e61cc5fedd750b9ecb4ae1865c6aa5c584a8246
za62a106ff5725092b41947cb32b1b32e263062a83119b9193f03a0a6398ba76f001f314bfa25c0
z6789f51e364f1d53c7c9fa7adc52cbb415ddcea489b9b0d0f6efb45b3f594c211f17f426e8f418
zf4a4285f12f3c6051005c989df198cc7ff346b6b0f5d9564840a2dc039bab52a4e1b34295da3f2
z77ef4252e5bc05e5d773c98117a343ac863f4f472e11f50b2572fc1ab76ebf7ecfbdd5b01d759a
zdc069ba99a46178bb4260d9532c24c34d137ef459f323725d1f7392a2f248628d299196bcdeb0b
z907bb0e829a3f518d553dd73447c70825464d93387dacf0092424461ee7cfef6270b88d895d639
z72140566438231fdb1537e41afa8823edf79461ba3a6940b55acef321fba8975125454b23b4cf1
ze5e27392aa5cc7448f55e428da71ffdc45355298392b8376ae285d5d2711c81a6b64ad955e2fcb
z4ee3ac4695c0d7908608d4a4cd0e99599d648b250998fb951af24cca589627edc79d860b44e9cd
z095d6475e8e302c332409c518d853988e7f481c7b3513cd2dc3c69e07151c42c8df1d36ae747a7
zca313a427d976f1d1bc79292519cd3427c345971134c86918d07832b5879ce2d7f640cd8e32556
z8045fa4705f73989a55e950c457a9f1f678ce2227ca6ae0ebfea3a605e4412c23733cd51fdaf5c
z3a10d2bae2ba97e703e3f6b726c7a67db36dd44034fb83ff022bbecf25420ee9c6912a4297b87c
zde74d56f694a3841ac5f537fcbd5fb3735bc1aed2a80a3aed0452b61712584cc7a492091e279d9
z829979e9efff873e608f9f0b14a23fbde881c1d34aa2af151f1a267c5da24e2d62f69776a6b908
zbb1d57a87368472ded2ddc45ee63dd8da5c769153418d198ee3b8b8494f527c2fcfa14d95e2903
z3179f62a3684768c236a1b732f946fe495fca9557bfce841647f27a77534ce520cbd8c66c9d8e0
z4dc150611492cb83ca42289607c8d26567c57541ab4d11bf074c95fdcd051b0d67d5e77be272df
z8010d3efbb6b41680a91d80ec85b14144e0280f78de97688b9c2fad20139b7be9fabe2884d6cc9
z6b8ab39a4cdd14c1dbfde5c8de1318336ef4e5de90c98614bcd0eb0d8e26f98f64ef0105f4b33f
z5a039c596543deef4b14fb56aa4553f5a550456b992dc6db29c7c169d5efbe3d9d3691d4e6bdab
zf7e86aec7b99a8cd1178ae7e3202debf0b58e453c99013d100339b5deb0724f8240c40695542d7
z0bfc3dafe041e0a3beb858e517d9a514d05a9e397ad5a02f4ca0b56a6063c0f1e57f23aee15230
z3dac8950d965411a7d5f1a558675361eac0c07809d33f0ad0b6fc37fc009cd3e3725f3662ac83d
zda5d81cae6990509b13f422b99ffdf0b645cda58ca090ec0b7b0819b41edd9904b0919cdcfabc2
zfb9802349b80d2646b4ed6867e8ab76363bb539a9a09b3f469c3942703331ac3f123380a9e8e95
z6f44c4a963de760226759fad5f0a83a3f532bc7271ff1b126a9b0239752a281b8db2de885b18c2
z2700af24c3597675059b44eb56332dbf2df4a5e86140a31e468a6c8180d1dab4a088f33df83206
zfdbade193c5e8ade43c3d1780bab22d1a2c69b054efb43d9175a19ea23f32f5979d60772a4f960
z3b5f5a56fc402f57b11938e90e39da9b2e959688308ed8ef2a1bfe67f4dd7751b0dda2b531043f
z6d1494d07da15fceee2c41d7a11909ba98fe41e416e2638eb200ab3e15cf974da71583175b4777
z7bb7fec6f7825831d78c39ee196376fe24b8fd0be276a08b0297fa8265da846c358b8d1ac5bddc
z029548e5c94cb2a337d1e86dd6d1150b7b5e0275d0bbf5925351014c6c36674bf8e2dce44dc5e5
z117cafb4fa30cd215d7e727a4dafa6fd56e40bc6379383a5766f3c7ce64e11160efaf50c34d1f8
zf4c04da6a0ece8ecd29571b4d6ad3f7cae2c0a90b576f34801b22cef6b735cfbdfaf87f0765435
z435e707f505fe1968cae01928b8731ebc1a34f0f14e7bf5a1cff5c75f616b332055d066a838582
z28c918590d76b4d8dee7c48b93c438d248e120aa6b7b71c48c442b8c9caf68ae5a8b5a2e45db65
z8fa3011afa3e5475f6ae7e0337656936c3ee4855445d2dbc02a11e9f16da5b8724807eecb91edc
z574372bfcc96583c1787bfe762b0d6da2eaad105fb3c2669162b5e2a9ec944693d6a278c49ada2
zb6a95c27a4e72fc40cc52291f44dff3698279e16645414873c6696d49806e381c64cd8509d46e6
zafa0b7d745f079e4ea8c7954afddff1b2acdc82dbafd276905f0919665f68c90bd2e04cfae458b
z15139728d8e27ac6a7abcc9d748de394dd7ba2ed15bcffdecf871930301ce5713ed77c7601bfb3
z1b6b5eb807ab25fc72f4ea7803bc756915f9fc4ec8ae8f36883987e2d05fffee9577011bae72b6
z2bd6735c581389d7d3c1220fa54634cf75b5bc415dd4008322f61abcdd12cf4d0bf0963c14961b
z75c6ff27517eef5129d5e42f1f435a7b1c3eb494fac0e8ac27c863892391453c9b19945cb107bc
zc5e8a5f19407730e6491c065c07e1333add7148fe797383834d1e48c59f8a07aca45bd34038a0a
z76170fa38482aae55211f331a08f673f21609892da1d3533d194738d11b3c54031a609b70f5abb
zbfde49dbccbf285810e5e736dfb06a21db92e15284853752382028a0083baccc7f1e595f3e728e
z0b2f576dcf16b1525e8de5466a15f36721ba57b8473d3d27a281b0f943d16ad781fa304160511b
z0deab3cb773f14b059e674c79d83f2fe93c3d2b4061156c442a05288b8c815f54458c646b31fd0
ze6016a0cffec8d55c5476f57c48bdd397f92eb71017d44a1c4f1091be6a37c7421582a8e68d60f
zaf7199ab5d631fa2f6f633404628352015453174309c78527160a5dd402b5b890eeb1ba53163fb
z1c78164d0eba57a10a217a83d862c0d41239d0a174c3aa0810ee6b7d8060b34a21ebed83531de8
zb3f5cdf8fc7fd6f280458fd7058a65ba7aa3b6fc9502efb11e17eead2de4eac0a922da83a3b201
z353d89d43c8376211cdd585d51d67a059c1b7a5a129b4bbc5645fbe4043c304badd581781e43ab
zaafb21aa4b0092d40bebbb3ec56bcbea4fce6de7a929975b06d1a73ca232c137a7f1fd2b817f75
z4c2219d7c180a31ea1b57d15e09adefdbf1d8e0eb19f4cabbe38835f710fb6d7bb6371e2b8f269
ze3aacd4a08820e72c7504ebee2de9115cbc80f0cb8899e9a3f1f1c94af2dbf66e4db9945edb585
z810f515c5b9d2eaec9d3ac64b6e3fbf6cc8cce43a6899a0b1a414ca5084aad7a89bd5e59896854
z6c85b38ca2a759d18ffd7309a35d4d4d502600c7d12224160de9e95151dc8d60256bb5e3131cf2
z0e36a8baa83685df8aa38ea3dfe5d4b13216ba41e312569c966dde47a0624b909d651369ae225d
z810008f0d9ba2661c6042a87e8ee602d4d4022907be728fbb6dd996827bc5320a35424fb324348
ze6b6d84aaa9780754992b49d7a41473514898f0f8bacb03d2c9c9c48abc1896238b5024c8c5cd7
z335c5051ed57b2094aceb366c990c9fc70b666e6f4ec1e92af5b20a0db46d8c198f37b8292ad52
zcbd72c1c1417272de13a7f161023053e08908821b628e1fa4ac33cc91ea2693669d9d56d0c4f6c
zaba523f73524d7db3ae9026fb3e6696a9c6283c49179abafefbb55fc732d05281c5151348c9e08
zbe2a1f709a9d601dd82383f5e3bc706289f7e0756b94d2e81bade903b7aca041f9fa244e89e9b1
z6533437f5f773eaa3d70fded7513ca9a7c6eae1cf7029ae5effbe4ce4c22df34bde3a348043106
z3329ec66d5c77eeccbcbf700571fa516f114a4b951ebfbbb597198cda0eb92df94f25b3faec3c7
zdeb620b526534630dcab2dbf4ed8e8a59689cab1dd4270501dd4d8c00c46ede7e2b03055e82a34
zba16a9f019241ed80aabf125289979c4ffab091f95b3091d24da15c54ce391d75fa72866d8a1ec
zb249b3bb2945b9414f2dab12317b4fd4da2ba508254d6c9da3e25218075eaff18182b69eb6117b
z963c6cff0c58abdd28f3dc60e9a529e41c187d31f1949ba7f241f1aef1ec9cc35cb845721815e0
z85fcc6b856de7f32b4b9fdd552149626f3b9039ed89e1a1346c80d3630f75df895f9ea15c8336d
z4311670d77c02e6ce47edc84839e13668a7e0957e8ac1578109c0503cb5d975397c72c817a5938
z74d574fd310ede2f9909b0af5638712d0e392867262ed6fcb9b032c38d3b0c04bdeecbd0159d6d
z26ba361445d34bf1919b5778408b629a9b47f42fb0da31bcb82758cdb723a9ba7250ce0623e301
z2741794f6427c58622ad92bb6b1d8bd0a1f347803d1c81726395b0c86582f4e23cd3f44d961174
ze2bd288cad4b5e11f9377593525a81d9a3970c2337c8fbea755e0859f592093f97bd2ce4c374c9
z28ccc6ff73ccfa0e6f1aa93d8dccfcab42a7e47b7bc7bc8c466c4372abfe0467d89ce00c20b137
zc59a8a8b6eb7bfd5ee59bc96b75969fdf35012f3b83b15d774df23eed2987d49b00f4a8c20e5c0
zf941adc4bf0c2b0da063eb46319f0e1abbb92fb906e9186142d1469a4ac0197e95da33b3515141
z667305efd6b5c54fd691d470aff309e26e88c4f37a5e3a442efc80c655d55a829a4aeb57f607d2
z286da723d6e0b66dd01aff63ddc3474a8da744746d395da89c7a718de8e3454c109b941367480f
zd5ac584bca8d8b000c58e280007bd3cda5a9fe4894a1d35871b9be2649dc77ead73a02dd18d41d
zd559fb0d149d5d986483a7c15de5ce6a8d64af52bd0313ffaf21123ffad0b5006274754c6d5796
z7702bbdbd136e643a7afad253cd97aca01780510de23e5d07ead3f11705d1690d36f6924914c58
zbc0f7f9b8b3dcdf825f718390d3e1988a43a4fa585b69709fea372c569e51293ccf65304f592e5
z4d849e658d56f27c34437694235d2a0c1a69e37ae87f0f29d0e3e84fda45c5152b26d7e9e19b24
z640c81ad344840324253ec7d48406f67cc5c9e774c8ebb77680442dc5f6b78bbed6787885a9597
z6a0ef561a671063edd1cc17c38b6a91f10bd33512e84c57074de3a39dcb866527f5757e55b3984
z47814e1d3c42d6a86761cbe75ab32b444ea9aac6cc9266ec6b052a6fc9803371e8e633bc1f06ce
zfba977865415be7bd7afee390d40f2d7c162335366cc3c8c46d9efd2b5b531a1460db76aa41d06
z28474b0d7e95889c38f6c7d0c8d4a15fbbd8520319067e3519ad00e831627dca35b3cc475126e1
z0d9b3af77feb3000c215c759c8247000272a11c2597b092c8ac2cf566c55abddb768c5e9b52662
z5b03979d03a38e90a13ca781d249ec8fd280a94f85c3175ff62de69a8ea4b633ec2dd46509704c
z0cdda03f196ade10d572bb82472d0cfd7a64d7630b9b576cfb29d35f5133f0917089af415b0a6f
zea040d100c0cc22bb161ca81b746b3eb214ec4c04bcefa82e800fc5f2a13b045352fa68ebdca49
z70574d702f99c4bbfe66560baea3d725f2722fd025bbea0c5bdd7960e2f61b9fce3e330bc3af6d
zb0e79e64d09a2191fca7eff4a25b43efd16e89649473db30101a1f7226e8867f8a3b7b33511667
z211ba7cb75414571e0185037744fbeae645d602e5753777aba7a337ccaeaabf912866c9279b84f
z70eb0da8d444fe7eb54890d8ec87c9cbb81a40101289bf3a525bfe13df68a40fb9db198ce46778
z4fbbb18e2338444da527c1723f8dc89f8c05c7d1232c7125c1fe7be1c94a599e0f1b3bbd45cf34
z0dd868bc2a0c96bd81acbb9d30c65c347c62c23caa5fe8210dd502ef073c72bff24504f28abf22
zd28f91ca27719550ddd79211cc5a356453b9c6690f49bfa559f0657c839b9b4dfe478b3179fa11
z406b5f9d330dbe8abc201177ab254c95cd223b19978a692ea0745dab42ef031afad27fec935d31
zc4b6a83a49ff2fa95ceb7bf2a563aa09c8b21f9a22876cf92bc00212bce9c043fff08902521b25
zbd83cabcdcfbae30afad72016c59118ee69b8bce22f7e7f99f70e91b3176b06f57dac179eaf27c
z248cae052aa3b3c9a928de7a235f06c1648b69a36358199ee3f777f3717f2d9bc2f8c3bc998922
z6476157384af17435b44a94088b09d30e528fba0c02d53678f822bf18c63d9417b7f99e776f259
z7041737b1cf1ec6b7f47b061b32f6d9e38ad3cfd840275f9d0d6b285e23d480da31fe3faa123c4
z01efd3b53ce30d3eeae3d63253cd9c83e4990fc433a7bd7a78081319f6dac42831c5361c5d53da
z1732998a30b3443f3c0d994b7a11be8087bade98d36ee13232628f97a142ba4f699da3e34209f4
z261d525d5dd8ee4529590efe5df5391e1b41a332710d2cb31983417b4998cff60bb9c40ffa5bff
z67c79662a50f549eb40548875cd27678b5f12570c7f4f0e4abeb52882b1a51cb54efcb2680808c
z790eef5309d8398fbb08746b646e235c8665c6ca7261c6160e8d73ed4a47eb10da071b1c4d8e21
z1a755c19979f078e01b266ffaae0352802dd690b458b48032bfeb495f44839dd2f0c765a4b2c53
z152de5a967c7298bce542bd35f5ec09cc22b5054c511b2e7c6b980d5cfb5b41168e46df926fb2d
zdee1986b7c34f3be6441bc5e35a792ad7b84457c464e989631f6f3252029ab62f1e61047d8359b
z45df2860925c4a777248554344afd3076aa6ac0a633ef30d6e3a8a31ffe0a4923aee77cbd101b6
z6aacf0b0287b6302fa71221e5e3972c14d2f6b08d18eba50d68195537ce1054d42722488324249
z7db68c229dd9d210ad967ed871370174a365f47fa08c6db331c4a7628d7b5a7741f705acf9bdde
z7553245243ef87f23dd6d10db676b290430f939a46307684d294361bd059e329a25828c30fc8b1
z35c4aa790ed5e9b16c14230e772085b72c9a6100e3aeefcec40c6b94c4b94c8b25eb9ccd91fe4d
z0bbf016532fac74e49f53c18c95480f49c2a274e556376ce1e32cdec7b42e7b549e8654fa9dc57
z971c23f5a69d39f6ae1e4510957660dd169104872fc33cffa8b2b39aaafd2168aecb1b0a6fb0ac
z669b95395e31ef63cd1000352a1f160b9ad553bcc164155cacb5b7dfab040c549f0274a442682f
zf76632f226c158ea71f40d43d77d13ff70142e8d394ea195ff6e13f795ea6cf7423f9764d6079f
zf2bc436ecb8d531220a524c88338ce0c08c05332bf2af8057df615556c55899ff9c463c48dbfb0
z80d9451e8d092f86daf717528ec708a170ee46742d156e964a73039a7ef5ebe9a5f86ad6768d08
zf1fc04c9e7cc8839e05875aebc7f29f6cc3915033837ded4258fe50c82d958debd32fc570d7e17
z5a4f28a1c12a8fbc42db2f49ac23c7e0ecf3693d97f1ef7df6130221fcb8055626c2837f26de86
z9a75009d43e81bcebf55f416bbc2bbb1ff69374951c910363e37b6e433b0ef38e507a7b73e1dc7
z8f1869ecdc15b2935e84c959fba1323448c9a4dadae89e39928ae59e30db2fb7424a040508e7d9
za8ff81600f816b71dbf1d4936cb1b84be9ed63690f7aa13d5e12254ae112d53d00c4bd454bb447
ze56d51bcd2432724a3d8601e86b80d6d146b177d440107752f86a0a4f459fca6f6a00a621de0c4
z65891d7fc8156d2ef3e69fa1bc550668ea1f4f9e091ace4e1a355d20945e259828ceb56f2e4866
z400e52dc99d9aeb8e2c7f92fce82a4e7afddf6f84d02af4354ed94b693be7e18715c76b459290a
z703375ea2ffe3572e7bc71a499e718464027311760d3ec3c76efef388690bf1c0f64a00567a467
zbe2781b35d90f07251646dab8c8af1c132c88b0856b0b0c88ee9245fb3c568ca3d50c7a50fabc1
ze85f02e14d1997fc6043a672f0bfdf9a5bac5047c777281fda5b9e130659f81177a82ea21bc0ca
z634dbd2b9fa01590c68f6dc3cb54f1281a08cac4f90e9cde6cf1cac6853e50d4047e840eca7e27
z46ad65ea0816fd99dcc820c5279e869fb0ab75f022c587e4f47215098734f7e7996971c798a3c9
z07311b9c758725d27d38098723f9d0ecf9fc860ab96c9e3be4886b373b9a1d1a7579a87ead025d
z2db342051ceabd5df090008af81ad8bf900ae3ce989882a2c7ed846407401b2671417548e8dcdc
zc20a78b3da4a3219f7e6dc9f61f01d840fc80b69377e941a2cde0062c64ce630c3b0b17f6a5000
z0ccc78f6453e3646780a09508545d38b9329df35cb845222801682d260381a00adcb46a36f9e49
z58bdd6a00f5aefe35b3275dc57be838ac3c26c5cd72ea844d4d7913c97c5f56b9e2d428536a153
zc9d592b00cb9e21677cb5e9f7aa64cb593f12ee13b2a8d289d0a979d24393d534d7c66ffdbf07a
z271b77e5bf75be6134272df180544231a7142350102a4f22d5ececf9a76740c7178086d4efe4a5
z9dd68e6d0b3b508b561d338056bde16eb475e76bdead26dd281e78f0335fdd5e5b9818df816953
z1cc4ff0bde1968f7b1bc1aceb58851707d8d74675c68d305e2469d1bc7cbf7bd91060fb0c9df49
z467f104293da5ec44a4987c78b16c9009e3e22ed27b1d303b92e4362a20e6c6102087e5c2de828
zaa7fd477fbde3f3f4b33bf756d6062fb45e8d47dad149262ab5368830963efe86ffd97aec48c7a
zfd355f29be46297727d4d9208351dd60aed1d8375ec6e6d8b78694c7f199e8ce910c787eb3cec3
z59a501645068c2a03c3bd22d538b0f79141c98e4d72a2cf21956e3c9ca4952ffc47be7875b03b3
zcc238ad605d21371d106dcdf8098964d75e5168c9c60e9d273a0220a9768b6422166573392d837
z1708c92323fe46bdb1b8490bdc76f167b2f54b89dc28964ce678dc41641e62af2d0f5668246d57
z577f59e2e97abc09b67238cbdcac48bc241d973cc14f814f38d6c27635ec77b8f43c88c074ea37
z044753a0a11d5578cbd116845878b97557f5777ba1d3495f59f4b43d2514967a81edec96f1b8cf
z0cd92585a6f90fd6ab4b15b772d6d9ee9275c5f4d0337eec4b8c3bb0edf422c63f0979687ff800
z193c32ab2179a3dfa51a41930c89db210931b0d1f556d329c86a8fc212d0295fac01758b554c51
z973504be632ee282f6add4a6e334ae0e13dfbd125e5270708e79067c22cbdf3499ca0c90cc2963
z1dddb69fb86d6bd74f8a7698c5654af174d6305d610230fac0bca6b15d5ccb611051cfac5dbaf4
z4118122ca669805d6c01bb914c0b175a59c7e07bd0531d17a126df06cee784755e562e4fe05b77
z94080fbd6c95d562a57a53fba9dcd3a418bca1f296b9ca1af4928c60575c992aed19bda13078b7
z78a5980e11175d327f02ea737885ea25a443d9888983e290625891e67b3f08b77bd6c2f0cdb670
z7703338865160e75d0ed30cc700493e7234585be226b15a1be4a9145c795b0a8bce07e973ed628
z2277b007fa165a5758ed9c3df14168675adc095886cabce151b8de60977ad94678f1496a98cee2
zc38532eba0089beedd395f9c031d92341c5148f904cee7a7f3765d0974c5cc9a248ec1147f603d
z8536dee0b6ce085cf82fd9181c2e2dd9bbe654e365cd4a8f709f890c863dcaf68970e18fa6931b
zfddf33061699c11a6dc3f51a1f70ea3e86437fe454f27958cb0c71a6d5bb2773bf35e02c16f8bd
z8b7dde800ce30739127b0c8312700d5e996d3fed849916a495eeb8d4f373e9489ef77e66d19143
z10fd448f60358478dc5a517b5e2e2ea2c6776a33cf3e2df4ec402036e7a5964178273ffeeb2457
zc714e5c9e35c76aefc88c6d8523ec997d89cb865a3247aac134e6f819d5a0e22cbebab7a7304b2
z4b13a3392f5d5ba6908bf48c572661d8f04c6489e7166388c99f6852469ed4f19a8123c8d13172
z51ea32eabefde26c7aadce71201fb333d3ef816341cbe782288c94df66750e310b435cd800a5f7
z19e62d35a084f9445114c9017f4693844e7d3b8bf67c2326f3eb509dd190587df06b60c8750e04
z23558222cc57db17f7632a2e31dd447808174bbf0a3f5e4cc55e9ffe83cd6fb6aca6e46813a74d
zb800ff5dd8c295ca80398385f0c9437c9aca279bb30133fab4f7d3c64e4fe09fa480577aff07bd
ze9ae328ab5cd9331ae67351d98373ee1f58bdbda08dd33fb9f7cf3dda4e09ca5b80e3b060046b1
z1128b61ff8cdf59e4fb9a17c6edc5a2ad72b63db6361d072be6e8f55ab0cd56f83f135c4958c23
z81699b83004b118b5a6ad09e1cca071dea7c80dddd588aada83974840e3c5d73b9d3e9b7cee79f
z8712ce8134cf84f4fe56ee41834eb36e1ecc46213f69a92211bf4e051da727d5254111991f510c
zaf419872d03e28c82848ddce0a880d0e7f440b80398e2984877b3d8eb999777aa6bb015258e6a1
za9ca3b9353dbfc37f8ece3ad2b5dfb45ea49f4166bca2c27095c01e8e545241a45f0aa01a01217
z8285c109f08f21f1487e5b3b52fcbd7080c7a655cfad6420adb655921fcb1d2139bfc523e0478d
zb9db501e1ba46401fc5a200dc393957e13862d4139c55c535b95eb3e8c2ed89c3e5308b23f93ed
za04f60c1bdaf1dcdecd4973e3fe0525f276e444b71719c71d4759e5c05bdead417e143eddc72bd
za85030c1b6a45936df094dd292a18896a72b83a84cc6fc1321f24701d8a3213415d26db95f2f56
zed0ddc3b6ae405b2a96ae430987fb7d2baf78698498e9d8edfa36e796bfbc41a5a0472cd315156
z77052db84afde663fcdb743ad2b3a13ad01fbf42cd4ddab34cfaa34c1194400e6d317fbee468cb
zf7d6f449b341926ae412fa33986b1c9b86c3f9960c6ed7dc8c06aa53173e56355c93c5ea533cc4
z7d45b43b96a3931d610bdb6496e7b163ab6310c3e9920f83cc1ee498dc4f1c3202287ee90b1bfd
z70860a88ee6fb420ee60098ac6a160b112df6e1bf2eda15a9c9169966e12a8ea5865be7b12bbf7
z137fd2878e0905ff080adf753ed629e98bf1377f02e1b1d1d88e372e8d16166612a9608edb1fb6
z4f21729ee95cb7891ee96932a1d6d2571e588f2bf6003f538c44b81285bfc141e9f5504d791c25
zf08af67c2caacabb651078b6126628586c2e2aaeb22fde2385e63da0d9832d201f7e6ebe99fd9e
zd88e0bd9deaff8a27c3c8a0637b096a7114d84762985f640b1e1bdec938daf46b7230bab98ac18
zae7c77a38a73c540adb0a4820f167f1272e06c530ae615b63f2fb5d0ab9e04bd26af5b6288b326
z768cbd1e2559bb98efb7f7ea844fb0d82a17b159a05f7bc8452d35fbaa44b76a5774b74d5d83cc
z5d159f20e87b85bc58339c78f64f0f0ed2e7ca4641ec6d24ce4ab00d57fad8ccedec6a21bc898d
z5fd7505e12e51958cc1673f00cce09c125b7b19c236df05b2afd316c7777122d06f9ecc704de70
z32abb3facfb65f8fbc6a22168124281e5c8d56335a0ca2c4b1040f785d9b6b5240c1b80650b32f
zff204895c3d0e266b05ca7133f53a42bedb532c207cff373f14992402b741a20ad42e21bfcf356
z1f83b8ba0bf8902dead7cd69ac868edf2b7b89f10684895151c8a25ee76c5e1f0d3cc2f1db153b
z8da840095ecb4288ff64749e0334c2648d9067dddd6297f5d12b2a12083a2f5b34bcc6edcc0a70
z21d492bf4f456ceb3e92770b4f9ef24f16cf1527057faa940f70830352f7b950df40a3bafc54fd
zfd1c61199f647acbee3469e7c59477741adba3c28cf49afe8c8e2e2250e4c446ca5aa8496ac346
z82b11bdd3aa683f874612350e09c20b12d76e184b83df861987cddb729fe68592ad1189ba60e3f
z65be30ff2b91c04ca64117b45606909e628be4ce36e1276da3ca851c8b46c6008a365baaa62121
z03a07099f504333972890734ba9e58d0462d8bcc952f48787bdeb3ea7d52ee0d6ccaa5388843c7
z30c41129ec93acc36fed900df623c0fbb85c986419a8cfaa543b047451149df243555a5d7170cc
za93a170c3bae0fcaada44350aab0bdb01e72df9c010759091136c3515f11a11269228b1b0c452b
zcd78c6771ce9b82a946cb52ae6ad3b1d5218a3410f1802827e5fb8148d46dbbfd5847483395772
z2b79c5a2763c0954ca7c81aacd20a37adeb8604ee8e8d5501722872cb924aeeca36a265fb37048
z4d52136491e9fb7e92a95d648dc3a5e5dfb9afafad9a3eb9357f0b63e45d48b8cb2966f3c6bf92
z63476cc46a18b9de41d386c5a35ef6797820aa0ec2421715278084455d7e2a4daef5d6c0ab35d4
z337d9571901451fd273db6d92423267249eac4f8defdacf18901d705c1a240dc3f037936f54eee
z0f89d3562c8094fb6cbc3d4d841611ccbf8b6e2bf0c073fd00ce08b9b925a74040157d4ac9d528
z332c32c5c36dd88cddd80102acbbc74037bfb189eeca2b427ccd0d527536e3a6067c8a77a27223
zf884c14199a15089ecd82c8ad66afa12a500afb272e4c0b77a6846a49efff1f36813a4828dcfd5
zf3e755527668a821bd9411bb369b637344110041af0e0d602e38526035d89e10f23a36d2b6f88f
zb4c7ddb0b60091bd555048ac4607052654cf109deadeae045cdbed3d3c142fa73515339cbe9707
z5e1015253cfafdd8bd6cfa08422f65c431a6be644114b103a0665249d5c47c296aee127b0fb4df
zcdcbaa2af2012882879ce24adfbb446d1a64e379ae2afd6107cce957647e6b6522fa227698de28
z560575bd72d02fdd85f2fdac35f0da3439085d41bcfb7a164f516094abfc588522cbc2e2699bbd
z0a2d4f4b51810651ac72bcac5bbc66ee36ae01c4541f6528a7c18278e658124c8e314a39128fdd
zdf5be4bc50a296eb42ba812184c495c65a32b44cf88badf6c85e72444c9a1b4117f7824bf3b28c
z04bc73b2c42ad0b5535e517b5cf03602f02fdec74b7059b720dfeef661838d90f2b355f8fedbd3
zba61f90609b958e4ea198dd02afcdd312455a792570e9c3deb5dc284d5f2e611aa437469d4a604
zd7dec148ffdc7d205769a0d42c4a1e021787076cb948cc12e0ca6348fe46040494f6bd1679d0fb
z3d19f87c0dacb4d9b2664d18019dc9b6aef14c7cda4434c02bba3c31ed7171be076abf8ed0b209
z4535c6f8b5c9d47488dab4066c3012dd24bd0322bdfbe4a0e3e3adddcdea18a3d6ec2a369f3d56
z2821d4f065196fd62f0602790b304898e801e85cdc581cdacafc50f6069cc741f7ced8f98b1bb9
z3bbc7a72774ef173642c765e07c8d954abadb2598e4855234f4eed13cf2f8d102465d755089e45
z67ba3236d57a5c133e0ddc643e05f84d5fa5dfe006afc1c959874f64faef5e1b78e4e2e73c10b1
z9570d9f3085e1f7b6927650fa4a78ecad4c0cca86ae39209b0a9614cd486a30b7a0db725118e8f
z67debd1f407aea65fbf909080dd2b0dec39a73b4c0ed904eb443adf4c782f7765da9e3b006f91a
ze51bfb376ecefb69dddc885111e8329aafb7a0fcea3605c84986924480ab6533f75d57081ec0b2
z9b56f2ab7cdf67a68ee917c2d85f8d4e75c966d6a6128bde3f1325b37dce2164a2ca357ada819e
ze00759b39cb75a59deb567462ad7943c0f543794e5f7b1f7850611a46e348eb3a0536c32b9ca9a
zb75a4f0bfc75a1d86b0c1cc60e551dfbc02b904dd838666602d51b68a643777d72d0c0ea3cd9fb
z8fc926e89134fc4a8e1480f051b9baedf3f8ebe1e26d4915a122a4bd43a53ce2ef2d9ed667cfbf
z622d6192d93cae108672133e7254c886f5415e73fbdf8781785cca70c21b3491e551c4a3ef9307
zf37f6030afe87bfc497105a1090990f7d1d59bb87092abeaa186a3275a219fd7e31c5d6081de32
z2dab04e5688954b10da2ea7511b8d6b2dd3728ff1f47e9d7d38366e1ed161bdc455f49b71e106b
z27fd8d6167fb2a0a8c3569690b28528c7efe7d3f52024f2df298610de7dbb25095c8036a1e942c
z039b6e6333d65486a4e1d0fda6851f8c041d28241e3d724b21d71727ab27c17d92f4e528fa2761
zfa614ade807d09f996c08580420bbeef2669f76d4df87998a727aee6b1585d9695cd0bc7d35b2f
z9f6481c1f33625aeab95a63237d82310633f7a24991fc7d6d0b0e3dff15f573540d71d9d9aea20
z1c8d136f39f1062f8dbe8195d56a36e014e67d891df1c871296e190ea6f6adfdd256ece054d03b
z8887396d0bddc3da314d3878dad52f000471e631b4e0fef99b8f64cc3aa723f87388846abc0f14
z02065778a2eb2bbc2ca905de25c7f0db360df0bee17f5878ed58a7826e7a3bafdf788fbf316df1
z0950c1ba02a62c491ae11fa1f368485f8f59283fdd275ff47a8d21661981e4639d3f68f8d4e239
zf866b031f36644850043a957b51f7ebfbf691b8ed0663ac17c7a9a0a236ab284214146cd5880fa
z1ec2459e5a5262dd90d30737a3761fb769ff63e823ab2f3a929f12bc388a6087204dfd31eff54c
z754853b04b15d84c4cd14689530dbb60061a5e14583028fb55fb3717b4a2fa6a61a4c665cc7de3
z47ed6eadc3d2c7f7ef1e2270e75ffd6a3e87fafae494ed97f35905c3dda45421fab07aec1978c2
ze55805ea3f606d61f5d420ebccd14d0d5a00d4206b40b54dbede6ed3e2c3f8c121afb90f363265
z151699112700284d9ed32bcde86dc439ae3dfe858b5b0ea29a29ee37c26738f8f61c0cf5d04b92
zd3c56240bb33def6a18c129a1a7cbfc7d2700b0dacd31f4f5d5eabecbe8c4ea5c3e102e6d71d40
za7f6fd07615bd9f54d73afa9ea58861528a4aabb977b577825b3668e6a6cb07673beed9070cddb
zbf9181a927cfa8af2b32bbf0090fb364eaff6779daad873f58aee9bb7527e1d050960b4f4132d9
z943919ba8663827827f5bcbc203c18ecad9f09c1e9a1ba7a9493bf7329426f7489d2aa0257284e
zdb6e89ab5106dd3e609aa9669543b3f89df728eea015f783ffdab859f79153ae863507645742b4
zc6563867355dd3c70098b3553e5c5f4c05805cb445376f710cc4ebae4493e8422ee8a3de730088
z703d07af5f499ddd2894cf7bdd94461e430c924d949643990badf8403aed195769c7c20847ba9c
z048c397350a1c8e7ee673581a5b0f455be492fc6e72223a493380de7e92f5b678fd6a390454784
z3f6cdd5a8304684fa6aa3856cb823e735021b57e296a43144ad639a3378ab539c523159f84407b
z2e6a2d1a3e201297c03be8b2b1efc0012fa4e0f48b4efcab7ac9a251395d6f31ac3fec4749343d
z75c071d9ca0687ae6a4169d02b4f9e994b5530aa7295be306a22f1a62df1a5c909e75051c2f5fa
zc0c712239d2382edae3d8a55be298e45f425d262323787568e5a9a9241d8d1e675e63540b42721
z67ea444a296cff256d93e1196e2fea44b72bd22b2bc9a8d8acefab6adbfb4c1acecf9b166ecc96
z031da961c5330e1e6f86f8590429e8ecf6ac175d778c58cb7b115521b0d0ade732186b24470288
z1d74a8593bdb4e94e03480e8ddb86bfe70e2d8f65a37ba7cb4bfec4c9d091f5b69d3bc5c1edb4d
zd255bed714cbd1231f547099be75ef0aecce74e4fef6372390ffad14b1a91d14e9708de707abfa
z2adb1c2317cdc7e63bb5b83f07e2d032c977796bc50da53645a1fd4340d28b7571b758ed5d5ab3
z403cf3f9346980eaad587828fb0b261987e5f5e58737a10c47e168a2a0e1dfdaea21fe698d92e5
zb718be15ed2cf69640ece92e9ec9f5c2b9f94867e543b1a36eb77869d723b115ce9549f9ff59d4
z91ef0de7142f0e65937c384862cc0a8f62f1d976a54b335eeb3fa745a82c3c3e1f27f5d4901841
z032f3ea0eb0c63ab97085d4786f88127617fc1626bfcd2513396784ee3bfefdf28c876b65a2c6e
z94e2723c8edb6c80ccbb1cc05eb357bf64dcd1b53a7ab792bc588910474af361122b7ec4072090
zc098e4d0feafd948cc378262ea0c0aabb689f767c6032872077f354f619551f8320d4db5209956
zb9cdff7af1a24319ce814fc9b9029fcfb8671ebf5ed998e0765b91bab9d75f0131638751c50057
zaba94d7ff3a424974161c712e08333f85efffaf2ebd646b6247897bbae1b84641c386656eae912
zfca5246d1eadb66b078511e0add08054e7a431381880beacef6861f96d3199c69c4f5f1cf7242d
zf4a057206676dd7a4b2054093b2b37f754d99833cb9a3396ae1c998a41e9293c6a9a926429fece
zfdd12249001f8318afc12d5b87325f5864dfe343fea8e80a4889c97a31143e6f27f659f3c06e4c
z54054dcf3971b808670b1614ffbc3b28946586dc709e60de6c331648e2b14ca46f537d06844fab
zb04f94f46f5882a905c764e00312a5eaeda89bd01d14e9d2d9a7ff17fdc2e0d9575966a5f383f7
z9b8f8370e72d1672af16ffc3f2bdcff47e2f44325cb4989e2500fb9c55a22daca1f1d77628a5d5
zba3a17b7565d0f0f9b99e0949c68174e9a33280330f238b806ba77d50dd5ee9e294894d6aed337
z489f703fa83076a3c62f4860a64fbb626fa1b28d36e68b4ed28e27a9d187162051f32e667051fa
zf6e9afb613c80ea18f2d34bba9e35cb9dd50b44b9c96815fdd4fb12b33eb5e77817da89c8e6965
z3906dcf871c25917cbcb620590099cf32c23f1e27bd81fe0da9749cbba9ea269a8446de3e59dd1
z03e137df5f935a17dbfa69bbe23aee1c1172ed708308ae25b5f756b6ac92a60f9c8cbb30cbe4f4
zc72928f056526c74d455ae88fb55f8105ad9ecc33538d44f2bdfc34c9cbb7e06a8ad0e9710f429
z4bf1dda09a1ea220fb6bce0c570598b39ee5d7115ffafe6df1ed6870c0bd39d73637ebf07ab77b
zf671939d92af888b5ed1bc65a9805a55426d2e84c1835546353938bf6f396f44a33b3867f9b563
z5588a5b4aaf4f2c1aa5238255dc16cd90d370b5597aaf0d80b9841f40c8516e21af95aec4aa80d
ze3e9b7907fb39d17f1f9bab32cb1632a19024ed8924236b0b7de674b08602e1060971dadbb95f7
za6adb599feec47083e8cf885ecb6a7212b07b076b1fa03042c9242abdbdcab2fd1188c42234683
zd53e379726698a68426f178398b6b981e4badd57d82a1704f635d648227b21b851cf4893a9ebc0
z60a96ada1d032847c072aab3263d96fd9524950e10b93f9618923009b8ed504e83cab2882c4690
z6506300f323561ef1ff9d5bb688436e6b98d65cd1a40dfc0c3c93114bf9bc2896e916bdf508671
z8f71296111789befccc4df379da8bef3e1cc35a9c5add918cbeadac0df4acfb993a7ed08865469
zd01a4a19e0452b1cd53f2a5cfe8b36d121168f6276ad038bbaf9dbce3766696e8e7ad540f200bc
z1d75f377d7ce5b7ae78f214decce50061db4d96c720d950c7aae7e11a40df588e16baf2f467f20
zf9f2f510e63830400f4fd300529a714e8ae056e499645aaad05d5a73fd57723ab445c0cbac6260
z2b4d0c22d19d4d5dc58f593e10254557f02642a296272f640d51b3afe498fd4711478178c673f6
z4da50f2a05f2bd6d31f5cc8d314c23b78ddef9ae80b1305268fe29529248715c9fb6fa80a4761d
z72dd70419e8c4d70fbc9d2fad95d680c904103d5656431a947c5697847d45bce60486269d38cd0
zc05542ab2c3f3c700614d9a2c6e8d1d1f1812846cd8d14b9dc103ec539859fb997d4897586ac5a
z2c1b7fe362c0abc3db05bf2d5e20dff463ed8be9dddb7b183ee568762b5a9d6838a51f216e33f3
za54e92a129a0e01814c564564dade50e2a328894129382baa84b0e280e8dcfed1bc81bfe28371a
za67ac0f1dec904c48db5bc6e2764a56bc49fcd899069e112ca35d3691e1cec4575999f49cd593b
zec8ffd9acbee9247897bab071f27fff0ade7464a5ae805c0aafb2e87ce31003840ce2aa40bbb42
z901a742268a4eec2a37998c098f3bad8684e4345aff24826461eb7e969e3d973bd06d2bd542dca
z3338be9d4e327cd3e1ab84fbcffdab25ecf158eaaaab4ecd46a527b222545f07d6fd1201ef2e89
z65160290aee70b4230cc9bd6e7e6d048b6c0b70e13886743810840a491f171d8e80c031b31f00c
z6b881656c0e0a98ed13860696ed105553687635ad79ec524a13a0c5a5aac488c18acf507271689
za23a9ff317b3de721e82aef1bdd1b1da0beceb61566949a8dd644d1523a630d7777ab471b35bab
zaf933f27fd7946a1bfd35230fee5e2223aaf79116908252880b1c07d66fef3811f1da72f0c94d6
zdc236d9bb52356e77f44f4558f12ee5ec922a7eaec3229cfcef61524f223ca1eb2d20a60219f2c
ze97e1e72b16ca161dd20a63deafa80789007170f5b67906ca8308233949411c95ba5153688f87e
z9ad9a3ee2437a4574b47800bb0851d22050bb38850b084c5c51a581150b46eae003b3cd6605495
z34ece41de39f594f0f476b2cd003b0f8b70006819b5d87d43200b76108beb79f29363eb4aff510
zea75192886f6ebc478ec094570f2836a8a5483a493f7ff8dc69dda75939268fef920722f6cf090
zd234e5886464d19d96a3ca8a56995bb9955c30a6e41d3bb69ebef9b4f90ecf19d055e514236c4a
za95ab073853258a0032de8c38950e6b34ec554e8a71013f797b59f5c464ebcb5aa728105609aba
z04fdfc5f8356b49b98ce8ceab570559595931b78b2957197b80ce93f107c5525c2ec3aa8dcff5c
z73b078d26bc0b09505c8b09a7ed037ed5a712b66dad6fbdb418d24c18ba827b832af7c91d43b57
z1a299b0e323ca7c64bc9a93c83916f5470aa303389b917c4c9fbcc682e01f1334a4a7bb9cb8cf5
z809446919e586687eb25cc3a054c9d25fc00d2d37e28ce37f51517a9d331f6d31a2fd6873b365d
z89f001be3edceeb942bc0b29aafefbb81e58ec9d57598352c623902fca6ea97f38429154f3f3cf
zc47f86af1c3e3e22b7c0a299f63eb26ea59374f0a1ba21ac1d3f369633db3d87fe37460f267c9c
z3d725eccdbed6fe890b6c424bea98195f36282c4e61283d4ada3fe7127304ded2b61eaa1a0d455
z56207fb8eef8c5f9b8eca510f50dcc00a84d835d27b5b36f69882ff7284b57cd2f62f6d034b196
z77bec1f9e0e2c870c7dc44d0375a9c4d7c61f2275bc0dfdde293db584ae7364e026eeeacfb9247
z8c66324e1ff68dd8d8ea8369aa0ac438b655daf700a6b1c9eb900a4d148679af752e504c1ec4f2
zd2dbe4c9de39901a806bbd9da3a3fdb0e5a5752dcba25907aa9b719cd0deb7a37b51aa8ceefdbd
z64092a05667bee60e43da8ce3d471b0839cb7f150ae63e95ce6129291776232004d9b105995266
z8bfdeead875ff791843ad8134e5b10ee7d85e1f5dc8540970d7af19d435ab01eb144b8aa748a8d
zeb55d669aeb77cb0ddb37b8118a5c338b8b206d98ee6cd598cda0b89562d6182e65311351b9d23
zce5a1b0b99d7bc362ca5814db32f2c8425392dbaca39d50c543dea7e8b52d7549fcfad24cf1148
ze5769a9b6d91df0dd9f3c77ba84a7adb9f4aa4db4436985ed51f7d9ae131889afb0f5991866f12
z2668b6b471eb64a5c26cffe363788400615118e63db118a9775335c047e194d2c6873ed3243539
z3b764592ed126e62454cacfc939836b2eba39fdd680e3d6c0808392267d628367102d9dc2f3203
zbe06da52976d5f0556dacfd360504354a064055b1e11df906f2ff30631c3b3dae78b60b34aeedc
z2a771e57de569d7adc4303b3d77692e6d5686d7e339b1d7d7f85b25f951f1d8542f5e55622e302
z1f6eee2237fdc5b1dca291a56c21de4069e14310754d92b8fdcaf4b51ce359843491d759de8c9d
z06f49dd59818b5ae7a55f9d3e7c496da878376ebd72374f070cf921f6b7d9e1c989825c8fe8889
z669d342f4336c0821fb1588b10894a18ca68ed5a2a7ab7dbe49eacc18763c49b7b1f250a2312f9
zcb87dec4d4446e09902836db80699f942c75fa13723412577c37c816f4f06d413f07ea63905405
zb6d24a70da68f920ba42a9782bda1223a69728d264cd90eb60499a333e1c4de7f2ce89bd0e4db2
z67b3b381aedfd283f9d13f338f5106e09d5751934bfeda63580cf081eae089aa11d7ad3344910e
z5ffe6ffd65dac5b276fd35b6a0fd41e25bb052967edee0e8168d8bd7bbf69e791099f7d8d5578c
z4952ee8b697b82e2f3437ff5cecf640b34169e6eec54d896c394de3fd06438cfda7661aacb7eb4
zb0aaa7c4b5271799a9b37c87ead96a918f1e4c35998c11b8148403d9ffc2dc511935adfb1f5604
zd8d8369e522760f7e1a782b8cec0b7ae5b92a437322d63d4e8ae4e0ea179a8cd2fd89cdfdfb645
z7f6f4c8bbe3b2d63d25b69bc6fe1ad67c7c863b976a8801fdfaed3960300415c66df31110b5ce9
zdcecd271fce0b3b78e2c6e106e822cd1cdb2cb077228b86bb08eacdd50f7919f87abc5ebbcf006
z6d9fc9b1e1ffcf9f6b7ce5ee90fac740240cb85671aaa9f16ccae0b396211bd75b9dec7966913e
z5c1e8e8183cd9f8340c59da9f2336c75758446f3645bd2c485fee774e768a29aa797630e8360da
ze33dceb4e52bee6615625ad52492a9eca2fa7e28a6bc7d3aa456883b8e5b5d2fbb8f77a5fd29be
z03e4409e251a77fc6983c7cc681e92e7156c73fbf0273b731e15d3ebbd70dba73959f2677fe15a
z22284acf6a95c104dd4c923a071a83d10b60830682025ca91a696fd85b23c392c22000e8dc1f38
zb9ce6ab998514106f645898f53837a6b71be9fbad6de78d1069b350fe88aec67a5bbf954050d01
z14d014f69f3ce53bcff3c39e47526a291f8c4a5a226e01b7c8253a08150ba6b7bd1f9f99dd8f48
zb6f42bdce672558ca82ba907847382c66853d97ce2dbfa7f65f3c9a4ec2bb87b0932c3de9ddc70
z6db3a7ee893b628720dd759b064b73a3ef40a4c31743413c7f3e22ed669a340ec421df6ab18528
z7b88e5abe2c6ae364e1d5db582897d689adc171dd5ea2cb11fd29254056e69ea3070f64f15dd05
za8a04083300a673ddafbb5acb55f25575bc918969b54cd7ee5af303e6529b1795bd7b6cbd78f07
zceaa459c2ab0ea14f07cc683395706ca175907a66c1dc0b06cf895d9b88743db42d53c1fca777f
za35933e7e82526706d7f7066204d58a8c195fa7ce58054720326229f487bf5175eea7d32584e70
z35be0e7aa719533fcaf36280245a445fc2f69195250c0b6515ef134961e0d3d74afbd32e653435
z2c1144c7e1476de3fc50bfd482e25fc112232a0fbc1aa417e68ad2a1329e2c778e850936f9ece6
zccb8f8a37d632db4480c705c552232863c8e8b95c4182e0c3a9eecf59435ac3360f1000e799382
zd0594068667a041f64362045e9317e73444ef705ffb088bd4d271e8762bb396ad917685299c748
z7a05aba592d8ffbca0d7594a28f74bd3067d046a6008dc42348178c3010cafa7b3624c10990aa0
z387b6f07cfc2035a62d526f811009da43a40bd901422eea6d0bc06524ff9bc19b6902239d9c18a
zfa5b420aa71e8cc9e43783eae9b87be4502bc287667c7038927a4357283b39fd7017e5be1e745d
z9cab91221771a8d1c80aa7cc45de50b22a9935c566c0d939ddf9efe230c361f13c28c41e803b21
z99e46e7a5303659cd2c20a8c9a2a8d01a56cb89c3b353eb59c241d01f4f299493c95a71a66bf7d
z06c8a1c95adb713a051418a186d146d2fb1c3d5f816d188e0fcb0b3e2224c449619861ca230883
z1de69512550527768bbfd002c16bce5c854113581b7926b5253c2314b182be13246bc0710fb634
z80e5de84bf2bceea872a527840a00e8775574579d7df2c368b2ac71ed89d29f615879095192b0b
z88e597d2663970c9a9423792fc22ceec7f8369d630cf0087f3eb53ee43c9d81f239352c8327427
z865732750cfab46f9e4c2b9fe1f8c98333617bd0c8c965890b5220effe3973c5b46dffd5d5bec3
zcc9e303a0b5260ea18539742e54def183e220089a0aacd6651e21e1c18fd5a3daddd41ade7a6bb
zdae3838e1ccbfb81282080818ad4618f2688de00a8c7911ec7263f6fe65f12b9665be341dd3731
z066418810eecc444ba2676e698446c27787b28eb82a599b2db114985f306c2fb1bd901f21e83c7
za996e91521e3bf1b4961bac67dd1cff8fd5d447c0ed10a91c1ba4ad5d6bb35477b438f404daf75
z611c971412541885c6e209491fa575a3f31c98153c7399917d0a3493466de236a25da2b6dcf9f1
z86c80ff11b5d837df4516b4213640822b527bd42e0d18688fe36f3c6a91bcee437d510a72256a5
zb4ecf933d7539e015b000d6261c4f7203ad9eed1e5930517a8658124788321bb3449487d9570fa
zb7f94c01426acafc5e7763f3d10a7ec629eb0ccdfef1727f45bfde839f4c20c5188d771e405d12
z759a9f401aa4ab934ff00a61a052b611016f41444f16d38b6f6b8bc8da8350b85a82a6558870af
z01f828ed4d3322eee3403a587d7ec72413d2d6a2fff50d9c1f2e4290205340eac24f4ff351ccd2
z0cc1027287dad710f54227f8988f177c3343ced0fe1d1dc9986b0974de9722d4561181e0a9d2c5
z8ac34d75d348dd229398d6c4cf03f2d0bf1369c1e21d44d826195d0fbfa42dc8f9959988b2eb57
z941e6ea721a94799d2d70ff920e15b927ab55e9c4945240f19e90529c706b4ab99f5360aeffbe0
z3fdb1041dfae971e89431be739c95cbab3a5001da81e54e250a6dbda43656399761630a8665aca
z84628d9f5fe94015a5bd50af6b79f4fb439d601049c886fd750a8e0719a713f481918e077de43d
zc5cf2315a6255ab60a20fa103135939b679404eb1234275f5ad5a85ba088a08c336e25b08652ef
z788e0c9ac0cbdd75a219d8d89781d6a3adaccf72caef7d904427b2964ea45e64c32337fb830718
z9a4b1e55e87f421cee4f31df0594594d5bdc4ab9220e276db1927aec60dac8d80138a0233a9dd2
zacb6ef63bb1c92ab762302569fb9b60b2414e9b4d414e3a1403283e3319384bc373b3170635aed
z2e1c0f18884d46b3267ae9ed28e5439b8b62bfa24b3b4373212a19165ec3efaae5fa6db82772fb
zb06976d085390e1ed8fce0e5d245a86ae82755dd3598a43092ea0c8eb3c84798e14840e627bc41
zb46efbcb9462f7cdec26541d7b1d97367c1f9c89194df83f119b3e1abb896c7ae484826cb65237
z4fcb382fae901f261b5ef583715d9e9ddc9a0d3704539f3da70e0e969c8ee3dfb55a836fcf9bcb
zdbcb14594f1b91814f43d3992a5719a5fb6ca1921065bfa9d9d7695a3270bfdb200be90b04805e
z8c8a5bdfceeea67ec230f8e6d12587a90f22f03f6fb8b5dd4b76f1baecf5cd1624ca90ff87087a
z91b702e8fcfa85aaf51bb6fe02b63f3ee01b64794110f45ca6e7f3029e54525d1a6f7f34a37643
z213418771732674353481c54773964e08bba73ebfe0343cd760918b9d91189b992f13c0bfde025
zb19a2508b4e5b03443dcd043c8e4be80e8cc2fe7a5886128ed89a9f8058f7e28980a837ec8c7d5
z93676680ef8261dcb40e67fe22e0718f365300cef009cdef63c8250619fcada3d59511af13f50d
z2ffe84b92df31f42127371dffe25e527628e09651eb4db96e19386cda161c8fd381539105826bf
z1e6af30a14d54c7905a8a16afa06b046dadc6ef487040fa71d25e4903e58243c9624006ee762ce
ze30b66619f6a90d8ecde0df97f2a51d83f55eab7436c7c5e63efa2feb469ebf54205e269734d2e
z13fc1570a01173414381ee60fa58ae8469a26623fcfeec384df07d5d92b137366ab52c4d1e5856
z6ffe3d141a66df4d361fcc529e11599964cadaef3e8414656a86bb0f61ae13c9f17985a79a5818
z84ad313bbb5b8123eafd1336bd181813105a76e9f926ab60ebca465222c616811edf1d0b877f46
ze8d0ae7af93410ef4c2c6bf80d0d8bd6a7d1dfe9194eac46659dbefe6286525334cc7deea1426a
z5b9544a9b7cca60016199a266866dac1432373cb841b70d600fca9f0996a8000ed677dee862f1b
z8766f37cce92070cd9cc2a9a58c5178510c59066a28e868fb408996ebf64554972306a4b192608
z27806723cb465b5ebb6cbba7a1a3f12e2cbbe366dc015ba0af9af015b61fbadba7e738ebc1e870
za918312cf82da96271d64147110d6de4cae15c3ea7806100654c235a5dde63eedd3c9280ae10f0
zdf19a427f18b5b7b48064e50690fd516c1323dba5dd85eca37fc4da4d15fa92d9afcd89ca9b093
z8f165f80ea570d0cc97076e6d1bf4fe0a91eb6f508768a1c3f7b207061b08ac7399ac20962eca3
z23f926d59e5bbae7d7dfc20a48db4bcec8d06169671794883965bca720e38458ad9633d0bc3fe1
z6e4824def7bab9e49e442b66a4171f3156954c0df37ea1fda5ec9422925c92fd916a8cd41e8e51
ze585eb6737d182e2930b2ada070a2962b5cfb506fe877bd95557ecff861d93a90dad473c211a81
zf12baadabab9b2297a55da9f58b111257bd5efa2dfb6c5094282b3225aeb86e8946d7b1b8b3919
z52addc9acb232d1b0c93f0dc4164d054962084a01e2219d08f812bdd93d331fcda3039e1874e86
ze4feeebca822d3c76059066a7c37fd8bafa1a63ffba3a135e4bf23bb0649355db27b14f0d7540e
z754485e8fbfa5a5d6b9632462af3fef7c0ba09550c13cc24d837c7edf4541b1aafd0145b777a0a
zb4d5fd7eed118c42016099f7f3f5c010cf4f3b19cd7d5e85620818f0c5abefbbd8f9bd81c22ad8
ze3c708f819fdc453468ae6b23b03061670333452330401f9bec8157f18c945c579103ab241446b
zfb0a59f7125cb48efcf2c382ab2bbabf2d0104f4d759b88c06bd56192cf0fe366949aa02f7069d
z0430f61ef3f944846357b609735eb42d2191f5a52ffa44243e2ea6aa671f82b80ba33b53efee2a
z55205d6e9e16b5f7d7e71d15d172fe00494fb22440fdcad334016266a3ca2989f3cbe16ff574d6
z6d0cdaab86d37652d7ac7933d9866dcd30361b06b82a355744ad5d526748e3592a046412b4ad03
zc9bc6479d59fea6974ca5458de2611c938719063720d2e2324d45ba0529bc561d0f846dd9ec2ee
zfca8ad3e9c5bccf8afe86da8e355bc5cfaff3bf98e036da9f00ac4bfe8eb1c3a126cfbe3b2cc27
zde9d82b1c5e7747d781bdd3e382b4b86eac5526e8dd215061c7cd0874613e3e7a7ea39ab1b1c16
z8902158861f8844becbbfc7c58a1b16c17dba9aa7abd760122d9461ac5d50328b5bc4a620e290c
z24b7c4dd9dc2222d3975dbac244cbb0dd9fb0fa90466b096d7035e231c8ba48ec53d7364eb8cd1
z8df64d48dd93459b6ac5307ce12efcc19d962fc0c1c02ee19c7ea65f5d8adeb514284d912213f3
zb05150818fac3944e5d7e7a02d20b02464fd8dfc95c618a23eff16ebb698d28ea72b5a7adbdc18
zd864d365d348170f2515144029a7aee4ed69a18d28487d6da024b929b818feb27b83a8f83d090a
zb130602158f076bb1b6cc200b06c80a8784125b5e9eee54890cbb17f08580b8a8fba49e6e48c4b
ze3b0f8c3037da3154cd2b625f0e8e5a1e5c9991df35883316e692327fb49154ba127476b909bdd
zcfa86c0805a78915c0111cb4dd6a7110028c3156811f723885f7d5c7d8064903bf68bb1c075c70
zba3ae1ab5baf3bb150e542a3de2ef970cbe7ebd8a912ad9e67324aedc437a1af369ace8133bf67
z437816a58b14c36bbcd1dca47034ebd3d17aed9fea05082ea3aa205f19f7400d9129855b20f4a7
zfe169552286be8ba14766b14a4979819e3e1fc2dbe08292f65d48268096ed2f7f0198e272dc5e0
z1ab223e2f8be70a3256f317ba01dff1d0c571982eca5c2c1acd6b15fd9b96667416be846cd5562
zc2363ffeeeb22f9713f21934ced8b3d598623bbaa3c3e85aa204d9fa8858699430007a6560e7f5
zc6fac8bba524e51a741267274f54af93b2163c5f699461513479bf257b4c6a13c975bfed82a3a6
zf2c18990c21c8eabb0d675714db228c5813c8f21e927383f516e3a6ceed0f5aae0e8b12e13387b
za475b71c87623d1fd00f6542fac5409f8d13d5a733203ce3cfa1118d3c7ccb177392861e95827b
zf13bd56abd3b13d5057612dd1aa27604224a006e436fd41257bbe0a7b6c1c37a29b63d1730db32
z611c343534e18817b5c6ac97710c1583ebe165e870195b767f781137a2f9c4e767a932d1c40a9e
z74ec92540b1952a8910228473d8db7c46f190a1a52622b3981c33943123d7d518247e210223e69
z07d7de76a618548321b3a81761e319c4455300b8953e3f61839649dc0c82e3f1b8e1a260d3f261
z41cc33f9ce39c3b101282677a14a5d7f9dc016192a7a7b68ce371ead95e7462b331317cb910aa6
zf2ff1ae19048079aae9738195f233f541a59bb8e8e0bc0626de47597199577cd7da1a37f72493e
z0aebe850baf5b132c5b34dc9597ee084d49f13464d2b3ece267020ab275a58fef1efc4d8dab5c8
z373f172fcfd09d5a419287cdc97ede583081c1e9ff5b6c314a1c250927eecc5ebaeaba626740a3
zabc8d4f28e3c3608c11bac0934119e0f917f6cb0a6f9cb06484118b2a36494b79e7a9bab1ac85c
ze5c0141285c46b4bfea79e9286952ae34180303110a5bd6eeba0b1e28fc0bbf92ad4b13563f376
z2dd1b756ec5a67859a26733a97d383d240d5540a6934d974126719b9efe57990dc2db453508107
z7c5582fc08914a5e28a2014c96c8c6f5bf09f5c8dd47c1fa5a2b5029d89f5fdfeeb001ef72b21e
za882076b8ced36c88dbb4a1797e1c3fe7dd77139d2314ab05055951b97ffd082efff9cb3ad9b4e
zdf9532bbfacb05a72bc7eafe8ff18486f57694437971cb8cb0f5f3b196124ca1f4b06144efd835
z72b26e03460d759a3ff1b15c0056f8079677dc73cc46ff7fd76fc8d20bae05cd7e460fa85e47c6
z512478ccb7c056e3e0cb0f6f1ef880a5c2d21cc18d61dcab1637da521197a3c467644145f2a60b
zb0815cfdf0e50573457fa6b9e5c922204d90a76009250ca2b66a9cf76776e4850619b30cdc2fa6
z876e3a3316a7087fb2f4419448c3c08855e9e5e6c4f7d634d3dfbdc136a19f8a18a4ce756462e8
z9734b7c55b568082a867c9b6ad646bff6d2e60e45daf3bf4ac4b8c86a753c84f7609958fda5beb
zc676ea5157d73a22e6d77d80efd920554e43030a54a420a05949aae2a2215dcf4e1f8dd4a0bb6e
zc11dd82a6b87da8218d0b1f1d7ed8c0d3c27c9889c720ca2e2d8960077feeb58e37f613b0223b6
z5224f8cdfbb9e3840f002c31be8561905e3401757d1c06c495542274ded4d2ef07d207c8663dd7
z0c75d52c4e8c4b34498ea65814e598202413e450a8e306323dcc7c6345c031a89ca1688b42fa7e
zb0a00f45dcb691247fc1e37005e8ed690bfd62c043d7543c112bea6723179b3206772031c77339
z82420243aab9c0c33c4a6c597335fc2a4cead736bfa2465aa3fb8e01a09f9132a10a693b5fe048
zf60162c49dc72da6aaaad034391a629548a805f41de68da32029d1d7e488a47b9b149463bae040
z36054247added775a9d8b3ed1bac8d4d8a0179918fecd731c1af38a44fc31cbcb1f295168e0f97
z5f83fd04ab659ba6d261c397aaa48405984421c297952c8d76916fd52f5e3af195bec0a9c58137
zec3f6bc48854c3acd4172ca95c457c626a2da102517aba7d64681f9057e294e036d9026821ac59
zefdb9d58083f2820f242bf9244d51306655522508541c517545e92ea389f931fe0bfd00235aa96
z05b1e2a57cc5ebc3ddd808dcb998a742f0992f438fa12bd05f632ca67be4b60ace04b36953e924
z426bc561a4d315010fdc25b92e453078d41995ecfcc9f68d2ada32800118176b625465754d877d
z4fc8f42a4571b17b62b8c93627a539a203c1bee80879f953d178263a162e33bfb7a8ba2e4bde52
z7c3c36e495c040016412380332811c1e795577927095d74497febe856b6484cb0fb934a0e8d490
zecd3405e614d43ae3b56aa34e81b885c9c09f6b0bf2d7f9d11beac93a70498cd727fdb9f40f676
z2fa19dea820efe5d2d301f0067f76c4825ebdc8754f5eb65952fc408b43ad93c177ca1414d8159
z12db744bf66d5555ab304c35d5b9eff3fb9c576a7a890fb68428d8fb7d189169a800453c3eeaef
z574811171c130a1ae4af75c41ed15816322c0b03e26e9ef5b6e11a61a8138087d86686f7fd9528
zb372e8a79a8923b3a022f489d26b323c0fd958aade1d7f52e9464ce7c6998c416f6ad3c995b7a9
z54cb9692de2dfca5415581c487bcfe4f830d1b17315eaad9fa767d095ff7e1416ad4d9500551b4
z1ae0c50da87dee02301fc0552d7302716b1e6dd79eb9000e96315d5b73971d0934feb16dcfecef
zff10ad86f9615359a82910292edcd64098cb6588d5f87583af13ec58380ba1569c817061a76f8f
zc6fff1977184d7517806b0ea81a93d6dde2e034c1c7fff9d5ca02bd49aed0932002e562d7ff2a5
zd5761c5a7fdc267295fe3b825a826b41d7749574a6671e036f7661af9077ffe396ba5d65673a6a
z49c2bf9deaf5f47f2a40dc9053e690eb9d5a176015b4b9f5df1d5960c5c1bc1960954cdbea1e4f
z62157c08ff876ea0475b2a8516b30a0533afa3f6cbe45a96e6cc6379c84cf889f6957124cdb96a
z6ab003313d41d471e0510a24da3299ff12368b64ce53595fef8bc80b072b0ae83a3c9dc8c7264b
z87f1c04f9476224886a0b30ae9ec35fd009e6b70a0afbc8e74bef142cbfed21f276ae3523b29c6
zcc96cec10f840ddb6841df268e1f3945e2de15a1bd0277df5006b230fc3c1a2481e8e44062f3bc
z3db955c55f30160ba530168f5ff80e35493d2cad221f603eefe898007daa078047543cf8bff76d
z1eb8ee688de4d3cc8c91b32f060f5083a93ca7af43c69c94cae4aeea8ed653aa6e8f210307048f
z18c85b5852c77cd31fa283609b4c7de411e3e46c1f3938539c3079502b87882381990745c2060a
z8cf7d9a7161e2e0ee105d9119249897c859db02aa11b9421b7526990c58489cd046cbc4a25dc67
z9f37a7ddee7737625026a69575498b518ae19a84117e0190a16bc4c72eed5fc960c2e6f40309a7
z2d26a2127135a652b1c039ed8bac843ea36d0f2b3de0482ae471dcc9b1e65d743aa77de46696f6
z0813a79e234424a9709aa82757404042fa5e288ea6e3f2a0353ed7b47bbfbf3107665cccab6bca
z633e1f5b5c32812bd30e82dffed2538aed8deaaf9ab69beb96fdd11c5e0c45fc8b8b7068b209be
z887fef465620db51c9f18e0a3b53dc06dfef555b2c471270e3ed5d5fedb9a997c327f24f1489ff
z11fea166d031526daf927e5c191e48c0cfbd69c537a3bdc080c9740b1b302a3bc41d57a4c33b3e
z32220a3d39d58314190cfe08f70c9bec3432c7ab381e8b97fc3089ffe2fb48f4eba3e5a59b99e5
z8d104d385cfefeb3b302753d2a30a6d1e19c304d7093e6096fee7dccadb4a2fc09fe8f79d8d68d
za83ec2e6f784ea25af906ea4fcd51aa71b0b366384556d7403d352f7c5cdf6be9fa7e80f05273f
z70197b5625126f4395b0cf47ea9c3c9e268866f48d86706857ada1b759d3731bef5cace6bbb25d
z83addd27b8f2e84253f49ae9194a16eafaae4ace6e1aee706029100e5dd8fed4af93ea07c9dd1b
z2764ba200cd5af38c325c74f39226bce992b8c91cda93aadd00e053ee5c11d27e57aefd419e2c5
z52bd40e518ef5f96b5d68d554b03786a0ca2fd374af7265eca81119cd72d43502b45af4ebd0f7c
z8659aad33726b386db982bc2ff9de354e21a0d903de99eb4eaf30bbe6fbadeec0c0eb7f09e159c
z2c92ce53c1381dfbe1f5ff60964611a4becf7a862c2888cd8c18e4a727a049735fdca8483ea7fc
z7990b6317fbfa345b4e0ade64340885d5bac1c07a341099243a0e3fb54943bca05815c2d9d404b
z5c6341dc5793213ae043bd2031a5900eafcefd0a886762ea7cdb7171afd33b65ad020a19605e64
za79fba51bf0e921bf90f145f0d6b9e9c26f3bd80b7c0ecdbcda281a9054a1db7211308cfe0d062
zc51c0d64ea25599468a53c4564bc09e00dc2c29a7edb95ae7b13eae105bc00172db84d136a4a10
z1bf5fa057b5f55ac78f080cc910a6f42080ed16db749a3ac4f83653cc2fc3e43575dc5a5abf0d1
zdd8faca5e02976c4057915130e66623266e3a722404aed088f2f4ffcb5df6b4969edf2a102bc59
z5a0fe7589e90aa73ca3bac37f5f380819b2d0c9fac22ef4e4c5ec2c7f50f2a4ea482f72460949a
ze68585b1015ef173b1ba0b8ae2a994b2fb1b4a27ce341e009cc353439f41ec3267a17182244c63
zdef4d4c48d7f990fa1deaf9562b9aa75fec1cb653b45329f6c4231d0b40de2e70fd9c6f21599ae
ze41e67c3b9244dd10ac90c390ef27bdc4966b684894b9c9816b6e1bb8c24a2d97650d8c6e27157
zd9e1dcf756ad4cb07aa4b8e38fe70e7b190b3037d36d963293c5658d39c9be2d31f7aec0a63099
zf1bad85a68e300789037b6ca7feb473fb6c6718cd0b9782a1defb0abb6d2a58e6ff2d3ecd30214
z304fa88b4c05f19a7c162b47269d7bc997d03521c6c2a4474880458306362d6b7ebafc12d9d4ba
z7139fe3380ebebb0c352c665e331ab6cddeebf54ef347670f5076fef41710ac13c2450646ca67f
za1ae051c32a8539e50d0be823069ea75132c5d42eed00cbc5b14262cd82f67106d01b69ed8ccc4
zb10a45429fe3c26967b65fe30c88dc9103bdedc2ab090dfe215696245c5ed2443fd371ee44f260
z7fb485a1cebef5d40cf9d732c4a7e8ee038236fe13414349e88d86a694a91d7bf9510e4f9e95b7
z874756c4bbedef0ceed81752b563c387a9dbe35a731760f319c4b059c78f461a56180d8b45fe99
z78cdfa8dbebd15b2e4bc4e5a551378c9dd1d0cea7d8dfd2e9e9e37f7f21cf9f6942680e0eca7ea
z6e90db0c2f6a88f1344469139f27199e32c3a3e1e8f89fe8ac8fda3c85aa8135d0d79afdc67c23
z49dd2a949dcb38d9b9c6c9b17f6d9c33ef1c6fb8996da10d5d1ba8fd42adfcf3ac8fd5bba5510f
z9352d4d8e91aafc4ddf6fef43605f22f411bfed7c92b51a167ec4caf557f5a03497c476ca1cbc3
zde841b29f29f2e7ee87ff2bcff6303ee8866676e1926639cee810dbbdaec2c9020d0c0e9fe161d
zcc9c1d3bead89225a99cf6eaacf770039fb4fd1e216ad0251db99b172b323a4d2644c6e7fda454
z16e2bc871bdd298a68558827f18a4a5d5d27f3df827a40efbb995d6399b6972d2b5522a8bcf86a
zdf97d80268be3b457886a2d82ff3e10f06f6e18bef6a9bf1a34ad935f3c7fc18472cfac089e9df
z25a0cc949d82d63534ef8989f94b61ab4290e00653ccc8e9c4bdf15dca7d5b5b34504c9e999731
zbc113caeee4eb46db9b5d9ad2eb358c4c81e20bae29f84c19312f1a2d13d3cda46ed2ded9010fb
zde24bba66123f32363ce96c9526da31cdd833da0a3227c532780dfb4f140a712122fb44ebae547
z20437ae3b7c152eddf4b166d2cb75cc9a029ae324ffb53b4cbd293840d5811f454960e7c5a61da
z43436d52d326bc5ba9aa567c695041003cd113e7f723ce87457f73b12b20cd594bfb169ba76c48
z1a14cb0be10e3b3911952de774f7cfcc863916c7f4024a3c5825c222f20a4ad5432d52f3a2a9eb
z0279cb5c47cac86645b60b9c908afe7fc70b7b05bae39701617962fb050d4b7f2c4a933cb1dbc2
z572ef4f417463116aa15a67d8f2c69ab78d2c254b4a45e554252b87c5954570eaaa78577a3a6b7
z8f29635966b87eaa34a2c5b7f505eab85a419c62fe029dc46ec76042e3056b67d11b0efe76dccf
zcc3c98c990a6f96f8cfe1c1a1ff4a786bf9fad81000fcedf7e8d3c227c74898af939bed982dac1
z83d4ed355fdd1b3593da714fbdb28f72d5128ac7e8865c985cdbc9f63572a70398f55d3eed134a
z4f13aaffcb83e19d9a6f63afcc9ba7c165ecc0b53010a3d4b550cc79ba7a02dba974ca012a8e36
zc9d573a778e05165a4a97d7bba21839ab13cf4b843940ce2a9ccd4714d7881271c8966ccb8058e
z12aaf9b5f5ac94a7a37dc7cfce384a983066103630026b7ca13c5acae7814bee0aa8b01c9cfd1a
z69fd3501ec6ecac90146e7dd16fbf1b14307c6db42bc02b83abe4ee246b3025fe5652c61281bdc
z54f3bb21dbbe26cac820587e2f3a196cd3d5474265bcdc4add9015ee92392a80b736930c76b8c1
zcd32ada52e3218225be5ad2d9d75deaf48ed5fdd51fce5002b12cdfb784e3b9bad2ffa7a10c3d4
z5519f27b302581c0966a9adde6a68f2d12b474997eafcbd2c5868cf7f407bff6069a8be9c32ef6
zc5e9ca1bd36065e7b99ad1dabebe40c3c34048a110ef19611e38c317f5a5fafb5b588ce57ed368
zda836801620275541ba50347bb87214abf24ddfce5356a4561a1ba74a29b30f602f9e5a3df8181
zc1a6187c11b70bd9a4016751d182fde296d2d42a982b2c14728bf3b226f11e76d4e5a339b4069d
ze4968389dd1ced750ce8e95de957a0e7ffafc1e6a113ba50451c766dd579b96bdc110ec60612ce
z74c98844d02790f56ccb06ff5c942be49b69a629ed13e0c4ba3eeeff58516f5a9458c5260be8bd
z96d828380b80166d0ee9e64757bef978e907179f5361da79fb7c2684b4a0ab6936f069e796665f
z61787d69ab506383fbc036f733a48a9dba49ad96a1bd1f07032cd1484c93de9ab866ad92034cd9
z1d0d98a67f55d006fb0e719cac083f38ae6bd73d06f5eeb0db9cea61fc093ec616d8121f0155dd
z5af4f61b35a51e19e1052ad0f61400a86905f7c415378cbe1dbff96d4ddc872ae3a660be7e78bd
z3af60a176ac618aa2f568835816ab8600b9f8199e96354ca7d6f91ec31b692976f1d7c6a2dc6ad
z2cc9f1fd78c64b59c021a5f10d419ff64eb1b99f1bc7988ed0f76193819e7bbbe75168baf9998c
z3dc1a8732c6d934887fdbb37b05efe49011d0861efebde50357b3cb4e0b46042e57b304912f7de
zfb7a8846285cea3abfaa6617cdaf21acb3e5a2eac16d0fcb643874bc996168d9ba243a7694bdae
z9fd6211a904a781c3c12ab15e94d7ea62ccad38a7161a1e04a2c2622084a8f3f61e12a181a4a80
z3981a60ab930fc5350282c091e7e43bb3ae8329c5e0a38b031057075717b572e981ac3cf684c12
z1977a41c9884c9849692c5a8359efe4d1f76c2524655cb8d2bd76d01e1f5521854bf375d705da3
z9e65caeb4727f2814cca5e48e60f3267df8cff7bc8147750a03a0fec45c049dcc7fcdac5533b23
zcd7fea032f1c5a849265a6e154342e39217e9bb918b9f719dda9e1e8824213a8f4e6dcd38c071b
zaad87eb210d59198a8db60431e724099af487910f45daaf3a65e34ae7425266a90d8c5790b6c9e
z564aaf74d4ccbbe11a4291d79f94d801e69ea918027e7f48b5909cff0ccb26e9aa066be244872b
z547355acc3b750afc2b3f455a7997ea22936c8ff2bb49f6c6b746992a6cfc1d26a7fbd71e1bd12
z3c0a571ceb758e52e085597d8bcb99a288bfa5183647f152401032eb49690642a5a8f0c8a90a52
z5901f55729aefaa281da05678d595dfb045a2c44098e010d608e5575bc571e393fb45c05b4c6ec
z5c736bf50067cb1449eec10421e1b1beda8f10b675d9768387462e9a74ffe48a3d365252bb3dd0
z4b18cf5e7289f3fb2b5c1b634a32558134cf11f8e3435dfe70ac5a0020b52e852d53539028df68
z54c196ae01fa12be367113bffaaee31ac4239ec85f87bb2b853834bcb027ba98a0e319695ee486
z8f7057edbfeca6837db258047285373e05732eab07f993d918829836effd9d75dadd33bcde9a9a
ze98b862bdbe69050eaa85f854599663b662cd9224115564d123c12743d5679958d4c60a9b7df2a
z4c96e313501e43fa27c81e7c46eae2e2c089d4d7e2dcf64ebb84f6ffcec48244ecea63a6f8acc0
z9779910bd243d3bb10dd13fe5cade39ea8468e1c6b5f577348c105356b3144d7e825aef4dce1dd
zd109e91c77b5d30ac87554b573ee08e006a2bb8f33708788e28b1eb4281e4d6fd1a8e96cf61586
z112f163799a2bc5513b6103599dd26eea07d3d1ef6f5c7d2456def5591657fce51fc7d2e1be132
zff891575953ea6defd973edb6b7c1c7ec6a47a615683eb41c9560df944f036bc7bca3de2400a95
z14c0f8dc8c713edf27e9632307d4fbac5b8f0af10a8dabfedd11912663bd21265545160f5a3df4
zca766a26008df416099e2d5b02013dae5b59569d8633e4c4a560130980658e992105bec806168b
zb0e5e0fbe3a63db8b517fda7d1ad64e16adb7ceb55bdaf3a63fcb7a0c1bd40c2e65f165b5d6cb9
ze93f665003c484e7c9b89dbcf7aba2675dacbfc6226bb4a2cd3dca7f84ad6b563dc493c522d534
z637063993fef440aab71210b0865624b821f4250800d4e6d80193babba3df36951e99c13053a2c
z81749053cf6c66a708978276a6f293b785d192dd2131de360bfb8929caee0eeebfe8b2c1029da5
z148ffccbf45c6d9bfa6c81c833a214423540f4b507e38b91a90ceed2a15a5b5a7df6ed8f4928c4
zaad973b4f70c4b8fe0f89d8ecefe36d491bdddc4985fba4e5a5b975bce924429f6477355b5907a
z8b7916c74559b7c2b4d39030176d3812af888be3f565fc8d2c5fa1dd19a34fbc0e475b58875bc6
z3abdbb35f7128f32086505c277c9988a9fd4e24c65a7f16da3847fe1eb693b89b4561011af0f03
z3b62c123a2e8e273248295e951bc0356497dfbb5be6cba6320fd7bacca84d7051d3e469fb70124
z964e64faa79fc6e4f9b794ac57b29a5af91b3116ee7377498a5edca264335a5b7386833131ba3b
z72ab9e450c6e438ed0743c283e8258aa4eb1ffba890edad32ee3aadc7f54897c2011adbf084fbe
zc049203bc201cb6fbae0b6bd220f76c7c9d013d13d9b2dbfdb073c5f0e7815b4f4b7b9f8db49ec
z89cb81023e1ff6efb58a43261c1b7066a68edb65fc56f5aaf9d04a4e65cbc1372081addd98e539
z29c2322da32d257eb7af9613b3a484851d5eb2e4add2aef02bc34b2fea5302703bf2e2b302c857
z3525f1f5ea30195cf84434539b114ced82bc56ea339ec72ce2e38ae8882bc17ff74b66129ddc7e
z6ad9fb641102bb05f60b00987c5008a8f54e525a31b95a0021820600a789f021fd5b017374c8ca
z8768152584a2e3cefd0a47d8541a97d1193497669165f4a4e1d604e958638455954f14cc90427c
zf984a2cbafc6510977119253cbb9cfcf4a89110b4adf6d6fcf1de20500f8040febc80ef3aabdf3
z0cbe692f9d0df2fa2471c40b25fb9918afc1f8cf8d23af0c2f808167310243355bb3b18d8195e3
z01e614deea4db0f180e9d340429489025d2ac9668cd6e61ddae47e906041c466c1b4a9ecc4352b
z8977dde83f0680fc2c2759ac53b43926ba0a8f7fda7ff745d5c0755c02a681ae05a1c685fa2042
zdac49e4de5ae8e3aec0790ae6ec1564563a9dfb4b827632b96e3dcb47c96f5ceb0c8864c089327
zdd275d2d212799958bab1964ea19aaa166100eae41702b8989a048303d417092a6c87100754114
z682f3833cb867ed0e0e80e8ea1c816afdb4c61b662d8b38c3dcca430d7d8ea78c61e141c8ae279
z759b9395fd3c32d5a38fada221a20148811500e53bb0b5e2e5c0c2697a63a50bf2777b23e82e5b
zbf6933281a6fb39bc117bfbc66f770657eb24110dabc20aedc9e2123184331a88b8facdb0677c6
z44faeacf022a36dcfa9a4277ef682ec399681f3a9658edd160a6221bc34065cc77814ebc6827b2
z942e4644d59cd71bc3affde0d7a6cc6bf99c379c6075f2df482e54b88f9247448660a0d1bd291e
z789f54616ba8e1f274d3cd8dd746b100ca30a1195a22e116515c1988c78273746028be6b7144aa
z0fe023eaf741c0d3e74f8ae8ab44f78e6aa6450e5028bc89cae3c9acf8eb947ff4f778fac0aa28
z4aed093c7ef1e634e2c4a25028f60e8badda7a8e3034b8455f0cdfe67c3c9843d793a967e3084e
zd109b47f5696b50970c219fc6951552fa9d75ba069cfda2acb03d0b8b143629f4ae5252e346d03
z26f87e3a4d6f8a202cd6f8905d7016e14d7e02e252cf20d4c9951d337790f51ab79314ee90546b
z076585d21d4a7e2dd7d33921c2b6401ceac2ddcf1e6f1397bb062a56723fb5845d7ce065e71f47
z4243adc3468aa284d48d1ad7ad4ce9f24371d40699b9657358a80406e9ceab7c3d01bdf489958b
zda61758227188bacd37130c2f4c7b84368e5aee6cf2d6767666859b4d4c445b5fcbec91db05204
ze67a0989682373758175a3637ed138b9e630902e836617649ba4be8fc7e9813010a13e3a0a9877
z53541e085788a31c695596b9d107dae053a4ae8820dc81ea8604ce7b4dfa4ecf39dcfedc98933c
z6fc4e2ee2f088ba61fed361b1eb4f71e638fdf9518cbeed5a7277d0fac0fb3f3a52e5cecff49f4
zf940f59bea215c2ad785d3c5e219b9a7ab153b4e9cb3acc0536db483f302058fd43f46d7c2446d
zd30fce6db8dc31bcdfe8cc53e5d88f18dcbe27a709401d87c01359d96a59454383322fa69727ca
zf5bfad95a8a110401c65f7962ce77fc6dd90f609b4f31b1e977d722fcaf43c8680b8ff5a79c06e
zc166018da5359d66d7f71f332fcff89e78a6562cec33ba9e028dfe0cf6c2ad21ca89ebafad4419
z2d20253a5ed6a3bb5b58d71c908381b3022f670b333e645fdce8ed4a26db0c8b1adbe331339eda
z0800a44bfb2e677808790d823665862ff63311396917d1f6ddbf8275b8a5a8d771308d9e509cc3
z031fe726fdc650157af8426d91ea3450bf230c400920e65883300e54c5371eaa3f0636e95b359d
zf1af870d18f8af928acc240e360cb1206d088f6e5a4fa28341c357996f1e4f5527a5e72a9393a5
z7f8ca5331b126d9d5664aa78686df3d6d0277f6d2b243e445b093fa96d7ed3b7cb7bb9530ea8ca
zc1ce1789bf138dafd79483d62c3cf8fc4e39f0ea73b6351641e99eb93ea09af707bda281e76d39
z05525c3065f231c960251e3a5d700dbf1b422fb862fd476d707db8719067d0dbe8d7d79f85426f
z41db0e078ab77154abbf5af55d3e67e3c510bada6880988f9cb0da300f22aabcc607d50cf9bf29
zcdea2ae67efa2197a8e1f0e5f2b96623481d5de7547851950b09b7d4ac9d32da82fa9cb2234584
z302baaaed7e36e6dba84b904e75186721e3271d20ce7f8f21f51443b82d5b5c962f8851ddba52b
zf1fe7836a935de1103fee7630379fd4f8e0a493034696319fdbd61be8237bdbfc6e802aed79365
z0bb2f3068d286a54898f6de1c5352c62de04ec6cad768795e9cf66965373566b711be2eb435ebd
z407e13723cd23f600fd46362590aa7a95005c5dcf34613c7557dec241f6dc61b18255745303fd7
zdda7a02977d22f701773d40d5cc08a51fe76b9782bc4bc0fcaec6539c9ddda8d5148e43f0f70ce
z71c0fafbec942d9974e7539e7c3222aca6f5465fd9c08e8154bb898b102933d87133dc07df59dd
zd898156e838963d9b97a046b848a4a6eabffe6fb1f8490a2245e5f39824c9880ba19983d0e306f
z489080ef9b8a48e915b5698ff365550ca08a08ff0d2832c3ebd305d9e83fa094e2d9ecda057395
zff4d7efe5361d21e45d2b0e199f60abe0c38c736496e8aacdf3603ef1a6ff60f47ce9062855e34
z1db4e0d60172e5f1f3120f9bcd0e0ac0515a7abde639fe6387b56228f87e7919a5db514d03551c
zb3a78c95a57b1cd5592c219f160fad30472138c695a7501b7ec812ec8f9785d4dbb24ddd74af11
z6522c2485ddf115f86f2b48831e34067ebea7cee23211860bc6a76cb046f4eee2399a79bd75388
z88948cd6256cafda0a3a0dd678ca0d51a7217fbdfe4bfcbecbc7a8e3db393301d3afa9eb616945
zd27d9a13bbbf77af79b3db48674d8fbad7381f922b97fc08c1266382af4a30909e2840719d7295
ze9340ff682f7e06c1d39a7b6138299b2404445b2d7cdfac16697a7dffc0bc5896f7be504acbddc
zcff9b47b72a704fadd87ee568a776bc6796fd749ae88b9e33ba72874df7eb667a4a97c9e56cb95
z81a8a2422e8bdbfbcae5ddf62dbcf489e9600f9cfc6e3a83a9ea62c780689266520d4989367dd6
z7acff9d15f009f0c4d01c73a6462674a0971a9e52d99dbb118d26f0618ffad7f9dce6ff34a337b
zd91539c8484a14b4522025378913aa63a0be6b31fef5a94ce53a9401dc353de69bd7d5f2435885
z47b47e85bfcc60fa03855f77155973ee2e9ca176f41aefcb8b2fe930e34afab47a4e977d917e1d
zaff4bf8d0b5a5a0b359b32ad5569423a77bf64d18c47f240e6be66308ae3f1f265c9cac208fbf2
z42f2e1a0daed9b01d39a4dae832595d93647854b08ca60933e1c8f4a1b6006aabb59202bcb51cd
z0b09ec5097358f6200969a7d7b146f46622f5674d8a9dc03977ec540b6fd765ac8a70c588dda35
ze39f8850933ea619af4b6525f004de14eecf0e844af9c7b0c2658c2633aa36e32525f44c5ce58c
z32f772b0e123aa3a280f7dc1ec5d6037003b927ba7038f52c5d2360111fbb46cdd30fc992ca36a
za26e563033dc1fe93da7a855f605b193135b60f25b20cfa83d6f237d71e8b54b93dacc2a1302ec
z70bb6dcb05cd4f6d475bdb8092afdaa29bebc92ced4101918e9e6ceb9fc0c68b9b3b3471c1243c
za3c74b696979b271c3a18ddef10a46f7480dbece62ea7d35df2944dc3dea76558ab029a35a4962
z4463939f1e4beeb108077cc377e1b19f896e6872bad39292bbfe2e24d3ab9d445b450cf16b5921
zd1d6c406ecd446adf5de07e2444a64c68978ad1b82d84bd47ae179287048ea621424e8106bbbff
z689a72e659865ef93c91c188a4a2f9f74049a1f6c304ce3b10aefcd417e2ca6a3b5925c8b182e0
z69b14a019ce733653ddf22e670097d2a4e62e9b6788a83830527b2a6542ff7c041ce08abb8c4f7
z8d3791bb072a46c2a41b9b944d8fe3fda9416e189c584d41c5de18c0c1d8eac3d1f731aeca962e
zcd0b0b9b79b6406b8f93cb30a304fb2c44d4081d4604679c64523af264cdfd3ddd9755ac3d5860
z1560d3d47198f5fc053bb9ad44fa335acafa0edbaec3848443563b319589e4cfdc4e522f2b19c5
z487a59f0baffcccf28d9972a5242a753ef2a4404f60ecd6931333cda557ebed86f8fa95199d4fa
zf0eb183abd38a2b5f8587d21767782bdcf4ef82a714c95e7c7d31260c5979ba81f396e567eac42
z72a995cb7ceb21763e89cfde86c6a65d2352172bc9ad92c39b9482aad3be21c7b72da3d6f7872d
ze784ed14d3c7ddee481dfac5f63f96d691383c41481197d8ce4192542f7c9b4457b6f0d922e642
zc201081a2835b6847a5a18c28b1ed91b8a6d7c538111983361a8186cd3c859db553b7d7aeaeeb3
z7bf5c051034cdbeec3ca0a04a562f530ecd041d9e4f14813badf2e60c7498c305e6af6aeb4fdf5
zcbcc2129e50aacb71945bcf97ba9fc66008fea01371c3db1e785c06ad83bf5158896cf6dd1f6f0
zfd59d8d7c54e865fd18fe464eae4f5a793ca1f99ed226839bcf63da68f67be9fc524da619f49f4
z730ac5d48d1c7a96b771983be2684562279f144574d933bd21067fde65334b19c4f31f3e38505c
zd9b6e3c646ab5a554a2946e59ad6454db471a922c7bd37b39458976d1e6ab39dd679d1c9283dfe
z9412cb8512ff918704b6438f3e1ceef6b10c0206430bf640c1925a95186ef72e20ff8accb817f0
zd9cbe4c9e77e1822dda5e3f3175318f2a9feb543d37ad947c845d9230cb0943b0d89f7359067b2
z47f47533cf07e1c5da257a9696e2e5c251ce0352cb0e11f35049202ab81dd41784d4a90ea87fd7
zf9733afc8fe5ffc5e3801593be081f0b728b79c8e996c3666278dc69ee9d686aa12e4fdd5921cf
z62ec8aedf8f8344e65b378819534940040d3a779419685565c4a83ae384fadeab8e60fde63b085
z97ed8d726a98ce97a2aa7bc558e9f36d9f59f43ad558f0b0a2a9414c3b3a0d0d919ae9cf5adae6
zec57352c206e00fab1a71a062dcb8af7a316ce2259f6d0173baf119be85ca55b17c18ad47dece1
z7e1f8b4bec1c64b4a6599b9da366177fabc4c0e3b8fc622ff94b0f6558e317ea78897c1121fe9f
z17f863b13db6566e79ee034f07fd8b73aa5b24396366d63b62e847c948925c0baaf17043ef19a0
ze60eee743bd47d653114f9cb56ca2e56036625177d4d8cf412e9484cfa48703171c12c77849d4f
zd74bed429e686c674d138aa6212cf41516608497f507317e7e2e32e08bdd27fec03160c92acaa9
zb63ceb40287242903423f58900420ac53f1f57f5fde051bc4c7cfd0a8863028acefc8da7a64968
za5be48341932919f2056d85597d359d55dd935ac5fdcec6a4bccfc66e9031f6ddcab42b57b0377
zbe0ec689650db0e9c345c716854c4060f416d12c72c281c9be6cd562284f3ae81f9b7d467affd2
z77c07cd84efa135b715b037da330a01fdb574f9688ee3e053ad7db1ade4743b1fb2dd73f59aee9
z90a5c1ae6db4e2aedad61dbb12b3300f0d37c0da1441676a55eb93c13ddb514c777ab072d4b4bc
z51e073cbc00a2cb6231f42212fb6af49216bbe53f4f89de0cad5d96a99a8a5d5aef41e1f97f923
z02474c59e6897c54e5c8cb2ee6c25ec473c265b0aa89cfe4a2c69d69c2334cf283996de16564ac
zdf8cb09154e621734aa4915346f85f8274d4b906c1172d774838bf0149268f46a6c6b320a9bec4
zc7a2ffda4f3a62e01ad3e7786529a3a42b0577092526d25558ddd762c135059842d211e6a941c8
z0844692ffd5d1a591d44d9f73d5b79b29321fcee93b0827105f4ae7b4cd6155a3fb223638d83ac
zbdbef1456b6702a7b7d4729cd1a46df29b6adb20cb1c7464a528465ed3d96dc44328b6d6dcab9f
z8525d3db8ea7d4d607861c6f90e0cb2d71d88f167ee3a4cab2f8e9010326d4092df1eae06b14bb
z66ca86368bf4c0ab2d3643bf5aacb89fa835db557bad6a7b86e732cbb6845c712ba762fd3d7d76
zcd5ac22e278a0295cadffd1d23e3bfe8362109d61f6c44f5fec16d43d80707fbfc75ab3515990e
zfaff0d7ef1bd78ca68b1c4ecfd7c3080ae29cc252a5cd9bae568194298a1fe6c84140dfc5201e3
z09cdd7c595133952cad7524b3e9ddf70261029d79eac49c7da9c9300a0fba06f21e68c06beb5a4
z5f82aaa1628390a65c437cb54d02183db4fc60d66527105fd0de4c96742fc7d78a023bdc4ef14a
z66df1b57f83cba68bcef4707394c49cf89f36f20cd48a0625a8368f05512443a444b3b288082c3
zbdc37c3ee1dec2e396d36ed6bf4aed2ccf636342c1759cb650a81eb203050ec483e1aa92e3a135
zee1f44dde443371182cb05059327bed70b13cc7aff85e32f72b42e51cbc4d563777d216e555d9a
z148929804639a6569283b91ac926ed600f257b5b7c3166b7d6f06762733cf72850ab85361a3e26
ze53162bc5bd5c8037e4f19edbec93f9a110feef48c655a6c346e51b73d05d9d3656120f9b5fda4
zb08adcc3b6eda51ac9992c48e13e61e16ac2175c81ca2aac7daa1b2cf2f25f9ee17c9fac50adcf
z07ae4bede922e34d5be68847f936526080e175b107fd5216ab73379b3b55641d80cbf62a735407
z9af5e50404bbb1b31f6817f5c4e534a872b995e8460763dda55a5664d69eecd3ec3cd93475665e
zc0798b9ad5b9e83dd7c62fd63829060dd4d95f5e42147b5e2b2fe1faaf535daf4bf943ffa1c13d
zb729414ae24401f01f942e95cd2a3f4e8e370e5b6d99f4ee173ee98fadebc75428da56a2ba0bcc
z2f4d13b76195955efdd12e2d19accf955796f43adc858071ad58da3b3c565970ceb85c15b6f7a4
zab372cf0cd316ef4eccfedc0a3a10ad6a7e3b5df708c2c8c73da8e49d5a35c8b0beb2f80092ddf
zd1bc1e47c4ecc257ac46c1933071e6d0bd415f9a5f240c3d5d6cd4e0cb67a442b3e213e25a7d7c
z35faccb2ce32f9afc9a75dc9f1166084855eff669684987c43fab8a9935432ef08db2d6e561c60
z6450474499ca0b0614e8d81b21daff665f7c103968594e25fce9fd4d03a9bfb61197c0752d7939
z2bae563f13722254c423993490190d9a546401ce0da5a78f3be1cd3410c28865a7b63616c97992
zfdc240931b2dfa3a3673ae49850c22b184b5e6ff69811b97542a6992aa0fecfadf4c233295fa9c
z62e88781d36923416466eb460f7a06a0540a8c3c5c3df64f1a1a5ff7be3bc26433e3b5026c497c
zf6523d247039ba6f03195197d40da465ff5a0ee0eeae2aabf819340add10d08e66216414dcb755
z757ffdd092bb5137ace8b7ef1cc9f9beebfa34809fd3d1d22868ad728cb5ab9c94ab2244cb4a49
z8832423f82618ec643c490a96d84fb298abc6058c8ec873e31f360ddb89d2bd5d5e9fca64d12fb
za1ea24dd289f9dac9b1df61be19fb02e91e117e6607298a0b7c4e52ea6d97cc5382a0de323b670
z96de7464ae7db1d0ebe7d7a46d77d4badf4cd714bd4e33004797dede26160493b5724bc169385e
zd346c53a5ecd9692c8c6f3f441fb347a6761de4301b11e2b3447f10a77fb32edd2ea83a4cafdc8
z42bc8f7f4a3e56c5a68fdecd369690769620675828d38234277b200e7a4cd9354faad1b34fd2f5
z35c718176f91d641b849f5055dba7fd220c0c52e9d394f0023785c345e1a03c58e0ff6db4f085f
z8bb38bcaf4e44d0fe41c500052333e5275ca21db96c328640b4e5978fee0ea3656cfeaaf5ec816
z9908324b7c8cc1fe7ee5d8b87ae27fa712fa0a090d254b4318a139b53b0922a9c32060f4dffda7
z3872e332a2eed3f245857066555e418c6e9ab0e6e4fc23a4d0594a2ad26f92cb4f34e6988eb695
z45e323589fef0a0b9fcd5b68bfe300a09849ca30e6079791da062b2602baa9717200e4416094f3
zfc3f7bc440ca41d239e1edb7ddf4822a9d71ff3cb47e38ec252790e67754c586561f6cdb3bbd29
zb5ed32e357c784689c04879fce3cf6c632129b5c34ca36a918b0fc9e8dc42b570618c91eb6be73
zd2c836d803dfb4d14f33d7100bd3263486282566fd37a99b2ccbe9f2f6749ea5aeb99d7631bff0
z3cbbbcb7b3fe222d845972df4fe6339c9cf89a218d5fb6504ec12b4f14f472a769e263cd4aac63
z5b28a7b005da74c7161596826efb63a85b484c9ed09a4dee4a05c077520e1fab927e50ac0d240b
z567a7378f906fd147c04d5accf434674136a81b75737ec23b6a7b0dc4d7f5308f72d458fea874f
z5e8a497528c0c750eb547f3199eb3526d7e8cc6e43f06695618d2e743a0c895bc79c60b730062e
za850061b3842cf67bd79cfe5bc9de803353c07d0e8a59555fb10260511d5c6d8848b59216572b4
za250c958473b796f03202619eb8b7799c4cd148d4548886d45f54814c9da29b017a470d1418e0d
zbf0a9dde95456fb6d23982ee24f45eb44f21c99aad1f01449cd97575a3195b0e99f09dfbb1878f
zd9fffe8c29f03acba9855088bbffb98a11713c2483319b3f247235e1b29a5d6e95c3987f749a41
z01a5eed0a2ea41b284de72a693dd066c024f11002c8d1c8bb0506d51069ccdf8b7cacec8180815
zbdc9b0915eff4b28fcea53d197bff40692a29c72edc1a8e39c99037a27f79fbd2090e59d918f01
z758ec1ffe4906aef00419d93710d15acb46e9b946a56bb63d0c348c0b4733dfcd7e918d5cabb5c
z7405eca917b7f47370f3a0bbc87396f4b57cbc79be50bcd3543a17ca9b070170fcbb76eace992b
zff6709125821db2da5f3bae31db7147bbf29c20b6cdb720ee4a130be067594c1f8116721d9d91c
zd23ef09945ce1aeff6f287c3040fb0c6dd5c77a0234ac49a21c9f1fc4f1d335f1bd5c08dfbe42e
z6e9dd6d34c64358472502e51ee0695119cee356f940dc049e63163889ba7156a576ec62414603a
z36881f7635afbb4ee1f75b7c1edf6a4202e8e4e909a8393f3f0ca0e43523ad9ea009462f075117
ze32ead68f40ae5c57f0f2b8ff00b17d803f9d7d470315d5991769eb1cbd892463ef80e24376ed4
zfcd504488a4e33d65b79c9002ce1dfa5eab917180cd0e3a9ac8aecfc4fc435b6008100c50c5e8c
za1356bc5bf172f60624bd1cdd64487926e2c8f13af6d910b1cf557e62309169c6ac912977e1125
z47cf84b3572855957462641993fbf9611927227199e865a9148ad2f3d8c13dc31eead5f0068d6a
z5705b9a705692825e4900899a77a69c84f7118e6301d2e37a416c89d1615274f68452530cc9f22
z81c5880afe0426396b2fe6c29de64c58adf55cf98c0b0f248ee570b116bbaa4abec91f1f544085
zc61639260d1f3374f52dbd3eebcc3bb9efb8fc4b9d5046cd2f4d8ac25355a65f611bec3d144391
zb243d1ac4354f8eb537fdb3631fe6e2124fd60f0cd1c96d7b5a763572b2d566badc4c2718494
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_master_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
