`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502626e6dd8cb1bda8666f0a8d22838
z9da05e6b2c0e8960a421266ad24bf866896df6da17e8f4c6c25ba42a15cf0a0eaf7abfc9788f7a
z218b09a59eebb34c6c8c4e09f350f6c502077494fd0bc7070ced08296572f336cab12160c9b04b
z36ef5aad1c3dd5fac9b7838eb84af2c2f850497eea09c94b25a33cda9e66a316d7a3c1815edadf
z2ebd906b71ced2d77774c300aed057f45ca42890a0dcae10bd776cc1a88f017d8ac37af63a5c9c
zb58e7f39058a3d1d760b41245fd33fd78e29ccac474485d863182785a2238d2011e11ff1bed9ed
zb3e284f701b532ceea0244c703c26813e7dea1b0c61a27f04ec32009816bda8bfc9c9f3908b58a
z7b864e11e504e843d6e81bc172956d9c9f9d199c385a2a80086d233f6e3e353226c5d9c7ce4444
z854882afd318b6191ba577adbf90f92755b5ae793d12ca02e409615240899a4b139adcaa1cea09
zeae3e12c5f77a6124c42ebe304026cf9fda881aba0f91ef292c84f54ea5ba47ce9503084f4df88
z00cb9d753cb33c85298d02528239f3952f942eb70c49de23702246fe7c0a54d4726bb8ec9c9505
z9cd7ec1f6c370efb9115939bd295159222194ff9b43dc14b706812d2d787410061564fd0fce8a0
z209adbd2f3477e1a37963aacd87caa187b5db37238bdbe690d192d31d48dbfc9704f1d24f3d8e2
zfdceabde93a01efedfb15eee85945a6fd8faa46273c9b844758a801567810d979ce29d46afe5ed
z7d00fbaf6f27b4dbb184837378989d89e9355dd2eb791e6904c43fbd81c550b390698384133820
z230911dff5f41604da05c5f31eeedd3d600b46ed6c0c015d0cc12f798e009e182c143a607934db
z03414221f92c1513e9120b8c993acc77230cc6f6b0a01ebd2f2714146cfdd4005b01f4e8120cf2
z49f1e5ea12969023634f42d7bedde86cc07f257bb2e4b6cb19935a10adb37912f372838bcec59a
zf21cb5fe19a5a2395cd15ee8d4d7edd14118a0ca31dd62769a03aa293eb1ced28090556e1605cb
z0ff367645cdc69fae4e90c03568a774aa24923be030a73f3c429971e9a9c14ab9af4faf6f968d3
za25380f9a4ca24c55110dd7492479cd6d8caea86eb72d4d7efb654329137c26f143ebf5e1f8ead
zd9c8049e40f9ead0e234fb09a856c28d68bad01cd846677110eb43f1e1f1e909440ced3a0c6774
z6f425b62308d8a18c941a5293b2cef79ca324dff91e073121925469ea2e506b910432e55e778a5
z673105f2a4adb60adfc732235a41965151bcf36a041b451c107b39fd1fdd3e9087f0b0e9e69847
z49c3cd634d7e57a4cd642685975f1117ceb9ad621fc93d597ff8ec3f805b438aaae58e278fa954
z470014f7c58988686303e39406d42cd29fc65a24faf02b99ff909934d9c349c228485ff1131970
z91644c3b44be82f88102f76944b0116054ce7c337d6209eafb6d3dedbccfeefe93076dfe8f0c5b
z200e0c8f35cb8612f4506e187a6e77a5799f6669225c5fa334782e9d64e37b2c24e0a5d9e0fba3
z986980f57213993f81c4c2f88692d761393a7decae37ccfb8657c420c389a9aeb0c0f8e09434e8
zb52471f4b4510afc64671afb8812c7e2a92241be0008ff94c2a7cb64378f3309c78fcb96638bdd
zc46f605b6ccf5c25b9d94be107743f66966f87e3c59f0e7d0dcf830654c66babca3a957acd285b
z679cfd798d73d0406e7e8431bd205df9ec0687429e855a04363f12cac25f0e3b483c9d3ea454bc
z358341549dd8dc01d06cb8f03e683156d68332f13a9480cd924622078bbd66a7012e66514cdeb9
z42351f7246a947241021fde421a775aea2f0f49ac0579e6c5e6b7ba4e1b2935618f828daca8364
zbee3343dd2dd66daf545c62dd8cc8415eb78f6f2047f4dac50a2945840ef2bd24d03fdf042df60
z59cea658e1ff2f233dea3588f1c5da075fe0311a37d64bb394629bae4c040be48968a97ab32833
z3fe012ecf1d6369bb2737fc8d138c67a729b3b0e0b6478e4cc4c78eb9951b8af610da402c0ebfb
z1deda839537afb2b33f8bbb85904ff467547688b40424a59243d558d4f70c386a1115ac40f0d23
z145e29135f2dc6beee836f05826fa511e0f5519d7d991d5fb81c80e3c3cf00b61a6270d1a00c74
z0a4cec107fd290e8187eb549f518faa441cd9ccaa2293c5d0ec18f56c89d8e3327bbf8ff2701d5
z3e2b03e9813af88d4622e6f4da414797a0da52f519f8c612899aa65cedbb94eef41f06cb2030d3
z019e926da0223183803071c275f277dab7094d11606bbc2447ff2a3e996a5be029d47095a3971d
zc5108c3150e7fcb7efaa6e6724eddb5f4abf8e14504dec857151c603fb1445987514842a7ab04a
z3197b1717894b31e7d81ac5a703daa203728fdf093a7bc243a50d804f12258bc017a698f427e86
z4628998935785e86d60629f4ff7c3e6be74428f9a8093d86c56fe615c72fac4274d10dad2e4eb7
ze032228d38644e714addf85c515fd0d32f5eae5b3f465047573df0d9f42270ac3408c82f7e9925
z6dc12947313ceb32b1331fe8eb1b497328fd20f480871eeb57c691ed68edb7d0d9779da88c7d5c
z8a063821c083f149f56a9ba4c7e0f74f12c3143523086a700f17941713da2418a6a7040db9e3b4
z90dec0c027d4e9052755ff1f665ff06577d7b5d67484d636ef94b89e39bee016292e7baf3ba0d9
zce4fe64329ee5e8af37a672ef0d727a639cab393fd26ef2291b35da4e4b0dfe6989a0ba612c2ac
za508717f43d4947a3951f149e5919b114f713752c93c5e95f698c03ab76a973adf376a31d0fea5
zb964a1c39d739f8071aca722ae9fe6b79d817ddec171a8277ab2c4406a6aaa878e70d36f488543
z4b0ec0f180eeb973c9b91364577efb668016cd14bac3f55a57628f08f758ae27388f1933c86383
zcc559ffd065a970a6aa9eeac080b6465238fbf97f53425e71fb27c7993facac2a3592a78c280d8
z9c434fd4fcbc391e01110a52086eaaaf63ff3a4b3fa3caa53a58947216d0e03ded1babce1180a8
z3946d58b134901b4964827704ef8f96988e9c63be3d36e2245b63237c3efd228efff36129394fa
zbc3356bd910505de06a83e7d34ada20d7a3b5a95c2e0eb85d201795e8d572e9d2f4f6d9666444c
za3db4bc10b6203948932a3cf7334f24478a38009af816184106f990b0d04b840ebb6677031d8eb
ze286115f81db2856dd1b6042be285f40c22f5c279931daa157a519eb658538cb2fc6b0782cae7d
z8334656cd10a224984e583b3d20288be4d35738aa59c2d8003c7c10f056a8346865b86f206f865
zdfde2ec3039d71f4d2c1927af898d06649f24ced95ac1db3a54b707d0e26f12766a75bacd35833
zc87bc2ef8b1935599e376c04b9270d7ba2affada688c6554a08ade730e933ea57b1076b775c255
z9277a55e37b66cdd518e318e8c31645fb3b9a9ed4cc3e1d8107c4de99f9b1d0b0eb05eec7d8e17
z74ee1f3e16e53fd18f163e5dfa6f203a60b41d936c541683129102bc2d14e54ad86fd835023525
z1b46f9d168b1b382438a59f4d9dc01014d335e628c32df0b37450b608362908475be0e6ed73e0c
zbda24f34d25f077069464c1fd2c7a4cc4d56112eaf192bab7c92b1014c333b691067038fa6e752
z5410027385921b4e1bdb949bbeab8df80dad0ba19659e5b88f88a41b0b102e3a37095f809f1ff7
ze5b04050077df6915527e918276c90666b4ba2bedb557c4decc4e79a84ff49e642f67dfd658baf
zd11ba418e431bb478ba8fcb074b5b540f5b4e747f648984b1644932814a742addf9c39dc7a25e9
ze2b5b057b49220f3a74c491f7d60ec9ecffd8ac92d10504e60b9633f800d6fc49b996fa1c3b4ad
z1e76182fe99e18eb32570db0c655399c24a4722dc240dd93c824c6224d133f5dd4407b10e52ce4
z90b2cb62b08eb954c278d9d09b1baa06e4cb5617db41590696f711c58121dcf2d9efa0826d1872
z3a316dc0fb69912d5f0677ee3fffdaf8e65af83d7485404e32e6f4ebd7e5ce2125472582d572ad
z97ee8ff922672dea38aecc94af784dd39ee6ff40aadf7e9dd6a7385bab2ca60a4c46b305de2182
z6b42276bd1b076ce7ad4a94534d14fd290da3c11a089964e614ae33e91fedfbca217369301657f
z9c46bb1fb0c49ecb541d0c4175a70a08f46371c75a7f3615f6a5b06876737d86ebb85204f36d65
z46f834e961596fd9af03ec473014935fcd4c59bc73db03051676326c58731bbdf9c163cf49fcf1
z7493ae37183ee5aba15a8297586b87811b2cd50f20686ecf5f010e070237b185717e1f21dc8498
zcbed9ed37dd2a4c4acfbf91eab68ddc4e13b174f29202cb826a3ebfd5e00aaf79a987c5c2ef9bf
zb9069cede27d5c12baecb5142ee5ee8d63c20b6f7e35514339963c8d2ed2125ad6b777674f5f73
z8f612e7cf588ed909dd215424ce4620c89507d158d604aa7a44e3587e73fcd02052fb80d4100d4
z67508a2d22df7a92d406e62a91f85e43e6a5a834404b917dd1a7a5f7c1550f15211bd8240de5fd
z8a6595d8bda522e195ce26a364e50728aa13da42807b8138622457363ed33f0ccd27358e9dc942
z5988e87043ba83199a7b953d07042873ed31c14549833046fa02023d2415a2415535445154aa6f
z877725afa6c453343350112ba6249d7266783ac7e7876a88f17993b0d09f3714abffd97abb1937
z642b19763017b0dfbcf872e628ef6786aa33af9f3a892bc237c74213208692c8344356455ad0f0
z2b26f44a147f207931db8125e657df47f96db522284e15e4ea6c6ecd9c4cb5f20cf9f313b2f860
z9e103df9a7d5119252eee9459b9ff8cc8f1080d69f2e1b44dd3a5f1115a5c56632a89799e23818
z50020a53819224435a3ea5ac4c6f0ba05492912a1d2830ac6af9ec5e5b43e136846243cedfa5ec
z715f67f5acaa5de5254187e2bdea735170c1db05b93c37ed02d8faee854a7846dd2d3aac31eda9
zc2f8b07563d6ddeb386ca3b5f6d840773cc4eb7a93219472f5a29a472c28c2c307aa4975cb3f65
ze6bbf63bc6aae392f79ec800ed6b1e411b85f7a6ce9544a7c1caf39e774fd96f52817ee584c74f
z21d052e80a7c854ebb9724ef2dea0cdd673cbc0e3a444a9c3565be315ced63762a0afe22ceebba
z6fd9fa541e888ee2e498b6373cbfa93de4dcd6567cc94af3542474f10fa232960d48622c2f67c5
z8c7314ef0c0fad6881ec3c77e4b5173706f8f285418770af5fdd875d29287760a47b750be6b88c
z0f2fe9df2e76dcf4ae522258b3cd23c79d6cc690dd80254c42eb142d3b22df5347bd2179b0d810
z1dfa9963446055baeab20e704a7b929483af297f6c91113a4624ff22fcdcff4a03925be35bd158
ze91a05ee2bfba38812c841d2d63238cb1597cac89d887318a55a796d4f2ced872d30eeb35d382c
z6977db9b8afd7c8cbdc86d8e23f60163e22983cd2bc426cfcf54820d0a3833ad80816c44a4ad6e
zfe9c89c8f713554ca4228071b56144d9327e35381e0eb5bd957483fcf481b82b7db21b23331fa3
z484a11ad2f188a564b65b6eb2f0c26638fbb4c63d21496cc7a17de37ec29ea46aeaf91c60e5310
zf24c1860f1f89125ba2630ba7b18b0374f2d28edbd4ca7ac5e6eef3c3e2b571f8f31c8f003b710
z91b62dd5213e7bc1701db1bee40ace0f5dee0b39f9dee8f7a8f890caeb00ee5192ec41c1b2dabb
z1334564e87cf3d77ee5b754027728f8dc7607c948764f46803724185c1cf51c8f37b91b1b554a5
zada2384a0b1bdcf9fa4750e86696a9d6d5c3b222032b7a4482cb87205866156a10b12b3b3c57df
zdbfefab3c902d52fa004d313f3ebf670868ddc4e954aac8aa17577c63b4585d861ffa4a13d1974
z0b0ffb4052f594170666d96a856778e0c92896a39da1d022c2767751055a9a227f6b348245be30
z42e8dcd002cfb85608a20bb0efe0b96dcf3fcf0bd0609552e2401e44ea6f96b2fa5738cb1a15ef
z7a86f6a9e1a3db31914675fcbe797a1af7f3051fc2ea716fb90592c66c9cc05bd9e42f1d0fca8c
zd376f5c6f004448d27ab847b810e00c69629cbf39c3baf676146788decd16312748f5e99f14a06
z951df591c04a2f53efbb2e68327f9b40c7adbb73190e16f7614ff6306e416d03af365bf2b8c851
zd3ab76885d9c056e28f0df8b0cca9b4d2c1f47e62dcda5735dd178ce4a322efebd7534f068e54e
z716c18d3b6046ed9e4c4821670af0635189363ef6dbce0b65f707c92c23d39bc345a86cbaa7aa3
z62ef94bdcecead19f2cc5c6e52b5a706a73694c376a5c8c8e6884ce3b601cd2ec35c16b6b36a7f
zbb1087adafeb90c8d0b9e17c69d91dbbd3f7848b5b68a197b062ec6f7bc120b44cb800811722e2
zea8012892908f1c4eac3d5bca9b52e82bb554d39e1020ecc37412bbfc63cd21a127bc6650c6779
zbc01e8e052254c0c87307de3e8ceac612c8d306b7626b6404cbaf219a3f799835b189e0f90dbe6
z63ad43f629000de240727a1b652af1c477e3739ceb63484c7781d02fbdb54cae5ea377e72b3669
ze814d09c91f39837ed1d5d2490effab7a142d6642ec562b01c18a7cc8ea81ec47e0f520c71bf34
z323c3ce5fdcb8b1980fe015dd50861804fc23d75d3b3dd394db00f9e55d305f2405699e2f763e6
ze993862711db922b3f59187018672caefc6d6b14c7ef99cdb718a1fe9764a635b2c93ea837d337
z06ae622ddd70fc55f64c9ad250111f4ef421f6d47c628c580d73156342dd8f41c2096538dcd4d7
za816be7b0717a4477c2a152e45938be433073219a905b5cbfbe5c8c540420c058150cd30c54c78
z0d59993115b7e3e14ad0b4c7a90084e5d284e3c8dc724e70c9ee52780151c0575e8aab0630b73a
zf368170c3c3d76eb5c1896452feca36cf23ed806c5a39cbb68238eb738b9375c4cac21f29f5a80
zd354f92d406c806c40332a655fc13d92dc75ab2d63211ebc4e22da7607d4fc2fceaa2948d9c376
zb5212d23fd1fd591f4fa0498ee69530352df6ce0a4096dbfbf5307f40d1f322c055ff6825e5779
zd87d642e5a4d0d0963aad7ce06543a554baa1ad56ae2c6eddd0f7e99d99380ebb8de30e684f864
z886a61cff79751efb7bc1f4b379df8f0ff546f1bc43d57da9b99e432dbfb177039cfc9980c00a3
zd27202acb0c98b554e0cbff1bc02a92e16f06baf04343ad224b87a86f2b52a3a37653163cded2b
z6246c4b777d5fb439794947ae9d9d5d9457316a72d9c23e5bc8b3957d567a5bd42be20887cc298
z7c5e4886d0e02d06b63a8f3838f06e27000cd93268ffe5e705dd2c3c88f6b5ffcb29cdd1aadce7
ze3e1c6cc1ac14d51c9320848bd7cdfc7cccd44e6e1d35dbf0554f8a4f759050979b91c48f0c3ee
z4fc251817851afce19e4b5e02336aaaa0cfa71dda6a208aafd796d467eba6ddf840cbfadf044df
zd4bc3e705e035ccf9c727f0df5ec78733d565d1a1a5228d5042aaf35482518308a05058e283979
z85f6def61c7a71d77a6ffaa837c30845e9dd3d48f0cd4d914733858a6486df860717de872afa3a
z86af09f85e18752537ba562755824c474060cf692980017cef6ede5d28d023864152f8e808a38a
z0f2b35aa1774b2a7738e441e8d3e911602a299fcfa2eb4c6624d5165cc2515a5f99c316a0415e4
z5335636fdfb7073ccafa0576fd00004eef6f27ba775396951a4876a53dbd6a7da4e3abf3a22051
z5169487ea7faf92f1030dc88786a157558f956976bdbe88359aac7b8de3c39ba013d2bcabed443
z6974befbf7477b19cded22e22feac92766d5efad2c10835247d1320ddbcdfb4411c4afe4b3b66c
z81398eb1e9112fbb4a1fa2bec0464b43faf05bdab57c69dd2b9e630c5010858071eccaea436c9e
z078e81056cd974fe9495e6289b50e7e9e258bf4e4d4232df162a1a89507a75107f682c02575239
z9d421464396dc4605dc863042ec12d955417a48f95ee1af3253b3f3d98a3a203e9b039ccf0e65b
z82e6a0ca83265533ce64b3f3040a82beb90e796fae26fa41e9043420620d0e8028e24a603b5e64
z5eda0a7bd6a85c86a161d8e6b418be5115461b88fcba63618fcba58fad75a15a4ee535c0ece93f
zcb88365574418de6a05ea7e79dab5b4e7470c6c17fce2cdd6f96085053ed7208c6aa5ad4426f36
zd1f25086902ef4f55ad7352c2c8a5d2da140ed149959b8a8643870044833d452620270b1e3c480
z1693117a5bde0f7ca419eda2bb9dacca3aed7b02a38165d670c28bb2cc495b266fbe273bc101ad
z24a2a853d5f7e71e3ca83fdf53516a99656c50ac3263d37070c1e3538d008e3198c57bac0d7a54
z0fb14c421a617d976ffd093314c4b00963f98c08dcd049dd866b68d745584a74c9e1006fe33b4a
zc5990fbdb1554fd936c85aa269fccf7b2c74f836f1c4b7f11a7c11d215171f4c8ff37018112da9
z571cff919d9f6e2f50a7a31a79f7f1a55716171ec1df90d44992879e091668dcd20924f596b11c
zb33b1a5aa58a29666fcfbb9b00efdc3c43c8aef769d6f02ba49bab3bedc55a5db08b9edd1ee2e9
zbc6f43cbf08a716d1dc5e102b1f8517b1cd48651f56fb5ecc044ac5643961db5b46b91116bed09
zc88c52bdd5804fef31911a66c57705089fb88a83c6313e6ee36f1751bdbc13f62dd9d83665ee2b
zdacbb7d013eae43a149f966995be25eea14522cb1ada30d8a831f3c8bc80d43071462dfe383080
zb0f5a1c0ced427518527a3c8baa0cb0d44a0022a521963308b30d4c60aac26a7ffae06492080b8
z24cdde86aeb18d2762b4e714c9318d7bfa1f3d494cf37dda8df82dad2591cc7b772dd6db682729
z7d68b84ecc26b1f512abb20df3cb1b54b696623a82a1f8b57852337aa82d0c8ced3cae337822ba
zbb4c24f18f41841314ae1adca11335aeb3680f1b5d8d184a0a532c823d0e10b93dc7e94cdd9e39
z429cc90aebf80dcad19cfa82bde1a703b250d59c72009574d9535c5c9689481a73edf3771db576
z8db318514092de4f1ab89aa743a0e43475541e15ffbd69ca22a7b722508aa5298423cdfa31358a
z29eff1b52b6fda03c0705b0fb6e13994dc9096fc183ebdb4a6917fab35c1529ac56ab45b9e8812
zb109e1d3ff6608b68a1baef812f83957ff5340f94a6c56f8cc7741aae506d47e92ce67c096ee74
zefcff1805aace3976871b6a22a6dd34b65a50bd91064a3db70f7d4da62a699a8ecf9ca43e6affa
z108f9b1754a18d64fcde497f8567fb87f9549eaecc982e8071ec877fd86e8b93c6a2f2589b497e
z48ba9528843557bf1984c4bf66abb247c361f60cbadb8dbc80709b7f46f37bb639c4de73a0625e
zcfcb441b34c53ebc71a1bc76f6ae767be8a4f979b349c37c53100281ca9402f92a47e17b9afd73
z6a0881d24ec66726a08c2e24ce3e123e7889d323015c854d3a3878f70f8c87d3653000000728b7
z7cc22424bde297c19f04f966d831a552fbc4c8de3150d34fa99c14b4b771a8aa7e9de594b7b4cb
z37e88f86d9d83710fd3a87cb55fe7178166cf30c3fe8224e0b6733a902dd6277fc0239540f4153
ze4f6ac843abe146afbe983259e4e1a2332c638d2a6bec0d7c995a3ffbca0fd37466dd66c50f3de
z49c5b0a4b044875c9c61c8eebec886e82eda6385d1be2bcc0281762df2ff7715a5b937d2444101
z3c0f5b509fce14b132831d63d681b30413a86d5bfcc1ef0a873cbde5aee88c1b09c7fd0a662a45
zeef2fb64105f3dd51e86fb892b3c9b42229180c2b8dc2584c392d93467fcba1a71c1a91b20d3cc
zcf054fa3a9382b35fa0c7bd9a982dceeca43814dee51f8c2c4ed4ca58f1453cc202734f5173ae7
zbf9ddd1c03d5da4d74852f0a29b1e3948cf816a2e71222da18a253e4bd0f98fc602d56d90256fe
zd8e5e4c7d14ac899e56bf53bbba47d99614ec4fec4b72097f9b6faf882b09de79dc2d53d92612f
z191927cec1413f2ae40c0357da86f2214d9b7021301670a2aae854f2c08d6425bd9193796a1cff
z49b8cf8d37a8aeb31f33abc2963d2149a1f939d317e743fc880cfcf48831a0233cfba728bc9c30
z2974d5b4c9cff43ecba8395251b1af4bafb8e4457bcb8ff8737845f229aeb33bc509426aafbe23
z26f56f71b3699dbbb61aa479a4f062bb0e42ac42489b6c6792b4041ecebd91cb880422f574abda
z2c00d8d9a9a658613fbfb8cc827e52a70093ca1b9174adb9cbf9a6675407f4d45c0a9ac6e76612
zb55a94d948ff17697acf332bcf619631313d44da010f6be04a3c10b0cadafe7718c7dfcd0ebd97
zb8c13b782103e17c3dd53a43b5f77b6ef4c128b6562b609698ddd5517ba029fcd025aebb261ab1
zaddfde820cdb61036b65b9e9558880e85f8139275f2a77d7c6cb0675ff6aa74530fa7d41c45c1a
z01226e2e173866009cdd4937e6bea8ad26de93d4274bfaad44506bae8649a172d49089613d0e37
z017cac0c1a3a935067fc64e6fa15a47d3ec253ca3861f4eaba7da8d5cd1c53098d96cd60289e24
z8cd6dea6a8ef098d195f45d7cb2a5be8cee56de7fe0c119db2bed31e33dbfa36872d709eb6100d
z98f8230926706962d4cd9bd576ba6fa44df2da116c8968f449001e64e713324312df1cafa92c20
z420e9d5c3ae329091da7690baa99ab49a4532219f416dba0b773ebafac20554194a02adc1d107d
zcec8947e57973219e88f21fd6da7b15afcbfe5843fd584321e083c4a6fb2d1cf570d6da5481a69
z76cb5ff6a151b78e61867700dfd54353a5c6b2f1f1934da5532245b3c90f6fe6780e0ea7fd5017
zdc6e9f42380c8a544b4ceb312cfad16356845c52522b40512878eeb71fb88850cae7ad563d268d
zad96b850b762616f4d70223f83d628791fcb976aa76e6b4e7245f65b0050a653339a3d3c5034ce
z91da7c1ea51b2699884ba893c1a6dd5e9c2087040ea416cc740adc177854f316b40a6a35b5ebff
z4d30430008f65ceb092d7eea19c6bae794bd6db640d89dcf96a0658a631bb4bcf7e1c31011b0b9
z53f00ad98981019a22a9b9c62894d445724bd9bf28dd6a653b6c7755e1b906babf68145a19682e
zcb81edafdef482fd55a7fc12be5ced3f4067b9089220ac60033d3190a80b0366a66e780911c228
zf05f80762c450b83146590c01f5121332d9ee1e98e4887eb6814ac8bc643aead447fba4ab5a8b5
z29196f530f4f136318aaaa8d18a029dd2db865cb7e3177cb99826a24b1c5f8360ae6e73d6dd451
z13f80e5d6e31e48110c7399ed98d97857167e7744a5b7d2a4bcaa2770c534f4fdfc858b5d33c85
z17457bdf7f5129bb7dea7c9b4367be5870c6ab4ea85f383e0b9c861facd831f88f0675d8ef0d35
zb44c9bde833b06a456d53c4184174e6c3005f04e2902e7ef04151178bfffa66bd5b153f6cec6eb
z8550d1e688cffb93687ad8914bf0b5d6f763aa337158cdcabc4dfafc8795ed4627817b24de4761
zfbf3a79ee6ab481cbb8eef34875fc6041520ba708dfdbae44f52a65108209e221bca8775026042
zb3851506792a481fc9155f956c5ae2a9c19c6779ce189af17d4444c27bca9d485b9ac5e715d24a
z705f04f71d69664948715e7476a0e110c2c3b99186b0dbdfd6144c3e141b7e1dbfebea482a6e08
z109af830f1e54222e2e249d6bb5c2c46f4ba092f70ab8b03c2a1823ca9f05948cbe89b2c9426ff
zf84452201b1da39fb27b3eeab249d8827f4a64426f026bd2ab553602bdeeef286766bee58c09d0
z5345585136b3ebe872ddee538f7917d6180e8a319ffdcf24d0352a804ddaa04ec9239e930afb20
zd967caba8165629a42beedfe7d423f1b202c16c03ab6f90f9e745aa24e71c980b0c4d2097f17be
z908e926d7e5b3c449fe16a43b6724ab3933214bc655854a3c10949480a1837761b6631bceff06e
zcc2c7cf684fadb048c2d9dc979611ed6e68cc45ff636aa364fd9b1c933f45169043a50c202a6d5
zccb49da24448674dd4ca827a95893f8fb6ae4869542662a2b2e44fe80e553093665830466cc11f
z0fb30db8d8e0152ea44bffb2b68f6a183f6085228e58cae19cb8f177d4031648f17a9698e7cdae
z6390ca455e2090194ba18f01b06ab81c6ead45e59510ab550515c06f1a78f9459216005108acb8
z142d8327e5b5d660ea8f44df8b3353c5b02626eb4e9863461512d773de3c9efa328a8d27e02276
z72e4785a19c08047d979b7318917b4f691945d0d9fd93f658ee5749f7d95b195256c95f6b7b767
z287001b7db6ff6154bf922164be8341f629ada14f0a07316c924e70a5e7dee986eea22ee36399b
z9c799e6f152a479f94bbd413c68f4d6ce10c2f0cd7613d0c649263da2d59b208a6b0f17269ee22
zc8035153920d4b35cde37737c5a39dbb6c613b41c19e562432a42d786e5370c9b19b4a1baf00be
zf926eb85cb7fab0e6d98d0b7d22f00fb5190756d5f887f7742b8e53fe5fc9e87b6cfe771fa39b2
zbe1ad07234aa1b2c9ce6e7e419b42176e376c9c80c36a67660b26a3290866efc624a8db71c8968
z12873d8727fdb565b375520149a2ae601ed470debe1b8756651750c31cedf8477ebafe2e595e85
zf3a87a4f6378844b861c331ecb598b6ea250ce4d6a30059414bc0419c40b87cb1bececf782bafa
z85641f581e776f294fcf298afd86cd5997ddd5ae46eff3abb233af4a55ee7d26ffe2520ad396fb
z55b6b2bac9000be1696eccfdbfeb32874403b43282521aff9e1f171385331539e487d482941564
z90d3ea9a0f87dd58115d4df4c8f8b265e0cfc06f9e43860694ee76f4845caa07ca34d1b5762545
z8bffd2defb1238b626d90ba33b5164e960e8422e6952aaac1e1791d8385ef0b33de9a914f90b9a
zb521f6a16a4a0240a6ecca9885ae6123fd392ff0ee9506e26caf226b37a59eceba70214654a4f0
z24014bfc9e84a0be4a3287f6fe176ac0bace118ab788b9acf5de2bc44545c6f8b3f032d353c89d
zfe4ca5a4df6db4478f4c113d8cfb32f4423a816167f27b711494d1718c0b12d0e097b08611fdbf
zbaa98b3cedfbc0f6f0b1f53fa7bf9afdb893dd30f92f0d41349744589c0a1fbbfb1bde5790b891
ze918d03efecc03de0c9011b330b514289f988a5dd7a5fb22cb0e00c25133ea45a3603fc046aa9c
z5751ad28c7a56929a17b2f424abb17ac11c6f7b36e1b64c1ea8c1c21b7064dfbaa2a02b7dd30b8
z4497e152f3e7737ffddeb8bd5ab595c5c9490b6b0d70bd1c19dd90a83f0fcd4f3302f44c2a2543
zc84ed6a9668e4a04b542f313625d9d2b154820daf302ce448313510b40476cc590e17bd3182125
z1bff6501e0e581abd8b9d42e6e89b56d2560af87688b5606f391421511367c712393fb464bae1d
z9e9ec4878757fdd154def5ade40474ce74dd469692d40ba2a43e04c96129b65e88ef2598c1f610
zcc8ff3f5e5c9c72f60c5cc94b80ac2d03799a6b276405e4a1cb75b472df7b6aa3440cb2426e66e
z75aebd5e67ed0c362da80ac2a6b6fb9ecb76eec591601ef16303bbfbf69abc562aaf90c8fd52e7
z28d047b2b9322f516c1edecc13d5962b63b4ece70fb03d0246ff0377f7d4a368d563361314f292
z62fb77ae9c5a84b6db1901138fb0d5d3923689d282a0eb5906892f12a5669966a36fa99133b495
z02c81bb271b3af5c62d7619437f72ceaaf4c110cc44232fe1692ff43c0bd142ad0eb6a6b613eb4
zccf332a587c93a3580f4827e701a27d85c250b4699d2cf45c8c5106b977123eabfb66d7ecdd9ce
zd4e3fc3c715f4fc8df380ee9d1cfef6550810dec1f74ac0ed6c7f7f28ede2fa3d7ee9784d7538c
z244b865486de4cca30fb264ba3cc4a8ba740c3a2212a1178ebfddfcc4122e33cf50bd8fd3dc685
z60f59acea556159c1183af153d9d59694eb96ea24aca38c7ca214113e93d1bd40dceb1153a8978
z98d6549b03bc602585c57d0e031240c63e9cfbe55b00b9bf9358d67d1f54fadd2e6f0eed94a837
ze02f57d05b440c1feaf37d2ff2ed15f39a5ffe1c5c32ab29e2146ed62c52f709084d1c9283f754
z63b23c9f98b5417f76cfa666cc8498ca00001bd7dd84b0fbefd4e9dc296e35336d501c4eff480c
z026054c5697f5e186ac239db91ff5e5947620abc9b24f0545e4ec40dda6b221b196a56aa44ce77
z3fb2eda07e7e8aed701e8b66094e0b909efddeec409b2118820353c60f2548854adb105d7a9485
z44de1865525d7d9004a874a800db6b518d3d0c7eec4d6114d2aa8245f9c56ff231aaa96c74ff44
z56819672138e683587758b101d6071845b74572c790d2cb25866ad7df420b67f19a2c8bde47a43
z333e67fac5063a26a0f918892edcfe8f5d5dba45fcd026e21997610e79ee07f10b693c1a7b1e06
zb5a2aa97f98b1765934573a40750b1c0766376f9f09716e53fdcbb4942fb88dbdf9161c633a1b7
zf031c2bad050769e75f25e40f7d0ec0a1d0a82718c889a36ddce96563b90e99a4ff21985ad1ecc
zf80f8c13771cd3e54a3716702e2d4ecd5129966a95f7dd2aed5040258264c251d0d9097d0abe51
z9b1396e4022d3ef6c2de45dd631fc47c63724fd3d901b03e2b23e6ef8a46680c323844da487cfa
z30c8a0a47372877a149c607aebc5c7b856b62d0e58da5c8755d3c8d45a3e704976b877b7d3a2f0
z8e642da7ffa3f7fc55d239dc4ad4f0bf783ae53793e61a560a8ec84bc3c00ddba784e4c28264c7
z8bb3b188156b023a1b106ee872e4a24b552624d7d7efb08e726bae67e066d34fec9332f97a4982
z6cb48ae67b0fe6f2ed0c888d9c53d5af5532c963bea75358365bf3897b00e41a649e79c2e73193
z6a4da845aa186ecedf51cbc2507b3defe3a953759af0d83e91158cde48eccbfed485839733f734
zb51e79538469f0be8ad3915d4a7b184e8f80b355970c024514e7eca0a0d95057097ab0aab81bad
z174f4baf57c19e8eaf759b4065116d01495ecd676209c0f151119b71df15bf7d4e26df84d158c1
z504e0537b62f3499898a8240ad5eb69f35e1298edefa70e26e339f6fe60b0107f71a5dd1475eae
ze649b074c61a072273bfd2e6624fe1253048991f137d0817d97cf43703e52c814695e21add3011
ze3394cd299c5190a5f681af0806a9fd8c517cee027c561c1c1604741513bb72da176b20e045f63
z405a393dd2690f826c85aa92f0fa8505f86e9795f3e65950469b30159c5e97851d72e4606c97c8
z91d5afefa8861255b44deb26a4dcefe4a7d8fde424e7c906d14774f37ef63539e437c215a04b66
zd61f3f849bbc0d57159f4fd9acb7ab796713ac39351f6e9734b68d59c245949e5a903860c08832
z8b4baf982ed3b2ab2ac64a169e1575055c629175796b12bc61ab10102f7588fef5fc99a1b61628
z5e2ee9c1763bfa2df39c4db2fbf8339f78e87761cc3d482580f3c4a1a011e59eeab8f63f076a9e
za5291a62f6fe573962819bcbabdd69af12ba9cf4448fd5cedb3b425c2c32bb177e7b9267e35e7f
z27530894afe3fb3abc7249697f00595dc5a71206aec1904bc38dbdf444e2afc3b33cde11b72f0b
zeb4dd91bb8f2bfe2e7c31bc93f8c37f0717f60ec73d2483771fcf176411806d526c9ef139271af
z58ec66d7925801b1005742188abee7683e94be83306842068ac43c32d71c3fe366c0e447367c0a
z6e08d4c1efdfcb69e13d93b55168fca6d84976683db20ca981cfe9224ee356c11cb2dcc9bb2498
z7f1a3dcbac90a92b5d5db15f24afe83fae57dfe85d97c42096a9cadf31af7e0765821cf5fefded
zb92e9c30b734766e190052c1032e40471fb9d6bcafd76cd140640db1c8f3a5a08dbf2cb0428264
z860fffb9b4720692a31e996941567183cdd2a6f38de1cdf60d889facddd4858ed1e6dc03996b25
z1ff9da2e48b6709ea29c8b78259ea86ee0f0a1688eca3f53c3a47657f8b537ebd6033a32239683
z2e38858e96781a8c61480bfe3f63bde3a8be9dcebd81bf731ca6bd33e775d2bed34ec084855f01
z5318efcf75abea13a2b486b5d346999a98910a26002798c794c305c9ac7e4387da373bb0423b25
z8f2b6bdff1778c6c08949655d1b44c5d2b2c9dde51504a8ae8e6eee46de891657b9d204a3c7d23
z21a1390c911ec3587d507fdaebdb484c8943f644d5a0e69d93503083a59548fc2f4bfff641ebfa
z6e1aeee8883a8252308681d1a97ff914566531e6fabc929fd8c3db845eb9d60739bc508eefdd26
z23a384f09e358ee7cd740af3476e36d47485455fa983e721d3f59c626dcd913f662adaccb14d3d
z740a22d963b1bc264b531d4cc3c7ecbee1fb1e595aebf4d4409f2e9ff4657672ba34332562a74f
z5cfb5993bc1cebdebca3ba9bc374d597d2fa0a65a0bdd50093fd8c34eacc9dcd6eebda27c70121
z671997fd7a7706623e4620b0c40a5a989f85d19275c4ed2e5e0c8cf9b42da65a9644787197fb83
z401d63614ded3142ad44f517751df9b4266280bac8c992527af81fea5107d15be8afd596626546
z4d1e04580ec685e44f8ebdbe9cb46a3727db50bbdc9dc195b3a9d410ea41bc9b1c906102aba262
z01ea2052ac3b5a6bc41f47a7403ee085492ac99ad0f5b0ee6ee232bccec849aaef23a2081787c3
z3d441c5517146b4dc620ffbcff2eba778d41549b339e13c7afc1733bb4a69ff3f852d764de91f7
z491ed8e509e0c712731b078309d3fbd32d1a4e1cab361b5b79df8112ad095f384efc9495ef944d
z3752ec45b18bfe383d0c052f0f442e269d89a8d1fafb060738f5953b9086557b4c459b5ab6a291
zce1d6c84a5033b098ce871d0cabad11334ab932001dbc3ae86c6cea4b9ef50e7ff68489541601f
z4f91976e03aa0aae8bad176378c116bcb7704f7ebc4ad4d5870036527154c192329c72db06c70d
zde37e881c2064cc2758d2966ff336323c77b6fa52180582b5c310bbf475c2576f60a9718796090
za454c0a3235409bea450896252818462e6194dd14b6ef2ef7abcbe3ee27d6210c76f7922666745
ze9ecb326f9665d56c4137cc2ea15f6c78990d72930626d68b78cca59c58c16903cf276a85280a0
zd9a82a4b9ce4539e7e649519658e4f925bf136b7d953364c0758dcd292954d5c96f35d47b0e4ab
zab294b5a7e8183a2c6ba7c676daf0dfe4114a7c47a07f25a8cb1e1c8572df1a3a28935edc4cb93
z72994b6715db520fe0e9870ea2ac83b78461c2dd8011ac86b784017cfb52978a6fe2b2f1423146
z0e110dfbd5e864899e270a7fc0707a41f600ba26418e13295f1625e14d3eaf66c05c2c22fbbd4e
z106e49ebafa6714cb161c58de32d03a2c0db97be41f38af28d3fc8fd8aa07f6cee815ff95ff770
z40f50f8ac8a25a3fe67d9580cb8ab5ffddb3ec848a138137bae5ae62ceb0c8b3161260819145fe
z1de1be58e957ae96b4152a2851a4fbeba835d2b0e642402ec5160308f4be3ac8bb8853ad3ab2f7
z00421b1ee29496d1579451ad70337e938196af13f9627742c75e53889e2d2d096cd6f1017a6231
zef1897f6ab997cade59a16fb356ce03b5cdd8cffb5b8c82cf6d3e9856d85a95ab3e5a53bedf24c
z63c50dbf63093384a974eb79e280a11d7545d0d421e28f61d9ef7751b2dd8ff14914cd11916916
z5043a4a2d02f60243879ac600b7a15cdaeaee027ed7171304192886bde25f4c14d3e8fa41ddd48
z9fb2b4ef46ce263290d0c06e49bf92a987809c0afaf5b3bf596ba7a3e0cacc64b157bc00713e03
z34acee8cb27ca0a40f3d03e6ca8cb237a4c589a145a995f46d42d2d788c8db5462142bae89d13c
z2ecb3599633992711b4aacb2a73f421cd1a427959fcb01f5ddfc77155b688a2a31893b18d82690
zecc3fa283373957a92e0474d5421d5878ab4de3f6c13b4422a832b4a11b72a8898213aef2461ca
z95907a2deca476b8d868509d4043ef0a24b5466ae805fc49f4a6793338f706bcf68876588bf266
zdbc5e9fbe2dbe1489bd08d64291481386787c9007e0c214c8f0af6df7bb08064f101a190e5d049
z9d74030859d4ea610cc32967e19d862e7f16cef1a25c23c89390b1c1aee6aa863f8228312c8516
z4eedfcb71db9e096d4887dba7bb4ca1c0812ef52a6e0512d4a4fd3c66a9daa52be342ec276d1bd
z66491489b6c306359fbb2f803750d85f7e1d0763a86fc7719b2b0819c647761493ce0d7013b47f
z67cf201e6bc983726780f852a5ff5f5917e0090765278c32ac3aa4378bcff12837ac2879e8b7fa
z1f1de43958dc4420bf34d6a7eedf040812a0d70a4a2dfc1e663e731351d4cf8cc574b32e5569d2
zf4a6925cc5d1ec61a0a8a868f5a6ebb404a23fb7096965b9feb5fd50d81ac0615f2db8b12e2af5
z17ed73be86810fa6bba0fe931d0f2ff75b78cd4b0a4d5ee149526b59195e122a1bc18a8cc21dfe
z0d7c3207d693d1d1d556e9d213e880b7f9474406541ddc97be926d7fdd148b63e9c46451c60862
z80ae1a52fc26b5545481ed8cb591119a971b39b7e6bb40b98b9419f992ea880d9ef8f00738399a
z66bbd5c53cb889cf77ba102214781016125e45044f17f74a07db952bdb7574584cf190820b56ff
zf6d1328b9dafe614a7675ee0eac399f6a37fe0a388c863288602e540f45e7b1ca0449728975e28
z44e1d92a28763f3eda97d72208a702c2314604e3485cc77d636a1ff2b7473f68937520f8b38520
z71f279be10014a2c098c0774b554023d37dfd295b9af1dd7679aa365475a46e1ee8b0fe4bba478
zed1ad9337a35191e9f917e9b3504de52d173157b7ad4e52e1ef097b12704d527f04de1542a8e1f
zbb847c279fbe60ba1f663364909b8fbb1b29b2ce4116bdf05af62abbbcfa2c9c91258d848e6d9c
z54edb4639a81bbd4c93b1881e807a8cdece8253346069e663d861d88daae280b4d2a8586f10b3a
zf54307e8efd7c1efb5694d894fe4a2083d909f0c64ed8ebc34627a057f15c31b68572628df6ae8
z1b32e567a44e1a6c3dac71534a127b04ef35c8141aa0b483c7f6132ecef97d489e05d12c1a03c5
z3382496c294500f04e0ca45c59789bab0f30b03939d9ba633dad394f74d4699ebfe253140abbf3
zfbb856cfee84066c0faf60d77ead06ffbcf5ca94fba9d43edb346d19c69694ab55547e12e0edff
z49ec398dd31a49f752e11149b2d27d8adeb215dde22e41eeeccbbe1a13869669121c1005331f84
z2cf8aafc7561d12cca228cc7000224206748a9a452aec8fa4cbd366b70ff2631bc8cff5631a8da
z0c7211297bd313a8866907e13e906bc5b162474f2b2b9c0bd718a5b9159cf1acd8960889edb801
zf80d70f6a5de30588e2d3ad3c31b67018181cb3113dfac8527759971eaf7f59dbe84291ba4c526
z35bd8e379acc9a06740c2172a468c8ffa4dffef6abcdcd83671476ce68dc313eb5bea4b5985d39
zdabe7da03a25cbfc89a630b23900a39908b1d777a8cbb16ad5c658b29603386e417e549fe95af6
zd38a675858518a0de8c7e499ff13bdcad2f41949f6ef55f39ac90af9a3ddbce6c51ee6fcb7d90b
z8f94c101bace4d1d10edb5834fbd47930182b9fc16134d1ff8f33f53c85b2da1eb114f7e2c90d0
zc777ed49557ab23348d1a47b6e01498fc461163da5cbe07432088aa4fc1a1e9665d97d2ddb7cdd
z6a3220bb7652a1f3abaf3856f1790a0c156de434957d82f593e3a9de7b6751c4103dd8c386094a
zedbde308c43bf40daeb59fa4be03424ee5cd3fdc876a0f1d53f037bf2e9a3c74e28914e41c0734
z46f6b68c6104b03c898fcd6c6503ab434076748ef23ed9a4bae60b7e835f6c9e25a76b07caa1af
z77b208c6cdeeced5389201d5d15b51c578c5f8de4b233919dfa6c8f56222b1ea5ca9fbf36f22d5
z24203ae13f976417429ed5735429b3e4aacfdd2a3a3f72fcaf1bda0b35dbd75d1899142fc1ed08
z744014f786be3a9d7670c7fc80a8dc5d3d0ced18f94bd88e2af04b4bb714cdcbdf00fd146311f1
zd6ad78edd233c66f04ab6c63ea306837d0494fcd395ca9d3578163b43d7fa7cd5746593a7e5770
zabd5e28d975614e6b5b63b849d649655afa0eb9a95dfeddcf0cbcf757cf006fca3d0805d6c6c47
z02e99def4f012e90a090e7367397511156410abd765894a2e98047276b57d2eda99484bdfb366b
z2625831adabc5e0d1bccdd606506b50be4d6750383be97ee771f8fb2db19e6a1de81c0d964053f
ze59a0e9655525f31d0a0a2558b175779de2d45eac4e36985751a434988acd9f055962d1d72ebef
zd8bb48098dd458672b13badb4439268760bc06f179c14eb6fa39ca7967d8f0f2bca20de873231f
z1b831c6fc01c30e2f40ed088feb291d05420c21e897d3c7286909fe56e2967a8cdc424d353cd37
z3879badd41ccd7eb6293b64322e2314bc12b7337ac488820d5a2cc31fa901c775aed0c955b68c2
z7548736de31453eac5a19ea1f0bedf2f573d3d16bf994e64885c5ab049a2112968f3fb92213190
zb759b113644dc271de09bbbecb3358932db1253fdb423525179b2851ee73c6914013cc7c1d98b8
zbb5613b6a38fb5b29ef1ee2f19d0e5a8538c8307c424682469a696d18e5d14e319b2e7fa0ad2bd
zafb7797535544e6cca5b1935bd50e62e48d7f6521e8ddd536a5c8cb32184ae66968bdc67186994
z1f9225e2a3c148feae1447b628dc05119aa4245997ddeacb0caa91d77b75ea0b05848420fbe864
z9a5ec957329cb7496f045eaaffe562dec0c4744fd716a28b52f389781ab323d7db67a90c1512f1
zafd8856887fd668a4594394d5ef768283a058ba0b79a62dcf5fc19acf18a15dfabd7efd6fa60ac
z80b1209c1856890c4175923ff4ffea4028e5089c8c95e467ec572744bcd152568ecf106a5e62c3
zc063391304a36ae8b48010c8f2974c7d5dbc651cd2381432e2344efcc4921709cb415a6cfd66a1
zb9a2726f6f248baa3550f51f12f46c9cb27bfc213bb7b5738da446aa3aecc938ffc5bb76c3aa6a
z8dda0e2aaff57d5129602392d5f89eaaaefcdc070e54b6ab9bf6b700186879a30f6e01b13ce8f2
z9f95be6bf85f6d8969481f2b7aa1f04323f041ed533a9f70fbec651fc64dbb6e04a7e31206af13
z324458cd77c3e2f61b97794648791fe8843c5f17c62b8af0f76888cb425cefc5671b086378c149
zd9b5947d28d6415b5d19760c3cb14cad7789e43dacc7084002e7281ad33e77224f1090dfb8b549
z2a524fc2c63e871ee61b01cebb4262175746928825dc316e53a42d11853c086d2e50dd14ef77b4
ze5c58546797e219e919c661f5a8670d9d167135e84eee0925c624f4124426b8ec0df92add75893
z1644e76cdd408e11b3c01a89697a80df21ebe27afe3c8a0b99c2bdc36a37590ca45dcfc3235643
z2a88ab95425efa39f7f7e2c5520edb9d6109903e16bae428ba1f3df9361eb73276a3597e73d46e
zab3da4bdd68ecdec45da16bd9ba713aa258e7ee6e04a1cad92edd542d18f2d775f4ca5d75cdde2
z7e5065f7a4c04133647bffcb1f7956c0428d52ef615e77b87431a0955f99e1379b30488f75a13e
zd6fb6b3edf3d92d58996a36c2224ff5207097227f16fca5a4146edb4a0e121f1fe59b77f9a9b36
zc12a7efcb13fa559cee9a1e3104eb53cbc6070fc808b524340e0ec396659f2076dd9d57412ea15
z010203113cb48df62ab9458d55f5c7f1258ac87b472ab9e62f93f4f430d8bdce8670b2d540e678
z1dd6eebe1c27db9b43c455bc2b749a7683fa3c75b5b3fdcdd0969cb17e51f076a0424b104de702
z564abc462e50c7ecc96ea8b8af995aad5585fd2ccb376fddba78d13117cec27736415969615886
zcfecd74791280f49b9e214845c93e0c3e23bcc117386c4e043d5db71db6b58f7a04279c4741c2a
zb56d3cc4937d8743442ae58d7fdefb401eba08cbf8da862dfa406055f7f36d42d56778003c20a9
zdeabe83c399e99add1af7bcfe341848001625c70408c8abceacb4f865463f1ac3f74f74c7564d1
zf0104d0989129cea0d31046cb359725fc32d36b9aa1e47b36269b3c52f40381c10ebf6dc16bf10
z05dc6bd46d4dbe38b3dbd4f2c2f6c6c9967d5a1272ae217f8fc6ed06d9671ab5b3319d9b7c8250
ze16e3b6d5a26000f0b0d41cab0cd740f78c0dad035c7185518cdb30227ce70de8529e35d000fb1
z7361cd077e689a8fabc12aa721450fc9e69c7d9d8f8c00012f2b9a871ec5c4200ce94bcfbc8072
z313def70b846420d0912c6fc1f94ed0fd4e19f06dff6569b14060d763ebcd99c6b7f5e34aed934
z1c3724ae913bb3e7ecc03f3bc9bfc801416bb81d3ed168078ce68315874f7fd06ff0a9c2dee436
z29c1fd525b652eed1398d8a88cc9bc0b42ac3e636f85d85f80d86edd283a4393015518d11e1077
z5774d4aa3202ad27b162093ae8bfc36c1e9792b41335c592736fb49846f5e799eda14e352433f0
zef8bb1889bb15733a87344b0055d01c38cde242fa80c7c0b3863f9ccb9db59a4ad8587072755b1
z9aaba51e4105011c53bc09dfefa083a722954cd422330108ef3b160f28ff997b408c668490acf7
z9371f6a773681e1fe3691ee5641f6bca09a028dfbb90ad15abeec0ed23a49b621fdf385e3b5129
z0f9e3f20ba148af9c0b100cf291da59744be89cd18ea3cd7c215cd978b0d88fc43a62a1052bdf3
zbf9629eb2e97a84aa65f2bdfcfbad6c101715130f45643d2ff15fe07e76b1808a4b255eb8a7bd8
za5f68b214e478e462b24b9f8138c59217e84269ecf16a38a0a79e14ce2bc4403361631d9b48f5e
z92c681bf64fb32fcd6963a012107659383370647a31fc6d7c7649d647e4164e917dab4e8e3ead3
z28233bd0976e7444ea0fd36e67720276894a9a4145f9bd3d72d9e52cd9b0ec029266ee42420a2d
zacc65e376cdf01de23122538e0509fb46271acc7334c3e6506a714fee48930e867b5ba00545d18
z8decd0f7283eb6fdfef807dc7936ebf4d3f8a2c617e8e80c4998406e35a75fc8a147099ad89b70
z1aab06980efdf4c3e987473fba13ac56b0a5e65824851448eb640f72f5731a2e24ef6b1bf513e6
z666b941c0c78d2e45ef00a62cc203b9da1fe1abc1f15223679578d81a4155813e284059809bdbb
z2d09e4523b90fbec27977b27b180e24cf5621a2d108213c4d2f336dd072b20d5cbc269f6092d07
zab6d66fe1d0173959250370dc17c1ac4933b7388f7ec25d7e2076c4d738c81f1988143e9327699
z5146376c420c2a0dd53d828698ae8c58ca16e65c33bef536346d614d897fc11df35c1eaf16f2cc
z3c37c5013bb76839d9a6e40c78148699af6b25d11aa2c29a2e19422fb7fd6bf52315f805c33ba3
zf39d8a69b32b58404aacffeb20d7c5c484d95bbed6233ae2586a67c764baff85f8fa04b7f96dd7
z65ed1db22170d501ba797540d890f48990d17103182b3286463a59754b9bbb0efc2eb81685a003
zd307556a91be60c1c95519ab8799d27b63b57f2bb55df4e401a85d305baa920e7a4692eb642cca
z4ff63788eac74d257608e335db7936d3accbe79c3935409d14f5f49cdbf4feb8c3f25c0b58b129
zac3c8062762182aecb7808b65c692fe5a29acc0ed95ba718cfb9a4416b05783ccfdc55a92ab78a
z1b5bc412e6c456aeb58423e3dcf372b8334407f1f8b7cdbee387b092c03693e513e0d5d5f6f25b
z1df9b6e7382d5b7fb7b7fa11cd87a99670e3f820579341fbf68c92355d926a9a97530ea46b5bbf
zeecd56e5adcd3b36ff519c872381ccec1cf6d3632ac8a3a6323ef9aa98a96002566a072c021d6f
zddd238d4a1ca113b0b7a3ddf832e92c977d6ef97a529cc9f94b7e98f62338038e98203b02a7e1b
z3d549dfa02b098991f0f3a661e6ebc043c8030e4108d71bdad8e1f8c758f40d3c2e3c8f8c3953f
z030eb759a3b8fd3b6147b78235ad12f2cba0a01247f9fbdf5864f324a9ef09af64979adb40382a
zc02732ee8aad5b60456cb8b2e89412e3c11a1acf506b0a71ee8f56edf9741f4eba86384bdd961d
z031cd96a15727f4514fa38c1633b31f155bd5b3d587dbc957ed14f18b58f4e4a3ac65d72f1d9bc
z43599343046b12612728da9a9a53adc52766f6e7c07d501855a75731e38e9a25a9fc187e9dfb2e
zacb158c469fbd8d88f725bf1a85ae555931677ae5dacae08ab599eb2a2218d97e3bf97eed6d03a
z43dbf587e3ac2c9b4de2e135b1c4374e3ffb14fbe052edbd483e82ee6af188597cf695b3a82216
z6f6160b4b9da20abc14d629479904d4c3bd862738ff83269292c4fe323dc64d8b488f3ac093824
z47c9fcc4ed8b70aaf6c634b1ba29394450c597f780dc093c5c067d9d7807a088e01667bd00f5c1
z940d06a36a1b0bcf327909b7ba8e19e8b713e86a66e996c1780d5b0e1104062fccc6dda94d3c11
z3ab9aea00ef39b0bd156d92e2f7f5d198795a064268037df796ee073e0504afcb0c1a2529953ec
z075e4b888a2b08836726811d2acb2171f78d6a966b536d5897044bbc047905d3616ef1bda3d69b
z88f8996777aca05c62bbd0ce49567aa03536d5a1400e3b02db0d49a59ebc4857a9602b849bf42e
zdd5e15d08c3a26a3aba1d24de05249944135de4859f549c9e51a8e0148ea1bc2590b3874ff73bd
zbc41d50306289821732b77d2f1c8aeca155d5b44f421880bfd5268549d209cff108759ff854d19
zcbb804672a823c8996290eb4957a9fc2ba716b3c91f231284cc91be58fc4c348f9a31cf313e54d
z0baed36b5e32ab64415027701e819710c81c454cd8e91cce1594a1ea000ac4109469e0f6a41a8b
z5d53583ca7f00002dc0f6af3b0d7d1da70c97bc60aaa1d5bc9d1fd20d4ce05a7fb378c223f9f05
z14aa43253a60729c3689f42ef46d17a8026e94a019dd6d5e50826a5e01fe8dbf22073586b538da
z30195fdcaeb423c4c03c624cb166c1a5304bdc24aaed669bfc33400175c5dd2b9c3270f4746898
z5ac0f63437c534c6fa4c21f3a61042647009b0271d476042e54ac2ecc40bb5d78fee311bc9412d
z5e6d5f923a3ac3ae1f5addea8c013e8331649c6b1bf85f65a30315bd69e51a8d9bbbb1c019dcf3
z55380831564aa0a304adb80978a8853cb4a4dc28b2f85485157bb374cc3e195e437572dca34208
z11f0b4259d86100224a5194327fc3e129b2247020035f25740b6db7a2d0313d676ba9f52f39a46
z4c60b99348487e1fe7a12ce479e2d8dbc0d12fc101cb550f7702738aa0df99e6457222c069f938
z97dde7729ad4f2dad347b7eb7158c6fa912966e4c8fbeed553ce8ddeeeaa8801b9cdbab28517c8
z36942a711781b4293b5808e1ce3d77936e923907983cecf28aa0e3a0954e607a0301d06a8bffaa
z9c5c87b6b16b1006b49a74900838a2130c4c35bbe3d8b61d5d8dea362a0504c3ba8fb0fe4d276d
zb773c68344f5bb5a7144d020ce362900a3eb63a0b25a063f70788f50313784dae3508402ac3ed2
z92cf1ce0ff8b6053e38886f83ea1b0f1cf948535f8fe3e294e68a4b112561a7773192286955c2d
z8f6c7f83181eb2ba4fdd8c82457aafa45df2a32c0cd27f87998a9cd37ad9ec9ff5b65c7bb552a1
zfdff2ee770e00eb8316ebf150bb08405026fea6b7d937f9938a7f6cba1ce974923cb05d9e322fa
z762b658556b872a336b4a0861343ad74b8fd465b89f0e10e28f798f3b0460dd69769c5b725c723
z869367392abdecd66dc6646b827aa8030be1d98bf5d6ada9f3c532b071508d6b1c67a65b8cbe28
z5c4dc2baeaa32064931091aaf015ed658217bf5a6900112230767b2d40df9bc5c2efcc54a82cd0
z43b28e4045b8c3679df72ed99ee5e466ba73d965c6bba3555e1c86fc3a207c59cbbcff2bfc4c0f
z87bd3083cb92989342dce64d75fc28fc997d7f7014131acd7a1ea088d0876dd2e7371dcf899fe4
z4768fa0f53b332ad13275910a7e6304e45527acb19833a780b808c8d8d1c81f0cd4326b5a8564d
z4fbdbc71d7fa76d5ac7b439b08534566f75c579e8505bdb05262ffd2ca6d42f710b4dd706c6cfb
z12593ac958df5c3f2a0ab412f6ba421805ece8d370e11cee546ad35b7431910013dff6d2af1200
z30710964cee0808dc6cc0fbc265b61a50e51e8501f0d3b1c8a40951edb27099701c050d28d2099
z5e0231eb901177bc33374ed5fbc01e16c506396d9fdcb4a771e86b7682b30367a45d2c3f7018c0
z78cdc743ecfc07ae559e1a355293e1636ce15fa4e205e5339cb7cc3367f0df68b3d76799eecff8
z6100d9874fb1040c76cd530d90763b3ec01b4d795a425cbbc47c3903b6de31ddc4fe62f9e2e2b2
zfca3c15afd6ee44378e24d8c4fafef990254f5b22fb618a38641e9f2da83078c4c04c366d01434
z2ab11964f86e4621491080a673af8a3c573a888d5fcb3692979c74af4880a5337d7d31809c9a32
z1107c0eb5290b70d112ef19a6735c25335f3c4ae8bd362c35bcacf56e04adc2a0724bff69c2c31
z175b2d0ad1d1d04bb95a0b6c768a1d55ca7d17eaa6afddb18a81ea9b22c89779f44ce14f2f3004
z12934a3bb22a37c01c4fe2970f65b8c94316e9ac5e4375ed17b1a9f546ba95d2d646978fe8f340
zb8936ec90b20d00e010b5fe9f815fbb1bad3306a87048662aa20529ca6893674d9ff6c44f39cf5
zb1db3868227f2984452a2f3968e0906aca62be9546300af612b72886482838fe014f80be2875f0
zc30ac1ce27dfc58bf833d3926ede81bd586e7eb5490c47667fc7b3b21d8ea823508c32efd6fa69
z613c5b9d1ca191bf007af07c363a48cd7ecba964f28c5d2e081059d7de6381d55a6d5c42ad742c
zea9935de1d4f915678e8d4713d399788e1e68b84f531d4351d7f1c7c772cff3de7bac5c4ce081a
z1fcb86dea8d16e6e0d00417f57b836b432eef5d5c60999fcbbc5b470c2f5781a5a4bddd6e989ec
zd41bad407699481f0c1e16ba099bbe1a8c47bb23e8066073a1bc662f3d85eeaa7daf4f39bb878d
zc30f053a4dfc90483cc03f95700cf445d6403848ee5bb39106ff952fc0fca22c1b8d0585bf2cc8
z1d034362126a276f5284a50de55c016aa40c0db883baa82e25cee27e0cb01762afac643a7e9602
zb3faf6e76f1299d0bdf3cba33beccaeaef9ee2e95a74643ff6f7f4a36cf383e3827cddccdbc007
z08371ba08b7ebd2ee97fe265590832bd3bd968a596e20a7365a777aeb6fd3a0e9ade35c38821a7
z2178b4bb70ff7855381cb35284a62b031dd89c8b48e83fd65fd7fff6ffe2ca83162f904fab68a4
z511de0a9358110709aeb159b9cd23cb005997491af32821e63ae72b0b9bf203c24a3d1e6ac7244
z5029aefd44edb6eb02f68c2395ba32342d4fc716dcf946b2e566c95651b819072041c0e41283c4
zaa803eb71fccbff6d7f1ea7f0e517cf45bf32541f3b410720903e69ad0e0afd47fb5a45184d01c
z10ca83995d16eda4020fc0963e85ab4f5aab0d05ef34f562c7a3c6c1280a712c0b76a0d77e2d50
z3dd387d0865bc864923998748b294b0432aa752b49fc76fe91fbf6b965c6e860c4fff66493a738
z79234d3528272b23c49ca45c3e3505706bf6195d441c808a73005b3d9bf071ed3b5290eca731fa
za614fd03d3f6e54d1a7c4d28e9c94cde173dc7a314fb2d9abd00d1cc5cf9960a38bd952d0c9e1a
zf5721142bbd3c90668f28be63587e3e2156e3f285ef6b70268c2d823593cc68ba1c7bd61394d1b
z52a1e70bdd7094c3ff1d2a5cb18d0af9b49455af87c2e9c867a7983ab28ab4a5ef44d2d4f1fecf
ze4d600dc5e43df25428867b7af66992b74dbbee8927786786c0ddad5ca7ac3a6b92e1891b8d349
zee86c2912bceb088ffbbca3a1777939b73a539c3039de9cc5c6db0a75b2dd06567fc9ab80cf7c0
z0e39745c518fb680cd947f4cbb1efb4750db2bc6c8fc7c690cc90816c12903ae14c12085d96b36
z74ea5fb22f9b27f90e10450ce62c6bb4fdc89d45ba90d90c51b042fa481e39a32a1cf7e3ef2f09
z55cb10f81db4e5402aa3492c51fba1149b714a8c55bec96917ca88d97833385134303064c291fa
z96096d040a91caef9e942a79c2b3ef487b5ad647a29a4535344dcbcff3e12d0455d4a999e9cf29
z364331635a2057289bcb0840ee157626b5e929dbe7532b0f5298fc2b21efaaf72cf8917ddc5a71
zc11ec66db2bd5ff0a1fb5a95ba1f420c69176facf02dfe253022968677393e4cdf6690ea58d708
z80540c122f2d9efb83455d39818da06dcd95333e26fddac4f97b852d4553777c619e33cf3f24db
zf6aed1f5762b9df546790a403cbcf2dd3d6b3334efb9eb8b317bf4d43dc7616993a38f9967518e
ze7ca58cb1be0f5266eea6c8b51d35733e65357f59539097fc4c6037c188643cb6288e319229bad
zc3b9d7bda79a635e89654f68e7006dd2dbf04dbdfee03f60df9c84111cd60642a5739ba1744f6a
z12879df1942fef68dd9a1ec1992966673002926aed80c2e78b91cce14bbb551f2073c73fe4fe71
z38f4380128339df7e58d160ff5e2434c475f2d66811477aa196f3eefd62bcdb842c31e948fbd75
zce80d225df49fc21cfa4eb2a3aee316e9116bfd0f85f59531ff363f8112e62950b11b143c5d35d
z40618209402c36021b01101b230bf95120f2ca960a626496b97db6a2e4e80005d116fba9ee5bfd
z8ee45360721b9464855bdd6be2221d00cf2c1e1f1aa1cffc1a41ebc064d67a20acf188d6a3ca79
z8383fb0909a5d2e929bd4d3b766504ec5de6ab84783849482493a7fa3336eee771515d26d90720
zb9279a91abae3865119e5219f486ec79cb8102bac80d3b2c5f1a8f68fc56f396d6878afd605876
z2c19c2df05920552cf44755e283d0c369a14254f6b8cb5633c876292efe0c438ddc31f0de6d131
z7593175482748239886381a28283e93bd4cb977ba04ab4d8b7d9fe7c22995003541b576c3a465d
z5313f43996cbeefd49be8f8903e45c8182cd247953fea6996f1144733bc0987d442747066f2959
z56396eca2bbe295595bda53096b848820a907b3b695c5390356ad3b0b3623998ec9a0b24e19c57
ze0ccacbcc481b0578c3a2ff661dbe3aec2330e275002a5fdc8831d917366f24b3116d5b8603437
z78e3f0a35320505aa358d6caf2c201d5b321dcd4129fdca4855bf110241ba7863e1374aec0ef32
zeb06608a0ef06446e565816674e5b0580bf9626b064d208f854bfcef9767bfe4ee966320075800
z800b16242909030f525aa5b0f0d2679fb4c552faf443ba839b297e667acf42ecebce3b1c80f79d
z65f09ee2668994650af4c7d751cc1871b159ba23c09797e11a1d527134758a210f9104ac8bb20a
z2291e34f640d6ce9e47aa330865f7f1e5f5cffaa28fc96963fd11655966f5752a39e0bd9911865
z76e4d3ecb3ecdde51cee2755f7f28a2188b76c61c286926ee62963c4fbbe0a4826a2b275af6bf7
z88e783d38f08ff5afbfc9475dfc4ed593276fb9151a063a3fef6e4df5d8e21380bb03b3e826cba
z63f239f3696e7aa364b24f283b3af3465b106908347caf27efbea651c8016348984597586b6654
zfe350816b3147787c1e3b6581b0d9395f2f4a62a185c6eba572d72ccb55f176af7ecc9e4a0a8e0
zb799f7665d9ea3873290d5f3dfa45ed638e71bfda39cc865a0f90cf474b67397bc62da81df1b3e
z5b33a6fd8f3c8419e7d43157aafd9ab82b2f435faeff5335a1206c2c5f1da483f4ec6e2c8ba3d2
zfbf60674f385b950d18f6b29c28c6fddc57362a402565b5f31c980d67b08319092e04310c6d619
zb91007a4ba1174c62a84295e7fe090c7707de63de28c25c19f8f7fba7fb1354cc6a7dafd29fa8b
zce20dd3f8ec14cb88ab6a3d86a30347de57444a4cd3e0302570633e1222c2e39c70d010c38d92a
z08b734f992c45b62c5b6ea2cc670f642d7b14ecaa9fc666af7af42186cc5bff73c7d3bdc00a068
zfe6d1ee17ba813f8cd4ba5e8daf25844a4c45fc63e0e2b9fe1fdafe2af674978be54b065a69956
z0ce6dbd3b880eab2ad490c4720fff107caf10f2da027300a4ec86d1bce71427baf5faf079ca034
zfde80f2e2cb4343d15036ce654bf668b7a50e598105ab00ee6b0228d7b01575303689a81643fa1
ze87229e7588257327645e82eec48676ab55c328865a138fba5e905aeda32b66563cf8c5c7da8f4
z84f3a15d29d69d5ac05a207de4c88e10bc26ca28fcbfce81b9e375742dc3d805bb4d25f9b607fb
z2c3776317597d21efa6f5c48d8c2256ccda39cf199d4b016c246d92c92619736a32cb582d88682
z4bb869bbc7d31733a7374a43b3ba871d720db8f8ce2be866e6add9173c14df059933a089d645be
z51ab3a274dc2811bac5a1aaff7b0274d43493ce92ec3f8afcb695691ef95f393d9f677dabd2c93
z13a0bdbdf50f4269f3b6d36b3e605ba608a9d20c74cc9a2eaf2feb1037a0abb70d52d8a3f1b091
zb72ce11a97fcd079cc153dc90c43bd21a6f56583f4b74ed2f4ac114fa0a785a5aa9ecc95b9401d
z07bc5b956abb8662df1e801f2ddb9bf42353e59800d90f6388ffbf29a697967d9d5ad1b120b64b
z057f82f4f708ba97ceb8bd0e72b85b177506db3debedb2a41caafb990a7b2a3feee860e847b216
ze46e98b3e19e0d76c21321f7841dd6c67544b1a070336fb88e4f5da66bb7652024a5d00305e561
za3a9b20e3a19449b9afcd2ecc59c4fedb103aaea46fd069f6ed079f5dbbb272df27bac514a7d23
z077a4e430880b96584025942639f9aa4d3de7d1a1036c81965f2d31f45603686e7d034efd3f0a3
z8aa207fbee0b9fcdad6a48e3be39a2ed1d691d178c3b6e455215833a8fa68d076639ff7e78fef7
zf7a868b6078b0cfe75117f8517f58763a149d24e36caa26f3ce1876ec65cb7e92719c0db3f963a
z9d13bee538e01459e8e2e612cac39d22f162f14d47b9d92399e2a1d5abf2123f8c297fd9f1e534
zcd8a69bd7d538a445e5815a33450f5883cc2c075703157f39bba218e3267196bda32ebaef22716
z55bceb6a87d9a1864755d4fea3f2e414c3b67936d6ba49a7ade9cfb77fa4acafdb82d60ef514dd
z53602e7af1251dac5a1ca98dd4ab91b5b793178ffc4c6b3f974292f8b33a9b1d792b1773f49d27
zef8ed014a3c8b1bac3a9585fdbe4e632bf71271b32f9b5b95f8c16c5b5fa26875cf8e7586a330c
ze840fe05338d3031ffb718ef7c8e015ccf9174153e25c21546be73e13809cc9949a39c67e49d6e
z72edc37c1d122a8d1f409e23c36c5e6c2a82e1654f26d2035be770ee5c79e943dafc32d04f014a
zbc86bf52a235f3aefff4557108e8fc152e3bac2db89dd4d80d6172369906ba007fb60920fe74c1
zb273010423f1222fd3911e5e2b90a0ed5418d7addc325a49d54aca349fa29aeec161cccc4f930c
z640bbc65ad29a8717d285972466c23dabc89f3a20dba36300ba814cc795c67360dde913b8abd40
zb014a5f44db6197519330402d559cd775b327f1ab37a85f628bcb729275a254920891b639297c5
z6e61e228e0c50451fe58eed92fc2ade8801499b442062957e7e7d3f711622cff7cbddaa5e6ecff
z7dddc62f434bc3c9db3e6b6bd006ffe169755252bad6aed8d77c67794c8a0c968c1bcc627b8f40
z31ca6a3e10088cc0d3d3931148f5fcd0bd273184d71308c6f6a37b04e4cb73f186b333929e5124
z20c4d35d35f0aedead159b5df09e2e959270324252252a7be8b089f5f705b82eba96f11bc838b7
z5b91e08fefb4174beb12041d44d3c47208765dbb912dbd61363b95eec8f4cd11c997cac42233cb
z1c908228a1e7df3b9e8ccf8f69a55d6ea9956a2aab6c965bcce353bbdea00f97b4eb8fb30ea16a
z2101d0cc53b1ad7fab1a5802e65a9e5c57ae88cce8505cbc8202521716caa1ae81306ab1807c2a
zef486d7b482f00726bdcf891ea9f7e6eda00296760cf052db5e8832984f12b4930dba26b722015
z84328d803bbb514fcfda8fddb7306677b75f7de7e1867f088693c0aacb463bb106796ad3873db8
zde4e4bfc46c92962dc12a64a8add03468394343cb0179067c405c73a3f897ff114a2c0d296c426
z1b43258165cabd8193f313ab4ab3fb9f684f245267b0f641d984d095a7db57275f051b7fc3bf52
z4f9858844f7d0afc9e27bdeb0ca5ac8871330874b0d17f637e5511676f401955dd9343c2d76e3d
z75165d66ec512c9e97d30beec16b60dea56924fe1659d6dc24095e5478e3ebb904824f3ec71680
z3ef3da5285c0d5dc5c72c7ad902822029693e8c24aedd6588e4dd9b096bb035b3fad01c29a9a07
zf317e6fdf1852705fdd89f02f7d255e1061956ab2485c35ed38a4c6661fe6826fb5f2acc84f7a6
zf8c00c93c7d45a31dcfe811fceca7e96a22977f3c5e24c3fdc9ec7268eeb02d3729ed6713f72a8
zf0f0e898499ebbbfdfe2bb1534ee0a0ab6fc9fa94c3518f5bf3c7079fdf36543343fcd90e13460
ze722dbad3d4977f59190dcac8d1bb68bfc599537f989a4cbcd0c8b14ebcddb04934de54c83224f
zc7394de3eeb6f729f1348fbf709ae5816465b1417e279833538f412a0cef348e0177704981b895
zb45ea966766beef21c0c13e5759db23ab2950d8295837b6be427da36f28e3d0c50a101e036c41d
z5d8041b8d6a36e0f6154893d5e89a75ade92ae6a73ccc19a9cfe3cf33d1dc3da12427cf17c27ea
z00aee9826325f9c36078c9e486b12bd2027009a071466c6d7b8585ba28e682e3cb0040c459e929
zc9305e180dfcff45ce4e6ea833f889b1e6f04e96702468d8eea58bda9be730c1dbc4701bed17a3
za506455b03748db59f3af817f839a818efb18e7acaa7cd53b363d2c2eb63a034631227817b1261
z103629fb0f63fd5ddf9087ea731038582394244d050053f233624dbf9279c04f5bd065a1392ee4
zdcef8dd30843e316a5faed89b53cc0ed823bf3ae7bf6fffae55764651d48414ba09f1f2e811362
z1b434f2bd8ecad0caf4460365c77da2dbadb687e211fa91f461078e66ba31c55dd29d3924d7a69
z4bb6f4d432876233f4d43962b9c5ad4661fba456622a706a558d5916167b773d35efb08d97f70a
zee4d9425abbd6ab3657a8054f670c7de36a756d53d9f175233256eda5e359ab774222556e7f99c
z727bb75c61392d9140dbe224a36006fd6ae3af367d39e7a6028b9d02032db4d9a5382b04aad51e
za8ccec003081ee7de2175a6c498b1c67370b98211a214319873c7846a22a055dfc9b7fb4260312
z700daf6f21e2e5048a05406bad8a4dc6194e456a835baf0c2c6b3b424803629226f657ace53b3a
zb38ab4598b736d0e64160688f53d3cabbb8dcdbaa8cd1d5f802abe06ee426d3caa14a03108207f
za40ee9506f45c28fe0ec4e5c1af6f4b98896686bf853a8ed1c771509491d97821a23a1fd6105ea
z4762775bc420570743e7532d4934830a7476786d0547867fa16909323e071e15dbdcb11d11dd37
z4a7412ecbbd62dfa5f191dfcb0eaa957a3cebd343ffce367a3910678618ad57a102b5e574023b9
z53f4d7ca614a71e8f88a0c8449ce6254e6856ac013b1c51d9b62792e69691d24e65539f039e91d
z4313555eb3fa4259e0624cbf1a3f27dac4b1a5e03a40ba3dfd030b24e6030f00a9b4dbe8d51b14
z68de3a5a7fc4bd39d70b8600ef80212fb4e5c46bc66fbdbd2116aec7fed14577e4e0eed45dec73
ze307f9a255f93375f904488813b8ae4a0792473f658cc94a6f889507c04a00662ef74b236c922e
z6c2dc6a9ffe9ef45f8e4f1e7360448e6334cd326ae4fcb03197d570e6ac1c28b12c9eba502ccb1
zce4265f227cb52990f76a4c8791000d7365ba445533047dc00c463bca2b929f6ac2d57d3c1b1c4
z0ccd970ffcf287212d3906f6dd874f91839c47d318e654a1f29a59fc4981a302880012793f3934
z2ce85931c90f5c778614e7b6d63a79863da61baeb22bff6fab86225a201e58060cb9ff015f152d
zaf310cfef78c7f2d97613b2a34341634e7f4827f8705e989d2ed71cc20f0decbe22c3f02922df6
zf5f1e9620d70704d6eafc47667e7ed40b5ac87b34844916a36fbf6467c85be7e77953b33990afa
za98b66a930e75dfe27554ce594966efd4800532f30bb7f2b5c39e92503c6eebff71b823a580644
z59baec1dcc3cd36a87e31e7d16fe6b888dec6137718a69e0b6434b9d528f4e9d3608916f8845a3
zec972ea7c4ebb113d9c72c9686bbdb9a7a864b60c009711dee8b5478d703c201007576b9b5696e
z7bacd8fddc7898a058c58fec287253ca5a465e6ed24984640a3190ced526f5c28e11f73b0f4bce
zb4465c849c9ed7313fefadfefaaf581eb898938ea3958dc8664ba7d56441af8bda4a128937ee32
z8dbcaf936fec01991ada4b23fbb0d7fd68f9d8198b65fac0462bd90733223fe2a841d0491441f3
z2160615ff6506e4ddbca4f82ce023efcf30ba1a0ed704878627ef31224b9903688091579bfa7e0
zd961ab9813b01ab774010eab0e96a656c00079248253b9d62490f97125ef39c180615067a4aecc
z0ffc85e3e707932625522c6b2ee55df1a77d3114267aabeb8634c713b48ed06aec0102ec9ee93b
z80259cd13683cb043b9cdc8e8920150ea22aa4f88b0286db7aee8e9c642f293cf50757daf3ee0d
zdf847f753a755f015f549d30e19b47406a120205b720bb16f54bfef01fd716bd61e4fac8694286
zaaf24ac7780fc6951171ebf638d8647b37baab01914a49453d46296fca920c81bcf2e5fee5b75c
z3bac58ac973fca02209ec1f1f048575ad4222c5aefe85ef0472b8788a5275a64e46e56e5cef115
z9a0502bdba936db94c097a9bcb09ba9a0da3a4db6d4eae6458345a00987e3756ab0568356a2147
z0ce729ac5d170daa48595c47360a81bc9a7ccc1f31c6e7198cbb6b4c9b261a4da407666bca6e77
zff337bba6d909fef3b8b0baa171ffe41b77b54ea10d684e937968ce2cc94dfa02744fdeb2dee69
z8075335e2e8541d655af2f78d71fc14fba3715a21633f88202600cb69ff1e8f146a989b2c9376b
z93a4eb359bbad5b72a9e974f3940ee712290f3aafa8575cbc716cf7853134358295a765e2638c0
z809bcd3ebddff4d8cc6faaac835eeb66b9ba8154aff88164b00135a570bacd60fd70ad28cbab2f
z8933eaa2353cf44dac310b275b61c0972d36306c520e28df1174e5ee1309782a7cfde9fffcd720
zf24845178457c7f0e8cd161a9cba83868b6022dff667de3a4367d37b7b20f61e0e5dd7e5c860e4
z5c1555ad27121d307066287f61f0277fa43995f74a0229f969507d2b7aa5e6275e66c01b46c894
z5636b93d88a551fb8a17d1de2aeee22ef5312de8de471dce925ac9366fc5278e6358b9717c1995
zdb01da320fae5c5685a45619cd15c5e353d98e9968c15266c0e5bcde3fa33945e2cebe0e266fcd
zb2fd070093132261e3d55b919fa610646c1a38fc568d60e2413c10740a7dc7d4e670acc46b9420
zc259ea59b99145bc906971cd549ff0fe3d803c21c7aab45da2eb410cc18f0aef8e20d0466fff08
zc84bf297b525626a43066a9e47afd9997f2ee6fcc2d0a29055ae49f9e4e42e05494b806f901cb6
z16108a4325437e022cdb1d4c252ced964998b204e76bb9ef69f1fad9fa950e8612579f26cc4e06
z36e7ad176c5008c5754c5b08d41f75ffddc12a2f3e3a35ad9842fa46e47bf2c88a500edc7f1bf7
ze2cba8ed3368f96650991d6dff7e2a391fabb8f7769ecc1db671bc505568f638295c55c77348b1
z5ec87fec77967e83ba22d7b70585b54fc4ced9caf8298e256141d7db82acb3ffa299881da95fb4
zd2bf377c7cad419eb0ad87888868406730d4789f8500cc57f1b5e3b7c11fb226d534e99fce9aeb
zace1b96ce413ed87e5e8d69bf9f6858bcb94c92a97246084e1c48a98ae6a31f5bdc329682900c2
z80bba958397bd3886e28cf5b34198befae3da25d1285c781e2c9fed1f11c9c83d33d54502de00b
z47e04a34d3392fbab823119cead433bc7a5920fc601e8202945a0e77c800c32ff132a2eb1ef482
z84f7c0dd1cd926b1c0d9d78acb4ffb32b574148ca21086bb4e11d24e3e042e71ae0f710ced6310
z08ebb70b849145a4952b6d99d0707c9cd93242ef6f53fc87f97577d7749c8a8c929e27a0af5bba
z3af38204bdda8f26d1faf0c33c683b51da5c9e455271744e215ffc938a9efdd62667ee53124e0a
z6608f0e9aa9bdb67655808526dd1186d1ada19d6f0fac7f2439c7005dc9da60533b491cbc70e44
z4be03b806a2f7a28d0f54fbd7724ca6f784e1dac812a705aed95042856b4e284bdb60e29b798af
z470fe63a4ca9b948f8f946f6a26702e0de28821356719ebda6c77d3578473c08555992fbb468c6
za1137a16457ac12d26a601aa6847e488f62b1ace10e9dbd15ab00150ea1d9aabfadadd73d045a3
z155c96b052781986f719581500638e7e16edb783fd00629457d918e0e37fe9ee7f88a582e1f40f
zd4d766d347fcb6802cb8b49a6013036db7cb3d42b562e60b0c39f066fa8b654f9ca7422829e28f
z3cae7daff3b9cce57a0ae18ec85947f516e66c80cbb65462f2dd3d5d93c668bd3c19a60ff2a3c5
zb9cf842d4bb9deec5c576670ecdeac2426bdc5ad7eb41bec8d6e2d9bd3e5752b67a0a3f8adcdf9
z065f238184e0781d86243f632f2ea9396e0c2ac3116f4dc2deb5095d2249af830738112a7ee1e6
zb48bc95c9b879644ade3ae67fad9b7af8bc9f8b29c71b8a55bad7ee72aa4666b85198cc2180ecf
zbfd1ceeb6fbb7499012f7225abc5e4eff71df8a5295c4438279359a1b9cf8466de8bd352361fed
z26b00cd5aae032bdd19f7fcdbd3dd3a80c67027bf5eb5c5ba46e469d5a24a2b79c7031d0cfeb57
z6c39d91222b7b2984ddac02e949ce07466d10d0dcaf6e42bb107b913bfc9a71bf2d4c5dd10f640
z6e9f4c41590e8d1ad700d364e4f101f1d5b17564e34d78c6a1fc23a8298b1320523246a0dfeb7a
zf38a8184527e3f2d1bee991a3d71066e47cfd6c6cc467f0df4746b7a930d3c3a1c95b9c05f0e3f
z42f6f7a834b43911a0e78c1bd4f9678b00fc2707adc79019c703a6a7b09744a5c70b3370d84c67
za3232f8250bddeae94970e4463af1e2a860c5818d26bafffb32a7325456e6c974b5beeab60cd75
z4c8e7b7980931e9212242d84cafe682f199eb2ee9eaafb748d5409cf4229690e6be7c71a9cc462
z9824ddc32307c4fd4a1dcf07620f61621a8677a2e3143e325e6cf04375f4d978d79d8fdc058e96
z48e400c34a93bb40b35d4469496c914968349b83fde67d894a0906e5854853db0366d33f627f54
z054d244ea72ab1339aafd65ccd825c9341373f28114a784239facf16b2bc0fdaf34e0a8402f78b
z4a1400d216c4d146fbaf3056788ce17ce22f2c34520aafbce57f81f05fb9e9e88815f6d1c6d63d
z98fd532f55efd8b5ead52ac5a7f44172a2b3af9b954e58274113c03dfb530474b3f0953f397b94
z197f4d458f1017217bbe2b878efc736bb9a2a1d5a3ec24c9b56692eccde73c527bf3fdbeef6457
z46bc4c5b3cc5a36749996bb9e077e4a5c24f0cd88bf8abefaf2ec9bcb64c5eee37d8dc003bf710
z57c9cae408c2f4e9a3b1de27e0235c8fa718bbc990bb4296f3115625b403a45b8c97c1c7cdeac4
z340f72e7103eec1a77603bef2b63a21bc2277b2d2211d958ab2d1934d6aa8915766b4463385d37
z9e97b5af495e1182d51c9ca6b210a62adccbb47e856b4c7e2a926408d84a1c9e1dd0b854091de7
z82c320ec4379af8297bc4624038c1f4bb1af1c6b2b9d8b56398f254780f596d9a588676f8c7eb2
zd82b07191b7b59ef8c26b13d243d4e8d77c04dd539f9f46b2d9ce0692c3a060329612cc5330586
zed06e3f79a91184154f499e8267db1c8a89fa9e0af2effb25f7b8e26dbedfe89c21a97bb1ffc6d
z186ab45033141b0cc92e8b37a6de188b7b2b1b272317e862920cfbc2d93a81b482e4e70241ceca
z81a7333488753fbf5d5c6d510f0f74dae8744ac9ce86edd43bab6b2b48333d8def3a3d4c7fda06
z1f975bc7850fba575382b45e4bd91d69dab50f556b822e5524bcfe1de9bd81a618303e82bfcb32
z882f58f00345a68c5a9d26442cf392bc6c1082be75e3fe2c43ed61b66fca1f6a2d26124964dcf6
z409976902c341328a8147fd722e0d02aca811529d830c09ea823675edec7d42e7833682c7be72a
za06694b926ff328f662df9c932484e86e5b048fe801aa28c303ead45a6b35f2a58ebbd526d31a5
z63e3d0e1e10fdf3871e5f9879ab6ea516b61b9d86b3f00434fa12584c62b2abe5019a0a3d7369a
z7e7296226ed253a64b8f518c64107ec7175ee33e460b6d9bc3da8297cc43fc4d54b1a928e28b33
z5c8f7a8b8f6cb63d26eb97888fd04b0df1fae1aea99e7b8fa62418e69791a25c50b0fa1f55cc0f
ze8faca9707a8c21b4301212323009b2913df1ef31eb36ad5eceb4d5b2af9936be6001e305695b7
z301130a9c64008a8dd38cc0828f6191ebbcdb85e6263dd71f7247d51b74e29d8f75490b8a75177
z69c559c38692af7450d33831c07c1a83dde1db36f4b635e2ab18a92d695c50e1bc0fa93cbd8e51
z3f54ea54226c79983dabd4dbacc54e5517ebc5f677c336b2ff0bb5734c83e9443cb714b38b9e9c
zd7f6c463ee5e880c7cec7671fbb585d0b7754d654d2654fe5f399cfac9906407a480db5cc30fa6
zadbc07401d2f0e33c74e45f0c4355c3101b7896bc0360e24128fe982c0b7ba2dc2ceb01bc097ed
ze1654cd2fc4823c8007d613d4c9f3ee39326c5ebd1993b404ba837dc598052a21bbd3ff1548f26
z02853435e90fe96c2914fc0166e27348a7d2d13a14e55a59e8dde7595d234cef098481b5e02b22
zc37db640731b556a35fd67571708734afb3c4d84ebeeee8ca8a4beb95aa6d357bf0fc7c0b8909d
z5f65a9358287bb4499fb095f2acd4c8578b55edb14634e5e4f0564c848f04939e9214a818651fe
z8db0d8ab4fa64733b3e271e75ca1cad911809a0bc0b6f5d11bf3f2b57e650f90fa8bfaec0907c9
z272f31e78eb131fc80fba71da5337b3f54780555c510f4db8531b7e5e507abbefece222b482d7e
z4f3d613d1cb76965a228126d1eccc267148877d5dc468bb308f2d98128a4a6f47b4ff61847bb4f
zfecc976c74b4ac67bff566a8dab646bc5bfd7e22698a2498b325703d505b87485bd4436a483618
zee3695074997c5c6159375e6161239633188b8154023621d807ad412258b575b4ba662a5d3b67c
z625d5b25b1cc5594333e2f7b6574505fd6ca4779715b4763eaeee0a9ccdd93707a8d9496c44be2
z95517ffa9bd35e247d64fe6875913be89a07ff234e866165e25900b0d5b2a10d133883bdda2f92
ze5913fa7f087c5da77b0e2708f6aada7c4b09a48c3db2da5db31061ac3183374e0adfc605eca27
zc76e322d085784e18b27ac187746fd3ec44b0e5fede26f8bc56bd05035b269c0e3f3d22ebdd43b
ze7f5bb99dfdc67bacff01fb8138b097f6adb66e49af5970dbd3f7617e3c7e7065ee32fab79cfd1
zf969bef74d6a6935f1477e78a3149064c4c278d7b21750c25e6eaa9b0036e57fb934217eb980d4
z0ddf0f9aff92a52c83c3e0800ad76e6105119f2d7a5f5d96a4ce5429c44487e29873367987fb6f
z7392b4e51aeb42683819431aef05a6a1034be53cca16686cfe73e3fcbe28fc29d92a9d1b8bfe9d
za77ce03ae120400ef277ba1358d3272160c7cc2a54aeee4910bf980597b956f2549abfe2533c07
z1c0798653391c87548317339c4c1486ab75e9b686aa49e9f9adfc5c80bee0ca8c4cb9b87c0a8c4
z346368f41c5ade47f561152bb69279dc937ff59c57a1e1830c6862abc0eff97635aa4dfd8723d6
z03ffbb14829b4935fa524faa80a0405e51e7937fdb4619ad012ff2a0326b7ff475037880d7e0d1
z60eba1012262776e5a23da0a8c375ca9fe4b06a6e6fe54640a513b649fdfeb208e6684f67958e2
z8dd613c82d7793c702dc53db060fe01b569a4deff5a89d8719635a602a07958eee7372c6c2eec8
zdf07a9c609947cd8b3bf391a308ea80575719a08d5063ac46f48b8951da25b60f8fcd497f925df
z1f3aee7f197a9bae0280912a500d46ef4627e8ebef4e0879b206f00e28e63c65d2a9177175e0ee
z4a708b1b61838b007158628f79692bf8aac2cc7b0a8e616540454c8763c1ee4c6cd32c66861aa2
ze0af221d767e27e250837c9134c635cfeefc85d2aee6cd043f1d7e0222dcc80819cb059379b2b1
zec55df7b1592bb94f9b7c8480ab80ed808aa481268b48e238bfa176110d1c0bb623954af88ddf4
zcb9553da3f5fb612ab85b7fd90d87103b28348a62a04bdb051318b8d3e6ab3ef2f0710f4b6a2ff
z5f06ffc4b1da0120193117eb729d5b92f4a9e2aae05f34f749488cce9d3abe536b46edf9a2a2ed
z1ec0e6f6650050b052b76927aa363fa09613907f18df47651cd8e790207d5314bef8b50554cacb
z86c4863d1b7f5371cc523105e10a74ef601b5ad38331d81582757519bab05771f52f7ae6933c4b
z3df4f990f07ddeeab08f470218e7d2591546f1f6a780f83b8f6789f8d1373b2c795b872c0f64c3
zd08d46d52a3f7f756aa5f19c8209018bbd07d926f4d3d08df74459c614c25d53b73a2027bcbc94
z68b0c5c8a37d298f4081d79f038b270d4de43ae081ba0179d4dfb4e422c62b3958203e667e8b4d
zb3e416a8a7d9f08a2f4f316d5b5013c09c49bb91046a809d200d21dd84ca45050bd14569e68de4
zeb44eb5f94ee3ee8527bf980675821e0ae6765ac723f1ae84d0bf2d73beef383505b9d0f6f081d
z27b631827706dc57f29f4e63b8a08eb8da2198d5ee9543caacbffa405d5273b9d441399f4a4388
z1c5b7f4d255765e0747468e4a405295a35ab9b4eec1779cbebc27e10c1f09631d8b5ad2cc347
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_stack_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
