module tb_multiplier;
// TODO: Implement multiplier testbench
endmodule