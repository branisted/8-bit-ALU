`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab30857016fc53a
za25afc8341302f0c829d94450c399b8ff9b0386c187cb854ee330605b7b59da379b1f26f488e1d
z36e675f0b1336408b3a1ad87d0723054f952fbefc8d5a33eaca6ef5be8f42bc59870a29a5cc9dd
z4fec09ce6e44cac279651402e7e1f590df88ce49ec26ab39f12b4a02855703c6f03b1e85c797d7
za357087d98e5b1f45502e45892e5823d6fa4b762932009620038c05d74efcea7c3fdb38901d620
z36515d0824367e48d1bc182335f158c262d396cada6b0ad58add4f945eee634c2dceadbfb5118e
z14969c29a743830a07124bfa78707f3952b96b0db7af7c9ff36f77137d8c490c4f79328328069e
zd7d5280e4f95742c9841340368b9764f0f80413adb175ecfbdf3c40716abca7b8cef6f7fe92ab9
z6bd2453f1aef7f7899c5365c5c83793cacc7795c269413f6cf0dabad14d40e9285afde8c01a47e
zb61893788ec5060288cabde8fb553f21b02eac61ab0b48ad3d54f4d1d76508b22f0c600861b5ce
zcb30ba708be817b1f50f59c0f6fce449203e73557b1ea4d25ee7597945d9cd5c651b4c2bebda9d
z1d3ccc0b324e139bf8ed0340e187dcee0635d170ae70865631bfd9f2e75fe56e4f78dc29771a71
zca75fb2316147d8f4edac39d595f05f42846c760552e35e976ebdfffb807b9e6fd3a3147b5ea76
z081208cfad8b034c5d384f986d488f617c81192535f4466e61c6753bb8eec0fa5f0307537cc337
z9ac03ad109b8115d1fe24ad740ea2cffb441aa5d6ee402b7a2c4fdc1bdb58d2f6744fce6d55e4e
zfac8f8f066c528d318565a219ae8a28e1f46ad3031f765eed3acbb1fbb4f291305ca0c62be6d45
z950e6e05fb331e796aeaf0ea01cdfc30561e050031296eccb3e5bdaf528172a8b854cfa3e86a48
zae26bbca163b1c26a3bbb86b1c9c59ee9e12d1c5012c398fc0ad9ade11c540f3c3a204ad2dd971
z004a340cf652a510531213b0f728b357c552983ed534805740567502ec97068f1551c0640c32ca
zf0b8f27ee616c093154c1cb4d9270cefdc93c179f5ec7be0e6fc33944e89f0fa70bc6f2774ed15
z57c69a680a05b7571fe2cceaf9e27b6b304b03a80438fa12242e5058056daba1cd6e85a4638153
zaeac855e7f64ca8fc043ef32b6c486ca03302dcf0822d6aaaf8825f00198906298c426046933de
z7ebafaf789dea6a508b34011d378b8c80f14e37b367deb0356388c13ecc0f441cfaeeb382b444f
z6d28d537015ecf41d174481e3f05c5ca908ae9820e5b35ad3506c605ebd7dd087d45cedb6e90c3
z271d9838be7a7d6b226086d6baad42d6bd19a2e94b46ba09a85d74181d481c247dc485a41631f6
zb84a73118b6e5edce329bd7b6494939265a0b4026e307e39201dc61b362359e5c164907544cea0
zc2fe1267a5d015190088d499bd43ab9b5b9c8966562ba773ad21a42ac18076156a100ba6ae33e0
zf76c7dd35dae3000719811d44ec3cf977f2f38d71c8b23095bbe5f462c24e7b3ffe552180427f3
zd9fdfca75a0a5c04bb243a1560cac73756e301c24595240692dd6d44cfca850d709586eb3c4aaa
zc526144a8c93a848ea593cf5683795a83acc12e586b2ade1017521f2d21c6434c31a8367b97d46
z71e7a79072143024bbe3eb8531d7d3a199c73885df1dc19208a66d2592f5c2e8143354ab2e5bef
z430a4e02b1fefc12c19431d8a0a46b179653ada230758645258a69c3ec79aac5f651f1b6595441
z7fd3de0504e8b59084e4dc204c37bc047a87b67010be776cad1f9bd2ccec63ec01be3e5f00761d
z084da289cfa1c39a572b4c1b4cd89b91f707ec571ead74d42098b504b013de548efd71ae1272aa
z96290e6a1a7255bf646d87cd7fc2a20c1b2e02e1e2826a73b0095a1a8fed85d5a78105e4df9e31
z3943b5c76144610ba72b9de9a0f60dea3da7854fe5abb8a94717276fde8c3aa36d12e8a3b7cd86
z77b22e7aca67684573ae6df3347bb2ec92eed2d6b9d3d4b1b6d3c3f05dd90bf7ebb4fdc6a02354
z664ed8e5f50faa2ed89150c33079babc07d4acb01e1622ce9d89a626b3854bf5f26440fe531821
z860161a6de467bc07261c1f0c5ab843844a7cf080b28ec7ad838046fb5c0ffff6cc603bb87999e
z3533acbf6f6a208a1d1a973d027fa911c73d87c8772474158c0f37e35c40bf7db1db3558f608ed
z2fe39af2f156ddbbe3596584e0d47140801a9950405077927c814488653927bfd46c476b4bae70
ze49a08f93511b7fb79c5f906308260b19c8ed8a59016bd8e5c61585145cf24ebec77090cfc2ef5
zc27c4dc1e02fbde328cfd20628ab04913a125716fe06de3c7f1b864d64809d1c6d516b6c28f251
z4555bb9f634bf29777c702e6357beb650365fd834d8d7d82cd2a2449c5cf5c117b83045f7c1617
z740f786d33aa84bcd38ecb7d3ac90565b0a98d1117598b6043cfd223b6b6c7d3e5e7606c376099
ze27b6f26ea45dddd9de6011f3055c97dbb71377702ca005557aea22ee7f03e6b33d8c7c3255c6f
z848b407876aa1048daed5beb2beeb7840e4f500226ac071846d5b7fdb8959f7cb5ddb6441ed347
z63dc3cdd79ac5d82b92f955fd04e5c75d692cf4b31a74a8bb4b4fa1468fbdd1b66f29ff715ad96
z2d6bc53f517cb88903973f6b02f06d3d1571a5f95594c89504ba3105647b368a6c419d4daa77cb
z6ddf1a568fb691525525484b0e84e65acdfd62b4fc7389cf7433af2f1206edad252bde23aba81f
ze4fb37b7425e0d5add4a1971acb8d7aba88f643eb02ca90b9f112a5e9a0e0b26d05d0e75d8ac27
zb5a231e381dc81f3bc1d558c7580b82b80c3c7d892d52f3cc13d7b009b3fa8f04852641d710511
zabee36e9d64244193ec8355291f054aac23cebea4ffdc49edaa7fa7012e32a14acec3b3e4911d9
z80d139d9ef302afb5bec00500daeb90b7710cb73c81f34b5dc98ed9113db61aa8d71e6f1d7920c
z1019cc3dd2c8fc17de377c6fcf42a063b1fe993c6e14177d146e4e306eb35cb45ba053e59230f7
z0e9f9a61ff857573e613298dac4d643cb56043f51b105a6b71d2cc351e838c941783f9727d6062
z9a95bd24e1cdce339ad74a8f9b7b312ceaf792e449fe39e4c01789b79c270748c6249f942b9e58
z88142dccfa3003ece5737d8d0072cf0c17d3a13cacfe2098e6e499310c40ab47dba29e6b106631
zc15cdbf01b15284e98ad6608a838b5a0475081c226a3b2575a24ae71b3f764cc4a355f4a4455f3
zab5d21d921da2a3714131234c869d301a3b144a88db320045053187a1e162df74ff5bafc1f458b
zdb1d467c7ab2c17edb56060a3da53197ffd607f58a127c8a5ec3192a30ebe2fcff15f00bf7c7ae
zceb066c85ac6d51a1e938b27cab81b042cde35fa8bb0a6496725cff8a7fe39e8cc275ba927f7d3
z5b28044f0b9417b5e24b456e51a568a59cbcaa958ac3f7424ece6da32425b922316ba19368d329
z52f9b9185ea58c216bc0982359915ed7c46279721aadc28a57aa24fa7a4bf35656713debf666bb
ze8d74ddaa50941706b6284206f63a30e1350d06d7886a0c32a52fe97fffaeb2275994cb4026ece
z39e9416901b75041aa0760f914e70de0a939ca79fdbb8fb2cd0cf30ba2b25663bdaf135e4e9b41
zd066f7a336d741737e362dfcad36c31e544432a060aa08488e31ba3a54b479cec905b33cc16fef
za1de01c05911a14feb9da10410cc73a4aaf76d63e3d120d921200254af808d5707a0a5c90c4188
z1c31e1d25252b3c7b26ac4f557c0079ec8ba0ac4072563fd60063dfee9e32f0121305660bba4ab
z0d18efaa67cf9f0363e5c4cb39b3b38d3376cd6f3e28de9f5206266e5430ef5d73d099bd32ed76
zbbed1305d62b0927240c65b557203f2295ec67e699671a0971f2823acd1555c1549df48ebe274b
z38e880b386ed2a1725507f3a5cde1c132def69114c4c4740bf437a9bd0e218c139c0f744e94d97
zd5cbbb427bab2b354a37f284f012fc878ae7e64a6e0f7482b7f41cb4979b6a694beff5d1fb926d
zd07387c3faa959dd5b11e875748b4fce4e45cf55da00c72ba0e2cdc17b469b2aecc2d981b02c67
z3fbf14deb2f38c96143bde0a9c96607534aaee1a51071502dec83b5f50dcac74c4b384a9ab57f9
zf58e356eb481c7584736772564ab8eebccd237ce36a3a37eaa1a906d076effc32bc36e6d893166
z6857563e816305ff731071cd3b0117ebdc6e75c37e97b152708c735c9b8d8a910148b0be7728d4
zbbe138c62bafdec873f7b3fada8eedd1bf6587756e5df1dd624ced0da3cc5d583efff991976e45
zf20e586dadd600865c6d1df4e7c85b5d080c38a1720cdfa8d0ca3636bdafd56a035e06b4058f6a
z1c7587c6dc6c550cc9073caaf67121ea4860c6e9df104b6a113325f0ae6413d60925bf89c13c6e
z6c43a6cb1ca7e285f384e7d12d939b1ac3577f8b242b38ddcfade2ff4643c1a4cadd4be4050cb0
z82854190541c79c05ddd69f3e4c1910f92362d843d24c1a2aba4f60822d9876ae1cdf05e0baaed
za73e6b257ee0042c552d7721d05f27b5e571dffe4a56c70eea487a144f0951d96ca12f003447ba
zd556993514d35241d0d8a1fd39ff63d8ba91d806f77454a435feb4182a9736c092daaa44e258cb
z88586e700e86b1b76c9128c76ca36579699a6e58d694d38d63aaf89ca5b130b08ba13bd4e4622f
zcd176b406881c3025aa1464ad6bd4f8c20a9c5d94f6722f4ee4e59a3fa199f824db7e1791f07ba
z57b8ae85bfbbcb18eed533df012369c7b19644aa9edd23829e87ebdf6807209a94202d1f0a0021
zd4fd441cd35c6a7bb6080d0c3d8d17f90d120ba5bd615a2ae9fdfa35968941c8d2834cf25d8bdc
ze1bdafede9f8a1fa0249ec9ad5ce00d0a2403083aac57082edc15c1e8dee9e075e8dd014898cad
zc5bfac27e1de69556e23959497d026bfca02447217d26be2414beaecdf7c26b3b6b13b9278d2d0
z77101c8463041f5915c1ede23b75fbbe1e6d6e828b292b3318aab1e9dd086bd7724bf522e6e36e
z5af557fa0b62603cfe5b630f16dae6037200f91767d001f9e7a02c78529005b11386ac97ad2c2a
z053cb2d7adfbee84a160de28619a67309cf04a4ed98916c7331b8da2ce2da59ba08f15da634e2e
z96930db8efa1a39ec73a70444ed53c1da34d170e8d36d2d74bc62bd05b084eaf9b3d0b042cb5cd
zd077370e864c2ff5f70ec426b53a508031858ded9f75595df757570f4d224af0d60a6a4c364867
z4fd2e805aa847f3dceaa9711855f72a9b16e65ea7a28dc0f262402a932e89db9e3116abc2fc432
z164a21b2b2c0dbf5b49c0c6987c451a417ce5e15ff7f195f6624ff434104a1d8aef4e39cc2c915
z5b0b003f726ea0c57b08aa79dc5cebb85be4923e069d15e037294114eec007ebf46c3782097541
ze094108be50132cbc0a2b87887e643fded98fa2f64d772e819947b9364484a64a2c6e6fcdc5f68
z5a15ffbbf53d336c9c6a04a2e452f0fe982f950c6a47bd00b456eeba7de41533e7e9957427dcfe
z8457d1042f6f5e522f2243a0adb447d85af977325fded9e0727b6ac3d725cb5ec02eecba72d1bb
z2e9bc8f2d067a8a79a798d37d34bcf935697794fbdf54898ed32a586ef7912ca070cffb1ffc202
z6aec0a8324393a560cfe339fa2f91a1dde079fe1883c3dd805fa3e49a76ec90ef8ac538835b76f
z399dbda7eb8dfc28ccabdadeea88d62ba0fef55e7cd16e4ea243a1c90b95ae9fa90480b83066a3
z2005c4b30b1318d9421de8c3e853219f285d8c42b0712cc775af696ccc469633d15f9f20c9d71e
z9e649df4926b2cdfba3efa99acb0ce1816896f7d65fd4bdbaa446c07a5c675109c4af8067051c6
zb9b83c5defa002f6c61867829a704ee9b360015801c2a3d3fa4212ca2b505e122a655fa9aa2bad
z41d67f8f6f9a6598b6aa5cfa0e8662c00c9cbcd35f0079f56e3c278e2ffa05caa052f60e464773
zd9f7379dff4448ef5172ca21dcaa2400b2ac8236f267b5c54f8fb946f82ed47a281b25f1bfc119
z8e033d666957c4f29a1d58154e8b90a83396c2ab6bbb224e8301d60bb4ef8f4260af5a82bb7153
zaaeb39bcc9e1c27e5cab89c43671e4e59bd927c74746e050bcbcb133f910a9cc325f18ab905c89
zf0fbf8240dcceaa2ce0508db35b55e96818f79de04c2a220a7f143e315aa1c8f83c542d1914a83
zd9d79ee3594fb5174027127a2252f868f63b1fc65c509fbcf44ede8ffe450325643e4ffac087d6
z623456db0e68d50350fd64b5f02605334e9c07a3f5eb8a726e011ed0c2f73c7a0b20f1a1a0b2e5
z210ad6c103ac05f57ee9c7442defd0a5bc1465004215cb67613afc6d5daa14cb297ded5ebec138
z7479b8fa74bb2e1584d912797527ae321b820b4b9737d4e15634410551937931ee803b2b17cc62
z44cbbdfe10486e7bdf052be850d6ccf511224f0c266a0bafdc265447c736aa597ea1c440e9fb3a
zef97cffa10159159cb96f9f97c002d5b27d298ba45ab80f78b35c2fee5a97f5c6f52525975dd81
ze0b9fa3fa7b7642b33459b005ccd5c7049c16f34f99cc7b605e08fa422aa68540b68a8b1e888b4
z30d0312641fc372bf25a74872c3ceb5dc78a4c8c09119fb3ae7683b7fe4b1017b868df78b5816e
za264344d4964d337045ddc297f5cd26f08a0732d49aa141a23840dc33af4df50c55f29e3441b16
z9748a11f035de3d20e60ff31956f5db405f15d78b4307942940e4d0b1282ada3e2b59ca0c88630
zebeec725633e1a20e90e41748ccfce8028ed22956967eeacd87643195babd9bf6143af0eaa5f20
z53d0d7423ae00a1af622c76958d6223e34e17bc6c4d88a3c34bf4f25c00f583096b272a4fa318a
z98cff733cd2690684f694a431cd64b44df661bc4c67b6ac92b4c68a2b984a3ab518e3e6ecf7d78
z27f10d7599fa6e5c90e4b23492891bf8d54b1106aeb1e72210da51a93f9f359969d09337a655d8
zeba4f291ec95f9bf7b8b3a1e7d0ddcf4a7e99d5acde3ad207f2ad063e28ea1db5d1797ce8b1ec3
z2a5d15f2ba9c9ec5aaf6b916ed9ee54b36a6c3cdafacb0752f389b23a7b8dc250ef34db5e94174
zaabd1d09f9695bb228a75cf3f8db8a3ddbbc453e465b6da96e20b04e3d4c8ba38905758e819161
z1f442333c386217307a8292408a2ecfe5e9e3f9fafa8328d794d33ebe4c6444957edc61bfc29ff
zf75e41f50cb9dc53741988f7148d31fae327c26a53ffc69a9754a0bcbc82b5bd7b30b58b936b9c
zfa91a49dd0430bfb34f513d8806982a504ea5710229e4127bd240559a6d70fb7f8d50ebff56877
z02d823c2a8b4ec5c22ea17846e75c879ad0db6a38d6c0d0ce9ef19cde1e2a9bf9b95809b1d83ac
z11ffadcf15eca8989c75a285b178d41e3c5c6ac12317833d2154383840f23d8cf0eee914f8bb89
z3361496a9ca6eda67c8aa510d30c47b6cc833ca624cc3655d0a9013d8f9ecb7fda8919ddc17825
zc557685ab458d3b6889fa9b401e0b3cfb576bed556b634c30ce22c5b2cd504f8a507d31510be26
z757fbc72aacd1a5bb94452d0eaf9f7f0d17920227d44555e6d76100d86f410a50f025cb1d60651
z3934e5a4111542d0e7f62cb8b33bd7a68801295ce0f439e3e2c074c340ca7396ea4a9406284915
z06d5f4eaffe0ced59c72f9d70f9a21ed5c8643f12e35ebcc6cc24f83a011e935758c3db6983e24
z4ea34f21cdecf20b35bcec2012e948c6d842a9d622a8179ff44bf95da5477d7a419151e61b7ccf
z4323d09336480dea34cdc7ca819f7c8cf5a746185352cb14cdf3ba55143e67e6063540bb1c1967
z021e20fcfed3648815b4c371d6f6442f6d0e97b00556c9d82dc6223cc215a5d3b9a18490103cfb
zd80e4fd03cab7c63d5e2a5572d4e05ebd5a979feb0367ea172e407cd0b53748058a57e3f4ddf3e
z482c56cb70bfb5ac37cbd243a84baa0995df6fbd00eabc6471f5e00d03ac88e1d3e5c2bf3e4407
zc5f5c4a729b5c790d3818644325143b94e14468de0c72a7dab5e08a0d38a279d8f9581aac6b5de
zb56195eb45dd45dff73f1db2fb5395f8f308ae90e6c69ef1a728465ec54edfe61f6d4f024f76ac
z79e3d6f08e7dda4b19fa2e41f28e312f182fab66245f56880d84cdc406c5b96e2a3ef891b2d05e
zd17496d0fa356aa99ca66b259f37feaa28eb9dab50c758faece743f90b2c54a030f0d132ff8204
zd68ad4248ceb072929bba54ce08108c795cc29878de0c8048072793ef290f53c03c4b73f074d63
z56a4be74025367c8a3f7c984ca75ff065f096a284c7c048a2c415d7543a10f17c7620ac0675574
zbc51de7870eff82c675b0e846031ff5485013e55634c4ea5c5d65c7a2a999b4672a4c8b7c8db96
zacead8cd5f6e325ee79fb69ff58908abaaa15e58d8cbe3f2b46b74b114abcdbbe837a057f0649f
zbb022fac2822fac5714309c77ac6bb1874a7387da0cfec4bab52bb8eb86249c6b7fe89ef00da22
z39ad5ffb99459a26cec830a78dfe034410cc4207e54e2a2cddb28f87d0a2ee85280819046ee32a
zb7689375cff0f938a9f2ed3b73e9d554ffd04c5167914052276d0b1da513deb8305646f7b94b1b
z71f0bb8e9b20648ebf27d25f76833e7b7f79c611b2b660dd456d67db42963d0cfe55948a7cbfd0
z701084ad78201306ead725be1b6289ffd08812bed649c101d0cd7bc76202b1b3360a22804577bf
z69d38a44ddc9186b20a18371a070f7acda2aedea471871e5179bbcd9dd476c6601bfffed059b9c
z0f710133676957d792748ed001469bcc9fb4205cf804ac2f4fa346fa461423acc6ccd485188464
za8b8e942d216d6faae9e2546e533b0b1f3b0ffc5dfc9389877571438d7b1a92644e33095965e79
zc0e6fc396f2d7c663f8670eb4ca2e867c244a66b199ecbc324c0a9025fe05eec30d5eb09482ff9
z0fbf06238b397f9a1b1388acf70f1f7a7f587b2b28f4506b4114cb156459034ffdf3038067dd94
zaaa77f07ffee0f3669f0c70fbe59ee5b21ec67a621ae310530079bd09e7776549916ab24201973
ze8e51b75de47fdb1ad3597ed5c91074a82453816d510508e9ce13bfb84dedfbd9da9e8ef8f8640
zfbe2ee88a098c4b5f82707050e22c62c108d05f22ccdf0c0de71c542cf4d6d06f2325fdd38167d
zcce8507445e8e6bf65999c57f88e510df17cb62e4fe95264a0200f79356de84b6ebcd67d6c1e7e
zc32b842795c20bf0d763630efeeee5dc575c6610e02c4c2bd3eb94c2daa25f08159ccc6d5b9789
zda558bb57a441ca06fd9af3b584bb187738da52b038b67ff0c0658f87421953be8e4645dd15dd0
z41d5fa11d207d409e7c111af79c2ad6d426e9c0662118527c8effe8e5bcee405e0daf626bcc2c2
zbd92e452477a08707f0edac835ef38334573a3d01efa562e32a27bdd1d57c6a136742c64907919
z4c4c727ece76bdb106ffb3d88200239baa5b135d68621139c8c65da69a1d3ad3bae7c1774e3be6
z30cfc30f308193ed36274f45b4e9dd1d5392fc61ea91cab444aa74894cdceaeee8b27778d893b4
z75f7ec498f8a83ec399675335727c507c14fd3604a41c9bfc87c1ebca2ef08f7a346c545b77e46
z375d9276d3f37b2402229d201eae691c139248d0a7645cdf488e2d37a9a6c9f2ebfb87d3ea40da
zee2453abd51f3722cd856911ce6e0dab490c391de5f2f37b2c9b5bc9df464b9cb1d1e28ec43db3
z7eb0c4c3a6237c33b9bf69589cb2ab6a0939fb5278fe29d1fc6cbbdde4f813eafce22c78cc7258
zc832f6f5bb150d6cf3e2abdefc725fc2495b5a66aa286d99facf9eea9a0d11b6136e204d9ae6d9
zc26a7d48a44b4fdf5b1ec3b330d9d8902bdc84a00939e24fbb0705dbadb3e99db26504fed54f9e
zaa83cbf5e557d42bbbee148e76f992f7a5deaf00dffd6645f9031ae62457cc951b2cc355cdb0a7
z5104baf16043cafb2feeb1840d36d2a027e9928ee31720b60cfff2452c1566766da2cf309844ba
z525a171966442c674212677762e39cc544da4bac5ebd77823a68ecf45d23681e1011280f463b32
zf3a8dbe306d3f903e15d073bcb7fffa4a2f5efaa511f0fe6fd45016bff636603514c1418d014c1
zf856c62cc369d525625b59dcd5fc02f81e83db871927a852c6e4c60ca81c90fe7e829df3240b4a
z7d865e7b47ba02c1ab03928772c62ab3482a3514635f0a4c1d2ecb87aa71779034d1428d0cee96
z3c9696d6abb484ea025443a6fcdb7c8e940441b757fd59ba5c77131024b8065fec6dda1c0e1d42
z2760453c60bc15f80e71a847f0b916277db5b7073f7101e13364428ff8a102b6dccce79883d666
zda1ee714e972b71b27bbb266377fedc87d8d130f741349a2e1ff2340c299b9e6b9b5e6288febdc
ze067bd45b55a833e38e6a1c3facbf3275b54886b0c10203ea94367a51c9c36345d89e2818acb11
z55e0d2523b5832824aa50d055b2459d81d944a954394d7bc1d42e94458d2c1f095780b9f00c9cb
z36120271fff504f546dc7d6741987a832767e68a0b23d08caddb25dd6b9c72f4642c1a78c512f4
z3dcf24c78587cac80b1eeca2b3161f636926309e4b00aa8e9c146f84ef21f9b69a5de7047cb553
z5cb9befbc6dd484350e42b526bdff589ca5d26587211d8cf73ef2f89f1df9a1767993db0c170f0
zed2293d63d6194d5365e711140049474303011240d57aa53bac45b81596751f0606adc62f072cb
z5e27d616f46fd8f87b3c34d23cccd75dddc600fa64849e814e1c213dfcb342ca9d72f11c64cdac
z1ee2c3e6289dd9418253a3b66af98352f898935ba9f1301c8ef8308113eb26dd19acb834671ede
zbf8eff98833c6c8662000aedf2cf8e467d35a9fe5853ac3c9cb8f1b1a2b9c5c8942363c2784bec
z91b452a1574ef2431af8e256bdad31c30a6aa90125731a5e51305820840063972f52ae7299b015
z151b6fe4224533dd206db55d4af1e97d5e003d1ffa45cd7fa31d00737b29e38d08fece190c6ea3
ze13256bdc4f6eff7dd2a34995927f41160620db1936726a8cf4354bd0a173fc02217fdc4f70a42
z3f04e2651d12aa270af70c70ad164e681e70ff9769cfec472aabf065cf125e68b7a8348ba68454
zf5c31adf4bdaeecff922c03d78a11866aec9f1728c623dc51efdda7fffbf7ed1c2549d276267f3
z1653cfa14c1becaff8489d9cdea43ab3f807e00578ede7eb8f853f5a0dcc0f5aaa732ace15c23e
z1916015378dbb07a7c114a073b1e2c4e7c6f970647818b0560c01eebaea0b212a552a3814dc3b3
z1f7f54f5b42ddd34ca9b5bf7878ad11031b1d1aa2a251a2da3fbf221db9c961a5af5fa87292e66
z2f884e3f067da3248b2e2f74030ea6c8def5cea5ff35010b2ca95ee616a84599ba91434615ec6d
z8cd4b58c35da697c5448d3668b72b8145d3d8661c63422cd406fcc2857697755530811a2a10f88
z78baa640dfb863141564a18d4651dd3cb63fcc82abd4d23361a343594350fef9f4117e4a6f2971
zb6c34ed8609dfcb9aee88c6ddd6aaea674323894f04a5a87571a53af6c5b3df12f3f20d9dba676
zd731c4dac04d731e67880ba0b6ff1cde7ac7a73d1e9edbf8834dcc012daaeb514d6d6d0ad00a92
z3424e159f42b5dc858c9b28b1919b5c492927076c7df731fff9f2d358605407926fd051e8d5851
z9f94a2a320363cf94d6d8dcded37cf5e48a05bccfb70e4bef5f4b6d155dffe151eab808682bda0
z058e4c08103cd0dd8f9ef4b0696f0e878266bd5077e74ac200343853a5abee337f0d15440c5526
z22fc2f3b864245ce2bbdc7888ad6b5fb2eaf2e244519dcb92c61d34db064fa2d7eb48565c64d74
zf2b633dda92adfdbbda3861d09e57fff1868243791ea8e0917b4b173c25ed9a16780be12ae08a3
zec1936420899ef8ecc1d8d7e0a30366530434dff3d93d63153fd33f7d60c206128decc4a4b4683
z33bef951424f7aa8e795ff2bbd932d5f257722d265b0ffde609b3ca8b09cca441d0f264765b2aa
zf815a4d2ac1121d03cbb793d2b6f7ea4dfff96615d01753374cf6a84475a60f5e7d1044f1ee7bd
z331e118cfb3c34795780d8d895d10a57bd0a0c154ebfcf41a34278514008674295b65a414abcc9
z7323b1c3ff25327ec034b2a78f26f0c8c5340c214aa25f13968aa9a8890bef193eba24f2cc38bc
z218161e86130db8cb0fdfdf26716ce0633ac99caaca25ee6c7ffdc08c183d22802778b08fa5022
z00800a3e5246d54a144f746a868283c0db1bcc6db6a36a3036dc4285d4a896eafb609f73d79645
zc883c4599a86fc7a018dcfb97b3d0b0edde944beab3962a2d346896f4f0dfbd069689c29874c2c
ze983930c39508ef9d1e7c06cd835ff08b5881b228e8ade935e995cbb95396d796f18df205c10b4
za3e0f774553a55a1bd1b77ab6dc1ca37dce0581c9ebf6006f80830023208fb0cfa8bcbc9a4bfd8
z1f7b34ab96432b61734ef40bee657e9dcf498381eb10b31346c8c61f407f77f31fc8fd5613e73b
z71039bfac0649e1ced1b73a10d12e01d00d7edf5976c334a4ab8ea9a81f2bb245a7f48cfb51f65
z5d0d7e49fb5d1260f2bcc055a37de4435df54a74a43906dc0f4a457f8d8e2c1f666bca243901ba
z3f1c90c964c3eb3818b6a96ac57b36e90fd35ab28568e94cb7bb7db72bd47fc606b89e5f7149fe
zb2c6e7bb37ce64e2e348d652bc9c2dffbb61dceb4feb9c7130a17341755e6f52e42ef0a6d71267
z59738c632e513f526ba2ce4222bfc63634283ab5989e703fee412cf658a2d2baa92e7a8702211c
z89ec313a1cd745b1a9d27d6a4e2a0da4ae4aad4d3a107ba28b7528667f3b707a9ff01f13fb324e
za4a12d13918972a85bbbde8dea86e63b99a394df7765180eb84c13c055c281f510680542a26436
z6f6752e20cdd83a52943a19d747c827ae0744d4f8c49eb55e5986dd76ff14456523cca388d83e3
z9fcc8a427fb1c55c462c6371171e09516bc550da642c3760e0d7e4c3abcac688ba9ab427c870c9
z53f286a34ca22b845db69d3116dbf3faae3d91f906a857e3e135b66fdaefab91b87b5138bcbd45
z013b4621ab911b23571fc72ffaff01d70d3f311800ce2c3db7f76a06c16fd410ab0604bf2f0bc2
ze8b0a332123d0808f8698fe876cd44a75b6a7db7655199f64f2b9307ab9911e7fce263f41f2b1c
z3ac6c15b4cf4dbbd62c7203dec0e021b3e2eef1d69096ff1f2813969c922213a27d9a3b2a31dbc
z946da3c0f777eeaedc547b05adbca208bf6b8d21816df4519757dcfa4900d229aff9a38599fdb7
z2844f34d6412e231cc665e4ccf062b583bd6a90e7df14a5d53ac16b45ee5079a02131ec34b00ec
zf23f081cc213e155e721abfb893425bdf1dae4eafda6af8741c53bdd643e3dadb9ce65cd9b74bb
zf7643f768344686b24cbecc50378336ee95dd1106d5489ea32b0a8421362182e7caa9eb3754252
z9ab2a8705f60da3ada7c21045676c66d58f90e89af0fe2d3c56bd430d730b5334d910ab0b0ab31
zbced878a36292baae4d190ea65c274685a594868e57262b8cc5207ee645884d6608dbef25eb163
za7cd9ff11c517046cc98dd818acfd7f05a615a42a75e0aa088d6d9482d48ed6b3080ad20f8ac4f
zdc3ebb5e6f97c282cd40042f3f74d4095281d1d002317f1b038326d8badce0635769c52bab92a2
z625fd7e57028b7280e7c581244f24d8581c081d6875ae5febff0ba542e33d1e506fa7b3f3148f4
zfe1148cc8ca9acff67614a8365fc533f2e7f247efe54b108d8cde14776bc9bd32651026a6f9623
z8d4e82521fe02f4c00523434bcee8ca38e2e74e818a7bd127424148c32f4d7b8d03c84d6e50dd6
z21075c3c2a8195593002e2932ab0084423878ec17f109053e28a2b61b7ee3c95a01b56227a7962
z119b7589bf464b29937fc6d14bddecde864c314e64c7695fb606a0c928f80bd39bd3bfb9c54a38
zd150d4043e3e6b4dbd95f3b43b716ecfa525fe163f7664a508f1d2fca152db0706ffb6822fe16a
zaf94e1b34f507013dbc887237dc6f4dda4ec92147a9418135ad36df9636c6bf45bbaaed0c85aab
zcac0760900c0b5d941287b9ff5dec5003372a7cbccda6675f0a51f583c9dcb54fa732456996001
z08135322e785b6ef3f58143782def6beb7b867142d6d6bc265e763e2a11f857181a466d3b2540c
zd6183797674514891fdfa011c4613c686fdf646ca77e67ffbde49794bf26ea1a1fbee161121653
z2d245e8ecbcd645db63a001d93b5c63b701bb5aa310e85ccf84e5ab6f121a71b0fb32157a53744
z8c49a5dee2fba40331f38386cb28bb3b96f40a7d85812e1eae153b941e48826a63ac8c4002d3fc
zf4fbdd7c95de83166f72803e58cbbb0f405dda1571f8cb5f3cf24cafd50238249a4cc11cb0018c
zd69314010e9d0828444fae7c167c937fe33a6a1e8c40c0067cd644fb936a86f905d5a91df368dd
z824290de16e91a13a2d267dd62645fc9a16bf6c897f88f4334a31ba7895ab99ff2ce012b750a44
z0043091579703d1e546aeae7f26d846ff217d37568c10ab58bbdd78293cffe15a8b572815aa372
z3e3000011f673cf75503199a8aa482f89ce2dd3e093e087cb386f4434ece8c9ab2352c4bbb359e
z77688513adad6628bf7bf1bfaa5b85f82226d4787348386d4d2c6abbc47e0094497605b619f5e2
zdc7b966dbfb57c4611547bbf32df621f45b7de50f1387e6d0782f1469976d944e810be9bf41ad6
z9613859de5e253aaffe8c3eb97221db358fe25b946fe3bd6f34880e5350a5e09e69f0f7708879d
zc3ad77c0ed185b013b6b86e13f03b2db9c9f5298470d12d78aff34f781308df3c34c1a6c2316a6
z624b30ef3e065e46fae98305cca707609b630be1489977830aa1a8eabedd234d1000f3727e985c
z958f1240c7525c3860c5f9d9c6be8d41f420da0327d79c13c559a364c523bc0105cf26b6926e48
za0c86bd66a6eb045c79dd6ebb579b8c46bfa5e8274e86540de03d881fbd29145a4b1952e66a2e5
z53f4226ef4531b034b41999023784d602a55eee61b6b97f036a1fcdf94384c4900fe3725cb4658
zbb4c322196c640a1e39abb27051d76b9e78a409d857c0495dde9193975ec5b9d984866c2ba5c9a
z1ddafffe9edecd600cd0e08a6bbc042186cf2d850dc40d2abfb37f0dacde63a89becf41bdb6d15
z3f6aea64086129bf9e58cbaeeaafea12ebc190f5d9b3a55758ffd7edd1dd7521af1c565bed083f
z4de58600686700d152ba52cb14b43065b865a63c31951107ccb9b1f12eed8ef7eb647229720819
z1671e65bce47025ada4fef395836bf80667571b60c9268bfb82cf1df59e6de87d8b76952c488cc
zb320076e2e695219fd3ee3fa567023a6c9dd3ff8697afdac3261b59726806b7cca9b0aa5c746bd
z213337b489c78096f78d749547633984ddce40c35348c4c9c53fb3c6117cf80c635e90b4774987
z702f1be4d719a2f7750f2393d53273bede9de277cece141af0ac3aeba3d696d9815229b7dd57a0
z9289a6333d0c28721ed4b43bde4e44b721da5a457a57acc3b715e0a51220c6595e359b5a9785f5
z40b360a6a226ab6aef30bb6457ad2bf1018252985d2d90b4d9aa80525d88d5d7addd9d010e0ff8
z5baa6beb9bb5a334d51c819223e8f4c6e1ac120b1919bd7ae940e69fadc409e33c30f0ef3bec3e
z814146eba2337478a96ddbd401be8bbc418eda70743bd53cde7dcc6c280f9fd67521c3642f5a80
z5cca09f5fa7419961b7625621e98b393620816556ef1a0db88a85b1dbe5175e7291cb1846f7237
zeeb64a8903a97c1847cc3d617182a361dccd236c3ef7c99f673d03fa56d1348ebfce644defa214
z4812ffab61d51c02b4bff6ec467b40a70a2956c27d0003049744d69095defbe83d00d44d888101
z5a8e2c6f765b6437d0678e542d1abe3ca1f41fb800bcd7ba3e8d0bc50bdc72eec0aead6033fa66
za323beb24d93a57fcdb88e9e7ba4d5be042d879c1e4a3306664ebd386d8804c8cd0a8d5b0e7bc4
z78b8f4437ab106643fe34e0ae8868e09320b71ae8899c4973d1308f0c6823997bb4347108fa0c5
z5db6ffc096f1f1afe771a5a75837031d7900b6a3332410c301d2979fd118fec36e0cf2cf1f190b
z11437e50d64d5193588e50ed201329fb8518c79b3180109f0524bb4991b0bf541aee598a5a6de1
z77abe24db2becbe12f78ad8fbd7bdf85fd6e9ffe52fba9fe011734182d2b0e6584cb21a7298f1a
zdaa7d88692aa56bbd6ff67dfb01d6b56208c660214f15286253f434c59095a6083c49f027d38ae
z8f499eb610c8928d33540cac6137b602f43e832639b661f06f886739ed4ba82fd3f25fc90ffd87
zfd9ad9802ec4832817c4050d0d25b27e2418e1dd4f47f315659c28e610f77a393c7dd1ded8004e
z5840ddf4e3cec1a233f5f7c7ae60b769d2a1777757dd0a5b21d38af151a13893af593539c70773
ze63effced5ce359a09e49a57487118a9221aa61926bf0b64b6f0a148f128020390cc0c547d1588
zff27974424653e117e898c0b841e0eb7ad3d47904436e1b894c7ce0b6e3a73aaf59b003e28e3c1
z77e48d0f15501e37d4ef06173de86939e947eb5780ba77efb4265f1733a332bd21784b42f68552
z5fea1678ee7630106aed99f174163bfd529dfdf6c2288fb4dd9468ccd061db9d7753f0ae222079
zcb96a82ec39b644591762a0dd8a18565c1d29bdf3d8ad584e8e241f001d83caab3ad95fe5e33de
z72eb5d930940816ee76eb8888c32bc8a1df83cff9f8de31fcd8a9a6a324666a0e209b71d499c03
z8adfa50a0869289c96a5c3642fa871c15d6b8967aa716f25d5ff97fad14448362269ca5c5854d2
z0595dd9dd08d9631177309dcd9c655d99aee84e1beee9daed905fe2710901bf8c9a324b245e573
zaea9d1d57be3d24b283ec9a131574110cce18769da61a951f361bb53eec425cc17541e77e74536
zb1ecfecbc5de1b1f1b5fb4f33db1930b6f8a7cbed2300bed117060ff9912cc37853a6ddb650ef2
zb865adc6efc39123c7a0b9af91cf845cf4e851e3be9e2222b152608b1084a16d7df4fbb5aa1895
z82b50bd5ef6e01dc1cf098bced9aff09954d07e607637de47721eadca7628aa79c9d2e577d986f
zacdbeb23e86e8aa313cb78a68dc04d0eec648bfe2b18cb2edc8d199e144375cdf9297a4a52a842
zda279107f335d461929ddf528e2b0e3f0776fd5fdf9b8e2abef1d3321b21ff55483671a6ef0199
z0cb0bdd49613f37b52f2549a81d52908bd77c6934d221de9acbc163a63eaf5a558d5fef0254ea4
z5524fe8c5389a850f2041839793951483c2864f3f708c32da88d2d85b2a0a519d756f6750013e8
zd277f56bdc8e5046e7690ee3e428c329b7484c75843030880b00a7cc694bd90994eeae6129f50e
zdb31d56d29a2705ba2cd8cb7d1a112b6d2d33258cd44133f56a1bdc06d23ae126bbe3029881adc
z3ddaacc46f184ee72c6bc110c95a462c7515fca6aca709ee2780b321ef86153fb3e9f8f99ab76a
z9110bc55dbe82597ef7abd23a58df3f6185f2feb611bd5d0a9df2b0fc56d337d424209ff4f5832
z64464ea70456212ea183e7f9170bc3dc357f9f6efd9d0b278d8fff6a8c9a60be204cd2b9564d6c
z747322eefec86557f3ff8722f6a4623179795164cacefa4bb9f97d78bc6389b5079f25626d9a5f
zc0697972d9ee27e44dd7ac2b15dcec40801d14989484a616bf7f033b3179e76619444cb83adaf2
z410547cf551982d85cb0537a755be0a1ef7a78202ce3115d09e9a40af7e42d3d22c409b199ba74
z1a107734ba3ecfc28354f2479154974929ba7901e2598858de40472010675b913d9a7e65c91d98
z093c591ecb25922b63f4658a3c4e2ddb5fb891d7f8872c8fb79a550b5e143b4331793935164436
ze56c545ef401151ac0fd1f9cd9ed6ebeaa1fa49b62d2f30d3783ad0981f791e464c6fe85f04356
z70165a42c5db250ef755ca78b863a963155174bce8431f675a3110793595f8030040c78aeb346c
z8ac70e2e50cebec5d29e8009b1de4e95c45ef25352177adbbd1231da4e8f733d9c4af9eb94a823
z916923e7b8320205a8cf27f69838437221b9d76cf8fff65ffe69e84f9e9da2871925937bbe4866
z26be795f30af8991b5bf44941c6d56949c704a6d67ed5dc3f27bda2a57314217334f3e4ce37b93
zb4c73894855200eb96eb4fe32654c5b4320488317492cd84d664036c2d8cb5413609e595fa5649
z3430f8f616f0a2c4502b6e33748719d201ed47ad591d3a15f4f78bc86e82bb70237d305cb9c5b0
z321fa4dfddd90ba810afe4fc1e1acf8710514272580d53fb6e7f75801494bea017351d9fcf71a3
z2beda701bbef0474949c9a70417bd8a3648db372abcc97c3aaaddb1b12924b323447b0d2c2bbec
z94ee33d9a18117abfe77e4cc3fefe44b38cb3e7cbd9f4493e378314d6d0bbbc6c32ec02d79623e
z9af4df4a517fc7f34b459b30887157a7ad879226cbef104ca06c429b1640bcc6cf223652ba4013
z2ee7c41187207b40c4ee6dbdb7198a6ac7460dac1c791f96c57e45976df4cd66670188ff0c5ecd
ze8eee53fd86ebb11a7c4f04476f9c61820af60264c5f7f861eec728afc7ba731587bbd254eda6b
z6acf4e889883dba596b4b51332e6fc5aff2d078d2108374a18c07ad9811cf913e11c4cf03e8220
z6123824aa1a9e0d3c9f1dffe2137319d3b1b1b8f6ffb31413ff62c7bdf8726ae2db4ad873056ce
z49c4df3278379a26305a8629a1a1ce50cf9b8bc72be1842e9dbcac94bda2122a11e12f8a860153
z77002981bd25311cd23a81daa88049c4cae99d4c6d517dc3d7fd3a987026a38003d03a17745f12
z08f036e999f6b2df4b3ed370cad1e6d96b3f1aa8e18ddbd627edba29cf16ce1e770dc6e3cef686
z4b7d4796193a87179d4b646a9c724a3c8a0c4bc05bfe7ca53541d3786aae60c191e059ded3053e
z1f0d306e84f619ec515736b6df8ff615ffc9ddb6c01efa7bd87181455f989054c08aaa1e99ed4d
z8047ef8c802444aebdf0ef2ab7f815ae20e4bbebac39b734036d4b9439d10ad7f43ac8b7444285
z8801e2b724079eb67ef735752ca8909a6bf51426bb7ad85295ee2a35a85b0a9d0c17148db5315f
z01bef47d1eb3624897b71a450b12ef57cfb450ab0afd5ab89100251ce1b75a17a4418fd90ba6a3
z4729c86e036bb243e668a80a00435aea940862e7589cab4dc67771b8358e6807d5279948ebd25f
z1247026ec26ada17dd2455f59ba4018e94f86d140f8826d2a004541a494fb860fb8836d8615451
zdc1cceb0feef1f72010d0779d857ce7762bbc5c16ccfb78da51fa1ecb2b38c8a386dcd191722ac
z05d5a4cf60792beb804e5623ab6a58d31a8473aeff93c3007d6a13e082c7580f2d812b6d657c82
ze16832caccf458c2f3847115b087cfaad447c3bbb6c7bf761b349c5686a5e5b043137099d4cc40
z893b460ac4a8720eccf09f9c484d615398946d6aedbd6efc87ea01506acba49e77dce7655e64e1
zc29f1e0b082c4e33024834d44b9f8b59150c1847d6d8de8014dc9aff4fa43dc1de78680d076a0a
z7518060e953dce74d6980295609c52afb4f1f6b976e51012305e4f1c161d64e567ae71b8c488d4
z08ee091dd78598f62c31552fa0c0fd7c88f494e641f0e88a80a5c42a9d87735356c23f3b351ba3
z1307fcf1c430f352257ea8466a140e303edf30ca92d4f6826e92fdbb16e2ff864c9d3eace202cd
z9bcc24b3cb26feff0029ab8d41a4a00023bbdbc3a7be48ffa6ac987184aba14c35247b2cc09dd2
za28c75a3ba5fcc8667e6c7e86d8dd71d35eed7b910372db923d6b62a0caf49432d224a3bd4a55f
z3f53cb254c472544372aa14f4dddb8c7a6949e95ae176d7bacd1b9df7b7a46047258b310d3488d
zc48f922054323a90990da490d2df55b8d3ae64bdc96fbaa796b66452d46e80a2455a1fb8ef82f8
z855722a70fcd818af938533e2865754766fe0b40613486a01062b1a34083e48165de299d0635f4
za648d0a31837e380c8c71037bdbfb9be4bf94fd83e820d1ed92ca241ba193b0f4067ce25f393d4
z80039d9c2f6b7fc1f2e91ff4c5ea9f17bb042fee85ecbe54729e783d4bc0785d3d39f4ac31411a
zaeda96b8b873fa166391d774a1ecf8566d1297cb700d62bd27490ba426530e86737e07b48a5fcf
z3394ef04f70d4a8c39812792beb04854327bfcc7ccf74c79eca341d466e0792f35cf2240ae9914
zd7131c40cd0795a984acf26ea33a71378e08fb777f3993418c029fecc83b2198a307b4331be757
z9838dc820a2b9259e1488defca2ea3e9a2ac407d271d749b932713f2e80914e2cb5aa2e495f231
za9d6c67ebe569716383f798f32dcfe5eaf79fb989babfd2356ab2366125d7460534b99aabfe5a8
z2b475bdc19459ea7003421eb1eced25c42bbe7f4ed9fda63c0836ab61444c2c4c5bcf5df1def23
zb1689fe1e8ecfd3618d704fd7a75e3f84d6ee49da49656877b441d22d45df119738a43c0ad7b44
zfe1511ea8512b466f4938289d9e0305cb4fc0e2818ce98a426a562ccf881458754fe4e690f966a
z4a04760e47f9592a0e586bc956048c4f1b733e531611e977430daa99b97f6e391129afbfecca48
zd1fdbdd46637e3785fdbbdd9e1bfb7d3d3bb548bf03ff4157828a2f1e86d5ac6f0b5cabf3635bc
z7a2836dfaa46429ad52adcbd86c425ad1ed3bd580760cb3be92e8355e8ae2ca4bf21647f644b1a
z87509f1b1e8480d4e1101cdacb2b4a90613fde9c982f4a12b23d920200ba0ff71e9f584cda03cd
zead75e5566f90013fa2791b4834cfc271f559b3edbcdb13c9590a5f690be535ec5fa49eb578315
z3815c30d5f68a076df7ea01a42dad4a67143d9fcd3a93c76b83e53f6628b7a8905922e93bbfc17
z0167423bf15dfd8195c652a5844e6bc620726c6017a7620d1a1c4d666c9e581064c55fa3b6d199
z64056bdaffb9014eec0a6e81f608426a5fa89cd83f552f2eb9b125042ee6aac84e66c7bc30ccb6
z12a2383d68d30dc62373d17c92818bee612b6af2d3b79ab88a995e4cb9a672fcc427adcbe35de7
z225bdaffd560e773fad7113b81da8c684b331a67fe3a2b72c36b9537f4ee87a619b08e1de083ae
z6313871324e3fcdee7d4fa0bc64fa0b5c24ee211f8b52d9708721a30c8b5540789d130b839e5a9
z9feca33d88a349f22a4c720c7e914cc4845d788f6dc588cd07a75968c19867271198bb83a9b57b
z19036b7a6a6490af14498b8b9789a4805befd9a095aa3882ec7694aea1915a6bd47f50ff9f00f4
zfa77ecaa5106de35569f39717b8e0047b5fcf07b394180a2dc2f5f0e1300b28848913582eed9bf
zba3600e280b10e21671190a5ac591ef9725076d03da3d8a4f47a9c598480192fd44c8b832717d6
z559496c00e943e369aba27842978d9d41b0b8f96846fe42583c48369627d3880c408867cafc7df
z083cbaa7a4faf9efebe70f214159c44d155c0675d53be4f13e985db870cafad8c4102e057537f5
zb9928f39ddb9669fea015bfa49ca67348c084109d2a871c2df78397fe0d774a63f4dd8558fae4f
z7e3d1b7bad3f7bdf9a94727e5c3dab568b2feddec2cee0e9572b3cefabbd2b42c574b9cd7be71f
z9a0f8cff3e591b585d2342f6084fed82ad48be6a424fc36152b56fd697c03e6151297cf146464a
zcab3bcc9e7a7f8a676be8fc0503fb55019f88a2263922402fb1a1f1aac11f1a98f7aca315b8dc1
z3621bd3c85bba68735801ebb354308a247407e78ccf2757ab4c2b0d42b85f4f18353d5e846202b
z973305ab8156bef01ea7dbb59fc7b7e5ed6db51020bb4da65c1d875fe113ceb5673caafa3f50a9
zc974d4a70b6546fe99e551ccb46bf38b3fc8558e71041d8c8488c371616ee6788f160c7d2afdf9
z6f90e7cdaf5febcdee519ca51ea2e55626fae79b05fb45ed04d970958af3e31ed35833b879e3f7
z612e63cc02a771ed74a2a79d23443b9d894ba845b29cba79f4e154870b70c755a9551d7c21d3fe
zff739b1d8983080cb5d7b84ab5965106a63014abb0e655a8b614b7ffcbe3896fd0ea999f1974a5
zf5de15bcb5288e71b3b4f726e0aaf309ef1ee3782cbb043f0052cda04563e2eef7c1c4b0bba8cf
zf7e55c5f4e964598cff0cd0606d123580e4a408695a3947fe1ba28d9eefc8866aaa4d545af5803
zd15757a93ccfd8cb674c44c8baf1a8098ef2eb2bd4be801d63b7287385914954665e8ab31fec28
zcd218ffb8e1aee2fa6fac2a1994f6702df23308deb9c3ea5d188b97b7ccc43d30823b6d30875d0
z90d047bb66d9aff4a72d6213b6cd1737d1b797f31320b3d460f90c4a24f9cf976a2e045675207d
z722f40de4c38120aa0cc4a26ca4ddc278540443157872b4944a2a2ed15c0c14a43e27c9a222b21
zb8f72989acc1e1a4b8d8eff6f5110fca4c73750e8d5310ea6489a55ebe7553ad36a59d789e3e3a
z2498eb586303bc4baf791e7a47f4f116990141c76dc647bd89ffaaffde49b2d59382b6370c3a0c
z96b12b7b3cbe3b07fd0766d9ccf64dda4047aed7adba9cd9e0a3b3a3c63fdcbbb699f951c0ebd2
zfab0a1ee7410c1ad8eaabe24a00f68e1d477f5a88a8ae6789a18b83f35a24af8baddeaef700c48
zaf6d5fb4aaa47cc0c4bb236c6abd2bfe122516448866ea362c81001172c657077131e02e3b8b54
z3bef63d99b17f51bead4f307bc78e72a0305b9083d2b1be01fd8975c0f47cfc027b35be910ed31
z897773c6f355f07779bde50c61d439b6b872524e0faeb6fcfac8d12e4fbe2296acaaf4629ce390
z60219b6f507676e16277439bda3a368b554a36bc0a22f67ebdafe712a57ba47dfb91ee516d067f
zdf52dfb207cd6e6f17a29714351498a16139992074036e191439d51a76c7f5b1c68407045ab429
zf04b0cb21c768307e361087559cdb81cf1c4f94ad0bc901dfb9f330a43c7003162036a1843a0cb
z7e5c859f0d414f1e222e64822e3d22f180755138740841f3937c18d36b78dddbc35e1cd67d622b
z344c3aac18eb312ef8743ac9441a74557b5dd3322170fc6f0ad837e0d60324338c205a0aeaab17
z1573198cb6d29de5e6d438ac6d3006270739feb37ca010ea123def722bd2f5d749fb4c489a03c4
z63884f06f2464dce2717f67675a89a7413b86a2dae572334a19139a21b0dc781f928b21c542871
z93c4c96605f1ae60b0cb46b1855b936c5928f62594c3809345a3c356c0913980e43ce658886f62
zc21c907746827d1d2c3bdb61f9d54f0b32aca933eb3cf4c52622d49300774acd4f9fbaeef3dc69
z1a3b5e68e7e653929e68e631ec97747c016c4419337f53e9c8160583723cd1b7b3aa08ec2306eb
z137b44271cb9f86f96b95ba3022fe623e1535656e5b3ae7f48e2c97879b4ad9b158206eb56a1fa
z72dcaa1f0bb807ec09788ce3b8f5f3985b262480ff1fea4329e26af632cd08fe1729739eaffc69
zb11ea65a791ae9c621f79e40bd7315e6742bde37265a01508ac53ea5a077a3d6cac73fc04f88bb
z74b95ef1ad45ac762c4dc5fd1390023863b464833f10287bf86f3d6e1b03825f0bf181e7595fd8
zd5bd103a66272fb36f8706a108a1ac21821850e494190cd8367f0e708da666a28b428fa3b9b0c6
zd75483dcafc7a9ab6e6c318083e32b8d9984687991477b2327c2a83fd6af6abfd605b23c661e6d
zc2fccaf96a2d92167840f92c7876498791a3eb188410457e5c2090d2916552142d49ae5059da85
zdcef12830eba3b9b6f9eeaee136d38fa99e2bf9a33caba621248ada23ef21ecc69fec741642948
z66cb25255baaa12ddec18693f326344dca448b54a0cc07b93259314197ff604178aee285e13378
zd5d30f47e5c7d0dac2d766e8317d34e5db36103d9e6db7c8c96bf55d5dd008cc39cf0f9f000b1d
zc54db733aaba35c40ff3d9e0d5814006d412bcc9607b6f5e1ec934452ccff33a0cb849d99ae9d4
z33177f0ed130e6e6c1dfe3050ca85a15ec4814074a7b3d8e45837537e98183d2dc4caec77e00bc
z55dec6674b01d92ae4bef54b28e9775976bf4801e52bc90b3097a0655e5bcb4a8d5dbb07e72404
z5198f071b3bbe8f0941c6afdc98c1eb29183c40274ae9e570f0cffd8587c5dad86266509310808
zad0a2bee7065d70ccf0b68c6a862f41e1203971a975633ff8d19892c44950d12dcc59a2e7e6e03
z31a8bc61d9595bdd51d43548186332d3e0b2cacf7cff45658d2305cc8f699c18269e715ad74381
zd7099b574bf3d4f222df4796c01b1c7527da63e87f368179185aa07c8c7dabf2e2a84c04aeabb2
z5fb99e6171b8a529766de3d6639023cd2ecac3b18c9c8f7c5741365f857104500d4e5d437fef89
z33b2d11b4686f17a1d7df422593f820ca38564565373301ad0e40f221c1fe82436ab83f544d2fb
z62f467d7a6bddd84a45bbdcbe2d0b6e4d3b0fc9927e4734796964c33e8a16e3e7578b8bb948b74
ze372714af353199a82bb52bf738462c0695360a022ea692b91f721e54d42f67873b1d7c4a95aee
z447da72fb90d04a1b7753d9fc5bdda2a9640f001a7b8da0ccf627bbc92de829d7331a59111b511
z3f8e817c8d40ef67ed67fbcd386ee6e6d9219238debaabcaed49fe232c1511e93afcd8c5ea6ded
z3877dc7f847f31f7495fe2ee5be321d6f80cd23a14e82d9fa03644e9e8756b7ba699c760e35f0e
z5cb9274e0675c5d960e99a885e1e55b0365bf8e1ac786f6ab2e28a49f8b9529ceb684fa0534491
z0413ea79eb0cfc7a51224b42c596dd30086c251c73cc0525b4ba6e9f440a8d36d0fbf63be21a1a
z806753b7f4cd9ed3be7caebb6b9f46360bed3aed8750b4edb3fec5dc4dcb3ea8076201d7575583
z228a17a8b9ac91782efd50731f0f5df52a705b43db5766f1ec6816cd02dc7ad0f59b8b43ce9883
zb85a13157ec05fa6812c66fa1f0ead088d3503cbae105595a932f943d790014891ba1f1bc5dc70
z112fd07ceac2953aa84a5a970d0e016a1d2ef216531cb9b8b1bcc1b7a9640cf4cf53844649c62b
zbfea8db88a74ac05a5bf57db4d75acffa36e7d7cb5f4dff2326395c75f1620e071c08e7e6b1dee
z91e0fc8470fb62f242bf8f9e60d1af5aea4ed67efd92495f33b7aeaf8fc259475ca2ee78dc2961
z065e73ede72ddb4874c0e12f3a994d86d69f6e3e4630d71276ee6acec1c184d42040669d13ddcf
zb242bdafa8126b0022512173e61c18e839dad28338394e89abcbe969251fa928a924263bc726f1
z61674c0fa77c89f1ddab231a2fb3f67a3f8ea095de3736037aee45b6427b01e42f39fee31c761b
z18cd02d7b24f38e96ee989c967623ee1fe35bd80ed971624e196f76a88f14e50c7a7e335818c6e
ze49e2221b1ec1024516ba0221311c3a2313758b3c5032aeb1589e8647ff985e02f04dcf3ba6d25
zdeac83e63974bafcf94d1d130d823fd11f4497dcddbc0f1cad6f0211d052adad5551774f895d25
z29f8b4ced2fb09a71b9004e77ddd0205edeb1b47376d355043f8a76200cfd7fb1430255b7f8b5c
za4fa988630f612268b30e0edd152195dd8234ab7ad89fd633f1b3f587f2c35d9c4fa53c222c41e
zea36b9a5df113018b252e1324d999bbc3f15e463bbcf02c9f10b21d7cdb7d9067c4f97e87e5d22
zcf5787ea91ee81546199f30d5f55b3457152c4b4185f3503b48c554511f0a653a81295bd13648e
z4f48c0be8c65a5d17d8744005ac5d8ce69cff0e9240585decc758be21d6b3274cc06af602cc9ba
za73865fab6b3f75edf466f61435e4fedbf4b978b911825a6f5fd783f95f52e0cd48fb244083b56
z47ff5147dcee94ab7e8519e075ca2910921bbc9f445ff87626a08c4d1d7de095110c6047b7b657
zb5268995ed2cea20e2581167e5b349a8c5f3da94994f6e50f100048ad2dad2242a34e97155089b
z069cea5dd2c64fe9d43d861b198911f43e008d6f501af48373b40d9253bc389e02e57c9ff6e70c
z8d7823131f1a049a688903a0270d85bb995a5034369229c266ff9829bd7506c058b7039d5688a7
z598f541123a797511177a92f7dd139e19e8300c160972bff67fde2abce7094606fe1980a77da2e
z8a8070817a9bc6cbfd44d7fda0f5a6111282a851d3bd8c6f7933c8fa710bcb61400c1e0f1ced0b
z6d208f66bf5c35aa011c79be8224d5123accd72230363c743f44866977d83725929a9677aff3ca
z272c164e14b4c7cd097254a13f9a6480a894f18bebb1ac1cbbef6fc8868acdec2bb814a35bc7b2
z8b02011cf09617fe0829d12acaf9bf4d5353d22e1d0e691a6bdae341d8f82b5dc7552f578f8733
zf8fda83fd44aed49c4c84a42d53e3f760cd7315005be5f22eb482e294522902bc2ebfc3a785861
z84cb9436b09b01e1556f0f0a2d0ae279158f6f08ee4ed695618059b404c2506911afc3bdd7a697
z22ab86809067a42257a0ee9d21ff1d8788b0a0a3474d0843b30c6e12ccbc88a681f2836710c7fe
z03eb2d218b21e9031b34828179ced653131a1ef55d0da18bc03bfba40b98b3978a7e790eb09c64
z0bfc9cbdb796f04b15fb73288cef951a04e56f9cdb3638bbb7dcaa5202f1053f55ed8d8da0f0d7
z8780991378eb2be31f27dbf862957e5c8cd8cbcd9af86369489f348b7035f6ec8cb07be8d58fbf
z06ef35d96a74a656b26f4b6b151bdaefe3aad7e79c1079609a1864ea7459637cd1bd9ce3a9165d
z6f8e06fe1efa1da4cdc3fde314c8f1f0456d51756177d491e46a95c1c62a69b1bfb1f99d9cdab2
z7902ec59b10e59c84de98f1c29dca56a8124b1d00fe42c46eb0e41604e1d154aeaa2eecefe0ae0
ze2b68ec26460310e400610914ed7bad5a759b6e00bf477045ed2eb3ed6fd1784ec1db8cc400315
z074d0efd502ecfc9158424f0ea5e74b78f8df4a3383242a4d396ce44b35b57c6605e2ef985074c
z4294df85d243baf8f0e6c9ed8a83beebf234f5e1f4cbc7875622839f1542f6aca5d845073744f7
za8e0bf74e613e3653a402c83b6a85a8f8d55428cb75201bcd641b87f7892d46f78ec223ddd18d8
z96ce1c319f520631ba91900b576b172a548490c5502a42e91441533aa4c2d2a50be5e1202b0eb8
z220ef89cf7d29902fe99b5cdb906f38912c172fc10b727fa8f609aea1a9d8381235191e4f5ee12
z06d31bbf4103e737535cf39128ba6a56a3c3ca07ec000087cdf7c7ae1f2b066a50a7ad883f99b5
z181b4234c4fad9ab2189ad302c25f95363f51c0e3bfaafb4b2bfaa7f2f3d4629bb58430a5f969e
z20f2e60d1f60119297f8ef692a475528a053fe7f9e158a3a4860684e1530356ba9cc7687dafbe6
z00bbf097715f84a73ad72ed73dbe588091605ffe9d12523a1d94a150601e78356843fd104efa26
zbb908d05c7a7f9e77740b9a54e1cb3ba3bbc1e0991c106cf71fe5127170e5140750010e3885e7a
zc92d824ba4e9a0da71f3882bacec83c41ec0448cbbd94fa2270b6f79618040c9821bfc42690a7a
zf9e02dddcd55d7067ca9b4c623a289bc04181acab5e124c52291feff806b399394e929a879ab57
z54d5240a2baa0e03b97c6076069c4eee878f10d730bfbe3bf8863eaf321ddac9acbbac1ee76b1b
zc5df1e54c0388653a185a9e9b69b9edfdb0ff0c0229ed358f41990ba9b6c2afcaf611e8ab96f5d
z6b874302c193e3c16cd7ac8d1baf1c3922fdc26f314d03fe9dca78d6b44251903d0541690f1c4c
z5cacf9b865dd815641fc613cf9b3798953f00687aeb8af36d49dedfa3747ae0f85573076e9d420
z5be699ffd37e72c73a746a9203e4c66f9045a843210249dcbe3a3f1eaac91b54992abd753ad279
z32a7e5bc28bd05690ba0a4970ad61311fd82acf97c9b5f13ae4333f41a8d0d6e86e2e97e659e62
zd65b46659d270600a363cc9d0c8f48109a5139343bbcd08ed3937a75d2ffe89cb4ef3cfe418556
z628f457bcad816f2d4968fcb72677cc60567f79b733259e1620b632ade2b61d7802d5125358c4e
z4209b41ab6f521c7568ce968e28c9ab0a8b62562f74c713e11fa4f4c9604e58dda70612c7d7dae
z6abe599991efd157959e9541641209aa0a0efa7aa25cab402fd1497902b198399a44fea3ea99c1
z2224aaf34e5494cc0d1ae9e87594c05c35237157cfdb8f442f7ee8d8a8800f011b7108dcab7851
z992544f18a1d4b864e91f7c4fa8cd5faf88189a532c8a101d37f5facd597923cda8bb1ddf6ebbe
z6a12c5a049ad6818e63eb9f113df6015cc992557b1ea45c19c091f0fd94dbb672ad9aada779f37
za787745e77ddb30f55df378f674d9a6162f5f637028cf66d36b3fe8d02a13dbb3ccbcd8053c7a9
z2bdb2b58abbbd35d0727d33063e221a3630ad8823f611846311cb0defc700c42c45cac2e444cc7
zd5702b29e404fdb7604f7d7e7f9dcd9931c4543f5155a83f81b3015c16c7d4aacc083ca457559d
z363ab68e1d577b3eade84662364c60822aae7c78b816158b1a626d86f5a1e697202dbdd2bd0f87
z58d1efd26d7202e9f7090cee87013c4eb6d91beafc702ff46f4638ab31c0c91e9afeb25e6227b4
zea595a78968b4f370fc7d94c70429ccc5f8cc96c2661914f2fb34d8f3f75e5dcfa0718ac142de3
ze3499c3cb2fc1900306a6fd049689ba5436054647a1d392e3886fe92f07abfed631e09a02ff161
zf44910947819e2867bbfadc4563f8d9a6baadca8c3a3cde78c48405d8d52aa4df08abf0326fb22
z7be7c075a0a2e1285e29352df00c66d8344df7e8101b045fa404c8e6425c1d61e134f4bd0c35c5
zde8d6b6489d587b7f3350e3bb1deeded071bfd284b70b25654db3158286a11ef7ce587bf157daf
zb810e8d77d66fa0f22cd1f7c46902b7484505da9195e2c3966e06a71080420dbc03cf7cc01047d
z8b90de7920ee906cec40bfe2d91ed17e3c84d09ea0905f8666b52bb82b4cf50001efe8b151a15c
z76408084261c463d71f127dd2964159cff37e6591fa76b58a92b5edd105e133e649a3b21f7600d
z8300af63b47656a83dbb4ed2004a3b2850118017c26db2be319291161e11b4a7350d7950d26fa5
z7574fe9d30ffb1a1ab009c35cab5a74a8839421296f314add91f379edcf168ba8625a1443ecc38
zc8881071b883b51f6e256edfad946c5ca7bdbb37981f13e3d72099ed504c3aec8e1dbcf2c00203
zc191e227dd96d3ec1d7a91f6282e9822db6178d598109d68a37659b8b7b6b6c58bd8a6b87a831a
zbd7b3f47e9b4c147458a3d09dcb017558deb83b65ab7913828bae6b72e45e87be889e0dcc776a3
z43651dfc0e92714acdea5723775574dd338710080d516df231ee8e82ae30b2248158c8863efc6d
zf27d9c2ec98407b6894875ed49ee92c3470f8616067e11393ff23b9f0020c6b8ea446cdb21a496
z08b7603ff046c4f01b3b91ec664b360ec6bf4e53c05ed88ab872429620503be3e63c76966816cb
zb2ca37cb29b9f218ee6ee1a2f37e10626e12114f4f69cf95732702f4b9cfbd51a2a188de625fcc
z94e71d2a57b5bd8dc1ec8de3d6f15d921e1d06295178e1ac605ee8b3db857bc3a0a0bf2032a026
zdcddf3c41053ab0444f57a974a49b457609cde183054695044a858dc6df57fc0d0c8676022b1af
z6b29d8e2e78ac78f88d6bda4861f5d4f32a4eee93a47bfa88b41c6e50414141ab5cc0f9d7f0e57
z3e2dc52594b7011b060ff355d6429e826eaf1ff95b61942f422ed88ca34727062414b431af83a9
zd4f48d7a94f4e65a5a92b229cce1b1a60daed9a2351ce9576e59bc63b93a44db39c3e22bb4dfc2
z163753ced06b4bd726ab8f1ca8e8917b97c6ffad9cf13889ebcbe99c0e2f04120776720cd38fbf
zc7666f39648be14089f4ccb5029a6392f7f29b55b8ae6223311d0d57cae5e249edf6c4041b2934
z8e8e564a72f7bf66413a6597c9b81950267f71f0b6cb1e7e30f327ca1a0fe1d003700b74ac0209
z89bdcc0091983728128e22157dcd8cb42cb058c9744850a990c33cc06824a3582670e65473d23c
zedba5abf917a82685a344abceea9dcc0d1d0750078b6b863f7747d2a261d11c619d34be36a9823
z4ca009d81b1f27cda212126b243400a4e6fcfaf1cf0e5e76dab4a5caa854b2f999f52239576086
zf1afe1369923427614602c592c90e8b6b278b9cb135bb2f0f1d59c589eb1c62cbe803669bba0d3
z91ef8c102f104eedfe8d43c4d0bfbbceb447b7f98dc2f1aaddaa68f6d1672884007d8d042912fb
z8eee2e865814abd98b3765e4eff370fb87d9d508026d3d5b228c5170906497f0c928ded0e4de1d
z50f7e44bb39323cb01e6ee3a5e046dbe5688eeab3d906befe2d9e3e76e9e2ed76d490c9e4d494f
z59c1e1407044bdd018126e5af62e85aba6301778162116f8e6e2a4dff10d9d1ecfc6186b9c6a1a
z3ecbe10b7cad8b3f11a4c97d761bf5d643ba558ff7e24c1f73d618878574e87f802230332e4b99
z9b7f61bd5b9ba1b55169c2e32e0d424b41fda5336bbbbb7662e6a03350ee890ad205f379d4fe2e
zdfaf3b047bee74220742666a7874d45a1879e6d71ae1729251f3b1e3b60ee535998e6ff3dccceb
z51488749281d27e667f5e958678a17543cabdef1ef14f1dea63bb18d1a6ff9bd5838a3c75ebf69
z474a167765103d1f54028fff0de69d55560463a373eb5eb532aa2f813d1da9a248ef3bc831475f
z377d155e1cf142bf918ed9a69988261df68f499a304b9a419d35199c3b13364e5f8bc2da25f584
z2a5bad06dec43dbd7296f1e118ed60a584a91c615c36dcdcf834a37b54a3af59ca12ebb754853e
z97a09d758490b002c34e5a765c0e128c5c6d747c5a0547ef83025f8f81b07d61a9347cb89d0972
z170a8acfaadd1c7e262471743991ea6833948fab1cfcf5d465fd4a6821f58c22be2f5ceb9bbe57
zdf544b5e837f1f2e113c688d27c1e41c49120b7f9fb5738641530f7be2c5231177d4b87eeb8208
z0cffcd213ddf472cc96b4d9ece1c1e9f1e4ed1f79c8746861ca8b20afd4f07a67b63adac9e965f
z9141a3a723852dbe319ee50929b7398c8ad3af3f678cdb17b4f4dc673a2eeee8277b8c2e46fd0a
z75af5c1f8af3966424ea0a235074bc4dccbf87c4d6af37446f215a4ab158a7f2d99eca25df412a
zb60100cd742abeec69fdd9683baa0d3f7e04d3ece804205afee739b1d6e1be8c634f0d046d3442
z74d365460bb18343604cf0ae5b2f3e4bd9d7dd502bd195c3cc0bf1bdcac24a5bb9edbc21ec2e01
z080930117784058ad30352f3531ac795e7228e945608f1ad3aedbe361a8511806eab2eed924355
ze3c827b680661840529e090c9c6b2e4d896ae5dcf42b331722cbd8b1f40390518c71f7ef32c453
z6e12ff087777b2c6f403380b02502d1609d54dcc93578945b5ea36249d7b4d92f3c2f859a7869f
z3dac24f7389a0becd615b32290888e5d4dbb8b35dd7b4ef4e60dc372d4ebf4bba7f7b534dbb799
zc8f6e867e92215e66c70c3fa3fdde5f1f5e95ef4cff86a189bae5ffe8e231f1e72dbe7cf507d3f
z698e0dd82f45f5d097e073ffed2bbec89d92a3c26fc4dbebace7cca6e3be077262c411af5c8702
z78ce5dbbed60c0127448e9379e2464c7ec3401414e0ece75431326d82a4fb8eb39be6d699298dc
z35fb86ae1dddcfb3d88a7fcead80206837d5a68a1b906b9d075f68c73ccf9f66071e3c5ed54345
z337752d999ef77e1ec399d60870e851b196aa036e7dc171084d6cb26b63df8ffdebe9cef4f85bd
z02e3de8ae23b8df7d62ba02d2485ddd2931f3e0888da326a3c184c364d30ae1f4753e08693fa87
z52eac98647bf485abe06f4167e3fc0989746769cefc2245a24c6335f660a7c59f7b1b570853aea
z9feeb7c830d93877e7a85a9d7a6cf185ae5d87dbff7998ca735e7229464c314409b2deb1692aeb
z8bb78554b274d31a68217f17e54980910b50e19cb3d444bd517d83f9505f34c751424005f43740
zfd248ccb11e5454eee59e7108224364deb558df6a3af7316c47b7797a27b7de4e73fe0c4901775
z28f74a2d6c78b24b602f3f9b6b39442dd0c51f9a5b7f20bf22a5491611149d0ec3547712309934
zaeadad6f4d30cda607ea35ae6fc9aa8111386ddac581755e57567bd14fa8979ba393319b4ff77c
z7fadd73052fa23ee9c527f2152431f242248bd798910723a8e7588d13137d69e8709f3beeb7ced
z2c0a1bbf121907c4cf06c687ba671be288527bb5c3747525c98bb4c5de57316dbb61142c734b35
z94835e6eeee54bf359bcc7890c529a1f52997c82fbf4184feec80fc48d3e79d57614747aee0840
zece5378d03b1c620acfd621a571ebc3f30f74f380e00f5fe4b562ff0bff93e707f84e3c2a5bac7
z9de4fd71dcaa779300bc656f749f6d41779c5c27e25c232a21cc91dc64c4efe380b3d2cb362b75
z9932a98b63b6f9a4bdb093b708040b50b8c1b8c6cd4e6ae4ca28a9d7cd78add3bd531fa01d8cf5
za336e043a4a186d17ee7218a2463c46bdfca7537d07cfd8fd82279a0efbb5f4dd0398634b38883
z9ed4f17388d2a2a70db458c2e54930d5e7c0ce72b6425850864ca961a527153551d09729577c52
ze7ea43645fb3538314a3b52043b7c3580129c3a1eb25c74d8b7e051666a07d0d86765d51b55c97
zcf24ff68f8495d984c925e68ce014a32753d54f7ec09dce5eceddcbe05f21f2fe5999cd29feae1
z9912e2bef9e41deda5370349696cb64015b9194f15aa1d2900b59fdd1a125d18f50304dfeb7293
z4bde09bf2f1774819f869aa2acf48ef4cd4174f05dc617eb581d7aad9395482d5dc8959522df42
z0dc53c758be39da0bf0cc8040f2f73113a39896f908072357924f881a1d82400fdb4944bc86001
za3645e95304d2ebe5b444cf0d146150c9d7d735c28dd16fcb28bb0d96d889634273c8c11832333
zeb67a083f0ce130597f7036c69f65143eaeeb7acbcdc82b209c49158b878bfa7fc33c1db459fe7
zba71c62a7a39516670667fcc351441ca56890da267df167e9f3be3c673994bdaa6a62272a5b832
z75c49e4bc7c21441288b0c58c88f11fc33b522517adae2eb80ecdec897a3a8e6211dd75a0d52d4
z1ccb86467089e09c67fe3f466480d13e37a952bd18e8b0e7fce216752a4daa49c7c3b87b7d7260
z860c161e60374f9c51dc1aa31f57c0d812c64ad3801395ed196a09099c0524c0af697f5e14fa81
zd91a96e1d390a7a448e5f8d9248c17fb7d40863343d42118c36566f9e271478a9f24dd4968b7d1
z1d5999b02df8ae8d73b8aa19ba6fac48a4abdf9458a69df4c0757c4d473bf6d119000186ec2ca3
z715c2fb3129d55327b71e23cb03886ee2ea663beafaee4040a413fd5f30903779a3f8c0d228a19
z982969dddefc3a624d8f305cc1268761d7bcc585a26071d9bf459c34d9468589b437ccd67bcef5
ze87da93e0d404fcfa34252e6628298ce6e33c6ff739327d95076cc4c39c0bc881e074b7881e156
zc780cba3787e7c6043fd13869f95185b9f5feb0aaf58e8588ae4444e59e94a7854624bc3c4b093
z3a38bae39d715982d96030aff7aec834d60e156d047b07ff2a05ce63193243d9aa3838fbf97ed0
zc059c9a4df9cf10915c3bbf10de2a38ca777e8369af77c27554698cdbaa0bfec4007eede80e59d
zf51cac4ad69774dc0d3fc81e7a8e86f255b2c3dcf440945e2e155ae0d686b24b8e8f4b4b33a663
z91de9625e8721f1d4e302854c04adf62a6208c48e8660aaa0fc2b425ef75b7460333575c423eaf
z7c5181fe97f164cf11fcda6def0c59fe420f0a893c36855bfb9fd545359a804a945f4b5ee65f22
zd349608b9a4f2827441d158ee7bd3a3e1492ecd63850b3a202d7a08fba26cd635688fab5533c80
z7ac77b68b20a6f2684aa463e633da12a3fab0b9ea04483e70fc9c6cf6ac119f0c93a57b18982fb
z26a669b06ebbc892343292e46a6659395bb4c16795778469620d183fb6a13528f7cf3daf928841
z6342f7c4bd6df926441e355cd8aea72687cf6e1da47d20193a17b3222220893f4038d1171fe0bb
zf6c857a527122accfe94f378cd3129378f918f827ff87e95740a07811434ad2180e7419ddb4cdd
z091cb83ff2539ec81f8d8ba4aab498baad29b91f6d41b5f3314b16dcfb49edc16c63e91db2e865
zc3ef8481fa9d3b5d7fbc5270827b6510535aba4a2131ce739109118b5cde295f80a6fe5c09126e
za9c7edc7875c60f73c94c2ad8f9f5b27426a46924a40fbd94cd4055dfb80888fdd9702bccfeca2
z2d3becfc028104471497aba2f5044bcda53d8bb9f36ef9d8af4d803cac560afe93c95421dd27c6
z3e287dab1fd161abd777f49870d96310869ff86d0f9669dcb82b515c4e4ee8485677389e5cd540
z1bb47b31dc1148d24daa326f28f81cf5f419152982666c325a27912069ae257fad587c5773667d
z5b0fee38f22bac9e40af080b29e707d88e34c19e4296c1c2bbdac43594fe633886032ac201911a
z4bfffcc7fb594b235917b23c66f8b73b3d0b10e1dec20e7220ae149bd31586e0597acc1cff98b4
zb2cf658ad76d7a05ac058ed2677b132acf643d289652700c1e44711224a74e3485b6bc51d51416
z23a18c3922945b08db76482f4a9fb932f730dc46f3012ef7fe1bb5bb2dc5ae4c12fe786b7394ce
zcc0378ae135e6c53149f12d89c58405c9670e422ba8232303550a38ba9f2984ac06ba1857b6753
zb525c0fa5daec971f5450aa7cf4d9b329ef2f0c77e22a21ac25c2a882228f3ca56922740c22839
z4b473edd902cd597e831136f41b8488623c4c6731be9e6cb684868d3cc3f99f6ec81d3aefdf779
zf57326029d775bb29dff05f6ca91406b4fc6a0bf83fce870da354f35c2c976e6d2cb4485728d8e
z790dabd9fc8ea880fc0b920a6ebcda9511e16d18be9d2a38f1491aafb86041b0b3b3dda3fd258f
z8524d5ffa35ef3b96cf3e5a26dbb2581545995dd1ca432f32538f1baffdbd718de180256cb56c7
zd5813ea4cbca77954c4d1d6a7894404d36b618238146d7b5929fa7cdb9b94a1afb50cd4eb44f5e
z6e37fe01c8c16ce534df279911da8e6d75aec6ad240f9bb4bcbbbfc1624d6fa18ccdb1c8f6d001
z2efb4f281e166d52b492bd07514820f24b38e9975cc06e7a01c43cd2d5158c3a607241207cf7dc
z6cea2f897de34c4b602490ddc2ff1beda9023c10f628cf983baceb2492b7eb8c057bd996941141
zc152114045fbec891132e27568396f6da63e1ffa6da9675dcf7c14bf7a4049e95c3b55d01759da
zd98253938b84b0a993eac138dbfc8951bb0ae338a108134813613581ff4b01ff828068c95f9a35
z6eb24cc42ed461312377231f82a1e2cda344ede3bf87f2dfa7cb037c01674c54372ac4e232e9f3
z9dbba69bcf6431c569259d01acd49f0f7968cc20419256a010b3357ab0bbd20a2c5178e4c8c3f5
z7096b2c2657c9215d362792a19836b7e2dba1d29d78da78faac29d1a62feb210384a9400efc8c4
z47829b076baf76c8ace3ffac300215c13b4f3ea723c0470a93030e4d1ed1ca8a3987c28cb45a15
z714efaa03fba457718d1709e25890ff9dee0cdfb58944f02295ce4f6f4d6e9e3dc6d1dd950e8b8
z01e927e8de43473eabe25a713f7fbdbffaf0699a8203c134249f62deac88b77c750ce6d99d23e2
za14c1d36b701517a105810ea1bca8141afba13d60598c55b68510ed1533ea45b85e11cab2efc33
z62a638e1a4375c2425950e6d46bf9041bf038fd1753d0a4e643f97ca2162b4fd781d92039a2997
zfafce191c443228e1916685e9131a21feafb13edb98b3b1a05472bf75359e3920d5774b69f6d7c
z6fb015fd7af4200a9ce251aed361a6c3abf83762fa02004f55a56353bf11e47a7f7bde7c141036
ze55b6dedb131cf87bdc8797c783b83e6fbba8f93462a3b1952731638227c9380eadba607e65222
z22323c9c3e831b08029adc318507f2588bd5ea94c00b9027370b5e304f18a2ddbcd1f640cdf1c8
z1e7c8315fea8047787d8ebab14cc64468f1277ba6c48f269ca83d6b80df70c844ddca7236124a6
z7702650437b5d7c6b0d14168d3fa225d7aa16da089ebcc12e4b618222a078aa8aebc3ed00bf9ed
z5407074bcfa76d20ad5f932d1e6aec9dba5a05913ddc8c7521e97e052cbb45febfd2c4099b442f
z462eb64c648bb1dd6d9826ced6d0ba606ea29f07826134a0abee65095300ca6009550587c86cf8
zf13d158aefd1d4b157ec97459842c7da28c116225ae57da702dfffef2b66f20c31a338484c16da
za5dbd5bf8fcf9da0f8f1442e2eef42a0d62756a9d362c20659781071fbdd211318a92840b14ab3
zb722e25cb57712f4372600b94f2f89adc9e4c6b9d2ed9672d254656031313288f63b350ec7c33f
z73185fe79a8cf7e88300954b46c255f154fb9e13e2f59473de47d904d69f49d72a4a75e4703328
zbab8062ed929bf3fee57c8251aaed0c1c34d73a475f1ac6b1d773fcc1d37e280c6a4cc7ae2d257
zcec035693748324a5501564912d6c0ab6b6e2b998a700ada283cc5d313fa6d38fd3b9c3a2a107d
z2c91f4c4b12600313fba641eaff6c56deffe47f7484edc73791e36941952538c9e0f045c23b8ec
z8080203c77f3ea1acc0adf204c1c76050b499f274f709348a2fa66df27f3c52a4a1a562332e763
z7ce83fd5a1d663a8c77cc745aaf8b2f66ff4da11c34c1af94acea3e4039e2630c742e79e60a5e8
za406dd69e1cccbd98e198b831bbd32d42636119e1d8229698e38e81591e6ce2d8880b2e7957fa6
zfe135a770bb1b28f51f2ea90e38fa91f52ced8f2c1b1c9ebf0f8cf84c242cfaf95eeddf928cd2d
z8859dcf597daae5698170a21f56465f4783023d6ddfbac35df9525e67fae528738564d8b0f2f18
zc24b80c4913119e97c0c968f48c84f4c26059534d1b155d87a29d0de70f0a5b9a99ea4640b3ab2
ze95c122929aa3b778dfaf93b6ac46660343bcd66f941d97792948eea3d94dcd4019881aa1876a0
z399705ab2bf8ae53f9a89fec09c2aba10638db54e195ba4a3a8cc4d327b9023dcf2a2a2c8e0b67
z9570359dee583de055b1c361d3704a28bb757d3155bc5210dbaca68db78074bc959cc26e530a58
z4ffee77dda47128b7f9974669a41984ef2fd79ffe60ae4a5eb8d9ead775eec66c75690be9f85ff
zc7385ca94ba75deabb0ecb724c6ec50431d919de92e889004a5e962e83fb675e61ef48821bcfcb
z3c0e1c07c00ea5f23bdc4352ce4fb26674993a63d991b8ad77685dca0208d35747409e2b2e241e
zdc3932a91c5ff01721e4be871393735d692912e5b9afbbb59a1d5ca383f23d7dbd9b8a18bc3acc
z3b523f39acae48e1bd98d0945bb9aa95d11381b9d768d73f1d387d8a98edac478ecad498043414
z6cb7bc37d3269d7c62703e311e2cd48debd7b00dae385f04c119eac54f9574fadcc0a57d601b7d
zf57db5ca14489e08ceaf0ca9414a5990ccc850022b072b2c144d84fb5a178314cd9208a1997e38
z1f3ef38014e394c3875a36f7b0b87449f05c820a51cf880cebf839ee09cf1f09a573b9f82adda5
z7cdcd752ecc07b3c215d3ca5b10c730261bd193fea18832dc37b235bdff9fbbab059f27f90ecd5
z1e7f8deda5b3a9ba7c1c63a88e7a45b4aee4fc4e5cb544a0bfedceff2175207bdf3967f9258d6d
z168360a7dac2f0b04602165b1136a394e5037636d2efe75abdf3dfb6508d13cec932276bf8a692
z822620d3b4d94ed9dec45f6dd65185be22e7e1b373beb4a2e2ce3cbd27d3ad66c1499901a58a70
ze1058346a86cbb3d72e68139f82bc4827fd47d0573cdc50f352708b97fe67c0f03fb4e56f794ba
z257e2bf0adad4737f4782517dc61d1459845172184fdfcf05a977fdba3282c55930526b6684d2f
zf09ebe032a2dda27e4c7a87cc4841ebbb6a81531b50e78dd2d46105d96ed1e5ada4301097c519c
zcebd8afb4c505324deaa9f0ce8205b1de5df8eb807a876841ba63089d086f17632106e3ef6d52a
zadb96f3c29423421249a77824f7ae62732a23e8351b55326bef34f1fdf554023bfdea1459760ca
zf341b9d0067c907d16086e5371dfd303806bd90e66d87c2bd6a4ed5c4c63c761fa0b9d7dee1539
z6ff2fffa2eac608632222e621a88f389d347a14cc9cea89e0aad6a9e143a3bc2e750452ca3372a
z499274d6dea5ef6729c4ffd1d771742b454f28b9ca0ab864cb3eea7662e4becac2a6347bf7f9c2
zfef3ed76ce70f6dee648e6752079d74064ee6c1456f32b404a930e6b1ba4bf1ed10256146ad87f
zd9f3a56709fbbed3423e0a434ab4bce3f47c07683f6fcd8189cb18710183d04595658f4efdfd2e
zb246b884103d92898f34c4a80161b0dc30a808454616c3524cd530c81e4da3a17ed36dd8f0d849
zc41c71a1cd540572508b25e0dfba3b74a3d7fc0705f9a7c612679aa17589802e9cc440dd7f744b
z0ac366acd8b82e64ea1f8c186e2353506561047f7d4973445f703d046cdcf923615a2049d8bef3
z67bfff4788ac6b9a1eb33b0e94467622c77fed44e22768cec7e02a7e8e7f1c64a4ca46837d84ff
ze729ea38c0141768fa286575234db6cb762e7b936fe80fc5e5c10a04ac3022d651c629787862fb
z17280116aeffe18a69a543bd2ce427dce219c3488ce04df5c7bb76a9553d111a44e4c77838a0f8
z3eeec4a815e12846c5aeca608a9620bbe36d2ed9329c81dfc5d9fa8a4ea2a8f49a4dec17b0edbd
z61b4c302cdec599c43b761fe701f5f2c96502d5dd9aa8321a84a42a682e9ad82255dcd8ddfd06b
z02896f55b77c56cea4799677367decc120efe12dc35f39ae7743cbd7bfc522b2b35a3b07977504
z964bf440a6b69ea4f33dd3f33a72628544142c598c7195229d044fe3d6a4653c9b8000ae4a69d8
z8d8b23591d99f9b999c312f3d6f3ca449cdb697ee02dad9fe19eaf622733d7fd52461c9a0c810b
z10ec6bf022e77a09e5c5b2802b9636e53215bb0afe27f4d0875ad2f649f62aab35de30c3050131
zadf3eb6192ad6d0015d9aea9d3c53d1e02839e0ac030573c9bf93c481ed659910a23d6faf30255
z68efcb3fca6656765bd9417f470ab2383c8fa54da6683d58fd66e0ac289b12a987c1db7e4dc01a
z9d0abaf17310fdf4f74ba6d313679f61912e7c2395f17310838fa67ac581a5780f51044d26c602
z22b44f7597346cf82d55705cdd04d5c878ae337bd1acffbb43ca2deb4e8fde7cab03c3603eb210
zb3e8db554559cbcca0036db52b71bd40d280b19e27d6bf68081a96346f9c832828f939239a9234
zc6690fc3e37af6f1395c15255b3e22c97b4727e3628c0cfe05be2b2d6dd25d12aebd5a718a3ccb
z139d1d3ec62b0b1ceb68151d0fa196bec665146eb75446c88ba4fc019c046883d6d283d065617d
z13e1fd2c6efa57369fc31e311e598e52a41fe93bfff0a00130da40ea0c29819017b1adefb8ade1
z9c7ee33baf3c3802c39a8f6eef4ac5cb9ce250a308ef36ea530fa2b4a6b183a7dc043d76986d07
zf077ff0831f77d5c231642743ce4abfd3b32149a2c2034a020354f113c3c8827856e34f14e2d18
z0cfb0e6229f807336351b314c655559f0174df6b5135a0b768d1f400d8da98f3c3db6ca56e29b7
z2361b6b650fb3a2073496013ee16a45140e82f205d7664c9b3b92b1485026c17cb5ad5df073994
z58c6bec7fb65fb067d749d43ff3f82b7d04f08dbf49063df2bde76efe442f302200c89e2c1a731
z0a5898072860e92721be7590085c7da46363fb519bba422bcdd39f6bf11ea46a80e60e3e5d5904
z1d84f845d2e1edb1cccce1245b55ff2a37586a3977b3bb9a5c5ff3f272e30266b66cfbd99128e4
z72c5db935c07c8aa29a65429ebeb499cdd2233747bb7370236bb20c56b7f82d611c4382498a61a
z83f100a53b9e0e4d05262378731d1527ffd1fed71af1d855b4f5dfeaf5a13faafba4444c21e969
z4cf4ce196afa70c757c2aac169e4a715273c79db0012534241524a44950f65d265ab0d5e4c6f0e
zc38a19c7352bb6c37621924c4efb1b68a5cdc9ac49ee370032535f508110991ec1c0428acb823b
zb8bb5d87c65b39bfa670248d1cfd5157ea4fcb478de50ec4765e545b14cc033bd1ca464171ebb7
z35384abcc7bf96a95f9a446ec8df70371bf087f92bc1706e374551aec5919ff1ce2ddc912e2021
z5c4d2bbc54a7e034392425e19d87687fb604994b042721bc0c533433fe76b3a4621ea17ad32b98
z21779cd34319b38635011fc0707e9c818b1f2991df88199e5fe1ef91d80d4ff7e2edb5cf262776
z181094edb79111fd4ed430f3c7ee68d72e4fa79bc027c9625d59eb83cdbca5b27147e857597b7a
zf48afc1c26de1e06fee0a3e29d0bb87133e85f5bcda551cef78fff9a00f72db862e62f29e81449
z0989b8217384092c967287c767b57e817e04ece501dfd20b9fb5c5899a3fb792b7b46f451cb44a
za6c69882f37be523b39e0d2991592dbf0a9af8a4259e50e3c4941500d412d95c8b29a8f29fa793
ze832cc768fd912c0026486974e04f753a4e1df2428c16d0a5f27f21d7d2192a643ca632a58bab1
z8ea393f5ff870c08b31e4a8ebaddbb5994af5790f5f224da4e11d5d874814421d48f02ec88884e
z5b836841fae92751ac513d9c7fc3630486171ae472c9c72d43cdb0a83d425bfb6643979b58f64f
z11499afaf36cf9edfd641274c9ae648c29bf3742cbe1ff8995c9de401d7208dbc8f98fe24c6b12
z4fecd7e1b30ab03cad40e59ad0b5786b22f71ba237de8ab9138167bcb7f2690df4b47daa12ac8c
zfac185ecbdd7485a673280a6ff88ec9da21087f5116041fce3cbdeaabb28feb9d6f4038c5d5a6c
zb7b7fe2bd675624f73f8054c277872ec9d8b31631862309522d6516610a2031ef0067c6ccfc869
z94962f1ba8ed43afecb85caec80982d4197fd4c3dd743986cb3d324d8228bc620b3966ffb45993
z4c4e3d3b6ea97df5ca96fe0016193918045871b6a219d3f141ddab3a05b893375920d295a7b4cb
z5ee2135712e9fe04db7f3ac1b207c8a0dfaf9fa56edf6b300eb890cdadae05eb996527c0d30849
z1cb09060b7c7f5704977f72492e668fc7e9fbd9784a47f65f9a3f3e0368b72324d4230dd07ec8a
z5f6ba93543e8e4d7411124ee7fc9e8592de852877d65df78d712da282a823388e818e04c5bea97
zf5823f5eaa64404b1a4f4838f8661df0a4edcfcd85d7a07093386b4a68550974b64611359217cf
z7f3142b806ebdeabcf62a4921fbe574414aa4eeedcce7abc0bbffe0357db97519e90cc1b21bfcf
zf04a245b0f460f6a237512b285ee44b7cc182aa57a4530122fe55630338655386ca1cd969dcfee
ze8451f94de9dd5171528eab2ba884be755878793ccf2d6246d1360fb49984fc1342b8f5060783d
z433d023c89d09bac4dfdff64333d803519d8a63a2086981b50d53425a31c961b44345ad6b7db42
z7c92c6f428808ed2a1c273af309eebc1a86f41f07264a8cfc671506fb9985714187fc2066c9115
zbcd0513ae9204c2185c525e942e2fce5588acf29c7449f8393e579ccced244b182f39b419ba2c2
z78879d791b9e4fce9011cf914b26dd1ed271dad2696d00b51783be079670a0c13e56029ea4196d
z065a4ac55686fcd123776308d138dd909ca048bf6a804c5825be494c51f6216123c0e7499e26e0
z44502d164d655195a7de209b9f6e10f2b57a7b0a690e8ef58dca100617bc2472ad7971bcc78b83
z5cf014a5c94c1d2ca9210613ebf32493e585a0a55b32a81d988d06b5c7cfbe844bf4d667f450b5
z507f097eb10b00e913ce25277790f55ac2530fe69235c50321170df1957ad0bb27dceab88eb46f
zb8b4eca318bb86fcafb13a28e114f0b536d76989f4e4edab3db92e24306f69af90bc34c63f9832
zbdfd87618aea2327ea78878f6f1d42a1da1ccdfdd4803323ae09f64774f82fb140c828aa16d137
zbc5f8cadfb1de6b3cb19daa01c9bec8bb56f41a696af6f2130b19b6ae9a49a3685d023b0174836
zd0e62b23fdff99441b3a50b0da8e0f7254935350af25e5f97df75b3bb3135543195f97186a4c71
z64925d326de2373beb696e47547ef9e29cdabdf64a837879f27ad61c3ce35edb8eddaa36a6a167
z657156a3dfbe9663080477ab81b523bb98869b3b4e5af66ce66e1c755438a63cc11c62918ac51c
z5b57962a700e0055485ba3e0c06509322592380fd2255ba11ec250b914d628a1d8cfaab23bee85
z9d7dd53f658d907c62b88ac532fffd5d6b42df2b4738365c55b98a10b4ecc7cbe15d8cf895a3c2
z265f82363e4cdcb81a49ec9a3b447bed6aaf9e0f03d1f3bbe3ad320bfe12e187f08127778627b7
z2397fddcd42d667e381cfe6b4b553db6377a9c27459b300a5706a734babcf707d629556955113f
z457d8daac078007fe98ace2ff3019465d03d2e8431349f00ecfa72319ff4bf71bfed08d2f6862a
zadb28d480e3db4a1ebfbea1027aad27006acf6c978633a9b5b76a58b30c5774d8ac12d17804581
zcaed98c4e6ac9ad44fb43380a58f8830cd880bf1bf8fba9a631193fd28fe7e37ff5e6e097fe286
z1f13521e62958f4155a14314b83515817018b2b607252cc9e864827f32d5344dc723dcade5dead
zf3a5261e82e70b86e50abf5fb12165ef9e1939be6f5884319ee236bbe8d199648c66c8945ac22c
zc50dab5adc2189b0f651a08ddca28a80411171c26d92fdbbdfe85f360b002c91d0bd05909d8199
zfab20bb2524ffa1cffcf13ec69bbf6fe3d1bd58c837a74b2bc5909af9eaa07103df2ce6831534d
z80de4d7a33e0b5e8bed191ba8463a0099810d291e0da1e60a7b55543b6851d00232134c14e8c96
zd5d63b964f68c62a355897ffe2a7322df2bd1489083a9fe4ab7ae61aecb0bc20788c27cbd31cd4
zed9c76bf5155db6a454c26a3b21906f2704d1cc61ca25d1deddd074c06e96328ea7cb0b81a8465
z488f8747761a0598347bddc4833c64a2f77164a8da361f7621fa3f5ec72ece185a2211d30bb489
zdbb55bc87337e033578eedf77898761a73dc9368cb1c4855a15f7e276c38117592566b7abc46c0
z89aaca589770f93049171d033171803f2fb44f1d4e7276f3b2b659bdfa47391a09794ced7f3687
z31830b3ac4e1effdf41ab1c997906766977104a247559229532df81c44aff6e1ac8e28721713e9
za2dd2fbb8b33c66e649e40ab5a8fba6b879ffcccfe31a2bde06bacdf589a65e053613e5b26f1fc
z6b9a16711fd8cc00c1beeb4044e250c514e9534de8ebc53a8afed86c2678cac16769c1447c247c
z20eeb2a988f0161aab7c976a1cb67b9daf072dbe6e01399e825a942ade9ceea462098de5aa2bd6
z59a16bd278be16f06cc5dde5bbadc599f717f94a1318c979d46e670766dbf331564e2139dd4e7a
z02e1ad106418c5c52a5b54bdb2a913876f5057dacbd15bd8dab2462e95ca3cf94388932592accd
z926373fdca46e27c8cb790c0fd4eea769c99edc6339ab866c4644025f69535c8d61159448730ac
zc4b0fa6d4989a710cc2e14d722e55bfa3ada5afc06fed4f3e78087d42dc06a4b7a29bbcf10e7e6
ze89b22fa8cb5ab325c502f0576f7e58c588d1a7a046be1e4a851bba21a1bf33987783330b076e8
zc9c0d3186766acc0182e90c39954f6351106085e1e3f742cd940ad03af211fb5b04c7b0d210447
zf52e1f56432352677d36a465da363bd598ef0097a20ba1f3ded0d0d6f1cd5847264665d3375fd7
zd2c7681090e3332fcc527ca0bea53bf8006f299684f3fcb55967d0afdcace989711fe1be0aed82
z10f37ac80da59a7e0016147aeea6576e781bc21b9117e4272baa46c1d074cc66e4d2d3a72374ff
zadd4215f8a231711843f3cde4f49bda19a535c31d4156a7d48f1107d283b9da0a8db18a3c4bd05
z43031fdb3b5a091ae1ba77ea33101b501b267978385874a23074af45935aa8fabfc6252e822056
z871173c3183c62c5790076db00eb9c395e3f4f8bfab9f733ae1d9d130bdb68ba9ea724ec24d94d
z0f13e1151c3f4ce3b197ca911d875fa9008fa5f29c51984f922f02052c4ad19e315350cc7b6597
zd40ba315a5afcafb658562fdd1b30dae232dd5d318e92832d5df402843cadd10e20510c20b1c66
z0dcc93b43b28e7e23bae96a5136c159811aed5c8453addfa5f29b0a028f6dc25ee489584a66023
z7faf8548221d7adddfd8296e68e0b6243fef68e27dae0673ade549f6ffe53dae1222d1de648329
ze40ad9328610e3c74c215af6e17458d509f16b97c82bda9aa22b95f70e43154963204799ad739c
zd85fe163727822ff086bcd01a93614c48fe98b98a0ca7ff9c9607fa4996bb5f519abc7e0154d2b
zb91a1685a8eea7d9c9a64b05fca584ecaa2b7ead4cb4f87b8b9c2b3d66e72cf4e844df6e829a8e
zd9bed64eb2351c8b0674734a16f78b58195804e1b2d50803de16306e98268e7d87bacf9653495f
z1a5c843838f253c5a912f48fbe095f614213ab83524038132d10c3e3a89215a5ba6ae963ae7770
zbe3f1216c6ea140eccfccc1bcc291748df8774b17561655c52b0077c32380e96bb948892b17879
zf0ea6ff6de66a09ad4c2392e4bffcb49de264fc076b107a6ec8706af48d3da845f4e188430b75a
z4aae3cb41da782dd41151390ec1c26c4e14ca29f986bde1b416a8987ce1d711a17eda28e2c4e98
z9c0d7011cc47616b335c29b6d58eaca859a4c039687e7eda4050867caa6568215e6c9e80b5cc47
z4eaa3b144ffbe1b816963a2f022b56bcd3c8c6dad0855f0872dc2e06c5cf5f830756ade9a1ce4a
z909be121d1ef570c6b94dd86360cb41b92bd965e4aeb8d2e1205917ca6b7156d7ed0ff50ac8c27
z31d40e6e598e91a79f4b3ec7f428940c4fd6db04e1e8f3aa52f7b3c83ad99ea667c660162b1233
zf750fc5753ae1af343da9c008df80d6cfee74cdcb60aaa652444741a94e1af7264cbd49b8b6dce
z75b32a2bfada524d43e6e1c436a9bd49f13136df8e30b1e7e755e28020412a1fef009af50773d5
z507518b100803ac2402cda696591b5d09b055996e60442e83117a7a3d375e1fdf8fb7752b953fa
z8400a8aa2fcecbdb93b271f0af0d006eede12e872edd5884d6f6026c1c205d50c4495c33c70fa2
z979025cd530ca49921b819a1dc4024d883e97e573d11e9d4a1204f8e12ce484f7e70afbf6a1f3f
z71761d72e5279c30abfacf5e4105f30a506217986676362eb4a2e629257645bc52809ba18eeb4b
z55293f9ff9528251775a4cb35833945f4bc1353dd619c2cf2e0d47dfbd882484ea733ca0fe9dff
z64dfbd05613e40e862012af6bf340c7530344ce6edca767476b4eabd8708eb9019f0c8fc60b4f1
zb218ba7049409fb58524681c07399114bde4cc5528aab006eef397aef119fcf84f78ebdb750a5f
z169ce2d195aad9e1c187a5f631a99320629c9869c6bf66989dd69abcd54d43bb076c00fa940d09
z59c0f6b3d81c3de5efa977f0610d3987d1733f6a6f36d0c21aa96d1adb2edeea2be32907d9dffa
z5a2510a2f66cbb9a74549653d1b53dd40b8eb5a49ef97d836c87c2acbebbb3f85713cccf60f483
z7302de293ef3579641340d9afbe1fda5a40448ea40c278a4d3ea2d067a10372331134da9a664b1
z385d6b4b133b6a651e25a68d380389b24e57d65c7e6b94d3628777bb124af07c7bf16fbe0dcb71
z5251a212c84c9b4ae88af5e532975bae982def428014f372c8e08b80f7c051086382d01f1d0391
z56baa3befddae5137de049475689f365a9585938401bbc69c97dad27dd7c5f78b9a5455215df16
z294481ffebf4d3f2ff51fd015c2e1838f1f24b973ccce5620fc470bcf272b1a8384b67fee22a8d
ze20944a0f2f9ac0d4f78f03f4cec22bfe281f9d983435258141884491355ee4b5c009ac76491d7
z29b603f22cfb4655bd306f52d1b10b4145fccc880b4a0473e745ca093c0c856488ab69f4786c6e
z802181041bf8865d6010f54587a9b8f8e88b0fc5e9e5ae96fdbe36f40f63f72f741b99ff3d31bd
z3c3379095d070c229dbc7b4b3f3003c797cb2e6f8bf47f25e97c335285941c546cd0ab5e13359b
zcb23fb29a3c17707212794d15ad52b895ed1089817e33af829961b825fa35a4c3d34cdbee1df68
z7244c152c6bd0cb8652a982b7687071f0873b9c3ce9926e7099319e8d8a6121dcd0a8497645d89
z8d3b77f068782ae318cf825c9ef2673fcfacc400cbf0c32494ebfa0c51084ef16384eb12b493b6
z185004e2e7885e7eb368417abdb04d6e69b8c282e3b52ec3bbfa627c659c025f5f2a36f3e0a7fc
z7dca2a728868f195d3a39c83dd87352c076a9e1ca0ab2c19e1221670a8994cbeae5cb77dd7b52e
z6aadd37ca792f74b1607f5cfa05677ece151b498f9b29f4ec2de25e99d937a27a10dc31f89fab5
z1df46cb8fdf95b3268cba6b491c9dd4d49fd15ec0a736c917b561f2cc98fe1b6f479a6ce5f8a4c
zb29ea1830575c608b09be5dfcd575609e8b43db388a8d94d815cd376713fe2b8a8ab624f037b1b
za043f51a009b036bf2e8021dfd8dab2a910876fbf77d31db8588eb2734cc0d002c48dbef6053ab
za80957bb5be3705775c3d048ebbf87587847717b4017eb6b3f8ca740d9634411a68c42af4871cc
z66746ac987ac8c16ca09411990078a2f5b635b944cfc756212d0f7e86469d2980803e5ba8d4abf
zc1cec63928fe0f24c34dac7380c1181c72ee7e3bce64e24b634ea48dd7601b727293b48c2604e5
za7dc79cf5d951fcf90569b766861348173185c3de4577055056b1ebf090af6ac7a8037a45466e5
z92929b9c655228303fcb104e80947bd893c51fbb4ad6b252b24286327bfd3e146937b4ed6f8aca
z180d73d0283ea12944c43e8199a0d7e564eab3214f791598cfcb8faa7bc6790ea019d03c0e3ca7
z7056fff5d5e9531134677e073c169ae28b937b223d3c4d1531476825730ea663131ce4c960e5cc
zeb32da0d2cc25dcf807bb0ea9919a3d8cfbb6b4885b2201c0bbd9bdc8f00410b62e364699a3fae
z4cd028951da506634d7f1976bea4d88a81528d4793365838534782dd86fc80764c4dbc70f6a9fb
zdee079a01cfb60647f077e93321b76ee7aff9fbe6d2e9c088ae337fac7f87fb39756cda032b27e
z1d41309d6a9b2feaf2acfbdfe93182723b53b9cac3574fdf15a1aebd3000037ac618c5a720582e
zc529188ff72a03fcdfd869a8faef843440ee97dfa30bdf50bca56dbaedf337a530300085fd773c
za1da5dc8612d423f299f78797665bf9ef13452cb90820901eeca25d3bc17f84db1ea7935a0e408
z4b4e18820640c7b631ab120bb4030fb436bfe88f7802815b8c4377760e864ffafedc5d32c000af
z01d7678889c554d9344798f0e53689374ced225a3b6d29bc60b4410df05c1228e6b60c240af538
ze135b4fc2bad91e85dbc7ede4d6a4d5f1f197176354e0995e860a346246ed90626c2b133362f6d
zd9f1cadf0450eb86d1a4b9c7bd43907e8c19b21c84bcf52cbc3dafa393a287e76faf800b5b8968
zadc37818b1bd5a6e94a6c36c8e72f3b9d464148f6aa9be60d454832a607e1cf03f62fa78553ebf
z1a8fa88f5f51c3926292ee778b06dfcaf43ad64c92d8929b9e5aca4a589caac853512c6c36b2b9
z65067d769e30823f2222bb7f821dfd58bd355ebef419dfa63a9e601c33dc4cb65d566def988fd7
z0593472afcf867fb59a92f6f51744f7372d1dc26cb91626df0bc4143aee35a60be5bed52d53fb3
zb21dad2d3891162de9a3226ac2ddecb638ab64b34fdfcfceceae36661f6ddd97fa39f6ab438fc5
z0f3405a899de215618477003ae00e29028e6c14555804d8745e060fa769c1f8dfe0bf1edc8cd41
z121456ae8c53e3b4b940a1b6e9b1238ec44ddbceed44363a043be5359f989296cad3feb411e389
zed43b490275ce9f1baf7bd0879ffa9aeec3bb388a948ead97afa69782ee53e772a2d12c770c016
zf3e676c698663775a11f9f446ce62e8c56807b1fe9fe32bbcf2bc17b988785c6f02e9a381896ef
z420f4e7ac88beed6ab16d51009649f908c8d3800bb93353969d43e8f9097be401bec02126a1196
z97a616b7acb0b4a6f96d0fe11ea83529a4ad3c2f1b455e87558caf0255059fbf720821bf9df8f2
z81907cdf09b1138cc97f26580ae98b2d6d06a3136ad1078c8b5e552d354daf6f0a070ecddf3d4f
z139d977f30a23b630fb69831e9933cab04f09144ac8b7c1460bff3a751a2a799c43503c4b58fe8
z32b6f1c79f5582ef3f2323b1041236e6ee54d472a2cded8c4d542bd3a72fc944f3692edb1179d1
zeb16dde1920dbff0be38e170d174e3c143016d7017c8e858dd82be6686d4a85ac85a14ecbc80a3
z3fa282b9a7360d5e37636be8265fa01fc72c3063de44f58048efc49d6d01c2917c2a78497c82d6
ze0d27962b06118448e35db7723981605f62b643250c1fdd1c3226fe22bcc0c6823647cf71165ea
z472836ec1cf31397be87b53b44033c87fdb77376db086d2c93cd380e20af8556ebfe929f84e056
ze61d06198bcbde020a7f186d7ca233789f9364dc47194fa673c9aa76a340030dab85056b92ac8c
z570de919c0ff569998dd96e8808f5272a82afa9622cce5335e1c9bd677543fd33f67f36b602dc0
z5a34f353213a1021d4b43eff0caab120416216620dd29d9fca5832a854468b1b757cff10d8e1a8
zef552d81cfa814de96486f7ed987af14584dd7652d07ead3d8d4bacc9ceadda6987543dbd00722
z09a25ccc0bbc389216d1363f1ec14ab857ebe2177cca202c7fd1b12220d2c94e0a2c57951da636
zfb529d83dc543c379a17be5cfb14d38e59ec930a6247b0803bd34a501e731bc7ece6dc0d476aee
zc7dd89d221189236544b8bce84f602c639fe9c58ab1db8e97f7f7995004a67ba491199645e1f3a
z65ba050f0aa8b83478bc57d3b0b135b781df382f848d8581c5fabf2c3c3cbf8a73fa215aa35b80
zed40e8c715db2da83805f9721df88839c1bf36f454db6f75b6998dc886aff28abe6d370f95e797
z3fb467bca09584ca5859515e3026a6f6c649a939a506d3b615e886223a75741119c4b1dc2ea8d9
zd92b97c86f0cf89c6176507217cfeee01f2b7ff2ecfb394625b49fd30d449473dc1326298defe2
zfc651efcee20077ad3ff3cc0f6f06fb91705878b0a6852bea33737455ab13a55f76bc999c0d27a
zb39a52ae2dcc1ee801a6b1b9a8c6d23cbb855750d004e5111d322e634b40ee0e37507460229ddb
z5cea3c0c02af25ed4c6683f1c6ca4ba69b3e734227fc196297e95576333420005fa2b466876bb9
z206342cd8b53c407417b1fa719cee2b377ad4165d88819320603d558684694832372a91157aee8
zcfd4136f940a8ee93c97d6921b27d38854f3b4b3801f26bd7bb0af88bcf179abee1b46bfd7fca3
za8fe3b0ea7854f48a83b04da0155cdcb877a0044de4eaf62136d5ba6012b011c06e4a0f66f5bb3
z798e5cec329b2ea5fc835a9d4d6326cb67c273eb0c444971bb4f3c0dbc382f2fe3c4f89d1c30e8
z2be3cac61aaf0959ecb061a80080201f8873a43a0b7244ba2a5288c9567faf9a2ec55184153efa
z8a4b934fd8a68ae07f9c8d3d821cbe1d573e4f195d75e8ec097c2bae92ca927a16a8376f09371f
z9daff6dca207b29620d56b9fde0e41cf18700c7979f4c5cd530f869100e3aa063a78c40b34c8a3
z6117dd4128059b05e196de3c3567acd46bc73fce3a0e1dea06396bae797df5673f29ce672992f2
zff126bbedcb32daa8ea0795952b915f84b48c47ca4b72926adcaa7baf68205e46eb16806184809
zc8926a9a26aa1bfd7fc38c0fa4b427dc49998ef756e2198e967db8bec5d261d81cbaeb9598da66
z273560dba1b82d747df32d56f87ab724f5bdfac832c618a91fa0c4d8148f598c01a9c1a40a46ae
z98506e987f3505e0499a0d407ed2e71f1d59d968701d84e30828ce1f0fae2ab69dcec38e0302c8
z1b126111011febb2d583e2245446bf451afe34a0168a82e98371476377c45324eb388f047aee5b
z77e5d962ea2a8b6df44ef67aa427ecd857e4d5817f170bd242f8a2c0bf7c9679c9941ad8cbecb4
z65e44d7799869115d94621a1c1e87eea0fdff01dfeeb658e50f4c10b9db44309949db51f964e27
zada2a80dac9ea6161fd524b9367f662119e8bfae847ecffce4dbb4b143e615dfbebdfa1c747fcb
ze7b02647237aad4422d465b42bbce5d9ae34d8da41a7d122195e8dd3fe82b5b1d672a65a0c670a
z8ec64ea1b3445e805390e81ae83ea39b310525f616a3eb4636f5435c732d39c738ff155205d812
z04f5a16ca40494e50b4b0b7579321fa65fd535168f5423b71785639489b2bd6ad58759cf8431cc
z6e9f30c3c91b7c21fb54e76ddfa0dc7909088620a16ebd61d39dec09b6fe91277aff3efa285762
zceffc84646842a85639250c22392412f6cba9d36896db8d23f403501909978a08f622676f13afa
ze7177e56557ae4ec2a18f5bfd74ef4a7b13a1a6b668f97e40d34d679748e553aac705476c349b4
zba292a300dec6f150f1bb9ccf6cdd0145c2270b7a97c10f0a79878cdfc0d00f8f50be3e4e483c1
zb51f64a15037ead1e3a6fdda1a9096a122db708c1464e51b1f68f3ebbe0b76143d61eb03f0d3e5
zf5f5595b1f17498866dcfe17b0c0828098d73926829e5d95231f107e7013a0a6f846e11a409948
z966c389d1b2ceeb3f0c331b3e8df1f57eaa9b5fcfe92072744dda446d9de53921e00382fb9642f
z09cd941672b1e4fb3a3f24cb8b3306067116bc081b679d2a8e0bf28c84c5ea49d69a2282e58067
z450d233f76ed9cbcb582e7c65ed5318bbb8c72481ecd5559ebb28d189201f72214ae48bf3ac3b3
z6fa72740b5a7f48398d04fe1ec9916022dae081a9f0ad4c9c2119450bd7978b7e566d60f48b49c
zf28e43f57f1c307c5247744fdd7cffe54e881487ba3cfd02150cc1eb9a9e7dc66657a60a528f60
ze728841552e52251202b962e2834a6b541d031cfdaa247716e7f652979f179b8b7d4fc10facd0d
zf6fad8a1fe50a3ba3d2a7050be1cab186287a6c0cfec3e938c96a220a7d3294fde0bcb7a8fc31f
z7214a836aee977fb3b79b8fe0017aa2c7c2b4f7fc3db00a64e916d0b6a1fff27d6745dc5f820ff
z73ecb845a987a5b84995b1280fee94a32ffdcf059266ff23a26aa56daf7577cb7726f5e4c5d6c0
z67c04e64d4850d382dbced6def9bc30b6127a34f8cde5562f277108f263addf5130a666509f027
zbdb2c1349b0d90397d5bd540bec85f8f2df772e80d1398c594c6c5428c0c023d0c7944d7c465b9
z38835a1518181a0bcacdb75f12a519d53d125bd9f174e63a1def090aebfc6eb17ca0a82fc91872
z9074057d21d49c3af97565929b9ddc6776a437548ff55ece3f758114f92246973c517952622847
z05fa2a8c561d5908aefb64550e7fdba2b015b2e42303bf3743626e5d01acb2ceaa1479ed7fbd2b
z465cec156c1b5d573c9601423d8368ecdb23dbda2473c0f398a7f312148fff1ded2915a84e2977
zce905bdacd95715c3a574ad172f0009b46d88074c7d71d85978f7c50b4b4389329478784dd5102
z816f81d6d3895504dc1250ef8486d6c54274ec852489ee7785c41a2edd24fe0d19bc15468c36c4
z4085b4f0457a73e59f3d0a13667a18cff4277bb2ecfa70001c6cd22cd7a69841a8bfdf532e6f29
z86c3348ed0f483547a3482111f700edbb2bf1a5510d5325a4375e811b4a73cd11decb1668f4b88
zb9b2f1a8bd70828d228eed26e48f9ae331c744bdf76cc41bb65587be5536bb4ff838f048531993
zfc7ed9452585a843109deced3cf1d9593f2e964d35a4b4c58206bfe544168891818fead405d3e5
z12f22ed830cbefad37ec687a2f8ce551646add13254bb73b850ac55c17c57c4faa54f0d52ccaa5
z74ff50aa9a4143d607177af90c8845e5fd3d55d840d2078ab099dc6d7e16739110ed4ef6f6a191
z20b7799a211a1c3a8a6a79add67ac4f61db322bb3317ab8ef839a290b3bfe02253bdb2bb077cbb
z756c5286688cdaaa5cfec6e87a2ae2436ddc99b597885538211b62db958d68f6f220ef01a140cc
z7927213b36c3387c39f06906d6ced5dad55cb2f7089f722901aa7de0ab1daf49ef43c826eeae16
z219e8aed905fba944b32cf973656941375320112dd64bd2851b6ab33ac3b2d0bf9cd7daf8b1723
zaaf24bcb4bcf01cad34775752cf1c9260957878fa03d234b2ae44022b8ea621f7de6bf12668466
z1a5cbd90b07584496ec073bed98f1e589217ed1ebe4f1723e0417ccc7676010f1651c00eb04417
zf61f319c7ed5630dd4d3442166708072f3c6fc6d2521e747e7e460c9b544bf125342b7b93a4052
z18659665e180090ced15b2bd3b05d35ba95a8b0c6209050f09ab5a7acd359aeedbbe1b5fc95172
zd09a59ffe76ccc1d45be077792f4f70d10fc7c62617e6bf1278b6cc80c43111c9301851456dd8b
z1a4e1141975a9b3e9ec1ffeaf62ae060777da7fc9df8fcb29366b847436fc230f88642d5dce7f5
z8c1362dcf5d3786a26c9e257e67f552424673da5d97948311f6b6315f54d6242344d7b8dd70422
z39611cc72d73b71721ca9bc67f17846e44a18b40342ee7928a9fd46a53426b183e1f962e9cbef7
z2e1b57ac200f2c903f051a16dc94db3420f2377a1197b8b0d31c4bf02b7c1ba3970ccb08dd5dda
z7668d2cec4b6089d0c5d030f9bc4ff2e26e5a4bb13da931dfe2e359c7e88e408c11c32ed56fc03
zfd2c2de0328265e6bc17dd3ad98cd92ffd0ae97ba24b773447b7b3d9084abb8640017547842d47
z4a3d9d9959d64e7c5a1a965e7e441e81cd1f630772c6ff61f1fa29756815be165527946fe0e5b4
z45487858299dfe3459817163987888eb6b5851af3e9c492491a7ae081f335b3063e925c5618191
zb66ea38821d4b8ff5d1ea085d9c033091c251ecfa3c0d1d0871a91d7f7b521a600139a50c82d8f
zeb5bd2299ba012d508416c5efb0be0b817c4791aad1055293eaba7e957500c7d1468e8727e57a9
zaf5019d624472cc17d6c4b36350273944c7268edf3369222f6de06b86f5bbd3fe75613380de418
za14294a93f5ca850255a00a6131ef1b0113aa0ccaf1dcfab4cf8dd793c7662ef3f704e9bafdd71
zccf292af32bb74da1fe0dc74f2ef418b6185cd3cfe8ce08e1af5e780f2f482534db982be1b57e7
z747e7e67b9c0f9788b946a19aa5589a58eef3b3c084a69b9474e1af0c3a11d1359136ea28199da
z5c11067ce9d6454afea4dda1ad65815fbb40acb021a5c0ec4ae930e232675fd9cd9d002a52bb93
z7ee648aa576da1d254769cf01c0f58602c88cecc8edc8ad3f87566325e45399c1ccb003f7b2929
z5ac12d47d4dc79bcf3b234bbaafc7bd65bd6c2d39b890dfc8805dd3a39a1453fe73ef68af488f2
z1d38d91c7046ca480f11323b56f0d6ced1e8cd3966a819a81b4d1e1523615a1cd30622f0c7f5f8
zf2d26728584e90bae302b5dd257dd6a66b42d06e7845156ca23f67437a119c73203549439299c3
zc265d52469a1c5f75b6a58396510d772d7434bec7d0feed0af50f26f6d92402664eeb13afa545f
z759d2e6591f096c634dcdcaf56b5f0f57aa6f94f4388e444906406c3e0ae0f2ff282c617adac62
z9079c6a2bc02ac4106d69a20f05860386905b21d82ff932704a855fae2aa5174e53247af85ac46
z67b90ed9f2e9d9244b84f8fb1e1b7c2e3faa1d1c37123f94a6022cea4801a04832c37a642fdb65
z2e2dd62c09fe48e6429ba2395423df7bad67568faa715ec00a3c5fdc883a3b090381937fc1d389
z9b4b8f4679a8fe7ed46ce0f37eeaa07dfe5af4cd30f935d32e459c228cef6511784e82bb1da25d
z2be2b450250744709bde8cfca8c46b05176a1f2508640fee8a20d70e0321746b4f2c695daadf14
zc304991697f0d1e7b5e73b64e97702bef7ac998d674fdc067283c9cf1a254e27ddf3d4db529d25
zc00e4ddc585b5bf0755553c2b0781e2f378701aadf65c79c23ccdee6605de55c65dd4285c5b68a
z0658e7bf7e878b1cdf16c3212b792fd18a84a85338365b6216b743ed08ca88bfb964f0a731bd27
z4858f8462280fbe70222d33b4056b420a1fb7a1a2b641d7940b641efd669652c73be069d03b6d0
zbc071c55de7f55421858e4d062502cf9766d8a407cc424bcaab1453f74a95c9f89941ebb2b14cf
z9f170cb4e1437224d750938233cb7ef21a94fc66ebbc451b365fe6ad08620af20ffa91e025de34
zc5faee874a9e663978bbbb3bfe903225ce2c5245ee18cc75bd2d1e0ed9f89739f6f2628de11ef0
ze2307579bebb1bff05f4a4d7b4cefeb086fe7be89714a8e7463e9660ef40a04271e19c5b29a361
z0ffd1ea344b0cec463a0b4bb622cfba7295de57ced2a804718d46c29b96bc44fed5625f2442db0
zc82e1e0cb428469ea0f19b40830061195184aede727c6b17782c8a59b43b0cdfb2ce616e804a10
zc34aa87a90e3571aa917255686104702283606bffd58c94cdee1f018c9cb69637dd045e983a43f
z04f636a26bd176c57bde6a436f03d8eaa8c9a926771d0b9f80ed156f1b87b23d1387291d3c22bb
z85f4ad5317831dbdb875af59fb192b43eeb6ec18f9730274c2d456e3174e10f6fe2f1809162150
zbc9fc3d64dfcc7dff149cc33c2a219eea2d7d29c65e0110e880b1e5338832ce002319ee8936dc4
z66fccb7de822f89d14596e83155f75f0f09c0464dcbd68842af8e0e0764da8dd1db66488a5f249
z86f9c7a1799053ccf706660cbac28b266ea1dda58d9ee9e79ad3f7df85470ea1f42a8ed840a1eb
zeafaca76b2da10e4998554071f3b18f3a233ac7ed54c3a5c0d085dc0c0d276543b4a056ee78547
z6bebae73c0aa3ee9caf6258ccf0cf3ebbb99731b7508c0d52bbd2886ce45da25c4afd4165b0049
zaa5ea88725bd982be9afa6c324c5902197bfd6cf043935dad9ca906d28430d2f7324cefe27d999
z7e115d235a2a4643bbe70f2495234a76c9da9f4ea00887d7901478993e27d5f52bd094ecddfe5c
zcde20a8301456b1814a93b0d61a931907eb1c5505d367279fd152511d51330cd0f16e6cd8d2d01
z267e4e6aeb9505f199fa1bb44790fc76d304ac69dc68de6a2932f658c5b98b713988c5597202a4
zb4d147ec5ca2cffc5b4cf3216adcb6eb6ac4ba1c1505258e545244c4f6172e1ba56ef7e088c8b5
zf97035c26c21267b10555234f243dff65cfd06189784b42206a5b023c01c7692124628e65e6c3c
zae8bb20db2eb65b4986fdecabcc41bea4977e0947ea7f2487b58ef7350ed248b8537c3ce15a63e
z1f1206add8b00d1e1b7a55a05b9c42634fa3e394105c2cbc773c4131d6e542cd70509addd490a4
z23e06f72e73d1658cbf3e5c280fb95531ea41202bc5f98ce2fc30cd03e585f99bdda244c779ef5
z92bf8f03c0758d39af81d65a51e07643162f210f71104bff6758e4a2fe09d79261d05ae61307d9
zb8a8904da0255cd87d1ae780edb1a045523fbefc1fa433c77df25bc7dcf57a756eb05d619384f6
zae4f0344d5d589f9911bad4f1494a697fc2e261874d30f369da73e094c6a3c51523a5b27303236
zd1899d2e97f6d29ffc5f5d500b3ec9b4561c097444767e28c973bd2843502157561a66bfc7d4fc
z22889c5db9f94ced4278986feecd59e0bf1ce013c8eb458764b820aedbcdc54bd1a735a404e29d
zab79950d47de5c670afaa14649cd7722835daa98d75f2047690e7cbd2891465a5696f243f25ec7
zc2bb45576a713bc5356ac862dc517381dd0f69640c1c1e0eb31d6d3b802dd1c3bf630a907a61b7
z867e67dd1f482d2ffd1e97c6a7fa3d85f8fc0fca8534fd01b04185a40d644f41437e767e0663a9
z533f66c804972969cb8ddc5b7f55895e2fb0999ab3c951828715ad3859f2e254e0f342dc8c46f6
z742caaf74e64c79521ebd410af00f6cfb4e58492519ee945ea28b2ca42be83100c9a95f4afc3c2
z7de2c8e1f234e80d4a23daeaa84323a93d28a2790bff062d05cc60f992f060e007eb1e9e109a04
zb595189336b7ed7f78b221974898aa7a44b08be02d3fa57c311095db520b9e06a474244a044ae5
zab81edc331df3680e76b4470b3662e8206c9063a5181df4801c73eec57fcfe5c54135233e25550
z0e0e70307b7c145748388fed4a2a973f6ecbe93f9e3069c06e8fd708892870540436fd689c8809
zcbfaf54e6d3c86ce8a76dfa243cb5408af9c7a804e9a857440f13fb3efad8d0e6f2dee92fd4a16
zc1c6c54e0e0f5b8c00691669974f3057da265fe2872cfcbc4b7b83c1d4af79b4e5031169c759e1
z760945b5f640c718d9bd9deffca8ccbc20e21e902d06e0a24c117e4669b1353a4172c25763d9ba
z51a05bda5edd5859796c62ad06612b87cd81f474c12fb7acbe75723e664694bd772160f49c5401
zb9169c28b359e26ab0700335467e1e3616d8dfc828f1c4504c6cd44329fff41df6b50901805784
z393067819784ac067b1acff7383afae2438a77c0a0c95519d9b6083471379f20227837af68a12f
z29efda2106d80042b05f5640b9ef25972d43c5e0e6e8ec6d45f26c8c31ea42910632b94ee082a1
zdd92a6dc91b23a114cf51f8b066388483e52ccd05bc857a0607a9ca4fb97b3ed6642d06e6df3c5
z03fe02285b6ee387fb37095e2ad9bd2ca7293f6d228daa0cababca93646455f9428ab7d463ecae
z4274ba0363c412ee3d3af60df0b697fed8f0f49189ad1c9ebdce207d99b7009f8c9a668679a1ff
z40edaa31692549236d9885a2250f58d63ea70305e54fa261df424a41efcdf51b6ea8f4c8456a48
ze53c84a71ed50dfc81d28c573fa988d5ba3077bacb8ce5c22a3999695ec5d519a55926c0432388
zbcf2ce3e4547dce2e77ff814ffd635cee6e1dada8187e6a5396b8f0a0096917dbf929c4d04557b
za6c16eeb94fc78b9d084829edb83974553cb49b40439216433daece627aca9931b20a58ec51b6e
zb35f5e94fcfc1f181f869e9bf4b8f8d6b38d24eb656364d44cd830bdf500ec1b49390bbadf04b8
zd75b8a0f85194105f118b047897a5d3b962198c8eab6e645259dea1b62e4af489b981e2e5594df
zffb048ee2e72327014227cf96b31dc943ae3a7a5f087bbd6d5ef0942ce55c7524f596ec009a7a1
zbd8b8728c7f2f76fc5dc4e90252702ee2639c319e71421885a0265f59f089ad19433f1df4a887f
z6907c9a7d14595d0d7688a88e807a5da4fbb543efc049524f10752b40c54008ceec274c97c6bd0
z50a8f9e0e05c75fbae64da72c26f5d92b1b00f80fec48d02b3afe7b9dccb828d31978a4f992138
zd2c7e7708735551da02e7f2fe5884c277494dda4eb539747074d6eaae296e7e6c9a670be4c85fd
zb931ab5c1af0a54a62035cb42486109e981631dc534288f3da4a874cc2b283d11926c00c3845d1
z221fdb43818dc15d440a55c2890685f11eabd53b1d5436ea0ddbe02d7a159227c599f55700700c
z9b6a326a9d1c0ea184dc548fbdd797eba096fd18bd6aea4ef7341b698cf92ee7d24874b4d26f34
z37a5b4b1993a7af14d634ca1e8d0cf48a7daaa23aa88e6ad4ec7d756d4ca27e994222d8e3cf545
z99d86e585e027aaa779e5a43bbe949f490203f8be67000556fe222016b76cac30de0ed5b72c229
z97459d0d89cc54400f456ae457ff63c9a78377331ddbaaf3387f5286be2b975aec072414aeb7e3
z28623ed308906329757f72168ee68fbb8883d29cd4623a762e566b97ce90b9349eb2be34feaed8
zb3cc220bd3489acf5ea73552b422682db7b5e86349b064500d471675ce33401a2533dce4d840b0
z76ac662109f76cbf76022d2b40bd978f55fcba060dec6654501e968944e54aa127d08b0d2ef5a5
zd7123cfe54ead8ffa21686dbbc4477e43bd0eb4af6daf664f114df97465eedcc7b6865114fbcdd
z4a1a52c678ceccf4cc00a4fea040b50e1ab79656fd4b3326cd9b04eb7821edd844bd301bc3a3f6
z11b0b7a63329504a49645f1f288053ee57d1f4cfca83892816dbdeca000b5ef829cf974c150b31
z09bc7f9181be60d1ed708b2b9571a5849a47a6f8b483ff75e9f8a06fe263d68f82d56028aad195
z586a81fe4ac60ed65975ef3fa1c85ee546eccfac77f17ebc524619fb0d39e32bb584aa29f585cd
z312e9c8315dfbed8691beccef27243e019d3ec0df7d74db97fa145b843e6aba1807129090911b5
z9b32d611153f79480b82aa51c6b0125d02c9581185b350aa3d38a285d49dcd3740ec239bdd5161
zfe3846f7d8a23e78859a4a26bdb46e573af2f81f576ef457c02a6746d8cc48824e05184e26ba30
zfae8e7ed88e3c0cacd604448a15ffc9bb3e586c988b542a956b36c64fb1732722d598d6a378321
z506d415aa3a506488f178125d182dc7a0bee0f327f82f5c4c9e7e06107d73919b5a623c44c4654
z484eca4aa5641e7ad005792c60fbf084eaedd9a4355099692d2dd5182a6ad9ab006e18e7881695
z43ea75decb7a11e0d2bc2342b761a5dacf0d1457068431852b5bf367d89a689b885d0e7f1e4fa0
z14320c0767e431af82f43ae48addd7372d57615b63c1148109fbb6c711a52161fa01a7b58203f3
zb56537dc9ceec8a05b4ca6009771fb94a49dcba96e6812f497dc9401cfbb4447b8d7cb26450d14
z4410952ee2848cfb954847085913e6bb569db1a3b7139e7fba536efc995fb61ddeea480dbc9f7e
zdc538ddf1c0ebfd1f25b4874dd08bf0b3f32533b88ec8bb5d2906bbc7cbfcb0454b2292ffb9671
z0ea6748113c3774bff98b560c41efe3c89791965ae7f6ae797968b5b576c7ca52bef4d1d0fc71d
z90f718b35ad38cd070faff06348ab727031e30df3ad6f9305454172d8f14697014a95d4ab92661
zf1011d9c0dcab794ae4dc232eaf15964f2054d13797b3c04901a4478591f819b1380d5b26266bc
z9b7ae0eab1a2d999602fdaea66c39659673eaca46c9d118906618c2c0060942a456d6976a9ff89
z0582aef4276a073bdf7692ecbca58f623dd6a43a6aae28757d66aa50421682aad23ccd89d5dd3d
zec277e0677b82b9db86aef31ff614a1a762315d062c5bf1b9eb9726d50dbe4000851b4818c457f
zddb41c44c0bd398a121b20af5dd64e7873039d6cb9d76d43afd6489504dbe551b71e9b06c672f1
zd733a69d9ded3686be59b067626d9b6f745ba1a76121db8fa50b8eb3e343d41ff37e5e9ca3d281
z78c87d63695459705e36dfcfee415324b789e19c1c77116e7310506cff7dfb95ac9893f9abca7c
z00f107ecb67ef28fd30b9482d8b9e2b6346e389da79077f58e62835fbd4503f9662a23f4a9e51b
z60269b5c9f48a7b23cf1e9f3ca374643e6e894a1cd6c2e5979a1a0519cc1e1404db4d266077e20
zcb33353f291adf14e2e68c65cf9a2cb9632b8e870f82a17f253782f3ad239a3aef7bb94ba17e0b
z7eb0225c223ddc920c5062c0430abb507b24a78879b76901e05424bf237ed952a737dc71589717
zaeed891fda14f46f84d209b4434f4382bb10bbebd6823733f15850ee9d87d48ddadcb38bc844ab
z3b931609b456edebff5ca79529e8c79f623606db4ffaef67d1e2ec565e5984df0fc01e4ac5a154
z2b7c2f2b3c79ed80e2e25a083b51fdbb74ee66d5649a03ac0ba852055801770afb9bc8f4c2253c
zcab334efbd01d9f4b9dd07ae1e24add9e8c3a4fb61ee1d8cc5fae699df84f194bdf39a67bfb106
za93632985e17d3b897fe3358d39778a3416a51604107dabd389864a65d4419d0c4a936d64d6761
za6a233d72a4b600d59e4356b64149b9af42a3ae47dce44f8f93ed3220dc5ae686638564b14da82
z24c6f27cf01cf84b7fc751d68605ed88cd98dd7df7c6db261ff71020f5ab3332be787b867e6e41
z11acd576bc5ac0a1dacef023313560e6beee32239e613d1962f1673fac863260c28399ac7caa11
z8aac63cc237a7db45d2cae0a196a54b028ba403df956837da9ca48d33881344208c7866d1b0500
zd9545d698809331a8c39740f9a53290d17d1bddafa09210b375b23ee3568048b054b986f588f99
zd60302cf22fcf42bd45fb8b7b614308009b61a2fb146ff207c976aafaef3a925eb4a10095ef308
zee8eea3f8531c5e65ba92cc2bfdac1d6a94d159c3d85d3f17ad5cdcbb6112a44981bc7fc38701f
z06331f50993d7b641f5c964f293793ae239320c83946f18dbbeeca30e892230c9f507fcd366777
zb418c55290c916f0911fcee919093e60f4503e3ca993a2364493ec7bd1721b45f2bcb87f575c42
zcff9723c21956d1c1b8814607238d055bf18f28b409d1a353df9d507f14bafb674b39de79f5904
z3fa56f7c8f2f8176f5eb0991e80726d0ed542ba5398ae5e836283408ef59b2c65c6658d4713874
zbe0a1eaf4c7e2c1be8a0eb8cee8bf761c7bbc35aca3cb5a379e72acf99a8abd41bf04234a771f4
z2f055a5c0022a9627bb4291b3a6641f029617300ffc82668304db3c5be64b5eef3dd37cbcbb48f
z2e04e3857ea9de78a82578eb73f7b1813f476ef28ffcf7268e2c292a50fe42476977e66f8a45ac
z7f98f7a2bc8d43cca403701c275f7bbffdd409c1f10db009d4d02bedd3ba2d8fc9a7c6cdb9a4f8
ze059f76e89dbce5496488f4b5b1dbd94c66f098cad87aa97a72b245068b378b77303db3bddd846
z3628f3af0091e344ff82b239a807b54694ff7d4afc27db18aae777c1f2c684068830d9aa8368a0
z74084f17a5f18979a38ecf0c14ae5583d4b8f2c8b3f2cbb1bd1349c167608879d665d3c5f3c595
zbe17cfa0b3a4049191e284092f5a612f88105d3c97d5e5da632a99e9c0104ed410226d491047e6
z66fce5cb00c142504a18605daadaf67ed9db26b8f0b0af0a6dcaf35ad54db9568678a307e4c63c
zd333d5671b2182f680a8a06ba763122a52ae61a9b154fff1b43931f77df22fb672cad4810c6d1e
z726e4d892a8452a7dfe5511503cd742e1d692b1a6ec4c024739bd27a921fe10835a33a65fa416d
z5de76bbc8e284c66c807a29812c4e3ad4455556e4c7dbc2c8f23e070d88f858fb6b505f250e967
z81529af767ccf1418326448408bed49d9df7746b5e366715ea4cddff7f2bdeec65f6175f871ffb
z83eb4cba0ed91a196d881734290af1ca0d3e710f45e109633c83efea0d2472a9ec0db60011cbc7
ze4c15ae11e3c657a0bd3b5d43036467388f51b264210473d29a25235c434a8d7e026edefd33d81
zc3e0248fb710b080ea7a9466348423b0b8c88fbd26d4c2061b8e0433497932dd204999dc9d0d0d
zf0c4b6b0a3bde01877c24194b7d0091578c886e2be6c67e7ee0ecda1ab9179c279d61de48522bb
z059d3013b423d65d1efa22d5f49659d66cd6b515a80a85e4a586ca38f3f39030c82ffe896f7c41
z26d7539fafb1f94e8fd729fdaf3d2a037d98d6e9dbbec195b833d0137045d2fe4a4cdcb8136651
z28c19a5ad174ce19120cffed89045afffbef68ae4a3cf358a1128a8157dcb2bcf01955ee1a1199
zd862094182f50d65e07d6b3294c2136ce7ba57a7c35cbf109e459547785cd5146c2da78f870ae8
zb86cc3c961e4a91ce737db0f40dac51bbeca04cf2b898d07c1ad5906599a4542e71bce5aef1a2a
zf939c5f2fca10dd7de7fd68d439d1554a61729e0c2188a7203ad53c4dc1342ccee2c0036e2e24c
z3aecc2f458952328811f8d78fb1d969a199502c37a68ff4495a2d030960d6927382c1ebcdab407
z9f9bac120f458e73d4c3c7b76676d62c4daae896a2caae3059a99d9cdd7e93c9884e16cff2e4a9
z47d007243aa938c6cfba4ea15272488e03a5e5a58300e04651a57776c37a96a6e6c0cc79076244
z69269137045e4273fe7381be7eb781b9fca4a7107bc587725baec90bbedde7cccbcd6f2f50641e
z2ea73d8143e49b9c86b659770e099200c90c7e2ec9ec0b7e47c29b232ff0f388d9cf6bdcd49172
z0d9e29da169dbb134efe579677dd269c68b8937e0ab772134e00e895e1f5a2f051e462330a267a
zc87a3fc8ac8fa2e188e1fcaad731729935e926732f8571dc5dec0ea1a86840c36568894bda3ec3
z5a12338e82a91f4a577b28b79fc8b1fd242f19f76c5afa721e137492ad604b3a3e24aa522114e2
z5d9d7ac5c0aecf2aa49bebf8ff1a5c0b32f6d9a8e422b80cdb8f329eb6bb0fdd5cb53535837622
za35e03ff24ac480666cdd427f15414c9d892e98ca47471fe71a9bc7ad4d20ea082b3c9491228a0
z03e236b0e72be7aaa92b33bb9b3878ee063dc215b3ac6e68773503ab3baf484e52169f2a80e810
z1fc820181351a78071b9b302cd09fb487ad667ca4ffb3c740c0373c5a9b79e337f49f360dc7d39
z6f3ea3658549ed141dd33e1c4450f0c476154ef3f3701230235d40527042e02a1a1ba10804fa80
z84236f0673e84974c1ee8a407be4b15f5c91efdf59a2489e7b6cbec89e0f53cfa61eab38c321c3
zbce36f2190f673e0e00cef5aec2988eb648ec1a73d62a8d8e0c4e9f7369bf966a59f766caec321
z2995b25908cec93ae56b9431050afc5a2570714faa1a82b2c6dfaab264ec2565e1f9e0eb8855cc
z55decf7376c1c5a92fd3039f2e965b262b126d7c98fb283889631bbd64c0c17186c1147240cf30
z03fe6aacd395e2e05fd2a76883a42b08a5f860abedf845e745c565f2e418b55373db5b08b226a6
z11aa0dbb92544d48cf0b0e484e21aca64db67451c03f9546523c27571bb2c28dd907a8c28a50c4
z84801d903e924d82041d6e2d1db1c783e78e8c0b9c40f0a12d4934fb2b489d6bb5419e10f2545a
zca8496c110f078b7cac2e9d05cdbb19cb2a1ff3c8f07f9fea096adb7d2e91495f8bf6e89b54162
z27e7d06c854172ef8cb8393d8834e974ba1e3d416debb62eeba1012646e1bc72751e54c9409659
ze89d0a7f6bb6a8771664a37581f0558b1ca527c05c1442c208b13e115efe27b7a4c07dd97f950e
z8c09931c2b029a02598fb0726215feae34a059315f7e93b050b21ca5e104f769b27f8c67f425fd
zcd055a3db1b434bed43e013fafa62b199d24c646efbc18bf114460071b904895c4b280b509f7f5
zd75513141e51dc262c4c09dbc21e19c75dc4388ddc2d8208bdcf23540413623840ffbd20a3b7ed
ze06c8242f64be18a022f54c3e8c218e3e544a98e942f0723fc501059c9da6e2c1a6971305ee687
z9397fb1f2739a5de21e3188402052ccaaebda9f60173addef6df5275deaa90d3b16702ebd9a8f2
z45120173fa23ec67fd69c881d16aa667c871d3876576099836957d2504ed5b6a867a4b852c01d6
za0ee8f7876f8e9890b53012853144d9a891d2b4736aaeeaeac7ac604a3d4193528b3f9ff1d6d67
zd839dadba42f873cfe03e1ae374b7c7ef3d17922c267bdf9d88df806639792b61e803ef1d72b0c
zc10aac7f79f47319c5d9ee857257064043e1a08186812e411b2c23535765622b0a3c79928117d3
zc842b1342f0ada37dbbfa9cdc2f35dfdb1fcb63f0cbe2f7d861a285c33361170cb2a5d3252bbcc
z282fad4cc098a5e0a72f49e77e2a90e7fa69be12b443d45fa70e293d65ac6f06d37c1262475e44
zd0aa435972ee15b80c6b4d9d53a16f13fff635863542240a362b53a09d61db6e8e469dbcb0d2f6
ze7a840c06147194a9e6b5deb9b946ad4bc9884a3a949e0dc0d7dde64d91d7a05eed7554549a380
z9b1780388db53c5bda69c90a9ad5217cc42142252c0c4b3d34a1bd0198e2f9e616d5721a96eeb6
zb9e10b6f22149543ec5ddda3f729868dce54383c4e49e0f4621f722bbc8e2cb5186dc62888f84a
z4cccd202ba327c293cda049fd509d864a795134c470ce62b4cd025d02f6dcf5f0eb75278d60167
z13ae0f20298f87b18d85f7873a2232e33155cb4fb29bd7dee3b6d297a65be3531b75a02786e488
z54d6ef0eec568d80d3428d32fde45407bdabcade48f9a9b2704262e81bc755268e7f71df5342e8
z5627b46aaaf562bd6c2535850c279a5fd454180a44be702852a7e50833e2d3582164ae905f0a75
z496abc6a826b63bcb8b188ab0a44ce190fef360f30857d5f117b28451ad4eb780cbcd1ed209072
z48460f94f0b8465669109fc17328f549faf71c571af4cea4ec06b8fc7e2267ae80e5102da80b30
z88a41a62b4cf0008ffac170349521a9a2badf56b29b19993e889044e1a00f955dc884bed7b29a7
z30616f2dbc29d28ea4ce60191cfe815b9da07c5a5a213a211478712b5b7c45c48bd0682b06f405
z84109d718fbbe5ba9f0e7b3fb43bf780a39fca8eb0776b9ad8e7337253642e523ae1cce7cd9dd6
z36f14d030220cd5b7b7480758bbc4621b80b678bac4f595484d732f038b47d3ef0a278e5074a6b
z425c76b574b0ce4a70a5e3e3c7177121700cabf7506d7b17374783bf74f15dafaac4e3e55cab6e
zbe411b851cb0aa46da256ab547eee3767910e821a50df8bb0be3166bbbd8abea7120222fb0ebf4
za25cfcb753c1e8c74b4d9886bff241c31dd97390071b13896b7a9dfabab377f6f44000368f439c
z3b6b17952ef5a4f9423abe5bf4e90e1f05d4a798e7f73ea2b54e4b8b2aa361a84ec9c66542a463
zadf4fe41b6891c757d1cab7309151d1cea2372ad3b8a0ad3de9f51ed3d9cf6f827fa54f5ea25e2
za2ba798b14886eb67b52bdd19f7da80198e1bff52763225191d85fd225bb8c6f08e55b59e51c49
z9b92213d2fc261aea61a6f40bf439699247ec4202ec6a46f434f8b54eac84bde0f8a7215362d7e
z41bd134e507315ee2aa193fb238a2de361255f9b26e28aea77a309db98e5b97346d767c87e5c25
z1a1545945faa5ef992ccc5d12203e979c63a47ce694218a44c86a0c8af73f51c4bbdb4e54978a0
za6c581bba806d2b6c855fe1e16b500e437734eb9791815b2ec23b9e3c2267e74fd24de9f822c9c
z9c21b3364ccb1dacf1da18f791c928949f32f0a60cd2e96dea81ca22dae1aabd2970c99ddefc66
z9099b3f651b0d7a794ac2088162286227933ce7b3a2cd6bda07de42d3d6cbc7a16d024a5dfdeea
z09873797af9fbf7da538aeb2dc225463abf4851447fd804d12076b5b0005ae97597ae8e4048988
z3943e144da9ca689c160775aab19882b82c78b54378ea67013afaddfb6816eb5500fdf59417d1d
z0ae161dbf83e75d590dad91c60c96490d5002334e6ec54c7119399f3dec673c1ed1393735ec7cc
z80020801450b8466ebb98d27f11097dab6978d7a86229e233fed5a62bc6a08ed98712ba6f418fa
zc13cdb2e0149e3362571e1eb59bda15f5486ecfaa0e8c1c5a4344dae41b2bbd2f659c529e9b983
z4624a3bf0b9398bbdbcec6d66ee2b752ec037ddeac682cd1c6a0dcedd72347e6c36e5a9a9d33cb
z283ff9ca667fa56f2ac1ab66bce478911eb870219823cf0f35d83f678c8ffbe07c18aeef437191
z95141b5d47729397e830e408ccdecb6173c6d859cad0434b9a0f5a1142fa883dc954026bb180d3
z615a18bdb2196cf59ca0548f65c4b1dec7e8f5550725fe4f0acd4e2a0085581bf79d31cc5f2eb6
z2b6be22cae13bae9c4c9f2ac104c828e8babdcd77840ef9630bd7161faf8ebd9b85ba1532bbf70
zb1ef59b0d502aa613d5c76832f1a770e9169aff3ae83e82a895485cd5c6b0592a4f28d866c6564
zba4f6a4a3723f4843b11ad35193f8f9a060aee39d3214003ab55e10cb0a85a2248a295edca91de
z8776f7a2de3faa8bc2db2f0d39e6a50dea152f990325063a5243307c047bdd04ca83de2a07f2e8
z60aa51c3dafccda77e96c5ed1ff0793177e3f099919975bc9f5d35f304b37f2a01da7c572624be
zb122926fff674fd1658871210461860a72b80d003eecba157b6e42e293f92fd32cff2290a28f90
za60e0103a5497b2ec6dc732a995fb056e9cc41e89c30ecfe8aae079b9fa3f07d4e5fd31e93c15f
zee75e6829ce79797af68027a5d8f7b284517f57bf8976389b47664a3a8fafae2208898c88846c5
z9550b94bc05f09119b0d02ce0e97e86fef1c06564a7f49d465bfa250aee5f2bf5ebc22dc857122
z3223e2243707a7b30cdb0800491f2325a2d2a7aa92092be09948c0185add9f1c0333591153f2b5
z6423a6c0198f6b3c57b5b9f836ebe73cbbca2b5ca4d625c5bfa0c05cda1304c98281c93d1c5df4
z9fcc50acb4b7014af12bcc14ea378b8b6bd78f0413fc34412cccaac65e1c411eaa1b3bfb2ec56c
z2412f30ccf65b90eb816317f7f8814c973fd4310ea79779fea612f8f9c925a32bbbd5bd3a1991a
z2e85dcbca046c59d759004ca5ed15e5afc5d4da2ca32a25a0f42db78d5be2165106554b6ec81bb
z2fb02b4abf26c976ad2605f03096ca7d23f1622debf9b5b11b618f1dd05cbd8f6dedcebd4c2292
z825d8f35b110b87a7b0e7b651e5112ea6b4e00b53ff70cbecf50292392128e8232e26353475645
z712f1d30c34ac86de9584c9b7077b16d999bbbd3261b79d1402695f5913b6e3f6bb24c71c1e8b0
zd6abd949726cd33c1f0a824cdb0fdb1d8b9841247b477e9ded6261e27db4510abffd4e38e81c1f
zf9e62a5a18d13631c58585623e3ac820d84aea1a67f0cae587fa2f814dcef7c830cc6d03d39e88
z03f98a207a5c63653aaff9d9add9ce7d290c5f54a95ba3ec8b8ad0b5b1e1063bdcb9922c1ab811
z9e4c22b48fae38deef209903ad74bd2b0dc9d3a01d204bbeb88aabb4411993a9c241f0483628cc
zb8207b0e4bd3c009e850418a4321362582051988e77ab14a41ee23422141cece55ede376e95bfd
z070d6c10fa2f05e42e51be08fe1fe777bc56378a0fd701c0b2f40855100ed9347b79c3bf83d428
z15c9aaf0b9e36cabd10620912bad9d0222e2ac2b8883d17d199185d7297a5a0ef4d555e2f607b6
z9130369958ca8da884e417933fc748cc1c3fd6993cd4b9947fb464fa17dc6db6f3614066f7adf9
z4aac83fc29b095dd605e2f2369b57d07cc1852c950fbd65e51688099e4ee0f2475e660a6a0a9dc
z597f358a7c1c414b75c0d79b254672fce4abd72ff0d773b56dcc6b4f1593d85013cb932a46385a
z762bbac397ebbbd48ec88256510e5a66bdd1836526a88ec71794d31ca95e7b96c02c55a1797215
zf66eef7952e76db44aec8c37fa865a450f28bc4c71893803a1712b4aca6fee2edfa8287d081500
zc40d4d990312d8d7951af2b8b38db53ca34b06b3f7bb59b945a897f62693f4c8806589a3767e95
za99002c49c37c9d0fba552d846c5f9939d4a68923e85193120a1e7e4b095c6ab6a9eb854e527c8
z6c018d91cf3092c5c51976013ae65251e5d443f9494301fc4cdedb744f09a16bdd0f7498ee2d49
z832af2f3c10eb186eeb55c61832229c07ab029c96119cffb944082158656522fad82f5f87dfd98
zaa60ed2281b075ed23e50daf7bc78b782cd0f43324ff9bfd2be6e79b85b0dbaa11404d7a896d1d
z09ec2148848b31fd3356cc66a2c10003d0fd3a5ff36189f63ded598bed1c245dac215dc22317a0
za1b98b3d11b45ba61674ae2392ca4c898e824dcab17ad82cffb40fab06828b46771c87b374aec0
z79b880ed9d9571c1a03f237b627eccc8b551d1b8edd530e7545dc09c4ccd67feca7f5141e60d74
z03362cad877d889f1e4fe6ddd161c6be49b1d575ac60d12a16d83530c62c1182d2ee99d722696d
z3038315d05e5134e67d22b915fe3b9faccbc70fcc18f7cd0e68d12a0e60fff2968c50de99d71d1
ze5dc30af39cf03302a65e2fcfef52887758244942134ffff601c477205194b1c6d476662564ccd
z355779bdb56255de13626a98695c47cfb58849f8f4f410bf3f9fbf75ffc08085562a74d8231384
z1f3aa54fda72df84ac159962cda4d3f6b5300e4fc02f6222bd0fcf30244b8d63ccc361fcdb717d
z0d4452266fefbd4047498a6cbacebdd51890793e1a5b91f766b798899ac62ab6d0c24c95abb5ce
z0b95e968debf8553a1fd88df8903043520bf2cc270bdc4cb8bde787395a24b2795b013753f88f0
za85865e904d5b0420b6997da124139e5de56cd728dcda26c619c5fc7158f589ce27c096ab7b7f0
zbeeac080c3c2cab6dbc84229f341654f21d0af25d9ab84af57e8d47449c40b557f45b01c6d066b
zc6a2fcdc566d48cb34225b07915d7b0152cc102b3879cef1c9814102244ba9312b35cb0747c41f
zd58c29db6be428cd1703520c88d283c9cfbd5e8a97337e40c15729f35e3f02b6a1612256cbe76c
z1a7856b1a0a617b2605a186775c8ad878498b2f1360e67de0132f75258591f4ece0ae025683cb3
z2106c9b3c90a3faf564e1233e47986bde1b3ff879707a83e06603885cffeb73caedb50a1ed2f8c
zebc0634c3443e61642ea094d3d4e42baece56bb840b802cc9640a26bbef2e12b00cdb2bfded019
z7c909c0c9c4a34f4d6705d2f50837c2091faaf26a78fd692fa22ad2875fa00a944883b5eece6f7
z746974997663dbdee8a4ce0f22969fd323525ecd4dd1ea16ec72e417107382ab7f76fe33541a7c
z2b747ddd7d0e574c09df6df7f7679bffdba2671b094ffc0ff84c74bf32410b277069d2742f3d3c
z2903c1756265d72dee557e02be897813d60f408990ae7b555b9339c762a4f44329c2cfa226101c
zfe862a90e37c045e3f0e26f955659e2e590fe6d6d525bd11e96d1f16fef0d6c90e96e4a88e9a9b
z9aca309b8df983af98ef52a5a798bd0933e5adf9f02bfe87ebd13959573e24249cbd54ebab3808
z67fcfa062e6abe23fbd6961763011d413a25517520f8b1d8cb37faf09adbbf166d942bbd564809
z7d026720c76e3f633bf67d60d34094b077cf01ed687ae2b4868af36a6c9a14538ccfd014e8cd9e
z51b976abae9a8a34c18dbac7f6fc35aea518befa4ee1f4476ba03e8b0bde76cba07b7fd7d3b2b4
ze9302d6d80b7cfc9355cdd8917e9a53ac60f9abe410ab5723edbf7db57f3fac558b8905208e838
z79050220f71d6ce871ced16a0abbe8625cf7a8f16ddad0595bb935a8991cc8c21fcd03f98e9829
zb986f5473ce72b2732bd1cc83b9d5ede3efd438a62734db688f1afe544dfc1adf8c7e1166fca27
z9ff0377e2a95241c3d94be8a64cde28882119d1f5986dd9fecc17fb897803f10a7428e681f5d4e
zdbbb93b81e64ee3ca902cbd8eba7f5052dc15bf623afbb5c2d570e0efc63c9787d12a0fd6d73ee
zf0c571b1cbf876d614e5900fae9c31b5e0c4b09be090b9098e43c2f5e2e0ae5ddfa2fe6e9ab18b
z9b252c130e34f94bb927c53188b9c87233314c01ea62ccc18baf34111c7cebcd6bd7741eb4a598
zc4499f34dcbd6f264b817cc67fb8305cda960b64ad328ba236af1277c5769a82d9173ef4855b20
z8b07b32edef9f79174795e0f6bb329ad03325bcc87b67df54bdf58e64802ab1828c062dc6943da
zd64fd655c8ad1606a6858d484bfa084cd7bc899c9fc0a2be15763d1790c98ec6e69fdc1396d2f2
z4db4e4c2341d5b8f9a55f48101a27a2156676373432ede26e41da00fd42b2bafe31a93bec9a1d9
z5dcd5dfe4848ebf8774d87af587f5595061c6bd28a53338499df6a61860f08c0e39bc7a9238b15
z26f73d7ff757b488bba9587c18fe3732732a565c076769d8700f30ddb4f7dbe6ad6345b102b0b1
z84d49c6e00ccee744d04f8ba4e828fd6d72fca7325d54350fa91d49088c86161cd32cb6a5edd3c
zffae197a8f167421cf396d53e3ddcc35ee5c1485ec445a9d6490351bec38cfe502341d5ad878c2
z03ef731d494f7ada8c3af2eec6ada7b68fabec108c45421e5461b43417347125da0065e2301b6d
zc82c4da2b349e1b48032183c8f3dd4863d1d48bd856ad9e542ba7dc36059c3e71bf71167c063ad
ze69940bf2cb3d60c383df598001e602593ae9833429caa81f4c45c3ee8382dfad4cd23fcc54ef4
z3ce53af09f64bc73d54ac9a4b4f5d2090c07da9acfab0acb71792fefbea8aeee4e2d2bc0ce66ff
z2bf937750b1bf313e59023ae5622420db644e4a723bb4ca9010af197ad17d843220433a2368006
z375e20cca9e61354b37e0719718972296aba38191ea1954d2d1b688608dfcb540851e682d54e93
z847706ece94127b6181f769a08ec309df86e185f43a71933cabb09809614733cf43cd85d371d53
zfcb1dd65c51048e89fc4beaa18ed0b83278a3bb2074b5f33c4697e850548fc984460aa9865a916
z43929c4bbb8860c8d08b5fd1f41ba078fb1cc7a8b75327255dd63f0f3c32c19fccd2a238ddbd49
zb9aa92285dd80c6de90812def7bf940454494ce5c598d13edd034aa851f221977887e3f20cf733
z4abc21209ab08043842049420f863f0b1a184583caa5f62071fc2b1d2e102b59bb7751911a4305
z359ca4379820fe4be1c79c9f4cad00efbd68e0933129fcc74ac014beade57689c786987a38f5e8
zb64fdcbbaa0be4b6739efb534d5e9cc399b91599a16a60e6003f0c23c85a14bd980bbd63a7ee72
zbfaa04d1d719c99c649a9939dc26be799c52ef8c86377a3d6f6eede415855d432e93eacc6384ac
z5a5179e90ed78cf3c109886f4ede0fbc06da03c16cc666bfdf9faee0d0e2be02738c9d367400a5
zefddc0f8a7fd7fac12746ea93986894421ff6e20f09dcc580afd90e7585465f7146c75b53842d3
z5badaa9f183f14ad1d59d4611ed381ed881d2bdf823636f6a118f602915f445c5abe6515ea7fc9
ze20662cccc790a5878c088ab5293939918f2b2d61137b9178b1b204a10e8c10828ca6b1a21c764
z9d6e404caf3f7964702c2f0add935889bd0d06166a03afcd1e1be32f5d1b3021cd6286aeeae8a9
zc32ab51ee8b6071f25639dc6b2e6b628ac15765b424a80e661f4ca515b6b60538ec59b4155e7ad
z77c07aeaebfd0a769092a47a1809b2d907fd8244499c4e4c85f3cdfcabd78edf4ca65b54f5e982
z409cbb7e0e77358dbe8ff54f08bb79caad07c2b0c4e90f3a38224f0e8b40585ba73acf9bffa162
z74e90c5fdfdf1595744d09ebbc4175441f7e3e7d6946bcc1061966b7c67da3315c081e4e625c9c
z92b12fa10d7c595a3d12b1031b709264cff31691c24bb954d381ac62fc4e5bb028db80392c1400
z19867c5baace601b4879c1fb14c030c8e2c895c3a9599b1084f97858191039d0fa345724331ca8
z8e828aea4097c851fd3437458194ee0775b31b2ddd4e6c9049221b65f0c80416cfd54b212bbca5
z49fe95f4ac4d671c3aad3f6f475af5794b4d5785682e899cd1a58a84733b763b5a4eac9a101fb3
zb0b0f41cc4fd059e77e99b88ee4bc23c8b92d85b28db07f4a7e6a353b95d405eb934ff378d7d46
zf788dff2f7e334caaa41b60becaf6ded53bbc2fc158416700e7ea271247f701664f96267bf6690
zb07c9f04a4b30fce0f4f9313ddf8ba8de8c3214f4a37b386eb5ee1541e299786d5766da1ea3d8d
z07031e86c4fbcf73e9ea4c4f43b6fa518130a139ca2a99444a1e529c120b23c4cd278685c21dab
zbd9c5e51c2a72ac417576e170713bac39bba6a6af3666d573554836b5f1cfb543fa9c6f5c85a9d
zfcc0a40518a50e6e72325a3f3c62aa12e50b484021ce42c613b4b049ce624d4ff13e3e658c75e0
z92c4a8146da66ce5d16024cb4d9f00a635a760843eabe0ad186a38365e57745700d759abac8170
z8fd1dd534d293ac4b51a983bba792c48f2b0d1b737920e621ab386f1a9bd3210ac5253893b32bb
za634af97ec591f905263abe08ec5d2312eb71c675348670f5a6c1d5494c0443585b2e4dc77bcac
zdd2da7c5422b98a9e2d0bcfb278139aa347bdeb3a3956a549ca9a0dc4bd37fe9355a018193da27
z22b58d2a75991239b14fbbaf5437466e88dfe711cd4bbf758c0aa7de41da6de708e19d8a11c143
z0cc1145431a33861fb5a206e0c6f30379a71c04ad334b9ece11db32c23503713b0614c181c1e5e
zdfd81ac16351bc8735c21aa1a6fb2ec32be1cff3ccc6273511d7416671022b6457fb8e82a69d28
zfc3c377c267020e493f6c286098fb88bcf5c72a0f8a56ba6a0d66b0a8d1373b8d5836ecc8312dc
z1416a68578ecb614f37f3d1f238ba3e708fcb5e396d79b6245c59824990e2855f1a53ef88a67c1
z2f083ed78229ed44db88bdce22f7fa8a435cba35007b9478cb83ad62ee98cc49d358a468125135
z3e65d6512cb7b6a4f727f0c89ed66904510347631a61d707c34eb8764883e90ecd32c829035e6d
z49a79906315a2196cebeaf66664dc8ba69f68e0cc22f34d10190ed790cb14ae7e2ab39fced7a4f
z9c2fec337348007acb3a2479efd68ed1b8f21e6b30c6507535866b6081bb85b04e915c97cafe1d
zb11d8a384ef6eaf041e0b45d2833bee9bff05494eca1bf4f8a7b437e343bed516c485aa8fc54b6
z9b622dcc68b5f07aee75d20e08a14d63629df407249be05c5b526d33ecfd23363d3d7c2be09f56
zad82be055ffc36737536007b169a712a2c860ccfceb8920504b0161e737a9d327c9d579db7c0f0
za0cfa1ec269df5659a1fe3d4abf5191844e9cfbaf9798beccc2cbc44ce980c83d23cd3a05052bc
z391cbacc2bf61c7ce22e3f38959c630d200301b09a946250d0f2a762c624a78bd2498dd26e7b29
zc792844397d18323cc0f3f146be921cf25899ee1466576822aa465c2c77e07b6633fa31102fca9
z9efd5bf1b7c824ba1924e11c00873ab75a6e2090c558f0f0f5e7bb119d59aaeb57eb57d1ba28d3
za888848c31fa6ee16c1b982b93132ad3da23eaf890384facf48aefc920059e3c39eb3b9c8c3fc8
z85a928493b6bf38253681bae3ca484e9c0347db9fa4d61f186867b41581a8c90808043d6fab0da
z66e3574f2aad104d587b7c3f9af2133fe783efce7b74aab8de33c37f18f66fc63fc8ed55905be5
z1382141c49a054a114742098878c445c68cd6b5525229b81d68d4f8fae3f687cddfa52f9012dca
zd68e6d9bfe5e10a971663dad2b55ce9edb2d05aa54163d72a0c0934a5d050652306b9cd650d220
zfcb0ea93b57136ca53bd7af869a91adfd8fe113c6e934f2a9ff7682463986430e9925aa2145fc9
z3829eca476ce931ba96de67c9ff875f83be64fbd1daf314b2c546985ccf99a3d90a14eba193dbc
z5ed55c19f7f8cd1e0526861e2d303828a6ad0d1b650dc779a7a51ce6f222589c58e359f0082351
zd143485ba88b05aae8399917f60ef33084928a99a0a67dfcd7e020ce1b64afc629e384b08006c2
z091a787e5074e4c5b9a379b11a002623ddf43f7f596558d338124bf2bb9be9a744190424b9b67d
zeb5ff953e2ec1a7e7e6129994eee2231e2d3d818e42451a86d5a95d384b276ed2ef157f19aeeeb
zd6ef94338f9f0bff9163b1ab27ee237d30f58760e366412e2f3f7f157253cde3a4e5097f4dbeaf
z9eeb6723db168b47e3f32d0de2a12e846e116c7b1f32a064dec3c51e5953a4fe261af4a9159ddf
z9ce27315e2c37d65ac644f63a4e4b503fb338a78615a59152b5b6bc1758cedaaa9b8ad6fdc3eb3
zbf94e823f48f8f884e6ac51c524bc8cce4a71d3978ae961e039844eceb5b29e5f3c1fe10a52911
zebd253e3a467f0650d19bf3ef316465d8c5774a25774824282a98b18cb78d579d372400df1e22b
z618cb344e8f68c321fea4aba25d3a8050d2151170a103577e55fcabcd226fca59b23de26c70bbc
z98888ea3d2f34534870b23e80b8cfc110b464c1a5f0251d1a95470c2ca78a7f472475ccd0615bb
zfac1d5b0be74f16809b0246d2c18011dd2a2c2f0615752b627517f77fae75cc22aa75f1e63caaf
z4396b2e99eea2b4a86d3feacf94a3f0167b0bb506e97e8829c008623ff82a0b5f0392c22253964
z26e281b906ceda7f2cf9a73d3950ee8e6fdab3bfe573bd488cdf5ce2305ba851ab65dea40fa622
z5dea34829b1ac586064f7118262007c4b339872681c307c6a9d9cd63f4209382f48f45211d1c86
ze4557540819ec0a96eafacff3f1784ebf4fe2d375cbdeaa8d99e2250fd3242ab7f1377ffe58d22
z4946b9f1e3a6d5f244cc9b73ec0a2c0ac00d29f78d2c0561018ada403676539baab3f1e3995383
z053b2f7baf267b92a9fb786382234d321275b76091ca6a2cf6b92bade8c1924ecafa3aaac23b00
z8e9f2b92d566ac0078ab4f4fd45024cac464ad7e666530f1a52c3b2aae6ff2b0d56aaade446d20
z71f3660434f3a8eb74cbfbf3985d1e17a0da10b19fff9705b08eb009b9312668bb470cd2f71a29
z3c556d88710ff0612087838b8dbe52516873cf82b3602513b4b86b7259e6c88fcf3efe7a5f0f30
zbc4d8921065b9af2b0b6b5e64509799bdce2a69e099799fa87baad2c4fd3c225ed92a7a12a1de8
zc49e9f73e8fafc29af6fae5ab8036c5a71f3948f7c2be10ff2a4dc2d8693cc0adf462e95feb82d
z32e435842bcd690aeea2852c8d77eb10b2c2de9da5270bd792b8ffa2aef89d97d0f1adff508346
z6d2aa46da786229bbd1ed93e8c119b86a8ab021c96240a4baa469c9be862031532a035d1d031ef
zf498935a671d329b72052900cf6abf24f74f64d857d92cfe9bf621fe458a169363d2ce14ab7e17
z84e38724bea4990a3352517183e287e1200acd277a2b88b6a6eb9f64e95d04d2a06f24b290738b
zab02ee19c43dc8f32a2705fd91f72dfa33a0652724d60f52560ec76ddd071862660caecb6636d3
z3405ad0537ecbef52864ecc11799dc0155db6051a0c59d4b85b377896fd1faacd32bd1fd751907
z8aa0ebcf57be8a8b6e9c04d430367113b0e739c175657f7eb9ea3a8961f10c0563ad347bf5b273
z1305986899940025908631c998addc7c27143209723b349380f45914c0864e39715233d6a08972
zba6c349c139b5367e16f1f611c33ee566c2922cf2907dc72f2b53b029b68239c4da12f277938ba
z39a862cf8216fc5dfb31e32436d39eb6af271db72bd4944ff9d98f1a4a7534056aead07eaccb13
z6eddc817d81a5957ef1820a4a96758854a688a766c593190fc8e7e91f76bc60a40f45bdcdcacca
zd0dfa1b03574dfa120a6bb7da890735cadbdc9928508d2f72ee7ee4f6cb10ed841a80fbc7e9883
z4e01ffaf95d161a7379130be90fc9045c9ee02b31a75a5a18e80213fbd3dd43b1baf2761df7737
z0b3c9f60a2910f6ab7285af14a369e030417057883a6525149de4a2d1fee68a3105c9ea29d6cc1
z68f0e472416cf61924bcf663c536adcf2e394001a1d13237e635d3cfaff24e969935bed8041791
z1c007f6a8cd67befe481609373f39ab15fee5e05e6e28526419954141c6d537847fb56ae1d09a8
za27757a4cacd182cc14608ee311ff312ae48d4d6d5a8c761860c8db0748c62f92d147feb76b81d
zcd14151c8ceb3bec2b90227f56d65de8749ffa873ec0540232975fb8dba3eca410be53d9c075e4
zcd3f19d546318e05cea44cf0e29e813510d692c5c1260df08f9b7c9ade9ab96d7ae004fa0e7006
zb7524548213fb013d19fd64e257180752a9d7b7bacfe8d3dbe3fe0bdf903fe768626353653cdfd
z05746132a4fbfc371f1f9292daa1f155418a053481963ebeda741ff4b816e4bd5ddffaf8846167
zd99314a990dde49805ef225dfbace12c2c1b741536a060ec701d20f501bb35ea1f0981499ad857
zff9f5f4905f225fdd4f5154fe6a202a2547356bbb738c2c3458178935a558ea2a09af4adfb7b32
z7047f36db7abd6a3b7305cf84631a755a6abc7baf98d7b9049c4ee60d084d48743e39725ff7a60
z4536e007d244fe312ca5b92a564987bb7ce3cee9354432b645616e0dbf3c4da32ac552459d4554
z55b0409b84bf8c673d96c6df426454e5c78f98fd65fdcd86e549c9c822b56115239decec5f914f
zbd2c1380a307b714e0cc95d99d937b4033e923c41c3348bc6eb1a0112fd0350df41fa5961100e2
z0aaae4e9416e4fa3a8e581ad92c02c3ec773c98c4314148ee9513fc4289b61f0bd32b2399a5445
z93ad10e66a49aae1bf9550e2572cc5a2c554cb03a3a9d671b1b4877f2fbbcd1f894782353b10c1
zb6dbd2ca7a6055eb8850f89632126b971109c92f0a98593dd1cf35bd779178c39e100e3d0e8bed
z9d5a4c702a6d2a0dfd0e872250f2842432ee5a96f9179a75d068614d8a65bb01e953304c2d308b
z3064685df535834abe9c38f3c89b8d820a277eb9825b38fd178c7b8d804a6ebd9eac40e7e05650
z214f1e662a6205347a8994e164b4a81e0c9364d7efebc6de63c40634ed3b0eb6761789555c24b8
z3269b79de8799cc925d125071fc0c5ac512b5035f40e5d1cd993584dfa5ddfac397cbece66bfe4
ze07d9ed85a00b422f807aa712cebdcfe1f83b0e4b7bb214481b2b70d50766358057db642aca4b0
z4d3471b707901c8c340a40e3a2bec4e11c333e85d0872a28f88c46fc8a7adcebe322b7095ac489
zbeb4eda3991f6c991c5296e00f8e2e66a29197f621d492719a4118f537f1a28778186205aec882
z39bb43a11b427d54243b8d3c8ec5e38a1b5247dd18fd5b0ad56a8a4af6d39e33d7e83135e83351
z4d55de0029ac46c53a6bde2e87068037dad9403d1ba83d09356a12553ae2af4e7d182a88a3fcec
zb182e857744f33434f260ecf7d5482891c5167366724b81c53b989757c7cb9b76e07d5d1861a88
zb3bc957762e1a91d64e683100c2710ae6cb1a994a97eb616c105e555ba02e1ae60054fd7da88ff
zb35a9af5e61013bcb89162e9b529eebb81e299b523a200e687dbd829db109e85bfe62b1bd327c3
ze28021244e9eb3400f2bdaad4232a57e133526148f225991325c6132fceebfdd1648c598600f9a
zfe684a21a053d7c9a06434251353d75f799c92de0c50972a6bda4606c98dc5d362fcb304178fd9
zbdbc27e12a84f2495a179a79d0661390ff56ac6edab8da4e2cae8070711c6d3b9acdd4c534bfd3
z44c638d21bfb633cfcd0577e5e660a41bb06a4d5753267bb7848ce30e5faa2a4b7df1b78c62061
z1e418e921ad78efba173d0d1d7b0a8c9abf0213d094a0b5ef9954d52d9d9ffbf08ec866f5e4794
z15daaca1ea0fb9b94d00769fe5c6be800df241a9c99d4f89b848d362ed56e8b32454fd67b0ab3d
z1930877dc1dc47bd80bc6c9a991c81e391e9d83af488d6d8ab1bb3817a229377b5c63bbba7a2c9
z3a523466bcc2403300298dd6311b9eeb28d012cf658f74d8e40e7c51c671a49529b942f5da307e
z76b07905d23574e3c52ff883e42254d95d72fb2e5011b7f8d20963598145c7edae5d8fbfd6eec8
z3ac7e8d9e7f5e1d18e6214feaa25d345697226ad5a4e1e993692d8842f37b1e01d53ed6fc98d59
z390821325c3ba4031cd3919d23f81532716dde9d4f896a22f45b62b9ceaa67b7cd06f965e6193c
z8f6e34882ae0599ef59e72f088fdff12cf30f884e9f2598ab1d2a26347a2a23726b0dbb8ac390e
zbd176ea9012e36e01b327252d4461ac2e5b0e42d5ce21803078c21915128e5139e08c4a03c2ae1
z2e0460fcd5f844daac6ef481e54f0f6c43f47c654b9af715f18413c5e74bf32a651130956dbacb
z1c864de443f48e25bea0705d2e285da7c9b7beeaf4ef185b99bc50d8dd927e6b129c45fddcb867
z7345d0142d0230a3be6883a882f79701972f02ec1fe9fdfaa454c03e5d7dcf8f5a1a6fd5981d83
zb131ec09b6352cf0fba173bc6dac924c21746197f425b96fae8de7b649cb9b2dcae9ed1ee48037
z6d4ac027390bd1c9fc64842981050ff088883bbcb42c176852bfdcc3b9dbebeadb2c524d06b3c5
z41f826dad6cb6351066137a6b88c31070d88398eea3d9324daab9c764c3ac545bf345e3f212581
z38d57400c8195c2d4c8b3d4b10082ec5adf0dcfd5e39e8639246fcc486641c981554595b77d17d
z20ae321c41391e3cb83faf900bbb9210140d76668f08f4a44dceac214b06df5ee34157a52b3717
z5854566de6e08448accf8c0213a94dac300f43e648ac43d19193b28fb2d4d5825cb853e7b36172
z842002bb58418b564049cd5634c2b4d2625a491df4942a4197f68528f0bf94ea6253457389ff05
zb0a65d10e0f6430dfec39bd3df755c58f0ed64021ab8395f11e7e104da59cb15d6dacf28720c35
z939cc77dc10b77319f52c6dcb57479c8e79532817c6f0b1c78485920516741b74df015c666f098
zac2ce2398829211580801eb26ca8c4e2311e5ead98169f8e96fc56cd5e0c3c5d4b5e5ee72a22dc
z519e3c540c0a27f16e2ee491da9b9037e9c13cafa500ae71678bab3a6406e4c565b54f4e5529e8
za80d6bb2e7b77a93be78b81addbe01402101d3f2faaf347f257feffba2798243b8b3285d4b1ca7
zb36d80e1175e6a8e4ad2f3154683382753e66516d4676823d9373fa2fdee27268a449488883c39
z11ec5dbbe29288501f2e7e8ed0dc8c41747382c5ca89533d37b141d90faa14a40ac28f7417ce45
zbdc3c8470f88b2e831ec1011ba3b81e0d64ef15b48599020c38adfa6e18fa235fa6f24b2bdf8af
z3a4c40f99afdd6448a1fdffe4bc81d6fdf11cedaa6f4a24558bf925ffe1f37ec179a4e7b7b70b2
ze69af46a45f94b1dfd03a2a8183f38d9fe2c8e0f546afe111c2433202cdd31382b98d624fb3c33
z7a9872292a615741c0cc3871403a27711ae4c87ed0c1c5dd369bf168ed03c666bb34c7c8894f5e
z1d32c3dc96e580fd7cd7b28c35466ecba8c310429a5639aa4da16f31eb1ca4c8cd041f572b2529
zf5f5086d95f5e22a7372cd687c32a4cbb338e034517117fd2c10cc776936a49272d2ece8bd5828
z6f29cb88fddea3903b30779f2eea1a1e3412d87820fd427ddfda00c592893d94315c3a20a99d30
z3da15f43d08ed2d598fb929e0c57f2d3019af5b83d893ed291f41c21a5f78320270f527b2dfd55
z86f2d60fd2c217dc13bc87d8ae07d7224113c6d88601fca26aa7f4a3b87c995bd8b5b5dbfb2771
zdc591149a93dec90fcae53e4f8603e5f863b1499becd01b81804c4e9cc9b6d4afb422a9854f6dd
z2ec467348933e05f08d7aa39fb9021b9c7c94fc7bab09f738a0b1da5a39e9ed4af56f0fdf3eb93
z33f98ecb56ac2a79984023cdf7701310ca2e8b91428850d45f25d2de6787727ad9389d760f5513
zecb379b9149468d15927513373ccc6d2011f02b86af917748b6a89c7113133e3f67dec33174fe9
z6d5b79ba20826f0807887d1b6b4953cf59782a4dc9f4d9948a7b9f14e03db56c37b19d2afb22a3
z0fb8e872ab8dfa9bff7cb77e4898698a4ced812c7fe1865838287c550251030f0229d026052cdc
z4664c2149bd2f63f2a38e61dce677af060288c40f95accb411ef344ad814e6b54c45234cd776a1
z85d2e0193987927f06e3c5712475ff2c2ffb94b54941f85cf2591f9dbec4da3e1210805735154f
zead812cc3c35daf6b145358b292fe07143874c723a769a9999a8f17c1663e1ad683fddae27e47f
zad9cbe573f10d3a312a5e7b9518e2ab98912f2bfca06f0d52cd4bc317bb641f992d4cd380560b5
z84bee5a3d37abaaa0e541fc266d5967aaf40893077966aa8a2150e47e72061e4172db81d03b8e4
z05fe65826b5c3c75184a3b4497db99dfdfb14cbdacd3486df9941e8a3e7d5dd737ae6874e16340
zfdc511ef69816fc36470543b93dd37427eb2c09396e6cb994492fe5ff1a0943d467f1d7d5b8b7e
z03aadd6adb8f37f9b789ab639a8558030017a9f42a404c29f417aacc19187abaf08cf2da6db87b
zb3ded84c88b023aa28a452adc70192a60dffd93d87fc60f4f11048de8f67d5aee5b09eb22d0da1
z61e8389cd95fd6783ff2fd3166d21b23e76382ab0db28215bfd1468b6f65c0864539827be1639b
z62716e22c62685fa08a280557087b0d08bd296e26fa63bf777089f08562a834abe6e8105bcf3a9
zb44f3c56b22b7410c3a5cff0a39fe7605f61da4057b14f43b3be2f6fd073a853145eff8e7682e7
zdde16654a7986eb60e0d537c09bd7f32e5a71234c2e1b53ccef3466214730dc105c507e0abd072
z958dd01e2357aa11896526037ca29d82391d179633a58fdff8a68b2edf8f45c11e69acaeb9c56e
zfd110ff7f673ae77861220cedcccf1b67cb00be1c300de1071d1cf6cfca2113bb14974194d9329
zc8bb278c8bb4039ec8b90fe4e4e6d97ba3a2df68861db06887cc736fc7accf0bd351b773047139
z3c9cc52f6d3059f36cf9c16068729b372e3e33d309034e02cfa0a33d1d020d24f5f649e8ce7b4a
z2bfa289d06ed2d418b075ea5366e4daf39c1f8cdf6028a67ac77587387b98181e013ee6a2c58f6
zf02078e015f3d2717b39fd005854d3d605d4994eca5adfc1b0397afb15add46f7407cb91c57f59
z1937d0f50300c7e37cdab3f52e9855eaca8072e27a542250aa62e405d79612e3aec4856579b4b8
z44c922e9f578a2500092b7e5dac29b70936ecdaf41d7d3fc3de777854d7acf99b64d0fa52742b6
zf78bc3c29463fbdcfb311935c2240678e1644f1ded9e048eb8817360bbdef21cde5746690b57f9
zf434c7e62a1d85a4b5d5f234e9b4d35cdb3533d313d1b1293e34dbaded8f5aa639ff50359532bb
zde68ba51d1dd75a4b19c046ec88cbfd14f0a4c789a9431b48deade29c095af0b863b266498a684
zfb427b7b54a8ad61f7bf5691e69c625b7a2a218e3d505e0bd51fc655234e73096217b9f4923932
z68ea37cd63a914efe2a069e2a64f624a27060d8eb63d756dfd130bd3a5dd046997cfcc51cc1fe8
z0eceabfa379ac26ae2639abaa74577b352de0b366637264801cefd928bd84d715d03fbc36cc883
z5338c502d1b29ed47d6a175254bb0beed81312ec8916e40eadb108808fa3f39e358a3691e7ff87
zf2921e0baa66723a6f21585f56a22c62ca6507821ca8ed2530cb75c5f72daab8e0bd171e340822
z6b42953d8272ef039bb8dc9ab114b399e30663442a516b2571965fdf5ddbe755e665c67f43f51c
z4ab2a020bd9e7f5f57010906f12d7c1c2e3590cc402199e9d2f5de951253007725b7febf3a4292
z1299e356fd32d741bd22e54e7b5a31c715863a30af936a658c09ffb278cababed4a1ed3fbfc666
za2d683e31f8dd03530b1607a7d8bf939bfbdcc01f1ef417a17c09efc5896d3cb4f57516de56f13
zc1759c9f6d0220e7500efae01ef937882fcc58fa3f864cd35caca8bb808d08ba7baef22a219155
za73a9e80ba22030fc17ad12b92f399d0225c49d97d6692105059636a00224790befa417b728ce1
z9357c3edce7bf4be7f5b4893a4c2d9c60687a23de81265f4def7109806aebd3100bcee8b014988
zf0a886639190f1000dd5ccd0f6afa94d6532b5ba338e8492578ba7cc7f0c3be5a5f4cd1f94e1ee
zaa495bf97b4ed6d3304390ca0bfee4f12d712f5681576ffa097e3abe3c42b9590da8e731078834
z3fc338d04bbc55824abd1650a3dc88713eecf06af30a30764565b45fc91693c836ab796ca287a5
z67a2da042b3e3b9adcc579b61b81152b930f4d6a56bd26a06cbff9423266979e299d82f1adb23c
zc64ab5de18056b1c2ea0458d43a8b3fe4d8c346b136d674eaa579ffea7a640f28d8035f3932913
z5bd06b6f60cbafe8604a28faf44e6ac63ce3952ddee3716fa782fbd923498db49d64d64c44abb2
ze6e17c619edf4b613d7878e6086ab85c9cdf926c51dd56c863285990dab8660bd541cf2d9c8f86
zf48d95d73df36bcc15f4e8ee7a0ab8b6b83b46957e262d85b84eb373c1495dae71ddd77a461880
zdc2c93f30df6a6e5295464209ca148dc72e60b340169e24110d749b8ac930b3c8a3e3b68f349e4
z61b2f8ae332e32c9284e35c9277656e4808d4ab5d63ad524351b144151fa5d1c07958b3ea00a38
zd288f897de9f17110444e0c6c4cc33c9096bf35d64f0133c3adcd4e6be9bac67d59b6a30930974
z5ec1f131cab83e02343026e4454e30ca20511ac942e8896269900b47486e8e93bfd0e0f0df108a
z1e1a56954a2c67fb4fc30c810148db1b281087eede68116b9d13e61fe5cc7dc075be568ebc2c0a
zb0404320919eb95e47db32561903930ad3ecd9e56d455dd88ee323e5fd244f544ded1c7c8d3f0f
z794007fadc8d3e3f2f911e3b76e574074a0334b85bee03dc1872dd56a5566dd1fc4ce0a183dc41
z5bc5124b59ba910219e078dbe43385110f8d13cf8d930eecdd216c90ef572ea22694624d5222c6
z5e303d174cdcf00ea7bf22ee3754a3bac353c82ac5492ae9bbad515e4ce14d0d1dc9fa07338c4b
z5c3ea97d106ba4c68d81caecd8c83f92b5db220db6146ce3e14e80e2b3753c0926d1316bac8599
zb4ce7829dce744292981d254d859c9f9ee0ebb429d5dbe46d25425abdbdb1ebd370c42d0fc9ffe
z5613ff32b900dd2e6495f797153bbda25e81def65fe9effb89edcdefec2d9b31f213c9664ecb12
z5e224fa57d3ad535b770f889d4819fa86704026cde7b8e8f5cccbd59fc390535f9f495643ba88d
zf2bec0b744b066841fc73c53e939c1a1b2e28398a13339616e0ccc80890dbdaf704b91c4b35cbb
zc93745831c2d80641c05226a5314613fa1e467dd77af941f833790e9b492ac547748bf7b535bde
z1c081bc315733005682969b825faf8e843259eeaa40712b63a534a42925449495ae4dc6fc62a43
z29607e99e97dca5c5cb15429fd1e3ed74bfbf7fc44c97ee852539bf15d598c3c6966dc27407178
z681275f8c08c991bb6574902bf2b263a6dd4e272ba7a04a60b10d0858170d9aaff601e266b8889
zee4d516094fcc41240b9c09e18dc6b6f13587faf36e6ea59dd0aaa310d7d8c0916158f6e031387
zb018dce87515f73fae3efba05ab4e6569c1a0007142acd70ecaed8ec7fb0a046cc26747fd7cfe8
zaf5ae07679723579ff2892b523a2aedc23e1f0227089f6a66eeeb8fd64f43f5b3214f816c34aea
zf04423d55a16f8ab32584db71f7bfd9a88be9728cdb28badcd9b59e8486bee7bc60da93cdfdcd0
z4a275f73ca80ccd29f7033b32960bfb0ac7ddeea0a47391ae51be758e6e9651e99d62531baf791
zff2f27042ed6ab6fc30940c719d746011901c8a5dbc696d4f54e4b5620711aaa7c0cf026ac75da
zc2ba6a497de74835dc50410350ef166a06c5dce9cfe7b05353517ec0fd1f7be07b192e97122a3d
z4aa9bb77eec07e1534159677644f1ee7b7cca6fb2ddae2013d5d0a62a36fb559079544bd23e15e
zae949508c1b31d43143429204058462432a4f3a5b9964426996771e89455c4a757f00ea60fea11
z216322ddf4ef6d132674dd29eadfbc0cdcd9bb31f3fd6128e7cf1e6e331f4364ba4270ff5a3c40
zdd5a089821411b919222a3600f6e9e5e97a2d6cfb1630501d9a06ab4cbb2e42f8742d8c773cd79
z5aaf3a1aff8a59775f634a0da3bc435e04569bdee890847ffa9d28551d26fce56dfbe751ea4ce7
z700a726a592a002772021875f2ac327381c508563acde33e4011da19d72db817a62ae2c76ee3ee
z666169e922b92a2ab5b812252609f5840cf41f4190b8835b7be14a9fd7c065fb7ad759b155f264
ze144e6f5803c8674ca01011601c53434c79aceaff94709fe73f25ccd33c4d64ae708cb61a7d262
z380e3a075ba60f089c0ee719443dd5f0038cec4e4ab40ec95cabf8d8874fe61b23e5d7b3c3eed7
z83d81a291d5de628fc4705f63e54322de811d8a691655c5765ba50e30170f563df87dda5a57f98
ze18c1d6a292b7f61bd73230a3beda4e245f2da852a97cd7d9a0c1c7879e9b8d5565c7abb8fd49b
z6c6daed145208ec70018bef517e2d83fc2628ea8e5e243311a1e313d5e9d1e209de4225a0b1d96
z3512cbff72b92f4b944914f4dd62d9c178986941f9481d5de80f47c40ebb89a557d8194f555765
za2f83425dc9e9b919e53e80cf70e63848054d957ed6f81c6f4aa71699578245d669a8db1cdd329
zb0dbf2fbe2e85afa0b9b30b8e4da10b2ccd88d24f9ac195e937ce176c5cc5bcf834a2b73e5a05b
z0d1775d1a202340e0b945bcff12fa81e5c12b4a8ee9ffdd97b01d39bfdb3d09945d3b15a62366b
z187f21c719f6737fafd5067c1db18df572f61ea17c94bdf1fc65571c0e43ac36995a6e649a1d7a
z275d5a68248f0989d13140f28eb45690649f895102d0ed2006d48bb9b79fb760859c928816488e
z05b2f19a617332acd4fa0454a0f2e97a8d8e5a9b6fa9edba3352e81377b8d3567c3b78f0f85e78
zd267c3e4cd1ed0b52e71e5d7a621b41b8ff859f0c8021966ce7a2dc8b1406b83b4f09312f161b3
zfecc45238ff83745734d3ff5eccd3e3c50ff1c69bba5cc65f0c653e4b79c5f03370627a3817ec0
z1ab43b667e192944bf1ab14798712cb6d31e7cba0ad0fad5f126fdc509da9d43dd6c16f8fa851f
z19133ff02f4a6958a1fd5ac30bebaaf7b5caa2c7d795878edab86d233731a844ff3e6501b05068
z13cfe11ba6c9464a498dc961d5d6ab7c840be154828be2989f46ce0d5d1d14bda79eab05b7e0b1
zc45a851c21f3da074e1fa9d4c9199e8e9b6269e052a421100ebf7a0a73b90e8ad214a430ef7c87
z8d87ca377c36044a388bdbd0f73a2c689013a6fd27c136b98957a4cda75f5c0f0809ac3977f56a
zb856a2cf886c5c35a55aa2d13362037ba755faa7acaaaeb2879b61990508d339487254e2c23604
z2d7b731e529cbb269d2d84ba25068f1271c6949aff332d68db75a59d80f5b81203c816228c3bca
z4e6aeff8c2142b53c049bfd6a41eef70de8bd4e20723640ea6f211683f9e250df0dd0ad93f22b8
z4c5a3a8d53627145c1137203deac9a6bc3b7edb5f75438177b5a3eeed0d3ddde207e27f8fc6641
z752f2f11a324a94e24811f5ad52a3aa64fa10f2e73866cff0fc5f73de496ba622a6687762d9af4
z3c0d4232a79b389005b755cad30a8704b6e9b00230c38202078d311bca4b1558bdf8d837ba12a5
z89ef4fae0dd72a1b7d37c6ab5a5708eeda652a125b6c33677e56ba9d10e1c7b6d5baaadeeffd67
zd1e79077b43314c4df7dbbab608429da5408508aa8ec90a4311b81490d6e9da1bb42823270ece2
z6e7e3a3cfd7c3acc01230ebe15eeb3495affee37f06fe83ca6a2f9398e887294457449e60ada6e
z848335ccbfc0546a423f5e50fbf84d1c7361f29325f9883c18b39033d2a512d1cabd71fd990f22
z4b6f6241e5357bb15c2c9d20e8e9909475b86254dd5ba0b579ea924ef400eef42920b0b06e33d0
ze379739c8f61fada1581bd2504c6d79ad789feabb7c6e7f690e28fc4cbfb551f49bce681e18cd5
z0581fae319c79edfe45bc7dff4f2b9213775ceb33a331c32e1be1e50a3e1a17364df7b497e231a
z4a582a223d4047628e3dd11f434f9f17579dac3a498098736fed3395c7119d14560846414f666a
z9526b6e3c087da079eef599e97805e0b9c1edf56954d2ad9c55022d48d854f34a4dc0f6ce5e793
zd22b53f0aa9318b1db187f52f98341ab46076969e81d60ed18ff1abfb0dbf5f1e7b7b68f4655d4
zfda9f64a4ff3d0ef8d33471cc4b0f75333561b2cc49bb898fd233afcdd296cf5207ccdbf13587e
z519dff8abead42f62170c2f8b2e6f9f7aff1f7e2a42be9c5008b4f9fe353b76ae0a98348cbfa38
z768363c65cda0bac202c22e41fa07c0ad10ac81efdf9bcaa327b1f1ee44c0b2f0c8e9018f0181a
zd032143057b605079ba60ccb8a5dc546fb2d26b2fde0f638ce496764a9eed08f26788b73636621
z69d37f0ac9744eabcce65b807d2c96d954cd33e15b642ccbf5512ed70b16ebbbf6b71b010382a3
zbd33a949c33ccf0179707be0a250f4a759314c7f37417e9d1e0d024f13414e24f7d5630d90ef5a
zeecbad3f409ba5f20c0d3d999b6171122c5cb5da70f081688b5f23369b07073c7397dc50ba8dfb
z2799f628dc5c94ddef007c4100a8c46f1790b4bc4cfd335f3f23a16fb74c5d2df763126ae0658f
z8621e9475f45c80adb83ba46a9472be38ebb97601fe7390fd63a1afdaf97be44f05fdc4b47c2b9
z39a79b537750833c8ec288bd2104d2ca6c2ee91d5b1db445c8708ac876afe1a1f9c674fab6929d
zf8d90c3d230b9ef89c1cd95f95bf882d5749d71ec70ac01dd6c5de91de1f00200fd6cea8193fb8
zcb4c31bbc56fd0febfb01f8b977d8e0c1e6a3157a51649c4edfe81aaebf3762eb20173eae4c19c
z8cd37f966b2a89d38d872ccc6fb51646b036771958f261808632a082a06b7fa6b4de31934dbff3
zc93bc0a626e3fe62e68c2385082862436225ecd26a8d0502c2734c98a6ef69dcf80e493e64d5da
z82e0b195e282020b3437d8e181f30e53d76d10e635d339cd9812cd84d66d2b4599f6a66442d3af
zc5abf4ff21de9c9acfd0948ce9bee2d7d8a483c946d9740d097c00964f7cd24251f684de3ade4a
z85b872fd7095a0e88f61c4c05b4236f4ed55a94b54e92d402212c5140ced9ed3dcd0fbf7f7cfbc
z5e5d07d17744042e23141c8bd35859e643f6ab5a1c59adb849b966119e9e297c01f02235afd503
z9a8131838e9ed2244a836546424324528ebc6d97cc567d4dfc4886575e4852719f5333472ee50c
zc053a9a3bb27959144c0ad8c912c169dbecf30333ceba1002a3e73f3e9802f3db6d34d2c0fef4d
za550e8700b61234bd142c1ad04471481e012a035f2634d8f9a3b5be697de11c016aaa80d8262bc
ze064a63b525a1fc09848f8ffab2033e9bdd5426d7d6605cfafdf57121d8656f0d1ffa78c614118
zebdd8011ea9e7ddf52d0a5326ce4bb67d694d9e6f6c49c4dcbf77eadf71bd0dada972d7e675caa
z7dd35bd73882651cfb9e69311fb2bde92ce3bf7e4503db984445329ec4f13cc6df73fc8a1f71b8
z741453c2f861d8115cc68392c730a477f8151ad78dc209c6778ac5c15404a7fe9e77454e9d6bc8
z80570ddf8344cbc4c0b6dfdb6a18bcf1d1d2200c282bcd23a56dde44bb5330c563e8bf4657e153
zec1b80d4ee9142179f6c18af60d2831b7d8ade6e4617d65230aceb9f1e57bd0d43dcfe388ddfa4
z82f6ab4be902e6f46b83579ce4d3be2690b2f79ef44b089bac335637c308ee9f332765f1f93aa6
z48852d71100ef80e18d798bce97c5361f4af1f7193ba6e3a4d37b203756b9519266dbd29968b47
zf5a85362b740917054614c887fb60c976cb48918ad526311b0a037cb24d0d7bb476026437468a8
zd65daca9fe26612665a70948b0bee11be62e7bb8d04cee67cb0b426f56d53c049b5ac0fda5d9c2
zabac07e0ffc90c7b7b356fe70861de21e678a886cd700b5006722352edbb7e0f2f5738d7dfa0ae
z8c0d7e73de5acb3c2f8e95bfdd897e74fb000eb1c6e3bdf3468e230b3a498e4f5266eae42af255
z8fbacc709861746d31bbc588f54f2d8d10c9894c9b5908e8f6ca017e602b49cdf8cab35c19bec9
ze75a67db058940c2d0d81cb65899ef7dc961a61c5437429cbaa7b7b63a1d7ab28b61b31c374577
z06a4cbb2425df9e024d3bae2b28b79a34e4088d82af4c84a93746547633db3901551e63159a870
z7fb3652f9735db6a932b39a36f3d73c6f6b76c7b81ea3cd22c19b42800c92f8a914746b5a3ec6e
z024bcdbb60eb4a18532c299c3d0a6d709875239aa5459b42eba7a870432993a33aa9f9e7bdb239
z926383c8aa70bca93577feed7876f264364644bfa91270c8c5972569d60a3d1a08a9c2e41825c5
zd60ed65e7860ba1b58046bc647e5c59d8d4b7c145aba24fd320bceda837ff6eabc6b17fa1a3885
z0d475288dff26e6f52aec8cfeed414e1adf31be714d0d51c835a360779dcaf1235e531ecd2e110
z62a141218a0bc807fef23a27bd9daa18396b028530fb086c7483197efcbf90dc87d7b7801bb2f7
z17a8e1eb861c0abd4fb9d653665792473d0036fa3a6d5ab713953859f92a13c5b7042c4cbf43f4
z26539daeeccf333f6fdd5500f9d73c28479001fde6889527555aff25d51ada5bec709b0ae99762
z33ec549aeb640647f81a81439e92dd0d8178138fee77198be88f8fb9c1d2f7500e16e76e8b624a
z827aeaef3ed7d5e51a3fe68ebcdbd16faa6ad1ac6239492e30547e48f14a96e088bc9e57bd9e21
ze1d4511d576f85885fd757cc310652ff974df0e77ff448704b104f8168f8a42d74945b33a74a5e
z39fda7b58bd78cd7c86a7f6a0f50a0b07ad83d157b2fdeac05d23b6a13a82115085b2dd628823a
z109e7a60e23e7d6d73f0ee98baa74161961780a432e2c0ddf191a9e805e5ec685f4d2cbbeea98b
z657bb709ed41fa83fed441b5982a9a002b3b119c018bdbec3ccc4fc583072df35819d53c15e8d2
zfb7e701b8704f7f0fee1bfaea1a20431981303500ba5fd0817dcc01e8c6f35ca4b5f7538a4fafd
za6dcef61dc3bc621a0de9bc2077ca7557dbc58b0a53f96fc58421b7d3cda2a7b043aa96e212267
z9404ffc9a2f0bcf3e99f435641bd884038d03afad0e9d1040bd77282f3f54387a645ce911c13b1
z70616f2d34530557da401e9213f0558d71ed5ecd081157223e7deb9224c07193f4dd6e541e7a71
z949947342a099617f0e85fc98e0e86b155f140ca11cc79fe344849f5cb7cea5f4a12b0f1002709
z232b2f0892b35a73299efde8c655ca59e0371ad14f0cd0679e772df2bb810dc5819205c5cafdf9
z1959718a1d4e0a57b3c3ea062795ac1475082d35945f363b5f48c18ba905c815f98f1e6e81c84a
zaf53c9e8ccf6d89b43f7ac8824d08d852f39e47811047bd6a800a0a13dc563798942a82dd248ee
z85b7070278aef6839b18feb6f88576bc90c811ec5ff80fbfc67f60f9df96b8a9017b8d5203da84
z3b2102f24ad0bdb334fece7a85c75e35b48f257811a2bada0e2e18ffb91269174573b2fdb6b733
z8c9c2c74f674fe7dd3e5ec9204c0e748e07cf4add743aba0f681787104b78342a1c8c1db2c5279
z41668fe6a1bb9ff475525682653a874995c4eb779889cbb66c37b66b63443340c049c23c15a438
z6c2c82456e869e26c94277b109cf65bfe72f3ff12f6e6a4ceaea8168adad888884ff72f76f6454
zeab40f792705edcb73a41f7db142c4983127338734a4a360d1a9ac514b6b61238553504d130251
z6f8a361edb1b0b08807d0497f3d497426604fab8e3269c087f52b50b5e9fcd7d39e5e47a6a19d2
z0a030883420c48e777ed1a3792e55c2a2da725bc2ba30ed3b103c3241eb781f031867eeb2af23d
z982d918eba391a348d0147d77cb7e0f75dd399457188d90dedf115b769084cd513b3c98df49969
z83119b8aca8ae62e773b2d976432d8f15f10ad4d055d552bb200c022392a9d860851db9c9c1474
z9dcadf7ead720a846bb553fa6fbbafb2db14bceb545b10c348914307218286f92219bbfe887a00
z3611f07a936900ecf86bde64a3232ec68c499a2e45ec3d0cb60a66ad9a58ab2aee3b570710a8ed
zee7a122f5fc38729acf9cc52568a38c0410bf1f44ff3441702b6838e67310e28ceed7c32826d88
zdec4fd831d582305f3b5132850762ac0739fd5b437a8724060cc4b3fbabafe8b2b41b239dcaf28
z502c1a52e4ccc4caa021f59ef7c6600541ea4e42bab993354ad676bd263898d46b689d5067dacd
z33fe128d3d4531ce6ceeb7760411dc157e8af347af1fb138f6eb1351f8edb5cc35ed853e074f23
z63041801f1c6d6464ac54ca208720ffde2054da00e0c7ee59558863f191370dff939581288ee7f
z1ea90615218a214e566b1e7b22e2b8b1735f3561f88ecc9fb4a7526f3c7541e4006ea65be342a7
zc1346a821dfc2cc78d79ef92bbe208fa52fb97b07c7e44340254281441656c9695286e782fdaaa
z3b599b080c8ca385eb5733360ebec4ceef7b734c6ad5b40283127d3a297d95191bd914116cedec
z91834d22aaa5e7969ae53ef3e5a7d97e1585be9aa7188e44c70c3f23f2b3c207869d0a99cb5f47
za815c8e9a7b6dab39342f176e63c5b16ada2577adf53979d4390cde8b01c352c8faedcebb22e13
za4e313cf1347c051b6c3fd844b74f16519988d0f9f7f2d3fdd5a2fbdefff2abb8ff13a8e873cb9
z4ccaafbe13c202f14e0fcfcad27f70461359542fcc1b86fa7d9bdc72e01a8f8ef4e5c6100b6731
z2e58ca1d0d94c332d2c8959d461b46cef86dcb0a6645a93985e8a62bca6bc603eaa84ea045abd6
z43b26d4ccb991c8f5680307b6da9f866f0ffa9f7a77590ad07f81fd59ca566a7b764c16f82dda3
zbc9e6e000f123d49f15538a6b0fd604b42f875ec3f921c8bc2eb35a9eaa17a24e0b1bb7181fb97
z5cbb4d91c20b0dded5130fc626782584a42770e6bceffc3d5dfea21108ea7ac89bc7abd9d7fc43
z23eb9f3d6a29f2d36a43d7ec67b367d2ddcbfc69496bc8e81582fd28b20931260f16747cc774ea
zbbaf5e6c26217a5781bc3ab9457e9ada78523906a5acc859895f395e36ae5331fc8aefd31ae2f5
z308fd99f6730b19e053897bf3a179900da02d2d35cece3d9fa65e9b3e26ffdfe8c44c687b69665
za58c3851f677bea9be68a3657fe889723ab02cd1c4877093f5a444465aef70bb1d71badd2764ad
z9d45abc1eae626c2fa5391b9213dafaf2a742e97d8781041e1bcfc5fcd440698bf40fc94b5840e
z8cfc2fc858be908216de8326eda92853a7bc4a462e596bc54cc2c81e35f381747dfa0925109142
z3557c5afb8d2c871a8eeb6c0df6a454c7f6a395ae00d08f26683ed7c50422992e96d28226d0e9c
za6d65892d1e5e9a326080f34cbf7e6e193fc9103f412ada5a66e2369a4d0f617b3c8eea4d7d083
zdbda56fc27247b657b65907718a668df97760aa8e6cb778173f52fbcfb0f4c6cbbd879d86db585
z1c83d68832f2184953d86608eac92cd44452c3d22c291ee1824bae2e964305585fc8321c2aba06
z37d6611284469528e5518803929b14acbd475e46bbc1b227b9060c6a060ccb494cbd6b2e51301c
z0053aa70759b8b458b194e6b0445103986391971b76f8062689971e4fd4b289fd14bd2ee865f42
zd4ef2e11c514224c84ec676aed74eb6ad646a61b391d5d71034585385674f024ff9b0e22782188
zb4e574ad9a5d45b8708345dcddb41926deb6fd8dc38bbb55c7521e5f7be23572e17cd73534af08
zc8b0fa814af3f47e62a266034925dd19e19f07df5dc470934af19fde7f9d852b94270a016dc488
z18a6c35ef2ba33d78c08f5c4034996a5eea16caaa855f4f7fd6d3ad5def80ebf1a5778c79c0287
z305a8a6b1c407efeb99b6f426b1d8e42d5ebd8f1ef4b52483daa30a03aa679461449139a8da6ab
zfd680b4c46d819f4e9545a554cb8b85c9d392b08494067f20bd4812b5277c2f66572316f9b2dff
zb44dcfcc28e1292898027103976b532b6015dad31d772a09eda6c04c48c95902a4b193ee22fee0
z62174630de1527982762ecbf84ecbf92754f6aa67e81e3457cf6ef2216981fe8d79e233725011e
zacf623495a10cf9947d4c580158f38379a064ece987f48887eae550f83ed81a8333d238a364d73
zeee238d9c5d2b877538e08273570befab87efc23e3bebec378d4e34a01f92d19f2804670ff3eec
z97263a6e37117bdeba991d8cfd75a60ac8f102313d731db6614ae4472d5dcf388fade62d37bc71
z71eee3cf10838f750afe9239ade5c94b34075e2df6e2af31f08a8e9c830a01005cf54c714fc58f
z0023eedf0a1587f300870f0345b80096b86d7fbc99890df9f493790402098d4507294d4f080b11
ze887a8739ffd63b1c0c3f27b200e7055775e6ffbfa6c0ad38f3fa581f8eba64f523c42936d22e2
zc6c5ba01b69fa0d376392ecf25eea891284f37c5f44d75d161fb424d9f277a97642600d3f323e9
z0516f2add6aa7eada6b854f08cc77b64e3892e84e55bf164cf42d23f335a9f6a5f8f5974f1f0a6
z64f55b9d84ed3c1957104bd13241e75b5147796e6c0d7473bfd4714f4877698edd76005864b165
z72a0749334ef3cf56a3b607cc1fadc70e40f17fc55e96ce076cbc5a5baeddb9f2210ba461724d5
z19e00070e9188689a4e9d7f836b201b48918c49322d6d8b3b06cfac9dc46ccff62aa019cb0c38e
zfc59576c1f416371dd6660b3b3128ab96c0f72b936e0e5906927f10f6afb1575e6113dca980190
ze1cdf4e719313a64169a8feff86b0c2f19dddfbdd3b1cb0735e78a0802f3a718703b8233fb847a
z1a09758de094dd444803ccb244f8df99f7404afc53eda3fd6a0a0a69597defa51e223054f8a1ba
zcf544d8334dc752f0de5671aba149c41d0c6cf1e6e3fefed2981133e1e563f87da8554c46809a8
z04c0efc21545f6aa2252f82e5e21d9afb2f99b94cc32dfb8dc18ceb83875ac3e5f882c83d52137
z798acb5c4510f2bb9313d5a9db532cd30cf3324979ff111eb1d0d53f6da71e2204d504664d8d3a
z91c724c13d4da2997df8c620b6686f0dbb9d75496023cd1349f039832c9d9755afcd6fd39c966e
ze3b47ddf0f1c671c0bd3ac215bc38327a70c4bc64f02dc6a3f374a03f6f5d7521cd9276d11618b
za7c2cb7d9f64fa1b37b0e8dd480c172fb2ebe82ed01cc1429517ff1ffcbe2ec9fa853815bd8c40
zd596f28dfe166d94f190d32490bbaf89dccb8669320a792a4643492c56c70140f032107833de63
zf45c05c28477c317dadcb838ecc9b82b8eea1742da9fb9cbd8ca63d9f11c040e4561fb9073aca9
z353ed8a8475c5158512338b78c8ec85266c5ff5f534ed13d6498088d4a8a3b05a10588ccf167d0
za64fd911b3c34ac280408795c559864cc882d43496e2de24e9c80625128e539e72cbbc8cc57494
zbefcf59a94c2dde10fd85f98151bd88938e2f41ba65924ca7b49eb2c4895a2ff6552577a2c1b76
z5cc4f1bf48766ace8308d216e913508ea8d2fce3517d457b529c7f79fbe547e684c733d4c8d2d6
z3e32e820afc3fbcfd0e8c8a7d0fb4c4ceff71a1aaed0eebc38cfdbe1a0a1d93341fae5a1dfde1e
z812f57a07043854bfb15cc2e30b4292e60a231e0ffdeeec02fa3220617183e60ff49c98c739b86
z36e03f4aa9620192cd1354e54f5881c72a0e476ad8e472691eef4f4f4da1562564cb548ce453a0
z07a120b9ad62c81a0857b3461faf3343af4d8f0bd168de5adfe144d3974c93bf05f4cbfd30cc04
z54d5daae846ed44d2cdf652e70e76e1377ffa2cbcf099f4b2feb3c51492e68b7c64c51bfd07c2f
z27f962b760886be441600ffe4d81087a40a6c12a8a0f87a240f387b93e7ccce87a263338c11c64
zd9d1758b74d1f6edda2fed0404d3ef39ff2a4cfe4a8ee971a57032a94fc65ed803d4976f4394b0
z4b552bb850a36ccd27dd8223e5526bad4cddb0d954b05f0a15a38d2733070d9417a531a61416f2
z73cfb9f43003ae2bb40d29c21ca1bc743134bf397cd61408c96017480cc0445f6b8a05957f36c6
zca46355405dce38698dde62315dec9351b11ceeee5509d1feb270ace9043a7564210e0ebc9703c
za8c60eed328af96daeed1f159022bd59b708bd6eb34e5a1fb57e3e69949b1e447f145f6f588f35
zd5f69ef9da2dc2f476226114c7c8b4f9ca0872479a8eec2f779e37f960225b54aaa91ace27b8ab
z91280ceb37df7a081a7418d1f914bf64b40acf063e562ad969dfb65ca6aa45d4390081408eeec4
z0efd9db13e8cedb741145fc52edd47d7e89745622a1d4181c44689d2576127571d63cde04d4751
z315b5065d46b247f65aed06423e7a86b7d2b1b2f7f9878c3cce227871a2ab3eab0a8fb5ddd9c2c
z1e08d5397588e08b14437a905ee1776aa70ed8b46d584166b5f0f82d13d8ff6c5ded52b1b4edbb
z0b3e471293f8c757307f1b9140a65274211e4df4b21f338fdea4b9e29b8940a73bbdd8c5acf2d8
zba58b6590b5d09d847085b3a4d6a3c929c42b32627e88d5fac6b5225cfaa2acc38d80cf3d3aa17
z09ac082bdfc3de22587fa31d21a81c1e5c08d2debbbde42a2c15c3854ef11abe6a8579050f4a84
z684670ccde0ebef6c5ba0a52778b3ba4ead28832ad17cfb2a1cceaeda46ca1a8a9a5ca33ecf856
zeb70a8003b3df6ba38efa7bbf56d32cfd6851c20b942e56f1914771784b5a2ad3fc4b2410e5015
ze49ae1842b4f6735cde65df6d920d1b59a36d1dab89194ef14ca9d2891e007c737f4d32624e705
z69f73bdf3696c0ce5045b89122a1e7cf8a7abc57207184581de00aa2ce237e56aa417553f5a56c
z59fa48b78ba458cad161ba2bfcfd1b4bbb5461553f5533c8d4b95498902c1234a3411a8d0efcd2
z3ecb68792ba31cfc5eec11b6d244b3d782518bed5d515edacc938d978946a3f95381a9da43146f
z62f05b4b8a57559a2ae869ecc1c78ddd1ed007c4278b299c5d14e443f8f4e5ddb7832b9e62c668
z6153289c0d84ec17b30a21a878d5d0b8cc62483939befb741fa0f1dee3287ecb787934f433df17
z7c5ff2c3efb7135ffa69f195655764461ea3654aac62abe7759f2b31da635547d7371ef704ab29
zda56d9dafb6bcf1d3f4945e4aa3df91c81f53505fe3cb35e3ce2433866a8e1673802899ce7aed6
z49ceeaa17197845166b3f1848861c26d2f0b3158e40f0033b1ecedd60eca38042accb986cec743
zca5e57c7b75958068a618994bef1cea9f6ff1f3aef9e205bd4fbcfa4f837c6a37c8aa3fc5bf3fb
zf553ed85baf925f8bd5be792fed6f10020b2f49166e1c69a25e614531adf6aba70f5518e63e242
z82894b492b988bb49bef7c70cb45e9940248f9282f34b85895d27d9a1c9460aa363a4b941418f0
z57c9ef9526b1a01fae9e4f4674fcef5261f8bc970935cdc2fcffff154054caa9c65f8f6c3f3ebc
zae3728750d54800b17e6dea7b4dbaf4e8c3a6a76b6f308c46f2b3861c0ca6837a961824bc76b7e
z20f7dad38509d0b9ec3fd9dcdd288b080ee35bd05be17e8f75be0ac617706bdcc7ff4fb0a74142
zf2c977d2b8a88dfc400c9d30b6838ae15dccd0e26feb0324859bfc29e67f380a985bad1dd6a9d3
z85769ff301ed8d3e9ade031cc940365fec108d2663cf9fa4e567d850289b1efe51654fa1f4d663
z9b8dece4734a18001318a41b0c780cd4bfcb275b5c2f69285c97f82a07b40150832b04839eb61c
z24b4046e7660757b4ab538ae7c98c189dfe4c057c407ea29c7624d4d5681358931549b60912817
zf4252af6bbd5ad1ddb19878b55d16cd6a1972c5a862655666e7dce03c8b32dcddea930c4a928d4
z62ca8779bd103d6f6fe75183be9e02259954b91bc5ee314471e892f665928fc40a53729bca9beb
zf0e5edc8823b9ccb0ad769ec04944715ef73de2dc7cdcf8c0073e4e5e8fb3ed999863864f5e968
z4ace3b80eaaa8879079303b045915a22b0dfa00e27e76b1bfc8e1061d862c7edbe4d8c3b3884cf
z32b383b22caedfbbf42f7d327342b4ee393501f2d899c8a6824dc078bb3a2e7a75917654052fb2
zd0f17490ae8f530059709396157e6a5df03729716e01d5fead13b7c1666e950b54d9f2ea6f707c
z633fc84b80caaee3afcf13b80d12022a875920ff1fcd43551cdeb066ded5608b3955ad75e5ec33
zafe91efc39d2adf422b05c7df56b294915a8e06d4b1a3114f7e67b6f118cfc92c5830d31cef2d6
zaeea9692eec7bf38d892a774fca0390f23e0347a8768457a688dc6015b0429ec8dfc5523c75622
zecd3325600a2f21bcc72b9f540a9ce0d323a5ab072fdb68a7e7408e4d96ba12505ac5f37f15823
z22e7010e0033fb24f950eb3cab82e0557753dde32340454ad31a60879967e4920e41bba1f8ecf7
z53c298ec612e5e8f3186f2977aaf0237504286a97ecd1f094f2228fd9b3d56d5f9a54c5b5aff12
z0893f1e4268494613963740be90f93600b4b17b229cb44722eb796bc722166098aeee826447bd9
z41b58504348d2e1277bf34997a71519dd681bc973255443c67aa3a1346ded4aaecee8f2de12905
z427b0825766cf22451e9240b98a46cfe645b96ab33e5f48c9353e6d79db9552db340c9331089a6
z730ba47954d7608cb724758ffe0f3d74fd5dc709d505eb5c0bef804f5e270d0ea04b0ff04f8f99
zee8317daa7d90430d38769554a08b2940fee3727ff00a225781979d5e34f23d13ed17d55e41a5d
zb90ccece828a571b6fc5b831ae9a023e6d11c7ed091aa7b8a40199e3b7c095248e558ca6d5eb96
z5fc86b9afe59974cf056a6558fd2a66f654bcc685f27bffd35a33e3f3abf4b640fa119a190bbf0
zabac30c4bbf76b92667d5dc76058d7dcf8f5ed2ce15e8e89b616a45c61cfbcf1e24c1a9222b7c9
z6d33095ede93d6747b2c56a26361d5d469104b82c4c4a88db156e204d94c5903996aae0c41e147
z5d7d8806d52129a9ff90ab18db903d614028976ff0147dd30d5a3f8759dcf00218619d3604e3d6
z2e8aa04091416d485da266e3409d6cf6223d8cd1a21185e97e419a10cf8f70f0529b79667dd24c
z97480b3cc26049908e1982732bc9fd89883876b5882f5ac17bf1a827e8bb9bc03e7e8113d4586c
zfff832c73995e5447dea5e7c78ec156b1b93084e0491cc5edc792d8d2e37fe33c787bf0c1de88b
z2ed101cb9adac191e7e2560a43966ca71f9b45cbd1c725e8b45cce98a96f6d077831663765dcf5
z0fccd883dde48acee74b938150389be29a84ed3462336378e20f54e05bd6769223313734df201f
z8bd7edb028d9a6502cd230bb09bdac9de19e9a57eb6adc9a653f2e4ac1f7113e94b8b2ece9b817
z6c49683a304049801318abd0e8567ac9aaa3a862a343c9f6fcece9bc64b57b8291ee5182ea858a
z4a57c8c3663e45b186bd1ba78b6e09f0329bf4bbb230c8a53a9743c3f0a12b4fd1d715f7c425fc
z85e5901d3553dd5ffd1c566a947d788a5dacab0725f0792e6ee2a70290c5c995213cfe246d9de4
z61e6c89349644beb286b5bb5f92da416efdb8e82c6580721c6b2d5562e8dd66ab616186fafebca
z6fb165f1481b6902cbcbe614838bb4e03d34d42ac11f016e29b9b917c06e587ab20e0e793932be
zcaaec1843b72fbb057012fe1229516f7e886130599a4e1c6af3931e6b4636b5713d2db686ab0cd
z1848dadf10f6d25c682ec89f3074122434314d4d28f019b6a45b8b82fa9ebd8703cf0801e5eaf3
zbb70cce4db4a4e38164067a354df7690763ef9cdae3cbf002b1909f20143e37b2f915fa2728d3a
z469e09c8849dcb3f91d731adcab687be300b58ab0c0504540d40e025687edfdb2834a82defb92e
z3be93aa81df11ae39dcc626b67345e493d7f1de277ab64368c8d718a277931e2e0a96c59edd20b
z5595ef0fc0981cb8205aec0c4b8487e742f9af1e625af3ecfa116eac8343b34639f6290427a4d6
z5fa08073c28482112647ce5d291e5c6652777fd11418fefdb4bdf032985cbc1adee81ed85b0de2
zec16adcd3a973b90b9ac022d46b4d43963d9c5e4d7988ea6301c84672528e926ad6e6ef9878bf6
zd1061e325fdec1b31c39cd0776e4d4c5fe9fed0d957bd9095111e6d3ca47ae1a0f93cf4afa8a1c
z4289b86d480f15541a439df3441b893acc53f4b94ff0a564d7972d5d142857200015eb2c71e060
zd2fe4237ddbb5841ce0d9881fbd847ce9956323a9db3740cb7ae1779994679328db75823297aa2
z8ef0e4fdbf1d37f508892893bffc8b73988a1fae43320406897ea3481bfe1f9a8f355db3a1b2b6
z989c000eafd35495649e48e05ee7dfc1a06c6d0c785c1a64311152056754b42b33e1edd10f94f9
z8edf4fef84f739f015beebac381c17679d76c4ee94bb4f6533e03d5e960a9df4e758928f9bfeab
zdb7743b0f249c70ea974d898bbc976933f6b187a9edb0bf2108c82fa038fccaf4e285127a3aaa7
z53ceae68170f6b9302cec029c5ed440d544b8f4e8664c273296ad309fe3fd8afdf2ee616871e55
z770ca705866cac314d8242800a2cd70b13566676b52ea1b484b024dc7a40b6d1efbb6897ce4d27
zb4c15eec82a43f5a10552c5f0cf6801c1c8d12a7fc2ffe7b7606859a4214ec4719f43ad28fa113
zd9ffe581045bfb101fffc6d114dbc1640e72b0398fa00359f8403a7914b24639ecba839712c55c
z86881f8494678678e741eabb13482f453ebb8beba69ad22843a4dc42bcffe9244de633ef4d0ca1
z463853be5949fca73a118c1bcaff3da7af5f0db5623472eba50f4396a7f087f4a00de9d153db71
zbe30e9f36d0780d60dfad3e064e72655d7525c69f7f693885aa87b7f670e22c24ddf1e23e65d87
z07329931dff18b68127e306cdc9d809b7868b0d66b2201c18986a6b1a3406e973dff4b7e47706e
za0ae90eac9ea1f189fdc4370bd8023ab5f8eb9198d4ce9d45d0dfb812163487ccb7f8d48bdf990
z6d490e9660db1a3cb2b545e821f7506984f9af1141f23bb0c18afb88c9d058430e301bd6c7e379
z84731cb2d67b79f15eab527f4d3463b4cb3f8a22e8129516e5b98ea24cf822fa9cd97e63b7a4ac
z08c1b2b2bb59ba51213806f17258cfbe974e48b292b6e9b9ca59314da58afb9317f8e18c3860d5
zc2d1fe2ad582697dd8328ded28228b09bee0336a59a74ced758c8d645a955e9466edd23d737d76
z7de538792a395bb78b305864da3e91709418897e2fd2cf58894b0c991d199ab46c01749962afd3
z22234bf123c69b05123f00b503013351ab705d1105a9129e65c285c207bc61138b9871768c98f1
zc6c3a848f765f4fd570c9dee53341fe2098d80264189b192fdca129c3b0405892e868c3666d2d1
zd86f2b1655a7fe8cc8b054c856623b7afa47142db8e8b22911ec6840c921d31d713b847dde768c
ze59eb912abfcd3b25424d222cd970a99e90882abf75023123b0c5234c6592aa4ae57d3b1a5c64e
z646afbc94357736828085363145447467c47587c11d7e748ac38644b44f4b9137866ab4d41f6cc
z6de52cf7cbc6642efcd95df4383826a38d8106fa55909f8e9188b242c23a7ae9085b03852751f3
z407bc647f1ef4054ceab2f30e323a84f1d47ec2e38ee67fa23283613a16f0de6ecbe3d9794a0c3
z1292a8029048ba67c5033873aab8d25e51fd2e5783b8444a23cfc300d2b88a52d081be741be41b
ze1b5a72cb93888c300cff39dcefc273df6e775231dc5e997ee1eb0becf94891f564791689436e7
z3cf21fed1c319cf18e3ef2f342aca9280fa6ebbda4ed750ed98833541035a60d798c8bb1059f45
zeb41fcc20d70c40d09d9acfc36a6125b99d6bcc936a8b6b8296967582b462af1c505b9f99e5d5c
zba3213913171c1b8f2e27fde4755427ab07b77f2110a9555bce80e1451c89afca6c0a188648807
z97747eaac45d5e0a9e0cd7bc3e0625be37a53b58783761d1c74a78a1f016c29484a4efe0193a3b
zdc1a98d3ac38a345fb537429a6bfaecaf89db6a86db4fbfaf0b008574676ae659afdd0ecfb0618
zb73c8cb2fad8141ea30850c9ca89a0df2dfb1c5cc1c1354fbd37109eba2c1dc0ffd534a2cd94cf
zf51f2293f236be9d08903b7f4db75914c4d030c19f829ce9c51e62c6577f5139337da7428cd9c6
z040b1c77f9a61bc71292f3735b540d4fc8b50879b5058aa305ef4e7e1584da90b94f2157ff1e3a
zbfbccb4e6514557e2a14c9853c5ca1449b4823d27fa5169c418e640427c1fb88df834016018dca
z13ba2e3dea16fb52389ed52cad7795059d60e93b10f0afbec92699e4c0df483e71bb94454b039c
z939e74e4e00f4a2a122936fd76a6a12d80a3599de4f7d52e8a73ed41da664de7619001b4ffc753
za6bf4b9a12ee782b0a26cd8548d5f5d0a2395664c65b6337688820174d3a52d459dd4fef86f0da
z2ea75ca3f999008842936a077b00d13bc555178cd051bf68e44c57c82aaaa91e95f4124e4e8699
zffc942a60904115065f099b6794fa44066c590fa1babaa7c48339f93cae4fbb815b543d2b5c451
z1982ec68ca1495a39d9a18929262e82c1e8641b2cea400cc61a19e8ce1e0d1f62b3648a3b94200
z98647941c0779c74e8d7360ebd6e9da91eff4344d2da4264ee24178da75fe908a83ea0c72a1c27
za3df2490e1b56f91a6aa8f9728feb9224d49fe02aaa057512b714512646db9ea5df58279a4cbad
z4f5398f6afc7d0169b5f522ac23cad45267cde84ca8dc63aef59c947cc5674a11ed8a477627ce3
z653b158c7a3eb2037ecb0df75a41c083143f457ba8ed42199499445f7de4124997f72e7b9061ae
za329c240bee365f873078668767f8ebe9aad0240e6eabf59dab608c0cb703dfb2f5d839a5f2ce0
z33f5bbf348e57b579a3e6dcc6365d3ed1d60ae6ba76ba472b5c2190e36365e0a005f10e41084c2
zc81ffc79b3105743861e4775227f8446e32337aba208dd384f23141628b80cb44ba1e42dc83d5f
zeeddbaa0ac99409b5e72cff8bf2b42be67007baeb2356b4e747cb6d6479173f7c51b251daec0ed
z26e24f4685a912ff448d872bddd3f383969ed8898b1ed415efe0b0f5d5a7635ac6320c3bdf3896
z0c0fa7e3f965606c22b388e7e0118f1ef3e4fe647644057352db1e6eb5f749a42426ab5536ca41
z50348a610125af2bcfa06ba5a6dd91a9b9cd5bbff5476d132ff9a1faa06d22821aa4a715b0ea48
zf236626d4af31759831548cb3dce2d48be6923fac7255601a4ce1fd450101a1c69b3e3239eb9f9
z83c291f7ec58c2cbd59ec1eacba233a30741523b592666dbd4f15e3e24b78f73af58a38e4093ef
z3d19eb1725c5a0ac678567b631019cde0b90008b217833c0aac04e155a7f92d4a35d5b65f04d37
z9449225d56c0b96fd541ef9f7d8fd53ea05b72fcc1d619be345f1974786ff260cb26c1041cb9b1
zaaa5fed03c0b3b596ff353c624c9e0bef71bd54357b9673bcfcb87517842f068fa2cb76da502db
zf7737a91aace788672a1cf443ddfa28b13079645af88e5e8ea198c4e2974c451e866533bcc07cb
zb3b6487903b0373f0f04311ca8bea40a181ef183b2b942ecc88117440ad30ee16aa59c15634d92
ze96c7bbd1dea0853d6390971b26bd62ac549fcd8952615e300c7d765124b588113407cf29df8ae
z4eee29901a2536b9ac32d0f1617c48f7d91ba1f67b8c402423a4b1881edaaf72ced06bdbe3ef0b
ze206adf6fa72a51ce409ed129546d3e071c52b65d8961eaa4c3b9e870f54d249abd4d5dd7732a8
z401807ebe46ea787df3ba42ca0cd28e0d36a590368005c0c45d59c62d6462e6d5ec8bc0b0ad778
z252978c27db26cf39930984886da2b6b08001bf7ea6d93b1178819c3f7ee48c092b3b59eb1a54d
zb07e3d8a283a8672080ce833eff8a87ac158b0e522dc972cf8953fb521570dd63dac2696e1fba3
z2466c5bf0a0a81c0fdd2d55ef3d5fed6099a39f06a13681b0c9cacf132fff5d7f1aa8d4cf04cbe
z6fdfa184dd4fe806bb1f6d02cf1f7f859d618473bf1f602eee08d8b28231170e822546df9f73ab
z048decba3212df8a217d2447f5328d8effbb794d0781f144d5db185112a3a2959649f7392820a1
zdfcc4458b384108ac2899fcc85e86bcdb8d07ee3209f0b466fb7d39feb1fbd00714e26eea67e73
z4561990a00af6d02559d06341cdb725496363666d9c3fa6ba4d47aca5b0a3d1ceacee8f6f3a0bc
zb2c02505ccf923c2c49ed129546e959268c4daa70162210e1b51820da4d361662baf49bdfcd1e8
z4175f4ed95aafa2b342e95bb0029208a55b5a421ef300fc33249de8587bb776eed910397a39315
z5bd1c7efed48d38bd4fd7ce1691f6f2747bc6adc47929b85fd5f3a0aecb1501e384793fde7da31
za1325459d2bc329e30ed1d9c67af7478be309b48e5f5de7a583008e357417a6333dee05f58f525
z6ebf59dafcc87b68e13dff10a5f9f87709e7637b21656221dfd7bf12a1c289fda78ad4068b8d02
z228f3ac540e7f179046889d041738d32ab979303224fad1d4d6e347aebf3b9918632f2924433f3
z63a14e3d3a09dab46efb91a3cfad075a0b23458dbafab3874a7f1272fcd286795a1774d4cf21cc
zac370596c8bf5d67177e262fbc96f82a3ea670c8dcbf0f600cd5344ec8471c0c738dcdcfaeed4a
z0319ac95cd0f10131071ad1d0eced9d6b63eb542ac5b461cd95b8cc4ef7abe736845f54c9f9679
z4516ee4b236af5e58ea51a486ab0a28b766aaadc28790ebaca880bd60fa5aa273c76e404a610b2
z7f8ec0e480e58a669082c84c0f0c7d64907fe326730d53ed9f56b38af8868991cd35dae80541bc
z99c858a7bed5495262ae85b375b534bf085c360f73c2f44ba2c3afbe3e464ae6c75a73d1e4f22b
z22b11936c9f5dc9f234c2ea7144629acf13cc86ae62ebc73829e5e624c8675caf4dc593b2e64aa
ze6c4e47563e3c2ae5bb55a1d9af23d274e81ea54c646df6cdb0f555bfd7835265d0f593dc9f2a6
za4c4c0d0ad96cfafb71df6a43b8c7572ff37009792c89adce2b7a9df0fac07f1a85bc5e4837eab
z42379128f0fad8224c099d5ce6e6ba25a3834603fd13cfebd275ca7f5a0836358516dda727b66c
z1cdd82919436e2603b503cfe005629591dabea0054bca275a9ca58ac7172859ff18da64e6c6c7b
z37532c0fd146af1d2885b6bdcfe3d1896eafb43eed92fdf874c4d1f20f50ff678f29446a608d5a
zc04c1adb11888a498e405f1be2bda8ed0184592ec13cc772b437c59104e8f3c135c676587477a1
z074871a75628cdb8521406d58f5302025e70a847630997dc7e9323c793385468b6104597a30d1b
zc23ca0439491cd2f95b82aed500e61e0998f7ffb1096ba1db8726120207aaee48608818fd3e753
za94202f74f9d7959926e5c283327187af39859d6ffa4dcdffab16fb6984e2f3860ed1d0673b454
z636d663db16a8e5db756d88a98e41784a5e09a79f7bf64c392b065f4c5a6eab9b76a3a67929fee
z901340c0f48b68d32edb1ba3717ed4ba3ec4c353a4df603b880969769c2a8ce7e5bf1454dc401e
zf1003cb811a58e32d81f335a988118a3e218a29836f3c18c6e19dedaf756d25c6daf5e50375091
zee9fe7df04dd403f544e4aca46cd19d1a3bd9ea49d184924d8c0274fa3f1f19464e93026120eed
zc108e5bd9298bc3314721be3651da6fca9ab314b16ca1116be33a477da2678ea0ef6b0eae53dbe
z2c8c2c68df77094d1ba2225f83be4b1fff14b40a7a839fa7a03816c91aa8274307936e3f9b251c
z49b071f85dd7470948ea3c92c1f5b41c2c39178c6fdb4b90a9e4db72013cd2ae39614e84651c76
z14c680cad2dd66c2869aaff45d78017a40cc9e32165518c31e3dc5d078fb052f39433af9ed8172
zf8ee97f3c6fc2972c7f3af2c83b0a69b9b10dfc9784745f3721fbe83f7c63feb0d7abe3dcbe13c
z7f78d836c63322e69a1bb8becd6eab0ff5f6f30334a151cdb46e9cbc4baed501ac841dfd8be423
zb7d8cdc42cff9a2725b5790411515938d7f475001f0feb22b8ee36050fb4b6306413833921f019
z0c205336dd9a9df4bc6a2d47b8b5c3737f659033aa3ec29e1ca71c01f25e9c31bf16bc94997a99
z64962f37b8d0a83f6e001ee2b49fde20f504689e6ecfc89b3b14c6b8d0c8c63698714e68f2ffc4
z7f44149dc375a81523d54e1f4c29b3fec350dfe18c93d5ed3be600954e99eb4391ca079c50d2c4
z117e8998c5d408269c111fdc60f0a2e8b2f72ffbe164852a25d122c64925eaa6d4bca6182a7328
zf4aa645a439239e99c5b97a05e03010bbfdace4c244468af2577e3730fb99506f2bd2771198408
z526d2df92eb10c52ac0b3db8bfec78e5be78cdc73bf015fe8253069b59cba5f86eaeea14b309a4
z5b22415db7cae1c0176671bdc7d25b6c587ddeebbdc8096ed69065062cada085d8ac32d8814bba
zaa8f1ce6ab91a06b259808ff11c8cbf188b74c0ab892d50c8e5cf75b8a47707c8f16b4cb1e7df2
z3d3cf51f503b23edac94e8f6a39b680e157ef683890cd6d9ee95511cf338ef56606754983c9b4c
zc385b8c9f444057b7a25b1845e7791812babd614eee1e50be4fa369b1c0329cdcc59074ee19ce1
z65b04403b939cd5d7979b592036f695a0904d5e38d7e104594eec208c4cda6a4cd33799cdca04e
z39c7993b5c8838ae0f388af4e0175b832783de78fe42dded411dabbc93b37668389a2d9ee5618a
z25c24311237f905160fa6a6e8ec6abb05fcc6cc648e31cb70ed2bbe0daf38074179561e7ff0bc6
za19adf97c464f8407b06822783077be03c72a6964a2b57a82ca1abb0a5f65059048d80b949d896
z5043fb16407157c7768a8c40ae3708f397e69dcd72626a2f860fae4072692cc88ca534fb38d60c
z9affffd16cb63cccd6d08626b05616c110c65cf804309f416b370fccc41d0393c5f34a4339abec
z773b73025c3cf3415e4f173650f6cdc424701b2c1ac358c7a16777ac440d6b894e4b0ae3008216
z16322078a3160ecf867673261543354bed5ec1934457c758883748a84e08673d0fefa4d19b748a
z90d823dde8c86de53451d25cade808aa8a55c2841428ce4601ca98e7925be56ca2a71dc3a374cd
z27feb74cbc1a03d81fdb4de91e6db1ffb42c66825bf0c5c4ce5f321d4249bc86b6af3f7a7da145
z93bcece14689d8b8b9af623363aa82cdbbad6b8a142f6144ced63740b1c5552112bb600a5dcfc2
z6ef879a0cd4509e8cbd58d5a0cb569467ddf6c838bb28a719192ce4bae40c8d1d049eaa1c4eb3e
z09fb20dfe8f7b4e7928168945b74e4ad1921a0e6b22f88aedd759c92ffbd9481ab0395572edaf5
z20ea95704301978c8d1ef7635236875b73e47f224e2d24f905db8a461485f038430800b724b1a0
z667d73900a51335b92e6c7eaae639bb91bffe61ff26e3fd2a4087c86eae3a911c8c29f0de4e570
zb7ce483f9442ab9f9e2815ca394dfed0516606fa2182ea21e2f6e785fde94cb11547bf5cc4430e
z638fb4d05b83761fbd8797dd5c04fd05e55d99067bc559f0c3c5bbd5c5963028b462401ae96dd7
z1e8efe10b9f56a21d1d8e7a4766eb60e13c028a1c360c9c9b66ac523f3111a4dc0c6e675f3bce8
zacb5e229934267f74ac471ecd4c74016b0cac8cb631287143a7a5290f1c0dfcc0ad561e7ce6e39
z30b334006a52bb012094c8614305b767160589f52c0a529a8120f0738bb306e8760a43e2cd2a87
zc7aee70d3b3f011e501058a525cc36db3c13ce9261e195befb7fa6886bd90b9a4023430c2a67f7
zb670d7ca1b79535aa7b78d43517781a369a71347f2e25582b43d6a5b651d9ca6fed4a4d95b1173
z407a3f72d40e74e05f39e87bd685bd700238b9c3337ac6c25e93493c193967403caa889f96b326
z9e24eb69882972ded5fbb31e5b828092d538617af1df390d174d39c3c2fffd3432e968dab8e376
z09121a517919a094a40ce7b5b813a787527178887a7666dfc068024aeebcd38f06310e8dc7aa1e
z74de3e26300a1bd5081e145398c154d4d7b77a157f0e3d8820d75c44a953c6688852d70beedec6
z97cb5ca67720782fa933058ebecd8511be6a3d103ea454252e6c7072417ace7590296313f35540
zde4875b8cb27031ad87afab1f20513c242e891d6d947a75fa140a67a3ed34ea64698f38d8ae1d2
z4d48ac340b4a3691f211a51ee92d13a12063761e665553e040fa5481c5f9904c93a45a12b1a8f3
z6bee8576afee9bf5971ec169c8af6b473b265dda4dde1151248e7cb7e1dc623f6f7e87648b8a54
z4bbaa3949fc0a13fa2a8d6b3fdabee58b1b5eadb2f352bca0396e63d0da5eb3040abe4c9cfeda8
zc47984e33be69b1bb4c40f320390c6587d27fa3775d1b005251fbe2726ef03df6e2cdb78099c74
zf1a386213a3d5df03e5b514c95674c876bda5bba349402c778d78619e97e2a02123f1ecab4b879
z09db6f28d79147615f432c744563d61c4ee122fcf4bf21bb952a2e81ecc01f20e39119e7175f8e
zf99afdd8fc7a1d53412c6dd92405375b15efe633dbee0367e1e835ac10a80d8aedd18ad73fb20e
za07d3674569ba168b49897676c8852f15a9117c71cdcf61c8d1d57fdf24ab059d436ae83c60cde
z4a63b047c7cc40af5777fc89399a9ff830b616b941d298a8366fd344eeaec26109cc3c033d69ad
zeb499ae7ea85447a497c9a7a2b130819f443f42819b5caa2a6d5d1f1645e0824bfc09b279de76f
zd4342158c423fcfd1818a6227180285714a4bc8156a41e81119f5761d103aff09b3a206d415182
z93ec27d601bc17eb1b7e724f6bd2a7160128879406fe3c5fa1b2843ed645ffe0d065730528b062
zda31b5d09ad5385a6a5e794405dfc97ce7d6db65c779ae9affaea911ad909e1f64bd7a99f52843
z12cdd3cbd86c899b22e5acfa002328178896c1953b2f9f78a1bdf193027a7777d1846834084eb9
z33af4d9df51990877cea956664daac07c20a977d4a45abf95d20f5dd54b981b22fc40ad726b3bd
z964e32e1293a68d7090acee5afee53d905be9ef193320dd12551c4e09b6373419160cad3fd61af
z712f9e7df83bf47c9dc80adfa63cec83e10a59085aaf97a1b9f7afc8807a113efe5f08e6f9aea8
z84b52377a55ff260f7a17fa124ddfde4dbed591d4e6b394ec9503eb000704ca5674aaa16f10683
z71ed6ede1bac7871d77775b59d8f9cebd53b7eb2728324c7b73224fff4e4ea37459d3848fa4d4e
z227795196efd388717a987c3cacdcbe434b6c8e90b9af67ae4631d7165ff808f1a9225faabfedb
z0f1ca11c11c70763a9f50dd335269e2ae272987c7ea48aa8c7c4121eaf07d90a86e4322ec4f9e3
z292e274053837305176e80b68de992c6e25c504c3bac330844d3906c87deba1bcea35ffb0f47c1
z81f152dd63369cfe96aeb7902874fcfdaa45a060a09f62b778f2b1947e884fc8bfd309b5e9779f
z0df4bc4dd01571f16382cf4d99e7a35b19bea8264430db32a42ed1a694f4496997b11129c4515f
zd2ad90bfa5d3c2172c894b964cd4426850b2fecc4c7d53eda71b17f96024c1f25dd687fe04aa12
z3d3c458616296e8fc3d19c3533b1c7055bd3dcfca6948719b1dd81ede3c8dcefb64972040532b0
zc1e130e99f0ea751ea92ba5caa47644f7a2ce6fc61d6a0c1301f43b83815b9b3da36f358bb7b00
z0c456f5ca1b4ea5e3103f6056433776c468fda186de9a7825b743a7f3670c0b6521b2881dbfaf7
z11c18c9c9b9a70ea9607ef98c04027cb97bdec38e9ff0cba4f8641faec78930c0d9e36cb9a696a
zb3b90759968e2203f37b1de7c6a305963f5a208005bd2eb8c56b4dca6edba92cd43b5bbab5a688
z6df50df6afeb1ff50d1402311b8ec756ea0eecd92edc8d6d3522398437484f8985d93368ce14ef
z758cd417d14cc087927f0f2ba87cce5d443aa732a08404c3dff9fa47abdbf6d8fa504142c7aa52
z5281daa2356fc1de438a012c631d2151c635fd789142f65941d6f0968daf6dce6c3d9737f7632a
z40ba28ab92218cab166c29c52280c06c50338242a8b52413b1c896678408510ab92b7cd4bb3d24
z94330ea09f171905921733ba2e0e53436dbfb135066ad8b9d06cf88aaed0901ef964d854d6a7db
zb352fb3eca315fa26ddb22d01a8842505071609ed03a80672e59a74d67311f1e326c1a4291a5f0
zf654845a319cdc7fb028187c9697fcc32ca42e78ee4aaf7b745984a81f81f68f3095f5cea6f156
zb15ff1d895dcb724a832112159f6b588d47c52550fce7b559e93979b79ee94ea7e95bfcf7141e9
zc8821ead42c7708517d59ebacdb7be54d3eed740738c5c9b139e9f4a8c1d8b6f221615ea5c6933
z7d2e065b35ac676b0e1c7d520ea8dd1b2dacaf5157baaa41a7799785a549cb6a2310ab49001d85
z3743078c8abc23d604622fc9ae70735408f2a8ee8c72f8101451deabed8ddd6b897010d77a58cc
z6191c87242f4b040773b7eed0557e57c9246bbb5c738c693bf360d6882e1dd0a8e44b6f2123f86
z854fa122594fa4dabacad4702c812db6d9f1e2d03c517cf3c88224c4ea8905308d4bab8beae533
z1a7d5a19700bd7fd60fc8f0ba531c14de488ee3f6b2ffca0698db4012d97d111fc97bf84439305
z1d8b0c93aa21fde01d583f05417a57b959348470bc8eca6386a1c53034be32e2b87c98b1167259
ze4258c4bdaafd9e2184c0a3841dca9432e8952c4d9e459bda5af4ddd6345b14fd9736d8a041e9e
z8668e65f1bd96d227c2fe6b07593c032b404772fa254c1b37145a76c6085fb36e5d400131eb779
z1c6e9efce1c882f52187b90b108e6ecc34d3a4815b5a4a77cce66d34bffede72f8cd20bd8a524f
z59a21339835b395530bd63fdf084b3c72ccfa94b788b4178361e6d99da406a807a63d15f5f7db1
z6d93cf3fee45ed9415c70040de6890d739195bb4416a224f2d95bdd62ac040449c8b180a64b052
zb6662ebe191140e3a9dbcaba095936dfa0c180add80ef580c467f886ec75e21ed0a8c9d44cb1ee
z3dd1c0d782d376242146e786bfc58dba8cb1b49e6da3b8481036dd27cbfd777b52673e81d84c34
zb0ba03fa9d7b1b73750406668f2cbc3463d68cb407e1c3db0d8b76c0799e0642e510a199493848
z1f231df3bfa9e19e513de2380fc08c253e8464d96675fa6010fd03d57bcb1b2b4e94a548528de7
zfe21919d24f082a1dc9977640fd8420262bad023a06c7f5af7bff07fe230ff9a91000edc29bfb3
z517d649dedd737cea85662241cf24962408bc4483c111347bc3d01f74fd3c4f9ceaa15254e7211
ze863d5a9f2bb03496253d79abb3dc36626b78c72e1893df930ab001204f6c4b4879d1cc7769396
z7094d34db849eea0ae55845355fea81b59378200725673ca3e66f37aaadb83baabafb58c94fcfd
z665704d1eda82241f9af72eacbe8ca9c202502705f0221b202640df90b2d028aba35afc2186319
z636efa529088122a7525a4d8ec1f45977ad8db8c138ae9e30d4d76a353598b3a8c65480ed84a79
zaf0eadbc6a1c03838993ed45600a9436c240323301a0fa830f720c05bf0978927c158509f2b84a
z885d64abc2eaa2480cb6d100f1846f0aa4631fe97e2bdc76c3bfb64c05f22d955bd9232c8c2589
z5d938365370523057f3051cb7e3a13c4c6e86910d43fd15b0e5c9acc7ce6b390230cf384899faa
zf27663cb4b2d11a1d52d203dd9e08e54b9177a4924a7f2df0ed90c763890c3d3ea4cef21e63497
zf57b91dc5dad52fecdb03aeb58e29e3839d44c75dd0e9732fb566e98b6f59eecb151ebdf69745e
z3c3d7f34f49849d04d8fab7fb35046ab35b6260fbe0708acaf771a9f00f5b897f2ca6c817b9d26
z7a0add00a13af6b9e39728d3d4208cbc7096a5e87eedf60d2c734ff2d1f0e882885fb12cf7ab47
z071b70655300078fd3df673adeb7e66ce160c59d97752f224b950cec2408737f6ecbdcf2826049
z09e1f3f74389fdcbdbbeb36e087526a72d06ae90c14cb8faf405061e613fbca8e94590016eef61
zce362aa56d1338f90c4db4286a28a060d5b0e0a6ed70f186066db59b5a5b225a338abe58ae09b6
z71153833eb7e02fc2d4f64caa256c5d007d03c1aa9fa37a5cc73c26c394c8f55680db18457cd13
z8ebd3f8f87c7199cc8be009d8e180ee632bb73cb4f13fd60c040bad67c788494b4393fcd8295cf
z44f148ebc3ab27269027cb5fdaf97ae5354d918f6225b2c5495deb22da74fd271888bddebb1d33
z95fce9a9e7e44a278f36ca315d63ba8d1f7c045235bdea78ed3c99fb81684a00c31f97abe9ae37
z32743fabc535979d20e00a0766584ecfdcd7312e34901c37830d9d570b50819d68c70336a2f0c4
z74ad2cda9de151ee10d17ba0cda435a38a6ef2db390a185d6a1a29f64d46ab4f1110f21227ebd6
zbf932e637fcfbd5ac4f26b02ba0d2ae0c120048f94a5dc7066de02f4663f66663035ce5032991a
z03d48ad118f4be35aad8ad06bd8ec83bcb5c7ef8c937970e7b0d8ff7897e824d74144460e8ffb7
z23e3b56f34256c5b9e7d6c6121a60b6a78c1008948993ca97ca99f6ac7f60ded1243013db93e6e
z8eac95b6d7cf243d8f44a2b4dc1fbdd3b0ab2921b97cdc278d0589f3127d985393e0f1154f10ba
zeaa7a9b2c68a2c0e009308861f09f8162b6b8528affb4311615c19303dd905f29eb9cdc38bdaf0
zb402c5b525d473bc418c605f6cba677c73c0cb4f753b2190668488284bd7a3f541a2c00555bb71
z1a133d5fce91ae1321ad7ba4a784c039d19a8ecb3f08bb98dd454320fcbed7a082eb28d2f0c0f1
z0b1234e04d835d68e762bb6e455c8015cf474d898d638b65d5511c68a5718ef8fba8eb083bb9ec
z007233a204f04d29dea15920ea9761e10bd147bcd89865bc1f93c692520a5f03124aa6ac4d26ef
ze3363eb9009718012cfb56c718305842069aeb3efd4db6ff91e527df3b01207aef48d1f163e18b
z94191dfbb99c623327f030595d5e365a8aa9d54b047734466669e30ff54b4f06dd9cb5900ab019
z536f83cef7498e0bb5171b51ff4ab217eada57db27ce7d40d44c2ca4d4724807524cdd2d4e5c0f
zf1b3226ae6e2c585490c10f4ca9796914822d6dfa9a8c606a9b10192cdfa20679d264fe4115b4f
z182d97c11833767b8a1c635ca11d4d5159c6f3381f6e99f8048bb60b4ac27dff85c411bab78841
za659a0524f7656fdee8cf9749c6e74571f73d70ad68fbe4b89f0fea3117c4878a8745024561201
z69402453fe145db0dffa5addfa850a9b2061409fff53a70edb8b1b6bebc3bc945f27faa322d0da
z89e1b202e9ac0aa359a4c76efee7dec3958d876d275b3c7552b4dcbc110d7fbabc57b1b1a878a0
z0d7e01d6a640e05aec1ace526d4d43e3f4700406134f907f73e8b1da83d8ce3f5ce6491975b37d
zfe1daff94fd849ab846794c552e9513e0dc59f5081b8ffad930bf66fb4f8284349c3ef118f14d4
zeddd5acc4f593ff672cba65b7a24304d8be5b3d23ec70328d66eb5b259cbb3a87ec50c6b0c2c44
zdb9ac372a6094322e70b196a8d0aeb146a4e4565925b9073bbecc92aaa9cf98b6f15f49d2625c2
z871e7ed505cfb607b4a0147b81c4187a8752443da90cb641d8722be4c1102a1f19e3678361358d
z558ccd607cde8e09bd8aafbbac14fa7eaf059830a92a1357d57379a6f8054d65bc6f0e2d959a28
zf3991d7448c0639dd4f96e7dd0c7c5f2b2c0d5b2aae5d5e4369c8b8bafcba3949dfecf696c5dfd
z68ee2ae191606518407735f8cdb09be2f52d956ac91ea247fe02d851ff8aaff7fe0c14ada93e37
zc999b8a97e7e89025ef106661e5f55b52c6ba87b708f2d8c9be7d2ff0da3c7fc30160dfe2eb879
z4158ab0f87b045180a2021ada74e0d98996f409cb5588894f40104363dd364f0c7e3df9475849b
z27c6da5c4988e358144396d4eef27aa40ee18e7491cc4986192840ef6eac26c40ea3d972da008e
z59ee9ae25c8236d3429258108134d41e5fd0c62fed76b486afab831dbb72c24cfb910b64fc8ed3
z037d07ff35c3cdc7e7bb0b7994f1ba18f55422702de060f17f0066fcc7e648ec3ef44c91cb18e5
z44d567f19a92fcb9a088fe8e4236741b04ef22ed7d1cacc93b10b5d6459bf1dbcc1f5ad078583d
z2bc9024572015af86ea9cecd003bd430b67d5c6985f43266db2bc44eb7bde67d498e3e54c40812
z0881b84bab05f4c7e198bda5dcf018facb72b3384ad5173d0562b35d4a5bc1daebd0e1e64493c6
zfd4457b551efa26db47cb8f32dd8629f5650bdc8dcadd8e8c90565c809af06c55a3308798cf7b4
z5f730870c0a7ef50f84bc492a83d116614f947afc1ce23a26621795c18302d60de0846938d9a78
z577c587d9a73c8ed5ef8f4f77573656d34e02ca84fe51e2bddd234e9777510078eb8b69dac7b5b
z26249225c99935fa7c79fe232c8f726dc887dc7004018eb7740c4eea92e6a5974a59d53a2e8072
z145dd8512d3e59b9b07b8c9a01e12036d4aa0bd843ad6b708deb3be475e98ef588afb8da403497
z55e6e2dff69506dd1260df5eefb16ce6b376c507c5b24c2d06f1d709cbee8cd7efb2c7dabe1a79
z4c7cbd02fda744fb8ffaf9d0d5dc53196cce9b0d0bf85507d3295e42d092c5ae5dc348af44532b
zecf7884bcefe6bbb68535fa8e2004d163142a2d4d11b7e60dbaccc84b56978c5610866af77ed83
z536eb0bdc68d84e53b146eb46181b68dd1068ecf9675f2a0d3073010208dac0656fb0f097421f4
z69043af0aa00f4c3f95d7a276f881cd9c84f69c27eb8241dc792e4e8b11164031f64734ccf4433
zf0d896c767d877e06380d9a4b8c803c763e4c79c57da89379086054dadee6b793e3d92d7783827
z68a0ab0c2846ee119a46ba2cf5487994b0d75f9cde187752ba9aa524a058a56b45a31fff5f528b
z18662fa2136b525f06aacf0419b9e0fd37c01b7920fc383f9ff69550bfba63a8d371194a598345
z4ce6427e1b2f5c0941d109f28382d493012cafbeb8a90cf2b7bef059bad75a0fa4af217fadd06b
zb1b09e6a14cd0297a13847be8d4498ca3343f82dd5d553b9c190d14c89473b6c9108e0257594f2
ze3f16f6f64b46ebf26b5d052bfc1886d90825ed41e2dc59ceaf7663b6dacee0d5b371f65ed0253
z9d055fd43008a594c9569d32081724e8aa9e81870e8230f8ab54fcc932f61c5342efaf9c7c0706
z9b0194de2414a623f91f34c06a5fdd2a89d207d79621852d83ae9aa7ebb5523e1e25b9835629bb
z547c085f35f35a646f5cdbc32a11af386165702b7d42cee7b57381928c940fbdc37e72e05e8a05
ze0dda3b3d958fc55e0bb4e6b924c3a8a300a9ed50a07b0acc18bd39814c2ee1384d55accaac879
zd3d8b79f00e3be87b296c2a2aa73f9329b30a1520c33139331ceacb506310c919e20e33b880ae1
zdca2638bb7eb7e8794d0c5138fda28e79bb32903c134dba63d4facd262955695ef3cbe91991ba7
zfd6b24b794e8dfea7aaf41c1a21cd46fa9f67039caf9be5be23a69294b0c5dc76fc92210819a46
zf874f44d3fd59a281e78336bb80f9db5166749c55d23b8a0ceced9702c152cf6f998a2225eb5f3
z567bdafb10f6c9faab4d69bb4458175bea7cfcf52b20db1397221c47345e1f7fe3ebe8cd91e104
zbd75c957b358047b4b4d19d30e2c5842d00d7b83361d43b673fc76085e7ac442c7ce9b3ee8ee3a
z59f987e916bb4767f4e3b0d8773e401433f02244d6114ddee8d876012005a8447312c062a48f9a
z997f1a5424883a57b8dabdd415804bf1a45e61ffa6d7964ae3cc652d4fe627b427f2bfe04228cc
z0f001eedf73a2ac915fdc2776ba152ff29cec4a352065ceca096b762bba63bbdc0d78e63292610
z86c9e60e71f6f5b272aab24ebae0edd0f4f04ee50e2c902f6ba43ec7034a8563ef7fdca6c6f5b9
z315a0ccf7e63d8a36b66ae8a2fd66d5e61a649ad9cc1f87c2ee2340d0fbad5d70be81a3ade42c0
z8f8055ef0f62e9997f85cc66d4e8bc8ad511db27cb654850131f18460b45702f73f3db32158754
z4587aa36292415783fd11d42d807352d73b0bd9c117e3ee11887cef7417fc79016d542b40f1df5
zed99437d1294d920a7ef4eb8018bba460f0beb57f55e1d4dafee86282d6952b5f7445c1d5a3722
zfa7edf9c9fea62ce1f8a444802caac6d2756ced9ca08dd8629b6831f8401ff8c9e1afbcfaf9d8b
z542a17fb4ca383d59cb47dae83f7835a8d3228aef3cb5809ddb824a7d5c26cb6996247ad5d8b65
ze1db382644a0c7636c935f1e9e2ccf240a7dd875db4445ab64ec25b874d5a775879bca75361506
z4df5205adb6aa872dd556ec3661666e3656552b05bc3e4f8c17c843c0e63df4cfaf1bfc7301f0a
z5e98f458ea63505e5ebd330d99d2b3643ba8273126794c6aad1ad224ab0d98f7326440725c3037
z06bc591fb63cc51db7baead330897cdda8c315b18bf3358ccf317a48218e7f367b224dc52a028e
z774cc5a5331986647d3abdc1e200279868d6bf30a697721b9bd0c75f603ef5ec96114abaf94008
zd0f8f8feb0949365ed32a6b51becea5d68746934c099deeade0f4318f9979491a195050ca07100
zef8c784819d1b24ac8035bfaaa612b08d01f1dcdcaf0287dd774017f0cb2262ce0911e1afb8f8a
zdc5e1f013cce5b9d4c4758a297d8e424fb001e43ae67ccc743135e24c3eafff58247bb6b1e4fd4
z2bbb80add723cd92982f5d63911c7124818233e90359583c77b5f35fa270f58909c6c6affe0c72
zd0c7ef288e6d1bd9409f75afba9aa219ca276b91df4691ae3580dd16f3761c12e8488b47c11292
zc8053cd84cac2ca5ba700d54a6fe916d27885d1bc9b6183f0398768ddbeafbda0a450fa1448d29
z7d40847022dd20a74caeea38326530e321ff839221d280f3adb435c14ed2706423742e2095201c
zf1c802d2134c9b915da70541a5e8d4dc31d300fd1132977e461597a14db3bc591d172325b72499
z3fc8b0de45556f83ed7328ea2115a5eaf01ef8388d028f9707972001bdc81dcf663cddcb60ea30
z5d12fdc0acce4473c3edc48d0d1a9e1fce52b6bcb76dcc8c8f3894cc8f300c8b573123919f4c16
z33b280da83b7b93e001524b4a409430b98cda51e299a84f6b5ba7491c888df51e9953e11c2633a
z4358b6f55b00c0170998b68158d51b19f61306c87188aad599febc4f3fc09b14b19c0a569f9f95
z5d21997822a623d8e0797e67c327276ab50daf34d684a051a8d863f7c1ee91d931c877e6d3dcc0
zb56a97fdbbc2eb811757bb99f30edd90e64f481a824763cf719a8e04ca6b0c1d8623ea5a57978e
z47faa7f416e25ede563ccfd5d67337fc78ae880e23f487ee10414f3f307513f9b9baf2d1ccd9dd
z9503305b824582f9fba3fe12d9292285a23c256a83295b25a8435fc9e5b8a4bcb09d326e05d991
z88952b9c9ba039c3a82a1c6e5cc94e827920db982be09727b5f99496814861d4f8ed692a6927fb
z0fff81202b04634ae755617463dea745c1a88e90347b35d5339e64eecf67ce90231a2c78fa3907
z97da3028c93603427c001294d725dc0246a1e07625ebe4b441222922a1795cf20f935eafd921bf
zb7bb59265273baf9fe1cdc299fd648c43034a7b1a4e247ec59fc72118ae9e786cb01bace4f6a67
z4d892be076a44d70392dfcead2221afacae242a9d57c54d49742de56276a0c87aed7b0808dd525
z60d3b84ebfdab075164186923df57762d4cd203fee7c55f034a854b8cf2bb27c841759bd21e39c
z9019a0867be9b10267844aa82bc3a14ebe9becace5ce4a89ac2a80b71ac32af5786d3b9ca487aa
zc3e323f88a7cde272df6eb7f7dd3c7bc229b9fce3645097963782eaa76e5492c6b01c671e03c21
z0af3495274fe264922feec1e3314f3e9ebfc20c15e0340d3a865bbef67dc2f6c32c297de71c1d1
zf5564d3ffe0ee68fd37de25dadc65fcf1d32e61e65d3d35d0c2ca8201803c57addfa3f0b9a7c72
z1c23f4ae0e15b51f6a1ca4dcb227f48dd4a8aa4da266e350e640795128d7273e60268fe74c7f1c
ze552024621ef24bdd6194c51fa10496334ecda3c29ae9fd447b788c0726772822fc36b8d74b1bb
z2f3b800da09c57a85ea5eeaeebdd41bfc22145c84721c5af3a28961d4d00d1da43c31dfbde555d
z54bdfb5a75960bd3f9e22d18e30af96607f63dfc677b503fe4d62672061400c79bd1939bf4dacc
z2cc5828c848b32d419b5f63ada064ab237a3a75f7b710d6f43766731d814e4fc61292abd4341e4
zdfabb2601a72fd508ebeefb211cf904ff20f9d65b85626a6b8070f3b7572c6f7bb33fe70433db8
ze8e2280831321dc431a4fee7d6339378b8c2520490f3ec162bd1e88d042230e7686b7800572615
z305b5d7b3a9687c539b1c240e2017d85ea1a627ae0fa57e105ed96819f450204783494f55c376f
zd2d1011f0316b84931c1a26136631d8dfcc6b5b22f8b256a0853bb26fb4e44544010cbad0aba7d
zdfcd9e89ace9f37e690c15b256137a888160f0c08d05bc49fd928e138bcb7ae3ca6566a3016054
z192ee4121b5ba9f95a9c272b52a0ec73f654a8bae056861a9dd0a6d718ccd6029ce0edc51a7fe2
zd622c0d6f34226cce7101075fde63225e836a81b9e29ba9d674a4ae786200997ee794fd969756c
z76434a432a8bbdc29e250c19df4310ac8956a4dd3995371aa1beb8e516eadbec18a8874b9207bb
z0cb8c5a8961f7ec957bd798d78551af3197339869ae5791bf05fbcb50314f8fb4488760d4979ad
zd654c2c96a02c1f85ff003c79ddc277e532f29be7d022156b093a79a13348959867cfa510de8d2
z0f0c9b478eac34f3bfe648f348b31eb636788ffd5f98d1a84747025ba2fb36b498e0bf59c8ab7e
zb9f9f76c713e26deda1a080518ea81c1f85f247a4eb0f0c3f9005ad9aa1046e816f5e650131b8c
zcbaed155d750699aa8b42d1ae44cfd168058bcb04fabed58d32a71645fc985d71d845c5a5a9cf6
z28762edb60022361d9be4ad63e6bb4062cdead1664c2ae27a7b34503fcf28cb5fc2332fcd4bec1
za82bcf4035e1b4508418adc14097f3fa1fd302749da044c28be9d7b0c020cbcffdbfac476800f6
z5150bf0298a6d60cc35692565c63640fd024aaffb6ccc5176d7cf0c6bc12ddf32d19b96866f8da
z01e7e14cb6c2234ee161b9b573a9350b737813a180b2c420d83ac65cb1698dea94c91dbc406a01
zc64d4eea7c42b1063dbfbfae9e3dc320eb4eb50640ce092381683e64c1c7b8df9272acab4d92d7
zc43d28f43f6d7dc4c8783d015e8c7d5384a952af06f620289c512cda0d825d579c1b38908766a5
zeb354d805ba83e5bda53a6714a1ca145ab9022caab145e13e78f1fd470e4d6e100cd86677e4126
zf75546a63994af993af4392de80022178a45845a55351e9522c6451913380914a16ca29d66176b
zf1040eca973a877b8a72cb16c2198ddb06ecde52a82a952b43ddcb359528ab838285f16c29e9d3
z269ed3e148e84ab67dede6e9088b27c4ca88779b0c30a7245212106ed0c56271f0601ec4c9df60
z0319fd23ea7db5428ca41dcf838dc4c79e7afeaf161a9060b0dc402687cdb5d8d3528c5c2f33ab
zb6b2ddd2fddf46f42e1d6c75fa3d0e3923b3698bd26cf75e206686623aeef0a74b86acf0e8d278
z684a20529cd4764663651cfd0ad6acb2ce252a4ea5eeade2571c11903801124799c7a82557e859
zbdaa1ddcd35be5b7125cf39d276bf15c88dbdca0d79e70f0f984289430db90e5fadec5c7d6f1d6
z9eb845cd8561a33669b11113dcc3162d9854c28281ec170afbf43303f8e2ca586b34015818f517
z2c9507c3c32780bd584f6aece3677e1db0a31cf23417d824fe1aa077d6acf284991aed8dceaf9c
z0b9792445f271a450338b66a424d0f3a7eaf266b66e9f99beb3323938a43457aac7e58714b7bd2
zfa9fb2fe5588191d8cbd44307c83318bba136d5555e84475be91dd6d9a1a0cb83c05e03e34947e
z7e3acb33d3623c6f542ad6e88154a95486cf8a73b29a06da7238ffb8d09369217d5b07994d7308
z58b5736d4406b0474ef3a393e8323e6ad2f8df9602e6a80555492cbdd7f4a08b6fa11d437eca8e
zdb78232fa2092577bce0e278a2058b3d7733ed66cdc645702b42e5c3e020092bd9f64bd7db7664
ze2394a6d7a78e55ce6f95a031848f2be1d40a7728e00aa140837992f3d3738d63ea68d42e11aa2
z017cbe4eaf6babf59e40afe7c19b3be17d8e3053de096b942fa0e36cb07be57063e7312a6245d5
z5d10c742bb86f808e729a63d128e3d67914fef549cc74fa07aba90f565507c82eeb6c824e10160
z6bfd7a2a5774903424be280711ca203bddaf40359d994d91a818d83f0dcbb536267285d0133b9e
z6ce6ad48341cbf96b9b22ec1786a43eea87e8b1cde24d297f77cec152e2cff470f47f2333d16b1
zab5730357f69866e999b4e7c1e2946076001d4a564af2dac389f25050447227ccc5bd5f865c0e1
zd6235189fdef8fec2adbe2a29b15d920ab633afb30ffb08ec8562f30e04ccfe1e55112d0b230b9
ze41fab8442e040a6f9a897206a90c5d1dac981bd1b535375ef9c8ad31959083ca87988fdd3155c
z011e7152b71beee0bdb9bcf850f01605dac353be3bfca2388d7bcd44c10caad90d8c193240d230
z9ceaaa4f304bb4921a4ccd14a2b4490a1bf11123491268bc57630120938bef3d95b4cba08c77a9
z254097714e710188440a978d662742fe1f9ac35d71d16c32104fa9f4f10837c9282e991936c9dc
zc047b3d09611653e6eba37a935aa97b12a19ab13b4f35e3a89bc9e8579ffe3dc7f1508a92c537e
zb665020ddafab6fb90de6290a204079afe336794c18ad992a4cdedfd4cfb400616be0871c00fd0
z8b74bc4a4254826e0a1d71c39f4086151c480588597be5157f35ae60eead10d6264fb5a8c727e1
z75d43b2031c0c0d0812b8bd5a759a56488326a8daaf052bd35c0c7f6c888b052006863a0af805e
z0fba00b684ee920fd8f41cc3ee9f87e284b64c8ab6efe4cb9ed40175f84eb35c1c0d23bc43cb3a
z3dcd7f15f987a2646cf613a76b48d5ef6384e5ca8e3cacff5dbff111db93ec613fa2e8c53095f9
z066a743e31981dd2b112592988f8642f397c519ea81f0bd4cf0210dd514f18be12c6e77656f9f6
z69ba30b721a64a0621db37522317bff5c8ed42ddf701a578af298e4135ef355cd7bd6e0dd9d8b5
z5999c8304c0e82652ae9f4292e52b93aa7243f873639aaf2067eb29d59be977bf2fe190f03f664
z631cd1ac59d2036bd91d5f961e3f408b24114a18e449c65fa4d20728ea408279aaaece0788d8e9
zcddb47914d39b12bc29c41a90ecadda086e2edeff7c33dc90cd66ad725e2103efd3ffede280966
z7789b272db5947460daaf8163f2e66af3de0b632523550f880888abb17d4ef710d6e1e00a62b47
ze7189f13af7e35075b37d2efc41280c41ffd44074ebe54e127b3cc0865db12112ec9cccf257667
zaf35291f0d35b4e1cf8bf503e732e5f5033efc74f488a82b400a0c1cd8f2fc5b66a061d93b7d99
z18bd5d9ba889de94634c52020b046f559e9e49381999935439cac1ab33f7828ec6eaa6ac5ce25f
z3d346ba695f2875bf2191c384bce58106df35cb922be7e99530911bd9d17828ee53d54f123836f
z4cb6a2cd3363d395cc94dc07bbf16cd7e2a43c9f9fdb1dfbac3ab360942b21ac9923bc10c019ed
za38df31bd17032aeb3a22073dca5709aca614cdcedb1e8b6a11ff021ad3e84f09329ebcf435d12
z1c8fa66b131fb8f96ccdfcb9673f5a5aedc745bcea465bec3ae73989823d91dfd50c4ed71e1669
z78f6fe33748a367b8d9f54b2b5106567fc69549bdfb88b2ae570a0a6f66021ac596414372348a0
z195051d903163a8645bdb76d304b7014b36fa77495d3c22aeea897fe9deb326fbed726a0e3a8d8
z72a364dbc4807e7c7b3a4e6fc9ad2446c4a1f30831230b079c0eb489889e7f1e1e602f2e19ca17
zca728c1d1dfd0930b6bcad0317f8938567ed52e1dbe7842acc60a2bdde68b50725c67ee1662bd3
zad07c702af0aa40056e07a5d75dc99b3ca83506387397bf6d35a75a707c6e9a012f61b0691b352
zd8c0450c3fdeabf01e3496dddf65792a6e9b68bb17072e505baf64bdf522abf7b067c38af5c353
zcb91adb358ee304fd81336828af97037be09eccbca16309edfc765188a9d0e0d89a56988277ae5
z3c8b913131f4a99b589490cfb006c54c7da55d5963dd79ba419a1320957e7237142190f1c05373
z1c47625e18e4d3cd771ffc9590da4802b537978ac5e7f1b8aa670d534f191a3cc3eb314ae46330
zf74eee3e999b1a04bcfa2dccc75d38f13468d69b53f12e21fbcc1dd9adbed9b349e65e693286f4
z206e04e6bc0ccc211d72bfd9d6efbd3365b3eda4fde1e6483022dfde5639741a86175d2643026d
z7094e4726cc962caf12e2730d7971f3f73bbb7ed350a983a4af87dc1278520215e18e3657da691
z0e59422091ddadcd92fb350c503dfe8b5360fed3c9774a962bead097b83e77a6e766d83eb578ec
z1d7fae06094a770403af2cde8c5c834d0b7267371e4483f618aeb505899fa807c3a0e9c00b4537
zf7763d374918e97c16c5602aec721be0c2c42d2654b224860148935a764d22c8d55073e53cdc0d
zb9875976469c284fc06ee0b59a99c2eaab333eec22f19b13f50e095c43f0acf694ef1c7842b36b
zae1185805ed7c5d7c8981aa7f68fedef6e271fbccc8f70109322da03030e2676b6036030f6333a
z390eff32582e520e7d1a928f9465fcc0a9b297460f2ea84d88f8b401d9eb102523f079c756f32e
z208f1e6e928560947bf7b404e2c046dd3d13563e4de6ed3a6e0c6bdaa77c8034ae81d0bc5f7669
z78316822bdb1478cfe55591a759d7da1ce42bb77e4f6d048d0f5ea7dd2447714cbbaec7399e948
z6fa1b816dd5ea98ca6cb17346d7124cd66539c36d3a7e5015bbf5bca50e928060b8bb2946d369b
z23c94bfbe183636956ca62e83a47c064f7cde1dbd947c10971a121dae464147a5b5e46bcdd7b3f
z396c53a5738babb39db2dc467c6de0fd2cbb28f30275ab07db9de6fac180d3417e8384137af15f
z8bb1e5a72dd4f3e8e0ed8581fa376398a5a9105863f1ac7b0f30374ce0ada8237d6162b50f9431
zbf11d3b7d4324e14d5377e38904a1b580d87351097ca0551c984d1bca6cb42810bdba95e37a35b
zbab7825093858c76d6b930b29091f7dd5c9972c861f820f4a223eaa899730b55a10545302bd083
zac89b59cb6485a1ed504c86a4c70a1e0a8796eb9717cfdf2892ada97a737521ec99bb7215e3580
z7093f26a67be154ecd6656c01fcaf91792b05198dbb1316a3a1a40b09ddc792054da23667a3b53
z5aee7a961167d8836aa67b92d980b25a64e9898cf6fcae45ce7d4c57e2b4158fbb25b976b442f8
zd347682f8a6f543d13a5612dade4be676b3e25df45f0aab441ecd6dac8841d24aa1bd2b07df0f9
zb448ec17e5ed318df43137a50b4189f275f4d381f32c87756791199aedfcd4f5f0d8e81e899b54
z9d488a0d3eaac31f69e01db9ad77c5df58410de54e68dc5dcb4f922c76dd8d19ad026d6fbaefa1
z0c295258efec5136e1dfdcc901636657d1736fda96f156c6d9f5ec7de80a9ed990bcaf3dd94c8a
z114bd3f92f3f3a52078a96f40735c3c8800c81d3ff6fb3609314e3f8eeffd613bf2aa52e4b6dbe
z14ce74364202ae2f0363222469141476a7f94b33a5424b78b23bd59bcf8fadfee32559bb243f18
z80440d494adc152b2889368cd00e6bf5d45dc44469ac674a6750f6e6083992fcd4bf9074e6b7cf
z4c42dd2495b989f2867fd370d32a383cd8b83375e959776e9712e143a1a650c760dda089f6fa29
z9ac93fd077a7ee4b68d63d5cf368ed49a85053c9f58abd9a08123f55eb75092475ecd3a99e7ab6
zb554e13945e96f56e488cf8e7752fba7d169059e1be262a9f74800c8ff77df5dd1777ab6f1e96b
zb27580ba8f36e674bcd0435c6e8878d85485a8d9bd9e3e2bfeeae53d3ddc26eb3355d2a03ac521
z4a1359f24e940ef45dc0a45dd552880e0190746639fca30d9457c948c95269c6e6264ce9b3a888
zbcf4dd62565bec780cee57e5dfb8d4a35a2977bf265d9bdaaa83c309e86e2a5fbb4d14acdb7b4e
ze276894fb23837066b88f7e9f41df2d667af5348a20543d00ff836f77102bae9a31add9eeb865f
zbf003ce7f5b5807521725faf6dc185ce0c1c47369f9afba9b38233a0e1bd9fea597f80c06007c0
z1e6377c477bd8f57d30bbfeb3cec6e3d1a9a59bdd3d91269092fde0effdf9e177e0b1be1131fae
z5a48077f4fe46f0afd088dd64f66a8c03fb5861f120eacc07c103d9e266345ed8435a912b04468
z5c3e49e2ff5a1e15deeb99e3ad1bcd443082152a911ba7e90b82138a5376fbbd844ca166314ca3
z9f9340120acec00e1eb5ae7eee40605847f297fed7486288eb07961e5775951d6c1db4bbb81845
zfc631547273126aad009ea7b0bbf5c69e0fa49096c847e572f73e793767fbe7df55c7fb348d5bf
z82c5123f09d8987c2ff5a55ab8bd072077adf1f0efbedc6cd0c8a34985ddb837d1d70c8971c4a6
zf9ec7610b2d81b884c5382e2d2ecd071e518718763b3cbfa99219addb2d366f47e2806b1743154
zb6c04ac87298969fee9820f978be03c17ccd413ec11b3790ee5c78431136a12200981fc9dd2771
ze79ff14e6b331bbf86f1dffe5812d5bdffc888a6790906db1ae3aaa908fb46de4b85e4173a247d
z0795199c04a1657def81b839393f59dff9f8a3fd02532e1d446af19564e37072763e2978e710c9
z63a73b9faa373954618e523c1f54d80b7377031d9df323a160897ccfab2c7a9a610cc6e57beb23
zbe70d35b0b3ab94ebef962929fbaaab294106456ba4aa35528dcdbc37739943846262544aa86ef
zcf4e0319a47c149345c25e8952da02bec575d3a3ec2aa19c974e67734c3d311251ae0b4028d9af
ze2b4cc33141acb5cc7be2d59cd15f2355d4b04ee71c0f89000778cc56db2132afde0c08e78a991
za45753d4a6f737b265bcf93f2489c2583116cb1c06e83f13bb63d622ff69d96089cbd4312787c1
z68e5c4015c28a9df4eef1e0eebeff1f05614cb35958a846fa99a4f48bddfcbefd00297dd9012cf
zd34633013fd491bd990c8729850e60de179ca6a788592a6f86964b27401018447a7afbe3e640ef
zc71dd5dcbde0e637947a018f100746a4f9e80f44b328eae4f3bc0f88cf851d2d867600d3a10673
z2d84766b85dc9c0fb0028717f5077d8ae0744025d0b6d2f006311690a5de86ccf1724e601f11d6
zf3bdc6a698e7a563047c4ed020fb5c64b1cfc8e9ee1d976e070cac9baa70eecbbaedbd5404e29b
z9da5d1b2831fe33273e64e3eada3f2e2d102f85182e3b96ffb546407e575a95e0be222a56a69b5
z026656cfd73c4f8b1aeaf05d515b67ebe099763f494a5cfcba1595c4bdda0511d07a9b1efe96d6
zea03f22a4de6156f03a98135d9346abf6bc661e3580128d6bdeee9182fdb67f6a214a7356b0208
z9518ef07d29f19dfde176cdec22e92239212ca06f3f3ee47403ce13c316d89cd0b8f12bde6e7b8
za1e809b7518befe7b2350638830f6f03730091dd1cbbf9c79cbf6f418fc7435293eb27136ae0da
z2ac94df02c7e554cd199ec68d83af9e2f443a76c6c8d8e081a834e5dd4f83928cb2a7ef211918c
z564370535a078004ce5379896317d88b5d112fc09f452bc40ef69aa61fcbdd02a231ecae147d86
z1167111f96087b81867df32cb3adf65a5ab4498b632cc6356a1b6ca73a42085b0f5a213806b89d
z485c8975bd289a0cb6e5b0e682afa87699c1d81709d77b2a9050b257d2d1d21a18fa16bcb4a27f
z07cf179a36ddd4900651bc62d656b2e167db9e32c1c60e1b1470fc541835919c4eba64736fe617
z9699e8604467517a5558b266fdd5fec87c20f9f9c4452228210224bcefced913a998175037a3eb
z8389011c54b620028c834ad1452f91de5a98ff33dee0bad470033839a20b7e2b7080e23764e8dd
ze55864bd753ca468740f9d803b9a8175be9a8659465815e7a13b70395c8a2243becc2dcaef9ccd
zedfc5cd6e92760ab09df5c16f78a4b2de6e6096a4458a6fd255ba0f29cff48a1f23ec538b0c059
z866a6fb90636c79432e782066e4cfd92680630dd1e05a10617542288b2abf907dac3e44dd464c0
z176b52a24847f4985bb8563d5eca0f4186b79db51b2469d18f11fcf350d40b5c219f7a385a7443
zed1cf2a7c1412c524860461829f44e2d60b8574759df212e23753187180095a76b919f339416f6
zb15ab661cda18acaadd6e993b0849d0b2676342528a8dfb4b5752a0c2a0e31b31cb245ce75bf73
z435a8e30e8bde08ca128bd9e8f0ff6d928dfe0c7622af55fe84b1766521d8367a2257eda7783ff
z708eaca81f145be85defb63674371b24569b5ef289f2d353c22ac3b0619fe4a3ab68ece965ca1d
za39968a7b32c97c4a0d57c3e456f0d3075033270fe5b2d818caaf8870212d5fd89330ce6f49629
z3acd6d1d7fc573bd429d64960a6e015bdd8502c18f3d4ec35044a606dfc49f9a7bdbddd23d9e46
z4a46bd81305f267005bd13e2d3784795b4126553b12a35c6b3261079caaf5f701d4b122163b427
z0cf09a54e153200e2b275530f9393a8f1b292424af9ff53e681ae712acb16bbb7ce0b38cb7d3df
z45704fb310b1fb9deec5cf572ec6f2d953db3f18f225a6f822a158814183a5543458d9429f1c7d
zf4e7b01b6ad21c5caed45d6735ff5a5fd8ba1f96b89be6fbe94b7e792d293b0eab0cbd30e4291f
ze2bb13ca8fb3582128d29ad3f71c51b3eb73cae13c8ecc6f58517a5bbf8604f6784bacffd77aa3
ze735eb5301c6df883232744ffdca1870d3dc68a9585c0d1cfab5751f0aa74c8812f0f126ed63e7
z9fcb1d96a5bfbfb58e5822501d1fbfe7deda47c9741b1e69fe76292c05bb2e989e8178d247f3af
z664bb51ea69fd4107785dd485f0f914984a1c659f8f4b9ba2500118114cdaf585277c55a78d8fc
z216f21eaa88f108a2340cb70bf7bef757077e63c0e38432521917fd77dd0506d87d84e134134e1
z0dd02f61e9e073341b57052dc65f07c108014cd01648419bee4fb97719602f7ae7cf043f5444b5
z6f3bc5283f6645d2031c1c9b031ccfcf90525450a0ac5a95f11462893ce759733686de6f5018ba
z3360fed47648439663094d88c7ef4161fcd457b9cf0c24b181bbaf47c6419ffa6f1f84e996c261
z52e37dbb5a8a6dcfc649b8949cc433943b0ca6dea754d5aafbbc92e725bfcdfb321d75faed9ba7
zb3af322e8b12b0dfa9f12925af4677538027a526138ce4715a4a4afdddf5796d7046377bfb7b28
zf5b683be1502c7c5b19386c6818af7ea8210401608f90e3d910ceeb75db8417f45b1b57b638836
z6414a4002156b0f57ca9947ad9609b2f9a75c008ba4af04972500df1f20e2141846a5826228cff
za28ddc41e2a10742851498e074be74634152cfbc4e85bcb2da64627d1542760183cba8c53ceb4a
z30b701692d5c3ac74454c23c6c193922a3f79489953dcc454d16b8229de0f5be175342638f60e6
z90bbe8c8e01ff09aaefefb7951d2b65058cbdb0e09891cd0413e4e2c6cc7780b50f6ce8f28d684
za4bac43d56443633d64ec3515874c420db565a7c5ae698ce9033c083a409d3a12fc19ea6e04a5c
z1ce3767cb329d16a0f975316577b7efb42f156261e1692b3abae96d0ada199e9721979e119f2ee
z79a2f733d4b133435d485a6779abc61299b0501810a913cc8b2f77c6cc6a08471fc1e88ee9b1de
zd3b0f21be96deef8ffe3296eaeae3e77dff3e0d844e9d66942407e289a943f820d325bd4733f1a
z4f34772a761396276388afcfc07a5d3557bdeb450bf8a8e6a24a8839e12c59e934a4efa4af0db5
zb8d50401d90df603a9fc6ff105006bce0a9dcff6e29a610a00b482610d9be8b890300ea8c8004f
zb20461ab5ff994355851928fedcc4da4f7c2c2fca06d63713acec9a65c493b40cb87b45cd3c492
zff47f17414c57a7ebe70807b9b93cd8fab2f4bba8253d4feef1b0fc81a2a3d9a9e1ea2cdb008d6
ze71b82b95ef16d396bc715b2bc0e2d334aa614d30fb39a7a04c883672d16a193c4e26748caef65
zf9d18ddd4909b9674ecce998a97671684cd0ba840a4a9c89642005c8ef642f0fb392ed434cd0ea
zf37ffdead981322445727cc6a7aa0f1fcfcb6e5e63e7f7aab7e6b4e5ab4d86ea5eb8ca3028a7c4
z9e131beae5d7c360166e6d1832fbe99d2fb4961435a0204d12a01eb901c6a68ae88e50909a0886
z731c6a43f666e36ed671aef39ab81d63e6214586d9843583f85aef9330fd421095028954b0e47e
z643f53e3fe012ee3d4b6b3bdee68ad237ff18984bbe50e36063d4e390da161b88f6df882fc5e22
zeab40ab0fb98ea7021119e5a3f29c3b4fa4a0881214a0f3037142f7eef5f9db49ee0f4b52ff7da
z50ab0edbd0f1a903fdcbf99b4a50857442c396c9bb0aecf2c0d8fe3afa59e48a17f19b8c507d15
z4cebba5799138b2b0cbd0981ddf746af7b599f16e28d1e064c01a5e43eb4b5bc90368ccee0063b
zdd44db2167b474d278ee9d5041b29a178a49fab5a503bbb0a76f771e65a0130be51d0528ce7edd
zdb6003cdebaa68147451e995f239632ef3d7d9c2c1533985071ae02a5525d27ef044fe5f38c249
zde7467f5ac8037ab75fdc63d350eeb7f63a560dc875e398ee7e660f2adc890f7d8543cc9480af1
za7638f84cf0c94b333bbc816b734c0d5b8cce91c78f75a9ee430e55c6472980e00669a297a0f06
zeaa30eee86b1e42e5b55375561b2ce410cde41228802bc2f50fd0a7c6a42967c6cf99d89a31597
z58c1cdbf0a1f853c6ad8bb46cde0c60094773fd79a83b39605c07d5330a1a1e03fa95bc89e009e
z3e9f20158be3411c769e3a951d5eea2dfa4a02a4b8dbd36223fc56a1554e24d0d19b2e78862502
z581761e55bfbd7a98879b747ea72cc81216f6c957cd4c02223bd5eec2991718077ce6cb4d172e5
ze225b06c17993798e4548c144c0e385ad162fe1dca6d58eabcabef52cf29524c046ea800ee91f9
z4c0aea1745551bff77e4b85b0d397775beb464553d7029981c8c40968047518486b28014bf3f64
zadfbdd9fd2332cf048918366df6b186689dd1daceb3fe46d6117b91b9b5e51d703703be51131a4
za420fa126e5b9fb5b5ac2fa64f277d3ba9bb5208baa1bf2eda7bf8e6e3dd88867e54e6547bd779
zfde792138db6276a411af2e3f44039cd10380855d727c4cbcd260dfdca9c1db36d25098276003c
zce8ad3892ed0330e006f8da01de2c5a5a957ccdd22c83659c8d90a729e3f1ab53fa2be53f8f255
z1ee35b2f64306ef7105bf4fe132bbd85394a1802e79277028342d798cd892c09d1f7a09c59aacf
z2ec17191c5e274bf195c8d5238cf815677ef76710757b968646b1bf2e110ba124b3360bdd68dda
z275d835699705ba392fd4b91908a5a98aa31f10580bcf2b01f3fc25649d07bffa1df04c0c1e39f
z4bce733fcc63949e600b04eb901716969648212d0a112b9300c7c3caeeeb6be5c9f9f8b18e1b29
z3bec5fa627d35cb8674648baebeee2f7dc04c35f963a7fae6045c2ffa13ef385bc828b07e5751c
z8ffe28401a673fbef35f6cebd1b56b1833bd7ecd0fd446c3bb2a408df134f697db76a459e3a0b1
zdba8e9a67cd9794b4fccc3dbfdd1f624dc4ca772653ccfa2be955043bb55535093ae0bd0aec80d
z0d9706432eb16e5f369b5b0e6fb15cfd3bc81c50faa298c4c32f56f8298143279b8d60dd59548e
zd48e66c7495574c22d3ad232842bf6815dd1c3c522350e5faf8d1c48b1f788f1549929318898aa
z9997c81591fd10187a6e21b3d8c81f15102d49d062c7ccda35baee70a219a6e8b1ac0d9a771ba3
ze38aa8e04160b027ea39bd586374f13c6b5e5fc1aa8d9a94f54e190e07141d0f2e948935228434
zadb342a1d1725193ea260509da662eb27eae9798bfa375e5cc75ae9d1b327101afe2a4b4058075
z6528ad3c25d8c04392f89a1e72c3b6a4cd614837b38433e5b6296b4f3a6cbe2430a3b48db2938d
z1bfa0a92627ff3de4b85112465316855cbf068ad468b0658d54cf8ea4bb202a8bedd694fb69d00
zc0a53799949d02914da0a321fb7cc3cec584e9820edcb53c72d1ed3eca21f29879568d6fcf1afd
z2b1e3a594710003d7fe05ba418126482eabf736fb795dc10744b2e8de776ae49f37ae132b9444d
z7d1961514f29a0c976e2c11bd6c0639c0d6cb263c70afb92f5e0881c57f4b44cfd7f62b136f18b
za7aef5650c09df68b4776de7db60e95226fd58d4e5036efdf960223e106212502dde61d5a111f7
z2def0b7123a7865f070a28f684326de685377b73d2ac6ceca3ffc2f3184aad3b0ea3dc83234942
zdf76039914cbfc8789c57cb987aa49f8d369544544d585375c7e4dd293af8b5d04bd73e208826a
zce273c9339e9caa9c2a952c431468edd2c4ce309c43082d1bd33e014223e32d41083b78fe18e88
ze032974029e2b98550245d061556ed695f309264b32daaa6d810cc6a8d6cb3df29c439046e1bfe
z535bbedd2d9e6b3bda269dd52c857d4948edc4f8ffa68e8d71937477819c8620f5c56c8cfb8a10
z9465648604d63211cfdbfe3c0027e57ba9a3c9b7066753c25bfae3e5b6d7b6b6299c34cbde3225
z6d4e5383a0d092f2a6fc38da5b7de3b9208dfcf3c99ad2b7b1d7eddd1527ba3ef59ee6dfd3c63e
z05408212ce2a6571c1a95952774af24bb67bbcc19795b1a1ddce00738e4d7b59c3efbc2a80982d
z65fd30252add3814c540d63564ad548dc6c82034ae0b50c81fe7d4d6cde923544b8c25f2b00a60
zc586b284cd3ceeeb1dda28230f5ea02577a6de362c6d74d58a5ad6de6e840f7dee2c24d2781080
z17d2859c867e367e0e0ba3f63eb436c32944b861e9ee953e5e22e5046fe9be5f374d57738acdda
z9ea307dae0c2c9d74c9123cf8f6e1d910ebead32ddac4aeaeee996691c16523b412c1f1d4431d7
z34db38d0a90f0651227fdb2eca2253e068c80e10c3eab5be7359d210163c03cbca76687d0e1e5f
z0d5d80b6aebf0ca0b03c9f5aa9bcf03f0a7e820e537b34badc8991c42534bcb189361bf0d144ae
z812566ef198ac15748a8be45bfc7428fea36cee2e21a34d6715c6caaedc6fec35d2ab7dbad99b7
zaad4155fe8f69f02254b5c5a6c2dcb8da8e43dc63d6128561e46d5b900ae30bba1eccce489c5bd
z7bf7c6b74bd92ffc6ae5640fb9ec917bd2f294699f96a6ee9125304293814454459f00233adfaa
z93b1263928fed4e8df77422bbc16c638a26b04e3d89bd4db2a358d073e7e3c5da4a8a4318a9f43
zc1068f97a8bb694f70a5d99183215991108680742863a8ad162b22103e064f6d712b2932533580
z9fa527b4b65138835231344dfaf78b5b5e51eb0eaf54524418575b34397ce2eba6398042da7991
z0800fd6979929c85119221185d4150e4d6b58e182e8da30eea84dc1c88832fbc60408b2df63894
z53adbb0ad2869b80268b7e87f2a591f292288efd493e3bd812262bc106bb35c57f1967ba089f8a
z78602431a6faf625ecf383f7235a1370369aa4eeebec3e92e793382546c5a1bd86db5db8f28fc5
z94639491e29563a16ee7e33517fb7629ad3e7eb2caf6031e92281b6866d9a836fe52c5329d5ea3
z412db1173c7c9579d06e024cb15696bb89dfe390e3b2ec953ba11b6471eb284923f2cd7eb2d21a
z81afdde673ea8d1ab8bf735b0bf597c923ccb8c6c5462ad8754846cacc0055cbc9ac54e2eb3e35
za6fc408a06bbc2ad9c74293ba141d89420ab545fa25ea6d8aeefa625bd01aa48be59cd10e99a83
z1ed201d996b610f8c13fb4795e98bb7e7d5c960b439b27f35699f472a72f0e764a05e8298d3592
z25458251c0f125e41453061f31972525f87124f0d47766b7493776b7057aeeedfe60915b8254d5
z8dd0db7ca11e31beccc83faf21353f4ff1bc1ba5a7f0a5b724c425b7dc5b86fafcce4f12aee8bf
ze98475ce94eb194e7b5226d05c08035f94aa2d254a717c9204f1cfd26b25607837545892822d18
zddb8e403403b4de4c52599d39cd095d70fd20f7c94fd1bec168f6698750e6af82284a7887bfb77
zd3f99a6c0f94a473635034676861329a356f155c4a301f6b1917a6abf29d9bdbd39583345d61af
z60cfc52fcd6eb613959a5f9a23391419929c299ca80f81037062b420c4ec364b792b0229894159
z742933f6c2e269b17ec91c5a15e0675a946a306265d85ea5e2dfb349fea9ba01ea625aa9474eab
zabbb9c913ddbab4fff50bd5b8d4d1812c4b15573ec7c907818acae7983c7c7cdd579fcb7daa05a
zec373885a230fa0f097a79d771345f7d0d7895d417c80061615e54c38e35da210f2bbb6a4ead7e
z89b26b08381e017a737979de1d990bb676d308d99feab4d3c517633f07b28ac67f31c1984b214a
z4efa19730c7e44ec18fa1d991156d009e1a104846b36e7427b5216545bd7dfc275cb17610fb642
z8d433c573e9cad1b6102e9d16b89f51eea0340986c1937b28a7ab3cb5fa6ea42033f65e3fb27d7
z0b7f7a2b432e1c1f8a0de83bdb4f46de74b71e59842ae218fee6dd579ee53e59bb2cef154e3329
zf95e5ed3c04aa9763d1716c57faa5aed802ffa51a74c2a16a76aabd221feca953b59cd59cb882e
z53aa8a2650b0bf152a604b8ae9030e9fcd8aee2f531b3eb43f24dac6ea7611b8a3f31572f02c70
z05f1a7d337d31fbf9f4734447a9c82ad754cfeb6115bf4fbce5d11c445e9ff56cb7278e8460835
z87730a2967095f2249830fe99ed71c8d3b7464a50515a04ed1c71634f82a394ea1c73c993b472d
zedc97621fb1e16ab7526b22ba54488965c9559df66c9b992c860505d4febbde32e097a64ed9856
z9437aa3ea4d606d64510c8308e2bdc4b878d7261b9b5772eb477f83f59401158178c26436386d1
za7c7ed617cd751e5f93ff47f36730b8622543e1b0559d9da4573371258594b3d08072ce39ad34f
z08b7112e75faa52b62dc7c8574f7f997aa240e658de76fb0eb72387f30fe5fa0517e333141b304
z57608d739805ce8e15cb3c3b16f2823b49b3b8a25414cb1d41396b24de30cba54384be75ce2e8b
zf2c7be4c152c3a73a199f7544f18d8f23d79143b8801d5b6128eec5867ee78d1c40672d7ae6f10
zff3d8ded96c5141efbcc699c41037179c0c3a100cc7ea23e3c54ea7a87bea428aa482228b9e7c1
z5fb6431a235ffcb354bb96eec7c526eff04c13143ec27fc8fa83965f787c09abe131c4953a7be9
z7292975b0e1fc44517cca006a3b8eca6cbcfa6812df09d61136acaa055f59a476918159a1b931b
zd58d111ffd32b5914e88df95ad53c653860812f5bdfc43cb1b7cad33b376d5874ebd55bbc3297a
zb103cc8c8e1d47ac108ec7425a42e29a659edc2d6e5762f39976b1f2c7f8d3763040d5fc2b0c88
z2847fe50da5ae5cb4b182923352ab6509340ae3c759de5949e89ed34d9c42f1a2606261cc3bd88
z210d2be67b43a3221c2aebda0ae25b117f4e948fe09ac4ca2fe12792734195172b9426857c6aa9
zc85a9cc6d719ec8403a9f4c85d043dfc24b2fa2045c8ed44d6ca75a3ee6512582e8d53e25d54c0
zd7ce096ca0719918171ab99e5da77daf7af0b07b99090a129c8a6b5a4eed6d7ac7389b6a6f721a
za3bdd11159c7f9d244fbff80232d3df46e97f135e1de05d1751b1ddc4fe2bf226080fa9beb52f9
zd4aca9c5fe9792b947d4b33f3dcc5a5b57793c3b159272117b5e4c10471153e8d33111bde8f585
z377560688892deffe02eebffe8b227fa7a50ebf5e7fbea200195558f194119b542079b52225dcb
z350b2216d3dc87be50dbd3cc0c767509539801d1953942e759e3b8b96c32d1e4678106599b2a43
z0016294d4284efca43f52e02aba9eb45d1ddc726d9052b718e926cc9166905988e8ede37b91343
z8292515328660c1ddf2f7845a1484644a38d2009af8aada0e3185094dcce46c4aa512b27934b49
z47cde2ba3b762efa5f91a1fd11c4c3d322939f9cba40903c73a8999800f953b76e6295c381cd23
zf717f1c3cf7350cd7b058fc1d2ed7720f10b69d6440281d13671460d2815d5b75d79fe1ec5c855
z45e32b24a9a277b5c7ed7a8fa4af3898a573c1e7456fc402d38a2d7a4412c7fad46bf0e4143e43
z0caf9145b9aa60115f4ad7d9a87a3f68d9f6be59446c20f071ff2cb6481defd62f339c48157764
z0b5b52d2bf8d460eb73f645e989a8ddfd763a69ff32b393f7ecf5108b912e5b371ee613695c118
z32d250a3de62dfc23f48f632ff616da6237bc3f78b51094fda76d4209e24416ae3e59bb2d4ba65
z8a473a87815d6360c6a634f3d0ed885d4b4b34b18e76590c1f1fb7ae4570a3b66258c2553c894a
z1ad93623e0ec79da612b1c288d298ef99a41d8002655ac51c3fe4a7579aab36cdfd83a8c268cf3
z0e41b0704aadef04f5a9a26d8c29b774470d86d617248f14774ab8168bc7d9cf2c952e2cefc7b6
z82c85d3c528dd0373890e716bbe0b7e26b7d1c6322df3c50ce3217c9298335ecc26f2be926ca07
zf892f4dedfc65b31aee024cb2ce88cc7117f5e980dd067ad954f6cc60dadf21668cf0902b59abe
ze9609ca44115214d60dab0ee34a65a770989bfc7518ea10566c310bddda4b02dd378e33c991507
z4ea40ebf0cd0af2b3ee0021ffac2d77e02299c55ede18be2715d45ca2e4b71162c428be9679ce7
zde78ffdf3bd33a6035a626626203f5466736e6b0a0fde2bdfaf336879bb63bb2a3b94a787964a5
z2740766f9c33680661092cba4eb70cb38173516970ab423eb5561874b0487559fc846f7564a170
z06eab40660920a5bcd5752a3bbfe0e33b41960e3de0b10e0d5e8bc39f37ea805a4d98c85b9e970
zdea6fd95206009a9564ffd2c24f747757453cad897f23139c377694aafefe0f44d7eddd7202234
z2cc7737192d26913c095d9bf42835a64c3494568755c594553f1825841ad92fc7d1f5f348d6807
z0c33aef52dedd3db4295e773821b56a90795829668a3382e7ff065e09cc840592d8d6f18ccbe0d
zbac2991284328024b88bc27186f9880d009eb26a6bce94122794114da671d68e5eb5635e320267
z31085e30f2b59fb0b71a8f42490606a3f3d886270e29fa6c7edb2107993f2dbc04b02d84fd89bd
z94ef3a8a95c39f3e0f1f2b32930b3d088e9a0cf9f17d540b87b352b3082fb411f6f3791c505901
z1917def1f0d7707af7d4ba5261a9949bf83f9b53c5b5b513e9ae57a8c0a71656a9b2eea8394550
z1070816f1bb55a150f0ad280ce9f755600ea822396de95f38baebe0f571a249474a0a62f5d0c22
z38ffe4d3465f3881189d092eee225d8efa52e06cb488ba3ee7702f380e0bd6ec8abe8efedcb174
zd8daadc45c802a1ec44a7add66b9fbf7eb28fd768edbfc2ae2cf2cd9cbcd3a7f5ebb155d184694
z5f4a2e6b4a1ea451036c2cd3741c5dbeb67d42b98202f5f973f7b9afa89ab740f60f6223dc9443
z7054156a65f00bcd90a1b2d839e9706e6a31c3f349b259621ead429025d3f0238ebb333cbe9359
za71dee42eaaae3802b90fbb3b83c2c078584bb6df8805ccc6ca5557d0998767504b714b6c7ae69
z4ac9af73665496fa3091fe7092e01698dd90c1ae7bda7db4e1730a399ee1b05226033a65f6512e
z1fd5f152f6702f942c432c2bdd4ce01f0773a47bf8e660a3d5938343ee01054f6dfa4a3c97430b
z6ad9c739c996c77fe5025cf8ba1cd8a4cc5b87c3a4c1b87eed149dc51627d5adfba576cfbcca22
z453edbb1e599d7c731b51bfbaf360513d15e3e027c921345efb7b7e17051b2b004e81b893e2902
z7f09ec4a9d57b75d1425c4108df10f5985b7a63e93dc1dfff38aae668308b4453a6167c1a50e4b
z208e269f0f7e11c586d0f63ca2a5fd906cd59fcdc5cb8c203921a2e8edc04ff7677f9258958446
z39d570d29eaabcf8a648ed5ef1a98ec6af7e62c0812cd6318e0fa8d03dcb03ee594eb5b61707eb
z6c0a04a66fbb951f3e4749d22cea5cd90682bf64823655deea291b90e860f7664b041338afd730
z933478616ea52e17b90712686dff43ec343d7639ea8dbcab99438a2feca2bfd26816c2185c0ea1
z7fab3e404d19925bd8af68199e4a22a4fde638b5317a63aeb49ca2ce3e56a461c600554af69403
ze4faa006aee021cf28ca5fa5dcd7024362d0f78b237bda2f4bfb29d4bb653e403d5f49521290a3
zb24c3cdc6778cc2b23c09f59b2b120cbfa23ae2ed2cc97867afbe08d6fda24083baed98fa3248e
zd6592b0032a2c495f7394bd50f12dbcb086d3d1978173d7e21d401a02721b39ef4c86e81a8bf1f
z87f317d588b174152ce81aa4817d55afc6fe6ea7ef4ca53e7f79d1825918fcc83775ba4e237cf5
zca0f94e9d2bb29fbfc5ec1ca4989e7fdb6867f3b512650262768d7425ee98078c0bca12a2bb143
z8b8d154a4fe90cea6d79a65785e12ddc3bc553cfc6125f0801fefa0ccb4585a6c6326e8c1f0cc0
z9e705de7d46c8b2c8986155117cf7842f61b97ba282af97a8a158912a784c55cded8d3d58f637d
zccbf39fc7fc8b6b230a459471c3ceb02aced22cd0c756e2cd44d4d00b7075b7e36e35db5d1eef3
z8bb140bca095181172867ae019c172ce06f6a34d96e7dae6795e449b1a6fca37745c1d2a5b9846
zf86f2f8c9d92842b883d5973bacdd8b822250d04b9d662d15b6c98781205aee8c5c9b7d8b1fac6
zeeb4b99e32b577b87064071dedbdf92f6108edcc5791e253d43af861095009a9bc261cd6628279
zd30e55bae236bb31a867f4b025a41c8e1dbad60911dbeb88d1734113b07a2261adc7cb26fe0307
zb584ccd2e9400ed255768a9bcbf5733fb4ffb102ce82dc3fe164fbe59b0c5ae2f8cf0596137a3c
z5a74264a5fa63ff4be2f6d474e8bf6fd0941d2d4b37db841bc37cc30158b5ee735590cd1db1db8
zffa7fefc3f6476435967b1f32f75a1e7d0468bf8f67fc12964f3c4bee15b9e44647943c9280e86
z5409d5e051fc9ed90c56d259b011ca0335a2e6e8076edc51a35575c76b5fa8cf36eea7d5f702f7
z0e4236af0bee4ac221e3ce96a35fd3ad7c40f02e4208215acb894fd8ed1dab4778b64c800b41d1
zaf0e1d02ae8b5373b600dd7b7c9d7fb2887fef6f1b9b408e80ba7982f5ec9b4167505ad0641e4c
z7a79fb3d2ddb99e1af0e861db94f65cf2676e409e0b6f9f09c648c164c9a709080656de8c45ff4
z835545c6aa052376e24ad1fbe33a6aaf88c511cf55719aa79e03cbf14bef964bee12396603d537
zbdc3dd66c0648b89edc9cb7d5e0e4793c7eb027655a8ede9e85fbaf1e6d43235ced108c818f14d
zc2da9fb54405226aafc70d6ca854528e0b5c77a911e1ec8b93103ac55fb2bedf94f2aa825887df
za23f68d9ae8cdc877b3336b88bea7849e86ad75e50a52182f575b2a9fdb9c7f574f42a7adf0955
z9f6f9cb4c8a075a9a2f2d0290046b8d7dd96b80cb1db9b9c33c950f9c35366bfac324c5ed53cce
z58a7efd9e97b2e04b1db3f7106c2706dc94b3b7862ac7693eb7b41fe97d1a3a11565bd49712119
z2db3a17b7117301a8ce4c2836a337bd23403fc5ec5b07c66e7092487035fe3f490eaac31f710ac
z083a02e859ceaae35c9650431ff45d19bb4d64d63d3a747fd706a7972b8fccf883d5542ca24d2f
z0ca35368a23bb5b9e8f1cf79adb4f3c2c003ca60aa0c8dd8fc15febb47f4100756e37f01a186bb
z54927eba2d49661d64ce9f0df4c6df3c662a60b4ddee823701714eaf963a9577cfaa9d280f46be
z1dbdbc2c1df2a6b6b3a3530cbd30f0286998ea3aee65507d7597dba2fdf2882d9c872648beac26
zf8fca4e2497d749e09f8174b5adb26de120e95b195aec92f87bb55cffcf7b24d55ae68446cefc2
zd868b8831c4035d7dfa20a32b760ff1a21a83c029763fa7b3f8aac1e606db74d6033b270a25e7d
z25ffaf6c483fd70019eca52caa0d5a863a22d4a22e4e21787153d509c4710322727186b3b51e45
z06ff185d268b32828b9aa4dd3fd4a2729ce2de9e6e35ba83037ddbde23ddfda5f25a98c0039d76
z1e383f192d93151526a9b890d6c185b31c56405ee9cf0a324cbcb184459345e34a2688139c398c
z307d02eac7c9990425e11e670c5b211f3ce87d68fffca7396898dd9fb08fca4b92d5f44b3c60ae
z15a87c84bfb9c04ab3c77e6923a40a87f43796369551a532867bd9834504ca6eb6141a37c6032c
zb8bcdbc946a14297e8192cf853bf858f4bff5f2147fcb77baec696e0ba1aae65292051cce7f512
z672124c1172ec4c9c28373e9378759ed6f78051a917f1deed225374cc255fca8bb8a81f8c6d66b
z787fdf7eaa7e0e75a5b681da6d4a721da088b3c6da9d0e89b28191907d240710bdda936b4d3976
z098b0f2e09f88ea881d713e1a92b80cb587615902765156783e3701a146cbedce5e1b11001a002
z3cb41cc3b2be0095ad28aacfa6afa1cd3e4a11979fc0b4c26126de59f8277d84b2dec4a4a64b22
zfd4d028a0ef01f9826ce261d793f9ccbd76ea67e9a93ad1cdd6eb6fb6fe5881fd09cc83d07f150
z99474059840f965c94a33ab6278427e8d088963d6704cd78e879df248d70b18b09ea945788323a
z052d164c7e6069b281e8b833c2f04b400a2db1aa1ad9344242f581db6f3e12bcd0e704bf76825d
zc54e7425fa56098b447abc0710165f8593a180a322b8e125e3aab00ce03b3057032433c4c0fea2
zc69b6676e59efb61d1ecdbc9e6c999820351e95a460c54cdee72c4222d2da6a5c941038c17331f
z9f8715b090cbfb0cb2bcac150ae340028c3dcd3a491932842676ff3e7eb570d5b25012a45990ac
ze7515174e9ee0fa30081eb0ba78613ff69c7ac33f55f60d5a5bd052d1f1404ff4f6c06858a89af
zf59358cd1aad2f3e918b5658832e5529c444638ad397608052aa26278712297ec25286c10e92d2
z8bbf792264af46654b6dd38cd05fc03b4b71fd11a203b369ec41598a01534565dd82f785b7b7b8
z2f9a312a1d155357aff441dfc90b263143b02b78c3976995c5bdd67d0ec3b6189d272c6ba79343
z7f368c6973ac5f7b589101c0d16f05166b4750c8cc79bdde08005fbdc8404b3f6820c7e58a5d4a
z8d8b8b754a0f09a4e4d6b1789bd478b4c6ac1e6713a5b43ac51ccd2bc4d3edadd756f81cf2155d
zf35876404554968af2e8b5c4bc9cb8dde74189218ea8a2f94cb9252cf0419fd5687c14613547a9
z1b92890792ca0a2450ce925facf8ac4e780499ccff0194a718f2cf16be064c97b7220231cc20af
za0f06ad4be4fcadcbb8f16fbac32110507293a3c430c1e8da9cfad786de099a7418de8cb966d13
z2e2acc7d55fd18f8f59e10e52a3e0bc1d820896f4bd3feb151ddc1e6a9f97d5ba26b0fffdd02b1
z9a4443a3077720733ee46557efde9b7d1065fbdd863e7cc345d8aa921caf3a015c9d21ffe85361
zff1801f451cb64aead6d461b4f7c240f129cf9d539d3233844aa9b1cdd5dec4fb1e4edc3517d67
z003fc194d88c2123d4c0aec77e620280a3dc406d5535d0361d0a0492bccc94fd7457803f87847e
z85bde453e36323846fd86eefa51f0ff64904a6fa64416127fa924eb7680243d6fc1d8491119735
zca83cf0e72fc6a9d7789c03fbb75df21daf0c48c31f146863b2e698367755e6b3fdc867fa493db
zc4f4671b866905b2fb036b17e347db3e02a388c7b9501cb6be72e93e424588edc967c69f1072d9
z2e080ff54a439214e36a974704464cc46263c3ad23439f6df1787ee2e40d22de1934c5ca44a69e
z089768c29ddfbfc8bd057af89f9652b102466ca2f3261b2419d723b61a27e439973432b3170373
z43e1648323e9bf7b2142e70c9ba0257c2cedd20c57751cbfcf2f12dfe27f5e6fd8c5cabece5738
z2cbe8800f39fedcf43784df08ad6469640cc48a086e1c35bbe0d68e56144d8a7ee85043ecdf2b8
z5c38789f1c3b4eddc50a58130133cf0e26db177c04ff2b276691c076e5adc4afb027f21859de15
zd6ae40eba0e574e87daf10e14b449daa75e9c206804fca3a9bdabdc8e34e3345c822c2bebe627b
z02b2619f36d59d9d831b796d498dc42e9c0bb06d87ef46c10e2b43850192b53eb4441e2e8be188
z70d0435c5dde13ada093a6b01aae6dd9d9127cbdfcfa6acc33e1e81513026b59024249bf94bb3d
zffbc5d388988e5188fb3cc66e48560428566c10b50cb64709d171d7fb14fc7260feda40e850f9c
z89915abd748d3a8836324570e579160543ed4487bcc1bdd7457bbeb7a57da5cea20a453b319488
z279a9cab49f825df4275713fe07ea4962c437cc51bbf3b0ebd335853be051eb14652e9336b382b
zc105cc52a29e71420607c2015dedd538784365102a5dbe00d13a412470f606ad7af4ea2b8d9cee
z6fd72b5cc4d30456d8af9d58d0a903275e8afdc03de86928ae4b5c2f3529ae665c0c930b91f096
z27987c43f7a34a0d853030d9bd3df7cfa43acebef738fe8efe5621c523b85c5a68a430769c2ffc
ze2f656ad9676418963dea3e914b2075f7bec15b244dcdd929939ef66a744249ef937f6b233e13b
z8eea057690dad76322c648507c9a792458cc5866238142b930043fdea6b10219ec6c15b74d1822
zd1840477898345cf9ae9af0c0cabd70722b5ab247c7d33beeb95d33ee528f17c45c70019040552
zb8869690ed4aed35b6d3ea3000d5ad4e06568ff8c177336e78c71c3bd4343dcae8113add1be5b7
z0c6fa87e1d77c934204853fced3cdb4ce7edc66be2c222c3f406ab5c4a16f5bd601db9559eb5ae
zb47c4b275441951eb8177512ba30edd5cc58e381d6c77dd0c34b04620291014abce66507fece1b
z58da35cc62cca7ae661ab94356ce6611527d25ec9410ebd1186306cd24d9cf123d5fe93cb9fa55
zb4635798986073c21a7809cdf1cfc6abdd3177ebc19868a073cfe88b14c91be050627757e9a9a9
zed14b9cdd58fe6b2dd6b435b8653ba6d60b3192cd0162fc738870c8384e4f72f87327490fdf2ae
z70faef854aa50eb58e8d47f9728f099a856b18d2e322e3464c3b3a37ebc4618c8c2447c4e796e0
z4a9a449d38f45f929cd69c2c9d34c5681fafd285de1ee76768a238138fba78c6b49ce8d775e1bf
z7d22379ba89b38b1116447dc0228cf5b1e1c7a04229b31f60c983b882d734b683dedddb2343d86
z09d0384465d634e022b0c726da887823f2deb71e4aa4fede68871fc9abb6ab75a9ac98f3b36dec
z00b5ee5a1f62e5bfcc114ca17480a493d3b9d5a4aea17f1802a2f54167fb6d47a3ace4e1826080
ze09b36140056a3fe63ad3e22a07d0f9a89cca58592e816d61d4e2c7561eaa69aa061433dc3595e
zeeaaa5c93f2283fd080d36cbb7760f61a208e0473945d06c693ce61e0f5571f9036dea56b877f1
zab3965694133ec9c83b160830c24d98052d67193abae3f9e322c86e69012a730054247e4b0222d
z7e9e1ad82cf8e2db305f97009e72ef7e23bdc937f2becaf214a2e72759590e97438c4b215600cd
zd02f2ee289e15a4951579f9ba158111f04c62809dccaa9fc45498f693a419f953758367018bdf9
z409336914eebd5481fad049f8eed9cf9b6a78cab8753776e500cc0f56419829382290c86d61ee2
z82b4ff6830909e62dc041ef05b59d94c413099747f24c77d51198cb6a63ecfe914c1cfe3bab02a
z1b581cf3fb955c13b39583cacadf3c2b515994419aa387014f488876b4283b1fd548a42676c95f
zcb81c7bead406a2b6d979102e6c51ec0485e14b6c0b10b9404e4c494ab6d960ae91fed27c74f68
z05afaee43d46e053605e184060cc914565befe69e11e9eeaf843286f8acbc77efcef35c5c56060
zbf1ce01d2e1d3c234d443b13979fa5901943dadf21f89b86665e4ae10af4699e4deb4d74db5595
z7c74bdde766284365bc14e653cec0819b419be43ab5915a3f573a35c9f182553bb169b52fbd34c
z00c8f6be729510552fa59f2e02962eecc45df7326e42d68c2953e2b71d61b3c76d77d9007e9c72
z55248e481ac01ff2539b141c444959ebad5a3d5af546cae99673f39c1f5a20938fe61cf5280683
zab07039330abc8397d1cc93d77f0f524afc366dbb7a41db8e6d424e66d5736eef63bea1bfe1b15
zdd55a26cb4d31039362d2e77a08fc74889e66a8c07e7b198e410a164594cb50e43276963b6420f
z28c1bbe73329ebaf757e9a8d77dd1d1de1d04fdcf908c8f33b0799f2200c04ac666db94ad93b67
z5a250415cebe1779e6d5e1e453a232d3dfc7caa84e4d48e81483e7efe2a82f845723422017a738
zdd2b41c69f3ad1952668fd6c130d4669e888d1e8d0cf326c631d8e7408833206640e627cb7884d
za3368d6b743f62f0da29354a296d3f82e970c993b37f05b9151493182b811b50b4a54bbc1b2085
zddda7ea1dca8778f15fefba4e67f6ce0e565830863ca7fe4582d01e0f96fff3f58faf5b2f42c24
z4df0b7366d15957f50f276a537a6fa751abd1b00063a756a05359fd2ad2abab72742584d64ff26
za9bb64e5ac5efdf2bba2ed7f0e24ace9635d58dc8d430e311b3b4d2f7aa610bc57c28ec2cae58b
z713986c9c1d284557c3d29d505dd73f29dc52734b940198a83dd2a72ba1bf3daba0631d906e33c
z2fb78b876d028ad35c9f88aa26206cf82ae1d5139983b5dc22580d6d937f5594e5015f8e5d121e
zcceb4c8753f5f9ae67ab59419841a383f85ac1c2ac258e48202cb4878225df4e94831777f03ab2
ze8e3600b4573da43d0eae785c5ff6458efb7c1dbaa3aaa657259ad3c789bc2068227dd7703a8ed
z506d765f799c5913c0b9e11c6004c92c21b6a05f74e592d38003c785aacaf2965dce879d9ee957
zeff30cba11f1f512b4f371b168b953c22207670b7a1a0f65d52414eae7e35fa8ae81f5f2884bb9
ze570036a0cd163160bd7d603d61198616a0d57c111245bce8a47f359bb1714a5e3b3607765f78f
ze5139fa086d7c7907cff4136fdaf9f036d06dc4d575a8499b4b90f22857c6b21249d3bfe65492d
z78e6d437aa465fff1c57bc2511d52a52a49ce3d5802ad4a7600758d46f3185010cd36a468eee26
z712510b88da141b7f207f31cd146513d8a010740fc998a7ed09bf0bae59d02efd4b4ad158c5f56
ze5634c46464e92a799e1c298922594bbdd11f06561667ea824feb8a1c7ce21a7de9c5db3b9393c
z545c9addc0a946a53c06f79fb47b1a3346f4ea935997a51b814f4bdb5f876ba8a299c15b8ea6ec
z96e5111991d340088e2ea433c3b86fd78310f7c3819720cdd8afb2241fca2c5a97bd8750edd634
z4ba30883e227fb57fe47a5e85bc363ce20c07dd56fc5bdfbcb3eac01103c6ece5c5f4f2f9ece97
z7224c92de662eaf4098bc6baccc456017c332c858b360e9a4cdde3e647c4a2b1cdaeb73da88ef6
za8c61a8442379d81390f98e757df910feebb5c8f9894097a423120703f9d88a7b01674faa4a511
zc818148cce1b12f5399e1dff88e1cd011fe296d77d38a4aafcc22026510e9d3646d789af0be426
z055d0e9b3a2f23729f28221e4412be25fefedba128bfad8b0bedadf0dc0ecb71b09e452fa37a49
z72452cbcc6c29271327febfb1a75cd73828b6a06c4e5d406ad9a965916b51594bcb8db17c0f7cd
z620bb1de4dae946719dae4de596f3e10399f4548e227e84dcd04d1dfdb44d3c7ddfa2de66503af
z6bcf07f40a9d6fe1973543fbecdf84daffd113fdf4e4c3ca4c7cde1e3a67935b163b0ac68db085
z3f5a5802df3b5f8bf8947a6b22c4c4f83013f9398ea892047678feec5dc4250ba42c1496462896
z25dec42676338cff4d1343d78dcb518215a461801a625c65702ea67e70b63388398df407916859
z3b98ed0f9eddc330e955796ef0bce1f2b914fc024bf5ba7021e497e9c929410ce73e33b7bb7820
zcb7416f50b763eb0e281964c04ac0829d49b9f2a2c325c01e8d3ff1755a2f9578c6b0999250460
z4808a188d14c59f85a2fb34ec6c9311a05a1cca22e66a363ff5d3659585e4299369d472bcdd5d9
z1f992606dc498750831c7c482a4d4faa8e37736c69ab2b96b2dd1c5d9fa0e0dea2e4c658cc35b6
zee28856dcafaada42057d1c53ec84df5ff3ed01c6ff1827929a71a44f12983087ef921c615a4c1
zcce9aa3069a6c4302202c33b2ccb74e843e3d529ed010e5845887dc42d8abbb31c93848a022854
z57ba4790823df29de68445679519aa9574ca44f06ed401c497ab85c0f11c6ba17dd6729efe505c
z1a7bbe2e23fe9573e3d4f9d8fe84d10620e5d066e56728cb24d248fe7ba237d645828694615754
zaba67ba1281c62d2cae04f0c95255f9735201b88e57ee0cc4a55b498e678595b8f0016a3c2691b
zc72c2cbe04bb875b50ce1de4f17b411eb083b3157e4fbdc3b4a76ff08b856b59c968a8c76f83fd
z92bdbc07b4be349b3583441b6927b00b2d876c0564168d482ad56c1a3b9711f0cdd1c9205a0ab2
z4ba616fc9df4b763e83a0399bf0219c09611efc14cbecc9d172832c7751ae81b22440e68fb60e9
z2d5e11f33a6d219ad9030d6d4acf1b4e47259489fe94e8a76bf4c16f0bafa6640a9cca6a8446df
z21ef2b43510e2231f1c16ec973e3cd2f36e7acbf76d46f4be301400630aafa609e5e7e597d4269
zd980d676d5befb34dbabb5cadbbf7c796b2c8bb289460babb30c29acaa573552e448daa2046592
z7d8c8ebc02c8f1b9d21254363dfe9940b4dbe2f2c10d7d291c2b20f5e1ebf64d639de0720d77ee
z08e116a17d22027919fa1b6cb5f17a0621be043bff8b32665cbdd3a0c4c5c7b10e1b4cc8fef09b
z082125c29721190b33c5f2ef8489665e3cfdf8bf46f4ea8ee993a75d48ec18fe9e6b4036333990
z14992def441d69444fe85f3943f3083f90fc8cc9441971f921329c41c33049b6070c63b5392c45
z6873dd85628f05dee6bb419ff388a7ce09a13f4879d084836814c921d0e2f8fa4955560fcfb453
z7bf8a1a9f2a957c6e189b79ff3053d32d7320c709c2f4356ee713ac8ebad5740d10f77ea8b0949
za0a76f96739f97460fc064705b62ac53389322f11df43479c03b7931d0ab0915b151c93136cb72
z0f6b4db9bf6f6ff8437fa3def25f60b5312996cbb5ba93894b1d5be27a10ae43f59afcc36eaead
z63fbb00b66c4216399591ef66f22ace193e30ce130c22f0d22e72f7a9f0b4d925abe79a0b05e09
z726aac6f1a423b953dbf60a1ca7aa028fb1368c65a818cb000a50acfedd56c5c8309a40a662ea3
zd02e834681cd6e7481c8e05267dd753ad16a0ed01ae2c3e2dba6bcfdd2a74c276ef63e671f1e74
z98a311c5fa1d1afb7a51f3327fd750fd80b7adbcb88b5abb1e6d2516faa685a19dd941e5794695
zf5d2d5f387b6f4179b4b691d58f609a016e54cc518de703d1ee4a59e58e1159902625c77c2ca02
ze5185d7e08c2c4392a2e454db0977a5c843492a65ef1ec48359ffbd9123bba907e8b71da957dc7
z84c1530bd43974c8f60bf8fc4018688ae012325a0b3c130534438ac58b347123d0632999202858
zf95541293d9128409be53c4c2a77645a9c1336943a3b119c66cec5821b49b1a0b762de6db3e15b
z5902102c1ba41aada14b8ed545fcf16f025511d6a992b469ea98cea5ea68714f740655d1ca6762
z3799fa997214752095712e180f87a314f8f93f7addedde51c3f280060aec9687b066a6ce50647d
z04308bf353af3e111c074ea12afe3f101d77d3a08dc2ee5ba243efbd05c3e033a14f6e2f55078a
ze7a2c78f68c77222f6299e8dc3ee3f3a65576c990fba41cf5b88e9b752588e06e0a5b25f69d038
z47b181f420635085004a2356c579de9d49e32f6243037a67e3bcfeba6c7d6e23a227515d012ed6
z86b8bc18e2b22707e762a5e736692e50bcf75317924f214c8d06986770f916c7eb3488ab1479c8
z811bcd8452159f464412dd42a32affb95471e7ade9fdb015c1ef8082fe04c0bf53f7d6d06a1be6
z3a1e459a85fdc25412b5626af2a57a0aba2a5493ad474a855fc9af435520d95bcb651f6adddf01
zc89484276a6d96bb0d9abe1019f37cffdeee383533b0e72034b3da07affce82a6643a870d15a2b
zcd4bbb74b768fc544cb64063d9eb39691fc0730c464c1dd02742398fb3ba0073d7840db1eef32e
z422c58c2c472a973a1bf16e053cceb6888bef385d9b4a520af366c2656c53834666f48572220d6
z0255c666372d6cb3f20943abc55239d804d13c7b5d81a04de849a6998263e5cfd9901144117401
z036ba0f2d1ba61539b338aaaafdbc3cf342b2289c627777a17de52f0fe8881269bbe4d75772d87
z78f8549aab575218b995b3a4839d3a91dd75f488840fda669ea83b62174297931e63c7a2a4192f
zc941dbdb3e35c26a36e6af473f2b3778c52aa51ff1a072ac720446dceb85f2b219b3daff0a574e
zcbfe541ee083c23424b146c41c2d04a0a6613d1f85bfff970b005eded32d5a99ebf26a57741482
z00d220107c3834185e91cf87c1420fdbe883b7946d16e3b51903389d790a85e78c2bed3f88be06
zf20125d9552e0f9576d958ab006021c173597b26aab90adb006b0f315d5e5f10928013ec412e5c
zfb929f92f530e18a15d3063368275223a87f7db60e72f9c8686e734a16d5e6e9ff4bc58fc160b7
z83e0e40dc594bc8dbb0a54d30e29a2d309939a25ee512a12af9fd508264ac9bcab8588ca668655
zcf7ef9feb3f78910f73af4ec3548ac534fb50464e55c3ea7640778779a95e7bff9fff61ad7974f
zd78ecce958c025c6220bb9c26249bb5a16fe9f537bd8560f50a5fcc4b47b74375bdc0a1f646ecd
zd7633c047a8d0fbeace7b6c9dd27ec76749b47cfed3687019177d5358e8aeac7b50632cf89b518
z5cbb51ceb3c40bc345d83a0bed1245c7c48664816da6451d911661ff9ed3edd14dc4e197469c2f
z310108cba57644f1f2490cf51c5bf87099c6a7f8531f41ce7dd67760bf1030c1e85bb2988dd917
z17a86d449ad0c184dc64cd4fce3a15eba92bb3752040f3a3c1e2131b7d3b564da0f863a2a54b9a
z7e70ff1617f53e0ff051df8282078271828e2ebd8b19f891dee273f4d1005557ff593ea6b3a973
z1c9957762c382e5b8015f300c484ced1bf0e7e59bbebb1ae327681c91e2be74fd6efab3223a996
z4319026f136af22f703a12a919711e8636fcc47134c49bef1180cd5da5014ea9b8a3ab299c9cba
zf6b2acf555757377eb87001044435d87639fe842d251613d7fee7e29baa6f50e925935388e965b
z9adc36d61823af645cf1cc8a95d3fa3af3c045dd64a58e780f6f9cc1ecefa9c9e5725f6b2f8fda
z85b5fa17b4fcd171be42b35a3379b6b2b3dd986893d537f08198f6e6c9bdaf9548610350808477
zc78939a03c01f542ce989494e17e04ed77b9f50499e7e41e510f6e257c16d3ae6882c44645773a
z28b498d38431575e0b877f986164e3f9fb91e939a901b3c83795444721ae0432621e586870f224
z46ac25deec0e5de8608d16cd5e44a18d0262073bc0c7f0ecb56e04bb5cb31e5f11bb1ce778cb37
z712951d6956e86b3b7c8b0ac23e69259d5b5415b3ac6f04ac20b7481b5f49879d2849875aecbc8
zcdfa4122ccd2f948f27c16ae20f24e5110568afed4aadc2c0383ccb198078aa7b5711b036e08c4
z8fe3d586498cc37f8dc5e5d5a81af8d6e0b748bc5f048a238366f36eaa07397b5d69686f69aa07
z6ce5ae6352feeaa1cac167ac41ae27c4e183c6cd96bddf95e9a4391bb78ef2c85891a0e5033e60
zdbc5597b5f02f9966c66144c11a9ed0ad21a7174e71ccc956bc920d9921073604ccd05d805462c
z529c38339e3da3f683ddc8c36e52d3060ded0250c2fa5158272bb993106ddc6fd11f4a91181faf
z7b6f6aed2accf636dd22106cdae80be19864182bdc3a7f77bed287c6a34c7df6f45bc739601c16
z532013698aec6c4596a6396b5ee53128bd723e3e52043330ba1d0af9a6de0964342b4b1ddc5f0c
z142f5d80634280bdb065d81bd3eec3b6a07d05444d3765870af7eb8df0d4d31d45171699311603
z56c0e1a5cddf54dcb3528b5f6217869a1d128a0e0965b692cb45184f81de7fdd882694929bbf5b
z8369416e88b03e03cf759cb035cd7935ff2e9ef68f2f3f42b5f4c43b0a9b4a9604cb6e66bebfc5
z9106f03b8e1a5df9385412e55c02c74eff271600647b93cb91ac293bdb397dc5ab30e271b1f5e5
z818e7b5675b5406cbd81fa321f328753c4439bca86bb27405cf74bc02536e384a97fb6a11954c3
z240ff681c304cbfbb9d2f5de0ca69a892e8a694828035febf80174ba9d019d966baff9567abd29
z8e330a55d42d68bc57fe34334d4676c54e217eb0eaabceae35d0842dc27705c4ace23f9120f63c
z0298f35f85cb9899b1b19fddbe4e2f4ddf37f39971ccd879fecd614378c8a18df5d56fe3b7affb
z39874726aa540edbd80de37efa843484879fbff49aa6dc8237771e26e222bf97cb1d9c6dc95ad6
ze7694271a9256677b5cb7e91cb1bfb4df06a164975ba779165e59a2ee7851f76bf8982d655d7e8
z59ee9df146b28276cf43de3bd50cbd5ced4996d0a53c9fe6aae6eb64d0e23266b66bc02832bfbe
z2ab64638ce0bdfc527755e077c5b1a4acd1c834ac7b6a7f61c004155efa9836643b79f44e4c2fc
zff9b4d33fe6937644ee7bddb20c472c630ea2531be84ef8c070cd9a5b388e2f4f2e5c03c157b64
zd63f35270c5c2d3b4848a27d6d9aa425b9baa3b9c51039697c956f23b826364a6b8fa7ad39c2d6
zfee0201633bafeb202f73cf4882e693da2859d4efa12e7ce5add57c8457876299271663b1ccebd
z0b5d94093e56f673623f59fbc644d73b79fa091de7cfef0a123531c9701d8dceb845fdeab43994
z0f6a52e199c5d1d6c1abc71b565d066068a4a796114752f04130d736adf8104888dc3c4de16363
z859ad8f5cbf9aa1cdd831aae3b77ee4769e7d68fd0e0bb314a1bca27e61908bd772dc7120d6513
zfad6b381e19f1ed304022d856dd404d2be9353cd6552a8ec35f26d58ce9c540c75742d58034344
zc485dc8748a4eaecd353ba42c2aa487adc793e0b6af9df65e6715c8a66206afcfd72062ca7479d
z42bf9c33a2c96f2197ea3b526c8b779a8e13ce1e1aa73e8f6d3cb8afc318b58e79b0d013bacc7c
zbce6679fa4b1ef08967f957e0099c54ca379187f57d9706551bb2ca62e82a02d9cd9e5f2df7b67
z37b39e62de13b37c8e23c697273f73c380b13eabddd84b56f3b4408e601ca9c42e09238bf54057
z81f26c7dc4837080c204e54ea7ae780630f91bbf44dc2ff148bbfb73c84dd541da427245b47820
z59b0271125a78781ba9cfe069d6bcaa3b991526aabea44eccdc7b4aa2ed083e77bfc4ff5cd71ac
z6ab189dec7d9cdd7dfcb31fe168d7e5c26ee2f30a4261f6adc410bd4a934d322b675c74e65f234
z84b6e69b2a0dda916869bea6b597873912d9e545fb94cd27b77250bf5fe61ef49f4b23ea529084
z0d9d92e9cd62f726b79a2b4b51353ebb1e4c31f25cf8efa40641234c2590add47c3b14af6e84a9
z5a9e2449d0a39b6ffb08484d6435956a5bd3aa5c5a8962dcbd43c2b02329a5f3d6f22e80e19508
zf8715720cbdf032883ce02445b829e53a281995eb93603734ec431585f513d20613907f6afa9c0
za4bec581548080801618651b6c6379287064909740d4c6bc79d00983b910f7721a86f1981e4f7e
z0ba456e74f0f81ec93de0759cc70cdec9dc8529d351cfa4eeee9f7fa9bed75473edba721f1917d
z0170fa29c6d342f24532ab501669aac5b2dd27dcfcf0e353ff69cbadbf2bd33bbe21a99d7c7be5
z0ca9c876ca672a95b6931b62f693955afc5b6f6b3de2e4e7a17b7710648a6a53369e148279ab8b
z762e51785ce4cc20f1baf3abb40f07071a9d2a71d048d333a10909f3758548079d88811b0d134a
z557bd66b70114e5d312c83db96d04da16ab124b5c65d59b84bfb2b76accf986a0282db4b19f173
z507cbc34df8f7198b542943385abc03399cd588f5e4cdc1e11f6700c536c9a4c205cecb88084cb
z56b8a0ee21f3b9d26df9bb19b101fff64baac995356c126ee2344d9aa8faf43844151324f39f0f
z8a81781a1540f76b31119a56029e896d1915e662ea14236057de463b7d7cb20e4ae52abf674631
z29c6c0b691b908702cce8bdd5f1ca6b9dc09fcfb49d942bb1800943dc2b59be9b5d19e97676b43
z9a858dacd968a94cc36893b1139e6ffd9cf65173bdfe5123a197b9ac589d642cb17802daeef2a6
z4401258259a0c5f63d267f4d33c9d3c8e62da79a5002cf099f890e0c3ece854c0a3497079cfff5
zebe2d38fb82d88fe075bfae16b9c3f2c5ffb7914b13020f9c1d557c6db208fb343821fc5b3c46f
za9302662b83d30c959a5eb6df62b9d16aad0e590010df315d503851daf60e0594bd329f1d45c0c
z7f0055daa1a372e7814f25d6f56babd010d0ea62dca52e10d868f3204b6a5436661319a616872e
z8a21ec83bc352435358344edc7683678f404b1ed11f6d4293e62c568228961a2a078ada75c6cad
z66fe971320afc0641036fcff80ab9f52dbf6157f29496d9742c99f861d3bcbe7ba86ad5b2da1d8
z98f4b491bf62c94736b54d86ef396a3a42f3cfba062bdf56c89ca4bedd3be59275eeb2076040c1
z204603d1121de419b1752d16c076980a2d7cd35be50669ef3ab5fa699c631d0dd4f039d1698f09
z18a57e00bf956ec5d20ac72aa57c7e8e336c8270f76873a83ca8fcf48619665e5a00cf4b4ba502
zb667d186e958080dc9a2c50c2e50fd67bbf07f955351b9d34ca13c529e055632bb9637ec403042
za8c68a4e7d320d2ad930385144ae48f27c7e6bd0a1e4880160b89c58cee36a742b7c2bd8c79d71
z2966bc04fa1b2c46ed8b7d8c7b8099e07c7e5bdb6fd55f4691da3bcedc8ffee4d94403c9d0a44c
zbdede739a0bda55b2638f1ce1b7e9fb69cec06f0710e8b759ecf1eb781c9fd951872fddfaa940b
z09c2ce89a41db72060a781bbbca8db4dd89fe4d8af27a0bf31a068db6642313bf650f77ccdc882
z73b1c99eafacd6b88b1ad3cd517c43d32d5dd2fc6dffb485f9ce92021e3c5d6c997558259a797e
z2f477511c558bfd547787866ed35b932834d70dbfbd0759adf1f1274ec099517d2cc1bca93c581
z47551bf9f3c6b149f062678b6927673797b9866f4c5ea66dfe4217b0cdacec25b37f0447addd12
z162b74c48a985bf6bcde63406806264a1a1f7e2c00c6e87b6030f546ee3be1adde34cb701e1f5d
z5772d7d61766363a30bdcb03a96d5dcc5f13a9434ddd1adc5d8d2d748e5890223e53e84029905b
z505ae6d118e07a171c5659867bb35fafc574b5fe4383c83fe319471686457fa40257bdf372bfd6
z4cd5cec40cb73411c406c66232d06df5e1492ae59efabcde9e3bced9904fecf4814d79c42fbae1
z060a77a24435425eda613f60639d6ade8740d7593cf067342245b630d3450996ae3c9dca9d19ac
z8e825fe8fa36b1255f04d63fd2033896316aa95f7c36b3d8cca6d8900fe708f50a1e8e27cbed09
z12490d8084e643c8c1ced5438df925d157fb078ed100f92765036e14ce6f28347d13bd3958a127
z6f86a00648f85bc37caa5500fcadd254b6729ed3932e5a8194c663ec212bf63ed4d1eb434f6da3
zb7e1a9dab4cd931beff2fbda301a312a87f5a72748a77fb38afbbe9f02c68d7bee0137d663907a
z936831e4c9285fef0881b8dd7ca8f27c993fffa1b0857f9ddb97c9c7e770522e49fdc0c9956ba4
zfe01b63627122f1a017f5d4fefd1454abb9644b849d32a10e356d8fe37137a4565e2c36eed11f9
z14f5300ff1737892dc42ae09f140b3b571a198f9ffd041407ed813f879f238b72e4951041735c0
z4bf1ef0b68a716ef4750ca95d79766b69027cae640d5739056359ca9b06a04639c2f74ff42ac3e
z477cc3c6314627f66a14e535ac58c7717a13e352fa9554f0e91b5d7f3dc4495e476b16c88f8935
z3568aaa4d5e25d780ed9069f0abc6bc3e2addbdcdb8c131c3187f49d1f2fc34034aa0629814f00
zfe1616cd1a3e6778cb32b7386682ea52cf671a35d8ee83847c7a0197b9e48b5f89a5779cf69981
z0d2152fe9945131c13f5455b810f39345171acb510d856d559ee92e31ddf35e03a13814a806db6
zb63b2ca7fcf16afe7686ff1c26e68ff2d2b9e0712cc35a17a048bf315fc941e13ed4c5357a0f0e
z25844d653d64517ca92254664f68beca606a87492f7af2ef1697827eb49c4a0bf3a7ebd42aa20b
z23813e1de9611299bdce9bc220637c27323ed41387eab6d7232d5d1596d49f23fa82d3d6d6d0c6
zb9850e6a6e9eba424df0e2a6d04d9f466cb275511267fbe50627ac8a2dbf2ac9446b3881b582aa
zf6c50e7b34e7e326b1c7da060dac1ca12195c8c490faddf868136fec17deee96527f6208c5eb33
z708b1c0f0dc234a0930adc0be7b2833c0af2b56d4ee54d571a1b6d3c2de3cb973310b0c8649b29
z612cb3660350ca6aea78a69b231b763fd1c7e965592b92b9b523c1c24b8bdcdf7310291bf1170c
z7f742f29c63bf2050a96a8d3e87e4ecadcf896478d8edc09cb2ea5fde87ea0bcf53baf5c3724f4
z43cd0a22c4cd6418eab176ff4a0ada872818a8a520daaac9b8cd5ed58d7b8964c2f0c19fcae0b9
zbcbe20409ecace875a574428f9dcd692303abf4467c00158590f850cc8353d8f0b3418a93e3e0e
z3cee1d36f833c80e7ff704dca794f5f64b8e0cf6eb1db3c45d21a9a472d037a2c3326acb8e4313
zf4d9ec1f0ddb9b39a7c9467e1e29f7f618f699524f109aff36bb6e483afc492b637421a0ec85b7
z1a41df4eacf76519b2bbaee985bba593b2dcc5526ec7bb902ec9680810d0bf64a4a7515b013ebb
z023f5c67e98b0a01a9cc9faaf540ed4ae3964b7f8b05f1270e77aa187c42a21cdb528e47ab836e
zff48eecf28e71aa082c84b2734cef3af6162649ef67a41a8bbe09c379fd90fb654a22b5eda424b
z182d56a0c1b566b37543ffb763eff7fd60e87ae56f72f0e637b85ac8e141f3e9147d8939dfe9ca
zeb3c1250a8891a5a325a102f13da03de8eb478afa839cd0a9c4866a8cea7d2e5eec47024149fbf
z406842d97fb07898c34fe5890cd8249264e604f4649de8885e4518c4186ff051e0147fe1c948c2
zdbc6b3b32cc03a6b7ad7442e66a674e46d80f69fde8569219eb30a2452f97ef9e97fd68105c6ad
z9f360f2cbbfae76243ae19e9f9661a16190ab15cc2c432f86ceb77f0ea3729a0bbc9059406f274
z9233bdcb2bb3ee2edb25e1c8758c329cb5db437b42239a80405479609c3857524b682880c72eda
z73e55b2287a6e64a32f22f33cf5516707a3ba67e8049bb34367b996fcbf40c6e11aec1343e1937
z9c51b467459bfd4171905372ce6265d0aecd1724c14c23d56129a854051b915f30f3424dee515e
z65e559b096b16b32bf3ce0185c12a8f1470e9b71968187a014f26c302dc1950c56dd1f4d7636dd
z64d33cab4b382c528e7dea13aa9ac1a1e6dfd2bf1a9a55953bb97d2158565485423285a1effc34
z2cca8f15e18608c0b53372e131168ace1486975d0e3111ede6916adbe17109d64d1bd9a47badce
zd8de6b08b49b2aae76feffdaa2ef2ebd6041065335f5dc62054b5902884f2152c054b74ba38e7e
z8959f17a38727959594a27f64c7901b1d6677ec0172a53b4238feeb578e6199fc5b213a84bf33a
z5ec2817ac8dadfd35f80a79d11de0a07b8ff47c41bdda88fac5559899e77db65c0c7b290a8461b
z0ff43a2d17f2ce30ce62298ace74ae90b4bd318b5e987429d62e49a1d2999befa858a782bb267c
z4d411dd89d5d6506921d81b6ac31a94094b9a82cba5ed72468af9ccfd9c4b9aeb94c871af86d3a
z2d24680678139dbf8d813a8a54bf7880119d5c03a3ea2cf912a5fb210f115e3060208f80ed3c0d
ze1b4f14d812a173891a9709f23c4d1bb74a7dafa0d53bdf426c53f4b1f2359a768817eb4526f85
zd059719654af3c1686b1d75829e9838d8256f94079159aba5729fc1eb92b75e9dc0886cf680693
z98af63f50dd126c1da502c5315b86419fe1ab9d4102baa75f4c6383259c376d096bb0882326e9f
z44e18ee38835e7f6b00400505b2de34c949bb3efdb59424acf75334bf551d855d98edd6411d812
z82d52c5fce00712155e7fb162cf73900ab874fccf2f212b5e71ed80089d664fe348d4eda6ca6b4
z271bb5e4cc169e3704d5614e31c41abc27619c1f91665f5b92014cd705d7102f0fcb11abf8fde4
z473a3d4d585113179356aef3718d0cc8131d2f26dfeaf9168c351f7295ff4875e861ec6d09130a
z9fa1403441bac1ca1aeb8e7f43af6672c796afa4b815b8a71a770b7d6cffed101fe86b6a7719c9
zcdd7257b9cefd373eb89563873369fe98e90470a72425acbb225f2c35f7d5ea7979d79461ee679
ze2d78f7c87439ff74d1b20edfce8059e9388617d23bb65b27c34ffcc582b5856a8084ffeb25deb
zcbcd3a005697dac6dc91daecb863b78a4f2c2b94a9607dfd060f98d58188778c666bb9342717e0
z2826514b4b94779e46cdbd963205ad6987228882d323e7ff09c00a3463b8521ff58ac3a9ed0fdb
zbad519115b01f3156b8ea1e9fe5e329c7348dfccee0c04915b1a9641d4de5808de73d5c046a558
z21a55a8b267490643974dce12183049c745c41d3847de6252e4c6696d417ec66c4b31b33118551
z290b146a40720352f026212da0f44a575a7d2aa58243a36d8f0cd9fcd301d5680da5065ce84326
z9374810e4dab2dc648c4171f1744f691787584e666119f63b432f2640a2a733d33128d3dbcd3ef
z431fd4c2ad80fb9a16cf28048a0eeda42983e252fe8811a6ea193ee5e147fed793a4408c8d34ed
z21c3ad578a305832703a6f3fdbd2ed2948bb4b353b864253b86e0c41fe10ff3d2d28ddc14e5ece
z50d8569c64d6c0d0a57bb746f9a1dc162d6b4fd79f5391c3200b0b5d7d3e2a6821029f673e835d
z97bff562fbb722c32282902927d559bb4f46272123fbd15fd4cc1fe91a2a7578f45df846fefbfa
zc842c628c16202ad2aa32d5740a85ff3b0f507f8c9acb958e0e9488cc074037d38bbe6f90be270
za417e6511ebf602edd2586f65368cb0d0e80d98137dda3b7a29665877edcc31a8017c8e8b6eb72
z866a770296d23bea3d4dee364705c1dc6adcd4f575884a7eb529ca91ec1b2bb95645483aa1c126
z6eb2525f6c9a9ce259c161395add70ddc73c099c7ed57de60171c49a37b67856502824c8bc2806
zb07f234729256d830175049a64638eb2e18d128d5aa15b0fd5c766cc6e5d95ac91c931387f161e
zf19de7d7539b1ab1060e30ced7323562f02cff8f0a889fe4e0a8e6cb46f24eb1d751a089a05507
z291cd573020893dccf44e2bb68a3f02614b456a1edf4d9cb7ed58e8a79ba1e130fbb8489c0dd48
z1bd7dba82033dc5e6f095965d7cda32d7a24b8714154d8fab0ac4808a5b3a664b0e2fd0d520657
z6ea32016f842bf6b9287de08a26f647bbcb550ee89a737f4edddb4a219e82a037ad327b847e9f9
zce9addbd6d50364ae519c59e17d6164c8681c58c9ccb8cf1fdb09d11f2e4002ca82ecc9a1abbee
z7f969912a300856b6feb7b42ef49e7336b63ce47d4aa79797fc4b28839d2045a60aa1e83a8ae2f
zec06353e00ea24fd608c8ae3f02a0868a3d393c8d325918345f7e6e2b207838eb99c75af2d0605
zdcf5ff36886870c2189c87b0494d05068cb517052618c68f2392dfaa780a63c96f2983a0388bdb
z47495d330a08ce7eee89ba5d0479765b231b80ad596ae39fbfa44c9812f764ce9b5843761600db
z2010419b37839ac7f91ce86524a2efacc9c22f6a1a7e614f7de6f89e7c07198ae9dd34efc47ab5
z7fd6c2e013743d250fb333da512f1511c381c029433120b3e3069f219c1422c34447a48a3ffc5c
z0042fa73aa046310c774a2c12d7cc2a51368421d11a74394ca9d57067ee1d7b20055d8eefd8652
z9e1cb877edac594350b4ab5a7b6f7409fc44cb174770f7a2275999e68d97c840a0cfae1aeb4fb6
z894ae0c668c848f15cdf870ea17879103130ef4c568a35968a729f4f538d2c4ec69854866e4c5f
z7d558a9de286849bd4e7f469b2d9d35c4109334d88816a4e779422f3870e2fce3177284a162ca0
za28a451401c7259d69546974e1a241d626c3ceccc4fe32776783d308e5604624dc2d8d4b04f053
z49cf8c79b6aa64fa142cf22278ca41565a3cd9f6c3c1372d9c3c1427a614cd26cf4f8e0c91f2fb
ze67ec7c599608ec09700ee644cab9cca562be4cd58d0536ccc13783c23a41b1f559da9865d6965
z398634d8b3ab2e1c085533e7f47c85bc38ed01c6e36128522d7426297d18a3f18f4442b0158536
z8d7c3c0f9e82af632197a58967b4221643874c8d001047b29715e18b7b4968ea0eac6ff39ab594
ze00852a645f7f1f0a1b85c88a5f33f69ce057e860999c8393372b837f057279e3283b462e885f9
z343d2603965d751dd6214486e09ca19df57dc3b750de9895e6199ecba60184a6f2f7d3527a0f5f
zad92f2edc432a04a5cb2955d15c6a7c0c868db0eb675ac28188a4347a381991b98babb488d2722
zd66a8cad4653d3b35c080145cdbadd927d3681224fdf5de03dc6259fa422659fcaaa6a09d77a3c
z98307e17d23b5ed38b8c79f59080ccf23035268d32b3a95ae1dd909a1775a3b152061bb1ceb661
za9de4e9c6d8dd0713a77641ee9938a67cfe82e5b871e11bc8cea987a6812e14977665fc233261c
z17d124a2ebb7ce8b5cb93ef1911d78a4f642b4f46462dddae85e3b6462b8bb883166f9bed7c230
za6a687cef988d07b9f82ed098d16836130885fb0c41571a81fc2e80b6678478636acdc13f80272
z913a3eb83b2d2484d126b570ca169aa5ac34306a7c60077dd9d6d217d2c62ea766a14131ede573
z51679b11cd5f89bc933f6d55d0078fc9fb557e95453ef0da0ab480ffbc1d1c70fc159d20ff28b7
zd50c1a064841193cde9ede038d8e43a6e019e32485376ef0cf1b461d6e96a9e6006b9a69930a37
zb90c270680556f4708239a44dd9e17011797d929342eec958afb3b8dcd1629a6c6a916fdcbf3ed
zc01394278b026f9d260a817a0d2027d4e883b9b98f65ff4d8da7031f700bf8a679c0e2ed3cf397
z1553c1dadd6404a529b562aebe27b7bd5f1c37cce11a12799a69b067aa0f7ddc357b761d6afe2b
z5cd9a07565610e52a372b30d635a4b3fc45100a05a9a73902c0562412c29af9b53ea8484497433
zbd924f3bbd70c99fd21aa73bf764f7928f0468f32aabd49f70456ed4f19431e7be9875280ad734
z05e1ab7ce1f04c928a355c72adaf110dc5b65efe77e7985551311002931ff6c68af9ffc7d4405f
z497178b1c3877a055c8678c42639d93c882bb7ecee80098f1b6c5c8bd0445d069635b9da07a8ad
z8f4174b2163bd2f673913efa8ca099aaebc189d4e6c129a4a4ef5a3d7f6cd16a29b79c73f87ea7
zcc92872b3d1908028b03de1b749be26af64a167656127a5073cb8fb22a01c97d038d64fd110c78
zc777c8ecfe96d252983e6beb2a004e6d964f63d2bf944f39bf80f57ef61b7aa10a71d1db9f3791
z7517cdcbedc8ff015f5ab7302043919effd5da43bd4bc726ebb5496cc05fbd6f27e512735d824d
z4745e9019368757d49e303fd0dc2ad3bbdf7e29b803ae6a08fd6777d74a084f14951fced77d44b
z96aa2baa902bff460265516f8ac20313798996c75f7e8c02330eee3c79bdbd20729ca72c5b47cd
z567873dd0cd86f70562ca603a00a09996ff3a6d2decc24b4d1c85817ac683f56443cc2c67fb39e
z736f0f8cc641f8ecb04522027b30209c151c9d3ee7659da91065258f226915b6849b2ec8b030fe
z2c7f28add24f239094aaf63804eb3905b0abc66286ae17375c47525ed78e7df4348b03defa6eb4
z98106e3f4c18c508af1eeef47f6c60ef8f4cb9694fbaf551d337689dc52d5e30e34d211fcafcec
z69b823f1c96047a22ee008ac1969c26f0a6dc0eb958a4a3630a426bd6efc2e6ad29623a4cd660d
z978275c1caec37770020439fbb4c73ed5432a0d31aabd1ba55aa376779feb8bf14346a061abdf9
z38b4ad8cf7086512aa10a870940ef87ea1a98bdef86ffacebd9caef3f1335ca273637f611914b1
zaa2c1752835eeda559f43088bf9863134a24de079d259fd2a7a1b18a65a1721ae5b53a746dba47
z9620ef0313730f76486e82dd4cad39452dabe7c74af5cd2f6289dd4a1a1c60cc771d9d43d90ebb
z38f7c92cfb09f9656192d902196c4b2f78d2fd802121745966270c8c1b86a54669e1c71aaeb0a8
zf2fbec407c3e497002572eadc220b3ae5700098e53a909d9cc554b73bb928ceb12387ddc0f80ff
z7ee7b6c58450f9a390db0ed63d2bf52a5ac4ef13efc141b340a3bc3503115d9cd8e4e49acc60cb
ze2f687245f5b901980459e25da72aede19680d4c0d32666f4e7867076a0a62880680f7f03d5e39
z91f0897d4688b87cbdf746cca79b31fca7a5d59a8f62ffdc28da6493ddea3bb79009bd6d37b844
zb593ef734b28913f2c8f083a28a3eb236f721a7e2e121458f91dc318ba6485dedc3eba2e87865e
zf0574188fcff27c4d2435fb0f7a33ce846fb3829baf012b77bd1d66ec332421395aed452b9f79f
z469bb0abb616d59dc7b6231671b0ad45434ab0b94c1f7a9daf8e6d8aa9348775b6940196ee54a7
z856aabdec19378073cbe78c8a91cfb10f5ed3224bcdbdb711c4ce55447ac8434fb8552cc094b50
z99a598832b062efd928bb4b8dfb96abaf493c956758653b22fe22863cde56069e87ae01846cb23
zaab7becaa548b8387096acc04536d6c3a569dea218037b056f5fcd8bb3afadf21d4b2899f87296
z7d21f2359acfee19be030c8e043cac2a0e1b4f020f28c6acc996283359f7a9353f4ca329138d72
z352541a09a3aaa3dfe43cd0ca6ba9161b9947de65d89ff6450388a0e628206de05677924381250
z91a40d1f8b7a070474b680ce0807fa9de1517c5c828ca09e4b34e8cddc03de1526a3e86fa0f9b1
za0f81b4bafc68096114b7f6f7b017fc025cfbf29846b3b87800f2d484b5757bdef83abe5cea93d
zbae6e1c48797ab9347b8a2c3ff527faa5748945a38d5770dbb417f7f296fe393156d0b4cf264f5
z3b8cd414a8e6f2e6c540f7e0d2f89e12e3761b2cca9a2a9ab3957925298831315fea0ef9d0c675
zc016884b4065563d78378d597b2d8ba4a122e7194b8e7faa3862d39a9dc06dcbe9e7c686049b1c
z7851aead7cbc79db30ebddece9ec4df627918a76723cdba2b4aebe9afc10a98f4e53343cc0b2e3
zf9886958e9f5e78cefdd7e7791453ddb373aa80923eddaa0ef7c26e075300b15627a286288c73b
z73140578f2f03210e9f86d2819dab44f375091ae1e1187a7f72008957c5fec02f6e7dfdc3fcde3
za8420f6509067b616701ae6f07411edd347d3713c6497f3c45152f3b9e5889c68854c41e7e9967
z118c6ccf9ccc685634851e3c3f27014080c113f6c2683fcbad2b5aa1fc8acf897a4f4858655616
z5c025689f0625bf3eeebfc358afe73ebe7cc93c94afb57e817d70ce62e0360664be2fd8721e527
z21c6b725f9053086a6c14f5bfe91f9f694365b5c318a152c070e66356583dfd6c479bc7a1a7aa3
z61eded5e6e6255dc621bb1c6f1a2249ed340ab865df5a0fe81dc255f70771bb426dc0680697bbc
z512b5c551eee446eb0a6fe111e34d25f07ced388fd4a790c1c74d064f172d7e672d7eb35e2bd0b
z9514322ce367ea36a68627bfca1478ec4770767bbb595e63b97f4a26dd9dae41980eaf10860d71
z4e25110ba371401fbd602b64cfe0c99fffb488089c24869f6eb660cbc456c66f25a73e7f86c78f
z1aff9c64e826b8a0893431048cb1d7f55bfbd58d215104a751f575f1ae36088a69e6260aac2460
zdb33c3cee07ff24bfcc7283c4961648c66ffe849dcab458d6fae4f71e4acc069c2b1d3fc97036e
zdbffc3a5f8d3e43af2dece5a344314934623c93c69434d3a1d0c4db70d129969dd19b4b6a1523d
z19eea115babd5ee47213d010e92cf882851372aafe34f52722749381fe89067fa97cc7ffc26c61
z0a61a0ab4bf2b6ebbaeb50d9e1ac9f7d509e0eeb36b717324419394a0c8f00a2d2349bce9c5021
z78c0abbc859e711a75ecfd21b826326a23432e94dfa766c092f8c765d2edc3e3b8eaa43d6530df
z1d642115bc646051b4458964852f3c74cd60f4f452a16350c7473b74ea67d5126409f54d42c8ac
z20af82d5dc96b1d41dc578d1da90da778e30ac24fc293d9db53e62aad1aa3fd5f6d96427ea6808
z4ff08f7bff0b6f099a5193f240588d9f5ed66ec02d3f7683bc7186ed43188bb277689381f3100a
z8017cb475d8a65a6ac95ff38111903178a9795b710dfd501d422f8968eceec2a280c516f6cd6b3
z8477159ac8c2b88583f0fbabf4418ec69d879fec4403b549735a80c96a8822e7061b6b01bf5a01
zb9c212ac6913cf7e14d620ede4ada88231de76712ed08e2952c52b88ef9dbc65b775e8592148c4
z43c07fc79fb287252a44aafe202b36db7698dbbc8faf2363b381ace98b7275b1d9e0c757db9345
zc525b8c4160eee6d94ef247fdade32459d86eb5e41921447f4b4506d6a16a80f4cdbb9a0650379
zf749828da3989f9b9cf5e82f3cc5142c7eb20caa65404a57fcc7efeea67837b76d2082899004fd
z7e34dd9cc525b021588ac4010b1a46ac1924cf14150f93509233d13100a57c573773be4e9c0eae
zd6bcc9cf247ff7834db7f007b151cea6a394ea91c7bacb5908e01cc9cb0c513e5c8642f312b562
zd9332baafb795a30c3cdc15b51be0b98fadba64ed63d3bfcd9fc8a244df9e3c09261d5ddc8062c
z257de20f0c7349d57abc5177c1a8ad35b763ee9085cec0845d11e5eb8b35a4c172a3c4efafa2bc
z8f43a193992b7974fd600781adfb13b53368fc30e6a1594ca718847401eed3099b6d1c7052bdec
z60f6695662289bbbd566483d00521fb42c63cd79ed0646590f3b20fb71bf4c357a8bcf5956e028
zb23263ccc26ad0ba9a01f80d5efb388e5c14536831ae1b94af81513c38724bca1d6c0c82f367bb
ze0613bfe367647381919ba922c2cffd3d890d0e069c8a4159a182d02f74dfd5ec57acc5751c218
z08644d081e5ef0d33ec4a006dd19854601c6996e57ec64ea2e44e079be7cdbda4303781de5c310
z4b247df272a23161bbcaef2b79a579fcdb4a2152e2500786a5fd63563b191098068679073fb157
z5f35de72a26b2716ab74ec447fbdd81b3d7948ca3a1b627990f0476c7a298a6d62b144787566e8
zfdbc3a320d9e9698c5e44ad554d5d4708493b04748c7e8dd89bb9cbbdd524bfab6e464bb453bd1
z14ca2e473a3c1e2c621285c4394bbfd86cfec49a30eba410a9fed621342f0052dc4983c65741c0
z8891b6ba28aa8965fc31b5a6bead1ed76102f56aff8be202e6a07f460e2b6a803e9228d6a86904
z0a4482126ec9b2bf07d90238de14477b4b6e48c4b8b5e8e73c2318a04553ed3eb65610c8095783
z24edd4504c24baf84afd6e5dbe6c8f503c02768cef1754ca1ecb8e19697dca2de3cceb3eb7b2ff
zc6ade973b8481c36f2ef18f44de1302913a0e533b223f90aaeb0c4885cac981cbd2913384b875e
z7bb9bc0a76a870efb640189f131ae2caf633b8da01c4b5617f6f83c9636215084cafb68a9cf81b
z9002107ceb634376d13b2a71a0ab323bc6d9a50dec94904da4a651f463b1a2d0b9b3db4ae3492e
zabd81ff5aa8d71914e7357d6b073932e44d790bb74a35b83e21f943b4cd2af6d717e390f2c6892
z567073c63e3c2277fe1dbeebf57ea276be439e799ed32740198768f26cd53572555eee3db7551d
z602bbac7c2ec34462476a57e57230d4ef5419ab36b1a340aa58f21d67825b76d3612c7c01cd61c
za91747c4dc33e3c18cfcd0ab3b54d82095a67bae861f229e09a2969db8c1cccf3df70c5b8fbc69
z0cf507d70a110a6aab3c537794168412e8b7d49b654824b4b4e4f2ab99e325bda89e0633d01f21
zee125ae441851d243f927465ea0d04adc9398258c71531b9bd978694fc95caf59b306d1c6eed2e
z099f5c16929107e9e391bd4b8033f8f840eaf3dbd9b5083140f060de1f64d66e33eeea05d86910
ze9a395780ccb841bc8cc3fef496b1e63615419b7fd5ce413fa5e14fbf31f6d7dfdd7435ded3cd7
z6a84e7abf634aae35460e9ac3dbcb3e6a77d89d282ec33c2a121bb0fbd45981453e38949d2ee9a
zc129a19e6242a08eecb692d2f63daa41647654f4171e1dfa86e4d54584490dea39d502590b11ba
z5dc89879898fbebd2b6ab0c19657e332017f3c1e17c978a2a6c7bdeaf2e033f36ec5819c7e1222
z4e2afdd9727d79336d8a193f17ca0ca2d6b1e06e3a05db2db22f8f62c73157ef0fcaf215e97cd3
zf3aff954da31bc3075446a318d88eff45fa81cb1e50391f64826fbe306863be9b9e39010c79402
zcd61bb4dc3eac96887c213a0025b99e9183b1970ad3c6e27a86d89331fe283bd2e82412535d8dd
z09732af651a27ccd7fa9aa5fe584bfcbe9a35117c02de75e4f4c51b168350bcc0e8075d2dc4189
z814f2a674ce837986bd0aa4c733e25d6a9c3e38ecfc50bdd153d12acab3749dc07575c9b52294a
z19edd20505101b58f009f68be7434547c0e48ffc7b207d191c74a0db857705bebb21a520c1320a
z910a2933efa7681259e9628f299b6933aae248345b7285ca706b15740b6e58c3d52d25e0dbaed0
z7535247c268327bd563c7439e66c676e854e33a94a41798a6f70ca6269a236ea4a58bc897a0d2d
z76ac54f23f20d6364361095e8905833a3ed27b47bc7f9d3f1a33ec0250d3977dfbab8fa76454b3
zdffa0a9abb4bf67f3508260a3ed0bc51c2b5809b9b851429b30ceb89edd09e73c667df41f185f6
z556ae8d8d8b86e72a87d4797f80f47d13b3ac30bf2ae79a090fea010ba53198228514fc3c4d3a1
z3746766b63718b4023808f08ad4ad1c4583fd53d80b89c5583a604e30c142590199c9eefa96a27
z8209a2a458fac3c6ec319a08cb5a0f39e7ab11875c8990b431199fa437b0d57d7b9b7124377ad1
z41ef18687b8a4e8bf792ba64e96144cac705dc85fdbfde7fd3cd9873becbff4d7ba99d96a2356d
z731690955c38487a7d46a8eeed84306b33634d3768c9f4cb44c31652c99256955f24e5d7bdc040
zfd41096ca0686d40c86e57ec4c4336ecfb7eeb2a1b4d9ff9a113e3e5502b59f6a6e49af7336173
z468758ef141906e18d26f826383de66526072879181e3a1cc395d447dbed13464fee477639779c
za8a0ab1676c4a882b4669a60293aad7cb569bce17748e816632b02594929a3a4a29d803a88f900
z23eec706bc3b0e93450f98a450ea74bf1bd82fe706d48245486363982c63e14dd5b3e8f5c40ff4
zc6132942370048e6a96634cfd8fd020aee8dc9ccbe87b3334e86eee89b7f1f7826a551fd431139
z7930a21f714e96cec2d23b352bf1d9b0b4eb1c67c521b78466bc31a8b7c37b3d98a0ccb07cae93
z60e719fc91a42fc3b24f030a0319c8befa8cb9d5a16eff0f57f5cded11c4dda06816c49b9a76df
z8b83219a2684977335190efc23db923f3549dc1847141220c7fd72fb3076572b67756dce4cba35
z23fddd649b43306afd86c0e48fdf94d16dad191e732051bb21134f9ed3cd9e83abbed1fbe03cda
z3c98511ed1e83c14b3b691ab28740430251038c2f6f2568213a3a506728b4b4a803d8025a3fbfd
z77c71c10dbeb0d472b9fb1cb11d3e29322faf371bfaa7cc37eae3fc9123f8e75bfd5da12814413
z34badec011f9c285d42cdc802a3e085b2610c7b32d594410815446af7f310f33be8b8e60793d48
z622c42a98ea3f0a42d8fe79a593fec197f82c749212840db97dd5a96323e37007ffd3d4d16a537
zf12efbcfccc4b612e376c78553c5a079ef0b2831a61a813ed0d062be96ba214dfaa17e425009c9
z65ad87518a850ef4f6d75f92833aaa0a2d262ea1516254de2b276c1516c8999516d9795ce67448
zba0fab78d0f7cc7582ed29fb1647e602fe1b4aa40a44acb5a1bd9fbf721a3a5760effade09d6a3
z10f43c2a026ced671f95cdc5198740eaf0323aa21c9de0e810d2badf2dd4b0926757ba0d41ab12
z298a0a75dfa59250905995a92a79b5e5ac851bb505e49f731bad57ea97aa5fa3361dd7ecd84c10
z0fa11c6aa8e3a731435f4f78282a303f10ed74945a3e0adaa72186a96d68daca9ae8104c84a7ab
zc21ce7767bebf2344cc280d91d2938364070f0f174b176e38c6f5398cc4ace1233b3f321468ca2
za8565da1577068296585b8ed99731cf54ea3afffd712f7b89c874c24a213b4dcff44d259886832
z8e4b975565a5f224460afe0156f06ae0ef428ff2d3e115dfe855f439572b0a7305b5b4d1fa2209
za8d766d8e4a7c6acd356375dd38cc471c3121bc34aaaefe2d997b8f145e52b1bbe10ec5aafb090
zba093a44c760a577fe874720dab2ac16d35a346e039d2cefc1c541f312e576dbc9f3d3e9250c2c
z430877927addc1ccc8840690c0270957919e7c085cd44895362b60be85b31db4551946c02b5fd9
z3b3b48c63b7b8d160fb1b70209816173704df3d070f0529b78f3f8f948664096d372d6db785d77
z907c7f09f44212cbe24525e437899b2639bb24642f1bf97536ee252899c3a4c7e1e31b50030c9c
zdf33b2219ea7add6d2672d7711ca864d338c2a19052925a4538dc3dc2f56909e83ad6518090f82
z6132008c9e0cac5716da35e5fccb4e104e0668fe14172a00b16c3a0379d534250a8beeb31ce073
z3d2e998401ee03097655148afea82a31e7727aae74aee29b4f7e5242b86c840ff7e25278e860fe
zdb335b4e0c122e5112a0fe68013f5c259166721299381c1d6427c567d943c3cfdd4c4e7b179bba
ze9b648ac295a6f3f6c446de4472d80b2c31d3050602430044fdfec8fb95c2c37e63f2d12c7c3f7
z54591336ca8ab5c7f8c3982d6e62402d0305b2a3eb1e7a78897abceac78244fde3e1dc4efa9999
z2cfe1a997e1f6d019280dbacdc31a8514d293c9fb055ffe31fc6ab1a1d49923cc2809b82b0ec89
zd472bb99e6c627d9680d55af912dbeb0da0c28ea882b3d2d140e67f59ec58455ddbd7ef2160821
z4386228d2df14ccb67847216d50ee66c81b7c0fa5fe380d81e97c7e9eaa5f182f6c17a320ed745
z9da283dd058d4dbeb19b1cd095b522212d634b8de921f439376d3fcd01434aafad43a18e9a0cfc
zaeff750e039c995f34b4ee15f84d58308ccce22ed9fb6c92f60dcd98768779315260dabb503fc9
z446c848b8a8a89098bddc9c980286853af0213333299fd68ce0f7cacada5d3b2a4a0b58e263d4f
zbd2d4e73717db8c0ff61a657a6bba20bd425b10c3b3c50b6c1ca68b18748f4305eb8dab405f668
za50427e99b6f132001c29fe3ef526e6b3c9a1008dc6595d3c743ceee6bf7d244d43d755d7132e4
zb99b07b80a34cb7cc0f3e974a7d7973771ad75b0fb13d05e3834d83664a26d6784890429323d77
z3091e74bb0c38ce281ec8b9fad97bef2505c27bb7b6729e457d596e5df4dd18d44c9a8fe43a548
z6788521a9287cb0ef4bc3514eab4b3809d2c51b3be152fd8f7c267f87c639c9baeee9630c2f64c
z2d75bae90d6816793ea2d691fc03731f2a3595f4faffecff4187237272c3318abe8c82d4291ea6
ze9f8f58e9f6a94f4ba46478cb540520010359292aa2ae100586f46208f54bdaf49ee9b2abd7093
zbb22ed34002ac4e1a4a1fcd6cee41d51c46172a6b0fe6e72320d776e0c42de1ef3c891dda9b9c6
zf3aedb1567c027725f6a6147c2850613fea58d08670b5623886438834ce37947463b9f251d7716
zde15fef6fb88e88e042433986eec166c1c9651f466b95b20a16a9905aaeed5fa40d3954704e5f0
z2d1045054ed2ad2c6d79439a12b18403ba967bc34de6b806e5d3bc69b72dc91ce9c59858b1d2a3
z44b0fc8b17da17bbcf27de07554dce1a35a37f859ba8a9b268dbad0f417cb4886645b0633ffe58
zfb4b269ebc5c1b6a0b0b4c19a273deb3325eb2fa3eda8d05289581287ae80b5a0e67476b276abd
z9a4134e8c5475bd00148b5d3deccb1e79419b179656c1f8fd37b8c2ccdafe028405043e8193732
z86b0c45c54896bf8b8b9fcff4e7a4df37fa1620491a51e6ade935e36c1702b224fb2fcbc7f8cad
zd19bdb77dd9e87fee2e2de93360756742c2d819d99efe342d4e7272e1dbfa85e54496252378fc7
zb8ab3592974aa87769116c152f28c5193eb630e97d8607637345cfd7b2dc59cb65cd6a2d18897d
za04d2ea8d32a2a8a1c0247c1d2de05f9c74559dd2f94b581a0fd686fb1f47dd198cfcf58311cd0
z376f33d2fc04ceb8617ad445e84f1c8a44fe4d46679ace37581ffa8e5b8a2db5464d7134aa4178
z6960d0af5adb457d4ed93c23f25ea006c6d342ce0d6623d559baca72ea670dfe3d7f01728cfb5f
z8f154e722f50e157adb51beede1534deaac4602c7b8a90b327c95585ff61afda60b26ecb18a343
z39b088921fedde30fca964a68888321f7dc215b1e0b83ca7bd007368a68a3d1f944b78e180e7e0
zae20a2411608c4c8df5e5db63d0a549e009ac7ef1d09272ee72659ddfdeaed4713caa77dde6dfa
zb2e66ceb8397f477147b378f1b39588ddea82e0dc75bc1347430c9be73c921c45777de69ffb555
zc01caf208f4ed962479b87fbeb3035fdc7e43314310cf8dd33c709849395f33cfc3fec11171127
z38c7f769e9b12d2554506d3f65f90f6a9639e1b0e763d4e45fdfac5e5af4f453645f3dddcb9e6c
z64611c71d1468c3da5f3eea124f5d13b9faab92474c5ad3263d572335cb7c36b71fd005a8db4f8
za1ff2009e42c88e735aa6ed543e656de23ad49d3e16a2bb52d17de6eeba73db4d37bc5c75eba83
zfb7f84c2b08f7a7d16bf3fb2c39738fd35be95042da4f82a189e3fcf57a6cef53b23023a3e0e6e
ze17fbb0083344ba283b87251765fe543c73cdee1aad4cb1f506083a124904cfb5ff730bb4443d9
zf3ecc5830ac2c9dbc7a56ffa631215d7009ceac659a044dc2c3396b64f0d79a47f9855c97edebb
z3234f23374303112e1b312c57464b4657806e59da37d5a73b4cbbc416f60a1ac209522be72c085
z3894724b2ca06e65fcf1f06d54fa63cf136b118007ace902e202d6d6152c0170fec014ba252187
z4c04adf768247bb7f1632f86711c4d4b94d2aabf9f7b0b043165d2b25ec9df2bb292d8c60c7116
z70841c81bdf00dc2cecd9bc284bcf092f48aab4eb89208fd72221e59612418049f58e30bddd361
z26030705c9d74c0c1a7439d48942303d2ce9484a2f08013ffcfe391a5ce7c7c832cfcd176289bb
zc592c2847c10bb0d02ddd1ac61b94dc78607bd5d58e00f2f75cf38e63b6470abe1c4bb847996d5
zc20953679a454e24cd783eb0c3dbd7e92aab06cca2f0aabc5973f9abf0f3b50b6d20d2440615a3
z0b348208ab31af8bf5cf971177ed2ec59911679ffa3de7ca317ccf3901eaabe9bc12197138296c
z4648759f85b7159aae92ab611bd7ef7543f4410337c901fa3a697695df6a14e5a7a9c403ed1cc0
z48548cda9c842db12513348232b41485808e84247101ad3973001217b2ed553ea942e83baef9fc
z8e5d08879f5d6160b21343d41224bfd50dc7061177481e43649efe0376eec7ebd00d749f57abfa
zd2ba8538aa3043311c3cffc903430d6de320b96c5bc89cc64ff2b4a37b9288e3bed8e8855aadab
zee890ebd64128dcc428aba5cc50756581bc85b624ac323395075c24d63ef15d07cc7e060226135
z42c4fb5fb91cb3eb45f5293ca7528a724ba7f911bbcfea2b74b3409af99ae33667a49ce087e99f
zec1d51924e0cbc6472bcc864e6bee8c7ef8c3e0e9bcfc4e28e141c22e63c8cb8ef56792f5d15a6
z208c1124d3471bc784b9ba1bb82428449c797801ed263bb3e1468b03aba5a6088b363ac76c752b
z1e9ef5aeb5073a53d69de17579b331bff10ed3dffdecbd376571073f6a9afa2ecc0c551c7538b3
ze4dc1dfaad1becd3516c75b31557abc4153932277cdd159c475b840ed1518c0d477c643c647f31
zfb6ad9b5093621df2901aa8c92f025851fa494f8f094c27ca731a85dcb122110910108dcbdae79
z8a7f581504212fd0d4521f5e677363d1c0290e84bf28bc88b97dea590c90a331b660e78167f2ed
za2444ae621bcb2ca8a025f5e91a825f58d069c2c5f51be43663d51b7ab32dd88e203dcb8873dea
z73d48790ed7e53b7731d428069cd158760db5992fccefdefd929379ddc0a661e8886cd4ef06ccc
zedc12c6772cd8848c905e753e0ae9491ecb0763c74041570f9c0a1ab6d474a2b2bea3c95a1ac34
zf3d7aaefc632602b12ab36b79c17ba22daebca8c3057e1276d7e2ae25919ff8eb8a2f97c008f46
z38d5a2101bb4e9bdceffeba7f33a055ea23536fdbe600713cc600c17896499bd3eb5272f4f94c9
z73377d28917d7e30f18974bb429a7df8eb4ecb7409bf5af9615908f6e907809998ee0c1960a7ee
z1b3034dbb2658f757fcc9e95b926f629347f5478cc97ea2c92552077b8f0f0c7402c5dbf3e8382
z7194397f9d26265312a8446709a0b69c447dad8b9ce6f16f271ce345a15451c1f434e457a04d3e
ze6f926b460242bc43268d6aaf1cbf60ab5bab33dbcd3d74bfa92190c1a2d2d58917e3d17cf63b5
zceca1f4db7ecb58a9342cf7bba7fa5fe6e56da52378f5153d6bae9803823c8a148bf6a8af316fc
z5769b344a9a0f4fc9737d13e8454f1cffbcd76527b74218f6034b152b42afb0839a1dd4d5a550d
z406104d7ed68c310707ca9fd12d0a866a3d425f9e1b274999bcfc0195e32a48cb441fffcd642da
z19b71e11c42b7cf8fde96072440102a12ea8ad99a1dc460d08094f091b3d61988a44c151aee6f2
z98f034fb6d8c2239076248b9c620d3960b8525d50622bee328b6fe1338117c2994c63668ff4cf2
z5f00a29d497c470142f7f7c4d5deca62c0a40e08ac7eff971ad6a61d429947f67cd963caaf6cc6
z13fcb61978be6a7b70942b419dae8574316960e6d196a90f78511cdf25e77e4520b235eb6cfa7d
z470f737c684288033fb64fb945d8ad18d59d41197f3e283b30633025595b52b405229e7b66ebc9
zb6ab067754850c4677dedac147f05c16625a29d30a2990b45e90776decfa03224d051063f229b2
z81e60e0eb831e97d791b75a9609387def4acdb0101038550919562f06dc7bcacf40567b43aff81
z6902ec534cdd438a61e6342106cad94d75430bc597c5d51340424fa4d663a63dd8082324434fdb
zb25185f77e23b92f343343f465cb864333cebb5e6aff3e89d218234c81ff5e589763ec7d81a99b
zaf5ea1ee2ae3e02eb42d1a24771106d69d528a2abd7861f729f5714f68c501a68b50f27e5b8d58
z7714d3d21193c5a5f310dc7ae915fd97c6ee939c7c15a7e29f97d1caa62fe21c818add721e7df1
z445be810926149f1f589ee749030174f7b92b27b0f49f35e324e9402471a0c9b596cd9ed96fe43
zebfbf4cc7680ec74605524c6a823673238ec5187f1f61481e0956cb36cafd4802d37da812bd2b6
za7f78a164bb84f2144c996119197ebfd82701b6b16d6dfe6d4c73a174a53ac65423bf65857ac23
z6c895486294b602cb089072a188a412fe21ad6f6d44a558655ccc6fdae381ba8ede3455d52a98f
za361d49e714f3a3c955213ed22f011f06d21f10beac0e0c043185b7e4b676064eee3ff799e06ea
zff5ba493e0d1d2c49ded3aeb9b4ef7b485830a4e90e9c8200be8482797703294e847e323acafe1
zb6b964ddb0288723fa5971dd6c3ff66f11e03b7093a5d219fd61f54289cb81f552415e3470f55b
z22eced5ae4f9fcf7fa107f0d579e482851af593cf859abdbd83aa6f56e4502d54ea2a886b47617
zad8c69e7d74c491683a964c8740bf5becc41b46cf887b707f19fc1ff3b20249109aece26338679
zaf0c8c84067186ec05c9e774ea4c5fa873c7863d07bbe1e033d7d5ba79dead7c5f8a9d3d0e71bc
zd35a69d7a00c28c5ac16ecafceca4b2ce56dff960edb07ffd723b2f44f463508b4ce06b359270f
z772bb34a46fdf2f8c1145cede6aa157b5e38585f5198cbafa80417036f6288abfa84bac238abfc
z7371dfaba331e9686df38d7cce10582cf5e497690d8bb710734c63337b298cbf23ebe4b7f91c60
zc4da8b0d5276115ec635194b865be2ea4add0b2eeb1835fa92096a6f785a80bc3094271a4c1e8a
z71aeb2cfdc44168478b8660bbcbee4626ff30703ecd7c8f13b3cee233b44bc54bc5108caa0e6b7
z356836ce9180cba709973c923b59c4974e4828c3990e0b0e96b2ae66415b0c7a94288e35069eb4
z8cbbe80e665a415d515312ec3b78fdffef03317f746af8b7ce70fa1ee1b4d8fb84b50bd7df80a8
z2bc08e2c9ea5f7537c94f89fb8b7e9d6cb716eb82098d56d5452982c938558c113b4fbb4024e7c
z17db44f33d192ae8034b46eb0940f063e7238e6a8817dae5d15dd25f09c72f647b1b761ceb911f
z1051164a74cd4165e26a1578ad0420e43980320cf0336cef2a3fd5e25578a476a5a12c87603f3c
z3993bb9fd5ba1f32caa39df4afe11784ad7a778400966f5cb97c81c051ae03bb799379a4653b7e
z95b80088606eb4364d7db15c2237f84b313ca2c22d62cc3be582530f75d6699c22b5fcb817a222
z6f2d5d13e1dff285676e1d0c5aaca51d2a7d1e85b96b970fcbbd7d4dcf5530b7396a249d2c2d7f
zee6fba9c62165b3073918a3a79bba32e46c87cdcc610ce14d7b7e7bc7e93d6bc55b6576606cae1
zcb3e44721717f8ae3b256ba48c90b3137d1fdb0b9c9244096d46e7c58ccb2094b254f4152d8c84
z11bdd103d6006935e33d540225afdd504f65b1acf327990a370d45317952cb8ab28f6a733b26b4
z324ae25af2b5f2093427a50eb8e6b0025115e214cb8d76be1a2e36097b3da9cb0f1cfb4f31f6c6
z3f192624f21e6833f07b4be10f6b4aaf9718d8d93dfbb8a974058bd0b7ebfa6285dde287bc414d
z363d3005914837b8e5bf92be0231acd6d02ee5ee69f053a8edaaa223991104db2301fe8ae8969a
z74ce739cdbf770cb7f9e5ba8f95d76fdc0e538d49935e4927a6525b28299c9723bc79c8e23c722
zf66d26c6a268641adb40145d7602322943172dac0aa7400e162b331e2ed4b1b5058054c35fd309
z3541c6f54c43024a439a22ff4c5d5b629405b3856e165125fc5a2e3f85e5b2c0452fdfc56bdee1
ze554396f380e77148bfffe4b0fef0dbd25521bb74e046bdb3a1f048536935d3886a0e1845775df
z67fcca6263a104a3a39494f0841b5c794608d5b2099ac4d33fe7509fd33be71695e71a7150201e
z8e0d4d137db3e64f24dd39ee8747f081b99a77e67fdbf0a963167c0da0b9e97a8ca335a79f34f0
zea14e362fa4d49ac8ca8811615c4b0e27275dc413862693c511ecb17e7a34904e3ffbb096b217e
z5d895e0526826ebbee9b660416d89d41e1cafff0af0e544076ca1eb4b02b4ee8fc10fda8a8e575
z0d86d535e231b2ddafaeae579148138934abd8b59b66c9a037cc1f0adc822f94f01d8f9aed3589
z7b4b474e13b2fd6439476f3231a1e2deadc4c39da96773e5436c33101d6a74a482d2c800ee7552
z4d4f545f1fa0700ef9d7a1da3fdf41acfe30e7cc155b710690d23cd920009524bcc2a86affc4f1
z743f07e9b8ec8b647bfd747b01e914dc5728a4f96be02613da74d383226099be48f0d0c1bcf836
z897408c03e2869143c89f2879d6e3f846db55e08444f83b4c6f56e3b53b28b92ee857d7490ff00
zcdba37c52940fb70d8f01a20a036751bb8b3d2f8c80ad162bbe5cbad214a034685e771756701fc
z81cfd8fe6fc73b97761ed4a3d04558674586f38d9225920b806a18d8f7e6034bbc6da8fa9f421d
z0e08fae14066a9cfa4ac44e8002e2608f7e331a40157af658dc08d296c5eb8d1e08b2ff559ffe8
z190cf15e3292e5f1b87da326ad5589e42efb98e1a26d8a4d8d2a9bb514d5b726a3406c4226c28c
z12471e168bc91902228ff6893becf18fdffdc5170c24a0d5cd59f15e0e35bb589362349dc18c75
z3dca4260a37def692f6fc5e8f46e8071a0968604db4595324b9b55cca9d173261a9676ab4ddb7e
z9f65888636194b342b05faf8371238bf1cdc7a20eee9e75e6144be2cf5af331678d196334054bd
z21dbb7cfb1421f9554ad907cef50760236d0831f99a26a7f8e9ca62219bda3bb80b0cc5e54a2f4
z86601e400becade29143678c45afe334f99ba6a076231fa9969a7f6b69d05d2e551c7422b77be9
z9140c7013e2cd9e08d08426e9d8c496acf0154fe25c62a7bf43ec2883632c3c89ed2e2d22271af
z8097042c8612fc7ddfa746b165b9c9a61416278c20ad5e85a6adc50e28445da6e8d713d19e6a78
zb645c9fea2b13d11a681d296162f956a928bb1726a115d40bc39150b689daf3f69f8196825cf6a
zef304564408aa7c7425e5515d39c4085448715f9b086c6af5c1e49093da5050776389d82eb9dbf
z7816ef519785a1ae39bb7029fe1c6cce1db749833af7b3eb7149d97483d1ae4bbf9f8e184fdfe1
z1d267d58a95a2d055cf6bafba0ce1f41d7eecbbf9dc853c7f33fe31de34f148b75dc64056d8773
z3cd3b1c060d742b8fd73459cfcf66c7fefbed01bd1f65f87d28c5f8bbc59a63b4d69441b330b9a
z79c772d5436c4def473d6c3ae0d219ee034b80fda78135df69b85cb8d6ac28d31e33e1035917be
z82d07ce54519f6dd3814a448d78f115083644e3ebf3960aed87523dde40fd953596dce31335f4a
z9cfb090add3c7602bdd8983374595c0bab4ca155695c5b29ae20feabfb6807499fd54d039fe8ad
z21086b4c201d2475c21725ef64d7639b218fd1b56ee0c646a4e3259d5833aacf172d638fad69bf
z7d52defab3bbe117ef2c5ad88af161f445145ec36baaa41d6813ed573e1cce1a18a16aed347580
zacc93abaf96ae98431f332d2bddbc1b3253d9bfaf7dcd96b11cc71767cdf1da8ac30aa6f1b2012
z65cb3479255bfebc9a108859602a398e4eb829ce051fdc51e705566cba94a60cb1763d8017830f
zb8aba09448937bcef1e0e2a68f776a18e759d825221187badf69c51ee8c22acb792b2793bc3f7b
za43ba65a8cdaf6b88c3c2bf9a29a666808ceaca4473cf4aefdd0fdab2216417c6ff35cf4b90edb
z634ccce12bb3f30a21938370d138b26c3d8e993d0a79e52d2b4875dc12e47553d228a439e4e01b
z75a818b6ecc8d936752833b2093aaf773dd40fe3636610164e424fdcaa77250433c60ec0c58612
z017eb5517f52190840683f98cbc030a5be0a30a65c8919fa1d9dbf25dc8daff60cfb2ef11500c1
ze952c1d57f0ecc9566a4d202a7e6d89f0e182fea9c828e8b85d2ee2bc5a1b711a4d85f6d537075
z1ccc4e86438925ae86d48eba4deb19199f5ac7f677d942e2f553363ff57f3f0f2c74ff3d98b6ab
z31eb16fb5fcb72cab4dddce05e6237c1e85c374ee8f105ce79eb887a31884748f4ad1162ecc330
z9830073378a9c8fba63fe9ba20199cf8d27bc485fabfeccbfcc120ac53b721d2b6a90f1162eeb1
z80bea6b5c9c9ba3a6fbeecb9f55906f37ff0afc628adbba5e8c16cb9c3d8b70ce4631e538942ca
zd4e3e1433d3224e25f766816ae9922fb268ef34958b399f2cba9602ce05f58c8bd73d4b61b06d8
z45ca496521dca530b504598800ea6b05110853d062eab13127777227242cd80185b6526bd8862c
zbb862fa7ff975174dfecbeace6a2c062c2595f779351abf1ab1272dd0175291080b26e921ec282
z60d83a7add83e4c331644a8176e57d84412b915dd7af1194002707812c3e72226b6ddb29e2ddb3
z402c221433856e98d735db728ee8c0993bb2f9bb5a3124fdb5dce858c0ffe858a2e02474c82216
zdb9bf8f185d07c9d14091b475146f5ef2accdd42373f67409b46a7ca0572366954fd47b4c87025
z1871186e391cf2c33d7ec5aa82449bbdab5595153d31ee2960ecca11f04e74a51a8560146732f8
z60745300755b2d8f1a11456b106de00c36cc876e5c677a0df23ab0d5a3ce5bcd22b073ab762747
z87dd65811f912dce0add5b530eb10db8047278f0f021b3e13ede01c3bb65defa01752929dde22f
z0e91a032c7ba205a4ba459052b2366877256d9b7aebd320f7c33ea7358ee4e75fedef71680b00e
zdb3729fd4784411204df4eff1775604ed6b7dde2fb999fbe5b0d47601cbc563113c0b268db7012
z19f55fd992800f60b885dbf4ce39ef6ff302767a3ed6c36c98be279143503fc874d976441c1d98
z1ccb0141e0649a11fc40635e531326e25b479830d4f183e8eefd900bee5b0c86f696651de9505a
z899e65e9ef7643acd70b578126b36d7a001998902c115aa8adcc07b69997304ef2ad90b0ecd22c
z9e1919c36f0475642d8c7fbd8bef7c4182683036eee828c7806f661ac5d0590a397042b89725bd
z73a267a2ab2e65adac8b6af2926c86425e8970b1bb78c59b2f43258dfd00c1e0310a387f0805ba
zb2432ca380247cca56c22ac3ea20beded8ce1de57c10278f7aca5f3035b573f3510172bce07782
z20ff77a8a63049e5068447362ddd9c75803cf824a9b0fb425bd2d4e0d57c37ac6f1d0aa70d90d6
zafde662b0cfec3562ef26d779d00c7aec4588ca750bc447cdcb80215b929fb2bae4c78189e23f0
zab9cd9bc62c863cf1e04797faf428729bdd58a6604243bd893e5eef4fe29e82f2c3a428f588fac
z47ef3f9b75704063cbd5710c87597d4182b42debe565af90c8f7847d801129b240ce9d42ff3843
ze8e6381ed8e96b3dee5025259aff4b862e529045d40243bed948f36f176626f28141b455b31c67
z05be3fbb746c51ed293231aa000701a65aa3f8ca68cdb9c4f34ec403f843e5e063ac2cefce26c6
zeca981d60ffd5b5b2ca9b070f1befa5443ee81c49344aba2da56bd01b211398d543f31be4fd57c
z17d7626b6059780623b541d6409abc748541c84e2508bf555e67f0f5639ee442e82cd0c3afa07c
z39ed4dd2e15159619575b4a4ae93af9cf2a807e561aaa4a778402483779056c6034c77ede8a34b
z45f549fc63366d72b87e67da091105d80ac62857eda185b59067fa6ad9b90ac60240f0e70e2d3e
z941cacbf4752fe69a0c3aa0488f9fc4b9b200497abea57455bc1ed8c6b6f0657e3974bff6057cc
z61e2987885ca8381517609143a5c1007a30b79e5185ce45a46dc516fe82933318ecd1e766f359a
z3c84d5e17e24f273eb9e91bab5482475b86288bf3c567dbe351c70f326e21d579d3fd8fc0b829d
zc6fdfb89dd0c17274663485104ed3f48e02cc0284b4c7f3815da5729da890a2e1f8effbb72b8f3
z60135d702d4142e1672a71dfe3d10cde3e42f79b82fd4f15044c5e216264a72093c9c1a12b3eca
z68a55b097625aa18ea1cf0daba770ae43125540d6a47800879945e39ed1e3824ff9e82d9fe969e
zfeea44bc2cc94196ea18af7bcffa50cccda3e239829520aa7e655cc514335c2ad205229d7ded98
z573714d9b8edaed5d7291515425cbecb7bf496632f888401765215ad1e0bc539473190991c7a86
zc8543947af9c2e4b8d82af327fcdceb5bb5785a7e0a16e6e03472064eef0ef6c5e657b81650b4f
z4cd340f453bf8aad1fe1d8e4812e46909d5ce69af2c09c96acd3ce9294840bf6d4214d683b2d65
zb0dd24e4da8af625af494935157df9a57953bca6049d6959352e505b5986944e4af73a11feae29
zfbedc519699f0be5ebcd427a55fba14d61212304e53d2c80ce1041e2887eec43a9599f51c06cbd
zbd37e77bd9ce7561dd9a6bd21be66e04c87d707f744c7e26e0631a7bea374f7371c942592544e2
z6f4e82a2aa7f33877ae59b90bd019eba2f8344308739d9897afcd1e7b3fac5daaeb0a9bf014240
z003683d0bc1e82f736f0ca934cbe4969a674bafee97a835ec55354cbaf77ac3c99083407d056d7
z0f294eed14f53090ea68b54eda43bbb8c007fbd40ba29846c937c4bc85597abb71721c7e799678
z2a528c170d742f4dfafe85d8e85a08d93e282d683477fd41fd28edf20e7d59b00edf5adf8918a0
zc91948010412bf6da9517c6a25d15e5a265b30b2cf469556501c619fa640009cdc5014d9835606
zcbc56b30c2398b1b120d69da034431df17dacb34634d6ca40e79be0e455073162c330cfd88bc30
z60745dfac05b1a8c3239a3e1575f740b9a7038042e53fe1a3de1aba9e1af8aafd88cc0c19ed4d6
z79b6965e65d75f8c2945fdf5e79d9fad6e1c4e1ec42fa90f2e66b675d2628acabbb627dbb8e6bb
z0dc1c17d95fcb9b3d53cccae7c8164461c92db0d64ad3eb854bc04d6db33d7d77cc8b315458e09
z3a7943f17c6a33b7f7c96f3562e34ece10721eaae2573c5ac7cb9ad493cd9f604bd4dda0aa12eb
zaa06a9464ffa2fdfd1019273beac6eb87ff6bb0189e345c327e00137f682e9175e92707aefdb31
z3c794bb0ea2611aa8f428e16cb8df97b1b3f4f524117f5ebf142f8d761f354f0f600fb4c5e2ea0
z058e6f89465a9070388a15ac260026ac23e9471403552ea63cdb2cb5be0cdf0ffed5ded69f6c8c
zf54faaad7216f9be6f530c3a2869f216e2b418b16f2127152fee06bbc7b2220d66fae681e564b9
zc9cce5f4e2cee9b1987fe6af35297f032e664fe7ea2a12a49c84d19c1adf9f42bb4343ad979acf
z54be7ed9a650cd54ae7d1c1ef51535f88032e6078dbaeb98f71a4db9ad54aacdf6b1d24158ff47
z2d4453bcd00d2dc45333179bdca44ce4c6fef8c3f651a11d6d17ed93abb1808594827453c6dc9c
za4719cb8ca66104df7d4aa9f2c9f87eef3361e6a58a0cfaccf7c610ab2de3e2c94c75c02208033
zc419daccf686c4a1c8b254f0f50655c035f0869dc206e1d994beda7dce28ba6a5e86a176ccad87
z59ee354460b8a722fdffa1dce935bf066111b7bbf10ed282085c72b41823d6d4481f8b57877775
z7455ea0c5f0b88e39d5ed1475a6f278abca322a3c9757b8f588527d2e91c7d05cda04af25f53c6
za9982e61a4982e9f95792bbef01da7cb241fdc9008dbb35fc152cb0f0ff6b494db566e5e5d4513
zd7b6220b5577e2b76da83462b2dccb034663e9777dc8ce0526e09ec101e354af17fb78cbe15789
z20a610fb5de5350243c573ce8c292480c1db45e254ab09c2c0009501e393c37332166b17074d89
z7bfba2180ff94a22f041a8f9974818199d650b63be77a2189c01c702cd83f281d1923dc2a34eb3
zb3416be48b49d8d0223ca28fe501446d8bb99c40de2bfa68ce60ab5762760db1661795e7ca1135
z7b207d866ea9f68a996330b590717c41779eeddd3107648cd8f327ddc09ccaec88f57fc7f154d8
z49e355d9b95e25ba7a30f9a3943151d04d6cf2eb9ce344828fcb9579f604adaa065b4ebd955178
z8895493fdae9313de2b8d3f7e9acedf8c4c809cda0f6638545df8c2ccaf211ed8159575bfb201f
zd31fe93801e7c1f75be298e3602835bcc86f4805b46557776fd132dfcf6c500fe7764ee9370ca0
zd87bb1c4e772771877dc98d4c264388964f09343b3c8744ab9752107aad0a808069fef9b87889a
zbf1f2887916d04a5ed62156a6704232a2278c9c503e19e37bea3c77daf893e35b767e37b5a5f50
z088bd55b78d74e7ac925896c8ccf2cdc40e0347fd08c28dbfabaa8b9c8276f8e80cc4b55374c6a
z0b98d7d52d69c5292c2c9242726a3ab937103fa983489bc9fb2bd72709c3efb7c9c24bf5b0f468
z145df8ea0db95747df5ebc20f13e6dcbfa834c56433f3014ad4534a9e223a477a5526ba07bb30e
z8018bc9d5e366f96cf1508a2c4d361e6a32739d000483238cc728829dc495589a81a4f355dda47
zae3a988b2c74bcc415d117dcbbecbd974c2a14c93af9726ed628f0288dbd44348624498bf1bb5c
z333695b2fb16ec92fffaad2d67e184a8151cbb19ce53e71384295770c07cc3122a4fce188e33cf
zba2068102589502d72802f1f8bacf6028de761104550dd3ff0a700be7b1e183ecb86e376512ab0
z9303eb1a61f115c2a8a0edf5d59affe488040fe7355cc5d68231cfb1c937a93913cc9ec15c2825
z4d077cfc59958f4c55d1c294a13068564fec7776e49370db102c50d2ab9bbba44ee2e868517241
z1656bfbcfd20249840893ca3cd1bc521685707480b8f5324e3e82d41fe0e5e16af9ae612e31f67
z7b06f8d1b161720ca17e6e8bc8affc39d56f20aad0ae8b176f19be14fcbf8a488501c261010b6f
z173195194c21a69dd4e015b4d0f1fea4c025f8328edf9bcc076f874f44247b8d1ac03064d94ccb
ze3a9e52d5c246b5ab550082c2018255a39809013e74629727552aa7d2824a7005538744ffb7462
z0eb44f012470e0194896ab239ed2f3f057687dcf257ec69397dbf589b26cd234a03d5cd3e2b96d
z0036871f67a9ecff23df85d93c879481c4bd85431305fb6b25b0557abd46e9dfe6fe833c190680
z6787750da6afceca0d2660b93ae2a279e27b48f4e4d256f968e1b298ee6bd3c668d12731e39f65
zb979bb29605f85ad0d9635aa8f424ea6d9f1adee1c52e7fe39d96a5a7e4fdbf506c3393a30d052
z90e7741fe6add16a278ea2a66e0de6f4543f9a4365c5d33303266ad7ad7dd2f8ee3f9b60bb24f4
z083eae60e034d680f82225980758c9cf7056e5865c3dd4d3bdbc559c806c12c82b3c44d6fb22dc
zd40ca0090b58c1e3f3fc8ea6ab331116111f55f015c9b557167ba30b6483838c3cc76e2167b372
zbaefd57aba3419ee3c3d97e57372514e1720553754ae35dfeb61c05ffe06e6b56565e66b0b0d44
z8c2ec4222c342dd1bd6f22b9aabcf4e0ecfa1fbe084fc46556b91eab0329eed6b5845a33166bb9
z2ea6d30e12ee8779e481b7be997b7a485a27718b5169c0931ca69cbf0454f7d4de0d45daba7d06
zaf332f0b730f0507a4a497a9b338ff5f38dfd40181721c40c0dee92fe0c72febcf5598c94c0b73
z20353adf4c205643c6c52f13710abf257031157ca0ad7ba63958d18daed7c017ed26815b49f726
za7f4f7e530c596d6c7fe7c256a81ab80d1110afd42efc28a9c8f3fe8454323e6cbac9d5e61a9b8
z3fa6ef8d3769f621b278e0358c4e7cef58c162259c3310660ca9163abd62eb96d95dc227c8d04e
zc7abb17ddd587abf223d9cc325a9727c9e63c9361bd5377d8cb3b2599913248c4983d910cd2a7e
z887a364990c5968ed0b5701eb90a46e81e4b02af1b70f0e86631cee8e6c3d6f7c311b1c3c13eae
zb89f9e184dea4a1b41db450e53bc5bfaa66e29abaca854a165b8e7fc8365df0955bb067055a2ff
z3f5407c969b05c89dc486bb5b190e8cd5bd7fe7c1e743262f2441c65a3651563c260bfd05a16b9
zf0ad13a08208bd22611cefc4f0b3b767826d32b3f86e5b0e637d7348d9393a9a03f135b0846f3b
z057a23d97e1bb63e0548e44c9f553a05dd5bc9323e72e560db894139f65ee5d2e7eb6056f893de
zb5da176e4b3e2f34f4459ed8f27261d465159c04024af3380d718ac7901ecbb17132985a1eff6f
z34e3ba837817f0d6c5e2d9cd828df12455dfd0cc886cf8d86ec1c8e392438bed84062c4fc60f85
zb26a417bfe19666a0a664d6f9a4537249318419a648de9c82d9b08ae7cdff20557d342cec95fe9
z467e170554b515b880f6b36859c7e78bc0778e73fe972e2911025c73bf8627ed89dd1d26d89da4
z8582646072b1ae9c35a764f13096acdf119dcb1e03705cb9859ec25c34ce23cbb4b1d25be2dc73
z07adf4c83b1f9262e6d18344617b0e83c9c1570eeb56ed3599212177ff0989d17577d9655d8644
zf422cd5920bb86ff3a153cf9b59d976edd92c6777f767b8f3dc2184066a51d87a429a11b5ed873
z69a3da12055c18773831fc02477e74cd32dff7ca2780c3047e66d14d9c3eaf0267f1f4941a9a46
zc9b83f4a0f03b125624da9e20770e584bcc75a996d08c2e45dedeaf1207d8418e88a01454de840
z81406fdd34e1edc80f33fe655d08ead1cb8e65fe1421c9244afbbcfa42b40486dc8b39f84778cc
zd7b5503a9b2ad7baf7c5b02e80e84401c768e2765153cc8924ffa1d1ea1e40425303b160f4f98e
z7d1980e5db9a197e5683166e2681c0d5812cf148280ada709fc2dde49cfdb18a8754ab4c6b31d8
zcc77587815bf764cbff86507fc0f14b00762d39b93771ec632ef2832a5bf4ac1cc1f6a86139a42
z80296f16b62ffac4e093e67189897c93bcefa8a18a184ef7bcaf11f1c1fba0272cf86ceb601cc2
z3b9ed2f2415341b06a7d5a946fb7d25c7068b0db1323c24dadfc1708c688422262fcfc9f66c748
zeb41b459ab2f87d2fd88f11757de51692fb477924d312524cf4373fbde42e26237a7b087fafbab
zae22dcfb6bf18b54010de7f9f88f1cd7d040a288f487d0dfc19fa6c3a6671b9b0f54f337352c84
z33d6896198f462838fb842a186084d41c091d8a77abc63f28f62372f25f2d4adc6098fe7e8068a
za45fcda4bf1db848efa6b9c378bf9c8d4c324292e933b8d3110870a1e7f44fd9d0f436faace807
z28ce621d44509d259110400bfc31890ca04f7cf59a0d3fe430daf82c5806d514c45cefd642019d
z73d4187e9fe1cbfb62fae7da9e3a7f3afa34b3b0ce0ba8bed90bf1b7adaf056135c2d5134b1d34
zd45a2453e90ba38f3faf7dad0cfecfc19f3c4e6b2607d795b7ad55b3a36ac0ad45ce488b62987c
z53e875b0bce70a88100bd2d10e9235cf0a44e5dc216b98362aeb3da716d0998e2a9a6f3eabba1d
z9ca9342758ecb211b9906bd5698e045fbb812a820663974fc0cf78b9a39ca4a8fff93095718586
zb772e2724a1c5f7b6debe34d7e1ac7c5a7672dcc285528b76caa0a5fb8250f6d9569f6a3d0a90d
z501fac806428a3925abae1a4672ab5d59b4c778da45eacce3b6a39b745f9b867ea202d2282dbd5
z0bea1eda02a157162abc7b581cd28b574d76158a7676167f398a2d3b0e9c39b896a296abb362d8
zf0f7242c6096f5ff5ee5fe3e5a3c727294938d6e3cac79ceb0a8f641a878d722637e53e3b86262
z43c78f7ade46f4b36d3106d9b8e9b220c5fc116762d7eb5d870b8f6376641b43bbf0db7379e03a
z1f056cdcbda309f35eaed2d1bd22a5df94a48875d98225b8bd2f272cbe48c5613db90c10e2fff2
z49ba0bb0d92d27e562faa17301dc9b2dc253f5fd3cdf77ee5a9c5d225373546b27af0f02ec8e8f
za9e90cc76508ab67ae98a549bbb0259dcbc6e6386e48c598afedef58ba818e9142e4ee7190e363
z3edf8dbce3062221013afe62bfff0a564a34bcf375b7f73b0a771d487df0f6254fc17257e950fc
zcefdad9fb76ff0f0687b17edeb21003bb8e8e9e4bbdb54fd768f9c4dba0014e20e29980a063d60
z861edbe35e5475d0c67bcf1df858c9771e9703598787c428b842521c2fbbe290b53a68e2707161
z0aeaa81f3bac31e38267a556aa8877d476a3dbaaa5237cd367c81cf63357fe440be66cb0a8dee1
z3b49fd364c7ba097968480f9b3bc22baa0c5ec46ca735fae0f6e2f98f9d780ba51df13c6c6519e
zc027dacd72fa0b22182ef6e162cdb872b4674713519a0474e8b9168d5a81096e6d90f6e9278867
zd3d0501bfa6eb0879285acbf79e8fc99f66303fddde8772829625d5fbb270c29afce48d4b0246a
z0b8a45e4c825618bf14159d61abd59f0614175d5d7d6989f8915390f5be9976d85849826f0230f
zc4fcbba73a79e224488220e61eabc30377b81b0314f59a61750ba2e2abd3428149202332b2491c
zfc8cf6697a15a8453f84f9f99edc1eb318833528cd2ff400805db3e82d654ec38a130cafb9748e
z6e6cd11d0063e6bed4813532c77714301bf575d9237f89ee2548c4024e41665643a2b63139a936
z1c98019b93a4330255fbd9bc166926103a7856732c381817d78de2b43a033eae9661d5a074fe5e
z9912e6eed2de87257ca2ac0261ce9b207aa6fd5575bde45a16a914eec933b164d3bd466b5b5001
zc416aa8c5afeceb84a6715100df5b8f04bd93be495b94e0d7eff9bfb1af2c54368edbc620c7a2a
zef2abdd9e4428c1c905b78b3c5da9993822797f8ad9967315cc8ba2263e83f2a4701eadcabfc45
z34fc71331c01ee4e103efcc4e9601506991e95d7b37f4a05ac136447217afd2f49a5fc7cf472bd
za6e0475338cedb219d77ca6ed05d80b084dfedccec6cb295accbd82e8372365551822e007bc7db
ze6bf5e3bf6200eb592d8c35aa014fbcab0de562ea68977569be66977f0565ac85ee887b4288e94
zfaaa2da1fdcbeeccee30358eca00308c2286be549cabace269638f1128546c58d9e8901531c985
z7b3b3a1cb328fce02df1ccbdea43ef383760ed9c345296901553efd64227ea913b2bda286aa814
z1f858c6924058f878347d48b87ec77a44f5e08ec2c00890779a1f68387f7aca286354bf90f67a5
z126c06f00b7cf026a21e8d63915a1f91c62d02f7283dbaadf1d49408068fe4b97af7ed37b10e68
ze6534b0af614ffb4e765b097e37b5ba73d13ff5b2bbec4a948e1b5809b05b5b064fe92cfef0ecc
zf463028514befbeb1f9324c0eb1ae8fc20c76e858e9e91cf751bb899ae7056c689bdeee0cb9929
z687dcac31d9647116318524ede970b2a38380ee4d27b2842912ec7bd921e6acda438e082d16ce7
zf035424b54d44d97ed7b51b3cc9407c2ef14cddcb44e2c1025ed0b3be7bd673ccfd97e8f75e5e8
z9027204a1da140c583d425e3883579fa477ce4dcd8f7aae555674c5d277366425e3978a3ceb364
z3cd18c232b51df88250bf1cf166513f47511943d4a41bfe8cc480f27d5c907ce3b737b8009d869
zca2e61463ea326148b46ba6bbf6f40a5b9c232f5c08a4aad8c388cbaaad4c16e9119781a17510d
z17bbc8bd739c295147c8a400bfefdeecebfaec218afc8877a38ac8098ed6546b788b8fbfab498d
z3bc01b175074c0bc0dfbe3ba316db0f3f603e69a3043576af3796872ef580b06e411d498f0c843
z4634d5272d413fda230307e92be4c7ea363eba32f6552499057df10afde48cd1fcef0e09bdd2cd
z9733220f7dec2afc9b60e1ea65b65c6f72ea50058703f891adada2cccb2a696ab6e4447b9541bc
z119a77f076b053655037345825214a1f16bda35eee0b6a0b32d46ce8c0ff9ca0d81b2a3478dc69
zd67d53b4fe0592461908ba91b0184ef7f5a55e0afd44920f6a3d4ed51284428187b8ba5d5cef68
z0431ec3f677a086d06c4ac17078f57c4c35d0955e0f1ff86e8044fb3588f3dc6ff3283070a9dcd
z5dbe075a97e4e21a4935596677e8f752d379a6ba762f702e47fd829efcdacb1c432f68796045b0
z6d15c58ebc582b36be0aa3c48ffab90a0a2b8dd3861f00fd7a0a3afd0127425410bc378c5f9532
z75fbc15db99fade2ee3a2b06271ae4b7f9b25411663b7f5782930aab578a25f9f9d2d0d183f6b8
z5976d854de101a6618e5bb740ee8a34aafca0fde0dc997c27b0db3a7dff3e91487b3cce178a35a
z8efdf9635ad6093dc708a95f1dc2fa961633f678643f12469e4c64fc30cb765d1735e68c86e2d0
zf470a872e07a7f7a48cbab5809aa89569d6642206614ada21ec3e225e05afa0b531aeb62f348b3
z8033630fd1fac1ce9f2a64472d83018e2664b0a3f3a7546aaf83db12520c47f5c27f4fc7986769
zfb5fa4ad114d371d1d1f0d27f6c868b704c4a16b3250ee8b9e8102000aaa7b1f244a1785888e77
z4f12de1b905d8c38c9ba550b05ffb91d48e82baff426bae2e0a41faf33391aa2405723a7542df5
zf46a42a10c537a51e5eda8543933dc44f1ac1103e66b705ab32c721f7d267aebacfa3ef5ac2b11
z93e2b5235aa9f71d612bb803efe1c9e359324d8fe95e1d321e63ca9236b3876e59491cf520abfc
z4afc11925b64e10c0dc78faaff9be11080c3f7818ebc9659160069b366c81398f4ffadcb8635c5
z61c496e8752ed9cadc1e13d4f359c39f305edf4a1f0d0d312c2162ab4a08be28d8844a3d9e4d9f
z4b645872d52bea71c76f35c858045e1d41e41a53de4fc4cb7a59932cb3380e6bea7b336ea4dbe8
z52fb375dff9b125ce685ec63b2fa910d4b8d3c0906ae4205e0e3cf027c1291c9e353fd72e6d134
zb7180821d0b31e7dcd2b86666a04245ea3057e689e187ddb2351ebb063a92093524b4423d72760
ze316ca06c277c0b4f3d2b68ac322d6b38b9b90d11b28bda8d6b2b9838b17ef95b00087927bf58b
z03f43b2c3873984d2a29cc978a2f1c5e0dc646d760245d0d3aed54ddcd822b9db287fa32fc33f1
zdce66b93fae032a10f0618cb566bbba528f3e0bdbbb6ed117dbb12f8344538f9094ecf6e552cc8
z6e0ac7ff380e5bb17c9a1a51f25b4a615ce61ae1b224740ff4153080689b29a9c6648015e4f7a2
z4ef368d546393f89f9350a8fe32e86ee21e795cf7942fe54c532515c4eca95917e0a08f1145971
z088ecfdac31489d8a7cb67857f166f80d9e6282691239b9b5ca860863031f847a885a90c8a434f
z22a68156aa7d46e28544228a9dd610ecceeb14c57b4ac92c4d0b1a13d9802d1678e8ef08862add
z5353db02ce70b2c75257589952c98ddaeeb1421da3beac1be8595a4fa1dc89f34f8f4dd097556c
z4eeb76d385d1acc160df2f4eb5fbf4f109713fcd8541c9909d3b09e0f91c00a61aaab6f701579f
ze9636598df8c0496569f8c221b33ed212e0399febc1973963087f798cd2e85360a1318538ee5a4
z7240bb3478f33ec12613ef74d72c7f83c257e4d8d2f8c8e563b2da35efd72682edcf5cdd6c318f
zad1a4bd9f287ae7056d60101fa423d5ac825d5e3f49f80797cd45620b41753dd5d161e83a8694c
zbf3dfcfdc55649de3368bb6cd8756c89e7e47e278e15fcf1c696e82ca79fdc8d513e9adec4dc01
z6e643b31c947347ef1f7a5dde855b97e2fd1ffcbfc6d6a4739e597fd509c4d5828c69204a8fbbc
za399d96af9d72eff229bbb38e87f53a8c0377f779018dccecf716e3f42c6f4b72e60670b115a88
zd271bc4c534bf48ddca33a2c1e642ac2d87fba8ce44ff7eef6e2707224e140c381837b5e175a4c
z2692338b69bd334fed0fc295a5eb8e90f09d2b0b77c261d16093f40ccc029439c6a598203200ad
zc255705c944711c87216c69b8cbd5a2b7f90df2edab510d80a8755c543538e76f003f232201572
z33fac3eb6a89b44e9d960b36c3e3394558a9dfc8bb7ef41626be8c10baf4fddaf0d65d24876714
z4055b20688577f4f7f12e461735f794e1ba82beb10e64fcf1ffc9a74e24802d3294ffe54090d16
z66c6236a36e29b796f08b6632c999af5f29ff662a0a37d221b29edc85f13f5037d9b76ba176aa0
z890efa69a948b50a268c75497cdf845e82ebb1f404a62d186f76941ef4f4c506db94d6f8ea6cc6
zbde2d422f6ef471a7f90ea37675d4a46e501c5f74e30a21dc51f29622cc5c2d4b1699ab90d37a6
z2756344475d6c7618e7cc0555ad13bcec4516752ed6221552c062aa42ab7598f6869e1db414585
z0b156aee31690cc5454b1ca1904f95323d6d8f8db48eb27867fb1f31edf834b07a7b0ed8b59db2
z2c6ad17b10175b91f7c11b242a39541ae0784dc1c7bef4f2a1066b4522c2dff54a86ea3cc34f9f
z92e63f4425ae859187788d9bdabf87358afef512fb0eef9d48bacb5736d116c795d781fb1e10cd
z2c0fe44aa6ae8cc7ccb92cd834f44c75616d265dc226049bf8205d936e9c2719b6da28c06538cb
z8644b550b2894e40da6a9f9c4c99e8208b6aaf44464c95ccd327029c952e1265a53b079b62843b
z5948a74982b86a05e6f706e77b8f7350972f6fc01ebc8f038f8950e0fe2e276a4f663c9c101b28
zadfdb43edbae791c67183e0e1698c6c80987389f04fa13a9cade6670c7c1a0882df315790fd410
ze4b1c9c2098e2b2244a43618a25b20be71caed154734f6dd6320fc1da1f1128f7f566fcd396c52
zc3c9123cdbd25ff4afaf4db073c636d20d88544313f1fe8d59c3fe8ad67ed1f42e6246b0228f9a
zec8f2259082719fda8a7cfba103164a4731ad4bbbe1ecfa0d12dd03499e2ec36fc92df97022bbc
z3564ddea193beae1e7ce31fe634cb3fc7d91ae7bd37cd9261f90d92af446a0d6451a77b2aede92
z8af2cff2c80509592c155d9950d7be5d53b697364dec7cf6728d061eda96d7aa7299bbdc31d008
zeb215a3166cb8987f5be7f277e45c262d09d37c8b2aab851203a7327b69d296516b4f370292c2f
z2f3470f2eb0971cd8406c632d0b53a531f141668c29d3e533791e98a0122201cb89136a31eed2a
za89e29a40a8103a9c5cb0db30dcf4db9fce37079fea483bba55280b4b335f7e007c1d6351c5f0d
z08b63d6f5ee097fdcece8a07037d8c95d22846902e6362a6b7e4dd49746848649aa2b31db64df2
zbd60c29a2834dc21cfd55c1e6aab93cb28daabf833615fc275e5d1c1b3fec6969cfe3e3adf48b0
zabd731e97dca7c79160ed7f13eff691e86e31c44aa9af4e9e7e3dff0a23f1d7bd1ef3db6952347
z144497a92a21882e8eb6850882c7cf96e11147c2e124f7c9c799f8776c6316c636268c8f9028ab
zb0f3a191b7745e38c3794555b866399fcf6bf3c2d4c34f5d0597b51b3014c81c8f6e072798ede9
z766533a0f221ae4e30b94935b3365142647aedd246d872a48b8f524afcb29d4e5d3a1b74d47145
zcf6ab9cae0e3346cc275dc71ac050e200564f57e5eab263437960bc20ac089ed8bf3a691e97fc4
z4bea13b013b57b2264aa965a28e4718b5ee765ca9a10161c97d079fde06dfdf280f00227a9c33d
zc094b886746f5c8e6de37732018bf87723ae3bffc5f32217f3355a042142ebc2122e53da73833f
z1df35b38cd4c8121a02448359536518e12e1100e30a8a11a0b66a2cab0342113c938cd9216e446
z8e0f3b76984e13317b3389ba2e5f5bda542413d7bcbfb63c2a3ad400e397f58844c051134807c5
z1079c8e7b9bd62c424216f0dfdd9f29a854737b85785d1fa24fadf16ee682930c764e878af8ad5
zc726e4df4fe8926d9278a726ed423c80a38ea1d69c62431ded75fc6b596f475731419b64743091
z922aeb01642248bcd8705bfa1d97b5112ee1d95de1a466e76ece0dffd2ca99ded072258be500ac
z844eb6e3f08198f691f3969d4ac0394c776fc94cdde7a67eca89997a48374b46cb02cf2e34c3b0
z7b3f1d6834772af0398e19501d5f6728205b921333b66a7439bbd7e042ae3a4aed16cbde4407be
z057e92988716da3d51908e9c9141b02f0a6cf56697aabb5fa4fad90cd581da05d65777670dd4c3
z61ccc6e026d80ab3a483b1832f6ac5f676beb4ed5a9ba4f8e0d41c8cb02a48795c557e122cfc30
ze69754954648e23cd2e0e828f667eb082f23147c61fdaf5e8a8e325ba80fdaa87979b7be6b3399
z654320871ecc1b501cd8f1bbe44f5ed7f01d79a6f1d986afb27a8d4699ec38e06f24bb90148b65
z7b3a0b206b8c25abae25e42c2dec2aebbebc3da2c488c2e0517cbae4af42a12fe0f6efa6d369ab
z6edbe21bb3216d7fdbf018c8f811d8419986b60c923b88849cc8b5602d359edcd844b1b8d7ab42
z6cc10b0b3de1b63bad84b6387e14ec0e4e26f3a6d26fa6af22a2be066d4482997ea363387387a8
zbbd827a70f97b57520af4da6e05e3ff2fd06415a445759527c049cf44c8b36446e5e2e74b6e88b
z7f7920db7b492cd22d5815f66691b78a06729b80cdc2c5a9a05badcc735ddec7462b14ee3c53ef
za0195066c7c8f8ea8c60bc0eec3737187c60c492673cd648e696c98fa21b2eb49f4718aa022eea
za9541cbeb2948028f49529bfcfa3b0036cab275a7faf48fb671d26e1b0e6f8c984870c045082c7
z6d1e875fc108e10eaa78ce396dfeacf7a4134357fe692dfae371a7ac959e9a8439e165fffddbcb
zc607c119a0203763b6b65fc731448fb7df83a90e3c9a1d355602548c44f664890c72da4917540b
zdd9b61939e193a92c48090a51bb858558029edca66806693cbf166c7b6c061eab90247eedf01d5
z7eb835905e95743bcc0c6821aa147172148b173a3d1a1b4776c0bc7ab23b0a6809a1010016b0b2
zead701e37dfbe419782f814f1df5b5f6ea1d4e39d43c86737cef1ad3e9a040fb4b3a4c4e9872e5
z94ce482fec8b610ef1aee0fed559571ec4ac8fa2a6bf2d36542e9109bedecba2f9e7b254c5c101
z782ca3e46f4078f93462c057bd4cffb5cbf26968240d4b7f39f6a6161882f6a6fa7f99d9ff71a9
zd73ebe645a0fa01501268ecde2f064d73bbb3bae7f5fe16ac0a5dc8f7aa2a8116bb77b9ad1a0e6
z8c82a2ea748f87bd0c0d7ea43924323b173064f78486160b922b02b4f889f6d9c810648fedd582
z89edd1bf7679fcdaaf12792ddd4e939697652f4c09a0152e9e4a12d911b0e23977917fa54cd119
zee1ab772b9e0c0c0af767979771e80b696f40361adcabf9cee30d5305ab747c061c6b8eadfb561
z5bfbd46b16683e0d58a7d22d39999032297f85a231bae578d5259780f5ae9a5191fdd0f0037906
z9d66aeb210950173ee7c6deb997df4fcb8ed3c46962f43f585487baf761959ff2e63c0a7aa37c4
zf169c59b0540a81c277ad78bd8da288107143c4cc155c8c1178563f7544a2804b3cd31d098e584
zbbad4073c324ab9caf1855b73b1c2411181104b864af17cd85ac54ac153ff83c82e12ca55ce929
z3ecc603f8c837a8abf9160ba4dc40f9f14e413eb1b1908a9e7786ff915bd0959cb1be3133c8a4f
zfdf46db3c9cbec25fab37b12b86da0c0ad705211c7d84f013981e4c3f529724a8a85f35ca916d0
ze065b1853f75ecf62a9f7d20e4ca1a1ff18f4ebbd74a764df0f07c2d6b4e77d9e2974044c1389e
z77f6755a94e99b084d6ffce7ba0c2bcb77659adbdd82f70840a904760c3ac153a4f187a62091e2
z3eb307f0021b308e66c9f9e4592c725221d30053f876ee5cde7cbddaccc9a649d79c91dc5b78f9
zb5fb77a1562fdf350e75abf581b1b9ab58941bb8489d230246d41d59f6f5af7dec728be1d01489
z7163b96178298eb411b000b3bcf77500337d677ed637491677ff6738ad803318669cacb0210974
z866c5e22bd8e26a4aaf5ebf3cb38cc2b9ace7b52cc68e51b58b7fb0e5f401b71c1a3e305ea9bdd
zc12507f06cfa98c3c975712ca3942cec6c565aae37b348d5b73f068cd3303626f3aac336811e68
zb28ce53d3f08faad93335e1828d36f714fa5038f6a5c3bdbebd205e77a58ac76a5f6faefa18c80
zc1832efd6c7cf6b7aa1d84c442cf2731d789358f40dda887b125253a1dae9b6ef1d2a7917a730c
z359b55fa542c9b454299b5548b22148a139f25780e87aeb7053da67fb8160f7f042098998dc400
za5c1109f529ce6b3cf6146daf15b3ddf72ec8d3442e8490262f6d0b2b9501a2d8f81024974127a
z3be94103f3aa47901732432995a021a571fa33e5f95515f0c110796b3ce5398250ef1be17e6c83
zfe22b4ab6af23580c19ce58f6f9374f1aa3b46ddd7dbf1dfd898bf33ac25fa7ee98214da77801b
za5aa04b9a907ac6629d8ac9398d36fdd6fd10b98f146bd4a51a1a330a08d5f4eb54ab4030e63c6
z2ee547c9f3f0783d6264c7ad9965abd8133b40c7c92fa5645b64de1e9207a5f7dc8d64f92691e0
z2174435ffcb4967778dcf0accb5a70c1762f404e9e5e39534e82ea2fe382c97e94f9953313b7e2
z7216bbe99f276aa2a8c694a479a53e70072550e6c53ed0c79b5d6a71c4b18055437a4e52f09ecb
zd8c8f583983aec63ddb6243a821df6ae16d48fdf59160ee2f462e4bd9686422932e235cab409e3
z13ca373a186db0436e01fb18c352a37c9026f3231757c7c2683d61791d7b26e866de268400a0a0
z1c152bb66d8034c00084c063bb6bf6f76ef8864119ca296a49a7c99d3fe717cd8ed6ef1043bf1e
zc87b4fabaed148492a8f12087595e0e218f8379fec72453c66483f0db17df16ef0dbe73a9d57f6
z71a429f8a7540d1f4d58614f4dc6658602d27b28a958f5cd7c52f0d76aa0d74d7b932f7ba14896
z454ef7722995fb5b6cbd6b43dcecbb0f98c96d7db467cd04eff1cab39763e0a562f1add73ef5c5
za73b69d9ee5bca6948c160b49922ef95413519f8e1064a0fe284258f6e28d72bfaef7535565535
z9e73541ea44c4d9b2dd26e00e6c9811407c19c5f93575aa7adaaf97db513480d524d656ea625bd
z120156207fb8a337efc20d83d995df5038baf22504fb76cb7f1e790eaaab42addbe54ffc4e7fce
zb4e3edabd728fbc806721e14800db25a890174abbb8d9157279ee26a5272fdedeac2649e107b0b
z6936e100c3b961cc0e8880989486737bbb46d85e28929351c0d78bbfe934ce37f9ab1627460a4b
z6b96a6626aefc4eda57d1e3247b3607b8c376bd8f2ce86c529d6b8bb96cc75c46a6442c9fa3672
z1c21850177ba0d3446df141dadafa43a0785b8588bcc06ee8bfb26fc8d9be9e8f366e2daedb1dd
zb3930ed8cdafd8f51a12362412d0a1f47abbaf6d53b85c797b0ae26d7663464dec8764112bbc7c
ze4853b2663ab7ace6a5d40677a9409829b2f58c4a3f69b5010dbfcf3f16ac2785a123f8b3facc8
z1c58b98a5de49b78ac046c950560699a952ed1c2ce9c3ae87bf0ad1db9fef4c02418e81c99b531
z96be92d14db2f4eee4365f3433c4b98b4f9ba0f1eeeb881a01c5a484b91571be1766d2afb51755
zec70d145e67b3f484f58f524f81e332526b6045e02f6d09fbc0dc31352c6746c74e4f9f57b4dfe
za0fe3cd477a3c0a03edebb073c84a97edc8254dcb600e868da3e9442bb122bce2b4eb96a05d3f7
z913479d5faa7280f09ee185b21b3a0831453c03a7f40a94d0477954c2bc9a9ca8eb000dbae376c
z95c9d7f75de927ecdf1802ecd59a1a15a0a3382d3f664dbc14d4e45ef36113fb35537105a3dc74
zc65893fcab6be654344200a2cafe99d638acbf037c531e50aaf3d075d72200145d650f6d2b9e32
z3731d6770f849e3bf1aa3c77fd633d73d4a28896c1f2bbe4426adec236fa0a0744b053f8611804
z3d5e407fca3acce113203c2791d309f629f2bd3d5cea7230feb9e2a61390e6aaab4ba1cdc77272
zf4389c18a7be9212013ae10acc4630885028edb9ebd2c7bc2fc6de9b7d37d55b13417fda2ad373
z32180932eddb6d5a66863288e146c106a42c64a754f45c582aeaa797716288a36f0941e8d1a3c1
z40d7af557f7ded738a98805603aa1e6e3a9cd7b28ccac294e4c3607aa15fbb5a8b36516a54f68c
z1573cb4df0118f37fd034a10e05990c3d9b39f388204bd381ffcca41b0f954b1868bcaa5dd9035
zad8d9d0b513ac6a2534feab64da6f870ce598448aa1df65950c05286965ea4e946ad072f2153cd
z253345c8993746806f90b7b90f6170501e9b8ff4021ead136e1f3e22f11be5c3757371b1d3326b
za20af22992def031402b9e8cce2d02e289d1f5335e80ba9bdb8af1854164369d7121324da4120a
z72c4a411d59f152029fc0c254c65b5e60ea1e3f83a47cc100a381e7e15e864294daa8c128e12f1
z9d6eaece89b905e1fdb2084d25e237fe5db2610f9666b2f87728a3077f3118179cfb1bfe3ca574
z0c5e9a3ee5cda409949382ad836b515c6f6af094dc12ccc5c77598570193401aab1ba4cdcdf322
zaec51b50d57a0238afced24c92636057a6b59bc5c17744106658517a9cc44f2bd3a225ce6d841a
z574cfc25aefb61a59256440f8ae258f5b12225790784e3b5dbabf7a0d19fb6fd6eb92f899b9485
zca097199f6f1cd61fc5a4ae9f768ff7cfbb317f9c612fe6fee2e771d0cfe5c89e5fa5136da7abf
zf9772ec03667041677a9a72e36b5569efaa0a12713d9bda78e874fa9ab5f4f8a9feac983d52f59
z6589d64c8473bdbea8570cbcd958e58fc472341cb6bf19dc23fa22cf3153cb766c09f55703e825
z2a66800baddcdec80aaaa1caf70d4c0ba1521d8d1d76745a3547f47207014cf4dc4d1078bdc7f5
z2b67dbc4c0fd1811ec9006d1e578e76477dcab07123fbb637c5d60b864e04ca9cb356b4c2b8537
z3261683464fcf68ea2801bc511a35e9f54e224b84972116852a8fa4332b6d6bfb4a17b1efadd48
z14741d803a7fa03987b303a89ff2229719b0e7bfa9ff33368362da187b39933a140cdc42bd8a9e
za2cccc1c620fc1b29c13427c17a6885935be31e4a0ffe140628a0d0542d0bf2be2f1d4b3051c72
z3b8f6d61d69378e8fe6f8005f0b0c5a0303123cd97d75f59109a9e61c8d3a94188ebdd90d2b63a
z9087b1b81956703602327fda7c8aa01889f1d32cacaf9e0370a43353efb80e8cddfa49e4eac798
z0a4d84af14d748551559389ed7291fc6f16997fd7ec47448426969b2fcbc4e88da35993ec30cb8
z8efc4ca7d9edba05f9fcfd24898679120267c4da38d616368c52c94f09f96448c9c0cf9f8d2777
z015154578f91e8729653174d1de5afa9010645009c19d2e5dea020464e6b264cb1e5857da9a26d
ze94f524b5e87e4f5adaaaf6e6bce71a2fda38abe754ce4b45dcb211668bc772d2a0ecb178ae943
z8137dce61e8e0f5d6a3ef66502b89aac5bf005ad572e4818031a31a44165dd244c21f7a980c8ec
zfb3ced810280e78f846475257f96129feae4e7f8ea260a0e96963f4ed0980a316ec770d74fc51f
z1243c15f1d37e91f6529e62ced5e252f636f094b34c30d72c5d1582da8c59390bcd6fe5ce15831
z0f7d384e361300032fb6101dea22713afaab5d3cbee9f1581410291b2cdbb38a608aae6713d9ec
z52b45a6a274340eb0959f7067433f989aee9c5bf04f8426924c694e544923012f8a6bd456717c9
z656f670c290282369fd9daca5e3ee12b6a1f7ab8de078d46655bef07f744c9afe8dcd999ec15fe
z749edd258d5160b14de4bfdaac692f5b902f5be45e411c265fadc104864705df6724351a9fc706
z645c03b15cfa4f7dc17ef2bbe6a89c4daf73c6ff0e6153d76c39e0689bac2b58fd98294e5272fa
z2a695375e79b2d90ad6054e4229370da19b39a4101197fc5fada11883fdef3381c59cfd27e0438
zc875ed72a757d1b7342e37c27d54cd82656ec9234981004db06cba5b1f1636d31c47dbe78aa2cf
z5e01e31cf75f17f48b37ad6048081b9fa0fc181e75174053463807fb224669fd93407c86916252
z602b133b34700a46f2f1b8605548742f77aad1d4af1268fdfb4358adf923e91e8722ec7f6feb04
z3fc5337e3a4246163a2e187af3ab8506e1c0bdefc69696b1d5d73a5fe65062e62d0cc39426dcbb
zc2d57daae997072ba478a4641cc2f8cb6ea71cc8bae2ce4a444192510d5f8b8fa4831cd48868d2
z303bc49c0ec473aba734ba1e016a3c3a326c61d535225db20bc911d203c5772ddd5957d47979fc
zd1ae5c75d7f6c9928c003058a94c8f506be3da05c3a79c592fb8e60b7ab7c32405d0de4bb5c99a
zb6bf02f0f53471051b931c22c49d6893db25d9d3ecb5e0a80ec11d5f46e9b37326c90d9fc59d65
z5bdbee50c9e80aa9b6ae01eb8e503f6f065c494ebfd5dc1f8e90d6ebbf755fac59af30b9a1b28a
zc77402cc4267874b90f817088a086882d6807c5d68b8dde8b92d38fab391c31efa21527c7a32f4
zdb2ac0cfce65d116d17e6ead2cd0ebcedb62344a9569ab925129d2f949818c1efe73c7a313483a
z35826a89654eb2ac9892d56267e3f5116afe2151173d7d0e21f73d57788240f32cd0737689c58b
z439e1f9cc3e433fb672d36cee74fda4e6c2b755de1c96c0521f03a5c7930633c60aa7a098f3369
zc9d6962289b2a9c00481a596d7b369b69ce479c26adac111251eaa19c91aa72b86d007439866b8
ze6c760826893943bf8879647eafc2e600769d4b24e9108384f995416589d936c3b3cc5930aa6ac
z43ae5232fd9f0dc17c1739f1c4b99cb4c28b19e609281314e2f2535e0c091ecbfd86a246fa37a1
z67829b8b9a80d915ba678a4230e452c957d156eeb694f15e2c790a04bc14250244e1d492dd736f
z12de1d7c65a04508981ca2cbc4bc3a570f71005f5c0e3215989280b7523c142bf70fe72ed97d8d
z82fb5dd32b208a4bb25c8a152e07d9188b42652d1adb5c79f0d6b58d7ef94e99b66be23c734f00
z6a2f9679ec6bc8a1d9b9cf0d35c4dac3b1d51c0aee096910823ea23d1aa5fbcf60b6a5c09a8a8c
z77d9112e65be6adc69fc14f508eb9d5bd7f097de762dfa89ba159161dc91fb6796330d6ee065a9
ze214b46d30ceff3659221ef7bf14e9624d5a572657d069bcf7ec170646b2d8bb303e49eaf5f123
zf70a575c9d5f1bdffdc126317b1de7e05fa9edc84450c48f6fcd0b5c8aed5cfec6c354515caa4d
z95d61d144997a9e64d9ca75b20da89dbf1769afbc1d2672dd6647a6949b5cc2124345ede5b7616
z2f5eaebd09eb1ac384e7ccabc424251b5e2c6acb04072ae9131d0f231caf61bef3b7dbae56eede
z396c01b21623d32e1c090da7a1f8cda7d1e3c38d94e20220d26065ea2178de6ee8e628e09078ba
z24f7624cb58d1cda712d32918778633d72d54962d40430e27b59ba7257368eee6e4ca1ec9de4d9
ze68a3b4739ac878b2ccfb448e6c6a2c43b733be494cd0d76c2696b18294d55eedb2b9ed9e1cb03
z552994af916107bb514141cdfb177230a2334f8fc650ff94cd38ca638658137db22e59bc2172e9
z4d0630575a3ffd331cc3781c1ad5528239aa3065fdb69e80883bed180ea3c1d84d70161bcc571c
zc0aadde155dba2a5edae6c61e1a76d55fccfbc371b52d0c8f65d02d1ab2e059787f3dc5dee5b09
z9a028a53e575ff633a7fb3b6f668642104f2868a3f8ba6dfd619ac3d2ab8de96907d5b56d023ad
zefbce2836808d2e06673eb5d5c2ba16dc1493d12976743c6016a3c81fac169937df63f65ac6296
z90e887076ab76fe160c1519e0e5f7b05fe90034da56f190d80ede0f9c6ddd4827abac806b25c2e
z1435b6564ae31795416ac4d220158082fcae6456be0abf7b7c22bcc8aa33f0c647641f6143d731
zed856531f9466d7b9d01eb4eff6317ae95520772a311cdf9c91cbb43a89e8d3544e106f4cdfdcf
zf2c1537941b16946d04666bbc08781b8d3da3820e9d54bf50afaadf4c9954887de7deea7a71c25
z2832771815642eceee222ec59610ee2d0b55aa44396f4737bb58d9e60c34f654dff0cfddd74dfe
z00f0d7492d1ab3bf1c9a0e2dd955a37fa56ac383c61189096f4435d4e3617ed6556211db8280fb
zc41dc71b4b79b916ac7006b85be2fcf3279c39c14631fe056d7107885879efdb01b09ea8cc7b1a
z8fd596a796e61e64534eaa7c247a36e8fee0538988c41cd69ddbc4c8fc18457d897dfcc2299386
zaee5e945fb09beaa9cd10fad54b1e16fd9fd01f0ad2cf9e25476e5c764fd85006dd3535f01300d
z12622a58c5607ab860cfb4c6ef2a3b8ce26cc96e845e9bf3f4c205fce6a9357622dd6d4ef3a268
zacd855a55c3a1953cd5f0e41bb5e34be79c0b484f06660dde5db173d48a3818893c5ed701f6e3b
z24068578e5d7d9fdfe1c570ee6d3e44565acad2a700ffe1887c7f4031352687b5356f9ad6afaaf
za5bca03d2258d3f7fb97b6036007304d609fd2d4b66c30d1f6a2eb6e013084d4026bf4d1a3e9bf
z054042d6bff72c67c48257723d22404f4a9fb814ae69bc8c88207ce4ea1ad1a890f1565c98f10d
zcf357e84e4e1a12f6c79946e1b5e71ac75982292fded92d70186d270aae0524a636830c59f1590
zeedc245808d27fba4eac3eec56561e0132408711ea0bb269d92c42a43b2fcad72dc1d7f164daf8
z2fc44afbebc464da402364b1fc3514d263b6ba9c1e70a12ccf802d0cdf56690416c0aa8815b76e
z1ed9ee21af61fbb27f680f7faa7b5173cea4e2e9307d6c3b29d581634afaa51cdd4e12f24afe9e
z73b13036ad8437e4f5c702701b9c2eaebd39fa284529b79fcf99d8726115a6554718152ff9d89e
z4bd99f50bef4fbb3df15530e28740d58caa66ff5532e7fa2988ac8cf9a8b5c8786f453c7e1e381
z925ca26370e641c0c22141d1cdbd222235ef501485aa8274dd2ca0ac2c3db592fac69d7ee26612
zb286d54537db6c8a234006d9a8402efab96e4059fe22f7ae19762034eafa448c3fdd9b12fc3f18
z81b0658a45cde402a045b18d325070077357d4192705bd9ba1510be9201018b3ab33c764376ba6
z5a04c2beee9de156429edc5e8693fc0592203b82fb0931263cd1655fa9383274b9762b0d99ea45
z876c2360336a090f25d8d72a437296f6d27ae729ed84539c685d19f98f128e4c3c89ad2f7228b5
zd586e155e2263f9a8f1e9086592030271fa72b2acadab0ff7df1f4873011234905944e49c3bbcb
z4c47bfd8411b510cc52a537058da717d1cc9c0dfc4c74b714d3113716140a508efd871f964342f
z75a8f9bb05929cf99c1aa6d68118d17d757464ae48a09aa14396c990ddf5d6f7df4a4d6d926ba4
z289c0b90a943996c98053261df9db74faf7a4d37da372f18faa2491169e9154ca2e3cc7dffd161
z5af962ceb78730dc229b8786ce5d3fdc9400e99b0c001c24139db031d27c675327205f8df56232
zc4fe1d36a5006f3826df323536d664416d546ec7bd0ae614b78892296b2117ffc61b3851a11a56
z812abae32f05892eab33652bc9c3bfff80736b870033ceedacff827cf23052c2467a5b728e2aa7
z9134ba87c948f2d2c76fd25f0963a92cff6904ff728b7c658dfb305c5abddb92e60aef7eaeeca5
zdfd1c02213869cdeeb006639ffd645a7b5648afec027d86ffa3eb6576d8d7c6dc6e29cf69312b7
z419e24b6b715391c97d2b37d81ea7d697a1ce04a1cbd70be0e38b52f81ccd25c4911db497f15e9
z78cf4d9887a8711c3fd7ed02d788f6c4e79baf01cbb189f7453118874aac11dcec15892c5169e3
z8577b570d8ace731ea8013e257f3575326cb02885a31c95825b8787e88fc51e61339b87fab6007
z6b03a3671ce1eadaae8c39de89fc15a810508de9419eef19aacd927830c34fb1fc8601ffb92094
z89c3e65fe2e63cce98c8cd91460cadcb2bd362b9182c128a09eabe8f08180fb7367bcf0867724e
ze139199c637ed40443bd2b0a7057eeeaf3a8d6ed3166f7e386bc43590d1eb5d24ccd19361483f9
zb995d8d13c4471c41ed52ed5876c0473f8f32dd1b3d5a60b316015546c2daed0f852d31e0ea18d
zcc9c4b65bd563530a448072d8a68218bec2baa249120f3c1c8d40251992669c1959c831dd903b0
zed94f8e56ad475f84b9c99ec9db39d6e5281ccf61d2cd3989e17600bf03567a70c9d185f63774a
z1c3d2ad60488ffac3a03efe0d4a8f4a099b4453d8914ef8f54423288c86baeeda4c9ed3842ae2e
z9ce1eccfbf8bfba0d5f6f5e338989dc6a783ed5f9731f58c7d91ea8c1573a07735845b86421591
zf495cb923d1dde01a462a72caf0e5cbc1a6a8a0f7e0417b16258b6a290bfc5bceaf44d7f706d7a
z4c3465f452e97549ed11abdebe6b36bd3b99df299c1d73cf042b53f0cef65bd4cfe15d6a03500f
za3d7f039020de8a5d5203d534940226296d64250b52ba0321c49468e8d493bbf605822a4e9596d
z858a2be2e8cee2d792beffdf24a97620d402bad4ad25a1d47d9a124aa5db57f98ac46c3ffb1ab1
z982aeec50b9c648c295c7176a7fc483d45cdcbc4504d67c8f2c9c32327026001f88ad6e4a1a968
zaf536ba74ad55fde5cc5269f394b7da6b8595a8852034e7451c6cbba997684b15ef2ac84c4170f
zdb763f266c6b78e23d824018cec2f64916212989e5363cb8b12eec9b077a22c436403545f77cbc
z46152e7c9927eb4d44fe51fd48eae45441e5417c4fa2273dc1db23332971cc4ddfe4a3a05b21b0
zfa51d7ebe3354cb4b8a44ae577f2f0486d1cf22864d9ef541521dc4c37e61c507500425f23d607
z5a25b70000689069fd24b6fbd859af96411728f3fa41a4facd5e5e66a347737dca646c8f6de3b1
zf79e993b2ce447c5e525b81ed796e08ab5a3f250c93ccb6f8630c80fa4eb420a638734ab0bd440
z2bbff0452ce78b9f5462553a59418ed7e68a4ee34979345e66c9239fe49881f167bff33a442450
z6180872f9a662b96330d927b407d17e49e2dbf4275c6f6610cc51228a8544172b35fa9e13192e3
z0da93be795c2b84e271f0ea027e265b0aaa942a1bc8661079acb0ef52ea1268a997b6370d6af72
z7cc851a5cdaa9f212e669ec9af736cf25588176a402bfb8894be5bf01528f9fdafee23d3ef5aff
z2a5358d2a2c8d60775e05b10354b13c02fb99155f7022135b9b0a54252fb9c6fcb10f120fe936f
z90b93281e5676ab78764fad6487768e176f62c6586588f19d6ef817adfcafb2e1804d43e94159b
zfed59d2d87d2f72231ce30fd2f16a31d6f909d136676a0f34f5d67152653371816eee0f7bcea58
ze59c5991603e5028a661a5ef69183b68164e35253c6c53713d2740c0a09e6656360a37cec5ad81
z0404b922b99813854a756f9b122fe5a83aeb643198cde96ad86a34b6019c56c67ede442d2de8b0
z539515b31043e1cbd094ed5975bbb00125b22a912764d575d8aacf894cac5edeadae9a5859c4b4
z79edd9bf9b705083cccf2956009ae36fdfdb82cb161dc0088dfb88a38ea561b716cc7a37658f43
z304feb17335a1bb50a57e5247b7bb7f21edb09b8c33d6bd0ba83ee7f233e260e29b10a448f4dfa
za2ff2e8a1085469bf691118acbb3a97afdaf768d2eeac6f233e094668af2e912baaf888e2b9f09
zffddf983ccb66516201b393aa58f1b551f75fa30025bc57cfbeb013c2b90f54bfc9b46a548f1b8
zbe9d7549f25846823246c77385af72d4d04f796ff4f45ecfc2f0f1b13414b941aef07ba92da2cf
zecc9467fc72c9e6bfb0fb9557817998e66c53ab3060462a165650d26d5b6a72b111ebda611a377
zf4e1ae831f7a951ee30e19c40a82e48811721500b8b77b3dd7a9bff635cf4c202b955b78f2c2d0
zca6cc7a57f424c127263d51ac187a24d835aa5f52f39a3ea06bab5583631673102c50a612f992f
ze70f332929e4fe7a6e6600e3d849ce3fe615d34e3b7809ba7cea459a7adc76ae60cc2f30c8115b
z7a327ffa7912f24438923a940568f3c452fbdf01327c65ce0626fa8032dff1d3c71b3f798c62af
z217e3b5d97fa9b7145071a2fc28e553c273dde0d78111b1ee799854e22288f484019313d61a240
z7432b380d150b29a0a54a269ef509942b2098e4a809ee20de939d74fcac2ba460e8aa6ca171e69
zd5453fdca09d92d65d89745994b4643dcae92ae5d39c2343563a71e3421bfe46a5c051aaf8e321
z00e74208a30bd9c809e7ba7ce3163592c8474b49eeba671830a7cce87b877803b74f4c7c175323
z4f9c7eba98258e557890f7621b245dfef994512b74adb4a0ddf80c68fd8f229b75468d1c31b53f
zcb057867fbefa6487ab926fe20482e0b55aad5b50a8a2289451ab2b32751e476e7676dd70f1647
zebb300774b8c3d9b6369f9824e5010897c1fa4c641a0e55aa15abace985f735f96c832c94061a6
zc1e9d304f0de47f79470559ba5339b3dd1cbeeb2f4c440205624778857fb5f37a9cbf2814cf30c
z14e2ab5d2565e2ec08598b7cef36b9491aeaecb0988eaab87f84e734b1706153d073b7976cd585
zd67872431d8c1714016a6bfbb8ec44fdcf6bba1020e7f650c4e469e1c3b852a875c1f0254e5913
z46f2876e27be9050c50d1041979698202f3945b6ad8093a07e387317e7b0640c5ea7445be2808a
zc62d312c55d0d8d579f9395aabec1b53dbe36e2dd1fbbcd45964d798ec476b8ba6365e004fa912
z9149820051a98e179fda0d64dd70ee34e53ef73006a393433a4d58421bc5537d54dc167aa560a9
z3798452ee9c4eb14c74dbaaa17d6b7bb02c0a87a5b6a1fa6725e11a59ba20370433179c16669ba
z6df88ab3ae612681e32044c5b6c408c87eaa608751eaa68417d7e82f3e88563d3869f8d5c5e334
z48eeb8a76bd85e429b5dacf93dabae31db5be2270f639743a6a6acc1b5d47dba60eaf8a853ae53
z8c8ca611dd52e199a9c1d9586205844bd4fca0a70cb23f9dc7dedcd183b03a406c8e2958389a7d
z01cfc63c342dd9734766c4d745ae710d8e09f850cb70d297c4aebd3155b04b8fbf6ead0b42a851
zb8ca4a2902a14bc93416e19fd36aec228f356e77db63cf9876072198676fc78c163a8b0ffd558f
z419734d0dacd1457b31779bed7812d37abc0741391d3ab3fa38f0e3d37aaf3fb53d6aa524b60a6
zab018a85a57ebc2baa239a885189ff8faffd71fe4e2f428048e92c7525cdb4e98cc2df28813cd8
ze35c0cec99a41b079f2b7d491cf3b25f267d4bed06fe446632e646cd29178893919a83d823a10d
z3105a70b9e439de82f1c626826470de1db381042b1dbf392c22ff924097f5cb001d9b53b732f8b
za7f7d811c89e506515dd60e4973f788fa2f4ee12eb44ccf0724ac76aaaea2dd8063a834bc8456e
zd41c8c45595bbf6a251aad91eeb696f93fc677f13329a59fbe1e300f5e16eb7a9433a65aad5033
z36b4246d2e0f0db7fa0278e16da784e39be009319cfe245147d10c4aa0177c4d3435887140bb3b
z873f39acff36d4975458dfb70736eb614860d90a3cff8c402bea3957180359031cb0eb474d2d23
za1534bdcfaee3b46bc51997da5ea3f77c2c7e5f9c48512b8e9cc092bbdc925eae66ef378a8c557
z20bb85750296ffa6a53b53754265b111c1d6d1d000540955241b747909f1d71059988aaf1bd588
z40abc13b0e3afe2d832198c4b0fe716bed6fcd26af5a4be4022b7704972471172812e6ccb9ecfe
z7f5e257ba641f6d1a14e54254c2f3b7fbd5109aa26a1f54b0cba4a5dd2062c57dff72821c982aa
z4f826a4190b75e27b97465138c2979fd53dc2266fc644dc11d03ee96cbbfa042ff9e01ed6aebb5
z20b8b634627b0f4087f3e3baf67669f871fbbcadd80702c167ebf060aa409acf1ecc462abbb49c
z2daf7816abaff7747b9b73e4e9e5fbe0300cd84a31d1a46fbd588dc90da35964c657d2ba92b923
z0f8a8686b53f85899b8be322134ed6d8ab58739bbb4c18a2a5eaced8720249517b0825edf74d4e
zb5249b1e4b6aaa6bc3af5cd878176d8332cf0d3b93b363b0b05c690276a185d2bfc673bb6a6c14
ze6ee4893f96c081b7d4c91b7899749adb3cf3d29fd437b0bbf5877cc4bfe659dd71c3099f700e6
z9f4206c86a92edd0bf38030378164f2e1683e847d1b938afbaeb0fc0508cefb52935edce73c79d
z108534a75723089e4ac82d9ec8e01ed0d0c21c115bfbda454040fce6806ca523f523fa0aeaf720
zde5e885475a227b03de09e8c58821cf021701b504dd9e9645dfd0b0a218b02a73a59fa974941d2
zc8ec1dc3761c5497539732d5a3ea00f8fe81968c5fb5d3b7aed2d7c039c19ce653113dbb028cd4
z0d3c51d42596cb5eba6d3c6a15834c181cb2ed9f4ba4e9023cd66e1ac8604f38db31d174494296
zb4905dd947f2253a60adc7fafa95157020a82023793699806e1f08a18fa64cc293642c7d999d9e
z75a4fc5714ba6e8ee2c91825f04707944105bef88ac609cb7dbf6078a2c91b708d3cfd4d0b96d5
z6ba2d25d2cfda1c781de9594af875fbc708935589109a825992b07b6d648163e30e1b756fa0f56
z6cf1589179d00359102a978041fe1042a52b4a1bfe48439ee3f9ab5decfe7caff1ccde0cdb7381
ze9429471b88f4460eee46799ccb69f6c5842b7ba28b76bab3a9e2a9e114fb724b538914880e374
zdd3165de188672438adccdf68bf4f47f46ed69eb905caec64fec8c113e4b572c46668f0134c01b
zc5036dd70c9e82535ee25a7dc5b5eed3c96d6096179c66643d57d0cd600d2445e8d5ce04515ac7
zf975da3c0aba5966e610ad391fc3a640f3bf3077c9a3a149ba241ede225cde1780b809b40bf388
z509902a49e8374e1e2dc134deeaf97d2aa685300514beda47f17fd8b3bf22c03f1d52e420a457f
z9dadebd536505a326cbcbf5d552cfb64442f33d27b8605181113f69b138bdf51ecf1d8a82943db
zedf759b9c94cd6e30d275af59da377925fe005feb8253530f6abbe3ef45ee468dc2eba00bfba6c
z554dcd1edefae78ec65b9ccd0233fd3a5e8700916319e88eb8c5994324ee0e2876c723acc344ff
z4711005f6e1ea8d4a236e8402f960f78c4eb37bca00e0bde19d1403169f91f4a21932568b4656a
z5bf2d3b94a0ee0777eae26e9be065117d3303300f75f8a419a45c53eee2e505bf78f92afcc0940
z8bd98869eb54fd6831a2a92f19556b84ab2d12c237895b5a65c5846af1b14fb181f2d30e0361a9
z4f373ad0d1968ebff1c8c17160e7697944ab6995dc849a99b693821ce969e24ecc365ad7b6a2f3
z50f61b66e048d2f8daee0d4ee0773f341e7c8cb6060ecb8efc3ce0447062bed9a9879e8f3c0c61
z2f0b7968ac2e541c65a50cb32912a6fbf96cfe26f2a912f8fda74056f018952b65c5e1aa887f20
z008c89005b6ff5df05366aa985aba8940df4e47924c800d330a78175d9f14b49a17458cc331988
z2b8e1f5f582a6919c73aee3651e70e6aef75aba74bcc8d8ae9b0f895b7589d15e89fe1c4561705
zd39c0b84bc08ee8b36d2ccb49e7dd9a2286c039103fbf57023225d8eb177b8bf2cf4bce83c7846
z1e9e25394f4d46929341f0b2c76bc51faefb99cab6f49a6dc763326a21e5e766933075611b8179
z2ef2b8b86027f72e16977bbc3273c92335234a5126be1265189f5b1470f0c252c834814eaff1a7
z09c1613ed8558d272b7f762e7afe31b4b61f485dc8e0edbda72ecb86c5cf7150503907a2db1ae6
zb3104c9e02010cfd477829d7bc2cbd282e610a849c6abccce2522c26a447d1b013aa616a3f09ab
zca6fc5af44e66526d2c891d34580ab47e1d82c3faf3644876d10ddaaa99a6577c3575dfbb8fe35
ze23ded462db536c3de4f72a748df6310ddd24561bdacdda2b1c097ef2df4b665390a593ceed66a
zf9faf903bd299f7706f0e799ef536d4e3ee447978ac768354ceb0776a214ee77a198aba2429a03
z25cf8739af39cfa2ed882b09dbb3062b877505eea7eccfee6a5512498a7435a92519986575517a
z9ac763a0a13af178f5032bb5ff36c3daf2c85c5c8147296c38ab1149c900a71a10e1936a4487ee
zcf4e465d9aaa62c7279d4d5625200222b0fb62efda48fb33d45a08185625b8a564ebd55af2fbb4
z04ad8cc7de4214da327747aedb9a7cede03098ffdc96bfa969bb7ae6620ba8b227a047571c9f77
ze07bbff3e81b73c4ea85c26ed183afdfc077e4fabf3a6b74872b0d0b6410b2d858c91026b962b2
z4504447bfa636d4120e290a9569ad45596443499affa21446b74f92963a28d2d10e11df7d50744
ze17f49a7e5d9ee6df4aff9b16a774afe4070272649c648414a3a3f7aadb35378837e0597236a52
z04d0b1a0a28e6f47e3003343e3b7886fd90c5f0c9bbe93f3a24d1172152c77c9bcf485a40bd5e9
z7e444d7952008717564b26fc3bd19def65f9c85e83d3ad0c361835099f7e9aaa3db11d502846fb
z2ab693f386a7ac0d0e9c94e43f3d3aedfa8f24a5fd689ef81de2e1bd2274e213f56c02fcc6511d
z02748d18950e28886cb2e4fed7425305ba6db84bc85c3e1e8be0676f1433ddd9591c52e7e05eb5
z350149ebccec7e375e7eba2088c00e21825069ff2d59625208f0e6951529feb36ef2423661a30e
z688360ac613d4221a36ff30bc4fdf29c5958fbc00e83fc06eadfd1196adc8b8c355440055cd3d4
z92910af0c1516dbf10b071a979c6cbb05503c684403c7dc7a30688638eb58250fd9c6645c3a15c
z80444771ea2f2977da38c74e3a5374ec071aeaed20fe8f498e158a681762b2021bd1c295fc36b1
z3272213ff699a3a08cd26ba9f33cdac3b46e1abec288f7620dc8028286f18c2be01ad82f24c9e3
z1e0fdbfc9bd7dbe055ca0516a16f2658c3f3116c3e74f32c736e1ca341d55af840c51506c4f2f0
zf441fa8fc8c269d02752781d2db5a4ecce7e5aab2e084289d57c8f1f61af6f4e0902c84b589aa9
za645b719e11b4005d4f636e466a1b2bc4ff7415eca5debc7804f0190cc4c69bbeba3f15a7ffda7
z1f418496fa2d7e498a8657fa0b3747681a39ebefd5e43c8ce52838295e7260d43625e2c0cca9df
z166dbe8b71a71b7994e356903cdb0fa6852473f14e368e9184e53ac486ce1c2d7d7241cf673d00
zf5049ebebb73a5aaa2a8ef267048c675fc631eec96ed06b451171a89c6a67f9e7c5b9aa9b4a20c
zff695609535cf2c5854347d77127a96ea98ff3c750b7308e1841d54e17f2758f847a1488902d47
za31adbdf502b7c2915eaa37c0ff68add24b55ebae15d1b377bfec25f31553c7baad6d19b1a6b98
z2d2bcf1d8138e61f663dd640b449be594932c3ef085de93afdc28929a79be61871fc13c4ac251e
z191fe469ad5e5b79ec1071bb08a4e78470dc3a95c5884496b24ce852f41e92bbe72cf41be2b6b1
zc1a5c9094603a744783fcc337937262368c94192da9809c0b4ed8e2c59dc703885ba4b034fef7b
zf08c3389adb1f948853e89704dc01e9bdf92b5784778ab7059272c5661358f288642131f9207c3
z103b45cb7bb6e2a25a024be6c2b3dbf36bb8e1921f589a2f4e3516254af7a61319c94fb2977e93
z2fb0da91c053c41e6af800ba5fcedbfe1c69e0c9da4490619f3717dddd846448adc3902b86973c
zae9929a817a71bc8a1516fdc46f0a4901bd81d2c22c1d4e7072c197cd49d99c202c41d10a04425
zbe98c02eb9e896cae55907a2e9dd1bb8e74d7f6ba68ee4416154c887ece8211c331b88081e24c3
z49d7711a4fa1cc7b61e335f4a813784c86d5227a37f042e9ada26c0ccb2a70178447841592d6ab
z3b6e771bca4cec074844700ed14132818c443f4ed0d17b75bc52656df21097ffb101deefac946a
z519172279f3c6b0eb315d348ce7412ff61f6586675d01c7abac4fa7aa9286cc2cf45fa0ebf826d
z60d741ffc851c9b002c02fbdc0fa928d6a49dc0a749cedc9940e6320fbce6e9e01e1350b5d1afd
zf275b32bd2675736d1ea9193a838f90f7441a7173adf099e0e72ceb263b29c14f690fd24d32083
zf71c44822cc07792b43a198eccfae56ac3b88daa9ee999bd2df240f4a353279b8c0a3ff02d52c4
z603cfb6162ee7d7c48e24f684fb836ffc779516c0a43c452183367e0657d6431c38b20d64c2fb3
ze00bcd6244d7f6171419f1edebed51416de88a50d93f937b5400c8c61b79b0e16448cd1ae71df7
z87d2c1d6ed664eb7688c57b2ee581acee520e8e439fcaae426eab77418fbbe571ad325bb1b05ed
z7f6d1479499880b4770b326a965d1d126085cbb0bc416a87edc84fa4706fc2c3153907ac84364b
zcc461ebbd272d6f91f5a16260260e284ff6d5b668dc52c43de4130b6d678f4b743a90be56c8ba5
za54d8b6e634f387c564107acd0319ec3508d6851810601fd3be11b79bd6f05e9dbe8e4f337d274
z1182ade3ab4ae9b883e684babf6bcb9aea9294fd57a3f7c0da41473d4c18c1cfbb302961baa67e
z52aba20a523811b58fb7160aba65c30dd4dd338ba9f6ce2aa75481d91af6ddb4fd3eeed94c6d41
z1381c74d645bc72d15358b35280d875f5bd0771c92422663326b3f73d862afb11f21e7760ed1f6
z98e7c66772c7e5f800125c7ce5cf177b46e439b3cfc79734316d2347c7ff3c8b290ca37b2dd12f
z9ac16ecb738303b2e1d824a0c4a9f5ca52210642ec7112715188b72fc716f40bd479cc70e74881
z14229548dab0d334e0bbc549f83345d1aac3daee29edd35e400ffce5a2ef672965efb4bca62a4a
zf4f13176758bce8b897add91ebd02b99fc99c65881a63406204997ace190a56f2290e75118f679
z035f154fbaa0a9167fc04062980608b8019107d9876b7d0253c830bd9e262aea675d7948800acc
zab3d51c14f6a1f487f46099bb2b4d3ba189fa0ba1bc227a7806af5926d7edef9c26ae38163025d
zde08135b1520db43bbf0a235ac6a1e537c272554b5c7f1b09de890e2945cf215e58958332228c2
zef3d733d467ca9f199a4e763fb9f84144972ebfcc80a64c48d76fd80a2de33d65f2994bedfeb74
z1d18770761095db4f6f6c5d1db2409a9cde312bb2c2a7d33a5363bb962ea557adf9066faacbe35
z1cb36d38449016941e8e2339bf850c886f589cd7b299ca2c8618419c8818547dcea8eb11ad92a9
z9710802d2442e6c4b510b77076ecb038582ac127fc67a03c15a5a887d9d90181ea95598944cc3a
z2f2aab2ff98806272c2208fd295824adb91a233b281d0e258307cb6644f06d66bbd3243f2f3ab4
z3e64e7366841b3b8baf8cec689024abc47e8ee3387baaaa0762cf985f5ce1e3fc45ce3ed467337
z979620cbde9fa88e60d57e421e5a6f9a023cbfec2214411727e251a508893adb97a12ac0334cbd
z846d1a4def7f4a463b17fab030b6ed09d97f358ca487601ab706e904bb49ac45340b0de09bf3ed
ze991aa20b09b4a7e6940bde01adc2ae5606edab1111304e54eef79a8d038c599b66c22778bcc8c
z5bdbb84ac49bf4ecfac6ad24b33a0c8f67c384cf76d7f4f3ae32a9445f81a7a9d57da04082e471
z5b650baaec8f227461792f2e13188e34347894c95d8f7df8e8d3d97d69584aa76487c6f1e6b02b
zd0f9baadbc4dcd9f265b6a80c7d3db4ced786341a0c5dba41d9d230f5560ce508417446bf585c1
z55da047c9fc56173bb0069dee4e792f908f489c63c314641a1496f64d5e2f6e6544977a9013e65
z8d2939a61fb510c729aed477927ed2334de133233ecb85b82250c91f76fe2498e9667ad1dede1a
zb43c6b791b55721b25ac607e36846007aae6bf16f1335903bd6c09c09921ef9de2be25ff87f9f2
z869b872bd8e0176a126bae9140bc62638ebb8d3d372b2c8100bd8a3412079db2f0de344b85055d
zcd1eee84ebd0111a21ed45d4d3e4d7437d971203c963d1a7f1f95843fcafdb702d7eb5ec4ea5de
zb318bfa488e047f8bfbcfc4c36f5335ef04f9fab00313244a67cff3c7530a25d5bc702f9ce9062
z58459553c4df355366a02b51644a0b5a72d672edca8e62c67ea848b38565d859fc0a369cad3c83
z258c3a42dda506b1ff10aa49c43e8d5e7eb98007941ffde314f594042cec4f43b3e911120f61cf
zdf9ad5236785ceaa28d26e29f0d21cfd482cfeef0ee836ef32f7c39a1ac36330a4d46e611a38f4
z2bb083e8574f84efb237df8c63b0817d6a9d79408adedd59355ebadb022c261a12bbf1971b0ba4
z8343b5b3bcfcc2cddabde2991a95a54d0858db5a857db5dc654d9cff323af345e72b1d8ca4533d
z77803ae1055b6245eb33f930b8e6ee0eae64ae06fe1ccf72eaf779f4df80bda5ca32be4e515de8
z82dc5cebb7af3b92039ec222dc7db1bced7516eeb93422799c9e0a8a00822c7fefb6ae2f4a6671
z634dba09c539a50cb6c200ab836ec32a75c16ace8181ae467bf0083bf17bd15892ce5f6d62a545
z285f93a6f91b2072d1de1191d9e178dade2639699891011656630e827da83de01780277ed3f3f2
z3756279d601098614d5023e8428b270277a6fdc4ef62966bba66b8d6f6dca7f99122c8c81d50ac
z831731f217dd07af42ef2b42f9a0940618939e49e1508e8d441bddd860560faff06aff526631a2
z33fa7394f9eb568bb7cde153ddcd12ff92947dda2fb4f56df443e45a121b9f79b68b1c3aa8e72e
z59e3dc67dfe8cf5358150f2ea2ff674235d4af38248b4a458f4e526e2623094d4c2496ce653276
z07a3cd911c178f639d8be00ad308a6b6c1a0effd95d8b5988d357c78bed43c433e59ab6e608b47
zc20dab0f7cb8a06785cbd17e6d79ee63fd73b2328988a32c856cc5960e5f0f5632fd5fe468022b
z8f98ba65321b1cacde7c5b57c6c5ca187b1a84f59656c4d5be00cbf2c7530da7bba6cff89f6252
z6cd52a5eaf29a6a4e34962d2b04af2704f5b10384980ccaa1fb9c04abd1fb5c630b161168d5d3e
z218a35f4d72d4725729ed84967a64617693d34fe73d60ce7c98e61435311b786344af3106f8111
z81dda806fc75f405c9098941509bc0949aed7ca326ead501915bdda8e0ceaa8e401963b24f195d
z8353599652b7d020466b88e3d734a672ced9dd53cb552a35e994114ebfc5cfc2d8e5b2b7262df5
za6368c32a37b63f19c5e9a15bbfffa8c489a724ad2026732800d7fd43d4c2fc6d4dae36119096c
zcaba1dd525df4348858f6e122ead12c9350b2ef4bc2a25017df3f3684495712c4ddb8ecd438da3
za353f204ea7bd1829e32a842c95860e153ae7d5bf9f0643a87ee6db3638dd1601df18b9d2f31cb
za63f6fce116e1061f6366df4328fcb9335fdd7b05fca98285b087a254dbe24a6c4978e79d38c59
zbf789450cdaf1cf01dbb09d6ac43502c69420f157f021668ce4c2ed1249b9d80d4eacf0a511901
ze93d2d164325e6357bc13d3fd318d95a5f4c287ad4f31f02dce7578d16b6d6eea13025a338a59f
zdefec3f73b01aafb775b6291460662572eebb4a825da80a1b5ec98a6d2f4b7a3a9c61961894006
zb1ea4f47bbdc9f19fba34a5ceefcb0613c434c3c61bac6e49c733c68d46a0f746bd3f688b99746
zfe2aab67e22731f3dc4ca45f2ab5a23e3a94e08deed7d5a33a565d060afb1e7d67dc19707351b5
ze32aa8a4059b3fb37887317a8d7ccc0398d08c86cd84de1f521bce2454633700935b03922445f8
ze911624a62018c6c834787c42e401a195f21f9ed2694189c7deb4237acf96ca535268bbdda46a7
z0eec1ce38cb1d6b18b8e6fd9cb2dfa5f3fb6616d9a0f51035e7204d66df5c01019cfbd9d7db884
z11a2107256cee7ea005953a69daa342acdb67122217767986f73b03c7764bf5379d9744bb14e09
z546233eb7940eb1d00508ccce931dc79fb308a6c4c2463f3747cdf7f53ae213c41578d0ef25bbe
z51cd5ea53a4327366bbd29d2cd6e45fb150aa9be65a0b8af731c744d56c1fbb734471e9e567a53
z61fa58ae48366fd31b84c625e1e2bc6b0061d4f40cd30d90a0dffbdb1935f32c12801b9752c6db
z5faa48610dd356266e682ff7c4ba36d69d50b674b1df67ebaab909d65d19a0400e84b5b909c6e3
z82190ee43367c8467d089113bc7d10b9421a9df0bb7f2ab49a94771123d852f20aa080a444e5f2
zce394070f80a3205e73ccd47e623486d554d50d833c9900f0a87cd0eb8f8ea82733686d5342e58
zbab34a3a06d8438a8f0b223ddbc6e512c93a9eb34fc91879581ad25a72a53087e2929f4154dd15
zc9f7bbe24a802c432432f551d3fdceb0b83397b00389bc644a118a6c9fec872c2e7262b2afac66
z78b248464651ebe453d296244b89e52ccd9eb8ff3e908af7b0f6bc81163e17f7d6339f349b3f54
z516225f7ba3cb21341579b4e30b8434428865506eddad7d76e8982e5dd8659ee604f0e83d0cf85
z2691714827adc31934b88fef849f612f057ceab56c8b3db6470df0046f3ef982998ce575c71557
zf538d97d896d70e097c51fd12dabc28d1f94553f3d99f41170e9a9c75ab5c19f290697021c72a6
zfe5e36c491d1112a2a41e69da1523aac98a2a532023ff9648216847e1e914c509e5f6362b3d430
z221ab255bc86dfad126aa8f16d2dfa6a9827f8fe85371f782dbcbd1fc113e5f31da5ca160d063d
z5a513a15047c83df462fb906e66bb9ff6c7dff5a76f7a826f8ccdbfb4c930fd58a4cffd74122a9
zb0cd789d74848af1a9f2f0f09b473ed073cbda015c6740c8aef4e4164c4ecd26fd2e2f57b1cd7a
z5634b814216f2ae506edf0dde45c972f4842d5f82ef7aadeca28528aeef503142d8ff9161996e9
z0a0a7240d19a3452480c4f8fef8f827158f696548360be55aba5df612af9dff31ca8d8c270ddd0
zd4e8737ea4cc63e833b828ac8f2b549ea0550d472b51877b1ae0d4e8061856a224efde84b3d566
zb522e7ae472bec2b12e8de48b9fdcf3064ad9a41c136c37204c191707f18867563c235c406a4f4
z597c1dfbb4e64f49c94b59e6f33cc78a0e2c9a841c199afb859aa6683504f4756883e34cf621e4
zbd7c5756100e2d5ff89d223374f5dc6b28f4da16af89a3d7471de112870f21fe94be589b26f505
z8496ee177baedd57a1456b76902616e9663ff07e5c4f57ad31fd6e7952d808ed1b89b3c6528a75
z37a396427e59cf8e2bdbe752e785600f90a9660b94778257581a6a1ab2286d225426646cc19f63
z61fcad86bd8eec0c588623de5204130ebe0005ce427ab189476846d182a6165da9ff7fb7cd9025
z6bcf054465ccecd7b9660033199b0779266c7dba86725d0d298dbe64ed6328a1ce32f3b9641dae
z0444af82532cab9dfd01c51a99b976cc9e696cc25bc9263e982cecb3d8fac01ae2130b8b390b6d
z4c84287fe832069f92d6941fff133aa491816f5d6a6a2b5df4cb99fe0129320425e6d5ff68baec
zf6be2b6307a51bb270c3cdf74580945737c6afd1f303425d1be78bf967218286ebd5bc366f4280
z2589888e198a19614b627fad9b1c390c714225ddf40934692ea1b2146f68e1cf33a87aad9c5549
zab63abb581db4cd5ec895d33ea8b11c2371f00d7b76a9f0548511242a5dfc5e0a448abbef72cb2
z6d32fc7de2f51cd1f2146aa4ee89f20635bf57bbc0c6289382765c3c89d5b8330157ffa206d287
zd763f94431f2889c0f0773b76c00dcc3ec69a8a8496f115ec019af3739cecd7bdc427a76edef34
z8b113bf592d8ddd025b8dc3cee05d63c0b6534bdf2ae9e459e1f38ec12dec0072d5ccc06df483d
zecf478769c77133e034b5f2a42fe1ec0ddc536c424d4795711c951fe3fed6ca14a1d59d3cf7f65
z78dda7d83372e0a124c89e9837997a8f15c43a9dbefb6b31c5a917714da9e97c2254231e00d4fe
ze21b139a90f36cd4f5fa708b30d28de7b07a0ceeca112e04cef1b4ec942e7d5a2a2ed52a21464a
z213c8729c4ee6b950e69c6c4765d691041709cde56fa5c6d7938d7202cf3d7590331494d3a6626
z350e0e46715713bebe88edda4a25a2c02978b419ec674e9f3fa2543de562e46f9540aa9154eadc
z0a7e116c5721aa74ad3d03d2714f3611d123ff6de7a32441478f645a7369be9e413b9a5853bf3f
z17f99059af37209e97d558cbe570bb173f21aa0881a1eeabd14ce74038e606fe80034f5c7ef5c4
zb89c927409b753acb54885543780ead361f6110387c637e86a3219dc5e460cb0580c106f98748a
zb79899cf4d0318596e7029a7521c0cd078b99b104b7511868e1a7222110e3952286c404757f394
ze1c89692a28834d8ce50ccf936cb00b588556509e8fff8496a2d3b5639850a42c593cbfb18d285
z360583434b185dc8d4adef281b13125534888a4d0ac8dd8dc0ea919dc338a3a7a0803587ee336c
zd03439a24557e9ac511181d8583f0015d209dc7f06bb2b1f56582026cbd2cce501b782e68a05ef
z6681f3fb2d89a150a87c492a25f3cfd67f3f517cf1520133be1183e57c059caa03abcc875b45b2
zd190a6879781689412fad57a3151ddc26791dfe376859863789d2c3c8671894cdbe1bc27942f97
zc4c800b0b7339c4fea0cbf443665a701780deb21272cdc7063bac254d8ec9093c008d2539cc39b
za5c3454d3bc51519dcb40c2146347ad368a8d68996a1211b81c70c6a3b22d2964a37e4ac73c608
z1ec1e50dea6d00ead69709e3322b51ffae536d22df3e759e6e2a3da8f423dbbfee0de8afdf852f
z2f9ffe9250dfecf4db1b7d6e1fbd41b07a42d09ccd05f253ac76a5babdca5ef1245b86865e0faf
z7373118567f0891abdfdad34f89085c5e030a96372c2f305fcfbaae11cad21256f39082becf3e8
z747311531eed111600667b27f5e4794ed3601503b5d88d03d5c9a0fa114f53e47624a7d3c9c06b
z117b6fa85dbe134a6392e63934dfe9bca833bfd325f333a50749edfe1fd8546f7b2fb4be26294c
z84a2d583f4f68d5a7aabadc7c4f0fb0f9d1b35e19d6514fcabed01ab41c07a5620386b32629a2e
z8a4790b36c063f258d1342928268a7a889ba08c07c3adb59f23f17e8bc1bbd80c344210518c683
z364deea6a18f036244da41371bc8697c4abd467ea8c2b8ac6c02ef18d1620168610a48d411c56c
z2c22ec6bdaf236864d5b6ef54d49e0f0a4461d21dc76b96cf2bf8231b2d3951a91925053274d20
zb3e1fbb00d86fb1e71001473d42749973d12c249a034b435d91ec5d5dff818da0b37bdafbda531
z7c405019c5766dadccdee9facae5c10f4bb940151d03925835b7428f4217aace17212941d26881
z7dbf3af76c256cea83d385b89f9bf079ebf3f0d6011530bf2c4b50278631a9d4e3c047edc883e9
z9b881c9d7e33b0dc1aff7403b05262440490f76dea1105310abdb62e047f3eb42782499a7db761
z91e43f30ee10ebec02f4d642e0cc299817beb2879d00a75d965693cc2454958950a5efbc4e3adb
z0218560cd45e853e4ad339f2f28c70a9af8e654131e89ccf7ec807c4ad145cb14e82f7eca08413
z35039d2d35ca5eb16307b769f384abef2ca2fa91660097d85706d994bcbc82b346f78cfb970aaa
z86c1200ec0427f3dfb9581d397becb6ecf0153cd703c561b253e0451a3bb8c12f94888b3986572
z98a9753c1897031a3896f8b837756605e1d5c928e4d06fdfcb867e386673aa72c590ccb83dbba0
zb8ea36f9da59b941bedee6884cfca8af37e47840442d580986ee48930ea3aff0370919650f7b0c
zb91136c64b38acb2b399fbe42d680633431595535b7d102da654fdbc2d7118b6d5c2dfa8a93352
za8762d8b28e600572e5b97d91190b7b97698be7f7177c3535aae9ff23d717da2dc409a6a686776
z2fc6d7a683a0a33153f863658d74a4cd2e39cce9942170b17148b1a5e80411194483909d50127d
z0e64bfeb934d36f6b830d8b96f0f89a96b123fd352c1d1d75862334931c2bdcc7fc0d10d0699a8
z4baa0bd63d548f7788afea9f83431a8e1e32b5a5c0104d727969e82b089fae0490912f45a6a74c
z6cedbed359b6a6259ad4ca4163f08ac7b96f6c8ca416e7876ef457dfb5718ba68eb11a9d4b4487
zab329bde86b281b504a01c5afe0d76ef083e5fe95f18170b15f28426078bb8f216886ba1fc6e55
zf2e8809887dad3a7f19072d7baa3b64bdd51084a15235611ea294baeee3d37f55bd3ce39c8d7be
z0d9ac268ffa49e88b0d12f888a71e21d305ffb77a2c8f7d794ee38129c2d6e0d12a9294f58cc43
z387a4fddfcf33c0942c5bca99498dce1fab70a9ae795e6b8b9119a4d6815ccafe6712f5e5ec9de
z69675ee64b47d969077b26d00f58a52ebce0ea94e75f206d079623ef090abb90edb27a24c7cff7
zf30c607bab83c22abe4969cec756b3a42447d8a942f2f7ec8c6feb8d35eb3368c1869a41db2348
zc0aef609a7ffefc6ea9827bf4a15bdb8e1389efe672e3f4a1e64c294d1c41cb4829464d39b7d9e
zb6b19ffacb8d5b547a0ce587a02b27277c7a0c878e85f43c55c6d7fb55d1daca90a82a7336ca63
z2cea6fb2b78a7e80a18816b02865a5e4be43423b3ccf3710118fa851d2524516b65bc7fcf7b75d
z8bc1272aa4c32f2bef640bb7257974d992b39c622d6868da43da22ffc33558c5430884715e1651
z876f91729561aeee91b41d288abe45cfcc41542f7f77c00304483326bd374726da112c227efc25
zee256823db7b29fddb955bf4b46a6cb3b969c43e5b300a65b5e4dffc13c0d4b3889af9934a344d
zb9f36c64657b2aab2b8a355558c16ffede9ea64ff1f93c4ea102d6a783f910c1452fce594469e8
z406f59127f96981153f3c08c84dd06a02c1533ee9962795791df7c48e7a3d0a1eee114510aa344
z95b4765029cd506073dea2951d7959dda680b670abe60d57917bce0734b18b96b06ec3384784fb
z1f9c7c17dae03315fbce26dd493673e6337d35a8add128db9d10a492b956f66ea4472b4ca1e3b1
zd6c2ba628f3b2ad6401f3d2539d5c2870a29248ed4f3af6bbe3a6a9857166d8898e2630f892b06
za4e41f0234c34219ee9502a1fe07538db51874fabde92df5ecd5e164367f9be67bbcb4a3a98f98
zb9a0d535498b9fa9867be280426b69be5eba1dfee4810ae6743d14ab30b78a6a4d4db1a8e350ff
z94260be1ed1b75f6e55637040117f76690d9fed6d748ef99d559c4bf57c9f8af528321d315748a
za4fafa4c5b037ed5e1334c3fc51ecf218948f600cfad57e26135886cae1ec6730c024e19a9daf6
z9415bd85e17e1dad22cd49f0304c6da02013622c2e382ae7faecefd83d4e474a3eadc15466c2cb
z37ac7d9e43c9882a094fffc493055cbdd5d5da254c0f9b265c7d8f1ee0e72c49a0fc0f316686b4
zeadcae33db8bfcf61c19f90ca58f11f47e512448738652ff6b17d03b723a6274287f0ba8086c50
za01eb5660071a0e35e7b2ff3b88013aac189c700642607c2c42eedb42e88ed66fc8707e3bc987c
zbca02053515507e18d5457d7d2c32b12bcd6603038b98d3810e725ac5ecdf5ec2406dfc7b8cdb1
zc86c22b8338f6758c4625b2f8f7bea250cf87c0e31e9466e5ca6650251d6f26427675eb08f22cb
z7136b4027f645a09a784c7f4cddeb7c63968255d447dd9513cbbff5847c108629ff8c1f68d9ab3
za948ef58119b34de230ad67845ed2cf70a0bcf02149b5d572f518881ae1b7db0692a984b9e8ed6
ze701d0b0d659ece7859618a2560451796a68963b5a19069c2d027d7d652905609160a09c4f2279
z1aa3243dccbfe669bc21feec8cc5a633e1f20a74f40c1f56d2b7aba336ad0d580404ebe27c7893
z0ef3ce313e949600a06445f9030cfafc38f9b13f9f090fdd7a11c9d12fea1e1512875118a43e49
zee1a6bf3194be88ea6a4dc09c4e11b42399329105e40134e26d435404e7abf96d596460a89d0be
z9e7651807eeef749baf127427010446bfe712144dfc78d4a1370337e873e348676ee2aead0d014
z3435a9f0a42c481ddba856d9df97603eb4e500472ac3819a69e54d6e670bf2e6db2abb91b96dd4
z4d86f7c3ee073e4420e3b3ba6aa9bcc9957d2583c1dbca84bc3c1dacaaf79f220637fa53a462ec
zb8d3a1896f8afb977705714d25fa5f70ef4feb142573d8255923d4cd5f9007d485d2a0cf1d9d7f
z411cc7b62870c23454be9e34d0133ecccca6179b304762c54766313ff439c38ff874bd21d315ee
za185afd0e9182e6acff486e8014aa006b838e263a9ab52d337eda61424a658459a5b767c762d98
z75a6a4186004bf1566c20f3ccbd1ad229c22ff7804afa06d31e7c1bad4eddc18832bce66b0f72c
z385a98e6f96c6f191a041206d98058bbfc2529c5d011a723b47522a4e6691c446c455a0a3b5b21
z8432b42924cb04aaece589aaaf09379d1f009ebe05ed3412b40a29c485310d0df43cde953be7f8
z06c379ff2d8ee85533247b825fb593578ea62fe6d766a867c9967fc366648d821df1810338e7da
zc7ce3a12bf4de20edea58d761cb7cdf9be09620f3c9cc80eb4d169f6c1db19056b372662b4575d
z459e25d4f22637ee9ef4aad1820e621413bb135e805983cf38705edd2617d5550ae0d49878c05f
zebec34e9a53afe9b8c777f26e5f4cf17f3e295766b612ff10046ba87819afa71edfe50371a1ab2
zb66ece89924184b087f8f06fe6bbed01d7b8688cb3c797e218f343565264618012054fc7e78143
z09584c9898789b3d39c050f0aadf3e72200f6f6ab7821b5f52f8c19d31945c3e0f1786b1c7b318
z32b954bfd32d6597ec11cf1c981d42c54b0a5d2de3a0fd977e678cc17f74f2c374686648420479
zbe4339e2b42c8dd74a3b4df76623028007945d6b71a06f66f7f7b615499ff2a606788ce5deecc6
z1448ac08803c33f7ca1a223ed5daaefc89a80096b4791b3ff046ced16abd424b3cf64e90529293
z615fefb7a22d34c86258049f2267a53cc7aaf01dc1dcce6b8bd034ed1208717595d854c5b189e9
z84d6c9f1e21205b1c2fbb2cd722a14179d635b3e94637343722683f976a5b4bcb1dd2ff92cb057
z565da9004d9766753aaef8e8a305e4da473cdb5daef048311b361abecfb7489b487e03ae7f33ca
z3bb219396785b1deca286558c7ed90639814e14cacb2c96f7996d2e7f03cee703a6c7e05b04bf8
z791ef6b0acfa989f3d01b543c50ed39071b174983fd290a8985c6fd1df0d47a754575703307fd2
z2db09ac83545eccb975fd0025cb70010281e6736779e00a71a1238d7b323d4f5917fffeeb66aed
z3985c81aca5610f62765930d065c60d92aafeca47f176b07b55147401150fd708a1a30ce261578
z2212935f0940490c87dac26cc6dc661ae1f95e1c6db757a4a842b060d1555e4b1aef7ae3dac554
zc28b1be0c880f4770ac273766f493823f8da5b829caa8377e44ab587faf02fc14a9e88f0bc89ac
z1d5afb240056610332adce0f748322071fb5463db7dfbcfba0b3717e9a82126bffcd2a496934f5
z34afb3ce3e6d3f04537df1dea0dd5d712baa52e548457db20c3c8003d2d9c5d458b9c5fdd99a97
z194d4a800a02b62d7ba8aadf7702d70f2383748aa57cfb98568034fdad5341bea5c6cacbdce283
z166fa2b793cfca9a052976ab0b7832d9e6a2ab4c8a04e70ffe3304d0739f71380256e4d06aff99
zde5b820ded2fb9c15e3b3909d8a0d2e1b575fe59fdcce5ed5f168c0b43d9d8a6ef61a70d03b069
z21349bec76896b3811beb75c91687862fc3de684d785fed44d2a917fa733171c10b18eb5bfa889
zb721e092ca0ef547b02071af04b5a480bd7b4a60a654d208032cb4cfd90519be87ac9a90011c96
zb33284f6f6985ad7e612273ca006e00175312af21da30b1a3c1f9595e8f40f2dab68279e146ec1
z74a62942b4a591f6ffe7b7748d98e2bcaa6ded9a2fa9d0fc0bce85b35c53132ae27dff5d2cd720
zdfd67229018f3094ea9a1df8f48749fbbbd30f2a509d709ab58e85fe37e6b23c09112f78eaa251
zccbd8198a498ef47b43eb93511216e079ec9d478309649b85a3f34110d151f81bbc4ea553feefb
zfbcb197a22b96c687e920469701c7fbffb6801863ce33413c26a6089d8a33847bfbe6769c31423
zb13769ed63e7800ce17f7d32603979942cfa198d8cc1bb04772e662fa6f57fc3968575006e8906
z5ced0c354a5ceb0ed21c9444f609867109da5a5d83946ba4bf835ace04ebf5dcdc1eecbd812bbf
z757c77b5b07fcf4905ae8e64a9ac38dd8263115d6de9c5e7e3101d50f200640281599fabfa81de
z59118e4926a2bd2fd5bf0be00115afec193e99e11a3dd7f35cc123e7f69845a2c4c33c53e07922
z114fc59665f463500e1a276578f63d9882e48f694c265ab008ecf01eb9d8d79a06b2da630f0a6a
zde6cdebf888cc7995abcbaaed91ebf3ecf62528076a86599556595181ad96525b665d0b901eaa4
z36fe2b91cefd241a4d5b956ef3678f59688f52d733652defcd18b99fb05b7ef0997775fee88056
z6882332e50cc6694b883e3a7ee48f3b0dba1b1055e8674b01b39034aacd7dcf70cb6a3443818c1
z49e68ea530e2355a807595d0162864aaba7346e28714d276016b8798e3e23e89b5920ec948673d
z7f18e3a95153477b15d7886a7e12a3e9b34f3d6f5317f04c092561a082e9765faef90dcf2c9912
z62ad79b51f92dbfec4802fec354b251295ca13621808e237d4e23dde9212909ddbb47e8d7e3aa6
z08c607ea8c935080ec68f43ea801bf33e7204fbed3dba66c3f786b8c664611b09fbe50a3fecc4f
z24daea9200d31af2c49be856738554364457a40b21c971937d72d8dbbf2f2221d0818e20436cee
zf472820a687a8277a342b9a0865812463cbceb5e6f1371d938fc5b28ed0af274b18325f108d8c1
ze1640183368ba3235c7c8c47b8d704ef26355ed89cc69e060dc6fdb793ddbfff10bdc2e9fc5c4d
z7e3f548be2cbeb3b344c998eb6c39c39e884a73ba8df17509e35a9189397e13081252ca877611a
z4a0a3fddd3bc213f428593b5823e2223158d567b105fd590d8fcda6d156320e5706e2f8d2de86e
z5b65edec35d847673276754d682f45bdecbfe088d250947b4806f065b52d3684892e0dcded3e4c
zb95975b9761176a279e223d04dbbdaeb78a3cb250f9d7ba23e362867a6c69c3312ce4ffe6be268
z355305bf78f7315308da217b543d4a6afa1a0a4acfd2849c1315d7fe3bc1f51b9481699aaafd35
zfd45a8f668b17b97d7a68e4eaa5d366f1c58058c79783c4f79cca4310d685e98a3c3803c34f3c8
za64f959f10d7696903c8fb4f86c9b758d2b23126a5662a9a8e794c0279f74fd8f405ed03850dea
z6da92a72281ff59004740e1b7691001e12085bbf71d4efcfd89216aa6798c6687a4e77c4132645
z92bdb98b6410d5e4f48026ca2a95e04c88c98fd4c1029c561c22c873c4c75e59ccc91f5068a447
zf0530fe426f99c93ce915beb21c675f3c9d9df45276c4f209957c163ee48751e84dd4c9f66f9ae
z5772d020b996130cf229b62ec526b709476f004b9fe3acf4592b871c64624d2bbfff649dc943ab
z941073a1ca42b251034153a919f725cd1a6841dad8c03b7a1178a862293308ea168c91aab240d7
za23f422c7fd49ca114280e2d7d9538c478b0a7b93b32485bc94199c084986800dfc935e8cef492
z5dda1f30ca39d4c988d6cbbb2afee773f91b3a82b2d69d237ce3061bdfe478356b04880edd5285
z352a7bc6d592429b246567a1c0a1605e0cd57821311432a8931393ba0d4232c190d31a01b7834c
zbfbaa67b27df10539c5236da3bd828ebb47e5f3a7d813dd8e1f35db32b7fe6c469f96711e1fe65
z7f7238c6df4c033ac3b4f956eceadaefbce86da63fa69aae3b9fde377662daa3417db1bbbaccfd
z20a8af9ca7b8c4dd1859db17ef5cd16227bd00fb8c37ea61c63b896227c75be4e09192ce642cf7
z5406258c8c8e67d5cb7554466208149b2c0e3bb0decb1cd6c0f9d8eb181534d2f6899ad6b4ccc8
z3a39d1722e31aa9740e25e562da8d2348d6967b74ff0482b1257f5055eae74b5b07dd86e194a5a
z118957c1a4d9a823ed8bf6ebeecf8aa9b9e2c2071b88011227c72a94f0f3ddddaab7bf59f5a7aa
z0813b1b4d638eabafe34204b105c025251b0705ff57b2c7e18b9d0194db47360880b44888e5b50
zbbf1e5be575f0ca7d30f4bc5dbb82e85e164a79f83b3521bfd5e5314e14496f6be053c2e8f3b65
z8688e487ccb8c7272e30461beff30603281561966308fba08b0e17959702eae8c4aa29bec3e597
z4aa4b6b5747b22f6752a6645e2e5f15ba9412e3d7585423f637be41b953b2b65103aacb9582aaf
z31cb6b4d934dc60e672cf25c6e45fe113d05415e0977eddd781cd151673bcb31b9bedaedd56cd2
zd10c9720bf10e1311991e234ef3ade98a99558e1bc9f70b42c09e9d2a784af30fcc71c6b1c6f2b
z56a6237dacbe2317dfd761621d7767ed05e5538f037887d79803a302e5a257c0eca5a39e5d1b6e
zf7756b205c5b1869a97de1ccff67c3d1ef40341c620678cf64db745de812a4cd8731773833c4b8
zbf50fcd8a32ef17b4917cb67666f9b6aeb7612b72a496861b3a524dd1f29c2532d5834683b9b97
za5e4c67b0052a77263c2bf26f4797a5d29e610df349db0e2c82d1c44e9a4727a825014a0e83627
zf54f5c21927699c80c9c6d84de69d6f4ecdd878c5d103b404c19ef67af8b3a163d7ffd80597885
zcf528033172e4bd462d8ceb5c22c96049b59b328207af415f784eb7fadcbad3f9f12dc894f56f1
z3e5f6d59dac515c2ded9934c70cfa373a702927ad9a9f3167af7e703eae1b66daaa598eea860d2
zff76ce4f28315b3bd8c24b62f030385be36a89afdf54cc93bd2c07f5ea657f28931e68d58de817
z90096160a8e62d958a2335a0087a1864ddb6bbe94a8cf47c2619127192d8f7f4ceb7f511b9ea2e
z818c7eb8efb1dbc1efeee8286f41a5047fe9a6a44383fa4b234b45a507a2047f6574d018effc72
za50ee56336e9bf82c208abd1430318b6edbac3ed5b7d56b8d8499b1201c895992f59769c482515
zb39774afe888bc1c8137bc79574b1750c25ff470bc9c9f6b22d40aa1138b4732ea9abf496ed940
z625f0ce7909f916246c1735dbbf3116de4b3819a361b1666076c5ea54259156d3bbd271947628d
z081a1b63fb05ae6c51dc0e96d6769950975b3eab333f97a19eb457da8c099bd50a285af1974ac1
z423eabd827691f23e6cd5ea642f60f4671
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gigabit_ethernet_mac_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
