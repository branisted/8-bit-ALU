module alu_8bit (...);
// TODO: Implement top-level ALU
endmodule