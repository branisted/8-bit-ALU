`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1bf3f153bd631387c118a296ca10cbf0349426
zcf2ea5eb241fa84c8ecbbf7180f10eb9ddd4966d421e6ca571b198ed195474578ea51160ffbd6b
z0f73216703aef2bba31d04f6d0877540c760cd2535de412f259f7ccb8f261f548081500194536f
z61982df641d53c7a2e879bf46dee12963675baa55723db72b3334fb3f3277a5def35d867003b3e
z96288dbdd29f8e098b1a338d244ce21565adc0e33ce2f3e05aea0c8b57e1c83ddf2fd204229b70
z8fc88ca804d08078a36a1561701b9949f0c4b5270a2440f00a9b1e69536428913ba706bb862626
zd17d468247b8ee68d04933ca35936c6223bbb01314b6ba7a88fcfbf7c1d0a2b197f2ef84b6ff5f
z28b98b5585c7440a0d9962a6b36d7444e52a9453dcb782d57a7ba27f6d0d5b8f36f34c5cd6c005
z3e1b09612c08e216d79d5d9d210a1ef37e2c70f686f5c87f13f96866198fd904b94c53c9a82a31
zf588301331b0d1e87b06e012eb5b44e7f2f7cce3f14a402e908b52052ae700f4fd4d9c1b8c34b2
z46bc0bc7363b762abc3a1f4873bf2c973d16ce19be961bf5eab9a61bb93acec0b909887ab4c30a
z8271ece745ea0533f984ce317c7827f896fded1c8f621ea493c3903a10d342cff044b181cac7ae
z2d241910a64ceeceb27cbc3510a350881c5ce3523ce5def32d2f222c056ecf68d70d9c90c1603d
z5b6db740c68549dc96273f519975341ac8c8cfd1e58d11e42f4569619e9745b65a3e703d94101a
zf07154c027349f759d119c978372b6c0e5fc899f1c5b285ee3444d8ce4108163f124471603a305
z003f1d13756624b7b461bf6f2e245d1d2102b181b8407028e7cfd85e10c5ee97665131545fb3ec
z5f69489afe52fd5a333a1f37e8a4eaf45b848298067525b0a4f08d6edc6ad64b5be7ce2d018655
z72b877ab0ab32eba326e905ac535737fd9019f455a293db2184b4a14ec35b2b5fa99b2f891b08c
z7172152f9bc1690ab9b0d7207c5e1cc25abec89eedb8455a23a66f51e458c60de26c4c9244a85e
z075ce8af06fa3eeb7dba7bcf9fa64838c9982ad1af77dbb96e752c93e753fba47581ef20380ff2
z7cbef6e344946ac3a20d205b0acbe5a9690016a598d3a1374aab52b3a280ccdf3363d2e213fa5a
z82ec4745576c86ac125ee2573d74312b4504dd3ed90bde14da44cfa69e48215bef6a94dfe0f2f1
z90d74ce361039c1f2f35ad5e8fb5a0ec2b523851da44bf1c7af7dab50a36d226fa768b54041162
z09fdf793866dd3439a54ef0f65c820b5d7926d25131b18f71ade18cf886410d788a16cc8e1b0de
z9bd324487d0892fe515f8dcedbd37187e92a91de50bdfacedd916cb0c3d583315f6d1c6b6215f9
zae847d47dfc2392c428a1f5fdaf861679b47f7e2716a268552aec55e50bbd08a95c25e37f3d23e
z18533a076c3542b5151070eb17e1727320c807e7e694a638a9a88902bc02f6767524fad802e882
z388d994a211a733eb4147cb37de913d61fb60b61fcd0471cc49049900e9f4ef0d5da52f1dd0201
z7d7fc65cb6b5b6298744cdc4e1db50d69c227ae12f57a413c5354e21cb41bc47c635340301b8fd
zdf6181065d0cc37c453fcb9da6e497e37f8c5f38213b4d1e0d24ce200c6fc5136f07451cc97514
z0b58320b818a38ff410c3505b6c052d8facd76ee162c73b1b764bd5785556d48c7c4308ef9fd5b
z692af89c59c3914fe4309848d670d31621f3336f2a01d90f051da13a5486af94995a735fb598d6
zac8f9d70e75fb7c637185b485dd441f96034b9db33c596324459e37397f114a503d29874a5369d
z3d2ac11c7331b6a5dffd7ddf11fc229b162ddb52adde3712142251acc2af27d60349699d5d485a
z91c0da3c881848fd1ed1711af325eecc26b141933b9cfa76f656a9add75ecec65ff83dc83fdd01
zdc952c2f75078e5e6c47135e7e45f9e68185bd8e0754f29b27ee4f4d3c567aea59ad8f09449c60
z1a79726a27ea8c41224968b082215de8633d4dfe29f74c5c5dda914da6badcee524430282ce7e9
zd73302623e5c1544d0bb14fe7e08cbbc07ffd93861a6ff281972d7c92deefd9caba97817bf980c
z82c8c952feb4e34d17362d58f486ce18036b8ddcaad29758c9665bc650c00321818cf38eaf3cbd
zeabf389d54e7d45e6f4c1339e65ebb54a7be5c78125dc2e2e7c7dc091b89ab23fe46de7cd1b5c7
zd6c85d4633431617168849a39463684375160e6ac8f0211e39faf4f5e34454ad578c5204a0d898
z9513bc6e806e200e13bdadddd694572bdc04c6f5bb2bfe07b3293b3160982e4a5fd05c09bd8279
z2a3f0dfc4a4f64846467abbf32335132a0acd2b81c0e82bb5c1f5f2a1a7a62bd914e54b85ab086
zf135df89afa571a95fc20168148e6b949c9ed91ea411febe84a21748b72a8c81c67cd26a27e6c8
zc47ad3b0523a3124d43f307efce486fe55ea4534e209cfff65c4607080774f545387fc63e6d828
z5281a08bd297dcc1e83c5be314fed9cfde488681e46d57dbecaea114bda44d603be984538f93b4
z7f47992cb1e46c1174645ea096c05e55e33470b2c992b7d0c5a6cc4bd48e6256e8f6b6e3fa1653
z01d01d02a9015b7b7b81a2c0fe938f94674577fbd9542a7bc99be7781b394b2c40d4aebb455b7a
z64dcd37897ef858f031dcd2311d93c054f7d5e32dd04167722a4575a2a6958d9b0f163df53467b
zefdfa37b8a2127df87aeb672dfbe17bd7505f8ea75e4d1912cd1d79853ff0a93733da1f3e296e4
z2f4c975b1cdf6aed2c79d1b8d62fa8c71f42280d7b9fe48e8dab741a1f5c551e66db2ffaead10a
z12decaa6c198bb12285f23488cb32ec65dd544a692883f67a3bb5480e0d63f193e853e3c414345
z10c2882720e6661fa21a029cc35076b552cd9642eb6226ede7e4b656014528e529766395124c47
zf94e6a76ba4dbc9a0b07174a9f00622e572f2637339580a090778ee543350b0fcc4a46245a117a
z31a930a1b6b7d5e47f4368392c27616a69e62e9759a69530bae5a2bd5a411c90285b26e6f86f3b
z8d7b37c1ad591aaf85e3960a2fce6cfdb73f35613b31e800a7131729534a29954ccccfd8cceb03
z56e047d27522110c0078387c35d7e29261513282b21ea8e0e59e1eb247a0a9a03a751a2fc9ed10
z3a87a53c4b88e4d61d8770fc4c6ec3fbeaf073f7aa7b959d7b29ec7869cc218303a27de50f2283
zbe20ed589bf6b7660c82a20ef1312470bf22f7aa4b6b6ac58a783b1e106ca37f972916c27cdb7a
z7b2c691d95425275435292e6b7b496b94d85a0b8f4b41af7720ca0384b3b385f7cecc8061ee417
z3ca85745317b97c09a60fbaa35fd7e069813b136839d4cd433432c9f6ad7545fbc8e3f7fcfa3fe
z1281e53ba01befb8f88b443cab3a01475ff0e7db5e559d85fd751c5e4a13e29a0403259c59d5f0
zf9c88cb9dae249ff290ea0b7fed37f7032b50bf4f10a507d64a3e8b5c08be94b0df59608137804
z4cc3298da4323d9db1f5aeb95bfc4f8fdd593a4a225f305fa478960f2cfe3f2f94766b5d2eda31
z1865b8e0f14bc70369d8bb09cddfcf7f1d0e45ae6b77a9f9068f251376e765e0d9558e862d3ffc
z356b2d95f531a4b5ebe182468601705fbea9cc95b0d9a87607a2c86e557124aab136a1b7fece08
z818752b290fbdbd464f7dea9e04fdbc1bb4880d5511fb6b7722f5011024fc69f91056b4bc79cc7
z15b0fd9396b8a4302f279d9f16d310af268633b2839ba3a694383a4177014ac6531afc17acfc34
z962522da090c6fcf01302e2e9a494b5bd9b31261c8cb149a4c5e8a36307228355f83687e3761be
z27724ddf83907108d117639da866b8d60c7a24998be46c2436d3eac9d08196d09bb8eb1454b6fc
z69d8e9213de39d4dcce515480017d6590cb4b98446dc380effee3fbf08559dff080dc1d453217f
z36357fb398bb98191f6bf8d07c80540143aeca4ee0ed47844bfe4e2212ff3607ecba9d59f93276
z904c22573b9acb95cc74b7a1c4220293a62b14e71efa1ae12c5e2d54bc81ba3ce4738d8f764cfc
z82bbb997acd18042775c2f0525626bffae98cdd838b7fd955219120b2b882e47ecf31d61992260
zc79264cc0765bb2530e08ee3076492309c3072e95a8ba8ed39480e183da9cb155344f5600f44cf
zc7eba9ebcc595656a6f2b932933087883bf46a38c2b934ff22715cf5abf2e2feb06abd79ce8de4
z59ea8e84d84fea0022ac85a51819955403107abc92ff0aadaee7f0b44ba0819f88065a48ba0c2a
z27d6270e115e5feb86af9fc05e434498b457512276eb89b8bbd128ebd1a7df7e7d37b0c03a0604
z16397f4ec64195f531b9c3c9dc867ff9812b274f6371315621b89c18a4ee48e55fb9e9cc24ead6
z662de80be8ccdfedb5eb69e5e742b73c20ae022adc5339c48a2be49b475c58f5888a39ee374a7f
zbcf8a7700537f9876a6c8263a410a3d1c9c7430e03207b4b54875a57ba6e250065cdff36a3e77c
zdce3dfbf6d3fe37d8e260f8f125060eb7a95f5d852d32f8a3e910fdaedfa291ff38308fc3a37cc
z6b1e7f74cfe3fd08dfb3fae83341c828c77832626fede2aa3093517e1b8b9cf632129ae739fb5c
z95cfd5dd49c778ea125357d284e17d160f93cdece0b3abc193a0648e381cc75129c85392cd71d4
z71bb81051429800b64e0cbd9aec1c51b2b7ef8d978452e8f4778e2563dff6a8cce6edc398da1b0
ze3fe4111afa576bd3f0e49c093fe82bf74a73d3fde75518cb7b8b6c5c1303108c3cd4361f2a6ae
z526ccf2ff00e7915eb263a2e9100c08ce515dcafcc78097c0e489b69aee8b8c26ec08cd015c7db
z90f89db3a1214c05b43475a58a51890063ef63025b2c9720f59c83542c86facc6d4fffbaad6d3d
z1d2cda0f9f85c63f46c2362f17800ff4dc245fb2be7a070e60ac1535ba2c34f95e71387ba040b2
z409ef523f860c6ffc49b6408a37fd3d06cf39968bfc775036f6ebcc08406a0802eb4a032c93515
zefd114f5aff092587912932ce08c43b3061bab9f3f29e2bebaa1df9648db4b0ebd43f13620a590
z95763eaa6524c7b8e4f6581eb99e69b65f13b7494e0cc486ca2c59ba31ed27439242b0a868fdf1
ze9e5f1543c0e4e2f00d2456f9dba246237c5cfcaca3b6238fe37cea7e5dd398e005edb5eb9f7c7
z2b319c44c330b57afbbed72f5dbffa19cd0b763f556adc9dcbd53b518a6c89f4d980d1b76db613
za21384767170fa71b335b4c237a3cda1ed9f5cc28676bef2af568630b18f044bcaf5512f18a6d1
zd81ace18d2dc50bd1785ef27f703264b60ae05e6cd776a2bdb0b178a28e04cffb8b9b6a727492f
z1c16f7fef4176f21f466a50b7b2ebad9b5167b378d84303ba23b9adcc10eab24aeb00a728f31f7
zb43bd18d7618ec5f4e5832687108960b521cb2858f06a7bb0c87c865f452c195883a2e605e6b70
z590a22706368ea74f22c6798b5a36bdc3f58c37fe72ffc491e788910d7429520729fcf168cd82f
zf4b41193a857c06159d8d31af4bd4ad00be820b61db2c67799e6fcd532cdf11653b841cf9b6437
zd1488e0b2312027e2fb0980c5106df58b718d203f51bfc9435ec8e46622e4bed60b9a3ccd553bb
z8cdab9bb363b7eab37667bdb03b21fe248ed2f93e0f91d56deb18352180f066e5a48babf274c2f
z0c75fc1eae0bf75f18d110231f37701800d3943a12d9b6090f92f184baa1ed4493d4b8efb1ba8e
zc4e22acf633a6920a2cb4ac532331f1e33c40496b2e3a3e31c7e293b52d17651d9f523d3be3c21
zeabc618255ef847aacb1d1b6efeb383284a0507bfbb1cb9bea5ef5dc0d28d7f2fea8df57adf506
z95cc99ba19958c3c92d0635f72ed47ea40042d86945e797109f98b7c068bb11754c43b351cd3e5
zd105cb2bcc1f4b88b2c14b549e2562acb1de77aacef980ab7c03c610cfc7709ec070f8849e8504
z49f74386b9a382c57b43ed0001ca9007dcd716a4a66fda28c69d04c26e6e308191627de2686376
z95597eff3e85d838e6e116e1c282f49f93d028a100cb124612c3c5bfe0709d5b00523e26b6e516
z7194d0af484db7af3b877b582d832472dc617b52ecf459680573d09843f22ca1849a3b2bb9228a
za6fe3dc4bec41ecabe3df9c2e4ed926cf57641a88954404cd6d88ff11a224f7c79e4de5dceb98b
z88b34837862059eecfa676f560584184884708522391e45a79ecabb8fa896d02ed3564167a9d11
z94bfdca7885e280085f6409161bea665ffc48dd3948d1f87e120d641a141befc6158fada32da8c
z4b28007146d53b3def4ffaa16fea5ecd8addf4827110fe5149d6042b87cc4b0258cb9d57c37a5e
z90efd6ff1fee5fff34189011373902849ab7f4e5415101196b52c4cb020eb2f9c69b613f1c1ef5
z2cd7050a151a3c73afdc802c5bda974bf3aa38ad9e5bf69d7a1cff6fffb09db852ebb942c7c86a
zf9581f091547816da363389a06859d78f5c99868801b22e7e1300e95fb1a59222b904b31183373
z917f2ddd8e2df8f0fe1d9987557b14463de5b1379f6d291a0826e0da95ecae76d3e87e0fb7a34a
zbfaf689deb9086317b507815a39fbb729211be71f73fd9d432ac05069f96ac290316ca5cc8da2e
z1dc65926e3f9f826e26366f1528dff04de7cc48bc4733e2d8ef59d66ab460699092f6e23ef823e
z0491139c688d69f6e421b7f224c5d2e36937bd60424a946c3d7dbdfcb535b0e174186179a3cfba
z017823623790c7b4fc1726e6bdfb2fe572a852cf51bc6679ba0d61389362742be9651ab0fc0f5a
z652e2419008cebc2ed10a9e04cc603e5a7062bafe2c5d28ebb3b91c38d43d848cc59ac7ec3998d
zd4b5670d003a5ca1c083401675a849da76621dd2234f9a321c0d8dc6af9e3d240f4c0fd4ed8efc
z0e93e4961a0c0b11ab44090946267833cdba4eff28296ee0e68eab1c20ebb1b132e291bfef79b8
zf1566a420cb8e8b30d8466c04127585113d7f8321bd1d6bbee671e45b6e747eea51b54d508b84b
zb8ec071e7cadd7d3353bda0b0f484ee271dd6b1b8d2d20f1a91219d963ab4fc932d09b32a8e510
z94ea111c2e9c26faee3aa80f2b7c4b9bbc664294ece582841d728ea3a9d2fcae9e55f84f571880
z25c36c3f79d7bf284d12be19de199414f8fe3a02284268c9955d890014366d23e807bc447bd1d9
z3d1c09fb48d88115273f012f14f5e8f1970e5e44b19452298ba0e0662fb961a037a2293be32f4c
z9f5f37437afed5e9795f11d86e4d7d2d04f4fc7721760686fdecd660791ce4b95a6913c9a4b076
z9745e9614b3c0348a39da26636ea3602105d162ac358a3aa7bc8d7e1ce1995b522b72fed3547f1
zfebc63110bbcc466bcf4a9201b167b87d13af35554fa5592a879c8b6779cb066a23df24ea57476
zba0724f99bfecdd207bfd324bf24eb5e3f46652687bde9a2db2e405698f1c0e8f3ca05e04c0d53
zf99b60528b321708a1461bf7dedaf0064407b387c536f7f1592d3e975bf3b3768636a7e87dc000
z57f709f59130253f573af1e870169a788f1a042510dde11ad15cf674987d7bf99a85e4c5fc5a91
z2bb38587a3e6f8627319421093797c3b6fa3d57e91db61f3266eff1a6dda842d75870ea943ea76
zcfc2b22dcd004a2984cc778a54b05a0f5cd2ec1df296430ae4612a6c32d67b3bd8f717da573984
z7a86c0d1a013e53c046b9600d9c6fb164f945faa6d63e5e93ee2c34354175b69776c6797a64abd
z1e597d6b29f4807950370ad915009b5787119c64a3e5d64da382377b2d2fdcc92e2fd0402de2d7
z8a9deeff24f997ce1ee0a1bdfeac1f7356c353ed58abb9ef629adc1797e774bb052cf14a2a8f84
z3fc4fe065b6815f6236e8005fa8b0e63fb16bbc5d33eac8dd08053c5691894ce33306c1c349603
z0ebca4abf8a4f44d79eaf35d987870c647512235329c0ac031b895d4f63956f3fe0b2dba8b1676
z11f54aaf684318414590544e06f62194ca6e0ee697b35956dba445fcddbf7bd44b4b2d8bd57ff7
z3e32edde00421670889d91a1218b0cd58e35eb40bf27bbc7aa141c5d9c54292627cd38b66e04a7
zc35a307fefba7644b2a4fe4178018adb132785a3c85a23fd8561e2afa061de4a8b6f31c346c3b9
zc54b3bd8d78c7cb36f1770803a6a7740942c00a0bacd3a81fb0cfbd49922c31a175b47f87b2a8c
z5495ef94fad6e630ff4969a6d630f1668aa7b205865c24153576af35b01ececc7c97644da80af0
z494678427e5a80e8d3530fecf8b7785077d3e9825f1a23bef4f92dd34d5ddfc1c90afa5f5ce026
z07c56a0e8a0f090a7c43333f97f8019e524d232ae8738e36b1eb80410d15a205e013d7d1febca9
z2df1ce5d3a4e0e1d2dbf5e82ce736c37ac16a680f699f7603e7e87c720a7b674beda15bb5ea471
z89dd4ef5adb0b9c6b1ec0a6ce4242dfa01794b2d110c300e49d5d4c3f2471601e6c404890e9058
zbda44ca86c1048bbdc291dddbb4609bc40c7053fb67ac6a4ede0e74b78b653d40f5d5ac539503b
z7f6a5741bff809eea9d6914976e3640dc9862acfb38f2aa58d5d6e98b6a964aeabe1b76b25c21f
z4414115ad7645fe8431f00e2ebfe6915dbc00ce2cb83b344bb1b2b2b602ee7b61dfd5892ac56f9
zd0dd2547a533a6277c430e55809189fcb702c3a1a3341508736419a613409bb3db06deef360e04
zac01e48ba7cb374a1d6bbdf59965fd680caf1be41bd5d2786a1b8f9fe0a24d659a266d1360f764
z05fd04dbd3c453ef30aca6c5cb978ebc484f0e366e8a7f03338e9039d98fd6c3e596b4079120dc
zdd411fe58172cf087ed140fcae53782d292f267568d26772eb3e448bad2a6fe34b46cef4c714d5
z817bc974ce56af8646134d19a36a52cc936ba07c773828cd0c9475efe22963d633961188ac7d93
zbe6a9ebf9918908be90177dd9614f267f3dc67b0a5ff927c996fb5d10b388167d23ccca449e006
z53fb2e2a2d6ffef2ae944a5a7bb853d7ff515dcc6fbf106dad41ed5aeed2dbbc2ba909eba33cd8
z98072e0ea98bc952b6616dd06d5b01141bd1dc87a2083e5ffb64f2229474e066e15c5483c42258
z605c51ca96d751e38406d6be20979eefa6a54edbd88a7f0aa4d06f49f72078578c97d2e8e0f93f
z02f9a11a02df0a681d01537d4c54a98a39603df85011e9807680dcfcc4422df1871c5093c8bb04
z40d334b927a54afc9ccf3f60ee98ba494173c56e8b9519cb2ad3246e4ab474a39890115238e111
z97a43c4208aea4a97392ceeffa04f8786f7c681b416ede2b447de4eda371ae023330783bed172e
ze8cea2a2c5b9cdf37db94dbed705689a612053153f78ad22323ce4fff35ec8b8e08826a79d2350
z1a261e7dd9b886f25cc815058bb000cab1a0d5df5aaffa158c1c2c9a1d18e1d9d860495e40b878
zfe4f61eb33969fdb887fb5a0449beecdd0b5915922c7b31d9fcbc2353f9cfa12f3d09d7123db14
za43d8ea85ad9f1742aa2d41f43f0cd8466d5b2bc8cca453b35979aba7e1b6e39cc523934a8b0e1
zca3db192b782851bcd0f062dd07443145249322cac8cfdc5aca0c019fc2ed057d3eaa7e743f6bc
z065534c45e322c481e884c8b0f4d2f36af2bf40f994783b909431ee11e15959212b7e99a6e7a28
z126fa054fd09bab1bf6501fae4a3d0142b070adf432155fd7fea8f1b0170372618021394eef698
z33bc352869cadc174416c2ead56ee553dbcc5880ad99b97b7326dc223cfc154dc0b5446e2cebd0
zdbbcd8356b79047ee3a5fcae5764e1937f740da233f50ab990628e4a46c6a34d789fa6957e3064
z2ac6081abb6667b818ac5d3714bb16cdaf48a2346a07ad1c8554d1693b9db1c9845c08564f742e
z4c4c5fc5408aed5f9f058e2b6befbe22e2472a252e208a3b1a814a121a5c44bd5ee8c8579a5e6a
z98226b67ee1df0c955cc3cad647025f4cc44b13349826d32af362befbdd6d52830265afa516066
z3a1820a0dccc57ea54ff683d3d90fd60b808e2a2fb4c3059411e6b7167949164d943bf2764e48c
z78216e072beb9d0dcca85e587e29cd547d0b42ecc58de57c6a3185c24299d90f38d126ada2f2d2
z987876c35508d78a6c424c46bdc4836d7748f7890b9b37318253ee10ef35886c765f5763a5ec8a
z2fabe5e86cc8b58a921eb6764b39addd7686c5a6680841fc89b038f465bc3c031e69991eb73802
z1367103824cbe41fe5f4c78fb634b053c36b3f81727e4c47dd15d675730efcb12bf6a3bf166d89
z4a93bdf4331559f20c293cd188560a4fcc8e7510a2879d73e3b3268bc6c147e88ef9f042d77243
z55e271247803ec33f95c8d8ba2464ae1a61c0fc1ee1c49d9afb6396cc0e5116159fdcff31bc127
z428a1272d7d769f02beda0bd775ce49e96ee8001c5325100d4d885a166f2a94ddacb1e85413a8f
z8cf2daaea5b530c32764990ebb5b0f2889610e87bcda262b9b115929b4897097858df78a1fc6a2
z27723bf7b9ec1964387a37e48f308b6d2198bd7022844a3b65094ec500e277851b36ad03450f69
ze4ce16b27f09bc2478d3a940d765fe04a26a3415bb3e3d58e2f887746d346b17b34fbce834acf4
z5c3f0e57b2d3b49c8417ca192c879ee676c0a102532a6eac1a2115292ef2d616a8e89922f903be
z3db753833fc98e1f654330b46c810f6aaaf9fcefe5f9368fe2166429469a99b6c1c0424d14746f
z6e9cf7ea1f06146b7ce9ac9c61678c4a2829dd9479debbf4f8e8cadc29473c4aaf0b5258d2a409
z3a702f412213cc4cbb746298b4b89eceab1ac787c9eb60ea4a08c72f95137b75c9915246b75d83
ze02b90ac02642b85299cd89df44205d6fc665f989af4992a0e56822177698135243f48ff5d66c4
z0f6e97fb0edf9bcb53457ce705f065c787bfff602bf9104100bc9bda013657f63954a15d42d30b
zb94901ad6720a31adfe14127a8cc8fd20553251f3f58aa58bd0cbaeed2cddc7a640ad5013693ce
z29bd87ff943d65ac41859e7eb38f02a04a311b880a1e0e3b393b14e23350c7368921d4b62a3a1d
zf0874bba9c3539ad8e0cedf31c7a568839a913825323be79252964258b8f56c6f665ff40b1ea40
z1a0905af2fdadaa6dcf0e110fb65ee75248b5bdc932a906ba7e22a01c6c1f4c21f78bf2b31ff09
z27061975472068a5540a8302adc2617960d4ec176db7eeedb577a96fb54287df8d80a82379f0df
z8a90ecc416e338e4c3e726aa45a0c485b12e13f4c2f4fe04876e0abcbdffda095ccf45fee9b7c8
zeb5db16b4aaf5add49d2fd409c030cdbb12c8e9802aa310653830410738d54f9f44e4bbba1d569
z47c88c57fee26b9fd910ac0321741490baaf93d319f6fa51fb3d3a4b326a635250eccc75c2e06f
z9ba25d731ae68f523cb33a8a44a74a56ad325b3459961ae24d9e4db1c63ddb5ea119283d0d909c
z9e13999d685213c1263470c354a1cc2c2b60b0c438cd33fa1d3f635f7b11bfd81b16f0a6979e7f
z0523f602661eebca13cdc980e01731638afb8037f0fbcb3de6860fbac0e89c1ebc672e80b3ddcf
zba96d375cd1df8b61ab184f34e7ed37f847aba3e12bbf91c8874482fe18370696c539fa6e65771
zd7c7a96ee568de3a761d1200e34bd5ba9b2c2481e5e775a657cb65505d8f0304d920fe43612bfb
zc7b2c0d8fd8ae8d7612942563cf8375b94f2646106b135f640f6035f31c5b08739a188cada53fc
za20ec076629fcbe50c62c1a5765bcb4e7ae413fed3fc35b45f423b395b448d5d12af10f059c4e0
z7abfb7f87acbb593f6e5aa87792cf1a2b60417d0ab521b11861f7e57e4129fe7ea0d200a694f08
zd593b20835dda72db0a00aafee7213ff2512e5e46b5c001823d17824604c8475ccbbcf224a1953
z43043bd065277e014a579431ffd928968adeb3abcdd5e5b9d2c410d6cf69ccda7209101eac93d8
z250321b7cb2cf2201a7ad0dcc480f334bb9094f74076d4d6e6971b6e743d6fb80bec242c335c33
z9929212ca0bd7d58f21b43a9c60d8dac22eb02548e9edd9a5b3bb142d284f9bcdcdf8f6916d672
za00b763ca35f4ed38d218cc3f6579049b4ac2f4b94c04632746f715c8f2fe895708446a660c022
z7590c220cc89879e4df71538319d7b9c437e7224bcee9b50ac7bdc1f5ffd8ebdf9e8c7f6b0095a
z725d49c8b609ccee8c1c1fd9719ff8c2dee5c96714a8593cb1b1c91d2027189ead6f92ef9b4b89
z364e79fa9d2fdf92d1285e66b0e3b9e116939662cf9dd2cfb683c37746ef8e6f847e9d01f5ab0c
z427a839fd3f9a921b4a11861e220fc638885e0a711a000e9311cfb6288a99f07f369e2438869f2
z1ccf76afdcdc7dd09bc31f257ccbc19b6fb9e834d135f5766e13b9e3de5362571f41aad5db027b
z17f37bfd173a04e1c0cc01d17937950ef9bfcffda522c303738c4f9401cc37339458852362de3f
z60261abb7058aec63bef66dc200c545d4a21e291e3ac5827a2a0066a9368edbdc74a70906159bd
ze087f26a519d0af33053676b5258fc18e21b77a133a073cdcb99b9cd0ea8cc4b83c6770280919d
zd08f5ef91f47b6a3abcb82dc755b59d33b468ac5b3a3734ca9659de65bcbc3ccb1a8881653064b
ze83dce7516f28bf802cb4a3a6d60075b69af7b85ee24e60c45e57aef421a73a25dae1cb7e87aba
zbb425e1159354531950f384d8c524b8ac21cd6fde34648b494c630f929d2d7a2ef815d4d96e546
z6adf7dbfaec749f4ab2b6c9b21da4e7a70632b696bf6def4db3c8a126b56b503c53c38ec8487bf
z30727c761345e5b8562471f3e2488f978b9fc83a72735ec19b3a52eca2541746e83554060c5042
z3d931603d66f7a30bd267d5a9c742e14ac20c0e97e7958572cfbae199337ebba319f91b310e480
z3fee5545bc4fb51aca8da37b98375e453fb052109293b0677b72c0f7c22805c82f45cc3d926626
z82f399b5fba50fffb471054bb8e1965dc1b0d76d73f5c15fae744659d0e5cc01274a76e3687408
z5a91b9dbaac4b1e2faac66f3f6748b8e6e08cf500802e215dd077db9fe246b801964ff1ad00d8a
zf5945ffcb3818bd337aebc7c307ada9e871fad2b1b24ee53677a1a22bbab09e7db42cda2dee353
z5ce3cc565bd18c5d499ab4be4d06e07b31d827b7ae3ef76fb135d5111944855ccba82a8a299b13
zb4960ab211f93b56fd06382c76693e805d413e79f260331094d310bc2bbe15854b7b85ca318caa
za8a86e7c2ac484992016dace06bf30c24dc07b989f681fd702ce0a88727550568bf03596acc4b6
z7a5d865b331abcf1dc625a2a2d9ae6a08bb818676c2a28a6781a29c8dfa6d002268b3ce5be613d
z09fb57910500dec04076c7c731f7404d1e8088e91e689709498cb724b2afdb2e36d2c44122891c
za2620eb5180a9c58253445007f17a79f11e9ac0300a25628846184dc3cc5f4acf974deee62d4cc
zb810e9fe68f6bc3783b297921d374414dc6f3b2dd28c4a5ca09dc2d974f8f6eb95c241692f6693
z9c5e3a1e7775db0e7a3d3f95f85e825d8aac1b0581001cab170b35ced3a7f42aeb9b51cb2d1ab3
z26088a80747f4136f4384ff889dc1ace886d2c8909d4bb02ec839a62d7f751cd50dd29bf1337fa
z0949de620130bab3b9a2d62478597ec67ddb4c00f44e192cda929cdfd386cc232669084ed7e4d0
zff7f56423d1583acba33b4164ecf8ec42109ec42a5c0a7d44566954e7c428f1949cb1c7c6f7883
z2280d319a12b71177cc2c19645d620c673212628da2b55be128f2258eb09649caaddebc497a92f
z7fc79bfa71a0ff8c229322def7319f769d2fbc71ac7dbb051d37957a35d0d51039e1c577212cda
zb7a4f7d98eb5434e33895bf8435a2f67e2115352dd3e358493aaf0e4aa159ef99627dc5d41aa5b
za3cad2dad381fa736e1407ad8df40301f661757ce8809f99a4995ba91fd3415ed01dffc9fc996a
zb3f938a055d580d1876e552840e173eba057f272f219bf794b78e2f547bb355f19ab7ef69d14bc
zcca200efe9e8f7286823ab36c3cf777e13891be9c602974f00d8ebf00a42bd0ac5edc0fd78f855
z44b5c67eef12f276d9a6c960c5d0e37012405efdf99487e66264b1130f0ec639bcc166c427bf46
z4ff92bc7528103f5f982c401a0c32c3c91aed73baf076ffef0297ec465da004fe05f646e9ff488
zea214ba09d9fab2279bca949231c6720d513543c6723177b601c104df8ebc62e8a6d8e26db538c
za23f3f4b7a68d4fd8ed6b4a0a23e16970a4be4ab7bea96ed8590e918d4affcc1570a1655271fa7
zb34d1d8aaa0d9b566b0901754674d95047db2b17641932749b00632bdb05df7c4ccc4254bdb433
za6ad649d4d87f2dc6a9e5af680f6b15b53f37a8bb63c5e874e71029cc4cd0881028edadf2523a3
z3feed89ae6d4cf3210927d323210ad29b56905dd24e2712e5d9111dada3ad3efd4160ca4d279ea
zf158764accf0b180280d34090ef392ca1eb1c63dcdf31afcfecf53611bce006ea3ecf95917c9b7
zdbf831d133553fcc8fa710aa85662c2333fa526124216cd3d4016c25c87280ab78a3d95bf494ce
za713ea6ca025aab54de49e0c79c86d3c4bc3de8db763286699ab60f1718f28d043ae61c5afaff0
zad926c7c83ae51b8a72ce4ce0a0fd5bfcecfc1e557006f61439d139169c3975677189dfa72a075
z293866e8f928eb20584f28ae4b3600318eeaf0d79366d3e4498b32a0f5da195e28dbc5d87b4f06
z1a52cbe063fee1a06ff6eb4fd913561dbd462456ddd2e4dd09a8907e9049ae8aea188aeba13ba0
z81ad797d064ce3f450136a82016a0e7aded28747f8c7443ca52e6e921386838f45d1524fefe0dd
z6627e43be6d6f57210ac1cb4f7f05d7615195074830f846278b62254c1bb4ee4ba90288e9d747e
z12c8fed9970d903c69d66089c2c4f3cd99909e9ff0da1126149dbf89e1c74178042e0d9242ecc0
zc5964c946342fbb1ab4bfc7006c3f86a46e3cd267abb157d74125a548feae762befa3862f8b4dc
z6a2a683a17ad901387944ec3aa4c8c88531b547ac2fd202e1d683e1f055cd683bd22193799bcd7
z87e350786c7645ab4504ce99e047e851ec8d7e7efbada9846178610bb6711db45ef432d53fc214
zbac714c1fdca2ebbac1520a3824d554824e07351199a66a264c6ca6c648c41c86ec577c1bd25ff
z33db3f71804cd56417c82aa4dd4bab8e548e31ff730fa73ee1772b4f0945cf04bf4d5b64bfb46d
ze45ecd41288179c867d8e0e4574d22fb5531f33df48591eb9b378ed8eac1e5f73a5e49038f8a7b
z1ff76e705880d382049d68441db02b81be8a985c603b6597dd843869f258a952e4fdc05df8bf28
z529b397781990e563a84da22abf5a8e845ad515eb958edb26832d043cc7cb0cb6a9dd1192d04a7
z6d71acd60f6081a6897c869465b90dfbf3390818dbcbdc2a02a326e85e87a02a5f26a81cd72ff5
zd6c0cc65eb6580519adfff2bb5853eb019754379ed5104385d5ea259c99ae3668418ae5435434c
zc7e05331e9a559ccc04355536a44e4cc928849af82cb5ecb4cca1c9be74fd45dc8bc0a66e31b86
z1b247b84caed029d1dd4604cc2b2debb274b074536d62a519263f3ef46d56c6a1138ac21571f10
ze4681bf18ae9a588c71db3b4e0639165b95177e666c140a3a00fa721f318d804e6239d45d85b4b
zb070b9baf02241e4e0c6bb946d33d603bf19eed6fc10870c891d4fb013b8b59640b33ae0f83c1a
zb8a1a3bf08b2ea5ac3609f3555b906fad9377c83af8e41b6f2cfd9f9e4c229423c91de97f996b3
z47e3e233f42ffb05b98425d03075a82a160619aa3af650390eebdfb51e237103b8b0ce44da20cd
z4346fe6fba18c367e1ab465eaca8a30a5e01b7740933c8c10e53ba32dd717f193efbccd34c6736
zc90a8203201c550f777e7d340342defe0e1690b189c241b923a3a78c37d41a8359c69d80a66a76
ze76c4d2f6c7d676dbca2b8708c755c654b80ea05554e12679ce233be69c739da94a06649a033fd
z9ade6f7d89c6c5b2cb6e5c30dfae94f3b28ffa4c1c36e3f8fdb641bf88c0b117b6eb241f8d5cc2
z8cd7375b8c86b5e7dfd93bad4cd724ebf94a4a2a566526d37c258ff547a1b6e1b49081269b6123
z77adeacb6cef3cd7fccf6634203df01a755d02822143088541baf3df6746360c3875554405bddd
z2fc63b368b9368df8f2e750914d08d01a56e31d4cccb59ad47b3d62b1d5f944d31d72ad277d3c7
z6c1312a98cb6971de9ec46fe9a0d724299ec313909912ccb1a377d1d073bcb88a9979d1ca15047
z0d5981572abc1e8436ab97aa95c7a4228838330c85c381b311e5b556dbd2ec52cbae1eb0f1f777
z4e0dd50f411515bb2b476d4795a823e3920acbddc2048e897702ba2c8942d64e23d743ac342767
zfcec301ae87fa88608375142d621d7f13a2e352d0faf3082fa1e8d3fb7b1ee234700c949a1fe76
z587a0e46d0e91f63aada753b321b148f1c3dcb890a823fa20e9a5cf6dc6369605da5b023b73c32
z9eb12c5ca69c5109cf4d626fd7355fdc9fc2135fb26a54622f63a4fbb736999c11b537cb32eab3
z9f91462568885f405cd59a919f6987d1be1055afad95e85f16c7b7aa4472a5eb819fd059f8e835
z3ffb0e6b2a239ed6a5c11e2c47e00a5af64360e7329d9ffd83fa93e91951545252d7715d94ab42
z265a148f1f9e430f8b42cc9f5277fa9caa2fe0c1efbc8b5ae18668930e7227c9d13f5b00116b3d
z601c386d50c6aa36a89a47f50edaf7db1b810f96b907fe71fe0ce64f32bd981594b4bb80c8883e
zcee1db7e04eb0283df79333fba28daad433f60db41c05e949fd91dfdcd338c0acf0a587f2ddb5b
zdde6ea910427aed03a05ddc35ac3456e40e1bf9549c36256c43d8941bab9dc2ce22552e1d4ed27
z8419ec7688e7e192bb970c55c87369cc119c078ea01e39ae379a6682e13aa15cb15986e2091fa8
zbdf8c5c1b72244102794e139fbc96461870ea4d3ac9f392e6c160f6dad6d2cf68c3a80796d161a
zab7ca6c8ce6d5b61a4b467cda27b5e7e75e61e1d38b58f3eaed9ed11fcf4c1d9ad47980f17750a
z1427788a7827f3c6c8466409abd28b1467cc40a05b49a53b2abba6fe28ade30e3bf1cc71ab69c2
z421c35770ff11b6918fcc8c769b6505dcab998ea3aaff2a5786f4b1ea61095ca2cd25a74338fb2
z04a0d3c30488dfcec5c5e9a0b8763f7eace91b08203639c8fc8e6fadddff1067b8bd98b98afd8a
zdb51e828cf3da360136b5c26281a3e3e0b7e0fc2c0d0bd840fb4377d9a52ac107f4a42c8af2099
zc1e506ec893c1ef934f44dd699a9765d3ed741065df1f03bdf2d5f02582430b76086c2012a9ba3
z4339d973e420685bc340cf51c8e550e50bdfa0b530ccbfaac664d55ef607422ada37b89e8de9ce
z456fcb19c523ca659ac912cf8a8d75eb6087ffd9067d25c9da6ab0e60ef348f5bc863899d320df
zad0f17c1e4e2cbabebbbfe04456bdb05b2ad6ffd50596df457f0ed9133f7f3003286d8cc4ab068
zf8d61468987e183e24359ab4e8be5d7f8db86132c18b59a3ea22ea5e0edcfb74a3b48264c1c4d9
z5e831dce58fe6c622861cf98846f124bc2331e2673d5fb732d190b033f1b2166434c8ee504f1b5
zb6d36c9f8b48bd1a4984d9401dfd7bca254c485e0417a29f65ee9e3622f7edecfd0cd51160506f
za8df00eafd29e905bea6c0475137b60cd6e3faf93f92dfb755852b624472a37cbaf126bc1ae07b
z17a16ac62be07c7885121295a505ccc04ed1e062d6554ada22a34f6cc63908e8609c954ca26806
z49b401ea0ddc6ce6e70e8789e1e8d29cbd5da75417df7db08ae00d0f6904993237148d4834ffb7
zcd8cb9a47c9688556de32e8442c7917585936bef91b3a26fa9611ea36a6d45fcd88e548d1d7805
z23a1eeaf4d2bd4a1137c6b6effd8807b4e0d4cabd334dfff5f3141d5f9aceba1881b5101f3e604
zb2df0e3013b2af1bf8fad3856b65fc18e06f71f9ceb68e43098f94a2ddb8b204902c3b953dc841
za895295750f6cbe8af8a24ce6ec51888cbea635122c05b51c7cae0455e567c276b220b6c47f803
ze611657214e3087638ab0e55c56718451bd9a1a0cb6eeff9631defdf2217eed6eacdc8ba0edf00
z5b7df031a4be55380db649c221ac898608b86b05cc13036696eec9e12bb7b3c1f90b0077fe3ce2
z1b50a03054fb5c12ada6c41df90d42a360c0cbfd1564a59b5168a5ca003c09defc26771f088576
z8423c91f1284e5647f7e15d984011b336a861ef2ea3e4961fd27574668ee1e441c639c180ef117
zeacc11d976f99b40d415d8c9a6605827b8925388f9c8f809c09d53cd35e7ce158d35233809d55b
z353d4d012a03db0d8afef0853a578e2191a49b7947dee3cfe02ed250ba7ba9157715b3ecc4b35e
zb40eded8db5db23c227d4f0cfc8d129a85a275b25cc1d3c8f2983f675c759cb85a7f17ad76b517
z9c6a5cb9a490be5e1ba46dbdf66d5f48c16c157706b347c344ac30cb58ae1aa72e5104fbb28864
z3295060c8a4b93dc26ccf8bbd80dcd4282d56d96a3f998593c4b54d3b5269605bff3a976001f1e
z566686264429e459a59dae5a110bf0b78dcf422a44cca455f42890b0b55e541194417be8599747
z39ba4c59eeb204dac05532e90b49d4d0f93ca37ab6972991324a9b628eb9ee39687be272b2c16d
z61e5b06cc0d5f7ff5835205e9a4da5dc6000ff41c856f23dc53be43183bc4b324bedb30373020c
z47e574b828ce9274f8b7c61b0508db32fa6d16f32ff52743513e4a8cb53edc0709919c3c0fc120
zad7238ec212922d7dc6f91af2c9e2a097096fdf9a9be7e1d39454c19dd6160666388c5f91ff4d9
z7b454980810e8c22268377a57cb5135f8e86673b5e99ac5c1edf57a44a2475845f12c87c12f754
zd1778d0d949a842cffd9256a313f3ef60645366e4e31cb5b1a70de643da94427619b7e92458ef5
z7ae2d64071b5f338a3b7cf03d2124e2acf5bd5ed9635c257c6fb22cb92e3e5db1fe3bd04cb64ce
z11a19ae33c3bc5fe55f77bdf646d9ddaeea981ce885fbc98e1ca4a398b5b6134d417c124494dc7
z44ab429ffdfad2c6c29f1d358950c5bb2fc73ae556132bd0a799c5d9d2f76984d813e1cc68c19a
z225c10a7f705626fad8db3f0026e951bf3a7d85e1218e474fe1949b8a039601e11aa34feae1334
z22fc5e3a42c223bf24e69f81424beed842b51e3383ed9650a397e217c60dc518bcbfccb079c1c4
zf2d608a94c7c34e2b14e8473cb9f066d0add1d90458e36211e429bea350cb7a51ef175e44cce60
z7756d7556014fc00e503f9b765cefce7578a58e9eb903ab4a145baa79a01c8bb97c886b6559444
zb867cdc2c52d2da608ec92bef1b202789fe23b8060cb9b927d49c32f2d8c0abc09ff0561fc8bbf
z26d6a2fc0153f18da787c06ac1c7cb67bd2dcdcc46004bf5f1f23726e5f1d55c889464af2d5e06
za60b1b5c5deb0fb93e0b8bb94b2c4efa956bc7a2355504aac88095d8bab5974d8f3f42580e0e5e
zf34245e3b2efae952f8bcbb0fb85b20d6ef6c9109da3bd6077185bd170ddb35eaf05bfa1454926
zdd888196cf40fbe2f6e86119d57207cc6b59da24830c92c235c31c2ebacd93cfb71184e3937b5e
z725f54adf810220aab7da5f4176d2b0bfc49bb3996e3a4f91d2d41bb3d9cd0c31a0eaf8f4e2b00
z38cde02d20004bd87e3f99afc0212644c1a46f9fc2168af8a39b5b9f0a46fc16c1ab3e037997a4
zffcad1ffa26a04a0175b9784e866811be3699a1321ad666bfea18ddde2ca8f246a81012846e269
zf38dc5ca1adf3497c6dbae8b78ed09ddfb095450b9229a1c96b8357ccc0041b2c4ccd5967139cb
z77ff73ed6b7d6d7e673d436d0503dfbfd7f3331d67b8e2dd95570e5c7913deb423dc123e9d7b2a
zd98df1ee9c018a184ff7120ea5d5a3d371b34c3c082316f1f85df52189c56a2d921583ea82008c
zfe0b15372e49881c149881a73c0ccaf6457ce1f9df660edd730f6bac5f642ca9ad18522b0c67e2
zf5c8fd5698e2f9c5b7e3f334f93a422430dca66009da6cb646009fd0695e2be5b74a1b14492827
z76a5fa7fe1590efabf669e86dfc611ad82c2562a04448f31db473c233ff9ec6c42f10a641e4fbc
z83a466d32b3f7b8876f8749c232b7cf7a6f43d8a64798e4ac8fa11d9245b5adb340fa7406a54e7
z4ce068edbe1a4c635e55c73a1931e73c41ab2546819ed90d4edc9093fb7d0b33acf1f867940e6e
z39d335e62a767973497e1b19e3d5c4cfe91353ac6b0f75e65cb0f91c9f2cbbd6094e9da04aa530
zdc8e819aaa114857834e6a24c83f4fabe4586f8bd0321551d6205c8b290b10a0d34cca2f94a678
z61da41822c6d7634e54b3672bbb3091aad8a0523461b32973ed063aacc41123001680c8d751198
z585bb72f0dbba3954d7a3722388a7b737458d39fd2281639585aefe826dca522a5035b0d6e553c
zd1410e659fcf84cb29ccb628f7dcb74b88b4a00f2d088aa53c29daa625665d20446cf7caf77b46
zcb42428919fc8a17be71c624e253b2965740b4ca1944eb34c8ef8131b0246bf5d34b93e1c4eabd
z023440a69bc52bd00ad44e882a6ec068eb0714f5c56c0346302953cdba69e70e457377bef1062a
ze13c40cc59de5d31697b717c0f2f416e45948c0e486c7a563b246047bb85bce415d585c623b269
zb4326c91abe3ce7c6f1096956822990bb837998634d7a1f8d84172e0c525c9ea148c54cf54e6cd
z98f37403c1625732d2cc2a52b94b3244137e84c336d39f3c64c7f3961a3dfb601882838be56a3b
z363b6a846fbf40b46caf9d40c873a205861c5613da5a3ed132daac305a2a245d67b62df987b779
z253448c753f3532f51d6022655b7328a7984d83b2e3bf9b433725a3b5cbffbd1374c62d31ad162
zeb6115b03753d6b29cdff313220cd075f8e3b56afe81ef295f6f3f9fcf09e128eba9ed18f1f47c
z58c4bb2d0d32b691df1ac25c402bd9bdc5c13cbfbd5739ae775dff4fdf9ed630dfa7f86dc26ba4
zf15834acb05eb7a6d106660e09a7b3595df588968aedeb5119b72514ea17bc1a3b968ab5e3e774
ze280b65ba1d2a14cb4e92e27a8633a44f742a1adf2ccd9ba00e1e0daf5b84ca23a16a57957bd84
zf39fcb37016f0e5889c699f8cc2bcbf04d74f75feabc927e11e7a162047ce2a4bb9f6aca8f7b97
z59cdb0f82f4640bd9ad94715882c21b168b35e47599ec0ab3a1f9e032a49f5a0d77f38be24e66f
zccc8e52d10f8c5b08f1545f1bd577303ca6d88a0083731bb19bd1e9fd1c7e57b2faf3f1c35c41a
zb8569448575182679bd4828ea8c4df872fefc3b96f0dd2cf9ffe4cc3b1b72d14962b155a2a729b
z1ff784527620a9756c0e6b8ee6dbdfa0311c66cca4eba2b59c900d03ca0fe2c4603dee3944d389
z4d756c3793e4fa59b58900d6af7b718b939bbae88ffe0f7a3d4c0cbe46486e0106efeefb5bfbfe
z471a5f2e3eca894aef57237e369ee973f96c8fda7965c9b84f83fc6d5bbadb8fc21c0ea914daa1
z2fe678b5ab180baa3d81f5b5ef4923ed04a83505cc30f6238d0b5df9552eaa9986a3c495d3c737
z0a957a3603282079bad4859c210d27525e5fec84de26e2152be7fefb73fd25282b2e4632f6e0a8
ze8de037f7c80b81aa89b0994ba19fa513c7b73ddd2c5fbd1131cbc911d8599ce4d18cbdff7cbe8
z0e64c076a73dfa21db478ccfa9065a3a6894ccc7e25bb230eba9bcf1a474f2fcfb2d68a1c5f232
z3a01651b53e71d19c49e7ebf1dc7898a70388a01100af4401bb66c180deb55fa3527196841e161
z41205c4490400cfc9ac5d2f1d1f1867bbc8610f43960cb6604db800ad9801f0cef48f29502cf7d
z63a557ceee968252ec7dd5b31596351c94e2a1bf14b71fa7b7b244b30b200b0aa5dc2a249c77c6
zec66f6e7bf913539f3617c2d9b7e9bcaa77d02775a88f373b10c248502d1fdcc19a494efde16d4
z753a956adf2257828e1abef733df19ad1dda06133958e557843dd6021e9fc9c6f37612e32f3f0c
z3e3bd42d8a2eedf973e8baa2e0e75e23034bbf1131e1e1aa4f03a904eaf62c78b699548093a9b2
z56c96aa4fc2271a3e13f4be9f434f62d3df9722a15b46e09758518ea8f34755f10ad4ad4af1146
zf5104b864c14a8cd4d059aa5d1fa008d9bef4026ee28768b0fa9d49635445d86490d975dcf940c
z7cf6ede584b677330d8b10c1c092173a53aa7a42caed832c67eeb92429d99fe0ca842e03861f3b
z51be079fd3080c8011b88c596d43ba001e495a5d2bb6a622c55552fe0b60133c9ae59bfbc1476a
zb7da80c140967f6794691afe3da5fa9f8ec05d15ea647420b32e0199355cef58046840b1b2edfd
zf08403c4ef43ca333584bdba972b45e339006daacf13cf31499befb92061be18a67b4e0db9db8a
z067611adb91c4fd37489b2aaac684b447f9be956e170045b6490a63225fb49f8155967696992bb
z63ff1f3296905febd42b1c70a4e33174af7c50b1d7a92cfb93951808910d45cc2e8d82a13c1c3c
zc32af2ed4a02443d16000e5e6e61978c1ad6f9225b2b4b947884161ed60151b7f1f0e6a7f83494
z3b10abc9e43336ec306b93b41bea827312a0d2558a64cf2c3dc9d378d616f95a868849b1f27712
z37a4628644dd2725bb758d59e58dde43f7080cee6dcc2255d7382c07163a18a6e15abaf553c3cc
zdfc19ac813223865d95121e55f75e787ad91d0d0b55301fa102605822f1ce451f52be806c0e67b
z5c3997796956b3b7983ff20f4d227a2e2823ae8ab006f222423ac45fe6c688a2e44b9e1d74d678
z42b5151891ead0b2d1ddfd24a4e9cd21b09d767f96494f44897034cc3a9445e7866192e4511c87
ze026ca37108aa8fed6555998a397e79998b40f03372e2634d448acfe2730eb40c6cc1e954121fb
z216a094e77e3389ac19a33a20eac7ca878b2a46726eb253a3394db32fb009cc8d0ea9c36111bf5
ze9a57d6df265258c9e67e6a722a7074e583e17054300bf501b8d99679c4f4a496832774be510e4
z0015622b94ded6db724b3d1ce93780ba028f35ea3101962ab6a18e0986e9d712df8b1ad77425f1
z8a0ea1cdc505a86f6c600fdde3ff71b3651fe8bbba4b8f4837cbc5f545cbb137dfa2a8b1c0a6c8
z4c90dbca177d93714752a0f0e9f6c6564498e1f4b097636aacbacf9aaf6d576d87b2798509a196
z487a4b22c67bcbda447a355d610c040be49c17be83fe4cdd265ac7aca5ce0d08446c7fcefbf1cd
z8167d373577cab0b7d0d1bf2f5b36829ee7ed7a373bf73e48e83e0a5b894e80e2d0dc0940e4492
z3a94530188bdf7f9146d051932a437a470ef8f94a9cf1e472282105b3bc18b883ced012d5a601c
z506400a54ada7333f0f83d0b69c1d8490ad141b2b631307a5229c29c74e4e0c5bcca43cb8962f1
za56de2ebcfe3992a369b8995a8caee1883ac28d1255b5343114ba2d061b3ab3a474ce751800fef
zdfd7b68f4bddf40f35b761940d1b1ab64a6f642d60135b55df127f8fba5e84b4e6998fed940869
zef34f0d0a2401843c204770321624e3770842e538252cc3bfe9c6383139c982e01e909f6d0c64f
z6de94524425e3de4b4d1f47534aa0aab6a5d051d16bebe2ee7bd202469b55d81ad94a5e88f8d83
z9962a8399f3603e1a0e4df936135882e81315c9f46042a57262c0973beec42f1b2a85024ae737f
z4051183abedf3c5fc5d072fae2aab61677a7240ca66405a78aaed66267465f911e552d55f54293
z8f0b76921011a606a234c939be0d31b6108188bde62d994d3f04a3a452a9477613f2c60ca94503
z14e40fbfae75600fd5df7a64d7a42b5aa095fc409987f3a48502cdc03ed1f9200b3857ae30da64
z584773274eff2759ca76033cb273d25fc11f13a8805d84b33a5c17665e8fb37772d78370d81704
zb78bfa1d2b09beeecf098377f35ee42f3cd5ecc754fe9f682ea815809703a5f111f76d1855fd7d
z02e42a87582868b72c76d722b5e274f9e1ca63a25aa5d04478c04bec65368698f15fbe68bf159e
zc61016fcaf2abcad498db7fb388a45a01ef4b72d64ea6ab8f7e76ccacc4d506e8cbc6a7b0b46ba
zd62aa7229bff4521d9ce70c56aa5577532ac77fa17a98b631a9b9a7f004934293885590402e98f
z11a48d7766a0f32151cd477378be05be09d60b200657df37c59094a8070d4af1997e8342896257
za067abcb385dd79e298306bb98bcf7f208f55cb670cfcb88bddfa733995525a893495c9186f6e0
z5c9141b9a5ae25c6a1d2c88020c053559a9ea802480bfe05b89ce097082ea66baeea367449a8e0
z246def4001435b275442619ccd1f0680aa1a221dd1c96ecf1e183f2f61a8c49a46b0daf2ce88b5
z4d6fd9b258fde6c9c9d47ba83601ec8770cfd6b221973b937ca329b6d99df0f215235fc4be84e1
zac5ed66b1a73888c42ae52a4c05e9710d00519d7b59540e440e44f1c0df200c335e5290c359324
z81953db93bb976280abead605b7b52b55c829e5bd7c387925c20d782434d0cdbf900ea67f375a4
zd4a5b92e4e93fa7a511a2575fc810a67d25d6e193a1bf6ba4864b70bd51a112745be5b7f99bbee
z6fde87436d82e77c14119600dba0be8c2bf0d7f83e64dac75c668d719b2744abda9208dcac30a3
z0f90ec58504029c95b53faece37d7089a3054b1eb4e65820441478a0b5305e172b1c0fd3667f83
zeeef3da8652c5f575d643bc5492e38c81f25861a96b6cdd2e10458b19fe51d475b2189c840a691
zcfe86f59019fe761ea9c01f3ab60ea07f637706553687cff22a4ef69005396b07dd86efd9d57be
zb873bd912fd190d536d9a83f7c664c36b25ce2be148b3771e41575c2ea0332d4fd5e32c6c0193a
z89e335a5d7246778e1e92527b7a1d170ead07ad2eba91bf7c06d15a97669fd3120140196f41b2b
zbf3fe697966343ae71d707facdb90bf7b677078399cea52be2ea14b408bec4e5ca3f37320a21a9
zb26ef2f0fc4e747c1a1e483637461a4aefaaa94c13e7b67f98f284642aae50c47a1ad2edf55641
zea87045f73a602f6493b8cb0ce859e6f8a6a795d2631604dc927ec5556354fb2495fe70c8a6c55
z3730e82dc81a1eaea403309e288ec8fb804ff337197d684c861a93f339cc27dc1cc4da8e1d20f1
z8d39647b8c93a8c3cb8edec889eceb9b2e74332ac68e6f1ddae58ff9e1be7866b86562f81ab142
zf2621f2015b7f73834e5679d2a3f298fb22b8dba41153c3625c4244d2a0ac9d24582a7a5f460c7
z1b0e561da910ee4014fb3331c777d59b98b3e3d5aeee1c502ef96126bf2904aee4cf756e705683
zace53f536144c96bf325dbef727ca67359da4ac29ef7b061312676604016ec7fc40a715c582f43
z4126e05d8618115731d1d6ebbc0d8580d2ced1b7747239a35d7c33bd147587130785139d2d1e7b
z5c4fd1b1d869b89ca6b788e90c4cd459e9c9cb5034e14cbc9115618d2e782b8e353f64071fd596
z433234f9aeb29aa743474a64425afc3a2d200511131f1adb05e971826d59d8638610027c5b4771
z38df5a5760f34cb3fe42270749d96079398ac5c93ba697c96708f093918d0f065e232a50a3d582
z47d394f3dc54c0df123d3a9c30d1eab089e9d6d812890c647df111adfc29137c3d1297608ddb25
zc979ad0253bf48a15abac8ab3a4cb3e0e0435308f49c9fd12b7308d5a10a6a6400561bc0d01ee0
z47aee51c39ce28f4fcb74f03cb269df06890bb7473834c075e089276665e26abc1cbe6f2396c15
z20e0ce9a97b6589d4ae11323b9bcb6d683110f5dd60eee6bf621255ca8f75cc51ce8f75af94467
z85949de9708c3fcfb3b7ba790932196b3cc9f657367ebd2d07aec972c8ee6568bc7dc3cb51b9ad
z5327ee2ebbd2e290043ac7bdda9f3db179dfaa97194ce5c1e2aadbdc15eeaed0675a705f7d057b
zafbee975da115ae7ff52fdcdb509756969b82efb1b8404b778bdc9a824f5e31aaf7ff2d5b7fa2e
z942b9b53168ac31bde0eb04c06a562cd3aaeabc11f723eff471d9912cd2909b8b3ccc36d50072d
z2635cbca16f988cf94c404fbde013ce6fb42c4e3e25c1e191733be14a8d0f9649a7a6467617847
zc9873ebf221cbb98e27faddbd8e99f3c2dc9b04b07d6f1631cccecc41733935160b5c91dd46397
z7f89d427f5bf8da1877f07b27f7bf2d333edc9cdb1223facbb74041006227cfe27f23d7615efa4
z69bed0095f95f1bad439d444c22af1f3ef485be30aa9fefad220cd9785feffae489e74c8fd288c
z922cddb819eb4f38d4f573ebd0b49cc61aa499c7db03768d7ceab772984a7f1a03729289eac721
zb192cf365a03bd1c8d68b0088f4354f81810c890533afb3426f4367fbd5c094d1fa56df3014a81
zc8ecb32e00c4800e7270fbea3c2f4ef6c039fcbd99c2b21be3b57880f981b8faa23dcf817b88b4
z644b3e3a3c62310a0153d99d461a7432d62bbad0861d5c2c34b878f5040a20a515373d02a2e10d
ze2ee886cb09cfbb187b781929fffae347de1a737fac1c84c772317426f4f52d12ec832651b6b12
z248599a08ec01df97b93338a99464602b593ab6322ab40885b3c436377048f03b6f8ed3d7276dc
z2dbfc6821fc29d4e37b7113540b54c9f6d386574db944e393ee8d5097204daca54e9990430950b
z7d52da79e88640575cf7d6f768e835d31330e4b00274c5eb8dfd5cfef34f40670c23bbc7b69b6a
z40a9b4d184c3a7b0f7156230c070dd5622b79538c9a5b4b4c3f0eb64f23768e05c7c07d347b746
z3ea436eac2e391cdd0a28a0d58a88d6f578c834036b4b83ab69899b50cbdcae4a66940063e88cd
z68ab759f1519781ee3c871d21e92b4b2b43a8b58d7d9161e507a03ed732de45203abb4cc7ee43d
z00c38011dca38407500d4bbaf570688b1b39027edac19de2553a9d573950c61449b5ab357cbc6b
z395bf16791564afc026a5d90f668147d1dd33570f99274e9334c6a76fab0805aa1ad33301729f2
z0844fcce34fda59834412a0c435ad77c540f0aaaa71ca82dc7a3353a6226e89ac2ffafaaaeaad1
zece08cadb3f16163ab712ffcdea1f5a4d5ad5b53cbd18c704986cfcefbc79c4c13293164e39d15
zbfc961d80efb537a345e009b4fbfc5019021472544b2dc971e197506d258babe57d3be6e5ac98b
z568c5f1de3ee35b96098dd4e8188c8062519a7fb355979a2bf36440a64a79bf25419c30b3d8afa
z67abcf351097a46a49801c2f3689242586f9d8532e7a3a9d0aa5a040ea53e7223a5035dfdd1246
z4104f715b9dfbae4bf742ae30d3a62a6d99d89ff3318d4deb6c5ddc84f6f65bc63d856ffb911be
ze0805617a316193388f2346e45356d05ab7fc6473a53381eec5dae710faff184e23cad840f0e2e
zeda39750f2ff1557e73d6ce468dbbefb47d6c067011ac27b48269c301aa690f3dcd7249f991078
z5a69523c48ef5bc5d4fe868aef3dfceee54b0120d23943de40ecc11fc36e1771701b55828dfb6e
zf1a10d5e0ba50a96414e37c7008bc7897801c42293ab99f53fd1d2729c2b71ca2e9e7618dc3744
z931e31d6494d2b71e906b16b71a81d3ea5eab3dbec51c6f89acd7035a9a6145d672325ae877a83
zf5fa2040467dcaa9d418503c1a1b9877438d661da5a7be54bf997b4d5f8763049f11e4af59f6d3
z177ce1abad537e8eda614615267355899df37b94bdd629bb72ce6e1b82411a8e1f6736a85f846e
zcc317f04c1476e22c6101775f83a134feb1c594af86792a06964fad372d45d45f9d9f61f16e258
z2925777571652148315308faebd38a859e468d904a5860eeb38bb404d920bcfbe6ad2cf7e67205
z5b19d4eb56c6718e9bcfd0115eb176557674b254f5d8eaed62d30d3983a090e1f2375f5d31a32a
z320d8fcbca8e2395ced1d11065e178ba2560a1b21bf684742ad1f18d901a7c5a56f7ec67c74faa
z1f20340c58d6128b788ef86b3f423c181809c9d1b95e9e24df86d3622edab8237d768426d72762
z3bab0c233b50b8dbcad3acd47cef68fa7f9e88f26d575912fb2a2fa2e8f1461f5e73f113b2a30f
zfc30fa3d560026e506d6366e8242585e6272816f4b857f86ab45ca36f1478f671fe5d026d424ab
z199901eb28a385c887ed27d4c87b08f3fbf2628eea6eacf0cb5b0ff6c1d36e364001821c93fa31
zcd961d0debdf3dc089002398c7b58afc7d7d130f2b99b195e5152002291f830f67d145a7ffdcf3
z463842a3e51225eec50409efdbf2ce4d69bdd09ad71fab172264b695d39ec0c76dc8718baedfcd
zd37bc8857af84755db2371eadc9ff0017a2dc571e8649f60aaf97fd5453b79f36509e0f5c8be86
z6b8921b605f4dfd7fbd733899d6e3fd671b46e535d57206c3bffd9ae27865cb0110fe31c5f5e84
z211925838e8bec619e396cf0da0af70c3708070a587c2c31648e3c4c6203b653435ce7002d1db1
zcae824db1beeff5d524eede687e81eb972ccf6eaa9819c04036fb6e3fe90e5d4043a31c93caacb
zbf6932f968d30e185ad4d470e010e3b58538d536ce3927d30d6c429347d61c93efa45b2cf4e3f6
z4a1f9bae66647aabfe6384ddd46d783271d6d765fd9d82ad1a9b91e0821cd1dec6c80020f333a0
zc04d07d5848c3bde49c7058be0b01244fe2f0ccee20b9f0c19727f4789ed1b26fd041887700eb4
z135713e5630749af8671a3968f460423a0986a206950400769a6ff9c773fb62bb8f17aa860aa6c
z3bfd32aa08b98b9e5b089ea36b22e62238589c23724f2111defc5278ebccccb6e40be3ce849780
z2543abc0e6435bbd11cc4075233dc2f017b1a2b40507bb2ea01fb4872c2193701f6a75183d00e9
z0ac9557a05f22789dc6a379e746a007ae4008b8361b8d926d9b394d245345aee423d56fd861f69
z9016ac8a39ccf909897954e12ab1afabbf720daf709e8777b67338ab9ff3b0362c7808a77a79f2
zd722cbf05e066e69f2e4fc6bab095d702616121f07cce000ce9eb468e2fd3bcc13b290b6e295b5
zc1e1e6afb084a952e291e63187de0435bee6060eb58a49c201b59d4cb054902c6c8e02d8c0e42a
zf4d735a3c144f621a7c49d2921d4616864761789195202153c5a5d10d8386ea7edbeb6afd23088
za057674139148fdcc4f8e12e637afb280b78c2cf165afa4d50ca32ead709fb7837aa1486729f08
z4d79237e8127edc12ba54022c7ffce0eaccc90af639677708d0e16a05f5994d13e80a0e1d554d7
z14de6c296948390e3a3a3823d2c945ca9402347bf2d08e70e116d44891033e5bf59d1990fc5453
z269c81d00a3bedf882f72007aaed0093bca0fff1aaba3feb5c02a45df5ee6d0c97d0535449d0ca
zbf1929fb120e83021f934a71cee2af82f5b895460efd39775cc53ed984e2311f7612913e3e9535
z3c560d0e18abad4dc46e38cf0d40b8acc9d6c690819cd5b82d7f4fbda9968b19be759164cfc6bc
z4eb9a322477e64d7de1e1decdf7b2a82989dbca1632ec76a998ad3fec7a3f31f515c13db17e411
zfffc5979732e8ce36bcea51997f1b6d7196e664bc49031d3f9fb94b3313d86f02abb27ceaede8b
zf89ada4e8feba6b74038f97d32b1a9d3754bb5ccc0789afadb825442d6bb9d9f98c54ef13b80e9
ze9c80e718b968df758c1bb5a28e7c32fe272f306d9220a4d5ab563c7ce98b6ec19036356b728c8
z541c067e4ce5e6e2338fb9f33a67ae45c0891eeb5a0abd9d6449a3151c6b6907570c889e05ff31
zac63a2b9a45735d10239e818684dd408ac251e056d42e830dc67c0e0a9fcbde8378ad905d6b6f4
z0dca793cf4f6a431c977d3a4f1e6ac7694ba1f03eb38441c31ed6c570f50616e0950448d045343
za1345ab781386a1fc7b0353cc3d0be6be75565953e9f919306fccd1e0b72dbf671c89f831ce6f7
zffcdbb2c90f676397ea5e9e3538476ae2b20f83a8d884fe6b79b9a8c607ab8fcee6a07f891b191
z5772b923df80bd3262bf28e98089bf68825a03089cf954fb0bfb1b1743b76fbd09e339516f6c0f
z17cf889339139ed9a5329733349d73d21cf9ed4b8880f9cd155035777c0401c83982802a8f1440
z0ed8fff6f1191dfecc5f96b211012b1a866517aac91350b2f4542e9be6acb938472a792183f8d5
z9b3008ae34fae55c23668026f42d673306ddaa3e1fcab6b24f7eed2eab4810805b019d78ec0758
z29c4a54711efd3740e8935bfbe66dc6af1d7238b92cf7459432843eb30b5f6b7a327bacba89b6b
z062c5ba561dc32ff3a9b2f6902b39a12a51a8d4181bfa0dc6e589e164b1849031356d9c9a7db22
zde9fdd3e4a68c97cece543185422370d9693897078ff225cd25d0107b5b7054269622efa39bc06
zc5e11a827337a0585242da2d0cd43ac722486ca7eab13ac0e816c198b1250568c8d74f95ecce2f
z736789d9d7d498c4265b2e3626a9b79f9116950ef8989c6ff02ed4de0e45eef961bde8c3a802fc
z6a2cc88f711ffcc49db191923ba07f856e9ad6f2d31adaee333cc124f15fddcb9df10002eedce3
z993c494e5adadd68e937d3ac2e848bda076d3a1552b379336eb3a041a8481323a8191e7d043914
zbc5272e3cfbfa869960a35fe47b68db2f30386cf8fea8267bdb0249fd6cb7b2343283f9e56d180
z18092b58cbd00f9ff474bf0996c6a71c38cf5d9b063a3d5ebb2f45f6821ed27aca5043d9af415b
za9997789f52109064e04b40832b3c1ea7df8389abaec9c3c719c0ec257d5916d6b16afea066480
zda5ef7a82b283d65057eb9b6ec622dbd42b5c91a6f87a9164fcc6ba15ff7128a06904468ea7a04
z0d93c6b14936d9ea8327107274c8baaab8e6a2243e09065f5d405b967aeef7db2c3bbcf7473615
za74d5ff7d37512939d683b81d538413b47a8ee1030d8ae4921fbdfd586412af9656993aff1f1cc
z67c3ee8929f43ed4c8cf4a293d8af6ed9642f6f5f86544d0dd77330b1cd8c0041b25c7c2aca54b
z256b858b50bdcf7ac35a969e7350b3530a22cf113a7c5607766b961cf3500edef5cea37f570f92
zfe6e870fb9fccc79a97b149e214eb1a02d81d520541bf7c832eb5a10edd79d2fbdf99a0aded80d
zb0af137e21fa189ae0db5210a46132188f611b7883f31c0b0976ea1f8c8d9dd9e8e9da3fef1381
z895f5f3b67b510f2cd8d06c20c463aace5ee29f982d6effb6353aaa4ae007493d82543c53b918f
z4a8b853418a432fbf5d451d0dad133e21f86c9f5e52638503269232353d6d7ff22b4a90d9a6adb
z43a86153298ad2847282a020d89e7d1b7459611c08f5199e1f19a8267260e433c2ab89f6d968f1
zfb1f9cb4488c65ded311240b8c9f72a5a1ea4978cfd54f196366684cad834134f603468f5f7fcc
z11389f564545511dc66aefc1e1f433d1e2b569c910b340e8d87ebc1ec48c3839e88cd6abd8829c
z50d6f030e29c670a9498c990709a04890d6b72a853d04fc7d0add943d8e07cb72d4807cdcbe7f6
zde833be434fae09f3fcc9292d89f4cedb4769be3438b04443317247d6e7a7e3b4baf79e4fed66d
z6953292b31c58a7134b515e7d33771abc9363a50ecedb5e329bb3bc592677394217b1457cdb58f
z296386c903ccff5fd16287402c8a676634c68947f25ba45f244cdc2d64e4657799e79e636666b6
zc5a1c82b2dba40bf8d39708a9880442c8cae6616a0d376f1f1ae83dc7be7a28b88032ee39a0bfc
z6a45a2ce3d436480f77e104e97bb958d12f95d499b0344ea9023d4dab76a956ed37c1d09122cb0
zd4e7164f095a6b5a7f760974fa6361c769e7153418888ded2d1db5cdf772b9c9a8c751e0101000
z8563c7ea70ab8353ad6645efd2578e823c011b45d93b31a838e96a3958fef258df1bbfd29faaa9
za5763e532b3d54ce4f6c863323dee37575d9ee4ee361a055c9902da15739f05c7392aed3a9b83f
z4cadf373798b8205c38d9f681e57c51a0b0f49ac6b4c5699c31f326ef6111fc7e2a864f2381f39
zb458297d209b32a78600df69384bd455ac41d2e54523df6ec525ab4f59e8a7cc3d49ad2a437945
zb7bb6c2108112e4fa4f71a3474092c9518b696b742bbda8cce527fd3c70e6c002cbc95d72b560f
z23085d306f40bc94ff96cb458da2771917e72985c55a9284c797b03fbd8a3aebd7496c29ce1642
z885b554c677d6b9f126e8aa89e679e8576091bcff35a8f139776c44c810d40e2d3e52af4c58ecf
z6eb69c7cebd97c01f99ce78c665a8d7cf38d603450a19ab62e63ad37f987c8f1c76fcdf05a5663
z7b548676d4d4c3e607a612716c85f22b532bf9f18fc64c6a03d67990433698053c71ee3c03c0f0
za08616d53547a3d5fde4837a5d694c38d9ee8d94708b5da3ccff46a8d272bb96679d91e1e28d5a
ze9649d45ba550cb1f4e8caef8ef3cf3f7a8e1571994f8b8f061ae84ad14d0764df2d5f7e4fe733
z906436c0cf2af52a2fed0dabfccaafe06a84b6cd7407da6138115069748da224f15d21f70330a2
z5c697191d40a0a2a9aa1804cfc5faa54d8f7d680de055a40ad30945e8b43903d2ea22a83429d15
zf55134263ef587ae80e253b7fcbe245ef220dd6a9300728fb0a70e9e7279fcb30506aa348aa413
zede2657679bd706e1114aeeb448eef7cce9f889214f4341d7d58380c23bd7a801f7b17569890d7
z8f2afd42b49733b6988fd39c41a85ca3a2f3fa56ad86022f69f3749956e9bc8ac66b6999120df7
zb2a75447c86138572a67cc039494b214f8fcb445a34e3c8d17dc783986a6088661f1262e52c491
z284e6e8c3846d4d162eb8fa2620bdac7e1668529103c63844dbddf0fb072220287e00bd7913b64
zfecfbec149ce90384f138a03b40d09f37257412e3084b4c1d49179e5de1aec9e0d9017765a64f3
zb66374f6d4e5714aecb6cb783b451be8e62f48d686d153befcdeb14c58a839dfb79fc4b9f56547
z957a7d2e524a5ba5ec586baf41253fbd91735a1e0966bd820e1a396168e4595f98493b154db055
z0fce02a69902311e98d60d1d5de27ab47e9d107aa6203cbfa1107f2c361a4716a04c925a775395
z0147deec148ac0e8ccbd9de2a2e9f659dbe67005468281b0059f6ca391fb085370df7fa0629191
z44183e6a7ab9461e1336cd8c6192e68d7949b7c1a7972d5d8d4965880eed9e5e4394bec7dfc3a9
z821e3e8ed3385151dd07cbc358bed7bb9e27a0bd70f71aaecd7f059be73809c3ea40d67b7ccc6d
zb85354349a9a86a0fada19483a6d131a613b083f98d0665c7f25c998bf3218abc68d9dbc789e7b
z612afdb70774b661632cb009718ccdec26545acc3a60ef7176ef80dbdb7769f21ed65d169ed083
zb8902135b3a477288993c7f7d5d7a272233f8209a48f6d27c4d5af10244868d5caadd2317fcf1c
z957926029f978b28f2d928bb369e7c40176dec4fa144cfe1363c430410439a806121933e3d2503
z3abbf1c2912a625439bb0f7b38937cd6c826fcce4a82145318e1a8f4dc2399568c6ef7987fa2d4
z16b375cacdaf3a7ea386a5e1a9d47f0568097c196b864611afe5836a2fb0371b9450464e1f9047
z8f7bc136139a6ec7764f286aeb55c67e99f8cafb9532fb4006a8fadd0da7f4ea36275e89415740
z8c4ff6775bcef4e6d9da75356958d7486ae92e14d8e439561a73f3ae2483ffe0ed1dca4e8784ce
zf819b22834fe05feed39681ef355e34c43092c89fca783ead1830e3f7480be3089c540ae211269
z06ad287bca8ef0c4d1f8b195696469d65ee4053b13773c24fc93269056bf713ef3002f2e06edd5
z552fec158b64a1315b17aabfd37a4357f1ea39a36777be4e56273ba697c1f4b3b17568f90ab1a3
zdc5fbe5fbf214e351c451d81b5cd8dac8e846eeb12486b66c050bcaf5a2dcaa9ff2f96135a85d2
z76da6454b046efcfb7f849449bc2a70778d14152d9dbacc153d545451f0adc0f4dfad77e9f5a61
z9710067df1bd98a4ade0565fc1344bfbf73a9f35e0bf66264c943433c1c5c8a53bc0da35a4b79c
z6d0127488acc5d78b4ed777bc456edfb29b407199d79c22f436d353373a55afdac93263e3616db
z26f815e3004364f5d447eaa1232f6d6a796a9e975dfadad38a0724250655981110d5bf58eba4fa
z1b8cfb85c13b1d49d9fdf03309ad90c522e53c07d0423638d317236b51dede35de8c0e4ac63581
z33ad3801e7df15570c76e87076843266a7d2256839d61f47bfee80661fcb2a16afcbee0a467792
z7c71d4bf21c2ccdc0bc7ad362e34ac25d4ab942c9dd1345704963d4aa82d064f6eb3f0796bf94f
z4453f88c623282738507689c4ed82b6693ebf5890dd6b62964a032ee4eb8c8f9e2b5ec96f50128
z0180ed93064c933b59de3c55fe7aab64d77421ad3fc74bb90499baf09d602bb5868921f755bfbd
z842284afc080b67cc3de53b443c32ead8b60e8bd8ef050a0d88ba1f595d234c89af331df804dd4
z0d65af4e70fdfc72d43ed831f776e42d1dcbc8f128f24d7b31a491980aed29821364b5aa2c3ba9
zf201a092747a543abec69e48294a70eedc70662f3f03d0c1500a2624548688bc0ec4441be69421
z1481c8a0de81fc458a3d00e3318916671f2c1784063047ba898feb1b61bd7d7ade9d8d2a48738a
z20a5139bf2d0595a6688fe7dd5ee121fc64cd8663546dbc25f466ab35d09805936735805c05a3f
z5b8bf100f654abbb8b769c06337c7d21e1f42e7d2a89a4f7089cdf7ab0284e32b1cad609316235
z4d2301441726397e8ef1ffcd954788738c6182a7bb400ff937b4d8df80028eb15dcf8cc0082bfb
zc5ffe3c56111267fcd5651e0a541f5355e252e5c289eb9eca3dff47a71935ec052d7fa42536fad
z328da8581d5c37250f3ca037420c35c926b73242318a7d5c2d3a333d55f14b96ff503d5a167d30
ze98a611831cc1fa27770712a0d2744231a799ae597a988eed50c4ef9f4d1a4be6ef286f3fc507b
z445efc568ab14829fedfa0612ef5df6c0d2e18f267886c963e3d8ba10e7ccb1a4b56a36d039230
z71e26a3bbb49cfd5d4d1a3639059a8eb54c35b070ff78f1fdb4ccf86a93098727268acefa05d53
zf29babe2a10d7af346cdd310052d935a52b0bbddc5502c184c738314d27100b1981a9c83d11da3
z62f9bfa8ec46298489eac1a3ae71024b79496ad5eb8d1545f9ab27dbbd3d2222090a4205d7714d
z51f44fd98e7dc5fc0c38b6962a6aaec3dd043dc32e5efce2324203ada0bafac8ba73a19d39d1a6
zd83bea0db467648bb1c5350e2fe73a740344a4cc51fd43f129d261b05144c0b103800ea96246ef
zd283b21e1203afabd27af76331ab7977f25ac44c91de9eb69ff533f07319bb9054d08d7c24c988
z3bbcf579f57a4340c42fe3b88f5a9f546a55d1406e82ae56198fc160b80de99718af429aed85cd
zd0cb2ada3a464a9ac9de4c25206163c4e66c24a0a7a1f57c39cf8806f55d7dedd715e586c94ed8
zdbfae74426b0fabf01004f896b802bc92023f24c946203762bf22910d79d083e1796d9e3bb0c85
zca82412433ca28ca450bda2e6f70294819fd2a19fa35b5a734579a6151f386a4a077c571f5ac05
z5dc0c32519ff153334230e7746c8c0dd510821e17e78a61a43bb1114e4940cc414d1f597a5a51f
z4ba7ba8b396735424bb821e35434d3304b17c6bb89f84d364291ad58562a36d0fb7c1855fbe8c7
z7a87947092e922fe1c65e3419a7335d39a43ac07fa612a4b6e444270988f80cd47c8efd4c755e2
z856fa18f1e14e217de09e9ca29a0768e496d779e90fca2cc8baa004c5c478259d1ef0959bff3e8
z32f86fab5974ff72e5dad7f96e0187d6b80fb2c7282b0d4960ec2a693840157bd6f0b610eb1529
za64003fb356d1d04d7396be0577e087bf51408c92da428d7206aa60949e4e4cb0bfc6961d2cfb2
z716e2a2f4d7bebee4841b288845f5590e2c3981dda252d69c58624530db506269f88f1810ac099
zc50cdee80acfa30586d3101e36dc757fbdae8e1aad78e90c25465d764c16cedc0f7ad8ac8a5d76
z9a39cb110a7a52c607c0101a3cd056ea65058b6614f74261aa17f1444bfa12a97b9d9c3f74dd46
z7bfe706e87733c6b6e1d630a756533b87cd8c1723a7bd71aa8fae8a7f4bc879721610aecce81f8
ze9a165a9279c7f6ab4815339962edea7750df32045fcfaa4a61769a78ece58197de97642d8f632
z20570345a0b591051caf6aaee7960ac58cbffd206a66a778afa780699071d90b9e3bc620670f54
z13868f7cbc83af21b4a5e76d53fb1f92f095120e965a3ffdfff42a04605c97e0eb8bd6b22cf561
zc5687ed970398718d0d694fc4d0bc4f0f8b43a69cd8d4cb017ffe8be75a79bb9eb0af395a3594d
z47a8b3f403ece479d87bb9798cba9970cfa1f2f2316e0f73239fe9475f7a2aee718e5a48b6f5ea
z732a37c81406111ba2f952f73e856ad5a7385eadce836d0284b1bba5a61f010e5ed8f9f2fef6d4
z09c2f49cef582789dfd53a63c105b98eecb0e09e400bfa5399933b2f5f923c357883c44557ebdb
za176be70f24c645f69e7f37e85345e7e9b9e1a70a49faab4674a5580ba1d896e37a4bc8e1c8f0e
z544be8167b356e13272c5d68b1e4dc65471495f5cb7026955368209cbfeca4d085372730669e8b
zbbf95b30e1290aa660be363aa668a03e219b46041b0b6fbaebc63ea03ddf4758f2d19d15b681b5
z546a49771bc247db0816f735ebf50f75028a19aa75a5112361d208226e2bdf90d6a744751b5f2b
z116b3c82152e5871507eaf66763327626d8097de749008c595aaa29934c1a9800fab5c6518872d
z3f97683eff32d3c95f06e2973a349537211be0d635f84586bd94cef3a94b8845747c65e4bc34c5
z1a182a1c8c2fc9270f5b55e4e7e141751a23a60f083742b472bcf50fd0a4e8ffcca6a7fffa0823
z17a56789bd00168d766b15f4fbe0bffd9c8edba4e9a8758dac9b63af3f96edd8bb999afa4fd66e
z29ecac2b30a00e052013cbdd54887e37e56763ceb978cebf168952a913a3e0b65759303caa99f6
zf72e2389a1efc2a01da8b959a67e8124bf64899706a177db6f6cfa59969979b18c70e06f92c1f8
z5a7a7c19bff9366ac77dc168aa5244b02b58cdd89164867cea11ed6ac7ec56ee5b6376b6a8a8c4
z735b83175f1c29e74cbb3a9121eeb4ac4dc16cb3ae91241a8d6bd370284b3de0f996e4471da080
z652c12b24cb034ea0fb806b6ff2b5c4cc424026c108d092c14770577b0e4241f2d37cac98c8e27
z9e5e08b68b1b49f34c1cf042c04e6d2578ef6032af08a48f4435f03beac85599e7de7b19f3661f
z9c67d405ffd1ebfab79789255841569f59e4d09df45b615ae597981d91593bc41bebf56689bca8
z4718ee514fbdfeaa92b9cb0b5f585f7e242c4c401fa56f14d7e805ca42636ed1bb5059dbb453a9
z29348d888080cfb19adc90694ed449650d8eb37f3e04e38ae32f04132e2cd71b70f9b7a0053e42
zdb9e219618d686c60e5585e7024d5dfb166339fee45fd99ab3974a0dc809a0a941193052fec35b
z8c9d39cf7dcc3b50590afd3315b4f7fc583d9ae3e237b2d40d93176f84e2f618a3f2913e11a16e
z5e305e875d458611b580d8e44745ae30eaeeba111620cb2385db03bec224eb850697c2d0bb79e3
z1520f8064ca8849ea1c77413873360d55dece93e479845d69d4930f65cf773db886ce7438169da
zc5ec6e3ea0fb71d2ed68db3db8ec605c3ee92181670423464412d41db767a45795a07819316a91
zf2d50649506352d65ef8573a879dc6029aa29e9c541e93f407d51b44ea20c79cb5825d66e75f84
z0ae64f5c4b54069384b755a470142ca4043bc1b0f904b2a4a167d2d01804e8c57062af5eae96c3
z99c574ebff3d45fdf2d8b69f46967e4ac16394384c513d7af44e8d888eb47409a5696eabf939d3
z677d2eb32b1127f3bccca9123850af9e7d488509ce2e4252682307090f50928eb53730ecaad17e
z9cea1d0e15027d9dd71d1c8561295c2303db9dc4ef66cf11fe56b8d152b8c3fa3652ccedec2ef3
ze0d7ee2fbb575f0f0b1cc93b5a9585579a4a9471dfe09f50db429a9bf6ea8c587d01f7133b5e59
z18f3b64fbe85b2248985968c57a1a681b709987264fac6c251fbaa1fde04bcf6cf8e8185cd8629
z314487d14ae0f5ef87e57d9c953d08b561469bb24f49e4cb0d332ec25e3127834c50d19cb48b85
zbed2e05a771027ecde76643e56cd80de9bc0e79aa10b0c303a7d39e43d0d3451f3d7b7263c1652
zadff683b7c4a56b8a9d43c5b15c75872b30b814aaaf8fa67cd95705caf4503e4d16901ee097993
ze28a9871f4bc071fdd17580bf2ce3df49b25adb0154b2b0b918694369fe0c1aef453a48b4e5fae
z1f9e5fc081121f79e1bb76ae8d6b8fac8211cf5aca10fa43abaf652b508f5c48e0c17d0534467d
zfd62abcac683b38fcb45861cce3cc94e7ecf48852516f7d8d78ec0f69cf3f915d56fd4862ee8f5
z80406cf18e437f210db593d0292d2ce0bf8be1e2e7535538d46374cd1a2d90436ec25a91dcfd1e
ze146a9362f8a543d8870d5289d5cc17b55cd9b7534516784e4d966785198eb2c2f1a787e31344c
z74960a964d853d6d2924404c6f09c8a86ef48c500e379ed0f14d9ac0144d2eddf0c70c155bdaf1
zea238f39caf8c149b082904f4479956991a80c4c47b1714723cd7f58fd0ed91b46f7ce75f6c14c
z69d7dd3896b1c8b95bf81d396b40983450edbfaf04a72e29d6e913e713728a0abdac578a964698
zd5d77340ee17207a494d60c05a27cc2a99417648940ebd40a7ea1c22a857924444818b46d19bdd
zd39a3333c9bcacf8f84731e49e67e33ad5234107e7be317f948b133285a2082045595795d2875e
z5450f98e271a523673320bbe580befa95197e15e1519024ab62472622f8d417326f69b70f5c0bb
zd2ade1f2ccbc006eac8b1899080331df1596fb1108b53cc5b36c259fa5aed92bb3cf1c43963071
z554d45fb62736f80ae6ce1dee732de8d8b956532c33ba0c26ec2224f26270ff4b0cef9a8c603b4
zc3b11151d843184646aa7982bcf2acc1c7f84b771b2aded4867ac0de0757e22c1259160f7e0677
z06f83b531934e4c9ced60a6abd1c105bfe5c7d34ea504afcba63490f7334eff5804989d89bdd58
zf81031eabf596cae102fdca6863e93c97e05b1314ae8a6bf17834d40ce488887fe097dab816a6e
z49ee714e9d7ab84c28273870ca11c6f2d42353aae6d2443a91b7f341209152f387162fd36c8a40
zfad6bc85538046e3814ab576785a132365510a05fe565e7803a6629eb2a1995868ad8f409e65d5
z9ee16cfd8e8c8a1d3c1f2ef5d984ddf97e5cdff9b1d5cd951f78828819f721abc22bb7efbd1497
z6aa05c1066619083cb819d4cde76a3ea14aaa324102394babe8b397638f55c62558b382a7e09bc
z58c057e02a56bc033ac4d02e1e3e83e3492efad8866e213d0b642fd60e2e057f0a257e8c264ed8
z7de95469daba4d8c260500b338bfa1ff79e0fb3a4d0941d976de388a4f3ef1afb98e7303cabf04
zc7bb5506227a8890c04f365a9a97f68c0928d6fb080e24255780e5550e25558fa2e52975f38371
z07948a9ef49708b27af92f0b98972ec55e8257b3b687036a9b5aed60580edd5f1d206cc1ab63b5
z7a367dfb246a2cb52d8b57cde56f41483f4e49d26b1ae56a1121b85dd1f7a69e9d7a7c5bae5bf2
z756ba3d00a8eaf8e60c42124f19442b0bff4922a7b58f4e84196b2f4a3753c10869271f3760e73
z8304143cfdbd079d62cf0318854a8a06fa9aedcab680d741a714f7fd5465e84cdda089c5333213
zd6d7c6b4f328c9e83215c6bc1bce5d4f5864382e3b0d7afe8c515cc34f9bc746013770bdc38772
z670e54eb9a4f1e7a15a2b8c6624fb3fbb28382777371ad0a1899c1507465a09fc1325816dbe42e
ze67ed78a9c77e46174e80e854355f7a2adf92d874d5b2cb749d962ba5765ea554c49668bb6abfc
z46cd0726ff5584097b0c9e134da57b287b31700c3d10385e84a14f68b0ae7a1920fc4f9f391473
zf1902ba2643f20e59962c01c3745452ae56104b5b174f929b1ba588bedd2c92ea6da55862628ae
z48913aabdb3c35d7c328282a078307dcce0b6e95234f9d2360c4389c654fc588f47136655b4233
z38f014da4f3fbabbfe0968e59c5174ad3ac79ae84db53ac68133dd0714ce54bbc8a07f8b0e0abd
zb9962a8f1748c196b8dc33ab472dfeaca4340972cec7219047b49aa42a64ba83358fcb02b8b555
zf29902c98cd41c07f15c895f4eab14fff0b13ff99d274157759f04e9abbcfeefb01cd436cd6ddd
zf3e198cc4c37344eaf855c494fef1ac4d6cb63b62415edd216bffaf6774e2859034c404da30ef4
z52cf38ddd50c004334a7fd134a0adab18dddb2acf423a9f2dad09816944583cff6201818704d1a
z88bac101546cf5ce2ea68a31b2f41e5e307abc717db774461c38df3674202ed9fa3412e1b382e5
z212b3bdcc0b7bfd39632c2621e1e75637aa2824f23e35ab1f6011d2cc7086f77f8ce84db648a01
zcd39e9a0500a69e23b2e2a88484a2de3b92c742cb9d281d0b1f260d6e11bbe58c41ff1ff125706
zc53fbe3c232f67182aa08dc710d53f858743f98516807a4169884d83a41d45e16dd0c6634ef541
z2eac904ec9dbaa869d1ff5c4a062b3029fb74864f8ba04523b985f239c0f95dac302c97b25ba00
z1acd3483a7a7a52650dbadbbb283dcbc268e7def7796d4d44e3bf553a75e78cbbce1547a0f8dd7
z864e0df7cbdba851648e4d7a774fdea3767f3124bdf86454ea2753ede1632514b384cfb1a80f01
z5e995c26c95ada8d6cca46251d30ab1fa3ff93a528a6d277aeef674a16bdf3680f1cc2e88832d8
za565dee7fde16e4ca33573e663a7b51a40e08e325b2b7012be69834393dd846132294885a5a61c
z10b091dc821a00a28f948dfbf1f1b339d91a6fee3e609f2a0a06daaf6e0a5ff2454b39eaa96edf
z8974d6457793331ef66fa3238dc3fcf2dd8843cd3463272f316395fbe09999008756af66be4f6d
z8a7ae18dc2fa6e2dcc2758fce266203dba118a69c4eefb360ba3f79e5a698e3ad8d3479ea3199a
zd19405207f5d3da0ec6a1f2274617b5282232737bcd3f3e0f5142509892e21c97767baf9efa77a
z9c3abca36f25b25ae8de8fba959ef505cf4db5c0a005e4ceba551dca2a7c8a1b0f8c9949c82d23
z5e76ef434ad94f701909cadd5db4e1b3f91451caa359d1c0b04b1e54aa3b391d81d165c2475b96
z3c5725a9fdb105cb148a6829be683b5dcb7bb82a7ee737db4d588c422915e0b010fef0cfd5933c
zb7ef00a289b9c174e878ed1a86138078974e2235ea21895d699f55037690d8f81aa1640779d150
zdf23e508b1b788ddb52a822341967bbdb6f234a0ae3adb796ce140c66655eb9784b01e2f80345c
za505bcfc953051bd496c0b10f91cd8694722ec8b15b0ac02d89d1c5d8620b3da1ef9f89d25559b
zed9e4c99315ac3e45c1cf07af22184ee31015680c49cc0b184a627b58d860ba95cdaea39de51f2
z0913bfc8bd449be89bed6fb944f22076f198b5d2fed15c875a23f7a2cd20a06d9f323476635dfb
z5a452f789569941ed701243a1d0595a0f8999ebfd2a7538426c063f67d97621b38f1421ac5f7dc
z235ebdbb352dd3fef88b50f17788c1b3e7bdce372ff1b72f9df6693ce499e5ea92544949070088
z340c5b4107f2e6eafaeb4d4e7e35e394b3cedb7c3b0ae6ccac229c4912925f88a211ba381d8120
z37b08774ce5f2bb78d187e824fa8bbfaf75fb9fad4461832c2e60f71d6e6b71c35ddc6fb762eca
z44e56cc0b000cad4cd0a9feb71fc5129276c262f7100d030fa02897d57f42491a76acd08eb35e3
z7ddc305c795a16e787c0c0bef0b55c3c550d160e108690da9a12f0f6cfebe1eba9bfad4a65cafd
zbbc857cd815eb7c40f581e8e7f2b1eeb0fb9955aaf3b14d1632106c48e11236a26ae7987c7ccba
z4307cdf9108a420a7f2b9bc830fe0df78ecca0dabe4f41dcb928408223908e09efe3d6ada48f4c
z4cb64c1064cb78c7a2ec1e62cae4dccad5ebd161ec12c458fbe15032311e5fa5630e8c2fd1d76d
zd633a95443afafb0d5adfe488c4b2f33f80aa3fed13ce0b60cc10e22905a43b5fc527772ba2e0d
zf829486e7b885613c457b60b393d90a29137c0b730843078d61cce01ed792a09b6a11eab7bd1b6
z861f1a29aa538c5f9f75fa1350919b073e879be7afa4e824c97e226689c9239f68d318672dbfba
z9b94e5da3391b9c412454cde56e593c84beae8173b80726341d2e37fb4d0e4b2a7b02c1572df28
z5bfb1f18b45f82304f7bd9f883d2f0c9b1474dc9ff142f370e0f87c1988678bf0e9654d41e08b9
z105caea0dca89e2c0a1336315978a2478c6fec4011b872ca10dccbf3c3311ba7439264f1be3c48
z25436e41117f2b3fa7ffbb6b8907f50f4747c85cc781c79c51098da4caf206ebc8b6f1c600a19b
za2ce71b89e0a369fe25185af11b9f6ca48c45f00956aec969b586e42b725dd90df00fdd37ded5a
z6005fa024ac5c8b42580ed58d59fff44fca5a8d6f0fe699fdfc68c19c8dadbf698c26439cbe815
z7c292e859c41e4a84aeece2d62a0442fd1142149dc0ee0c4fc0c91abdff86bd0cd2314c5b86696
z50a1d944dc498bc0c6a0c945c1f0d02a7b41d27609e6e9c2164484a6e68b1c6fde1a5132f1b46e
z23d6d9afdbcea9c44c07b0953b27201ffbd884b12f8cd7a5b034401aa5435fa7c3b2f7c0ad8d10
zaf40ac8dc1baeda1915bc29cbf210833a63fdb5d98541eed95c67001e5e769107accdd3e01a9d0
z3ff971c8af0cad1754959285c8dcce2f7c649245511b6e01578e3b15ff3242029ca8475d812b4f
z2d549ad78988ed13301eb10d0f18c7e29842400f223b21c77822ad9bd595ac240c34787ce297a3
zd83d408e8cf5ecaf3fbcc76f2683531f5db656bccc0433f50dfe13b1019898b0ebfb67becca9d6
z661f6c78b8f75b1681b5ea804a73a40b8bc11c58e3c0978e32f4b29968f24912307cca511ba482
z888bae42691c6eae511352cfa669736b553d6e3d6fa969234180502292e4eb0dc35ba3c23c153f
z7ddf0b4aaeed23d7de448a015387764735f2cd0b3592005f2cf866d17a214bdf01dd649d92e043
z4c5379d7fdbf2ac3b66141616bf519ac514175246ee6e6bcb3c1b6a44efed095a25ce718d55c39
z5b4efd523200b8075428b4fae14df908082259eb87ddb5e39df959a4c5e27ef2f1b79d69bec498
z7c185dcf74b7c7993854bc5e714fb84d201fe4a1469332ce540ac23a147f81f11e4c048a3fb235
z733a6547e125c81ab4ec13e85488a1eadea8f274f533ef92b122a0f6b88f0167a357dd0f252e34
z678221266ebf6f50967723c553fc21d7c30bb096aada3e7c0e0df76c9d2afb1f947abce49f3b7d
z419ebf1442b326985b32187e4c891dd05d8230440c563984b44617bc59a01860ff53522cc489c1
z5c14ebb3d056aa3b091114de3dffde49d8f54da60415ee83126c4767c5d860d612920ea8954d4a
z94402fc387b6f0d8aaf46b0b1f9ec80a739cf84c6a734fc391b92aa6abbe05ece126ea3d71a9bb
z718dbfed063e9a031c2e3d0f29abef3757500b4402281f4a62fd15022f78b4c0fa5de7a8d08a1f
zd2d758ee556ac4a946e3c5af6f39d035fe14e3855339511836f08d8f130490ee94b064e6ee2b3d
zb805205f51340955680425ad1681665928b551b82e6485e86349db7d1f4110e635262477ce4e71
z169a27cebd0099113964ac46b3a9197e55745b237a01524392e8914b1046d565488ad098f9e625
zdb6f19426bf56d8c319d0c4bebbf033369c6dd7bed87db6a43f1e572bc8b6829118f7d459e4855
za70c4faee87f90078c5e652e94f25e3c9a025a303c867d72fb3cd781d3f325e3fc760246f67e2e
z6a8613d75469bf368ab9481984418864a402c45f71a22fc2c2c2ccade415f3ddebacb655b18a7f
z08685bf487a86fe1fc213c467d20aaa0fdcd577e838e9e664682531a23138c0313d805578fe67a
z7418765cd5f19af25341b5139c169e28f5d1f0ee48dfe82a47020eb0987990cb767ce3db11a10c
ze7ce12aacce73fe2b69e367c2b95b39773bddf93aec9623ef6cce14e8fb20724112761e48a78f8
z6823436eb7d0200232932a134c4dd70c00d61f6d923fa163c1cebbb9e9ef76dce3581824576ba4
z5e10d70de16a0330122c3162a2f8c1e8a5c2e7358b01c33e21bb880432848a5b8292d45f1acb32
zf06ff6f930352422846b6df53f9317b2dcfb6393525f0ec7f298c68b522b568b36eaba18ec8a67
z8fe3e8d109323a6352bbed96e6f9a219b1435703768c3cfb4a2d8cd7cede6093c01dcb5d04f5d8
z754992d2ba8870fc58b1f5557db58fa9efb40909e77d8a69f59d8cb860f09779825f4e7d2d1041
z7a1a8cc9928c2d31b827cbd3392492ca5762aea16ec100939d53003e62b62f4a7fca55ebb0d886
z4c1a2a202e51d3df6dbae2442b2742a02e1558a54796d90ac7fb52cde9031c8c6ce8819351ecb3
zfa23a001e862ac687596f4a712a985acdb6e6ea197084f5afc4246ef11cb3c3e6bed00a1cd913a
z156faab11e0a16e01f1f9b95480e2d9d6911f173982abdc0898067611866314ba0e24b1d6e081c
zef1a932ac7783a0a3bf8dff42fb950f1e5806809762a28ae35ff8d9def4ad09ea9cc43e9cb5ff9
z6147e91891285ea75af129239a283720845538433b4e206bc2fe835e6eaf1a78d5f67f6c0f43f6
z0d7f7cdda733af991d23378478ce7e889cea80db661852854411397e0e48dadb8268f96cf669b0
zcd58c0370dae80333840a9f403500666a4435ed875206de11a186bb3969f226539dca41db25bfb
zde4ad744692507bd993fb2c67142e965108c547d0701978159d9e4bd6b4556f6e4f1efebbddf2b
z9d2d5056c6450df2da34a5785a0c7f1fee13e6ed6718128a90ad191aad0ae3100c3bfc6eb432cf
z6414c2daa6f84f39b682df622d9b6003e283dc010076c5c9c5d9fe5711e4946dbcfcec25bf976a
ze7afb3213f982bca2da80037bb9f57fcfeedf17470aa7fef58a6db7a2628a4c5057a0424f814e9
z1f82abc51687c046fb940dfa4a00efb96e1bccd893e526f1f6679d3500c93d2d8f23b62eea0988
zf7bc3b410d80b93845dfc61fcd338df2d4165d62965d9cf93e88c51b6043e55b563181e6c25fc8
z3362092978a339fedd1a6832d834801e6fd08d03065f5ca2468185a1fa9f229a2c4562ffdf71e9
z7c8b2e31c0cb4aa7c9ac259cd0ed4a5d2ba1ea98a7dc1a8e694583c58e27dda31f7be38ce76a45
z51777aaf1bfe1e9cd36c50be03f94762e259ba714f151bbfc2c260b4f3f65c7352273cee0b1de0
z99649e947542a6157a6ddf129b0a8b032b5dc818fddff46e0fd868fd8403d36cb28f5e80dd57b9
z7e78a27e48ba30639ad8b001ecc0f7fd590f1e586db8cef3d7ec697b15240cb2f201e7d720d246
z396ad0f4efbd7e57ae78eb9a6ee59a0abd4342445046bfff31a6df1fc3907f66c4498352dd0dd2
z5a5f9345bcde6629b29a9c19e52b18d7175e0f3fdf605c4c2cf63ddf10f2b0290fe11a005c99ad
z817acd1545226baa35805a03ec9a8a6300ac79e287dcb1283714510fd02d6b43fd395b07415c73
z848698d9ad27b7970a4adb43429e46569960f26ffac4a8887996f8280b45a3972ffc5a4897d878
z6ebcded975dee5d2596f68c22d9ce7c1128e4d1255006d32c315e6659e70d32fe6aaab72a38f71
z5d57aea9353bccb1923f31003fef11480f0efc565869fef011283fe95e674cdbaebd27eb34fc77
z9fcfaefec2b928bf0bf9126cb6d5819960707af042ae1370b8479a628fee6dcfa6136e28f0dfbc
zf9eea177671af2863b8e7f244777e6abe6e3dccc34fa14066ca0294e9f4ed5d3545b644fd210a6
z77d820fdc7396ceaa73841f67c2f9599319681b4454fbae60ec50edb88c55e5aa998644695293f
z157b21e72fc9c707d1b82a50eca2a516d990532391a724b6f66ca12e0a51ea400d65b24a9482c0
z5b591c81eb29e00f371aafbef3da71d3724e4d770385810d0e5a7b91156897f76339c4e04633b1
z862f85be18a1ea2b0120a92f271013e0900ecba7e3fab01472a25096292d14a9093a6a7736e282
zf459c2ed449dbb16b432656f0a23f603d4c33a45e67e64053fa39b8acc27895d120b85204971b6
z29b3d3e16072a1d7581b93080c4ef844e545183f385c4360cdd62bfae0e651681a1cfd6c12f115
zf4d83b213f48cc5b73473a2b5649913c2fe953f38dccee419b4e428408a9448f2473a6864493be
z2a64e35825866e08fd768ddf5952fd9c594cd44bbf68a7f0cebf4d3321715466a574788369f21b
zcb85eca7ea85418409097eb1915558f42c82466ffd3545c69907717727a8fab70dd3cd4c09d34b
z16a4430d45de7f16e8261089b969f9edc774d31ffa32693a494cff8feb1343a0c620b078f68b0a
z563d9faaa4e53282ab699451cd706b80d7c470771bca7b9c7b9b73903504934e89e1523312ae5f
z45c61f46be9b3ce90d99f51995d591e8c8447ac4a9aad7d7269574ab2fafdf543d3e3ccb15c7b1
za045ffa2849ca6e45c096f28a6b42363376606ed451af441e4179e6a571ec97daccc4c27b9f0e9
z83c58212b271587000cb4d1231fb0964d37257bad70c5e76fc84e85ec1015f67c2d62868c41c6c
zd2e25de0f8af309085f1a694546b3a728f70ec8ad768679ed3195a882f002c4bd7bc5339b28fc7
za40aa3803291982e4be1860470679cf61f9d90ca54f156fb9f0a5e9b07cd633433921b2e0ebaa2
zda40c9b066f9ea7711ebe4fae58ccfc31d1caa1e0df2ccad0e66124201198a5d729ac7b8abee87
zc49ad4bd2ec8ea270473c0d4f8dcab70e01dba526ee04f685d5faad4b5dcbda563f09c82fd5540
za79a0ea1becfaef847ff7a1b260b0600ba3482e8cbab18101aeab454ac46dffa61c891a01276c4
z4e1980e29d4135985ae4f46344be5d6f6d69e89549bbf4e7673e4fa1e465bed84684db476d5df0
z97aa817ead157f65bd45d88ceb4314d4d9ecda6a3a6865cd1a3794b8066bda9417184df1ef96c4
zab9f22e5f9baa9b1eb8ec001cfff9dfa5478a0fc87872b4af53bf12f8b9139d4d28ec5a0926cdf
z590cde6f91f5932b2bb59704e78ff6923446b3565282902ecd4e366fa8f56c055f75d0f69e22ef
zfa13eb56b8923530a70ea2aafebecd5f529ac06949da6e4b3b6cb5fa64ff376f95268b7a81360b
z44d70c48ee61bbf7ac90ec3a72c4432dedb3d4203f09100b3f0dfda2869fcf8dfb6afe838bbc35
z3e286b74a0bec38ac9ea89947d41921bd319510647ebd0f020e33edd2231361718ee1af1c0a520
zc64b764ce34789ea33c12389cb9064e3e2ed9aec91f5c17ef8a227a9cc700c3eaf0f7a3600c3cb
zf9a933d3774c78ab75c5775f503462be31d37f8ea00b63c8c23f462f9029a566bdf8c54580babd
za2841e78b76ea6d4a71c805fd3c090019aa9f8707c9f557cb07a29e7db310e3919bf24661df0b1
zb8a3611fd693f465b9a745d61a1817431507aecf246fcfd869d8bdb30cb2f1f8c827acfcaa38fb
z955b00efa4451b38c5bdbde5f16c9573a7b9973d8299515774a4365c1600205022d4986c80be61
zc93c2e6ef5be50db1bd6fef4e5b09021c502ea1b81c0f3ebadb7140ef3299d5db11c885d719381
z26e07f6e5002bd327f76ffaa87646ea6f808ea66597daf7c0c5f29cd831080f1b349ad3240be31
z2f490c73ca8b4f208137ac48ee079a5c28a405f09d0af024289d349d5dc1ade4a84e4fe2a19867
z983f9babd0f8ceda57db61e4d2addaaaeafe29372b8e6b8a0f5af490a9602f72d2fb62bb98b99d
z7fbc9e6d349680272c28f5bb543ce07bf280032f5e7c23ae1652befd27ff0dbefcad22e5eee057
zd02a5217f4c6f34aa55bf0fa096a3dd6d1a263eddab1254b3142c891f3cf99575b87becf726c1c
z0ddf822f150c5e6371999807597b6265cd5fe70c0ab628c4957ec0e7be896983b03d057ce19b70
z9f8bc8656ec7e2eeda98aa5ef2a79611aa2ec6786e64b76f92b97b6048ebda335a088ac9d6df4f
zaaa7c9602ad3f312a26ff91364b84db64867261a729ba2736648f45cb1e114e5f347135c109ab9
z54eb3830c1a43e6b3d5d360bfd34369cda7f30d1b61d978edc51da0e7751266e0709a9370e2521
zda736f5cb2d6b8372e10dca3210f5dc44c2e6614acbd285be67308d1968bd5ee64f6c396182c7d
z6b9d19d6e29f5c1da798c142d6636317d32d88f6cad9e49ca0960ac916defa08a0c30a93d7b514
z6ef00d805ede854b297b6e5dda2954d079ab5d5e8d0ebde563d6293252a2e70af0da9088299dd5
z5a342e1f551fd41a83ea445157de21f8fccc96d19e6349614aabc4a41be4fce55313ae12db7ecc
za9790622e418bca14c4cc0864e5eb350b946200a2235aef7f80e048c57637b7f3f754cebea64b8
za4e61fd7f9a20b7e0d4975f6eeeddad2db3401dff862868dd4ec69c8eed93b9a5568c2ddbc7d7d
zf1a0dfa86fbacec06d79346edd9445d1b36a30d0f58e1054f065223b110e07952180d71bf4a25d
za447ec490925fa55f14d13df12216af56decb786325769a1a29434e33776e2cce3f9876f344764
za1ca8a3f79b0510e527795d8af9ddedfe0d0436da651bc2cb5544aaf87bb243738d273e2e1c8d8
z92e6f5a697afcf9e05fa4bc6cfc3cba35259a2a26fb8b481837148a32c4e0f7529c868c90d77b4
z06ab4fe8ea00c9ad38265f930afc32c9aed6e5d3e6e53baf76cb9367b521da1006aa016005652f
za5c749b776b3e1443384cdebbb95eaebdeefd55ea80a96b8ac21eb6824e8538401dfa74278c820
z90c24301444aebb11a64435478d66735ffd149c0cdd2d5166e2f974dcb6ea49edea230d43927e0
z9cee631636b4e9ddc7693226d7d3d24af940f87f1711c686b486a9d117ac019b82c93718e92bf8
za87f1d07ecf321fa613e381bd9bf5129a2315c33e77dc331c380b1775314cbde5314d5ac78706b
zb5dfb4297fd06f39e1c179006c3e0e3ff03739f3e4f5609676a0d92d762716aa00e76c340cfff1
z3af7232a9abba97a1b8508cf19f49042487063f36e08d6f5c2718dcbc86bf8025d7a567516764b
z82ca23b13916c075aed3e058fb73e06ce0bbcfb9754392f69fdf05f4dd92662f20c46ba2966323
za3ed3bce2daa866c4826515801b153d671d64ea824ad83f1b6145c34c6381f25ad21648352b4e2
zf8a663d2e474a41d8bfcc3f817e905c5f7a93045c610e7279e4bd0c4821b60a744f852246653cb
za8c1c1ae620f461c0a101404b83ac971b1d66badfce2b88c240d670919b56a51bd360b449cc7a8
z59510aac69cd2b006b5f6d290cc02ec87ca7deecd44b110da73c140f2a45265fe8b700d5cef5f9
zd3494c481c8077a51dfeb12a031fe8f535d9e0860e895ce623ea6cb128fde2cdcc6b42c5c3cf9e
zb722e2a72695c5db777c252bec486e216a33a2e8212e1f124620425f5ef0ba236865e1dcded172
zcd55ef3914ccf363c0fdce63e793551859cc1a770e670d6878c416b444ea27f5ce4928745f36cd
ze3601e2046271948126e05b79d870497a4aa1763d96f4b4dbbb5fc9ba54d3fd28cd0298c0c7a17
zfd5fa97fca1e2b27756ea3f420762a95bd9c6f8500e069a80f1bd1a99726714c1471dec5ceb01d
zed6e25e197f54f6be97fa2917c8de156fe02af5ed4dd859bf0b130b704675afb3150a12c639d22
zea037d796e370c682530ceed95c3e55e908c52688bd258a7403e4d2f7867e899fd678a3d157805
zd1bdd3851cacac383e6115a9d15c5b822ad4182a12d45ba419640cec91c86135bd2c0060681686
z069267f214f6c1337bea597e60759b85b43bb91b4131432705b12f7d89e6c96818a09af54b3a65
zad5745d335dbe69225b61339ba01e57a34402fa0a2896c428ecf31871de1f7739fa5597537ef09
z0856657f869bb686fadbaf86134ebba31158a9fe6d3dc9fd4b2a1f84e2b99331ae7c06631cad68
zd134e9da9331e408f1513b82c23696bb624b34fd4df1ef091cdaa4409e60313f56d60c8d86a13c
z1ffd1ef117429c10a4e7dc5ba6442a19f5461e3e44ecb8fd0bb760156cd24954ee0480e5d2d8df
zf0d45b7131146861d4846edfc448b0869452b13a20e388e0528a228aa3bb0915aeb5c8ea77a103
zbb2c63161ed2da2fb2acfb630e0eabfa734057cd213854c2ef12b4441b80596ad99277db1efba4
zdfcc7e8d0056d7d2f996835829bae84ba0894cb84240c66c66e31f757ce741984a22350644e5b2
zde3828b77ed49bea094617b8e667198cea74eb397e40d7300be2b256c4125bf9be4c7bbb0d42c0
zb85756233ff1d7c3b3b3ae0929acad28727cf5afc3b891dd0f62652435827105907776a4655700
zbbe7d8ea18f53cb5da28075051b69a7cecfceb092b1cdafc70cd0d9132cf04f3f793d8927c0f78
zad37f4892421122107e3dca34a031d210c24836a40668cbdd5999437ef7b41d47e39cafb3c547f
z44a5138cd2b857c8c6500c6f222693b0868d31a8d51b746c5b26af11f4aabf7b52574af4cddb3a
zce23fe3039afcc0955febae57fb647b9ecd2724d8b705d90b50555529a42a7745b276f6017b017
z62c5130b7d38dbf5c41bd4a9588a3ff141fea8b555c698e99c1819560802d406ab915b7a752178
zc655c1974625a2e3e2b23d3f7bbe12462766f02a3de63466d0bb2103ecb7098bc831574d0492e7
z488dd1a706a754f8ece9f2188f33ed2307f86c84b079af18a880fe7af5f78c74328bfdd25be19a
z8fb9e7f1c0c8188fd1b9450e5c948ea02ae8371d4520ca878b830be16680115e19d3f1230d6822
ze0a578ba2d0a676db2abc40bfbfa2b6f96e772654834cb2a235fdfa6afcbfc3328f9967210aba2
z223b1c093c949da916a0c2d5a0b7e98f2f0c48c0cacfe926306c0dbbefb4802626675c0ab1672e
z7b4786101d3068b5f81c770c9c7defedee23e368fbcb875ca0c39b1dc838481b8a55ed4bd1ae2f
z735563d4c9c63c21c163603cc96e70e9a35d956a392c950e476626c6d60493552c16d9d343a760
z7a46eb4143d1468bb74107d3984e66c075f6f64b57d4e8712600a49ae72bcb646576ddf6d2e029
zc1d76edee076666db11c318f4a95a770e0c91756f8ecfeb5fa95d21575aa5cab13066ca0638768
z5a85dd3efdbc5868f0986fba08683120bcb5859935d9cb0cddceec6879a1e3753a8613c700f9e6
z761dc61f481bb96d7153d9029be19b6666d17141bf501a003a6e30298dde5aea9871b8cec74693
zea852555ef43816146c999044aee4f1b653e449d52a4c6fc3a41466fb9fe5cd8b694ec5bbbfe19
z06cc39816ec723fa6b9f6ba3310368c4ad2cb273cf735645aceb68e181d9e8682d325fb93e5f18
z37bfc1047aee6672fbf703e593a06e5501de52aeb756b632a5a7ac5438d40e7bbea7c8ca69471e
z9700a6f184cfaa607b49cf4958d31716c620194e7150372d7b7ebe1ff7d434324ee706eccdb4ef
z1b406c2807ea1d707aeae633ff59a362fd42c40d774ab602f6b36aa9983cf8213d7a4a17520fd9
zc2438fd23a73b774fd0519504d3be6d04d9a4c178b7150d0b8eda7385893d70c2c5bc485124ca8
zb7dd3259c718e5b16356efb2f69e9361ab59026cf25db5386f5582bd168a1b9599ddb3ece8381e
z1fb655a6e0180a5995d14e97fbc2beac93d888b809810de4de748cfedefe2322ded08db5e77772
z1c17b3c43a9ce74e08020df30f5a1260b0c525f9106ce955cad91853caf82c55c79ff55f0550a0
zcddaeaa8c8ee95322628accd52a0c3247e82f9c9ae6b6913c250e254e13e7dd9f416ca3e3f9bf6
zdf88df91f332f6737a3c89dc54d080e8a2eaf44205ba7d16f9ff056936a60d8f3edfe41c77269b
z2475d407da6e50ee3e826e2d56e6f207cf5b366782cd4066c5a754352301e06767f762464e88d5
zb3986529f63c35833d8457133621a87add89472c49f0acfbeb95d5338e0c1232ae8ed4386dd902
z5c7c3b9f41c057eec6c6f31bba01ecda524ccab28573a84dc3ed0c042707972e744c19071b581a
z964fd41e93ed7372d098df8d73b39b53c2cad154a94b45831361e4d6c692f73d1799c32161c7ba
zef33ed948ab14d115cc81376772bf4212bf9c515ac4f897bfcbbca4e5e171dabd7dc7ed08dfb85
z70e29949467fe781b6b5cd93d17ed68a649985a96a6d1168e45ec4ad6ef0b5fa3ebe3f84a8eb2b
z203768f8abea6644c5cd3b615060fab94115ee8bd885e1269ab2defc0e90c727904e8d0281c1d1
z2a519b0ecb2f4e7906647d2f48d7c27de9568d94babd01e4ec2d7f8df5d239e3f1b53bf7d8d592
zaee5844c2836c261272013988af6ecdd0b38db7b7b7a94076faaebcf943f9e3c66f60ec1412eed
zcb4ded37fd0885b22fee9f192d824c93e876cefe2b42c4b8f53a622de3ef50bfb8088867e88042
z4a95bd3cb2ccdf378e46935c5f12e521cd7145db5d1b131c23d74a1b149692d9c23b8cc5099960
z32cd25fcdbec28e2d47fb4d4f5b8e8e659b32287fd54870628722f04ffa70a87e11f337538ed43
z3da0abfbf5eceb553eb75612040bfaecf2c9e09f433090dab5fa725647387fc40b59a790c1bb5c
zbfd7c2e8301154a267629f28e7a90f3637b3c2f0db9090036726a2394a74a443fb51d10c6c603a
zf80804b8abfd9e4d2ab505616582787bcac8b4b7aca675b788195a286128dde372017b33adb01c
z3be2f948c3cce1fdc90ae411ecca9a1e07a75ed1b1b6e4a9bec3116c59fcd78d812554a149bc70
ze73c5452778308b9b6e9a32581b285f982d21eb19166b44904a4274a9fcc0bac387e7913b5b456
zf220f10a7aee7c41184b836b37b40f221ff27b11ba9c779416a384fcd987f54e6bccd37e2332a9
zd0a3a96c074c7eb0be2c5abecb110858833d395f9b11f1f5524624887a1f7d017fe80a468ab254
z709ce17ae2c4bb053436c1770c494f20bc019c9dd9f5a2794d2761c080832e32014ee91ccdf3be
zb5dcd46260621a84e0e4e4689b63a15913fbb66d9cacd302c1e3b43642426a87fd9138a06cb422
z586189719afb4c1350d096c99d71308650d289a52a32d920fd769758cad64b0bd0d31c2c296d7a
z16a209c3f82ebc7f54ec16515e2fe2af7b9bc21873d87ead7399c813027daaf2ac551b4136064b
z2f620991b2d99c501a2df6f29fecb5d1a4c5ad85f07befeb2c8ed5a0f25b768ff3cb1ee4bf0cdf
z5cd996c65b415ff9ab919f3db06cdf7737deb50c4948edbada17ce8508a07b105bf2119a69655b
z91ecc3fbd10aa9c9c970bf612ed6d48291fddccbdcce1343b38f98558d8194e90d7baeb9158bab
zc1239fcb8a73fc1652170c11f03ffe5b9684b3fc65e08319f0c4722dc5e655680334b00ebd11d9
zee28ee54ede106d64ad9d60c5f499ad749046b5f98fec8d1a077d811be1ad7fd4560a7e1a8bf27
z0fff7dc34708ac3f2386c9e88c20f35a6ec7d8d5f2c9aaff4cf78739fc2686a8bb03c33e6d8d5b
z40df6177827276f644096aec865750986729a834b11533daa21e44cef22eafa9dce6fbf2bf0547
z0d7133cc2783ccbfb93902608388f68568cf579433a4edfceb97cbf4301e38a56142e61b65e9b7
ze74a99a3c3ebb1fa69ceebc6c7a5605dc99f8d5301030a165a842d345246333dfa6fa46edebca5
z063f03ab97161446de524722db2e2f5c5acb594c024a69a233a8383c63148f21fa3320b8b2e989
z1f6691ddee658d33227ea19c56a25aea58bae6f5caf4d6e22891c9f4a4d8736b5f80c9cfa0f4cb
z64e7202546e06c3a7a5d4b0b482391cf9b7a47f32928bfae3217837d03b8a6da41b66c6886c2dc
z86fcd591136978d2b5cd980d81c8910bd1228c428a1e351270d332e8f4bb632b331a7e0fc51f09
z987211978ecf758dd4194b130e3d5a067c052925cf0abd84ff87f9f90284e01f2f07c5effc71ef
z84ddf87537f044777e2cc0f41689556a25a88fb35e715311f0f904292f0390bd43e6f749402e1d
z7baca8f0f04646dc6554f490a04986374fdfad8cb0c0d814ed61d3bbad6c7714ebf6fff8b56740
z078d9ddefed7dad1d97e4de1e8e59dfc16d342acad876e8717a3815d520df7f8568e9fdf46582f
z6eae2ccce721c9628a1c0ac062519bd5ef53248040074e42f4787f60eb630cffdfc1a594f6985d
z3fa86b6c6bb866c474b1191cc57c32f93e0c7f9a3965d6a6f4bde4362766fe29e046c082830925
z3a4a6123d959973a4477cdd3f7c06bd27e2ae155e75972de33971868f666dabb0828e3a5d151da
zf8de1a9ddbbf1d3333fac4d3d690227ec87f4d1729113ae4d9a8147d96f0fde0bd7acf94849441
z015cd7e1228e6d206772859121fb30768ef5c58c877a57f7c956cff202affd33d98d6dc3d6fe81
z03948fdd38c913473ab19a0d36852ed0c174896365ad852f2b0e5619a9b125b7cb9c718d6b00ef
za594aa954986bd4c34247868609e77d432205b2470250e0e68c4e27ad30c28d9b052634e87b5aa
zbffdcb3f497f0e6bf800f53035d12925b689ea5ee1590639b4b87d63bbcc3a0e2d42e19c67b47d
z6da7155fb35fd0ee12c5fdf07a7ed8570aa0aa3fae69713362f1ca5ff0ccfd33cc3cd7e7c58079
za64091cefbc8a79193fe304bc7b3435b7b9195f6eeb5afdfab3c22275f72d747727c480be6fa6d
za8c8e374392ca2292a90c745667d651fc8e3e7ff60bc57f6ed33cff692eaac16e5ad2f3f4ed1be
z2a0a0dea9b2ce5c0388ee7c5ebbba937c9a6f16d69f2e7722f9fa23ce1c6975d353eff1b60d6cd
z520fd1c3cb9a7b985021b88b409b7317541ca8db23f0922f363a81617463cc4873ae95c9664a87
zead7f3c54ef3ed56f1e391776ebeb9505a37e10f60d816fb3356094a5858a229fa2a00fe0dea71
z52f05d73a059874dc48abe10e0379ef51b0b5feaa2a6e9880dc1ae037cfd56cf39a1a6d939407e
z38a6ffea48ba8742745fb219a03a1329257f30fc2d8c00fd70766f5c68c9cb0266f1542e8854f4
zc00579698db97c1765152d7cc85a4be1f301e62204910e4836c596fa6f672beb05e064042f052e
zcd99a3aec60fac62aae71b40f5f6ebb7cc96846064e5d0fd874bead5a67c8792b6c81cef4a2712
ze45cf48d2b397a9755ef01a637d5c11f94fa6e84986f963a472e3b0be44f11f288af7549de0dbc
z10093173cf824f4e065ab9aa38e28bdf3deabf5a476ac90b8ccbc48fd802837238b42f8857649c
z4be28ddc3a8272bd6c353029d6bdcf595af3e72846fc1676b466917040910ad64a97eaef15305b
z16630919ef161d288b9ef7a77d8a08fb3079a0cf17ee8165d0a4b1ae376eabae0286739ac92666
z342b04d0e0eb708c5483668ced6885d8f647ce844da7af3262e22da5adf8763a7c87499cdec561
za12623cec02391d84e55ad1ba6b9df652b8daface56cdf0be5672e0137084c8c8a73a76d2bcd92
z671a712e33090792049c75872ca0753d9371d46ce3a8e491d63b560974accc0aae2f2d8b598402
z587ae4598636c0dc33fb9d33d82636adf32f49bd187c6f3e4348190de2c196705988f2f3993da6
zd41e2b297e851f9a97da4f16c4cb90d1cff497d456c4690cfcf1102d58d805e593e9fb0e101e3d
z85265b7850fa027e0f0c8ed1a57102c65bab6884ea9b61685a1c9af93fde5e32fe3069736a9c7b
z56124bd0f22b82132a0dee3fd72758708c94df312ffbaa403ceab3a5ba3dd393e1cf2c798ed594
z1bdadeaa008813217aa2534b19dd3dc6516e1063e482c7f51bdce5b055a0b557687ca621333ed2
z0ff89ad66a7fdaaaafa0ce6d2a0099e4561e7c22ceace8f3fe8980a8d239f6664b3ec4c8713826
z11b7bc80446d90b393df891a1cb3651fa7269c0d0dc734bccc98a84f8eb79dda3f6f143ed57e8e
zdd7c9e96aab3236478b2a0c008ae7f3998f8325ac9bbc1af8ad6a11cd4a38d9dea708441f29b9d
z7bb4517008a4ead69934193b9946213348c50fa2e97feef5cb777692091e056e096ee4174d43f2
z53ca4ea0c445f9e07ac7204a75a2da46ba10ba3a298bf070f212ff8bfd13beb1954db8c796fb51
z38134382f4f13cdd02449863d077c03a37aef657e08000826d7f02274e0e97d15912e3e6ddcac7
z85ac99356ebbf8558bd1db840db61156eac8943ce2fc8f8baf4abe3f5fbfb31b687b2a4a87f949
zffcc596e6162b792bffe4c5291b9f602184f09b66e883f78347f996c0da1434843b70dd4027950
z53dfaf77adf0dbef90f8e1071721673c067ce50ee05da5bbda4332e4772f9d4f22740476096830
z96f68ce8887ba8c58ae24f175003ab04793216797054484c802c7ae24de4f3d15fe10a789daef7
z7532e6a2531ad1e744ac9e1ffde9a49c0af9a25bbe89cd56db207fcd30596366b5311252985f74
za3cbd4e4f7db18c577b9165b807c36aaec9f85c64ea70c84a20e012437454e57c0256185733ee2
z2f2669aab7afab4213ef728f739f55106fd2f84697e70ee3a0bbdcfc2f2a270c20e8a3c720061a
zadf869cdc966f385f54ee351690cb1243c79823f8f3b6f50c3b243dc2d23040e201fc26bbb42bd
z5a89183c69aef13b0aa2370a78d9a842dbafa6cdd5338439dbb6898c9f4f166cd8e29e029655ca
zc1f1f1c06d3ceda3d12035c0c136c36eb422f9cd18a46328addc8297ca3b68592444d08822912e
z8bf403663d3d2871d68ee4c62498f2ad729c152f9161936bf70f851c94cb2215e818bd17a85c65
zd236545dd8f891e12310fa66831eab3eacb80789d34e2a304cb7cd0ee4ba8a00fa5393814af0b5
ze5f9cc0f149a6b6b4bb61d550269d2311c6e0a9ec9cba6e7dc14486db49a7a77cc9d19aa6b4c30
z945750fc10262fb7eb36cb653b902af0f0ad7c9c8fc0dd044afcd646dcc33526c6b20c358dd7ff
z62b1775d473652a0edc315ed5accbb9721c0af1bf4cdfb29571c6964cc00002bdf05b5f143c7e6
z7489231942e95adf4f577bec908940d87361771699d115ba69db2484a93cf99fdf0193b3a686fb
z7f18b2074d750e452947e2679eb5c2c29992603ce3c980babef3554e76d9817b4122f35020f0c0
z209baf606939b6c62aaa677a9fec8e0dfdc518be3bc8fd87bbad1445ec48c96e2cfd6ff5c5d204
z414548f0436457f35fc60b4322829cb3ae1323aa8506be815de563dc85611ba00c957db9900587
zecaa335b1e6daa06b5ff5e2dac894f3f0e9147237a37908a15fbb2b07353ea5f199c97e08cd542
z55711a9347c45728f578c110e3525305d4ed8913ce64c60f262960db0b551d41530adb21deb69b
z815a10c442c949f0d1e0be99a1847fd19649a5d8efc0bb54d97d73d3433b35bf9d16e5fafeb525
z12801277cb15a65394d8009ee7cae784bee25f77aa746a56069d115da2073b66fc964194de086c
z59b133cd0a505db2825db362866c23584946db0f7aa3dc5204a14f563b8a6b84faa9fccde4aec4
z9259ca0667df089532ef2ea79b9929d599cd7a47be86dcc881d8225da04dee65a24d7e15d2f435
z8c21f754de27eb2136bc50d0cad3792d2ee2aef621f2ff0d3ed586d1e0b5e122e6b8a0d86d38a3
z709c0daa479dfa6200063858c53e3a4152a7ce036159f42e08ae031b978d504be02c7f4718a136
z7f034fa4abd1a31d33f1c2c6458cfaabc2528d51057b98c7d35997985d6315a7fdc57d8ecc1e9a
z1dc1a3fc67269c6ca7d0a001b0b8de775c75cfaaa6793fd7d7d6512a1c680db43cd67360b9cbbb
z6dabfc3e6d440d69e744ff3a12b1db4561e33272bccd92422ab6838c0539bafcc0d6fc513fe1e5
z913781b4dee1c5f222e2a43460127390decda850c520d0bd51e167d8d0ea179593957c3ac93ca9
z074dfe04fe7de73df3835a16e862d7ee68dd6c31f984139041597ae41a56d1cc32016fb04e9dd9
z783352b12e2d13463a17bdc1e789571832f310c7a40ffb8fb96b2a9455dcb8b4d23a4e6a318ba7
zac0500eb723b63a565094c491f95e12635bbb16d68306c84fec998d41e7f8b6b116a167eff79e3
z5c49036eb74832e56c60d9d343645e705aff78186016dc9a09d0007e81f794accb142bb55a2567
z81b7aaa8616233933085433849f754b1f387d5abfc81392c0ab623111656cf85a1bb81b79543f8
z26badf6574d6b720d9a3068ff74642516ecde40d083b7cb5c1dda7bc8b27bf8a528efecdc3e64c
z8283e74dd812b01df94a225b598484083b1a54dd1dbfdb099310c319868353f830c55983e79075
z70098f494c3f23a3f6302b910c763a3978596ad72ba142e5f829faeb2f120ff3da520049dea5c1
z046175d12d7e8f56af981a43ed4baeaf63a626cc4e286f6cb5f74cd7862150d1a8eaa873a4187e
zde1253af2c915c4598af6075250dac0832eccf73c354c0edd777c483d494437910f71385559998
za5f1e6ba95f40c30145672efa82f0f35d4d4e57f1016cc279d05c15d14e077da0320c7016dc9ca
zbccd43b5cc2f595b9fa86994801744f2ba0561bd83b66a7bc69ef15fabb8e6b2c87bb8a6879087
ze23bc8435c0e8d6b6c8984e1832a77cebffe87573847bc01d802bb951dd602d1607c3feb02a320
zeddd3a06c806d657aac1ee8a71a8cf13d109f973eecf988f647697cf95445b2f285207cae1ee7e
zee5412ecbaaa8d2f4fe99326e23da39beb535db5c13bb5ef23f5e8fadb94f2ac0672e9ed8acbb0
z85c57a316a662a497b1405faf74c68e3bd1cef44d70816d2b02d2cb5891b92d6db2a7a0d335e4b
zff5bf3a4084de3a79a1bfa5bb0270b3a46c014b15e7374f97e63abc091d9daebf434907e0ada86
z369dd98f8452556bc03804fd3f83ce69d3c17bfe5324ca168f9cbcf6ae08c8701379a7034ccd38
ze2bebf98159cbec99bf0a490c179dd4147f83ebdac36ceaccff74cee2b8819c70896c2ac5edd12
zee5d26f89342e187a59dc0d3c2009c7df1d8c129ccaa9e0c27f71236ee0809b581e0d09e52590d
z505b03a350f8fe857f84c8516c1802b02b14b3697c0cffb6f3979c696138810a3d76de16f3b3f2
za8cc127e660c605a1ddd7cd4404178a23294b5c928029410109554abeef72ffc4e9f7f98cb6967
z5e58b8ea2231f8baeda48e3cd37df927235d2048853ddf4081e622ff85a8be52b731f3da1fd53b
z9a17c33c78a18b2031a607ac6f51e123f1340eb56dae823d67d5d19606f74c31b88a46deeb46e6
z0b26abe647209cf5da3d1a73028b54415791a8e1038c2129c4393376114fe73ac18a91267319cb
z635c5ea0777d241b0837ff4240719135447a988bcf12774f812daf6b639ff3d8653f464ba61009
zb706643697b2127d1a0f69447f297e19034e889aa8742f001acec39c2f430c01c93e1557b91b48
z0f130bbd20027b6ade9946448fe9d57b7e7ca1f720c79f442ca40c0b4ced65d554d264ccd15ab9
z562471f4c3a80d68164133a8d3ae4be1ee402c928aeaa4a459f2b3fe2ad953fbd79138e498bd0f
zf7691bdb2a92fa8d632dc392f217109bf1ec1b97b3deb63ec56dbd96f0db57e2c46eacf2dd18d7
zbe02786e7a4e6f5a720ecc251666ee168fd88ff3030c86827654ba6c70d740ee49e118480b797a
zcfd35f5efd17b5e6bed549f2432eb8c1a2a97dac2c3d34a5b0a001fde1d0c928a0782f2aa0c9ed
zbf2b3c05f1d4ccaa3687aa53627b8b58e2dabb7424dadc4d3eb422f55718dfda6e2463154fdcc8
zce7dbadad2f1d06cd67d6c979610377976d800525fd8a2e6466382eb9f7917b2d44fc2e599cdf1
z54b274abd6e4867c218af2445f1e50c907202620b4fbff3db88aad7101bda6948426bf3098022b
z2984426a4f7f1c88cbca14f7f4a4f2ebfc2d563b133f7961cb80b9909550f890ec5b4a40fded24
z60c3924a8e9a095702e4ba5311bdd5c0b2d5891703e4abbf0fdcf32c3ffe4e9a7a6ef7d2b5d376
z4db095ea688f60e3ad87d5606cfbc4a543ed95104001703effb6426a34db2a0994187991fba672
zeeaafa98713c71b0cb82ae82cd66ab1905142ce9a5bb0a670c102b6beb8c3e8250683358d2108e
zd5b652f2ab32a463809bc6f3e173cf32430585dcec381759a5f5107907499ed0cb96a4a3cff1cf
zafdd5e6ecd694ff491abc4c9b0f3353f6d9c0db94f84bdcf938dfc46e4212373efc5067bb99285
ze6046288eaff7a9716a81163e517631062efea0ffecad916cc23ec14a542052ac9093cc310eb00
z567af28269b7cc1c619e655cd68eafc30beb77106ee9812bbb081e58936ddcf44fc54a96696931
z01b6212dace16e0f4a2a389ef3c97dbcdcb666f112ab3ddbf2d00d61a667ae7679f0b48bc80053
z4d599cc3bca2e5ee95636820beed096b5c243dd7c76a689dcab79105d5077bf3c87e47b71065d4
zb857e92859e1582dcece14ada1040970c4cc3fc5fac8ba9dce83e00aa8bf1ee893e7b11dd0ab65
z9b9a3d6d6ff06aaec36a96399860be79ea4c928d57edbbd230f48a13270c50b5c4141f78b06619
z333721198a7b02b157fb5a707524fa491e52bbcf78b2feb0af0d770b2b79331438922a654a4ed1
zea6a604bbdd42158508ae71f2f89b66d1aad8a047b0ec94d974c845e5ccd8a9e315b1abdfb084f
z5cd82db231830003d6516a1bcb2dd60e5667deed40bec750e98c420c7a5f4baa59c84fb0e8239e
zeab392f8a576b8bb805581e9902e24c0b1f523fa132715498895c4bdfb14277cb29d2836f6493b
zf5db1bfac00ddddd972a8d403e24fd9001ffce742d8797f164ec66a598e45fc830b6ddabea271b
z378bad3e3c542973ff0becd0b7e643b8962f5ea69d93cc8e6d931aab4740726c337bd49cd2c05d
z1c39f3fa6bc18fe120b752e8f27180cf8701a67581ad96350f0543e13b48b59d738af9214cf6cf
z5307b77ecf66427a852f135a7c33afcacbb1e4b9a466e1106970bdd10baed2e90bbc993d78e5c0
z7abf85993c4d6a17144d73191a37292637c0c6c0fa440f2d6b67aff3ed2a4b0e69256714d982ea
z0df027873eb97bddbbe5123d578e6f2a576d93ab772f1115e88a2748aa9088e811fc95a6ab1362
zaa08d748714d82c4ea2c8f305fa245d00715eec65adf3da1f27497177b62abdea884a2da0b50e0
z0396e033e516c9ac11ff572683f7512a14f8d350c4b6e427db47eb156d65314e71fdaaca75ef81
z855637d8b398f57f0c04a771a3b44e81608fe3efefac2ee37175d09333d63582627a4146ee5162
z7ec1ac7a807b54ae116370939a7981e06e8c35542b236b95fdb7914c71d69f1a71cdc0e04154e5
z8491b2288380f3d2c11b6ff600d5561e025bcf99734618d9fd7b23d3b6006fa45b6fee77f2defd
zba9c6ab37b21b770084681f2f762d01178349defd2b1e723efab9f113cd65048d8697ccfab4874
z2029fe904d2c56ae972679f287356431a255dba7e29ba1ad2c01bcdd1fe48cbb20717b61183378
zfba150ca097725f6687e4912b93b0b6389e3d88f25ccd4317e313c02ea5dd6d2d000d6e0e2dfd1
z0930cce7b1c1996e7a49ef1b5c0993055033ec01e9777c76a1c6e5e64f6ef0457cb4ac43a854fe
zcac10e3b93ba60205c5ad0b5d2dcade78a653305119493ee8f5183beb667d6c8f98cdbfce7f1a8
z67084236d8d3d2b629b5c5e4ccb3c65fd0648872e643d2a16b0c52c967ed2d4f0cc23b07250ded
z593ae208091e83d18b618b1254c556f99216f36d202dc92699f2ee5670555f0181efe4a0f132dd
z5764173727ef0b84d05ddb41242e30b6ba094573722f0e7df7e7ce8687cedb50fed2bb8d779e46
zead3d8731e7dc1cf7acc4ec8728605cb6ca694beab86c91a5b910c044ee0fe9ac7bbcfdfe92267
z95fc6b2b0b9531fb06fac3512a57979342dca94172c8efc8fa36a0124c47d03a1df0aad36836f4
z854302322601aa70d00244ac6e26a8a3d16eb14630cf0d0e696d2345a3222a352dc2ba44af5e75
z68778c7e9beb68ae191ab5823c1859925916c21466809e8ae7cabe9daadc49c64e9e77a9550360
zf3a24313468fd4f2b7f7518b0124cbf5e5f04b685847bb9981a4608266fcc98e2bd540128770f6
z2fdab5bb6f5777ae1d89b06f335abc231a5678af78003c0cb70bdf768ad5fc1a09a9b8d3a12cf3
z19953d1cddca6e3e83cb3e7ffd3c4718bb69c889dcd29a1182ec72425c90da2b2354d24cc6dd04
z32d474fa518f7325fc5e4707effa5cbe4cd7e6143a70c52f07dbc6fdb1aeea3eb8d7f3a9d77d10
zf07f92b61e0bda28a83ea8cfd9d6cf2597230f3b1df7e5f8fb5474758f894921b88a43d18c6990
zab973378c6ded63906d35bbf627602b210649ff443f87f9c55a322d1149edd939fb33a16de6529
z62d7336b8def3cba83ecf5fccc55897cc986c75ece73417fa2913343437e01d1a5944a32ac820b
z74ec6e15a5bb96404c275492d73843c8eb85ee5fc6b3beecc9fc016671b7c79b3a0833a3ba9472
z7cb4f12d850cbe56798ca6642ac7371b2d0fb9f7ef1449e280b777e8a2f2cbfeb1f7129439c91a
zff6a6a04b3692c87abd7b0271db7afe300f528ef8ab27db53bb13bfedafdfb7826722e2a9c0fc5
za98d3cb58214b77d134eaf16c663df0c594016d9576660104ff390776887ba743d2dd6189561a1
z2afbabf7d3319250cab7ef71b0f0fa6a97e388a0dd5b28fd38e48e84c2b1093e5ab79b47c61016
z835b601f1d110611a457f7b0150125e879463fa0550ee40cb6c30a68004ac2da6306e1cfb51498
z211f9a4f96e69a13922ae6a31323a84b3e49ff2901c6443e3c19a9b953a85389226b858d354694
z3490375751a4c8087208c37efdc825942d763a75e3931fd80fb028dce10792ec6097861d60282a
z011c84c2e3230a8e4a4e1f4299ed125a374b6263378d334e8ef002a45045f1c3bb1c6c0a966ebf
z77b886420b0957ffd6bd5e84a9d3cfc1840e45603eae7ba6f7bcaa2971d049ef9504eb308688bf
z422c503cdfae6824257bd4b4ef8f6d3295c530eb6096382bd54bfd714fa86c4f862ccedf1a2046
zd54cdc7c43cf1fe76c86bd2723b59f57f385d378c05819f7a2ec54b94ac77a1208659f920afbf4
z0455dbe5741d3ccb2719204259a316346767fec7a7385c3aa0d84733d6d7ac148945e89a44be82
z8a4e4a1bc874ec31099c32b69936b5dc1c5d62d4431871cfb95f41ebd6bed02e1dd2d51a6ba8c0
z90afa10effba925252cec5ff090c674175223337e3047bdf7ddb7064bb6cd588f87a6f8d444ac9
ze58e9d064ba5272681e97400fe5d396fc9d09e11c16df1b378b550fca447ad6693b28421c4f0da
zbe520c08e9dbac626b1db096eb8b394b76b9872f4db058f46d05f23eae397049c43eb9b9b6311a
z51e0af7e7916c860cc3ea075f4782c0991b773affd3d6d34474d19e5784e78d6f12ecc6e236180
z50ca36418635539519888f3e2ae2eaaa58f612faa6be9d4a64a95f2a881db3b803318a7ffdedd6
z6ab497274856711aee444e130f222523bbe093db9011d76db0a3b869057c16719ec1d906a4345b
z5cf7d6c34206bd26ed89d01c63c3bf039e5d11fb5d11451d204f4ce5444e354cf577f0222b2c51
z9f543b13f352f922d8f7f0c4a59c843989e5ce24281e7b165d9f5d5f1e274f0a2d558bbd813402
z2055e6d3ad221ec91a3877923f2b68fde3e8bcb237da75c68e79498a641dde66ae4e5adcf01982
z0509f717e97b4c91925d939ff7048ec6df88285e75aa6afad9ab87ce864990b10a658b5f7e6203
zbae9e71d6f63d58a53dee78cb8fd1ef1b2e82f7be665a615ed710a811f7b7ac1121e722a4de4e0
z9aebc29e35f8483408aca35e59392bba54b43da5abaf4418606f7ea04a4868994cb216f8459faf
zf004f05fcb62d46a1f61f782f3ad8e92c8d8452e19e0292c97661a043dd0a936946914bfd20827
z169bc777948c342d81fd86190255b1381e87fa06bfa8fb1d9d63c205816d6633176e1535f228c0
z8a12731d433dcaffdce340afaab5bb6b87e74411eb1a891c4af799a3182f0d4fa5ad6be2e5c018
zf293741e201173d572ba47e08c82580001a61f3fd49cb9cd7b8ceec334857e7cc1a5acf3408801
z0c6745ebd997154ed721eec70f367d1ce2689d4345653755f4728ea8a66b17a336a154a80f8439
z5300c1e870f74439d3de870c31f7b4e79aea485c352d06023c331ed935fec4f61d1536db0bb961
zd40eab9b3c827243400fde894d27deca642dfc53280564c4c8946c528f6b105b78ff7c78767d0c
z431c55015fddb6afcc47bf92bc76a256d86ba9a2cb6016e35306d119bdd51f051909633f36e2ed
z59cf784afcc578474a4c9a771d09022005fe8df45a88b685b4826db0c5982e2c3229f179e6ce71
z50aedc62553038d21866fd76de4f1f57ff51d6499a561029f1bd30295978df448ad7a07d93e900
z603cc7819f5826cea75599b11e0dd60fb4745ae8f948e13c5a65c9094dac2e019345ec6a5885ee
zd65f0809ee14a90279bcd0d4521f95efed156bce4f99c2d69c19f9c63745aaadd6b3127b11d8f1
zb59839656cbd35204fa1e3f43988b4b5e7df85e3dacd68bfdd68919a8a7d1c232352e05a249da3
z0269a70fb69af61412e6ce236beb2fc3f16a2dd65a1508843c1f35ce365b5be693459e405e7997
zc2efba49a56f6449ade0324e678ccb8f115125a748ebd8e69e7fb3952f64b1f4734b958c3c4827
z2b1d4df7f03d1c7ba743be95b837e53eee928d63d37614f7c985ec6503731f2dc7707ae6ea3c1b
zd85189c08040ed09c32a69272b02f4b1c8f9587a166beee55193438987cefccca16f4a5e35f790
zd8db81ae287fe8b0d57a06dec03aacdcf429b8100115ee40b8ad6c017f44c93236397b38d1da9e
z3270f839fac0711efb8a010144167f3ab991704fefd331d82c5dca5dc01ee79d4d3a8732f8ccea
zcbfe8d334bc7fe5e5fa232f8f8987de7f16f61216edf76fec0c4187b6de19d93a6429bda81e6f0
zaf55f4ca484b2edc3d54e6a97991899d9493a3ca0a1742b3888a08beb16660abcb4da88f36161c
z4440174701a244a3a331cac375ddc72f02b96747f263968ba94521fad169259548eef3c2507362
zad0fa3c6b22ac9dfb55b0ae7ec184f9d9df29c7c1d810f6b95c1da5a50d889221e7f2fcbbfd8d5
zd0df03e9cf057f7109e92307e1375c78506c21d95a1b53085bb2f6c2bb3041288386e09bc1df39
ze95ead4b1c94296a2802d5e76e4f96b458c485422379513d7d43d7f731cfa3fe1b5d60b1824ad9
z9b2078c3bebbf5a37ace9419bab8043b23772aae2bf92e4903f70965c37452a3b3f519276ec555
z5826585a086480b0f0d4720baa9677186d4b9d4af169c17b6659db3066f54ecd58906c58d64493
z02e3e9034fed3eb59d7a347dcbab6cd09284366ee68e0d32c0560fb59241d3846142e1fbfa81dc
z1b919e230bbb2a4506f8d667ea3884051a209b2ca6f10448ed7d203b031960a49b6e48132737d5
z38497110d7ddad9f10fc86150f0f4ec642b53d042181522c6faac7eb6014770dea7b59c5579982
za2d6ee982c34c0fc60fc5837e23f04b467def22d1575cbb79a75dff5197264bd3e4f4ba7dd43bd
zcee0a5f175d2bcdf7a1639af5a59aa796003bee77ff39c20f42474ae83c5c3ff95af27ad2765a5
ze55f0f73883e8041f202aa1fbaee02be3886ea7a69ff8bc57bb1db61956417269a6b5e7e9f6a29
z3f69cf892fb3fc0db04ad1a4a46458d6a823b8242993b8f81135d7b36bb6873b1a485d7b653a63
za316470d02a8179731aa770bd574db6d82c993bb620fdae8722637d4ea83b8d71ad26381d7c075
zbde8b1914f1cda34d29267284dd9dce31788ee00e7a1e98e803ce0c230992d992ed473a67ad82e
zefe447a0579ba6d09a556223428aa77034a1891c36615bf2a2c24d0f2791e28cd74de9fca9f530
z8816782099e760d06fb1878662c105b14c69d9c164d7c221fd43545f50d995b765fb998874dccc
za5853690d5bd1bcfc3aac5c195d895e7c24c135d0e65f7370be90db0c5ce13b06619b8d5116fdd
zedf16e46a04b31ede9d4ddb57291ac66abc3520ff5bda644bc79e867068a4e1b23357ff59964da
z0b212149618759ffbda2f113b42fea3b72f0612abde22d6dac99bbbf2af47e98e6d3a03efd98b2
z7df0a25677dd45fc798458b3a36782be712f6cd76b30363f1c0edccdeef457bdaf24a23fee0708
ze9c1124af7c13e1c99c8292f853b8d25cd9a6a5a2c21a89ad57522561e5ade0dc9bf3ee256a7c9
zf087597f53ca3b06e6c49d4ffaf0e0c131f8392c0306c488283f64eaef09368d84b031b9954c19
z091a559d9d83dba613c6d827106053f0ccb64b14fac3bdd173b27f27f645561e267aff49aca336
zb5fbe552a92150129653f4c79d6845d07ae24bbfa13812d25092d96327f34b23ead16f37532219
z5b6e9d20217f5c1ba1aac5e0dd08e86eca6dfde3010c1bd3bb0094ff315bf1194776bc47291f44
z264271099658b0e3358d8a79cb8bfcb841982065628e4fbebdb68df6705aa3021b245c92ba8e93
z6d63938e8c8f55503620d3bd70895f6137d146c2ea48070079c0d7212f2c0715e067a8c4a62c59
z22a0790af01ca0f4e42eb8862975977948b28adc9c99d2598627c1cfc26e034445e72813ca9807
zecb77c1e58644dbe023faefc349b8e501a7a63c3d7df1d63c7643dc967130f19f4561639909e35
z276cd1b6a0138f4078f10f23295802410e62702929e9f4792138b1ef2a314124e48cfe487368c7
z2d1b28027fef269c68a6b480ac52836d1ea558d630905a3c3ef332246facb78e85654c72bb73ab
z5de21225c56e3287c7242a2dbaf3d787c53374ca112cac98b719343e6f4cecc63a23868c2e3779
z50089a3fb9fe2d0c204558268f7a78cc80cf05a35401090381ff395b89985d9f0ff0567858ee7b
z3d57fab8e4b4aeb5ecb6bda60f244d85f628b0dbc56d90026b4757decfb3bb03b55891a0b8f867
zbe795d9fb86d40a1c2d4b5c7ffd90a6ad2f1e9f60a3d14c940d29a2bb49353622fd4e70b588a14
z333fba2b8e63bc6a5a724462262dcfdbfdc0aad10a10d72eedc44d070525f1007facf7ac68e9bc
zc210636cf4e97d8cd34b8cc843fd4373936d66d36442e6772206bdfc6fe15939724cf358b0baa5
z0ce604e88df5513268ae22201024bde63b61dc821e6d7e534f30a9807df0917ed43ae65418c9fb
z9cf285a6efeb1ab6d3de618a830a7d529f798ac2f373d6ce6254fb13bbddc19ef9f2f629226c40
zafd7fcce6c4162ee6d9211d0094f89937e468fb0dcdf6eec775ccf2e2d7e1f062ea996e62db9b4
za33a6f50961a5a308d963eff41244d14d4e081dc469aa4f180346747632118075573993ebeddcb
z30df7977464fe25b36de74024a37ff5dfe6dcb51c58003e1987032ffd6dad43c169cac9f16ead3
z26e11c39652487c6ad997a4a2a02fbb7612bb81a51ed556f2b1ac95237ad34ff87cf13f6cac8b1
zed8892aca007be38d65099cb97d6f792be1d2e445d2672e9a9d1301349a1eb84bf08355effa6bd
z01a24ff44cd971616802f589c29105b4008d27fbe8d8ad5eabfaeb58b52882bcb2c444961c6d71
za3a4d5465118ea2492907490628914b0ddc68ca1643d9f13bae26ed2a776b5998726eb57639abe
z15dbc654344436df6272027d182ed0f57f8a55aa3b55dad8d7e8f5d5bff8cdd042855ff52799cf
zbba1fea1d6050a76bd82f48e5a66d5550729b6523f74f2d7bccc3524deb565ec2699985d6d25f3
zf7a08ad021c4797586e013bf3b80c1a0211e6f28eb8a15c67574376e3d07901ba8a4ea5f825ab4
zd1db47232f38940af24ddd46803e271e728d3c5ea88a489c4e958a43b0c51e2f6deba28459e8cd
z2b5e1a9cb6bd8d7dd5645db00c67845050e3108792a629a54ee4314822e706e028eda7093bed20
zdbd1c82a53ab6748284bab7684af7d32f11a0b0bccdd69e7f73a7f2b110e97905b0ced607b11e5
zb9a0c7a79af9f978740195c40ed0069b38c7113042d2ba1167c88ed7ee6e1751314e347f7e0fa2
zeb84cad06d9da64500ed8c21b32d22a9af520b1e148efa0145af7cf1ca6bdeccff777d923193c2
zf6e4da08aff21b06ec4bb89b9456f187ee8e028d5005e22a20d8c36d1c7728b9674cdf916f09f5
z2d65f8bd17ddd7849839b46daeee5af0fab23f548c018da3a86f765edc9d9469edfa5e2f5c74e3
z9e6895ad95e6c95feb464fcf16222e46615cf6e8046c3242d7cc60267eea43a4765fb44d4ddd4d
z743aefd61115995b1e1a7b90b7f0bea46bd06a2babafb54f4d595b573327a6955ca835c9d14106
z313f98a360c6f866fc75a381302a95c9cd5dad4b32afbe329143bac509872cf986096a94c80b5d
zdcd2813d93b9b72105fe9f93c120488d7f32cb1125a0ec42b7972e358c31f885c903043b4e0520
zfd004f2b189346fa218aa42bfdbf232bf170f68420391a2bd20d6d040422e1a21347ef9637e486
zf51cb8d83cb87bceecb89144f265a40f94a87eecd4c8cb377e954162e2c631ef34249c4814ef02
zdd1611210fb0cc93c98bb51132d3dbaa53399f47fa4f2c97019e848f82282089f5760222c653b9
zd2ec45c36545e3c0f8c1dfd39ff88212cba015f1f0a5e0c4fef1fc2cf166eb57e8160b864a81c8
z8010384664a4cccee401c61bab0905f1f76bba0d6f5207e1afbe3ec69590b6ab4925d22426e8ee
z25ddd010a018c786a778cee42f048169ee529c3de49c238fdd7634ec2a7156266b9e5fac9ad720
zcfe79f79288fc5c2b961a738fbcd17b023f1715e443d42939006053871e0d0064c092279c6be41
z9eb72da5781007dd9b97639b442b1788d8befe6147a7ae935eda6ef2491fffdeddbdca3612047c
z7c244a5bffbb79e6127c7e2a0a457fa16eee058777dd9ee29f2785e8661f210e6708e061bdf73e
zbca0f65d67cd1fb463662e56343815cc2e14aacfa0959422f59555988e0574622dfcb31782b2b8
z44a053bb17417e5a414433dcc82694b17c73638654ed1184469a6764f3dbc1af4c10dc14b2f4c0
z857e7c68f418c419f9377ca0d13e8f6bb608a7b8f3728bda0d053d53513fe09eb12da10feff85b
zc22e4096232d888d6c796151bba6031e155ec131349546768b2f06c07a9a27624ac7cc0d73fc78
zb3c52c6a7b7fa065e94fe7ad14a84937cef4f8d3af33abc6d7a25d6d72c7130e3640147403d3b9
z635ea01ec6c1f40a7cf2138de0619150634c2cb547ddc064922032bcf123a1502066753cca11ad
z82675d8b5dbf6e2128981c134bd4b58790f712c21e4e4ce2929d15343ac41e67933d50bb38b92a
z3931685ff94ba7cb9b5ba9e1927dea7074b739cafcdfd949c2b5bdfc1353e5fdd99c81f0454a66
z97f2f846b8abd9d2065e159552a4e793bfdaebf83b24eb43c2fbd212934cbf507cddcea4691e36
z41a8d92b6c13b1970871f1a3eadc55c496ccacfe65fa0d70a698fa6865c8d8accac55c20b9c8de
z04aab9a915c6f7f6fdb555ba3373de7929cc61c42ea22344ab1860b93f729c474297e7113bf8e9
z000b30c3a6355adf428445729629a26eade4f8e1e6c579a7e9d0d2d40004350596fed1d5dc3979
ze6245ab0db20e7cdf27bd2ee4150a48dd5ea9fd27de200d916270b9b54ebd3f791356ac77180b5
z54aefcd7d913fc274eafb58c4611b6adda12e164f7c70ad8a71ba8eb7643dc18b447b0e30a95a5
za7fc16b734fcd3a75fbf61e0650ead772b4b64429fae104fdaec77fc23d5a50075af9684c61cb9
z4f91fe00bbe5d23a5acaa06d497da3e614fecbf440b69a880fe9075581e0746f9ef15517344d76
z1939581b077827ba3541f76f1a015e8362728352fcc10a4cd46c23d1ae14224de49f7ec9ecd82c
z2341872c85afcd9b3f3b380bc43a9c2a8f67bf3a619ac6b48f89e4582619759c0c831e0ea87008
z1ee879b4ce8797607931edbfc10480343d33047b89205fb3b961e0865e846031d4438c30ae5bb6
z2df13d811fb48eb2e0d11e3ec1ad672523034dbc2f1d119293b03bd1539795337c89edbd2fa620
z5f1fd22a17fbee285204b7d696aafdcb9a7a3b5bec8880f28f69d8f14b9c872d5703d34115df9d
z1f85677cfd807e3c3ee7b4ea2426800fbbf69058f5eaa71680e3f024d405194b24d91f0b6c99f6
z154ab3ab28466a17956f5976c3d726e9ecd484cff2e89989e3c400e98ab5deb65da96ab020ca0d
z75c292af9e40f88321051f9603fdedd114b63558beda3509f862697540eeca8d15a31c60617457
z340114f9d06c7b2ce04280e4ab456d9e2acb8a00cec2952e26b748962fb3c660677093eec210cb
z1dc3e816fa21798817cdec59060cb8c6756fc5a53ed57945671c47596a4defad81c6021f23f00e
z4b8c8ad77764271cfd371757fb048a5e2e25d027c41fa45b2f0c935b52a3ab9311b0dbfb3e23df
z00a0cd14fe2d3e2697c6996d065964ece3f617d235dbbb0e3595ae22dda0c0271bd3ddfcf2ee31
z7c96da1254708b9183ff27b1bdd392b193e6ada2fae988432bcbcf8b6c3cf16edd39548689368c
zbfccc2759b26966c38156cfcf280f6dafd03d463f2a7f014ce26286002a8ce12c7c3242a16b996
z5f18a191cfcb77ea4b0571b78e0292b376db79f1b11ddeb109643ecda2f07b099089b76edc808f
z0b6b44fc4401492db3509b3a8b546e59d6a5a8b5f27b3ec3307f4ca7d65f3e7aa94f1781ac0363
zdcdf72dc5ae69ee455e9bce79ad519b33d2c8f319fbd6d6b0ea7ee22c4e57aba57210553c84fa3
z841055d0f9db59b39b714933c5edb3d1e84cb35e5c3ec104e41d6bfbed76bd87e8c5fe38e159cb
z5032ca6fc0d4b3928c3383cc3ef4783b408a70f686336af080984cfce557a5e9e3d0ab075d88da
z69fe3c83b76f40c0d541478e5f1a1a81f9cfdafb01d7669b0f98d2043426a29560d53e17feda0c
z1cfa81d6e5527386886e01e5c11aa3864bfa6cde840d5b7b9b05daa2b3297675a02f35a9db02df
z8d7feb562bb820c11fe9d64719e44c72a76f677b8640781743adbaf9bb4f706cd53f1c2dd436cd
za9e295b236540b39173c4ff4e1c42352535ba40c20c8e4cf977854a92a33f6b323ac4345d356a4
zb065ae12acb410117b3d7791d53d19b52c3e53ba4c94925e761919d5aab1c751daab765f24f188
z0a7f8aa713d4b43ab63a5a68b0fbaeb9844f364a891e1120be0200fbc84beb64de01b3fcf6852b
z7091a52430f7b96a35cd1693cc6ad8049e96d6e9f32bbf71eb062f4a59ccd8a10d5908756dc8f8
z47b1ae2675e19b1e850203e77db8333bc72ec1c240c663280354cdae73310f37a45c1adae36ae2
z0e9555be597352c6b5a78011d840b716e2ae38899b8be14e5d4b64ff8cb5dd1c0257b612cdd0de
zaea6e06adfe90bd5f9c4dc77374f637c59cf94a2049b9ca44688e0ff508e058eae4566b60985c0
z7406f1dc971c66e3ddba2ef4c2179629969dfab829def96448c5a637c2c3f46a473fc892c86931
z0b32abbc33eda9d5a22f6997bf0021449f70ca7fda829eaece72ba89653daa3b22d8baadce2fbd
z4fd4e26065f139e9a21365ad2bfcced466ffc89b9e67637eadd4ffabe03f7dbbc9f39b5bbbb095
z7459cdd6aedc3c65a7bd8d7d78622f38513d89882ec3cecf7cc988f054c82133d3279aa2a2a3c6
z8a33fcba0acb27fa06d756cfaca6097bb37c5b9e917c60f7f2820698dacf61a47986faf5dc93bc
zd42d92918684109f5c63a0d895e7158b207b8dadaed0522a4e531d8d5fcc5ff35f286dc5d0497e
zfcea7c76f7b63a59fcaf497499c451df35542a4f0fbae3c35acf17d1b90adbbb94c6a420c13bc8
z5fe575e905359c3d3a5ffc0e3c4a81635b95c9c5744b0e92084fc47c895c9cbd80a2ec5f528bbc
zb5aa407029f711fc2ff01dc0fdb279b417eede86d8f61765a18232706919256c5766c67c61ca2f
zee3b724cc5884b6102ae43e1410e228268a7564ae16c4a81d61a0677761b6fb1c4b4f1c8eb67a2
z208d19fd5494496ec664e846291a55d03e4e3903db8d81f6b4a510a1349077a70ecc70588bb1e1
za6aebc90628abdfc9bbeaba6f63dd4310e799612f84256a8f398dc997d8588533170d18ef0e91a
z05139bcbdfd8e99f63279be0d7ab497daa3bbe02c947aa8bc6ec94c348d3e8d8eb5346d3fe0f54
z6b2efa45f3539bd5a243c875d4a92611acaf0ebc8d6d3eec4cbb494e0bf002e577cbc6df9bd01b
z0780473e49ae172b91f2c535736e6f329f4bb9afd8e06e53a4cf23d4d4cde75d5bf54a8b1ed419
z2e60a31e489ffd7b32f4dfc47f00997eb53c291038634d5797fa6114f78f0abc4e4c0f2b9c4c9b
z976b14906be137b79e0df298a9d2f65efc73423b09c3c89731183de37b5c2d1dd7f0de2c2588cb
z25ccbee4aa07b04c3a7540fb36ee3a2c6833e9e37027eaa74dab94f443bf9fc4b263f030c4fc39
z9e24592889171c990fed1068d75fc3b88da18012d01042aa5d604f0bba397dd05eec2fd4537be1
z56110da14e3d97434939c70faa66bcca929f88098395dc14061f2afeb67bee278e5e60c8a4ae85
z108ed1248aef730da146e2297d9c41a61dc8ff0e762459d685c1692c09f5072aed80fa00af4e85
z8de8f580642c12f8f8c1e04d5607eb44416062e91efc20a25fd5c0f090b1c0942d89e1fb78bf16
zb6265880e2748bf7ec7dc0856b8b02b745c83317075130b2f38f557781dc25873b4247f9065d3f
z833a980810264b57d6869d2f9c6bb906b11dea920a92b29f73f6810e6f9a49b7065aa59e9aad71
z3763de359085a434882d6ee76a96a037c3ccc7d71ebfbade8c7b331d7e35c06cda52e90eda08ee
z1844f609626885b83ddeca6703ccc660ceed55d805a1a0184a14b450cd18d55c7fee4285a1a47e
z382101bdf05056fe202b4cb3e9b4df5461b69e9db36994182f4ee9bcbfd40d6882f9678a2fecc8
zbf4db809559401712e9a2da26cc318cf3d1780e0d3c545af5a9dc361a4a9c1a82c2f2d1781d1f4
z9ae06cc9333bfa30ee36ab436a8c304f856800c5023664c5138141ed8afcd074cab1558608c4ff
z9cf40a8901c1fbff9c14974e387681edf9e5f47a77148b0b33089c43f765623ff162ca588e0ed9
z25c460f0472dc560c6ada7e25add29e2d1a8ee7588c53690707db7c5467687a56be6de428fe245
z03d1828f4cbbbf39fe922e0bcf4c882de0b490660ba39c1cbe3405d3be739ee088728f44b3c006
z48cf54fb7865c0dd730cd94e0c7acf6bbf640af204d67ad12c8e0cd4bc4e8bf170cefd3ba509c8
zdebf4575dff9ebc1cbae0dab48b196221e10317827826af1afe8de715f05b6b3946955f1fa9860
z8f48cc5285826e080a8e1d952fe6f24d0be6feda82ff618f5fb56ac98105ac46a1b58623bc9a15
z59c905547210ad65964d1e7614c3651262facd124e167550d20e5b0ea04cf5cbdbde4827bdc12b
z3dddb85193ffec1a668b01b9e2a9898c4003e6ac38b55777d2dc6b881d92b66ac46feeb602ad20
z2f3a3d169ea2326926b889b2a368217e0aeaa56098ca908be9fc62f8fa6c9ae797e47059cbc218
za8911c1eeb1ac205195e028d2829d25a4f7569383f4a7fcc345ed5b8990ccb7342ba24571b9cc8
z7ae4857419e719037f6ab12ae374b57b0e67426a1e39ba6a88705b031a6484e29b59dc5446b4d8
z5d6de67a50f03bda0a33694d7ed3ede55d9f200ed9a6aec2e6f3183fdc36849d1e05dddf188fd8
z042d86ac8bf2439b04d37df446b6e368cfdc1b4a6046f85fc2a851f9df265f2d61fe7d52b5b35e
zbef602f375520d05f015fcd97d7a0a012c7f72904db6a5e05741ee94c6cd4fe0fe8757728424da
z6598761a39f6351c5656838e1667d05f3a41b6b67d22e677e9846cb52707cd8518994265d3a0e7
z61f0c6123ee1c08978e42243128e53072bd67f15a6f21c32a69529e3c247ebc2f973eb626adf9d
zed6f2b70ecde60c3b8c75dd6946b9cd6da0185965ebd5aedb86fa82b03f693efc67f4d1c69e424
z46adaeaf9212fe5600015435a48d4bb7fe8fadbcb2b484ceaf56acae1c76503894d8f850e96e9d
za740f56b73a9bf609d152cca052f34678e4261df5bfef3265d78815e35d2a1b3f6381c6dc5f09d
z140ff109f71b0c958dcfabf4c25def1a48d9de5621c09f1a7e2492d674fa8913c65a1eff2498e2
zf4c386d0f40f5b21f024e5b063cb983ed11b71d6a1a113504cac30672974fe351eea63bba969d6
ze4b30688940d2eff6edf34c2875404c420ff324e44d4a83c4b15fc093dd00723f3646eb237f964
z9258a1627f2e4e4ac2b10fb2077cb1133a8f5ec3172d238d9fabe5ff6e6b37f19db19401bf8d26
z82e74f72bb6fe648f88227df747bca659dfd1bbbe9477f1497f2100e73293dc2ff3ddae9292b2e
zc039f8f9e705d267e77cc88bc75794e9eaae4f5610d950142cdc9a9db721efbc20400e215fc5b2
zd645d3d9667c23ab157b24a8cec19cf595487493b02ef9fb6d093d810df8eee0f614e3d9dc86a9
z864a3c5eeef44e5f8b7b936843a88cca2235ee47ff5dc13ca16c7df8f534da177478484bd3c10f
zdc1012472662bcf215ef7a999a052585ffd0552bb5583d57c72d4765b6ab6237954b87bbfbd984
z7ee2a3ac7eed9752361ada79d38630c8eac84909a3d6d4447f7d3e32f986f655b3f998387c9472
z8c733fcce6a95e115855e36f083c2cf9f08710cf6ac66b756dd9864a96b1d4793541d7013a8452
z704c775a0218de44009fac989cbe9f5adc71b2a588eadf5f54356723c5871c56ab260cde77bedf
z53c6c84290cdba027def12d2a7f1bb32a3a87db3890bd76f0b6abd19de8dcb4d6a2c1316f75416
ze479806e6ad6de7268fe2d7521b0346c1e00abbff7868743e52c9d567297e72ea1c4bee8f98e6e
z5cd3243dd17fa3065e1a333df13e140f93b8e6b1938fb6077aca9252d86b97d3dfa40f01172ae5
z89fe6306378c0a79520ddee7730d3d65d0c5ca5afee1a5e74783130572cbd3859133628d474c56
z68f789978ceb5f44e450d64564c9f92a858dba4a6f6601dacf72633a23034e1584c2323ce5f26f
z184501f670da863b18a60f52ffcae7152cbdc29743f6219b1216de7ee5d77ae2c1213e2718c24e
zc6aeaebbbd365db6164d3ebd2f6332ec80158d683eff22ba5a8f1fc5937b6b5c0774c877667a3e
z44e545296f5d2a405150f226d4144e71eabb368d4d6fd99ae58e404167d632103f1e8f8a2934af
z41c52aa49b45844daacbe7bfd87af5b07f2a20aee047bba477efa13dfc943133406babf2f90060
z7c2bc320380e40a494fb04c6759b7f0db7df3dd5695cc1fd1719d174379d16f5883b22bba8e91f
z3ff427305c99131e5aa7c68a1a381750a626dc4df5ba38c3ccb9ad06af4f0e17fb100690cce0cb
z7561324cb384e9d9a91bdbe2b10066757520038b66264fefd19c380433a22f50a5728ceff32199
zf07fd298bd89970b6a4d940283e451327ae3881b87b2d0357f169baa0adb29a686505b70ebc3c5
z69615794bd1e254a41bec305a9679556ae1623b838868c2cd54113536d2d12f4583fc714e08271
zcf2893f50cca6aa8c15b63238604581ba744d57a8d26d9c4c724cb3827d264240f5ed8c34d0621
zbfbe2c757e40cc9dd066499fd0e7e17d2108bed370b53d56547915bac18ff9f14a3c66b6800f20
zf306f4778aaf99c1268310c5e533e71fc22da07580d4b9e6f7b0c38d97e718251dbc5e6fd8b610
zb82e0074fb19d0ab0cbbad4bc7eb2185c0d83cd934e6113311249082d8fd9d88615449b9fb17e2
zd1a6c795e8c8555cd44eb7282c229241f61cc7995c54d3bfcf73938501f4dfb06ef9bd2c1407a0
z12cc25d4dbd134019924b4b2af78bfd0c212e1d1261ba74440b1312ca132677df0c8adbb40d9d5
z6e1cc76cc0b962cec2a1e14d7fe34d5582b8a3457b68c1ac066f82ac780dced54d2aa515a4b63b
zea22d2e01726d656fb72579048495dfbb83e944f11e9a5d125fbecec149ab040839ad91529e4a1
z3bbec2c6a5feb42ac6619c79dd623a056ddc16b0a7d652ba19a7217db151da52daeb92ff086d2e
z14bf915d6c6a9ba47c458750da15e2dd8c3cf4184b5921138b9da6e55af082b376991c7f5059d8
zad0595b384afa9ae28406b9197aad2e30c4391abe6c2448e460366104ce101cf65d6d570ef80ef
z5d6cce9baf5b0191190e0e727a37336d3fa619300937281dfcee947e5a33a886dbfe9245bd18d4
zf9da503a2fab0c08ad44f067f9fa7f1f90008c09301c5bcb4a92c3c2ca7dd1e0ce0e4b8c5f5d3b
z9d1f3d996bf5e98110632ea0ef7554fb101070b8580464e18b6bdf48e0386a7b7a40e626941228
z2c0cef463032d87d7c063cf8bb280018a2bc38424d7ec0332ad585c9ed0f905ca4177c4c158d3d
z33d836102a0bc8f9c5fefaa99b565de47f04f9c97ebc5bc04199928b8f4d7f39819e252c870e7a
z9217f4b7c387b42cccf000939e6b00a5009066c314fccfbfba359f8a0ffbf6ff229fe183ab6b62
z0aa232db11a89183de5cd4a5e8764a83786d9246a563845a5d51920abeb4ff00a0cc7c84cc44fb
z3896fa6a65298c0261cfae11abaa02e240a8458eeb086ede2d8f3349949ad3f4e708b2d483f815
z60118443936c15382d9ba468a253f36c3f5ed35be318f5777d90104007fc66edcd2f0499e1f4ac
z6316da96f40f48631931ec939bd0a49bedf4f10c39876496bb2e6dd7171c20607703b9b53e63fa
z335ae5b720159a5ff751b57bd6dfe7c09b30e65c430396a1b5bee50ba68b20dac6c00a499349e5
z2117e52477b3cd8fd19652c4c2df2eac6e69b2f517ccb5559dca83458119d1c5529173dbe3c245
zed9cfd7803f2ea5957549077281aedf9f1a2519d0803010e5640f1d6165d81495e2d235d505649
zdce67f1fa40925a7bf3a9f1fdfe75eb548ba24da5ee8c78b12b06830a8351f7694295449097f50
z51adf34bb3599e329ff428067252b7e7c32936e970959b71867c32010aafe46a4c22f4912caec4
z91549bd7aa55fc7b53d8e3876ad03c793bf51e8ce706d40c1bab298904b1f042244b9446e7add3
z2d95ec7f0560aec57992f72dace0a47df9601cfaacc2dc4b1cc3c4af44d2f8be0057d0a8085e99
z5395d50b1d3003b2aede59e58f843c1c42d68038de2ae26507677b7cbbd18b8edb0de8d4b64c64
z55fbae51928a3fd952c11067c43fe1765e23c724a5920f70b8ec6383c950672153b90213336998
z47185dada3acdbb6ceead3615de35109296203422cc6f7627b7332df533c61184c74f79f193c13
zb74b8c227c6b0dec4eb251be60be8383645ed6e573c35bfc9b9d5bdbea457a3aeb733a637465a9
z24cc94fcd699b696a346c9444153df5f3678be89e5670fde9fafba8f5d97732af0ca787287d4c4
z5494cd7d4d3ec6dc9e6115477f31571f16591aacc1611f16fa7fec73a4ef43f7b1b177aff0914b
ze74d32ce2a86b0ed54a85b243a29f3e48f0ea21c4a5687a1b970259ec355077e1884e7798f01b0
z3aec0872d2302d03c0768c7c993dafe5065773b23e1cebbd454a44a35d2adc0f2adc2b6d31d9e7
z65982bb478dea46dd0c97397110115276b50df3fe9837b792a15897b5c64c9f94b9ad2bee2f9ab
zcca402a7919573b4e7e748723c38d0725660e0f48e806b028d9c987f12b8be8d83091b512180f6
z09b203fa3fb4ab1facb0dd59361489bf3c14c65b4f40678edfd290fe4b0f8e624c4f32a866192b
z0d9bb85c56d6205dda94a73d002923c2388b704f607b04943a66823ac7f011a93b3712ac8de401
z25ff80a69adb195619a9db995cedbe24504f3f90c27f36d82361a10fc3570f562d4511ee4507ad
ze5bb386f4e80e42391e58779d2ae6549b4a27d8292364dc62fe024820b76b486c1f99df7db16c9
z226e9cfc1a59d67ec9de8deaa4fc3e64a3caacc0cfb06ee348c4e4110dc91700deed891fa8d88f
z13102f5b68460ee1f0d492fdbea990d638e98341c2dd69d86289c441147a19ef83d8f1cc351e80
z999f5c2cd58aa98772f28b3f05ae89e922344d69bab69165a0801c898909b78cb04a37227519cc
z41997b5ac9e5fa57ba39009fd37629b21495d21adddd2b44c0f9b1bc694ca319571183a77a1724
zddd7cec0683159b3073c6933046286064fb99f72de1d6732847ed1a2db345bb5a7b8807e21c75e
zb7b222e697c6f9fa72aad379fabb03a680c03a5886b0bf9eabb041aebe17f18c8cd5c38385d202
z490f3970cdc7021a66932f1e23c0dac8917d3a0b1405f2de274bb958966b1b986840867a06985a
zdb3052e872eaa36cc151890418b0943eb0ffb99e3bcbaeda1b298372fe59760828c745145f4217
zc7b57730a909283117f4fd87a532cec46fca0bd09cf5b31122987c1079e83b286ab0f51223677c
z554e73bbd13a357ce3d1971261b1415a8d4a983a37367bd48a25e5afcd685bd9ef4be66ecf76e1
z250122f1237b6617cc329320de4dfe2acd2f78ad7f883d0fc3f000524bdda4549d6d8603946323
z9c85c8f59c328e6516e684a38d0de1b7d0ea370a00cddc503ac95a218c525b27975b1600d19561
zccebe490a6a86afada9a84bbbe06146f506dd5903a98aef4bb578ca33e3c51094519e9290eee39
z5b9ba4dc9f1929e77f910a7d893f9e5a96037de8f198b55f742d41ab1dcf72b863264a6436c549
z9b820b37ced5ca2a8db273a6d5b0e2d9ce0204018d6653b9ef21bef7a5059ebf412dcd9e7f1680
zb616c9533c80a16fc8eff99073e077b67445f4681aff30c1e31e65945815e5c5a7daba193aa31f
z9b511f0fe1037be017bc57e3f00ea4371490079c236c7f1adf9c59a1cb5e0e7c51a51dd8680583
zb8eeef615f422741a5b5576fb1e8f277e457b40b6124341406c10c148739edd35954f6273fbaea
z3a2a12f216abf1fdbc11c5a00c171c938665b9426f959ecb6be2a9d07164ca5fc879c8b8fe981c
z8f9433257b23c94f3b2335f1307a974a21c2f564d6b00280a260c03f6a16482b5cee1f5b9ae2e2
z7290a561efae0fade06057751aa934578606c2360c0dcc2ad3b8423b4191dbacbd3cf7966cfc51
z5772da48c5b37747308bac1db2cb9ed819038f831a3f53044aea58a13d0c00205b15e8a772d19d
zf5d533ef7f4fba70e6d1e0883c2ef1f801fed8e570b186d84f550bef18a69437a530db75effa62
z57b3e456bc9805b736cedb8e1bc39aa05a781e75384f68c52bcf9f204cfadfe9b4ccd062cf7194
zd70bc9ef68301f4caea717dc86ca0716234711c4f2ede426357c567b5b2776f3fdda9f5d467a9f
z57e5e8fd00523ae7385661cf6bea923fa64b8a209b922c2942c16948394ee46a376220bda1949a
zad6594292e13ec5db794701cdac2017359854406d7de3987a5972beb20bb5cb2e88716794ef31e
z058e213debe9315b200492b5cae8f0178506fe3e628891a7e5c76d05ad29ebaabe6b9b3abec942
z925a4caf437d34b036ac97dbaa14879a159a9b3e1822d339dc395c110ea592e6823c28b144bf04
zc7924aa4b3fc157cc9ce1f33a70e93a3a0b8037662764ac6587947eff3a19c355eeef4f22adefb
z9eae99aeb8622226742392f385a80b41857a21a563c58f736fe7286277a99ee084b9028b3dfc5f
z10db05d283251b51f7b4f32fc9990ad3fe60300cbac30ebe39d8e748d02b4625b7abc1d9341803
z8c0d145cb3f1c068157cea2237f40b2f786b2ffcaf5a5e4ecb811f595b7bd7314c0f1a2bb27de7
z84ee07dec1c8998c241d7d4963368e2df42c1c57c400b44c5519c5f01e1ffbdda37f81e96523b6
z3d02d0821341f521265a8ed658f22af9179e299213f6750a4516fe64c091bfe466409ea50bf5f8
z1667ef5399c62f7999871426c1b0d05da47980e6f8507286cd32197a5f422f73087d8d0a714325
zd3af9dedfca25991a682b5d5a102599ab0e4fcd45fe51e45927be2033c83d73d34481c7d5fe1db
z4d7323086f64e82f0387cc391f30e48f5811bc667cfb14efac6485216155b22eb9e872cb5fbef8
z1ea35682dca741a7abe71f8a4d157067afdf8db41f920eb7b6c0b108297c5081db058fe52e8592
z188b741de46afe2474032078b56f86621e91907d990dfc6ccaae629942e2697f7c1f6e953d995e
z1d3f3dfd0b1bed42cb1579f9813e7a69830d5ddfd3dbf0b18232027e22bcb41cbc5db5d78b96b4
z232fb7aa238f965097f90ebb2630a82fdd399f51ddf97490fe63bacbfb824b6ea0d45c309deb49
ze67b9ed61ffb823719c4f004dd3611988f4348beda992721f2f0222182406ff0e08d05db7286fb
z71070c638fcb46f018219ed91b6ec8d4c5169f01d77dda4bf7b048a88c22d632eb3f5ff43435b4
z36e0a9f56f241f9d9619e41b921a5d1fb46e55f16a6fd1b9321c9ce3500bd622750e44c0f79366
z6d49c410afdd59e08a90529ad8462dcafd620fca9480d3aa52fe5a22a502ee314d3cc87ddffb8e
z986aaeb134e6c2a6dec068424a2b35e3d39e7447902e42446f183ab095b9721d02c51a3afb540e
z68af0845780fd516de03265a07515a7c0f9491b00459f802a25e32fb8c0ec3e478ace96dc26d97
z030f75686d98b7b11206d1dc8d4487fa4b99a855ced78c96cd0394f29491bbe294a5d822461780
ze46b4bec1f11e71ff17dba8b6df5e3a718dba4f1f44dcecc3f964c0f4d8dc8699b1ff3a62a5610
ze336e72fe0d20089bcdf025940bbd091af6f95aa829eda70e64c646b1f08ceb4f2b1c8c23a34cc
zb14d1f037fffafcf306c97deb9c140059628b783229eb88ae47ee893840a63b7503b4d11632af0
z686b09bc00460628f76dc29504269f84e21b1c9db3d62b67546b667d5f9da08f5a1009d1327cec
z9b638e63d394a7c984b6f4a43e8b08a5af7df11ef68b06ae770c75dcfd6e77446a48975fcb308e
z31fae0a289a2c900f9394ad92c79cd593b34d481c2063b767980f40fe36919cd8113a3238378f3
z4d80681a145258f3ced56ab422908e943a8c7f59e0bae2f15a38d63e6cfc4fdfd0e2d606d6a535
zfafd7af4023ffb863a02b06dff47e9e71a630365cb0dcfb8f6fed6d223df193d0f7eed1d5eeb51
zfac92ae776e33390afe72b5b9babf6df3d5e21aa971deeda8022875d50d921bbdabdee586bf43d
zc0b8d746f53aef86a0c5a7c1f374a9953e2b7714f34ca820a662ec78bec66ed73379106a57e0fe
z4f9562f31684e6490865e4ace6aba6b8cd4965213fbc62f20efae8ac317801c14868653f05118d
z59dee431df6878a3a22a92b4e4f57fd1ed2f38be82d3e5335f33722a72012923b20daa182ab726
z88803f1f9f1918acd5ca2e650f9f532c3f5e38f48fa447d1545d114e3030fcdf5b886a8beac64f
z21442f9f36bd7dc6f227688c89250e7a0e64e74c3c508893681cfdce92147f27451073e89494cd
z5598ed37aa6fe5f70641484e4e92d97a1e2243ccf2c77942d730ab12730b1e6c36a375b792e678
zcfbc8889eac5ba8c83eaa2f2376946b06f3aa8a30f3f92c77bf05183f86944b5114ad0619627f3
z9cb06ef51ab888c8e7fece0cad70d85d369a04668bae101c6d38da743720588674ee3e2a675577
ze8e72f4b47ee02eed4ac6f387bcae2d99b25e68b75a3f0cad342f39208520bca8f7352e8086526
z3e37a5086b355f20ba969c4b3678f11fdcf7b8e1d291c6b5ca27a008af7e0ba7d711d6595ef1d6
ze4a25407a27fc0cfcf69ffe1cd775174366b5215d94116ff1e6b32c2aacbc69be7dc4a11caebb4
z6e3f0b50f651926550ea76b1c4b6f6b97ad840d1fe58f7152ff62aed52a06f63b727dba101c50b
z77e85494f3268eea54f0734ea698689da24f9c7b73b82951bd8df0b4389492779822e7fafe294a
z1923c812c10234d8d580b6a786cedbbb98e880f6beaaf7f12b369d02744e0846875624b36786bd
zc4f569bbc8ccdf9df2170e5de9087f9bde51e745070719f936d3958dfdc30d087295837aad17f3
z25ba7ed67c414bc3f72c9dea06b32e03004b5cd67b7a4a36868a666c644217b22dd308a863e5cb
z663a2108ba6870ce6b7da4e60fd37ec85e2e884afdd4d6ddc0ab2750d7259111d74a2ed6127ca5
zcdb4883372d5f31829f0ec6dd83b4c73d5caf412080df04aae9886164d086e8c2ff94eb1aac47c
z557c8e62ee1dc2910d7aa428b3259bd03b2b5088fc65f2bed9dfc3ce1172d7c180373b66ceecd7
z27ea4a29c003c9ef1efe172083b9e45eb63bb6de427e555b0a3b5d6cba90e641e7f359b12c0b0d
z50a47d2ae39972a347256121bfe57984e21dfd04c2a12dc356595c2929d3179491825916e8e61b
zb06acb152a7daf55397f7c6ac83211037e2ca0de426f3f9ab87e6390ba552d742b9a4add2c7b43
zff8ee708eaba8b450fdf03c3b31d44c9ac73efcd6ac21dcb4cca8ed792ba3bd24f83bac8711a08
z47cb7c7913d68d0c0c128b20359b5b74a773dd618723029b4f441e5b30f1addfc6a1137fd0684d
z1c300eb55f65d379c5a1cfc6e210505ae7cb901c112afa2e7eaabc1aed86ad68acc3b62d623ff1
zb4728b68a4284f7d7eb4f585109c85ac49208dc031737a097502112e69c03e5d2cf34e90a3b012
z57eadaf0ded2b826af8e749e95867e77b9e3aa6395ef3562adbd69a2a59bcedb24bc46380890c8
zed91931408a4697fd5916a35b60471288fb90a71e01d19a1623788b0e9a3f4da0b540c3b21fbcc
zd9e1309a09328db45a167cab38e6768c98f044c8d7dc2ae73ba5bdd7ea3902f83bbdbf7a909cb8
z5a016d14725749e48a184682baed47c6b0e97a0b5b5c7459984a7a0705bd3d6129c9df40c97f7c
z103ba747959cce40d81751a6b5c9d7431ed9dd8457ad32013e1c2658b242a16df68bd5ce398191
zcde252a18fe8ce7135a097adffd4854b66bbd0a05b9517a57e4bdca23e0971b9834e8738f415d6
z2df6dd11ed1e8e1e912835b6c7dae35941ad3da7175840ff985a06584170154730783c72f0b97b
z482398e6bd25ec44ea07ca06e73c7ac355c1382a6ea151cf9e1a574d67337ec59bf0663ed04d35
z5ba9ea5b71c3183d095724a119e5bac33933726aac0c7980c16dca6a1342f27aa718eac425755a
zfbdd58608c17468ad097252838b2aa0e8510a58d2ec13d25ef914bb58e5ade49d560ea26481bd4
z08dfb44de06fbb9b23400851f76851d2bd9e97ed6f7d00c66b687779686b801b55e1440fea0652
z19a82a9891bb401d0edba2eef22f67dfe6c60759afa2005d3a9b1dbbfe0e55043e24d6f525ad21
z0dac1cf8d8abb99168fd116add31c85a2a0844b6e39acc01189be10889349171bc6549a700ae06
zba9f15e5cab33d088d25976278769d971665609282785e8f4789ea35f58f7c8f7e8444ea08c2bf
z28f408949c15f5752070d55f28a95d2957ae8a24cb010c65377b19065ad4ddee4745c015e56600
z9b8dd8b7462c41c0af3672b1d121b1d8ba148749c75a8becde59db6f6f2f619f6f2c6203f678e1
z8cab8bcc47b5f7c283c7d70a8b1e7988b6b4f6c76f5e9b47300c64c02175f58700aba5ffc3a498
zd1cc3877fa2f85417672c0bfca853c0b845f8673b42b073ff5d7bd009e8bf3d82cd0a075afda78
zb5d776a85cfdd8620ddc3752066995c38bdbb7dd1d0f5d8256f96b3093f4f7fdfcdebf053ad26f
z4c5bf22e410c69d4b379fca2d0e50f3a094db8b460f93f60bc04b02523c3c19672b47ff52549de
z62e16392d0fd18a6f3a5ef2796d2f9cb47068edfba21218e8fa226509f50fc8d38a2ab74261683
z41059966ec8421f60675e622b9a46cda58c0c1eacedaae81d3424bb13f9fc9c481ff689e2d5ae5
zdfe20a2cf854194bd8b89519181f4f178bce7dddcfa16a6d9ef2cebc9b95375afd14632427ff43
zba19289c181ec8148c353318710d7a85bd7172539b73bbeda52e22e766ad5711e427bf9237849d
zeb68a3a251c3aaa9ef097827cd365cf2048b09f916b58cec0bbe7241e01edb085afca3370e9b97
z551fbd82c44324c9471a66029a64c528a3472ea5cb89d0ef1cb9bd00729e5419bc1f7331eb9c93
zc4aa0dc98c7a29c0b99fd939c674154fd2b602ced2093a373786131ab2c71d697b49324357b85a
z6eecab6f82d1eebc4cb5b58fb77e3949c489df63b6dee51cdd005689025d5137128b15ebfd5dde
z263ad46d3bc238516fb30497363cc7f24f89f12c5709962cf8020cb77fc02c07d66315f6ac8d19
zbe6dde9282138af43e9f1e16ea8ab4cfbdd14c727c11abe2d5a9fb14ab1807ee249e67dac00858
z782eb548fc543cb7254a85120e47940e69112e1e6581cdc29fc696486ca67000007a25ede491c8
zbee936d22a2e8090f8beb5ccac4c8d822555bca90847216f285ba90626c9e908cd95b009ed0ca2
z487abce6f9342db8867d603ceefce46874bfcc157e8303b2d729e3cf5a01c0738ab244264d33dc
zae695ed95e7a6870c77c862b492eb0fd0e7029ac367753a8c9a14913edd6397d65c7420e00058b
ze40fc6a9e1cd67df554da9495a09cad48ef9a8b32923d9b107cc9702492cbc4772292121cba65b
z072e8998aa2150f0d173f40393f4170774b6c5d422594226a5b30d13a7cb0f572279c83e43777b
zc3c7f6f6673f9b83e5ec095533cd7bbd5b0957e245d7430c2ffe88016b7ebf9b49f65b3d93deb2
zc3eb5fca535cbf52ca9113c5b4145ed2f4b9eaa2397a800034e479dae50f386520866cd8da795a
z383afc156c5adb298c705c42f12c4ea0da68cbc5fdb0e35bada57bbd4650867cf02d0b1924c8f4
z6f989b8dbc4c9bb1bb038df1bf19737daf03859aa6f6699f300cce5b0e199a2515b56817b7e3d6
z4ad6951af42c1c5b9373f5f46f26607d5a26a21dd02d02f4b1f8cf8d62f888d9783c53a6d88490
zc8201b5adb7260100a530c8d9f35ccbfb5c8a820b76d2ce3e05693d2ffd4853696fc3752aaf67b
ze421be3b4133df30edf7ad7e68fe2b9f15c78001adb081cf95d1cab09e0cdf675f3bc287fdc892
zf21a41b86fc49087125fcc987202b21f8c206ac4b27256e81f5b445249f720fe16ccc0df1eedca
z5079557cc87a4dda02b1e3e7a16cfd586e6715141eaf55049393f16acdf4f67f5f4999438e27cb
z4a42f54d6b4bc44f7a3867ffa7f1a83bbb46c5a5d379593fd9c5cdba27a131925c52f7e6160902
zbcc00eba7c83b164c6cfdc80a41fc49c2779380f8835bb81eeed4e624425a04cbc4923beeac86c
zae1c56a64fe78e8069068428bdda347c998e06ece56a8d4ad8143497aee5fd9475f7854014b2b7
z6b6fcfe3233ae543bca655128ead9a1f289c650988ffa29c532f99eafe7decdad34f10f18b2526
ze6b0606667016b6a9a86256b64fb26e1677b310455128691d4c77b56af7eebef04098e6b8b5acc
zd6667adf4021d8fc5d70cc9a70512601fc0e7ed8437ae5d5548b63e721944f3ebc2794497f6d49
z7fa163276f32257a69c3172851ff6b7efb7e67b947a53ab75eb1e972c5c8acfc0dd59f83f2d8eb
z671ac20c28d4354b2e7e100da46d27f42c898de2bf2a4cb9c22cb0d2a63f70497c8e790c85f27b
z78da9d85ca841f6a7c51ba4ad9e4099abc3f1ba16392f6b4f69d12fc1afa86b3ef525dd2ddd25b
zd3cc370591bd6eabb522ebeb7c79c69099cab223d1d54af8670a916a85dfac1cd0cfff1f7152e1
z801c858476b712728fdb804e0251e7e73401d2f88a57cd20de7ef5ffebf5c59f619e8a7b69908c
zcfe93f6f60a462e1f53037a10391d25bf04fa847061051c62e594e62d7ec77026832acf14f4b19
z0742a1e6fd936e70fda137b335096948b9928bd629f35854f70bd0deb32948cae6fccf39ddb53c
ze915a8620b745e824867983c5ba16c195a5455e679d225782448ebac20d48ff2dc5e8a89d53359
z7463268f41de8a7574d37f658ea1e6df650688dedf3b019bce3b5a9a980b104731114726d9bd7b
zdbe4df58a5737c12be7866e583ea9533a8b89428dff160b13f66ed2e960663e92077101c379d88
z6384747ba15be997c234cf8e4a317345915cf1c056c20c7bc7aba513f6031817b0d67792650ef4
za5d48e740db669bf8dbb16fb32ce3f60b3b262b559738f4410693db9a31a29fce360d43e402a58
z36f3adeb89d8aeb94b9b697c25e6371bffd6b757ec09369c30642e998a88e83e310b0049a905ab
z570328a2e65c4e1f61b9037e190aa037f3a91e9f8b80aa51404495d93cef5f788fbb75f9e5a81e
z59d1f690b8c863b3be7aa7740db6334da973e6b6ec7c4a63e891d4d593d340cc77cb9d916b2543
z8f545449dc377426aaf8905ab04f00e79d3f32464289c20f3e7c9a8ba51d5e20f4b45187017e14
z5888b8cab3ffa85a267be32ca549048b06da321a9f9ed24fa3e663eb1133f967d0ac50039178e2
z0adb1f648b0702576549c82d4c09d46bef95fa9a01c67dfd3e90088a28d4b30c2f90ab3474b08e
z6eb79749657311d14c2873e61aaefcc656994cc625599e589c0dcd95825a6f18dddb910a60941d
zed91037754dcc3143e5249c580b62bc628e3201287864dbcc0fea63cb192bedc65524da74b77db
z84628b0bccb91cd2658d451a7128f905d08eed31e6a1a28e01dadcba168f64d0b9083d3d5249a9
z5ce574ca4a3f3b0aa662b29feb521caa7cd17e26e54229ecf437fd2f043bf2032d887d54f5ff14
zc48a10273420c5ce77e18c8012806e594dd678413fb4ccac687028c25d1c3a9778a6ffafe6be1a
z373c50b4a5d1144b0fd3b50fb8266b7b3f5d4d37931f432e504b913dc1c94e3c69262417af6d25
z0b3ac116b8a23bf852214a7f04a40813f45dd54eb632b99cd2662324cd71e23e94b900bf66e370
zd8e8ece070d598299c602946217b072c27ae0e40f5b61eac22c6df963e61568152df5f19e43dfa
z5a56b22e27fa8a435a2a36521663dcc3f16913d2913009f4db3c116ecf50894cbbbf1a6a32384c
z90ea6963b2cfd32d7ab977e95d91fb1c0d27514bc792eda7fbd8ff5ed39cb40f15b16e081cc523
z1f14a3bccc3bd8099c5234b81f2bd1df86db9a3ed074d3d655255d116525a538ccc86599a3f1ab
z9ff286dc22769144abb1bc71164ebe5d7a1216b4904b24f745c33b9762e177e65e434c2283a09e
zd4d3c7abb175e0d3b934b251a39417e63bc5b2c0c82195d77b876757757bc5a6b04ecfd17faa31
zb0c3db92a5080c1563c33488bbea7d83f10c211a8077f3010ac45150aa5c113585a176024c80d2
zc1884d8e198a412067989d13a8024cc8cefec2bb9d3bb8ad698b26ef4bb7887a3af12915812269
z950001d42ad42b91467748a65728392b48dcaa4926da43a840fdfa7275ff514959cd241eb87be1
z260f22c3faebb096fbf11ce0b0b1813c33bb488778db0131bd1c5b0c69f09967c5a4f87d145895
zce13b24834b84f1c54283fdac0724e2be33b25e313a426af53f941f06f222ca7d26db52e6e4196
z2b729c0348857c1fc0f3540e1b48650c9af871431f4a8d6595a55c7e1ff41bca000952bf0479fe
z289f413a8a16bc9fa1e32587bb801e8588eb9481b83b5abf49b0722b5f4817d81e3477d902d5d4
z721d9518b0bc15b55beb00d38ca3bff1a15a50f2dd56446442e19af857e204890880b47c2f71b5
z1e11cfbcd66ccea7fd305c6d7bd7ea21b5958e01cd77128c15b6d56109860c5599ebec16d0e718
ze216ed663641dbbc57b33b31c558611c16e4589c7b89bde34af7ad7e6c0b2d711b2c0b52670fb2
z201b7e13539ecf41655ccf8432caa0f1175b995d8ef3bbfc2b63e71d46033be49add7578ef9738
zc719c39ff3a0103251652ffb3050273edab8e2eb77b9d288a7a7f2a90d2ee53e66ac2c9424abb9
z9533234633cd6f974fe90eb0d077200ae76a016e09ffcfe4eda630252c92961d085ddb37e68968
za9c98ab0ea19fd87c329d926df2c034ac9eaab0f1dac918c94d69a6f3eb345f7ea0815c3a00cb7
z38acc1fdd18fade469d03bb6f4ba0d649eb1a598f72788ccfce061a53d125a76926d0e19ba353b
z5f6b0576c42cd458e15a6a6046c6a1a1d8f79feb560f06a89bf76cc3dd6a1d12ba3eed22e1aaa5
zbd4b7a5dc1931cb076acc7c70ed61c380599ecac7a3d15e4353ae6853c1bd9b49d06515cf94d71
z9e0c0c523918a2699ffd3476aa0fbd461804dfee8437e2b503b9f3a0d9b8b0df97e19fd3c27fa3
zf627fb5e21fd7a4c77e0e63ffc3f9c0ef746695a4bb0d42b0b87c8ce9478265490a83b79ffa7a5
z5e18854970c9441d9fd7f7b4a1225d5e526aa646427885f6d425516921c4b9b2417a7a00f5daf9
zb52cb40bf37cefeb34cceccf409afdca0567d3199c68b98e38ddd508d4687ebed8e021196e141b
zac2b08314c3ba6e07e472bf0c6bcdc57b16674f1206d6601e22f70d47e483fa21fb6ab401142de
z6d0d0e4962fa44762cb7c065e6e1131ac61012bb8b81aad94127d403b43dad1d96fab3b430f56b
zf0568bf90122907707b57fbc76994dd6c5178e8198a529ee18c548ae5be8fce35623fc90e22e28
zaf8d7d8b7e624c3cb449594942782ab1b2a5a9a880b0b175948f8d575383b222587cbcea99c402
z803beb0b8b8faf19bbcec64a59ebb4cce0b77282b17b97bc4f5c84fb0db1d528def400173b14ae
z9cab57e0d3c223b9540a086243f6062ee8a231633afcbe6f25c9ec5cbbac94d14cf875419b364c
z89e932d7a6c6710e3b3fa05b41f4e27ac2554a078317419037715aec0b66e890445e5f4fa49561
z295252c02d77e41d9c5c7ca7feef288630e494c7026438113c232adf0efbd1cdabb01b39c7c9d8
za7e1e63d9afed8bf8bb03aa95cf5abdf82b5d75e66175412feeb75946fe72fcad82ba95e1de4c4
zae5e07e3b79fcb7450720e99e60a8190a614cd0ed22586ba896f7044b0e8b6da8586bd9f62a36f
zd26dc6e24294d238633319b912e101093eaf77c57af2ece420251597bf95826ccbb35810bb2d24
z5b6999e2448e5a239cc3b7e1219127a2d82131eabc934efab558349639f490ee82ea7ec8e282af
zab231a6f3891cf12cb9681668b3df21033ed8c194ddb16d9345a39cfb7c9891433a9dc3bfcb226
zeb076cf83bf3f9522b40a4f6cbb6a0d047c57ac939a8bf890a3dc9b85d698d8925fe1e79871cfa
z564a5a571b1632f9fba76c534c1790265111afbb3eef2bf86d47f9ce55e3b1c3700d27bfc60480
zaa4fb1ebcb766cd5fac680cf238f342a788fa4013211726ea8ee0ed6db8f3d190c66ac90802730
z7ffacce23de39eacef0e18a889fb0ffcc8e668e75ab18d41e849b23b613be7bde564739b159cb7
z7edb3eb5c298bdae005fa34b3d786cec5abc4fe3d28730d889a0d796268ba418e01edd58d082f1
z142bc08b1389173494ecfd83b9d0165292415ec163102bf5056d109ac3b99595d801540520799e
z97257ea6d145f06ee2f983b79780dbdb120081aa2fbdf49e66b2a9b9e07a35e0418889cab06a7c
ze8853542c10e6275c7d26c9300777100fbb77066a74ea46429217a6c9d82a9127c11d8b9de1001
z41c8bba6291cefce2586a66ff7a426a56b518e1b881fba62ec0b44c14342fac8fbe0f55c670f6d
zfd0fb533faf4146cf5254b8392558791c6b2112e2e67993c5cc6d70f14eaf0ebb288e094156d29
za7cb1134c70cd3eede426b6b0c2ffaddcb4fc9e5f0e3fcccba1fc71ee7e29040d3dde2abaf45e9
ze5e38867a7a65defd994f1a8b2fc1be9abffc596e272f846d3ecc57b46036220a5c05da2531ba1
zd545f5ef577e60250d496590c0612454a2d4fed4f5b60a61a3f73a03508bd60a8592b867745a4c
z5cbf337f95e3d1b748b8882546d46e6f754316b093dc22737bd527a3ed0b7c914ae212685801e0
zcb6c8d9ed5ee4cac6a1f69158113d253926d9e6b581163e30626145e8c98d529c0b8f604437e42
z6cd09bc8479f3a0226b8a36f090aa4eee7c443199ac1d3be0d3ecb08c010d0201b9aad053497a7
z5ec02adfb1901ee460d889b3af2232c550b23278a1fcfb3e4de5f70b8c40c9f3ea3a8b68293ac3
z28b14deec32155e40bac5a79bd0ebdf52bfba90e66030c1aa7b917524ee1529fa272baf141f335
z5699c556a37458963c17640505dc66f634567e347d6061b8eb9b3c7db8bc4fc253049b5002a14f
z4bad2ec6628d922ab4d6471c35511dea8bc5942aa6a3408fbd25be78928dca5dcc884f71827519
zbb1483801b46bb4873700027dc02bf0da811cc4ee7462ba2294928c286199a58a5520fa483d076
z3500c712b27b3181ccd140aa3a3f29c3ad119ee1f3ead65114a77ff4a30098c1fd5de601b6f602
z43476f980690cb56c61f16803ca9de09f675a1545882e82b6023b28c3f57e81917cb79559f3c96
zf421d4bd22a5f4cdab8a27a92b4f1f45c0d8532b1715cde3dcd4b1b10ae87909cee0e03b574636
zf56b7845274935c24c30cf611f18c2bcd70848843a64d38edd41f9b214b08907a5e3f0e3b6132d
zb5c71dd297537289300bd4f7c3689b2d9a2d9f535a782af902b856958a80927d0cb571786ee348
zb2da2895ebd23445737f4d273a0dec587f0b0ee6d5cb59289db9e1a26dfdb14fa984c9b9ac4684
z18e1855840d4336e5ddf4fcbc29f2ba25cfe2969912e94f4abea529b38ba063d13474af41ca717
z86d97877c4c9e42c73a47ef7cf67aea2e812a79f5f54ee280a090687bc945608b00621f5f5e0dc
zdd3fa93f7b517f32e371e81cc62ffbaa6c37621c6b8033a81b534466a827cf3ee7a9074255448a
z115b0724aeaa7f168eb51f37a024d97eb0ea15bc64fa2eaa1ade8adfef40982770c949ca1d21fc
z86d442b48e876e6fb90713ce0175389b2f824290addf3b8b9fed33d5c97adc975a985e3a227060
zd4ab1836996449ea402cddc36bac63fc3d1bd07d052348b951c7d676443aeeecca6a9c2aa0da14
z5ba7765e9705c85f3145c446ca3755cb4bf6443e6560baaf09ed2e5697889e8871fddfc6eddce2
zbf5b99a4100328a6f5ba87b5c4aa260e35d2a4c713369020b92aa5468d999338aed7ce08d1b419
zeb178218b4b8126b2bace164b6ed767f95dc209ef14ee2deb85f09fdcc181a6d317ee03ec04286
zc00c9662525432a30ed20a55691c1185f25a0d02a1031b51cdbec8507e1ae681fdd1e635dee4fe
z92b24ad0a54feb53bb8b18814563e7311428ccde36ae5f27b52d0a0d07390725d33b426de4d079
z7b9a55ddc50af28feeb2f0988fd428cce6838eeed968b7f6d5a68478d73dd60f9956d48ba6c968
z7a5ef2da4bd8374cf99f0b74ddb558734a06aea47c86855602cf73040d3db9102478dd0942ed00
zb9ff260182d115907c2a08421dba21203fbb0548c790996f622d288ae62d84bbd3a36e61edf511
za47a55840dcbf0e33b6cfb5fc859a0c91a3f16274022214d487639acdcd860493727ec73814aca
z1cabf2786021e08a35f2fb63600bd9d169d3a88c7c5f0094800ec058c009a8e64ba91f22ec4eb9
z379b1d570dd970ae9476db390f341f181c0fa5fa67705db1de67919d87c30de4535da8f5ed25b1
z7080b6f47c6742efd91ba39b5f18faf9a9f7e603ec510986322ac967586d3b25580e5de1fdb01a
z4e9745189bbe5247149f97bdbb586db738e1d4af49750819fe27cfb631ba58a6441f0b9e28baee
z14da2e3f93462cfea9b7609530dabfac7e407f0f7d5bdf189088a2b52f6a1d1014b3e1c0b25ba2
z7e357def9474b709e513c6ef8f743b57691f629dc3a4307cd25f74ed94fca0fc319539ad430c30
zcbc530c1a1e43f6f376cf6597b415052e5a94ff28e7503aa5d563a84f99c85299dbf9888993b78
z4e55b48415a6c8024f64ca4fbd436628c742d896db1ae299778e92a97ff283f88275e52b1f8c3b
z4fa0e9de0e83ba12ce88d052e2a8eaf5c10d0f93e0fdefb0b14b84113f27c24b455b417d9a618e
z3a513675e4784c2480e30e0aeccfe6801f815b137b9488ff3cdd3b51e74e8c3686449e7c26defe
zfeec162941c0a9a17c1f63715ecec879f3527133877bf8ca1e849512dad3617805b7ba014051b6
z08089d80d533699140daff6655cce5684a6493c4ba2d96d42d3a038d465c10552212c6935df056
z210d37eebfd9aef403928fe79e8e66bbb89e10b0d27ac8888ee24763e7b92ff118b0aa08d428e0
z1918dca5b161351117aac009afcc3b5d8108828da13b00f4f572bdb80923f2dbcea1f1071e150e
z5587160f9e9d95c47eb67332d4903bdb7e80e0417cbc0143f3f8be604697166dc974e83d1038d4
zc50ce41182380f3fbf4af1d941d0c7535708c79cb207a78a56bb1f40003ef30a3f48934bf93d35
ze8c6397e1ebd730fb4e5be683cc137677bd23083bc4c1f95c77815991ccff31c4b954c050dba37
z6680a16a1795a2ed8083f816436130f7ff121a0f81df3871d4fc1dfc132f8432d346fa6d66eeaa
z4c875a572591f93ca9ea447c75167ae2dd57b24205c9f3fe2cad5c7390fe614fa6bec84e2c791b
z40d548a06ce34f994f429c309d9f62bbdbc0bb77aa8bbfceab0461046ae8b6dbf7b4ba6f1908f5
zad4db97f051bc3c20edef5161d4cfbe85904bb111ea8fba13672ae65319315274d6721a0a6fdb6
z913d63a6da334ab5c8779eacde3db15e5b78218130530632ee29e44b8d44814937e438603fa54d
zda2f0aec361e6cb88a2b9a3e297a4ba292e4f3929ebadd7bd733c11224aca1f4bb4f68f03fbd12
zff0b618eaff8edadac73f299f7b552056522e3c3b0f6c88daa5f8140453e614c08d63a757974e8
z32f643c9c1a4e587ea965b2fcd72c0027088d1e01470713b756bb3d3b210b0846c0f2e110537be
z62b152378aad8d7d37714bb2de32bf3d0e0ceef5bd9279c1fca84b1cdefce80cdc6ab62ba6c512
z6ad7461bebbafa821d69e7cd6ab55165b533af5d36813ba00aa10ebc847a6e4239a7e52e64a3fe
z020d4f6f43a890dc28b8a403f9e38fefcd05a1149c2b69d8ae6e876b5d14b4d0d72d8255ec28c6
zefe8f98cc9ddc5fbde3a11219a200b91956ea1fd18f101695feafe553240782ca126687da74d60
z5872a7e4395d3679cb6718ba49ac40727ee0e6735d71229b231e4f1bed48c1d37c23683064a46e
z1e4407f7936fe0be0cc3899b029eec14bbd9464c5d20fb7a3723273ef8ef613a451192ee544dfd
zea5de10325da1e6f0f4ea7d6043c857ce6c5b93a98907f2bb6331e0030c3dcfcc3f63fa9eda38f
z56e5cac5699698aab8b09ece95217a9f08f3a3ad3829b69f63946ebf39b74ad3a84ef238ad748f
zbcb71ebaef153c2c3830c7ca5e5dd28cf253f51349623bf2c6932a2d746547e231f7d6f2bc7a5e
z4e4887a3e0e7489baab6358a5182458bbfdf969ac16ca959b21bc079fa7239825a433c3a46d35f
za4b32c622f1e58cee0afa37f7cb0ae967e7c62935f0f828911f61c17771748dcc23116dfe91f19
z8acc315099f130bf78e5c7b36ddc011dd83219381fe1bcc743aacb9467713eff2a5c2f78101b6a
zf6ef7b71fe7b79b9ed1f0bbc04f6a5447a65e1680b4ab5a50b680222fee001079a54e89ba4bc21
zd935000329ae433eaf731d94acad1f4da77efbd1f8d03ee8f42bc55268315e2fd522eaf40d7bc6
zabd7d83c00e076070b854f4f8504107962e830d7fdb6642e803d775f56c3c58f2df60a6e570bfd
z71d1b739fa27dba7ee2f0a9e410c3b249c0bc49e100495fb3fe1e8671f42fac17f289c94a34e21
zaf202006337096dd788663aac6c8264f3000833f8547aec8f70ec25ec4cba6c56ebcdbe373d283
z23b6b4d5e30ca505c77848457f7af9397fdd12696693aae3bbfbd166a59545ed1ea62b110fe5ba
z85609fdbed2c604b54154a035f975f73b2743cf62b912d3b8648cbae6a3e0114f6c9a0ca2ec55d
zcb45b29d38980e50b381399c7766d93fc056dcc85fe1f61645ea278df2fa3802c506af99ba4954
z70472f3416d878743582b39907b07264d2d8a1385b2b61e953f6558c6bba315b212783e7a7e301
z8435cc7e629c5d2277273504d65421036fab6b0828fc756635d519aff7fa4361ae6d6741a412b4
z7979b9703a9bb1bca27b1310738935c7df6aa4bb45bdb97b791e7de0bde03364c82adfb9bff832
z35e2b11f319db77247e207b96158de07904069ad07ac105b6aedaba05f32df61e1f141244f1455
z98a42db80206db78fc888f5694f737cf0b0e380594be6b81ae0eb256b38767967903a7c3c89130
z5878c6bb1f087dd251a3fb485187464bd8186755e63935ac125d69b75e545fb1edb972b2ac33b9
z5c0012f5b448e48f1d5cde23100eee6943133613c9eb503038704b6693981db05187af1fd8f905
z17320030d5a57a9091798f9d0ead86bc565553eeccf94cba19f940d34d8a67682208cf06e36984
z3054c78bbf324b349e09e7579a26c01583b52ea2bd3a7e83962429f8bfd750309cefbb73125506
z2f9c202949ec6cebefcd1a5b9e4b9fbf4c5f738547e2f00e42562a48357f66f7f9dfec853a1e40
z3693541558b844afee597c3e016c96de5301ca5db5b366a3110d84a63622fa05d7444bc7c73cba
ze08eb600b28df4ffb3f41583e538e855a8f94a9c4ade24940d4fbc3caf32cc466e0c17ea7591fb
z4e9b46a0be9b3b2983ac822db38a9d3ba47c3756e57f73417884557fae5cdd836915f9e68feab3
ze5f41b6f945c28dc413205497997b66f439de603c54683710fa51e13e663006dee283144ec0b87
z16fe35ec088d414e8dd60b38c9e3252a87bc6bc8e4b590be95b762fd4ba93885ffcaa6d0f245af
zb69e5dad26f8fdd26bf5951f06595ad1e40d44839e4f6605d3ec0312117332214d3c707c4d3d1b
z02a7ed8e7336f10e2df64b6a5c2fb00dc531d034a5e305a60312d2e44794c3309e6d79c782f233
za7fb183ca1609b403470baf5e2a4ca0d8ec26cec10ce7792f4adb833de0e96d25dd35e199ec7b0
zd4373e12e071b2f8ca236ec79f3120538b1ca3a1a9078983db9835f5b4693635fd7e0a6f1c7e46
z4c382ce86e02b952ce6a1fb14a6990843271e05c7248d2702ea38badcc6fa188051b56e321584b
z9b2498ccb5fcfac5c8f700cf61cfe63773c64213937cb8394dd3ac1363787aaa3910f5ebd9979d
z2bd3cc0878a0c0bd5d23f9cb787784170bdd9571676e6541e960a48ed7b5a886b655ff7ce876d7
z0aa77438166184022e7b94373a88873fb2bb529e5788960abab366fccad948cb9ceaa22ee87e0c
z7654d678a87a5ebb61aac2dc973acc3d7ab242d7fce73b1701f93eb7641c37102352cacdb9b977
zbf99d928c9b70e8af30604c2a424e38bbe228e6142e15d0d1c97d7d2ee2da65dc5ee4953067283
z67e58c37a7831b0359b60ef162364f9e0c1aab129cb649b32e08ab2984480cd9fb3d5afd8749ca
zade9ac4c4d7f5f8da1785781a0236af82b0d7ac435596c462660710adf9653062ac2405553deaa
z96ca500adc75955b8dd259581b6fe3d9df85991fc3f3c9d117a924379c7adc9233d4f928b0bdb4
z01281b73c40fb4e49eb78c6c45526f477c4ee77ead90ea927e5cd46a00e44373e3075f5a12e200
z456f3767deaf8d2b30b844521a5fe8af9744b3bc76170a7ad41fa37117da9b651d1511c3b4aef0
z1d7a93e7ba3ea0868c061daeec3a76665a7162fada3d9986d8dbb86a03e441101e3056a81e66f3
z700855ec2a5070c1ec768932310fbe0bde73c400a133c5cfe43a0cf54b1d84eb6792da1c5bcad5
ze2a1aecb42a18c21c399c3ece3ab5992bcfb92c2a80f175173ddb5e1e9124927ef598fe4aeb49b
zb274fa097f85178fc85b7703b86bc75bd9e5cd5ef49b0a28cc99b0be4dd6b69ac970d0c4407bc3
zf2ae37847cbefc1825e8d50b13e7f0cf2170ed1a4d5ed32ee068a83b6cb34344b871c58ece6cf2
za3661633b635c0ceb895c119ba6fe42877e9db2aeccd0d32269b70f432eec27cdd6ece5455dc2b
ze01db1aaed40c0a0ab52a81c656c4cf9347c675e9a61c0caed699b205d4f34fd4f4a9a7a5674f1
zf39d330bf3fa07921c9c71fcca74af5b3ac9dccf26eaf6b4cf7bb209d60bf68a8d244588382e68
zdc06b2565bd210aef137fe5d19f5a3c9ea2881b2c3dab370aa7944fca5d6a318727affb8e5d4d8
z5bc78399f3de12e185fc8c815f2c6702dfa7c54f2e783b47404df01619675d5046f7e90fd35e40
z8f6449895e4b9bb09e536177d87286a8c1dc9f36599aae09c71b8b63e2b89ee4847f73a273c69c
zacab83bd9022939c08acbd3497c18ca4a96ec17db7c667eff9827dfa5d964c259e91d9b598ff18
z16f7706b897ce96daa759e15910831a1460b6cb279a485e83536d8c4b84a284c99df3d4cf1da6d
zb1f7b96b2aac1f6be2bffe9e8d1c39a974d52145e95fc85e2dc025c511f7eea03e2366916b1ab8
z317753c49620959e598e274647ee781eeb44a3ad2699d1fdf9413ce46b5f0971c6721957a0f737
zf93cb85ba8997a85bcc6f9ddf2222d258a1f47f580f22e9cbe6882224458bc0e3e1a4b68800b5f
z787d7e10fb482f454f1c095f605f23dba164d213411a749a51d022a741af4bcb92f3b9fa7b5715
z4edb8157df6df7f89a3b116d918c729fbb6182b32795ff588e6f5e2b23e66f4d45d7ecd70780f4
zd16e7d1f0adb295746b4fbfe7473821e3bc5cab7bd4009c5059b55345f1c204629fefbf44fb79b
z30a5971c018b1dcd4c259d246bffd6be20f1214223c329fdd62a71bdb8ba153f27c75b4c909d98
z589a77c9b1700a472f264c3dcd8cc34f75a4faa392dddea2dfc9fc85abefe27ae8a25b8ec24b38
zfbefface7253709561943a663cf81e454d32a229796fbfc0500efb11b387e63e42d0d09d317793
z2faaa9dd4b778c27ac982e08ec7645f7ab72df1529c10ecd759a3350e952833e3daef279d377b8
za136d79421df8c97ca4bcd78681bb8c87d16b2211b29e4628e9ea5f349c94825e0f1727b796ead
z18e6f69b2908e0ba1ef48381f5bbd0134ddf5d07efbd7177d81fb4630864643f59106b6b5ca4d4
z1570fb2c5165e1f27c6ba27fffe0a8576c117ec484d3a1d64ee98fdf8495ddea5aee501af94801
zc6597902733b48782b04b7486b3fa3d99319d28d37edbcb649c6f5dd7feaf026670ed6136e3fc8
z6af9f3b0bfe08575818a5a4c59fa4c8a88f8ca052e8b334565754c69cb9e8c5d9a5794fa24a3e4
zbe417f0688879f08bebd61f1d06351db25baf91d485ad729cdca5f16dfe545d9c25734b71c8784
z7fba84ca4ae60ea63bc4d6f7af06c836611ca0a9829660a05be09f4f6d15b90375604304e5fdd9
za962796e7df0ce9e532bf794a92ad675f729a574672794ea8cb23002a34fcafe954ad27facfc04
z14dfe1adea45343f54c4079511c0dce9cd0be99509265763ac86c523100f5b1b3d0cfbc554258b
z7c99aa3ec0180dee23e8546604c96f0d8e7540ea30807f459fef1856fb769e75d6ed7aaa006fa7
z376b0633a0b4886deb1ae47cba1c896e0759a155039712e2fb8de09d57e903aca59df58bf34711
z8050f6a6472d2fc3562642de6ebcbe8b0de4dfc5e1a1a17f9debb916a4861db67c5ceca4b8eb6d
z113f05340d293d5ea416b2347378449ddd24497cba9699fd5616d420b53340e8d18ea0f0348422
ze26392c7ce67ae874c55fc4347a82a2b6515befce852d5e5d7d7a3cfd6c876c3a3672833f6ae0a
z871900f757f6fd7ccd86f6a671bce2d1bd1f28e5ea996d93b5d97cf0b3656acb42ba84f42f15fc
zeec05662a276c3c2810fad96a0b714a7cae487fb2daa7ca09408fc871fcda7df1c8d0a8ff5c17f
zbdc88dd5349c02119bb165c09e572c8a1398bdb0b85caee7cb2a607d610e411291f3476e398259
z3dfda06ad2d87b0081f2a380a66f42b85b1a0586bae46e8cf11114516f5b7db935b16111791fb8
z314e7a84cea04282158c93b2a1c74441aed7b89b73ad1c43cc4c97df824371e4a630587376b199
zf4da28e0e2888e62b49cd4e491597faa7ef12bce45284383cbdaf92475b37b26b7d888df0149f0
z2d613737ff08a921375e82b99d6782a719c446f347d604bbec72c1855b4cad8a4058a8863a39d4
ze45dc5eb118027002d071f35cde693279192986438407b604cef6b88ba4ce822b85461e0a239b1
zbdb2758cffbdf3014438561fc9b54093d534977fa694159810b88ac13742cff83417a48ddd235c
zd766c8583f7d23a7886a07750b3b3c73a7e19595cde1054ee7e3c941e2f2d283d9882b3fc564e9
z8a0d82eb58bf13352d3ac7a3adbfa0b9e63156bb4019c51831272f249085d8fc5e3af60f158e01
z597c80d8161a6aeac74a509ee87a3b9bfa5ac5fa5328fee352da61de7ffb9e0086d3385a205831
z607d13c6c4c9d8d18d51725729da933f2f361274fab486c224d846444a4e52f70e4f00bf289574
zdf265baa9e3334165dd7482ad74258b08eba9d99f8bddc5da1db01eece26fa36ba4d1bbbc95308
z38b0ecfa6444ff509f744e663acd6d1b144b0e2b037b69619a358e81fd348bf58d3480bff89200
z4797893e02a7fde042534e6b4b36fce2de54e98e517ad941289ec4350de59c6c02647effa375c8
za5aa06384bac1812e0eb7176779f078b755b695dab6864c77626541ce0fbffd53d4656142f584d
zba3e8541a25ee3fa9b749cbb7c4c1dd3bb5a3f5ac2009fb2b713f63e38d4e7e7d493e690723805
z0f97671912628c378669b4a77f70a2c52784899896ec9ee556fadd6c8b3fcdf980681c48ba3b3e
z95e4bf83d7d374b340e840d870c970220e55e5ad1974b865db77fee0ee9bca0f25fb05fbe23c5e
z712af335f1716039b9b4091098390bb48b1a97da4a4c01190385344f4cf0996c4a8dd8a6488bf3
z728d2d8eec644658775a6bc8f14cd62d7bb88e1a839e8f2071055d508d453e0d03f5588e4e957d
ze36c395e0bd7f6fba51de92bc246eb28f572985a06dbef936b689e66e2923ff64aa371ac3584a6
z3228bd74efe4a79c4874511aa43b51ec72b7a984ee0c2c74482216a8b96e0baa93e27ce02459aa
z4152816706e9ee8a7f142d3e83b1271c15c90c31811806c1b151ef160d2403c2c4f4e049f16cc0
za88ec20013a447e64a344d5166a55ec8a5ea45ffd097d3f1e5d34638c2d9a99afaf98ed73dd4fa
zd991f6c3f987c89814ade315982961d752062f74b9c98871491c296d95e0f7fb40aadee33b96df
zdd981c97ae0d22488fff414721e6b7e1018598d76be55aa4990fa94de6e1d5f6e204428824536a
zdb92671fbd9fdd780eba4b9caae3b31dfe744823699e94111bd3021350f5c0e744c31f52cd38d8
z42296831bd90cb48346ea2aae9566ae110a2c743ee1c0ed8eced8d1ba3f42d16c52f5357dc5da2
ze1c65a0bdaf508a38e0955ae7bfde9d222240524e5b4ff000d83ddd38721a1f37d71bf26e90234
z83f236343c196e88b334486579c2da496ecb4aa0fe7f65c441d7db5dbb8b2ce7e6e244c9f71da8
z57bdd55226fe99c21fbe154f1a512a68d18c41d6bcf82e8415ed3e482fffd57a1cee75ae7141b1
z5b0e8a73021a31f7cd0073537489d5d04d3009fe93873ba3d233d79e9120da30286ef1aa36c1e6
z7e35a64c8c30a1267cfb0cbe5124247b9ba9b59ebbe2d1a84a617dcef65de170e1a5346369dee6
z819fd73a9d50b005fb6177d28a015cde02f98eec2fbc268ff3000da639e30cc5ac34a3f48227f7
z6a1372db233f88f66b4b8eded384e2620eb26cfd29c384286103a23d19d859433b267466508b9b
z934330bfdad8a42629fa25baad7c70a2b99c2e9b0d6bc2bf6678a1e3507130b51d860b1cb9d945
z5620309d1041fa5e0e906222ace133cd16a3a1d074f6b5238f22cd5eee72a2255918a1b9cc6b7a
zd7c835cc31d3cb945f1fe806c92df5c394c03bf666ad406a682db53c86bdac81ae5a495758f1eb
z2028c5817a5d03efb9b63d07d391a1f538151e0a70658c9544f8d0388d08a582f1e58bab659426
z5e0edd18aec299058f1725438f6c23e3a600ff3e0a375ad20c8ab8ba941ce0006805c093bba65c
zb50064821e21fb1f314ea0ee91ee21d35bcb87b1ca043d836da437bec32ca74a511f82b6f33359
zd4034e620138a1285dc4d968643f4022780de32d121db69d6edc175ba29836cd1351f3986444ac
zb57cd58dc070386056f6bed4a7caf919c3e05950693b3be6d7c53674d4ae486a1d84871fc00a17
z9762404662fbfa65ea8a65312c4743dfca2addb9d691ccc0d2b4601af4e1df293a4fcb37446b02
z8220d39ccd6bbf0bfb87ecdefd1599ce9ca7fab96b5f54bb2f72faf8947b7b76fe1bea519c0072
zf342441ae5bce8ec9e974894a32aa7fb74a540dd38003e96edde08021d5bd09b52edd2af3608ab
zd95f6229858e5f8d1560b4f41beabe563cf47fc328fc22820dc1759109bd5da59cba27ee35fc81
zbfca429f6bfe15ecef9cc0fffa4654ba0d075849823977f7b333e2faece62705183ee7d7c88f85
z5b72e581be3ccc83c80446ba85cc3c43230d2c4e459a8e9abd5ace9f7f66a391e23a9f353638a5
z0e6b6f0361ffb3149a4f81ebba483148f62aa780d3ae8eac7b1f2b6b978201a7c8bfab44a2816d
zfcd899a97b1b2515775a783d994df67dec2cf7d98a046b610dc22250226dab9762b598ee53919d
z27ad3bd13d2f34fe47658706d760e64b0c4d05209ec90bb0b6d419eef2dce8c5844dfb693d1daf
z45403c9fe8e1b16d317bfd9df399c59197b6562bd3964ff9546153f4a3da409a0cec0dac2fce8a
z74646f24eb636cd2d5150eb53870a07365bb3d04742b309f4b5a0cce99f2fb8c0f520cfd9f3785
zd7c78207dd9b37bf33c03329ad45b3301b5a01d6624d7ef98dee8adde985035e46e824af58a956
z84d58c3cf1428fc8c880c2903b6d758412f6555eb91e50ef12d4ede2d649ea798e785b7c2012ff
z4582d54761a97a392af364ab7e75b000739e3c96504c50f4ac09ccd014563654026291dfd92d6b
z95ad7f0a2f1b33febb0484cf3b3b8ff56885a27fa0794b0abc20654eaf8cd2e39672edef0c6203
z4bdde9b3d84f733e35a6f47151e0d4ff24800ab999790322c43ec8965cbaa37e1b259988499cda
z5603e74432d130d91f92a4ffcf9e30b19cf371278d489c15105a2af404a315a7e51496124e7718
za2d7b5c51de69ba587d4ed063ef5ea4839d740a39a523a7ba0cbc328f60b4c58fddf925093efa3
zad0f7751059766930a034ea57d4ae31f21e109e65ce94a5e970ae3e1cd6f62578135ceb0b4dee6
zc350e52dbc4be3410c62f929b3ca2c19ff7126bb45f3f7134639091be78f2f6d11e2e3003c6117
zcf3fb6132fd43e01bd596302fac879ccf56e2ad0fb38d08b3f253a9c899fcd7e07a930ba2c67c6
zc6bf2e25b78a222565cd154a254bba7962ee1b62e20696ab3e97f9f043c15bbf440dc024357a6a
zb99aa40e6976a9fc3ed7b0cffc9479447c0babc5004903815fe1c16d85f7bb50b5f674d200f871
ze56c8cccd8c146bb035ef8dc686f2b4206affae859edb44d872ad1f489428ccd3b1f25adea955e
z5d229c6bc691975b6265b9bbe13ce652b6a60170d800fee3381f2c33f1a4ffc205eaaab86df0c7
ze3f83482a9952f23a134897be4f984a1b56a72ef0b8350999b036600d0273e49663d0f09c845f7
zb69d0b63815fa391ef45f73b454d557bbfcc8a0b9b20c850ec6efe2109548d29b6f9cca3785af6
zd27c0f0ed733b206674256c4d621659ad16c9d8f9d183df4897035b62af9eb9accbf564b1f64e6
ze74c23d30f352e7b60178d719a4ad05414c29d3d49d9131d52aab4c976e82862c37fea8b40b45a
z99ff6fe06d4755c9133b6bf3c96519877e98b67bbcd70d7643b01d83124544b1cce84d52e1a7ce
z1353067118c900a87f5deafe0ff1c2a6bf73b0fc900526025b704a5bfce6a0b8a16b5f7b07769b
z763503dfabb9ffa8fae0e7a2b86b18ac4820babdf61aa6f103dd650c1036ae458c0ea6c6996617
zf5d46d685c9843969965fcc017d6ec34ecc8c2fda1db34133d470be20837f8d9f9d8b96771cd41
z69698100bd3c819fd4983e265391723668c83c3149e763e1f9a6ac07c5b8f4f8d18453456bd5bd
z945dddd47cda3709d9d250e33b9a4301ffd2268e0e38337d34690e6df8f79f50b531fdcd9a7558
z9e35281aba8054ec23bf8cafc72c74d3d5c7c8e869673e25ef2eaf108214ffd3af6038603650a5
z2907ee6538be9cb69ecb77e44078b1850bac2558db9f66d7a57bc791143c6b1f4cdef80ff2d846
z19c897f9df649dec4ae4052a5b995503e5c6f3076092a37837b2176f574480cf4fb9ddeb9f9930
z8c13a72f5bd2515bfd1bcfb86282f171c05445b3a5015ca3de5d22598488c04e0eb3a12dcb5e87
ze0c0752b84ac68483646ce5c219b9a49753a8c70fdf3cad4263fc1cf6c9f0815833206221c37f1
z5a6323d36826a817092da487e0770e5861503ca05de55c002ffb8a86a12a43a76dacc069394c8a
zbbffb03e7f874bd4e863d632dd2708c2b18416efd64a17fd749dbdb365866bf6f343eb6d70a5af
ze9a5ea6c4a2508934a20874faa875df7eed1243cf2dd43eafbaacff92dbee958c03b7b132b802a
zec884fe8dbedfbce13705ec3631a84689f3f36a2cefc3deddff7fe061e04c126a89d749a25e889
z1e9e6bc43f8257f667d00ce1e218888ae7f57c4094e9714bbe80229f16875d59ebb18e6a72133b
za4682da25ab4d54c33ea675477345916c78866d3f6ec2d3ceebf0e3012687f8ab3fb48a0a7a3f6
ze4ea55b0eef87e6bce8f5a5d6357c882913f3317f1fb246a14e32b2aaff3210f88baec37b7d19c
z417a8e39b26682af71c03ca1f11a67b4504ca6f26f680b3347dd3416547aa2bf0cbc3d021c6a73
z688d44c1cc338c75522745a086920dfc57c000b5f5aa2dadbe1c7fd6a823be601e79764385e00b
zca1fdf2c5b240fb11ef206125ef1903284c07d195337822d9844d4828882f76d1c606af6616973
zacac755f94fdcab5d99862b8f56906e94bc09833ec0eaad76b3441371925d068683fe662ca5611
z757e5320588dce6e7e06889702336442c2d905d8e189f99acb47fc6ead0f6526196b8e5161f2fb
z6828a8d44ff147b2b67e4c0cf812c533fb706eb742b5844591417965e9920a815056f62cc69e21
z94c6bf42e8c8278255d05c0074b02be8ba73a7df92cef771ddcdf3f37a9f4bb403d35a4aaab239
z07fbb1319ec40a2e646bfe78fbc3a5a5d51bd51f4a3cc7dfaadd7bdaf9d524d2dc5dcc56270796
zc30b40925802ee5a1a75560ab084b4e6f2e7474a51ce6321f5334d99a3515a663b83d7288585fd
z1fed6166fe29617c5568ad35a71e6ab7d1e1dc9d17c5be879adc6d73643db522ee5b1c283c3415
zf2c965bdadf0aa8243dd310ddb90210c425bc2eca011561a53bae33141c9c49d9333b288fda74f
z6985911477dd422702dc5849ba9833fefdd4aa8c5656de5369ae37f4939b635fc5edf444ed9228
z2df1fe7cdebf4108d8288fc6d4715ba57a1d38b12692dd9382c583b90d5a0c2b85d81a1dcd58ca
z4929363232504ca4b4a8a7a3942c6244868a1226b6ae36dd93ec9750305b8645648756455d66a6
zc01f814928e12580448d94b4d84adf79c0f4ff028e36a769c4df19fb2b79584a4a6a3e855af60c
z12c91c67d7d79b42090be64da3d6c16e140111ab9729622ebf32b1783d1d14136174f3065abf86
z4c52c193925b0345e3871bd17fe6fe97d05701ece5c6919e359bfdf4e1e5e5cdcb8faf6439a187
z2ecd84dacdf7974cd60082f6b39979fe8cc6636a32cd1bbfca03ff86d1adb116ce33e67e1c476a
z5eaf1751bb7a04b296b5a016f414534c835cc355ee00c60d9318e7866922347aa40d6c40d05bc1
z2ba0db45941a3c954414b7c14b00c9e4f9fd5afcc028cda4811d944fde220181c0c1b17a505032
z2f252014114701a881d8fe5cd5fc8d6adfe33d05be471a350c6fc83ce1e04172d6719cb09bdc7b
z6fb822f11de3e1947ceb0db2b37aa94baf860d18ae91e610434398fd051b9e67cf2999c972e5d4
z14594741b4a69351ef990e648056411385d47581f43380a1403034abc367f0db588918869ef63e
z9452af481a5fe743ff5774a332081fb24d082dd99bbb6d6cacbaaffb5e81cbc8e7b1d498764ad8
z70300340c4e3e2041d54f537e898ef251e75a828667e9a865eefb2f01937d9d7d6ced94013244b
zf3725d3fba8b392aeef353b11807581a7e313d5a7c76ff77c3a67cb035d744799a6b6a018e50bc
zc8feaf2a38466f6cd385b771da1bbc8f435ac65b7902aabb3f059e994be7094aae6ebf2907bdba
z0fcf36e5ef037a0cc0288432c7821063a0874f203ae125abd0204b6ab1ba44bb0623592b638553
z9a55a8e3e0b71763fe390c441bad6b01b1300acbff68b2d63cd7413649bd9eee65f5bb3ad74c7f
z4c831ceb9474cd7ef52251314c430dfec658689567f23c15489320bdd7408b00a8fc7173ea4c94
z2218aab92724a90578ebf0beee36c31921c2242a6f81cab72bf8009eaf927e230cd49d555480d9
zdc42b36a524b3bba9897586aef3f7d9d4bc8f6724a3b9b2d6e49e000f8d0cad7d55d66bf945ad6
z1d5c93f57fd7f62bf9b546e2de8079a6e1cd5694db368f17fc5f0b30ab3d1abb840e3ed6201534
zba757890e7e1f1136e7bdcec9fa3d26094bab0344f6182356006612d24f6427a29876bd2bba88d
z62d12caf5b3e9d185455ab5870c178c8123803703cf2c589f400c3f56f354260352e5067cf95f9
z6d87e86db6e97adf8d4ac95b870371aa5969f9de5458e4dff3c74220ef10c9659989220cc3e8a2
z31c9920e6c4e44f9c7fb529f2f8608e4debc87451bd6bcb6c8634c5f5ad12076d4ce79146efe60
z86aa5b22305cd00450f1772e03dee41c2223a54adad6fc79f7ff59234e8d398db8a4c83505f971
zd23c94b4fe2b41d3500e5a71893015dcf55959d6208f01fa32cb8c769a5c81407c296a32718cfa
z4b5f6096530bc54a44e3d9df614b2ae04b489719bca885bc1c408949350b9d3321f69ec58fa97f
z7a08b565a8d28338de24c56387781f93cd931451be0603c5b2226514f379b22202fbb8c2d68532
z95420299c607c41b52a684749c43d9fe4ad711a23e0a7a9a6df5dc714e3815e9001da8045051f1
z0a157830e13258a00686889874e0d53786cb980a2aecd539414314d7adf43977b1fd7b0fc4416d
z6b90abea1e0614499b56b2f8c476bfd7f930764fa541686e98caf49a1cb0d6358c59d90e7d6478
zaf7c0d54cb15dc4e891e261abec7a85fff5d7c6bf8d9d4940427c5919e6e442c9e10eac6c1811c
zd73fa413892e433777038782600498ba495780a5ac4c5ab61426cbc0ea6df2b4e137f481b3d033
zfcdb498a723c9070b0fafbd701ca221a1205f10cc63e795c613ce064b758e96c8f573a9e09afa1
zacff6efd68c926c3a2dcf3c8f2db11ce2f59b0f082341a7dde3828409dc0e81e574100488df6fd
zbd839d11ea32acc8d5e1aebfbac0f36a5a33ecbf00faf5db9d53c8e21faf9809ad670fc5a4157d
zbe206ee3e2e438a3af1dcdf45d9018a24a983e1bc92b6b5b9040e33f3aabd4ac4e9499000dedcf
zf29904dbfa2dcb83fba6fb25baef38df415c8ee5b9dd6cc4a65ce3e7c85ac885cea572fa247fab
z06566b421a50be78be9d0da7864fc2964c8a967b280e13a667f55ad7354efc185925c6bf39c3e5
z18f9245e374eb6afa62962fc040a0543bbda01d2623e5f5aa0ef5931a240808b2b7c1ff00eaa50
z2956254340a50de30e943d8a03f566facebf2e72ac54352b770a9a236ff4c8a3e539b4756d9d02
z36b938ad70716e7de4007220fdd8917802edde129a4726e9ea3b87af3e4b697b52b00c78cf7f72
za9a7133fca86f069aa4a132a04888e7b0880097269f10bc226056c34e9198c4e9d6c4c492b10f7
z0239f2d3ed980c42fb275c8612fde2b47af39ae0d6fda15043e9c5f313f6716ac7119ca5ffc508
zed1bc284150ab0349e2f27facf472636593fa0f5cf838eaad9f8ccdf0dfe9d683e46b6e685f25c
zc03588d9e74af2997ba0598c3d6da51a5f7ffd4f6680c79acb56463011d871af2a15b0a98ec38b
zc97fba86aa6308144bb5b612f06c4b9a67d2915159be62dbe0e39b96ecc54b26001ec8303bc087
za7ae8c0bb59d831a0cf84d86e10900235239cd91c424857e62a1f2e52945e41bccb70df1387160
zb48e81fde1d8410191a0c9cabbd49a9e2dc8a42f3e6268936c0088598c1216efe8557256319c74
z5b747bf9f585915cec193ccbb8626e377ec96c7356018c809c7b2d68250bc92ae33f2a54f302ab
z639ca6d5391c0557e0120e1675929e17bc4254f43761c52db31ea1361a9c19e969d588ce56302c
z3a8267a342af44368f75055d97bfb934f2963df8fe1c8d4dd2302431a1a7e58a73e8965ad7b1cd
zf8e9ea44343b3aa03af33095d072c92a406638fd13220939d45273b640acf7e4e4f0bdb8769eb1
zadf3a159c2364ea5116d7e3732cb87a1513ea8b828fe6f87e42d0ecf342815ba37aa14639d3f49
za2ada8c5169755501e97b6e32a0ecb26417566c22158b7f2bf0f01dd749585b9a28b25200222b7
z5e95b1586d4538d1f4f0c6cea4fd0f7d641fedca92d0641a2387ede3f1c3e86d52334763253314
zd80cca78e48075abfcbe87f027e2352107ff9017d44706a98ec93f65794b684cca139e60af938c
z46cbd2e67311c0d0e73b29586764f32583047cbd8263cf67efe3772fc06c6406caa9faf4b46858
z9a7e51adc3936258b192873b98fbf603c4d07a6f21541c35aba169fca5602700f22d2acf510af8
zb3fd64436c4762da2340eaf1ad9d8b47791f3336078903aae079d11d3d5ce3c8f25b0dfec2c356
z7a10b2db9a773b5e5e0ca17d04a19973599211a2d305b5b0c3a432618e8da68ce3b8f9e344c1eb
z85cf34eb87ce6b86471bc521ed0ab5e7d515e932c0d8690d3bd0a40c3fda7825d823e8ca202e43
z65ab5c422a8a2fbad213e052bc825c93ba11373e207f989b64af2459baf1839cc08d344e11ed4d
z9863b5891bb1742b94421cd1724df0c890974107d7ff4561b335ea2738eecd615f004f3ee35262
za70226615c0c8a81d1b02deb21bd1ffdf6d48c16e8aa95a2ffc023f397f984c9656d7399d33fd8
ze5d95239a129e3154cd6d02583c833a799bc1cbbc6b072065e16ef50d485ef7a28af6b4346b197
z3522c1ed1a7c5a3b99b39491b17ba1ae13444373d6acc91d789be7aa7bbaa4426532dbb683be4a
za9c23f6986898e5a344c26aba99d0b93a1db0352a4474aadee0a2fc50cdae065b186b56622f9fe
z978cceb64d16c16af8c4909e824f9aef8df2a91f81762bab24f2e5a63a5ae5350f073221a5b831
z590c63f7c37f6cfc463fbfd2f0f0250f7557bf926e42238fd2add4d698806dbc8266ba0bc89389
z9fbe680afbcfa7893c248dd7b40a8211a17e101ed5bcaba54dcdf022e6d0a4409fb0d15a6415f6
zfd965fddb7b2a6f6c8cfd820915a342c8ce6ad4d2090f5640a66e847d10162f73e10f24b6c37e1
zea6d7b65a52ca9b7139c62326dc230ec8a5f9adc4e13eb0bfb24ee584e844c1a911e570a8c445b
z06074e95252e584ca28309a9dbbc0b5bc7e88b7c4df9f1fc0ff9e742f12672637e9c196e0940df
z00ab5c78611214db4065776150f3b39d93e6cd9bf78bec43099dd1f75675834e9e90435d2f3fb7
z0bd141e828180ec746b909f41e59b38045a89279ab4aa28fc19c01822ac0f4be255004693a0e2b
z8c432f119ccf96d58d498a44c36edc03121b3427c3a7c8801b6d08f12fd2abfbd57731fe34fe19
zccfdc69dd3cd1930c1fe71bf813917a0133d53b52eb47ff3de053ebee0d8710bb1f4f11b6cf606
z3678d1ada077e2ace5021c8b16c75674968955956b7e61ccef92e81a7e87dd621130295a45c5c1
z54c4e0529cc961f37873c8cdde227e10b7631f8b134bfe59d75f123e5cfc99e37c02337b860e52
zf10e23342626e831a86c2dc79aa3fbb8612347745f708483ef782b70837c0a297052c4dedb27fc
zaab608a69d6afc37f0aa10fe0ae022a1877b87258ee6e3ffef6bf68e9f9aeb5f046e509f917374
zd5a447435cedd3f8298eeadc3d6b27a1fb25028e24812930e02903f1511dd1c52712e426f5fdbe
ze22877e56acdea56d698419d1a65c0e0f06dd1edbc1887f168320727c35197335d3acc0d66ad70
zb42518589da64741e8b4c02f08a1d4aab7a15d8f076c9101d727143b194cc070043c2519d72359
z333708778b34ef785233edb1ac946b84589e466febbe3de7a96d7271cc6ae6a578bb78430f1459
z4a7e4d711b23d508a32915ff096ab95388fd52f4c5744b8d624fb6f6adb26c3a3baac93941bfc6
z6b6aa1e3c9cd5fdf55e7bdb35960bb14e7feca4979bb157662cb3b09d867c4e76729d137b150e9
z5d456cfc35bd86e711a1742fdcdd41e94ffdba851fbc4f7621ef92b00adab1daaaf96ba69c9d83
ze336d28dbb696e6fd47dc22df7ac792a7a4aad1fe179cd57d38e0d838c02593f1c95d315528c00
ze010a48eaf2df703c9adb57edf279dfb4579087f0dd342b0ce243806155ddcb1d2bc2132af526b
za8007a199d89d866f0fec14cfd7015424fda52f09b39b7f6b30d29751727ea8dd4654a89fc45c8
z688faf72e849bf916872cb079cba1aa6c4bbc8507827d1d8893df4d45ded8e48e45bab27b808f1
zfc16e03fdaf739b0f610e1d23933387486174486875dc9116664c36c087342a04e65a1c1d25d27
z37db8b8e8a1b1698b52f602b4cbe832f11623c6230fb74e48cf0cd44ac09a3fb6252b4002aebb5
z2268ec8fbee957917edb0067c2a0836697a170c94414b726ac33b11efeede74149442a8871bdb5
zec17efedd1096a4f7cdf73d279b99a1d40713d6b512906c8d5ad817ce968838f29ab9facaf2cee
z844f17c2a886871aed6a737044b8cbaff9ff94e8c3af56e231805d4fb8a8ed48ee0a4022c94bc6
z319f52db08a5ae17dcf1fdde881001d162527cc065d8a029dcffb30e2a9c41b811afe64a034b2b
z3c99a6e8047ec89690dcd8ca6db6a06d45e6f9cb9be5393fd9dbfd20c7b86a7e098cfa18089380
z45536dc74b57e7891838ad287f00b76e49bc66c40fd26b6392bd7183f0e16f788611e3c45c6244
zd59ff65352442a89b1714d81abd54a1be56c71247cf9032beea0dbf1a7845ba2caac4a801f56cb
z4ba9233f9ad2d425d9e8c182169c34dca3d393b272c45e356aaac584493c101b5e7b3ac10a7a19
zcab10cc17287609c28abbaab0bffe3d566250444715d67d8c5044fa65fc9d9c72eec53eab3890b
z6c5175e1ed46293d948690ac1894ebf290b2bb128415bc7d2bb951f1997a79fad7ec3b554e0c28
zbe0b9826db6d2166d3b2c2f5d8fe77832b0867a3995055731f21e3883e2740dcddbe4d01742f5a
z3d4ad95d10a264d763a67b2f7be7bead9e7200ebca1256b4c4d17caaeb4f40ef84371d06f77046
z40ef037f6728a33ad1e37c9fd53f9a0b50c9f88b33b17364d5530d316bc03653ce74899501c550
z0af4ad370227906797c794befa41da2fcab4059729f698c3388fb4b4839f48b191783a2ff73d69
z04fa0c93fe7623ee6cdd97d94caa0db439ec9d1eda28511eb3faa823790560fc2accc9a2094221
z934a2b7d7e53144541b8b9e777db8835dd53643779e95b141dccdfd5323575120eba5afa134883
z7d64cb3ebbc00ee5d1911ebb5deffd496acef2a828e08a0a4b3ac42cde3df7a64bc27736c80c88
z4e7d47c4d8f6b50728b9a0b0a76322ea509c39728435c08a03493caacc3bc07d1cb75e61d0750c
zb41932d227526a05864f15baf68e1e5f0bd61acdc069e2c9870af4450b62766a2844f20350f69c
za6c83c35c949dd00a3a35ed6ed3008abd827a5424937f74934c38e04018edea5a15b3026a1b0bd
z3b492397583b4eaffdb2340d539dd484faa11bc0efc344b6be91dd8b18087f742d218bd48ad220
z35c3d10a0feeb0dc3c07d74d039bc65f2e0126d7a87eb89b35cd94471ae30c9f2a872fdc379b51
z9dfbfe0cadf23a5eceee6d9e79bee360acd19ed53c1c694cd027bc4321c4fa4f7d59fe3c3e5fab
z9963f6af2b668791d9ce978b3cbe17f6478853939d7d1f29e07af433d209b74e87e2110b9ebf92
zc78ef9fd60066b10f74a22ffa01b1bbd9e3aa91c471a8a6ce2f24b6f16949d1441d233117232ed
z1bdd226d85961acc31eee32c59038d3ee9dcd48767bd9f46659e91ba544564a03858460378b0d4
z6958bb1eedea3efd872aa203c8a75777f22749007e0c34367af0dadaaec3745666559df83ea58c
z166897f01724afa87d453b175e93f4c874d84f90c66760ca97c51cbb10201f0640805011ccf300
z62baca78f79e3563eff32511995759e600a1d3f2f6c7330965a7a011219ddde11b97bfa8541fe0
z9b60b58fb345b4378229ca2746d330f5dfc56271b3c5ab4101cb3fb3af6e82160a9ccae9179813
z012a2cfed89cc517b87b219d56df59fd0b54ee27912a9be5291b30596b231cb6a378cff6cc3668
zd3587b25d4716ca26283527efa617467d403a232437266adbbaa380b780b11e5df79ae61aa553d
zb7fbd4623e7c17778dae3e7cdd330e81b33c329e84614ae61414086a292d0696725a0264937288
zefe26a1e599278d5f11ad8b4e964d07cffb7c1ddab0b01e26dcfe5072ff3d7561ae92427150f55
z0251cccdf6c1b186d4648e19a50db1ffd2947f7e3fe6d6ba005757c576a3510c607e8e0b254d9f
z06f8fcc42fe80fe16e5ffbc007eae452367af2af4500bb2363c07c880fa27269476305f5c078e9
z5e683627d9b9796ee02d919087102ad4759b3c1af26b58d29f9ff8ca5a584c339153fbb388b70c
z2060fefd5117c03ee8043df8c66a2216677f7d7e79de44e098962fac0c834461f409f810663790
z75da88071666baee9b939d0198e7d64c9e09105becc27d555e4ec568f595d4217cf1172580d418
z44a94c5434aacf2ad5d631b188636c8716ae88c410816c288c792e0d0b2d00d5217f7ffd850ffc
z43c72df121a79be6546119e66c344374ce064e720728c4ebc902badac81f5891f02595e47788c2
z0ae378d35d054007b20013e4fb02629c4aed6d8b457d30ffd00af3780ec45ad076afe6a1562386
zb3b5e084c81910a07a3a401c60e3afba27b4ae1e738c40b424a62ee97737818d7295614d95e1ee
z9ef7f9fa36f6e02a4b8f2e91eeb961fe7e2c6deb46842a1c9dc34b7deb1a123e791d4ab86877eb
z4087bb21b11e1ed178a3ce0a954de7f4b213a63a819fd6ea87563fa7ffe732d2e2be73c4050fd8
z05408b6b9a3bf6c9953819e30e23b37ebcb1fbceca132e718f42f728aeaa6991f045d0637625b6
z79abf3d7c17e31fee1ab755c453818a923f34aa7759f16df291eeecc1048493fc84780a4615bab
za47ee9e1fd20c9180eadeaed26aaf893731c462ca891c35d7ea2d0780597f1abd0a8552380b828
zf1f55ed8f968d6f045f12bc1a0e84da2ae0854017482130e81570961741ba87dc8a91835a31d48
z21a3a34ba5eb4634939e409ecfc15c8dd32666ef7afd80f6d9f04f7df620bebc2ea8c3bfd7cb05
z8b7566661338c2c3b698a232af81f8815543f08e9af83e7e934d772345b508dd934e4ed3642b45
z05b1474281fdbf3e229974feaa773b51dab076a7751eeb78e5ec1163ad7d83948ac825ca3789d7
z7544697116e4e9ff0281f500b66267426e475a5d1938bc3d8ef6ade8020041d6275f5f9f5ca6cc
z4e960bdc3250e6df5c13c2b4d71075ea6651764c96289fcbda0a11d3a6f504955519ffb0e3065f
zbaa131aa6ecc4733364bbe6f40e652a9b50638a43b50d8a3150f8a10970374f57500c9082878ce
z4c469020780e8cd776751c216182348e7880f7b6b4d4160b7102a430dfdf115c6f86ac18b7f47a
zf37a1bda5ead1cc98fddc45b989fbafde8fd04739f4223656928b21ea1a5aa4ae9e67d22ef2a80
z0a0c66f3ef6bb16f36ca87c55ac3a2fe6acade5946a650fc88edf0b5884d03830b6b24eb0ed9bb
zf0a0c36b25a6a0d029f4c9d7c50750a9dc23e368aa0143904856b274d08799192a5bda62f0c064
zad5eaae422042c6b1349a72bf7e81214fc30e25ca2ec12932be668527bf420dfed345e1e5c5373
zf5ca9a9c6895d3b8b170a4af41f248e28c32224fdc188b38a210cd58630e23afce74e031612964
ze62dd47373cb3ba3cdaea63347184d45fba62eec1893aa21562b34fac4f91df80a4461b36a2186
zb5b429df71040a601e8b8b21d1faae0209d1a120b97c03135a8a24cf648ebc1c111c8461c73508
z385fc55a4afbecb1e9e61de9dd9e272d61e0556f465d8c5ac5c17b8fe1fb672d32cabbcd7e1e71
zd794d59222921e2c17b21f20ea80cba4b4dd81ec05798f9f908372a38201bf2e037bd7e58af348
z9c22d5945466908a6267be3d9f143d6c09a4e3fefb0d5a20a5cd503da7d8686a0b5b4668ce87bf
zb213cd8f47e02c08769db358388512cb6fddf52cf5b6aa095bdde2b27f21af4c704ec92ae98193
z9f153ffac44bb38bf3ffb97a997b54f9477c8c902e9a8e8674c460ac97c3e8f60652c9ae66c354
zc9234db6471df054fa70dd514d214e697a3bab1481c33296a19ba40ead7b2240df8eb3a5545611
zd81403569c9b601d46257de4e00c95f9b1ac841cd7e4d7bea48d42f45e2ec2f0808fe123903950
z413ce448a91327c7a5f8c4676608552b21dae6201d49fb36eab763b193fee3a7ca8d0cf75d7537
z25fe7cff7a20808538378eac4601304008472f6884f22f7f4a20ab9503ca565808d86f89758240
z1d0722263d88a63c7b76bb63e2fcb5e96d6fd3d69bb23f1e5764bccb01f3e53036f293d21427ca
z120724ac5b7f34ef11bbeb59fdf92f9162a21660d854b743f40c7e1d09861f514ed927b8125a86
z0475098883b37f970c7650b3498b1956ff97b2ffe6667a37a40070deaf0d66c009d4340090a94d
z7d0ba3cc27b408a76d1285811bba502f7b7620be059728f3de0193cdfb2dcbd30d4cf07a3b7ca9
z9f8f83eaa315740cc57262d7a56a6cf5b8dc9dd51b66ac73fb88bf65bac31ba9f6e486345c509e
z8197f5c572e110e087c4f582e851878d8285ef5b86909ad600e49ce7014f750ed2440e8c26e692
z0504ccca2b70adc163ade4d9878140938ca68c90560bdf5b3f124b2a83a78ea6fb6cb7b4f3abf2
z41b75369f8ff759bc7059e35c214a5735285219efe155bb9ec4b4719487d7aed391abc5c5c2156
z82513eb907e93c9fdf7eae5f4ebf74bdfc291c43fdd61f128e8cd0bad1b881c6af16d656c53647
z204c671e07ac5751cf18f1223d6fdbb19df219441da38e99b1caa86de50b67bd350c2b7dedb201
zc9aaf8ed269c0f62402c555e13d29e9ccba383b7b2c78ecf6de80036296f45e3422cb79e47a978
z81e5c6ea2555473d137545180fd1111296a9965363fc9ca7353ab170384c54b8502b69012c1298
z68f139c07a00cb45f3e757a22c83302c8ebaad7f218cb0b85c33b7835be090caed094b12ca0146
z4d04fa128a6ff342c88634cdb33c1bfda0f38aca0cd507bcd4f7d3738a7b9b5b85b4610aac293c
zd156455afca033e14d6fdbe7dca48633a11d74c464556fe8dac8d788bbf4404fc9533748e41a5d
z008960aa5aa86e95aab7a0691e18b8456107b56f46f40ca4eb0791d145983368ac9ce9ef39eb5d
z48125f196e177e187fd224c6df3b47c06291b0e194e920f13667661af7a3057a4edfbb2cfb4bf3
z2e5dfcb99af50c8b9474d815401ea8ba76a8b30900471356a1365a8c056a1e64f255ae7126d326
z50d1fc0089c07584e969698d990b678b4663c825c4f6037f48acc35ce95e6acbef0f39ca2289b0
z30b07d4641e1f434a7b9bef08e9b319252669361f7823e3203667dac88a6e33cdfb9ac43773ef7
z90abfc609929972866046ac4fd972f77f7b0e55145a2edba7edb44bd931db2c436415988970f52
zaebab4d380e80b8d8ff8bcdb3d9cb174690a4d43144f2467ee405a8adad518653599ffb4a049e9
z66f7b08f05bcd2632eb030ef13dde68851bb82e0a89c11eababc09d92a164395a2eb6e70a2774b
z865f4c8b331e01edad5c62d79d6acb359c68116633ad5cd4e0b33914e26ef7dc8f07e2ab467ad6
z71100e1d97064151762300a5d6bae06750f92ee77094a7c5be99fac9144104d05199bf1a07530e
zd600e40acaa573f7c84df1b92f54ed436342bfe8d6e81f427ef93d9ddbd17f78961e392f600c65
z7543a630fc63d8ff9d4e42416766fe0e3921ae7fad146076a1a535948ceee9b4eb673255212887
z81de26f0e4593cf4c9673aa27dda144931688eb814cb9dfb247ef28572dcd8885dc875fc4eed1c
zd0d205e2a1b99d01cd858dcba22bc5561612303fadc8a31bbb1df8e16455c35a08e3631eebd82c
z4469218a5144fd2c394c4f86b20f480db83e477376c5bbbd0a68d4a4ca2b3877bc7ef7d426abaa
ze0dd6088dd897f55cae0b3082d525f0f96a440a97404d1d44b6086f07dd60c19add2fab4229124
z7dc16ca6944e19a466682488bb3435afb18f658d1c414846542331f206b725e0504d308f03be90
zad82d7f1a349cdb00da0cbc3155923995d83b652ca46e5858e625d5f34e37005f7b0a43a11804d
zb8e4cbd2fb0f642cf3abffc144d30598bfdaa9b50e849d2a2b6b8a8214f2392bf27a1821a9c5de
zc3c766d60b0da8844ca25aec1ad5cacc232e718c8df71c954dc876e49ec967142de047023c5892
za7ffd5b140b553bca596617cd0e6534d1c4fcfbd736d599f421a2675fe58c9311d46ef9751a14a
z392c14a1f96d3f8a1ac64b1c00ea44d1500d10dea270f7032830156a7dca14f103607e6740393e
zdedd61a6ef5841150d9adfae70460ccce78fb43b2dcff152d75673d4d9e57f8f6a6d2f0924e831
z3cc4887d391913f70268d8769f72335d7dff558ef4cec2562d218d0c4674daf1d1ece74c948642
zd406c8adec43eaf9d834c80f2f8bdf9b43728ced5c0b36b45a0777a451345571251ccdc2b9e39e
z3840f1d317affd9abc26b6f4eecbb95f7673d88894feda53c5ffd5f46910a5623361961afe0017
z563ae2684b5b76a3dc562c30238b57c18c4d877790846db354cdd104f65619436f4b5bb972fe30
zd796088dff86387eaef98910f85f08b084e7b7f653c5626c823d2b3fd1428f9dd716ba239cf6a6
z60c71a6045bb9322cbb4a3e9747328ce1dfae1975d598983250ef5b0f16c0c9f2cb704832b112a
ze95dbe151a0ff7f63317bd3ee631ce80a3be57af3e5b99b005ea4df06c74ee97f790ae09dae918
ze7fc6f69274e4f6909d1c67b50164a58299087b3200c430332e2c576d073c82895a92ff9912d67
z767acfacf2c43e0b76df99e5974281f08b82e54ba6b123816f3935e024272ff38d2c892e72eb69
za73e8e866c499ad10a9f80437c93d2b8e24bdf1e9c7c7b512340ee50571b36379a916d8c05c281
zbe042aa473b18d2cbd64d73442dcfd17d1e0f9c34a2c2e4cc3fa9d2a48cef34e194100aacb1cc5
z674d2ae0fac309828e31e845cd92a1ac877eb3a37767c82ebf8a93da4d847b6437e3cafe125899
z74af4cae6867f70328adbb2a7e1f52156901ffdcc0c1c257b2db54366756dd1b663d389dcbfb84
zd95d8e5a9b1d9c65f75699bba993dfd2f93eab9a8a83136973f7c07436b30cc0b466a30a9a8652
zebfcd514063fc7cc18c00ebd68565a69d841f97247bcf8c42ebd1b661d01cb9ab07bd94aabce3e
z6f20387af15b2b6936b6d8d6638ed5b9063be074c1fe52a2ca8a00ed12cbf66a7818285f9c8264
zd1db7a8b9512891e537d339fd7d1feb2631de6e9c3106899ff9bd8d9d27982434be3b8111db591
zb5e697bb88c861e45bcdb77f8d68802ebfa71149d150a659426195dc289acf0b9ba3b1c6a51516
z87c851824f4ccbf998e4684ec48a3a799adbe761e9fc6972b2779eae4fe992c78ebe6af09aa9c1
zef32471d6bbe4bc897d15f232ae3bac62b139463f2f6ff73a9e449ab201ce6c447535e1a5c815b
z184d3596f0a06e4edbf40af9c0b8d1a0bcc301b310671dbf81f7729c80645057ef3ec1de519f33
z1d9352c07a4964e4f9952f0298ebef72070dd537fa1eadb0de7715c1dbc96fe31c1894db080748
z0fd45b6bfc98f1b2f0f6a5b12283b4fa24ee419f63122602c910eff051a913d45d7215ee29b218
z857aac3fd803e4bb49a4a4f7bc7297110f290155a81a3f8f2b82519d33c3cac872360d1d8c0714
zd3af110cd3c5c299f59b22f6e5b213d472e3bbfc470029f0e97896c46b7c9eb2697e036c5e6a0f
zdce3d907cc462ce9908c8b830595a9158c3ef6128dbc13d3918ba2f7ddee1f8f181c81f0b42222
z1848727f535d6010e30fad60ea0aada4bee8fefa0bb70a2ae334059d56812a6561c2725b245232
zf248a8ed2f3fcd14cc7acfad297f38f1e6a30f9771c3cf9cfb2cc48aa4bed16e61326a5283547c
z26c2726afd0599e769139bdb7e67f4860c510db05a630848aef2b1265465a36071174b12b9cbd3
z0a804b017990467cd5a3d308af645cceb645bb8d4b5a5671ae4d7c362e0f552f14949085e91de7
zf3f017dcbe8846a9884e1270724010aab9f2eec1c2174dec98c424730b19225089ce7cd154e657
z98ae7e5b2f4e2101fa139489a1ddc13ec24dab87d47ac4b800b48284ac7421a94352a2cc8614af
ze2dd969be1d783b95b0dbca674c043e7fa1f987cc7f55fc64b7a041ed486695ed48b9b1e99cfb0
zca6de295d428ac3750220759d70ce52df033816ba0a077fe904760ec582ad6fb2a76bba4bf0e53
z4e41f4737e01701dd0b4fcbe6f40e0cab2ee0803c18148d22de6d548bb964c85dbc4e53111a17a
z2721d84826bc92e4a869fa992e52d3817a0db1e0f656ebcf7f25f8dd4bbb7033d9b9793f784375
z2b65fdff0ed6226bd87152b4728c6fa72e6daca02328428d5e6cdf1572289a8917c1c4e8c2f59b
zd54e2c50f350ff5b3b3c388aaf536b19705ec66e17f4d25e7c6b2908aa02a7c956a21a874edcc2
z6828aef87687c4df65311fd5b354d2e0ae442639c3838978bd0dce053ae37e367369da99557b62
zc7efc795e7f14df5ecf9664c1b7c02bce6d112bc5cb0d39332bc7cf6bd35a8e0d652774dfdc19d
z629494f6e3d96e35060204f5323578c3393756ad5d12eb0af86ab5c36114e6b3e04e9b920e7027
z0a73ebcc4615e20c9fac67aa7b556430ab1105cb3c4fbb98f486cd9cb3da59ab9dcf3dce678ef8
z6c55a93b5664406dbc4f8471d7d35171c57c23df48462b5a4266e8a0c974c4eb11241f1d5afd79
z2c3de0ce65148e1d6b69a3f651eb1d5a487966bd97cb7e1dfa14638983d1bfed06f5ee4d49689d
za41dfabf25785e80055b1b573fdb75a89617f7295d351d05ad1796bdb120bb0c76a9b1bbb2d3c4
zefa514ab843e593278a7a97451386ea9c5fc3fff0c104d408ac63f74b42472d0133a8b8003ff92
z5bb7b7ab6d21f77d22fbe221365c4511af56dc7fb0fe320c688a046d8008d97ce640d516656431
zecc9b4b0ae9ae5b86de957606a5c1a30d15ea51227589b2fe8c651baa8e073eda21fd266a9a08d
zb64e2abf9c5b5c923418f25459c011db0cbcf40426a46b3ce92959484e0f301502b4ca5511a87f
z109c20a993bc3b64005711e1ab9a6e09678aa43879f97524b86b1caf7d2dd50e9bfbda12573d5b
z9032ab09ae676d65fdcdd2772ac977d8a9f5039f2170e8eae979e95cfe842551972b61fa7e2dd8
z202618e231f1009b36ef4782368c4c396710666197a055ce0b903e425164313326bcf70eed04b9
z6134c6a3df00beee67088af24bd685e65d9ebf4116bd8737a895d0312ca1873b5a2993e332841e
zfed39d9d5f987a10cfb303e9e5e17f0f96600350e5afebc0ec4e3f50ef6523b7d76409007b3bfa
z76fa641ea7ca0da8373607137505c82f63b40937537db8a247947603721a984fd1c7a0051fc43b
zb49cc03343c48c696a7ddebc4d5a0a6c1d3c1f10cca7b1306f6603ea71dc28666d51ff192e8de6
z245a40ea39f2c05232b8f0240ff2126f0321c1cd1bb008c8e8bd007df290eb1a1e4b95a18c2b03
z0fbbace20a1e6bd11e6dd3cd1e3009b45a4778d29090683d11de00a6526809867498fbbe71b9b2
ze8187fb6b59a0cc30660d14707b9710d961021bd683c9e38521152793711764fccecc69d9ca11d
z09cc2f631c1a7eabae11dba1c674bc5264b6cf2e5be713b6afbde839e8333ad5e5511e395172fd
z0ccfd8ddecd3f3666c04fb2a92e23d02a44a3d38bc67e84f7267efef8cac7c84a4b416eff1d029
ze13b5422fa4599d0e1296fcc9f7965b9686c5d10ec198dc98165933d15512896a71867b367fb4e
z6daa0ab99254d777161aac84a2377892f395a413361378fe13946ff3a9670cae5151866fb706e9
z83bc293b0b384ed5d619ff84f7af1108cd799256b59d7efd135ee6b318187ac1850c866c53c438
z2f9b272e1d24cdcf00a56b4b35b3f5721e3185490a0fecc8ab2ed158ce12cd5accc06f591d49e5
z38a962d3a77e6d5d0eb559746693e744dcd6c6c9d0cef92de4786382487e8ce3ce2353e0c62e2d
z51d36533008db1ac1d18d2b755fee9a044f0c2f7621997e307988a878f16d9c8a4994fa8da3a3b
z8ebd7b49e67a5e66904e1f31959da2a769075efa44066982f5dfd31b0553d63456c186668f33ed
zfe591c1b7becd00e6d4c8cee9a973690b99ef2364f55f44305de2fb6e2686ba001254c4b751db9
zfe601428969f635bf6657ad8b24feccea187fc57f4010a18352b74a33d4e971ba5cbd25dbcd637
zcb80705c64d868a8cc11a6541f52adee95fe8e0ce1e3d3f73db411a53ba33b55ea3ea743749482
z51e817820b2d7847345280b2e3c54945e43af5b9bb6d0fc1bfc00050a9159008cc50b0d67d206b
z02a87ebfa85b67cc023becede49b08ac60af27c44b1a22d444e3af31d2ce7d0281a631034383bf
zc6bf98631e254f8d7aa07270e5d7eb14989877c70381106c0b95dd141d12eb302f212e29de2eab
zd1c8c2f2ba3202f9c8aca8104bef40bd4f56c9f7e0a2a4ead1da4764b7b70c883ddd28199a5229
z8d3b8a98bbe461d7c310798a273b61cbd40e2eccb17b21c445f698667dc23414f5454fe67d18ee
z69c51ebdd585b43fcf79a999d3f5e4c72f34e8ba0f56ee11a027505c442407d131d3b5ecd285f4
zacb5b56cf54651f7c6eb55ba1faa591322f617a0d57593b18af7b568c6d8fd41234ac1095b3f96
z347651d9dfc970d16d8c61a995fcb7b27e68b30ff3ca6a000ba646b8420e81a542ec26abe452c4
ze64ecb1163ef1ba6a61a7196665c19079b2b21e21fd609a800d328d7f93a2f1299ed0559ebb12e
z339762651fe8f1a38d735ba864480988a66b349220650461b8ccd69804367f6f107b539ee43036
zed74710c7cf6c4b222c223c2d449658eb534bf0ffe712b940c12bdc63bb987bb5c9c72e044435e
zb1492d570549c39c0ab2c06082f6f4abdf3761b3cc77e07382529fd8d852c695b32571297538a0
z64ea2413309235d012395696581f083bdcd67e34e63286e7a433b8d932f505a784de46e869ef48
z13c37e9626e042cc48ee22210b6e17691642d00015fc281814c0a15ef532c0f9e496688a78fb56
zce32864d2e37b101c43ca37c847dea9798c9b60d6ad249032e0096f83dfc25f33cfcbf1f7f0949
z97b0b95da922898eaa8f3b660b213581189f381a753d33b1aae5bbe115e5ffe2672ec0ac0d9a3d
z91fc5118b8bd7e2828c4b979b0c1c6e83f6b126cbf3e23cfb3734bee3cb97d4866a07d14b860d4
z0ca7f5037bc3cc98ea2c1d00e0bde6841b22e86d5a6a6e671af11b1c38f63be28f8aaffc09a9b2
z89fab8cc1310cfc29e51ca39ea2fd1dbaceb6a195c5736f5171cdced0e2816106568357f7fd8fa
z54f7d081780789232225873ac4c3943aaee42e0afe80a4506fe9b2fc4414ac55cd9b7595a7f840
z9b5e42ef00d3922881dcf44b58fdce4cac9a96ce1c9037828062f32de45a24ec44359d3edb9bcf
z2c2efb386b7b12e9f3c1ca7e374eef657dcb954f3930cc8f035c6f1eacf7aaee88471dc082fb1c
z04f526cb807d70125ddbf0f4201562991c2a050c0f03d5530afa7f6e642db77ea121760dd5ea44
z616adedee62b12d241f5355176d55d206bd2610bdd1e862bc63d1f56f96212f9a657ada6cc6b23
zce73a1874a9fe6e490f5cbfb593f8755151ef3d7793fb802ab42790ab70c13fb85879dbbba5a8e
za29ac8e7ee32c432e42c152b964792cbdd2d2a5d563922c514f9f2e34607d09d5ff5cac916954e
z1f34715d6385d0eade5ecc72d6defe2c90034be43604fab2aa841e769246e63f307b6ea7b3dadc
za4e35e1b51e4b06c6dc88c48231c4a256415cf3ffe36c9f2920f1d34c0174fe5b64139678004e1
z0942cb0d55077958892f44af4d16d0a9eab6f6c90bf92b7251ac18b77623653e9c2fda5065afca
z596684bfba0dd8395072490e3fb3ec99f88fbe18809745c62976f798b7c8dd87aaf5ad5009f90c
z8579db9899f2495a0c25e35602f7fd6f382738cdcfb7b4cef6b68b5afa7a851d57251f22224a61
z953e44755289c61ee9652c94af86bcbed343a7eaa685017b9e2bc68f1b6d216f35964c801989a2
zed653a4ce197171a5554ea824a463f337ecd4b6af94445e5213167ddeeda3af1e9cc28b88ee353
z8bca1a6dcdd33a90f466363f7a167954caa36466a9b99020e80a25bc5e9e9ecb820e52de99fc32
ze95ea2e5c3a56cf8831b128813e6d55fb539b3c3a73c86ef1ae716b0b343c3c3469324373cb371
zc5e8d28414370da5cccadd07a23b14d2086768461b4c6d87a20041cb811f9540cb2df7cc871e19
z4a81bc19216cc695d7cec3179cee93fadc73395cc0081eedac7aa2380e23cd367704a58c400cf6
z4c8fb25647906bd8fb0fed91a45863fbedd8a47293584f3a65f408b7ce24694b5489637cb21224
z916d99eb9a97212393d4cbc0f6a36fc6daff37d583b1a60b56b5d5a6548c7ba73233c06425ed62
zcd6f00c78abb37b64876a7cf31ff668e6f7c1723877c517bbece92bfef3c6abba7926cbe69c09e
z3bd08dabc1e2ea42d323d9a13c6efa2066ce4fef62756ce5ce4fce67176b084cf73b32bf970586
z0c9d8e5318fe226fa0ed2caa4339b77f957ef85fe705d7f9e6a078b87cd68cc76a0a570b033719
z996cae67a340f033f1d215ffab8bbbcd2be547836ce02710aacf9bc73b34170ef8e2f01568a9d6
zf942b41123ef9011de394d4a781be3d8fb275ab1efd8273036b25a5c6e88c8f97975acf37a4041
z7ea31bc9c9998d053287e5a2ab5b9fdbb354a19e1274e53480346e67b8c11331b1ccfae1f31033
z900e16ca7e2cdbaba79b26e281e498f89c5cff3282bf0a0d43b00eef09fc242f0b779cd68498cd
z9eb0ad6eae847c9e4a67d5db35decb4a4c63903fb924a52147873ac40f4b7b41ab09b9221fd4c2
z8571cdd30d4e512309c6bc0c0b9bde75441f04c45d8cb8b3b0ca174b7db2835a4627f0ceceb8f5
z8236d3f8bd2d0e6d73502420fe639bcf82e330d67fc61c8cd6bb7376a643b81d9bc647e2248dc3
z03df6d1dc428d35a4631a1b6bbbc2da00113a98ecd7302873006c3aab693b4035535c6b5d9d0fc
z1a5ade96fa8488091884d13d9658b32dffccf7a33114e9557f0973132943e68fb5f5f05226845f
z00f265a6f604c1dc80ff86e8ed6868ce884a1b20b2ce2284a79cb8253de94147f996fa8a783418
zdf632ae8fee13c6438f8a2e49e6617cfc9a0381f1ce759a5b95a98e573e018ee3f9160f5a00eeb
zff1495f6dfc7f1b983fe8ef317cf3eb000b7d9ac6043000ee7cd410e054371addd9219544cf807
z20d72b8734683d42be4ab8768eb3a90dcfb272f929b6c602e1b894220ce16bddc4f621e5564cdb
z0c5df5cb4e596d2fd54e6039a38aeb59ad30082e4f936c502ae188158b959ed456c7f543fcdac0
zf5a9fa53fbc3ade99f65e9f9cafe44a9936ed711820f267537c46f47f9587a495cf05fb065fac6
z95a9f2c30fef9b72783a0eead6cb68f8cbb67e38ae4e23ef6282f128fdbeee926a78b2e7806dd3
z96e72726cc8404fadbbf78c9638156c97c6f4e4c0e54b775f9f235c2b002e60e6900c93ab170c9
z6354877a9fccac319b1fc85c308da7add40a18a194434a6255ffab6440e578408264775afcf988
zbfce1e8afa0ca6a9cb7adc1cb1e10f02fe965ca86a93c8bf0ccc073123c95fd44731f3123b5995
z10571056798f2e89fb051291731f208fefa0a5ab68a3b00f8b4399e4a4a368fa94d74174d3da2e
zee1da455df1c99234633d16a536f6bbfbbc59c778816273c88d9d3499a6c0ed308cb3c4b9516a8
zd2a15b25113876f7bf57c152d6e10ceb48b1f38401fd0f78274ba0d77d698f8b3e40c8d810e422
zc6045660ef8fde1bb6b0b4519fb3768acbe81fcd6fe071ffbff9099e2bd7cf7d56b8cadc498c74
zeb79c635220ab9ca7cb151edad9dadddea8255af35e013699a28dcedf9340f4fc8ffe6141d91fd
zf739910f2f5b731bb7ea74c55bb14fcf5d4a94ae327e055954a78496a73e14585aa79d4a69e916
zfaf970d7dd43813d6602596a7041e1f569bc6dde4f099591b4e4d3c5ef76d038e78bcb4f14056b
zb548cb1239cffb42c08646e41b8c1a667869276cabc6d98025aadd660fdd61ddb2695508144baa
zd7986b50a6844ed75dfbd1fa8b8d33d9baa831abeb68bbc6f3fc6f7bacf6602eeb630b62de13dd
z88a2970a9c081de1155a6ec6ddf079c872588a233143946e5201d16578acc3b873b19a3d31e7f7
z113cd636ad658e3aadf9b30e4ece4bff2ff81efb45a3e6acaf00a0ddb39c974b5d5a2c7d668693
z52c56a3dbc3c6a02d8acb7f9e8a70e8096345c6531f6dffb32500aec4040bcbfa464d81551af2d
zc4c4d062a8424ecfd8bf776f9e7fa3281f6962ca19fb6e02f5127ee07cf869c3e023ed9a5c1916
zb1d8d7c136ca5c0f8a73ba169d65304d8d625d7b272ba8eb6b0f2b465a402dfe6880877353a1bf
z7dbcc4cb8ecb57f2ee41aa2af554ea01470968a46ba5fb68cb20d21536edfe1061638739174d10
zdaf099d933b532b95a976247dbcdc8e91d6528d1751719212ee8bda404a90b72f465527f8079ec
z467a4cdf649d117567d595c06768567e98695f6bc354cd2c2a92a03f5522f77f424cba6126887a
zaf38ac07b4212d0342e6dd767f01da61e9498d281e4c9bc3d6236c701507623382f8b7519c652b
z18c7a2c1ad1a1f159009ab96b7a7c966de6d4c5b86438afaba9d232738db6e5b03ad9d9b57380a
zde51e200857831fb624852611e2bdcfe89e75fc0c7c78a530694d3730c7e7eec636e97f35417b5
z2b2531f44856ad51352afe3b530f5ae81cb1d916dbc9d85f081eeeaeaa9394817b0edbee417eb2
z9c92e43a3fa98f18faf456b75cf6e7c7340f71e0ceed6d1d419eab39f800686a154e76fe7f4764
z2305cda82e123679f08d255aac2fa70da9e31f25edc7b7b82a0fb8c0a34a6b6ecd3da9e67d4a10
z7685acab8c0fcc060b1997a961ce1007e4562dd61976a42fde4023d9d61a908982eb1d60af8f39
z8aa36feaaaca48981b324c5d70c72f2d28de9ab4f3388e7487ecf9e3a2013115a7716d436cfe83
ze497373e4d3f83f1ce84cfb06b9f51fa6f8d2a865a381ef34f29dc743c97f6972e1a85eac569c5
z53e58d5e4c0a32ede1169789a06ea0303db2ed0aa36153846ba795bf74a43234ae10aea435c924
z7633be9cc71e09a94ae2d35b1286d3af21765fe7be669a6667df01eaee02ce5a7c54ef7dd3b34c
za81466f3d56827bdc75cdfec536ceea04c08e71ba173270b346159bd1ea23ef1886226247c6c2d
z14ced4df18c24df2bb2aaf23fc521bd23bd411c206341d84b94a8c49a1e3cee1056030d4cf9d5b
zcbf11869aed174d838f1f180024b097d063c1c8d85a9b74d53f82382681a6a900e84ec67bf24b8
zc31aecd10c7fdab66a832b95452f0f44f1686a8857c24e6f6c396cde67d0a0bae0d1bba5fa3366
z1bcf164511a9386943819e70f541b48e14c9e5a810a0da1f0e68aea45a6f461ddabdfc2dcf5a73
z2bd561b32aa4330f484d57cf88c1556282df00672775bdd0a3030416955e28109e596bc720af46
z1398a91f7027c304fd63e646fde6324ab2e6200969c53a2531206c55b4a1968bd404094809689d
zf64d76cd568dda22b0efe010ba5ec81fe772367c099ae791ba76bc44f350f353c766dd3cd9ac49
z1684a370655b56053da201573c2bb5280dcfd50036c65a42da6b6526599ce7290a823c91b82f3b
zf64fe9678af658ce81ebedce2642903aec956f68302222ee38c7d9e87cbc55d2afc394b8f2530d
zcc1d7ecd4cca617de0363f24e3ed81cde456936fd6c701ef6b1ec7bb8fca640993d512f3f6f525
z1e98aee9eab9c718447f625d3200b173c20a929ebee4aaafcdb1149e0c3597a4d2c954ad109da2
za0e54768b75b7e507702acc8dafe4886e2dba15b8b3fc23bc42e22902ad2625a297319c7aae66e
z67aaa2e4193ea430af61e0ce1c93bbae07814c7beaab2f598b559f57c0e90096d2af5c7edae2b2
ze37370eab10a7540694895537bc494278e10d7a5db65b1c382d706064a52244e6046af6cfde604
z8ecec16498060492ebea0f3d40e706a47372c26a44c9f54a3e04a096883cec2826b3fdbd48a2f8
z9fe9a07c8f471d38233256ae0eb4057b0ae7f24b75237f93747d662a8c86c3367a65013d25d99b
zff2bda09e3a66b80dc34adbd4d65ec73a29a5c36fba2a84005dd5acfbf9dd4aeafa4e1f8998eff
zf286565afa6aabc127436e29b5577a87826a3a0b4067c688e43ca719507fcdaf6ce8573fc95096
z47b0d1d2f193fd0752808d12a11d36805983745d8cfb9be47562f85bb49e7387790c125c32f345
z72734c351587df8604e45b505d8579b70d38017c2f5283f812e981295b070387b76a4c6bf0b18a
z04a6964b4b4d6480cbfc1621d29fbec8861412a60864a71e559b2dec57269b19a091978e7546b0
zae514a3dc6473bb4443f170d0dd2ab5b13eb6ef1c9b4ce6d1a272961aeb8481dddcf4db138bab3
z6bb5133b7800ee6e72a812401f558a9900992b9ad15fbfabbab694fcf3bc05d7b4f7682e107866
z4553c5cc6e2040179efe12d21a2cff27d13c3ae5236508424156ec58cb639cbf5d60a0b700bb82
zc24c9a04068f8ba9f3b92215dcea69a5d22e0b525e53569a4d563ef3c6c34dba7cc8975c609985
z262280cbb078d106402a287549d1bda8676bca872668859baf93df747e3ac25187ad93371d3a14
zafc2570cfc597e1eea7ec1717dc49a00f0394de5acf1b8bb976ecb33c548ea5799a322722d6d67
z787b77d4b467d547cf0ae281a208698a2eb46c94f3c0469c63c7c928c973a33fb2ff0d02516ec0
z70be31223ca8dc3efdfdf600b0ea3823de1a13195486b82c1bcf5b35dfaa163ad154fb6dbbaab7
z8dd2e891f47d1fe52eee7ecfebf63a83cc2c21e295a76240acb30b27b9abc199626b78a946c036
zad8f63d6cb7b8a69070dc43d7ae1719ca84b312ccc1a40863d3414e3642df3a01f47bc747eb095
z1a84a67b938fe7dd04adf84ae0af336640274b5f2c10c0cc51a8ca18a9576c127adb85c331465c
za8ef9c2730474d43bdb061b5b17595536015ebac140b0155c724cb9a8bfd9d7e16a5b7543cd55c
zb90706a02320186377ca69ff24a1d17038d71f879eb0d0598bc43689134b53775f8b2b975d3d82
z434ae3e4a4c16731c39ced75747620fd20f93be9644fe3d35de87623c18e89b37cfb6bd1272a42
z2bcc49ccc8b453daefb4f5156d67fcc0a9f80e11a56955fb3d01e24ddd3cdba323de0d5c711bb6
z18d6a9070feb123cd2b5f1e3a0a764e490c6431dcef744a033dc860fb04278666d78178e0bd1b0
z202b6d997b68ea501aaad738c713689454472bcc2791039d7e317ec0f29d89509442acda218895
zb72eee57ba311cb66ae4208a40831589e5bb9c6147feddd6a4aafcb879635feb3467e8332751ab
z352ac9ab86cf7c06dcc458f41809f21e7fb1d73622e5f6049e5765d2861dafcdd07292c56f6d3d
z01a09fc0b1ae872f98042c6a126b542e20aba414eb9126700d606a0c1716f7cd881bf73b4af2fc
z69c89dfbe055cd4e98580b635535de9e3c7a7b0faf2cae21f298fde4614137699b9f96a6df833d
z4c2ad1116e855a161094559be019db9e0b5aa4017945d3fb466994f2b719367cd8eaf48dc3edea
za64b7321cea01175bbdb1b9905fc8254484cc9bccf2dc9ec1c78e64f42769d31bad1b44bd62d5c
zb9e7265e82b86c9d5ce4b11ebe700181a762bf52220aef16cda1f9db5dd662091f43d6aecf73c3
z12cfb10d752b1d0cc40046f5118253f1826597ee5ff61553e3229eee6d4774faf0b642312eb5e6
z587dc571aa0afe3f2451fd3d0e13c23f8b9963e43c773ae8390860e902938fd1027d3b0d5319f0
za3a2d97db832ed0d42bc81c0d21f7cd2e82f1733d372726c9d31e7e824bc015a29d0378aab8a5d
z51c31673ac512387a391bba63de718d3d0a4437c9f29cfcfef0a5a8169233491708168910447e8
z91eb4249b3d50bc5a1e4191f04497146ff8282b7c4871513461654de151264005818990905b11a
zd7a9b324b492430459b7e9119dd47297f5751c9f888a175caaca723e8f8d9727593129484402a2
z07ebbd6bb12c85c9ededdda7c3bf7203178273da74ee1d5a4c4c1f3cdae601723c04365255fcd2
z3cfeacec70703658e069d5a2b2b44af50459445df16438dd0bc60c09bbcb9982ae06a15c07d036
z0bb5d1959bf2b8c262064f26e414a6339fec952ce8cedf335485ef7fd0beb2d7e646c77bc7aa5a
z4d2f1737aed0fd5c7165a8388d1616c216abd6c4762fd00dd0f23a4421123758cace3967583806
z3f60a6bceab1a4c8954204ae30ef28adbc62f1101ccc2d910af06090e18fef2de2c543f903b9d1
z02d10e3b2f42f3ef2eed8f146ffc93b6fc61dbd689ab26f0db7fd5b452ebb8a3ac70c5779ecbd2
z0e051c3c68627db4d71aec7f9641b56fa769fbda8462de7520496b73e258f472a2f5339fe6bf73
z9b6c8d9c6d6231b93cecb31ba17b3946b6ed18f8d3cbd4a3505c3a8ec30c405c580fb44f1ef316
z08f9d73457fbd2a6ce89caff0676492dfb55cd431ce61058c6759f630c6d96ebbc595ba88c51b6
z25a9b97a0b13ded9cadb7c94bb7483a095469533be5f53a87445b95e9fdc5c1cdf1aeb6fbd608a
z4df2ff5d73534b7de6c828fb3bbb0ee6d126eca86adf3c9aaaadd4deb77cc08c025124e9e44c63
z2fc25aadf51bb92d0a3612f47abc8307a220a612c257388dba86c62bc0f67fa80ef21bc044d43a
z685d32006c64381f6b25d352f14b86b1aa6aee7325f4210b549f6fdf87927d4b701765b36d7aa0
zdefd2faf39bcc05fd8cdfec2b263e9c080a54c42aed0715c8429ca2765213e33da7fd4a7096701
zc47068028a26d3d7114cde8fab37e5e6ec0e00c418b5ca6c161cefdfa987d9922f810a617ff6bb
z82e1f5b862412ed6e5060fa75d2a5f9f50b44c2574ccbb01e332d6778be79ba33fab3612ae618e
zebc000cc334694b57ef12879edcc0309e08f46341b462651dfa399a052f2a03e9659e493738428
zc7c313e7f81904a0b060754785d0a5bedab6b44c5d7b6f05fde14927167faa5fc0a6e0baa57dc3
z6ccc7ce57c08075dbeaafbf4088d626d7e397ca2fa483eeb2615147bf2fd3a9062d346b623ace3
zc0d6e0fe2f05bf0c8b5bca6c1ab2aac005bc3e235a33ffd3395427c11604efbeb0155783a68b01
zf3e1bdc64d9b7af0bc7f5cd61c40dcc4400f2915f4a2026a6c49544a863ff6beb1dcf4d5368b86
zd166c1da0fa65b0b52ac69fd1a82af7bd109832ddef31f66a7fde514ecf9019c686315956cbf8f
z61de5beb17f9a768c04e3bcff435df142d123df6921d420ef36c97a52eec959c656c7d7ac2f20e
z994d526df7850c4ee8367f1ea9613504504f03f37275c18681a74eb3bb061769554f127aa12388
zd67a10f531adf2b8c3df300f622120d4a01eee657c870d1d55c0328e8f59ada5c75b8b6fe2d55e
z308e0d7674840f44f86be76f5ca00bc2ff3302cfa0a11e474a783c0aea34862ca3b3cc955645cd
zbad6d8b35c4793521db5ba77c05442f9776bf29d979959e6e618eba46a6617590b45b75f22dc66
z4784bd18554a3b58b49c4520c5e4e553aae43427474de1a76cbe5a60d0d9e347a1d6a66a2264a9
z7ca1f544166b6d7e0c11be7bc9ea9857d9164c7eaca12d4c71d8f574feb8a94ab810fa994bd306
z54fb2c22e8eabee9b4a6cb5d36646c535d38fa22b330cd607aa588c35c3e47830d42b61715ce95
zfc2848848778014842a864a55569b29ac770c9208e58874c58e3c9ee64493cce9cba6704e5245f
zcaeb0418459d842caadf694b8ebf4ddac374e3450741cd10332cabc8b94895f46deed0af52f98c
z9e2f1afc66a9de2b0cf0da57b428836a4b45d7638d04dfa526a2ee1da5d7075d014bde1169e424
z5b2b3264f7f38bcc835e4f3633ebf3dcd8e7927245d4abaa5431664dd23f3fffbacacff610af12
z6f9f1766376085eddc0973396ae02c812ab64ae8dd7e17dc2213014336204a9174b4ceb0e48705
zd0ea94c6e11af3073e132533ca0c18379fcdaf723d74d7d0de41f59dc4f0ad34c2f64ea7412688
z499ade81956f7ff78b184f8af659e9a60badc522df4615ebdd7160aeba38be0520892df2d8e380
ze073ab345436c5ce627b9d0a72ddae52f5ec182398af6c6bb5938d15c42d4f2ce22df28dd6d3f0
z7dcbd9cd5265d317f9f90e265e005990ca6e4e4f44941839dc0d7065c2502c11f443dd9a1551ef
z476e0e359959ce89e8a121cb6f6aeb5b1227eb832e32fbce10d89a92a42ad07af96f0cedb7fd21
zf0cc32585b0262356f225fc50ba8422572567bf2b86bd80f608dd7649a9a5240687149c3318d99
z0a5724b93834d2690fb141cabc0ebc64c0144d6ca61add101bbf3642e85bc814c0a5f6637915f0
z7ba7973207fd863013020fddba3c91c92cee45bb621ccb3868756bb8fed917f4bb2c55244547ae
z91536e710ef1b8376820f77ad2574771041479182b1d1074688bd9fdb7ea17a4c917c60030e988
zfaae368f3e1096000d1135712042c59ed334d7bae51381516e1197f15827e90d26d3e277e0fc71
zb2345649cf8af6445e7227a4d8e58acdf656b4be8aa68a887d282d7b7d16ac52722afd8e2b33c7
z24c244317e6193c9e946edd6d39c0d8ec41d0d299a1e960911324c2f8e0a82e7f7046b0c44531f
z6e878b4ebf9b2d2deff6ac569b9949baa97fb7086881d635b4c21f973007e4671c91336862fb27
z922892e44f571b528b6d7d14df8771b1732d4bdb15dc1c295f356dd9436761d897612354764dd3
z68269cbe5ed8d495fa36a3d887ec33c465d5133f863410928dfe5b8131b1dd6870445212e4cabc
z6a8e48d23eedd8d4a936e5cb4f911adbdacc20b4bc5ae64ed87ea59a1b802634f12f7aec15839d
z67fdef30ea4dae459689e7a72bfb3dd26eaad9bdf88692e126edab3fd2c3b00c430b5ff3b7c00e
zf8da0852cd9087a1c3d6f6eaf1a9e4d93c471648c83e1a77ab51b46ae33e5dd038517f312aa667
zabb3c286ecd8b023975351cdc370d061130df64e07fd6876573927675ba1130d828c3c8c078c43
z250f92695f98831ba1a1a2c0cf25b7ed4c51cb11cd01b32827879b421a39be9263f18328aa04d2
z7b7267c33995d0897a12aec1c8efb90068770be573e8fe61ad0280e6400814d4e275e3695ef08f
z3cdc77af78397c22d467d567621b7e6b52716e6367958c1cccf26dc99cf59eaf44a43569178a37
zbb83c2d853acd403ac5fd4a82d8046679c0215b08a24ecccd163c191437d4159fc83fab10ed369
zd99f40c0aaa8590fca679e6d23bb2fc11475f92ae7534b1783047330109004e1d7e756f530d15a
zb6ffada566249a2b21a48d3f690489df5c778ab2d5fd8a77fe7d8a7129d8961abbd259449c95b9
z069627adb85d05e0e0afe2d2c89ec97fb06ba4daf09e388f2359f47cfeabb06503c6c50d7f6749
zbd380fca22d2ca1da3bff27047cf1bd4facdba7f2ed42c4f236c7bcafdaefc3058a83636ec1ae7
zf5340b0de4e3d98e4e61c498ee7c4d6da9fe2b7cee63c99ec26a72ef6179ac4444029f3b27aef0
z25652f8cc64eca928e50987fa9c3d65be76b965f0630f2cc2cbdf9c4492400a7cad7cf922790d7
zec4f5fa578ebe5bd7aa3740c642580f459f98699ee55ce8686601ad5fe1fab001441e016adf2cb
za55946a60c7961351d98b3ca34787e953c5aa0888f187dc78add42be07fe17972f92dd51f75bdb
zbf60c5b636f8ea08dd0e2a69e13ed3060ce4c65b0b287a6e6d6a5715a2a37d26908d68811485ba
z62b01d19bdd112446e8ea9ec56cfcc985993c8f10c880ffa542d48b7a8fa575c74136dfb18bc1e
za4a6713898a47bceed0551822cf64f44b2003456b0185e4bfb61d61c45bb49560b193ce7679432
zf6c12811ccb598ac00bf96ff84cda8e982787cee560018153683063babf5ca1311878733e24533
z65c6f8f3caef50965c76fec516ba125dffd65904713ff0a69636e8b0f00bba2e8c310dadcbd5d1
za44e8b820788bcb27ddb0ca2c42b724af93ecfd46e8878f092fca5574abc3ff2a6d249782f884f
z291a4354b283251f0f4571f12599d645e49df9831d790e2831a48da09179eeb8a4db3da2244d6e
z95f8030c2496b0a96aedf9792adc2c57d083c1a30c1ef3d78fd4ce21ec9635797a69817c77ceac
zd0bfd5978c9868b26338112fa73887474180dff65af8c4b3a3a83b334af6773865dc4ead42d325
z436bc0044ddd57a0091d8bb0c80bd948a0ff929ea82fecb2515d7ec932918051b867e05c56ce6e
z7cfbd6d56ab8c0ef273b05240a9a2e710cbc501f5df7936f6096e8b164a9b634cea2a00590bccd
z68ac02e1a40cfadf2fb3ce98a73b88d343977d0cceb9c3bd0ec6dba2f0bcad694ab9eb108922e8
z86b3d9f6ac6988958106315b79088fc6e79c2a69e4a6c1268d03cfe88a73107023d8f7e4e23519
zdcbc5e00bfd145b7f22c95de70ba9afdfb44dcfd08d51ac7cc3fa5d4a958b0a744f1b397c25007
zb469d149dd49f89dd71d468dfa52926f9a376c80e89fda48d1f2b2c75b45f86da640fb324b48a7
z5b89efa182fcfaff2ea6d1beec93c3d3ff2a0774bf8ab29da4178949ddb0976ddc93dd7c901697
zeeaac86a74d766cb4b806d95fe06866db2e0e118600c90cfae9978e0cb9fcd34636c2aa8b69078
zc7f8d24899dd000beb4f6514cc9751a22bc0c20749b7708cc02cfd619c17240cacd7f1e1204bd7
z22d01f08425c3a7161ca2af92c2afbd8575c0e6f2e018c0fb569a1ce555650b0922f6ab7a4cf22
zc5e7aada6f5c8f369f6e7d0f25a489a254f3f23fc1834f165c58d999dccc67fe82797f1e33aa87
z972d4f7a99583cc5ca3cbf1c673cbdff130509970cd5734b9621354d3f09d300ad26d8e3a3e06b
zc36ab91b3bc4a8b8a1d5e3d821a38306862306888bf604e4b90656f2f504b3578659d2ff82df82
zf0e695669df0a27b660dadbc778a942549edba6cec3c4e403a4999fb9125c3501f3690941e937f
z04250630cf75b5fcdba1bb7bc5068521cc2f7af7383603b9d3642e9cd9a1666692356e3a34f63d
zfdabe0fa7c9684f4fd2f3eff28ef780123e60e1ff6e1c6feeafda07512af9809e2813af2390cfe
z35a59c2e854e6a42b451c49dee5fe6def2e40d2196c20e18865aefc5b4874101760d2c9459b9c2
z77967ae792abf665280bb83c2ec571b8a19e7fa08c0b4de35afc809b1e612c516467e89d93737c
z4836092baca755198508b6accde5c82f426581b9fa058b2adf725d03b6c98939d6518f0dae281d
z693f52d2d5d713dd161e5ae16c9c46a1c0ca1657f357a88105e772433aa9e1939c505b1e79d5c5
z64511a19674cef9a91c47cb6125a7740210c5cb07dc33255eb395dd7e83868206d277f264e21da
zbeb85e1488b1aaec5feec0448b1a800785a603a0fc5d9eea891bc1d5e85e32fe0f91de837fecde
zc6e7b072d82ec709d247978b0363c37147162d6821d62b30f9d05938c56e2f89345043033b31fc
z2b7911e0249bf93941b4b502813bcb709c334e89e67151b90936b97ddfda35a15951ee73116a35
zb6c92ec6f395613cfc1f0a9d46aae57764ce5570cef94503a11787c97ae571bcd8dccf6a0efb05
z41d52b294fc84dd0f00da0f90d1e4a55be127a748bb1d95e56deb122138947a17fe3b3c4e7b4b4
za01448ddfff5315726d8445eb25aeebd300a07ccb8db59c38d70dc0e5720415d0d263a091e6baf
z3ef8b3721887451ba71fd23f3834833d610e64df05260b31d5e571a79830c695b41bf97e38c271
z38d2b90b7a41dbde5ea82de7d06289c0d4817a828ee2915f07fd60dd9900fe5c3e9582a4d81ddd
z9262151ab145818a3837569da0787e30472100585051bce987edf045698b59454dedab8c7cb3c1
za6402f6303312493cc35be57984a5a35e117e3047d370bcb419d767d5f231fb59e6ac55fd680e2
z87145eef1547a7bb99c5a360a1808b91fb21c106974cf45716a4e6d14587fefaab62d07229f8a6
z3a6dcaffb8f3d9ceb4db1e46f1898eddcbd751a84633e029e44169837d97e2dc38148239a8128e
z42da80996a83ada200f4681f3ad791c0b86f22364e30adee7053d40e2289c595564d4bf9cef70a
z5019216fb928b39c8c7ad1e6766a13ad64249e7de5d1ba90d61b995e820bd107d0e6055312dede
z5d43f0662254ee91135ead5922558d331ad9becc382c12023e4fbdfc293b8c44698866d2465ad2
zcffe3a1c41122667c6c041154238ad5ed16b797a91ed935b7f85dc6b8bc47c02522588acbc10cc
z6e1af2b401f61060e7612c75ad9c8d2a777e41d65c2edd442c51cc8b92f8c0d09d528a3ee84063
zd5572185618980fdecf7473302cc3d4a2613dfccd39b00c65cfcb36cc29a8bcc4936b26eb04d2f
z21e8adc95ce1eb1b9eb15509ab3ee9d753147b929ea3af2a1b26ca4e750bc7fc3b0b3359c63eda
zd5172febd89ad905cba060e86a2025ea77b8f8dde83d4888b5bd28a45a5640b65bf9ddb17dc038
zd52e806c66196fbdf0848c13d708d332eefe30f89bcd056bdc8b94b2932a7d2c5be2745a50e066
z834cfe9483a0ae7d012c9b29b41e5d8031952f3d124cad11d2387696ac1926d6223476d801d6ef
z4d547e16c32c193c967d11543e1dcf264e55d1fdce23c6debf74fd39ed9c9dcccf43a0e799e254
z3dd361a9b77430e2a6773649e9fb5749a8c604dc3579934d9ee545787e7262d815bf40ed21c9e4
zb3b657546d6abb6a1310763088e83c145ca0d8d3036ed3ebb86124c99c55a0a7d93c3214e5028d
zd489b6eb932211573dd01e16a816ab25da1bfb3c5d5e7cf17060485705740863ad0f72a7e9f861
za5cf063e834d94662027604fafa803bbb06af4746385f23bac4118b745f399a777d2e787f8dea7
z6d2136d545b46da0f9553f13199c45e2a49284dfa44bc0dcafb3bab3fab4729c8bee52309f0407
zc68e6cfca2505d5bd07b71a32f4400214998b4a3cabb108ff885902c0f44daf499d72c02603416
z0634044198742d42f24693f82d52dd7dc8972871de72ab83969502b2e00d81f80e92d29e805c5e
zdf1b7bcd8afd7d434561d97b5faaf81c23c88e0e0be2a813223bf0b8b052f0cebfd4730a0b5d0e
zffc4f257edcc91497739da5bcb33149a5951fe4fee120e128fd1da6139b4f41c13325fca2f3147
z3316c92b9623b4110e3a7a89ebb6c8976e13aae5b34a95448a5e56c6c0c2bfe87eaa1b477fc28e
zcc830880b038946aa5121d9c8a292edba50eb13a4fddb6e68e91d482f45fcfbafa46c472f2b0bc
z7fa1589092318c1709646bacd0c544c76b0e41730fa6b98edd4d1103ed099bd607747ce11d5791
zde1af02ed948eeb897f1829161f4ffff4b61590275c4122aca5e3466fa891093470607911fe362
z767057a16835daede73deb1c69e56c35ca3550292d1fd36a073d003d459f625caf3c8db3fefb32
zef5d80420fcdf3eac57f19d3875aad7318516ce0b461d0f1b98101d5455ad05c471d3d41925426
zd8c3bfc75ec525b3fb7324d8af717b1d4df94ef405d9271e7ff3ff55f13ad6ffd9f143768eb52f
zb1824329aa9b2c28d94eab2656dd9bd27e95b896d273d78f02cd57400f84d473e306214e08e614
z94e5357379074a86cce2ee337b9fcbcbc1528dc9c7fa541d7d72f138506fdf95c0af84a1dc5caa
z7ea1f52677a13139987f2b8dd1508426a4f23cd853f902c9c2b9d7eaae2e24a136e446058719d0
z3c2c2b41debc7135dc189b0b5e44947d2b6f71ca319e8ff6309752bb1d90ca1aa173b9a727157d
z6bb709ffa82a55b7ca178452102e166c4bf26f9817e0cae5d07559e85099606e62b163310a25e4
ze68d4a6c140798f81777235d2d7c9302fc6581a25d2b200f0bb46bd890e677507c4641e8790dbb
z23ab34fac38c87f3651aab37794bde25363f7729cfa4a6d1dea3d9c2293fe7ea3a9b7707f27495
zdcb217dbd43dac8f3e1a53d125101e158d08a30d5c135aaa92a70e7b804142d0b6c747ac8e8fd2
z5838f495225ee712e65c7c9df235c0a484ea07976247379674dfe72e948e6b44b6bbf73531e0c4
z9e498c0a894c6f946992e676cbdf4cc517e31c2d25bc022c101fc80feb6078648011523ffb217f
ze76be68746f3a2e933233168d22729a068d103489ad0f924615b7a28856cca9fda698ec091c716
z5fa21d08e7b781bb8cdb44b5fc2bb4538238daebbae35d27d8cf7a1711aafffb290ff058501161
zc5b97d1a9e6c5d921a51837a8c92df0ad27f76a78f7bd2cef2b2de7e12b5d3e7e34394c2a83dd2
z509c375a13365c83f61048a62fff3300bf8cc62d34f8d2150f48542307a3d3fcbe926a33c8e139
z48e5d138bcca55e10681575062d915460d37456279cfcfcc7ff77de068c4641bb45cf224f5f2aa
z3b26b3dc2500b2a767c9f4a216a85df29c5853243266ececbed64f141c4aea3530d4995c7051c6
zdcba02fd36ceb5adc8191a24929e9c764f8c78f16ba14b9075049282cfca8c7394b90f0b6cfba3
zaea72763b96dd9be589921993cdbd5fba534aac6b2f1a6829b85f840f14e5ab68f45853660241a
za7a04c1a433c648bbf5090e131656124263dd1784482f2bae5adcb2cedd50953928ff3ae2a8d22
z076511b47c975e53929e65c4d3c9b5ace630e8307df7949dc2bfa3ceed122e6a4526ab9fb70f2e
zc0414c2b32344131ce3aa5060c92dff71fb392abaac911f5e2212cc49230975b441d861e2302b1
z43136bb7a3c8d08f7ae940111927fc5fa469d753eb7892d14d05354b6beba35fda6aff074893d0
zb21b49262fbae8c7f32351cbb0df908162199fbdc8181d0819b20a395fde6276f3445ba9c03f8e
zb25be0b68169584b95691b27c8e1ed09b4acab9f5e424109543bb1567713d06c478e7a89954d99
zcd0bd8b0bff5f11bc6f4a56f8084cf78fe6ca85831b7111b68684a1a8d848a1d0c0264514217f0
z044f084e80c5b2866cbbc70d9a35c9d823488a4fd54fd668801db28282741c0c6633325d924873
zb23d56bf7243b5edcc7d1578bf2a942a4f069f20b1802dc7650d2e9935b1ff88a9d068706b8f9c
z3e5fc491932a226876aee449d337e353dcd929e1028d4bb8eaa010099e910ea4b390ca5b1b3d2a
zc30dfca898c43f43ad051ae4651a384332b28ac1949801b1228557ceac2b437441f80d64c686b9
z75fecbc74390e3c37dd4f0292adb4651fe64e06fdd2b2f884bff5f57859066c0974af9a22bd9a8
z2b988b7af47e758c35a5ec1f35f48de65fb6ea8bda6193dec750a98aacff5bc519f6b4812e39bd
zc7b89b5320c8aa20b30e382a52d8b4eb15244edc46181c9c3c21913f374af668925cb7ba68ffd2
z1be9691792b444a42ea592202f1c465ea78178fea9dc589dc39fc654486952a5bc70641837ea7a
z53ee0518809166307ae420c7ec1cfbec64c0d056fc58802503deae53b6bfdf9aeb62fd8704f5c1
z5670a0aab7352881f2448d3a068c80f51c881f05789f30cfaef482eb7cf664a76304b511bcc059
zbe99ca92cad4267bbe2cb7c10375ff2184f72871e8e1a6d5c6ceaec40e44afb905da652db1c28a
zd836a45629166d64dd08533f66ee16b723d8ec21ac651e0c802a7a0242628cd3b98ae20470d3de
z18d75ae08cf68cba5f08d6afb9d86b7b9cc15d3b86258e928c866575b60299b5b91c07618f5bf4
z4224ac7caa644873ccc1696bb335344eb09379c021bb351a8179b4311eaa29ec26fbcb1f924c5b
zd44df67433dfc21d30f317e170eba3723d532c439f6f6c5493be570e10e9f7a2ecee64f07d4dac
za9a409128715273302a0cddb3b5c7beb8cd38b72ca626508c7f21ce9307fe6421a85964db31e32
z36ed04ecbd7a4a29b628342cde9c86049a4f14661dcfc58aeb4bacf6b8c4f932ebbef445070f20
z09133c896078ed48fdcb644c115023f41b0308997cac2c2247ee41f3ede04905c1f1f9b84b8b5c
z925ba3f58826fcff50b7672ddb4da1177ca4d366c609451f85493c92518bdd8398609c2cd57105
z4a49187f9dc6d306d07dd2a3cf5e95229b928ddce0abfccc73d88095ed8507cb38d8a00d3fad99
z4145b7c509722e42d1fd795a0b9dd5567d6ecabd71df48bfbe4f11d8cda46b61782bba855be88c
z95523d88e95aaa23583a4e475d6e15eeab817d1fe95e96b711423e6b89d3582872d6b868e3fd69
z93bf4edd5606ab01225329f102f5dd4872f9a226f87b4a06989c5ff43f939d6998ad0494c1044c
z6af0db35ec13f861083034d4723898fe29363f057ece40561608ad0049ed951749028115cd61f6
z57b500823142681262145fb3e319a5d3b04882ab54e220acd3e44a885b8dca47ad7a9c317b9f86
z2b9da66ebd5e3e62791fbe0bb633a44862a41818879cf9d12c4ffa3d296c1347586154002041db
z2f6a7c3d4b620248ec24ac6e62238b5ceb2f0e9e6c4df7acc286b5517adba1ae6ca01ff2a43941
zd6a5da1e150fbf946485df9ae8471b11262016f6e3acf551789028e2dea61ec1c8a68b0d4171c7
z158a59f6bdc685a3add87108873d5bd4d982868ececd3f3427f92ef21925430d720837a650311d
z56eb6c4bb4a41b5deff235bc18ff9f365530072aca8f3d6e7dbf66ee5ec6c7b86d563d55c12b92
z21c636229863564d2aa6431670c5c27f2c5851ca197728b4736057ce269487e722473a6797d027
z60e50d4cfb637320efedbf59f5568122bd361f4541461355fac2c80b434e43df67ae8f2bdfbc3c
z47baa61c812e1e461f83d8157482ce745c67f48362443cf89522e6df056d2f107aba6a0080c384
z8f031d2845e909843b537ff59ee372e8d92da9becad439c958eb433b593faca2ab4e50ba7ea5ae
ze6abfc0c0abdcf8990f2741f9e4d77d2e78375625629de1f7f0221bde4b732dc5dc70724eeaaa6
z4af2675486bc2aba4f1276047cef69b2a9a436a03e157becc6ad4f2342d320d832ee523e538e3d
z9748708594a554c9ad3f9f1a5c44ced3364b8aec78a3f172c2fefb5f8e49e3f82592a88864fbac
zd168c1ff4d1cf96832285458759c7928c17e05f9c94ac4acb2c4785434bdb07128abfdc3f2fc28
zc19ab87d08a8f130a741c0ee6426ada7272f310bd3204e30746e1c2ebf155f64a1482cfc1206d5
ze5fb0058cafbf5fbc7cf4be176dbc5bad141990c4c658df3fc82e6c541765716d8b8b62c3d2108
z9727dc519b3bf0f7edffa06da3fc763598ce9f077cafbc9055013b7bba17f23d8274aa7ad7c6eb
z94a3bcf00467dcdb8695b35be3c886c1c7c415d59cb3f8628b0f867bc64b2064d0f57bde092f9d
zbb5c3967857f54b743b1177a50205ed56f91621bcba26b0a9873105acda8d1dbc0e43159a9bf6a
z34f327e670cd7adb3ec99a0c9aeba5d096148d33a9c6cf63ded3548dbc23a9b5bd5a97c82cd0bb
z551aa2d58160e61abd949042f16630a5e9366222c8041630f077399926cc213f07e5d3488a95df
zd3deff9ecb03a9485c3bb4bb73d101c211609c985f059554b34d2415d9b37d81b4dd3908e02c88
z98ec6c02c7f39d918b58e38805474dd91b79cbdedca79c3f74f597e2b0851eb5d35d6d8bc34a2b
z416151e40c46e5bb0c32e6ee6fd1bfb34853be164e702f3c18ab54113f5ffb84de4cc301ce92bc
z72183e495c6f4c632554b5517456fa1f8b70e4a4287f2a713d0935914aa4aae9db2f8ce5496ebd
zd648ed071cbe502203a44df8ca6b4ccdb9c464b7a8b4320c24456cbc0986538ef90efd912a4837
ze538b4bcffa299ccaf46e9b9851c88c5c4e6e4f53e5ed515f572338ae6cae114df39d91d914fda
zf010535ef2db7e027e35a3463a456a78c78ec646099b6806abdbecf729426191d9f8ddbe4b66a9
z64949255bba80b7d1e7b9b7bb846e3bb574222c978167aed25216327c3db8b07a89837aa064b09
zab432845e382c720ac7bd8ef72fa8cf1786d096102cff9769940afd2ef88ef46b9e87bd7f9022e
zbe07f5377c9739b6ddcd69af2c3d0af817b1999fd87947b058171ade97246b71f61b6eddb82edf
z96637203ade7d9f74e311961ba241d117bff5a6607252889f99947098d80ea368325539adfaa34
zfd07f86b0a51788cc51b7cdc8b62c805e823f651ec0c2e0e05b18ea79191ffd7860361e0018850
z6a559d1225a96eeb5f31aa673080e010f479dc90bbee8880b8c88d1691e9c513b6bf079313fc54
z6271d3c28c9d0a0f8c1529163b40eaed45cdd099937f64caa1825efeb031584e2111112c71675b
z3b2e5081455696a9906cdf38f82c5bc0b5866370ec83cd474b4f46f709339ecb7f7401acb12f2b
z13686184b9c1360c97a94ff5b4a1162f799779acbf8d78c5924def9a058892e9bf938131181f2f
z2f5139e2325343646bcdc2997679a15115cecb8bb3608f8e25bcbd74a4c1b0b0804dc8b4ecffdb
z4a61d627d04e2503c0f9e5d8e33918ce90342421cf33243b91e08a46714159bd84fdbe6f5b9d93
zccfc5f96c0899a8cb530ced8192341057666e6ddae43813dcbe77b5a73634c48ff32f9cc894a2d
z19e1e51d7e8b05fed4e0ef6454597bc592b81c2751ac382a00fc50c8af6573adae4b99a9d589fa
z40253987b0e5f39811f091d5dfc7ad3090061dd37df69f63f786a71ab8f5c5933c6bf0c587a7ec
z56e82a612314fb145568113cc5e15a45e0e1883e622b69f551e28214b10895938c742688834f27
z906001179691e5fa2f6b00b44accf573d082bfe8a8f0bba1a554c1b60a3687869ebf524f6b0ae1
z6e58599ea36670e9f90b5e4557e2714f0ffb8ee69b3812576ae9710f2c334301bbdb0502b84bdc
z6027eb59bcf9828398b3de477859b0930a44cce38e18521c027b76162ff7f942d5419a3f688dc2
zbaf99b219b9dd1d43039dab6e6fe91f530a1356519f73795e8e2397dfc6cbcb4cfb4b20eee9113
zd9923a7ebc9807e0f40a3303f41ee73e92f3de01ebabbf706d2573b66c025ec9fed85d3c6e409e
z1e3395d4e08029ff48c4bed75858b4b4494006bb6f75452587fb174cd3c73c83beeab08dcb787f
z54b755ffbf61d562dc3d28caeee254bc63ee8845f22ee55ec32f285e467fe6f8471b92a0429b7f
z966739985e2c61580e65313972d9643eb7bf05669991e4e69657e8c6d20b6dc62e093c97632cf9
z337b9f9771a0105e210a4b228c372e63c54ad0a93a7dd1601cb9676b667d5e6ef6360a726947da
z16b9442982a02eb08811b7c085a1a57be82efe49573bb96b5836a15c36bd9aa3cdf06d9f00d3f5
z94c283ccc8a056ede464d27ad043243ee346025476ad91f583c468cb1e8b9767a39d8b141030bb
z31aa95d9f586197faf5481773aec61f07c3ae68b0aeb6b0b5fbaf7bd1f032c199c9e78de11b7c5
z3bf225aa27ce882c4dcbee95a45d2586b9cbab1871b63869241030e9703cd823d207743eaf34af
z0bb260fcdfc621b7018b9462309ffce6813dea0bf169fb8e74a2cf0646e49133f865d17a3f3418
zecfd3ac1da5605855c863392ecb196c79636d3b40cd2c53e0f9e63f4249170642201500a3a8865
z042968460b45e7ce42f3ca894c14f6f008107681f83b4eb0d8e810f3e97428a3f1daa12605b039
z2e3fb73f885df24ca228d4afdcd8371850650f1953358094bbf457e976221c78c14c94dcb2942d
z125474d0598c11891ee87757c95ba67a3c148e054b997f7a710386f666cd1f1914f9a35ed2d850
z2161eb44f0244b5e33233cd712db43904f68e01de775ccf63cbe559f32776ada97640230d03ceb
z724b4132f80b420a38475061a0c16df59b6ec71782f820ac185d386ef7a3caef7e5e3618f4ec46
z93f6575611731c14bc2a7825ae54057f87b30c6573edaf32755c41510a22fd7e685a607c44a432
zf8b2621e4ce4e30c26f2b4d6616f08945d26ee845032410b0a5f46b30286da0c668f1e35430610
zcb6fc60c6eaca924eb9709f08e8ba9a92df88a9715808504c6695eb7679a4ff7d75a5e7b2f34ec
z92a535137d1ca6ce7063a9db04085916047873ae3c54ee6a8282ded2ac58b8d85269a5cab40291
z580985434222bc03e94bd228ca81946add5d86b4af58e4c150bb75929c09aae66e3a0ad7fee674
zc65fd408b1e35d544a23508011aa9dd6d84df031b5e370cd8f390d762b5880c7e09155d7b9ef5d
zc5cbb21703851ddf7bebf02b8641af961eadc89a7490dcbf09b6ac968b58a1b6e7aaa6d0373535
z50f28dd24a1e8d46a01c5cc4b5603b76067497c951f1f649af7605878df7b9fe549cd3faaf9076
z15bfd3665ee358b499ccb5a2f3eacc9e898f42ede56f2a1c25f747297e9a329ed17064cacfff05
zfa35d1808a53e0958019cd45301beefc1da54219deaa2f7632657d4428668192d5ac1d964f25d9
z520dc5617c479c7d509cb9d88e1b10ee6085bcfdd06b8db673b06ce53e95d78af4774a67e6188d
zee383f6b2eff478c3b544e4821b42534b0fc580524429b7d180b0d086840faa52a1c8f32b62f49
ze02784d8a545ae717eddef8987efe929a7a501d2fe1644c0ed93973e4a6a0918221290861f3ee6
za0a6b35048dcfca969c46f7892bec67b095c3659381780dff7d20e990ed5aeb8abdc2e3f9380e8
z7ae6d43c97fc1f556c5ba486fefd40d8e28e4e255cd2505b58c9d4079cd8eab4b6e582669e91d1
z72c732bd971b7439623cf462534c26e47313c483dba294c0da8b2b68f1bdc2a9f585551a9fc781
z80795c1a60ed047e2f50eb50d648bc3acd60585fb9987402bf989fb8c39fc00d6ea548e8d39207
z121ed92ad650030d5a631ff13bbe1a3d20db400bd32caa8e0430ea5157e590abb9b62278fff096
zbdf41a53e1651d21cf9a187465a9483524a6a218793609c5a3bf7867a70454f9e2271537ce2965
z00dfcac94126694bede95a20ea28e641b235fd27c64a02457b8a7e9ed5d7cb1395b43f250eb2db
z2efc3c3e99666a13e090c6b0173cd873354d804a1cc75ff1b5f76f49eef4710ebd3eb671be7f50
z300414610eca0a06c8af93e4f1e74d1a9deabb66dfe8a1ccd63594bdeaea800c6adae035934489
z01099d7b679c16b14ff0f42feda62a03338d4709c83b9238b60334881287d44d099375d2d67e4a
z3af5e351c180b61b2a81643894b877aa8390eac6b7c6da15752660a6cf9023f31f975a43f8d3f3
zb4ea97be9fef4af43ab0ea91ee3ac0bbc305adf59c823388bbb30b01bb971ee33583ca22a6d3da
z77b57f4e2aa30c40fe8c8e31cb50bc071b779ecbf21afa50e730ed80d2af0594b46f10d3311b69
z496a12ce64c5b9660083f1d83cd22497de552ef107d9793c8e9d70a93123d26cbf18aa60dbed40
ze8c980aa6052dab1a0ce0106ccdc1e4203db3c7cc6a2179956b414156f66d131069fe8c618fd99
z2a1fca5aeae8d15f3df105bc2b627500f9a697b0454005a561af4bf5feb276efad3c4e744c264f
z5d28612657ad66c372711040abe3e6f37441483073c30315b59de7f4f112cbf1dce12194a69a69
z3414960d57d9eee3af9fd13273f5b9ab45905a5c1684a204b514831288ab3b729048138d8eabf2
z13b956ab41cbd22b3fa92fdbc8e89f2129ce197588d1f4029961bf9216793d51119ac2bf72beb2
z39cb0c75d2c950ad13cc90dcf51cfc67fb930fae8423da0c38e14eb6c3297decbaa3e1d8f7ea74
z99bcb67ccc5d25f9cc422d2b57fcf20c2713f09218d15ec3d7b0ab5f9dffced41d91a317df9b46
z23770902b1109ee2baed646cd9cb1bba1b1165619afdb807964245642c86338ae5cf3631c12f9a
zb7176e0e4c0324e3fe4a9dd3383356b7a88ad4e894a148151fcaee88513a534574b1b754f6c365
z60689b4a46280ebbf526ccc96fd472debef258e2882c988308e4c5bdb4399fcf2b9fd34ef02dce
ze4418e6d4870615003612ee6fe050ca8787469d6fc985ee4650e5d9d111171590c8c0863244e0e
z854f32eb5bb08019401f5cc51377cc575935f90eb11334addaadba31293642f1936fad275adb7e
z4ce67dab589ca3cd68f024cde3d7ec0dae7ab21ad8351b379fe618218eccbbe7eab3fb3a42acac
zcfac93e01b15fa5d495f26b2478226b4d81940f3c7ee556efbb231d1a208a569815aeaa00f7666
z42d3d89102034f5e70928d5ad747cfcf2e02b765dd3c3fcd8ce998c5253ad369f64fe62870a6fb
z59d2d484fba7a4a1f0b3d5d240b1c2e964740aa8196b4c8f6491e646085aa6ccd1dfc7f36aca41
z162e1003d05dd08c81c5d1a704cd142d3f5401190be017263724f3243cf748491484e612353884
z5fdb88d3b45cb305e7aaa18b346073aec7ce90b988533f1f4a362f86f8adf2780d1b653547637c
zb75f4602a27af3b9da410f591eb726d1a0b46a570ecb7f2772620816e048f508ef815159e757d9
zd2d304191297707d65341afe033aebc221e8c430d5e6c39ab0e7d08a519326f8f5c8bfe114f19b
zaa41730d0da6379b6d0e3e80e2fe7b22fc68a6c30f358c2f56f9afb5cbed87f9536bcf6cb8725c
ze45bb7b78b5938fa69713c86ee7243d7b20d126c2b64997bb74e8798bc8751ce9027dac9c97d63
zb07dc6b912810c91663e6b1b33e5f720b961eb07f6046987df6766f56f1a35894398978e007b18
zaf05d8fee011569920d034aa044440bca4f91bc6aa690a31217f8c13357d0f91cdd727d4b43fc7
z3e39544f5d1b2ecf047b7e0060f7641be8240ca96399a4a5f35b4b2e82c6b97716692e8158429f
z27b348dbd9db6c95e6029359a699a30a643fc8c699d26cbc7f7924893d8481d1a72d2b45eeb2b5
z90b1fe632640ebe0404cd7e6e268fe940ad81f83dea3b053361319ec0cab74044c4d06899c92bb
z71e7d72db61ec2bff414eda5cb9462cbe52206898a541749fc00d86f9c79700db8af063b34e081
zc7607018c2fcba5b8c95d224623ef512a7d219887ecce47da3944ae43b3e73e98f735d314ccfe7
z8622e2d7a3f0804d4cbd36d3fd9fc9dcb8dbb185b7fafd8a61a7168610149dde70a2ef6a7f07bf
zaa824af3b96d441ea28b8bf035833b9cbd6df52401d1e05bbda03f96b09cfa2b245cee68b78b5e
zfe29f25afe5ae94a115ec04f0eb4f3bc359ddb508b179988e6e67e4353099c3475920b036200fe
zd9927d1caf43e4f25b9437f4d59de833b74b80e4c18b58c9f90f909998a050d78ed818a4c8c54b
zb1b3c15ba668d6a4f5cc43492495baf705963eeb5cccbe4d33fc308932e51ef24ba18e5cfbf348
z2736cd0cc7751cdd10cefb90ff11c644f45bb03ea43b1b63bf9be56ea52d04c489136fadab95c0
z1c69a71b5e1fe0369cf6e499d21c950e1d0e8ad58c800f26940508c78ee6d8dd75195ff739f09c
z2c802acc2a534ba6aae553036a6d211ca688ef84ee9970d6276466277a1ed7e9d3c43c68c10eb5
zff2bb870fdc633e60c30610e2bd5adfd4196971988820b3881950f929e53a892e7d3f5c327db4c
z9c2093e46447ddb4f6353d3523eac9d418dc430346e022c0f7b65b9de4d74e1ebd949c762f0d4e
z84786b1fb8d300076da119ba84026edb1c6df8ea2c589da3b949c19c643a495bd3560ef601a640
z958ce8bc5114f48163e71877f0b891c45dc17d6b6177e74f9fa13da52f8fe5fba535ad784f83d9
z904d46d2929498ca8d6c657bc2f83a883b5c34eb5da9191e57cae3f0d7574a180e3e4c855c9513
z4c550bbc93fe5baa28d01a90d23c7915ccd8813da9b86a30dde496a0e14e3fa5df34c8f44693b4
z836a5a0d2ab2a07a96321ba3a425e6db788f07cac3373e91d2edaedc38a9ef46d56f5a812edf44
z2e1b1729b317a9253b30200e182c6c654b9f85012f7e66dff37804819c06091fa3de722d6da2da
zf7674aa0bb01fc9bb3266a72b47dc88329c683bdf8202971571363818dad223c1aa6b30f0f5b5a
z9f5b6433eeb889f9e1b27afddce0f02b2c52a5191dd4c89db808793b03cf1a2a94bbb129595345
zb347ec6c1c192139d6e7c6933110d4493b94244e2f4107a9b4a796c9dffb106053f67a262d1e4b
z552aabe47e7bb3104a11684797de799a9cd4b3a197c23df7e1900a7ca287010ee25e630d0f75a6
z960d36815f79ef0c64f8cc8efee6c6bbdfdbc1f054f2654af271e021da12b74344666bb8809f79
zd0760bd8fcb640e83c17c6e2a8c896136c6b15e8465fe9b8f678274c02c974ab699ea31d68a93c
zdc1ec409d78083e6f72dcb9db7dd8fdddd795b4ae4b115d43449bd1848986b1ee1b960a98139be
z8546146190d712fc7b75ed4c5cc8640691e3d0944afd6166aa5ec96e79cac8a01048b5733119cb
z4a1f06e2810cd2eb0b28e3ffe82489dd7808a7839f28a7f3b7dd77f7c9017d18256321629ba967
zb90d19e104246af535d534602d4ccdfd0a1c49698585dea1f4b122992638de92f36dda8952b067
z76d42f4a75935cff40ac9fa38c4d18731ef4af5d7e1f7599391a6d24657342b9d28495f07f4bbb
ze1f23ff7c5d56c7bf6dd648e2d3949de7810a18ddda18e312950a4370dc3d27ce8f5a047fa9102
z81d64eab9e39c72e46e125ff50f32c09f97be2c6663203b1b54547fdc21c88d81d71eeba730e08
ze639d7f8adaa483a870a1af3aa9e3f23fa6b429849b92aedd27e74a9e526eb63374971fe6ce263
z54013af6548c1ebe6cd1406c406c03d27048853fdf09b232e96f1c26eea780287f5583b5eb5da0
zfbc1d5ddb81728626886bc6739b28909d575ce0ec9c55c5c88d8ef0a143fab086f1b42c25140c1
z654fdf84d06366d106f9d87b1e36780b442eaa0cc423b9d3946afc203883246968f01744458e96
zd0c20cb173ac7765d19d1ee8a10b367dec77bc1460efcff2bd7968c5b8c7581f353e2bb43ea9fb
z12bc72c6d03d2f8d9fd0505b5cc80754b789aa50f4ba9b06604ccc595f58b567da5eada41b31d6
z5b88c27e1303405ef5cda487a6e06478b4d5f445753c4f3133ac0c1794aea39455fdc9fb25609c
z087f1aa98b589debbf5b57e57f0a2968fb013dfbe7fcb912d384f7f904d2ad426b64dbded1c314
zfd51d58e90529f15bb523fc3e8384be9d03ba11e4b2a54791bdb5aa55e6fa086e343a704fa06a0
z4c06161cc00c7dc4c1227cff539fd759147b7ff83ac1df140ab0c7f4bec72d951da7e80fe4161e
z547f25b0b9acf3b738bf48f2f1a667f744cd052a8bedd2bc4ce118eb6c3a6b0250bdde8214049e
z6d78f3b3bee96f46ff6cf120e3f98b4afec74d49cad7891a504ea5f9967044966b753b92405fa0
z6fb69ce894dde6b31c4f0eb761bd8855e2bc94e369badb2e74fca6691d58b66a637fd695f2e6d9
z02c824768dec52f14a25ca24f6a7aad648187e4b6ff72886a6cf4418c1ecf17dbbba90d63b1498
z603e147bc97e811bfb7031ed64a3fa184bebee6cab6714e9548fcebaf40b010d36a1a692ca7269
zb7a60df71816f6fff508ff87af0c87156ab07db62977ec210120f7c107134c3f12174d3d57f447
zdd854eeb60f38b70db4ed93d14bf5ff77dc73718908fcf2644adb0ed075f2eed0dd0489ca525f6
z1403b1fcc28821cfffe59856c42c9a64433725df8f7683823f46fe5f81fce987e318290becb6f6
z9f1f0bbe2b9c7d126168d66e26d447d8d89735a8aa7027e149686474ab7c92a2f173e551ed1ad9
z8ea7f11ab8f121fe9598f98fc69ecfaf3c2dadb043dc2578e7f871d081fe3eb7ed34671cf23a91
z6988e04eecd19251f1201cf6da53fb7470eb3cf078a8ac56a8f988a57f056fab483b1a6bf04b71
z5653aeb43a679d0786c50d610e937ec35caa8c8f043d994c5a1bd1c1141a41082338d8ffdd2dea
zc322470188c23b44421b28668b48c2aec7acfd4adff414c28b7fe0dddb536bb48abef9acb816e4
z85d077114c27ba03e16bf13597e4c07076c5c15e4a03c1e53cf182b00e5d39abbf907a709a750a
z84b78f1aacf916a1eb867575f98cad5f86d9a32ebbdf4c1fdf864b2d14ad9ba8952d08940ee001
z3c711c7d7b5e5a30f181875136ea6f8f8ef8de53d29ea042286489af860c53deccbb98b6058824
zc43254a571a6cc7f8caf21ca8648b9df756a71b699d1b95102a4e2d378c605189b8cf62ee40aa2
zf00f7f67ff0fdd712a9c02b1325504fdd5e8caa4a6f3a8b5cca14fe25828e8584fc2de67b89bf3
zb12edb1621e8153f09af3e55e63af96bf94a95dd4e422966e28c3c0cda565b005dd4fa03abcd6b
z2076599b611bf7065c3e2c73c8eb8a804daadc094b5b148c2c24bf1487126307e2dc22f28b7f72
z965e02b36a092e5366b18c516b5aacd6d0e72bc3ecc54faaeb0bda881f3ce2412662f01c040670
z911f40f2f0190a827e9ea846de4654f3ac4a8ccb925fa3d18de7139cf80e18332aa2fb6669f791
zf15862a856c7f650c729477e1481cfbb2eecc0304c6ac4ed18ae28536eb082b519060f8ada06b4
z1863c586aeaf4beae6c905956146ecf676575ee377d7c2f97d7267f8c0b04106444c79df797ef8
za65bd3c1eb3ce735c244a5ceb352abf1aad92011704e3faf117d161f78c9d1e0c2d42bea841e5f
z63342afcd18805ec8bd373554883d77252b67d87271fb4635f1663b70b73a3f9c99d1ae01807fe
zbb005a96fb15e11e516f9a7ddccf5dd86f94baf12ef7faa054e5c54bbc9fc1106b094bc346eea4
zc5528812aacc9b456010825b2ed0ff77fe0a11905fc82b38cfa323ccc95e6ef3ca2793d82c73f1
z5a932a1fe6ebc001f18b9deeb62744b0470a46cd684baf960fa3ac4b13628707deebb521f1f250
z1bc0dc39fcab89867ce1c4adfd860a95c0340ff859442837b26002e16fc92d240eb05c076c0af1
z574faebc8c0ad782f886018b3215377a123307816868237499352c0d21b206816e01ba20aec9d3
z634301e717165ac9c0115fb487d0c4c7af05adfb86b2448d1f27bcc386f48e1f995b6e7f5e3604
z78c2d877369812e7d58c7608c80bb35cf638bd77607200c44ed0f02c378cc46350965c09213ad6
z0606bd878939544fd1fc4ece99cd50470de7a8faea7bfff94365da40a5b7e0a7fe8e29cc4b6227
za93f9c5a5211c8a6c6c9d5a448eff3adfbf20394f884748885dbec693c766447975cfade0426d5
z6c20b1efbf144e4fff454b2cacf17c605128d7e855d3d711dc276fdba67b4b376984749792cfa8
z5cbc607ad02839363bc2aabb145958b24b88e6ec512696146b0676ba7208079c0f9badbda48e98
z52fae944f7d34bdec3c71e75a4fde0e83a7ee594085a1ec8627a84edaef5ff1597439eadc8f4f5
z0315ab672950dfb28c295ceef8d58bf82e10031864b564dbfc351ac14a59348f4548095a168502
z02821361199b83b5d9bbe36e4fda0d5a9db1ae59c8444266626952bff6ed725eeb167911ebf0f9
ze60eb196b42385ee3206e022dd10a7e2027cba2d3eb73614a0660147106781cd787d294011c4aa
zacdccec3e7d92e2d8743deadbb394a62ceb204d930bd3a4d35444499bf9ad14985fec9bdd2472a
z21aff17f964700ddfe1d0e520886540f8aeea7b06359fd04701e3208193710527fd337be4c7b02
z7a38d4bd3177de95b3bf6834188590c02dc79470de4f18324bdff61d581be05a78847f074a1d01
zc469a9a583f6e1b7309930b976ecde0d7a2919444f8f95221dbc4449f4f76e64a246b8c4566ec6
z7fc0171280ab62ab4a5776765b22dfac85be153cc2b86833629f71c7b91fc9b661e5da757e4d57
z01a3853a9dee1782e42c920fb775bc941dc51b26ac8f76b1f89f136d7839865e22ae5d494d7957
z157efeeea6179414e3b270f3ada6edbaa3121316935cec37dbe91b16b05406833e8b4bfd22adba
z1a30461fc1aa783c65daaf299df9451b07ea80b76b38ee746f8a8031e4debde5cee042ff55e706
ze3ea3b3e49aba29efa58f9e85628cc6540842e3f26eee9c6794e7c32e911c81aded76f8586c74b
z726cc56ed385ea1685a408bae75388b71f43e8b0c1010de4944afd26b8ad4691c2003a4a5fe0f8
za782a0f6507f9f21ee44f5706591ef48d8709050aa5285c8c83d3735be1137ae2659d80821cf60
z900fc8bd30e772ba75aa2e9bfbd57313ec9a869f7ccda49603133f3ec2c2935e3dbc55a49b398e
z0ec70af3c6cdffdd44a53ebb01fc96f9d017873272d15c3e5fa27fe6ab1c6aab8b1b90d2047230
z274c1c11edccaaebd2c31aa54b7b6f1c8389d96ae4e9736238c8a82716c536ed988033652d53ab
z8e979fff7b719fdfa7776eac81086a1a423745aa7cc165685cc627cc3b8903267ed62c3865d026
z621fcc8d411536b11595fac09688acb048a5df6638f49c3a3cf852b349a5daa37d01ebee54a4f5
z96824eeebe86427bd49471ef241c77e34f918847f5773c3e4dac2abe037485145f75cb3f8c7775
z21651d50b3bfe4ddd8b1584bd20196c3b20fdff094b9b5fdda0af33c2cc662cdca02d2cc6069df
z480d11921bb09b0f8b4b590b36ad1430511f32c291fd9bbb5f5635ab48fe061e34842dc14b6648
z3c1ab4b55e55181d68b60b1c54d5473e7ffb44e984a7ed0ff21bf3f3f099532d004d5bb8ff03be
z8badb99a76a27af01495ae7affee63e40abdc356bd4b8f4af01b7d566005c165a0b68eec202746
z0e82de39090fde593a50aaafdc109319589cff83292601ecbfdb71d69aae97508deb1f1840ce22
z04d9a5bf02376d84d0c7d00e84b2318112071df98caf750fbd41ee801cd5af6266db55e92837dc
z678096b2af351bb6bf4da8911a8287d1a744ea29ca8d081b806b1a247702c5355e530b70cace1e
z9ba1fd1a742a7a97be9289775fd19dd2699e2a759d046c613e8bf7f26451628a79e51a21a66168
z64656837a38b582f5998055d347e83d9efa9639fc9f7247e48cc7f6d3bedfa805667cc65803d6b
z928fa27b1a5bf007918cc24546bcd725612bec433c14359ebbbbb98980cd897c4c348596f5d0dd
z984562cbcc991d111c8cd10d8730f68ab1742ddcf435a03f73535b7e72c476c1a37f1495258992
zc22b04e4bb914fbec0190fcc623e6bd32c0b5c3d07197ac766fd00aecac6205600ec06f3f77c72
zed6c3e51aff4718a87a512d3d3cd9353c829777341344dea72e4179d86673b69ef20788119067e
z1542e73c05a818192df9f7fe63eadd7906c1fe77f8971e84559b6929bb78b8ddc7773810e4d2cf
zbafb90813ca3c4fe6b15e32408df0fecf57ef680e1b2dd66f19a5e1c2b0734fc63a986bdd65399
zc0ae7058813225eb347f09bb287e67b9581a7669f7f012ad4f1b2b518f2d5a856d29453b80b13f
zca6adcd2a93102a559bded31de3c1b94a60c9f7ec8b63329f8e2d0a6ac8c561c220e4aba083cfd
z865307047610330b246b021284a77969606ae3ecf4e4dbac8fefbe896ed9cf9d8b7d401095695a
z7dad8bba02b08152fdeb8c794ad06fa09e5bc2bfc074a8e72df3eae254f7f76010de7d6c456448
zeb50a9c91fc955ca502a7c7370430ba634301321d7d62215428a342e292e01eb30533144331f01
z3db6f0d5b24e946916ca24b19681c2d96a34308cb1fa9f3a7db237794bf80f48133af8f1146b46
z13e2c2de2a2b4356b2b7da2bbdf3d9daffc2b02532cb0c3ccee5af21ee935966e770f7cb537847
z457fe2681f67c8305f87c44a7a05ec49d281c96892b68dd5166428206f54c674e7f5bf453247eb
z4c5ac7980d1438497bf97639b64af2d251774048c8647e9cf9fa37f2d1d5c4a50b2ec9a5f02c5b
z77918b448e2f8e2c2a6ebc1fbe4ff0dde1c390e36d9354f1303f642c2da75d13bdbefadb8db5b9
z454d50e19dd2569df81b1080b57ee69a29d5bfbc0c591bde309765b0b96821e2da973e9bd753ac
z4181bfaa45a69b92ffea3815508e902612d58b296eb62407ec00fdd0ba1113d04a4268c723a56f
z77a66ba9589583d5d3c926557d41f447a9e300aab638f82fcbbb3e6df5e477932322d7a3db1236
zd1b8a33242d2f5acb47c867b6249889d129e80bb6d9be9c64a5bb7eddee432b57a60e94b566e1b
zb4fa1d0978e6a201b144bbb3f0c2839b7e3779f99d1f52bff886539ddd24ba93dca0d71607e2b8
z3dabbcebca5bca39d14ceedfffd1e4b253a30ce91cd0d79d2d33b0ea18f654e207fe2967f74bb3
z6ef987f9c7755fe4d30710cd7200a46e610bfe7aa05ce8e0dae82193da1e1f9b19f29e1064c355
z4ef84ad4b655181ab66c7f639a11ea8379aa49b4f36d182d4e0953976079209a0eb167f441e94b
z6538717e783b57a4d66c85c36d45e682c1d3b12d504082611fba2d61d8be369e9c0fa34693f066
z3801924ccf56905fedc94e1c712cba3b0f63fff5094cf0bf5cf0157a36b2fa971715b84b13a9b9
zc19f5fbdd41fe1beb26d8fc646e18a62f1719c7ed794d22ed2739f49babca87fb37e4efbdab913
zf66a1d4dd4f4853bf76ae15180cf7f66277b5ecf3489f0e9ee181b5c8e3125a43a80243a3b0297
z3324d037c96b3011c65b4417522c8d233220794a7e54a51fe96a73fadac9541f92d65f492e307e
z77843712e50c32537dc62d4351b79a09df0c0cfd8881c60b3a52edd37c56fa602b9c1ca2d6ff1b
z2a13ed003d7a9dc0563712da92e735d5306900f65215937af3b288c040b0851f5250e4ec5b61d1
zf33bc91930c363259835a2536383c710b26cd59a9efdb7c1db276533bcd63106311cbf0edd3e0d
z5e5cc43b61c73a312bf50202db63c1fdef21984d9c413ed629958cf26ba897a2d0fd754c18e84d
z2a21106dcb6553ccc48d6150a4888951bc8aa3f21e8f81761ad60f967573fbeadcab416201b45e
z9af883d8feba44215a077c6723d0c6d61c08b182a59ec98c537ba6062794cbd8d0d0bc7661287e
z3f831c83deb71540b48593fa646b70c222332e2d545b174b2f298691d14a3e58f6e2d26e4fc7da
zb7038b1c7eb2c4ade861527a93ac6fee45a73ee39fe66b4e793578096c53c0f40c34ac2169c287
za29afce17495346ea23ddca4c5d007ee3dbf7e2a3df88795c745ebeee2699ea9bc21e7771cc03e
z6c94aeb4ac2c9f76275aadeb0435a897cfcb3989c46ef145dbb5e10f8f3e00b290a2895a0213ef
zfa813c38a6055d20cb96a0950a85febe771025e5e304d01f2ec634e3b8b16725ceae00abc1819e
z4be759796d175fc97e24abb87e93de146cdbeedca5c0a840242dd283f8fe44147ccee63024d862
z39d8136138c9e5468656614f4dd81de1306a9e673865c49a794fc3ece73791898f36d251277099
zf437c3eb343cfc9442f48a9c64b29988ef3b34bef07be67e1f842f796b607f4d5837abe78c13a8
z5a094785a85b5bb971817d957a3ed5e25a628a2cea843f26d882717262ead9214e2881eef71d54
z80af18c56b0e60a00a66200f1b829c4382777cf8d7fe222f278bce045b430d829ebe29966ea947
z7c4fae91bbd459b5e54363dd8e30aa7c063dabf1416d0abbb0736421619f2f4c19320af40f3601
z7551899e3ce0dbd2f66a63bd35400baf8a2ba5874a4363b738f37876338c02a205e6d55b8e2fe9
zb079ff1cb7edeb15bc4f075d66546d2527eabbb28dfbf57cc198b5817f8540fe79616a6e6cb3cf
z37381d4926590b8ce2a78a7f30a9b822158f91c5218c9ff57675c1ba9d1344dbd60edd0f74025b
z0ba96a80fc1ea43f79729b883aef8e2c9876d222c7ed7e4833304a50a854ef79225b2536c98dab
zbb43ea295acfbf3999cef8a004c5904479f4536b688b30f5be86078b19d42234c650493f87b435
zfb0a36ee8cd2c3c6167f12d703624918d6b08a9db765b8cc215a07b874033ea5cedf919a2f650d
z2c9d972f208f1b8a2870746876495b71e00f20113545eb8acf0f314208a92494d46dc76db3266b
zcffb68ec8ab8ca3139e823d347ae96b2af59235d0cb1c00c69fec10b142e067df2235345b1e96d
z9619287d4308c9a97f6477c6c6f091a415ff287ac9e799be439d3e80bc3b3e86bbfb362dc931df
z1e4dab478e62df612c35d98bd4336761dc64f6e0f052445f80e09cd58aa9b1c40f0f3a2f870a5a
z8525fb7e034b93099edb62dfc232b9634042390a2f3111f09707566f189b3ec9c7c5d72e8b3d66
zb338c0a0179d1eda06962538cb4f30dbe98ee37fcd971ec80be7e796ce43c98c4c8dd67481efed
zb6dc5cb8c073b14d94e07c89bf14a444cd1dc40f31ca2c47d46abc75767558ea5e320a10668649
z46d1cdf5b6d7314579d3398e7cecc8f9b1a314698b0138f99161e6215a4bde3995cf3142e51f53
z2d3b29b436f42951590a5a2c3622562a0aff243c8115ff962fcd79ae45dd2d78e170264c30005e
z0ea4bf2473e28837d74ab8993895a17c77205638da10d1ccd53e6bf3e71cab541aa4a7fb70685e
z3225f0b7b95e1b91756ada8c84fba8d6abffc06d86003942e54c03570176f35017e88226670846
zf67ad750b43b4fe95477ea8b49afe5ce1d78626af03176e9be413e6075ac30641080ae66dc3cce
ze01909ad3a5fc2c716cfe8279bc4cc03fd61d7f4ad282018e2c68c8814805dff4907f30fd5ef85
zf0c85127cb197268503cf48c2765d0ecf050a4247ee6fd7ed4c30fedbf6a97e796b89050ce8c39
zfd3e9087efa90f921899cf6d5be01142ede4f7536fb843218d54bb2fed42ca25a67155add8bd01
zeeaaf8dc86c0c453f560f772c97ad99b4eee872d33876497d5cf6c3a75f9988a91a3d84e061aab
z5f5eab7591da8bca1a83f7dc6d7593c1353ea95445a6e0b178efd6d49461d9aef94d2fce368c60
z14dda947f22a9d1c55f6c832f1fa5b69ea20a57257c8efaa71fa34e82ab74d69c15a28cf4a91ee
z5c110dbad1fe3be9190364ce8ef3935c6fc582f38a25f93a92073d91f1cb3a366545f2a1ded0fc
z6a095c25554e36bd31c4587b9ae81f97c5fb387ced83e91d4d3d8dcef0607cebc5bf0fea95c5bb
zfe52399e8bf71480362204914c8780c7d73d9b738ce5e4ae299763fd38f9a905974a1f400ad8e7
zb67f77cd5aa839a729459b8fb0bf2b104f5059aeb851ae4ae4e86869bcf97a83182b5345c7e9e2
z55dfd0224125fff3ecaf486c4b0bdda3843a05711347852747cc8a5f20a285f59cf3cc8bc69398
zfb5c9cfecb1085c24d5df68cf8d1da7c513944bcbef93a5a13e0d69c5969329888c7f0032cdc67
z9c97299aaf9390841304d759d77d1ba5359a5b9b380b02254c7bb125be3eed56b72c4cf9265a93
z674f8f7aec3f1339836d9a9057464a267be2e75752575f55ee405abcabe130dc1b7dd33a3ae5a4
za898af8dd64ad534b2f99f40edbb512b00425e16d870f00b4463c117f15671f0af49979b032811
z8aef10074d3f192eb9a9899db78e14a69cf65718c86abbfd317e4579108f2382b4ebca5f267f5a
z5e231fb8e9715791d795c801ae7515a9c5030006c02e8470b8c3d5bd35ce851f1b5393b541f610
zf9922c9e44a86df16bf4f07b3611d5ed7fd9acf1046919776333f500bfb312fa90027c855fe93b
zc09310d82a32c591fad1827ac896654d1cb549a2dad482bb218ff466d85d289df3453992f1f46e
z2447c68c7972a50d4daaa47bb510866bd2b7ec486875c96a92e1b0fb958328058437ea5c3bf799
ze07492f1242dcedd91a7444b9f61bffb182e81293efc89f329c1582223c0a118e88668c5221f53
z4918cda16423d34f555468395e1c3e54a7ef9d3f48ce474747b60da530386b6510cba5f1711a73
zbdac8ccf5d9d7205136924b90ba6d439b5fee2c3b9589b2ae40fbf9a5395e759f4685bb4d2df54
z03f4afbf8f6150dec3bf4d48d6a8a29d321d59b0052c988971574fb095b9ac36fe32f5d5474b7c
z39cbb0e823a9bc9e8e561924d7ec1d01d55cd9079bad3aaf6b6b2043c6f6a3993c2f3896871016
zf5455beac16f2d26f3690abb333105a36e9d0e8ba11b1b886df09866d4957267f0a25cec357711
zadc99d8ff7be3cb1564d12872bb35bf49e8f800a778d06b91c07e4b60185af7a28785d94a659eb
z382e896be752a5be52986bcfa63079819c2c8051f09d2a5829987772f3c0ae33e67b49ac3a7898
zbda865555d08065c04371c04cd4d017cf02d3b419bfcdaff8466155bf250626668957acc99714c
z2f6498c24e21e1c38a46f65c4a24706b2f41a98e96bcf7f4f2b69a5861dba5ec814eca396b08f3
zdc3da4535d17e50e778beb1404a4b3ae033a50740d8e982035ef2b8ab67aa4895d70eddbff9593
z13fa73fd14b6e8e21a80a6eca11dea82a607897e02a5b9ad508829624ff760e95f496018fcdc74
zf5721576331740f8453c6805ec9c14d1b1e7204ef64524a3247642546e505c40033cc22510613c
z02e6c4da2857313574168e79facea561e072def1c4ff0ce0867151a06468b4ae4423b7700a7c57
z7422d43665c796bd27c9e57e485eb4197e9464cbe3a8202856fae93b943f85931795f4c5a85342
z695618fe7d704ba3892f324aaa5ced6eabab710f833376c63dc64663badae704fe37f22958467e
z97e477b583a430089a64961d8a0f55c5b6282f46aeea39b36db2f2361557dc9e4bc749d7876339
z94f534cee3098583ca0eb32b33ff21426f03ac00458dc097446317d0b7fe8a3b1d6bce9440ac1e
z47286baa471c7546068fc76b9f3158f2d963c3442f234c3e205a16e840db15a88d9d7acfdffd91
z61b7cd4fc828e887c1994fe66198d0f118da7bb387d2c8f63078032eea3e18fb333df66f703e78
z18ea8d68e4cd12986f5bff25e4c73368a57e9e84f31e3c12eb341f730ed320c4408dc8f760a60c
z85328366ea18f380b28c83b584a0425c95e296e242fced9c4310a3d9f871d0959f9ed5ceae862a
zed3c2aa76697ef4c5a6180d7f82747bf76a39ecebef9d2f789016994e3cbc0dd35af34a7681b3b
z404405003fd695d99b7dc70a7a03c247811dcf5d565527f426754ef676d9de040bdee55718e916
zeed2f77be3319a83b0b380ffab6374f2716dfad3cce7f4936f60ee800d11860a95fcfaea62dab1
z899b5e28372fac2211e9fc7247d113bfe4d4a2c12a78420cf0ff2c06a86864519a5e801266576a
z764886eb32248728ff07be7ed010e62780f5a75a6f54ea95902d3fde43f997dc92068e85e47b23
z627930a943ddc25439d42802b24ae1297e60edb00419aeeb959537a3f476f0543ffe3d44f704b8
ze493eb9823fe1c3913b5e12bc2035b76986da6cd52597b1ad56801d2d23ec7f4210b16c9f53c27
z66ae371dcbf2141e6c9f51598814a9c4c05e525c61eb6f60f216b36dff750f3f573b116368332b
z66641cb3498070e3d41639bfd8ea2d7908b8e07dd5a60ba4a096423102208dfb427d385d5dd8fc
zc5c75adb189a387b27edf1fc98a22290f6b2ef3c34484b2f351a544ec76ebbb16f5f6b1c563e06
za4643b7cc31d4e61758986b18c67750780c8c730b1665c018ad656549ab79250c38da1667b93e8
z870345791b583d6f1030bb0830c5b7681240f7239b1ab854f9a46021c5c4f7221419798b6e8472
z6935be200773e6ee55875919cd64b9d54138b191b37bfc061941925892e77c8c2d067cf2af9c02
za9302da49e522ce6c579b668e701fc14701c7a71bbc7cfb862e4fe93e3f0e3f7d529479c0e743e
z1f8dc56de57ce6b704fc201eed5e1f0f982367dc8802653e34d64d0687e64313fedd1a0f476680
zc13cbacf5ee1a8d15055020ee5c46ee211093b06075f16e4f18444d5b61841289f5f09d78c70d4
ze3d4752ea7eb555e4ac0a0179921cc3853c2a7a7068b84434894e34e70af7784477b907f6d0aee
z2e73c17e0d7db75dcbbf04a9465e93b678f721560bed4e414654f268eaf2316950107e4d6e1edf
z13a694b4b18230f860ea7bcf3650755d6025b32d72fd8d59a4a2bbaed5d4810dff8799d5703017
z27a59d52ef1017a40f2d05aa5769121f96d24c310de2d083101a65ca4aa3da814d081abd166b14
z06be1021cd5e6e0fe535b477f39469ab0a4cea878fb623c9c71bf7eabcfaef1f5fffaf79427008
zfd458d564937aa2adc7702bc73019e11a2eba0d996f0e157aef2334106d51581ea23857e70feb9
z64139cce770efc7c695d3643b4e47077b7aaac3238ed75b7c1716edc39d8eb7d169c1a192e4463
zb0706e3e5d0ee6ad27f5ecf73c1f1f88267488518b457f83cac394e9615c6677a8f1dca0ca7612
z0b8405a81407b0f5ca3a44ebceff5af33f63761b68ce968e0c7dce6b51a865585f414c1bd2a605
z04785cdfe5adddec65f76d895886b3d9f2715f22f91f56b1d1833529db954f8dc239646a11827e
zd57c39caedcfbea0c84d0fae6a8311923ce1426642a9724da57db315c226be2f7daa2388cadc43
zdb959e96258c882109ff8dac0aca05fc07f59872b9a67185f3e7484a85ab26a32131a9f68664b1
zedc1568c8ff49a0aa6bbb3542a5d66ef68976c88eef9eac6a3786ed20d36b63fba0c45e3cca2ee
zc6c53fab59166040d2c019eaf4af2ee08080d1b93b087c053506fc5b5f3b3e85762177691ec12d
ze77eb120374bf1bf7e40e23d475df363785bf5b65d2e414d7affc328fdd388198693cb873b06a3
z507fc48beaa9780c6464f4de9f84c159f2059560e6e4575dac6e85837f1de9cfec1f851ab64849
z3ed1c67400d5283b8798fdae8b89dd4f0cc3bf869f0a85bcd812016775505df22501d2047d3365
z2258cda6d7cf5f4c13a1f48cbe7f5bd9f29aae00bad3458707b29881ec2fd8cb3b2608e2708a3b
z78d1c049951ba54229213305faa35427abba5ea0637c5b7a6614ce19ddc06bfbf81c4fa06888bd
z838912b0069807e9f01ad1330290df23509850cc21f638a9d7acb5606752bedd0a727660238ddd
zbcaa2401558b3d6e0f5a17df7d1bfc7fec95dde1b9dc693e37375d9e3adadd1222c3ec0ce0d83a
za13c20dc5373933f9f70789aa75eefbf64a86c250d25076ba3f30c83cc072190e3f3230e16fa95
z086eaf6fd6e37dacee558a26d0c47a57cddb970f6856306bbaa7529ca6104a8aa0740000d15594
z63f513b352427157dcd665c34438469798d3c825f4fc19fa3962df6c424866f1dd1d3db42b1a0f
zcf1dd17f9c290d10fa995dd0d363212a5d7a5b493326907982bb3021b0ab7adff8d6e1a79adc7f
zd71fd3986ae7d2ad1dc2903de0f2c82267c37ccb307d9bbc16bd2f1b555cf10e518fb7ee0ba793
z87a8e599c8640169747d26bcd6c553707d3716105ca840d4c07d546abb05ddcae322f8b8ed939d
z2ae6b9f47a519dc83729e488819e92fbf27d7dc11ded768b9bb80b62e5253a68c472417a0ecf7c
z0a9648b7da7dd31539147d606b7a5f2eb14c9f0d8d8f3203d4f90d92a1a2b7e91452e8443565fb
zacacb522b81553d820ca944599496a4a43cd4d53647841dad9620f71bf9fba6fa85f2e319e2104
z060b1f321d76ac563be08309114531e1d01e231ff2e91819b295cfcc237edb42f2cac9904127a2
z749dee5bf2e60db80900d84ec2fd4a1c967d13feb4246ec7f7626a0b215fec5c1c05072ea67640
z7d95cf8cfc1ba2c4024df7031a57667ee22b63fa833fabc4f15d39d7698f332f286c4325531f3f
zdbd4a5c0f85b6190edcc2e6b9e7f2719ee0c8b9ffd21ff0e5ee4c4c0b3366538f27906a184ec87
z14c1d44a6934183886253d306a4bbeaf04fd9107da44cbea23aed77f8cf2d038cfa6214a3c2223
zdd83628a411e87898117bf2ee0c7616398c6f8ca52e28c939295ded554dd3da3f47c6bba70b7e7
ze54a425218b2838f2885ff1ad94c0841dd9cc149610415317f4ed8b7d12c8b19cf7594a840ce5c
z12c3870de9f98e7685cb8c98f958614113a8147b72c618f82e5f92e7883271bfa35f1b77dca383
z3d8c945a18c61530123413de30cb5acd5b1b9d6b29271807eee7844391b0e93568a7ed6c9d795d
z6ec0697cdf10111972874fd683d90431c154417e351a493dbd6b2acec48e836a70fa4ee926bcfa
zb2f1204e18d1c5147cf289b1e980b71bde2e9fbf886ccd08f82e245116e00f8df729d20ea16780
z8fb43a77f2dade19e9d93eda1d52cf365741a878793b3b43d3d7ca4d55b0d23d7fce5ab09d5411
za8567225253507542af7c23d3de6df56553371729c070b7584f4be49b676a4d857d3b85b9312fd
zc8889e21d411bc312c75c0bac6973c3dc6a051345b22bd19196e896913823e1f1607f3e51f80c8
z00206959d43f89da33f1fafea69895f4b60453125819257b12d74feedd0c09d27fbad6b2999ac2
z6f159471faab23d194ccabda68165c6844c98efedeec16ef814e3402221d2f762a8bcab924f42f
zfe0911bee5c079ff599fb3913ebecacca6bf273f2f1f5226a4608e35b00d540f39795edab15cd9
z84194490873f756647b721e0396e94fefc751d76877c956ff27e3013ed4b1d1708337facfda36f
z31467a928357bbb96bf909ede24b4bc3147b46f9868117a19f72b8e2d974ae849c1052a7ef055b
zb5789bae2305c7a278dae82ea7de1c47089a3a097a17c10fc048190739d15fb047369b8b36ec5f
z64e481d5b368d231943403cfb21d05c5be6c7a9ec59cb8c5bc0b2c0fa849f282aa10ff527a7089
z9be24f23ff0abd9140bdfd2b9d3063e5c6b346de7a25ccf931f91133f9bd713c046d8db43dcfe1
z6e48d53d56cd532fdc59df44b2591ab3dbe68a540052ef1da60532258a952f7ec09a29fab453ed
ze471f471adc62350a4044e46358dce97493e1f2eea80712ff09079f37e66471360a29891e21816
zef4d2231f460f6eb43d37a04ae469f245917f8203153f0b10e15ee4b729475d613ffce2e454d74
zb338ed819c8887d2c8cfd7ebb94d8d5786f85679b3b97297c471e2f287dd11a5b9fe47af02cb69
z014b8cc576289ec8c075242e545b944f4a95eb84f7d63dab624dab8ab5add949dd11830a48d5a6
zb621aec78c1c231050927fc4298fa45f09daf27065ea47c3f3b399619b59c718617138457dd32c
zff936f548031133ccde1fbb2666e4c313bd77de43839da0b37c8c604c2a600fec385f3d8f519e8
z2263e87e936a959c7699eeed6adc3910e268f54dc385651b9265111b60acd074d67aa4d8ef8352
z189e05e8319c421e348066ac780633cc287270553f2ad934391edfa6ebb470857b95513c511afd
zbb44de223310ef01141744fa830171d41574d07073a563cebbb830cf06c8617ed28464d620c9da
z36220ed3ba0dcc6fb3143d114a4a9f09478d67889c6cf625eddd44018b8a08717e9db1c8b51c9c
zbc86136083edd48ee947659c8ba9035d2553c1cc2d2f521654674e4324378ff33bf81b417bf1c7
zd81961a0869f5cb22ff13ad92e8b139af2d3cbfdd729e9772b9a941ffc8a9313be9a5338652c7a
zcb64e334d4629d214d509e5f292945ea498358630042a16aacc0255cd09dbd704bcb5c6ce88711
z43c87e6a02d2b35f59cf3d36121af656960965b2aa1037a645815c6ed509f4776efa544e24ea3a
zf169027bf1d2b6d44a39810b0935b503ef8aece0bf6b880d06c5650f550e4f3047fd99f15ac74b
zc66dc69846cc88084a7bc33503b14b4518ca7743e4fe6eb84ff0b8f3880ae1b3297dcb18e2b167
z20b3fe27061e3afd02c33d1bc37bd19f281cebbba851822edad542b27c568e41d390e9b96db097
zf63259b4dddc90095f4393af51b3ca8f94dba192014eee9cf733f6c29995dd21e47077da6d9ce1
zcbccf2f65238f7848b8eb4741a56820b8bca38262cdebb8df260a4ca91baa9c569199db469b615
z156a07ec5c95309c25e16a91af39a8559d1ca24e489ff8d16d07cfa63f6ce07e48f38a6acdbe96
z55f72e69e2c82066b96ce66b6ff164acc88c618e3fb92dc4a7441dd3822f6635993bda1246e08b
z672640fcd3e7079b894ce8fa67440500a8a26d0f4f7219bed2a4e9181154f28eaf201b01bcc627
z4bc91c7d4e2c9ef361daf9efb3d24ff8883002b8fde31fe7af474bbde743842d23a78ee7f22d83
zc6a9c1a0c9e4e5d54a710e76376f3a3370b5882700def3015e1d51978e4f15ddc3f75d1c644ed3
z0b357a73d47b9e053d3c1f382396d2f9e3fee99d29bdbaf2c7c16a89ba6a895789676e846eda29
zf62e07aaa91673287d955b2f0af0989f67381c8c4b423d2b722e7ec684ff9ae11841620290c000
zbc52541323e2823fe998b79c3096071349c19ce4c67e2d01cf585ec5710d8b7fd3ab1d5ea998a6
zd044e493b4c025856455c8568c85c0068178fb07d41ef1bf8084fe75919a4c1c0da6a1b13813e2
za8d23413e6c057743a11856ade224c56b9d196cb2f5850c4e0b362f6bc802d5f31c784ed56c635
z1f85ecac8ce3e3c511e27bd54c99279d306f375aed52eedd1a2bad20ef1528504b54a1c0a32d24
z0e61cc4c001e4517e376695d90f36d7041bbcf08b5cbbb09732970764e84f88cf428ef142976d4
z5c8a3ec55a09d258e8385b824bb0609ec9ee72796d22fa4cbe4a628244929503cd0839ce193a55
ze937de153e3fbbc4bb24b17bcb1443ecc1fc9e3217d5d17ff66b04822c5180345236ed1fced874
z86b49c97191ae5be4deb7148158258521e51431e7955e739fc869c6189f4f6f87f64644a162f62
zec026ac0d328d67539de14f858ecc4a9370883a9777f67de2d7665f0baa2060ee81055014c4cbf
z48a79cd6f45f7c565a839ad49b2733caaec2a2963251d229f93a449e6d01552466c707d3a45901
ze3e38297e02c23623c3e81b97f162ff7888ebc6f74b4b384ac2dca9566516b9d08b8254f0c9fdc
z3be7d02edfec352c33369755743fe85a449c40f831f153b7c4cd53db5be104336eb256bf6142c7
za3b1ffa2c5f3bc5c221e329e86298626f54f195052f16b3d2d57cb4f5b409df3a02292023244b9
z18ee0a894925ff23171db51d89e7a448ea132ca8c479aff593180b7de3bffbcbadb19bdd5410ea
za9ba817b12215f70b51b2c4085dc2ffd47be2057df37f6524d90fbc97a6aabc79f46e8e0e5bb43
ze4661ced092ab3c1b893aba2bfb6a5370b355a18b596b41498d3411e2755f06e88d0a713bda42c
zf2e31ef069998a1e020f280f5b941312dba4f26285f86a3a796104f3e10b649301d44728581223
z4dc03010bd05a3de1c4ac2d1557745634e34f331b55651a97e76511273bed563ab89b89c223ee8
zd620f7ab636d6f0fcb0c13def9c89182b961efb96cb2d816d57af21abf0a12d9b9383371e6776a
zb219a0d6cb401d771ff1caeb192961bf7df2dbf517ac11da2cea17ddfa7dc7b31262bd271a06ff
z1fb9ac0cf7c9a3a7f69a06f76fd3ad272ab82e272f9516fbcee248bcd7c078ad44f209e0c51a7b
z40e6057a195d3761ceb82ddb317094d9498ca7c13c377f8671200dbc8d5a6bd10757fe515d42c6
z3f15a3367abfdab07ae4ca475ff4cc607919ffb23b6217848219ebc7b81f46f3710529bb06dfd0
zd30904578cfe130f51133b2d2e04a4ede6ca515aefc1e56100af83737527c8fa0e62d5c0cff384
z3ebd159eb3cd8267a0078b26f626af94d04aacf1b09bca2bed01caf0bf20c42fc3cc7ef74f6bf1
zfd8096e6c90a32412ca2c1dbb19d7210501c453485cbed1306f743adff7b8970d0ccd8b52fd75b
zb951bf5b75adbb3566ae6c05661ab395190d89e2fe5922b06ff1fd84964f67702b874f2b1483a1
zc4ada343e3bb90c9c4b69e0462f8b81e04ac618850c5b7a7c98c91d0f21000a6f423fa61fb4d0c
z6548f50d1b1505f6e2968ae3e408f6165ec8bab7782527850ac7a47f921bbcbf2126f9fb584f8e
z54b89d19f9086c9257ffa35c049ed527059082629dadd26e2a1d29bdbd19be62041c6c4f31f286
zde00ce3586a1b0e9cf658b29dbcd3c159cc8f5a1daedc273e59a0f7911905dadf02bee0c554006
za415278c3574b04ae6aa0ef226a39b7baad80a1ae3ebbde0149d199e9be3e1fd7a2e9e31f759d7
za41306a8a073209fffce7cfafa0348b4783d8d1e47461515428aef966418f1de577e9b79ea6375
z4177b5e739f9e0419ba9763ead6e7b1159c71ab8444e61a8484a0aeb7b60c8c95946d286a2eb6c
zee1da207c10bb04bc690c0c718ff8fd23ec6ac40ef053643aad5544e8652840d1c2fe2383e061a
zfa7b0671566d63bc9b1cd60c911e9f3957f7964fd324258287a227c6c42c2b913faabfa6e4ee79
zd73f9656e4a08737de96aa06d781b87122fed69a49d28495328f7be34b90507900784810b24ccd
zca355d106432140c22c6ffdb3919ed1867978f1fddba1430ec1e1aa1eee41a1affd1fc1ebd4849
z718ed35cae568cdf5435305480703923a8ef4754cba71296b9153147bea6b7583842d923b93790
z04a5eabd082e4ff47b9ca4d595b2c9f9636dd582fde4590895e02a1a6eee89ba272ff52ee322ca
zae24fb0a313d8e2715c92446d41c51a99a046301539ba35187c5e897fe7abda4ed5a9cfbbefcda
z2fc45499e50030dc31bb5b117e2c31cfe65ae84838021dc83289007b63fe17b3efa31b13c2508a
zc4f25569837f078a756dff5f355b1996263a2dd919d26f51901414fd51ed4141a0f744923d9365
zbe851a08596ebd074b0d05e00f096ec351194bd2b81f1b2efc07b4a99c7dc9756e3a83f946e0f0
zad64d4446cff2d2087e906a2fb3b5c6c45f5afb58459b61f34445dac3f8143bfc1eae1633e6331
z158ad96ef9246e3c069f8d2761c5e9ba389b6c0dc756f8a43349399e63931ef431e895b879938b
z37d5cba6b7612e9ff6bee0c8422288f653d9279ee3253fed20124af23fb088795e165a2597dc8b
z87df4c6608a1d1e6886d707303fa3cd41e6970b53ec2387538ebb74d37425e3e934f0149db3b61
zb4b68043c5dc7043c403458e46641e6cd49aea28731c57240ad6268383ed4d449f115928774c88
ze0af3a1ba0a8137477319f2fb84988b71f5f4edf37b561ba767e1c3490299d520d1a484780fd4b
z6f5c6462590d51cced718f8b3a5c74780fc4e51bb728f864a03f0377f6b6ef84f6db8664df72e2
zec81be27c8c873756b64a74f111da2c89fb0ceaa75ffea2bae802b2b1d2b9f3c24c782a9e6e9a6
za7c8b7e11bdaed0ab0b8889ed4e99e526cda256f90e02e95f339dffd3c1b1936b9ac27f312ac27
z5d18425fe5c4e002fca626a55a351c643a302fe463e11400fba2aa349123c21e476a173ca43316
zd77c5f6cb7c439be43227b11c3cf30b1ed01ba94a9395feaea6c02fc02b38a49bbcd201890771e
zf623282b30151aa34753046a58b87c93c8da2d2190c7ad159f35ae2d1f060dac9318affc9e2e23
zeabecac66987372870436521c873e4776628d3c67f40dc93f57cbcefda1c40fea8f5a71b38641d
z58ea5ac69eadbef30c03b28d1db8161873045b7ae9c12507c898656312613ec9fe34a05e51493f
z1210d730a42e469e7e830b55572297bf3bc81b4d9b98c2d53c930148734342ef07b881939fa24e
z760f237722fdecb4d29d1f55dcf24ebc73d26a97cf2a88b22a894ea9992cdb921bd802f6da7335
z61caa115b146a9b4962567c8174644ed55849d50ee3b0887c58139fd6433efb158cc8ac2ed30fc
zbdf0a7c251baed1f77eec5f70c79676d6aacbbe27ac5280ad7477ac3847c24ae58471aa2076631
z5929666449605ea542106a136ca6a4096456a8f4eea2348af081cb710550181067230d9ba82c8d
z263dc1bf21564344a356e49afd7a38fed57a12405f4ef8656aef950f721d36b6a50c0920bd6983
z4dff823d9fe8ded5923a4390ac570714df04e08ebfadd58022674a3a40611c5f459f20a7109292
z3e069eb645840e88f8a94f864f36cfb71593fd9f5a20225f5326c6cd036c1db03dded6750b864e
z89e3b8835599571c1d73c85c1673ecdaebfc751166dfd9b721a7e1f2df36024e355691afe69dd2
z493317de710f008fae6be6fdd999a142391b614652631cea531ea100ba1a339695f1308f3c41a8
z684390f5723e658f3b8ceaa8a6b136ad71492285c62aa2c736bec8d24d6a4cf7433595bb6ddddc
z0741f5f0296b57b326d5490ca3515f0f0e251427b937740df2506ab30eacbc7f865dcd8b8c78c3
z88d405ea00c81d179c7d37c1f14dc2ae7fbfdfa0f6e7cf774244633f55d83efb0265df7a47fae5
zf0a8e43dc2eb63dd62649d4a29d51dc26ce61cc5f6add0dc6bfb33e98644e898f149072a9c9000
zdf696a8a2dbd2ef62ef324c89046a02cba297508854ea8d569f090d1b22d9fd3dff2ccf5c3f5ce
za224a9f0cf9878e3421270635edae10c603a613fbd2c96dddb0fc208c2641279365c4152aa4474
z3dbb34927ee8540323645c2da59d54d8648e8ec2ecba4f5cb1c8bd7f5696f545f9c92b6e127316
zad01daa191630966263e94c0196eaf42fcd500466c23cee0191e615fccd360a9a3f1367999b1f6
z8ccbcd5f54f98fe92e367d9ea07271474a1197b32731a4ba9cea5be8516e2c58ba42923429e224
za51b988073dc2a6eed283941c7220972ce82dfbfc2ea26ffcfa343519a81c412b411ec4eca90b9
z2511be16f5574563d7911aaca0ed43d4ee6e66c5181a5195c2a90bb1e67a5fabb1ad5a19a84881
z3c9f1cb8089fd74d3d99ef03c12ea5588887890823e337ea15d3fa341f551c600031ae20f2e03c
zb4a416a76551bd9c3ce02bf504a73c07880396118ad1d8dd904309ffb8aa8f0ebb92568088fcab
z7695a578596d6b480b70d30da08abfb221af0267df6e2523d012ed238451d15524a2c9d5248334
zf1f93392991743fe7009663259d49339b916a0979da5bb12b5857a8c64b3e6209d34f853f50cad
z2f50f53b0f57864c67cac3994f345ee6880e6d29a6867bdc5415d6c5769238e959c7fff88b739c
z60229377968d9c8aeda61f85fd8275fb04d0945187817de3b7b3d415cf471111358661b1a1a4f9
z0f7bc258f4b53283ca9ab702f08df7775efd9e007625a902c2bb21517797a3ef5c2c6772fe3cd1
zffb6d5e8172d3edd4cc0fa891bfcb98355ddaf76377a081fd0b642ce2f38ff8c2ae05a2221906d
zdba65e87401ca811f405b87abe8a9bcf6ba6dfe4644b9eccf63961ae767ccb9bc8ae333aff0ef2
zb80bf3f04587b532269284375cb389cb2281e180bd5b7fc193920d493b21a759436584c4ebceaa
za7d86b9a4ea81196ce6a0fe1f94d14b2db2b17c99462a9163c878bcae3b9273fc6aecb507be681
z31c2bc8e369004d784c4bf6ee0a0966e0f78aa11adfc3338426eb7225091ea079c249c8b46d90b
z0ed430acb4ba6d0bd2075d8c0cd5e53059aad8a3a0b3dbec045db25fa46f37f49300ac3102e3f1
z49be92a4ec6a9d16b8d042a2b767f74b11d236da8a006d2b481a82550ac5768f97c3ef81fae103
z84ce371d14407930064839872ac4fbcb29f48abe5efa121864832ad24aee4bf85da30425f6fb05
zcff5474f5bcbcc7f20212663bfd6b0b555a33e830247f966d707d5c30e82ed105bba0c647ccedf
z24c1fdd24099fe9af826242060d672cebba7b0ff0cef1d67ef8108b7c67c18bd1c8205390b8e8e
z2777ba44bf640447e6eace23fad628ba311bf0a6777bf7d9bed9ce040778d3bfe3fe44f9c393ba
zbd294e3a184ed9155270d5858c6cce7528ce47cd17021040eae8e1037ed6012e6bfea085fd7ecc
ze000f0ee585c78582af9eba397e43c7109491bf91ab324902c3d7c64db35105409dadf2b68e14f
z8c0e32489b60ef9e3fa9380d2cd714058a9405272293d284bc97656f8dddfd327f153c2ec2fdfa
zf97bf9b24e7dc27c37c2e187077f7288b2c6e470c23852293e2621492b2856ded44927a13cb868
z14232cf0194616c0983ff5cf6fcad191392ba4ab8bfe3e83c641daa8a87e9e936a4fb6f84ec2ea
z87fa503cc82bc7d5bdc16c411efef8b41706ada59e0b4da5ad56e6afb327bc3a924fb6c4732e73
z76652b1b03664075d72864f7f4c9c4c2a3ada0e6c5db3f2ea9db04a1f259cdf9c37b4f2cc25fd6
z0e2fe511a51f9e5c5c0eaa784537b5f00f531d17f21d96113f9d82855cdba74b2e4894c9521101
zfabf1f69548b8d0321ec18165a0cfb010182dae0d5df0dbe8fbcb17e14870c822fdd8bbdae324d
z0491e2b51d3a4eac9a888c3c81826858d09a5056db850b80feb446056af1b0ec75cdbc0a8f4d4c
z80069126b6f8b5b58ebd17de02cd2479135607b806ef8aad662193ffc53fc93ab627eddda5cbcf
za50e9ec544e1a63f0d75bc22f239fb2825556f405ddd86948126224c7cc9d4b951bd63023308a6
zf8e910b89d02b688b0c39e043763e5e4a2ac7983526be26a03c659ece56746d112ab53fec56612
z56896f07d170bf762dd65e782a378f3499dc0d626d23338a43580881bb2cc0bb71d97bbc4c652f
z10f4e4940bc2297858067c031d292df5ff76ca0ac2b48d15856f210ac3f9d5921b7723ec23b3d8
z7cbed6f3caa2cf002af50a6186ad7e96dee8c03347ca3a05a595f315a10a26eb5473b8fa596417
zd81ca06a5b25c62d3f4efeac601b9d7fd86d7af8e3686750e1d078956d97377b602d24fe634152
z9ef1da5617f660852942694d21df66ae5590d3610172dcee95d0d30d5cb43e147d5e218f62975d
zc9f5cc0c3cc7c7b68ab30b7020f4d464153559fab2c396c2d2f79206fcbf40a6d3e17db080960e
z07ec23ed6543e39c29231b69c1334120417234d1756084d11129ed02ecc6270f3fb589a0a70f03
z361a391218833be8be43df177367160f0245301b18e4ca259841415078b1743511f92baf8b121d
z141716622e448c05ccb93ddaa23779f33fa233a2042e387e697bdb2b077bd4f269271b4e2fb635
z1853b74f52178a06007906d3fc10a78b9285d74f4972d9de581856678e259dc97048dd893f473d
z21410a9e4182730b13bddf8ad8f79323bcec9aa5569e1bb0efce2aa2a9d0017e1acc0f0513a491
zfd0cb02182b838615f72c637e2cb8934c5ae2a117688ec4ac6b37081fd63094fcac58653bd954e
zacdccb17298d5cdf230d200d1afddda46ace3efbd243cb6eca79317e0c489de63ce3e49c4b1f62
z90e14e06cccbfbf14baa200a976f2443dd434f6c456816842e3df5646a9541c95a9d8a0a8ec1dc
z9fea91ea1fb09a66a317ebaef71e8b3d36c48a0092417df30d03024d91b6de2c30dc56874d1c86
z32f7b0794569692e0d36d24079621a355832e8f70dc5a42f8f9187678a015b2cd8b0b7e5eabeea
ze1636dcb07830bf3d8ea778f71fd75ea48014a314fc2dbe9cefba830f77f5d0ff692f987c7db41
z25ab7571f84f582020455b518d0bc656d69476ca5637f0fff9ded2594ce38c45871cdfc4484707
z1693c963d7bc8e99e844572ebd4e83e2cf20eb139239756049e827fe96b9a331a879381e7bed31
zcd8818a8521e8636974531cb4fe6b473a78f53f2f8ce5e0512c1b629727920a4661008f6baa124
z82a7a5b800852ec7712063f48e1442e864ae492dd325f280b2965ec90bfd0211a8d62444ea7134
zd7a00338d465523d20e43f0a8b39ed07a6363236450e8f104d89299e52fc0675f652f2f34e1841
z3597d0140e2202f6ae911c3b2418910e78335977005cec344e0e8fd432a511609c48ef5f38ce7d
z3080ec391dedd697a35c0fae8ee6e3b3e922ed4752020eb7d844055369e939ee92b4f2d1322334
z9c413aadc711bd191ae060c4893206b85a1f592d1e41795d42655d7c2876db81a3dc377534a623
z40290981ec2821c31a5ecc4ec47ab4540acc487b8ace1458cee9b2814ae8fa587a792984635ffc
z3a02039c21580fcb1a46e2303a70bead210b2e267fb9443a3433e67e01182eb9a2d7ea74106acb
zb56bb655e5a006c59d3b1e38caf6a74a3495b1d78b93b858be1f95c70590fb769de7fb093e7425
z95e121b5ebba84287d6b75366b00e9157298130adfd1a690cdd6972c5acbff099e849abf28aff5
z8650840497ad85fd747f926c87fa4ad31286316b3d76d7d1002026db9764a73e7b15ea4c8f3129
ze1ccbdc27069dd5eb8b1924a16c10b35bc5fbacbd01e0dba8c3cae52d0d96286d32faa234b815a
zae6d82e2745c70b6463e3bfa357eab179bd832e629e5e16db768f9b63736e1bbc2bd1b7ac6dd9b
zcaf604d4646e2ce1447d29898561636f546c4b401b17936b035655f661d6f4de7cccb5d06d696b
zafff0d410cf68574b226baf9f24311ee6fa83e69b866278cc5c4867be5657ab879ddd466400e43
z88dce0a34d1c18ee858393cd58f74afde62c287e747bdc248d43a28d92c6bb8f7d017f83b5169d
zdf0ec01e38940536eb4c99a7a9ace7d8a049286d67bdb3e2b84d4d7ad1b5ca40c7e00b7447fd49
z8bea20e1086d67aeb0aa8739d785cb6326acc246dd795d7d6df8ec0df5b0728c37007bed789a02
z383c100783a1b072b778f4e05590ff93958f34a85487a22e04ecf575ddbc13fc785cb8e3cbd9cf
z9215cbc02b84bebeb2302bf18294acc1dd7df8fd78caabb5bb2f7a57a6246f03e165e39c3bd7cd
z5d82dc1d4328850914174174025d00441832f8166441bfa2040822c02eb51c5316160309e61ce4
z8e171340b36fae4f584ab07fb15482e38c0fc7eb48ac74035a5ed9285f54ec2369b8b80a20f25f
z100d7a1b8833e2b21e7c1ce183862cd6f8113677ab8043243e2a184f16a2b42c84d406193c50e2
z685a6b1d5d7b269ebb5b53cd7652810d87b179ee9fcba4f148004dbfe160f3a59101143acb37ed
z27011c46dc5fc89bf59452427d2ab67dc78ebb024e6f1226ebb0046f244050bed97379d9875d48
zf838fac5e2674694b25e022751b49169366517b850cf4ffdff3ad2d555b4bc952b6dce058ecb65
z1903cfa901635b4285314b39bcdbef79b7d01c3e8d3650eff90741e4e186db5c39c07322898d4e
z14fa33d6968d957c7e00431c0eaf53184a3a2730dbd5574e3d146aa512adddde2c7efbc4c995cf
z80b9908ffccf4dfae7957486ae816398f9cc74ed1fec155bdcf3d89dac7e480ecd6d6c37ae896a
zc86b36d96deaa8a6ef2a5484c17724dd4ee7248618983fabf5f83108572a1319b79b1efcad365e
z598b76eae985d0be71ad61052443c4dc47713dc368467225bc097b0f74c75e21476e7a6e993164
zf8136f987977aa0e596d301c638ae26f2f517a765f6d5ecf45666a685500248e18ed8972bfab53
z52f4a8b382d4a79187e21970783a75ce2bd6503cde5d443a5a6180eb9ff9655323a643fa3a4255
z1afec72dbba4cd40c66652d98a591f25158c92517f3468dcdd83b1594e888f6fb76f2a3a1c3943
zaaf866f617a13d2304a13ba84acfd0ea08c82b0d3d3404d03a8630da4882cd400def01b5484cbe
zade63eb9895de0edb1d09e893ed11493575490f98471060be8d304d307866853b6229b3ec062db
z9272145c79c4d94f87f8c8607d2a7336b40a71b94fc908f15c3a1182803cafa5884ba91c64a8c7
z40d7d36f91f7e9d354e93e8a0dcf29aeb2b7b63027b11ff433747b88007f391afe93773bb4ea61
za07efd6fdb754f57304c1d19a3d952ce4f58bc890a8718e596b31cc2bf8e9132e4d21bf8e53329
z753f0ebd577466f52905640238765f3c30610361754900a311d52e420891461cd7cd0c2e2f4f04
z67dc70a2457c4595bc7325b744db7c70bdb93aa1135682020bc61063b46b82869689bebf1e0430
zcd5f6c1ed976db2255e35867b035287a524bc45a6317fbbd4e534e9ffa9c150f216b02f1116033
zf43b2bc2f70ab1527fb3d45786af359cf0133dbe4af126a6503797113026e96a0be9de8eb7bcb4
ze5ed21a4c6013399724dcc2dbb9f7e9c5970d7e92a66674edbb7a565855691d7658d03077ec23f
z06abfc05464c9808ef3ce0b0d73bb32cc1249f34d1c4751db40a293263347630bf1cd76cdf2ce5
zdf78122adecf2890d64ebbb95b182937913997d0ba018d2ef18e7c547954d55efda1ea598c2c93
za6c972f160eef910e9a5450c76c0a2fcc3a5937feb100671fe80f8378df6bff4afe4284bf2e32b
z4261a3d40dfebaf33bd490ed5c6cb771cc821aa7a4122203368d3fb8db352552041f688188a34d
zebd511e075305030651f71f78b2717e6a1a63716615fe663aa6bdcd0d00e57ff72ba5ebaab561d
z6e93f008f0f3d794cc1f092420dd24c9db48be7f610a28182b8bfd86842b57a0fa4ae6e365d993
z02f3c32314834de2bc811cdc001f9f1ef1c96506c7470ded818d053af88b711628aac47357fa9e
zb2ab52e579d972a408c4424147c7ef78231039a6ee89ff66c319675eef7b4f5f6c8a4e4e0ad4e5
z1489431a276a53bf939a0f0ceb09fb082bb017d69357689c729d9b3056fa05c5f71a70fb13d8da
z33ca0167c94926c34ef6927b9c2cb741888f60ec17a62061ef2c82e411032dbc4c3dc5a2f7bde2
z141e8a3c1f941b0f9ef78df03abba7350a35699d253f052f4ea7b9983244697d9547844764dc9a
z5c1ccfd1fdf0bf8aafc0c591f2f50df032e35953ac5de165d9f27f8161cca90f44c562c43cd9ee
z38d7f985bae46f67f291d523b04feff2de49b51b7f009100dd40254952c6c5584e05cb7744c74a
z50e9911aedd6624a6a5d04fa1ca64d73191115a3bc094aa9f64d537bfcb5848c7a704bbefe9563
zb3627d588600e3bd673340ea8b8a4005bde01fca95916a41091ec97f2045ed021b788ae71ca412
z9b4ba351fc325b606f32a5f731505707bf3a71125087859fe4dea63034b090dbe180b47c410761
z4b95e8edd57f01f96e012413782b9fbb20a65017b36ec592842e8041fb1b298fd1a19676bee121
zd0f2f7857e954d43a408c26cabf3b880236561c6758f8f3a49e1172da765463439e6a79a8860aa
z96c3fc4530ac257663c97521888b99fafcaa50831bf6cb7d2b851dd968eb94a60b13f24feca2ec
zf5b2253b97b503a272d105dba479882b48689f1d9b7dd730d22e621c380b9e692c7b142eb8f840
z4dac3b1921c6498fbdee33cae472bb8f2bb19482704357b2a08c2fbfa23b9fe9fbd2ef4c390433
z9d60e5ff5bf49c1b6bb4b3e45d8c6e272585c125e652522c9ab7afc05fc266cdb73e6a280c13bf
ze79dd80657d993eb239a5a944acb97e3562b30504495b8191e3bde5491202ba138aa8d2fec4608
zea209c758a1d48b4cf776dcb130234859f8588b641d6957fa33f29a02fe3c35f767b3ba78834f1
z484ee93b0fadcc2c9f5c17440937d44738947d5d785b5d148e5aa117acee1dbd5f5a1c8f84462c
z6d8b55dd79fa760629b606f8176da717c861c9136bd7aee20f235aefa553d80ce84fb1b781fd97
zef99a398a9f601b08f7ed1e948fb7f5db66049b740964bf1cec676f57972793e5267a29da7a83f
z330636a227fcb75c939b39f3ad0567900aa88b57c942cf91cbd09438d4a25654139e2a6346abed
z8672b11281374afdb452e8662de9d7d3bfe1333eea29a01784473a27ed92c6ea342e43d10abcd0
zf06ef79725f8e08a1728e1b7d017a6f9b7113e97dd9d8db94c502801819f35b31d3cbd20a8568d
zb74143b9eb611be80d4ab0504bf48a6a240557b0036771ad84c2594617ec7ed4194fc716db5bab
z0a924b901bdba1e04936653598872a8aabc9920aa9959655ee2646b86320646053dab4f08fb08e
z4d7db89e3930fb7149d5347b80f9b6e9732df3447892e7be03655caac083234bcd98b7d79a1221
z1acc46f3f88ec25e9fdd56fd46dea7ed51d4a9f93b6a8528785565c3874409c2af4811fe7f0781
z21deb9bea9530a987cc7e26a4cc2c4e78de4f73d24fac3cfbf54f00a41f4e82e9047c8b9e0a329
z40d262f8f5951b8e501c9db405cebde8aebacf1dc273436d13c60fe3d163146be759bce3e77829
zdc7b5600911ace342e90956f8e46f2e23f3d143f877319c3cfde9ba11654dde818a6b3a8baea0e
z809896ab0f7f81f551a4c4a82a8639a0300d11b21b1d2da54fa8c3a4d87c7010b68f51eb13825b
zcad7f58c54e3d51cb04944524326347d06daca3589db5303311aa9ac41c8b9e78efa8e5615344e
z7b701346e4f5d7fdc8bf6b83497b98dafb1f7722811318759e58a6ee8337d3296f9fc9b718d362
zfaf38239378cf02b40ca7ea5113ac631424d019698258836fe154dc54e21fe0e3dd362f3965460
zb0273b8f2ad2ba3e3f5c3dac18e34031ef4aeb85f7d22bbd949f85106448ce45df53a955976f8c
z0f5b4c6c73e6395296dc65914ff254836614976ed6f62579491162f72394095a657df22869f395
z9be1b27ec83bd84a9c61092e3fdd9be5bb43b47871f205e7b7526ecd88d53cf68df92ddbabcc92
z12be2490c428f4734a5a3969743a842f45a37add11f8135029d7b2d6e55a255724ce449089253b
z71ddb830089c7662acbf663d10f648bd8bcdda0a789f4b67f1bbed568fc9274edf8e36c1d3941e
zc9db1a5cea0a6920da495e1804553d5fea0fe1d9a1b297398703058b6c46e98d58194447417f63
z58fca7286a71d8eebc584f41ef9c3486283aba72a256baceadbe71647cf851de160cc05337b764
z21573628b0018e4476c1cf42fa0d4e8d0634ff5504747c22c79c3d7e5c37a2a16ac526a9ec2acf
zc3dfcc068faf0a10907e4e8f1f09dacffac69cea1da04e9cb94ed4a2e7a43d5fb0477001725fb0
zf6a8e52d5735532eaef4b3c1e83e24c18146b72c643633ba739cb8ff3bb181b741f6ffc055ed07
z9b0d1c01877b1f5b3813df9455c682767d58b6e31da59206534e3a8900914ccea3026abbe90701
z0b98bb5c0e28cc311fbc05a520c9b2277d793fb74fe4cb85a43e923493ce5248c202436f4c5cfa
z166ae2a601c1a917d8126a595fd83987fd745a8ca996f1bf3100995202fa39be060d9c764b81a9
z235ac85c425a06dfb84c1a842b0006ba59497b80acbdb1c6f4ae3f0d91ef8c6e18be17d2369f0c
z5e0dce5c6319669a4a2c744959d4970471f53594b1b0f87199a87f7220f0d8b713a0fcea1bec0b
zf7f38c2cee3f469798af88bd5e32c8844bb19f6992e6f30a6d960ebdc1f1a99d5c5c00fc781730
z527b1a4eb65f05c81c5b0abc3da5765f6ab64c487da0711e4032f81269b68ddd1024cd1037978e
z0dd568670f949d320fc767fca90e994b209a267db6b0820ca0e8ff5fab20b0d75ab3819e4ca1be
zc7b5c2680b9e8a9d786d5860150bf1164f7d439ae347f22e14b0158ac51b2a944678806c78d338
z026b94291c1de50c5f6aa8e9fc64ca89b0a6d57a6b92e5f930d533260b04df381650a37c0b0af0
zdcc5d5dae273a83e6ee5376627afbbe3e89e6edfcc56b4f5dd4d220141d824ab764a9f8c9610a4
z998c5fc7fbf7954eec1d473efc816a058a6f2e22068c35af39703594dc74fd9541b489b7a68b76
z466b93a820f408238754c856e9fe8322388184fad350ddd2b32e929c2fbb4f396c03a52e2de249
ze8ab4d15b45d25527abc8f425e5632c186e0a5f2f63f9e3975f2c7da90d42e60b1f6f483618d50
zf4fa099d7c448e9b00ebe7b1a9216f43e52944f657fb4257955f8ad79bf0ed9028aff1a227a57c
ze9210745be18e7f89df041bfda700d4e811d2cb2a4cf91c3dd05dcc639b0386f2db9897e2de7e2
z6b14125a9f7e3070478860706df277465221bf83ecd49efe752b66f061f276d26ee317bb4559a5
z20776d4ae952e394d3233f80e86a25fa113f0d30281ddb9b7e36943fc69dee8651d68a34f66575
ze3975efa7b887984fffe07a8d5697cf578c4be885f75492fd969ac13128e1fc0d413b415fd8ea2
z1f839bd69e0d7c5986c21a7202d8f4f914940fc2eeca65e128efac14ab2d886ee4735d6fc20bb5
z2a0151817ff6bad44f436a314787f60c325e89a7930f47cbc9a2c2e2946ee91694d05c8e3dbae3
z3b19d4cd21d411d3b3edcc20c62a912a7197b2d6ce5696bba9ced58fdbef868ff7b005e0b2a138
zfdc85c5b2466b87064aeca680e081ccab009a11f3d614038752d61ba919f6cb945884ed5a83f68
z20d1b440f8bc85eaaa75d233f2c46e2d34a128c78cc0c04580d368dee376d8ed0276636f55e5db
zea5525ff26882f80df403d0626fa3fb1a2ff116a957cc530fd537009180091b65536ac815ebe28
za60c8f2fa0481275fcd1bef5c2b6259663ba746cdaca5c9136a8c55f521da075af53bfa8215e0a
ze20e83338de1765fdc74fe499d18adc2a4e7fc343264d7d9530b17237b18ea3754568501aa7e94
zf2a202db2dbe0bea3746841b529af23366bc9459eb45fe98f8dab4006903f663d0e3cd366477e0
zd5ac8b893bb55e22e5bd8b5850818ed4b6cfa09fb4e248e121f88ee8dc8127ffe0b02c78cedfe9
z235cf1af5fa0ddf789ade5e250bab743031eb1c18831b156e3cd2295769d810083f0f21c7fc747
z369b81afcac7906aa59cc1504f885feb653cc66926c2d64e7c0800ab8be617a24a104f692c347a
z002d962cdd2f74ce04d840aa19a218c82c3f4785cbe3f3a73efedc02ed27eb5e8d8defbf9556b2
z88e0bb6a0e3abd540d546b541b03574435040ead2fcb9af26408697601487b373307d7ee0f4f77
zd07778eb9579b105d0daba5aa6090db5bd4a4590e2bf3de4e8a77aae7944dc3e595695a52f4fd8
zeebfafd83fe7ee8a743908c01ee3353055bc9d27349f6849eea11486de549b283ed157ab2b9552
zf4f7df11782796b0b7746e2322c6a6da6dea72fe7810b38c140a59579be60f43e7c5921bb312c2
z44fd0f999c5b70b6e679e9ac5117a693a8b4f62386072fb655da4e7e037a075a89758e05c11331
z2e3e08038c65c98964b5c2dc94c1ca4c6306c4548a68d54be32fe86316caeb3bc9148efeae237b
z9f92cdf92b71a84aa7cef18399e4ac36f48d35c5fc0145df172c3f6eecd6012c7f57b29539032e
ze18a33b486fd1061b620bbf48cb698874b317e10b526d4f93975715c212aa63e08fa7258637004
zd386566377dca1ac665486af06a9123db5efa06cfcd45585c2afbf7dec2beb5565fe5566edbe83
ze384801111bfb11809311d4fbfdf212516fda341ecfa42e8d310860c79179c9529aacbf299bcd3
z94ec864f82fcaa7f1020a5c677ccee512e7765dbe4b8513d1fb8dcabfb798e92685dd9e8ed3737
z7b9e911b59b70e43fb3ae20eef6887bd6c05e784eb326e56993366a19181bc2443c45f404b25f5
z60ab81376543f14e64bc442447611936090741c045207c893be30edb04f5f75a7bad6700631351
zf73721622a55d9174b5d82c5d387d3a836cd42c73b8cee5b75b11d368d52cedf3df75a4049e5e6
za027ee9348fef25c6940d87710e494d55251225af9cb5fcadb9a0817dfb48ca0d47b17885708bd
zf96ee5edff830679a597a4bf4f96e654b9cfaceb1bcd158d5f00f41b70f4c74e878339b2bc3a54
z46cd12be82776ec197895b0a13c6b4c084e5c4bdf08d6e4c1bc2d5d2ec0f28d7d5f887a9bf6116
zc409e2d867d0ffdf3af77f8b64a99dd3e65750324435210467dde96fac77cc8a001bb54022daae
zc52cb6f0b5e208fc64ec1f3d5661d6ade31e723ab213c39679bd68bb92004bbae23e21cab6ab65
z20752b3f1f044cfe38486ddc4e7845b1244e11407dfa68ae98e620a7078972595c56c8eeaef3ae
z683a3d310a13f47014d18fb8797999fb8b2a71a12c197f99dfdb98092896e94535af1217541e01
ze121ddaf31ecab40325407104170cc24ec2a2325ce2d48ac0da98e825646ac6def932dc508246e
zdd747a17c3f8c297f7d365beddd5b05041afc9af6bf3b7970265b34fa2c7b1548e36179877403b
zb5d963c428ea2d1db41846de08114dd76a9dda1ffa1b38d91b8ffe19b4a496544acbe348de1423
z7b69c00a4d6567636e4672b7686905fd2751219048b875d85ee643cdd95d1ef434a5abc5a750e0
z4a4c251bbe2e0874e13352c78d0434afe16250dd3e8146004a5d89a85e88803c1aa269e5149a09
z078e2a6aad4eeccdf1070c3c3cc6a22e07ac6ca6aa809423363da27748a8e514147dc6676cd9bd
zc9bcbe802a07bce9174ad167eef4bab118d12a1efe791c7d273ba3fc25b551b58203287e0e94a7
zffadb186a0932dbab3b04eeb6678a919e144afd7cbb78fbae44f00f78d3ecda4ce1e3f8c1ed631
ze36b41c0001a32ecc7540d47f8f179046a7ca2739ff86492437b73faac71c6b081707e08ecdb09
z6c25e1ca8df565cebfa1fd9882946c8a9fa3622054ffea1f87132939aa7888b85dd1419508d87e
z0f9ef7fea8b1a6af52b84c5a197f7feb84cc708b45c8e5001db4793770b4863e1bd1e4ca02d76f
z9b3ce19150dfa7dc0e77ec4f8d005d4aba2ac20ee55f8cf6245cfd369d44f661036f05227e32de
zd0e1ee69ecab45a65bf0559b6b438b24f190031865bfee7f827e4670282a9acdae554c65afd58f
zd6c7d0f0cf3f8c91f7d81537200fe033f95534b54eb266736951c608e17ac61c90598f57a7d865
z9305b7747f85f18c6c9ede2901a1fd9788c47289f9122c4739c23c63bee9762861adf24bef3ea4
z490bb932707dd4a2de7162059ef8849a819ab14116de30705ae9393f4941357645e07d0da9a47f
z5279d89127e704d80971fdb9fa643d347e233caa3941124ef87032ba5f7f09fd356da56d8a68cd
z89967ceb8c6b29c2d27e47b35cf151b227f96430095e117ff4d36cd5e6d603c660d66a04934beb
z76fb53bd4eaf84770ddb48d83c72797daffffcd67909aea2be1b5094dcad15940cf191f61aff83
zcf13b388e46eef1c2add25fbfa6939a3c0cf9cb776be3dc9e14fcbb2521099a2fd1ef33435ade3
zf4e601ebdf51d1e78139993452e66425cf9d7234ba8cfe1f062a9d6450d5a33bb247ee9d351fdc
z38a6dcd1e6a60dee457ed4f0de3888ae728bc095d4a2b8a93e95fe178397257820bbe309e84418
z5abf435355da8578c589ffbda0197da9ec096de5fb8ae393d7b0807a7c386cd6f43ca3847d5574
zd1168b558384cce0f646ea7ce86fcf0da430d27d6c72e87974cd6b6002f0b3f691b4d9ad6e7c57
z225cd897c750a9d85eca4e25638e57e2226fa37be0d4eccf5f54fa4b0f39ec76add254b5ba3594
zbfa8efa61e00624fa368dd6187435fc97fcad61eab38c97d1802007c94a60c292597ec677fbbe0
z49d8df8d03bd3447734e5b8c5507626b59154eebd4777ee3cefbd3dcb8399e574d03908f7fe3f9
z188dbcd14bde7157fe1170c47a18799b7d5bb585a5b12e5cc1f3805b1e747e0332e84e50c081c9
z5c7e4f2fe2c6f36ea892143ea83fb4b1f5de9b2a321102bd38fc8741ee45b81d0b37b495b9bd3d
z65b73c190b2d1d25821993a79c71222c102a885e2bfea0325615ebfecd1c5fa15890a63ad86156
z3f91b795ffef1cdca8f4e58e12f04b23c827bc5c24e56aff0458b4553d8092cd043afeb2aba41c
z49943cb5f3035ad4202e264c6a606a674749efeb32d0512b282f58eee9eb08211e4b291bec6e85
z49fdee6c26c7074b0a0915e7b786a12cc2a60f6a419439cb028a8943665b47dd1139afed87534f
z65bbc3bf7e11d0eacad1e88bd9cbae6a231da36daf60348313703d1ed940db2d237e73f627d155
z43a6e1fe13bd8bf1dd5eef6081b5e987eecad320233b598d635abc639b84ae7786e1d088294e57
zbe1e21f252a24a36ee847f300810a95ddac6b699aa56696ba9b0fb650770958e82417575e6100a
zb3d43bb4b09d40e286548942cca4c003426d15263badb8771fc86c2a5228b5517c2ac3552c02c7
z0708def08ee8ca1025c4ced2ad2120ced22062af6d36cd613a09fac83d86893a9f147037b59439
zb4f0d8bd99487b641e08c8f617988c230062c4ef474e19b0f4e4ed08083e3d9c39e6773584c1b9
za6931a1f9f0f37b9c42c4fbd8122490c650ed87f1c01558d81f8c91cb53900f439c945aceea59f
zfbeca42618d5ea8a8d89f3833b700bbe278a8cbb12078f271ec453c89b4f01134c969ef1e9c7a6
z7fc3435b3684da678807913c1cbdd31118dda38273c9012c5f391aef90a6c798c80fcb135e9809
zfcd25d3cb84366e3159edd3e8bfb805c48d9cc08c4d67d0ec687c9eb411af884c99d35313202a3
ze6a739f14a6747ee3c523077dc873a12c04ae6fde133563fc6b793c0fde1f8a7583833239f4066
z90c071dc5791524209aee45fb721027d4bcd086d880d17864094580f3e0c11a76689189628116a
z7df4b8e438340a8ef989e705a16a09e751993dbfdbbaffba1e377c3437411e20d92584b164348e
za01f72e02891fcc0c0223ee65a7619a3dd87e904a295b4a6d0862e0706f7a5f34399f6b881c25f
zb8a067cf51817b15d5a13ad029ac3a61c60caa78e630ed011950e8eaf4e5c6404e5b853031f0de
za8a800d40ff53f96bd3e5e6e753241d29a7baaff0c49feaba779cbfe64b9e2929f1dd06e765e37
z4478904e71fe76d7f5ebdb8629a7160fef28f6508328f2a0bc8077da49207cd970eb4b4a7a8a2d
z72a568f61b919d2f6b1b40903c427ca782d2b739de0589787d6fd12abb4d0718fe1ac4989617f2
zcf5c1724ba917681929e5a9a84fde944bcaeecdbbef1053fc33dd9edb3410226bd4fe44be2caf2
zbbde54a55206576dfae89d6630f0f76d6e2f363ff28a483bddb9b46093c9e29e979720d98708fe
z7f6f530b3201698641adf616a81261c9ff314bae101457afc381c8825281a3ab522918bb2d8f65
zc2397a3d2f479619ffa1faf4bc48fce4261d87cfc8e0a180dc6cb9db6fc3a77e9b769d1be41513
zaf8faab42bfd51c3cad0597246c7cb75743c8444ed741eccf29fc60e362353cdc93193659a515f
ze511a49e9378cf2dac817f085285ba943fdb6e95658fea663b7e0ea7ece779500030e8349d0c11
zdbeb627b5d05dbd3fbea045328b7e9ed9c975b88d7c81571d364b56231a03e1599ae3ba4c5f2a3
z0f3d68612ca4e39a407144899edfe0ca8aab2d4ab32dd8eb6bae0c6b810329adcea575cf55c5e4
zb3ad7e3c15241c2f56e8249234ad76be92ff88ccf3239e95c080edd71574433c7100ee13306431
z83005208249958ee4b26f13fa52c8ab11c2caaa9b7093765f0863557baa8bf8dbbea54a653e698
z9185da34da9e4467e6051173ff1e5b4e56691e32c238c033967b9df6e6c97cab9cc5c2c47e9e28
zcc7c9178b75f844f50c2e3ee1b3d470c3e37ef04ed349970648c682407e1e36ee39f1ba3187f4b
z4b0f82bf66176dba520bd25124cef24cafffe006558d7ca838d611254cbbafe3cc212633b30648
z5f579ba1b5e2ab7e532ef2ddc94ab3b04507b092e07609786677e3cc4a785f260662b6bff3a874
z5aa69b3b6d6d20b648e21ed9adc4c8fb429984d0e6214b32664a36e1fdf957a70897a192335fbe
z3e94411ff31f781c6bb0c5878beb1bf2c2eba6e1a8b85d11479ec9a81ec0b566a7525b8a754b5e
z7abc7b3e8a788fcf1470d1af6d12683c7515c4375c4b8802099ee6fd510354a1dced031997a244
z4b083ca4c2444f164dba6910a33fe68967328b0c032ac3f86f7d4bcd083a347c616b9343fb7f80
z0962a351d9574c31ca0e5adc841337a3b79503944ad04246efd60d62e4e9cb89a43bd5e186340f
z48cefe62d18d7f26d87c7a3c07f64f2a3350fb104e15132ee7e7c644bf4431a0c0dd1ba4fd2928
za7360586823b41f0895a07c993f9b55b9cf565d3c89800a128c7f8974780ff184ffc6ca51cf532
z5db7c208c691aab6f0cf141478f6ebf4be6e38feb497e1d4a1d482b4c3c4f4d2a60e8be3f78f8e
zd27cb68019eedd36eccb8445505c1471c3783a10c7695a14d05b654c0a183f1fa4cce717038764
zf46c92ac52845b7ec8b2009f778bbd502501f51a5747690010af5f2291758a7d2f639d80bf5c72
z07a9ba49b77579bdb4f4434924340b6c73c9ab9baacfc16aaf2771ecf5ea91e4585faa5f09a105
zc3ea652bb09569872bf4a4831d14c0474873c572e1104e40ea6a76386b6fb2ebe68968703d68d1
zb1959e8f9d2bb155d7ab82ad499b999c6825ab29271ca0712a7422dbc67b08b905169ade3e80ba
z66cc3b2310f3d072a6e182caf4ff8964f5c7676b913be17d55abe133cb38e19509a2263b28c240
zde8426b727b75a16f02f3f08dfc2ec5ede4dff901433f29a7ed266dcd4bac7f5041f98a9f4ae0c
zd5906492b140483fb6629a8c4669cab34310f3fe2e60c31ee180037d9bcd6363e4c164c4cd41fb
z6e65a9128f017b060a27da4917e60419d47461617b9ca4ebd7875fac676877a1ee814fde98d499
z63670a26a0df3e32fa48e652a52ede2e3e7b5517963ee6d7c208ec0c8280f5aa3d418b8f14afb2
z67af3b72eeb5d83b97ef4d4239b1e6b92157189b068b75fa8c9b8176440985735c72568bad3e82
zde01cdb65c3abdd2681ede052cfa1cd430947137bb936ac79721d34bdb3bfa5f541f71ad3c4e00
z54b161123a7375e6b0c34ddec4e5491ac06a83cf30126a48f74033b74c58a5e9e425779ee98e4a
zb5b425cc1d04f37c22c7b33ffc240496cd793b2583277481cf2eb6ded57f11433640557784aab9
z14e83b95a7a22577ff242574d01971ae900e0a0e194ebe1e7683f7aa845e77dcc2513f47956414
zfb35398b9cca99fb0678d4cf5e7c487bc24f32fe1452ba324be259f23503245ea5712602ca9a92
zde2d16d54def103be7e56c50f835d201d6277fee1e8f7c2d957e9a129e559a1bf8b7fc34370562
z649c55f06c6f3ad50dbfe26d188755fe12d564972b22564ce28a8d5739bd9e40870566bfed49c1
ze8efa376c804cdff8f2cee14c7236cf7fde14bc050c1f3b1af5e256ea3ecb80b36ebf5a69450c2
za368441590af4483e6a64b0466916f7f90e22c996c7f915e5432fb58bd5d5f5c60cafa73a6f05f
zde444891c3db24c44f9f8a06fc345b494a2f12644c660d2eba47d38ffcbfed5cd6bf9f7ae0744f
za8a18a7660a44ea13c8fdb814da76dfe875cb2933033896caf6b4af02326e54d05296da1e6cd54
zaa3a03b858646f3ba3cc3a4721011663fd1460f97b95c27f8f40b16ae3dfee3ec0fd8ff3fb245e
z9d0cc13c40a9e19f88b5575e357ec52c9525535c8cbaa9f4dc2af9eeb1f5c3ab34c7d6a4054a0d
z8394f1ee3f68afecdc94591898bb266b70ab3f90c99742b84818bb139ba627b21450bace69f96b
zae4f95f4e30a0097b3905e1eb34de1a458b542374aa8a656f6f9e8c12679f49bc30829ffdb867d
z6ffe7544ffc9eeeb860c093695e033f2a06070a1164506c1f17340ab44bb0b829059ea430da21b
z39155fba019495aa158b2faedd04cdb142105b09ab3611152550ec728f0c2407f8374b86b20735
zac7d10834c6ebce017179ede7d04ead7192a65bb6db1a42779fc3c55a22393c9f4c29a695904ac
z7e3b8ca7f872dc2642e5cb04d09f2a4163c6b81e4cffa10e8e05ea1045f569f37e4f11404f6ef9
z9ec11a1511934a229871fb74f90d832406f101593263c57539db2df56723a3d7d26d6c234550c0
zef2701e73135d67ab053c98df3f8e86ad669000ba70abb7bea57d90a11a1aa7e8762fd80e6cd9d
z21ea62467d1f5f74cab6c496ef642d7c91597959f53a9e05052f8e1b80295b6a463ef948124965
z1b01b8754c84913fbdd86d63f068d6bb0d1372f8e99a926aae1f7ea0eaf394c88b299a5d7fb997
zdae8438f8d98dfcb4206672b00c353dd15470593775280bf06c6573f15bad1a50513d5f53c32df
z26a96fc8a5893f28e499ec7be455811dbadf1da5869ed6e71fbb8324a853357cbcfee8494d1f82
z7c778c794663d2c5b32f190e092635a131c283be986214d337c40fef0ee764aa93ff678d6df53d
z26a0f94eb894e1606f0b084d15bd1bf6bb816cbbbcce1f15118d5c8024661a6dcbe716d1df64a9
z50f7f794c0cc96eabc3cb18a3eaf00598a7a9aad6cd4822483a6e6868d3c9a3fc3054e1468bff4
z7b6814bdd6a7049d222581320222437891a49d4c2991faa1929ba49f673330b40c4539ea0888a6
zf5972d1d52c412d87d0df56e3444b99bf0e8c764ca7e3d16a809c11fed813895d07b576278b8fe
zbb87b4d6af09e4b6e3a16f39d2acd13e5adfe8e6eb9aff6f53aca1c535061bf525706acce34d5a
ze7d5da04cedd10681f7c6506920825b8f3dcd275385d02539aba2ec484054179bd471a7b393b36
z6dd51080b393ee1da8bac70467f8f5ed0fab0e8b984078f7f8cab9782a2b9a7e3fb0917cd53412
zefc01054942451ffb1c34b2c8ef18994af74d51e5bfed36f0408b36ad5a25b43e6a87ae5b00f4e
ze9a0e842a5cf1a5a449985045c53de79addb30b4c3f3b76a310be72c2b9b374054f83393a33e01
z62fdd6a44b9b8c8b216c4577cc0870e19d9edab9981dca500b907dc2a5ab86712f06dc0365efd6
z112f21b1d09f384a729d9e40f514231804887742c57bb79eda0a100c4cf6318ecbc98e554db643
z2b6840ab2416cb6782c0590d9bd0fb51a25854a775c83045fc9f5003f68a9b0b9925ff5dbbb114
z0df364a677539969032df4696b52ec848be83bcb9578ef22fc8100a068b2c7827028461da8349e
ze5a95327b332eefd57726a3d53d19826dc918e0be4fa528396dab13b771bcb7637e1632fe1456b
z7849fbee59ee98795f9dd25cee0a07b2be2f659fd268a8d53d32523cfa15a83b6f016faa7ff37c
zcd53cca20b6298e2fbb282c9fdeef7853d44319ccc20d5bcc9ee06b3c9c8db41025ec08e45dbd7
z335a4e76d64fafc46e0ac26a794f6d22cbfe9e3920aff2e030fcdcd632b4fcbf3af93b831a862e
zd8850a5d84a4e51f8cb8f2df7fb59d201acc8c58b9e01d57d6edf9ffd28f4a740d090ebe11a256
z3e9620b58ae3b1965c9f6a64ce1c77ccb269d8674ace34f937723fff6aa84574ad1875d855416b
zc23ff8e67cdce6229b0f8eeb78d18a2bd545f8b467624f9c5fc3a7556d4375e2900e1740ab2ca4
z8a18e8a0fa5769b9b1dc010ef366fcbb27341f0d5d94701b3dab2dae5465e545a03b0159cb79c3
zf2b6e524fffb776a965c610bde872322045e63e26eeaf1c9f9b56dc8a5a4343a0a40138238cc10
zd82d0c3caadb7fb65df113839333bed7419793a0f235ee8b26a02cba2c10279c308f3b4d093dd5
z987ceada827d8ea73ff49403997f838d5569715095d922cef65369631c7bb38d3fc5f709278cf0
z5e3bf492eba77b2169649cfe5626352305f0f24af4dcb9adbe193ce17cf18135c32ac5d50e6193
zec29e3f189893f61272cf8a96461c1054182f62289f3cd109984e80941426852fc956aa00dc93d
z111c7e05d3795100fa0bdd867f23099e2673fb7c745b6d55420f7454f96d522a0333dfc79a4980
z2557635b1d064b70e0c416fb48a4803ad3ffd92b2464bd16dcd995db602da1d306f1f53d30b575
z16e99210fcb48dc0247ac0979d7b9328371bb9f52a94818f2e57fc3a315a0fe46fee9cf1fc7c57
z814f5ce8a7e4d5083e273310d2637d77a793da8a8f74bd63943e6da188e87663d91a274fc0a897
z6e6ba76b464b8f0988a609c8a4a0f531659a780132317ce0e709aef0b81c15b4f49ff0e2732519
z8ea6cde4001eeaf87a83d5fad5522f4dbfedd77d2688f2b9b2909e3e1099f7731d442ca55f781d
z95c5ca6c4c8088367f8b3d0e653377de3bdf6650334a28be7a414d7e10a06f98303c299c7628e2
z2f3a0927598f58e51e170588756a8365404c083af07125fee84a222752dc85c012df0955d1fb84
z7158fbf8707081ea7623f9c51b45244facf41515215813ff144eb60ce990d66b77f5cbf533904d
z2c3480d8888180bf7ab25f7f2685c8f6728d146cd1eac4ffd329b328a4c2bc089a1fb5f50f296c
z62618b613d8df400676918d63138f8d735656c52d56af318501dcc5c0b511878300ddac6dd9368
z073caa37b0d338bf658af9fbeecb0e6325b2b88b765941e6a58de78dc6de3e854bf2289af85017
za9e103302fd9733981554528214c2745c1ec83f39d25ddc7d38a1446d1fab96699067ff3d25ef4
z7fa3d951810f9276fc859a684d1357a15a99e5035e5da62316f3176b22fb124d1734d1181c9cf7
z226ac22d7708b47f0bf779b9a4f11914294bf3cca52f94dd878666f9465e69242b917ac3e45ddd
z0e15f2d72aaff3f64ea2ac7109f2dd05bf28025004df6ca8d6134cdb8e483f985fdd64dc60926e
z7cdcafc8e89534e65a0147a81fec2012c2ff2705140810955e93f9699814454123cfebe169e0d6
z13a988eea1704e9512b7f5e2703745edb598c625c4dc78eabaf09216c4f793fe19c0c7aeaaeec3
z88369909c5fa1e00eb71c298f5a261bcddab6ed5fdad195e394f54f71c8ea852f0367987fecc55
zeb91810ec6395c0657fa8242b7fa23a62373fcf933648bbd8ac0bca245c9bb88cd4e06a2e1e8bb
zc605b97d8d948148b977fb02070b8695afdd64d9279fded190c5de8aee3ec1b0e6124dc0cf4652
z06d0cf127e0de6e2e715c55a48430446f6917bb35b81998f81053223c60fbf55a139c6a0900e02
z8e4d7d5dd19f6c7d4920d0503155e4741e2827b17a8222d0cd1edc17780a07a79f04a5badb4906
zaf560afd76c2243623c0b82a3f021ac51e81746259b804906f7365ad91c20643017d8030047432
z701c49ba2359d8824b05233af0c72da75f9fce1f25d77cfff904a400bc6bc211df1a21a3a87e1f
zf3081d28a6e55de5ded30c8127b45a8d2da7eaf4852291cb028132914ed82ed75f7097d0704e79
z084b40b8587991f98ac931413c6ec2d6f2477b18bc2549466581ed11edafd1ed74d39f394c4a70
zaf646ba8b4cc0f72dbeef0143632cdf9c1f5ce583de24c9269abf19eea9d5c7cb389d31eeca618
z1894a28e0d0ff204d56b83c0f0e9403de187e5690dd6c8c37d06ffff6544427c821fa65806c2c2
zc2e07aed8d3fd038a75630a24244b4c5a7f4ed733066e8481dc5bebe2b714ab8489928a82ebb4b
z5f34ca1c819a33640274eaa634208e287f6df90a0f51ab310c3472efccef8bfc2c488a02ff9d78
zfcaf73cf8b03409333af9b74e8997e4108546bc9d761e29a29516d5ae23b4832b89b70bb47b495
z8dd57b0d5538ab81b82c995147437f48b07255d4ee06e7b36e7c113ae440ebef1d995c36a8d19d
zbce094bce2b9c1092fa745733d243795d7b58a19837333a8d64d601f5395a53169e7a7e95206c5
z0bd6b6acf59d24e67137dca6b6fc9e1a598dc75f2a8f429b13015e627ba182935ac8a7df44b19a
z88625c1e8c8dca53c078966d41a850f44ad697828b9bfe906c23968264670569120279174b774e
z3948f007fc08ba4d7ed96048b96c42372a0e2daae102e307269a011efb3518660ac7f5edc99125
ze83a07a09cf6562555a3258fc3c8cb757ed31326651c067e68dcb919d1e4ea3be48c1d7bf62b79
z9acb1265ab6b50cc3c3643f3df7f19fe4437d2a1daeed714742ca8001821f29a5ee4be1cd36422
z8a14906bd074d2de879d97542ff060bde3ac30268eb44aba6200a718676667ae8c7a3a05ab3851
zcf13828acc589d5d154a0d90dcc0cc10a0b0564b8d6e609d447c207d8ac8351ddcd9cc2f9b22e6
z75ae8bd188afef6cad2d73981d654983cbd378150670293a096042c54a812c1fe0254b22088dd8
z0cb9a3cd291f4739cc269b245042656aace0aef7d06ce1d31d641a83f1fd9ab0ca621045fab3d4
z1868b40e2ec7a0ab60fa8fb2d50ee94fafcbd0b41e793e094fe8353b6bfd643b39259bb6853066
z9cdc8732f60e9a03fbc169288b93b8ac83e6129e45441292cdfb6bb14ba197db167df788ef87da
z8d0c2a71376432938e9c661f034e9e4b3ffef7b4384b9455c74f621bad2946caf2cd60570ccbec
z68a019c28966973c679341b02bead63abde21f99f3440c784e593e7953541354e1b32971b0ec61
zcb9d18356f1f9293b33dfca53c40b127d1064a2bd6505710d0632107918e0505fbcfb1c756e7a1
zbea82e85e9160845b094eda47a657343c5574462ef5d2da05b48d50074adf2b56c1423c35f6e80
z616cf0ed32ed1539a94ad718fcfc6029854625df95368460275182a8635af9b8cf72261b9b5a66
zceafe6c7a531233fc30d9e2f6fa5c9d1cb7db5074fed5dd3c77b71c8f2a052426cb1e8f7d3db70
zf648ac67cd87da7f69ffc606230bc4d1b65736a8afd49c6ab1ce2a816182521440fa559d695eb2
z53755fc7f26e461f0117ea5ff0e49c4dc26a269e8738246fc26d71d27156790d75e55ec8b30f5c
z8067b1953ce723168eb78064e83b0a993eac12a43c98a41915738a90ad5c19ee00650fae2994c0
z3b13a6218ded9b43b9b36aca0037e531ca26b79fe4337acabce89477b9a45756832649f540ef10
zd79dfc4115c743e7fc4b408438311493d385f29012267f20ccee7649708890b57171da55afe625
z43fe2d3d097bcc400e9a62d5c35cab7613981e2cfc897c6ea188c1de1dcac4fab942a0cad6f479
z1c0b8deb9dab0ded9db6b5281e297f94f00a738199cc3823e4eee913a560cf725bc3e1ce2eb545
z313f7558862fdcd220079dd41bf0580d4764187fe36cb6a2a541053a77808da4d19ed4cec8f699
zad97efa5ab0b7c5b1d46798dfabd21802a66414398eea474765ea54aad90eb2c3b48d9792d8d2a
zfce9d02b68aef41f52860c5f39843fb85160b2c6f7972010272badd3ffdc0dab52d896c0c13b75
z89504af66b2749db889911e9a3f91a77b039c8dc09e1b71cd10502151904c780504fd624f1e9eb
z1e8d9b7ecd627a44504019a94f59aff301a58c7d17d6b4f334a6a31c4d5bbdf70f41f88252a483
z273ea131f631ce4efe134bc510876c8a312767879eea53fce097aa872e6cbb18b5d1db7244aadc
z4f9a283da30d0ea38bad20ae71db5418672c022c5854cbdb6a292a3f1da6b2a138563a412cec62
z4a6c1f59c4753400a77f6df2bfdb33a7d86d9c1a96069edf712c2b0bcd79bc157944f1ddccc07e
zcbb5984502854fabea96ae60eb096c048704ad93d916078869017a47df07409d6febadbbf02872
z312cc92a95d47d6c30207d142649659a40e6891b9a72a47e3d399fdc54c7e8b9332a10c9e60940
z9fa9e714aeecf30ec9d87e77399f1f1ba6dc6548b60149215155453f76c797adb2044c42f5c542
zb1e41aef1244df4fa40a744f2a5aa5fb7f550975a9262da75776d038e8f75b3e8cb891403af44e
z91ce0854eca95e1a394d4e5d31e1e79da8a1078a4d43bc2305d78b207816cf3ff8963b0f43df79
z0db10917e4fb50a7c277849b95127793a596a5bd11f96277120aaa14ddd985047db79ab7035b44
z149946287c31f54cbb03af3e7d2dec99fb44b0f2ac2d5c13e137916bcea3a25c3d0dfa5efbfa12
z19ae36d08b5ee9b090d0236cad5b0e5030690e2423e9b2ad281817ab3ffa366b10881911b8f8b8
z098d1b2f90202e5a0977af3aaea2ea1e5634ff2ca6a84645c3053f57af8b4248b828e663817e9a
z5c566f65aced94c1085e3559cc3307620de4d7530ae1160bfc3ef37fc234dd6b07369dfd179c8e
z7a03c04508d481e24f97ef2ea443c6238e197cf6c411986476a632212b76ce5524b395edfdbfbc
zc0c291a8f40934ef745e5f083ebb2b2e13e1e975a2583f3f0983190410e8e99b5fa834871e5423
z4e94772592ca24711b1ec67889a69ddd232670357fb4265b9170532375a6d546520866adfc0512
z5d8f8f92ac0bdfbf384f4a924ef44c084efde465790e22b21234a5ed6bab7546481f2fcb02da46
zd64bf659290457b6d1258ab29e3691b4b398fb6c0bb0003dfc91750ff6ee7f99d8905ca29146be
z02d23c0e6d98a49052b16a509f1de729ce07365e4631cd85e030f3bf9862104f81e03f8cbf8535
zad9823b696261b46e74c17a4d4b449a89b0f261da756228e45b5043d2dd058e1ca3bc4f307c944
z1e6a5cada50eb920033013c5514baed1d28d06a1681f139c3fd2e9333c80df9e40c9f08348e41f
zc6ed3931a08616a4393179b858cf78b7c5fe71cdba0122b491e7eb539cefc9e599bcb1f6f741d0
zdf50a38b8ecadf2c6cdc86a06138c378c1081eeb17ddbfcaace75e41f702b15aa366e25b3b66f1
z9e5c81ede1d2d42993e2649a8facee85577707eeebfcab7974aeb7ef699d3bf59106c241635bef
zd94a8526f0bc615ac5200cdd872d2c56a6887c33ec7febfa555dd4bc6dd3ce417109480c16936b
z76ba55ce3f0e1ecd488025e0ed3d7e00224059aec00a123db420eac015f9c5433a5ee6fe48ab82
zb1996b70abce032f38e12d9abacec299d3f3218fff48882084ec27ba967f637fc6613c783ff83a
z67d1b1514f62e9c7c5a25c0b20c1c7df6abbc7d922826a31494a93a418d4c490eec5b5dfe5b977
z05bcd61ca646ed80acd2161b45d98a05ba6c4746433fd265a4f1efe3c38a3b67e2ccc75016d902
zf72921926db971e8849e77eae448133a53d8d09a25b329ba56cd03dfe0ac949c28ec91a8953dff
zde0cf07a3136c82309d3acd1fc5aa39630c8b7d807e8387854772aeddde32ed0594c18aa0e14ef
z8d76a31b32bc71e0cfde593e0c1524ff679548b74f3deb5d6d124ae6e762b9794924481be08ba4
z02513df8fe8008b713efba3d7de46b084a289fd1b959e9af2cb6aecf7f22b74fe55960e4847b8b
zbfc5024c66ef5379d444eda09829086aefce88badaa9f3c1ca617b643049bdfdb90d7166d8627c
z3c5cf18fcd8d0258e5e4254191bc9a5eb0df39bdfd483615ac6014c7ec264829028487504db798
zc877185e11992b1f1aa511899350d390c818b5ef17cc099f2f7559c6ede16d62cc70cdfd9973cf
z6e36628c28a32169f9ab6132fe181ef9bc2ffd46a58e1898dbad0accd41f1d90d02ae947d22e9d
zb0a2cee4336ba825089f4787d42a7dd41272d22d9bd87e12831a9d734f134df21f9b6552daa1fb
z28e1f002bc829abfde7d650b6a7b4bdd5211a74a105b0c259710b3e802c60be0b2b21963179bd3
zb1fd5449753c57b993fcbe0cfd46a2c22ffc1591b9c4b0f9ee073fa885ded90e31eeda68c8aadd
z188f3f2d555f332173f2059f2054e588d28e3d55424e96271d62fb90087265021d6998c20716d7
z765211fb43950071c3107b64fd40569e23d774dbaaa118f6d2f3049dfc6c0de6b26e454428d3b5
z7075091931a87dba4d0ebb810f7dbd298b32b741e73687a87467a96caf5d58cd13c534b138619a
zc893a0a6fdfab3222e6170c2f9833de305f0b20dd7d69095b4506f57865c247bb09198230b5700
zbbd6afceecc68855c225db15f0cee7a5381d78e95b38d6f2dcff09e4041aeda827c44bdaf84333
z7f6e3ef0173ed8eca6c573d83219711d20dcd3b79aa6fa5cc2d35fdfe9cf8a2f74a106d1612c25
z131524c089e1360c9d79232d35f1cda25f7d578c170a9b86d089e88a54a2cf24a25a190d27c7b1
zec9313805fdc13af5fa30c480ea9fb5e239ccc2ba668791801d0ace5434d16a93a7505edb429b3
z0f6d3f919618397b4bf4a4c5aa5dd02b7a3dcf583319d12ade0aad3b3a104f27ba066bab9e7584
zec749d61c31b445fac6c81ac478cc510c2649d723d82877dfc174b9f6773721f51eba99955afbd
z17c8dde6b0e4ab0efec0df5de30b0f2f8938592cf3302ae1aa4ee3bc5f20f7a0a7d4e480a32b4e
z0cc1f1011c8ac74a42eba5385ca903e5ca6955976cc24893143c952fa352c43eb3056de355880d
z8d915d6f391f6169f1121373fdd9d6808fcccb19c6779a19b5877ed4211bcb990a4cc9ff6b6a81
zdcebc987978fbd839abbb87a7f0bdbdad5a17784199bb5ae022ddcaad77e50644bde470483aeb9
zcd64fa3df5f3c97132cb95cdba8577ca1b1f84eb302299875d5d11f1035bb7f22849d81465bc90
zb5cd037094ab50c2bfa056cf054ee7f528b70d60c6909c58d148ebffac2cacf817021fbd3389ff
z0bbf5bf47966a51d6603e6b2bc4f8a277d7528e08d4e5a85412cbf2be10c6d0cd18f6d166770da
z5eba2b914dd8ea4c97515d68147f98fabf95fecc83dac0fcf5fc9cd7b3c1696eb6444d98fe2bb8
zbbf28b6634f700d01dda6ae1c0320110f61f278aa2d40531b661e2edc5f0615e0c89a03b006e61
z79e0e51217fb0d7a5451e5aba0826baeb9e263337c27c1da28d9a0464f35064f4dc4aa2bbd4e3d
zc86ac6f26f781f0f8a73bf42441710b1818289c7ccb81c3e239eaabbb628875a951b19f6f728d5
ze05b317c3eb7796751511c58cc8ca6d27a6116bcdc2d5ab849db22c7fd9b710083979f82dbf580
z7a733a187b74795e249f5aa71b1f73e814b4af443a225a9a317c14de998e0235e2ebecadda5898
z20c0453e7d36221d226c542f2e91579100f269aada26464b23e9a64c1dd9bd7bf50c57bde9c94d
zafd6d9c7673960e5770f4cd6f48b4d4d02e1157c3b50959c9f5ade09a1bf3a03623431a4140fb4
z99b015557a95a07bd3e18dca43373bff68cf3144ccb8f02771e7ba96fbb916cf31e0ea4b220fb2
zf66b44bd432b54fb5e90f9f94e453690a50c7061faf239c59a76f6469dee5b10ad2fba77ae52ef
z98cd27a7ea4650b019975ea5320be794eee600c0778eadc88fcf042a984be1ce52b6c860d5a402
zd047841fe268226a5438eba8cf4fb54cf382cf8f12fa242a28304cf9baa837a64d910168c012d5
z92f8c298fe05b24ab04b92165e67638eb4cd2aaaffe7960c2099409442a5fbfb9fb9ce9fbab13b
z502fdda5d73dbf871b66d35422b75bff0f6c8f54efa35c73d730390a6c975378e37c17ee26a2bf
zcb3a05a805e5e69df7bb1efeb2bf15a61706177988ea2f585db369a8b04ee6b724bb6b5b807a1c
z4669a42f3fca5b91376852cfdfd9c650f1c6ea1607d7ae69a28e92aec495f9546e92e9afb96677
ze2f66dd6398c824f635bcf13187e25dfe67426c0daa657f775cd1bd716f7d0794b47c525b5ea32
z841529b633d9e44eb0b50865f2563da54121a11fcd16b87f6325afb5408d3711a2e48f8db2bd51
z2bc0d447d8a27d520522ec595cdaf9ba2e622244bec1bab13e5739e7a7d64ea6f8e371b03909b9
z96a154c8a86bd56768071ef72f65fed593e5744d28475f9e01f572b6d3ffeb669ec9460ac91aa0
z0fc2fa92861c18e246a3597a62c6fa710c8803ca08a8769720ae88625ca7717bf005e4062a8535
z6d765a69d4ab70583b40b886f5e827a12982353d6f230bb669c8cbd851974ab4707da90b98d2f7
z77c8fa4c608de29df564f3eb7852655a6b676d6b32ac03170fae2b1e4744fe79612a0f181cfcf3
zba4cee2fe9ecf01dedf23c76e9dd80bed7f2789621d2a1ca84a7e6a9b5ecdb0201347a6fa54f57
z5e4b01139667af605a37efe096e0a32e4fcfd565dc6ec093a9e3ccfd0fa2ad6af6949e82458f7f
z8f2d7622ca0f099496dba9d0eeb0fb998373aa559252e5ccc16261ffbbd65cbc0ffc391a189a30
z7bd2d26f100c15680e3eeb5bc2ca7f4db0ef5bc47277fb818adf187a08759727a27b0ef35fbc4f
za48f49eaf5321afd9b918d888f6e39f9a0efc59572ac0891f5dfda3703150bc0b6520099c14573
z3877b06144cb40ce86653a141882ea84de81edb5cb2541d70d7caeed2af9c7102d6e75709012c3
zc5b1a9d4f2b59c19390b3b6845d0713839069b6b98fde03207436058c3f9bd346fc6996937f127
z671391aeb99a48d94f48829549b89cf36315e6004da491ab1fe7bcf62dbf0e3c745a8517b5821a
z1d16e59763299d8d33b55357a2895442240f238f0d18481d57b683feaa4cb18586c175dd769882
z6092cadf088a6258f7f9e8b0b9db992597e08dff1fe54d7863224072a0593417fe22e34522aec9
zd8ea8443121c7ab3f810dd2e92472c80425b1de7f6760845381fd6affea25828bcfa18d0fb4ac4
zbcc7720477fbc552f30a0eff75f61e1e6deb71d63929cb80a5042c1b9e1a6c5497e3653261310f
z695f2f64c23331856b61a0d5c2b8087257c11d3eb5cd34c62ad8502a08052753df7cb7355ecb7b
zc8c52339b9448f26c5dcbd4e44c2d4bdaca3bcb82d6b2dbf0286362bb9fbd6a0b6264b037ed0d5
z89876b999c37609fa7cdfc2c0ff4de31de744a0a45fac569b6cee29572ecac4251d647fc6a9a9e
zcefeb3a947e6559860ffde0960f974f2e8f043db6ce3f03ca143b48e299b1e71c5451ee6fd0424
z3ddd199e6432346bca551dfe175127e8a4e82cc73675ba9200a38a0414588658ffef4e0f116a6a
zcb4787f0a00d785f198691ddcee8732254f276bc21bf90ae3839c24553ebc4e1a702f5dda39d0e
zcf67076ba69f350facefc7a702115341ddf7d49d9b84dcaa2707c9bf6c4c579f99659851d7b78f
z7d65c9a7e06aac2f3c32dc4d73398714282c83f267d45f73f8b934f357b49ab8c9056725e62757
z74c7de19498ecb0189a687eb31ca6cf542507265c3b88ecb9e2677a223453bfda430dd05539140
z6c5195a56736ea4b0c117d0ce4bc1ee1d917cd6348939c9edc8210dc157a87074a3ec1998dcc5d
ze15cfd5aa4090e41e258061a0c55d350e0434c2e90b63b09c2d3b861366c7df775db455ff50967
z2d6d4ce58b3ae2d717755641ef0b9d4b4cb1222f88484a19029d70a3f2fc06d0446f7c88085f22
z547476cc898cfc0b2df4bf0e113067ab00eab75023fdd00f0678f5fc3f6881445b91c56f33ea0b
z47b49971df87bb4562286811fcf10da428df9aaf9bbe914aa54cc1fb1e33425c89ef835490552d
z52ebcb58b9eb26f09f078e343bff3b46a0001d4001649bb4cf2d32020f125f78507142b38e8bd7
zec632a83818b085bf64c10b444af3cba18befdbc0c6e524d023f07a8fa8234b4bac31a1c33e602
z245ba663144a1251b99e3c38ddd54f394e0db7d646e13a3ef66c87eb5965f25cc6e91ac3f1ff44
z446c65b67a1183508b2bcaf026ab827960beaa40d8e7ba93cea7946ae754a9fa814e95f02c2938
z68640fe5927ec197133d103e5feadb2c5dbd998b6e9a3a4fb6881ff018e9e976a6271a3c5b4a0d
z03da97223ff1897da2249572f116aa396d33abde292392d8957cf05f4be088de50785d9ff45244
z63eca641c10455d3ab194cb61ff582fa0e54fa4824bc9fccc773b4d850a23c7c4b16b648769d9d
z25a3be6335f22ead28892087f766c05841541cfde1f03d80da82107d3567823c47dd8441d28d7b
ze63f40e35a758720976c51fb0ebc809cef2688d99b54f0fb64a9f5dff772ff726ee79621df813f
zb3a02c20dd0de56b1bb9c2e13cb750800dd7c36448ebf3d113cb68aa35d3bf7a356ab9ed470b8b
z7072d1028d75fc81e6c38135c86dbc5189ff9638714783ba78497b4530ff2fe50a495a30b2581d
zcf9d2d23591668d7605898c37af15367d3179863c6c669ff14cfc1cda191d9cbf73b3f8b427527
zef16fa57502391f098cd828de86711b82bbdd2e652f683153c564e9d67bd1ee6659d18f990308c
zce1b9e66c2db49e186f68d348cbecb6a204188b70a668fd31ca4ff9f1418e5e600fda357217acf
zf7db7d51fceed610953294d8e6fcfcc978544eb0bf12b9b024e111196cbe54e567c60eebd165dc
z7e7e753ddf68d2c71bc75cf8662dc0c3875ded1c7ee2bdc2e2f16ae0482089d03d78c1213c5922
zb2ab73fbf7125e219f3ca031b73aa47be467882f9358b807974e5a8ec1703deae99ec9a307e64b
z997939f3965f94ec4f2feb957ac8063bcc130198a2f1d122d131848aa062da3c7f613e772c0ef8
zf7d841a9358764344e9d2dcc782682c7743d5189a42cf8d57ae4f12007ae19c64015247a4c5084
z2282b60314ebaa4c9e0f04e2fc8ae5dc5f21c2325e36619eddb8ffb053ff23585934cce289dc53
z43fb2cffa26b33bc71d49678552f78852eb7193d16c8780af2b20f689d5fc0b520bc6dd0e6d762
z375dc6437880469e6e7bab2e21752c8f9b8727c5be5e48df5c819a1ca872fd20c8dd195e27bb40
zd86d2aa473443675345692ffba6419ce61c1380d04c27602aaf711edd642f30380fabeeb94b953
z31229b70ac2530c180b51cfc4fb6d3ca1247b15b542130145cac0de551591aae7efb49a47d3c25
z2d94a6b2bcea78d979d6143f2eb4438cc9a75bd8f302dceb3e7b1bddea577b13eb3f307629e79c
z2e05e552bae89d9c4159837f7024b3d03337362ccd8719805a418a8e1eb4261974af1ac876664b
z02aa8f969875ac18327ee85738b8480c2bf483a7b23509ababc3d86ef6ba927016ce05b1eb4007
z9f3126a26de5ec787e3f61373ca32f7753f81a992512d87901f62c968407da7896b7a0e5178e9f
zcdeb967ca37274f6868652f7763570ad186d43f933c27d2ff767788591ed6408d5ecaaaef7c959
z4a6cefec654346f3fae4ab5c82c8e8ebe0c3646fb2af6ae032cbd031ee738e16f707b74185b18a
zd162c96c8e7347fc7754941ba239f94bef5067070c0689daaaf6e488272b95b1426338a9ca98ec
zf678c141c0d5af0c38c697dbbee67e26e4220fdf8a5bf8c2b4ffe0b1670d8f0506d3c7ca79b631
zfe8ec6cf75dc2efc81495cffd1b3423113ac9703651e135df8b53571318bfb6a0b0f3d6a67df0e
z77612ea01f3654f32585bd3e46b99faae0d55a0a58de24ab19910304842ae80c27c5254e81e08f
zb422c1f0807a2ef8a7dd50c4f221827abd7bbfe3e145b119d0a452cb5a6e7528729410b43e0904
zd6205a27185f424650cf7005af496367d907020364b8a40f3116de7c9fe29b195de1637bc1cf97
zb68a09a1707a667f6b37b0327768e3a060bf903080351eff9d525178e4634367504c0dc2a632a2
z4a7c4db5b383774521dc47f7e180f6d05b998270dadce4ddcec707e514cc5422514299b2b243e8
zb42827ab71ea9af406124a3ccc0b0e34fa8a526e06c9bc889eb1d4c1ec14b2c9d1a89919775623
z3dd63cf675de974228e8466415f4a1bfb92d2168e3f0920a26f326a0a1ec3a507728e64c91ed50
z6fe4872048519d49d253a4adcbf632710f1ab8da140c3ed3b694536a2a98ad419ab4752ec53b40
zc7c56f703718eb2bb4027995a57a0e6f2bf4099204468a406a88c3737dcc2992b13f505a154c4f
zf7d321bb8162d3032b83e7ac766b2826b06a3015aa6bb13c6fa4e3c4934415cc514b6d5bb7cfb1
z3ac43d4a0aa6ad0b659a3a93d0185a2592333c0b77c1384d429966e13f8d5bd0c20a2654e87a17
z70252b65721b2335e2f9856ae97952e19cc436395684fb88a71181e3989ea035b4f7807b1d2859
zeb942af9da8e02c7d0781d142763982898423024104f296ab0c6bf35b5167245377c6c078c346b
zb4dd5a8d865796a93ecc37a58d49f90b035450182f91145e6697d4d049c63b747068b51e7c34aa
zb4acc3fe9342676d522f8f124db93d23fb4049190b1d63a23774e53c0378c5b145b6e636187071
z5721324bdd96f8738e93ecc5553e0bd0aec8a20c1079bb7864a6b86200be235cefd7a709222cf3
z23c0c0433de62d28750a76e5da3fefcdc6a32aac5557190a1293091d4f5d43c1523328a104fa60
zeb599686d489c4c1b6ffd88c9ab2dedc998552dd3254415c9f474d7a6282a0de73f50a49649293
z0e036037b2666e814a34205e0ea2df2fbbb3bc43075db838ea330dae7a912e4290dbb297ff77ac
z9f7fb3cf8c1f915127994b67fb5539a06c19c6444e6a0977648c7fa8710979bcfa599acb846ff4
z0edb525711405e4e22dd3561465e3567fa440519bc0ae9967620f9ac79b21a2e4171eb169750f8
z1902b460d17f523a39b22eea026e6310ccc347d0e8d56f04654171a65e2c2d10567d0a8800ad9d
z285f6be4e53ea3e2a6a4728f05a7d5acac8af7e2c4386a5b890bf0463d5c0a228b0f4c3c2fdd70
z8c5c3a89f9a9be6e52a178e264590784d8783fa7dd49bcd346b618a64bfdffac55bcba28ad1612
zbbce290631667aae569be24c383876653df23ed858f9c6bc561ccbbdfa4c530ae0a9c85f0729f1
z3820eec5a714e825a2f3b07c3a7aa6e3cba9332d38be08dc20ddcadffab9c2b742e94d58c3cdc8
zc8dc74e09e3449aa5642685949d5dbc4af9e955b157ab850cbe513fea4ad7a64b70ae39e410c4f
z6d90bb02982d401371cabcc8422fd6bf62aa4a9068c5b68e40baeb03166aa4a213a83696e4ea0d
ze43799a9008a21f34707053317694a36e7bf74bb88414bf6ce901a0c9d9df8d0b2b3556b60a590
zf298533f6d390f166782815e8af73e15018b94a85037caec8e4684e9f3b15fa6cbd72cfbdad1a4
z3428f7b6dfd68e5eb3973d5e980d9b1659fa4cefefaae5c5787919e4e88dcea940a3c5ba46d5df
z0e0c0a4bd5019add1b9c4865678da03182aba3075376e0d4c0cf8db4c447c01909bad2ba7981d7
z5e475d08732e18feecbda43256ebd29ae7423254326a8d17306beb19dd487ed25da301a2fde171
z6453bb2348b3df13537862ea9f22fd3fc496d2ad79ca759490ea18ad91bf82b6b110d7ff0c26d0
z4764e2945586d0403fd7949b61afca228c871496dd77982194ce1520739dd74821bce5b8d8f248
z320eec2294b1bcaf844c52e829b89d0caa1659496f471892f23aee406e4a29cff3d7f9d21104bd
z54187f5e1e81f8bd0d1a58c0ae4ad10c3970fe961e6bc72f5f4c6dccdc6c64ff5200783ba62c53
z72e2e324b52d561c0ccfe89a39d727368e399ec5480252b47dfd2d4531b84aa366f0c54cf427c9
ze2e836cb5f660cc113932fefaf030bb8893610cae9735dfff5c9216ab67a0ce9956b3fcdfb7172
zd1aea00afd35ae1ebb3336ade1cebb1d555ba29b978380c855750fd291e7a215a5d80b549e0378
zd84dc808e0852eb2ef8492b50d0ab96b83261f7a4cbd2703e1593790d003b30379ca04fe51def8
ze6fd869b510029b78ffbdae43b1d3a89a83280938bf23ac6a4ebb95f1f9e75c5328563802faddd
z7e9b744db37abd886a9b3ae293d2f4cfea643d308922ab3f39a3adb08d6fe84f0a698b8450e64d
z056baa80af715b8c9e016a0bb2c72b2025320a31de452b2a49ad92f5a15dd673d26ab6cfed1482
z32ba7384c9d0c982a894afd724286bdfd5d515eb33d178f9f4b4db33bafd69ae12ddad8bb4f1e4
z24a4155f3e97abee5d5b9e9c6b3f90b8a36c836528a8758d2b14583e60a34de1628e7ad69f4ad9
zcaadcccf06c12933ca5da0c0c83a499f1d947a528c7edb1883051d9d752afa1f0765bebd878088
z83cc7ffab40b0544a117d0f3ff0b8ff3a2a4d88d5819b55537309b3aea8233e01f7e20babf340f
zf379ce33be3cf61e54ba2785181aa8904c4789f77c4f017000c527b378f47914205f635fc94da7
zfed7fe57e36cfbaabbce80c69ca7e2283435d5700ee0b790b20b0ce1eced4c4d1b77ba9ae53d9d
zd4c08231b001c55a99f9825dbfb22e5c70eb168e3abbcde33cee0f83443325278d020274b2bf1f
z155a11c7b8e9e46d55110faad40f77d01301bac4836dda6a1aae5ed823247ec8568561e7a9f3e0
z0afc582f5f3a0b953a6d0d4b907d28664f8da09036e8542fa5e8008e0db519e30f3bc0175ddad8
z01790dcee560c233e6a492aec5b38ff1b029ea5b54202992226ed9f5de6813b8e2d5a44f676d5a
z1cb7b917c33a199178c0d2d57a72b1fe4b342c0198822f986206ed6d543dc0615f03db4be41d23
z1f3628172387d01db22035a8bcc2779cf2eff1fa05955ec1a5a2e2bee902e01b50d570b017d5f4
z7e03310b90acabd903aa92d9ec2bdfe91885843d1819a49329fbe43374275f6e04ecd4b59e2642
z073e6ddf12280f785c238433b158d64c645c91aec5d531f3472a024996c798c1cdfdc51d1319a9
z426f6bcc71e475448e52fd7163501e59214c358330a9014efcd27227d659e48454fcba238c61c6
z970ea0a4a7e15f4deaa416b63614ec2ea095fe0558153d618799f9b385f3bffad269191cb67471
zff232d038b24eb360792f62e2b6969c8f5d78116fad82b8a2f9582e83a665256d520b12db68479
zab791d9275c0b08849a4b5b74f420de310b66c6166fbd76b4cf318c9991c9034eb107daca46ed2
zfa86034a16eb75c33b1dc2df5ec4bbf77cc1cad3238358f1854295c4f998fb7509e7a3f41383fc
z7ab0501f9211142f978e9cfff35d4b665c8b95eefb16437047a3a73d72fe7d80446efc5bce9284
z13fbc39059c7057c883514272ac54fd8c40f25daeccd2f618199ed66dc7a9cc404c0841239227e
z21488921db07b26e254c905e2e6d45c4b06242402ac00f3d6f1d270a423df97c64253fbbfff698
z018f23381682727786ab8f4c1e19ce86e50cc10d57e884f47da2c6fde91d34e3ef8ac41439be94
z6b0e4fac66e0220597a68a3b58599abf4965aa0c0413cdccbd5cc6fcde475daf10ff1845c8e2b8
z62af69008267acc88b32c9ad8dc10ec22a0b313728364dbf77fcd92fac89ed49c52dcc8aa58c3a
zd4a67bc4ff0b02f34003ae43b706ea30a8924e3bcccaa21965404ce1c5c6d1d39c83bf987cd8da
z8bad4804e12bee387b2665ccf4bd4f7e89804f28cdb6ac25daf201292945e3d08d0e2a26ad8bce
z1a7712de43e3a2dc6227587e0c2b1eaaabb06651b995ab967df89ac9cc17a6f6681aa35d5b4833
z9c342c823edc3a1e1fdca2ebb931a50b1b7c66b3ef0b75e0b847b1c359b077fd50e2cfcfaba649
z7271e25d3d11cfe38b5c8c706243654a798b7ea5c1a52d84f94eb42f1ab0e693765e1359d0fe82
z3555c9197b6149d241a523c9917d8f1928d4a44e6d39d8bcf8e981c6e3ec8d34dadfe01ab5d45a
z11ac16184472bc7a1383c6ee512a2c2029835c57d8a918a019988abc0f6cff779dbc0e1952ede6
z62789bed2a4f53e46fc458656d29e0f05803ffe17d88b5845515b1f7026784f48bb446dfccf98c
z78a56dafa06056e5a9e9386d9f4e9beea911a5f1e5c6888053e8f2f3df6221522c8935369d44cf
z07b0e4b46273fbedd085c5e7fbfcf8f0ecb25f23db5c8d42439962d3484447549b7017315215bb
zd026348ae642cfa29827a0f7324149c3fffc402d7b78fce786f600a3b1fed5bfdb206c8f4da0cf
z0d5d96ca22a111b22c79896f447996e5a1c139aa29417eb0061fca311ea807b931770ac97b4937
z3c7a27b5c7ecbca4f8d3af60055534e00fbc06c899b94b7d47849a1e91f651df7847eb1bf57170
zc48d8e511d5657d0db4900611aa571121cf0c7f0e485e66cabe778fab0e56b11504992a12066ba
z987d695d778a00c1ee3ec387fe5841d3e46b57ff03b65c4453c87542522d9915c786b67d81cafc
zacb773dfefceec269feeae29d0020211ef72d793421af193511ab8ed8130240f1f295a7db2c29c
z1dcd0d5c47b63341ba2e53bb4af16dc76f2c7d90e16090130ad30a1f8d32e36633d5a4d4142b64
zc661af04a041915117c499ce9e261c7b9354598999b3ba8a1b15f457445202113271e9e8312565
z4560b736ba3e5108ab5a1c3b6837c41581ac84c7b6e5ed7abacba46c23a1f9d24327685199bfe8
z9a1b744c9f9e44b198c1ae11078d033b294e8eaa53d925912f8dd240b7ff36f3d0d644c143d587
z851f29305d49a75f0d59a79438318942a5debbc0b35bce125262cfbe952a935437390876647f88
z2da07de55a6e9ac9a9fecff6cc77c71a9dff1deb692ea0f3929e5d139d82e7bf92b965bafa951b
z0cf471ae2101090721f4e891e2c419642b6a7aafed0f3537b543beea9ee73f1cb3aadcea0d2dfc
z5204b23a6b466ea5fc98f2cc4e5664846ebf9ba7ce31286df21e17095cf83015b2b24d82496130
zd3e29113b70328b17a665992d9d1120417f9dbf3d3abd554627c31335a6b3ecac0e8a6c7fa54cf
zdc9f805234e9400f73d1a3addd70a7f436d39aaeedb2ca4eb6026f97159c4ebc6d725db7bd54e7
z99deb11fc0a3ca7002da607293687242df70d0f11669073d68024f2d6f62a6c36c9b7307a17486
z2b9190434766bda6c51e57554da63e638089114c28702d40e059ef908275139b66d9f73361909b
zbefc74fd3cad066223b614d157e1d6be2179d652b04713c606a6c718d0d6b23bc79954f3da1033
z5a6260e8f6806bd1d5f3a1aa4289874d10fa29066ad3617d783a0e6fec196af33e5a30b2c4d12e
za5d69c9f8d1a5520dad4e4e4fd4072f469c4ca5d8afa0e44903cd05bb7d3b310babda6df7ba625
z0dc17e4d9ed71f605e2ffc8eab229c11c46ebd26f3f6b4cac2b47724facf8d23c927b11efec571
zf836905f545998a7dd67afc9c83c3bc8dd3f5b46e9436b6c770ba2f0ea88cd7b3069e09ba8b708
zb03a45e053aef512d7096e674ef82d70b932ea91442152988bdef088525248e8dfc52d08360eb0
z749bd7b4428b4df45b98b088e0472c334590cbdf0573b52365abd99fda69b0fe10da159c3edfa2
z99d223c15935e57853c010dfc964fc01fd3fbb9378b0543a60d2690da24e8b2024a0de63fb3fa0
z5e261f33e2e18a39b62fb2606a4f83babf7a566d3b4cb1b49495650e40ea4a009ba89c4a812843
zea7f54ea77188af9c99a6326f5f60e4f8d26cc40da761485f54139538ffb061fd3cde7542337a1
zc24a58100b7b0c0b9eebae7bbedc5316bfe26a2ac57afaefdcb8f754d9dd035736141ff3ba17cb
zc2c02d79008ca391eccf2ee467df9c70e0c5a5f31beb50f6d42be5256a44cdf358170464cb8786
z042f67f83efe9890cc1d07c0678c8d921c67df7d41dc45a47e28a9db91a39363f0717ad52be98e
zfcb8bda1b22c4a4bcb52b6fd6bf613602a1b316e3cce8c6a17ad2b1cdb4033796509e1fc6b165d
zbc48fa1239b959f690433614b4e75f832be8819aa01fa52b1c0d44f4d42c70080b85dfa22116de
zc84c19dc18dad842b16c0e49da4d71991384e1ceb32b1a75db7876424368a6dffb826d31ca3543
z497918c0f4989d4d39817436c910cf7747a5bd288bb6842ec319f7f7d3804d8ada6e7da8189413
z13d6f3470f303512e79815d190aacae2fae4e1249782a6774ef17bf42bc085c207d7e3c915977b
zab80737e80895202c072177167f71d40a514881fa01981b0707a5fbce72444c5b060bdf485d1de
zf50227648289313f5512e3584da0ef6f509528dcf88d6e3d1ec64eb1b8819e5838fda797a2836c
z8ff5f90825a21e075e724d3640bd95dc3d732eb979ca56fb823bbd0bea1cd3dd464c2b0debe108
zff6fe18c8702739ac07555c8007260dfc208498339786d685c06deef48255436f1171106ec056c
z6ed3f977528e97e0eafc54c5d603ec1e66b29705e3d666979d9d50c12aa3d709f8edff9c0a7a06
z2e44cc10ba6a2142ed94e23b40df1dfb4c8f72d5706a906378f228fd4fd6ce060d330da98efe3a
z1fdf2b3f999e3df8056c746797be7f880c7da8639fd540d2e4b242e6bf587c2b29895f541e3b80
z9c1be06a4832bb29ae3ebc4a756dc3302ad82f85e4ab4d7fa369b0842e1ed38315cc44f85960c6
z2119c5c43abbc9fe69807fd41415e339609151b1d619c5c97b571f178422a3b94036366b32a2c5
zaccaa57c503b9f96665affdbf21caebb6dbde5df473457d3665c49750491d6b2cd240d006671b2
z0bb7158cfcbb4b35443bd837eedaf89084d2b9f663cca10187c0da8deb3700062ba7f99edbca76
zc6ff7f18fc5720eca9cc88295fe9f034127f13efd9b01b1db535bb17459dfdbf51106771e4bbfc
zff8ff5a32a510c003a090c8e93740ec3b55c9d5af4fb4e1ac2d5ec37caf196b31fd32842e6d52b
zc0231c8bcc5c7e7448a820a3d1d7b926c391ee265fed43ac9b06c880c8ef963480d1636ccb634c
z6a1bfe56c67ac2f695a2db458a4b2699f92782c46010a208fdd552368cec7b9d3dc9dead5e86e4
z730352f82c10ea445c86a21389b6098ff813b6dbd25e0c4479ff91bb606c861ad2ac96e2aced1a
z7b7d9939202ab6f07a1598e6ea77162b20c3b981f941587c414f1bbc2967cd84288c5dc68969f5
zac720495c5d3116ed16fc71190c7ef92549bc33f540d8b07701412c7f1129b33832bb6ccd9f03f
zc26ec07326b115d0e0acb640655b95b248300cbd4751d5a9b4e4a34e583fbefe79914a8bdab2af
z675b20d2634674085c37a898b9998d1ae48ca64cadf104d701db827810e0cdff641f9718895a55
z5ae786bf42ba18992d5fcf47d25011ac707e15d1f493f8e133298a5626ec7fc02950d95ac48f1c
z12852fef33497bfdf9ce56bfbac9d38b6b9a62be51a41094567d936f9b62426bae2c6275c47f3a
zc273fa17d980215e87b1974b24ec2832407e9aed4efe53bf890d85cf682ff564f5d7785aa2ea9e
zf435f4c738def3dc64c3de18be05990f826d4c6defa2e2e72f89fae3a9166e6a8ca0934ce9e077
zc1efa99859c07f3d3f97d4d5b71a120b9f63b5905ef40d0b9fbe2638ce607b82a1df305e4d6f07
zb189363b4c0bfb126f7331718e3d0e95326e14d29a3f58ff6dc1a163655244d6a95a2280ff3a4a
z65268c18758fca050517f64a0c361cf0fd87507a43e528578ef60d1e665fd7c35b80089da26dda
z995f0a5f90a3735a6df9e8d7d4e923a87a37e05a452b2b65c38fee85dc3904a5627b5a512c3a24
z35183158760b79129c67789f288c4b399ea904087b23fd60d6c803ec6a6d511b7b24d6c24fac4b
z586d12baa648621e3de9724fb6860a48b22b56b817a9fcc7479b25c98387c7ac73d6259baa5eae
zb46c0d9bb599fc78242186c7817c75158a5338449755eedc3aab275e3958ba83eb86b4402e21cf
z64047737168e4fe67f0fea4eb5cedd9b3c58a68ce28c5a0fce3f81e80567e491228bc8828c0991
zc11ed9a9f58d17035e1d8d9a5099cf700ec7985c3a1e11606ab75cc0e7ebcca3e3deb5fdaa7aca
z18b4aa11c4e24ee019abe19beb86fefb078eb53ac309f2f24ee0d88464c1e5640ed508229a61ee
z4d2ae9f311b98a4f0d9d68b142ae7ec783a4ab548dc125b893ed5ce10e59408ac3f5d4213b03b6
z1366410b2364e111f4d1f15cceac05037bb9f12fb29d8313dd4bc168261cf5c3b8c4b78556f12d
z4b8864a16cfab69a90d1039ebcb7edbe236c05bd8186d52197c7ebb4fdae912f3de3c0f68d0bb0
z4071d93f991c2cca777e38ec97e7fefadffb443b8a7caa6324b78f69d2cb9f9def77a642d9a34c
zf57ab19fef19d114c5be84fc47b01f62d28411efe1ffc290a9615ffd5ec8ebabd60a1bb4505c08
z441511a0d884fc85177ad8fa78588a6136bd4bbab8d57553878b748ac4428004856acdf55ccfb2
z26ba73cf75d447c7014421f0b4dbf22b3747c5cc72672a40b08c09f30cc1078236755dcb1660f3
z238c324963251e835e710043b771ce1b50ffc800ca1320f589db1c53ddd0a6604c2a9beab17a68
zd06283e684f4fbdebf74d1bf299380a501460312d8b1323b2a509cc8aebea0e4e045764552e10e
z3728c56f2aadbe71864f846026efeb387a205c465b787c7886a0a9ea6acd6d38342274e6a36c48
zb7dd174abfaf138c1bc8823077740ab74cef5ac9e6b92e8903d211f227b07f3dd27c729e4dc7ef
z3ba614851ce88d48ff4599dec136f4b5521e68e2dfc4496d32091a6d80fb1fe89d95ab8828e473
z9234d21d8170119f5bd79242b9faa79f5248b3d09a1d46bccc1569fcec1fa1891897db37568d7b
zb8c7ce943b806aaf97c0dcffc835bf49ea77a878ec63b6b3cc6fa0a63a476d653adc84ad0b514f
z32942e2c85df01fd364b49ab63347e5ce6e91639f8f0dd775db99bbdfe398b8fa42531ca7944b0
zda2219206ee5691b57941a25852f188d44b97b6d4981f3a3f8dac33431bfa41d892feff6597d12
zee574127116e8acdcaf852947fd38580424ed4913b0a5e2cc226c6d1eeb530212e082f36269524
z401111a0427a7083c0b1bdbf12e619d9cef99554ad5d3b99318b0dc5322479acedba997c11d78c
zcf201c75998f209389ee1e11bc5ba7eb040f0a1980c4c6618beb027c443629f63c707a583ae902
z2a92ce89597caf851d7a8c4920505900669676a9388064483838f7a7f65b8e6df50f28973a6c4e
z70b60baacd364811616c1506108b5053dff11be30c2b1c742cfec0f15f64b9ad90b338c6c8afa1
zfb89f5a0b2f9f3527fdcc9af4b4a9340990471ec354aab2b099fabfef60861b95caade713c5fe4
zb490fcf67c9b96721619336ebd8c4485a645908fc228b94e596ef6572a2af35e7b0fba0c205cf6
zb2f387c54fd6ce5c0997f8e69cdd9c683f6066211b082868be6c0b90fb67876204e1488a7dc8be
z53e9ac860e52bbf4b1dd2b42889c4196490c235534b30118c8343283f6ca27713916e50a53be43
z75b52de250529ae8258d06dd99c6a162049801b3a46b3e86fa2a961a29b05e28db2b7ede92b0e3
z7f044de23793d5bdb035db7055f133990ecf4332d35b2b9e4b77c18e132b4a67f8abcce381a81b
z67223632b265a42530494c347c045ab256e1d606993fb7a9e952d2743134b3a4ee30770970dd0a
z436e57246e2f89a34d10cfe83e194c115a650643ac9356639c6468978fcd7e30d823ff37e316cb
z630eabade48857b176169f5a322940ed10f519d55685d462600b9eef9865e8262917c0f121ad5c
zdd1018a256e21cbd6e5c44ced0697b3108739a010d3878118371909db4b59ae9eacd6df1e59743
z7efc2a402bebfc201a23b0e0ab5c1db0729428b30b438b41ec971da0457646f925eed70a24c09d
zdccf2c60039321ef0a522a40cf030a2f00135e289c1f0232060f98d274f65f9d9be12a422ed8ae
z69c0c545866e46395e615b9c2e2fbfb72c403a999785a45231932c26b61f6d3779381491d7cb28
z9a7197c0b14927be165ce256ab147d9acd5e18017da3d00c1fa9a4d3fb1de52b5d784fe2f57bc4
z9f3d795924dce3a7509e6fce7c1f470329e681916f5330067687fd8e1ed2fe11fb1a3cf5a67e00
zd0c463e8bc48fe6cde839cbdc10f138c5cc08568fa9320cd71f27a1573c0a9384690ab73f44fbb
z0d50f12dde714219443d21b73ddf626a83ed2420a1d885b70228b60d32a4cb6fdb3dff157f2e9b
zb99ab47993b303507577d9a2444b8c8e7fc4bb34a0020d110d3baa75f24c84778580ca8a801358
z50842b421d88a3a510cfa447e8c55df5cb75386d30bf17fe0769170718b4974b61f91747048dda
zc07473f1c544f65d6d3a50fd9973ea6547d0254e59d45d0f4eecb85af52e5fba42c5e85b47b2e8
z690b1ca3b0a296c5c19e286598bd0936ca1b1fd7918facb0547d8954903a319d5159ff3cd783a9
zc2c09ca93a9d0d567db71a1ac4c55ccb575b1acc7aed4576d7c2fa175bf94fb334f63d28898d36
zad9507d6137d62818d37f2057377229258d16a1a57bf5af610db910a6264f84907c5815020bfd2
zdf2bdf1f5dbd7934f9f09063bd694b811ea55b43d85d9b608edbec48c709c83a40390ca2aace09
z041b3ca4ec3abbc73394ee29f0effc881c578f2f5e4a6357d0fff0b005403179aa5e5c8086d649
zfac887e3816b406234c8fe7758cac09d8a44a98ee204f83d55cb23c047cb0a398ff28cd6b1f8f1
z67658a6403426a61e2f13c645d7a0390cbcfbc921da96610f56447f76989bf9f23e8b527e3181e
z5ad9166c369cd8fbc440d1c4be0bd0dbbacb7602606f83f83d29e140f329f5da25c0eb91ffc2cc
ze59bf0b5567402a999b1bf9068d3569ab976a5df01f1c74560c5ba067e3f2c367285adbf2f27b0
z977af8e2f0fcea5d04d1bb9bd916426dace3ac7663f5fed42445751b8ed3616586f34c1a9dc84e
z936c74300d6e46a3fceaa6a6f5a066ead1879e2c917ef87865cee680518fec44ea6f693c5d3213
zbfe2cc666b5698df7b0fad4275d00b9156fbbd005896461c6c02ea0303b7378c9addcf23367378
zd7cc50eca39d417e78aeddcca46bef49938407855a57a27a0a37d6a33b1bc4cb846ce133292b29
zd90a87777c958ada9d9979d323b7f257d7eed6a1920face2dbfcd1a0c4ab3d52dbdb276a325401
z486c773607ccc2f0b1aa0184ce203ca0fe441a19bdf8ebf90d6880b1392e70ef7f6a329cd6fd3f
z2d06508b1bf908e84efe139a7cac749b84d1db5dab18969a1cf653d4f299103782f0cac0d52c0f
z7e3f824c7e19971d8003424c4f73784c82493af016f4da4847d6c593d3dbbe2df7b248f46a24a1
zb8831abec9eacc749feb19cfbf583398a2e0788b8a575f93a0522010e8f7cb084cbbdf7a8be047
z7b3e3deabc0ac314096f0b4d14cbab3dfa82fc26c08d3a990f2a08e85d3cf44625e9e34184e66f
z934195347dfbf22a48173f7de12e4c670a38d4f1b3c8862a7961a73dc21598fe5897fc2194712a
z58486b0d78c90a9a672ddc3db28e1774eb44eac69f43a5bc719ec24e8a1160dcc6c820e3d08fd3
zdaf44e2fb0e972980d7016e64f794e697ecb855b05a950693bcb077671b1d00f1bd1f55a010b01
z60b3d4184264d372b04c6c0c3186b2c571f9156eb87f69f19e2076d84225c9b45a0599da19aabc
zbc3b99de55900fc69fbe3d9f38f2d11c0b6d7a4a59781a536049fdf15151a02e2de01169ca165c
z78911d0f65087c317d69a6f7270f40d8aa302a10209f7f4b613218dbdefefb2c2486c4ae8e07cf
z3f2c618f5f636ddb7c2d55638488354ee4711af989735a09966b8240e7a68808b42124bd5d8b5d
zcaf266c02df6fb6ecccd244e83cb82b23ef2cea20fae569c5a8ec099cab3e48ae3ea977748fffa
z92eec85f9291dd9e4895f6ce06e27c9d6b08f0aa89f0e2db091caa1eefc7e1eaa82855fbc8de03
zdb33a3a09a19ce5e2352a2f45e2d2318b359f645abec4f7aef296883add001dc0cffaa1a522d09
za5e9116c93980175dbb560dfe077ab0783668f4c39964d177ef86ddcc39759cb7cd3d96800a17b
z06da99d0ba14de718c7f8417920c3758e463e3eee071e50d9fb7df65567365ddffd55c70aa5e9f
za5a77ee9a37ca23d1e36ce75240a3352579384e26fda049942d8b44daa7315d4e635b2bf33763a
z1111d15338af054dac9234162c3a03ad30442c78b71de854b8df9369b44338aa99aa8f7f9f645c
zb95bfbd4b55228baa8e6f60b1d867d8a8bae288ab32517b9fba2f95acc62caa5434e3dd10ef520
z88e71763725d82043693a00b71ee456bb847ea87b036f298bef05a51ba4130c707553038d82305
zcee0b5ad8ab51881bc04e81014756ac5b70b3836286e8054aec1f04f3ecacf09dba41442d7393c
zd37c788bfc06943989e051e90f8773da53fe528ab8c80952c6bb38df63039eb34f285061e684a7
z76aab9b0c1cc2b799872e65f27ae27f8ea19f887ec7dacf2220c417a02fd5e312c96461121fe12
z520235db231a59fb5b8cd3294fe0ebdae614027b283339d6d828ef2fa751ceb4b6028c537de3f1
zcedb7f3a80d9291eea59fd9d36246c959adc96ffe71dc27685ed0ca2975a49673ccb6bb14e67fa
z588425f2100f3726cfeba7680a48cfa08a24b4ab67c157543619479ba3821dc8510c7f239ab254
zef732548d3d96c7bb4550321a8042524c0e13f53f33dce7483971766a05cb5b3913c98efe4ccfb
zaf19a672652c156c20b929be2fa246bf1c296ce45a2aa62ef4f95d64ec7088b6d9c197b5ffdd9c
z8db3adc20db3c107cd4e0ef7af9f4a8f145cb4e87bc7107a787368eb86f61ec5ce91a6b42dfd58
z309cb203ad4a3f17f7241f68129e0aa83edefdc738a21288db66773481ce6e59946ba6b18526ad
zf9d4d5cf9a9c70c30ba2b708ba2165816469668ed25b365fafc4e61ed5d6ae704b3d1830fd8bdb
z60f761f9b2aababe378656f27ab29d4af3ca6b765c7bcf39bd7ec82547f4289d29d7011c37407b
za03503b7da3631760e468df7fd45738908882b9aef43b33a8be5bfbc6b35215427bb4781da7bc3
z56aec9b76582d6e757a7fe5df8404582118e094bac041ade9917efa036aa6060edf95f9ee9abd9
z66a9c76fa01e157da257774762a651dba14974f4c2b7e6b38a81989bf7af05660d091641865a81
z4a10f39560fcf13b9310fdae05b5aefa9ce856e5abd1a464b6e4fca8c65257aa07b94ce0055c62
zd77a8252420f42306cbfe4d211197cd630063df54650693109ceadb214b5420d0a2684067ae305
z732eb5ea2221e0baddaf65fad8eea2f1eae1fa020efc31f2533c3fd4840cd35906f72b7f0e5a63
z94b06df70618eee3bd5348917371b935ce7314bd3271b7cd70ced1ae3c7c1e702658204cd45673
zeefee58b96d9972db5416c1ae34a66b4803a640791ab3cb2380c073ca8e1ef274e1ec9c9457cbd
z28337708a38a1987890511569e73ea18608c9600fe850ab39852f4ddefc350044f59f42a7b000a
zd0d59fdae9d33f4c0663ec928df7e8fc997e6f3958818250c111dc70e412918367b0ffe7389d38
z98c2b2f21e118829bcc77b900d8db549fa93b266994e692094b1041bae0309630f25620c5e6c18
z70412184fcff39c6462e47b6e1f1c0455ed74b875dec24bf27e50b853696f63c38b28c498519a4
z72e37f4ea7b79da45657367bf8f1602c234ab7bf04e24c8eff6ce2cedb9a5cec60bdfb49f9dfa9
z9f499fbebd3e4ff4125357a91579039810dfe1ca4591f64a0c27f0b1a47af9b8bbce3fbe74bf3a
z6abfdba35f02442c0369af21ac771e870a540542864f8f5f05d1434e709b8584506b2af1b75d03
z35a4a26f36ace2eb251f1cf3d6b7b7f048a515a2291256b0d1f98717d35d009564d6a05d7af500
z1495e78d0de009808c6f353fd0a3f3cfa1cc39fb9310c5d78decd8ce39421883419c96d5699061
z992f92e07fd7ffcef74576f8c1801f664e5c8f2e7e6bf485f16d86424120e43059b9988935f24e
z8c9f3add86be920b37a2c33f9ae44fa4b31798626d54132489b220013e92bf2fd9fb0d19b33bd6
z029d6612fadf7fea4ab8678eac368bf4909dc45736dba1c2947b825b25d5cf63e21a62502c14a4
z67b87e5dea4033a30745503e1a5e0bcbb25a887866fb3af018fae6f88462c9aae2908602112807
z34a0282684d37defeb985f03bc5d68a253c9cb68b6d640a8b2782d2fe046a818b776aab5b016e3
z461a6f3cdebd18a44a5f32e3c96b8e62e413bb6431178314361a36676b683b11acf448ed86918d
z2831f540ab0f2720857be138872d5efa74239a790d0dbf471bddd6104290cf9906d279ac1467c7
z3b39742ce5276496c7450d85a54da3d5020ff0a5bc8dec63bea46ba98618ce9a254a1b239d5282
z27916cade7bc44899636a2d8b0a46dac793c9a0bb6a0cda7e9beac12a2579efd9cfe711f342678
z13d63d89981e631a3a5c154ab6ca2410c057220257c140a98f14a1fa70101ecbcd69e71c01bd48
zae0921c39f1640f0b8a625b45793c4210c64039bff3d8755b0e1a367e12340b2a88372acbbd9a6
ze55b8c57e03208e881147079614ec19a0973c54a3b153f2c1bda87bec2669313e158a0329949c4
zf8878f6b430ae88e95cef4584b62fd5e6ebc19de3a89ac9519f37e9d7aa1a972ece2ee31a0ab29
z2f91b1bc223c0dcacdfe526e4591879779193c04bf184f73ecb59d1ee5e5be5f261377e8249dfe
z36bbec37f240287972e1b0e82f5b90c07532637e5d1d52e7ec2ab69997445a7d34811a3cd1b8aa
z089165f2f6c0eb162b9cc11ffcbd3ebced73e7759ceb82ade93040f8f9caece0ef303b04141c0a
zd124dca96e939931e0ed979d81134a675842e6e0a72b91524dfdde24d247ef59ee35df6751ed1f
zce863fd03467f21811c275d4b3ae179879a94202156103ab4ddc65ea41e6ca735396885b1db251
z287c21fefc81042c878f0356f7b199c30ae48c060ba59ae65c534f6bd15895fcc688de2b23e1ec
z1c79b310e4eefa1969706e9a337f0ea3e9f4154628b946f707cd03e74c5d8c48bcc15d06e52122
z6e187b2b5954995206ef3288b5eb73d0f32caf22fd47becb02839cc85d7bcf2cfc540b823e775a
z452a7758f76fa327382282c89006586ad476cd44c6b673d5065d021a83816d21fc8458ea7f983b
z3f5b95ec58c672fb94463b9d3d3672fd7892de15a094e6a9ba9693aa58c50100bb1bacca8296d6
z8308687b9ac431f10e036246d39d0c5849be6776a63940e8766052b9ada3bd8a7f3646f214d51f
z8e1348712518e3afe92be50ab80085de8e8d507f469ebab3e4dada03c1fdc3fb47e06f26290787
z19dc612af506ac6431da80bb990787f716e454d7c681e9ab09be3394b56a7ed8ed2b59ec80f446
zbc10387763ca095f1f4d3522db2f671966a02a1cf4896d0281fd561b85d64e1a609e062826b799
z11509cbf560f2749376b1c7a3719c08db8e28ae577e02d96386d840f30085818a560f053d10cd0
z6f2091d7b83326c632039b84be1fe8d6adad54265dae7de933b36e01ad53bc66f1cb4049650e11
z57252a800f96946ddb1d7296c57f7edc4bb31afd2fbc149fae8e60c2af9c1c1ab769ff975f0097
z08fa373aa02033f1853618596044f065b2a224c8921217a74d0fdf4778c91a308112e737b0b509
z68e89b087a0730c03a41354c10b93ad44c3c2abd8d0613fddb2d8a0017cad539b471c8ff5cbbac
z778af58691053e3b5927421b95b257baa48c2d16fc1b2f438cae3663a685f188e3bdeda8848935
za9fc729e0214c2f3cddabddc18e309592ea1d644bd8621a61f0b487ff929de0b588480b71cffc9
z2197887d4e7c9571bdbfce3b49e5a268bc4ef72f28041919e9671d637af9c22eb2357d813d0c76
zc2d0fdd086e2cf3b6d7bf2ffbdb828898034e75d761a92d7ae8480665e098cc2389b22bc517c73
z832ac0a624d12acf6dcdb7a1167a2f43aca8e69d0ee6612be65d4f83e6ca442aec97ac764a9197
z24a4c2d13f241bdb692d4d36c35aa234f59c2a1cd6bdc03e65214de9a3f202eb85444039385847
z9cd432c0f149d419abe32a3b13d519e0187a09b9c6af0dcb41e8b9010d3ae2898964c073495e84
z09513b7fc8205c11b2b363aee8a7205d030d6eee0c023ca365e63b047b0df9a751fbd4d1a12b5b
z57ce79c80067513af6a3c444b35e57618e752325068c69f9ad5685b6c942a4c024672af47ae600
z1d10b3d1a17266efa970473ed90b2f304bf64da5533259125b14c6eac155d687f82a34428b347c
zfce7585b846ceab8a6a3a8e33b4d8170afa2a758b5539b236cc66d812d2561c99555024a031801
zee5352792874a180a74a80888e3bc4bf1897282e003719de549a03d143e4b35203f60286e699c0
z09ee9fbd3258cd5ff6550cac9bf807365458e4e87e8ee50207fbeaea75c81bd3597e244ecea3d0
zbe04610c1b9d317ed30829f005f8c14bec9b6abded5d093d71a1b3a129dba39ad61e841eeebff6
z6fca1b3c9864d082896a7541252c73a82319a7546eb18f6aedac7b62cd5c76a7d00e34d8d30553
zfdd6f716e78f0d3e19804bbaa6c1cfbfca0226b305717211e6fc56b00eea4ca354a8308378db18
zaa56a7bd6b733b5bfa3d09115a854e5e59a38dd4807289063aeb221d3d0783e3d528d119e3571c
z311c848df4d5a64735719898e252e759b3b25d9e68159f171c81bf98d17d40b38350f8da5e69d8
zdcec503fd3158055834a1727df61d21b09797166c1267236023a287c8cad3b5d183b98aaf0e19b
z00c3a6b2ca8a213eafbe54c988aa52b547a77ba3e89dffeb4eaae1ac051b172546955a6de2b3d4
z9610e935dd377521333a941e87a4d824f3d47bf0af9db427859cb5876c5be78916394f17011760
z467345777efcdcb30fae4538a88b9f76bf934bd016b3c2e2b462e1ebc7f4deed3a0fef4e9d1dfc
z9c185a7253dde6b70940dfbce7de8880c8ae0298dd0cdc6a2a018063a619a325e9856c7a81eee1
z79c88502b7f273b7000c37723957f396582981038c8b0a9fef42dd9d5e5f4ed6c1046edd59acdd
zd6928812dea1a9381a666b7f084b790b0eca5323a807655526d467f18452066a6fab1881db241c
z7f21ff547e44755758bc8e5d9d8e1f016d37d012e8d6bc72776d2b4a01d0487f7c98abbae301aa
z1dafbcedd6b6d97953871070acd137de7cf0ee76a1e7e90d91d4da7f92ec4ddb89a971473a4caa
z40e2361fa191dcffa44d49beff8ef6421f0ac4ae10d1ee5b156d718cfd0a546b61a1b8773a468c
za5178e69f02623e2c8f340cb488a7aebbb201199661081eccdcfedd16a023db0ba82fb1f0aa42a
z977f2f22f806e3e2362af0448678056514024e7f0926f4c953d506b0c71464d5d1e84fbfe9aa1c
z31afff04fcacb2c63e9bbf370431ddc4113f1bb44c388407a14f9a0a5823842976758fdc41fa4b
zc2e5977e22517247ac8929ba5ccd73ccc4f8ed545895f6942c57a3d89bf891e82925c522b5ce0a
zfa06268c95c8dd5c66476017af0f21d95bf135386ff0c96c7feef6e9536a19588f3f750c622939
zc51f8f4a9f34c0d719759f8138168b2a1237ed13d51ed888a3d506c45d4d159e257f8758d0254a
z17248027a095bb10726af830fdd9ab51b38fc91ebb865380e6b653cd48399384f23d6f18b49bba
zde3d1722351edbf2379330ee290ce33772132a609a0b185a192d26c26af8cf3ce6c1288d77f208
zfe12e6bc6f3272056a671f25f0f434620478d55ea28d0616ba900a4ed177ec532e4454b57258b7
zfeb0cd4b7a48816b7798bc50e53b440d0bdec67125ff8e1851fc4b5e94f8e7d33ab4d7da8d1798
z5090a888fc440fc7dca2f9b85d2d926b66e6f5d3dfbca4d32807fcc9b35d7b3373f2d2a04d6840
z34ef941a6b8d4075d552ae188d519dba27c567e8d1fa1fbefc1e26075adddf189f194f8c7bb6fd
z75df0ea0f6e8b16099b6b7b8112e2eb9f16befcf3176f0dfd3d05b446099a3cb0bcb6d61469fff
z303fff33241142ef05d7d384b077ab458d8519413c8ecd0bfba7cc55a4a2a4a9de0a9e00a0f938
z24236a692774eb0c546e71a7640a88dbabb2e598a11b7c76e5231254bbb19a73b9e37e9ffc2af3
z198075f4fbf051324aa744b7af252c81c91876be03a3777710198903f651041e488f67d154e956
zecf7e92459fc037be9c83df0b671a149499e6af9e915916fedf835f547686caa29af2d4b5ff50e
z367e36a7f3aaa3f2f22a2c16d4c5c6adf81852f66cfd08c0e8afbfa662984181a32d22ea77ab9c
z7ea470f42b782dff9a21e1979950c16cfd5854ceb9730cfa589fad18cb7445027b95c69fb6b655
z9ca9bdf3d4585f8db14fd68978d639a439e48565d77b3894b031387e34caf17e2806ffaf246167
z25e1860b58d2cd6621eae284e4a1072f399148e910ec8a6f71aba8dce20e94ca33cba7cd8ef6c7
z83507c5bf27490a242dfe0c2d436285b93f3f05a60a6a244d73cd01796b8b48fcb67ebd890bb12
zfe8ddd0dce6ef327a79f4da1b2a3dfcc88313f48874604b9b2314202636ea1984bcee9eebce8f2
z3c461af9c97f0575709ea6966df2a8e9582f319a7e78c67240437855d4f94dd0625d211b84408f
z3bda0008683fb4ed7875605904d762b8a331f18a5710ea922b5b77ad426fd6e4ca8d68b34c96dc
zd0d6e9eaa540b5c9daefe34c092dd095c876f44eb23f2f511754874dcb760fadd3060f4f534894
z0fb9e5103118bbd7c1cafa9e57a4d7a029652384d077064cceb2d811e6783edf693ed4f30681d5
z36a2661e398848f299bb704ee75575fafeeb0828ba502a3389319b7cd3ba3a67135bde661f0c06
zde828c4daf5c15c17e77e396bbf378b971909588aa930f30c298340a46ef0930d1b30d9d645105
z35c02eacf59258f532657f255903bd8534f5d641b8ad475f6aa075e3abec92df334efbc36dfbb7
zc6bf375ddf34dbbfa4bbe26d7edfa5bc579b1d920365fbc8e32ba85c0e55f1a08b2f3aca044da2
z39d53e26b5a0cefe314206b6c09364e57d6742617365c15ab7a2aff2a388523280b974d3948bce
z1e6dba1af8b046257d9e84e55bfe6b111562306428caf6e2a1bcb89bca5ad6c9f4d59cbbad6286
z4a20260e43a097a3caf19a08071a9de41cc9d8ae3b42a3930307d21e53437724ca886686fa71c0
z1fdb0dfcd1ec6543bf4801f48c25e4670787d460b2a5579ea0a39ebc2d618fce72680a43ecb2fe
z5da80253a96b7c79b04ae34067e4dc8f4e1c5b263b481278723c557be2f4edd6c46c95eeeab9b8
z098fb08627df108d0aeddf0b9fdd48bd95c61cb0ecafd1153c13c93d6c5d03430ed6ffc276c1da
z795021f33c5febea7dc26c8e7f88491e9fb03da71526f647ca908eff0507a1d1027e122c2eb586
z557a05a6dd4d4f7bf89ee6fd9b217694c9143d8c609836f66b3d34d12d65ed1ce5fcbf4065b8b2
z7021c493b69df108506530f468f6f8412fc65a8813fd9d8010b0284652903b4997798f44ce11e0
z8ff1c922d5f9de3a83c494ea3c5238edf98344ae6104bd656865c0df3da466a180146c45c867da
zcda5638f85454631e9c03915b5215d0569bec01348701bbf6b1e11d4f9d56762954b431430d0df
z360b1b6eeeb9a65808a4d83348c1c147c69d0cbef314e7dbc5c37aea605990c948f8591e367401
z0de6c991c019f0fc18786ac76e7aa59b9aa792df39307b5d2d0c944e521595b7e75f12e4c5740b
zc65778ee9b15bff08de5b8c1bab2a7ff6d0466d315de4477f4b9db6bcd8ec21060fe5edf26d1be
zabce4512d86d2d010bf3b5395ab7a945fb6cc38ba0ccbb70827317eb5f9839f790545584cccd0b
z8236ef554a983f2cb6e58466dc66373cf4647dd6f7e6b39de7fc76835d30307bc3d1b4481b1db8
z0a1b4d4400f6592a54180c8e2fdfa297a12b4722811b5eb995c4b4c433de3f1a37da8505020b4e
zc25e6d2187dd520d71167d68c021128f1e863e8a87a39e51aea064b5c809cdc320a8bc22570dae
z88d6fe757d8bd9dad7bf8a651951782e882dca61379f628726061f2159e697af2065c0b8e7f876
ze298afbd6978ae52d241ad323c3ce9b7a311b030bdf8fbc2966412e89c0172c5cea2e76f847f95
z9c4f75851c4a8d0461cfbb53472c66fafd2b4ca3ff787725e6fb37d16291f9bf2add5cd9b02eab
za99db46bad4b066b597828109c4c95b11bdd63b307d1cbd072a232618d217e8c5526a9c3377755
z29f44a47f77b5e5e052b36288705c1becb0f7c60d55bb5ff1843dc3cfa65e54420cc64be93fc6e
za9dacc601061906c95866c0370e7a62b6e61e770e0e2fabe591b131f8d53c22e74f0902e051507
z643162287c139e7ceadfb7fbebafc12b9bbb9e3aa74cd640cc812abbfcfaaf3d31e57ca419b73c
z9612b0bf12976ef4b2296338b53893991181a26f88d1466f7c943f3894d8c488436e5c51aadbd3
zc4956894696d97618b13a45fa0a94f01a71478b6377d8a676103945a6764a4311765a5632190f8
z7cdb43264a6650c54eee68e06ce09091e3c9698380f172a7fc4848a2ed49833a2235d7b3fd856f
z113ffb8c855937a03d36b98c6d9b3f6bd2184a5f6d560894687479a59bd1d3742c6a6c83675792
zf1057326616caa7d2020ece99387b4cbb0644aab355181f543b17df38546104df3bbd4770ba664
z2ab8407daa2a5b7322fb693c393e814fcea5b0b6ffad8171f482a485d1445e7d1c78497cba2c21
zefae830bd7ceefdcf933d49dd4b51b7d0d2ddea44655771ce850685d75e01cdfaf500d811994c0
ze4bfff23fb1a4e1d9f8d48106153001ff1e47028c542a87b65b2b57ad92086b6c414adcacbce5a
z2586deac7c103a17c8be3b7c677437da5d63b44a79510a8dece85a48ab9143b534823e973e9ac2
z3f8ed07d903544f35b43b48b5ae4ea4dfd33e471934ab4b61a3791ede6225b23de5cd47bfa828d
z84f38a0f3c1cecc7f2e7f9ec63dce2c57dc7ccfdaf2256cb3194abd9ec00c3f0257d2f502b7197
z9a1063cc2e1e22b2174d7345c85b8d5c2bd5d878421263e5706f7ec8607d2008f08311e5ca698d
zf852360d0162adb6b1426f9299ef8b17f8b0e39aabd25a2053db34d28145daf5b6af65926c319d
z7af70ea30a3b2fa3d0fbff36edf710e01c986806504cee9e81f9d3ef0115783eaadfba7e42f0ca
z0d41a44ae9327edbe77a68dbbed0d06a7638eaa5f4b1881335e6965e27d3fd1d543fb04ab03aab
zb12bd433ec123f5064af3a2a8cb2e6ce31e9775777f96db874e01ad72363abd83240a6b03905ef
ze33b7a7b55acf770b0ab3f4fc3593321c5e75474a7beeb8e572cb1cb79d37a601eba30bfdb5fe7
z61a44a3a804023bc517e3b6672dafa9f8a6d76e0ae4f99f69f5d07e4ef28ddf170e4d22b2a2063
za8226a1717e624300e92d8adf71b05913aff080607e767e44027e332bb672852d7cb85c8175616
zc044cc68fb3166a204fe9555213eae739f49918441400fa5c1bd657988b32101bbed5043adf333
za6d8035218638e50a7f573a21949338b53ba9508778f1db0211301f74e948b439251435751005c
z99da8952b4443ad6c3128869ab0f69345b1d2d3f23f26eefdadf37a3f134622908dea6ae8e26c3
z4cceae59b4101564d842c8cae181702e1182781a10a4f88fb0520083490e0eb1c6f4400756bb0a
zea40eea38ff6a86bdb65c9943d589a5be28155c6a0c18508500e55152c726c5a015c6027b6d58a
zf3545722a1630453d215102a92b2064c313627686afc5161a039dcfee2827ba52c226e37b84ae2
z9f55cb25b7995e63bcd0666e19a2389a915498854454d2683dc84ddafef031f17d528e995d2cfa
z59f6d4cf96d7a32ec4cebfb0b31bf9e028ede38117584aaa58a230ec0be171cd5530d568270f09
z48e9715bf3a67e32f2a648f91d08f7a74cbe2c3de81bdb0e207074d58a934edaf7f68828ab820f
zc964da010fa0c4a23052c5409003ee839bc13e5dc215520e7101a092a41cfc7457f42a2159ef64
z2a39c34381d3cac817f4f87d8352828d2d82ea3ff2484331d1a3276eac4a2cd2ea1f4fcf34f1e3
ze83f0a47ba70329290e0a49ccd80ab883bce5feec864a32f80fb9c0b2633e855fdd180c243b69a
zbc9f5abf8fd38554c9f521c4c85fb5ddfa6b7c45ed8b25d32f9b8ca6291792d3e000b03b40d7dc
z91a04c80cf22c0c33e958dd36ee78076c5cfca5bc8692d2f5a3cf6f9752e0c8225bd98269b747b
ze5664186dfbaf7ffe1a8fc924610f07aec9ee83cf2e892d16e0ebe97000213dcda18ff47c03638
zf8820e7a44af96984c3ec9d0ea575e9e6ec16ba90d7f1318c086126bb3a469cb95fffc5bbd2a19
zb9d5bb9327a5668fb3f4a464eab5e8681ff647a2ea5b65eea5476891d532748ea021f39dbbb3f7
z21271fdd6c77b5d8f28eb6c81bd4e8a38f75047fe1d679a4307c38c79c6730de766403755d12ad
z9d5d81470ee5833212caa24833a30f8868adef76b3821def9d4d6ae576d49d05ea0300471f1000
za5a2dcc3b5ecc60bf6bdc22512edcf97ad2281624fb4fc999495bd3cc8996df325ac39d6aba547
z31fff4d0ae5460af3e3d2ff35052c53c9f02cbaa9d88208113b6a9fdd1f3426c7581eb5334e6cd
z9b1a0d6b02c98c5c7210cf188595eee87ff37344c21c6eb9cefc7e6637afd3ba879fe1a4cfb7f2
z0e7b7eac2a9213cf7cd37730e64c7b78d4cafedc6d756b9dceb58ae5790660798affbf297e9a68
z044936ab91fee80ccddc6af58d0e8135cbc45fad5dafa0bb669bd564e197342b928e2a3154839c
z3d5e2ea2653a2d9c4cce002c1c2d06b06320361b42e4703ebbbe930f6e0f28a1fee386b4098e2c
z4ad90a46a84407556a2f20847a4956612eb8bac38a074b00933db7a787e2089f2c883783009b3f
z105d24e7c84298afb96ba4a10ccf76c5a7296e907e5bc6ff077700239851be9b33757a3fcada82
z93567debef13e2a75af61737324b70d467f65033169177b5968b40111c0fae62acf8bf88d643fb
zf1f792d5c44dedcb951f7df9ab348b7cc85c5281a89a4ed2f91ab5ab0e054b43d0d6c03f088a60
z49cad77a8ff757344cf643225de36657966c1787c538f646239f566ea7986d0736c59639672465
z84ca3f658c7d5ebc13c618ec03a5743cf7cc9e2db483be7b581f22ff3c87fe13855083665079b4
z275ffa507cc4e42e66409088bc0f748413adc4c9da8fa5199e4e80a692004b148e417617086416
z27f0b9918ff3c715a64e1741be11347d02e8fd37759ad7f52ae4c446dac53449683c914c72aae9
z200bd85f50a15f408eed4703b83beaed3d91921639ccc6f007e09802c6febcbc3a438b473318b7
zc2fc6d4f845e2123c2ec0248572c37e3abe6bb9e0961996c6db77fa8fd599218f87ec9360692a8
z5eebfa0e98ebf04dc2b1ca12e515a1c3389afe2718b2d0f2e734d57284739f0cbc56de4a59739f
z0ecb26051ad189149a77e14be648457f860f555b464745dee1f3a3bfd3a5fda03253133a86cd12
zc9ed5faf3e0ee8186157f7d378af415a9d81647b55d13417effc232d024bbf74362a27d785b5a0
z1399d2b41c38f938c2d7705c157b7f1238e4ff85abcab2eccbc327388f3136f9a7d967e67ed251
z7a694dd292980e57f16388e9248e7f1e59220e780b9ce89651fade81b8a15d283d6cbfc96729ba
z718fcee88a167ad062abcd847e3fcb6f1eb1f389c6385abde14ab0447c7baa913c3cd51378176c
z912ba2c9050c81c867b81e6c350c75167d9a3885d2aee8bd04402308240bad1102fd7c62297f60
zf6c1497ba156c8ab3046a65054181ce0daa5fab377131efc72064315daf7c931c4d7f7c5f6dd2b
za2bc5f3fee313be1484e8f01d65f16e3a261e2e630e69f45bfdc4cb6aab5d146e271f97e1f449e
z6e27ede7bb89c5165c3013331ecc4f6097c8feb71fba46fce199d606570bbf595a9b2240cebd86
za53b483866b8a14ba0618b7bed01106333770d5e083f2c10c8cce9ce7c55793aaf00f3c60b447d
ze2ffec6e55b924e82b25661c3d1571f283a18810fe6afd375551e867e3505769281b5afd39b4d3
z2a8575554db42766e914057c057260ad8d06d41049c526739ce58cf6c09c2fb4e733784931c2ae
z30b52672f595ea9c45548fdffb1cc07712b373e52ff30f3e4a357fbf4090fb2dd1d9ca3f31f533
z3877e2c7eab097a91808af661834bf7e6c68e5d1211d3d9ee4fa1124e3437454bae8605e016fc6
z651bb0769a5ed1b8658882bb3d28f28784037e520b4b2d13eedeee973536f02dcbf6bd0321ca86
za9506392683eb74a83e0769e4ffe5f6bf7e60b52b03759276e65cc1418ad47cad6fa502877962a
z3e6bc4ef4e997c429cc33629c2c3785b8cf7133ee43717987856cf29eff7219236fc5105a55409
zdf06a344597cd0efafca075e19a1a61cb6b4e5daa46fd9a4998e07d8cd50ee5f12adfbf036bd60
z1d0a12d9f08eb9886815a66df5bd215c04f1ffa393c15fe65be56ce8530ce0dd63a6357e1a1cb7
zbbea541d3496b0a852117d7452742303fb5ee928d4dfda093d5975bfe214352b2ecfa1259263c2
z37321bf1475b6a563f20eff3ac913281c35dea5500f6bebfc3fc5fa6610a9e5af675ad9b5a8d89
z6d4b82ca755573ae30861aca888e04d07f7f25c2a910a52cea9497298a2f8ad269c9be76fc3fba
z6c20ad22a51cb838ed5a6883112614934e54ce8b1ee169179de01b6aa4aceb54c0c62952e093e0
z9cd7d7c9858d13acee32c737aa154127478084e4e894625e4f2911cacbf8ea08d962480eb171d0
z192a0b25ea7b11fd6c119becc898ee77e3d5f8f0ff6130f472c3f53d105544aceffcf3a17c6231
zef2179781c3f74d94677ee3be6cb107454db5cad78240a6e7929cd324836547b5a892249674f01
z7137fb414b25b55a0dc328f29da1bb7df6c7b0c3b2a22b9ceefcf1508a38d786406f2ca301af07
zae9133ca454571b10111fcf74ba6518a482801f2521a62d2e2ec4f74af5618c4baa218d4580ba7
z0e16698223f21d2a70f30a723d7312f86ea218dc9f7944667775ee9a54cb40e936c6a8037e7781
z2878d33506348a1965a08a71029f4e48c3bb40f30e538142f58bfd8462dc9fea860eccc700169f
zcad021e4ee56fdb54871f6b12d7f334fddc756e77a488b5d069d31fff85419475a47db507798ff
zc6b818075a354222d210a1c7df626eaa5c2ccc0409c2b46781c76793c9af96edc8810ad86803da
zdac02168ee18180d28f7d29735d1dd9feecdd77d597f706ea41113ed48895d0f0441676d3bd10c
z81e08a547fd48ea52f293eb7c0e6ab4f500f72f50f7d2ca846a5a4854094c459c0b54c8f29a728
z72474ed94b8d1835234eb4f0aed472d6f3eba3c0e81abee6d4fb80ca46f14fad313a4227c977a2
z943f9392931b080fa25f49c1367724d08dad846e791f259ee781c3bd3e62bd43afa92e48a7c1e3
z4c9558f88c77dcaab0ba4051d4c9368410eb112d6015622070d81d77ba0021bdad989f73ee1d22
zca591a8cd87faec1043ee585ac9d4acf3c01eb5aa2af5ec05aa95ac6639029076999cd0ef94a12
z7ffad7b44bcb3b95642435294b6b5494efcdbdcd1a22da7cecb04e7b1f1ed7b27bc4b482aae9ad
z2276603303c908a6c7d7621fcb593e538ae7397d665495aa6283435676a35330d7d6888195daf8
z865b69312857f608ff9035f87e5f0a4daf0edb034539ab0b9f61d3ccde631ecbe6c94ed23a003d
ze2530df2b07af2b1195346a5fa9e6d188ff008bf226649fa6a2de28a289e735cfaeaeb1967f5bd
zc04a9bb88c29496483fbcf1164f47597f255559b7c165cb3cec316634ce581233c07a93c0e7742
zfc8dbf637d18f86a69f485504ecb87cd46546bae206d9f9cc2dcae12f473b31e9afdb8ffa1fc7d
z56f12bb8df722c8fdd87c20f1e7d8364759949053ce38aeb8caae4648d3b54d0a64bc984afdbd5
zaab562c2172d47a00a23c49a868a2050890737c2b98aeae23e71da274baf6a8935e4d6f3aaeafe
z4b69483dd35b6f1f654f941cc4ef99ba3cbf5c677fda207a18a619768e3eb2001f84c7366056c8
zd92643bc2debea0adc8589cb958069d4b3ce4ff6fde29000f5e8792f054f4ce2dbc97012cb409d
z1437b6b4c2cb86556647a426e00f341322f0e44c1d23e0b8c9ba42cb62e876e4dbd253536de99d
zb2dfae6f61d39f3ef6e81b73ff289ccb2b2c8d24f8b12ed00e80efe37dfe58e498ae837bea918c
zb27d7a60444c7f1440e1ec22e2f185200340f861d86cd267c814b7c7f192cbe8481e1f3e16842b
z1e9c16fdcc8a9af2cb0b2a65f1715368738736a4d7e5fac98bd6890cd4e71883b7edcde1afd094
zf09995f29d4c2c719f9418fde823c84b0d9bcba4a5b1ecfa73797369413a2da3a95cac384fd8c8
z3543868c7bca9acb8fde6aca33860aba5ad49606ed3437b0daf75811376295ba6901124b902a8c
z8b68ccc64aa040382d5befa7357d134abab03a4041d2ab2f81cc5907c24d2b8778f05a77b18d8c
z6c4054793404e71188274490ec7021ca0f8d580396fb24e04506de2b93b2628a8dfef13dcd5722
zc7c059e9a36c85afe93a5fb3d5baca0763dd189c54125268d5684afc39a507bc005010ada223b7
zbd2d4172320d79247c8dda57a141d4685af667aec41d65b8c13dc071ccf7cdca3d8a9061aab3ec
z76c7e649a036f8b2539fa4a0dc0f82e9d679231408737e6dbaba68f88cc247a619d7b9158776dd
za6fd4e02359c8fbdce363b57c9da3641da65f59178ed99fdf08b8d6c7ccca7aa8bfe3e530ab2ab
z2bd1fa640d523129a4d114ff8f6e8c1036460769da54745046e4ed2a85b8ac220a84cee43a8d39
z50eed017323f3e33949eead7e47512ba331ddd7988db74629357d7f4a567c9becdbe25e4d0b262
z70b5db55cf4c3bd11576f1ef88636cae7d4c4e2bca6a38ee2d881090d81ae02bb434d302434f9a
z5a01616d409133d0c2861fefc924e2cb5117037856bfd204dc23b6e6115a787caf21f3f8d07e76
zd48a6cac5c08a67efb0236aaf3ca59d3a8baff3cd031f74b584987bbf12b3cc19a3492bde1db0b
z684518d6ab3733e0716b61f5f84cecf28b86f6665b656dbe40507f03b6b11c96ed1e514126ba06
z6a687f9a64858840c29ae265c4a988fcc60d5130fb1cb0acea61ff1bab8534145ea7c28168712d
zdf2b28e90bf67a7c843ace84b642b825ae7102f4004afaf0658bf844f3d36bc8e3416cddb5f9ce
z7b0d2361efb6cd0cfd4bc46cfb7049c1b376a52623ea583e7db48fe6a281d4f69706e98a7fee2e
z52a3aa9f09af6af33928960b53ea6388730282b1352d56f9ed203309830b0305139d98ed9f1d3f
z66e9210dd4fd8816689e7fe9cce1513acc1e1e1f21c16276c1f908cf99f66dcfcde06e97c7c6e2
z186eb93503201a83aa4b4aa18e71ee585f6c32757ee9b893d2f73dd6ecaa7c731d58a968374883
z5de42fda8ecd7cb7f66131e9222ea99656ba828b0962fadf65876e5546237b6fedbee1e4de038c
z4738eee6b2957a12e2dfc8234250e525bf60770e2736af67bfc364b943222864c00b78037d55dd
z4d32f6a0bc6c354c8db0180a64449b5091eee15e2f67c86a3b40372e997022423b438b8fae19be
z6969e7dbabb7a5fa08feff268ba3a8fe30757c8f3e25362d7390b3fdaacc0bf5d88f267a3ea957
zc9b8b836b6049c10622faeec11e358ef600b9a338861e98d3bf35c2c9a7ffe7cbb427320528a2c
z58a35c43d2ce0d59ea9903f7b95ba3f361fd3e82d04baf941faa97f28fd2951b179d38359757ba
zfe007c7eed7c9d8d4d3308656c7c81073cf3bf401c2af16fe44a68af9fca0fa721898e5e3c5c70
za981f5c847f8457030be1886685523895dd866f876947a2bdc762b12cbd73df64864887c718a5e
z279e9ea5bfb0a779c32b76c1561cf6a98dace9d0fabc38933f81ebcbbbe6c72716e48227d3921b
zbec463e34882cb75c398201f554d609c2002a90f14798a3f835fc01c784c7b4f79cc439e4f3697
z12f3a98e08c743f6afe42ecc291803a1aa744de931854da487d59f5216d27fce43d3f77c5e5c01
zc77cdfba629ca504a48214639d52c029b217bc828206bb8fb66051918c94c77f83a4dc8714681d
za7cef912114bee2fe650994bbf22c13e53227f413603de110118f8efc9bbba7d552d1f3bd230ae
zbf2a5badc7f1986becf1fffef79657e0afd9fb5217a27fdbc856fd3cfb1625c93e249071eb279b
z8b2f179bb07881d8c7de00ca3314af6d8936964ae82e71abcd8660834a8d7d7125460768ed5844
zb59cf82ed9acf6b6a926bb89685e5642ed2839056e178d163b1ff17f428e41f7a803b3011fb35c
zbb9432e797c90ef26d745f3159c7303e1ca23a2f136249b3168ed2cd9c5be459c16f8258c088b2
zb7d7f1a5e10706723b1de43e5943e2dacaf5457f40c10be0833f34362322c28afbce70b2c4e88e
zd821ab4f006201f91d440e14b9e34b01a6403ce66239a0d51d5e4ae5ed4431ee9887bc3598e02b
z89c762b338eed366758ca366ad79c00f5177a832282d29c9fcb2e1b1c170159007463967b85150
za4b13673c120fe109a2a12dc97ab18ae5c64da912b92bffefea7b0e794ff41a6f82e44659f964c
zc073c2417f04f083db7e0a06c5bb32f28a632b45026ec8f52e3f496b0f475c4942e830543271f7
ze2a97d0487042535261548bd2b0158493f20dda9a2d7a92affdaf4b08c0429d07c9fd2d0a85fdc
zcadcfa3af9223a7ef13b6f02a414b1e586e044d9fda1c4127237c627258200885c9f96eacd4d3a
z1ef1b7571a69364b112660f6f99a6fff603d751735ec312b41050cd678099b1d5ac0dd300c5f02
z36620e39cab01137e68d3e05da5622994f9c1c8f320de357d6d99b5c31fe429b12967947790a03
z9019a8d075de49e33e7fba2bc0daf59a43d9bdc0ffd723622c00b64d406e64d26e893a152ae98c
z9590afe88d5ff0baa3d5c94578024066fd4c65d3744fb5e1ba2d30079d40171e9b2c30932e9879
ze2e0e085b90ff4bf6c14a4095664def280f25c31989a6ff2b26b55051166402f49774bd67b3177
za6e4d9dd5902b575ed659b7f3e699f92ffd8307dba76db2c8dc16878c7730ec7c03110ff60ff1e
z8cca542d03bb34792179332e431db8e518fc79ef000d54ed18578d7178187879bb76b783a326b4
zbaba8ba473a832ab4e821348a017019091648f604d9993ac168e05946f31106973562f5bf0bdac
z6b1dddf950cf05169b0335e5b1f739a68916acdc6e2881f00814f66b4209c2e9ce89572a8d7518
z5e20d03cea395343e016e6494a7dbcd223e9710dad54ccc49e4204aa8e19ee9b00562023a93289
z88aa7685a514bf00930840d48d0e6a6d12e00f7d304b82c256bac82e76906401df94a7c1369a86
zf447a22ef4d349bd53b069ee9131c428b62d7717913b3e352c3549eaef7f2879b19648dad5588f
z8d5dac8530e0a7505772a28a31977f238acde688a42d83c27a4f72ca5988cb072713ae67bf3501
z774d6ef5044979a3855109db7b3f73123a220c7f85624bf04aafc4c700536207c88f944c16eb60
z43a71b71d2bf60676f2d978b832e89859d4b89fd1ab5095697dee4bfdf206cbafaa26dd2862410
z8fcc56ed6fe49fa061a45c89ce4ae503ac4f6a5157348b8bd12633cce1761afee2ffcc9378ad2b
zd6ad38f77a0cde30f29cd467b1f6fa762ee9109fcbbd8d4450c516ac20a19b2fcd0fe3eff5575e
zb234802c591f6fef5c5838a9d1fc27755933950a77830d058940744dc0c8e952e09a3ce3425377
z1931db7f22764dfec0844cba0c8f734e5d27b2d38f93d0d4d7260137595765b97217d71885967a
zf39129882c64c6aee4ff096caeb1d9644801dc882a508c4378fb0d77ce4798b72cf4ea3b733955
zcd1e463fd3ea1f4c92830b831f5fb5b7c58b9d1ef189165a51db83187667576cf7a7330e90daa1
ze92feeabf095825a4bf267a78748ecedeb0cbb4eb84e2d847ca4f18f7f2014fd6631fe72fd588e
z28fd1a8ce17e2028dc11948c94896b334bd742d9dbcf45595a72b2ef02113161226664f77ff0a4
z7dbb84b050a4742c5ee1961ccb9e5608d8bd429348646be1a848b4219932a47ad39a37a6ecb583
zb902c4758656f37da7e4d868177ce4fef1c7d2d9fe0ad1052efe22e14b54fc6edcb6d0183d8ec7
zc932d15863b6aa11a2d23d9b96be63bf9b4bd35302956d6f9d8c225e1e3f1e12fe00fbba605d71
z1fdc48dc88b65b41b386aadc3f71aa9249449838586285a393d0551227458f17005fa06d956a7f
z47f1f3e0a983c26dc433bd8b322c44149dbd73b7402258e21f71c5acf609fe494f5b57d8605173
z5b507b3b5d1e211b71f8a583bb33570668c6b27eafc533583e7fdd38820db242e79c1846fad3e6
z7c16c9d3833801813891b700735268ba7b5276b222788af6f81e9f8b3932ffb0698a214bdf482e
zabe31e4ac509970bb72e08829c1c9ead2e387a1957d3d9f221be0896a73cdf32cb295d52676610
z5210f2b68665337e8d48cc1867be30c42242465cdf2ae8793c0c7c2f357533a45683525ac85eaf
zbf47133413061c3758159454f46fe20f3a1ef69ba2e6370b40b4ca22d9ba7bfc82a12335d4d44f
z1c8b196ca2c7bab41c61036fa9cf9de127a1abb7df94084c0e708f60b7683c8b6ca3ae15554270
z56ea5ca3ab508f982c7d218e5f5761d4f711e1d81dbece37a43910ee62426c216148af3e674af7
zaf3f93e521a960bd061a24be7858b75223fbe7b3fddc7f5e1ec1bc80b0758bd91855ebc15f4772
z8736f774a18801efa1dee31e88abad765c9adb14db7c562f5261f2e5a431409b3abc4cc5524505
z41a48ec11a90e818ab8bfadef81d1d506c10cce2b1750f7f382289f7aae484fc0ea308d149e37a
ze8d7adb16a9821c1419f6e1b8e1b1da0658620181cb6778c3635fdbf7d4e1fe15eb99679c7b6a1
za5ef698955a920c05d8b0790488852be1b1ea20501a312180751a28ae3127a4d00d08c263ceb5d
z9b1714e781048c9cccbf0853500d6428be84a7c1f23277c1b09955459c40cb29e6674c34a5a7cb
z9983925b277393dda6a368a7690f89dd66f9d2e466b8e912e65896c6b08f4319e07f2f1e091ceb
z53754c0f2feeba2a937257f67a3520ba0586b19972c15982fbd759e27dc69cb86c35235e7f288a
z20bde2374138a6bc8d0e432234baca718693eead792f1e70e2003b189340bad48c4ff17b52865e
z47b38ac3b2fb284e6bb0a03deed41f99673613aa18dfd96db89099222b1c98c373706e9a548193
z7b5dc442c4958629dc7351f6ce82992093a702facccda42ab979f29b797f47ddcf9c1c41fcb907
z66dce1c5ff1f76b737bcb193eeb041561286a63b2b249132ce65152f2b879a036a17fc67e406a1
z9f05c72fd625df5a7febd980d434460e7b08f3b06ea5810190b4f3f2a879a5b22abf0792ca9ea5
z9f8977de82a624cca842bce04a5bbf068c51e2fc6f36314d34314ecec8a60f4614dd6d8b002c70
z3b15f980f7a17df62088c9d44e721398e4cfb765016fc744efa3a35a34b8906376aa1ac0f932e0
z6d13b0127f5559ac24e73de4e5c47071a999c07c51bd80bf39ab20fe4ca11cd9019c565587836f
ze5c748726b36178f1b668ec755176bf7bd61ac320a051b6735bf0e12bcb4f5ca0bbc1367ba623b
zdc65ccad3cfe8ff5d3c7efd02a9256815a42325ced81efa11f8b898e0014370249969e28e056e6
zc43d01d769a0514deafb1ebf709066800c8048f3666a000e1ca5b6bfbccba732b6dda33a62933f
z26a4c00bca1931a5962f21ae0e107459f7d1745bd490dbdcb87922f19657b08652a277c3a9c89d
z24963d40d7c7568ab0a38b48c56f9c527c70b94fe43056c623b3d3d6efe82119024ce3e4726fe0
zd989857c1f1e044961801b36f1b511b20507c8bdfb4247daec2ac25c71415fe6344c536f526f22
za1ec71d06452e5949ba634c8aa83a8d8dfa7821790663173e53b2decccf5542adaa3d76f16450a
z034d0f769181c3e2aef990a24a7e4e4a8cc2f4b6a78f6cdd2d633ce6943dd1c3e2de65623921b2
zc24250804c0451cd4661e367e57e3fbba772301ee227788916328253923f5f0d2d34778a502d70
z4ae3104ebdf443afe82e02d859d3835d02dc3de119542fdea358677d68778bb284500eb9c02089
z898edecdd9474d2c8f5baff460d190c5eb78b54ca06921b9eaf7a721da4f219c0190cef8ead1b9
z08bac8da7fc624454637dd23cc93cf93f89956f76d0060db63bc029c2df5ccb6972283fdd226c4
z9fcb187ba977695091caef98daa09a601f86afbb0b126430b29a7aaf826df89cf50b001102cfcc
z0f0d21e5bc23f76fb142a47acf7d26df7c643b966e95f0a88d6250dfdddc934d5e8da2efb4f7a1
z8f497c956f87ff15b6190b361f71a564127eefe7c2c10d9df2c400523e15aa5565d9d9206a6a3a
z8027f5cdd00ebd00d5f276c42a5a9c7e9d46bcffba4cca302fb51ff4de094ab45aa9a417a901b4
za2e33d3980c0f93883c5d399d4c16aef5566d122882403488f39ccea91766adba191cf57f91d13
z8079e4d8deb41b63a7e8e45c1a35798c1e9bec917c11d40e40103ab3a11c85fa3f756cc755f972
z9622fd5c3de6e9883ea8c3acc717891e6ef12a233429847b85a25b0689548ba54c3a310b1b52e1
z1296eef67c8de7d681e980b64131305d012fc2c4b7dec74cb63cddb3e18f98bc20682f06dd41d1
z2c563c3d366e27e698283f3ad4c1ec37f80a08c9868bb0ed47ef16172f1271caa3288ab7e8b33c
z3759ea2c961d359cae54f20f9da4edb19650dec882259a022cb70ad1911a6b0bcae1b2411ccb1e
z69493a56b412d36a93d13e08528ed4319c4ad0a72a0680d5e2ad36a9c51ba7621abdaa297a9178
ze42d14dac0ef40a977ab78c22504e59b86ca6930933b2ecc09645bc92ef9b330cefe7568a8eee7
ze0aaf08a125123d640acf908385b40d3fb817ad19e18af3fb3dc586f4679b81136c5e2c94bec24
zcdc098701b4274014272150f0da59c3df94076944a93065f18edace5e29eb8f7cd3c2810aefa21
z4819e3d75e3d101e6e12ad4397d2c03bdd0c926de163eba86f9ba7315bcace0c97cd60df27221f
ze2baebc271867cfcd8ad7624690afe37f1ea927407928d027926c279b88e14f5f45c884fc9c3bb
zc46267c7d4bb9b0477d023062ba448c043a331d2d6de716b23d9760bbd827fa5c6e99e8f0607e3
za724a721beb00a023fd2a3a28f5c7141b5ed3c737a65a7e073e9b27c94fe0f7475e22c8f8a201c
zd6e2c804bc70288380e27188c24ff55d4bb886f102aa749c0d44f04ddfe28c807bf0b287e43bb0
z2af79d313fe8a82b53ba83c2d9eb8ba7535d66b823c222fd012d47179d4f4173cb94f601499bf6
zd6c517fd631e50e9d75bc5bf65357bc693d18f1dd8bd79227bbbbfbd9447edaf1e456c83604348
z8813a4f212e1eda0fe96d879d0d2a494947482b4dabd402f3c211e80e2b04e97963428fb132fdd
z123623ad8e8fe5ac48b681b4843be8d9ca6bde900ab152863e981ffe06b6539782db09d555e640
z6c4fdd427f1067180043b9b80c4e2f607cb5fe08b20a9ed90eba330191df59add18b5ede96368c
zbc84c7468b2b0960fecae8432034c5733f56fbc5c988af0e1517dcb6643c6d9bc6143c1ab6ed74
z59c99b04fc8a4682f28ee02d2999714d5937df020cece7b7a31242c21866bc2f88291fe8cf43ab
z945a2169af02c332712be08e786bba81aca90b61d85426e9e91b6fa101bed37fca747e8459726b
z68412c7f586bfd54bad841444075097a80f0025d268771fa20d3f735a97cf25ec22bec97500804
z0983158f1a2e9cb62590d9b96970c548ef0c975ba947b7625fff52463207828cf3ea0df28b13ae
ze1a3d032e77f3dd6d4e645da2d33d3c865f1b498f4ccd1051e9a7a7dec73bdc5ecd4535d243bf2
za54c095fa0cb327ab8477216edadc158bf2e822dffe9049c8beed8f22a3beb835710dbf17b7167
z21314e50b5e9a3bc728df1678fd03d1ce41336b99008ef3b5ea5e0030df4cdee8d253fb06e82bd
zfc09f0f77ded6e235d6bf7ba681a5553b8ab238813f5d6bfcf51730558edc91937a9d01ac20812
z3a3bd8ab53d60da8dde197085c35cb309863eb6d962963d1d203fc5e495d79a8594cfb6697bdc8
zdb785f5d5decb8d55c559ba18d1ad1254df88405b924e608bf223b6e1f2d74fd7dbccb70ba84ff
z0f7a72997266d5d7d1906508123f29455626ee056d66fbb178be82a98659d48c7bd4a4fa8c4ff0
zb15af5cd076ff090ce7afa7441dce2a25aa84c7e00e374db4d07ec009aae7e4132810ab7b81912
zb3ac43479dc85d07b8f45b0ad63556976d9eef022be2f69a87b00e531f442d6ef2a03e81033392
z1dd81569b1ffdc21ec64b0f3da059ec47b85762f03dbdb80777967cc677e8b30e5565f7306e38a
zc50b1b49383dafa7d1d12237e2acc0fa3b0b444b76519ec79268747987ba813ff38fcaca75ac5c
z89cdac60f8c40d9789609aca8ef70c623f663611d89594a62423d7aae0c1bd88ad426a051f9bbe
z7d3d40a33b7155591f704d7fe092fddc074b8e31775c15a4a26901af12b4d5deb9b97d4ce2a462
z09ba61d4e21d8330ce6e7d2bfebe36bf548e59170aae66ae0ea1f2ec2fa2fd0274515af27286a7
z3108e86486fa314799b346446da0b82c40718040069b80c4cc950e3c2a37a49cd574677afa1fd3
z34e1d971401a41b6e2afc198efd5c1ea2a45515091b029ecc21af9fbaec0d0eb52d8f36d8e6df3
zc54f1c5801a75cb55d5848f7386a1d290b6aed0d341c87d89862a39b21afd31af775c573419a43
z1fcebd076e76302968fa9de94b8e89698f196f2f344d7a31eb79c0906ee03f65a62b88d94240e9
z0bcef601fa882a147bfdb60767d5e156d91be3f3271186241c29ac0c18e4157cb15f39ca32fb07
za3856d1a7043964e5a270c9029f465fe7e4920a7ebe129959710ce29e7fd5516eeebb910066f06
za2696fa45dcfdd80cf4a3108b7c220111903360baa633b869b7a4057b67c7fa75f0834a4de9638
z75c5a1ef04a933efe0d6e09b6833bafef001be00719189829baa72fb58ac38a17f29cc5671cb9e
z4443134c74b37d586a70870c545a9e8d1199bb4c78481e26314f739eadaf298da8f1489de17d31
z650db1e20f2db9f302a3eab9116779f2fd0ad935efa2a54a31eec740c4ea89347388ccb8f8c3dd
zc86d0ef518408a5e4cd18999c7abb0f9018883de2e4139ed5e16c2b1b2ef4ea25bf5c891c21c44
z98d92d8950988d587ea1bd0e26d1e79e6f6e330a75349f7032a22230ca17b8d689e583e83db418
z59d513d6eb47747ad2416891fa8e7c5dbc75aac72a966a74af84bf287ece981a93a5b44cd985b1
z67609db8644f82f0d450ddf2f00e643b4dee2e44f2ac8cdec4211f95b4e0f1e70e4b2f47caed2a
z548ac2060fdae2a56579c12f7d91725427475af1b35518c5d07104a8bf4ab7246471b08382744d
z8f831ff0b89eacbc2b4188953b947ec94a974c57eae61daa442029fd1e8277c9ad07406f9eec3a
z880944174c0ebea1e7a83c0760e482f28594ef7423b0462d69eb4b427ed54eff677dc2c2b985f4
z6844d078f3acbe74eddbe19e1eb2c1228dd97483f632ed24994613041af7387c598bb4b22719dd
z57052d0e86035e34e11e84b1cd6060287447244314d153ea9e4fea2e1b8a5b35df1fde0d82d757
z8bb144e2c3077ae2ee352fb8d25dc99ed5bdfd879cfaf5c1c110d76c05f714dec9656e78b38022
z751bbcf720bbc5efbea760986588ee74d82f69658d28c7b7df831dd39e2b56086b076d3928587e
z11b7b07728264109c4f82e54b8b7b93cc14d0b9e188eb0aa292af8a695cd854d027588aab16cee
z819f62a67baf4a1d9a8ef0d96b1e8850f320ff5a7e71530c2932c87732c9f3172c045a5ac8d950
z8ff6a16bc3239f17a438cf1677e03ab41af5827677735525ad9206dce0237f31e3a6ba5a622251
zcb6345b701b2703eba4ebae87a2d3f9b71bf6384c5df7512e99d31d57b40320c15187906a72f7a
z71aded6fafd1039f6f8bef4bf801e54c12c4c39f788c05e742b1a1796f321a9012afe4c6488860
z0dcc3a64cc4e53ed0a24d61966b3d9eb0aa8099e126ac907f3e2c1b08f70ca13b3a7528feeddbb
z5e80eb5fb6f05f9ff06378c652a0db209010f1b80adb3b3d66b0d6756341f001ca298ba1374120
z03ff2b45a1faf51335fb2d81973af4fc7eafd3bca827e832307f38707b54c82b93be3a4ebbf769
z4fdef14c1a02b2bdbaba8fcf8f6b7ad6d7cacb24ee17a560b640cb1b6603b1e1890443eeee6f71
z592af3cb42c218e16d412a5da6f10a90d648aac97a06f95a44da8aa3012e5e0d0254a0e0921a4f
z2363ebd47f6c93bd206fc6bdb60a88383af95740da3f4bbcf87d591577b977a4af469c8ba62399
zb7fb0f3ca5802bf794cb6cd17822cffce2260d0bc945d0f727207743431f6e1cb10a0f10e49b3f
za9d9402d17145ffc5d86d1daf0fedc82367165c6098d0951e59c7e69be453821436801b7eac7c2
z74a269925987374d233093cb962f7be9fc266259e4e9f0fcbaa2cb11c7e722b4b1585b242abf6c
z3a26cfea55e24c7763b11d5bc4233cd558f7929215c595500e4970227a66dbb80ede169185768c
z8dfe48ff8e9a4795e59e94a279175b870408522aa062f2ebd7e5374243cc9fa1192550c48bac6e
zea9568cb3757cb803a9e0cf2c041845dc25eddcabd0e5f786b7078bddde0fdbabd5ff5d7866b42
z027529639e74bc8dc2da1cb80148c62d60e435fd1ada2b7861dd7b04c1692d26c7799564a407c2
z0c46f9a70c78dd1f366cf03e8f5d0d6ce9c16923bafe57079320acdd2867e75f566cc3455907af
z0e28973e59b0b6d0deef2ce1ac92bbe0c625c8f29bfadcac4392e0855119dd2a7a25e73fd4d729
zad283b1082c64ec975224b2c154bbf1668e930ee76dc425c89dcd30a634a552fb37ec359e710ba
z9988ba5c686390328a991acb68278873b862693dcbc3bde8b8bd553550dda04a8ce2802c49f5fb
z867a9ab55d82be05fa8ab65442872ada329f37b1ccf47f012081ab21f2d772a6ab0eba71430a26
z37e13fb2d3299001d730e92cf94fdbe6f2a2b2869fe219f8f032ee988d7dfeb93187609e19d876
z4245948aa3b00d9fe2b86243065531b15e17de25fd0b6429f85e285c9facaff4dcac2937ff5f9b
zc42e0a0b13c8b08dcc8a465ca6eda35fb9a226ee84acf7559a389d204ad6bcb42f82744cf1b0a5
z093e21cb3146db2d86b22633f9fabd8baa31d8eb8f655149fc400617dd4bbc022efdbe31748c21
z42aed681840bb8cf074fb03ba9e35abdfe95bfb5281d3f069191c0d54bd85445e9b069005fbcc9
z3e9077379d25999ece7614b04a96f18e1fdb2c5a43d7fb773a344429674e8fb388899f1b0c40ed
zc180895c81612c8ddb1d36ad3240358351115cd10b88ddd0acf53c1dcc2193d634b42f489dd90d
zbd3800384d7295ae5c165644af88bb912aec88017d7fecad19aedc18d21b53c2809de0fa53f5a9
zb1dbd89ceba4da842ac38ab0d580464152553f6e57dca01cc57568961f2420368ff9aeed5f12d0
z050c46c5b7c3a14886c3d7405ef9785e3861e5c2d7b9bae0c2a25464919b13d0cf79e193dd260b
zd1ccbdcb7f0f6a373dd1c9a60c9ecc2f77387bb293befcbe5e635da9d6d416134205aec41ee76e
z1bd416f9b29f51e3dd9e9471ce070509badd68d92766bed14c53214a4d803553fea5164adc0aa2
z6f0ec95ecc84f7c5285e14f19781a4a3151a87b14d0b11cad0e7cfc6716d76db301c895a016375
ze8bd4ca755c4c0e20c4e91c4833b1e4fcc5e982a7fdd112065552d52cc89bf28675a9d2e93a937
za2f46235
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_usb_2_0_packet_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
