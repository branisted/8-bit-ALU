`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623157de5a10b769d98151e8110a
zd367efa3a3230248de2b9d0f01c16b4add6efa9819de33062944baf87f0e3f8c5faaede23fcae6
z5f92ad4df9eea8cae8f047478d81547b1a0c1c71f676c7f2bd9618da9c3e23442edcc9b65c1668
zad199f1d02bfa540c02610d048ba2f60ca4909b9d418890de14dee0f4bf4b9d9fa4875526e6ff3
zf3ce252e3691ba11e986b706b39c4a87ba4e0d6194504612d2b113aae4d95c24254f168fa5984d
z64aeff60ead3889fbc850156c7efd10a3f91b1a8268b31d766d9b3a3cddfb3f3e5f3018e05d863
zb25c1b02709b3f4839b99983d4d15ca56904b6e9344e8e7f1df8ba4b21f2aebb065d8fe82ca81b
z9b88e90330e044c8d3dd5bd278b7b0d700030fd487609ebcdb635ac3c93865a125aeef65f08b86
z44c9294297df5506d4dc43fcea3c24eb1522c61cb5d3b0bb1ac1ff00e52b72e8178bfa5a6e8fcc
z19f89f1b9e605964d24f57428a723aa9047098a2d80f5b2c3e3bb17785becb26e0a5c5216125ee
z17d14ae4af5a4408a0d72265add22ca664e34ef09c72e9d158c89f1fc4c4d5494b11eaf62650a7
zc33241dcad763ecb352099fb702fc6c21b1afc97e8fd456a1152eb0ca057887b6e335c9049a700
zda57bc96466880cab2e74bf2cef5b92afa936ff845ee77c6253d5de1d7f0521a419bab09ca2c17
z6fecbdf4915d27854ff06c8778f8dbbc2ab8847ed5be25f5ee6dd2c75131c70f53a19bb9b68f79
ze2866fd74fb1f0a60c60b3d1ce5b45bf347df65633d5307f492471d6c261a1272c9c3ab9789378
z61127a9aa827e2637ad0770018c0edf54ed294e0dca4c1fa76954485f043206b7f0761651afb7b
za54ca687a5294016223e40516bf459877c0d4917e6ebbaeba38ace6b596f76dd3ef45bc395cb10
z706da16ef6f56b0c7c2670b4c3ab9595faaf837ecff31b8cdb518a0ce30277d5bb2ec8a6bfa143
za131da42c32657fe36f2bf33f291b9cd855a3a02537db18b7c3b95d81d56730b75d29b093a0de7
z4637e25f95e8337a3efa6863f22afe7e5ea6f155303f066a9d1aa2190d112097e312b94a7968c0
z4affe7af42219803c7722b53c9e0b2c8ec18ae510a718e6bb54a52f0e75b3406f5faabb71516f2
z7ea6f000ddcb968c442617eb3ef746ab0e4f12924b146a95f8910b79f292224ea9948e36ebb152
zcf2568ecdc08b06aa1fc374fe5d142e5a034f019d815b5b7e4ff5c994791087869ad0f06c8ac68
z4aa34ebd470129ce9f9e82e03d47cb845a3d4a4c8c9f6807f04927b9a441052f2e943dc0b94d9f
zf7e022460e638822b6ef81892d195354aca71a55a868f962647c67172ea5126648c108343ce1a7
zaaf1a0c0899a5da3d1a01fcf30c481b53074b614a833b10f493689a12762103951be38be677635
z527d870a9c545f0e570995e481a7f03cfd5c37733805581e533822d48ca07fd52c91ace8bae308
z0cd9767105765b23cef605163f40cffa029b850cdba37d719be608ad9e360bf06080531ffc38d7
z1af3e85fe9cfa7d4fd30285bebfca6e40dd0d64584a55a968e42bbbbfdb4bd3d3a8ac1c48d8573
z96ad79b3f72ebbb159fa3ac705d9242cb0ebd9f641baa0f0c6ce7feb746ee607ea226fcf5ca2d7
zdd1d71aa471f9598ceb0d1f8f3033e49ed7b6c362ddbaf7379b6041df1ccd16630c69bebe98408
z9281b468a367379fda71121a0891f0852a1790c5e05a222dea4fbb2ebe71c817edb2353a33b769
ze6462255f544549bf9ad8eb59ddfba9eac543954e4a235a98866d3629c8f9da6e59912d41fe153
z63faaafa7d5fc8edbccae9a453c1ac225847d6b247801673f47672c4284b00cb01698c8e621740
z0ce3a9b7c7c255f6ccf805f73052fa9549b2a1f962cb387e5f762d9c1a341584fa6453d9193602
z9e92642b652128471e88404d5b0d2aa1718128b14ab54351fc66cff265d487691e6c8eb8dcb8b1
z6a88ae14cdda78dfb74c4943138418a3185049144252dd5f040d1e4241f90d24386d0aef561c26
z9129641bd972fa32ccbe302addce7e2234baa0408f7cccdcc2c90d86a208eec50e268c542403cf
z04a19175e78f2ce7c248fe4fa87de69cf3eddb32272f8ec7c999541da92cd5d62736ab33d3e4fc
zba1aaa71b7f8f6e4396ceb2c41d0ddcb328f35c0f17ea40d4daf25ebf2bef03a2882afdc90371b
z9ad78534ae3f83607823d466cfca2583b09540eac0f472997a0d0b856706da261013f4dfae65db
zecdb7d9543db8d7d2c0a147890b0f14185da0c07081a790b39934f7acdd182327345a99ee9771d
zc17c62f1c00247239e86c535553fa30e5cebef8ded77defaf536580b6937ea07e0c7f2a355526a
z93ac96ebeff4cfdb5c32b27bb52b3dbcae7ef6b7e9537199182982b85d03803587498ceae85720
z9054b5044cf7f65c42f8afc77b090b8df5137dd51983e85a1acb68352092098bc114a54684e37c
z34c3d78cc270064e376eea69c02920cb033effa1d3c2119baaf198283d3fb21325dc182524a56f
z4289b7abfd88b7b24214c351363acf1092709954a2c2ff53c4ccd859083e1bf71f517ebd4a00ab
z9981356abcbcb8bb43a47d3679a9b6360b9b97786b46c98cb87e54ee5635fe46e20df93cee5684
ze75c8caf38e187deead124fc7e2495a33d044682bbe1b75061416dfe37a41dbab751d725987f2f
zbf05fedaf95a8a0ae3655c8f922175cfd65e4f9a2e9f3d095eb610dc13a5f707345bcecba89632
zeb6822e005a1dc3054f3fccdcdccb737e024ed217c8fb0bf786285b0e623d5cb55edffba656417
zf00789cd8f3775df5a98f246128227292f3d326ad69b79f879ce00ecfd21ae04c094253b1c1bfb
z46697f007f506127d985fb742050fa95f342543998357aee406772afc5f6393c97fb2b64322bfd
zc9afd0d45744a15840bd8bcf7c846debbbd6fd8b64a1b3a7e624915dff06e89a62121c80158a8a
zadf96415b471bc9925f3dde80aa8374c0c3f6d66bb0d0d8aa65275dc4582b75924f9c783e71e29
z6d2c5e56b7a1974005a90ad927dddc2fac1010d32cb590c41b08e1028fad6a69c3ced8115a6675
z8e4f1c791b34392d7495c1aaa34d198aaf49548f674830f17b6ed5b8c450390873cab8a461ebec
z6a8d10559976c32b44eb4290bd577281ae73b392ca7e7248ecc94ef5f42502303373643db115fc
zf86148b9269779289d951b2a2101d1d2fec8f839a9312c1f1f2d162bb55daa406210d87c73a4ff
z95551ccddb6437caef91094d506e00a27820409124ed70f0229d370b03c7f48d9e46ea03786f80
zed49dee51327ddf5aea867d9e8e9e4d74934fe3ea2f51f803f8e045da86abdbd09e967dcf80dca
z77d6c7f8c856a7cc41007c66b06b01c9f9db31bf98db31dffa02f9fd92dabe3d2b95a2b61217ee
z7016c2e0c34a19a60185eca051778f22d6362738becbfe2a7fc53fae93a931c31004287114c12b
z4a660655b4051b297a4197b2ed08a9c30aa69fe9010adbeefd3f265e4c19dfd06a836e68300bf7
z9a8e5494673c14376ea63c51340a3fbceda0ad6f4b391d5689c94e2a98ed72c3f820ae06436107
zba6ad88ec5308a844a26ae5499308e7e944b0f96779df67ae6af9a7c14901a781bd0e6d9aed40e
ze081de004663c2f3c86d7ffc63036d3d1419d9a21c259c6969b698593cfaff07aabc1871a26de0
z69a5d7420c9bb52dffc3d39ffd5450b89afff4219eae2592fab27d5209498c8255c23a68ccd2f0
zfeb3eec0e3eae41b17e0bcd388fdabd19e8a79f3bb1f8fca7266a0d8fe42543afb9415ac8db43f
zea01d16f75d1b4bbad7dfab8014f68e67c9444438937b9a792a2967b8542676a47ce3533e3e743
z58e2acd90b9cf9b6533ac20e623e386221054ae2a736a6a41baec5c936fdfe54f1c78abea776bf
zc09a29fd69bce72252ea1c46cb3bd723a0125255f47749a679eac673bad0a39dec064869402cde
z974c0258f6fac8c0f36b8268dbd9eff66d5ee10c2c58ca72ded69be7e54de7b3babc123ab7d8e1
z755aa37f4dd8f21fdde0d9c2edf090fb2f90a9f6a6644da22edc58390ebd96f006592b3d3fc9cc
zd93c4262b401eca265ac9f5e29c7c40cf8b84450df29abba573dd9f0c71ccafe0386695d223167
z43e4767074f33de51f1fbc9ed68ad94172ef5e47fd9065a91b51e60049cd09b553b9171d9bb335
z8e93881ddf1ab590f1ffde191402ab6362d40b2b96afea7d87ee275b93c98cef9eec7a9d11e436
z24274166202155bf8fae1e0cf1900a542a90b3b1f54eac2bb1d04510e6d39c9ec61ed841c66c0f
zf1df8348f0a224c2a03f5f8c47af2e46dbbdf4bbd0b26fdf2ba0074b526fdf1fe44bf27d94dccc
z6fe9a279ed470898831e0fb625870d84afc0f42e6d249dffe66a287a411fb6d869f512be442923
z2c2e2b998e9a7a556c2cdf4e2c77e4cdc6bde302c61a5719bc256690bd8f90573bb7efa4c6072c
z51ff748d6e17ca36d871f6b2fd7488777892aaac8292a4ab551a15e37cd66c2929b014d210591c
zca251cb22150b88d2ca9082779161295ab20462b554ffc11cecce4670de381294183e9a0fe98d5
z5d753c742f34829c5a0a28c865dcc8785575dc9dcc5e253f1d21a2f6d2aae774ad270eabc60b96
z9f107c77592bc608548cddc08ea6d35bd817faf2d7747f72134557b3a9264dcea48626f35de090
z60155298bfdb3af4e593772254110965fbad80a57fa16b840912a321ce2d98bd945c15c8bddfa0
zfb03acfbc8998587d10377724ad54690d3f1a7192d422a0aa1c5886f4f7bf0c23776efe1e874a8
z4f1db6cae432f10a9417914912e07ba548a73a395ae9fb1391edb64505554db660c84784d9fa95
zdece836052bc007a2439a1a1d2e2cbbec73f91f767fa1dcc13b5f45515400c687e341997b0a93f
z05a989499bb8500854999cb6388bb9d30743bcc302792b975f13e3240dd19e995724d9d275bc65
z282bfa13666bdd4c963424599f6bcb7449cca10af0c448593ac712c03221121e5b579a969b438e
z7adf872119860abc02c19384ad2a7672891f70bf09db4ec425d0cb8eaeae34fbcf0c2c226c8eec
z47c6882916cc12339ba9f7972443d5babfa1af030ba7167e42f84d40be8a7ab1fd1796d374f514
z5152e88a23714494d4f460055f65008b8f8f9fd3118abf547df387baada2e45c1747183827fe3f
zb6b454eeddd752a470c1478eaaec99109bec055f05f19de28bd66017124a56be56f15a4a5f35ce
z90002ec38dbc8a889f5e50f29ad3708d387d6341c0e057fcb692866af3f68ea4cb24f26741ceb4
z71aad136db05fb72bbe99a7248bf4feebe029488507ff36dc5ba556be2771e044dcdc2082c7526
zef4b686102070885ed820ae61f880c2174625f82f4ad4f2b46289d4cb6d54553493dfda41d08ca
z11c66614305af5205effe7e4a4bd905970fd241acce41c4dc0dcf2a1f68c3a76e7cdb51651f531
z8237b5edce386c61c71b07b269896b3438e026336d37ca9d3db0e2ed28264cf21a43b2ad880d2c
z7d8dc53a1b4efe8701ea7dd5e103e24881298d3a4d53e75e220751ca56e1548d016c790297feb7
zcd80ae504b7ec548aecf4373b63fe3a59b51e0abade98f0234d50d51e8325f9b046d72827487f7
z40cb72c8866d79ba597698cda1b87164e5aa219f9f7b7a09c725391a47613dcbd9eba4a66f952d
z996054b1274df170ddc5d0864bb95c7402acaa7067162c8a28dd2520677268a4c897f33be5c998
z200794c853191ba24a63dcc2e2eb0b9e81bb1a4da53920c046e3696fa3a8143bd23ff4b3909bc6
zbd9006f218c2fe7d266c0707199222f83706e27b6169415e5b2670c5220afc0525adea30e1ddd8
z992b0eb5062087f6c4f676c0acb0a5901cb548d2e5441ecee23c7acb5c6536785c699ce1a361b3
z89417ee8d3938cbb085dc7c42ae40571e48e369efd2481d9a9e653d05c838660ef8b326c8c5094
zbd5a14e985b7d3a4e2bb69d11cd78e361075ad7ba91f56cb72b4a4e72cb65039667ba493d3f8da
z4d8d60eceb3af35bdc5c57055711358f2abd6690ea3a605863306d14c004b754d49cc4b9b5b868
zce13484bdb884d10eb2ce2129a9c61ff499a22ed9457f91c5c5de69d4cd926a952d3037db05714
z4524c82abcf1639a7579dceae1fbee699cc471385cf1a3752b379865ed095576786d86f41aac20
z0459640b318d18c4b430b5fb0ab01c2a6892dd945d15f99e0522037dd24b35f1284edd72f497bb
z9d7cf7be4064d2a457de9ab451725adaa9cf133b96ee8ba19cddacd311975a71e37ef066f8972d
zabf49731104f05d8b9bddc88f4b593f638cb72a8c740dcf136d938cd012114da1cd30a760a8722
zed6eee19e270345092ff223b5de1ae0dbf014900f3d6b73498569ba0452fd10f2f80a22ec9d24e
z029e99fb6beb9875a8df91267aa5887b10170274765b353140f089e09a4f785f848a6d48afbf9e
zc8da470b9fed0dd8662891088d1a3a3e7b310493cef79c11cee409735cab0351af56502c75f8c5
zb9c8187c4ddbaf7f6c6afad4e36109e7e24018af260ce6c154116f4f65635e4bc5bdc91cb2968c
z80705d4f3d87a4a903d8623dd58cf268cf36a9d1a55ab4c0d4a5ed5b50443bc45f3491ae80af95
zefbe706f1e216625ca93b35bd4d29335eb3dc0740c5f7a1d6345f96eb2a740b4a57d7f2a56b494
z18143e0e373281ea102af6478ce3e1713c248818610db557be777230341c50d0a2f2ce6bfbb1f0
z9795c87c269704cc6d0ae2e18b0082ebd0d48c028c13e5d4fe11edb79e164930a17c5ee41ce5bd
zcfdbfbb7057c760383352d763f0744b8d0963b66d67028f81ae92507c710e3137dee94ac7abd42
z44ab150ed24d766a00e77c27baba6624672a4fd19acc23cd6c8c0198f3c771d92f2a9ff5129d76
z2f7fb11d167c8437573f73e40c8c5f362bb7800ec3335ff6808c2090ca1995a96703e33ceb9b94
z462db2e185ed6ff0521623c8bccce466b2d0806f3282b3a428b479e2e7c21cb1e200ad21895620
z0305fde8bd6d99a49f818fae3c7eb64e60999fd39fa85ca856ed449eb8d1a619da87099f1cb305
z372fb68f484c3d7738dade28d70c0f23a86ac6157c842d06085e1d4465576b3972302d87d503ce
z44aeaf30f54c5a1269c8de3e6fbded5d58d958b90c386e3ca6c92d34815b5a34ac45b69cbc1cc1
z6858ec187c331055c79aeea530a9d1d7673f71243ec19187c02441c669fc96b25d7646d5d2a687
z265671458d068d208514af35d681a51f9ce2e0b07cbb9c588c95c8deee901ca56e0eea568c3fdc
ze4666446662dc2de3f5586cffd732b07c025ea25ada05bcd7908422562db789e63d68d3dca0852
zb5b60ba38e6e97a403164002665a2455fbfc50ab654d8c55bbc205689120dac46a8473b392d856
z136dae1727f389de5cb84e9cd6c7faab71add8615d173e1449aaa69b6a6a65d77fdaa3bbaf63af
zd60beab78b4afcc8ffde841479ca3b6e55c04b44508b71e73dae8592d9cdfb359f7129c56294b7
z3d75e89104adba2eec1b9aca01e0cf46532c09a80cff52a8ed3e91ac8067031bdd5ae9f4cf3963
z2f231cbb3ee726a878908e7361a2a2aa999714d7cafe118be82908f43afe461e6bf7daf60653e6
z4d04fb4aa79d2d3dd7ec9406de7bbcc3014b0b4c26df1e2b7c11d0cad4ee67fcedb7e49d1c1fb6
zba58b06564ce8645131c7dce80e75c2d3d81b7f09453fce44a22a0e075d6a190c1f5ab42a1ee79
zd096389e83417d39c761b798bedb28da0bfffd3395b756179231ba592c0126dfe76e89d2d7e815
zbb937392e469670aa9d48e376959ac47fcd1821900c05385953db6e09fb4f8a3772b912049ac25
zbcf4341c52c65cc25e6e41314816925c1ee103575ea4f4c6aa4ef836620701b8a878c6e70fdddb
zea4e064638c9704dabb58a55a2ed59e5ad6e3f4c34deed25cd4186071ad80377af976f2fa242a8
z9740d55363be7a1043a855abaec8e03dfbdcbe1c5c09ffde59704e96eb3d2f3c772939309e5c44
zf1ef575b259b3bb8044676d99821a85508675a9eaa2931d0788299d391273c4b29ce19f7b784c5
zf6011d8568501a2aa14571b053c492eb7d3f235c980237020ff464219c5be7053e5313830d51cb
zdcf49e4c801c08757d8f093428fded7647a1d9ce8d98ded27f33cc3601d8cca94fcf0634c798db
zc283a0d3875c03c613a41f3a5781fcf2ce12bd3ff340f421834e15be4ce7ee5ade7022503c95d7
zb3a6d07d13c684e7943fe6c822b18e5ba1444cbfa03abc8bba06d1a95d1daeca91267cf53365ea
z3a194b4b7ee6843ba1f64a669c8006eede189015128ef957e0defbf5786b5e225b56395f5d90df
z5c0db4eeecda92b641c4c1fa46d9dcd6b1df98c76099fd61df53706100f5264784c8c360eda151
z3ac021a3191041311aa46f944ea5f211a7891416ff63211734736da15b8e6ad8fae011b17089c1
zea7168ef2d5d441d8a6260a2560d561da74fb69e21ba556a471aa005c860a1bbbe871b54ce28ba
z5ec6ced6c9076430c1d40caa4d6bef3feedee74e228b455680bce29c0188e4cf02a9c00c1cadc1
z6b30dea105d0fb9c9ee6c7e1b7c51f22b7f91847f22b522d73248a200db30b03f6f9826e11e19d
z396d0a5b53fb4426018b36c3f5351526e81afc0db7d5b3cd8e72aff38004e3bd35d4c5d434d34f
zdc2b33e8d73c513332b1878a8486e0591ebd9040d6c75cc8c3ac68673bbca971ad6e29057ee932
zea438c36937613e17ca8fd20ab1cfc487ced3969d01ad60a78a5eac96f9634e04a7d263d5c04fe
zf880bc7f14a03e3695ce135a6becc2578b96c2285af294fa2c1125c28c0d2dedd1f7f49433d714
z7232abd4876acb5e0f1272fa1ea1bcefa38d7c9cb6dc23205ba273b472449085caa327afb28554
za497e75c55eeff4355007e0c1149289a307dcf381a65b0418420e848d0fbe7afbf59e819363ae9
z86d6dcf12d2d4a58b7278d0883dd248beb7f669085060e30c5c50809e0bb4fa90014241d75f340
z606919c1dc71e5b7605c8869392dbb4bd7007ac4fd2b247dda166832584a5634b9bea32b70fbcb
z554b10b04b324ba013c75c076e338dc83612f34be6a8960638422f36d13eb3594e33063e0cb8f4
ze260f73c0a3ff8bce8ab4b51c4720bd189c4c85a40a82dcff2ff48324059f3746dc726b19907b0
z35ab6a9c3b89788e49319868ad5edf7b727c05ef5a8db997eea9d247b823acb26494209ceefa43
zab5c591116e9b5ae2a811b1f63760126ff4900cb80d4857636141f476ba7b71c0b8f05ad345aa4
zf6e8603e2d233758e7b30e181aa5628b1ac30db30c6a3adf10e167f6ed9fc4c031cd6930e79790
z09043bebd9c75582bb47fdd83ff5d9bfea81ad48083433ceb51d2cd381ab6a4644f9a2d7f48e5b
z55e534c726284a9daa98cd4cd4a88194733f176e07fb5c16ee6bf3a9b07c00b8d2671e366dc6dc
z9e3d76cec5b80448574114b7122dd1873a2fd7fa604b32d8972317725492583416b10f9c473391
ze52dbcf1a0ced5fd4ca3779e05d5f7a3688f0d9eb66b41f708652f170ab774461672a693a825aa
z1b8e430c97551364a0cfcf26053a3d6f321c44c9ae58507130db86a3277de39af71ba78df36b1f
zea167ddb93bd861fec0f776720e61be1f8b9da449f410c978cece7c022307b310b1af5fcec221b
z0aaa3a40f34bdca2467c4eb38f718d781794dfe0833dedb3d22d9d46d9fda926333d93d011e859
zd930804b8f33d7054841e2e4dbd79ea6d0f8bb628900a31a848db9155666cfce28372b6deb5367
zabcbf3c00155b2e068966c8919d0c6ff6537c195a730e89e809dd0ac03e5a65b1d862cd771f102
z223d41d8119418179d71d2e7cd3a85b80e107aed8f5c3c9fc89dd46bba2d0912ebc7e8b8afe079
z0595a4d9310a08dd0dec122bfc79d64548d1a443a0b55ee32c68c7099dc7ab02ccc1a78941f341
zbb51a67a2d092525fef7c16bfa64ac6be17834522a2ec9f995c5507e844774fd33ca9b5c9c3abc
z9614f8deb955eeba20519b77e15b06985945e174306f6e0e537bccd2c355995ba98521f5b9ab13
zee11bc9d7d695703145c21c631fe7ab08d6ef9c0e1ad532d201466a5cbe31a56ee10d6bef59d75
z781543ab5728989a82869585b05542af18d079001145ae38f9113312c13e43108c8d83bcc02632
zcf85
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_xproduct_bit_coverage_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
