module tb_alu_top;
// TODO: Implement ALU testbench
endmodule