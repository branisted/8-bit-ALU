`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026201628cee5aae21fb892db766c4
zb5b1406e11aebfd6dfacc9da5ec03b70c276807a3eb15e28ec7ab1dddec42388b9424ea285623a
z248195c9f894b36317ca6e59c86f11031163f5f5e0af432ad71a370b503d5afe29967480e0ac49
zcf7c756f92650aa81b43bb5505acefc12a9333c15090c386c323f8cce4e7934214caea9fd9c42b
zdda79bee782f6c797ee18b17b0c257e45bee7908de093c385d7e8a753e689ff7fc8a8c9e7ce08d
z05cb3d56bf84f1fb3473afaa2d473467ed0a852501771349b43fde42b4344a1328f0b9488ef772
z0ab2e71ab13ec995ee041d04202d900d95c299a1c207aca6e4735d4f3857211f278f025542d047
z1120c7526d7c7aca9b4535ac2a7c89914a071ab6e28ef5a017369bce3e9ab2a40b1045e640a03f
z1eac01f38537c460592b18e6569eeaf3cef2c2394144d0b4682b5a48720ec74e4d0b2c6180f2e3
zb86b55096a5ef9be48293937fffbe514105bba4c72b420bddbaff7c98716faace082ce2b7270d0
z082943369f9adbbf070172be89ab7354b521930c5a900dc87238b1766e67b7a0e1191854639319
zdf1223e075dde8a5cf288060271fb236b0645c68e01c0ec3232b83e1cfa0e95b47ff1652160747
zecde91b28ebaf7a1a398cd45bce9bdfb59d8a39c019333c8c70a92757f3498ba94a1700a22cdc8
z871aa793ad3267f5ff895ad9188610226db47921a6b2373776668a9b2bb5daa92fee02383d142c
z8b55f881e25ed88fb59ba9c730d78bc55a0757a3afda6902bf697868acaaf20ee3ab8a85200ac6
za186225ff0211433acc05f5df1c2b0c330e70a04bdb8ae144ddf093ff61e1e143a2dc7814f5445
zda60f461b3cc96c31c3ffe91af592ab64af298369479c6402812a8f0aef1298bf74b9348aad66d
z7096e30f35ea4205e6181575b95d59b1704055c6530760412ce718eb5b1e106fd6a179f4165d39
z8b30846ff76b49c610f1199062e473940596e20516e2a4d93413f9b79c94cad57b5fab211ed856
z7548faf36b57164d3e598195148001d10a1ee6944d21f69599b7b4002edf2846bfb91c88304bfc
z7c2ef11e4a5d4955d82d2f79e0f61ce32e3e1a32d73c6aed2779ce5d7057401c0b53a1ce86b67a
z14dce24a1141fd5577a376b61629ae692164d11b92077cd1cf211a69967e8e2507bbb7b018c668
zd3a4c8bd78ccd7e3256918367dbf654b6c0c31f9fc3d170253249aace4f7db3b1940d44f44c9e8
z4a1c5b5ca99c3087c8b889dc4e453c650040afa921ec3bc79711a8afad1e6700c6508a487142d6
z1b495436115e5ec58141e54bbb74297e058d57b8bfe505d384b0857689cd22076b5212bd3ea481
zd881d2594bd9829b0183212fdc49fd49b234b87dbaacf31472edcb89d34babfece7ca2050259f7
z9bba58c8d989b4e472092233d94b57dca47dc69c547969363949ac4e45dcb38c20478ad0f76e52
zee812be562af73ed06cbbd1afb19bb37840e41305d5169047d9842b7f850acb1cc71924aa55fca
za56ecd97d5d2fd19bad64f8e43fe3326b6e2ae877a910982d87bd0d607ebc539576f81096838bd
z032f50eea83ce5060df70f577ce5163a92a2bef3b59ffa4aa098c7a00b39ed48748b7c232b4e43
z1fe32df17673251debc24f699efb28168714094231f3a47a9cf70fdccef91cbc3882974cb5a59c
z9e3e019bf96b1dcb63c025425e149b13932511123c2fdc1b697818a84f23c4b899f717dc37633c
z71a63f60774e9a418056c6156492e7fe7f8af18daeb5b3c81a2bb7263f7545eb66317a0b216bdd
z1d7fda29344c9dc228f16f133333a1c4e471f1cc04aef3f90884acefb698424bc6c87b09217bd5
z868120a3b350c3742543ad1b3960b15b3af67bacdadd7fe47bb8fe41e96d14524b97a1e88728ae
z25bd8a4f76309d1ca4ce35f4c4d8d78ae5411bce4f761323b91412ff88ce7b34795f25e9f4d30e
zf4133861f84353669d9a81c7dca7ee2b306a62de23f17632d7792479c2d5acf9a6316e0d5d93e0
z765be2fb1eca748c2a6645205af4c8d9d7c8cc9a840ec8307d02118facaba0388f05df3223d6d2
zf2defa5dd5796e268630731f48d471fd9f16a9ee151b5825bed1562dc5160424ce35fb74015be8
z80db3721076d61e2ed644ac939344ec61a33952e45998f621994ed20760b49849ff1a3deca4abf
zba334e4ae5dd7d794496b458e2e9ddd582a41d0ecbe5e45069072a209a08cbbc5ee4e5e6f5512a
zca68a86293df4bf3881f737a33d8954583ee4fc46fe4e7ba3a8867ed88afe153393cf470ac4d67
zefe5cf87a143e7abff710ac12309084361b46170d540780dff3fbf21312bd3a28048e618cf27de
z9f1807d2815755af6079fce1c2a5531fc98f51e91092bb8dde3f55e9832980b40a0f7c0875fa25
z61be7d40d9b4bc160cb8d3cb144d916d25d3548123059a183d79a9a132af804a02cc548b06452c
z63b3aab32df32f3e74e1c677e54cdfe273eed1856eb8c5b033752423c57ea0c4a22367a539d0fd
zdfe2a4d751a91c0ae87ce35cec2e1c8fd636a3fc922712a799e9ce96485d9dc975d64b1f610c2e
z86aed5cd184133dc9c19c446fb2d293e67a11d04d84fa9cfec363992da7d601a362c43dff8c467
z4e159cf9d05011d57e18051dc44689d8451d40d1c3df36187feb3f77a08643779bb6a11068ad81
z47b4c6ee2d0ebada2ae266464ebba1e4383f6731460493be17493696aeb992ab5b8ca735154a4f
z58a3bacff7fcd22d75970d43a1bb0b1c2af32768c979667ad2445198ff998d16c50494177879e3
z1a7d0e264050fc7395ef8206b590b8ab6cce2ca633c1b2f123d227c33da2761f99ba8b83255075
z4e658ded24e3afde7f8378d2058bdb094dc9e9f8262121fd556e616255ecf65af21a134d41b4e5
za221a31670ea5a00a43772533f91d1e4dd6fd2b007c28c5a53351960febde743ab7c70b47a23c8
z237ec7eb3f584f34abd35a42c8f45bc822ce2e891bb5d9ffd43c6de71a4ec488b06c558ba64593
zedcdb0d596abd40489882279abf38933962072aaf6936640e20714196331915253e92c8b0827cb
z7751a3a4c6563783a7cc669abee44fab4e178ba0e0ec87fffe5f8f36769aa528668bc37aeb2072
z120f0cbf6dde0591b0e334392e6da44df36e7793244017c2b8c7b2585d3a8d3cf9f9ecaacfee1f
z65e0f131f4fa0e943a1543499cbaf5cf4b63749fdffdcd757b154eb9cd147e020583a3717e4e08
zb6ed41f7bf249bb21843904694939075655b0608c63dfd08d8a29ff1cb3b0f46d96cbb350b9872
zbf2dde0c225fa45f242e4becf4476649b54a78cda685c5ad86f5c5d1d9bff7550fb2e508ad8211
z7ab7e53540ef3a15a044672dd652f6d6c8ece1e7ace5cd49e73de7decf4442f9257d459b0085f8
z83bbe6d5f6f3edd894b57e97d44188653972c61df117c1245db4a22a39d25f210590d078ae28f8
z633952c85bc533201dc7e96c4e8b257580c2e6e50141eb926470091530ad0469e8bdc6f6daf9ca
z01218f849e1cdd8632ba031e7a27b80a793672d6a37798548fd79535d518231b6efc99de64e112
zf2325b5ef6a821abbb71d3a4639d677911f4381fbd73660a415120f4935c20e8134af24fd7c723
z3a341669186acbdfa50b066b650e10515edf29445eb172b500f3d2ccb88d323a28477334d5ad25
z0d3e63c306d01df2b67a07182602858736b5d2dae0d2a4c5d463eddf0607c3d52fbf97e15e7b47
z67b07a30ad33105c3e8c0964ef3c3243b7760f251ecaa768cbe4856eb856ddce46d0f43213439c
zacf5d803ae4004f6b04afb777ab5f063f70b80bb6f5e6cf8e8b0536dfd2138366c7c3dccf22be0
z0f147884d0b8def890cbafa609482aff6fbc2ebc40784b56701ca796d1848537af4b87f0dc65f1
zd2d74ea1b3a6e3ee87b92296b9836a1022c7bc196004c96adebfaf0f87ea0fb52af1a56e536ef7
z11f1dd01ea9e1b696c3c6186884697054a2e41208164895e9ffeb47e7e613368d17b74ca396e85
z1c7a095b336b22b097777c1c681f34d0ab22ebddc6b0da7447dd755d7c941e541b979fcbf91544
zef74c354750498fea2a61dad8d39041c91aa57cf30f2f883bb93ade04943eee32f942758678424
z6996c64f043faf459443d2c95d5a628ad37f9846ab230c6bd07c4c21561b71d883ac58c651ff5c
z4c1ef7b6d031da343c3e19e9801a98c98eb836cb807bbaaff743e7c2a6e31b24353b19075793f1
z4b44d53982beeb7882fd6aab888bcd92d7a93469ef9beabd07dda7c6d3bbd0f929f5cf97b88029
z57cb87634f33ceda3485c798b1eeb89294d74b103ef55c716e9a2c3bc05e86bc80086ef39a6233
zbdb0ee3ea839be2e7743c815d6308ec8cd1aca4e7c7f9c4dc567a092bb66a14a6072f7a9e76d3e
z37784a1c07bd06e9d34778de2676821a502057f646e0170e3d9933c963c5f67b4e632426c41b48
z7eac3a33a3593fcd4ed1ac70a060c839e3e7a2e1f5d71d64f7816a434a4e905898cd9e1542e9d4
z3f7cd9970ad77d68dce25381b4f22f649dffe6fced267d2408493b191df8e36d05a9384874c681
z4a4a0a7430d77f0e57fb1d40fb328082985803b27383405cee11e10c32763506434bdd88094711
z5b9a351b652a95d06b9f13737eb7995efe1075b9b06f89a7ae9367759c384a25a91280e439057c
zde5d1e72425f9eb4f967289520d1ad781a4d4058bbf25f74d1ab9640e7b59ef3eab0efa984bade
zefde8dc5cb9c003f79e8a266c8a7f11e5aae3e9e3126c3bd85e6ed92869b07c4ebce25f767581f
z1d9afd87b6f0bc5dff30f3b838abe836bfaa073a8f80d25bc00db4866bf7d6da72cc2aa55d47e4
z612a03a26d491b0f60d07b83616bb3a73701c69060cd3f6dd1da9e13b3c8d04a379038c64a4754
z8e284b1851692d4cdc5fb1a1e4a4a930fb57708ee599b9a4da4e45e840e98197ce870ac3d5cf33
z0de1a920467c7e423f66179e0c6fa242bf2bb20b0455b9759440867bb5699121b7cfb119e3cc49
z4667cad81e1b754a280d3cec210265240e325a2abb6adc2468c5e00bcfffaa0027bfe7edbe9e7d
z8db0963d9267e3c665e11292b4c48a7b2e80fe738843317faba854e0f6981041d9f8c986937093
z8643612dc873f7a63089e8ee33f806c684f73a0dc298877c7d0ad603e7defa19071dc61ff911f6
z7945202d6b2311eac7da0420c1280c3bac4b8538d5b8ccfb7b466da4309e7351ed45ed4ead2984
z3cfb53a928305df4cd501fc370496a76511e190cc94f76956ff6c6cd941531b84c8e1f56ba9a1f
z329a2a4be97abf928840fe57ee4ab5f672e62fa8585bcc425b72389b9faed58be3fbb842be7a8b
za7a5185cd2833b1ac44b1dbbda928e80429c223a037e16146b7ca8e95c4ae7b18c10b36f372420
z2b916fd2b5a05ad39618e9e5aaf1364fb0b90d4d6c7f76712ec829d8dbd4129f49c76809a8cab8
z33ef9bbcd435033c8129a7fda6f9142850f6e2681a63007f6b6da835c37e3d739134dd8703cc6b
z1b195233e7e6e42f09addabae97341f77274e0f03b9cb9d4ba6fa595a64328a97243c43a8e7a3f
zc30a3b4310e8bd40472d0915bdefa01fd87a88dd385ccca0e60d36486dfe01a46a40c2310d13bb
z697a96552f603d6280dcf58bb5557e8e4a1c54cb85ccbb8a2c9ce81508f758fe96ad7a50c4314c
zeca5979e01a91b32b3ce06ea8cf7742aa4bfb2275a5838e9f4d6e21d37d538d6f4e5ecd4ef9015
ze21560014aa46e7caf5407dd150bd0fe544107db6cba6ff85a13a73f7f3931d036608bb36b1b65
z6c4d99de3ee2430ddefdd64dbf6dcd90baa62171f03bf9990d20f4e880ac49747a15f44ddbc693
zc6b901d036dbdec597067750e71c0c8a2b6fb6e0a9fd2b2f60ca7cbb4b5aec4d05b938f7e2d814
z6f576735cd9fcc9fe900ce51a62f6a016bfda129876c451c97b6e23be295271d83d9a7c7da5e8f
z71453155c97f63cdcc61b3be29e1025dcac93355a6bc2ed1597365b09ace8bbdfed44a8edb9499
zbc77dcf6acc8b03bfa1527e5d298897713611d64e402c7deb26767713e4271f7ee49ca05794391
z69f567873043baef1c225ebbc64c1df88ec097e2d7a1b2e525c234080b9c9ecd89038b1fd5b2b8
ze83e017552db1b37ff5a7902cf6a2097d2ff4c9f1aceae1a96a8ff410ad09c6688e6df787e13c4
z1d8703e0f7c5b298870dabc85477c5ebf7a3c1ba6bd983adf4f0d32613c298671e757acf8be50e
z0e6f0a431e701914c723bc1bcee8ed1cc88d9c38d223c79928610d64be0e4865e20f8dbc30a2c9
z631c7e746531c93fe1be84a9ed5199b1dc8eda2190d88cf9b7f97f3d6ebdb34511e792cdb0d998
z72fae93d2cb07c668894285c8901645d571ba8176d71f54bd6afeded47da030a88188a5c09090e
zfcdf95a467f37b91456409003036ed86844f9373e90b76c5d557fd9827ed53986ee41cbd3ba057
z1d548d80cb6052ce59f4c14b53ce9c9a6ffd621abfdf112686f0cb72c0cf66ade4a5178b88a0da
zdfc5c863e9d273d2f7cfee7f3a0577112a9cb013f940a5890d731a799dcebd483438248c07ec39
z16de4acc0a4d6f36ac001de3b9e2bfb75218638892c35057c95cf733105e95ad20c930da27b367
za122cc8032a6ca35f89fff30e5926079794bb0553bfb9cfa99e6ca166cd00ac127aee564140606
z49ac7395c24a3018850130e8687f8e47d01dee395bfe9e4505dcebedf7667fe4deb4cd776685c8
z3fbeff8bb4d0f6cf95a6e4ae3782408384fe04981ae11b185818ddde8f28a89eb4e0a2b97e0c16
z39b67c5da52b51c0d14835a0af2a3e3318da179428b798f72b8b40b8034de583d2b53760925c5e
zf076f233a771fcd5aba6fa98ffbcdb261802158c31e441d907e2b6ce998b57570cf928cdb94bee
zcb7afbb0a1d9c76a09b6ba811edd9bfb947d78442869a8228f95a00b7dadc5d939e2a692bc6757
zc1611298bc400cb0fec6afabf220ad11beaf6f47afe6fbd0eb61299dd158690a16319edc076f21
zcd8cb712799ce79eb9ba38bc04ae03b4a5cf109d50b848d945b9ceeb66ad4ba2a5161c4a70f96e
z1fc45e13b585b8c4db4e41a87f9a006de237cbbe304d392c510ba6e323d9eafb337463f72a1518
ze53b705651fb15ebc33ac8f0e6d9a3809e772acb105b054feac1abd0e1e781aecd460b5e3c9c55
z631cac3265ecd02c41c893745a913a54916f6b30b5696053dbcebce8f86898b7e7397a1e57a4fa
z0bafd3ea9be928ace3dae336a256ac84d8daab10de732267088f2677b9347fd5163843bc3f7ed3
z3ebd3964e146b6a9cb2cb72e53fd9e55376ad9f5a4bb2a75f0108673962776398c85cbd77538e0
z5137bed7296440db873bcf1d1d853ec51dad1541ab3e7576a6d2937da56f41dfae67baa6e6e31f
z2f499ee70fba2482ea2853ddec33cd94cb1211b540dd18754845de4554d49903790a8d0274eb46
zc0fe9cb8e8ad283a6158bb0edbb16d8b24bc3d8c109e1479bb96cff9e9f1019a72660b9c65dedb
zbba24ddd7f1608cc665e5780c9ea7b92e7f403224e2b023d753190b0be1cd145f15799237c1b47
zd2d1a57fb9403d1e0aadafbe5ca285685ff5f9a00ac2443b91afea2d34e8407aa4d09da516757e
z2a86f326895ca0bb244cf64199944a94238d6a3affde372431e69110cea7f4c148397b0066731c
zc59d17ed64130f818be1500b974b3b4edb0a54e29431161b3f38be931e7f140f88f752eb2f3787
zb4e0e679bb612e4fc81bdfde482e6167e960bc3358aa7a5054714308b76afe7ce1e9513b24b99e
z52317191bc672780094c044b92fa752462bcadc52920395ea0e7c1873926d5e3989c72bded3646
z41e7d0c1f85ee93bb6b5e21fc833ee97ef39c8b6b5d184113ea2c5ec867e69cefdebbbe74a7ade
z94f1d42a2d7b91bbc12a9e9d0739cfcf26ff744f6dcd3edeca8a565ac46f47f1127efbd445bca5
zc919b22aec9f81d2acdaa7a5979b8b0893918f7059b89f01da6d2fd61302e037becbeba926a8f6
z5a6a3b4d352cd93723ec6d8b19b901c37175764f7b5ce7c14e4d34a879caf2ff406a3ffefff1ac
zf94a735d8edbb688638b49cd10b8ef25f4ca812818d2ebf509a7316938e36f25737d48e8cf5df6
zf487ddf0fe62c3e5761edbdb2677b3c236a050985e1957323e8b4a48f728f0020a5aea79925931
zb1963777b0181d3455b4ee42d9cc08786a6db1586bca1463dfb91a661d41d307eab8db34c4bc32
zcf504011ccaaa0087cad6da76ce5da19c19322dad80ac7e70f2ce0a14c14c73f69e2a0919f79e1
z82ec4d76449ec6bbfad2244eefcc4e2e390725395d9f06b052a1db04d4caef1540cb185844ee53
ze1e4c68810a8de4e759ed95c2999f88ce173fe9bc3cc3ef445e24f8fcc550b022a5039475db2aa
z8eef8f15e83cdac0825f7fab06e92d15818c1a9d5f398ff235789f10f22fef04ffb5dadd60522c
z73fd0758ceb7f3b9d46310653db44ab82c3bbfb6b1a85c95745548ddc1842d87b620ee683e14e7
z41111aa141ceb8d29a0fa68f9a92bf85a80d0270441792c6d89287d4fea6a4bdf492c5949ce1ab
z7b7d55d0d9687a2b005f174ba1ae555fb5d55fbb93eeb9cb3829841c16525efb57ae709f226443
z47c4cc7422fffc04f1dc01ecb711fedab750d8c8a99de9489c85ab18308ca75ac4381791d524bb
z9713231582adac9c72f6d8cea342b5813e223ef9601005fff284d8ed0a79929c592e3ff90cc511
z43eb9a681c0f72586f9f54a9d2b91b27dd3efa1ab077ce0842d89d84ee9e4127449c5da07fd678
z67b3575e4572b55fb006120bbaa901e8c108fb54cafb3688c2fa30d8e24e9175d557a0b120fc5a
z59786c4d12b1a47b4f9a07eb9ea727f864ab8dcbae778e183350e6fe0344eff251ce1679514588
zf29431fa40c9d466cf593ef50737e438df110a3579393b66d810d50ab61ad80e2ff58f15de4a3e
zdfa040488c653e37854358ca1050edb42b7d1460a906c1060d7d68e7ccdf265e707ba5cbebbe23
zc2add59387d12c553b208ebb3e89254e1d2bc2fdf57afcf6c8bed3e7d3500ab4b7563bafa0ceeb
z21aaee5ddc6fc16de974dfddf886e069776f8d394b0d7bd19dd27ae8d10c738eef0b83bd4b34ae
z03e199609996e0a72feb74386a031344e2dd722a23be1ef853244a1454b1927d7c0891e5f70a13
z153120e6060e05710afd5aa0b1b51c97b97e66d519601e54235ecd9d551aba062653a8604f398c
zd526d5b0f55ad62e73446f8a81c173c9ebc5d98b1538ca8a3d238087b7138efc45a9c287c8ea10
z5c736e0b40e43f80d3886f7c41aa20eb88193e9fc0c93e7b1c718413f2916e795657631c219caa
z18e5e9617bab1f44640cc5891a29eda97bb27cb423da61ce179855201e7a421706b363d2b64962
zd173e0f6af417fc59467515565de686009bd66ed4b9d578d9d10adb6ceec65db68239241cb94e6
z8c2ed12541aaeb295fbbf900b40796fb300ed5feb3284f918b7e4a9be45db7a7451583b4bb667f
zf5d7516c85f1644fd4af63b8a59776a9bf6f226c55d96cf585d579f781b0632c06031701c3529d
zf969bcd55e2ac459f4dd85879b24ac321526e7ef0a69913b551961196fdbd79478848efd73c6c8
zd1d6b01dcf91bd024119cbe7987ceabf7964c957c936ed55b8ad9dce5e5f0f6c969b718a4f7874
zd41dd9d46bdd5ff5b8e789686c87ae05feb109db7e83e765d579125b0f6efa5d1aa9de1a31ef24
zedb83e74a0fb5460e5a8d69b7f67ac055c1f1cd841a0c98c230fbd2e968827daaee65b0d1c825b
z759b5e8d4c102ce0e0e07dfc2925c634c7bedd090900c4d183d3dff395891a7af13ea19b0e8040
z75b8e082bc904ca18699fd2dc4771674738d787bd2ccdbc7427c274cc1b0baa6dd5484920ef25b
z23abc3131fd000929eb2ac4c23ac59839e0cb8aa8abc8a3746b536eccad507a767968d3b8afa75
z964af57148905ebaee495369a845d573cb7893efa974cfe0b24a0f168c711e55df10dae602e8fc
z6a2373c5a5e70f6f03d69fcbe22ce1b484b7aa46e39442066aeed5901de7bcf39b4cb8ff645d9e
z7b101f9c80f193566d99e6949734c43a180527b64aeea4e898e299d44bfd6591f4abf7f36d1592
z5e537b8856689e2af1d516740c7e823bfc93c284c9a55580c1a4bc98a01f1e2cc182d16924f77c
z7e25a298061a4c77c266ffc6f291162f2489dd0955f571e30bdcbfdf1af122b8f742993d2cf378
z27a702a181e64b88e577f9770b17234f61a72e9bec7b016563ff5d62c0e5f625f2b8d660a55d39
zc82739780991ff81c4649c421e95a0b4de1a28fc89566562260a8909fd00a7830d21825d160bc2
zb7af9d9b10d09e6742a038902a01cc980c4b9de67c09007d0d2e0cb86e24665cf1595272a604d0
z963695198d20e6ecd7137e87d6ae8513c71b04321e7eddf82244c0cb15ca70b64f22a104b261a6
z60af8c5c48f5ccca39548d4508d810a31cd770408552e101355d66da1ae1c15f5382a885da63ea
zdfd202fe907e041c31482dcff21adb1bdde718ac37df53a2a7f37359ca59ac899c44c7daa861a2
z6af9e30770e4085468904431f4ef8f28fa45479cf63af35d9a88fc1190444e1e3463531fb9f5d7
z924b05dbc1b7ce8af6a4ccfc64d5117b8533f16978a8f5156318dda5b5a4d106ad3ced95c3c57e
z39dc4566c6fb3cb953cefadb9ac95f17e21d9f811147c2a4c782f6e1523cb16d33eb2750ee3b1b
zffe732c0bda34e4c79d2a33c3643c96ebf21a0f550cbee0e57b9a4a5f18fca4a9517b2b8a61af3
z116d446a734f734a36586097dd0f7ac70a3272768235a32673222499aabb3ae805e71f3ce70aab
z41c51cb5601acde1f7e8735618dd1a9d713af1e0350fb0bed3acdb1f7557b33fd1bd47bc6d09e0
z75d8249ebf30bd113b45798a3346726eee123b8f59ed160f89c48c1160904c9ba5b2a9cc549281
z520748166a1e71cbcd90ded5995da1c1e79c143493aa3adcf2384c078ec1c53f80cf3000ffe8a8
zaa0ecfa094b922489399344b338dd1fd600bb93f69ebba66635bb0f7c487a5a24f28ffd5575b8d
z735977c5e96f4befe094abe24bb442489bd1e209277571338946ee65fd2a121fc9fd9c4a66563f
ze3c1bda040949b467451094295c0f4ffd952940bf0b4c68a71b7032146cd004d238de8a5941272
z65d76f01c1f49c7cfc0f6f55ce19aed87934e619560b6040a7b74c7e2dec30e691c72d0f46419f
zff7309b77a3eeab2881afefb5f548e389cd26afd6a41bfd32e263c518c1b4bdaaad8bb58a63bd8
z6c88bcf1e3fa53fa02cdd1f6bfd8f8e7ec706e01e3b1b09265d89b528a21c57b78015e361c1170
zfbb8d15a485427b67873ff3a944035e313378428b9c5f73b0e9c2be8666376e8b1d66c5a1cee19
z22055e39709449b3e7ec18b9a2d291d168bdf46a1dae1e842f78d3c26e0ec1f3061895dbe8c557
zba4131d906c595fed911610e31e695204dc7750f7084ca94dca2c3e64eea093c1bf7ecbbf44561
z51db8bb2145ed5201287d52b80b0482f07d665a4730a48989e1ee28fc74be38d3ff546cbe78eaf
zf03d2d65f192ad490c71fb7f851392d1c243814b9276b65d7e9f54d2b3e7b38538a90698003ce0
z8432bd94b20cfd56602036bdc9d1934d3f42d241b7b75b8ff1bde3d2fe5c873aa2b3bc49f05cf3
zfb67317566b48820c74a6baa6aa9b912136ff88bd3ca061a0015f08ad7d1369a5792a5f4ca0415
zecce937057600075458cc375ebc2b85401d72ed090ec374b651743830f3e03a425151104f6220c
zfc9a0bddd124333e72de3fd46f77781e6504783c241ab8af5832d740f16b41943082c00ecdbd1c
z4d84e7fc6f0fe3a5131261273088efae70d9803050204bd19545fb709a27ebbbd85bbfa2aeabaf
zad35ea07ab4573ee53fa56ec8ef33e4a7788a808bbc7ebf7d0fe9cba00083e0438fb898d03a7d4
z3b40f4a91035d36a455002fab5f8d27ca0c1bc7bc9de9195c12242ec0190ebce7fad7e850e5b80
z03004a25187ac93d3c9ffd48a0b7e1501ecb13d1e03f16427909c1ad57d5515e0d3e886574c8dd
z0b94e4144bf7e15c032d37ccbfa5911bcbe313b36e9e256baee90ae5d0f9b88beee513210ce420
z6d7d5eedd4a374ca6b73098905da9f124d16eb622029e7c2d38ddbd2f174831f88eaee36d10f5c
zff817f924561045a30a11b73bfea9b0430f5ac291c1dfdc63f13221be3f3b2816cdbc62ba55334
z239f27624b6907ee12100461aafe38a3407dd7eec0dc6261a8c97f511056188e057542b81ce966
zae29e235e121e3247ce526b1dbcfa537be1631c19b3a2584865018473bff3b346db29b7c0c18c3
z95d8f55d1c9a8d926db39b493b6712d7c788a73e58379b6a95e0e804c9f44702feee60c7e799a9
z9bc72d2e3625074f4a5fa42177665069939f69e0bdcd9e2022bdfd4702a89bd6b133d239c0b403
zc893ed641bd6898eb4c8e6d860f267a6febb210604f85eac2997ffd8d05a74117fe3714d64e7a2
zc00b67bdcb5bfaaabf49ed4c22e40a2ef9d935acf6df32e50fa405359d62df524f494b007cd02a
ze6ea61385d094b034fc4cea8450e1bc35a2420ac6d133cf75b25a78ed8b83f065e73eb08480128
zdd16d30cf62ad6045b41f10688f5e7b7ef92c8aeeb77a41e8eebd77c7debeb6e94aa6a2195ffc5
zb45e8c2cf244bef37388aec246cbca5aa9606d1e51749948fcadd8ee6e44bbbe3df70809a00cfb
z8d1f8ebb83e9492e4cf876cd61a2cafe8816332f3e8ac1f396c771613b905b3e45161c185a2652
z1c383a56a44eb955119d86f26aedd43ed87c9e45b0a4077bc6dc8e9f07c384d069689cf25d9c0f
zedb897a011c1e5918a7f599bbfbfe8ea0922495296fa60b563bc26d20209d4914325a291135103
zd0160762a564ba6c077722e599502ced3c0958ccf96a199696644230891d116ac7c30430971c27
z8fb1d8ff0fdd9f7b15db75faa6fe945276791d3a1d4a2195e8ce588157c4c8cd80a575cba08ac9
z904b65d61acbeaa940915087293a753461c54bcb1653208e36e6071321d2d740b07324e4f0310b
z39c99f01956988f85ee7a720c858c95dec4b32b2cd219ebc02fa8e1f273a25c9730895b7ba4aa5
z1611b6db80fece00f72cbe1b1b2ec2987e519789b1002da50e4b42683393eb8516db0bc20173f6
za49a3956bcca4c3fb1f3e2da5b4e0e67c49b8c711eafa9e9f173bef4b769e861d170cf615a5530
z0c12f25a545f75907e3408d9d5a36814a59eee43cc03fc84de4cde36c081c5e802ea559add48eb
zbfee58574d1c5d4608159ffae2c728f9f8b7e4cccfb3b629ccee9ac2d66c2e98f6293a143db5a6
z13dbb25b789719cda2d6156e678b50dbef9d410476d70f2c5ab93e6f77aaa534c9ed2b5a4ccecd
z8142f7e9adea9a2673c42d7a15e75aa0ad0d140cf2da4652d334b12ffe8e9815ae29f4c6170907
z6daf47549eb08a1723861d811160b32b3716c17aeae3f7c4d3a6722e33f50032fb3dcc7f2b39cb
za1c6fcfa12cc20d589cb92d674082eca0bde3068486f9fc03b65a4c037aaa757619d4947a4144f
z2c6a82ac2b0c954d0dfbf702f2648039493b75fcc0e3f35e9fbe9eede0056f0f253b799ccc4c70
z13d3ba3ea4932c08d07bc86b88a2a222392e6ccd9d4053d2668fe9ef750a0c5537aedc2854ed2d
zb79f11dbe28e50ca82ac6da7c7d77bfbb3b536812a9a82b0a58d5bd0beb31c7d325edf470c23bf
ze194bed5b108aca768c23e073ca564c535d923afd0daaa10abca1d917da48eaac4e59d3774ed47
zbca9edf78658555d865461cc935f2ae6e60c2070de50e0a3f9d58bac962f63fb96bd848759b88f
ze3986aabc0a7a38e802fda8a190e31e49372dc7e53a35beb9749abfdcc982221e22f5960a41c87
z6015205dc5c4639a12c1ecf0485c20966f172f5c44591fccc311507871a010b03478e82e26fc1e
zcd516e169cf82f9f32c572297a17020e7a5c57e43d50511c419edeffc5643a427ad0f6efbdeede
zc76bda56d75d12f8cac8059f5a7fe1b68770f9e0a03c29fffab4d6aaa5936b4fca371fcf7cd5d9
zbe168ea695d5f201b1ee2a222a9516cd5c7eb74a5cb2e4f6dd26a72df2ce8d578b014f121daca1
z82d6d67dc6c5247679e9df1676eef6ca0385eae4497d76fbe2b9959ade44df1b458ead219ef1fe
zd32c6ea17f2d613a97db932a2c09766c65bf6db7de2bbf4e73d931a429e92ca6a91fdc0e6c83d7
z3251aaa8301e786b6fd3c457d7964fc48dd5ef312f06fe8274840941063f4522a1ebcbf772be91
z3390f539532236307bee4f229ab44b82159bd470207f34b73e94adc2a66ce5eb1a422e3c975873
zff4ac87c068848b9d7355fa4faedf921ec68661866e2f7231ff3b942e16b71facca8dbe50d1056
z773e705d9af06ba12e09d0340ea6044ff78d820c5b5fb4f517af8f4e6ed53cf69e2bd95c566ae7
z32d6be780e546b7a2f7a65d6527668731ab4e9d28facb8ec199767d325e23182e69c42dfe01979
zb5545941b8b7e8adb0858acdd9bbd3c30a0a7f32461a016cc2869e356e95ac4c8df89ac737c860
zde2234269d06bf6ca895a24fe8b75981e633dfd43757d0115b863d207328b39092738860345041
z434d21bb010492064546712ed777c25c6a9575779fe14edefa50e021c38df3d2a239be6f4f581d
z289e65b2cdadd26f1a3b8485d583bddfcbea9a2a1c35792741ebe494062543673768ce78cbe74f
z9f0f92b7dac1e14bbcb708bca626fa02a6bb5905209cddc16f3ef2901ecccb4526ca71f580ce97
zbdee345bd4a08fb317fe61ca79d0eb43623b1cae5a9837b9f3ede0382e7821dcab2b919ad911e1
z16f8fde84111c80970c75affa3fea11381ac3796cae00135be94d0ef6739a423e6c85261cd17e4
zb16046c942f140e42407aa2d5af987eb01862c02071d058164bc52001dd498b3a52d1889434005
z71ab6f8040c4519fcbf62dd59f59503b18d8c757ab0110e00e7a454fe218256e6e8374a2730723
za1264902b75a0299b5aa12dd90bbfff73e5aca7a326062e983fed840ba8e5a215441fd0a3e7f22
z1b1ac567097c103e9cac17a3914f1dd6d1e9962dbdf82c7d415ae251a19a6091bc4c288bdc9cb8
zc4944721cc739647e8ce884a1e8a9abbdbd74e1587c7ebf855e5fe187af94006e0093e59178d7c
z78a7cb2fd264b371c13aaf763927429cafa5ccce24b44d5c131912e2bf1a443555fef47d736082
zc5f1c576883baf4420f78593cc24bff93edcc4961ffb4941eabf7f23de34cf83ea5ec8a5bf0fae
z6631502fdc4245b8103a7064077dae22869cd83693483af27ee1c2962f2484f942bec135d75ef5
z910ca5ef106a3a20910dc3239f87cbf0a7e61aa6223658c1caf1beca99b36967e99b1f5f7370df
zd797ef7d65adba697de6e4369ad9dba0dc3b5719b41c509df5a048989f7d54dd9bab6c267af54c
zd59547bd7729d4202babc44ff2cc2776087d53e0ae878a1fab6cffd68cc4b750785bc25a677f36
zc7ef874b214d2917e9997dc80e90ac78bd862568c8b4198dc96adfc911dcdb5baad407b020fbc9
z1701159fcc1f96c6ae8c52c37ed9a53c2bfb2ae40be820d4404347e936ca808e859b5fe3298b43
z566447779fed3d9b7564d3776d7c74f73e3f9f3c513aeac20308a60ed62c1d4347840110858799
z12a3fd0135dd9b9e89274faeb7e6082652039a133d1601d2a0324fe9dc8ac902819f54cc2a0caf
z8b5475b21756284807ca27a727c8465a4cd719c1b6ad115316c28db69f001f7a95ef785f00542c
ze120f9fabf3e1a8abcd6ebfe6afce7d22ef8c33d242c6c52f8af884e5cfad2b19dee92bacbd905
zf0af731b3db4c8c55e96537044e1e2e5b770a0d7d7f1e9023c7fe449e7db1529a47cf3a41f8ffa
zf72510a56221fb7c1ed3ab18d8d954ed28b353bc406ff7466cb949b12d1d2dbd90be45d29d0af2
z5c2d08b44eb70a307eceace36f7385092bd008d9fa3e3be414576255411f6b668533cb1da54842
z652f60cbca49380490e1991dd21fb286c6a58f13c774598cf450f61e581e9955fac581a129c103
zc5202597fd8304e3fff9407128e1dc002ea1284c018dd859e322e2503f78684bece693957813be
zbf9e6f01cfc634219ba243e99f139aa83f03e68898678fd31b6cefbffa8bcf39f8f6c3e5229e92
zf140fc5cc9e515566d3a56f8ae3b31d03eb654d8ab5e5ee8455d48115f3a275a047dc5d8f22e6a
z3f6ae42e9dd6f0ea92bc2fc2b3b5206a5f124be1ce589e42d8f7e1f9e3fd5c726b68d6e4868fd2
z298445fc98fdbc19683874a1430d0f7a3fa32e85cfb27fa9c732a95b59e8d7af2a24f4f68cac01
z420e775cba9d8341c26d05ac637d8d61dcb820b0a1c2ee259a6c53dc65a300431c965731ec0676
zeac0272f6b03e95d34d00e8f1ef5a61c740cbc346e98b0bc929d21a2f30cc537ca884606b05e72
z7c062b79a1b545275b3a6987c75a0c0e78d64364dd518e652fc744802ff97811241920b523580f
z098ec226a73c5f56ac4ea8325c121a582d7dd479cf180140fc6e5f7829f624a8710b1318a04cd3
zfa0b588fa9daf8924d6a967dace7f579e3658aba5caa4be0e33b6e1dac552f2e651d67b13eb5c7
zbd737c8b3eb2f84aa0d6506b25955a387662600f01964f9cb1f47d5c48634e988a5a91227f5bbb
zdc6a7faf4b136841a806590eb4b8324dfe5353d9a5922214e6c3ed0dd427d1836c5ad740746f67
z246678a9457b1dc481651c9fd54528c272b588de49d382729b33e26adff61a19d2db84621a059d
za9765952b45b346a68229547e8b2db2b073762affb066c424374b0a8003b465aeef5fd6f16ce17
z4adbe0c40ab6fd453a5a0973217a69bcafe1498558f4301055ebd88ba38402d6e802d97d96ac5b
zbcf126a13de1a5dc4eddca2950cffcb391ebd3c16327375419b2fa9f77fd50a7c5ad192082acc8
z60953b2d6f6f555eb09788c772d3f302716f4f9b5de0b04e7234be146faf1a3aba97b1574ff73f
z0dd8b7295ff6316de53b9c7697647d87bdec0b7541565bae4ac330c0777e986949ff575410653d
z4984840cf67966403145a270c39d378e39c861231308446377f2b7de1e66e74a41c3fac07c5cee
zb35359f1e7f025667783b6db30f2eab294fece2dd3ee7b7241d883063f527bf72f948c5dd83b39
z3ba563a067b383667ceb2520d72fd28f6680d556b0ec62b777ce67f29ccb2af7a5e42fdb1891cd
z9ed83575a70de2a179874e155f1d9ee4ed71cc70a3efbf2614ee182a045132a7f764ed91d7f9c0
zbdd4c61c124f947fdb001f122bc42fdc1af931862d528a7a8a3b93078973963716ee94c431c38f
za83d6cb48d20d1b091e9d05ee1c1d85eb8d88fb04787d19566d3c4d5edc849c2acc6c203c084c7
z65ae62412b8ad777bfc5e616f92d18ab1e2a83d37b77cd07c0083929705118ad1b20f5a42198c8
z6d00d4b9d01ada53a12d9300c08c27f538e759540beb2cab069f7733113a1b5cf5c10315527f66
z7360d47c5656e1567020fa82c2a940f9e0a3eb420aa6aa30e8112d21202db9ee297442b117f149
zfae4c06ffaf90b593f0c6da80c51a272fef3d1524e45563b7399fbffb01906ba1c84391ba086c0
z48262cd769bba0f77fae9d31f43dad743377081eeb75cb78a0dc1ccc41f197e37def881eae6a28
z4f508c7ee916e2b31303567f95a6d266982d59fdf4e5379d2dc363fb41ac6e830a22de31292771
z61e140857c65883e15dc4d379132248d6cebd7e88851868b94b3530e4efb33845a48bba1abd0e8
z9ea4f48daf939aeb874c993c72e772874c1ebb9942e4adf98cde6015dffbac7985dfd8de391804
z9ea02dd4e36aca55be168b4b5a3a8044152eaac39e2b21f68e9b39aeda38588d6e367c753e0504
ze83f3c3e5ab1bd8cb832ef6736b67cc624c0b0e5443fe59692f8b4f174a430ee3da6255780152e
z75f1035e668930e7b7fdceae4df640c11ce89c3de5ac9a104131b457f181be4b8d1a34eda4c9fc
ze25b57131b6afa67ffdd59fabcedc059d310fbfa1bd14e3f318f721cbe20d09341b8a88da9710b
z884fe37611f4622caac74c756eabb77634d60d11351c56bbbb0b3158d80c011007d4457f5801f8
z468b77db4f773f56f2d8bb007c2b511ebe516f16085bb73e36e46d0d496408caddb3cea9a6e160
zdfdd8c72d82bebb82c13277424c44e41f3f4d29a8c8b2515baf8cde3bbe1f0a1bd662b593b0850
zb70b9a19f5d2e3785b39aa413d3f87df428c5c4018a3e0ba6522a1ffda57f8eb4c40d295363fc3
zd5d35398435590552c601d4b59900fc2d4c6bb4de4c33946b0366196630beff9f5ec8f1901f133
zdbef37a43ddd27738b84faa81b674aef0dd139f721fee3c732dce0ae6fcf564c3b65fe8dcbbcfb
z001a9a2201cc1788be032dbee4ea1f1c95fa2b6f9164f48389452500118d462bf4370cc140ac93
z397577ee3027bfb165cd6947da8833bc6c9806de88163c05f9fedcfa5e336a171a50d888f03c7f
zd6e28fa3cadb109d4fd1044c9e1e9332396cb90bf51c9ab46f853f77c61a78c492df56903c75b1
z89895d75e6abdbf3551543cf9d58a70abae14970ac0245aa4e94fe37d771fb562fd6cb47f37c75
z2126be99a200498e5cb1de1e8dbfa5b86549eaab355bbd5b74e6382d5dbbad2fcb282ab66b90db
z26060127f7d269eef933c68cc4c767168d9e92e98937086669fcefa87ffa7e509656131188f95a
zc3322df4bd2494b7939d7ee0310448224dd4141379988d92153949c4966eef4b9fef5d395b1ec4
z6a09b54ef56bce2118dce5f8bed7b6971a462e3873aeaa20f95bca27caf8460d55a7c87a8a18e0
zd8fa45d01447ab39176c061314843974c4bd26e4c08bd783ca61f99f270c7d3f10c1b3a7b523b6
zb7fc647c6f159795658a2d958307dc83a611cda0ac0381d4cb7601ef89904093f736ab22067726
z7b4c3c99dc695f1831cf5aca41ecbca0b787ebc5b2f54889e6a0847ba607ca81ac0b9544461e6e
z23d0df43d6f9cba65cfffe74de5f1160ec41977940083598593914577b303b3dfa3a54f6af37fd
z2839e47e01bc1462378874a8578e015c08260a3cf5289fec8813bfef13c8619ec44c18fbe37ab4
z86a4e8025693225c9dc35daa972cf3f525b3cf1a9f053261667d9bbf6e10e4b515234ff9e0b029
z70d0a0199ba9335fa97fcc4d06907a6a852a91f704f2469f97cf22b32ac9459d28a4564d1deaa2
zbf766ae7d4b7d46b7bbd2c430a9d7e02bc167998b2082b45d26c999d55bf0c52cf973924fa86dd
z8977d271f98d99aa183007faf7919b06d92e1f8080bc55b596fe538470a9fce32d572d329591d7
z6d7d00dfe01deb2b918d655e3a12bb3729d61937ec54d3242d6c4b83e514b842d1335f80a9aa9a
zeb5d1ece46c4b26b6b49aa08627f8a99a8fa2b9cde19fc558feaffd52a7f09125cdb6d88b38bc0
z73562981bf62948cab0c0f52dccacfb1dec012c4873f3baa351b3a09cdcada760c9ed56c8e9aba
z0db5748397682fa715cf5d0cf0cc76f45a808167f49d7973e43d9ccae0024e74378ecadafd71d3
zcbe188a762c4ab824007fd34bd453c1b021d2c3255983aba0b3ef1a5b1e0e641b992ed39d7382f
z38a2242c1d42141f33aedc2d6025ed8d90ad05a6322ce827a10df50e5c7c6da2f3c57d85449e69
z6f21c67fa1bd2983e0f6def4de079931c7a1a5119c65a4bc99de5d5f93539ae9c51bea4ebf4968
z898786d5dc9a73bbe10d81c4f1a902f7c2b4ecd8230384f91253aa2a4f149aeab8b28212dcad88
zfe2029da6073de2e03c901d566ac4117a7b92c06943e446240a6233bdb29262ffd333e7b4b4b8a
zeec865f735f0fcc9dbc0ef23cabcf9ca5929734f8e1d1ddf0c2148e6c1889772add6625e7f495e
zcfa7a7872fd8f967777ff2dac1c514679b0cb41d99d18b55805a6c8571972dcbbe3347a935c6b6
zf7ae48758e421bb0c3a15456e10f3845eed42d0de5a034ced6621b3786c91af09942ff9809e465
z171bbc219984ca88e23581179f2761e46cf356d55fbb9181d791060311d57ce9a07c163e4ca488
z553311058aa6941cabce2faa08dcc4e2907489421f146d53b97ae42562f7e5cd18eb353c5759b0
za4420b94fc57325c38c1238ae4896e30805a77c55f01354cc3a163e5ee259d50315fc0fda53d0f
z961386126551b04110038cd65793c0bb98a234e78bd4c6cecf4b8bf5dde293a591e43a3d98ef56
z13b4275732f642ea1677568b2b536aa3424f20c6b4528274dd1945967d475c98197382c8cb2ea6
z6fa12ba4366ee1abbb59ebb96edd14500711388393f4c600f901ed8e718e3aabbd4cb3129a59a4
z9fb3d8d47270b1c69488eb9d70cd0d144105dad72d28baf19441469fd8d3db5efc109e4aaab3e0
zdbc666d9e104b3546def3cbbd6a8b09270a8d7b682de64e65bf22c9680002cec4f794b4369a93f
zf81a015ff75dcf8973877c7363bc43655ad15a9e6af3f31a77d9e62afdefaac261fc1f50cdede4
z76f1c112155b61c8c6ab41fb7bfc7e9885a68f7a08f3f41ecb449e8e9d872a983e1a7dbfd3944e
z2dd77b4ca46e0fb3e2313460b88e4d8089e583b373332eb3831ee3f6fa9c694e0da14ad8583411
zea4f30b9102a0ebf13102e0c22f6a9a3ddea56ea2e4d8b3daf91179961238b47622eb8394b6df4
zfc82d9fb4f8a4f4336edc232156d94293b5dc031c45f3340376d91a37fe45090bc0bed6498e7d6
ze81cca25a054bad3eaeb6959eb1a80da680c1ddd53fef450720309f0bef973c4c97ca01c6e7873
zb05afd0fabc53cfbaffc88338ef5c8f85d18a05f6295b576254952c58713b8ba75d6e3f6fcd0a6
z10d75182a00f0a493f32b5dede8c356ea2c8fc07e6890518434e45067d27a0db6a7c2512b2a775
z80ce2e3801ed3ce5f8b8fedf3c51150bd6389eb8edb710c06a5a4b34c23435602da00c00157819
ze7758fe3d97d0678c014e594e664656e034e909e3b827972cc5f8f71f6d09acfe4c9d8cf678044
z2f25b8333eaaf0d47ea0ef839dce6974b24bf6dae8944fe620cc4f1fcd3c37c5d06484abc3a787
z5f1fb251458fa24eb765c9990c21f5f108563999757bafd2eb6750ce19594deb0336e2b15e0e6a
z39d0b4d0a43e90f1e573510aed4b4871854ba11a4f785a3275278df61ca838c4195d1baafb2523
z259db8452678aadc5233c8701d356c5360ffe29cb4d597293b66437a35fb19cbc05fea136fce0f
z682f88a316720611eda47f19b128fd90b4bf471310f303ef8a4349004b129f7b73e2ce712a33d5
z5ccaae83497359e98b7be5169a7c93611908c3749706ae22c918378432505c1cc12fe6c753d5cb
z83d7842b16749798e0ea4ac19e3ce2f679834f479f56cd2dacf924693d7b7820f18503f13e6d81
zf30925fa9fa1e9fecee06a7a959e85ff52e3e39412e8fcc46c40c312056e018424c819be4bfa94
z922000637e1899f39de854d75f3081d07344b20c41084534aa9a2a94eabcd7805e7e2cdda842c7
z4b23a063c1335ffa4541f1a0fe8e8072beee5c1c4cc5df752a92df81bb06ed8481161193dbc0a1
zc68d4bba22343a8391f210a65bd1848d8ad058278e22b68bac8b3d2fba0477b3655ae0449a6d14
z9c651b763a994fc993f058467bb342c1c55f0789f24c8b909289b8afa520afd936ef163130ee02
z5010cc5ba39711b2335c6a8934c8bf05b6c6188ffdeb1c76b963d58afcbd8b1ef3179ed6f7c0da
zca614737429560da54ba15786ebdde371a40d772cc8778bf3e90c4eb837825b5b04cd2740c3350
z45ec19dcc10793603a652cacfd30f78ec6832eff6b0ae87b6d4a40e0bb4c303bd4db82fddb81b2
zeeaa6814703d0dbfee0544b954dbb7d3d529d5553660f68cc99136fab91622a57e0e5d8e71ebf5
z300f954d690e26c5ab544d02746bc63645d97f10153ab3b8d0a1cdb92cf56fcfd66812404922ae
z9287224578fbf5f488203781f5078c07d0d084da1730865bea218480177930d4c3d137e55ad668
z9f09fdd339738057473c78f945256dd5c53a7f9ea71ab36b30415ad88ac66c39ef9edbe2ac12d0
z4aa8efac557a1e4e0d8cca7083a823fb7e25d085369d1fe6e4adbb7388cd05ab216c93d35a541f
zcaaa3740daf4936943a759fe43beef401b758db35f62b4017086c9d5546b94571321e10ddd04f3
z92eb7c7e18e05fbd19a822439bd71f9752f88a63c62695fbc68680ad91b6410dc4c9c82d274a9e
z087f275c06ecc7dd37cd89f3420dc50f4efcd760748249072d2310ee037ade2856e9ec080b4583
z01ec855ca5b20fcec99fa7bf05ec7255ac01f38c3cd4674411880f62e11d0e89380ffc7d06fc07
z9bb9b36de0cd718f548a9b309c8deb4b499010716442402001d73daafe34330d962869b8f1d816
z8ad8e54e4f15429bf353c0eb89e58d3bd9415c4293a035ab1f15187f250b7e10bb3a06f748044f
z3ba8a5709c4c1261f0b3fa36e01fd41c838771c21f89aa790694ea1160a6b7434ffb34b11a6944
z16557b6c78b63672ee0fa8304a66a16cf78987cea9f3748f593fd1ec2dfc421fb8ac6ba5affa32
z1c2add274b2fcfa659a982db508620b2ea4f64961ca7f7fd3b7b6a327ae32377364abc679bfedb
zf7e71b648ea67bfc90d477b87b2f15f40341c9e02e893c6fb793dbfa704ffec674ab2254331c04
zaa26d888b41e601566102f048f1b4d4fbf5002270916b5ab2fcdf1fe8ac82b825d6b3e35394335
zaaab6d98a1b3a31bf718bc0fc716027655324f9f9fca8e43db3f095f60b3beea5a143167100398
z01614e0ee4f6498f6be6549051f4eb7d8f55b076ca0ae66cc9cb6448727297cb84e452872c4fbd
z20954ea4bfa3c3cb52d6e6bf1c4a5093a9e0e42ba9d0e540984d7d2aa12bebc810d1d785a9fe25
zda3f0739ad7d27f0589597256530d1c2651b025f78fb852f00551e54234bfe3a99afe739aa2e7b
z3a729459f093070f9fa2d40d4b5901b3ac8e8c6dd237b69cd0bafc4102e57327199582e678b1bd
zf670897c306fa1e90ae3d5ecf7819535a017c0a08c9ffa2a6f1b84d6196243650667df735eff9d
z226dde205e42ffed3e8750eee15818fb4f4e5587282be75ec4d24d835187e5ebf26942a81594e8
z33577fdd0c72575debc1019bf43d53c433ee0d17fbb7c5aee2ef50edb1867f448c75a2ce94df61
zfb9ed2fbe43083c05dc8ccffd6efbde0fb71246b999f989a7bb0905255cf848eedd58e1acd78b5
z08d01cbab5a4a17a86488ee07ed62bcc4bccfbaf8ffcadcf86eeb9a7392b19a697c13842c23591
zb2094a7f0c39a5f7460a6e7b511bc39942df5a10d68176f9f6ca0dc1565dff0e02ad22ff5339f4
z8c3c31984520fbd8716abf6fce32e157dc4cdc13891ad8438071d9a0bc4516a9d622c7ab2774c5
z3b01a393a013aef61ca7cd9a40d53f6845079ad28e2eb84256f8dad9aa020835c5516976610857
zd8c843d5e297ed1a006be04f24fdfac5573d9b8fff515f1d28521892a247d700c5382bdb760548
zc66667720b541111e40d1941fa80fad81f9b4241dfc325c4b8c859db2e648ce802112e1a7f625e
z48a527f3a67aefca65d00e7083e7899594b80f96443d96a8b976160e1f62d2a550316c4eae2e07
z0613c527ed9b126a41b96b8403197c65529864d8f411c78dff533024fb721812a175d45a825fb5
ze58fc436f67db22985af032ce6e14651dfa064671aa5a5ad251c13af4e3ab21eaf3f471984c801
zb5ad8e7722c4ef17872a828ea8f42a9132331cc454eb2aea310c4f0fabc1730452154477fc28af
z6ceb983397f037b0be2200af200d2f558c1335be11a090ef84ef05e0c29969d91fb42ebec87596
zf28c78a6b485d90f7013347c4be42e4e45623dfe7fa5b0db6822e37691921538ac768659366ef2
z09f750f37de8cdda777cb80fc1468561934643f541a659b95938f843dd043212062c2e50315167
zbb27d8d3d7580cbf80797e4895a53a993721a161140980cefb329d83c1512c7f8d3b8f6611a202
z673054d72badafa117d4dfe60dae9d4d60ae6061b53c093ef5bceb0f7f360f08277a9d4dcc4dcf
z0b5ca83e7aad360a65b057bdee64fbd5b3cb0c7064647f27ec296183781e8e6fe03219b106be99
z2cc7bb4f470bc198fbc3d62aea63fbf9e4a7fd69cb4627b3e1cbfa7f127ae72623d7e10ab6464e
zd01ce627f2a9b0a404515058a6d30946044f9b3c89006f60b8b9d4d5ebc713ee02fb01eebb8f4c
z5e99402c39bd9aeb7baf17712bc395f08d46ec47aa274cc4e626421102fa8ed26005dc185a313b
zf7e7bf7536b137f911ec0dec07ac20565160d0c548a14c631aa2f81e4c445f4add8662d21cc27c
z1d4eacd38bc956fe2e8a8ab7495907454a67c8ef260dc42723eb7313f77ed984f1787b2a496dc3
z9d47171236cb5cedcba49ae92179aa4451d2fa8a98aa7c488b3e9976973c27ed16b520218f327f
zfb6efe039a75b02e33583d6ec1f9604efc1b8ae01a27875d3e748920aeff4fdf549e3872ff266f
zc16a5f65c790d98761f71fd8207870a7a2ce6f6cc4bd3cf170955b6a4d765dd723860b3e7645b6
z27a5c3821ed512a65835543a368b612cbd49a5238b7077a076b1e9dd4ef982eabcf7e3eb146a99
z6a08657f1d95cc4869ef84342533c5557e9c65167ad6510e7c292717b89f6a471f864e92581e7c
z3bb1ba8770c7db735d28a43e102dbec5d2f4570a972eb166e23ddf960fc6b51abb788defc058ce
zc61ba4fcd1119d2f6e3949a21fbfd61508ae28462fef38d14fe37f401883193bce3c0db7922b16
z39a6b44078f39afd6aec7c0e09a3212a69cb441b1dfe1b8a9866c48a905758950271034d465795
z76281d107e05c908a234d4d2c09ff3d770c4bcf82d852c2ac02f9b6441d2953a4f356d056805f1
z0fc68fa8b20292a2078c948163c8c07d9fe1e4e671146408b31b17c729136cc9adc808728e8aaa
z207eb0c7f53bf71170db44935df3fa09da115dada0e5fffdc625cf5991ab6aeb562fc473b73c80
z14fe87c3e320b0827f37e29a1ae4e32d28becb28cf995ee8ae5b136398bf3c3e76ca957eb45fd6
z63b04cc96e353af53382d1ea527a264da33e6d6b459af9da0c0862bc7950e9bfadcd863a009536
z346c6ff905e9eda5e975c8da86a6e3af0c05e2fcfa9c5e741c211ca6fa00bdf205bc0d42f769e3
z20b83baf8a2eebeb132212c30f2164e3d17fb4c76d715bb1ed252517a742b8fd70a6f5bb4dce9f
zaf5d2e84530167c08af6f52291a1363e36272bb3a85e1ee34d13b4750571b31628b72ff630609b
ze002748801899d55031b8a08d40c24169cbf7d11498f406f41da669a94959cdc16f2cb02d5c3be
zffe90c112d2b2550a1d6e5a96862e512ec4adc2b0aea3c2cf056057a45b68f54f70c0a8ec5aacc
zc1d01c1e4a9231e8c503d6e54da3d014e1e34f733f4a98b739e1320a21bd159a74a5ceb0e1e602
zb7205e31fc0ac92745c8b43b20a63d8a55d243b1dfa9ab09c575047c10a297ad8e46602675717d
za13449c89f5850be6ed8e74f749eea156e0b7a79e06ee57b04371b77813b2cd0f5e21f5fd869be
z93d8b4432344ea44e2071cbf359eda5a957cf654735b898cdc02b9b0d3a4dcda7964d9914c7379
z1c419fcc33db7421f1c9a55af082878757ca84905bc3a4ba6083443c78580cd7c1088161054394
z2a94962d81baf5924843d4f635358cb153bb96a24d456f7b089f65ac61d8be79fefcad19e831a8
z60254798f9adf7f784e7359fd6d485b90946c1c44597e15cde513390f9ac41baaa4c66de7464c1
z404528521d1c4f722ad00296b84589bf07f4ee8bcc967967051b0728fbf1f100f24e1c91c867c9
z881f5bf5c35775565d2597f467cd3ecdfd31f78e1cccbcb7248e9a408b0faea0be37acb7abf982
zea1326794e26e76bca67b0adfd1a31ebe4898d6a11f9952419d33a0838b1921e3a365f003e2611
z624faae185a75c0b24ede1426e61afe8f0bcb005f2e6762d946f1629db6bca4e8228aefca7e078
zefce835e528800ad382f1d475c220ae95467d26a8cdafab2e66ba7d3ef2f553f2f093422c67e92
z2ff972ec0605b7387a2866b2b17e83a84d2b0ae82dd0aa51e578167f4e688cf045ed5f49bbee17
z7923e7ab87e8e2839909a8bf4d27b12c6c6a483189a461047d1bbeb290edb5a3ae557181534b3d
zfe4875f7f8b66159092c57cdfcf8926f2584b4c3e167f0c72e6e5addedc0631f2b924e3e5236f2
z50109e5eaab549ac0201a122f73c3105a08006f1dd386726d0ecf8cb8d889576f3691028134f96
z1f1b70c41cb4861104f16043098519bd225b0923eb507f640c39aa8a15006b4b95ce4da033fa2a
zfe2b12904d969079c63d57dfa6a1d7c3d51a2516b3a9cffa8aee5e13403c6235c7ccb7564c74b5
z91b227d4e7ffcc386ade931349a7dc61203653017761a2821a8cb3c2ac2633919ad9fd635cae08
z18378ceb1dee21bea9a373869a9aa6bae512d15cedcc2656c12903c209d5c6b208e487f9ff0267
zc69e54b56e5a5993a3dbf0f5a7ffa279ad200224a81da00e7f85f2c6861d3194b39895d111f408
z4ae9ea4b899fed42c4e94b257442f9ccfa9ea919a501a60e8ab6ba8f943c5be1c5153990a41b5e
z9a531691827ebe187e4e42c31ff31507d6abaa862d603e2bbddb54036564eccfeab16cf9ecd0a2
zb9a8b282d281bdd32c36bda5143a3d94e6f703bc077684715596d33d731d447972caa28a7f6955
z688fe423afd32dadd6984ed9695660ad7fd3293d9d9e8e6893dda2ee94a427054d66b387ad06b4
z71d80be2f3e4ab224f99e03b8da31b68a876b41e4854e516478f3a7c3067e6408f8fdb05c5d778
z826e02c01df0a3697d62b0f4130c792a52847f83b4fb6d51ec9e6390f22d47791225b344c40980
zcd2e54a7330c4dace0fbbdfd0b5a4f562af3319a82dc2ed3a83f040fb31a9bf7d86923472a095c
z91201798f9e72a33498517b8c7d12cdc763bd8e3fbaa7494fbd1d6cf6d116c24d605f1a1f45d6c
z7cffbf89b7d7ba45c45b72c31398c820f9b90dc20795e2dc877603f8843d3354eaf4545c8d3d53
zdf3b1365914070e9403a5a6c1e03206a67c240a7079cdddfcf5bbde2f7b86d6893265e64aeb35e
z2251108d9b3f60b87c7073823fb3a55bd4f56e4dccc79eb9517e3846045b4e7ed68100b85904c0
zec3ff925f0ed091fe68c1036416c4d6b8e8eea9fe402fa3743da3c92734422cee6349bc01a9752
z6eccf6707b64bc4d7b8c665f14c7faa373797603f829d5ff68f82bbde1e6f2ec0ce43713029267
zb4c6698814d41d8b85797d04e0d910a2a4fbca616b17e3037e5887f4c0e220941dcdad74c8ab8a
z68a9b5ff244cf59cb2bfb584cc111fa600ae53cde1c5ac49aea4fe345f874331bfca3ca7f68326
zbada9c508c82b4fada700dc8928d9e6928c198d27f128f8ad5f24b9fc1d54780aea7ff995e15f1
z625a4eff22d53cdd84e1c24846a7227c654cf6e6ac358578633905036f78b515b6b6fc6d0dbbc1
ze8ebead8e41a19cab58f25826c9045c9b064cbd8f3b29bf77c68d48a7e4eae339a3bef570cd2dc
zb54ad559bd219674b52f6cdb8adf577723a8920f0c42d3bbc664d2d690be43cbb6b95a1a54a999
zb9f17f48bc2b1b31585dd3c97b056ddea80e5180dc48fcd8ac8d780a1665aa362e00ed7d5a9c3f
z9612cb1831b1238b37a9e9f97495a18402e187018dbda35a7b59db8402f44d4276fe4169ed93f8
z03e85d415a0fa2969e0ded197345d488d11f6760647dc60c5318ae0e95177cf97469c821b24275
z495c9b71fde7bcbdf5fbfa1d82e599935a515242abcb841108cfe8412797d05c24eee48d4d0bd5
z7c94a836a34bfd8add5b548f974bb61ba498b846bb799c78f1697e49614116a4a8fb12a458ddea
zefc3371df5604e246542d95f306221cb75471ce92e23cc2a771bd9dc968c081876382949c5b6eb
z132a141f4e24b14282b55f2f4e8832a5c7e4571fefeb639adf2de39a6929075d2bfff51c5cc3e6
z50ef812770b975b9943d80dccf283d833dd34799682a6af586cac6b015b413b4c3ae1a09d1458c
z8d29de8abf1403b89256ea09b04598b93eefe8147b276206edf019504bd7d16a4d3d333e1336d2
z5b14a661a55f16c50b47751e5f7470230117c015195fdb3fad2afce312ddc893af6b7d6308003b
z6fbd379c141fb84b8295fd104bf89f77a4ed845c17c326c4686f8cd6786d583fd764f95d8b2cd1
z2e2380d43028117225fceba42dbd7d9a7392ed4b45fa685094ad8237c627695dbf9f311e9bcc37
ze0660d2ab3c11bfbe35e5f171edc21fd06551e2b8660dddba94067b4c21359819f468e3c62ab48
z4cde724e10008b1c3f559ae22c76948ae7ea952433ba8c1041c02d4d859401676d08079b111ff1
z1d5846795bbb2f2b9664b2b5550279d0f7b386baf91ce1ef1a4173f7ea163c758eab0c54d92925
z26a1ca8f248312f36ea77c3617b28aced58e3bc44d50752f7fa018d6a62b6fea7d8bbdf41841b4
z118fbc86b34a64c06124c0940e0af35aba05fa98401b80be92b8877dd5885c8fdb6a2fe21f7413
z4157b790e4a86eb9ef794af2983300ed9d7310706c71060f3141309ade4008e889e659b5097517
z885a7fe8b84e8fe14f43b6633b5534b36761e95bd48acaea05f45e069c693f6fd188620464ead4
z4f3cf67a6459c63a287069e09ef1366ec79bcb795e8e05ac9ac9c20f0cb6f55ad18f212db5b0b3
z98f136ee6b251df0e2fcdbb1c775d24bb7dc690a4bad0da60f620aa597fdc52387444c2753adfb
z26ee63727c055ace949e96c30570e8f809338e303437c3dc37fd9eef6e5c8c912cca7c8439d33e
zbd90b3a14f7ca547259799f6f8727454a6dec1334edcf10a94cd36adae75d94e33734e67a0c319
z494988257ec5829934e5b1e330f3a8da32dad501b34484cd9d2d57fe65b10cfefbfecc9e7313d8
z05232317bd73ad5cf797940feb523e6da08aa8d9f118ce419acf275715f827d4fcd1a22b81fad9
z29b3e0094fa9c1a743ffb5e5789e3d008c789e068e58d0ba29ed31906bdd021522dffa0afc0c5b
zc41c32c61e2a225635a84b88e9a6552c18a032969fbd1ad48adc0c03c07a4cad03e84caf464fa7
zb1b889d6599e4fa7cc7a33297723fcdc3866c1953374d2cdf5afc2d7989ba96147565c1d53cac6
zaae870f7bcdc5fd847f0d9742e219f7dad9934fe39264160e4b1da420e7ad72b56bb0d95e9bdef
z55111c94c81da5e4d103240600f73abb8118d889a7f3c95f8e13fc4d1efa95cc0d7faecdb58f22
zf97fe92dd0e6151a28c0ad266b3f2649f6d599c899608d1732223f40d40ee49c91ea7d6d103430
z2fe0ff6d3fe0be7aa7d74dddb2ae34cfde719dd576714908b060835cbeddad9585049eae695837
ze1819551780ef7a6c3909018fd5ca24fdfaafd88b08279dbd27dd839ae1a085e061c2afb9e192c
z21cbe2b85ae7b079d5f6d6562274e14e3c556bf52c2af7315efe9f9f796f7828bb2efee1669077
zf3a53ffd6608759dda199a6a0f5f30d477307a0805c0b7ec7f826e71a493a1960ffd75a6f037c4
za6d758387bbe2f12cdacf2c3f8f846ba81d8df07a4f35f939ca1c7e035f995b200b203919b150d
z87e9f5c2dfb09b5d4eaf2cd24286e906c123a7aa9fd38f49863d76c2abd5a4f0662ffae6c43e70
z37251fb6113930bfb6fca1570d2c81e3b090f0e6277a11fe0bddde019b81d1399e990d087eaa5c
z8d0a555043b521b2864eaca224ce01fac05dc1c15b7f054ed4f1ecb3f44a454805df24e24fa282
z5b444e3ed816341493a0516b5fcab299bf8315eed285fd14a27cac392d40a03cf270986e46c92a
z9fcd7e360dccf07244bf2084e4c9b03e7912c41b14397ec98832b8d718304ff8400ee29ee7c417
zcc7d630af71199ded6f6fd6bce9ba653562f920a622e9b4666a01af38023c97c2b803754798e0f
z08ef758c94d2825a11d4b325501d292a5397e07d4ad200de84bdbf7f4e5eede83fff792f802a48
z7cb69e63aaf7a245585424d44c5415618ce4fa4efa3047a4d865c4c2f4b7a718483b963f1be297
zc84b683420bed86da7f407dfcf6a2e6a1ed15730430f25ca8ae25bd32cb53a8c7d9b12c0e28367
z14f43c3e68f0bb546fed5a538b7fd666f76138cf96e2f8e545f3e49655b33da9bb7b749164dd21
zc43a862f8bfefe2fb5617d27334a41f5f8c48d5c28b46d0afc068eea5c85bc8be611c7eec80bb3
za599dc5e3cd9021a807eb59d9f01e497c5c53b09fbcdd7d5f924fc368a3191441745fe9779ca25
z33286d590fd3cd839c79c3dbcb6525461dd28736b3edb9b5314c0abd9abbc8d396b97751995ef0
z6892f8361a812571a4a5a575ebea553b266d5f973f06d2af77ef6d92a1f1cc31058ea1b47aac31
z95bdd6b54eead84f91231f661bec839a4a2749f3233f4215e8346b47069b763fd092867875e587
zde2c5731724b5186433c6143f591e4781b7eb3dff17162a69175ce0e391ad856020c02f3ab539c
zdbfc2384c652239e80a0bcdfaa24f14b3707d35afc709bbbd990ec27a1d83e66c39008f7cbc59c
z95ef0b554fa444128e6b16ec1786855ecd03c4d088257b02d53cc15bbd2961caa4eef3cac83367
z46f0c4cc34378191cfcdcd545a1ef90c3336a8310466ca4d78834ddfd23812e21e170be113d152
z8d4932ffd835528b7c978f48891907cc227037e8cec3da945a103ac21482c4e90e6e1517590f00
z3a16bb9ca9f1df731c29117a2a2c54fcdd423c0afffb810b2eadcc948e7c1a2f13b5eb7092991a
zb18baed4714e9cde236399b74bdeddc525fa36bfab2bfb267772b38db9e276b5b809a7e22d59c3
z811bcfeb5a754fc00fddf802d1504777bec596ee9b440a0b6d433151d0deebdc2611141632bb8c
z18d576a2e2a150972d25d34b7bf47f0124d6934a4ec5a5e99bd60f6fa790c3ed6220cc533a19f2
zef588e5ffd2458bbf6bc50e59e8db25950cfe1902d081d73b579fdca08b3fb6f9c0836d758d36f
ze27d732122c1abd60ccaf9acfcfdeb76d29629e35432f276e90db4e479e275ec8655555e46d9fa
z76d5dfee0bb618b77bbecb2517167e42da5a4a39f1cb3696e3101ce3650f0cbaaa35051197c23e
z92b5c6d22b79572d7284450e2e7b0eaa83dfa943786c22c19c89525c839e33d1416e9e884364e9
zd88a00946a138ddfc422fef1a0d351d407b2d515ed210cf1f05c1984e095bd99ab52e0cad69516
z5de5d66ce3b291029b3575b389c01f11244d20703b8c089ed14894bd0d2fb0a8b50563de0919c4
zf6a01765117fd861250d04d27a986b690e1c9695c078311b41dce9fa8b8101bdb579a5ae817a12
z001aef70d70178e017fb7eeec5afcd15782dd398a32cb11b6d9b33a9f42af968f8ee193017dd47
zfdb8047f2f68e066ae00618ae593c289efe80cca752c80880de3b068a8320bc8e79ecf085ea50d
z7fc83518ffc9c451263fdc9b510f33e76a23d1d76bc4847e0d9c4432dc571fe3d9e3ddedd1bddf
zd0f61d88782020f48049c973c737e84b760ba3ac0c1a4673355d1cec927c7b6350752eeede2d70
z9f241c60533f1428602399b5c1ea4785a0d58fe003fcc95194ffea7abdb4612072325e95cff0ab
z7eb7d875c710f1ba0733d5d3cbf7c427979c09c834c4de9ec8ac87c686d202d3af0d490c7d33de
zf0d206e7de5d4940c9bf07de2f55a353574bf240f1a9d5ea137d220b86f81705ecd2f438e90cf4
z94e4da9be50467046cc37cb83f611a7350510d342e5c7a979b91ae5d36c6f12be02d11440bffaa
z0abc63223dc2604f188fbdd5d681525b4e4a4d6a4364ca5684c41eafc0ec4b232558287c5db17d
zc3a299b95a9b406212ff39420a8a708b950683f5b6790ff341307e82f818931748e8ba936ab23a
z55179f307f103deb0eea98e99d1581ff3af9b4e0b41481888717bcc85c8191ff2cf1369b4b9d70
zb995335f701f3af33c74978074a72c262cf00c616cf981dc227b1f62ea584488e2656fa3f00afa
z5477ee46d2bb56736779499f34eb9a8ec1e53fc1e242e46d17e9309cc19c166132175c6abab817
zfec775f0b04a949bbef6a094b923902e94d0dd6d3dda60d0b545f3bd78f60e46fcda285044d4db
z0e9275adb716f398b6b59b2b82e0c99262056a65591a07b11d792cdc3153481e062c305eeb64b0
zdd841e58b9543792785353bbaa2758149f1b2fc5fb7ad8d8c43048e09a4540bfdc9948ab8559f3
z24904cd7da5eccc983a28288d64d907cacfe589063ce125f9c48140a1ae581fb9d1e1898bfb574
zd644d7387ae277250892f4084167d380f0bd533b5a273413cb9cbd5bf8387c9c71d8cd4df954db
ze93461d8e25fe245455dd32bc070b3ca65109dce6fa9dd4450b844a3b8e67b6b1681aa73a96cf6
z398d2920fbbfe6b6d92859dbeb79efee2868afccf5a6cff538a1fdfa3ef265b7387cfaaff26378
z6e060e85a2a83345a236e73f160643108c140c4e80bddec980550b0219804caf65c4729b820283
zded143facad8805cd744895f1ce42e7fc3933d80d8d47857f6caa1f63eeea1f162bde66d08b867
z422fefd1e49bd6c360d7864749153005bfe59dec2bb788e43fd1d7ec1324939781ce0e7cef33b6
zb76206637f768aa0d5228b8b34c9e861611d473371cd3a868148eb36ce458bd0f928d9b05c5f96
zc7d5797b79ed83f6781f0bc00d115b5b5892c828ef238d67f956ee46140c8dd553f5c19eaba7ca
z7a2fe0a87a1d7c4296e4a7d7712d2ffd72501e6e192e7e15cf9d06dc03f840db23b3998895c3b6
z7d7c043ef6f38662b00249fe1127d9e2675dd673e3b309cd48fad51c699f552094db664c125f50
z5e2ebf3453c6f17b7792723a6a9b21fc92197dccf3f58fc4f18ed6725bc118adfb8d3522903c20
z41aae394f5d0ceb9433d64ede321303371602739e3d62cdd478d4e568e78a841ad593dc72d3f55
z455ec8f2db92120e75578e622d3e964a0ef16cca501fa68a5f781963fd09fcb21555d7a757675c
z811921b94259db8eb68d166d68e84d681d49f3034e599fb73efe1bc3dcedac16489685a97a532b
zf9db5d3035d8caadb8824deb351359df6d133c07ea50d951545c16521f5068e2dbaaacfffbf27a
zd2a4dba892fd1ce6f76df87d93d365f3029fefcbc5045d0532d3c5fa893f7004c5b5f34660cdeb
z3b3301a96c9bd6ce7cb69275f54855559dd31bc025a553815ec9e61777d68ce741b3e87d6321b5
z64af6d6b7dca209c42bbe7a313c1d143f90cdde8f1b26d00ef2b55000a1d4a9acabce7fbe57873
z0407cf4b207948cd6486cf8fa6ddbecda25a56a539804c93cc4bd61270444bdfccc4154c2b5fa7
z9e688d84da258d0dc0bc083c647f56a572c7bc70df84df0f4ae85e79361ca9db29c9de4f9c913d
z40e24e9430598cf64c928009808c4a9742a09da8a6d5a335e1972d9bf26a0baaee22375680321c
zbd6be2b50be101d46addbe65ea18db6a47ae4cf48ecaf13318de3f66b9e46a4d8ad3ffde4036e1
zf384e4babd6910e1606a07412d8c0d0997caf0b62dedecfdf7875c1d71f54655af5c9fbdd92fc0
zb5f08f4089b0bbab30beab5736591239b085daa8e38ac7b6c7cc4afd8f6872f4ef1fd16684c99f
z3cdd8be7dd48a2bdf9659a2b12f8ffef040fc17af56fa64d1489b653bfcca46cce8ddebdd2d17c
ze9170462a9327dbccc5af8a8b080343de698d061afaef60eea281c2455dff2dc2fca9ec6aa6cbf
z4a4dfbd0f345611dfba41e444646569f607eff6766978888c0585bec05fa471bfb069977482d83
z411b1099ac9f765d8f8a53e0524252446acca94dcda4a129052dae5f1f552a86ed8ac3d502da65
z52d5b8494b03bdf4a025845023496528a64e3b80106668092d2862cfda2af02104c6559c18b9a4
z5881f21d1b795f0b6fa8489a5796ff97f12cab306a055080f7132ad5c64eda3587c03d55e04f47
z705d3059d2b14ab0de9759844192267be947d7679de2456b3958ebada192ca3c274c26824ecca9
z73d08986392c1ef89c8914762e00774fdaec07752e22ad70ef4977ccf1f1dac1ecdd363d8fab52
z963023e255977ee7170ea50ed94e8740e98ba4c5d572bc181b2e61a3fb4aac389882de1f4c6b34
zf06aed913c96b73a7732fe857bc50ce01989282ccd3cf7175dc54e2057e5e8f5679c64d1713c76
zb7a0096e5752df33ec3bb116773ff828e98f7ba78c55bce84175f2819ee81961cfe028a1f6b6a5
zf41ad16d536bc792c639f04d2f44482d53b42b1a769404284f953b321e9e605c210cd503454ef8
ze30781f751f66227dbb7977c040b431b3fb9bf6af8a9092ccc0f40891c967afe798cf108eea021
z0cb17bf432650752210b3dd875e58fbc74a7b842aede776eca8d0fe49d27777fb14870e2c12ce3
z30b5df3b7dbe5a5a9464878f88cc47bb8e6f88c3ed042b59b848d5e93f11dc87b318c7b421a931
z6ec565a7019904c704d8add1169cb82b10646b367d0eefaa437fe75106693f2c482a4ee204e88e
z208adaacb8be2a04df00f89fbcd63729296cf7adafa9a337fc8b05bd4512f8306ecda3649cf414
za202c57520db49a5ba18eb0d6384ef6978ee69cc7cf0f3089b67dae7c01a4334c4fd699ec138ea
z56ab6551cfc56ea9b781b6df3a385522c72532908293cdf79e7510f216d15635625d5e54a08228
zb57bcfb5b599e9fbda1aeb5b89bc24ecadfed27c43ee5f668e410d21e09a12a9eafaef7bffc6a9
zcd702cb100b83de6eb826fe9e3a1c672570e6da8eb5c43e5791a9724995e865567f8c6d200af7a
zfcf359015c11b918514b1941bc706a5edf890d5848580557f252b17a33ece15c7c85b9da7086f7
z6b075578ad6ddd1acf4714acde7c46ee0bb0dc88855b8645ac3211eab22ef0809e05cae1421f01
za8784c1e6c3e64f15e75235ee022d090410ae3fe45435c7611a88e25831e44dbd7a91f61338f61
z36d5c468c9052acf6b91c746993474ebba89c9ba39be041ebcc5222f712822997996bbd86f62bf
za95f0df6b2cd8af4a3f93ec18e500dbaad8fbb69aeb5dc96af6df56e0d944f12886d7efeeb2adf
z148a2da622a8260ee67bc7177abf9c19fc32ea12f081a80bae248424f540c91c29ecfd31c51297
z226d646a46dba3d90875833795ba47c2407ac062673e0709e8a3f9f37a13c45fd9b290699cb62f
z3bb01652f1d0e041931931e83f328964cbd639de93852c458e531249b2adc5ef6f77de25823ca4
z2ba697efd89894cfeef77df9c97ef5ea13532eb599e267edcac1bbfc932fe7fe3fb548d89c7092
z8cc815ba5a430f0086534e25d8a0716eacc9016903fb7eb9fa899fd203b705c614c115e0d1fa59
z07ff150493b0c3d828b7c8fadcb6458d5ed660e8e2e54a50abf5e67e2448d08c61f439e4151352
zf294672689d2c93332cf9fb03d6b4c572ac23d04db17a7315a6ca528200232d403db4414f67f67
z49d5711763515016586530473a2383c6aa2bc1f2df4acd923b2d0ed0e0e77171980fe6fcdac4da
z761bec5039c4d6c710f119aa16b4aa5709975a9506c2a87b996cede542997b8eac79159bc247ae
z29227170b3c8b0e95a4bd0db420e200878a89a328000022f8793ff1d4bf151c0dafc17c2d4a510
z081809382b2902431f069b3ce41e8ca5fae2311faa749dbaf0074c61e28b9bed24a1c040f9224e
z4b5e21e4250783fabec24d5d91a9efbdd6e4c0f6225808db7412799eeddba09fdd4a913b87a0e9
z839d0538d12b26e1abec305c45045d5bfe2ed4eb736412d3f418b4e778f3348c63bdfb34052c55
z9ac8cd792da5965f998c77eb3f49206a19900fc4c9046f7776ffec3572aeb0ff91b1a70b9ffc94
z33c25d19690f3dff8e92a2e094867cc156bd0ed00f6e8165cc34b6ea91d428507ae0aa1cc46cda
zc475196166bafccb5ad7d2ebcd5a9b0812f3721488f167f864a4e3376413ba1c7c9ea1c5e2fcb8
zeadcaf02d5ddffb6dcac3ef69293292f7a75bff9770a3e36a8a4c0a82bc7f1f52c6674d3349e44
z5d72071a1abac5159c87de57f95da80433b67b65be39db6c07aee6605aab42f0886b8b1297618e
z73192330efafca6243641dbdf10788c8113c4f358c96a9d67a35679538017e450be2877197c729
zee100e45b636d5499fda489a633d0b2029bca173238ff4007e90be811359543171128bc67a21e2
z387f64fb118165507e890a9e99d13ea5c6324e009a5038d5c8d1dc4dd6a72f19901f33a5336b09
z76e82b85597f706ad7b69f7f15fbb028bc128e7682827c11a14767e13224b1ffff5d037ea121d4
z0dc1d1f37f5c4150c5b76139bdb198a4e547d71514f8d1653e2aac0a2e8b92d69c52974c683597
ze79bbd77d120742b80c79740e0664d1bfa6676dcb30d5cd9712b49688098ca6a9bbd5bef5d1cdf
z193d887b3e18ec2c43c049002bb1a87467c48dc4ff55e19bfcb3049fc01e8c66abf48fb399f295
zc9d37d5d8227654e925b8faa25960c821d0d0908ec372a06e47be06540eee653508e250d474e7d
zda23647599e8d7fc106db736d82cc8885c88ec3a021bef5a9c6ef0a1c113e46900d5abe1618b6c
z606a115aee41304285d17f086738a2e2c1336710e678ca74a3670cb6870fac5821b7c2b89c8656
z67335339ba800af52dcde5c594147dd1cfdf47e269187ed6e512f5e28535cabdaa96d74e05f091
z9be10bbec3669745b8e09fc201dd16054012da5a6cf34178e67448b910ea16ce00eb99142f9687
z36a97aa65bbaf682d5cec23e6689f5dbbbfa526089c98e3376bec8a68de1d74418ef9a6a5ae496
z88d14fbfe2e7918a41b3f0178cc0c8c63aede4f61e67679c4df164704ae72b6b7fb8679dcce6fc
z8137455aaec31bdf67a1a81130e0f5b12d1d3354deb66a7a760575031f4c689a5e320ce8df257d
z1b0367ac519f546ad7c3ace46959dc2c9cb9a561170eea2ab9c494c76e53c0c84ae0977a239419
z6b6bf0c9e2e042bbb155193bede37e0a2cb2372d55259f84a8f32ef29380e48a92c1cd53f9d678
z7a6d6523168f4a851e94195393eb8365943a1852f895dbba708521874f3662f98229dc8d670ecc
zcca6cc27e155aa7cb8093aaaa2f5a4248ad9871931d00a28242b3eef08d7cdaf6c276e19544e68
zf73f28c062ec1652f70f3529a83f505b23268b83e54c58a84f65b443a51a1ea0f9fe41b32e6700
z3f53d72f06852f7990666f8e24cb42515b6a8f89c309787b0267271bf7d1923d23f3dcad148d60
zc88a114a0b39d71a3e9c509f6d4b8bd7606dca70018c5354419f81fd6a0635d3aa8682ecf2acab
z7c28cfb9eab24a51f5bb22b776e3570f03671156c6c82b438b73178bc8e6e36dfe61bfbb5855b6
zf62d507523c0d81058febfdecc0aeb3c0a59501bfb44ed5b4bc80eccff15adf1460ce020021901
z83298df6ccb97aa96e627d774df9340ac60c36b7c7471f250685ac7a2a8693d9d9d3672759ce3e
zebe3b57cb35d049efd3dba0cbf9aabf031026de4e71ef83958e6646c76d5c93a61f0038d4c21a0
z218d8e6a8944a88e125e70197c0739bffd4aa2aedf192c70ce1f2606ba5e06384ac4f7c5734707
z31fb5fb78479e460807451d09007c6dd8177fb03f0112547b5ab3093e30fe082abaed389826195
z97599fa675455f1474e733dc1ea2794ea18d2f5faa053b8549727cf03bb59ea4c385bb3f4a9089
z26d8bdd4a3aff963e8d12f14a886f40831a038e6c3a9ae66f191bc03afa9f7af53a6c98459e646
z20ff6f67af7a8af0deee4d1800917f5b6c0360f323c1d7c8559d12532daf1840d3ac2b5d151c63
z1af6e79521da57a7e76b202613714cefe2b92625e71c46d654c0f1ec5ab6987d42c228eeab3730
zd6c147fc5c0202964bf6bb49b625ec52faa983765dc659ee174b055bf4c6b79795e8b060c65abf
z141fa73671e6266b5f71c536a8362de55054df62b250d90376fd314ea714748cf23d141a8ea409
z5f7bb78cdeffd37981312fbdd9a1af31ed49d8cefed160c876b777b82a73dd5bf7a400c6b3b8ba
z5221f4a2bf8d3057eec61eae9d718c25c9920b13bfdd1ca67ad652b3fcf7577a1adf5f46a468be
z74b9761c172f89f014ff9d02ce98b18ad2e7e4191edb01a6ba55f032fabbcc9c8606e7ecdf6326
z75e620b453438f83b3d95f958326d7b891561418fb93b94f3a6e319ceb7c7506c0f939a891db33
z121b7c49efe1aaee1db608fb5508423fb994c7e7509a22cac4c1dbd2c17d08777d0c0c4bfbc8fe
z8e2f6ec7278f78d444f777e2d6300945cc5c77acea518c1c936b7b678ddc4f199ab517b0c2de0f
zed20b714b8fdd1c054577e75
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_i2c_slave_checks.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
